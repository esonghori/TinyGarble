
module Lite_MIPS ( clk, rst, g_init, e_init, o );
  input [2047:0] g_init;
  input [2047:0] e_init;
  output [2047:0] o;
  input clk, rst;
  wire   N24, N25, N26, N27, N28, N29, \PC_Next/n311 , \PC_Next/n310 ,
         \PC_Next/n309 , \PC_Next/n308 , \PC_Next/pc_future[27] ,
         \PC_Next/pc_future[26] , \PC_Next/pc_future[25] ,
         \PC_Next/pc_future[24] , \PC_Next/pc_future[23] ,
         \PC_Next/pc_future[22] , \PC_Next/pc_future[21] ,
         \PC_Next/pc_future[20] , \PC_Next/pc_future[19] ,
         \PC_Next/pc_future[18] , \PC_Next/pc_future[17] ,
         \PC_Next/pc_future[16] , \PC_Next/pc_future[15] ,
         \PC_Next/pc_future[14] , \PC_Next/pc_future[13] ,
         \PC_Next/pc_future[12] , \PC_Next/pc_future[11] ,
         \PC_Next/pc_future[10] , \PC_Next/pc_future[9] ,
         \PC_Next/pc_future[8] , \PC_Next/pc_future[7] ,
         \PC_Next/pc_future[6] , \PC_Next/pc_future[5] ,
         \PC_Next/pc_future[4] , \PC_Next/pc_future[3] ,
         \PC_Next/pc_future[2] , \PC_Next/pc_jump[31] , \PC_Next/pc_jump[30] ,
         \PC_Next/pc_jump[29] , \PC_Next/pc_jump[28] , \PC_Next/pc_jump[27] ,
         \PC_Next/pc_jump[26] , \PC_Next/pc_jump[25] , \PC_Next/pc_jump[24] ,
         \PC_Next/pc_jump[23] , \PC_Next/pc_jump[22] , \PC_Next/pc_jump[21] ,
         \PC_Next/pc_jump[20] , \PC_Next/pc_jump[19] , \PC_Next/pc_jump[18] ,
         \PC_Next/pc_jump[17] , \PC_Next/pc_jump[16] , \PC_Next/pc_jump[15] ,
         \PC_Next/pc_jump[14] , \PC_Next/pc_jump[13] , \PC_Next/pc_jump[12] ,
         \PC_Next/pc_jump[11] , \PC_Next/pc_jump[10] , \PC_Next/pc_jump[9] ,
         \PC_Next/pc_jump[8] , \PC_Next/pc_jump[7] , \PC_Next/pc_jump[6] ,
         \PC_Next/pc_jump[5] , \PC_Next/pc_jump[4] , \PC_Next/pc_jump[3] ,
         \PC_Next/pc_jump[2] , \Inst_Mem/n1984 , \Inst_Mem/n1983 ,
         \Inst_Mem/n1982 , \Inst_Mem/n1981 , \Inst_Mem/n1980 ,
         \Inst_Mem/n1979 , \Inst_Mem/n1978 , \Inst_Mem/n1977 ,
         \Inst_Mem/n1976 , \Inst_Mem/n1975 , \Inst_Mem/n1974 ,
         \Inst_Mem/n1973 , \Inst_Mem/n1972 , \Inst_Mem/n1971 ,
         \Inst_Mem/n1970 , \Inst_Mem/n1969 , \Inst_Mem/n1968 ,
         \Inst_Mem/n1967 , \Inst_Mem/n1966 , \Inst_Mem/n1965 ,
         \Inst_Mem/n1964 , \Inst_Mem/n1963 , \Inst_Mem/n1962 ,
         \Inst_Mem/n1961 , \Inst_Mem/n1960 , \Inst_Mem/n1959 ,
         \Inst_Mem/n1958 , \Inst_Mem/n1957 , \Inst_Mem/n1956 ,
         \Inst_Mem/n1955 , \Inst_Mem/n1954 , \Inst_Mem/n1953 ,
         \Inst_Mem/n1952 , \Inst_Mem/n1951 , \Inst_Mem/n1950 ,
         \Inst_Mem/n1949 , \Inst_Mem/n1948 , \Inst_Mem/n1947 ,
         \Inst_Mem/n1946 , \Inst_Mem/n1945 , \Inst_Mem/n1944 ,
         \Inst_Mem/n1943 , \Inst_Mem/n1942 , \Inst_Mem/n1941 ,
         \Inst_Mem/n1940 , \Inst_Mem/n1939 , \Inst_Mem/n1938 ,
         \Inst_Mem/n1937 , \Inst_Mem/n1936 , \Inst_Mem/n1935 ,
         \Inst_Mem/n1934 , \Inst_Mem/n1933 , \Inst_Mem/n1932 ,
         \Inst_Mem/n1931 , \Inst_Mem/n1930 , \Inst_Mem/n1929 ,
         \Inst_Mem/n1928 , \Inst_Mem/n1927 , \Inst_Mem/n1926 ,
         \Inst_Mem/n1925 , \Inst_Mem/n1924 , \Inst_Mem/n1923 ,
         \Inst_Mem/n1922 , \Inst_Mem/n1921 , \Inst_Mem/n1920 ,
         \Inst_Mem/n1919 , \Inst_Mem/n1918 , \Inst_Mem/n1917 ,
         \Inst_Mem/n1916 , \Inst_Mem/n1915 , \Inst_Mem/n1914 ,
         \Inst_Mem/n1913 , \Inst_Mem/n1912 , \Inst_Mem/n1911 ,
         \Inst_Mem/n1910 , \Inst_Mem/n1909 , \Inst_Mem/n1908 ,
         \Inst_Mem/n1907 , \Inst_Mem/n1906 , \Inst_Mem/n1905 ,
         \Inst_Mem/n1904 , \Inst_Mem/n1903 , \Inst_Mem/n1902 ,
         \Inst_Mem/n1901 , \Inst_Mem/n1900 , \Inst_Mem/n1899 ,
         \Inst_Mem/n1898 , \Inst_Mem/n1897 , \Inst_Mem/n1896 ,
         \Inst_Mem/n1895 , \Inst_Mem/n1894 , \Inst_Mem/n1893 ,
         \Inst_Mem/n1892 , \Inst_Mem/n1891 , \Inst_Mem/n1890 ,
         \Inst_Mem/n1889 , \Inst_Mem/n1888 , \Inst_Mem/n1887 ,
         \Inst_Mem/n1886 , \Inst_Mem/n1885 , \Inst_Mem/n1884 ,
         \Inst_Mem/n1883 , \Inst_Mem/n1882 , \Inst_Mem/n1881 ,
         \Inst_Mem/n1880 , \Inst_Mem/n1879 , \Inst_Mem/n1878 ,
         \Inst_Mem/n1877 , \Inst_Mem/n1876 , \Inst_Mem/n1875 ,
         \Inst_Mem/n1874 , \Inst_Mem/n1873 , \Inst_Mem/n1872 ,
         \Inst_Mem/n1871 , \Inst_Mem/n1870 , \Inst_Mem/n1869 ,
         \Inst_Mem/n1868 , \Inst_Mem/n1867 , \Inst_Mem/n1866 ,
         \Inst_Mem/n1865 , \Inst_Mem/n1864 , \Inst_Mem/n1863 ,
         \Inst_Mem/n1862 , \Inst_Mem/n1861 , \Inst_Mem/n1860 ,
         \Inst_Mem/n1859 , \Inst_Mem/n1858 , \Inst_Mem/n1857 ,
         \Inst_Mem/n1856 , \Inst_Mem/n1855 , \Inst_Mem/n1854 ,
         \Inst_Mem/n1853 , \Inst_Mem/n1852 , \Inst_Mem/n1851 ,
         \Inst_Mem/n1850 , \Inst_Mem/n1849 , \Inst_Mem/n1848 ,
         \Inst_Mem/n1847 , \Inst_Mem/n1846 , \Inst_Mem/n1845 ,
         \Inst_Mem/n1844 , \Inst_Mem/n1843 , \Inst_Mem/n1842 ,
         \Inst_Mem/n1841 , \Inst_Mem/n1840 , \Inst_Mem/n1839 ,
         \Inst_Mem/n1838 , \Inst_Mem/n1837 , \Inst_Mem/n1836 ,
         \Inst_Mem/n1835 , \Inst_Mem/n1834 , \Inst_Mem/n1833 ,
         \Inst_Mem/n1832 , \Inst_Mem/n1831 , \Inst_Mem/n1830 ,
         \Inst_Mem/n1829 , \Inst_Mem/n1828 , \Inst_Mem/n1827 ,
         \Inst_Mem/n1826 , \Inst_Mem/n1825 , \Inst_Mem/n1824 ,
         \Inst_Mem/n1823 , \Inst_Mem/n1822 , \Inst_Mem/n1821 ,
         \Inst_Mem/n1820 , \Inst_Mem/n1819 , \Inst_Mem/n1818 ,
         \Inst_Mem/n1817 , \Inst_Mem/n1816 , \Inst_Mem/n1815 ,
         \Inst_Mem/n1814 , \Inst_Mem/n1813 , \Inst_Mem/n1812 ,
         \Inst_Mem/n1811 , \Inst_Mem/n1810 , \Inst_Mem/n1809 ,
         \Inst_Mem/n1808 , \Inst_Mem/n1807 , \Inst_Mem/n1806 ,
         \Inst_Mem/n1805 , \Inst_Mem/n1804 , \Inst_Mem/n1803 ,
         \Inst_Mem/n1802 , \Inst_Mem/n1801 , \Inst_Mem/n1800 ,
         \Inst_Mem/n1799 , \Inst_Mem/n1798 , \Inst_Mem/n1797 ,
         \Inst_Mem/n1796 , \Inst_Mem/n1795 , \Inst_Mem/n1794 ,
         \Inst_Mem/n1793 , \Inst_Mem/n1792 , \Inst_Mem/n1791 ,
         \Inst_Mem/n1790 , \Inst_Mem/n1789 , \Inst_Mem/n1788 ,
         \Inst_Mem/n1787 , \Inst_Mem/n1786 , \Inst_Mem/n1785 ,
         \Inst_Mem/n1784 , \Inst_Mem/n1783 , \Inst_Mem/n1782 ,
         \Inst_Mem/n1781 , \Inst_Mem/n1780 , \Inst_Mem/n1779 ,
         \Inst_Mem/n1778 , \Inst_Mem/n1777 , \Inst_Mem/n1776 ,
         \Inst_Mem/n1775 , \Inst_Mem/n1774 , \Inst_Mem/n1773 ,
         \Inst_Mem/n1772 , \Inst_Mem/n1771 , \Inst_Mem/n1770 ,
         \Inst_Mem/n1769 , \Inst_Mem/n1768 , \Inst_Mem/n1767 ,
         \Inst_Mem/n1766 , \Inst_Mem/n1765 , \Inst_Mem/n1764 ,
         \Inst_Mem/n1763 , \Inst_Mem/n1762 , \Inst_Mem/n1761 ,
         \Inst_Mem/n1760 , \Inst_Mem/n1759 , \Inst_Mem/n1758 ,
         \Inst_Mem/n1757 , \Inst_Mem/n1756 , \Inst_Mem/n1755 ,
         \Inst_Mem/n1754 , \Inst_Mem/n1753 , \Inst_Mem/n1752 ,
         \Inst_Mem/n1751 , \Inst_Mem/n1750 , \Inst_Mem/n1749 ,
         \Inst_Mem/n1748 , \Inst_Mem/n1747 , \Inst_Mem/n1746 ,
         \Inst_Mem/n1745 , \Inst_Mem/n1744 , \Inst_Mem/n1743 ,
         \Inst_Mem/n1742 , \Inst_Mem/n1741 , \Inst_Mem/n1740 ,
         \Inst_Mem/n1739 , \Inst_Mem/n1738 , \Inst_Mem/n1737 ,
         \Inst_Mem/n1736 , \Inst_Mem/n1735 , \Inst_Mem/n1734 ,
         \Inst_Mem/n1733 , \Inst_Mem/n1732 , \Inst_Mem/n1731 ,
         \Inst_Mem/n1730 , \Inst_Mem/n1729 , \Inst_Mem/n1728 ,
         \Inst_Mem/n1727 , \Inst_Mem/n1726 , \Inst_Mem/n1725 ,
         \Inst_Mem/n1724 , \Inst_Mem/n1723 , \Inst_Mem/n1722 ,
         \Inst_Mem/n1721 , \Inst_Mem/n1720 , \Inst_Mem/n1719 ,
         \Inst_Mem/n1718 , \Inst_Mem/n1717 , \Inst_Mem/n1716 ,
         \Inst_Mem/n1715 , \Inst_Mem/n1714 , \Inst_Mem/n1713 ,
         \Inst_Mem/n1712 , \Inst_Mem/n1711 , \Inst_Mem/n1710 ,
         \Inst_Mem/n1709 , \Inst_Mem/n1708 , \Inst_Mem/n1707 ,
         \Inst_Mem/n1706 , \Inst_Mem/n1705 , \Inst_Mem/n1704 ,
         \Inst_Mem/n1703 , \Inst_Mem/n1702 , \Inst_Mem/n1701 ,
         \Inst_Mem/n1700 , \Inst_Mem/n1699 , \Inst_Mem/n1698 ,
         \Inst_Mem/n1697 , \Inst_Mem/n1696 , \Inst_Mem/n1695 ,
         \Inst_Mem/n1694 , \Inst_Mem/n1693 , \Inst_Mem/n1692 ,
         \Inst_Mem/n1691 , \Inst_Mem/n1690 , \Inst_Mem/n1689 ,
         \Inst_Mem/n1688 , \Inst_Mem/n1687 , \Inst_Mem/n1686 ,
         \Inst_Mem/n1685 , \Inst_Mem/n1684 , \Inst_Mem/n1683 ,
         \Inst_Mem/n1682 , \Inst_Mem/n1681 , \Inst_Mem/n1680 ,
         \Inst_Mem/n1679 , \Inst_Mem/n1678 , \Inst_Mem/n1677 ,
         \Inst_Mem/n1676 , \Inst_Mem/n1675 , \Inst_Mem/n1674 ,
         \Inst_Mem/n1673 , \Inst_Mem/n1672 , \Inst_Mem/n1671 ,
         \Inst_Mem/n1670 , \Inst_Mem/n1669 , \Inst_Mem/n1668 ,
         \Inst_Mem/n1667 , \Inst_Mem/n1666 , \Inst_Mem/n1665 ,
         \Inst_Mem/n1664 , \Inst_Mem/n1663 , \Inst_Mem/n1662 ,
         \Inst_Mem/n1661 , \Inst_Mem/n1660 , \Inst_Mem/n1659 ,
         \Inst_Mem/n1658 , \Inst_Mem/n1657 , \Inst_Mem/n1656 ,
         \Inst_Mem/n1655 , \Inst_Mem/n1654 , \Inst_Mem/n1653 ,
         \Inst_Mem/n1652 , \Inst_Mem/n1651 , \Inst_Mem/n1650 ,
         \Inst_Mem/n1649 , \Inst_Mem/n1648 , \Inst_Mem/n1647 ,
         \Inst_Mem/n1646 , \Inst_Mem/n1645 , \Inst_Mem/n1644 ,
         \Inst_Mem/n1643 , \Inst_Mem/n1642 , \Inst_Mem/n1641 ,
         \Inst_Mem/n1640 , \Inst_Mem/n1639 , \Inst_Mem/n1638 ,
         \Inst_Mem/n1637 , \Inst_Mem/n1636 , \Inst_Mem/n1635 ,
         \Inst_Mem/n1634 , \Inst_Mem/n1633 , \Inst_Mem/n1632 ,
         \Inst_Mem/n1631 , \Inst_Mem/n1630 , \Inst_Mem/n1629 ,
         \Inst_Mem/n1628 , \Inst_Mem/n1627 , \Inst_Mem/n1626 ,
         \Inst_Mem/n1625 , \Inst_Mem/n1624 , \Inst_Mem/n1623 ,
         \Inst_Mem/n1622 , \Inst_Mem/n1621 , \Inst_Mem/n1620 ,
         \Inst_Mem/n1619 , \Inst_Mem/n1618 , \Inst_Mem/n1617 ,
         \Inst_Mem/n1616 , \Inst_Mem/n1615 , \Inst_Mem/n1614 ,
         \Inst_Mem/n1613 , \Inst_Mem/n1612 , \Inst_Mem/n1611 ,
         \Inst_Mem/n1610 , \Inst_Mem/n1609 , \Inst_Mem/n1608 ,
         \Inst_Mem/n1607 , \Inst_Mem/n1606 , \Inst_Mem/n1605 ,
         \Inst_Mem/n1604 , \Inst_Mem/n1603 , \Inst_Mem/n1602 ,
         \Inst_Mem/n1601 , \Inst_Mem/n1600 , \Inst_Mem/n1599 ,
         \Inst_Mem/n1598 , \Inst_Mem/n1597 , \Inst_Mem/n1596 ,
         \Inst_Mem/n1595 , \Inst_Mem/n1594 , \Inst_Mem/n1593 ,
         \Inst_Mem/n1592 , \Inst_Mem/n1591 , \Inst_Mem/n1590 ,
         \Inst_Mem/n1589 , \Inst_Mem/n1588 , \Inst_Mem/n1587 ,
         \Inst_Mem/n1586 , \Inst_Mem/n1585 , \Inst_Mem/n1584 ,
         \Inst_Mem/n1583 , \Inst_Mem/n1582 , \Inst_Mem/n1581 ,
         \Inst_Mem/n1580 , \Inst_Mem/n1579 , \Inst_Mem/n1578 ,
         \Inst_Mem/n1577 , \Inst_Mem/n1576 , \Inst_Mem/n1575 ,
         \Inst_Mem/n1574 , \Inst_Mem/n1573 , \Inst_Mem/n1572 ,
         \Inst_Mem/n1571 , \Inst_Mem/n1570 , \Inst_Mem/n1569 ,
         \Inst_Mem/n1568 , \Inst_Mem/n1567 , \Inst_Mem/n1566 ,
         \Inst_Mem/n1565 , \Inst_Mem/n1564 , \Inst_Mem/n1563 ,
         \Inst_Mem/n1562 , \Inst_Mem/n1561 , \Inst_Mem/n1560 ,
         \Inst_Mem/n1559 , \Inst_Mem/n1558 , \Inst_Mem/n1557 ,
         \Inst_Mem/n1556 , \Inst_Mem/n1555 , \Inst_Mem/n1554 ,
         \Inst_Mem/n1553 , \Inst_Mem/n1552 , \Inst_Mem/n1551 ,
         \Inst_Mem/n1550 , \Inst_Mem/n1549 , \Inst_Mem/n1548 ,
         \Inst_Mem/n1547 , \Inst_Mem/n1546 , \Inst_Mem/n1545 ,
         \Inst_Mem/n1544 , \Inst_Mem/n1543 , \Inst_Mem/n1542 ,
         \Inst_Mem/n1541 , \Inst_Mem/n1540 , \Inst_Mem/n1539 ,
         \Inst_Mem/n1538 , \Inst_Mem/n1537 , \Inst_Mem/n1536 ,
         \Inst_Mem/n1535 , \Inst_Mem/n1534 , \Inst_Mem/n1533 ,
         \Inst_Mem/n1532 , \Inst_Mem/n1531 , \Inst_Mem/n1530 ,
         \Inst_Mem/n1529 , \Inst_Mem/n1528 , \Inst_Mem/n1527 ,
         \Inst_Mem/n1526 , \Inst_Mem/n1525 , \Inst_Mem/n1524 ,
         \Inst_Mem/n1523 , \Inst_Mem/n1522 , \Inst_Mem/n1521 ,
         \Inst_Mem/n1520 , \Inst_Mem/n1519 , \Inst_Mem/n1518 ,
         \Inst_Mem/n1517 , \Inst_Mem/n1516 , \Inst_Mem/n1515 ,
         \Inst_Mem/n1514 , \Inst_Mem/n1513 , \Inst_Mem/n1512 ,
         \Inst_Mem/n1511 , \Inst_Mem/n1510 , \Inst_Mem/n1509 ,
         \Inst_Mem/n1508 , \Inst_Mem/n1507 , \Inst_Mem/n1506 ,
         \Inst_Mem/n1505 , \Inst_Mem/n1504 , \Inst_Mem/n1503 ,
         \Inst_Mem/n1502 , \Inst_Mem/n1501 , \Inst_Mem/n1500 ,
         \Inst_Mem/n1499 , \Inst_Mem/n1498 , \Inst_Mem/n1497 ,
         \Inst_Mem/n1496 , \Inst_Mem/n1495 , \Inst_Mem/n1494 ,
         \Inst_Mem/n1493 , \Inst_Mem/n1492 , \Inst_Mem/n1491 ,
         \Inst_Mem/n1490 , \Inst_Mem/n1489 , \Inst_Mem/n1488 ,
         \Inst_Mem/n1487 , \Inst_Mem/n1486 , \Inst_Mem/n1485 ,
         \Inst_Mem/n1484 , \Inst_Mem/n1483 , \Inst_Mem/n1482 ,
         \Inst_Mem/n1481 , \Inst_Mem/n1480 , \Inst_Mem/n1479 ,
         \Inst_Mem/n1478 , \Inst_Mem/n1477 , \Inst_Mem/n1476 ,
         \Inst_Mem/n1475 , \Inst_Mem/n1474 , \Inst_Mem/n1473 ,
         \Inst_Mem/n1472 , \Inst_Mem/n1471 , \Inst_Mem/n1470 ,
         \Inst_Mem/n1469 , \Inst_Mem/n1468 , \Inst_Mem/n1467 ,
         \Inst_Mem/n1466 , \Inst_Mem/n1465 , \Inst_Mem/n1464 ,
         \Inst_Mem/n1463 , \Inst_Mem/n1462 , \Inst_Mem/n1461 ,
         \Inst_Mem/n1460 , \Inst_Mem/n1459 , \Inst_Mem/n1458 ,
         \Inst_Mem/n1457 , \Inst_Mem/n1456 , \Inst_Mem/n1455 ,
         \Inst_Mem/n1454 , \Inst_Mem/n1453 , \Inst_Mem/n1452 ,
         \Inst_Mem/n1451 , \Inst_Mem/n1450 , \Inst_Mem/n1449 ,
         \Inst_Mem/n1448 , \Inst_Mem/n1447 , \Inst_Mem/n1446 ,
         \Inst_Mem/n1445 , \Inst_Mem/n1444 , \Inst_Mem/n1443 ,
         \Inst_Mem/n1442 , \Inst_Mem/n1441 , \Inst_Mem/n1440 ,
         \Inst_Mem/n1439 , \Inst_Mem/n1438 , \Inst_Mem/n1437 ,
         \Inst_Mem/n1436 , \Inst_Mem/n1435 , \Inst_Mem/n1434 ,
         \Inst_Mem/n1433 , \Inst_Mem/n1432 , \Inst_Mem/n1431 ,
         \Inst_Mem/n1430 , \Inst_Mem/n1429 , \Inst_Mem/n1428 ,
         \Inst_Mem/n1427 , \Inst_Mem/n1426 , \Inst_Mem/n1425 ,
         \Inst_Mem/n1424 , \Inst_Mem/n1423 , \Inst_Mem/n1422 ,
         \Inst_Mem/n1421 , \Inst_Mem/n1420 , \Inst_Mem/n1419 ,
         \Inst_Mem/n1418 , \Inst_Mem/n1417 , \Inst_Mem/n1416 ,
         \Inst_Mem/n1415 , \Inst_Mem/n1414 , \Inst_Mem/n1413 ,
         \Inst_Mem/n1412 , \Inst_Mem/n1411 , \Inst_Mem/n1410 ,
         \Inst_Mem/n1409 , \Inst_Mem/n1408 , \Inst_Mem/n1407 ,
         \Inst_Mem/n1406 , \Inst_Mem/n1405 , \Inst_Mem/n1404 ,
         \Inst_Mem/n1403 , \Inst_Mem/n1402 , \Inst_Mem/n1401 ,
         \Inst_Mem/n1400 , \Inst_Mem/n1399 , \Inst_Mem/n1398 ,
         \Inst_Mem/n1397 , \Inst_Mem/n1396 , \Inst_Mem/n1395 ,
         \Inst_Mem/n1394 , \Inst_Mem/n1393 , \Inst_Mem/n1392 ,
         \Inst_Mem/n1391 , \Inst_Mem/n1390 , \Inst_Mem/n1389 ,
         \Inst_Mem/n1388 , \Inst_Mem/n1387 , \Inst_Mem/n1386 ,
         \Inst_Mem/n1385 , \Inst_Mem/n1384 , \Inst_Mem/n1383 ,
         \Inst_Mem/n1382 , \Inst_Mem/n1381 , \Inst_Mem/n1380 ,
         \Inst_Mem/n1379 , \Inst_Mem/n1378 , \Inst_Mem/n1377 ,
         \Inst_Mem/n1376 , \Inst_Mem/n1375 , \Inst_Mem/n1374 ,
         \Inst_Mem/n1373 , \Inst_Mem/n1372 , \Inst_Mem/n1371 ,
         \Inst_Mem/n1370 , \Inst_Mem/n1369 , \Inst_Mem/n1368 ,
         \Inst_Mem/n1367 , \Inst_Mem/n1366 , \Inst_Mem/n1365 ,
         \Inst_Mem/n1364 , \Inst_Mem/n1363 , \Inst_Mem/n1362 ,
         \Inst_Mem/n1361 , \Inst_Mem/n1360 , \Inst_Mem/n1359 ,
         \Inst_Mem/n1358 , \Inst_Mem/n1357 , \Inst_Mem/n1356 ,
         \Inst_Mem/n1355 , \Inst_Mem/n1354 , \Inst_Mem/n1353 ,
         \Inst_Mem/n1352 , \Inst_Mem/n1351 , \Inst_Mem/n1350 ,
         \Inst_Mem/n1349 , \Inst_Mem/n1348 , \Inst_Mem/n1347 ,
         \Inst_Mem/n1346 , \Inst_Mem/n1345 , \Inst_Mem/n1344 ,
         \Inst_Mem/n1343 , \Inst_Mem/n1342 , \Inst_Mem/n1341 ,
         \Inst_Mem/n1340 , \Inst_Mem/n1339 , \Inst_Mem/n1338 ,
         \Inst_Mem/n1337 , \Inst_Mem/n1336 , \Inst_Mem/n1335 ,
         \Inst_Mem/n1334 , \Inst_Mem/n1333 , \Inst_Mem/n1332 ,
         \Inst_Mem/n1331 , \Inst_Mem/n1330 , \Inst_Mem/n1329 ,
         \Inst_Mem/n1328 , \Inst_Mem/n1327 , \Inst_Mem/n1326 ,
         \Inst_Mem/n1325 , \Inst_Mem/n1324 , \Inst_Mem/n1323 ,
         \Inst_Mem/n1322 , \Inst_Mem/n1321 , \Inst_Mem/n1320 ,
         \Inst_Mem/n1319 , \Inst_Mem/n1318 , \Inst_Mem/n1317 ,
         \Inst_Mem/n1316 , \Inst_Mem/n1315 , \Inst_Mem/n1314 ,
         \Inst_Mem/n1313 , \Inst_Mem/n1312 , \Inst_Mem/n1311 ,
         \Inst_Mem/n1310 , \Inst_Mem/n1309 , \Inst_Mem/n1308 ,
         \Inst_Mem/n1307 , \Inst_Mem/n1306 , \Inst_Mem/n1305 ,
         \Inst_Mem/n1304 , \Inst_Mem/n1303 , \Inst_Mem/n1302 ,
         \Inst_Mem/n1301 , \Inst_Mem/n1300 , \Inst_Mem/n1299 ,
         \Inst_Mem/n1298 , \Inst_Mem/n1297 , \Inst_Mem/n1296 ,
         \Inst_Mem/n1295 , \Inst_Mem/n1294 , \Inst_Mem/n1293 ,
         \Inst_Mem/n1292 , \Inst_Mem/n1291 , \Inst_Mem/n1290 ,
         \Inst_Mem/n1289 , \Inst_Mem/n1288 , \Inst_Mem/n1287 ,
         \Inst_Mem/n1286 , \Inst_Mem/n1285 , \Inst_Mem/n1284 ,
         \Inst_Mem/n1283 , \Inst_Mem/n1282 , \Inst_Mem/n1281 ,
         \Inst_Mem/n1280 , \Inst_Mem/n1279 , \Inst_Mem/n1278 ,
         \Inst_Mem/n1277 , \Inst_Mem/n1276 , \Inst_Mem/n1275 ,
         \Inst_Mem/n1274 , \Inst_Mem/n1273 , \Inst_Mem/n1272 ,
         \Inst_Mem/n1271 , \Inst_Mem/n1270 , \Inst_Mem/n1269 ,
         \Inst_Mem/n1268 , \Inst_Mem/n1267 , \Inst_Mem/n1266 ,
         \Inst_Mem/n1265 , \Inst_Mem/n1264 , \Inst_Mem/n1263 ,
         \Inst_Mem/n1262 , \Inst_Mem/n1261 , \Inst_Mem/n1260 ,
         \Inst_Mem/n1259 , \Inst_Mem/n1258 , \Inst_Mem/n1257 ,
         \Inst_Mem/n1256 , \Inst_Mem/n1255 , \Inst_Mem/n1254 ,
         \Inst_Mem/n1253 , \Inst_Mem/n1252 , \Inst_Mem/n1251 ,
         \Inst_Mem/n1250 , \Inst_Mem/n1249 , \Inst_Mem/n1248 ,
         \Inst_Mem/n1247 , \Inst_Mem/n1246 , \Inst_Mem/n1245 ,
         \Inst_Mem/n1244 , \Inst_Mem/n1243 , \Inst_Mem/n1242 ,
         \Inst_Mem/n1241 , \Inst_Mem/n1240 , \Inst_Mem/n1239 ,
         \Inst_Mem/n1238 , \Inst_Mem/n1237 , \Inst_Mem/n1236 ,
         \Inst_Mem/n1235 , \Inst_Mem/n1234 , \Inst_Mem/n1233 ,
         \Inst_Mem/n1232 , \Inst_Mem/n1231 , \Inst_Mem/n1230 ,
         \Inst_Mem/n1229 , \Inst_Mem/n1228 , \Inst_Mem/n1227 ,
         \Inst_Mem/n1226 , \Inst_Mem/n1225 , \Inst_Mem/n1224 ,
         \Inst_Mem/n1223 , \Inst_Mem/n1222 , \Inst_Mem/n1221 ,
         \Inst_Mem/n1220 , \Inst_Mem/n1219 , \Inst_Mem/n1218 ,
         \Inst_Mem/n1217 , \Inst_Mem/n1216 , \Inst_Mem/n1215 ,
         \Inst_Mem/n1214 , \Inst_Mem/n1213 , \Inst_Mem/n1212 ,
         \Inst_Mem/n1211 , \Inst_Mem/n1210 , \Inst_Mem/n1209 ,
         \Inst_Mem/n1208 , \Inst_Mem/n1207 , \Inst_Mem/n1206 ,
         \Inst_Mem/n1205 , \Inst_Mem/n1204 , \Inst_Mem/n1203 ,
         \Inst_Mem/n1202 , \Inst_Mem/n1201 , \Inst_Mem/n1200 ,
         \Inst_Mem/n1199 , \Inst_Mem/n1198 , \Inst_Mem/n1197 ,
         \Inst_Mem/n1196 , \Inst_Mem/n1195 , \Inst_Mem/n1194 ,
         \Inst_Mem/n1193 , \Inst_Mem/n1192 , \Inst_Mem/n1191 ,
         \Inst_Mem/n1190 , \Inst_Mem/n1189 , \Inst_Mem/n1188 ,
         \Inst_Mem/n1187 , \Inst_Mem/n1186 , \Inst_Mem/n1185 ,
         \Inst_Mem/n1184 , \Inst_Mem/n1183 , \Inst_Mem/n1182 ,
         \Inst_Mem/n1181 , \Inst_Mem/n1180 , \Inst_Mem/n1179 ,
         \Inst_Mem/n1178 , \Inst_Mem/n1177 , \Inst_Mem/n1176 ,
         \Inst_Mem/n1175 , \Inst_Mem/n1174 , \Inst_Mem/n1173 ,
         \Inst_Mem/n1172 , \Inst_Mem/n1171 , \Inst_Mem/n1170 ,
         \Inst_Mem/n1169 , \Inst_Mem/n1168 , \Inst_Mem/n1167 ,
         \Inst_Mem/n1166 , \Inst_Mem/n1165 , \Inst_Mem/n1164 ,
         \Inst_Mem/n1163 , \Inst_Mem/n1162 , \Inst_Mem/n1161 ,
         \Inst_Mem/n1160 , \Inst_Mem/n1159 , \Inst_Mem/n1158 ,
         \Inst_Mem/n1157 , \Inst_Mem/n1156 , \Inst_Mem/n1155 ,
         \Inst_Mem/n1154 , \Inst_Mem/n1153 , \Inst_Mem/n1152 ,
         \Inst_Mem/n1151 , \Inst_Mem/n1150 , \Inst_Mem/n1149 ,
         \Inst_Mem/n1148 , \Inst_Mem/n1147 , \Inst_Mem/n1146 ,
         \Inst_Mem/n1145 , \Inst_Mem/n1144 , \Inst_Mem/n1143 ,
         \Inst_Mem/n1142 , \Inst_Mem/n1141 , \Inst_Mem/n1140 ,
         \Inst_Mem/n1139 , \Inst_Mem/n1138 , \Inst_Mem/n1137 ,
         \Inst_Mem/n1136 , \Inst_Mem/n1135 , \Inst_Mem/n1134 ,
         \Inst_Mem/n1133 , \Inst_Mem/n1132 , \Inst_Mem/n1131 ,
         \Inst_Mem/n1130 , \Inst_Mem/n1129 , \Inst_Mem/n1128 ,
         \Inst_Mem/n1127 , \Inst_Mem/n1126 , \Inst_Mem/n1125 ,
         \Inst_Mem/n1124 , \Inst_Mem/n1123 , \Inst_Mem/n1122 ,
         \Inst_Mem/n1121 , \Inst_Mem/n1120 , \Inst_Mem/n1119 ,
         \Inst_Mem/n1118 , \Inst_Mem/n1117 , \Inst_Mem/n1116 ,
         \Inst_Mem/n1115 , \Inst_Mem/n1114 , \Inst_Mem/n1113 ,
         \Inst_Mem/n1112 , \Inst_Mem/n1111 , \Inst_Mem/n1110 ,
         \Inst_Mem/n1109 , \Inst_Mem/n1108 , \Inst_Mem/n1107 ,
         \Inst_Mem/n1106 , \Inst_Mem/n1105 , \Inst_Mem/n1104 ,
         \Inst_Mem/n1103 , \Inst_Mem/n1102 , \Inst_Mem/n1101 ,
         \Inst_Mem/n1100 , \Inst_Mem/n1099 , \Inst_Mem/n1098 ,
         \Inst_Mem/n1097 , \Inst_Mem/n1096 , \Inst_Mem/n1095 ,
         \Inst_Mem/n1094 , \Inst_Mem/n1093 , \Inst_Mem/n1092 ,
         \Inst_Mem/n1091 , \Inst_Mem/n1090 , \Inst_Mem/n1089 ,
         \Inst_Mem/n1088 , \Inst_Mem/n1087 , \Inst_Mem/n1086 ,
         \Inst_Mem/n1085 , \Inst_Mem/n1084 , \Inst_Mem/n1083 ,
         \Inst_Mem/n1082 , \Inst_Mem/n1081 , \Inst_Mem/n1080 ,
         \Inst_Mem/n1079 , \Inst_Mem/n1078 , \Inst_Mem/n1077 ,
         \Inst_Mem/n1076 , \Inst_Mem/n1075 , \Inst_Mem/n1074 ,
         \Inst_Mem/n1073 , \Inst_Mem/n1072 , \Inst_Mem/n1071 ,
         \Inst_Mem/n1070 , \Inst_Mem/n1069 , \Inst_Mem/n1068 ,
         \Inst_Mem/n1067 , \Inst_Mem/n1066 , \Inst_Mem/n1065 ,
         \Inst_Mem/n1064 , \Inst_Mem/n1063 , \Inst_Mem/n1062 ,
         \Inst_Mem/n1061 , \Inst_Mem/n1060 , \Inst_Mem/n1059 ,
         \Inst_Mem/n1058 , \Inst_Mem/n1057 , \Inst_Mem/n1056 ,
         \Inst_Mem/n1055 , \Inst_Mem/n1054 , \Inst_Mem/n1053 ,
         \Inst_Mem/n1052 , \Inst_Mem/n1051 , \Inst_Mem/n1050 ,
         \Inst_Mem/n1049 , \Inst_Mem/n1048 , \Inst_Mem/n1047 ,
         \Inst_Mem/n1046 , \Inst_Mem/n1045 , \Inst_Mem/n1044 ,
         \Inst_Mem/n1043 , \Inst_Mem/n1042 , \Inst_Mem/n1041 ,
         \Inst_Mem/n1040 , \Inst_Mem/n1039 , \Inst_Mem/n1038 ,
         \Inst_Mem/n1037 , \Inst_Mem/n1036 , \Inst_Mem/n1035 ,
         \Inst_Mem/n1034 , \Inst_Mem/n1033 , \Inst_Mem/n1032 ,
         \Inst_Mem/n1031 , \Inst_Mem/n1030 , \Inst_Mem/n1029 ,
         \Inst_Mem/n1028 , \Inst_Mem/n1027 , \Inst_Mem/n1026 ,
         \Inst_Mem/n1025 , \Inst_Mem/n1024 , \Inst_Mem/n1023 ,
         \Inst_Mem/n1022 , \Inst_Mem/n1021 , \Inst_Mem/n1020 ,
         \Inst_Mem/n1019 , \Inst_Mem/n1018 , \Inst_Mem/n1017 ,
         \Inst_Mem/n1016 , \Inst_Mem/n1015 , \Inst_Mem/n1014 ,
         \Inst_Mem/n1013 , \Inst_Mem/n1012 , \Inst_Mem/n1011 ,
         \Inst_Mem/n1010 , \Inst_Mem/n1009 , \Inst_Mem/n1008 ,
         \Inst_Mem/n1007 , \Inst_Mem/n1006 , \Inst_Mem/n1005 ,
         \Inst_Mem/n1004 , \Inst_Mem/n1003 , \Inst_Mem/n1002 ,
         \Inst_Mem/n1001 , \Inst_Mem/n1000 , \Inst_Mem/n999 , \Inst_Mem/n998 ,
         \Inst_Mem/n997 , \Inst_Mem/n996 , \Inst_Mem/n995 , \Inst_Mem/n994 ,
         \Inst_Mem/n993 , \Inst_Mem/n992 , \Inst_Mem/n991 , \Inst_Mem/n990 ,
         \Inst_Mem/n989 , \Inst_Mem/n988 , \Inst_Mem/n987 , \Inst_Mem/n986 ,
         \Inst_Mem/n985 , \Inst_Mem/n984 , \Inst_Mem/n983 , \Inst_Mem/n982 ,
         \Inst_Mem/n981 , \Inst_Mem/n980 , \Inst_Mem/n979 , \Inst_Mem/n978 ,
         \Inst_Mem/n977 , \Inst_Mem/n976 , \Inst_Mem/n975 , \Inst_Mem/n974 ,
         \Inst_Mem/n973 , \Inst_Mem/n972 , \Inst_Mem/n971 , \Inst_Mem/n970 ,
         \Inst_Mem/n969 , \Inst_Mem/n968 , \Inst_Mem/n967 , \Inst_Mem/n966 ,
         \Inst_Mem/n965 , \Inst_Mem/n964 , \Inst_Mem/n963 , \Inst_Mem/n962 ,
         \Inst_Mem/n961 , \Inst_Mem/n960 , \Inst_Mem/n959 , \Inst_Mem/n958 ,
         \Inst_Mem/n957 , \Inst_Mem/n956 , \Inst_Mem/n955 , \Inst_Mem/n954 ,
         \Inst_Mem/n953 , \Inst_Mem/n952 , \Inst_Mem/n951 , \Inst_Mem/n950 ,
         \Inst_Mem/n949 , \Inst_Mem/n948 , \Inst_Mem/n947 , \Inst_Mem/n946 ,
         \Inst_Mem/n945 , \Inst_Mem/n944 , \Inst_Mem/n943 , \Inst_Mem/n942 ,
         \Inst_Mem/n941 , \Inst_Mem/n940 , \Inst_Mem/n939 , \Inst_Mem/n938 ,
         \Inst_Mem/n937 , \Inst_Mem/n936 , \Inst_Mem/n935 , \Inst_Mem/n934 ,
         \Inst_Mem/n933 , \Inst_Mem/n932 , \Inst_Mem/n931 , \Inst_Mem/n930 ,
         \Inst_Mem/n929 , \Inst_Mem/n928 , \Inst_Mem/n927 , \Inst_Mem/n926 ,
         \Inst_Mem/n925 , \Inst_Mem/n924 , \Inst_Mem/n923 , \Inst_Mem/n922 ,
         \Inst_Mem/n921 , \Inst_Mem/n920 , \Inst_Mem/n919 , \Inst_Mem/n918 ,
         \Inst_Mem/n917 , \Inst_Mem/n916 , \Inst_Mem/n915 , \Inst_Mem/n914 ,
         \Inst_Mem/n913 , \Inst_Mem/n912 , \Inst_Mem/n911 , \Inst_Mem/n910 ,
         \Inst_Mem/n909 , \Inst_Mem/n908 , \Inst_Mem/n907 , \Inst_Mem/n906 ,
         \Inst_Mem/n905 , \Inst_Mem/n904 , \Inst_Mem/n903 , \Inst_Mem/n902 ,
         \Inst_Mem/n901 , \Inst_Mem/n900 , \Inst_Mem/n899 , \Inst_Mem/n898 ,
         \Inst_Mem/n897 , \Inst_Mem/n896 , \Inst_Mem/n895 , \Inst_Mem/n894 ,
         \Inst_Mem/n893 , \Inst_Mem/n892 , \Inst_Mem/n891 , \Inst_Mem/n890 ,
         \Inst_Mem/n889 , \Inst_Mem/n888 , \Inst_Mem/n887 , \Inst_Mem/n886 ,
         \Inst_Mem/n885 , \Inst_Mem/n884 , \Inst_Mem/n883 , \Inst_Mem/n882 ,
         \Inst_Mem/n881 , \Inst_Mem/n880 , \Inst_Mem/n879 , \Inst_Mem/n878 ,
         \Inst_Mem/n877 , \Inst_Mem/n876 , \Inst_Mem/n875 , \Inst_Mem/n874 ,
         \Inst_Mem/n873 , \Inst_Mem/n872 , \Inst_Mem/n871 , \Inst_Mem/n870 ,
         \Inst_Mem/n869 , \Inst_Mem/n868 , \Inst_Mem/n867 , \Inst_Mem/n866 ,
         \Inst_Mem/n865 , \Inst_Mem/n864 , \Inst_Mem/n863 , \Inst_Mem/n862 ,
         \Inst_Mem/n861 , \Inst_Mem/n860 , \Inst_Mem/n859 , \Inst_Mem/n858 ,
         \Inst_Mem/n857 , \Inst_Mem/n856 , \Inst_Mem/n855 , \Inst_Mem/n854 ,
         \Inst_Mem/n853 , \Inst_Mem/n852 , \Inst_Mem/n851 , \Inst_Mem/n850 ,
         \Inst_Mem/n849 , \Inst_Mem/n848 , \Inst_Mem/n847 , \Inst_Mem/n846 ,
         \Inst_Mem/n845 , \Inst_Mem/n844 , \Inst_Mem/n843 , \Inst_Mem/n842 ,
         \Inst_Mem/n841 , \Inst_Mem/n840 , \Inst_Mem/n839 , \Inst_Mem/n838 ,
         \Inst_Mem/n837 , \Inst_Mem/n836 , \Inst_Mem/n835 , \Inst_Mem/n834 ,
         \Inst_Mem/n833 , \Inst_Mem/n832 , \Inst_Mem/n831 , \Inst_Mem/n830 ,
         \Inst_Mem/n829 , \Inst_Mem/n828 , \Inst_Mem/n827 , \Inst_Mem/n826 ,
         \Inst_Mem/n825 , \Inst_Mem/n824 , \Inst_Mem/n823 , \Inst_Mem/n822 ,
         \Inst_Mem/n821 , \Inst_Mem/n820 , \Inst_Mem/n819 , \Inst_Mem/n818 ,
         \Inst_Mem/n817 , \Inst_Mem/n816 , \Inst_Mem/n815 , \Inst_Mem/n814 ,
         \Inst_Mem/n813 , \Inst_Mem/n812 , \Inst_Mem/n811 , \Inst_Mem/n810 ,
         \Inst_Mem/n809 , \Inst_Mem/n808 , \Inst_Mem/n807 , \Inst_Mem/n806 ,
         \Inst_Mem/n805 , \Inst_Mem/n804 , \Inst_Mem/n803 , \Inst_Mem/n802 ,
         \Inst_Mem/n801 , \Inst_Mem/n800 , \Inst_Mem/n799 , \Inst_Mem/n798 ,
         \Inst_Mem/n797 , \Inst_Mem/n796 , \Inst_Mem/n795 , \Inst_Mem/n794 ,
         \Inst_Mem/n793 , \Inst_Mem/n792 , \Inst_Mem/n791 , \Inst_Mem/n790 ,
         \Inst_Mem/n789 , \Inst_Mem/n788 , \Inst_Mem/n787 , \Inst_Mem/n786 ,
         \Inst_Mem/n785 , \Inst_Mem/n784 , \Inst_Mem/n783 , \Inst_Mem/n782 ,
         \Inst_Mem/n781 , \Inst_Mem/n780 , \Inst_Mem/n779 , \Inst_Mem/n778 ,
         \Inst_Mem/n777 , \Inst_Mem/n776 , \Inst_Mem/n775 , \Inst_Mem/n774 ,
         \Inst_Mem/n773 , \Inst_Mem/n772 , \Inst_Mem/n771 , \Inst_Mem/n770 ,
         \Inst_Mem/n769 , \Inst_Mem/n768 , \Inst_Mem/n767 , \Inst_Mem/n766 ,
         \Inst_Mem/n765 , \Inst_Mem/n764 , \Inst_Mem/n763 , \Inst_Mem/n762 ,
         \Inst_Mem/n761 , \Inst_Mem/n760 , \Inst_Mem/n759 , \Inst_Mem/n758 ,
         \Inst_Mem/n757 , \Inst_Mem/n756 , \Inst_Mem/n755 , \Inst_Mem/n754 ,
         \Inst_Mem/n753 , \Inst_Mem/n752 , \Inst_Mem/n751 , \Inst_Mem/n750 ,
         \Inst_Mem/n749 , \Inst_Mem/n748 , \Inst_Mem/n747 , \Inst_Mem/n746 ,
         \Inst_Mem/n745 , \Inst_Mem/n744 , \Inst_Mem/n743 , \Inst_Mem/n742 ,
         \Inst_Mem/n741 , \Inst_Mem/n740 , \Inst_Mem/n739 , \Inst_Mem/n738 ,
         \Inst_Mem/n737 , \Inst_Mem/n736 , \Inst_Mem/n735 , \Inst_Mem/n734 ,
         \Inst_Mem/n733 , \Inst_Mem/n732 , \Inst_Mem/n731 , \Inst_Mem/n730 ,
         \Inst_Mem/n729 , \Inst_Mem/n728 , \Inst_Mem/n727 , \Inst_Mem/n726 ,
         \Inst_Mem/n725 , \Inst_Mem/n724 , \Inst_Mem/n723 , \Inst_Mem/n722 ,
         \Inst_Mem/n721 , \Inst_Mem/n720 , \Inst_Mem/n719 , \Inst_Mem/n718 ,
         \Inst_Mem/n717 , \Inst_Mem/n716 , \Inst_Mem/n715 , \Inst_Mem/n714 ,
         \Inst_Mem/n713 , \Inst_Mem/n712 , \Inst_Mem/n711 , \Inst_Mem/n710 ,
         \Inst_Mem/n709 , \Inst_Mem/n708 , \Inst_Mem/n707 , \Inst_Mem/n706 ,
         \Inst_Mem/n705 , \Inst_Mem/n704 , \Inst_Mem/n703 , \Inst_Mem/n702 ,
         \Inst_Mem/n701 , \Inst_Mem/n700 , \Inst_Mem/n699 , \Inst_Mem/n698 ,
         \Inst_Mem/n697 , \Inst_Mem/n696 , \Inst_Mem/n695 , \Inst_Mem/n694 ,
         \Inst_Mem/n693 , \Inst_Mem/n692 , \Inst_Mem/n691 , \Inst_Mem/n690 ,
         \Inst_Mem/n689 , \Inst_Mem/n688 , \Inst_Mem/n687 , \Inst_Mem/n686 ,
         \Inst_Mem/n685 , \Inst_Mem/n684 , \Inst_Mem/n683 , \Inst_Mem/n682 ,
         \Inst_Mem/n681 , \Inst_Mem/n680 , \Inst_Mem/n679 , \Inst_Mem/n678 ,
         \Inst_Mem/n677 , \Inst_Mem/n676 , \Inst_Mem/n675 , \Inst_Mem/n674 ,
         \Inst_Mem/n673 , \Inst_Mem/n672 , \Inst_Mem/n671 , \Inst_Mem/n670 ,
         \Inst_Mem/n669 , \Inst_Mem/n668 , \Inst_Mem/n667 , \Inst_Mem/n666 ,
         \Inst_Mem/n665 , \Inst_Mem/n664 , \Inst_Mem/n663 , \Inst_Mem/n662 ,
         \Inst_Mem/n661 , \Inst_Mem/n660 , \Inst_Mem/n659 , \Inst_Mem/n658 ,
         \Inst_Mem/n657 , \Inst_Mem/n656 , \Inst_Mem/n655 , \Inst_Mem/n654 ,
         \Inst_Mem/n653 , \Inst_Mem/n652 , \Inst_Mem/n651 , \Inst_Mem/n650 ,
         \Inst_Mem/n649 , \Inst_Mem/n648 , \Inst_Mem/n647 , \Inst_Mem/n646 ,
         \Inst_Mem/n645 , \Inst_Mem/n644 , \Inst_Mem/n643 , \Inst_Mem/n642 ,
         \Inst_Mem/n641 , \Inst_Mem/n640 , \Inst_Mem/n639 , \Inst_Mem/n638 ,
         \Inst_Mem/n637 , \Inst_Mem/n636 , \Inst_Mem/n635 , \Inst_Mem/n634 ,
         \Inst_Mem/n633 , \Inst_Mem/n632 , \Inst_Mem/n631 , \Inst_Mem/n630 ,
         \Inst_Mem/n629 , \Inst_Mem/n628 , \Inst_Mem/n627 , \Inst_Mem/n626 ,
         \Inst_Mem/n625 , \Inst_Mem/n624 , \Inst_Mem/n623 , \Inst_Mem/n622 ,
         \Inst_Mem/n621 , \Inst_Mem/n620 , \Inst_Mem/n619 , \Inst_Mem/n618 ,
         \Inst_Mem/n617 , \Inst_Mem/n616 , \Inst_Mem/n615 , \Inst_Mem/n614 ,
         \Inst_Mem/n613 , \Inst_Mem/n612 , \Inst_Mem/n611 , \Inst_Mem/n610 ,
         \Inst_Mem/n609 , \Inst_Mem/n608 , \Inst_Mem/n607 , \Inst_Mem/n606 ,
         \Inst_Mem/n605 , \Inst_Mem/n604 , \Inst_Mem/n603 , \Inst_Mem/n602 ,
         \Inst_Mem/n601 , \Inst_Mem/n600 , \Inst_Mem/n599 , \Inst_Mem/n598 ,
         \Inst_Mem/n597 , \Inst_Mem/n596 , \Inst_Mem/n595 , \Inst_Mem/n594 ,
         \Inst_Mem/n593 , \Inst_Mem/n592 , \Inst_Mem/n591 , \Inst_Mem/n590 ,
         \Inst_Mem/n589 , \Inst_Mem/n588 , \Inst_Mem/n587 , \Inst_Mem/n586 ,
         \Inst_Mem/n585 , \Inst_Mem/n584 , \Inst_Mem/n583 , \Inst_Mem/n582 ,
         \Inst_Mem/n581 , \Inst_Mem/n580 , \Inst_Mem/n579 , \Inst_Mem/n578 ,
         \Inst_Mem/n577 , \Inst_Mem/n576 , \Inst_Mem/n575 , \Inst_Mem/n574 ,
         \Inst_Mem/n573 , \Inst_Mem/n572 , \Inst_Mem/n571 , \Inst_Mem/n570 ,
         \Inst_Mem/n569 , \Inst_Mem/n568 , \Inst_Mem/n567 , \Inst_Mem/n566 ,
         \Inst_Mem/n565 , \Inst_Mem/n564 , \Inst_Mem/n563 , \Inst_Mem/n562 ,
         \Inst_Mem/n561 , \Inst_Mem/n560 , \Inst_Mem/n559 , \Inst_Mem/n558 ,
         \Inst_Mem/n557 , \Inst_Mem/n556 , \Inst_Mem/n555 , \Inst_Mem/n554 ,
         \Inst_Mem/n553 , \Inst_Mem/n552 , \Inst_Mem/n551 , \Inst_Mem/n550 ,
         \Inst_Mem/n549 , \Inst_Mem/n548 , \Inst_Mem/n547 , \Inst_Mem/n546 ,
         \Inst_Mem/n545 , \Inst_Mem/n544 , \Inst_Mem/n543 , \Inst_Mem/n542 ,
         \Inst_Mem/n541 , \Inst_Mem/n540 , \Inst_Mem/n539 , \Inst_Mem/n538 ,
         \Inst_Mem/n537 , \Inst_Mem/n536 , \Inst_Mem/n535 , \Inst_Mem/n534 ,
         \Inst_Mem/n533 , \Inst_Mem/n532 , \Inst_Mem/n531 , \Inst_Mem/n530 ,
         \Inst_Mem/n529 , \Inst_Mem/n528 , \Inst_Mem/n527 , \Inst_Mem/n526 ,
         \Inst_Mem/n525 , \Inst_Mem/n524 , \Inst_Mem/n523 , \Inst_Mem/n522 ,
         \Inst_Mem/n521 , \Inst_Mem/n520 , \Inst_Mem/n519 , \Inst_Mem/n518 ,
         \Inst_Mem/n517 , \Inst_Mem/n516 , \Inst_Mem/n515 , \Inst_Mem/n514 ,
         \Inst_Mem/n513 , \Inst_Mem/n512 , \Inst_Mem/n511 , \Inst_Mem/n510 ,
         \Inst_Mem/n509 , \Inst_Mem/n508 , \Inst_Mem/n507 , \Inst_Mem/n506 ,
         \Inst_Mem/n505 , \Inst_Mem/n504 , \Inst_Mem/n503 , \Inst_Mem/n502 ,
         \Inst_Mem/n501 , \Inst_Mem/n500 , \Inst_Mem/n499 , \Inst_Mem/n498 ,
         \Inst_Mem/n497 , \Inst_Mem/n496 , \Inst_Mem/n495 , \Inst_Mem/n494 ,
         \Inst_Mem/n493 , \Inst_Mem/n492 , \Inst_Mem/n491 , \Inst_Mem/n490 ,
         \Inst_Mem/n489 , \Inst_Mem/n488 , \Inst_Mem/n487 , \Inst_Mem/n486 ,
         \Inst_Mem/n485 , \Inst_Mem/n484 , \Inst_Mem/n483 , \Inst_Mem/n482 ,
         \Inst_Mem/n481 , \Inst_Mem/n480 , \Inst_Mem/n479 , \Inst_Mem/n478 ,
         \Inst_Mem/n477 , \Inst_Mem/n476 , \Inst_Mem/n475 , \Inst_Mem/n474 ,
         \Inst_Mem/n473 , \Inst_Mem/n472 , \Inst_Mem/n471 , \Inst_Mem/n470 ,
         \Inst_Mem/n469 , \Inst_Mem/n468 , \Inst_Mem/n467 , \Inst_Mem/n466 ,
         \Inst_Mem/n465 , \Inst_Mem/n464 , \Inst_Mem/n463 , \Inst_Mem/n462 ,
         \Inst_Mem/n461 , \Inst_Mem/n460 , \Inst_Mem/n459 , \Inst_Mem/n458 ,
         \Inst_Mem/n457 , \Inst_Mem/n456 , \Inst_Mem/n455 , \Inst_Mem/n454 ,
         \Inst_Mem/n453 , \Inst_Mem/n452 , \Inst_Mem/n451 , \Inst_Mem/n450 ,
         \Inst_Mem/n449 , \Inst_Mem/n448 , \Inst_Mem/n447 , \Inst_Mem/n446 ,
         \Inst_Mem/n445 , \Inst_Mem/n444 , \Inst_Mem/n443 , \Inst_Mem/n442 ,
         \Inst_Mem/n441 , \Inst_Mem/n440 , \Inst_Mem/n439 , \Inst_Mem/n438 ,
         \Inst_Mem/n437 , \Inst_Mem/n436 , \Inst_Mem/n435 , \Inst_Mem/n434 ,
         \Inst_Mem/n433 , \Inst_Mem/n432 , \Inst_Mem/n431 , \Inst_Mem/n430 ,
         \Inst_Mem/n429 , \Inst_Mem/n428 , \Inst_Mem/n427 , \Inst_Mem/n426 ,
         \Inst_Mem/n425 , \Inst_Mem/n424 , \Inst_Mem/n423 , \Inst_Mem/n422 ,
         \Inst_Mem/n421 , \Inst_Mem/n420 , \Inst_Mem/n419 , \Inst_Mem/n418 ,
         \Inst_Mem/n417 , \Inst_Mem/n416 , \Inst_Mem/n415 , \Inst_Mem/n414 ,
         \Inst_Mem/n413 , \Inst_Mem/n412 , \Inst_Mem/n411 , \Inst_Mem/n410 ,
         \Inst_Mem/n409 , \Inst_Mem/n408 , \Inst_Mem/n407 , \Inst_Mem/n406 ,
         \Inst_Mem/n405 , \Inst_Mem/n404 , \Inst_Mem/n403 , \Inst_Mem/n402 ,
         \Inst_Mem/n401 , \Inst_Mem/n400 , \Inst_Mem/n399 , \Inst_Mem/n398 ,
         \Inst_Mem/n397 , \Inst_Mem/n396 , \Inst_Mem/n395 , \Inst_Mem/n394 ,
         \Inst_Mem/n393 , \Inst_Mem/n392 , \Inst_Mem/n391 , \Inst_Mem/n390 ,
         \Inst_Mem/n389 , \Inst_Mem/n388 , \Inst_Mem/n387 , \Inst_Mem/n386 ,
         \Inst_Mem/n385 , \Inst_Mem/n384 , \Inst_Mem/n383 , \Inst_Mem/n382 ,
         \Inst_Mem/n381 , \Inst_Mem/n380 , \Inst_Mem/n379 , \Inst_Mem/n378 ,
         \Inst_Mem/n377 , \Inst_Mem/n376 , \Inst_Mem/n375 , \Inst_Mem/n374 ,
         \Inst_Mem/n373 , \Inst_Mem/n372 , \Inst_Mem/n371 , \Inst_Mem/n370 ,
         \Inst_Mem/n369 , \Inst_Mem/n368 , \Inst_Mem/n367 , \Inst_Mem/n366 ,
         \Inst_Mem/n365 , \Inst_Mem/n364 , \Inst_Mem/n363 , \Inst_Mem/n362 ,
         \Inst_Mem/n361 , \Inst_Mem/n360 , \Inst_Mem/n359 , \Inst_Mem/n358 ,
         \Inst_Mem/n357 , \Inst_Mem/n356 , \Inst_Mem/n355 , \Inst_Mem/n354 ,
         \Inst_Mem/n353 , \Inst_Mem/n352 , \Inst_Mem/n351 , \Inst_Mem/n350 ,
         \Inst_Mem/n349 , \Inst_Mem/n348 , \Inst_Mem/n347 , \Inst_Mem/n346 ,
         \Inst_Mem/n345 , \Inst_Mem/n344 , \Inst_Mem/n343 , \Inst_Mem/n342 ,
         \Inst_Mem/n341 , \Inst_Mem/n340 , \Inst_Mem/n339 , \Inst_Mem/n338 ,
         \Inst_Mem/n337 , \Inst_Mem/n336 , \Inst_Mem/n335 , \Inst_Mem/n334 ,
         \Inst_Mem/n333 , \Inst_Mem/n332 , \Inst_Mem/n331 , \Inst_Mem/n330 ,
         \Inst_Mem/n329 , \Inst_Mem/n328 , \Inst_Mem/n327 , \Inst_Mem/n326 ,
         \Inst_Mem/n325 , \Inst_Mem/n324 , \Inst_Mem/n323 , \Inst_Mem/n322 ,
         \Inst_Mem/n321 , \Inst_Mem/n320 , \Inst_Mem/n319 , \Inst_Mem/n318 ,
         \Inst_Mem/n317 , \Inst_Mem/n316 , \Inst_Mem/n315 , \Inst_Mem/n314 ,
         \Inst_Mem/n313 , \Inst_Mem/n312 , \Inst_Mem/n311 , \Inst_Mem/n310 ,
         \Inst_Mem/n309 , \Inst_Mem/n308 , \Inst_Mem/n307 , \Inst_Mem/n306 ,
         \Inst_Mem/n305 , \Inst_Mem/n304 , \Inst_Mem/n303 , \Inst_Mem/n302 ,
         \Inst_Mem/n301 , \Inst_Mem/n300 , \Inst_Mem/n299 , \Inst_Mem/n298 ,
         \Inst_Mem/n297 , \Inst_Mem/n296 , \Inst_Mem/n295 , \Inst_Mem/n294 ,
         \Inst_Mem/n293 , \Inst_Mem/n292 , \Inst_Mem/n291 , \Inst_Mem/n290 ,
         \Inst_Mem/n289 , \Inst_Mem/n288 , \Inst_Mem/n287 , \Inst_Mem/n286 ,
         \Inst_Mem/n285 , \Inst_Mem/n284 , \Inst_Mem/n283 , \Inst_Mem/n282 ,
         \Inst_Mem/n281 , \Inst_Mem/n280 , \Inst_Mem/n279 , \Inst_Mem/n278 ,
         \Inst_Mem/n277 , \Inst_Mem/n276 , \Inst_Mem/n275 , \Inst_Mem/n274 ,
         \Inst_Mem/n273 , \Inst_Mem/n272 , \Inst_Mem/n271 , \Inst_Mem/n270 ,
         \Inst_Mem/n269 , \Inst_Mem/n268 , \Inst_Mem/n267 , \Inst_Mem/n266 ,
         \Inst_Mem/n265 , \Inst_Mem/n264 , \Inst_Mem/n263 , \Inst_Mem/n262 ,
         \Inst_Mem/n261 , \Inst_Mem/n260 , \Inst_Mem/n259 , \Inst_Mem/n258 ,
         \Inst_Mem/n257 , \Inst_Mem/n256 , \Inst_Mem/n255 , \Inst_Mem/n254 ,
         \Inst_Mem/n253 , \Inst_Mem/n252 , \Inst_Mem/n251 , \Inst_Mem/n250 ,
         \Inst_Mem/n249 , \Inst_Mem/n248 , \Inst_Mem/n247 , \Inst_Mem/n246 ,
         \Inst_Mem/n245 , \Inst_Mem/n244 , \Inst_Mem/n243 , \Inst_Mem/n242 ,
         \Inst_Mem/n241 , \Inst_Mem/n240 , \Inst_Mem/n239 , \Inst_Mem/n238 ,
         \Inst_Mem/n237 , \Inst_Mem/n236 , \Inst_Mem/n235 , \Inst_Mem/n234 ,
         \Inst_Mem/n233 , \Inst_Mem/n232 , \Inst_Mem/n231 , \Inst_Mem/n230 ,
         \Inst_Mem/n229 , \Inst_Mem/n228 , \Inst_Mem/n227 , \Inst_Mem/n226 ,
         \Inst_Mem/n225 , \Inst_Mem/n224 , \Inst_Mem/n223 , \Inst_Mem/n222 ,
         \Inst_Mem/n221 , \Inst_Mem/n220 , \Inst_Mem/n219 , \Inst_Mem/n218 ,
         \Inst_Mem/n217 , \Inst_Mem/n216 , \Inst_Mem/n215 , \Inst_Mem/n214 ,
         \Inst_Mem/n213 , \Inst_Mem/n212 , \Inst_Mem/n211 , \Inst_Mem/n210 ,
         \Inst_Mem/n209 , \Inst_Mem/n208 , \Inst_Mem/n207 , \Inst_Mem/n206 ,
         \Inst_Mem/n205 , \Inst_Mem/n204 , \Inst_Mem/n203 , \Inst_Mem/n202 ,
         \Inst_Mem/n201 , \Inst_Mem/n200 , \Inst_Mem/n199 , \Inst_Mem/n198 ,
         \Inst_Mem/n197 , \Inst_Mem/n196 , \Inst_Mem/n195 , \Inst_Mem/n194 ,
         \Inst_Mem/n193 , \Inst_Mem/n192 , \Inst_Mem/n191 , \Inst_Mem/n190 ,
         \Inst_Mem/n189 , \Inst_Mem/n188 , \Inst_Mem/n187 , \Inst_Mem/n186 ,
         \Inst_Mem/n185 , \Inst_Mem/n184 , \Inst_Mem/n183 , \Inst_Mem/n182 ,
         \Inst_Mem/n181 , \Inst_Mem/n180 , \Inst_Mem/n179 , \Inst_Mem/n178 ,
         \Inst_Mem/n177 , \Inst_Mem/n176 , \Inst_Mem/n175 , \Inst_Mem/n174 ,
         \Inst_Mem/n173 , \Inst_Mem/n172 , \Inst_Mem/n171 , \Inst_Mem/n170 ,
         \Inst_Mem/n169 , \Inst_Mem/n168 , \Inst_Mem/n167 , \Inst_Mem/n166 ,
         \Inst_Mem/n165 , \Inst_Mem/n164 , \Inst_Mem/n163 , \Inst_Mem/n162 ,
         \Inst_Mem/n161 , \Inst_Mem/n160 , \Inst_Mem/n159 , \Inst_Mem/n158 ,
         \Inst_Mem/n157 , \Inst_Mem/n156 , \Inst_Mem/n155 , \Inst_Mem/n154 ,
         \Inst_Mem/n153 , \Inst_Mem/n152 , \Inst_Mem/n151 , \Inst_Mem/n150 ,
         \Inst_Mem/n149 , \Inst_Mem/n148 , \Inst_Mem/n147 , \Inst_Mem/n146 ,
         \Inst_Mem/n145 , \Inst_Mem/n144 , \Inst_Mem/n143 , \Inst_Mem/n142 ,
         \Inst_Mem/n141 , \Inst_Mem/n140 , \Inst_Mem/n139 , \Inst_Mem/n138 ,
         \Inst_Mem/n137 , \Inst_Mem/n136 , \Inst_Mem/n135 , \Inst_Mem/n134 ,
         \Inst_Mem/n133 , \Inst_Mem/n132 , \Inst_Mem/n131 , \Inst_Mem/n130 ,
         \Inst_Mem/n129 , \Inst_Mem/n128 , \Inst_Mem/n127 , \Inst_Mem/n126 ,
         \Inst_Mem/n125 , \Inst_Mem/n124 , \Inst_Mem/n123 , \Inst_Mem/n122 ,
         \Inst_Mem/n121 , \Inst_Mem/n120 , \Inst_Mem/n119 , \Inst_Mem/n118 ,
         \Inst_Mem/n117 , \Inst_Mem/n116 , \Inst_Mem/n115 , \Inst_Mem/n114 ,
         \Inst_Mem/n113 , \Inst_Mem/n112 , \Inst_Mem/n111 , \Inst_Mem/n110 ,
         \Inst_Mem/n109 , \Inst_Mem/n108 , \Inst_Mem/n107 , \Inst_Mem/n106 ,
         \Inst_Mem/n105 , \Inst_Mem/n104 , \Inst_Mem/n103 , \Inst_Mem/n102 ,
         \Inst_Mem/n101 , \Inst_Mem/n100 , \Inst_Mem/n99 , \Inst_Mem/n98 ,
         \Inst_Mem/n97 , \Inst_Mem/n96 , \Inst_Mem/n95 , \Inst_Mem/n94 ,
         \Inst_Mem/n93 , \Inst_Mem/n92 , \Inst_Mem/n91 , \Inst_Mem/n90 ,
         \Inst_Mem/n89 , \Inst_Mem/n88 , \Inst_Mem/n87 , \Inst_Mem/n86 ,
         \Inst_Mem/n85 , \Inst_Mem/n84 , \Inst_Mem/n83 , \Inst_Mem/n82 ,
         \Inst_Mem/n81 , \Inst_Mem/n80 , \Inst_Mem/n79 , \Inst_Mem/n78 ,
         \Inst_Mem/n77 , \Inst_Mem/n76 , \Inst_Mem/n75 , \Inst_Mem/n74 ,
         \Inst_Mem/n73 , \Inst_Mem/n72 , \Inst_Mem/n71 , \Inst_Mem/n70 ,
         \Inst_Mem/n69 , \Inst_Mem/n68 , \Inst_Mem/n67 , \Inst_Mem/n66 ,
         \Inst_Mem/n65 , \Inst_Mem/n64 , \Inst_Mem/n63 , \Inst_Mem/n62 ,
         \Inst_Mem/n61 , \Inst_Mem/n60 , \Inst_Mem/n59 , \Inst_Mem/n58 ,
         \Inst_Mem/n57 , \Inst_Mem/n56 , \Inst_Mem/n55 , \Inst_Mem/n54 ,
         \Inst_Mem/n53 , \Inst_Mem/n52 , \Inst_Mem/n51 , \Inst_Mem/n50 ,
         \Inst_Mem/n49 , \Inst_Mem/n48 , \Inst_Mem/n47 , \Inst_Mem/n46 ,
         \Inst_Mem/n45 , \Inst_Mem/n44 , \Inst_Mem/n43 , \Inst_Mem/n42 ,
         \Inst_Mem/n41 , \Inst_Mem/n40 , \Inst_Mem/n39 , \Inst_Mem/n38 ,
         \Inst_Mem/n37 , \Inst_Mem/n36 , \Inst_Mem/n35 , \Inst_Mem/n34 ,
         \Inst_Mem/n33 , \Inst_Mem/n32 , \Inst_Mem/n31 , \Inst_Mem/n30 ,
         \Inst_Mem/n29 , \Inst_Mem/n28 , \Inst_Mem/n27 , \Inst_Mem/n26 ,
         \Inst_Mem/n25 , \Inst_Mem/n24 , \Inst_Mem/n23 , \Inst_Mem/n22 ,
         \Inst_Mem/n21 , \Inst_Mem/n20 , \Inst_Mem/n19 , \Inst_Mem/n18 ,
         \Inst_Mem/n17 , \Inst_Mem/n16 , \Inst_Mem/n15 , \Inst_Mem/n14 ,
         \Inst_Mem/n13 , \Inst_Mem/n12 , \Inst_Mem/n11 , \Inst_Mem/n10 ,
         \Inst_Mem/n9 , \Inst_Mem/n8 , \Inst_Mem/n7 , \Inst_Mem/n6 ,
         \Inst_Mem/n5 , \Inst_Mem/n4 , \Inst_Mem/n3 , \Inst_Mem/n2 ,
         \Inst_Mem/n1 , \Inst_Mem/inst_mem_reg[63][0] ,
         \Inst_Mem/inst_mem_reg[63][1] , \Inst_Mem/inst_mem_reg[63][2] ,
         \Inst_Mem/inst_mem_reg[63][3] , \Inst_Mem/inst_mem_reg[63][4] ,
         \Inst_Mem/inst_mem_reg[63][5] , \Inst_Mem/inst_mem_reg[63][6] ,
         \Inst_Mem/inst_mem_reg[63][7] , \Inst_Mem/inst_mem_reg[63][8] ,
         \Inst_Mem/inst_mem_reg[63][9] , \Inst_Mem/inst_mem_reg[63][10] ,
         \Inst_Mem/inst_mem_reg[63][11] , \Inst_Mem/inst_mem_reg[63][12] ,
         \Inst_Mem/inst_mem_reg[63][13] , \Inst_Mem/inst_mem_reg[63][14] ,
         \Inst_Mem/inst_mem_reg[63][15] , \Inst_Mem/inst_mem_reg[63][16] ,
         \Inst_Mem/inst_mem_reg[63][17] , \Inst_Mem/inst_mem_reg[63][18] ,
         \Inst_Mem/inst_mem_reg[63][19] , \Inst_Mem/inst_mem_reg[63][20] ,
         \Inst_Mem/inst_mem_reg[63][21] , \Inst_Mem/inst_mem_reg[63][22] ,
         \Inst_Mem/inst_mem_reg[63][23] , \Inst_Mem/inst_mem_reg[63][24] ,
         \Inst_Mem/inst_mem_reg[63][25] , \Inst_Mem/inst_mem_reg[63][26] ,
         \Inst_Mem/inst_mem_reg[63][27] , \Inst_Mem/inst_mem_reg[63][28] ,
         \Inst_Mem/inst_mem_reg[63][29] , \Inst_Mem/inst_mem_reg[63][30] ,
         \Inst_Mem/inst_mem_reg[63][31] , \Inst_Mem/inst_mem_reg[62][0] ,
         \Inst_Mem/inst_mem_reg[62][1] , \Inst_Mem/inst_mem_reg[62][2] ,
         \Inst_Mem/inst_mem_reg[62][3] , \Inst_Mem/inst_mem_reg[62][4] ,
         \Inst_Mem/inst_mem_reg[62][5] , \Inst_Mem/inst_mem_reg[62][6] ,
         \Inst_Mem/inst_mem_reg[62][7] , \Inst_Mem/inst_mem_reg[62][8] ,
         \Inst_Mem/inst_mem_reg[62][9] , \Inst_Mem/inst_mem_reg[62][10] ,
         \Inst_Mem/inst_mem_reg[62][11] , \Inst_Mem/inst_mem_reg[62][12] ,
         \Inst_Mem/inst_mem_reg[62][13] , \Inst_Mem/inst_mem_reg[62][14] ,
         \Inst_Mem/inst_mem_reg[62][15] , \Inst_Mem/inst_mem_reg[62][16] ,
         \Inst_Mem/inst_mem_reg[62][17] , \Inst_Mem/inst_mem_reg[62][18] ,
         \Inst_Mem/inst_mem_reg[62][19] , \Inst_Mem/inst_mem_reg[62][20] ,
         \Inst_Mem/inst_mem_reg[62][21] , \Inst_Mem/inst_mem_reg[62][22] ,
         \Inst_Mem/inst_mem_reg[62][23] , \Inst_Mem/inst_mem_reg[62][24] ,
         \Inst_Mem/inst_mem_reg[62][25] , \Inst_Mem/inst_mem_reg[62][26] ,
         \Inst_Mem/inst_mem_reg[62][27] , \Inst_Mem/inst_mem_reg[62][28] ,
         \Inst_Mem/inst_mem_reg[62][29] , \Inst_Mem/inst_mem_reg[62][30] ,
         \Inst_Mem/inst_mem_reg[62][31] , \Inst_Mem/inst_mem_reg[61][0] ,
         \Inst_Mem/inst_mem_reg[61][1] , \Inst_Mem/inst_mem_reg[61][2] ,
         \Inst_Mem/inst_mem_reg[61][3] , \Inst_Mem/inst_mem_reg[61][4] ,
         \Inst_Mem/inst_mem_reg[61][5] , \Inst_Mem/inst_mem_reg[61][6] ,
         \Inst_Mem/inst_mem_reg[61][7] , \Inst_Mem/inst_mem_reg[61][8] ,
         \Inst_Mem/inst_mem_reg[61][9] , \Inst_Mem/inst_mem_reg[61][10] ,
         \Inst_Mem/inst_mem_reg[61][11] , \Inst_Mem/inst_mem_reg[61][12] ,
         \Inst_Mem/inst_mem_reg[61][13] , \Inst_Mem/inst_mem_reg[61][14] ,
         \Inst_Mem/inst_mem_reg[61][15] , \Inst_Mem/inst_mem_reg[61][16] ,
         \Inst_Mem/inst_mem_reg[61][17] , \Inst_Mem/inst_mem_reg[61][18] ,
         \Inst_Mem/inst_mem_reg[61][19] , \Inst_Mem/inst_mem_reg[61][20] ,
         \Inst_Mem/inst_mem_reg[61][21] , \Inst_Mem/inst_mem_reg[61][22] ,
         \Inst_Mem/inst_mem_reg[61][23] , \Inst_Mem/inst_mem_reg[61][24] ,
         \Inst_Mem/inst_mem_reg[61][25] , \Inst_Mem/inst_mem_reg[61][26] ,
         \Inst_Mem/inst_mem_reg[61][27] , \Inst_Mem/inst_mem_reg[61][28] ,
         \Inst_Mem/inst_mem_reg[61][29] , \Inst_Mem/inst_mem_reg[61][30] ,
         \Inst_Mem/inst_mem_reg[61][31] , \Inst_Mem/inst_mem_reg[60][0] ,
         \Inst_Mem/inst_mem_reg[60][1] , \Inst_Mem/inst_mem_reg[60][2] ,
         \Inst_Mem/inst_mem_reg[60][3] , \Inst_Mem/inst_mem_reg[60][4] ,
         \Inst_Mem/inst_mem_reg[60][5] , \Inst_Mem/inst_mem_reg[60][6] ,
         \Inst_Mem/inst_mem_reg[60][7] , \Inst_Mem/inst_mem_reg[60][8] ,
         \Inst_Mem/inst_mem_reg[60][9] , \Inst_Mem/inst_mem_reg[60][10] ,
         \Inst_Mem/inst_mem_reg[60][11] , \Inst_Mem/inst_mem_reg[60][12] ,
         \Inst_Mem/inst_mem_reg[60][13] , \Inst_Mem/inst_mem_reg[60][14] ,
         \Inst_Mem/inst_mem_reg[60][15] , \Inst_Mem/inst_mem_reg[60][16] ,
         \Inst_Mem/inst_mem_reg[60][17] , \Inst_Mem/inst_mem_reg[60][18] ,
         \Inst_Mem/inst_mem_reg[60][19] , \Inst_Mem/inst_mem_reg[60][20] ,
         \Inst_Mem/inst_mem_reg[60][21] , \Inst_Mem/inst_mem_reg[60][22] ,
         \Inst_Mem/inst_mem_reg[60][23] , \Inst_Mem/inst_mem_reg[60][24] ,
         \Inst_Mem/inst_mem_reg[60][25] , \Inst_Mem/inst_mem_reg[60][26] ,
         \Inst_Mem/inst_mem_reg[60][27] , \Inst_Mem/inst_mem_reg[60][28] ,
         \Inst_Mem/inst_mem_reg[60][29] , \Inst_Mem/inst_mem_reg[60][30] ,
         \Inst_Mem/inst_mem_reg[60][31] , \Inst_Mem/inst_mem_reg[59][0] ,
         \Inst_Mem/inst_mem_reg[59][1] , \Inst_Mem/inst_mem_reg[59][2] ,
         \Inst_Mem/inst_mem_reg[59][3] , \Inst_Mem/inst_mem_reg[59][4] ,
         \Inst_Mem/inst_mem_reg[59][5] , \Inst_Mem/inst_mem_reg[59][6] ,
         \Inst_Mem/inst_mem_reg[59][7] , \Inst_Mem/inst_mem_reg[59][8] ,
         \Inst_Mem/inst_mem_reg[59][9] , \Inst_Mem/inst_mem_reg[59][10] ,
         \Inst_Mem/inst_mem_reg[59][11] , \Inst_Mem/inst_mem_reg[59][12] ,
         \Inst_Mem/inst_mem_reg[59][13] , \Inst_Mem/inst_mem_reg[59][14] ,
         \Inst_Mem/inst_mem_reg[59][15] , \Inst_Mem/inst_mem_reg[59][16] ,
         \Inst_Mem/inst_mem_reg[59][17] , \Inst_Mem/inst_mem_reg[59][18] ,
         \Inst_Mem/inst_mem_reg[59][19] , \Inst_Mem/inst_mem_reg[59][20] ,
         \Inst_Mem/inst_mem_reg[59][21] , \Inst_Mem/inst_mem_reg[59][22] ,
         \Inst_Mem/inst_mem_reg[59][23] , \Inst_Mem/inst_mem_reg[59][24] ,
         \Inst_Mem/inst_mem_reg[59][25] , \Inst_Mem/inst_mem_reg[59][26] ,
         \Inst_Mem/inst_mem_reg[59][27] , \Inst_Mem/inst_mem_reg[59][28] ,
         \Inst_Mem/inst_mem_reg[59][29] , \Inst_Mem/inst_mem_reg[59][30] ,
         \Inst_Mem/inst_mem_reg[59][31] , \Inst_Mem/inst_mem_reg[58][0] ,
         \Inst_Mem/inst_mem_reg[58][1] , \Inst_Mem/inst_mem_reg[58][2] ,
         \Inst_Mem/inst_mem_reg[58][3] , \Inst_Mem/inst_mem_reg[58][4] ,
         \Inst_Mem/inst_mem_reg[58][5] , \Inst_Mem/inst_mem_reg[58][6] ,
         \Inst_Mem/inst_mem_reg[58][7] , \Inst_Mem/inst_mem_reg[58][8] ,
         \Inst_Mem/inst_mem_reg[58][9] , \Inst_Mem/inst_mem_reg[58][10] ,
         \Inst_Mem/inst_mem_reg[58][11] , \Inst_Mem/inst_mem_reg[58][12] ,
         \Inst_Mem/inst_mem_reg[58][13] , \Inst_Mem/inst_mem_reg[58][14] ,
         \Inst_Mem/inst_mem_reg[58][15] , \Inst_Mem/inst_mem_reg[58][16] ,
         \Inst_Mem/inst_mem_reg[58][17] , \Inst_Mem/inst_mem_reg[58][18] ,
         \Inst_Mem/inst_mem_reg[58][19] , \Inst_Mem/inst_mem_reg[58][20] ,
         \Inst_Mem/inst_mem_reg[58][21] , \Inst_Mem/inst_mem_reg[58][22] ,
         \Inst_Mem/inst_mem_reg[58][23] , \Inst_Mem/inst_mem_reg[58][24] ,
         \Inst_Mem/inst_mem_reg[58][25] , \Inst_Mem/inst_mem_reg[58][26] ,
         \Inst_Mem/inst_mem_reg[58][27] , \Inst_Mem/inst_mem_reg[58][28] ,
         \Inst_Mem/inst_mem_reg[58][29] , \Inst_Mem/inst_mem_reg[58][30] ,
         \Inst_Mem/inst_mem_reg[58][31] , \Inst_Mem/inst_mem_reg[57][0] ,
         \Inst_Mem/inst_mem_reg[57][1] , \Inst_Mem/inst_mem_reg[57][2] ,
         \Inst_Mem/inst_mem_reg[57][3] , \Inst_Mem/inst_mem_reg[57][4] ,
         \Inst_Mem/inst_mem_reg[57][5] , \Inst_Mem/inst_mem_reg[57][6] ,
         \Inst_Mem/inst_mem_reg[57][7] , \Inst_Mem/inst_mem_reg[57][8] ,
         \Inst_Mem/inst_mem_reg[57][9] , \Inst_Mem/inst_mem_reg[57][10] ,
         \Inst_Mem/inst_mem_reg[57][11] , \Inst_Mem/inst_mem_reg[57][12] ,
         \Inst_Mem/inst_mem_reg[57][13] , \Inst_Mem/inst_mem_reg[57][14] ,
         \Inst_Mem/inst_mem_reg[57][15] , \Inst_Mem/inst_mem_reg[57][16] ,
         \Inst_Mem/inst_mem_reg[57][17] , \Inst_Mem/inst_mem_reg[57][18] ,
         \Inst_Mem/inst_mem_reg[57][19] , \Inst_Mem/inst_mem_reg[57][20] ,
         \Inst_Mem/inst_mem_reg[57][21] , \Inst_Mem/inst_mem_reg[57][22] ,
         \Inst_Mem/inst_mem_reg[57][23] , \Inst_Mem/inst_mem_reg[57][24] ,
         \Inst_Mem/inst_mem_reg[57][25] , \Inst_Mem/inst_mem_reg[57][26] ,
         \Inst_Mem/inst_mem_reg[57][27] , \Inst_Mem/inst_mem_reg[57][28] ,
         \Inst_Mem/inst_mem_reg[57][29] , \Inst_Mem/inst_mem_reg[57][30] ,
         \Inst_Mem/inst_mem_reg[57][31] , \Inst_Mem/inst_mem_reg[56][0] ,
         \Inst_Mem/inst_mem_reg[56][1] , \Inst_Mem/inst_mem_reg[56][2] ,
         \Inst_Mem/inst_mem_reg[56][3] , \Inst_Mem/inst_mem_reg[56][4] ,
         \Inst_Mem/inst_mem_reg[56][5] , \Inst_Mem/inst_mem_reg[56][6] ,
         \Inst_Mem/inst_mem_reg[56][7] , \Inst_Mem/inst_mem_reg[56][8] ,
         \Inst_Mem/inst_mem_reg[56][9] , \Inst_Mem/inst_mem_reg[56][10] ,
         \Inst_Mem/inst_mem_reg[56][11] , \Inst_Mem/inst_mem_reg[56][12] ,
         \Inst_Mem/inst_mem_reg[56][13] , \Inst_Mem/inst_mem_reg[56][14] ,
         \Inst_Mem/inst_mem_reg[56][15] , \Inst_Mem/inst_mem_reg[56][16] ,
         \Inst_Mem/inst_mem_reg[56][17] , \Inst_Mem/inst_mem_reg[56][18] ,
         \Inst_Mem/inst_mem_reg[56][19] , \Inst_Mem/inst_mem_reg[56][20] ,
         \Inst_Mem/inst_mem_reg[56][21] , \Inst_Mem/inst_mem_reg[56][22] ,
         \Inst_Mem/inst_mem_reg[56][23] , \Inst_Mem/inst_mem_reg[56][24] ,
         \Inst_Mem/inst_mem_reg[56][25] , \Inst_Mem/inst_mem_reg[56][26] ,
         \Inst_Mem/inst_mem_reg[56][27] , \Inst_Mem/inst_mem_reg[56][28] ,
         \Inst_Mem/inst_mem_reg[56][29] , \Inst_Mem/inst_mem_reg[56][30] ,
         \Inst_Mem/inst_mem_reg[56][31] , \Inst_Mem/inst_mem_reg[55][0] ,
         \Inst_Mem/inst_mem_reg[55][1] , \Inst_Mem/inst_mem_reg[55][2] ,
         \Inst_Mem/inst_mem_reg[55][3] , \Inst_Mem/inst_mem_reg[55][4] ,
         \Inst_Mem/inst_mem_reg[55][5] , \Inst_Mem/inst_mem_reg[55][6] ,
         \Inst_Mem/inst_mem_reg[55][7] , \Inst_Mem/inst_mem_reg[55][8] ,
         \Inst_Mem/inst_mem_reg[55][9] , \Inst_Mem/inst_mem_reg[55][10] ,
         \Inst_Mem/inst_mem_reg[55][11] , \Inst_Mem/inst_mem_reg[55][12] ,
         \Inst_Mem/inst_mem_reg[55][13] , \Inst_Mem/inst_mem_reg[55][14] ,
         \Inst_Mem/inst_mem_reg[55][15] , \Inst_Mem/inst_mem_reg[55][16] ,
         \Inst_Mem/inst_mem_reg[55][17] , \Inst_Mem/inst_mem_reg[55][18] ,
         \Inst_Mem/inst_mem_reg[55][19] , \Inst_Mem/inst_mem_reg[55][20] ,
         \Inst_Mem/inst_mem_reg[55][21] , \Inst_Mem/inst_mem_reg[55][22] ,
         \Inst_Mem/inst_mem_reg[55][23] , \Inst_Mem/inst_mem_reg[55][24] ,
         \Inst_Mem/inst_mem_reg[55][25] , \Inst_Mem/inst_mem_reg[55][26] ,
         \Inst_Mem/inst_mem_reg[55][27] , \Inst_Mem/inst_mem_reg[55][28] ,
         \Inst_Mem/inst_mem_reg[55][29] , \Inst_Mem/inst_mem_reg[55][30] ,
         \Inst_Mem/inst_mem_reg[55][31] , \Inst_Mem/inst_mem_reg[54][0] ,
         \Inst_Mem/inst_mem_reg[54][1] , \Inst_Mem/inst_mem_reg[54][2] ,
         \Inst_Mem/inst_mem_reg[54][3] , \Inst_Mem/inst_mem_reg[54][4] ,
         \Inst_Mem/inst_mem_reg[54][5] , \Inst_Mem/inst_mem_reg[54][6] ,
         \Inst_Mem/inst_mem_reg[54][7] , \Inst_Mem/inst_mem_reg[54][8] ,
         \Inst_Mem/inst_mem_reg[54][9] , \Inst_Mem/inst_mem_reg[54][10] ,
         \Inst_Mem/inst_mem_reg[54][11] , \Inst_Mem/inst_mem_reg[54][12] ,
         \Inst_Mem/inst_mem_reg[54][13] , \Inst_Mem/inst_mem_reg[54][14] ,
         \Inst_Mem/inst_mem_reg[54][15] , \Inst_Mem/inst_mem_reg[54][16] ,
         \Inst_Mem/inst_mem_reg[54][17] , \Inst_Mem/inst_mem_reg[54][18] ,
         \Inst_Mem/inst_mem_reg[54][19] , \Inst_Mem/inst_mem_reg[54][20] ,
         \Inst_Mem/inst_mem_reg[54][21] , \Inst_Mem/inst_mem_reg[54][22] ,
         \Inst_Mem/inst_mem_reg[54][23] , \Inst_Mem/inst_mem_reg[54][24] ,
         \Inst_Mem/inst_mem_reg[54][25] , \Inst_Mem/inst_mem_reg[54][26] ,
         \Inst_Mem/inst_mem_reg[54][27] , \Inst_Mem/inst_mem_reg[54][28] ,
         \Inst_Mem/inst_mem_reg[54][29] , \Inst_Mem/inst_mem_reg[54][30] ,
         \Inst_Mem/inst_mem_reg[54][31] , \Inst_Mem/inst_mem_reg[53][0] ,
         \Inst_Mem/inst_mem_reg[53][1] , \Inst_Mem/inst_mem_reg[53][2] ,
         \Inst_Mem/inst_mem_reg[53][3] , \Inst_Mem/inst_mem_reg[53][4] ,
         \Inst_Mem/inst_mem_reg[53][5] , \Inst_Mem/inst_mem_reg[53][6] ,
         \Inst_Mem/inst_mem_reg[53][7] , \Inst_Mem/inst_mem_reg[53][8] ,
         \Inst_Mem/inst_mem_reg[53][9] , \Inst_Mem/inst_mem_reg[53][10] ,
         \Inst_Mem/inst_mem_reg[53][11] , \Inst_Mem/inst_mem_reg[53][12] ,
         \Inst_Mem/inst_mem_reg[53][13] , \Inst_Mem/inst_mem_reg[53][14] ,
         \Inst_Mem/inst_mem_reg[53][15] , \Inst_Mem/inst_mem_reg[53][16] ,
         \Inst_Mem/inst_mem_reg[53][17] , \Inst_Mem/inst_mem_reg[53][18] ,
         \Inst_Mem/inst_mem_reg[53][19] , \Inst_Mem/inst_mem_reg[53][20] ,
         \Inst_Mem/inst_mem_reg[53][21] , \Inst_Mem/inst_mem_reg[53][22] ,
         \Inst_Mem/inst_mem_reg[53][23] , \Inst_Mem/inst_mem_reg[53][24] ,
         \Inst_Mem/inst_mem_reg[53][25] , \Inst_Mem/inst_mem_reg[53][26] ,
         \Inst_Mem/inst_mem_reg[53][27] , \Inst_Mem/inst_mem_reg[53][28] ,
         \Inst_Mem/inst_mem_reg[53][29] , \Inst_Mem/inst_mem_reg[53][30] ,
         \Inst_Mem/inst_mem_reg[53][31] , \Inst_Mem/inst_mem_reg[52][0] ,
         \Inst_Mem/inst_mem_reg[52][1] , \Inst_Mem/inst_mem_reg[52][2] ,
         \Inst_Mem/inst_mem_reg[52][3] , \Inst_Mem/inst_mem_reg[52][4] ,
         \Inst_Mem/inst_mem_reg[52][5] , \Inst_Mem/inst_mem_reg[52][6] ,
         \Inst_Mem/inst_mem_reg[52][7] , \Inst_Mem/inst_mem_reg[52][8] ,
         \Inst_Mem/inst_mem_reg[52][9] , \Inst_Mem/inst_mem_reg[52][10] ,
         \Inst_Mem/inst_mem_reg[52][11] , \Inst_Mem/inst_mem_reg[52][12] ,
         \Inst_Mem/inst_mem_reg[52][13] , \Inst_Mem/inst_mem_reg[52][14] ,
         \Inst_Mem/inst_mem_reg[52][15] , \Inst_Mem/inst_mem_reg[52][16] ,
         \Inst_Mem/inst_mem_reg[52][17] , \Inst_Mem/inst_mem_reg[52][18] ,
         \Inst_Mem/inst_mem_reg[52][19] , \Inst_Mem/inst_mem_reg[52][20] ,
         \Inst_Mem/inst_mem_reg[52][21] , \Inst_Mem/inst_mem_reg[52][22] ,
         \Inst_Mem/inst_mem_reg[52][23] , \Inst_Mem/inst_mem_reg[52][24] ,
         \Inst_Mem/inst_mem_reg[52][25] , \Inst_Mem/inst_mem_reg[52][26] ,
         \Inst_Mem/inst_mem_reg[52][27] , \Inst_Mem/inst_mem_reg[52][28] ,
         \Inst_Mem/inst_mem_reg[52][29] , \Inst_Mem/inst_mem_reg[52][30] ,
         \Inst_Mem/inst_mem_reg[52][31] , \Inst_Mem/inst_mem_reg[51][0] ,
         \Inst_Mem/inst_mem_reg[51][1] , \Inst_Mem/inst_mem_reg[51][2] ,
         \Inst_Mem/inst_mem_reg[51][3] , \Inst_Mem/inst_mem_reg[51][4] ,
         \Inst_Mem/inst_mem_reg[51][5] , \Inst_Mem/inst_mem_reg[51][6] ,
         \Inst_Mem/inst_mem_reg[51][7] , \Inst_Mem/inst_mem_reg[51][8] ,
         \Inst_Mem/inst_mem_reg[51][9] , \Inst_Mem/inst_mem_reg[51][10] ,
         \Inst_Mem/inst_mem_reg[51][11] , \Inst_Mem/inst_mem_reg[51][12] ,
         \Inst_Mem/inst_mem_reg[51][13] , \Inst_Mem/inst_mem_reg[51][14] ,
         \Inst_Mem/inst_mem_reg[51][15] , \Inst_Mem/inst_mem_reg[51][16] ,
         \Inst_Mem/inst_mem_reg[51][17] , \Inst_Mem/inst_mem_reg[51][18] ,
         \Inst_Mem/inst_mem_reg[51][19] , \Inst_Mem/inst_mem_reg[51][20] ,
         \Inst_Mem/inst_mem_reg[51][21] , \Inst_Mem/inst_mem_reg[51][22] ,
         \Inst_Mem/inst_mem_reg[51][23] , \Inst_Mem/inst_mem_reg[51][24] ,
         \Inst_Mem/inst_mem_reg[51][25] , \Inst_Mem/inst_mem_reg[51][26] ,
         \Inst_Mem/inst_mem_reg[51][27] , \Inst_Mem/inst_mem_reg[51][28] ,
         \Inst_Mem/inst_mem_reg[51][29] , \Inst_Mem/inst_mem_reg[51][30] ,
         \Inst_Mem/inst_mem_reg[51][31] , \Inst_Mem/inst_mem_reg[50][0] ,
         \Inst_Mem/inst_mem_reg[50][1] , \Inst_Mem/inst_mem_reg[50][2] ,
         \Inst_Mem/inst_mem_reg[50][3] , \Inst_Mem/inst_mem_reg[50][4] ,
         \Inst_Mem/inst_mem_reg[50][5] , \Inst_Mem/inst_mem_reg[50][6] ,
         \Inst_Mem/inst_mem_reg[50][7] , \Inst_Mem/inst_mem_reg[50][8] ,
         \Inst_Mem/inst_mem_reg[50][9] , \Inst_Mem/inst_mem_reg[50][10] ,
         \Inst_Mem/inst_mem_reg[50][11] , \Inst_Mem/inst_mem_reg[50][12] ,
         \Inst_Mem/inst_mem_reg[50][13] , \Inst_Mem/inst_mem_reg[50][14] ,
         \Inst_Mem/inst_mem_reg[50][15] , \Inst_Mem/inst_mem_reg[50][16] ,
         \Inst_Mem/inst_mem_reg[50][17] , \Inst_Mem/inst_mem_reg[50][18] ,
         \Inst_Mem/inst_mem_reg[50][19] , \Inst_Mem/inst_mem_reg[50][20] ,
         \Inst_Mem/inst_mem_reg[50][21] , \Inst_Mem/inst_mem_reg[50][22] ,
         \Inst_Mem/inst_mem_reg[50][23] , \Inst_Mem/inst_mem_reg[50][24] ,
         \Inst_Mem/inst_mem_reg[50][25] , \Inst_Mem/inst_mem_reg[50][26] ,
         \Inst_Mem/inst_mem_reg[50][27] , \Inst_Mem/inst_mem_reg[50][28] ,
         \Inst_Mem/inst_mem_reg[50][29] , \Inst_Mem/inst_mem_reg[50][30] ,
         \Inst_Mem/inst_mem_reg[50][31] , \Inst_Mem/inst_mem_reg[49][0] ,
         \Inst_Mem/inst_mem_reg[49][1] , \Inst_Mem/inst_mem_reg[49][2] ,
         \Inst_Mem/inst_mem_reg[49][3] , \Inst_Mem/inst_mem_reg[49][4] ,
         \Inst_Mem/inst_mem_reg[49][5] , \Inst_Mem/inst_mem_reg[49][6] ,
         \Inst_Mem/inst_mem_reg[49][7] , \Inst_Mem/inst_mem_reg[49][8] ,
         \Inst_Mem/inst_mem_reg[49][9] , \Inst_Mem/inst_mem_reg[49][10] ,
         \Inst_Mem/inst_mem_reg[49][11] , \Inst_Mem/inst_mem_reg[49][12] ,
         \Inst_Mem/inst_mem_reg[49][13] , \Inst_Mem/inst_mem_reg[49][14] ,
         \Inst_Mem/inst_mem_reg[49][15] , \Inst_Mem/inst_mem_reg[49][16] ,
         \Inst_Mem/inst_mem_reg[49][17] , \Inst_Mem/inst_mem_reg[49][18] ,
         \Inst_Mem/inst_mem_reg[49][19] , \Inst_Mem/inst_mem_reg[49][20] ,
         \Inst_Mem/inst_mem_reg[49][21] , \Inst_Mem/inst_mem_reg[49][22] ,
         \Inst_Mem/inst_mem_reg[49][23] , \Inst_Mem/inst_mem_reg[49][24] ,
         \Inst_Mem/inst_mem_reg[49][25] , \Inst_Mem/inst_mem_reg[49][26] ,
         \Inst_Mem/inst_mem_reg[49][27] , \Inst_Mem/inst_mem_reg[49][28] ,
         \Inst_Mem/inst_mem_reg[49][29] , \Inst_Mem/inst_mem_reg[49][30] ,
         \Inst_Mem/inst_mem_reg[49][31] , \Inst_Mem/inst_mem_reg[48][0] ,
         \Inst_Mem/inst_mem_reg[48][1] , \Inst_Mem/inst_mem_reg[48][2] ,
         \Inst_Mem/inst_mem_reg[48][3] , \Inst_Mem/inst_mem_reg[48][4] ,
         \Inst_Mem/inst_mem_reg[48][5] , \Inst_Mem/inst_mem_reg[48][6] ,
         \Inst_Mem/inst_mem_reg[48][7] , \Inst_Mem/inst_mem_reg[48][8] ,
         \Inst_Mem/inst_mem_reg[48][9] , \Inst_Mem/inst_mem_reg[48][10] ,
         \Inst_Mem/inst_mem_reg[48][11] , \Inst_Mem/inst_mem_reg[48][12] ,
         \Inst_Mem/inst_mem_reg[48][13] , \Inst_Mem/inst_mem_reg[48][14] ,
         \Inst_Mem/inst_mem_reg[48][15] , \Inst_Mem/inst_mem_reg[48][16] ,
         \Inst_Mem/inst_mem_reg[48][17] , \Inst_Mem/inst_mem_reg[48][18] ,
         \Inst_Mem/inst_mem_reg[48][19] , \Inst_Mem/inst_mem_reg[48][20] ,
         \Inst_Mem/inst_mem_reg[48][21] , \Inst_Mem/inst_mem_reg[48][22] ,
         \Inst_Mem/inst_mem_reg[48][23] , \Inst_Mem/inst_mem_reg[48][24] ,
         \Inst_Mem/inst_mem_reg[48][25] , \Inst_Mem/inst_mem_reg[48][26] ,
         \Inst_Mem/inst_mem_reg[48][27] , \Inst_Mem/inst_mem_reg[48][28] ,
         \Inst_Mem/inst_mem_reg[48][29] , \Inst_Mem/inst_mem_reg[48][30] ,
         \Inst_Mem/inst_mem_reg[48][31] , \Inst_Mem/inst_mem_reg[47][0] ,
         \Inst_Mem/inst_mem_reg[47][1] , \Inst_Mem/inst_mem_reg[47][2] ,
         \Inst_Mem/inst_mem_reg[47][3] , \Inst_Mem/inst_mem_reg[47][4] ,
         \Inst_Mem/inst_mem_reg[47][5] , \Inst_Mem/inst_mem_reg[47][6] ,
         \Inst_Mem/inst_mem_reg[47][7] , \Inst_Mem/inst_mem_reg[47][8] ,
         \Inst_Mem/inst_mem_reg[47][9] , \Inst_Mem/inst_mem_reg[47][10] ,
         \Inst_Mem/inst_mem_reg[47][11] , \Inst_Mem/inst_mem_reg[47][12] ,
         \Inst_Mem/inst_mem_reg[47][13] , \Inst_Mem/inst_mem_reg[47][14] ,
         \Inst_Mem/inst_mem_reg[47][15] , \Inst_Mem/inst_mem_reg[47][16] ,
         \Inst_Mem/inst_mem_reg[47][17] , \Inst_Mem/inst_mem_reg[47][18] ,
         \Inst_Mem/inst_mem_reg[47][19] , \Inst_Mem/inst_mem_reg[47][20] ,
         \Inst_Mem/inst_mem_reg[47][21] , \Inst_Mem/inst_mem_reg[47][22] ,
         \Inst_Mem/inst_mem_reg[47][23] , \Inst_Mem/inst_mem_reg[47][24] ,
         \Inst_Mem/inst_mem_reg[47][25] , \Inst_Mem/inst_mem_reg[47][26] ,
         \Inst_Mem/inst_mem_reg[47][27] , \Inst_Mem/inst_mem_reg[47][28] ,
         \Inst_Mem/inst_mem_reg[47][29] , \Inst_Mem/inst_mem_reg[47][30] ,
         \Inst_Mem/inst_mem_reg[47][31] , \Inst_Mem/inst_mem_reg[46][0] ,
         \Inst_Mem/inst_mem_reg[46][1] , \Inst_Mem/inst_mem_reg[46][2] ,
         \Inst_Mem/inst_mem_reg[46][3] , \Inst_Mem/inst_mem_reg[46][4] ,
         \Inst_Mem/inst_mem_reg[46][5] , \Inst_Mem/inst_mem_reg[46][6] ,
         \Inst_Mem/inst_mem_reg[46][7] , \Inst_Mem/inst_mem_reg[46][8] ,
         \Inst_Mem/inst_mem_reg[46][9] , \Inst_Mem/inst_mem_reg[46][10] ,
         \Inst_Mem/inst_mem_reg[46][11] , \Inst_Mem/inst_mem_reg[46][12] ,
         \Inst_Mem/inst_mem_reg[46][13] , \Inst_Mem/inst_mem_reg[46][14] ,
         \Inst_Mem/inst_mem_reg[46][15] , \Inst_Mem/inst_mem_reg[46][16] ,
         \Inst_Mem/inst_mem_reg[46][17] , \Inst_Mem/inst_mem_reg[46][18] ,
         \Inst_Mem/inst_mem_reg[46][19] , \Inst_Mem/inst_mem_reg[46][20] ,
         \Inst_Mem/inst_mem_reg[46][21] , \Inst_Mem/inst_mem_reg[46][22] ,
         \Inst_Mem/inst_mem_reg[46][23] , \Inst_Mem/inst_mem_reg[46][24] ,
         \Inst_Mem/inst_mem_reg[46][25] , \Inst_Mem/inst_mem_reg[46][26] ,
         \Inst_Mem/inst_mem_reg[46][27] , \Inst_Mem/inst_mem_reg[46][28] ,
         \Inst_Mem/inst_mem_reg[46][29] , \Inst_Mem/inst_mem_reg[46][30] ,
         \Inst_Mem/inst_mem_reg[46][31] , \Inst_Mem/inst_mem_reg[45][0] ,
         \Inst_Mem/inst_mem_reg[45][1] , \Inst_Mem/inst_mem_reg[45][2] ,
         \Inst_Mem/inst_mem_reg[45][3] , \Inst_Mem/inst_mem_reg[45][4] ,
         \Inst_Mem/inst_mem_reg[45][5] , \Inst_Mem/inst_mem_reg[45][6] ,
         \Inst_Mem/inst_mem_reg[45][7] , \Inst_Mem/inst_mem_reg[45][8] ,
         \Inst_Mem/inst_mem_reg[45][9] , \Inst_Mem/inst_mem_reg[45][10] ,
         \Inst_Mem/inst_mem_reg[45][11] , \Inst_Mem/inst_mem_reg[45][12] ,
         \Inst_Mem/inst_mem_reg[45][13] , \Inst_Mem/inst_mem_reg[45][14] ,
         \Inst_Mem/inst_mem_reg[45][15] , \Inst_Mem/inst_mem_reg[45][16] ,
         \Inst_Mem/inst_mem_reg[45][17] , \Inst_Mem/inst_mem_reg[45][18] ,
         \Inst_Mem/inst_mem_reg[45][19] , \Inst_Mem/inst_mem_reg[45][20] ,
         \Inst_Mem/inst_mem_reg[45][21] , \Inst_Mem/inst_mem_reg[45][22] ,
         \Inst_Mem/inst_mem_reg[45][23] , \Inst_Mem/inst_mem_reg[45][24] ,
         \Inst_Mem/inst_mem_reg[45][25] , \Inst_Mem/inst_mem_reg[45][26] ,
         \Inst_Mem/inst_mem_reg[45][27] , \Inst_Mem/inst_mem_reg[45][28] ,
         \Inst_Mem/inst_mem_reg[45][29] , \Inst_Mem/inst_mem_reg[45][30] ,
         \Inst_Mem/inst_mem_reg[45][31] , \Inst_Mem/inst_mem_reg[44][0] ,
         \Inst_Mem/inst_mem_reg[44][1] , \Inst_Mem/inst_mem_reg[44][2] ,
         \Inst_Mem/inst_mem_reg[44][3] , \Inst_Mem/inst_mem_reg[44][4] ,
         \Inst_Mem/inst_mem_reg[44][5] , \Inst_Mem/inst_mem_reg[44][6] ,
         \Inst_Mem/inst_mem_reg[44][7] , \Inst_Mem/inst_mem_reg[44][8] ,
         \Inst_Mem/inst_mem_reg[44][9] , \Inst_Mem/inst_mem_reg[44][10] ,
         \Inst_Mem/inst_mem_reg[44][11] , \Inst_Mem/inst_mem_reg[44][12] ,
         \Inst_Mem/inst_mem_reg[44][13] , \Inst_Mem/inst_mem_reg[44][14] ,
         \Inst_Mem/inst_mem_reg[44][15] , \Inst_Mem/inst_mem_reg[44][16] ,
         \Inst_Mem/inst_mem_reg[44][17] , \Inst_Mem/inst_mem_reg[44][18] ,
         \Inst_Mem/inst_mem_reg[44][19] , \Inst_Mem/inst_mem_reg[44][20] ,
         \Inst_Mem/inst_mem_reg[44][21] , \Inst_Mem/inst_mem_reg[44][22] ,
         \Inst_Mem/inst_mem_reg[44][23] , \Inst_Mem/inst_mem_reg[44][24] ,
         \Inst_Mem/inst_mem_reg[44][25] , \Inst_Mem/inst_mem_reg[44][26] ,
         \Inst_Mem/inst_mem_reg[44][27] , \Inst_Mem/inst_mem_reg[44][28] ,
         \Inst_Mem/inst_mem_reg[44][29] , \Inst_Mem/inst_mem_reg[44][30] ,
         \Inst_Mem/inst_mem_reg[44][31] , \Inst_Mem/inst_mem_reg[43][0] ,
         \Inst_Mem/inst_mem_reg[43][1] , \Inst_Mem/inst_mem_reg[43][2] ,
         \Inst_Mem/inst_mem_reg[43][3] , \Inst_Mem/inst_mem_reg[43][4] ,
         \Inst_Mem/inst_mem_reg[43][5] , \Inst_Mem/inst_mem_reg[43][6] ,
         \Inst_Mem/inst_mem_reg[43][7] , \Inst_Mem/inst_mem_reg[43][8] ,
         \Inst_Mem/inst_mem_reg[43][9] , \Inst_Mem/inst_mem_reg[43][10] ,
         \Inst_Mem/inst_mem_reg[43][11] , \Inst_Mem/inst_mem_reg[43][12] ,
         \Inst_Mem/inst_mem_reg[43][13] , \Inst_Mem/inst_mem_reg[43][14] ,
         \Inst_Mem/inst_mem_reg[43][15] , \Inst_Mem/inst_mem_reg[43][16] ,
         \Inst_Mem/inst_mem_reg[43][17] , \Inst_Mem/inst_mem_reg[43][18] ,
         \Inst_Mem/inst_mem_reg[43][19] , \Inst_Mem/inst_mem_reg[43][20] ,
         \Inst_Mem/inst_mem_reg[43][21] , \Inst_Mem/inst_mem_reg[43][22] ,
         \Inst_Mem/inst_mem_reg[43][23] , \Inst_Mem/inst_mem_reg[43][24] ,
         \Inst_Mem/inst_mem_reg[43][25] , \Inst_Mem/inst_mem_reg[43][26] ,
         \Inst_Mem/inst_mem_reg[43][27] , \Inst_Mem/inst_mem_reg[43][28] ,
         \Inst_Mem/inst_mem_reg[43][29] , \Inst_Mem/inst_mem_reg[43][30] ,
         \Inst_Mem/inst_mem_reg[43][31] , \Inst_Mem/inst_mem_reg[42][0] ,
         \Inst_Mem/inst_mem_reg[42][1] , \Inst_Mem/inst_mem_reg[42][2] ,
         \Inst_Mem/inst_mem_reg[42][3] , \Inst_Mem/inst_mem_reg[42][4] ,
         \Inst_Mem/inst_mem_reg[42][5] , \Inst_Mem/inst_mem_reg[42][6] ,
         \Inst_Mem/inst_mem_reg[42][7] , \Inst_Mem/inst_mem_reg[42][8] ,
         \Inst_Mem/inst_mem_reg[42][9] , \Inst_Mem/inst_mem_reg[42][10] ,
         \Inst_Mem/inst_mem_reg[42][11] , \Inst_Mem/inst_mem_reg[42][12] ,
         \Inst_Mem/inst_mem_reg[42][13] , \Inst_Mem/inst_mem_reg[42][14] ,
         \Inst_Mem/inst_mem_reg[42][15] , \Inst_Mem/inst_mem_reg[42][16] ,
         \Inst_Mem/inst_mem_reg[42][17] , \Inst_Mem/inst_mem_reg[42][18] ,
         \Inst_Mem/inst_mem_reg[42][19] , \Inst_Mem/inst_mem_reg[42][20] ,
         \Inst_Mem/inst_mem_reg[42][21] , \Inst_Mem/inst_mem_reg[42][22] ,
         \Inst_Mem/inst_mem_reg[42][23] , \Inst_Mem/inst_mem_reg[42][24] ,
         \Inst_Mem/inst_mem_reg[42][25] , \Inst_Mem/inst_mem_reg[42][26] ,
         \Inst_Mem/inst_mem_reg[42][27] , \Inst_Mem/inst_mem_reg[42][28] ,
         \Inst_Mem/inst_mem_reg[42][29] , \Inst_Mem/inst_mem_reg[42][30] ,
         \Inst_Mem/inst_mem_reg[42][31] , \Inst_Mem/inst_mem_reg[41][0] ,
         \Inst_Mem/inst_mem_reg[41][1] , \Inst_Mem/inst_mem_reg[41][2] ,
         \Inst_Mem/inst_mem_reg[41][3] , \Inst_Mem/inst_mem_reg[41][4] ,
         \Inst_Mem/inst_mem_reg[41][5] , \Inst_Mem/inst_mem_reg[41][6] ,
         \Inst_Mem/inst_mem_reg[41][7] , \Inst_Mem/inst_mem_reg[41][8] ,
         \Inst_Mem/inst_mem_reg[41][9] , \Inst_Mem/inst_mem_reg[41][10] ,
         \Inst_Mem/inst_mem_reg[41][11] , \Inst_Mem/inst_mem_reg[41][12] ,
         \Inst_Mem/inst_mem_reg[41][13] , \Inst_Mem/inst_mem_reg[41][14] ,
         \Inst_Mem/inst_mem_reg[41][15] , \Inst_Mem/inst_mem_reg[41][16] ,
         \Inst_Mem/inst_mem_reg[41][17] , \Inst_Mem/inst_mem_reg[41][18] ,
         \Inst_Mem/inst_mem_reg[41][19] , \Inst_Mem/inst_mem_reg[41][20] ,
         \Inst_Mem/inst_mem_reg[41][21] , \Inst_Mem/inst_mem_reg[41][22] ,
         \Inst_Mem/inst_mem_reg[41][23] , \Inst_Mem/inst_mem_reg[41][24] ,
         \Inst_Mem/inst_mem_reg[41][25] , \Inst_Mem/inst_mem_reg[41][26] ,
         \Inst_Mem/inst_mem_reg[41][27] , \Inst_Mem/inst_mem_reg[41][28] ,
         \Inst_Mem/inst_mem_reg[41][29] , \Inst_Mem/inst_mem_reg[41][30] ,
         \Inst_Mem/inst_mem_reg[41][31] , \Inst_Mem/inst_mem_reg[40][0] ,
         \Inst_Mem/inst_mem_reg[40][1] , \Inst_Mem/inst_mem_reg[40][2] ,
         \Inst_Mem/inst_mem_reg[40][3] , \Inst_Mem/inst_mem_reg[40][4] ,
         \Inst_Mem/inst_mem_reg[40][5] , \Inst_Mem/inst_mem_reg[40][6] ,
         \Inst_Mem/inst_mem_reg[40][7] , \Inst_Mem/inst_mem_reg[40][8] ,
         \Inst_Mem/inst_mem_reg[40][9] , \Inst_Mem/inst_mem_reg[40][10] ,
         \Inst_Mem/inst_mem_reg[40][11] , \Inst_Mem/inst_mem_reg[40][12] ,
         \Inst_Mem/inst_mem_reg[40][13] , \Inst_Mem/inst_mem_reg[40][14] ,
         \Inst_Mem/inst_mem_reg[40][15] , \Inst_Mem/inst_mem_reg[40][16] ,
         \Inst_Mem/inst_mem_reg[40][17] , \Inst_Mem/inst_mem_reg[40][18] ,
         \Inst_Mem/inst_mem_reg[40][19] , \Inst_Mem/inst_mem_reg[40][20] ,
         \Inst_Mem/inst_mem_reg[40][21] , \Inst_Mem/inst_mem_reg[40][22] ,
         \Inst_Mem/inst_mem_reg[40][23] , \Inst_Mem/inst_mem_reg[40][24] ,
         \Inst_Mem/inst_mem_reg[40][25] , \Inst_Mem/inst_mem_reg[40][26] ,
         \Inst_Mem/inst_mem_reg[40][27] , \Inst_Mem/inst_mem_reg[40][28] ,
         \Inst_Mem/inst_mem_reg[40][29] , \Inst_Mem/inst_mem_reg[40][30] ,
         \Inst_Mem/inst_mem_reg[40][31] , \Inst_Mem/inst_mem_reg[39][0] ,
         \Inst_Mem/inst_mem_reg[39][1] , \Inst_Mem/inst_mem_reg[39][2] ,
         \Inst_Mem/inst_mem_reg[39][3] , \Inst_Mem/inst_mem_reg[39][4] ,
         \Inst_Mem/inst_mem_reg[39][5] , \Inst_Mem/inst_mem_reg[39][6] ,
         \Inst_Mem/inst_mem_reg[39][7] , \Inst_Mem/inst_mem_reg[39][8] ,
         \Inst_Mem/inst_mem_reg[39][9] , \Inst_Mem/inst_mem_reg[39][10] ,
         \Inst_Mem/inst_mem_reg[39][11] , \Inst_Mem/inst_mem_reg[39][12] ,
         \Inst_Mem/inst_mem_reg[39][13] , \Inst_Mem/inst_mem_reg[39][14] ,
         \Inst_Mem/inst_mem_reg[39][15] , \Inst_Mem/inst_mem_reg[39][16] ,
         \Inst_Mem/inst_mem_reg[39][17] , \Inst_Mem/inst_mem_reg[39][18] ,
         \Inst_Mem/inst_mem_reg[39][19] , \Inst_Mem/inst_mem_reg[39][20] ,
         \Inst_Mem/inst_mem_reg[39][21] , \Inst_Mem/inst_mem_reg[39][22] ,
         \Inst_Mem/inst_mem_reg[39][23] , \Inst_Mem/inst_mem_reg[39][24] ,
         \Inst_Mem/inst_mem_reg[39][25] , \Inst_Mem/inst_mem_reg[39][26] ,
         \Inst_Mem/inst_mem_reg[39][27] , \Inst_Mem/inst_mem_reg[39][28] ,
         \Inst_Mem/inst_mem_reg[39][29] , \Inst_Mem/inst_mem_reg[39][30] ,
         \Inst_Mem/inst_mem_reg[39][31] , \Inst_Mem/inst_mem_reg[38][0] ,
         \Inst_Mem/inst_mem_reg[38][1] , \Inst_Mem/inst_mem_reg[38][2] ,
         \Inst_Mem/inst_mem_reg[38][3] , \Inst_Mem/inst_mem_reg[38][4] ,
         \Inst_Mem/inst_mem_reg[38][5] , \Inst_Mem/inst_mem_reg[38][6] ,
         \Inst_Mem/inst_mem_reg[38][7] , \Inst_Mem/inst_mem_reg[38][8] ,
         \Inst_Mem/inst_mem_reg[38][9] , \Inst_Mem/inst_mem_reg[38][10] ,
         \Inst_Mem/inst_mem_reg[38][11] , \Inst_Mem/inst_mem_reg[38][12] ,
         \Inst_Mem/inst_mem_reg[38][13] , \Inst_Mem/inst_mem_reg[38][14] ,
         \Inst_Mem/inst_mem_reg[38][15] , \Inst_Mem/inst_mem_reg[38][16] ,
         \Inst_Mem/inst_mem_reg[38][17] , \Inst_Mem/inst_mem_reg[38][18] ,
         \Inst_Mem/inst_mem_reg[38][19] , \Inst_Mem/inst_mem_reg[38][20] ,
         \Inst_Mem/inst_mem_reg[38][21] , \Inst_Mem/inst_mem_reg[38][22] ,
         \Inst_Mem/inst_mem_reg[38][23] , \Inst_Mem/inst_mem_reg[38][24] ,
         \Inst_Mem/inst_mem_reg[38][25] , \Inst_Mem/inst_mem_reg[38][26] ,
         \Inst_Mem/inst_mem_reg[38][27] , \Inst_Mem/inst_mem_reg[38][28] ,
         \Inst_Mem/inst_mem_reg[38][29] , \Inst_Mem/inst_mem_reg[38][30] ,
         \Inst_Mem/inst_mem_reg[38][31] , \Inst_Mem/inst_mem_reg[37][0] ,
         \Inst_Mem/inst_mem_reg[37][1] , \Inst_Mem/inst_mem_reg[37][2] ,
         \Inst_Mem/inst_mem_reg[37][3] , \Inst_Mem/inst_mem_reg[37][4] ,
         \Inst_Mem/inst_mem_reg[37][5] , \Inst_Mem/inst_mem_reg[37][6] ,
         \Inst_Mem/inst_mem_reg[37][7] , \Inst_Mem/inst_mem_reg[37][8] ,
         \Inst_Mem/inst_mem_reg[37][9] , \Inst_Mem/inst_mem_reg[37][10] ,
         \Inst_Mem/inst_mem_reg[37][11] , \Inst_Mem/inst_mem_reg[37][12] ,
         \Inst_Mem/inst_mem_reg[37][13] , \Inst_Mem/inst_mem_reg[37][14] ,
         \Inst_Mem/inst_mem_reg[37][15] , \Inst_Mem/inst_mem_reg[37][16] ,
         \Inst_Mem/inst_mem_reg[37][17] , \Inst_Mem/inst_mem_reg[37][18] ,
         \Inst_Mem/inst_mem_reg[37][19] , \Inst_Mem/inst_mem_reg[37][20] ,
         \Inst_Mem/inst_mem_reg[37][21] , \Inst_Mem/inst_mem_reg[37][22] ,
         \Inst_Mem/inst_mem_reg[37][23] , \Inst_Mem/inst_mem_reg[37][24] ,
         \Inst_Mem/inst_mem_reg[37][25] , \Inst_Mem/inst_mem_reg[37][26] ,
         \Inst_Mem/inst_mem_reg[37][27] , \Inst_Mem/inst_mem_reg[37][28] ,
         \Inst_Mem/inst_mem_reg[37][29] , \Inst_Mem/inst_mem_reg[37][30] ,
         \Inst_Mem/inst_mem_reg[37][31] , \Inst_Mem/inst_mem_reg[36][0] ,
         \Inst_Mem/inst_mem_reg[36][1] , \Inst_Mem/inst_mem_reg[36][2] ,
         \Inst_Mem/inst_mem_reg[36][3] , \Inst_Mem/inst_mem_reg[36][4] ,
         \Inst_Mem/inst_mem_reg[36][5] , \Inst_Mem/inst_mem_reg[36][6] ,
         \Inst_Mem/inst_mem_reg[36][7] , \Inst_Mem/inst_mem_reg[36][8] ,
         \Inst_Mem/inst_mem_reg[36][9] , \Inst_Mem/inst_mem_reg[36][10] ,
         \Inst_Mem/inst_mem_reg[36][11] , \Inst_Mem/inst_mem_reg[36][12] ,
         \Inst_Mem/inst_mem_reg[36][13] , \Inst_Mem/inst_mem_reg[36][14] ,
         \Inst_Mem/inst_mem_reg[36][15] , \Inst_Mem/inst_mem_reg[36][16] ,
         \Inst_Mem/inst_mem_reg[36][17] , \Inst_Mem/inst_mem_reg[36][18] ,
         \Inst_Mem/inst_mem_reg[36][19] , \Inst_Mem/inst_mem_reg[36][20] ,
         \Inst_Mem/inst_mem_reg[36][21] , \Inst_Mem/inst_mem_reg[36][22] ,
         \Inst_Mem/inst_mem_reg[36][23] , \Inst_Mem/inst_mem_reg[36][24] ,
         \Inst_Mem/inst_mem_reg[36][25] , \Inst_Mem/inst_mem_reg[36][26] ,
         \Inst_Mem/inst_mem_reg[36][27] , \Inst_Mem/inst_mem_reg[36][28] ,
         \Inst_Mem/inst_mem_reg[36][29] , \Inst_Mem/inst_mem_reg[36][30] ,
         \Inst_Mem/inst_mem_reg[36][31] , \Inst_Mem/inst_mem_reg[35][0] ,
         \Inst_Mem/inst_mem_reg[35][1] , \Inst_Mem/inst_mem_reg[35][2] ,
         \Inst_Mem/inst_mem_reg[35][3] , \Inst_Mem/inst_mem_reg[35][4] ,
         \Inst_Mem/inst_mem_reg[35][5] , \Inst_Mem/inst_mem_reg[35][6] ,
         \Inst_Mem/inst_mem_reg[35][7] , \Inst_Mem/inst_mem_reg[35][8] ,
         \Inst_Mem/inst_mem_reg[35][9] , \Inst_Mem/inst_mem_reg[35][10] ,
         \Inst_Mem/inst_mem_reg[35][11] , \Inst_Mem/inst_mem_reg[35][12] ,
         \Inst_Mem/inst_mem_reg[35][13] , \Inst_Mem/inst_mem_reg[35][14] ,
         \Inst_Mem/inst_mem_reg[35][15] , \Inst_Mem/inst_mem_reg[35][16] ,
         \Inst_Mem/inst_mem_reg[35][17] , \Inst_Mem/inst_mem_reg[35][18] ,
         \Inst_Mem/inst_mem_reg[35][19] , \Inst_Mem/inst_mem_reg[35][20] ,
         \Inst_Mem/inst_mem_reg[35][21] , \Inst_Mem/inst_mem_reg[35][22] ,
         \Inst_Mem/inst_mem_reg[35][23] , \Inst_Mem/inst_mem_reg[35][24] ,
         \Inst_Mem/inst_mem_reg[35][25] , \Inst_Mem/inst_mem_reg[35][26] ,
         \Inst_Mem/inst_mem_reg[35][27] , \Inst_Mem/inst_mem_reg[35][28] ,
         \Inst_Mem/inst_mem_reg[35][29] , \Inst_Mem/inst_mem_reg[35][30] ,
         \Inst_Mem/inst_mem_reg[35][31] , \Inst_Mem/inst_mem_reg[34][0] ,
         \Inst_Mem/inst_mem_reg[34][1] , \Inst_Mem/inst_mem_reg[34][2] ,
         \Inst_Mem/inst_mem_reg[34][3] , \Inst_Mem/inst_mem_reg[34][4] ,
         \Inst_Mem/inst_mem_reg[34][5] , \Inst_Mem/inst_mem_reg[34][6] ,
         \Inst_Mem/inst_mem_reg[34][7] , \Inst_Mem/inst_mem_reg[34][8] ,
         \Inst_Mem/inst_mem_reg[34][9] , \Inst_Mem/inst_mem_reg[34][10] ,
         \Inst_Mem/inst_mem_reg[34][11] , \Inst_Mem/inst_mem_reg[34][12] ,
         \Inst_Mem/inst_mem_reg[34][13] , \Inst_Mem/inst_mem_reg[34][14] ,
         \Inst_Mem/inst_mem_reg[34][15] , \Inst_Mem/inst_mem_reg[34][16] ,
         \Inst_Mem/inst_mem_reg[34][17] , \Inst_Mem/inst_mem_reg[34][18] ,
         \Inst_Mem/inst_mem_reg[34][19] , \Inst_Mem/inst_mem_reg[34][20] ,
         \Inst_Mem/inst_mem_reg[34][21] , \Inst_Mem/inst_mem_reg[34][22] ,
         \Inst_Mem/inst_mem_reg[34][23] , \Inst_Mem/inst_mem_reg[34][24] ,
         \Inst_Mem/inst_mem_reg[34][25] , \Inst_Mem/inst_mem_reg[34][26] ,
         \Inst_Mem/inst_mem_reg[34][27] , \Inst_Mem/inst_mem_reg[34][28] ,
         \Inst_Mem/inst_mem_reg[34][29] , \Inst_Mem/inst_mem_reg[34][30] ,
         \Inst_Mem/inst_mem_reg[34][31] , \Inst_Mem/inst_mem_reg[33][0] ,
         \Inst_Mem/inst_mem_reg[33][1] , \Inst_Mem/inst_mem_reg[33][2] ,
         \Inst_Mem/inst_mem_reg[33][3] , \Inst_Mem/inst_mem_reg[33][4] ,
         \Inst_Mem/inst_mem_reg[33][5] , \Inst_Mem/inst_mem_reg[33][6] ,
         \Inst_Mem/inst_mem_reg[33][7] , \Inst_Mem/inst_mem_reg[33][8] ,
         \Inst_Mem/inst_mem_reg[33][9] , \Inst_Mem/inst_mem_reg[33][10] ,
         \Inst_Mem/inst_mem_reg[33][11] , \Inst_Mem/inst_mem_reg[33][12] ,
         \Inst_Mem/inst_mem_reg[33][13] , \Inst_Mem/inst_mem_reg[33][14] ,
         \Inst_Mem/inst_mem_reg[33][15] , \Inst_Mem/inst_mem_reg[33][16] ,
         \Inst_Mem/inst_mem_reg[33][17] , \Inst_Mem/inst_mem_reg[33][18] ,
         \Inst_Mem/inst_mem_reg[33][19] , \Inst_Mem/inst_mem_reg[33][20] ,
         \Inst_Mem/inst_mem_reg[33][21] , \Inst_Mem/inst_mem_reg[33][22] ,
         \Inst_Mem/inst_mem_reg[33][23] , \Inst_Mem/inst_mem_reg[33][24] ,
         \Inst_Mem/inst_mem_reg[33][25] , \Inst_Mem/inst_mem_reg[33][26] ,
         \Inst_Mem/inst_mem_reg[33][27] , \Inst_Mem/inst_mem_reg[33][28] ,
         \Inst_Mem/inst_mem_reg[33][29] , \Inst_Mem/inst_mem_reg[33][30] ,
         \Inst_Mem/inst_mem_reg[33][31] , \Inst_Mem/inst_mem_reg[32][0] ,
         \Inst_Mem/inst_mem_reg[32][1] , \Inst_Mem/inst_mem_reg[32][2] ,
         \Inst_Mem/inst_mem_reg[32][3] , \Inst_Mem/inst_mem_reg[32][4] ,
         \Inst_Mem/inst_mem_reg[32][5] , \Inst_Mem/inst_mem_reg[32][6] ,
         \Inst_Mem/inst_mem_reg[32][7] , \Inst_Mem/inst_mem_reg[32][8] ,
         \Inst_Mem/inst_mem_reg[32][9] , \Inst_Mem/inst_mem_reg[32][10] ,
         \Inst_Mem/inst_mem_reg[32][11] , \Inst_Mem/inst_mem_reg[32][12] ,
         \Inst_Mem/inst_mem_reg[32][13] , \Inst_Mem/inst_mem_reg[32][14] ,
         \Inst_Mem/inst_mem_reg[32][15] , \Inst_Mem/inst_mem_reg[32][16] ,
         \Inst_Mem/inst_mem_reg[32][17] , \Inst_Mem/inst_mem_reg[32][18] ,
         \Inst_Mem/inst_mem_reg[32][19] , \Inst_Mem/inst_mem_reg[32][20] ,
         \Inst_Mem/inst_mem_reg[32][21] , \Inst_Mem/inst_mem_reg[32][22] ,
         \Inst_Mem/inst_mem_reg[32][23] , \Inst_Mem/inst_mem_reg[32][24] ,
         \Inst_Mem/inst_mem_reg[32][25] , \Inst_Mem/inst_mem_reg[32][26] ,
         \Inst_Mem/inst_mem_reg[32][27] , \Inst_Mem/inst_mem_reg[32][28] ,
         \Inst_Mem/inst_mem_reg[32][29] , \Inst_Mem/inst_mem_reg[32][30] ,
         \Inst_Mem/inst_mem_reg[32][31] , \Inst_Mem/inst_mem_reg[31][0] ,
         \Inst_Mem/inst_mem_reg[31][1] , \Inst_Mem/inst_mem_reg[31][2] ,
         \Inst_Mem/inst_mem_reg[31][3] , \Inst_Mem/inst_mem_reg[31][4] ,
         \Inst_Mem/inst_mem_reg[31][5] , \Inst_Mem/inst_mem_reg[31][6] ,
         \Inst_Mem/inst_mem_reg[31][7] , \Inst_Mem/inst_mem_reg[31][8] ,
         \Inst_Mem/inst_mem_reg[31][9] , \Inst_Mem/inst_mem_reg[31][10] ,
         \Inst_Mem/inst_mem_reg[31][11] , \Inst_Mem/inst_mem_reg[31][12] ,
         \Inst_Mem/inst_mem_reg[31][13] , \Inst_Mem/inst_mem_reg[31][14] ,
         \Inst_Mem/inst_mem_reg[31][15] , \Inst_Mem/inst_mem_reg[31][16] ,
         \Inst_Mem/inst_mem_reg[31][17] , \Inst_Mem/inst_mem_reg[31][18] ,
         \Inst_Mem/inst_mem_reg[31][19] , \Inst_Mem/inst_mem_reg[31][20] ,
         \Inst_Mem/inst_mem_reg[31][21] , \Inst_Mem/inst_mem_reg[31][22] ,
         \Inst_Mem/inst_mem_reg[31][23] , \Inst_Mem/inst_mem_reg[31][24] ,
         \Inst_Mem/inst_mem_reg[31][25] , \Inst_Mem/inst_mem_reg[31][26] ,
         \Inst_Mem/inst_mem_reg[31][27] , \Inst_Mem/inst_mem_reg[31][28] ,
         \Inst_Mem/inst_mem_reg[31][29] , \Inst_Mem/inst_mem_reg[31][30] ,
         \Inst_Mem/inst_mem_reg[31][31] , \Inst_Mem/inst_mem_reg[30][0] ,
         \Inst_Mem/inst_mem_reg[30][1] , \Inst_Mem/inst_mem_reg[30][2] ,
         \Inst_Mem/inst_mem_reg[30][3] , \Inst_Mem/inst_mem_reg[30][4] ,
         \Inst_Mem/inst_mem_reg[30][5] , \Inst_Mem/inst_mem_reg[30][6] ,
         \Inst_Mem/inst_mem_reg[30][7] , \Inst_Mem/inst_mem_reg[30][8] ,
         \Inst_Mem/inst_mem_reg[30][9] , \Inst_Mem/inst_mem_reg[30][10] ,
         \Inst_Mem/inst_mem_reg[30][11] , \Inst_Mem/inst_mem_reg[30][12] ,
         \Inst_Mem/inst_mem_reg[30][13] , \Inst_Mem/inst_mem_reg[30][14] ,
         \Inst_Mem/inst_mem_reg[30][15] , \Inst_Mem/inst_mem_reg[30][16] ,
         \Inst_Mem/inst_mem_reg[30][17] , \Inst_Mem/inst_mem_reg[30][18] ,
         \Inst_Mem/inst_mem_reg[30][19] , \Inst_Mem/inst_mem_reg[30][20] ,
         \Inst_Mem/inst_mem_reg[30][21] , \Inst_Mem/inst_mem_reg[30][22] ,
         \Inst_Mem/inst_mem_reg[30][23] , \Inst_Mem/inst_mem_reg[30][24] ,
         \Inst_Mem/inst_mem_reg[30][25] , \Inst_Mem/inst_mem_reg[30][26] ,
         \Inst_Mem/inst_mem_reg[30][27] , \Inst_Mem/inst_mem_reg[30][28] ,
         \Inst_Mem/inst_mem_reg[30][29] , \Inst_Mem/inst_mem_reg[30][30] ,
         \Inst_Mem/inst_mem_reg[30][31] , \Inst_Mem/inst_mem_reg[29][0] ,
         \Inst_Mem/inst_mem_reg[29][1] , \Inst_Mem/inst_mem_reg[29][2] ,
         \Inst_Mem/inst_mem_reg[29][3] , \Inst_Mem/inst_mem_reg[29][4] ,
         \Inst_Mem/inst_mem_reg[29][5] , \Inst_Mem/inst_mem_reg[29][6] ,
         \Inst_Mem/inst_mem_reg[29][7] , \Inst_Mem/inst_mem_reg[29][8] ,
         \Inst_Mem/inst_mem_reg[29][9] , \Inst_Mem/inst_mem_reg[29][10] ,
         \Inst_Mem/inst_mem_reg[29][11] , \Inst_Mem/inst_mem_reg[29][12] ,
         \Inst_Mem/inst_mem_reg[29][13] , \Inst_Mem/inst_mem_reg[29][14] ,
         \Inst_Mem/inst_mem_reg[29][15] , \Inst_Mem/inst_mem_reg[29][16] ,
         \Inst_Mem/inst_mem_reg[29][17] , \Inst_Mem/inst_mem_reg[29][18] ,
         \Inst_Mem/inst_mem_reg[29][19] , \Inst_Mem/inst_mem_reg[29][20] ,
         \Inst_Mem/inst_mem_reg[29][21] , \Inst_Mem/inst_mem_reg[29][22] ,
         \Inst_Mem/inst_mem_reg[29][23] , \Inst_Mem/inst_mem_reg[29][24] ,
         \Inst_Mem/inst_mem_reg[29][25] , \Inst_Mem/inst_mem_reg[29][26] ,
         \Inst_Mem/inst_mem_reg[29][27] , \Inst_Mem/inst_mem_reg[29][28] ,
         \Inst_Mem/inst_mem_reg[29][29] , \Inst_Mem/inst_mem_reg[29][30] ,
         \Inst_Mem/inst_mem_reg[29][31] , \Inst_Mem/inst_mem_reg[28][0] ,
         \Inst_Mem/inst_mem_reg[28][1] , \Inst_Mem/inst_mem_reg[28][2] ,
         \Inst_Mem/inst_mem_reg[28][3] , \Inst_Mem/inst_mem_reg[28][4] ,
         \Inst_Mem/inst_mem_reg[28][5] , \Inst_Mem/inst_mem_reg[28][6] ,
         \Inst_Mem/inst_mem_reg[28][7] , \Inst_Mem/inst_mem_reg[28][8] ,
         \Inst_Mem/inst_mem_reg[28][9] , \Inst_Mem/inst_mem_reg[28][10] ,
         \Inst_Mem/inst_mem_reg[28][11] , \Inst_Mem/inst_mem_reg[28][12] ,
         \Inst_Mem/inst_mem_reg[28][13] , \Inst_Mem/inst_mem_reg[28][14] ,
         \Inst_Mem/inst_mem_reg[28][15] , \Inst_Mem/inst_mem_reg[28][16] ,
         \Inst_Mem/inst_mem_reg[28][17] , \Inst_Mem/inst_mem_reg[28][18] ,
         \Inst_Mem/inst_mem_reg[28][19] , \Inst_Mem/inst_mem_reg[28][20] ,
         \Inst_Mem/inst_mem_reg[28][21] , \Inst_Mem/inst_mem_reg[28][22] ,
         \Inst_Mem/inst_mem_reg[28][23] , \Inst_Mem/inst_mem_reg[28][24] ,
         \Inst_Mem/inst_mem_reg[28][25] , \Inst_Mem/inst_mem_reg[28][26] ,
         \Inst_Mem/inst_mem_reg[28][27] , \Inst_Mem/inst_mem_reg[28][28] ,
         \Inst_Mem/inst_mem_reg[28][29] , \Inst_Mem/inst_mem_reg[28][30] ,
         \Inst_Mem/inst_mem_reg[28][31] , \Inst_Mem/inst_mem_reg[27][0] ,
         \Inst_Mem/inst_mem_reg[27][1] , \Inst_Mem/inst_mem_reg[27][2] ,
         \Inst_Mem/inst_mem_reg[27][3] , \Inst_Mem/inst_mem_reg[27][4] ,
         \Inst_Mem/inst_mem_reg[27][5] , \Inst_Mem/inst_mem_reg[27][6] ,
         \Inst_Mem/inst_mem_reg[27][7] , \Inst_Mem/inst_mem_reg[27][8] ,
         \Inst_Mem/inst_mem_reg[27][9] , \Inst_Mem/inst_mem_reg[27][10] ,
         \Inst_Mem/inst_mem_reg[27][11] , \Inst_Mem/inst_mem_reg[27][12] ,
         \Inst_Mem/inst_mem_reg[27][13] , \Inst_Mem/inst_mem_reg[27][14] ,
         \Inst_Mem/inst_mem_reg[27][15] , \Inst_Mem/inst_mem_reg[27][16] ,
         \Inst_Mem/inst_mem_reg[27][17] , \Inst_Mem/inst_mem_reg[27][18] ,
         \Inst_Mem/inst_mem_reg[27][19] , \Inst_Mem/inst_mem_reg[27][20] ,
         \Inst_Mem/inst_mem_reg[27][21] , \Inst_Mem/inst_mem_reg[27][22] ,
         \Inst_Mem/inst_mem_reg[27][23] , \Inst_Mem/inst_mem_reg[27][24] ,
         \Inst_Mem/inst_mem_reg[27][25] , \Inst_Mem/inst_mem_reg[27][26] ,
         \Inst_Mem/inst_mem_reg[27][27] , \Inst_Mem/inst_mem_reg[27][28] ,
         \Inst_Mem/inst_mem_reg[27][29] , \Inst_Mem/inst_mem_reg[27][30] ,
         \Inst_Mem/inst_mem_reg[27][31] , \Inst_Mem/inst_mem_reg[26][0] ,
         \Inst_Mem/inst_mem_reg[26][1] , \Inst_Mem/inst_mem_reg[26][2] ,
         \Inst_Mem/inst_mem_reg[26][3] , \Inst_Mem/inst_mem_reg[26][4] ,
         \Inst_Mem/inst_mem_reg[26][5] , \Inst_Mem/inst_mem_reg[26][6] ,
         \Inst_Mem/inst_mem_reg[26][7] , \Inst_Mem/inst_mem_reg[26][8] ,
         \Inst_Mem/inst_mem_reg[26][9] , \Inst_Mem/inst_mem_reg[26][10] ,
         \Inst_Mem/inst_mem_reg[26][11] , \Inst_Mem/inst_mem_reg[26][12] ,
         \Inst_Mem/inst_mem_reg[26][13] , \Inst_Mem/inst_mem_reg[26][14] ,
         \Inst_Mem/inst_mem_reg[26][15] , \Inst_Mem/inst_mem_reg[26][16] ,
         \Inst_Mem/inst_mem_reg[26][17] , \Inst_Mem/inst_mem_reg[26][18] ,
         \Inst_Mem/inst_mem_reg[26][19] , \Inst_Mem/inst_mem_reg[26][20] ,
         \Inst_Mem/inst_mem_reg[26][21] , \Inst_Mem/inst_mem_reg[26][22] ,
         \Inst_Mem/inst_mem_reg[26][23] , \Inst_Mem/inst_mem_reg[26][24] ,
         \Inst_Mem/inst_mem_reg[26][25] , \Inst_Mem/inst_mem_reg[26][26] ,
         \Inst_Mem/inst_mem_reg[26][27] , \Inst_Mem/inst_mem_reg[26][28] ,
         \Inst_Mem/inst_mem_reg[26][29] , \Inst_Mem/inst_mem_reg[26][30] ,
         \Inst_Mem/inst_mem_reg[26][31] , \Inst_Mem/inst_mem_reg[25][0] ,
         \Inst_Mem/inst_mem_reg[25][1] , \Inst_Mem/inst_mem_reg[25][2] ,
         \Inst_Mem/inst_mem_reg[25][3] , \Inst_Mem/inst_mem_reg[25][4] ,
         \Inst_Mem/inst_mem_reg[25][5] , \Inst_Mem/inst_mem_reg[25][6] ,
         \Inst_Mem/inst_mem_reg[25][7] , \Inst_Mem/inst_mem_reg[25][8] ,
         \Inst_Mem/inst_mem_reg[25][9] , \Inst_Mem/inst_mem_reg[25][10] ,
         \Inst_Mem/inst_mem_reg[25][11] , \Inst_Mem/inst_mem_reg[25][12] ,
         \Inst_Mem/inst_mem_reg[25][13] , \Inst_Mem/inst_mem_reg[25][14] ,
         \Inst_Mem/inst_mem_reg[25][15] , \Inst_Mem/inst_mem_reg[25][16] ,
         \Inst_Mem/inst_mem_reg[25][17] , \Inst_Mem/inst_mem_reg[25][18] ,
         \Inst_Mem/inst_mem_reg[25][19] , \Inst_Mem/inst_mem_reg[25][20] ,
         \Inst_Mem/inst_mem_reg[25][21] , \Inst_Mem/inst_mem_reg[25][22] ,
         \Inst_Mem/inst_mem_reg[25][23] , \Inst_Mem/inst_mem_reg[25][24] ,
         \Inst_Mem/inst_mem_reg[25][25] , \Inst_Mem/inst_mem_reg[25][26] ,
         \Inst_Mem/inst_mem_reg[25][27] , \Inst_Mem/inst_mem_reg[25][28] ,
         \Inst_Mem/inst_mem_reg[25][29] , \Inst_Mem/inst_mem_reg[25][30] ,
         \Inst_Mem/inst_mem_reg[25][31] , \Inst_Mem/inst_mem_reg[24][0] ,
         \Inst_Mem/inst_mem_reg[24][1] , \Inst_Mem/inst_mem_reg[24][2] ,
         \Inst_Mem/inst_mem_reg[24][3] , \Inst_Mem/inst_mem_reg[24][4] ,
         \Inst_Mem/inst_mem_reg[24][5] , \Inst_Mem/inst_mem_reg[24][6] ,
         \Inst_Mem/inst_mem_reg[24][7] , \Inst_Mem/inst_mem_reg[24][8] ,
         \Inst_Mem/inst_mem_reg[24][9] , \Inst_Mem/inst_mem_reg[24][10] ,
         \Inst_Mem/inst_mem_reg[24][11] , \Inst_Mem/inst_mem_reg[24][12] ,
         \Inst_Mem/inst_mem_reg[24][13] , \Inst_Mem/inst_mem_reg[24][14] ,
         \Inst_Mem/inst_mem_reg[24][15] , \Inst_Mem/inst_mem_reg[24][16] ,
         \Inst_Mem/inst_mem_reg[24][17] , \Inst_Mem/inst_mem_reg[24][18] ,
         \Inst_Mem/inst_mem_reg[24][19] , \Inst_Mem/inst_mem_reg[24][20] ,
         \Inst_Mem/inst_mem_reg[24][21] , \Inst_Mem/inst_mem_reg[24][22] ,
         \Inst_Mem/inst_mem_reg[24][23] , \Inst_Mem/inst_mem_reg[24][24] ,
         \Inst_Mem/inst_mem_reg[24][25] , \Inst_Mem/inst_mem_reg[24][26] ,
         \Inst_Mem/inst_mem_reg[24][27] , \Inst_Mem/inst_mem_reg[24][28] ,
         \Inst_Mem/inst_mem_reg[24][29] , \Inst_Mem/inst_mem_reg[24][30] ,
         \Inst_Mem/inst_mem_reg[24][31] , \Inst_Mem/inst_mem_reg[23][0] ,
         \Inst_Mem/inst_mem_reg[23][1] , \Inst_Mem/inst_mem_reg[23][2] ,
         \Inst_Mem/inst_mem_reg[23][3] , \Inst_Mem/inst_mem_reg[23][4] ,
         \Inst_Mem/inst_mem_reg[23][5] , \Inst_Mem/inst_mem_reg[23][6] ,
         \Inst_Mem/inst_mem_reg[23][7] , \Inst_Mem/inst_mem_reg[23][8] ,
         \Inst_Mem/inst_mem_reg[23][9] , \Inst_Mem/inst_mem_reg[23][10] ,
         \Inst_Mem/inst_mem_reg[23][11] , \Inst_Mem/inst_mem_reg[23][12] ,
         \Inst_Mem/inst_mem_reg[23][13] , \Inst_Mem/inst_mem_reg[23][14] ,
         \Inst_Mem/inst_mem_reg[23][15] , \Inst_Mem/inst_mem_reg[23][16] ,
         \Inst_Mem/inst_mem_reg[23][17] , \Inst_Mem/inst_mem_reg[23][18] ,
         \Inst_Mem/inst_mem_reg[23][19] , \Inst_Mem/inst_mem_reg[23][20] ,
         \Inst_Mem/inst_mem_reg[23][21] , \Inst_Mem/inst_mem_reg[23][22] ,
         \Inst_Mem/inst_mem_reg[23][23] , \Inst_Mem/inst_mem_reg[23][24] ,
         \Inst_Mem/inst_mem_reg[23][25] , \Inst_Mem/inst_mem_reg[23][26] ,
         \Inst_Mem/inst_mem_reg[23][27] , \Inst_Mem/inst_mem_reg[23][28] ,
         \Inst_Mem/inst_mem_reg[23][29] , \Inst_Mem/inst_mem_reg[23][30] ,
         \Inst_Mem/inst_mem_reg[23][31] , \Inst_Mem/inst_mem_reg[22][0] ,
         \Inst_Mem/inst_mem_reg[22][1] , \Inst_Mem/inst_mem_reg[22][2] ,
         \Inst_Mem/inst_mem_reg[22][3] , \Inst_Mem/inst_mem_reg[22][4] ,
         \Inst_Mem/inst_mem_reg[22][5] , \Inst_Mem/inst_mem_reg[22][6] ,
         \Inst_Mem/inst_mem_reg[22][7] , \Inst_Mem/inst_mem_reg[22][8] ,
         \Inst_Mem/inst_mem_reg[22][9] , \Inst_Mem/inst_mem_reg[22][10] ,
         \Inst_Mem/inst_mem_reg[22][11] , \Inst_Mem/inst_mem_reg[22][12] ,
         \Inst_Mem/inst_mem_reg[22][13] , \Inst_Mem/inst_mem_reg[22][14] ,
         \Inst_Mem/inst_mem_reg[22][15] , \Inst_Mem/inst_mem_reg[22][16] ,
         \Inst_Mem/inst_mem_reg[22][17] , \Inst_Mem/inst_mem_reg[22][18] ,
         \Inst_Mem/inst_mem_reg[22][19] , \Inst_Mem/inst_mem_reg[22][20] ,
         \Inst_Mem/inst_mem_reg[22][21] , \Inst_Mem/inst_mem_reg[22][22] ,
         \Inst_Mem/inst_mem_reg[22][23] , \Inst_Mem/inst_mem_reg[22][24] ,
         \Inst_Mem/inst_mem_reg[22][25] , \Inst_Mem/inst_mem_reg[22][26] ,
         \Inst_Mem/inst_mem_reg[22][27] , \Inst_Mem/inst_mem_reg[22][28] ,
         \Inst_Mem/inst_mem_reg[22][29] , \Inst_Mem/inst_mem_reg[22][30] ,
         \Inst_Mem/inst_mem_reg[22][31] , \Inst_Mem/inst_mem_reg[21][0] ,
         \Inst_Mem/inst_mem_reg[21][1] , \Inst_Mem/inst_mem_reg[21][2] ,
         \Inst_Mem/inst_mem_reg[21][3] , \Inst_Mem/inst_mem_reg[21][4] ,
         \Inst_Mem/inst_mem_reg[21][5] , \Inst_Mem/inst_mem_reg[21][6] ,
         \Inst_Mem/inst_mem_reg[21][7] , \Inst_Mem/inst_mem_reg[21][8] ,
         \Inst_Mem/inst_mem_reg[21][9] , \Inst_Mem/inst_mem_reg[21][10] ,
         \Inst_Mem/inst_mem_reg[21][11] , \Inst_Mem/inst_mem_reg[21][12] ,
         \Inst_Mem/inst_mem_reg[21][13] , \Inst_Mem/inst_mem_reg[21][14] ,
         \Inst_Mem/inst_mem_reg[21][15] , \Inst_Mem/inst_mem_reg[21][16] ,
         \Inst_Mem/inst_mem_reg[21][17] , \Inst_Mem/inst_mem_reg[21][18] ,
         \Inst_Mem/inst_mem_reg[21][19] , \Inst_Mem/inst_mem_reg[21][20] ,
         \Inst_Mem/inst_mem_reg[21][21] , \Inst_Mem/inst_mem_reg[21][22] ,
         \Inst_Mem/inst_mem_reg[21][23] , \Inst_Mem/inst_mem_reg[21][24] ,
         \Inst_Mem/inst_mem_reg[21][25] , \Inst_Mem/inst_mem_reg[21][26] ,
         \Inst_Mem/inst_mem_reg[21][27] , \Inst_Mem/inst_mem_reg[21][28] ,
         \Inst_Mem/inst_mem_reg[21][29] , \Inst_Mem/inst_mem_reg[21][30] ,
         \Inst_Mem/inst_mem_reg[21][31] , \Inst_Mem/inst_mem_reg[20][0] ,
         \Inst_Mem/inst_mem_reg[20][1] , \Inst_Mem/inst_mem_reg[20][2] ,
         \Inst_Mem/inst_mem_reg[20][3] , \Inst_Mem/inst_mem_reg[20][4] ,
         \Inst_Mem/inst_mem_reg[20][5] , \Inst_Mem/inst_mem_reg[20][6] ,
         \Inst_Mem/inst_mem_reg[20][7] , \Inst_Mem/inst_mem_reg[20][8] ,
         \Inst_Mem/inst_mem_reg[20][9] , \Inst_Mem/inst_mem_reg[20][10] ,
         \Inst_Mem/inst_mem_reg[20][11] , \Inst_Mem/inst_mem_reg[20][12] ,
         \Inst_Mem/inst_mem_reg[20][13] , \Inst_Mem/inst_mem_reg[20][14] ,
         \Inst_Mem/inst_mem_reg[20][15] , \Inst_Mem/inst_mem_reg[20][16] ,
         \Inst_Mem/inst_mem_reg[20][17] , \Inst_Mem/inst_mem_reg[20][18] ,
         \Inst_Mem/inst_mem_reg[20][19] , \Inst_Mem/inst_mem_reg[20][20] ,
         \Inst_Mem/inst_mem_reg[20][21] , \Inst_Mem/inst_mem_reg[20][22] ,
         \Inst_Mem/inst_mem_reg[20][23] , \Inst_Mem/inst_mem_reg[20][24] ,
         \Inst_Mem/inst_mem_reg[20][25] , \Inst_Mem/inst_mem_reg[20][26] ,
         \Inst_Mem/inst_mem_reg[20][27] , \Inst_Mem/inst_mem_reg[20][28] ,
         \Inst_Mem/inst_mem_reg[20][29] , \Inst_Mem/inst_mem_reg[20][30] ,
         \Inst_Mem/inst_mem_reg[20][31] , \Inst_Mem/inst_mem_reg[19][0] ,
         \Inst_Mem/inst_mem_reg[19][1] , \Inst_Mem/inst_mem_reg[19][2] ,
         \Inst_Mem/inst_mem_reg[19][3] , \Inst_Mem/inst_mem_reg[19][4] ,
         \Inst_Mem/inst_mem_reg[19][5] , \Inst_Mem/inst_mem_reg[19][6] ,
         \Inst_Mem/inst_mem_reg[19][7] , \Inst_Mem/inst_mem_reg[19][8] ,
         \Inst_Mem/inst_mem_reg[19][9] , \Inst_Mem/inst_mem_reg[19][10] ,
         \Inst_Mem/inst_mem_reg[19][11] , \Inst_Mem/inst_mem_reg[19][12] ,
         \Inst_Mem/inst_mem_reg[19][13] , \Inst_Mem/inst_mem_reg[19][14] ,
         \Inst_Mem/inst_mem_reg[19][15] , \Inst_Mem/inst_mem_reg[19][16] ,
         \Inst_Mem/inst_mem_reg[19][17] , \Inst_Mem/inst_mem_reg[19][18] ,
         \Inst_Mem/inst_mem_reg[19][19] , \Inst_Mem/inst_mem_reg[19][20] ,
         \Inst_Mem/inst_mem_reg[19][21] , \Inst_Mem/inst_mem_reg[19][22] ,
         \Inst_Mem/inst_mem_reg[19][23] , \Inst_Mem/inst_mem_reg[19][24] ,
         \Inst_Mem/inst_mem_reg[19][25] , \Inst_Mem/inst_mem_reg[19][26] ,
         \Inst_Mem/inst_mem_reg[19][27] , \Inst_Mem/inst_mem_reg[19][28] ,
         \Inst_Mem/inst_mem_reg[19][29] , \Inst_Mem/inst_mem_reg[19][30] ,
         \Inst_Mem/inst_mem_reg[19][31] , \Inst_Mem/inst_mem_reg[18][0] ,
         \Inst_Mem/inst_mem_reg[18][1] , \Inst_Mem/inst_mem_reg[18][2] ,
         \Inst_Mem/inst_mem_reg[18][3] , \Inst_Mem/inst_mem_reg[18][4] ,
         \Inst_Mem/inst_mem_reg[18][5] , \Inst_Mem/inst_mem_reg[18][6] ,
         \Inst_Mem/inst_mem_reg[18][7] , \Inst_Mem/inst_mem_reg[18][8] ,
         \Inst_Mem/inst_mem_reg[18][9] , \Inst_Mem/inst_mem_reg[18][10] ,
         \Inst_Mem/inst_mem_reg[18][11] , \Inst_Mem/inst_mem_reg[18][12] ,
         \Inst_Mem/inst_mem_reg[18][13] , \Inst_Mem/inst_mem_reg[18][14] ,
         \Inst_Mem/inst_mem_reg[18][15] , \Inst_Mem/inst_mem_reg[18][16] ,
         \Inst_Mem/inst_mem_reg[18][17] , \Inst_Mem/inst_mem_reg[18][18] ,
         \Inst_Mem/inst_mem_reg[18][19] , \Inst_Mem/inst_mem_reg[18][20] ,
         \Inst_Mem/inst_mem_reg[18][21] , \Inst_Mem/inst_mem_reg[18][22] ,
         \Inst_Mem/inst_mem_reg[18][23] , \Inst_Mem/inst_mem_reg[18][24] ,
         \Inst_Mem/inst_mem_reg[18][25] , \Inst_Mem/inst_mem_reg[18][26] ,
         \Inst_Mem/inst_mem_reg[18][27] , \Inst_Mem/inst_mem_reg[18][28] ,
         \Inst_Mem/inst_mem_reg[18][29] , \Inst_Mem/inst_mem_reg[18][30] ,
         \Inst_Mem/inst_mem_reg[18][31] , \Inst_Mem/inst_mem_reg[17][0] ,
         \Inst_Mem/inst_mem_reg[17][1] , \Inst_Mem/inst_mem_reg[17][2] ,
         \Inst_Mem/inst_mem_reg[17][3] , \Inst_Mem/inst_mem_reg[17][4] ,
         \Inst_Mem/inst_mem_reg[17][5] , \Inst_Mem/inst_mem_reg[17][6] ,
         \Inst_Mem/inst_mem_reg[17][7] , \Inst_Mem/inst_mem_reg[17][8] ,
         \Inst_Mem/inst_mem_reg[17][9] , \Inst_Mem/inst_mem_reg[17][10] ,
         \Inst_Mem/inst_mem_reg[17][11] , \Inst_Mem/inst_mem_reg[17][12] ,
         \Inst_Mem/inst_mem_reg[17][13] , \Inst_Mem/inst_mem_reg[17][14] ,
         \Inst_Mem/inst_mem_reg[17][15] , \Inst_Mem/inst_mem_reg[17][16] ,
         \Inst_Mem/inst_mem_reg[17][17] , \Inst_Mem/inst_mem_reg[17][18] ,
         \Inst_Mem/inst_mem_reg[17][19] , \Inst_Mem/inst_mem_reg[17][20] ,
         \Inst_Mem/inst_mem_reg[17][21] , \Inst_Mem/inst_mem_reg[17][22] ,
         \Inst_Mem/inst_mem_reg[17][23] , \Inst_Mem/inst_mem_reg[17][24] ,
         \Inst_Mem/inst_mem_reg[17][25] , \Inst_Mem/inst_mem_reg[17][26] ,
         \Inst_Mem/inst_mem_reg[17][27] , \Inst_Mem/inst_mem_reg[17][28] ,
         \Inst_Mem/inst_mem_reg[17][29] , \Inst_Mem/inst_mem_reg[17][30] ,
         \Inst_Mem/inst_mem_reg[17][31] , \Inst_Mem/inst_mem_reg[16][0] ,
         \Inst_Mem/inst_mem_reg[16][1] , \Inst_Mem/inst_mem_reg[16][2] ,
         \Inst_Mem/inst_mem_reg[16][3] , \Inst_Mem/inst_mem_reg[16][4] ,
         \Inst_Mem/inst_mem_reg[16][5] , \Inst_Mem/inst_mem_reg[16][6] ,
         \Inst_Mem/inst_mem_reg[16][7] , \Inst_Mem/inst_mem_reg[16][8] ,
         \Inst_Mem/inst_mem_reg[16][9] , \Inst_Mem/inst_mem_reg[16][10] ,
         \Inst_Mem/inst_mem_reg[16][11] , \Inst_Mem/inst_mem_reg[16][12] ,
         \Inst_Mem/inst_mem_reg[16][13] , \Inst_Mem/inst_mem_reg[16][14] ,
         \Inst_Mem/inst_mem_reg[16][15] , \Inst_Mem/inst_mem_reg[16][16] ,
         \Inst_Mem/inst_mem_reg[16][17] , \Inst_Mem/inst_mem_reg[16][18] ,
         \Inst_Mem/inst_mem_reg[16][19] , \Inst_Mem/inst_mem_reg[16][20] ,
         \Inst_Mem/inst_mem_reg[16][21] , \Inst_Mem/inst_mem_reg[16][22] ,
         \Inst_Mem/inst_mem_reg[16][23] , \Inst_Mem/inst_mem_reg[16][24] ,
         \Inst_Mem/inst_mem_reg[16][25] , \Inst_Mem/inst_mem_reg[16][26] ,
         \Inst_Mem/inst_mem_reg[16][27] , \Inst_Mem/inst_mem_reg[16][28] ,
         \Inst_Mem/inst_mem_reg[16][29] , \Inst_Mem/inst_mem_reg[16][30] ,
         \Inst_Mem/inst_mem_reg[16][31] , \Inst_Mem/inst_mem_reg[15][0] ,
         \Inst_Mem/inst_mem_reg[15][1] , \Inst_Mem/inst_mem_reg[15][2] ,
         \Inst_Mem/inst_mem_reg[15][3] , \Inst_Mem/inst_mem_reg[15][4] ,
         \Inst_Mem/inst_mem_reg[15][5] , \Inst_Mem/inst_mem_reg[15][6] ,
         \Inst_Mem/inst_mem_reg[15][7] , \Inst_Mem/inst_mem_reg[15][8] ,
         \Inst_Mem/inst_mem_reg[15][9] , \Inst_Mem/inst_mem_reg[15][10] ,
         \Inst_Mem/inst_mem_reg[15][11] , \Inst_Mem/inst_mem_reg[15][12] ,
         \Inst_Mem/inst_mem_reg[15][13] , \Inst_Mem/inst_mem_reg[15][14] ,
         \Inst_Mem/inst_mem_reg[15][15] , \Inst_Mem/inst_mem_reg[15][16] ,
         \Inst_Mem/inst_mem_reg[15][17] , \Inst_Mem/inst_mem_reg[15][18] ,
         \Inst_Mem/inst_mem_reg[15][19] , \Inst_Mem/inst_mem_reg[15][20] ,
         \Inst_Mem/inst_mem_reg[15][21] , \Inst_Mem/inst_mem_reg[15][22] ,
         \Inst_Mem/inst_mem_reg[15][23] , \Inst_Mem/inst_mem_reg[15][24] ,
         \Inst_Mem/inst_mem_reg[15][25] , \Inst_Mem/inst_mem_reg[15][26] ,
         \Inst_Mem/inst_mem_reg[15][27] , \Inst_Mem/inst_mem_reg[15][28] ,
         \Inst_Mem/inst_mem_reg[15][29] , \Inst_Mem/inst_mem_reg[15][30] ,
         \Inst_Mem/inst_mem_reg[15][31] , \Inst_Mem/inst_mem_reg[14][0] ,
         \Inst_Mem/inst_mem_reg[14][1] , \Inst_Mem/inst_mem_reg[14][2] ,
         \Inst_Mem/inst_mem_reg[14][3] , \Inst_Mem/inst_mem_reg[14][4] ,
         \Inst_Mem/inst_mem_reg[14][5] , \Inst_Mem/inst_mem_reg[14][6] ,
         \Inst_Mem/inst_mem_reg[14][7] , \Inst_Mem/inst_mem_reg[14][8] ,
         \Inst_Mem/inst_mem_reg[14][9] , \Inst_Mem/inst_mem_reg[14][10] ,
         \Inst_Mem/inst_mem_reg[14][11] , \Inst_Mem/inst_mem_reg[14][12] ,
         \Inst_Mem/inst_mem_reg[14][13] , \Inst_Mem/inst_mem_reg[14][14] ,
         \Inst_Mem/inst_mem_reg[14][15] , \Inst_Mem/inst_mem_reg[14][16] ,
         \Inst_Mem/inst_mem_reg[14][17] , \Inst_Mem/inst_mem_reg[14][18] ,
         \Inst_Mem/inst_mem_reg[14][19] , \Inst_Mem/inst_mem_reg[14][20] ,
         \Inst_Mem/inst_mem_reg[14][21] , \Inst_Mem/inst_mem_reg[14][22] ,
         \Inst_Mem/inst_mem_reg[14][23] , \Inst_Mem/inst_mem_reg[14][24] ,
         \Inst_Mem/inst_mem_reg[14][25] , \Inst_Mem/inst_mem_reg[14][26] ,
         \Inst_Mem/inst_mem_reg[14][27] , \Inst_Mem/inst_mem_reg[14][28] ,
         \Inst_Mem/inst_mem_reg[14][29] , \Inst_Mem/inst_mem_reg[14][30] ,
         \Inst_Mem/inst_mem_reg[14][31] , \Inst_Mem/inst_mem_reg[13][0] ,
         \Inst_Mem/inst_mem_reg[13][1] , \Inst_Mem/inst_mem_reg[13][2] ,
         \Inst_Mem/inst_mem_reg[13][3] , \Inst_Mem/inst_mem_reg[13][4] ,
         \Inst_Mem/inst_mem_reg[13][5] , \Inst_Mem/inst_mem_reg[13][6] ,
         \Inst_Mem/inst_mem_reg[13][7] , \Inst_Mem/inst_mem_reg[13][8] ,
         \Inst_Mem/inst_mem_reg[13][9] , \Inst_Mem/inst_mem_reg[13][10] ,
         \Inst_Mem/inst_mem_reg[13][11] , \Inst_Mem/inst_mem_reg[13][12] ,
         \Inst_Mem/inst_mem_reg[13][13] , \Inst_Mem/inst_mem_reg[13][14] ,
         \Inst_Mem/inst_mem_reg[13][15] , \Inst_Mem/inst_mem_reg[13][16] ,
         \Inst_Mem/inst_mem_reg[13][17] , \Inst_Mem/inst_mem_reg[13][18] ,
         \Inst_Mem/inst_mem_reg[13][19] , \Inst_Mem/inst_mem_reg[13][20] ,
         \Inst_Mem/inst_mem_reg[13][21] , \Inst_Mem/inst_mem_reg[13][22] ,
         \Inst_Mem/inst_mem_reg[13][23] , \Inst_Mem/inst_mem_reg[13][24] ,
         \Inst_Mem/inst_mem_reg[13][25] , \Inst_Mem/inst_mem_reg[13][26] ,
         \Inst_Mem/inst_mem_reg[13][27] , \Inst_Mem/inst_mem_reg[13][28] ,
         \Inst_Mem/inst_mem_reg[13][29] , \Inst_Mem/inst_mem_reg[13][30] ,
         \Inst_Mem/inst_mem_reg[13][31] , \Inst_Mem/inst_mem_reg[12][0] ,
         \Inst_Mem/inst_mem_reg[12][1] , \Inst_Mem/inst_mem_reg[12][2] ,
         \Inst_Mem/inst_mem_reg[12][3] , \Inst_Mem/inst_mem_reg[12][4] ,
         \Inst_Mem/inst_mem_reg[12][5] , \Inst_Mem/inst_mem_reg[12][6] ,
         \Inst_Mem/inst_mem_reg[12][7] , \Inst_Mem/inst_mem_reg[12][8] ,
         \Inst_Mem/inst_mem_reg[12][9] , \Inst_Mem/inst_mem_reg[12][10] ,
         \Inst_Mem/inst_mem_reg[12][11] , \Inst_Mem/inst_mem_reg[12][12] ,
         \Inst_Mem/inst_mem_reg[12][13] , \Inst_Mem/inst_mem_reg[12][14] ,
         \Inst_Mem/inst_mem_reg[12][15] , \Inst_Mem/inst_mem_reg[12][16] ,
         \Inst_Mem/inst_mem_reg[12][17] , \Inst_Mem/inst_mem_reg[12][18] ,
         \Inst_Mem/inst_mem_reg[12][19] , \Inst_Mem/inst_mem_reg[12][20] ,
         \Inst_Mem/inst_mem_reg[12][21] , \Inst_Mem/inst_mem_reg[12][22] ,
         \Inst_Mem/inst_mem_reg[12][23] , \Inst_Mem/inst_mem_reg[12][24] ,
         \Inst_Mem/inst_mem_reg[12][25] , \Inst_Mem/inst_mem_reg[12][26] ,
         \Inst_Mem/inst_mem_reg[12][27] , \Inst_Mem/inst_mem_reg[12][28] ,
         \Inst_Mem/inst_mem_reg[12][29] , \Inst_Mem/inst_mem_reg[12][30] ,
         \Inst_Mem/inst_mem_reg[12][31] , \Inst_Mem/inst_mem_reg[11][0] ,
         \Inst_Mem/inst_mem_reg[11][1] , \Inst_Mem/inst_mem_reg[11][2] ,
         \Inst_Mem/inst_mem_reg[11][3] , \Inst_Mem/inst_mem_reg[11][4] ,
         \Inst_Mem/inst_mem_reg[11][5] , \Inst_Mem/inst_mem_reg[11][6] ,
         \Inst_Mem/inst_mem_reg[11][7] , \Inst_Mem/inst_mem_reg[11][8] ,
         \Inst_Mem/inst_mem_reg[11][9] , \Inst_Mem/inst_mem_reg[11][10] ,
         \Inst_Mem/inst_mem_reg[11][11] , \Inst_Mem/inst_mem_reg[11][12] ,
         \Inst_Mem/inst_mem_reg[11][13] , \Inst_Mem/inst_mem_reg[11][14] ,
         \Inst_Mem/inst_mem_reg[11][15] , \Inst_Mem/inst_mem_reg[11][16] ,
         \Inst_Mem/inst_mem_reg[11][17] , \Inst_Mem/inst_mem_reg[11][18] ,
         \Inst_Mem/inst_mem_reg[11][19] , \Inst_Mem/inst_mem_reg[11][20] ,
         \Inst_Mem/inst_mem_reg[11][21] , \Inst_Mem/inst_mem_reg[11][22] ,
         \Inst_Mem/inst_mem_reg[11][23] , \Inst_Mem/inst_mem_reg[11][24] ,
         \Inst_Mem/inst_mem_reg[11][25] , \Inst_Mem/inst_mem_reg[11][26] ,
         \Inst_Mem/inst_mem_reg[11][27] , \Inst_Mem/inst_mem_reg[11][28] ,
         \Inst_Mem/inst_mem_reg[11][29] , \Inst_Mem/inst_mem_reg[11][30] ,
         \Inst_Mem/inst_mem_reg[11][31] , \Inst_Mem/inst_mem_reg[10][0] ,
         \Inst_Mem/inst_mem_reg[10][1] , \Inst_Mem/inst_mem_reg[10][2] ,
         \Inst_Mem/inst_mem_reg[10][3] , \Inst_Mem/inst_mem_reg[10][4] ,
         \Inst_Mem/inst_mem_reg[10][5] , \Inst_Mem/inst_mem_reg[10][6] ,
         \Inst_Mem/inst_mem_reg[10][7] , \Inst_Mem/inst_mem_reg[10][8] ,
         \Inst_Mem/inst_mem_reg[10][9] , \Inst_Mem/inst_mem_reg[10][10] ,
         \Inst_Mem/inst_mem_reg[10][11] , \Inst_Mem/inst_mem_reg[10][12] ,
         \Inst_Mem/inst_mem_reg[10][13] , \Inst_Mem/inst_mem_reg[10][14] ,
         \Inst_Mem/inst_mem_reg[10][15] , \Inst_Mem/inst_mem_reg[10][16] ,
         \Inst_Mem/inst_mem_reg[10][17] , \Inst_Mem/inst_mem_reg[10][18] ,
         \Inst_Mem/inst_mem_reg[10][19] , \Inst_Mem/inst_mem_reg[10][20] ,
         \Inst_Mem/inst_mem_reg[10][21] , \Inst_Mem/inst_mem_reg[10][22] ,
         \Inst_Mem/inst_mem_reg[10][23] , \Inst_Mem/inst_mem_reg[10][24] ,
         \Inst_Mem/inst_mem_reg[10][25] , \Inst_Mem/inst_mem_reg[10][26] ,
         \Inst_Mem/inst_mem_reg[10][27] , \Inst_Mem/inst_mem_reg[10][28] ,
         \Inst_Mem/inst_mem_reg[10][29] , \Inst_Mem/inst_mem_reg[10][30] ,
         \Inst_Mem/inst_mem_reg[10][31] , \Inst_Mem/inst_mem_reg[9][0] ,
         \Inst_Mem/inst_mem_reg[9][1] , \Inst_Mem/inst_mem_reg[9][2] ,
         \Inst_Mem/inst_mem_reg[9][3] , \Inst_Mem/inst_mem_reg[9][4] ,
         \Inst_Mem/inst_mem_reg[9][5] , \Inst_Mem/inst_mem_reg[9][6] ,
         \Inst_Mem/inst_mem_reg[9][7] , \Inst_Mem/inst_mem_reg[9][8] ,
         \Inst_Mem/inst_mem_reg[9][9] , \Inst_Mem/inst_mem_reg[9][10] ,
         \Inst_Mem/inst_mem_reg[9][11] , \Inst_Mem/inst_mem_reg[9][12] ,
         \Inst_Mem/inst_mem_reg[9][13] , \Inst_Mem/inst_mem_reg[9][14] ,
         \Inst_Mem/inst_mem_reg[9][15] , \Inst_Mem/inst_mem_reg[9][16] ,
         \Inst_Mem/inst_mem_reg[9][17] , \Inst_Mem/inst_mem_reg[9][18] ,
         \Inst_Mem/inst_mem_reg[9][19] , \Inst_Mem/inst_mem_reg[9][20] ,
         \Inst_Mem/inst_mem_reg[9][21] , \Inst_Mem/inst_mem_reg[9][22] ,
         \Inst_Mem/inst_mem_reg[9][23] , \Inst_Mem/inst_mem_reg[9][24] ,
         \Inst_Mem/inst_mem_reg[9][25] , \Inst_Mem/inst_mem_reg[9][26] ,
         \Inst_Mem/inst_mem_reg[9][27] , \Inst_Mem/inst_mem_reg[9][28] ,
         \Inst_Mem/inst_mem_reg[9][29] , \Inst_Mem/inst_mem_reg[9][30] ,
         \Inst_Mem/inst_mem_reg[9][31] , \Inst_Mem/inst_mem_reg[8][0] ,
         \Inst_Mem/inst_mem_reg[8][1] , \Inst_Mem/inst_mem_reg[8][2] ,
         \Inst_Mem/inst_mem_reg[8][3] , \Inst_Mem/inst_mem_reg[8][4] ,
         \Inst_Mem/inst_mem_reg[8][5] , \Inst_Mem/inst_mem_reg[8][6] ,
         \Inst_Mem/inst_mem_reg[8][7] , \Inst_Mem/inst_mem_reg[8][8] ,
         \Inst_Mem/inst_mem_reg[8][9] , \Inst_Mem/inst_mem_reg[8][10] ,
         \Inst_Mem/inst_mem_reg[8][11] , \Inst_Mem/inst_mem_reg[8][12] ,
         \Inst_Mem/inst_mem_reg[8][13] , \Inst_Mem/inst_mem_reg[8][14] ,
         \Inst_Mem/inst_mem_reg[8][15] , \Inst_Mem/inst_mem_reg[8][16] ,
         \Inst_Mem/inst_mem_reg[8][17] , \Inst_Mem/inst_mem_reg[8][18] ,
         \Inst_Mem/inst_mem_reg[8][19] , \Inst_Mem/inst_mem_reg[8][20] ,
         \Inst_Mem/inst_mem_reg[8][21] , \Inst_Mem/inst_mem_reg[8][22] ,
         \Inst_Mem/inst_mem_reg[8][23] , \Inst_Mem/inst_mem_reg[8][24] ,
         \Inst_Mem/inst_mem_reg[8][25] , \Inst_Mem/inst_mem_reg[8][26] ,
         \Inst_Mem/inst_mem_reg[8][27] , \Inst_Mem/inst_mem_reg[8][28] ,
         \Inst_Mem/inst_mem_reg[8][29] , \Inst_Mem/inst_mem_reg[8][30] ,
         \Inst_Mem/inst_mem_reg[8][31] , \Inst_Mem/inst_mem_reg[7][0] ,
         \Inst_Mem/inst_mem_reg[7][1] , \Inst_Mem/inst_mem_reg[7][2] ,
         \Inst_Mem/inst_mem_reg[7][3] , \Inst_Mem/inst_mem_reg[7][4] ,
         \Inst_Mem/inst_mem_reg[7][5] , \Inst_Mem/inst_mem_reg[7][6] ,
         \Inst_Mem/inst_mem_reg[7][7] , \Inst_Mem/inst_mem_reg[7][8] ,
         \Inst_Mem/inst_mem_reg[7][9] , \Inst_Mem/inst_mem_reg[7][10] ,
         \Inst_Mem/inst_mem_reg[7][11] , \Inst_Mem/inst_mem_reg[7][12] ,
         \Inst_Mem/inst_mem_reg[7][13] , \Inst_Mem/inst_mem_reg[7][14] ,
         \Inst_Mem/inst_mem_reg[7][15] , \Inst_Mem/inst_mem_reg[7][16] ,
         \Inst_Mem/inst_mem_reg[7][17] , \Inst_Mem/inst_mem_reg[7][18] ,
         \Inst_Mem/inst_mem_reg[7][19] , \Inst_Mem/inst_mem_reg[7][20] ,
         \Inst_Mem/inst_mem_reg[7][21] , \Inst_Mem/inst_mem_reg[7][22] ,
         \Inst_Mem/inst_mem_reg[7][23] , \Inst_Mem/inst_mem_reg[7][24] ,
         \Inst_Mem/inst_mem_reg[7][25] , \Inst_Mem/inst_mem_reg[7][26] ,
         \Inst_Mem/inst_mem_reg[7][27] , \Inst_Mem/inst_mem_reg[7][28] ,
         \Inst_Mem/inst_mem_reg[7][29] , \Inst_Mem/inst_mem_reg[7][30] ,
         \Inst_Mem/inst_mem_reg[7][31] , \Inst_Mem/inst_mem_reg[6][0] ,
         \Inst_Mem/inst_mem_reg[6][1] , \Inst_Mem/inst_mem_reg[6][2] ,
         \Inst_Mem/inst_mem_reg[6][3] , \Inst_Mem/inst_mem_reg[6][4] ,
         \Inst_Mem/inst_mem_reg[6][5] , \Inst_Mem/inst_mem_reg[6][6] ,
         \Inst_Mem/inst_mem_reg[6][7] , \Inst_Mem/inst_mem_reg[6][8] ,
         \Inst_Mem/inst_mem_reg[6][9] , \Inst_Mem/inst_mem_reg[6][10] ,
         \Inst_Mem/inst_mem_reg[6][11] , \Inst_Mem/inst_mem_reg[6][12] ,
         \Inst_Mem/inst_mem_reg[6][13] , \Inst_Mem/inst_mem_reg[6][14] ,
         \Inst_Mem/inst_mem_reg[6][15] , \Inst_Mem/inst_mem_reg[6][16] ,
         \Inst_Mem/inst_mem_reg[6][17] , \Inst_Mem/inst_mem_reg[6][18] ,
         \Inst_Mem/inst_mem_reg[6][19] , \Inst_Mem/inst_mem_reg[6][20] ,
         \Inst_Mem/inst_mem_reg[6][21] , \Inst_Mem/inst_mem_reg[6][22] ,
         \Inst_Mem/inst_mem_reg[6][23] , \Inst_Mem/inst_mem_reg[6][24] ,
         \Inst_Mem/inst_mem_reg[6][25] , \Inst_Mem/inst_mem_reg[6][26] ,
         \Inst_Mem/inst_mem_reg[6][27] , \Inst_Mem/inst_mem_reg[6][28] ,
         \Inst_Mem/inst_mem_reg[6][29] , \Inst_Mem/inst_mem_reg[6][30] ,
         \Inst_Mem/inst_mem_reg[6][31] , \Inst_Mem/inst_mem_reg[5][0] ,
         \Inst_Mem/inst_mem_reg[5][1] , \Inst_Mem/inst_mem_reg[5][2] ,
         \Inst_Mem/inst_mem_reg[5][3] , \Inst_Mem/inst_mem_reg[5][4] ,
         \Inst_Mem/inst_mem_reg[5][5] , \Inst_Mem/inst_mem_reg[5][6] ,
         \Inst_Mem/inst_mem_reg[5][7] , \Inst_Mem/inst_mem_reg[5][8] ,
         \Inst_Mem/inst_mem_reg[5][9] , \Inst_Mem/inst_mem_reg[5][10] ,
         \Inst_Mem/inst_mem_reg[5][11] , \Inst_Mem/inst_mem_reg[5][12] ,
         \Inst_Mem/inst_mem_reg[5][13] , \Inst_Mem/inst_mem_reg[5][14] ,
         \Inst_Mem/inst_mem_reg[5][15] , \Inst_Mem/inst_mem_reg[5][16] ,
         \Inst_Mem/inst_mem_reg[5][17] , \Inst_Mem/inst_mem_reg[5][18] ,
         \Inst_Mem/inst_mem_reg[5][19] , \Inst_Mem/inst_mem_reg[5][20] ,
         \Inst_Mem/inst_mem_reg[5][21] , \Inst_Mem/inst_mem_reg[5][22] ,
         \Inst_Mem/inst_mem_reg[5][23] , \Inst_Mem/inst_mem_reg[5][24] ,
         \Inst_Mem/inst_mem_reg[5][25] , \Inst_Mem/inst_mem_reg[5][26] ,
         \Inst_Mem/inst_mem_reg[5][27] , \Inst_Mem/inst_mem_reg[5][28] ,
         \Inst_Mem/inst_mem_reg[5][29] , \Inst_Mem/inst_mem_reg[5][30] ,
         \Inst_Mem/inst_mem_reg[5][31] , \Inst_Mem/inst_mem_reg[4][0] ,
         \Inst_Mem/inst_mem_reg[4][1] , \Inst_Mem/inst_mem_reg[4][2] ,
         \Inst_Mem/inst_mem_reg[4][3] , \Inst_Mem/inst_mem_reg[4][4] ,
         \Inst_Mem/inst_mem_reg[4][5] , \Inst_Mem/inst_mem_reg[4][6] ,
         \Inst_Mem/inst_mem_reg[4][7] , \Inst_Mem/inst_mem_reg[4][8] ,
         \Inst_Mem/inst_mem_reg[4][9] , \Inst_Mem/inst_mem_reg[4][10] ,
         \Inst_Mem/inst_mem_reg[4][11] , \Inst_Mem/inst_mem_reg[4][12] ,
         \Inst_Mem/inst_mem_reg[4][13] , \Inst_Mem/inst_mem_reg[4][14] ,
         \Inst_Mem/inst_mem_reg[4][15] , \Inst_Mem/inst_mem_reg[4][16] ,
         \Inst_Mem/inst_mem_reg[4][17] , \Inst_Mem/inst_mem_reg[4][18] ,
         \Inst_Mem/inst_mem_reg[4][19] , \Inst_Mem/inst_mem_reg[4][20] ,
         \Inst_Mem/inst_mem_reg[4][21] , \Inst_Mem/inst_mem_reg[4][22] ,
         \Inst_Mem/inst_mem_reg[4][23] , \Inst_Mem/inst_mem_reg[4][24] ,
         \Inst_Mem/inst_mem_reg[4][25] , \Inst_Mem/inst_mem_reg[4][26] ,
         \Inst_Mem/inst_mem_reg[4][27] , \Inst_Mem/inst_mem_reg[4][28] ,
         \Inst_Mem/inst_mem_reg[4][29] , \Inst_Mem/inst_mem_reg[4][30] ,
         \Inst_Mem/inst_mem_reg[4][31] , \Inst_Mem/inst_mem_reg[3][0] ,
         \Inst_Mem/inst_mem_reg[3][1] , \Inst_Mem/inst_mem_reg[3][2] ,
         \Inst_Mem/inst_mem_reg[3][3] , \Inst_Mem/inst_mem_reg[3][4] ,
         \Inst_Mem/inst_mem_reg[3][5] , \Inst_Mem/inst_mem_reg[3][6] ,
         \Inst_Mem/inst_mem_reg[3][7] , \Inst_Mem/inst_mem_reg[3][8] ,
         \Inst_Mem/inst_mem_reg[3][9] , \Inst_Mem/inst_mem_reg[3][10] ,
         \Inst_Mem/inst_mem_reg[3][11] , \Inst_Mem/inst_mem_reg[3][12] ,
         \Inst_Mem/inst_mem_reg[3][13] , \Inst_Mem/inst_mem_reg[3][14] ,
         \Inst_Mem/inst_mem_reg[3][15] , \Inst_Mem/inst_mem_reg[3][16] ,
         \Inst_Mem/inst_mem_reg[3][17] , \Inst_Mem/inst_mem_reg[3][18] ,
         \Inst_Mem/inst_mem_reg[3][19] , \Inst_Mem/inst_mem_reg[3][20] ,
         \Inst_Mem/inst_mem_reg[3][21] , \Inst_Mem/inst_mem_reg[3][22] ,
         \Inst_Mem/inst_mem_reg[3][23] , \Inst_Mem/inst_mem_reg[3][24] ,
         \Inst_Mem/inst_mem_reg[3][25] , \Inst_Mem/inst_mem_reg[3][26] ,
         \Inst_Mem/inst_mem_reg[3][27] , \Inst_Mem/inst_mem_reg[3][28] ,
         \Inst_Mem/inst_mem_reg[3][29] , \Inst_Mem/inst_mem_reg[3][30] ,
         \Inst_Mem/inst_mem_reg[3][31] , \Inst_Mem/inst_mem_reg[2][0] ,
         \Inst_Mem/inst_mem_reg[2][1] , \Inst_Mem/inst_mem_reg[2][2] ,
         \Inst_Mem/inst_mem_reg[2][3] , \Inst_Mem/inst_mem_reg[2][4] ,
         \Inst_Mem/inst_mem_reg[2][5] , \Inst_Mem/inst_mem_reg[2][6] ,
         \Inst_Mem/inst_mem_reg[2][7] , \Inst_Mem/inst_mem_reg[2][8] ,
         \Inst_Mem/inst_mem_reg[2][9] , \Inst_Mem/inst_mem_reg[2][10] ,
         \Inst_Mem/inst_mem_reg[2][11] , \Inst_Mem/inst_mem_reg[2][12] ,
         \Inst_Mem/inst_mem_reg[2][13] , \Inst_Mem/inst_mem_reg[2][14] ,
         \Inst_Mem/inst_mem_reg[2][15] , \Inst_Mem/inst_mem_reg[2][16] ,
         \Inst_Mem/inst_mem_reg[2][17] , \Inst_Mem/inst_mem_reg[2][18] ,
         \Inst_Mem/inst_mem_reg[2][19] , \Inst_Mem/inst_mem_reg[2][20] ,
         \Inst_Mem/inst_mem_reg[2][21] , \Inst_Mem/inst_mem_reg[2][22] ,
         \Inst_Mem/inst_mem_reg[2][23] , \Inst_Mem/inst_mem_reg[2][24] ,
         \Inst_Mem/inst_mem_reg[2][25] , \Inst_Mem/inst_mem_reg[2][26] ,
         \Inst_Mem/inst_mem_reg[2][27] , \Inst_Mem/inst_mem_reg[2][28] ,
         \Inst_Mem/inst_mem_reg[2][29] , \Inst_Mem/inst_mem_reg[2][30] ,
         \Inst_Mem/inst_mem_reg[2][31] , \Inst_Mem/inst_mem_reg[1][0] ,
         \Inst_Mem/inst_mem_reg[1][1] , \Inst_Mem/inst_mem_reg[1][2] ,
         \Inst_Mem/inst_mem_reg[1][3] , \Inst_Mem/inst_mem_reg[1][4] ,
         \Inst_Mem/inst_mem_reg[1][5] , \Inst_Mem/inst_mem_reg[1][6] ,
         \Inst_Mem/inst_mem_reg[1][7] , \Inst_Mem/inst_mem_reg[1][8] ,
         \Inst_Mem/inst_mem_reg[1][9] , \Inst_Mem/inst_mem_reg[1][10] ,
         \Inst_Mem/inst_mem_reg[1][11] , \Inst_Mem/inst_mem_reg[1][12] ,
         \Inst_Mem/inst_mem_reg[1][13] , \Inst_Mem/inst_mem_reg[1][14] ,
         \Inst_Mem/inst_mem_reg[1][15] , \Inst_Mem/inst_mem_reg[1][16] ,
         \Inst_Mem/inst_mem_reg[1][17] , \Inst_Mem/inst_mem_reg[1][18] ,
         \Inst_Mem/inst_mem_reg[1][19] , \Inst_Mem/inst_mem_reg[1][20] ,
         \Inst_Mem/inst_mem_reg[1][21] , \Inst_Mem/inst_mem_reg[1][22] ,
         \Inst_Mem/inst_mem_reg[1][23] , \Inst_Mem/inst_mem_reg[1][24] ,
         \Inst_Mem/inst_mem_reg[1][25] , \Inst_Mem/inst_mem_reg[1][26] ,
         \Inst_Mem/inst_mem_reg[1][27] , \Inst_Mem/inst_mem_reg[1][28] ,
         \Inst_Mem/inst_mem_reg[1][29] , \Inst_Mem/inst_mem_reg[1][30] ,
         \Inst_Mem/inst_mem_reg[1][31] , \Inst_Mem/inst_mem_reg[0][0] ,
         \Inst_Mem/inst_mem_reg[0][1] , \Inst_Mem/inst_mem_reg[0][2] ,
         \Inst_Mem/inst_mem_reg[0][3] , \Inst_Mem/inst_mem_reg[0][4] ,
         \Inst_Mem/inst_mem_reg[0][5] , \Inst_Mem/inst_mem_reg[0][6] ,
         \Inst_Mem/inst_mem_reg[0][7] , \Inst_Mem/inst_mem_reg[0][8] ,
         \Inst_Mem/inst_mem_reg[0][9] , \Inst_Mem/inst_mem_reg[0][10] ,
         \Inst_Mem/inst_mem_reg[0][11] , \Inst_Mem/inst_mem_reg[0][12] ,
         \Inst_Mem/inst_mem_reg[0][13] , \Inst_Mem/inst_mem_reg[0][14] ,
         \Inst_Mem/inst_mem_reg[0][15] , \Inst_Mem/inst_mem_reg[0][16] ,
         \Inst_Mem/inst_mem_reg[0][17] , \Inst_Mem/inst_mem_reg[0][18] ,
         \Inst_Mem/inst_mem_reg[0][19] , \Inst_Mem/inst_mem_reg[0][20] ,
         \Inst_Mem/inst_mem_reg[0][21] , \Inst_Mem/inst_mem_reg[0][22] ,
         \Inst_Mem/inst_mem_reg[0][23] , \Inst_Mem/inst_mem_reg[0][24] ,
         \Inst_Mem/inst_mem_reg[0][25] , \Inst_Mem/inst_mem_reg[0][26] ,
         \Inst_Mem/inst_mem_reg[0][27] , \Inst_Mem/inst_mem_reg[0][28] ,
         \Inst_Mem/inst_mem_reg[0][29] , \Inst_Mem/inst_mem_reg[0][30] ,
         \Inst_Mem/inst_mem_reg[0][31] , \Data_Mem/n9744 , \Data_Mem/n9743 ,
         \Data_Mem/n9742 , \Data_Mem/n9741 , \Data_Mem/n9740 ,
         \Data_Mem/n9739 , \Data_Mem/n9738 , \Data_Mem/n9737 ,
         \Data_Mem/n9736 , \Data_Mem/n9735 , \Data_Mem/n9734 ,
         \Data_Mem/n9733 , \Data_Mem/n9732 , \Data_Mem/n9731 ,
         \Data_Mem/n9730 , \Data_Mem/n9729 , \Data_Mem/n9728 ,
         \Data_Mem/n9727 , \Data_Mem/n9726 , \Data_Mem/n9725 ,
         \Data_Mem/n9724 , \Data_Mem/n9723 , \Data_Mem/n9722 ,
         \Data_Mem/n9721 , \Data_Mem/n9720 , \Data_Mem/n9719 ,
         \Data_Mem/n9718 , \Data_Mem/n9717 , \Data_Mem/n9716 ,
         \Data_Mem/n9715 , \Data_Mem/n9714 , \Data_Mem/n9713 ,
         \Data_Mem/n9712 , \Data_Mem/n9711 , \Data_Mem/n9710 ,
         \Data_Mem/n9709 , \Data_Mem/n9708 , \Data_Mem/n9707 ,
         \Data_Mem/n9706 , \Data_Mem/n9705 , \Data_Mem/n9704 ,
         \Data_Mem/n9703 , \Data_Mem/n9702 , \Data_Mem/n9701 ,
         \Data_Mem/n9700 , \Data_Mem/n9699 , \Data_Mem/n9698 ,
         \Data_Mem/n9697 , \Data_Mem/n9696 , \Data_Mem/n9695 ,
         \Data_Mem/n9694 , \Data_Mem/n9693 , \Data_Mem/n9692 ,
         \Data_Mem/n9691 , \Data_Mem/n9690 , \Data_Mem/n9689 ,
         \Data_Mem/n9688 , \Data_Mem/n9687 , \Data_Mem/n9686 ,
         \Data_Mem/n9685 , \Data_Mem/n9684 , \Data_Mem/n9683 ,
         \Data_Mem/n9682 , \Data_Mem/n9681 , \Data_Mem/n9680 ,
         \Data_Mem/n9679 , \Data_Mem/n9678 , \Data_Mem/n9677 ,
         \Data_Mem/n9676 , \Data_Mem/n9675 , \Data_Mem/n9674 ,
         \Data_Mem/n9673 , \Data_Mem/n9672 , \Data_Mem/n9671 ,
         \Data_Mem/n9670 , \Data_Mem/n9669 , \Data_Mem/n9668 ,
         \Data_Mem/n9667 , \Data_Mem/n9666 , \Data_Mem/n9665 ,
         \Data_Mem/n9664 , \Data_Mem/n9663 , \Data_Mem/n9662 ,
         \Data_Mem/n9661 , \Data_Mem/n9660 , \Data_Mem/n9659 ,
         \Data_Mem/n9658 , \Data_Mem/n9657 , \Data_Mem/n9656 ,
         \Data_Mem/n9655 , \Data_Mem/n9654 , \Data_Mem/n9653 ,
         \Data_Mem/n9652 , \Data_Mem/n9651 , \Data_Mem/n9650 ,
         \Data_Mem/n9649 , \Data_Mem/n9648 , \Data_Mem/n9647 ,
         \Data_Mem/n9646 , \Data_Mem/n9645 , \Data_Mem/n9644 ,
         \Data_Mem/n9643 , \Data_Mem/n9642 , \Data_Mem/n9641 ,
         \Data_Mem/n9640 , \Data_Mem/n9639 , \Data_Mem/n9638 ,
         \Data_Mem/n9637 , \Data_Mem/n9636 , \Data_Mem/n9635 ,
         \Data_Mem/n9634 , \Data_Mem/n9633 , \Data_Mem/n9632 ,
         \Data_Mem/n9631 , \Data_Mem/n9630 , \Data_Mem/n9629 ,
         \Data_Mem/n9628 , \Data_Mem/n9627 , \Data_Mem/n9626 ,
         \Data_Mem/n9625 , \Data_Mem/n9624 , \Data_Mem/n9623 ,
         \Data_Mem/n9622 , \Data_Mem/n9621 , \Data_Mem/n9620 ,
         \Data_Mem/n9619 , \Data_Mem/n9618 , \Data_Mem/n9617 ,
         \Data_Mem/n9616 , \Data_Mem/n9615 , \Data_Mem/n9614 ,
         \Data_Mem/n9613 , \Data_Mem/n9612 , \Data_Mem/n9611 ,
         \Data_Mem/n9610 , \Data_Mem/n9609 , \Data_Mem/n9608 ,
         \Data_Mem/n9607 , \Data_Mem/n9606 , \Data_Mem/n9605 ,
         \Data_Mem/n9604 , \Data_Mem/n9603 , \Data_Mem/n9602 ,
         \Data_Mem/n9601 , \Data_Mem/n9600 , \Data_Mem/n9599 ,
         \Data_Mem/n9598 , \Data_Mem/n9597 , \Data_Mem/n9596 ,
         \Data_Mem/n9595 , \Data_Mem/n9594 , \Data_Mem/n9593 ,
         \Data_Mem/n9592 , \Data_Mem/n9591 , \Data_Mem/n9590 ,
         \Data_Mem/n9589 , \Data_Mem/n9588 , \Data_Mem/n9587 ,
         \Data_Mem/n9586 , \Data_Mem/n9585 , \Data_Mem/n9584 ,
         \Data_Mem/n9583 , \Data_Mem/n9582 , \Data_Mem/n9581 ,
         \Data_Mem/n9580 , \Data_Mem/n9579 , \Data_Mem/n9578 ,
         \Data_Mem/n9577 , \Data_Mem/n9576 , \Data_Mem/n9575 ,
         \Data_Mem/n9574 , \Data_Mem/n9573 , \Data_Mem/n9572 ,
         \Data_Mem/n9571 , \Data_Mem/n9570 , \Data_Mem/n9569 ,
         \Data_Mem/n9568 , \Data_Mem/n9567 , \Data_Mem/n9566 ,
         \Data_Mem/n9565 , \Data_Mem/n9564 , \Data_Mem/n9563 ,
         \Data_Mem/n9562 , \Data_Mem/n9561 , \Data_Mem/n9560 ,
         \Data_Mem/n9559 , \Data_Mem/n9558 , \Data_Mem/n9557 ,
         \Data_Mem/n9556 , \Data_Mem/n9555 , \Data_Mem/n9554 ,
         \Data_Mem/n9553 , \Data_Mem/n9552 , \Data_Mem/n9551 ,
         \Data_Mem/n9550 , \Data_Mem/n9549 , \Data_Mem/n9548 ,
         \Data_Mem/n9547 , \Data_Mem/n9546 , \Data_Mem/n9545 ,
         \Data_Mem/n9544 , \Data_Mem/n9543 , \Data_Mem/n9542 ,
         \Data_Mem/n9541 , \Data_Mem/n9540 , \Data_Mem/n9539 ,
         \Data_Mem/n9538 , \Data_Mem/n9537 , \Data_Mem/n9536 ,
         \Data_Mem/n9535 , \Data_Mem/n9534 , \Data_Mem/n9533 ,
         \Data_Mem/n9532 , \Data_Mem/n9531 , \Data_Mem/n9530 ,
         \Data_Mem/n9529 , \Data_Mem/n9528 , \Data_Mem/n9527 ,
         \Data_Mem/n9526 , \Data_Mem/n9525 , \Data_Mem/n9524 ,
         \Data_Mem/n9523 , \Data_Mem/n9522 , \Data_Mem/n9521 ,
         \Data_Mem/n9520 , \Data_Mem/n9519 , \Data_Mem/n9518 ,
         \Data_Mem/n9517 , \Data_Mem/n9516 , \Data_Mem/n9515 ,
         \Data_Mem/n9514 , \Data_Mem/n9513 , \Data_Mem/n9512 ,
         \Data_Mem/n9511 , \Data_Mem/n9510 , \Data_Mem/n9509 ,
         \Data_Mem/n9508 , \Data_Mem/n9507 , \Data_Mem/n9506 ,
         \Data_Mem/n9505 , \Data_Mem/n9504 , \Data_Mem/n9503 ,
         \Data_Mem/n9502 , \Data_Mem/n9501 , \Data_Mem/n9500 ,
         \Data_Mem/n9499 , \Data_Mem/n9498 , \Data_Mem/n9497 ,
         \Data_Mem/n9496 , \Data_Mem/n9495 , \Data_Mem/n9494 ,
         \Data_Mem/n9493 , \Data_Mem/n9492 , \Data_Mem/n9491 ,
         \Data_Mem/n9490 , \Data_Mem/n9489 , \Data_Mem/n9488 ,
         \Data_Mem/n9487 , \Data_Mem/n9486 , \Data_Mem/n9485 ,
         \Data_Mem/n9484 , \Data_Mem/n9483 , \Data_Mem/n9482 ,
         \Data_Mem/n9481 , \Data_Mem/n9480 , \Data_Mem/n9479 ,
         \Data_Mem/n9478 , \Data_Mem/n9477 , \Data_Mem/n9476 ,
         \Data_Mem/n9475 , \Data_Mem/n9474 , \Data_Mem/n9473 ,
         \Data_Mem/n9472 , \Data_Mem/n9471 , \Data_Mem/n9470 ,
         \Data_Mem/n9469 , \Data_Mem/n9468 , \Data_Mem/n9467 ,
         \Data_Mem/n9466 , \Data_Mem/n9465 , \Data_Mem/n9464 ,
         \Data_Mem/n9463 , \Data_Mem/n9462 , \Data_Mem/n9461 ,
         \Data_Mem/n9460 , \Data_Mem/n9459 , \Data_Mem/n9458 ,
         \Data_Mem/n9457 , \Data_Mem/n9456 , \Data_Mem/n9455 ,
         \Data_Mem/n9454 , \Data_Mem/n9453 , \Data_Mem/n9452 ,
         \Data_Mem/n9451 , \Data_Mem/n9450 , \Data_Mem/n9449 ,
         \Data_Mem/n9448 , \Data_Mem/n9447 , \Data_Mem/n9446 ,
         \Data_Mem/n9445 , \Data_Mem/n9444 , \Data_Mem/n9443 ,
         \Data_Mem/n9442 , \Data_Mem/n9441 , \Data_Mem/n9440 ,
         \Data_Mem/n9439 , \Data_Mem/n9438 , \Data_Mem/n9437 ,
         \Data_Mem/n9436 , \Data_Mem/n9435 , \Data_Mem/n9434 ,
         \Data_Mem/n9433 , \Data_Mem/n9432 , \Data_Mem/n9431 ,
         \Data_Mem/n9430 , \Data_Mem/n9429 , \Data_Mem/n9428 ,
         \Data_Mem/n9427 , \Data_Mem/n9426 , \Data_Mem/n9425 ,
         \Data_Mem/n9424 , \Data_Mem/n9423 , \Data_Mem/n9422 ,
         \Data_Mem/n9421 , \Data_Mem/n9420 , \Data_Mem/n9419 ,
         \Data_Mem/n9418 , \Data_Mem/n9417 , \Data_Mem/n9416 ,
         \Data_Mem/n9415 , \Data_Mem/n9414 , \Data_Mem/n9413 ,
         \Data_Mem/n9412 , \Data_Mem/n9411 , \Data_Mem/n9410 ,
         \Data_Mem/n9409 , \Data_Mem/n9408 , \Data_Mem/n9407 ,
         \Data_Mem/n9406 , \Data_Mem/n9405 , \Data_Mem/n9404 ,
         \Data_Mem/n9403 , \Data_Mem/n9402 , \Data_Mem/n9401 ,
         \Data_Mem/n9400 , \Data_Mem/n9399 , \Data_Mem/n9398 ,
         \Data_Mem/n9397 , \Data_Mem/n9396 , \Data_Mem/n9395 ,
         \Data_Mem/n9394 , \Data_Mem/n9393 , \Data_Mem/n9392 ,
         \Data_Mem/n9391 , \Data_Mem/n9390 , \Data_Mem/n9389 ,
         \Data_Mem/n9388 , \Data_Mem/n9387 , \Data_Mem/n9386 ,
         \Data_Mem/n9385 , \Data_Mem/n9384 , \Data_Mem/n9383 ,
         \Data_Mem/n9382 , \Data_Mem/n9381 , \Data_Mem/n9380 ,
         \Data_Mem/n9379 , \Data_Mem/n9378 , \Data_Mem/n9377 ,
         \Data_Mem/n9376 , \Data_Mem/n9375 , \Data_Mem/n9374 ,
         \Data_Mem/n9373 , \Data_Mem/n9372 , \Data_Mem/n9371 ,
         \Data_Mem/n9370 , \Data_Mem/n9369 , \Data_Mem/n9368 ,
         \Data_Mem/n9367 , \Data_Mem/n9366 , \Data_Mem/n9365 ,
         \Data_Mem/n9364 , \Data_Mem/n9363 , \Data_Mem/n9362 ,
         \Data_Mem/n9361 , \Data_Mem/n9360 , \Data_Mem/n9359 ,
         \Data_Mem/n9358 , \Data_Mem/n9357 , \Data_Mem/n9356 ,
         \Data_Mem/n9355 , \Data_Mem/n9354 , \Data_Mem/n9353 ,
         \Data_Mem/n9352 , \Data_Mem/n9351 , \Data_Mem/n9350 ,
         \Data_Mem/n9349 , \Data_Mem/n9348 , \Data_Mem/n9347 ,
         \Data_Mem/n9346 , \Data_Mem/n9345 , \Data_Mem/n9344 ,
         \Data_Mem/n9343 , \Data_Mem/n9342 , \Data_Mem/n9341 ,
         \Data_Mem/n9340 , \Data_Mem/n9339 , \Data_Mem/n9338 ,
         \Data_Mem/n9337 , \Data_Mem/n9336 , \Data_Mem/n9335 ,
         \Data_Mem/n9334 , \Data_Mem/n9333 , \Data_Mem/n9332 ,
         \Data_Mem/n9331 , \Data_Mem/n9330 , \Data_Mem/n9329 ,
         \Data_Mem/n9328 , \Data_Mem/n9327 , \Data_Mem/n9326 ,
         \Data_Mem/n9325 , \Data_Mem/n9324 , \Data_Mem/n9323 ,
         \Data_Mem/n9322 , \Data_Mem/n9321 , \Data_Mem/n9320 ,
         \Data_Mem/n9319 , \Data_Mem/n9318 , \Data_Mem/n9317 ,
         \Data_Mem/n9316 , \Data_Mem/n9315 , \Data_Mem/n9314 ,
         \Data_Mem/n9313 , \Data_Mem/n9312 , \Data_Mem/n9311 ,
         \Data_Mem/n9310 , \Data_Mem/n9309 , \Data_Mem/n9308 ,
         \Data_Mem/n9307 , \Data_Mem/n9306 , \Data_Mem/n9305 ,
         \Data_Mem/n9304 , \Data_Mem/n9303 , \Data_Mem/n9302 ,
         \Data_Mem/n9301 , \Data_Mem/n9300 , \Data_Mem/n9299 ,
         \Data_Mem/n9298 , \Data_Mem/n9297 , \Data_Mem/n9296 ,
         \Data_Mem/n9295 , \Data_Mem/n9294 , \Data_Mem/n9293 ,
         \Data_Mem/n9292 , \Data_Mem/n9291 , \Data_Mem/n9290 ,
         \Data_Mem/n9289 , \Data_Mem/n9288 , \Data_Mem/n9287 ,
         \Data_Mem/n9286 , \Data_Mem/n9285 , \Data_Mem/n9284 ,
         \Data_Mem/n9283 , \Data_Mem/n9282 , \Data_Mem/n9281 ,
         \Data_Mem/n9280 , \Data_Mem/n9279 , \Data_Mem/n9278 ,
         \Data_Mem/n9277 , \Data_Mem/n9276 , \Data_Mem/n9275 ,
         \Data_Mem/n9274 , \Data_Mem/n9273 , \Data_Mem/n9272 ,
         \Data_Mem/n9271 , \Data_Mem/n9270 , \Data_Mem/n9269 ,
         \Data_Mem/n9268 , \Data_Mem/n9267 , \Data_Mem/n9266 ,
         \Data_Mem/n9265 , \Data_Mem/n9264 , \Data_Mem/n9263 ,
         \Data_Mem/n9262 , \Data_Mem/n9261 , \Data_Mem/n9260 ,
         \Data_Mem/n9259 , \Data_Mem/n9258 , \Data_Mem/n9257 ,
         \Data_Mem/n9256 , \Data_Mem/n9255 , \Data_Mem/n9254 ,
         \Data_Mem/n9253 , \Data_Mem/n9252 , \Data_Mem/n9251 ,
         \Data_Mem/n9250 , \Data_Mem/n9249 , \Data_Mem/n9248 ,
         \Data_Mem/n9247 , \Data_Mem/n9246 , \Data_Mem/n9245 ,
         \Data_Mem/n9244 , \Data_Mem/n9243 , \Data_Mem/n9242 ,
         \Data_Mem/n9241 , \Data_Mem/n9240 , \Data_Mem/n9239 ,
         \Data_Mem/n9238 , \Data_Mem/n9237 , \Data_Mem/n9236 ,
         \Data_Mem/n9235 , \Data_Mem/n9234 , \Data_Mem/n9233 ,
         \Data_Mem/n9232 , \Data_Mem/n9231 , \Data_Mem/n9230 ,
         \Data_Mem/n9229 , \Data_Mem/n9228 , \Data_Mem/n9227 ,
         \Data_Mem/n9226 , \Data_Mem/n9225 , \Data_Mem/n9224 ,
         \Data_Mem/n9223 , \Data_Mem/n9222 , \Data_Mem/n9221 ,
         \Data_Mem/n9220 , \Data_Mem/n9219 , \Data_Mem/n9218 ,
         \Data_Mem/n9217 , \Data_Mem/n9216 , \Data_Mem/n9215 ,
         \Data_Mem/n9214 , \Data_Mem/n9213 , \Data_Mem/n9212 ,
         \Data_Mem/n9211 , \Data_Mem/n9210 , \Data_Mem/n9209 ,
         \Data_Mem/n9208 , \Data_Mem/n9207 , \Data_Mem/n9206 ,
         \Data_Mem/n9205 , \Data_Mem/n9204 , \Data_Mem/n9203 ,
         \Data_Mem/n9202 , \Data_Mem/n9201 , \Data_Mem/n9200 ,
         \Data_Mem/n9199 , \Data_Mem/n9198 , \Data_Mem/n9197 ,
         \Data_Mem/n9196 , \Data_Mem/n9195 , \Data_Mem/n9194 ,
         \Data_Mem/n9193 , \Data_Mem/n9192 , \Data_Mem/n9191 ,
         \Data_Mem/n9190 , \Data_Mem/n9189 , \Data_Mem/n9188 ,
         \Data_Mem/n9187 , \Data_Mem/n9186 , \Data_Mem/n9185 ,
         \Data_Mem/n9184 , \Data_Mem/n9183 , \Data_Mem/n9182 ,
         \Data_Mem/n9181 , \Data_Mem/n9180 , \Data_Mem/n9179 ,
         \Data_Mem/n9178 , \Data_Mem/n9177 , \Data_Mem/n9176 ,
         \Data_Mem/n9175 , \Data_Mem/n9174 , \Data_Mem/n9173 ,
         \Data_Mem/n9172 , \Data_Mem/n9171 , \Data_Mem/n9170 ,
         \Data_Mem/n9169 , \Data_Mem/n9168 , \Data_Mem/n9167 ,
         \Data_Mem/n9166 , \Data_Mem/n9165 , \Data_Mem/n9164 ,
         \Data_Mem/n9163 , \Data_Mem/n9162 , \Data_Mem/n9161 ,
         \Data_Mem/n9160 , \Data_Mem/n9159 , \Data_Mem/n9158 ,
         \Data_Mem/n9157 , \Data_Mem/n9156 , \Data_Mem/n9155 ,
         \Data_Mem/n9154 , \Data_Mem/n9153 , \Data_Mem/n9152 ,
         \Data_Mem/n9151 , \Data_Mem/n9150 , \Data_Mem/n9149 ,
         \Data_Mem/n9148 , \Data_Mem/n9147 , \Data_Mem/n9146 ,
         \Data_Mem/n9145 , \Data_Mem/n9144 , \Data_Mem/n9143 ,
         \Data_Mem/n9142 , \Data_Mem/n9141 , \Data_Mem/n9140 ,
         \Data_Mem/n9139 , \Data_Mem/n9138 , \Data_Mem/n9137 ,
         \Data_Mem/n9136 , \Data_Mem/n9135 , \Data_Mem/n9134 ,
         \Data_Mem/n9133 , \Data_Mem/n9132 , \Data_Mem/n9131 ,
         \Data_Mem/n9130 , \Data_Mem/n9129 , \Data_Mem/n9128 ,
         \Data_Mem/n9127 , \Data_Mem/n9126 , \Data_Mem/n9125 ,
         \Data_Mem/n9124 , \Data_Mem/n9123 , \Data_Mem/n9122 ,
         \Data_Mem/n9121 , \Data_Mem/n9120 , \Data_Mem/n9119 ,
         \Data_Mem/n9118 , \Data_Mem/n9117 , \Data_Mem/n9116 ,
         \Data_Mem/n9115 , \Data_Mem/n9114 , \Data_Mem/n9113 ,
         \Data_Mem/n9112 , \Data_Mem/n9111 , \Data_Mem/n9110 ,
         \Data_Mem/n9109 , \Data_Mem/n9108 , \Data_Mem/n9107 ,
         \Data_Mem/n9106 , \Data_Mem/n9105 , \Data_Mem/n9104 ,
         \Data_Mem/n9103 , \Data_Mem/n9102 , \Data_Mem/n9101 ,
         \Data_Mem/n9100 , \Data_Mem/n9099 , \Data_Mem/n9098 ,
         \Data_Mem/n9097 , \Data_Mem/n9096 , \Data_Mem/n9095 ,
         \Data_Mem/n9094 , \Data_Mem/n9093 , \Data_Mem/n9092 ,
         \Data_Mem/n9091 , \Data_Mem/n9090 , \Data_Mem/n9089 ,
         \Data_Mem/n9088 , \Data_Mem/n9087 , \Data_Mem/n9086 ,
         \Data_Mem/n9085 , \Data_Mem/n9084 , \Data_Mem/n9083 ,
         \Data_Mem/n9082 , \Data_Mem/n9081 , \Data_Mem/n9080 ,
         \Data_Mem/n9079 , \Data_Mem/n9078 , \Data_Mem/n9077 ,
         \Data_Mem/n9076 , \Data_Mem/n9075 , \Data_Mem/n9074 ,
         \Data_Mem/n9073 , \Data_Mem/n9072 , \Data_Mem/n9071 ,
         \Data_Mem/n9070 , \Data_Mem/n9069 , \Data_Mem/n9068 ,
         \Data_Mem/n9067 , \Data_Mem/n9066 , \Data_Mem/n9065 ,
         \Data_Mem/n9064 , \Data_Mem/n9063 , \Data_Mem/n9062 ,
         \Data_Mem/n9061 , \Data_Mem/n9060 , \Data_Mem/n9059 ,
         \Data_Mem/n9058 , \Data_Mem/n9057 , \Data_Mem/n9056 ,
         \Data_Mem/n9055 , \Data_Mem/n9054 , \Data_Mem/n9053 ,
         \Data_Mem/n9052 , \Data_Mem/n9051 , \Data_Mem/n9050 ,
         \Data_Mem/n9049 , \Data_Mem/n9048 , \Data_Mem/n9047 ,
         \Data_Mem/n9046 , \Data_Mem/n9045 , \Data_Mem/n9044 ,
         \Data_Mem/n9043 , \Data_Mem/n9042 , \Data_Mem/n9041 ,
         \Data_Mem/n9040 , \Data_Mem/n9039 , \Data_Mem/n9038 ,
         \Data_Mem/n9037 , \Data_Mem/n9036 , \Data_Mem/n9035 ,
         \Data_Mem/n9034 , \Data_Mem/n9033 , \Data_Mem/n9032 ,
         \Data_Mem/n9031 , \Data_Mem/n9030 , \Data_Mem/n9029 ,
         \Data_Mem/n9028 , \Data_Mem/n9027 , \Data_Mem/n9026 ,
         \Data_Mem/n9025 , \Data_Mem/n9024 , \Data_Mem/n9023 ,
         \Data_Mem/n9022 , \Data_Mem/n9021 , \Data_Mem/n9020 ,
         \Data_Mem/n9019 , \Data_Mem/n9018 , \Data_Mem/n9017 ,
         \Data_Mem/n9016 , \Data_Mem/n9015 , \Data_Mem/n9014 ,
         \Data_Mem/n9013 , \Data_Mem/n9012 , \Data_Mem/n9011 ,
         \Data_Mem/n9010 , \Data_Mem/n9009 , \Data_Mem/n9008 ,
         \Data_Mem/n9007 , \Data_Mem/n9006 , \Data_Mem/n9005 ,
         \Data_Mem/n9004 , \Data_Mem/n9003 , \Data_Mem/n9002 ,
         \Data_Mem/n9001 , \Data_Mem/n9000 , \Data_Mem/n8999 ,
         \Data_Mem/n8998 , \Data_Mem/n8997 , \Data_Mem/n8996 ,
         \Data_Mem/n8995 , \Data_Mem/n8994 , \Data_Mem/n8993 ,
         \Data_Mem/n8992 , \Data_Mem/n8991 , \Data_Mem/n8990 ,
         \Data_Mem/n8989 , \Data_Mem/n8988 , \Data_Mem/n8987 ,
         \Data_Mem/n8986 , \Data_Mem/n8985 , \Data_Mem/n8984 ,
         \Data_Mem/n8983 , \Data_Mem/n8982 , \Data_Mem/n8981 ,
         \Data_Mem/n8980 , \Data_Mem/n8979 , \Data_Mem/n8978 ,
         \Data_Mem/n8977 , \Data_Mem/n8976 , \Data_Mem/n8975 ,
         \Data_Mem/n8974 , \Data_Mem/n8973 , \Data_Mem/n8972 ,
         \Data_Mem/n8971 , \Data_Mem/n8970 , \Data_Mem/n8969 ,
         \Data_Mem/n8968 , \Data_Mem/n8967 , \Data_Mem/n8966 ,
         \Data_Mem/n8965 , \Data_Mem/n8964 , \Data_Mem/n8963 ,
         \Data_Mem/n8962 , \Data_Mem/n8961 , \Data_Mem/n8960 ,
         \Data_Mem/n8959 , \Data_Mem/n8958 , \Data_Mem/n8957 ,
         \Data_Mem/n8956 , \Data_Mem/n8955 , \Data_Mem/n8954 ,
         \Data_Mem/n8953 , \Data_Mem/n8952 , \Data_Mem/n8951 ,
         \Data_Mem/n8950 , \Data_Mem/n8949 , \Data_Mem/n8948 ,
         \Data_Mem/n8947 , \Data_Mem/n8946 , \Data_Mem/n8945 ,
         \Data_Mem/n8944 , \Data_Mem/n8943 , \Data_Mem/n8942 ,
         \Data_Mem/n8941 , \Data_Mem/n8940 , \Data_Mem/n8939 ,
         \Data_Mem/n8938 , \Data_Mem/n8937 , \Data_Mem/n8936 ,
         \Data_Mem/n8935 , \Data_Mem/n8934 , \Data_Mem/n8933 ,
         \Data_Mem/n8932 , \Data_Mem/n8931 , \Data_Mem/n8930 ,
         \Data_Mem/n8929 , \Data_Mem/n8928 , \Data_Mem/n8927 ,
         \Data_Mem/n8926 , \Data_Mem/n8925 , \Data_Mem/n8924 ,
         \Data_Mem/n8923 , \Data_Mem/n8922 , \Data_Mem/n8921 ,
         \Data_Mem/n8920 , \Data_Mem/n8919 , \Data_Mem/n8918 ,
         \Data_Mem/n8917 , \Data_Mem/n8916 , \Data_Mem/n8915 ,
         \Data_Mem/n8914 , \Data_Mem/n8913 , \Data_Mem/n8912 ,
         \Data_Mem/n8911 , \Data_Mem/n8910 , \Data_Mem/n8909 ,
         \Data_Mem/n8908 , \Data_Mem/n8907 , \Data_Mem/n8906 ,
         \Data_Mem/n8905 , \Data_Mem/n8904 , \Data_Mem/n8903 ,
         \Data_Mem/n8902 , \Data_Mem/n8901 , \Data_Mem/n8900 ,
         \Data_Mem/n8899 , \Data_Mem/n8898 , \Data_Mem/n8897 ,
         \Data_Mem/n8896 , \Data_Mem/n8895 , \Data_Mem/n8894 ,
         \Data_Mem/n8893 , \Data_Mem/n8892 , \Data_Mem/n8891 ,
         \Data_Mem/n8890 , \Data_Mem/n8889 , \Data_Mem/n8888 ,
         \Data_Mem/n8887 , \Data_Mem/n8886 , \Data_Mem/n8885 ,
         \Data_Mem/n8884 , \Data_Mem/n8883 , \Data_Mem/n8882 ,
         \Data_Mem/n8881 , \Data_Mem/n8880 , \Data_Mem/n8879 ,
         \Data_Mem/n8878 , \Data_Mem/n8877 , \Data_Mem/n8876 ,
         \Data_Mem/n8875 , \Data_Mem/n8874 , \Data_Mem/n8873 ,
         \Data_Mem/n8872 , \Data_Mem/n8871 , \Data_Mem/n8870 ,
         \Data_Mem/n8869 , \Data_Mem/n8868 , \Data_Mem/n8867 ,
         \Data_Mem/n8866 , \Data_Mem/n8865 , \Data_Mem/n8864 ,
         \Data_Mem/n8863 , \Data_Mem/n8862 , \Data_Mem/n8861 ,
         \Data_Mem/n8860 , \Data_Mem/n8859 , \Data_Mem/n8858 ,
         \Data_Mem/n8857 , \Data_Mem/n8856 , \Data_Mem/n8855 ,
         \Data_Mem/n8854 , \Data_Mem/n8853 , \Data_Mem/n8852 ,
         \Data_Mem/n8851 , \Data_Mem/n8850 , \Data_Mem/n8849 ,
         \Data_Mem/n8848 , \Data_Mem/n8847 , \Data_Mem/n8846 ,
         \Data_Mem/n8845 , \Data_Mem/n8844 , \Data_Mem/n8843 ,
         \Data_Mem/n8842 , \Data_Mem/n8841 , \Data_Mem/n8840 ,
         \Data_Mem/n8839 , \Data_Mem/n8838 , \Data_Mem/n8837 ,
         \Data_Mem/n8836 , \Data_Mem/n8835 , \Data_Mem/n8834 ,
         \Data_Mem/n8833 , \Data_Mem/n8832 , \Data_Mem/n8831 ,
         \Data_Mem/n8830 , \Data_Mem/n8829 , \Data_Mem/n8828 ,
         \Data_Mem/n8827 , \Data_Mem/n8826 , \Data_Mem/n8825 ,
         \Data_Mem/n8824 , \Data_Mem/n8823 , \Data_Mem/n8822 ,
         \Data_Mem/n8821 , \Data_Mem/n8820 , \Data_Mem/n8819 ,
         \Data_Mem/n8818 , \Data_Mem/n8817 , \Data_Mem/n8816 ,
         \Data_Mem/n8815 , \Data_Mem/n8814 , \Data_Mem/n8813 ,
         \Data_Mem/n8812 , \Data_Mem/n8811 , \Data_Mem/n8810 ,
         \Data_Mem/n8809 , \Data_Mem/n8808 , \Data_Mem/n8807 ,
         \Data_Mem/n8806 , \Data_Mem/n8805 , \Data_Mem/n8804 ,
         \Data_Mem/n8803 , \Data_Mem/n8802 , \Data_Mem/n8801 ,
         \Data_Mem/n8800 , \Data_Mem/n8799 , \Data_Mem/n8798 ,
         \Data_Mem/n8797 , \Data_Mem/n8796 , \Data_Mem/n8795 ,
         \Data_Mem/n8794 , \Data_Mem/n8793 , \Data_Mem/n8792 ,
         \Data_Mem/n8791 , \Data_Mem/n8790 , \Data_Mem/n8789 ,
         \Data_Mem/n8788 , \Data_Mem/n8787 , \Data_Mem/n8786 ,
         \Data_Mem/n8785 , \Data_Mem/n8784 , \Data_Mem/n8783 ,
         \Data_Mem/n8782 , \Data_Mem/n8781 , \Data_Mem/n8780 ,
         \Data_Mem/n8779 , \Data_Mem/n8778 , \Data_Mem/n8777 ,
         \Data_Mem/n8776 , \Data_Mem/n8775 , \Data_Mem/n8774 ,
         \Data_Mem/n8773 , \Data_Mem/n8772 , \Data_Mem/n8771 ,
         \Data_Mem/n8770 , \Data_Mem/n8769 , \Data_Mem/n8768 ,
         \Data_Mem/n8767 , \Data_Mem/n8766 , \Data_Mem/n8765 ,
         \Data_Mem/n8764 , \Data_Mem/n8763 , \Data_Mem/n8762 ,
         \Data_Mem/n8761 , \Data_Mem/n8760 , \Data_Mem/n8759 ,
         \Data_Mem/n8758 , \Data_Mem/n8757 , \Data_Mem/n8756 ,
         \Data_Mem/n8755 , \Data_Mem/n8754 , \Data_Mem/n8753 ,
         \Data_Mem/n8752 , \Data_Mem/n8751 , \Data_Mem/n8750 ,
         \Data_Mem/n8749 , \Data_Mem/n8748 , \Data_Mem/n8747 ,
         \Data_Mem/n8746 , \Data_Mem/n8745 , \Data_Mem/n8744 ,
         \Data_Mem/n8743 , \Data_Mem/n8742 , \Data_Mem/n8741 ,
         \Data_Mem/n8740 , \Data_Mem/n8739 , \Data_Mem/n8738 ,
         \Data_Mem/n8737 , \Data_Mem/n8736 , \Data_Mem/n8735 ,
         \Data_Mem/n8734 , \Data_Mem/n8733 , \Data_Mem/n8732 ,
         \Data_Mem/n8731 , \Data_Mem/n8730 , \Data_Mem/n8729 ,
         \Data_Mem/n8728 , \Data_Mem/n8727 , \Data_Mem/n8726 ,
         \Data_Mem/n8725 , \Data_Mem/n8724 , \Data_Mem/n8723 ,
         \Data_Mem/n8722 , \Data_Mem/n8721 , \Data_Mem/n8720 ,
         \Data_Mem/n8719 , \Data_Mem/n8718 , \Data_Mem/n8717 ,
         \Data_Mem/n8716 , \Data_Mem/n8715 , \Data_Mem/n8714 ,
         \Data_Mem/n8713 , \Data_Mem/n8712 , \Data_Mem/n8711 ,
         \Data_Mem/n8710 , \Data_Mem/n8709 , \Data_Mem/n8708 ,
         \Data_Mem/n8707 , \Data_Mem/n8706 , \Data_Mem/n8705 ,
         \Data_Mem/n8704 , \Data_Mem/n8703 , \Data_Mem/n8702 ,
         \Data_Mem/n8701 , \Data_Mem/n8700 , \Data_Mem/n8699 ,
         \Data_Mem/n8698 , \Data_Mem/n8697 , \Data_Mem/n8696 ,
         \Data_Mem/n8695 , \Data_Mem/n8694 , \Data_Mem/n8693 ,
         \Data_Mem/n8692 , \Data_Mem/n8691 , \Data_Mem/n8690 ,
         \Data_Mem/n8689 , \Data_Mem/n8688 , \Data_Mem/n8687 ,
         \Data_Mem/n8686 , \Data_Mem/n8685 , \Data_Mem/n8684 ,
         \Data_Mem/n8683 , \Data_Mem/n8682 , \Data_Mem/n8681 ,
         \Data_Mem/n8680 , \Data_Mem/n8679 , \Data_Mem/n8678 ,
         \Data_Mem/n8677 , \Data_Mem/n8676 , \Data_Mem/n8675 ,
         \Data_Mem/n8674 , \Data_Mem/n8673 , \Data_Mem/n8672 ,
         \Data_Mem/n8671 , \Data_Mem/n8670 , \Data_Mem/n8669 ,
         \Data_Mem/n8668 , \Data_Mem/n8667 , \Data_Mem/n8666 ,
         \Data_Mem/n8665 , \Data_Mem/n8664 , \Data_Mem/n8663 ,
         \Data_Mem/n8662 , \Data_Mem/n8661 , \Data_Mem/n8660 ,
         \Data_Mem/n8659 , \Data_Mem/n8658 , \Data_Mem/n8657 ,
         \Data_Mem/n8656 , \Data_Mem/n8655 , \Data_Mem/n8654 ,
         \Data_Mem/n8653 , \Data_Mem/n8652 , \Data_Mem/n8651 ,
         \Data_Mem/n8650 , \Data_Mem/n8649 , \Data_Mem/n8648 ,
         \Data_Mem/n8647 , \Data_Mem/n8646 , \Data_Mem/n8645 ,
         \Data_Mem/n8644 , \Data_Mem/n8643 , \Data_Mem/n8642 ,
         \Data_Mem/n8641 , \Data_Mem/n8640 , \Data_Mem/n8639 ,
         \Data_Mem/n8638 , \Data_Mem/n8637 , \Data_Mem/n8636 ,
         \Data_Mem/n8635 , \Data_Mem/n8634 , \Data_Mem/n8633 ,
         \Data_Mem/n8632 , \Data_Mem/n8631 , \Data_Mem/n8630 ,
         \Data_Mem/n8629 , \Data_Mem/n8628 , \Data_Mem/n8627 ,
         \Data_Mem/n8626 , \Data_Mem/n8625 , \Data_Mem/n8624 ,
         \Data_Mem/n8623 , \Data_Mem/n8622 , \Data_Mem/n8621 ,
         \Data_Mem/n8620 , \Data_Mem/n8619 , \Data_Mem/n8618 ,
         \Data_Mem/n8617 , \Data_Mem/n8616 , \Data_Mem/n8615 ,
         \Data_Mem/n8614 , \Data_Mem/n8613 , \Data_Mem/n8612 ,
         \Data_Mem/n8611 , \Data_Mem/n8610 , \Data_Mem/n8609 ,
         \Data_Mem/n8608 , \Data_Mem/n8607 , \Data_Mem/n8606 ,
         \Data_Mem/n8605 , \Data_Mem/n8604 , \Data_Mem/n8603 ,
         \Data_Mem/n8602 , \Data_Mem/n8601 , \Data_Mem/n8600 ,
         \Data_Mem/n8599 , \Data_Mem/n8598 , \Data_Mem/n8597 ,
         \Data_Mem/n8596 , \Data_Mem/n8595 , \Data_Mem/n8594 ,
         \Data_Mem/n8593 , \Data_Mem/n8592 , \Data_Mem/n8591 ,
         \Data_Mem/n8590 , \Data_Mem/n8589 , \Data_Mem/n8588 ,
         \Data_Mem/n8587 , \Data_Mem/n8586 , \Data_Mem/n8585 ,
         \Data_Mem/n8584 , \Data_Mem/n8583 , \Data_Mem/n8582 ,
         \Data_Mem/n8581 , \Data_Mem/n8580 , \Data_Mem/n8579 ,
         \Data_Mem/n8578 , \Data_Mem/n8577 , \Data_Mem/n8576 ,
         \Data_Mem/n8575 , \Data_Mem/n8574 , \Data_Mem/n8573 ,
         \Data_Mem/n8572 , \Data_Mem/n8571 , \Data_Mem/n8570 ,
         \Data_Mem/n8569 , \Data_Mem/n8568 , \Data_Mem/n8567 ,
         \Data_Mem/n8566 , \Data_Mem/n8565 , \Data_Mem/n8564 ,
         \Data_Mem/n8563 , \Data_Mem/n8562 , \Data_Mem/n8561 ,
         \Data_Mem/n8560 , \Data_Mem/n8559 , \Data_Mem/n8558 ,
         \Data_Mem/n8557 , \Data_Mem/n8556 , \Data_Mem/n8555 ,
         \Data_Mem/n8554 , \Data_Mem/n8553 , \Data_Mem/n8552 ,
         \Data_Mem/n8551 , \Data_Mem/n8550 , \Data_Mem/n8549 ,
         \Data_Mem/n8548 , \Data_Mem/n8547 , \Data_Mem/n8546 ,
         \Data_Mem/n8545 , \Data_Mem/n8544 , \Data_Mem/n8543 ,
         \Data_Mem/n8542 , \Data_Mem/n8541 , \Data_Mem/n8540 ,
         \Data_Mem/n8539 , \Data_Mem/n8538 , \Data_Mem/n8537 ,
         \Data_Mem/n8536 , \Data_Mem/n8535 , \Data_Mem/n8534 ,
         \Data_Mem/n8533 , \Data_Mem/n8532 , \Data_Mem/n8531 ,
         \Data_Mem/n8530 , \Data_Mem/n8529 , \Data_Mem/n8528 ,
         \Data_Mem/n8527 , \Data_Mem/n8526 , \Data_Mem/n8525 ,
         \Data_Mem/n8524 , \Data_Mem/n8523 , \Data_Mem/n8522 ,
         \Data_Mem/n8521 , \Data_Mem/n8520 , \Data_Mem/n8519 ,
         \Data_Mem/n8518 , \Data_Mem/n8517 , \Data_Mem/n8516 ,
         \Data_Mem/n8515 , \Data_Mem/n8514 , \Data_Mem/n8513 ,
         \Data_Mem/n8512 , \Data_Mem/n8511 , \Data_Mem/n8510 ,
         \Data_Mem/n8509 , \Data_Mem/n8508 , \Data_Mem/n8507 ,
         \Data_Mem/n8506 , \Data_Mem/n8505 , \Data_Mem/n8504 ,
         \Data_Mem/n8503 , \Data_Mem/n8502 , \Data_Mem/n8501 ,
         \Data_Mem/n8500 , \Data_Mem/n8499 , \Data_Mem/n8498 ,
         \Data_Mem/n8497 , \Data_Mem/n8496 , \Data_Mem/n8495 ,
         \Data_Mem/n8494 , \Data_Mem/n8493 , \Data_Mem/n8492 ,
         \Data_Mem/n8491 , \Data_Mem/n8490 , \Data_Mem/n8489 ,
         \Data_Mem/n8488 , \Data_Mem/n8487 , \Data_Mem/n8486 ,
         \Data_Mem/n8485 , \Data_Mem/n8484 , \Data_Mem/n8483 ,
         \Data_Mem/n8482 , \Data_Mem/n8481 , \Data_Mem/n8480 ,
         \Data_Mem/n8479 , \Data_Mem/n8478 , \Data_Mem/n8477 ,
         \Data_Mem/n8476 , \Data_Mem/n8475 , \Data_Mem/n8474 ,
         \Data_Mem/n8473 , \Data_Mem/n8472 , \Data_Mem/n8471 ,
         \Data_Mem/n8470 , \Data_Mem/n8469 , \Data_Mem/n8468 ,
         \Data_Mem/n8467 , \Data_Mem/n8466 , \Data_Mem/n8465 ,
         \Data_Mem/n8464 , \Data_Mem/n8463 , \Data_Mem/n8462 ,
         \Data_Mem/n8461 , \Data_Mem/n8460 , \Data_Mem/n8459 ,
         \Data_Mem/n8458 , \Data_Mem/n8457 , \Data_Mem/n8456 ,
         \Data_Mem/n8455 , \Data_Mem/n8454 , \Data_Mem/n8453 ,
         \Data_Mem/n8452 , \Data_Mem/n8451 , \Data_Mem/n8450 ,
         \Data_Mem/n8449 , \Data_Mem/n8448 , \Data_Mem/n8447 ,
         \Data_Mem/n8446 , \Data_Mem/n8445 , \Data_Mem/n8444 ,
         \Data_Mem/n8443 , \Data_Mem/n8442 , \Data_Mem/n8441 ,
         \Data_Mem/n8440 , \Data_Mem/n8439 , \Data_Mem/n8438 ,
         \Data_Mem/n8437 , \Data_Mem/n8436 , \Data_Mem/n8435 ,
         \Data_Mem/n8434 , \Data_Mem/n8433 , \Data_Mem/n8432 ,
         \Data_Mem/n8431 , \Data_Mem/n8430 , \Data_Mem/n8429 ,
         \Data_Mem/n8428 , \Data_Mem/n8427 , \Data_Mem/n8426 ,
         \Data_Mem/n8425 , \Data_Mem/n8424 , \Data_Mem/n8423 ,
         \Data_Mem/n8422 , \Data_Mem/n8421 , \Data_Mem/n8420 ,
         \Data_Mem/n8419 , \Data_Mem/n8418 , \Data_Mem/n8417 ,
         \Data_Mem/n8416 , \Data_Mem/n8415 , \Data_Mem/n8414 ,
         \Data_Mem/n8413 , \Data_Mem/n8412 , \Data_Mem/n8411 ,
         \Data_Mem/n8410 , \Data_Mem/n8409 , \Data_Mem/n8408 ,
         \Data_Mem/n8407 , \Data_Mem/n8406 , \Data_Mem/n8405 ,
         \Data_Mem/n8404 , \Data_Mem/n8403 , \Data_Mem/n8402 ,
         \Data_Mem/n8401 , \Data_Mem/n8400 , \Data_Mem/n8399 ,
         \Data_Mem/n8398 , \Data_Mem/n8397 , \Data_Mem/n8396 ,
         \Data_Mem/n8395 , \Data_Mem/n8394 , \Data_Mem/n8393 ,
         \Data_Mem/n8392 , \Data_Mem/n8391 , \Data_Mem/n8390 ,
         \Data_Mem/n8389 , \Data_Mem/n8388 , \Data_Mem/n8387 ,
         \Data_Mem/n8386 , \Data_Mem/n8385 , \Data_Mem/n8384 ,
         \Data_Mem/n8383 , \Data_Mem/n8382 , \Data_Mem/n8381 ,
         \Data_Mem/n8380 , \Data_Mem/n8379 , \Data_Mem/n8378 ,
         \Data_Mem/n8377 , \Data_Mem/n8376 , \Data_Mem/n8375 ,
         \Data_Mem/n8374 , \Data_Mem/n8373 , \Data_Mem/n8372 ,
         \Data_Mem/n8371 , \Data_Mem/n8370 , \Data_Mem/n8369 ,
         \Data_Mem/n8368 , \Data_Mem/n8367 , \Data_Mem/n8366 ,
         \Data_Mem/n8365 , \Data_Mem/n8364 , \Data_Mem/n8363 ,
         \Data_Mem/n8362 , \Data_Mem/n8361 , \Data_Mem/n8360 ,
         \Data_Mem/n8359 , \Data_Mem/n8358 , \Data_Mem/n8357 ,
         \Data_Mem/n8356 , \Data_Mem/n8355 , \Data_Mem/n8354 ,
         \Data_Mem/n8353 , \Data_Mem/n8352 , \Data_Mem/n8351 ,
         \Data_Mem/n8350 , \Data_Mem/n8349 , \Data_Mem/n8348 ,
         \Data_Mem/n8347 , \Data_Mem/n8346 , \Data_Mem/n8345 ,
         \Data_Mem/n8344 , \Data_Mem/n8343 , \Data_Mem/n8342 ,
         \Data_Mem/n8341 , \Data_Mem/n8340 , \Data_Mem/n8339 ,
         \Data_Mem/n8338 , \Data_Mem/n8337 , \Data_Mem/n8336 ,
         \Data_Mem/n8335 , \Data_Mem/n8334 , \Data_Mem/n8333 ,
         \Data_Mem/n8332 , \Data_Mem/n8331 , \Data_Mem/n8330 ,
         \Data_Mem/n8329 , \Data_Mem/n8328 , \Data_Mem/n8327 ,
         \Data_Mem/n8326 , \Data_Mem/n8325 , \Data_Mem/n8324 ,
         \Data_Mem/n8323 , \Data_Mem/n8322 , \Data_Mem/n8321 ,
         \Data_Mem/n8320 , \Data_Mem/n8319 , \Data_Mem/n8318 ,
         \Data_Mem/n8317 , \Data_Mem/n8316 , \Data_Mem/n8315 ,
         \Data_Mem/n8314 , \Data_Mem/n8313 , \Data_Mem/n8312 ,
         \Data_Mem/n8311 , \Data_Mem/n8310 , \Data_Mem/n8309 ,
         \Data_Mem/n8308 , \Data_Mem/n8307 , \Data_Mem/n8306 ,
         \Data_Mem/n8305 , \Data_Mem/n8304 , \Data_Mem/n8303 ,
         \Data_Mem/n8302 , \Data_Mem/n8301 , \Data_Mem/n8300 ,
         \Data_Mem/n8299 , \Data_Mem/n8298 , \Data_Mem/n8297 ,
         \Data_Mem/n8296 , \Data_Mem/n8295 , \Data_Mem/n8294 ,
         \Data_Mem/n8293 , \Data_Mem/n8292 , \Data_Mem/n8291 ,
         \Data_Mem/n8290 , \Data_Mem/n8289 , \Data_Mem/n8288 ,
         \Data_Mem/n8287 , \Data_Mem/n8286 , \Data_Mem/n8285 ,
         \Data_Mem/n8284 , \Data_Mem/n8283 , \Data_Mem/n8282 ,
         \Data_Mem/n8281 , \Data_Mem/n8280 , \Data_Mem/n8279 ,
         \Data_Mem/n8278 , \Data_Mem/n8277 , \Data_Mem/n8276 ,
         \Data_Mem/n8275 , \Data_Mem/n8274 , \Data_Mem/n8273 ,
         \Data_Mem/n8272 , \Data_Mem/n8271 , \Data_Mem/n8270 ,
         \Data_Mem/n8269 , \Data_Mem/n8268 , \Data_Mem/n8267 ,
         \Data_Mem/n8266 , \Data_Mem/n8265 , \Data_Mem/n8264 ,
         \Data_Mem/n8263 , \Data_Mem/n8262 , \Data_Mem/n8261 ,
         \Data_Mem/n8260 , \Data_Mem/n8259 , \Data_Mem/n8258 ,
         \Data_Mem/n8257 , \Data_Mem/n8256 , \Data_Mem/n8255 ,
         \Data_Mem/n8254 , \Data_Mem/n8253 , \Data_Mem/n8252 ,
         \Data_Mem/n8251 , \Data_Mem/n8250 , \Data_Mem/n8249 ,
         \Data_Mem/n8248 , \Data_Mem/n8247 , \Data_Mem/n8246 ,
         \Data_Mem/n8245 , \Data_Mem/n8244 , \Data_Mem/n8243 ,
         \Data_Mem/n8242 , \Data_Mem/n8241 , \Data_Mem/n8240 ,
         \Data_Mem/n8239 , \Data_Mem/n8238 , \Data_Mem/n8237 ,
         \Data_Mem/n8236 , \Data_Mem/n8235 , \Data_Mem/n8234 ,
         \Data_Mem/n8233 , \Data_Mem/n8232 , \Data_Mem/n8231 ,
         \Data_Mem/n8230 , \Data_Mem/n8229 , \Data_Mem/n8228 ,
         \Data_Mem/n8227 , \Data_Mem/n8226 , \Data_Mem/n8225 ,
         \Data_Mem/n8224 , \Data_Mem/n8223 , \Data_Mem/n8222 ,
         \Data_Mem/n8221 , \Data_Mem/n8220 , \Data_Mem/n8219 ,
         \Data_Mem/n8218 , \Data_Mem/n8217 , \Data_Mem/n8216 ,
         \Data_Mem/n8215 , \Data_Mem/n8214 , \Data_Mem/n8213 ,
         \Data_Mem/n8212 , \Data_Mem/n8211 , \Data_Mem/n8210 ,
         \Data_Mem/n8209 , \Data_Mem/n8208 , \Data_Mem/n8207 ,
         \Data_Mem/n8206 , \Data_Mem/n8205 , \Data_Mem/n8204 ,
         \Data_Mem/n8203 , \Data_Mem/n8202 , \Data_Mem/n8201 ,
         \Data_Mem/n8200 , \Data_Mem/n8199 , \Data_Mem/n8198 ,
         \Data_Mem/n8197 , \Data_Mem/n8196 , \Data_Mem/n8195 ,
         \Data_Mem/n8194 , \Data_Mem/n8193 , \Data_Mem/n8192 ,
         \Data_Mem/n8191 , \Data_Mem/n8190 , \Data_Mem/n8189 ,
         \Data_Mem/n8188 , \Data_Mem/n8187 , \Data_Mem/n8186 ,
         \Data_Mem/n8185 , \Data_Mem/n8184 , \Data_Mem/n8183 ,
         \Data_Mem/n8182 , \Data_Mem/n8181 , \Data_Mem/n8180 ,
         \Data_Mem/n8179 , \Data_Mem/n8178 , \Data_Mem/n8177 ,
         \Data_Mem/n8176 , \Data_Mem/n8175 , \Data_Mem/n8174 ,
         \Data_Mem/n8173 , \Data_Mem/n8172 , \Data_Mem/n8171 ,
         \Data_Mem/n8170 , \Data_Mem/n8169 , \Data_Mem/n8168 ,
         \Data_Mem/n8167 , \Data_Mem/n8166 , \Data_Mem/n8165 ,
         \Data_Mem/n8164 , \Data_Mem/n8163 , \Data_Mem/n8162 ,
         \Data_Mem/n8161 , \Data_Mem/n8160 , \Data_Mem/n8159 ,
         \Data_Mem/n8158 , \Data_Mem/n8157 , \Data_Mem/n8156 ,
         \Data_Mem/n8155 , \Data_Mem/n8154 , \Data_Mem/n8153 ,
         \Data_Mem/n8152 , \Data_Mem/n8151 , \Data_Mem/n8150 ,
         \Data_Mem/n8149 , \Data_Mem/n8148 , \Data_Mem/n8147 ,
         \Data_Mem/n8146 , \Data_Mem/n8145 , \Data_Mem/n8144 ,
         \Data_Mem/n8143 , \Data_Mem/n8142 , \Data_Mem/n8141 ,
         \Data_Mem/n8140 , \Data_Mem/n8139 , \Data_Mem/n8138 ,
         \Data_Mem/n8137 , \Data_Mem/n8136 , \Data_Mem/n8135 ,
         \Data_Mem/n8134 , \Data_Mem/n8133 , \Data_Mem/n8132 ,
         \Data_Mem/n8131 , \Data_Mem/n8130 , \Data_Mem/n8129 ,
         \Data_Mem/n8128 , \Data_Mem/n8127 , \Data_Mem/n8126 ,
         \Data_Mem/n8125 , \Data_Mem/n8124 , \Data_Mem/n8123 ,
         \Data_Mem/n8122 , \Data_Mem/n8121 , \Data_Mem/n8120 ,
         \Data_Mem/n8119 , \Data_Mem/n8118 , \Data_Mem/n8117 ,
         \Data_Mem/n8116 , \Data_Mem/n8115 , \Data_Mem/n8114 ,
         \Data_Mem/n8113 , \Data_Mem/n8112 , \Data_Mem/n8111 ,
         \Data_Mem/n8110 , \Data_Mem/n8109 , \Data_Mem/n8108 ,
         \Data_Mem/n8107 , \Data_Mem/n8106 , \Data_Mem/n8105 ,
         \Data_Mem/n8104 , \Data_Mem/n8103 , \Data_Mem/n8102 ,
         \Data_Mem/n8101 , \Data_Mem/n8100 , \Data_Mem/n8099 ,
         \Data_Mem/n8098 , \Data_Mem/n8097 , \Data_Mem/n8096 ,
         \Data_Mem/n8095 , \Data_Mem/n8094 , \Data_Mem/n8093 ,
         \Data_Mem/n8092 , \Data_Mem/n8091 , \Data_Mem/n8090 ,
         \Data_Mem/n8089 , \Data_Mem/n8088 , \Data_Mem/n8087 ,
         \Data_Mem/n8086 , \Data_Mem/n8085 , \Data_Mem/n8084 ,
         \Data_Mem/n8083 , \Data_Mem/n8082 , \Data_Mem/n8081 ,
         \Data_Mem/n8080 , \Data_Mem/n8079 , \Data_Mem/n8078 ,
         \Data_Mem/n8077 , \Data_Mem/n8076 , \Data_Mem/n8075 ,
         \Data_Mem/n8074 , \Data_Mem/n8073 , \Data_Mem/n8072 ,
         \Data_Mem/n8071 , \Data_Mem/n8070 , \Data_Mem/n8069 ,
         \Data_Mem/n8068 , \Data_Mem/n8067 , \Data_Mem/n8066 ,
         \Data_Mem/n8065 , \Data_Mem/n8064 , \Data_Mem/n8063 ,
         \Data_Mem/n8062 , \Data_Mem/n8061 , \Data_Mem/n8060 ,
         \Data_Mem/n8059 , \Data_Mem/n8058 , \Data_Mem/n8057 ,
         \Data_Mem/n8056 , \Data_Mem/n8055 , \Data_Mem/n8054 ,
         \Data_Mem/n8053 , \Data_Mem/n8052 , \Data_Mem/n8051 ,
         \Data_Mem/n8050 , \Data_Mem/n8049 , \Data_Mem/n8048 ,
         \Data_Mem/n8047 , \Data_Mem/n8046 , \Data_Mem/n8045 ,
         \Data_Mem/n8044 , \Data_Mem/n8043 , \Data_Mem/n8042 ,
         \Data_Mem/n8041 , \Data_Mem/n8040 , \Data_Mem/n8039 ,
         \Data_Mem/n8038 , \Data_Mem/n8037 , \Data_Mem/n8036 ,
         \Data_Mem/n8035 , \Data_Mem/n8034 , \Data_Mem/n8033 ,
         \Data_Mem/n8032 , \Data_Mem/n8031 , \Data_Mem/n8030 ,
         \Data_Mem/n8029 , \Data_Mem/n8028 , \Data_Mem/n8027 ,
         \Data_Mem/n8026 , \Data_Mem/n8025 , \Data_Mem/n8024 ,
         \Data_Mem/n8023 , \Data_Mem/n8022 , \Data_Mem/n8021 ,
         \Data_Mem/n8020 , \Data_Mem/n8019 , \Data_Mem/n8018 ,
         \Data_Mem/n8017 , \Data_Mem/n8016 , \Data_Mem/n8015 ,
         \Data_Mem/n8014 , \Data_Mem/n8013 , \Data_Mem/n8012 ,
         \Data_Mem/n8011 , \Data_Mem/n8010 , \Data_Mem/n8009 ,
         \Data_Mem/n8008 , \Data_Mem/n8007 , \Data_Mem/n8006 ,
         \Data_Mem/n8005 , \Data_Mem/n8004 , \Data_Mem/n8003 ,
         \Data_Mem/n8002 , \Data_Mem/n8001 , \Data_Mem/n8000 ,
         \Data_Mem/n7999 , \Data_Mem/n7998 , \Data_Mem/n7997 ,
         \Data_Mem/n7996 , \Data_Mem/n7995 , \Data_Mem/n7994 ,
         \Data_Mem/n7993 , \Data_Mem/n7992 , \Data_Mem/n7991 ,
         \Data_Mem/n7990 , \Data_Mem/n7989 , \Data_Mem/n7988 ,
         \Data_Mem/n7987 , \Data_Mem/n7986 , \Data_Mem/n7985 ,
         \Data_Mem/n7984 , \Data_Mem/n7983 , \Data_Mem/n7982 ,
         \Data_Mem/n7981 , \Data_Mem/n7980 , \Data_Mem/n7979 ,
         \Data_Mem/n7978 , \Data_Mem/n7977 , \Data_Mem/n7976 ,
         \Data_Mem/n7975 , \Data_Mem/n7974 , \Data_Mem/n7973 ,
         \Data_Mem/n7972 , \Data_Mem/n7971 , \Data_Mem/n7970 ,
         \Data_Mem/n7969 , \Data_Mem/n7968 , \Data_Mem/n7967 ,
         \Data_Mem/n7966 , \Data_Mem/n7965 , \Data_Mem/n7964 ,
         \Data_Mem/n7963 , \Data_Mem/n7962 , \Data_Mem/n7961 ,
         \Data_Mem/n7960 , \Data_Mem/n7959 , \Data_Mem/n7958 ,
         \Data_Mem/n7957 , \Data_Mem/n7956 , \Data_Mem/n7955 ,
         \Data_Mem/n7954 , \Data_Mem/n7953 , \Data_Mem/n7952 ,
         \Data_Mem/n7951 , \Data_Mem/n7950 , \Data_Mem/n7949 ,
         \Data_Mem/n7948 , \Data_Mem/n7947 , \Data_Mem/n7946 ,
         \Data_Mem/n7945 , \Data_Mem/n7944 , \Data_Mem/n7943 ,
         \Data_Mem/n7942 , \Data_Mem/n7941 , \Data_Mem/n7940 ,
         \Data_Mem/n7939 , \Data_Mem/n7938 , \Data_Mem/n7937 ,
         \Data_Mem/n7936 , \Data_Mem/n7935 , \Data_Mem/n7934 ,
         \Data_Mem/n7933 , \Data_Mem/n7932 , \Data_Mem/n7931 ,
         \Data_Mem/n7930 , \Data_Mem/n7929 , \Data_Mem/n7928 ,
         \Data_Mem/n7927 , \Data_Mem/n7926 , \Data_Mem/n7925 ,
         \Data_Mem/n7924 , \Data_Mem/n7923 , \Data_Mem/n7922 ,
         \Data_Mem/n7921 , \Data_Mem/n7920 , \Data_Mem/n7919 ,
         \Data_Mem/n7918 , \Data_Mem/n7917 , \Data_Mem/n7916 ,
         \Data_Mem/n7915 , \Data_Mem/n7914 , \Data_Mem/n7913 ,
         \Data_Mem/n7912 , \Data_Mem/n7911 , \Data_Mem/n7910 ,
         \Data_Mem/n7909 , \Data_Mem/n7908 , \Data_Mem/n7907 ,
         \Data_Mem/n7906 , \Data_Mem/n7905 , \Data_Mem/n7904 ,
         \Data_Mem/n7903 , \Data_Mem/n7902 , \Data_Mem/n7901 ,
         \Data_Mem/n7900 , \Data_Mem/n7899 , \Data_Mem/n7898 ,
         \Data_Mem/n7897 , \Data_Mem/n7896 , \Data_Mem/n7895 ,
         \Data_Mem/n7894 , \Data_Mem/n7893 , \Data_Mem/n7892 ,
         \Data_Mem/n7891 , \Data_Mem/n7890 , \Data_Mem/n7889 ,
         \Data_Mem/n7888 , \Data_Mem/n7887 , \Data_Mem/n7886 ,
         \Data_Mem/n7885 , \Data_Mem/n7884 , \Data_Mem/n7883 ,
         \Data_Mem/n7882 , \Data_Mem/n7881 , \Data_Mem/n7880 ,
         \Data_Mem/n7879 , \Data_Mem/n7878 , \Data_Mem/n7877 ,
         \Data_Mem/n7876 , \Data_Mem/n7875 , \Data_Mem/n7874 ,
         \Data_Mem/n7873 , \Data_Mem/n7872 , \Data_Mem/n7871 ,
         \Data_Mem/n7870 , \Data_Mem/n7869 , \Data_Mem/n7868 ,
         \Data_Mem/n7867 , \Data_Mem/n7866 , \Data_Mem/n7865 ,
         \Data_Mem/n7864 , \Data_Mem/n7863 , \Data_Mem/n7862 ,
         \Data_Mem/n7861 , \Data_Mem/n7860 , \Data_Mem/n7859 ,
         \Data_Mem/n7858 , \Data_Mem/n7857 , \Data_Mem/n7856 ,
         \Data_Mem/n7855 , \Data_Mem/n7854 , \Data_Mem/n7853 ,
         \Data_Mem/n7852 , \Data_Mem/n7851 , \Data_Mem/n7850 ,
         \Data_Mem/n7849 , \Data_Mem/n7848 , \Data_Mem/n7847 ,
         \Data_Mem/n7846 , \Data_Mem/n7845 , \Data_Mem/n7844 ,
         \Data_Mem/n7843 , \Data_Mem/n7842 , \Data_Mem/n7841 ,
         \Data_Mem/n7840 , \Data_Mem/n7839 , \Data_Mem/n7838 ,
         \Data_Mem/n7837 , \Data_Mem/n7836 , \Data_Mem/n7835 ,
         \Data_Mem/n7834 , \Data_Mem/n7833 , \Data_Mem/n7832 ,
         \Data_Mem/n7831 , \Data_Mem/n7830 , \Data_Mem/n7829 ,
         \Data_Mem/n7828 , \Data_Mem/n7827 , \Data_Mem/n7826 ,
         \Data_Mem/n7825 , \Data_Mem/n7824 , \Data_Mem/n7823 ,
         \Data_Mem/n7822 , \Data_Mem/n7821 , \Data_Mem/n7820 ,
         \Data_Mem/n7819 , \Data_Mem/n7818 , \Data_Mem/n7817 ,
         \Data_Mem/n7816 , \Data_Mem/n7815 , \Data_Mem/n7814 ,
         \Data_Mem/n7813 , \Data_Mem/n7812 , \Data_Mem/n7811 ,
         \Data_Mem/n7810 , \Data_Mem/n7809 , \Data_Mem/n7808 ,
         \Data_Mem/n7807 , \Data_Mem/n7806 , \Data_Mem/n7805 ,
         \Data_Mem/n7804 , \Data_Mem/n7803 , \Data_Mem/n7802 ,
         \Data_Mem/n7801 , \Data_Mem/n7800 , \Data_Mem/n7799 ,
         \Data_Mem/n7798 , \Data_Mem/n7797 , \Data_Mem/n7796 ,
         \Data_Mem/n7795 , \Data_Mem/n7794 , \Data_Mem/n7793 ,
         \Data_Mem/n7792 , \Data_Mem/n7791 , \Data_Mem/n7790 ,
         \Data_Mem/n7789 , \Data_Mem/n7788 , \Data_Mem/n7787 ,
         \Data_Mem/n7786 , \Data_Mem/n7785 , \Data_Mem/n7784 ,
         \Data_Mem/n7783 , \Data_Mem/n7782 , \Data_Mem/n7781 ,
         \Data_Mem/n7780 , \Data_Mem/n7779 , \Data_Mem/n7778 ,
         \Data_Mem/n7777 , \Data_Mem/n7776 , \Data_Mem/n7775 ,
         \Data_Mem/n7774 , \Data_Mem/n7773 , \Data_Mem/n7772 ,
         \Data_Mem/n7771 , \Data_Mem/n7770 , \Data_Mem/n7769 ,
         \Data_Mem/n7768 , \Data_Mem/n7767 , \Data_Mem/n7766 ,
         \Data_Mem/n7765 , \Data_Mem/n7764 , \Data_Mem/n7763 ,
         \Data_Mem/n7762 , \Data_Mem/n7761 , \Data_Mem/n7760 ,
         \Data_Mem/n7759 , \Data_Mem/n7758 , \Data_Mem/n7757 ,
         \Data_Mem/n7756 , \Data_Mem/n7755 , \Data_Mem/n7754 ,
         \Data_Mem/n7753 , \Data_Mem/n7752 , \Data_Mem/n7751 ,
         \Data_Mem/n7750 , \Data_Mem/n7749 , \Data_Mem/n7748 ,
         \Data_Mem/n7747 , \Data_Mem/n7746 , \Data_Mem/n7745 ,
         \Data_Mem/n7744 , \Data_Mem/n7743 , \Data_Mem/n7742 ,
         \Data_Mem/n7741 , \Data_Mem/n7740 , \Data_Mem/n7739 ,
         \Data_Mem/n7738 , \Data_Mem/n7737 , \Data_Mem/n7736 ,
         \Data_Mem/n7735 , \Data_Mem/n7734 , \Data_Mem/n7733 ,
         \Data_Mem/n7732 , \Data_Mem/n7731 , \Data_Mem/n7730 ,
         \Data_Mem/n7729 , \Data_Mem/n7728 , \Data_Mem/n7727 ,
         \Data_Mem/n7726 , \Data_Mem/n7725 , \Data_Mem/n7724 ,
         \Data_Mem/n7723 , \Data_Mem/n7722 , \Data_Mem/n7721 ,
         \Data_Mem/n7720 , \Data_Mem/n7719 , \Data_Mem/n7718 ,
         \Data_Mem/n7717 , \Data_Mem/n7716 , \Data_Mem/n7715 ,
         \Data_Mem/n7714 , \Data_Mem/n7713 , \Data_Mem/n7712 ,
         \Data_Mem/n7711 , \Data_Mem/n7710 , \Data_Mem/n7709 ,
         \Data_Mem/n7708 , \Data_Mem/n7707 , \Data_Mem/n7706 ,
         \Data_Mem/n7705 , \Data_Mem/n7704 , \Data_Mem/n7703 ,
         \Data_Mem/n7702 , \Data_Mem/n7701 , \Data_Mem/n7700 ,
         \Data_Mem/n7699 , \Data_Mem/n7698 , \Data_Mem/n7697 ,
         \Data_Mem/n7696 , \Data_Mem/n7695 , \Data_Mem/n7694 ,
         \Data_Mem/n7693 , \Data_Mem/n7692 , \Data_Mem/n7691 ,
         \Data_Mem/n7690 , \Data_Mem/n7689 , \Data_Mem/n7688 ,
         \Data_Mem/n7687 , \Data_Mem/n7686 , \Data_Mem/n7685 ,
         \Data_Mem/n7684 , \Data_Mem/n7683 , \Data_Mem/n7682 ,
         \Data_Mem/n7681 , \Data_Mem/n7680 , \Data_Mem/n7679 ,
         \Data_Mem/n7678 , \Data_Mem/n7677 , \Data_Mem/n7676 ,
         \Data_Mem/n7675 , \Data_Mem/n7674 , \Data_Mem/n7673 ,
         \Data_Mem/n7672 , \Data_Mem/n7671 , \Data_Mem/n7670 ,
         \Data_Mem/n7669 , \Data_Mem/n7668 , \Data_Mem/n7667 ,
         \Data_Mem/n7666 , \Data_Mem/n7665 , \Data_Mem/n7664 ,
         \Data_Mem/n7663 , \Data_Mem/n7662 , \Data_Mem/n7661 ,
         \Data_Mem/n7660 , \Data_Mem/n7659 , \Data_Mem/n7658 ,
         \Data_Mem/n7657 , \Data_Mem/n7656 , \Data_Mem/n7655 ,
         \Data_Mem/n7654 , \Data_Mem/n7653 , \Data_Mem/n7652 ,
         \Data_Mem/n7651 , \Data_Mem/n7650 , \Data_Mem/n7649 ,
         \Data_Mem/n7648 , \Data_Mem/n7647 , \Data_Mem/n7646 ,
         \Data_Mem/n7645 , \Data_Mem/n7644 , \Data_Mem/n7643 ,
         \Data_Mem/n7642 , \Data_Mem/n7641 , \Data_Mem/n7640 ,
         \Data_Mem/n7639 , \Data_Mem/n7638 , \Data_Mem/n7637 ,
         \Data_Mem/n7636 , \Data_Mem/n7635 , \Data_Mem/n7634 ,
         \Data_Mem/n7633 , \Data_Mem/n7632 , \Data_Mem/n7631 ,
         \Data_Mem/n7630 , \Data_Mem/n7629 , \Data_Mem/n7628 ,
         \Data_Mem/n7627 , \Data_Mem/n7626 , \Data_Mem/n7625 ,
         \Data_Mem/n7624 , \Data_Mem/n7623 , \Data_Mem/n7622 ,
         \Data_Mem/n7621 , \Data_Mem/n7620 , \Data_Mem/n7619 ,
         \Data_Mem/n7618 , \Data_Mem/n7617 , \Data_Mem/n7616 ,
         \Data_Mem/n7615 , \Data_Mem/n7614 , \Data_Mem/n7613 ,
         \Data_Mem/n7612 , \Data_Mem/n7611 , \Data_Mem/n7610 ,
         \Data_Mem/n7609 , \Data_Mem/n7608 , \Data_Mem/n7607 ,
         \Data_Mem/n7606 , \Data_Mem/n7605 , \Data_Mem/n7604 ,
         \Data_Mem/n7603 , \Data_Mem/n7602 , \Data_Mem/n7601 ,
         \Data_Mem/n7600 , \Data_Mem/n7599 , \Data_Mem/n7598 ,
         \Data_Mem/n7597 , \Data_Mem/n7596 , \Data_Mem/n7595 ,
         \Data_Mem/n7594 , \Data_Mem/n7593 , \Data_Mem/n7592 ,
         \Data_Mem/n7591 , \Data_Mem/n7590 , \Data_Mem/n7589 ,
         \Data_Mem/n7588 , \Data_Mem/n7587 , \Data_Mem/n7586 ,
         \Data_Mem/n7585 , \Data_Mem/n7584 , \Data_Mem/n7583 ,
         \Data_Mem/n7582 , \Data_Mem/n7581 , \Data_Mem/n7580 ,
         \Data_Mem/n7579 , \Data_Mem/n7578 , \Data_Mem/n7577 ,
         \Data_Mem/n7576 , \Data_Mem/n7575 , \Data_Mem/n7574 ,
         \Data_Mem/n7573 , \Data_Mem/n7572 , \Data_Mem/n7571 ,
         \Data_Mem/n7570 , \Data_Mem/n7569 , \Data_Mem/n7568 ,
         \Data_Mem/n7567 , \Data_Mem/n7566 , \Data_Mem/n7565 ,
         \Data_Mem/n7564 , \Data_Mem/n7563 , \Data_Mem/n7562 ,
         \Data_Mem/n7561 , \Data_Mem/n7560 , \Data_Mem/n7559 ,
         \Data_Mem/n7558 , \Data_Mem/n7557 , \Data_Mem/n7556 ,
         \Data_Mem/n7555 , \Data_Mem/n7554 , \Data_Mem/n7553 ,
         \Data_Mem/n7552 , \Data_Mem/n7551 , \Data_Mem/n7550 ,
         \Data_Mem/n7549 , \Data_Mem/n7548 , \Data_Mem/n7547 ,
         \Data_Mem/n7546 , \Data_Mem/n7545 , \Data_Mem/n7544 ,
         \Data_Mem/n7543 , \Data_Mem/n7542 , \Data_Mem/n7541 ,
         \Data_Mem/n7540 , \Data_Mem/n7539 , \Data_Mem/n7538 ,
         \Data_Mem/n7537 , \Data_Mem/n7536 , \Data_Mem/n7535 ,
         \Data_Mem/n7534 , \Data_Mem/n7533 , \Data_Mem/n7532 ,
         \Data_Mem/n7531 , \Data_Mem/n7530 , \Data_Mem/n7529 ,
         \Data_Mem/n7528 , \Data_Mem/n7527 , \Data_Mem/n7526 ,
         \Data_Mem/n7525 , \Data_Mem/n7524 , \Data_Mem/n7523 ,
         \Data_Mem/n7522 , \Data_Mem/n7521 , \Data_Mem/n7520 ,
         \Data_Mem/n7519 , \Data_Mem/n7518 , \Data_Mem/n7517 ,
         \Data_Mem/n7516 , \Data_Mem/n7515 , \Data_Mem/n7514 ,
         \Data_Mem/n7513 , \Data_Mem/n7512 , \Data_Mem/n7511 ,
         \Data_Mem/n7510 , \Data_Mem/n7509 , \Data_Mem/n7508 ,
         \Data_Mem/n7507 , \Data_Mem/n7506 , \Data_Mem/n7505 ,
         \Data_Mem/n7504 , \Data_Mem/n7503 , \Data_Mem/n7502 ,
         \Data_Mem/n7501 , \Data_Mem/n7500 , \Data_Mem/n7499 ,
         \Data_Mem/n7498 , \Data_Mem/n7497 , \Data_Mem/n7496 ,
         \Data_Mem/n7495 , \Data_Mem/n7494 , \Data_Mem/n7493 ,
         \Data_Mem/n7492 , \Data_Mem/n7491 , \Data_Mem/n7490 ,
         \Data_Mem/n7489 , \Data_Mem/n7488 , \Data_Mem/n7487 ,
         \Data_Mem/n7486 , \Data_Mem/n7485 , \Data_Mem/n7484 ,
         \Data_Mem/n7483 , \Data_Mem/n7482 , \Data_Mem/n7481 ,
         \Data_Mem/n7480 , \Data_Mem/n7479 , \Data_Mem/n7478 ,
         \Data_Mem/n7477 , \Data_Mem/n7476 , \Data_Mem/n7475 ,
         \Data_Mem/n7474 , \Data_Mem/n7473 , \Data_Mem/n7472 ,
         \Data_Mem/n7471 , \Data_Mem/n7470 , \Data_Mem/n7469 ,
         \Data_Mem/n7468 , \Data_Mem/n7467 , \Data_Mem/n7466 ,
         \Data_Mem/n7465 , \Data_Mem/n7464 , \Data_Mem/n7463 ,
         \Data_Mem/n7462 , \Data_Mem/n7461 , \Data_Mem/n7460 ,
         \Data_Mem/n7459 , \Data_Mem/n7458 , \Data_Mem/n7457 ,
         \Data_Mem/n7456 , \Data_Mem/n7455 , \Data_Mem/n7454 ,
         \Data_Mem/n7453 , \Data_Mem/n7452 , \Data_Mem/n7451 ,
         \Data_Mem/n7450 , \Data_Mem/n7449 , \Data_Mem/n7448 ,
         \Data_Mem/n7447 , \Data_Mem/n7446 , \Data_Mem/n7445 ,
         \Data_Mem/n7444 , \Data_Mem/n7443 , \Data_Mem/n7442 ,
         \Data_Mem/n7441 , \Data_Mem/n7440 , \Data_Mem/n7439 ,
         \Data_Mem/n7438 , \Data_Mem/n7437 , \Data_Mem/n7436 ,
         \Data_Mem/n7435 , \Data_Mem/n7434 , \Data_Mem/n7433 ,
         \Data_Mem/n7432 , \Data_Mem/n7431 , \Data_Mem/n7430 ,
         \Data_Mem/n7429 , \Data_Mem/n7428 , \Data_Mem/n7427 ,
         \Data_Mem/n7426 , \Data_Mem/n7425 , \Data_Mem/n7424 ,
         \Data_Mem/n7423 , \Data_Mem/n7422 , \Data_Mem/n7421 ,
         \Data_Mem/n7420 , \Data_Mem/n7419 , \Data_Mem/n7418 ,
         \Data_Mem/n7417 , \Data_Mem/n7416 , \Data_Mem/n7415 ,
         \Data_Mem/n7414 , \Data_Mem/n7413 , \Data_Mem/n7412 ,
         \Data_Mem/n7411 , \Data_Mem/n7410 , \Data_Mem/n7409 ,
         \Data_Mem/n7408 , \Data_Mem/n7407 , \Data_Mem/n7406 ,
         \Data_Mem/n7405 , \Data_Mem/n7404 , \Data_Mem/n7403 ,
         \Data_Mem/n7402 , \Data_Mem/n7401 , \Data_Mem/n7400 ,
         \Data_Mem/n7399 , \Data_Mem/n7398 , \Data_Mem/n7397 ,
         \Data_Mem/n7396 , \Data_Mem/n7395 , \Data_Mem/n7394 ,
         \Data_Mem/n7393 , \Data_Mem/n7392 , \Data_Mem/n7391 ,
         \Data_Mem/n7390 , \Data_Mem/n7389 , \Data_Mem/n7388 ,
         \Data_Mem/n7387 , \Data_Mem/n7386 , \Data_Mem/n7385 ,
         \Data_Mem/n7384 , \Data_Mem/n7383 , \Data_Mem/n7382 ,
         \Data_Mem/n7381 , \Data_Mem/n7380 , \Data_Mem/n7379 ,
         \Data_Mem/n7378 , \Data_Mem/n7377 , \Data_Mem/n7376 ,
         \Data_Mem/n7375 , \Data_Mem/n7374 , \Data_Mem/n7373 ,
         \Data_Mem/n7372 , \Data_Mem/n7371 , \Data_Mem/n7370 ,
         \Data_Mem/n7369 , \Data_Mem/n7368 , \Data_Mem/n7367 ,
         \Data_Mem/n7366 , \Data_Mem/n7365 , \Data_Mem/n7364 ,
         \Data_Mem/n7363 , \Data_Mem/n7362 , \Data_Mem/n7361 ,
         \Data_Mem/n7360 , \Data_Mem/n7359 , \Data_Mem/n7358 ,
         \Data_Mem/n7357 , \Data_Mem/n7356 , \Data_Mem/n7355 ,
         \Data_Mem/n7354 , \Data_Mem/n7353 , \Data_Mem/n7352 ,
         \Data_Mem/n7351 , \Data_Mem/n7350 , \Data_Mem/n7349 ,
         \Data_Mem/n7348 , \Data_Mem/n7347 , \Data_Mem/n7346 ,
         \Data_Mem/n7345 , \Data_Mem/n7344 , \Data_Mem/n7343 ,
         \Data_Mem/n7342 , \Data_Mem/n7341 , \Data_Mem/n7340 ,
         \Data_Mem/n7339 , \Data_Mem/n7338 , \Data_Mem/n7337 ,
         \Data_Mem/n7336 , \Data_Mem/n7335 , \Data_Mem/n7334 ,
         \Data_Mem/n7333 , \Data_Mem/n7332 , \Data_Mem/n7331 ,
         \Data_Mem/n7330 , \Data_Mem/n7329 , \Data_Mem/n7328 ,
         \Data_Mem/n7327 , \Data_Mem/n7326 , \Data_Mem/n7325 ,
         \Data_Mem/n7324 , \Data_Mem/n7323 , \Data_Mem/n7322 ,
         \Data_Mem/n7321 , \Data_Mem/n7320 , \Data_Mem/n7319 ,
         \Data_Mem/n7318 , \Data_Mem/n7317 , \Data_Mem/n7316 ,
         \Data_Mem/n7315 , \Data_Mem/n7314 , \Data_Mem/n7313 ,
         \Data_Mem/n7312 , \Data_Mem/n7311 , \Data_Mem/n7310 ,
         \Data_Mem/n7309 , \Data_Mem/n7308 , \Data_Mem/n7307 ,
         \Data_Mem/n7306 , \Data_Mem/n7305 , \Data_Mem/n7304 ,
         \Data_Mem/n7303 , \Data_Mem/n7302 , \Data_Mem/n7301 ,
         \Data_Mem/n7300 , \Data_Mem/n7299 , \Data_Mem/n7298 ,
         \Data_Mem/n7297 , \Data_Mem/n7296 , \Data_Mem/n7295 ,
         \Data_Mem/n7294 , \Data_Mem/n7293 , \Data_Mem/n7292 ,
         \Data_Mem/n7291 , \Data_Mem/n7290 , \Data_Mem/n7289 ,
         \Data_Mem/n7288 , \Data_Mem/n7287 , \Data_Mem/n7286 ,
         \Data_Mem/n7285 , \Data_Mem/n7284 , \Data_Mem/n7283 ,
         \Data_Mem/n7282 , \Data_Mem/n7281 , \Data_Mem/n7280 ,
         \Data_Mem/n7279 , \Data_Mem/n7278 , \Data_Mem/n7277 ,
         \Data_Mem/n7276 , \Data_Mem/n7275 , \Data_Mem/n7274 ,
         \Data_Mem/n7273 , \Data_Mem/n7272 , \Data_Mem/n7271 ,
         \Data_Mem/n7270 , \Data_Mem/n7269 , \Data_Mem/n7268 ,
         \Data_Mem/n7267 , \Data_Mem/n7266 , \Data_Mem/n7265 ,
         \Data_Mem/n7264 , \Data_Mem/n7263 , \Data_Mem/n7262 ,
         \Data_Mem/n7261 , \Data_Mem/n7260 , \Data_Mem/n7259 ,
         \Data_Mem/n7258 , \Data_Mem/n7257 , \Data_Mem/n7256 ,
         \Data_Mem/n7255 , \Data_Mem/n7254 , \Data_Mem/n7253 ,
         \Data_Mem/n7252 , \Data_Mem/n7251 , \Data_Mem/n7250 ,
         \Data_Mem/n7249 , \Data_Mem/n7248 , \Data_Mem/n7247 ,
         \Data_Mem/n7246 , \Data_Mem/n7245 , \Data_Mem/n7244 ,
         \Data_Mem/n7243 , \Data_Mem/n7242 , \Data_Mem/n7241 ,
         \Data_Mem/n7240 , \Data_Mem/n7239 , \Data_Mem/n7238 ,
         \Data_Mem/n7237 , \Data_Mem/n7236 , \Data_Mem/n7235 ,
         \Data_Mem/n7234 , \Data_Mem/n7233 , \Data_Mem/n7232 ,
         \Data_Mem/n7231 , \Data_Mem/n7230 , \Data_Mem/n7229 ,
         \Data_Mem/n7228 , \Data_Mem/n7227 , \Data_Mem/n7226 ,
         \Data_Mem/n7225 , \Data_Mem/n7224 , \Data_Mem/n7223 ,
         \Data_Mem/n7222 , \Data_Mem/n7221 , \Data_Mem/n7220 ,
         \Data_Mem/n7219 , \Data_Mem/n7218 , \Data_Mem/n7217 ,
         \Data_Mem/n7216 , \Data_Mem/n7215 , \Data_Mem/n7214 ,
         \Data_Mem/n7213 , \Data_Mem/n7212 , \Data_Mem/n7211 ,
         \Data_Mem/n7210 , \Data_Mem/n7209 , \Data_Mem/n7208 ,
         \Data_Mem/n7207 , \Data_Mem/n7206 , \Data_Mem/n7205 ,
         \Data_Mem/n7204 , \Data_Mem/n7203 , \Data_Mem/n7202 ,
         \Data_Mem/n7201 , \Data_Mem/n7200 , \Data_Mem/n7199 ,
         \Data_Mem/n7198 , \Data_Mem/n7197 , \Data_Mem/n7196 ,
         \Data_Mem/n7195 , \Data_Mem/n7194 , \Data_Mem/n7193 ,
         \Data_Mem/n7192 , \Data_Mem/n7191 , \Data_Mem/n7190 ,
         \Data_Mem/n7189 , \Data_Mem/n7188 , \Data_Mem/n7187 ,
         \Data_Mem/n7186 , \Data_Mem/n7185 , \Data_Mem/n7184 ,
         \Data_Mem/n7183 , \Data_Mem/n7182 , \Data_Mem/n7181 ,
         \Data_Mem/n7180 , \Data_Mem/n7179 , \Data_Mem/n7178 ,
         \Data_Mem/n7177 , \Data_Mem/n7176 , \Data_Mem/n7175 ,
         \Data_Mem/n7174 , \Data_Mem/n7173 , \Data_Mem/n7172 ,
         \Data_Mem/n7171 , \Data_Mem/n7170 , \Data_Mem/n7169 ,
         \Data_Mem/n7168 , \Data_Mem/n7167 , \Data_Mem/n7166 ,
         \Data_Mem/n7165 , \Data_Mem/n7164 , \Data_Mem/n7163 ,
         \Data_Mem/n7162 , \Data_Mem/n7161 , \Data_Mem/n7160 ,
         \Data_Mem/n7159 , \Data_Mem/n7158 , \Data_Mem/n7157 ,
         \Data_Mem/n7156 , \Data_Mem/n7155 , \Data_Mem/n7154 ,
         \Data_Mem/n7153 , \Data_Mem/n7152 , \Data_Mem/n7151 ,
         \Data_Mem/n7150 , \Data_Mem/n7149 , \Data_Mem/n7148 ,
         \Data_Mem/n7147 , \Data_Mem/n7146 , \Data_Mem/n7145 ,
         \Data_Mem/n7144 , \Data_Mem/n7143 , \Data_Mem/n7142 ,
         \Data_Mem/n7141 , \Data_Mem/n7140 , \Data_Mem/n7139 ,
         \Data_Mem/n7138 , \Data_Mem/n7137 , \Data_Mem/n7136 ,
         \Data_Mem/n7135 , \Data_Mem/n7134 , \Data_Mem/n7133 ,
         \Data_Mem/n7132 , \Data_Mem/n7131 , \Data_Mem/n7130 ,
         \Data_Mem/n7129 , \Data_Mem/n7128 , \Data_Mem/n7127 ,
         \Data_Mem/n7126 , \Data_Mem/n7125 , \Data_Mem/n7124 ,
         \Data_Mem/n7123 , \Data_Mem/n7122 , \Data_Mem/n7121 ,
         \Data_Mem/n7120 , \Data_Mem/n7119 , \Data_Mem/n7118 ,
         \Data_Mem/n7117 , \Data_Mem/n7116 , \Data_Mem/n7115 ,
         \Data_Mem/n7114 , \Data_Mem/n7113 , \Data_Mem/n7112 ,
         \Data_Mem/n7111 , \Data_Mem/n7110 , \Data_Mem/n7109 ,
         \Data_Mem/n7108 , \Data_Mem/n7107 , \Data_Mem/n7106 ,
         \Data_Mem/n7105 , \Data_Mem/n7104 , \Data_Mem/n7103 ,
         \Data_Mem/n7102 , \Data_Mem/n7101 , \Data_Mem/n7100 ,
         \Data_Mem/n7099 , \Data_Mem/n7098 , \Data_Mem/n7097 ,
         \Data_Mem/n7096 , \Data_Mem/n7095 , \Data_Mem/n7094 ,
         \Data_Mem/n7093 , \Data_Mem/n7092 , \Data_Mem/n7091 ,
         \Data_Mem/n7090 , \Data_Mem/n7089 , \Data_Mem/n7088 ,
         \Data_Mem/n7087 , \Data_Mem/n7086 , \Data_Mem/n7085 ,
         \Data_Mem/n7084 , \Data_Mem/n7083 , \Data_Mem/n7082 ,
         \Data_Mem/n7081 , \Data_Mem/n7080 , \Data_Mem/n7079 ,
         \Data_Mem/n7078 , \Data_Mem/n7077 , \Data_Mem/n7076 ,
         \Data_Mem/n7075 , \Data_Mem/n7074 , \Data_Mem/n7073 ,
         \Data_Mem/n7072 , \Data_Mem/n7071 , \Data_Mem/n7070 ,
         \Data_Mem/n7069 , \Data_Mem/n7068 , \Data_Mem/n7067 ,
         \Data_Mem/n7066 , \Data_Mem/n7065 , \Data_Mem/n7064 ,
         \Data_Mem/n7063 , \Data_Mem/n7062 , \Data_Mem/n7061 ,
         \Data_Mem/n7060 , \Data_Mem/n7059 , \Data_Mem/n7058 ,
         \Data_Mem/n7057 , \Data_Mem/n7056 , \Data_Mem/n7055 ,
         \Data_Mem/n7054 , \Data_Mem/n7053 , \Data_Mem/n7052 ,
         \Data_Mem/n7051 , \Data_Mem/n7050 , \Data_Mem/n7049 ,
         \Data_Mem/n7048 , \Data_Mem/n7047 , \Data_Mem/n7046 ,
         \Data_Mem/n7045 , \Data_Mem/n7044 , \Data_Mem/n7043 ,
         \Data_Mem/n7042 , \Data_Mem/n7041 , \Data_Mem/n7040 ,
         \Data_Mem/n7039 , \Data_Mem/n7038 , \Data_Mem/n7037 ,
         \Data_Mem/n7036 , \Data_Mem/n7035 , \Data_Mem/n7034 ,
         \Data_Mem/n7033 , \Data_Mem/n7032 , \Data_Mem/n7031 ,
         \Data_Mem/n7030 , \Data_Mem/n7029 , \Data_Mem/n7028 ,
         \Data_Mem/n7027 , \Data_Mem/n7026 , \Data_Mem/n7025 ,
         \Data_Mem/n7024 , \Data_Mem/n7023 , \Data_Mem/n7022 ,
         \Data_Mem/n7021 , \Data_Mem/n7020 , \Data_Mem/n7019 ,
         \Data_Mem/n7018 , \Data_Mem/n7017 , \Data_Mem/n7016 ,
         \Data_Mem/n7015 , \Data_Mem/n7014 , \Data_Mem/n7013 ,
         \Data_Mem/n7012 , \Data_Mem/n7011 , \Data_Mem/n7010 ,
         \Data_Mem/n7009 , \Data_Mem/n7008 , \Data_Mem/n7007 ,
         \Data_Mem/n7006 , \Data_Mem/n7005 , \Data_Mem/n7004 ,
         \Data_Mem/n7003 , \Data_Mem/n7002 , \Data_Mem/n7001 ,
         \Data_Mem/n7000 , \Data_Mem/n6999 , \Data_Mem/n6998 ,
         \Data_Mem/n6997 , \Data_Mem/n6996 , \Data_Mem/n6995 ,
         \Data_Mem/n6994 , \Data_Mem/n6993 , \Data_Mem/n6992 ,
         \Data_Mem/n6991 , \Data_Mem/n6990 , \Data_Mem/n6989 ,
         \Data_Mem/n6988 , \Data_Mem/n6987 , \Data_Mem/n6986 ,
         \Data_Mem/n6985 , \Data_Mem/n6984 , \Data_Mem/n6983 ,
         \Data_Mem/n6982 , \Data_Mem/n6981 , \Data_Mem/n6980 ,
         \Data_Mem/n6979 , \Data_Mem/n6978 , \Data_Mem/n6977 ,
         \Data_Mem/n6976 , \Data_Mem/n6975 , \Data_Mem/n6974 ,
         \Data_Mem/n6973 , \Data_Mem/n6972 , \Data_Mem/n6971 ,
         \Data_Mem/n6970 , \Data_Mem/n6969 , \Data_Mem/n6968 ,
         \Data_Mem/n6967 , \Data_Mem/n6966 , \Data_Mem/n6965 ,
         \Data_Mem/n6964 , \Data_Mem/n6963 , \Data_Mem/n6962 ,
         \Data_Mem/n6961 , \Data_Mem/n6960 , \Data_Mem/n6959 ,
         \Data_Mem/n6958 , \Data_Mem/n6957 , \Data_Mem/n6956 ,
         \Data_Mem/n6955 , \Data_Mem/n6954 , \Data_Mem/n6953 ,
         \Data_Mem/n6952 , \Data_Mem/n6951 , \Data_Mem/n6950 ,
         \Data_Mem/n6949 , \Data_Mem/n6948 , \Data_Mem/n6947 ,
         \Data_Mem/n6946 , \Data_Mem/n6945 , \Data_Mem/n6944 ,
         \Data_Mem/n6943 , \Data_Mem/n6942 , \Data_Mem/n6941 ,
         \Data_Mem/n6940 , \Data_Mem/n6939 , \Data_Mem/n6938 ,
         \Data_Mem/n6937 , \Data_Mem/n6936 , \Data_Mem/n6935 ,
         \Data_Mem/n6934 , \Data_Mem/n6933 , \Data_Mem/n6932 ,
         \Data_Mem/n6931 , \Data_Mem/n6930 , \Data_Mem/n6929 ,
         \Data_Mem/n6928 , \Data_Mem/n6927 , \Data_Mem/n6926 ,
         \Data_Mem/n6925 , \Data_Mem/n6924 , \Data_Mem/n6923 ,
         \Data_Mem/n6922 , \Data_Mem/n6921 , \Data_Mem/n6920 ,
         \Data_Mem/n6919 , \Data_Mem/n6918 , \Data_Mem/n6917 ,
         \Data_Mem/n6916 , \Data_Mem/n6915 , \Data_Mem/n6914 ,
         \Data_Mem/n6913 , \Data_Mem/n6912 , \Data_Mem/n6911 ,
         \Data_Mem/n6910 , \Data_Mem/n6909 , \Data_Mem/n6908 ,
         \Data_Mem/n6907 , \Data_Mem/n6906 , \Data_Mem/n6905 ,
         \Data_Mem/n6904 , \Data_Mem/n6903 , \Data_Mem/n6902 ,
         \Data_Mem/n6901 , \Data_Mem/n6900 , \Data_Mem/n6899 ,
         \Data_Mem/n6898 , \Data_Mem/n6897 , \Data_Mem/n6896 ,
         \Data_Mem/n6895 , \Data_Mem/n6894 , \Data_Mem/n6893 ,
         \Data_Mem/n6892 , \Data_Mem/n6891 , \Data_Mem/n6890 ,
         \Data_Mem/n6889 , \Data_Mem/n6888 , \Data_Mem/n6887 ,
         \Data_Mem/n6886 , \Data_Mem/n6885 , \Data_Mem/n6884 ,
         \Data_Mem/n6883 , \Data_Mem/n6882 , \Data_Mem/n6881 ,
         \Data_Mem/n6880 , \Data_Mem/n6879 , \Data_Mem/n6878 ,
         \Data_Mem/n6877 , \Data_Mem/n6876 , \Data_Mem/n6875 ,
         \Data_Mem/n6874 , \Data_Mem/n6873 , \Data_Mem/n6872 ,
         \Data_Mem/n6871 , \Data_Mem/n6870 , \Data_Mem/n6869 ,
         \Data_Mem/n6868 , \Data_Mem/n6867 , \Data_Mem/n6866 ,
         \Data_Mem/n6865 , \Data_Mem/n6864 , \Data_Mem/n6863 ,
         \Data_Mem/n6862 , \Data_Mem/n6861 , \Data_Mem/n6860 ,
         \Data_Mem/n6859 , \Data_Mem/n6858 , \Data_Mem/n6857 ,
         \Data_Mem/n6856 , \Data_Mem/n6855 , \Data_Mem/n6854 ,
         \Data_Mem/n6853 , \Data_Mem/n6852 , \Data_Mem/n6851 ,
         \Data_Mem/n6850 , \Data_Mem/n6849 , \Data_Mem/n6848 ,
         \Data_Mem/n6847 , \Data_Mem/n6846 , \Data_Mem/n6845 ,
         \Data_Mem/n6844 , \Data_Mem/n6843 , \Data_Mem/n6842 ,
         \Data_Mem/n6841 , \Data_Mem/n6840 , \Data_Mem/n6839 ,
         \Data_Mem/n6838 , \Data_Mem/n6837 , \Data_Mem/n6836 ,
         \Data_Mem/n6835 , \Data_Mem/n6834 , \Data_Mem/n6833 ,
         \Data_Mem/n6832 , \Data_Mem/n6831 , \Data_Mem/n6830 ,
         \Data_Mem/n6829 , \Data_Mem/n6828 , \Data_Mem/n6827 ,
         \Data_Mem/n6826 , \Data_Mem/n6825 , \Data_Mem/n6824 ,
         \Data_Mem/n6823 , \Data_Mem/n6822 , \Data_Mem/n6821 ,
         \Data_Mem/n6820 , \Data_Mem/n6819 , \Data_Mem/n6818 ,
         \Data_Mem/n6817 , \Data_Mem/n6816 , \Data_Mem/n6815 ,
         \Data_Mem/n6814 , \Data_Mem/n6813 , \Data_Mem/n6812 ,
         \Data_Mem/n6811 , \Data_Mem/n6810 , \Data_Mem/n6809 ,
         \Data_Mem/n6808 , \Data_Mem/n6807 , \Data_Mem/n6806 ,
         \Data_Mem/n6805 , \Data_Mem/n6804 , \Data_Mem/n6803 ,
         \Data_Mem/n6802 , \Data_Mem/n6801 , \Data_Mem/n6800 ,
         \Data_Mem/n6799 , \Data_Mem/n6798 , \Data_Mem/n6797 ,
         \Data_Mem/n6796 , \Data_Mem/n6795 , \Data_Mem/n6794 ,
         \Data_Mem/n6793 , \Data_Mem/n6792 , \Data_Mem/n6791 ,
         \Data_Mem/n6790 , \Data_Mem/n6789 , \Data_Mem/n6788 ,
         \Data_Mem/n6787 , \Data_Mem/n6786 , \Data_Mem/n6785 ,
         \Data_Mem/n6784 , \Data_Mem/n6783 , \Data_Mem/n6782 ,
         \Data_Mem/n6781 , \Data_Mem/n6780 , \Data_Mem/n6779 ,
         \Data_Mem/n6778 , \Data_Mem/n6777 , \Data_Mem/n6776 ,
         \Data_Mem/n6775 , \Data_Mem/n6774 , \Data_Mem/n6773 ,
         \Data_Mem/n6772 , \Data_Mem/n6771 , \Data_Mem/n6770 ,
         \Data_Mem/n6769 , \Data_Mem/n6768 , \Data_Mem/n6767 ,
         \Data_Mem/n6766 , \Data_Mem/n6765 , \Data_Mem/n6764 ,
         \Data_Mem/n6763 , \Data_Mem/n6762 , \Data_Mem/n6761 ,
         \Data_Mem/n6760 , \Data_Mem/n6759 , \Data_Mem/n6758 ,
         \Data_Mem/n6757 , \Data_Mem/n6756 , \Data_Mem/n6755 ,
         \Data_Mem/n6754 , \Data_Mem/n6753 , \Data_Mem/n6752 ,
         \Data_Mem/n6751 , \Data_Mem/n6750 , \Data_Mem/n6749 ,
         \Data_Mem/n6748 , \Data_Mem/n6747 , \Data_Mem/n6746 ,
         \Data_Mem/n6745 , \Data_Mem/n6744 , \Data_Mem/n6743 ,
         \Data_Mem/n6742 , \Data_Mem/n6741 , \Data_Mem/n6740 ,
         \Data_Mem/n6739 , \Data_Mem/n6738 , \Data_Mem/n6737 ,
         \Data_Mem/n6736 , \Data_Mem/n6735 , \Data_Mem/n6734 ,
         \Data_Mem/n6733 , \Data_Mem/n6732 , \Data_Mem/n6731 ,
         \Data_Mem/n6730 , \Data_Mem/n6729 , \Data_Mem/n6728 ,
         \Data_Mem/n6727 , \Data_Mem/n6726 , \Data_Mem/n6725 ,
         \Data_Mem/n6724 , \Data_Mem/n6723 , \Data_Mem/n6722 ,
         \Data_Mem/n6721 , \Data_Mem/n6720 , \Data_Mem/n6719 ,
         \Data_Mem/n6718 , \Data_Mem/n6717 , \Data_Mem/n6716 ,
         \Data_Mem/n6715 , \Data_Mem/n6714 , \Data_Mem/n6713 ,
         \Data_Mem/n6712 , \Data_Mem/n6711 , \Data_Mem/n6710 ,
         \Data_Mem/n6709 , \Data_Mem/n6708 , \Data_Mem/n6707 ,
         \Data_Mem/n6706 , \Data_Mem/n6705 , \Data_Mem/n6704 ,
         \Data_Mem/n6703 , \Data_Mem/n6702 , \Data_Mem/n6701 ,
         \Data_Mem/n6700 , \Data_Mem/n6699 , \Data_Mem/n6698 ,
         \Data_Mem/n6697 , \Data_Mem/n6696 , \Data_Mem/n6695 ,
         \Data_Mem/n6694 , \Data_Mem/n6693 , \Data_Mem/n6692 ,
         \Data_Mem/n6691 , \Data_Mem/n6690 , \Data_Mem/n6689 ,
         \Data_Mem/n6688 , \Data_Mem/n6687 , \Data_Mem/n6686 ,
         \Data_Mem/n6685 , \Data_Mem/n6684 , \Data_Mem/n6683 ,
         \Data_Mem/n6682 , \Data_Mem/n6681 , \Data_Mem/n6680 ,
         \Data_Mem/n6679 , \Data_Mem/n6678 , \Data_Mem/n6677 ,
         \Data_Mem/n6676 , \Data_Mem/n6675 , \Data_Mem/n6674 ,
         \Data_Mem/n6673 , \Data_Mem/n6672 , \Data_Mem/n6671 ,
         \Data_Mem/n6670 , \Data_Mem/n6669 , \Data_Mem/n6668 ,
         \Data_Mem/n6667 , \Data_Mem/n6666 , \Data_Mem/n6665 ,
         \Data_Mem/n6664 , \Data_Mem/n6663 , \Data_Mem/n6662 ,
         \Data_Mem/n6661 , \Data_Mem/n6660 , \Data_Mem/n6659 ,
         \Data_Mem/n6658 , \Data_Mem/n6657 , \Data_Mem/n6656 ,
         \Data_Mem/n6655 , \Data_Mem/n6654 , \Data_Mem/n6653 ,
         \Data_Mem/n6652 , \Data_Mem/n6651 , \Data_Mem/n6650 ,
         \Data_Mem/n6649 , \Data_Mem/n6648 , \Data_Mem/n6647 ,
         \Data_Mem/n6646 , \Data_Mem/n6645 , \Data_Mem/n6644 ,
         \Data_Mem/n6643 , \Data_Mem/n6642 , \Data_Mem/n6641 ,
         \Data_Mem/n6640 , \Data_Mem/n6639 , \Data_Mem/n6638 ,
         \Data_Mem/n6637 , \Data_Mem/n6636 , \Data_Mem/n6635 ,
         \Data_Mem/n6634 , \Data_Mem/n6633 , \Data_Mem/n6632 ,
         \Data_Mem/n6631 , \Data_Mem/n6630 , \Data_Mem/n6629 ,
         \Data_Mem/n6628 , \Data_Mem/n6627 , \Data_Mem/n6626 ,
         \Data_Mem/n6625 , \Data_Mem/n6624 , \Data_Mem/n6623 ,
         \Data_Mem/n6622 , \Data_Mem/n6621 , \Data_Mem/n6620 ,
         \Data_Mem/n6619 , \Data_Mem/n6618 , \Data_Mem/n6617 ,
         \Data_Mem/n6616 , \Data_Mem/n6615 , \Data_Mem/n6614 ,
         \Data_Mem/n6613 , \Data_Mem/n6612 , \Data_Mem/n6611 ,
         \Data_Mem/n6610 , \Data_Mem/n6609 , \Data_Mem/n6608 ,
         \Data_Mem/n6607 , \Data_Mem/n6606 , \Data_Mem/n6605 ,
         \Data_Mem/n6604 , \Data_Mem/n6603 , \Data_Mem/n6602 ,
         \Data_Mem/n6601 , \Data_Mem/n6600 , \Data_Mem/n6599 ,
         \Data_Mem/n6598 , \Data_Mem/n6597 , \Data_Mem/n6596 ,
         \Data_Mem/n6595 , \Data_Mem/n6594 , \Data_Mem/n6593 ,
         \Data_Mem/n6592 , \Data_Mem/n6591 , \Data_Mem/n6590 ,
         \Data_Mem/n6589 , \Data_Mem/n6588 , \Data_Mem/n6587 ,
         \Data_Mem/n6586 , \Data_Mem/n6585 , \Data_Mem/n6584 ,
         \Data_Mem/n6583 , \Data_Mem/n6582 , \Data_Mem/n6581 ,
         \Data_Mem/n6580 , \Data_Mem/n6579 , \Data_Mem/n6578 ,
         \Data_Mem/n6577 , \Data_Mem/n6576 , \Data_Mem/n6575 ,
         \Data_Mem/n6574 , \Data_Mem/n6573 , \Data_Mem/n6572 ,
         \Data_Mem/n6571 , \Data_Mem/n6570 , \Data_Mem/n6569 ,
         \Data_Mem/n6568 , \Data_Mem/n6567 , \Data_Mem/n6566 ,
         \Data_Mem/n6565 , \Data_Mem/n6564 , \Data_Mem/n6563 ,
         \Data_Mem/n6562 , \Data_Mem/n6561 , \Data_Mem/n6560 ,
         \Data_Mem/n6559 , \Data_Mem/n6558 , \Data_Mem/n6557 ,
         \Data_Mem/n6556 , \Data_Mem/n6555 , \Data_Mem/n6554 ,
         \Data_Mem/n6553 , \Data_Mem/n6552 , \Data_Mem/n6551 ,
         \Data_Mem/n6550 , \Data_Mem/n6549 , \Data_Mem/n6548 ,
         \Data_Mem/n6547 , \Data_Mem/n6546 , \Data_Mem/n6545 ,
         \Data_Mem/n6544 , \Data_Mem/n6543 , \Data_Mem/n6542 ,
         \Data_Mem/n6541 , \Data_Mem/n6540 , \Data_Mem/n6539 ,
         \Data_Mem/n6538 , \Data_Mem/n6537 , \Data_Mem/n6536 ,
         \Data_Mem/n6535 , \Data_Mem/n6534 , \Data_Mem/n6533 ,
         \Data_Mem/n6532 , \Data_Mem/n6531 , \Data_Mem/n6530 ,
         \Data_Mem/n6529 , \Data_Mem/n6528 , \Data_Mem/n6527 ,
         \Data_Mem/n6526 , \Data_Mem/n6525 , \Data_Mem/n6524 ,
         \Data_Mem/n6523 , \Data_Mem/n6522 , \Data_Mem/n6521 ,
         \Data_Mem/n6520 , \Data_Mem/n6519 , \Data_Mem/n6518 ,
         \Data_Mem/n6517 , \Data_Mem/n6516 , \Data_Mem/n6515 ,
         \Data_Mem/n6514 , \Data_Mem/n6513 , \Data_Mem/n6512 ,
         \Data_Mem/n6511 , \Data_Mem/n6510 , \Data_Mem/n6509 ,
         \Data_Mem/n6508 , \Data_Mem/n6507 , \Data_Mem/n6506 ,
         \Data_Mem/n6505 , \Data_Mem/n6504 , \Data_Mem/n6503 ,
         \Data_Mem/n6502 , \Data_Mem/n6501 , \Data_Mem/n6500 ,
         \Data_Mem/n6499 , \Data_Mem/n6498 , \Data_Mem/n6497 ,
         \Data_Mem/n6496 , \Data_Mem/n6495 , \Data_Mem/n6494 ,
         \Data_Mem/n6493 , \Data_Mem/n6492 , \Data_Mem/n6491 ,
         \Data_Mem/n6490 , \Data_Mem/n6489 , \Data_Mem/n6488 ,
         \Data_Mem/n6487 , \Data_Mem/n6486 , \Data_Mem/n6485 ,
         \Data_Mem/n6484 , \Data_Mem/n6483 , \Data_Mem/n6482 ,
         \Data_Mem/n6481 , \Data_Mem/n6480 , \Data_Mem/n6479 ,
         \Data_Mem/n6478 , \Data_Mem/n6477 , \Data_Mem/n6476 ,
         \Data_Mem/n6475 , \Data_Mem/n6474 , \Data_Mem/n6473 ,
         \Data_Mem/n6472 , \Data_Mem/n6471 , \Data_Mem/n6470 ,
         \Data_Mem/n6469 , \Data_Mem/n6468 , \Data_Mem/n6467 ,
         \Data_Mem/n6466 , \Data_Mem/n6465 , \Data_Mem/n6464 ,
         \Data_Mem/n6463 , \Data_Mem/n6462 , \Data_Mem/n6461 ,
         \Data_Mem/n6460 , \Data_Mem/n6459 , \Data_Mem/n6458 ,
         \Data_Mem/n6457 , \Data_Mem/n6456 , \Data_Mem/n6455 ,
         \Data_Mem/n6454 , \Data_Mem/n6453 , \Data_Mem/n6452 ,
         \Data_Mem/n6451 , \Data_Mem/n6450 , \Data_Mem/n6449 ,
         \Data_Mem/n6448 , \Data_Mem/n6447 , \Data_Mem/n6446 ,
         \Data_Mem/n6445 , \Data_Mem/n6444 , \Data_Mem/n6443 ,
         \Data_Mem/n6442 , \Data_Mem/n6441 , \Data_Mem/n6440 ,
         \Data_Mem/n6439 , \Data_Mem/n6438 , \Data_Mem/n6437 ,
         \Data_Mem/n6436 , \Data_Mem/n6435 , \Data_Mem/n6434 ,
         \Data_Mem/n6433 , \Data_Mem/n6432 , \Data_Mem/n6431 ,
         \Data_Mem/n6430 , \Data_Mem/n6429 , \Data_Mem/n6428 ,
         \Data_Mem/n6427 , \Data_Mem/n6426 , \Data_Mem/n6425 ,
         \Data_Mem/n6424 , \Data_Mem/n6423 , \Data_Mem/n6422 ,
         \Data_Mem/n6421 , \Data_Mem/n6420 , \Data_Mem/n6419 ,
         \Data_Mem/n6418 , \Data_Mem/n6417 , \Data_Mem/n6416 ,
         \Data_Mem/n6415 , \Data_Mem/n6414 , \Data_Mem/n6413 ,
         \Data_Mem/n6412 , \Data_Mem/n6411 , \Data_Mem/n6410 ,
         \Data_Mem/n6409 , \Data_Mem/n6408 , \Data_Mem/n6407 ,
         \Data_Mem/n6406 , \Data_Mem/n6405 , \Data_Mem/n6404 ,
         \Data_Mem/n6403 , \Data_Mem/n6402 , \Data_Mem/n6401 ,
         \Data_Mem/n6400 , \Data_Mem/n6399 , \Data_Mem/n6398 ,
         \Data_Mem/n6397 , \Data_Mem/n6396 , \Data_Mem/n6395 ,
         \Data_Mem/n6394 , \Data_Mem/n6393 , \Data_Mem/n6392 ,
         \Data_Mem/n6391 , \Data_Mem/n6390 , \Data_Mem/n6389 ,
         \Data_Mem/n6388 , \Data_Mem/n6387 , \Data_Mem/n6386 ,
         \Data_Mem/n6385 , \Data_Mem/n6384 , \Data_Mem/n6383 ,
         \Data_Mem/n6382 , \Data_Mem/n6381 , \Data_Mem/n6380 ,
         \Data_Mem/n6379 , \Data_Mem/n6378 , \Data_Mem/n6377 ,
         \Data_Mem/n6376 , \Data_Mem/n6375 , \Data_Mem/n6374 ,
         \Data_Mem/n6373 , \Data_Mem/n6372 , \Data_Mem/n6371 ,
         \Data_Mem/n6370 , \Data_Mem/n6369 , \Data_Mem/n6368 ,
         \Data_Mem/n6367 , \Data_Mem/n6366 , \Data_Mem/n6365 ,
         \Data_Mem/n6364 , \Data_Mem/n6363 , \Data_Mem/n6362 ,
         \Data_Mem/n6361 , \Data_Mem/n6360 , \Data_Mem/n6359 ,
         \Data_Mem/n6358 , \Data_Mem/n6357 , \Data_Mem/n6356 ,
         \Data_Mem/n6355 , \Data_Mem/n6354 , \Data_Mem/n6353 ,
         \Data_Mem/n6352 , \Data_Mem/n6351 , \Data_Mem/n6350 ,
         \Data_Mem/n6349 , \Data_Mem/n6348 , \Data_Mem/n6347 ,
         \Data_Mem/n6346 , \Data_Mem/n6345 , \Data_Mem/n6344 ,
         \Data_Mem/n6343 , \Data_Mem/n6342 , \Data_Mem/n6341 ,
         \Data_Mem/n6340 , \Data_Mem/n6339 , \Data_Mem/n6338 ,
         \Data_Mem/n6337 , \Data_Mem/n6336 , \Data_Mem/n6335 ,
         \Data_Mem/n6334 , \Data_Mem/n6333 , \Data_Mem/n6332 ,
         \Data_Mem/n6331 , \Data_Mem/n6330 , \Data_Mem/n6329 ,
         \Data_Mem/n6328 , \Data_Mem/n6327 , \Data_Mem/n6326 ,
         \Data_Mem/n6325 , \Data_Mem/n6324 , \Data_Mem/n6323 ,
         \Data_Mem/n6322 , \Data_Mem/n6321 , \Data_Mem/n6320 ,
         \Data_Mem/n6319 , \Data_Mem/n6318 , \Data_Mem/n6317 ,
         \Data_Mem/n6316 , \Data_Mem/n6315 , \Data_Mem/n6314 ,
         \Data_Mem/n6313 , \Data_Mem/n6312 , \Data_Mem/n6311 ,
         \Data_Mem/n6310 , \Data_Mem/n6309 , \Data_Mem/n6308 ,
         \Data_Mem/n6307 , \Data_Mem/n6306 , \Data_Mem/n6305 ,
         \Data_Mem/n6304 , \Data_Mem/n6303 , \Data_Mem/n6302 ,
         \Data_Mem/n6301 , \Data_Mem/n6300 , \Data_Mem/n6299 ,
         \Data_Mem/n6298 , \Data_Mem/n6297 , \Data_Mem/n6296 ,
         \Data_Mem/n6295 , \Data_Mem/n6294 , \Data_Mem/n6293 ,
         \Data_Mem/n6292 , \Data_Mem/n6291 , \Data_Mem/n6290 ,
         \Data_Mem/n6289 , \Data_Mem/n6288 , \Data_Mem/n6287 ,
         \Data_Mem/n6286 , \Data_Mem/n6285 , \Data_Mem/n6284 ,
         \Data_Mem/n6283 , \Data_Mem/n6282 , \Data_Mem/n6281 ,
         \Data_Mem/n6280 , \Data_Mem/n6279 , \Data_Mem/n6278 ,
         \Data_Mem/n6277 , \Data_Mem/n6276 , \Data_Mem/n6275 ,
         \Data_Mem/n6274 , \Data_Mem/n6273 , \Data_Mem/n6272 ,
         \Data_Mem/n6271 , \Data_Mem/n6270 , \Data_Mem/n6269 ,
         \Data_Mem/n6268 , \Data_Mem/n6267 , \Data_Mem/n6266 ,
         \Data_Mem/n6265 , \Data_Mem/n6264 , \Data_Mem/n6263 ,
         \Data_Mem/n6262 , \Data_Mem/n6261 , \Data_Mem/n6260 ,
         \Data_Mem/n6259 , \Data_Mem/n6258 , \Data_Mem/n6257 ,
         \Data_Mem/n6256 , \Data_Mem/n6255 , \Data_Mem/n6254 ,
         \Data_Mem/n6253 , \Data_Mem/n6252 , \Data_Mem/n6251 ,
         \Data_Mem/n6250 , \Data_Mem/n6249 , \Data_Mem/n6248 ,
         \Data_Mem/n6247 , \Data_Mem/n6246 , \Data_Mem/n6245 ,
         \Data_Mem/n6244 , \Data_Mem/n6243 , \Data_Mem/n6242 ,
         \Data_Mem/n6241 , \Data_Mem/n6240 , \Data_Mem/n6239 ,
         \Data_Mem/n6238 , \Data_Mem/n6237 , \Data_Mem/n6236 ,
         \Data_Mem/n6235 , \Data_Mem/n6234 , \Data_Mem/n6233 ,
         \Data_Mem/n6232 , \Data_Mem/n6231 , \Data_Mem/n6230 ,
         \Data_Mem/n6229 , \Data_Mem/n6228 , \Data_Mem/n6227 ,
         \Data_Mem/n6226 , \Data_Mem/n6225 , \Data_Mem/n6224 ,
         \Data_Mem/n6223 , \Data_Mem/n6222 , \Data_Mem/n6221 ,
         \Data_Mem/n6220 , \Data_Mem/n6219 , \Data_Mem/n6218 ,
         \Data_Mem/n6217 , \Data_Mem/n6216 , \Data_Mem/n6215 ,
         \Data_Mem/n6214 , \Data_Mem/n6213 , \Data_Mem/n6212 ,
         \Data_Mem/n6211 , \Data_Mem/n6210 , \Data_Mem/n6209 ,
         \Data_Mem/n6208 , \Data_Mem/n6207 , \Data_Mem/n6206 ,
         \Data_Mem/n6205 , \Data_Mem/n6204 , \Data_Mem/n6203 ,
         \Data_Mem/n6202 , \Data_Mem/n6201 , \Data_Mem/n6200 ,
         \Data_Mem/n6199 , \Data_Mem/n6198 , \Data_Mem/n6197 ,
         \Data_Mem/n6196 , \Data_Mem/n6195 , \Data_Mem/n6194 ,
         \Data_Mem/n6193 , \Data_Mem/n6192 , \Data_Mem/n6191 ,
         \Data_Mem/n6190 , \Data_Mem/n6189 , \Data_Mem/n6188 ,
         \Data_Mem/n6187 , \Data_Mem/n6186 , \Data_Mem/n6185 ,
         \Data_Mem/n6184 , \Data_Mem/n6183 , \Data_Mem/n6182 ,
         \Data_Mem/n6181 , \Data_Mem/n6180 , \Data_Mem/n6179 ,
         \Data_Mem/n6178 , \Data_Mem/n6177 , \Data_Mem/n6176 ,
         \Data_Mem/n6175 , \Data_Mem/n6174 , \Data_Mem/n6173 ,
         \Data_Mem/n6172 , \Data_Mem/n6171 , \Data_Mem/n6170 ,
         \Data_Mem/n6169 , \Data_Mem/n6168 , \Data_Mem/n6167 ,
         \Data_Mem/n6166 , \Data_Mem/n6165 , \Data_Mem/n6164 ,
         \Data_Mem/n6163 , \Data_Mem/n6162 , \Data_Mem/n6161 ,
         \Data_Mem/n6160 , \Data_Mem/n6159 , \Data_Mem/n6158 ,
         \Data_Mem/n6157 , \Data_Mem/n6156 , \Data_Mem/n6155 ,
         \Data_Mem/n6154 , \Data_Mem/n6153 , \Data_Mem/n6152 ,
         \Data_Mem/n6151 , \Data_Mem/n6150 , \Data_Mem/n6149 ,
         \Data_Mem/n6148 , \Data_Mem/n6147 , \Data_Mem/n6146 ,
         \Data_Mem/n6145 , \Data_Mem/n6144 , \Data_Mem/n6143 ,
         \Data_Mem/n6142 , \Data_Mem/n6141 , \Data_Mem/n6140 ,
         \Data_Mem/n6139 , \Data_Mem/n6138 , \Data_Mem/n6137 ,
         \Data_Mem/n6136 , \Data_Mem/n6135 , \Data_Mem/n6134 ,
         \Data_Mem/n6133 , \Data_Mem/n6132 , \Data_Mem/n6131 ,
         \Data_Mem/n6130 , \Data_Mem/n6129 , \Data_Mem/n6128 ,
         \Data_Mem/n6127 , \Data_Mem/n6126 , \Data_Mem/n6125 ,
         \Data_Mem/n6124 , \Data_Mem/n6123 , \Data_Mem/n6122 ,
         \Data_Mem/n6121 , \Data_Mem/n6120 , \Data_Mem/n6119 ,
         \Data_Mem/n6118 , \Data_Mem/n6117 , \Data_Mem/n6116 ,
         \Data_Mem/n6115 , \Data_Mem/n6114 , \Data_Mem/n6113 ,
         \Data_Mem/n6112 , \Data_Mem/n6111 , \Data_Mem/n6110 ,
         \Data_Mem/n6109 , \Data_Mem/n6108 , \Data_Mem/n6107 ,
         \Data_Mem/n6106 , \Data_Mem/n6105 , \Data_Mem/n6104 ,
         \Data_Mem/n6103 , \Data_Mem/n6102 , \Data_Mem/n6101 ,
         \Data_Mem/n6100 , \Data_Mem/n6099 , \Data_Mem/n6098 ,
         \Data_Mem/n6097 , \Data_Mem/n6096 , \Data_Mem/n6095 ,
         \Data_Mem/n6094 , \Data_Mem/n6093 , \Data_Mem/n6092 ,
         \Data_Mem/n6091 , \Data_Mem/n6090 , \Data_Mem/n6089 ,
         \Data_Mem/n6088 , \Data_Mem/n6087 , \Data_Mem/n6086 ,
         \Data_Mem/n6085 , \Data_Mem/n6084 , \Data_Mem/n6083 ,
         \Data_Mem/n6082 , \Data_Mem/n6081 , \Data_Mem/n6080 ,
         \Data_Mem/n6079 , \Data_Mem/n6078 , \Data_Mem/n6077 ,
         \Data_Mem/n6076 , \Data_Mem/n6075 , \Data_Mem/n6074 ,
         \Data_Mem/n6073 , \Data_Mem/n6072 , \Data_Mem/n6071 ,
         \Data_Mem/n6070 , \Data_Mem/n6069 , \Data_Mem/n6068 ,
         \Data_Mem/n6067 , \Data_Mem/n6066 , \Data_Mem/n6065 ,
         \Data_Mem/n6064 , \Data_Mem/n6063 , \Data_Mem/n6062 ,
         \Data_Mem/n6061 , \Data_Mem/n6060 , \Data_Mem/n6059 ,
         \Data_Mem/n6058 , \Data_Mem/n6057 , \Data_Mem/n6056 ,
         \Data_Mem/n6055 , \Data_Mem/n6054 , \Data_Mem/n6053 ,
         \Data_Mem/n6052 , \Data_Mem/n6051 , \Data_Mem/n6050 ,
         \Data_Mem/n6049 , \Data_Mem/n6048 , \Data_Mem/n6047 ,
         \Data_Mem/n6046 , \Data_Mem/n6045 , \Data_Mem/n6044 ,
         \Data_Mem/n6043 , \Data_Mem/n6042 , \Data_Mem/n6041 ,
         \Data_Mem/n6040 , \Data_Mem/n6039 , \Data_Mem/n6038 ,
         \Data_Mem/n6037 , \Data_Mem/n6036 , \Data_Mem/n6035 ,
         \Data_Mem/n6034 , \Data_Mem/n6033 , \Data_Mem/n6032 ,
         \Data_Mem/n6031 , \Data_Mem/n6030 , \Data_Mem/n6029 ,
         \Data_Mem/n6028 , \Data_Mem/n6027 , \Data_Mem/n6026 ,
         \Data_Mem/n6025 , \Data_Mem/n6024 , \Data_Mem/n6023 ,
         \Data_Mem/n6022 , \Data_Mem/n6021 , \Data_Mem/n6020 ,
         \Data_Mem/n6019 , \Data_Mem/n6018 , \Data_Mem/n6017 ,
         \Data_Mem/n6016 , \Data_Mem/n6015 , \Data_Mem/n6014 ,
         \Data_Mem/n6013 , \Data_Mem/n6012 , \Data_Mem/n6011 ,
         \Data_Mem/n6010 , \Data_Mem/n6009 , \Data_Mem/n6008 ,
         \Data_Mem/n6007 , \Data_Mem/n6006 , \Data_Mem/n6005 ,
         \Data_Mem/n6004 , \Data_Mem/n6003 , \Data_Mem/n6002 ,
         \Data_Mem/n6001 , \Data_Mem/n6000 , \Data_Mem/n5999 ,
         \Data_Mem/n5998 , \Data_Mem/n5997 , \Data_Mem/n5996 ,
         \Data_Mem/n5995 , \Data_Mem/n5994 , \Data_Mem/n5993 ,
         \Data_Mem/n5992 , \Data_Mem/n5991 , \Data_Mem/n5990 ,
         \Data_Mem/n5989 , \Data_Mem/n5988 , \Data_Mem/n5987 ,
         \Data_Mem/n5986 , \Data_Mem/n5985 , \Data_Mem/n5984 ,
         \Data_Mem/n5983 , \Data_Mem/n5982 , \Data_Mem/n5981 ,
         \Data_Mem/n5980 , \Data_Mem/n5979 , \Data_Mem/n5978 ,
         \Data_Mem/n5977 , \Data_Mem/n5976 , \Data_Mem/n5975 ,
         \Data_Mem/n5974 , \Data_Mem/n5973 , \Data_Mem/n5972 ,
         \Data_Mem/n5971 , \Data_Mem/n5970 , \Data_Mem/n5969 ,
         \Data_Mem/n5968 , \Data_Mem/n5967 , \Data_Mem/n5966 ,
         \Data_Mem/n5965 , \Data_Mem/n5964 , \Data_Mem/n5963 ,
         \Data_Mem/n5962 , \Data_Mem/n5961 , \Data_Mem/n5960 ,
         \Data_Mem/n5959 , \Data_Mem/n5958 , \Data_Mem/n5957 ,
         \Data_Mem/n5956 , \Data_Mem/n5955 , \Data_Mem/n5954 ,
         \Data_Mem/n5953 , \Data_Mem/n5952 , \Data_Mem/n5951 ,
         \Data_Mem/n5950 , \Data_Mem/n5949 , \Data_Mem/n5948 ,
         \Data_Mem/n5947 , \Data_Mem/n5946 , \Data_Mem/n5945 ,
         \Data_Mem/n5944 , \Data_Mem/n5943 , \Data_Mem/n5942 ,
         \Data_Mem/n5941 , \Data_Mem/n5940 , \Data_Mem/n5939 ,
         \Data_Mem/n5938 , \Data_Mem/n5937 , \Data_Mem/n5936 ,
         \Data_Mem/n5935 , \Data_Mem/n5934 , \Data_Mem/n5933 ,
         \Data_Mem/n5932 , \Data_Mem/n5931 , \Data_Mem/n5930 ,
         \Data_Mem/n5929 , \Data_Mem/n5928 , \Data_Mem/n5927 ,
         \Data_Mem/n5926 , \Data_Mem/n5925 , \Data_Mem/n5924 ,
         \Data_Mem/n5923 , \Data_Mem/n5922 , \Data_Mem/n5921 ,
         \Data_Mem/n5920 , \Data_Mem/n5919 , \Data_Mem/n5918 ,
         \Data_Mem/n5917 , \Data_Mem/n5916 , \Data_Mem/n5915 ,
         \Data_Mem/n5914 , \Data_Mem/n5913 , \Data_Mem/n5912 ,
         \Data_Mem/n5911 , \Data_Mem/n5910 , \Data_Mem/n5909 ,
         \Data_Mem/n5908 , \Data_Mem/n5907 , \Data_Mem/n5906 ,
         \Data_Mem/n5905 , \Data_Mem/n5904 , \Data_Mem/n5903 ,
         \Data_Mem/n5902 , \Data_Mem/n5901 , \Data_Mem/n5900 ,
         \Data_Mem/n5899 , \Data_Mem/n5898 , \Data_Mem/n5897 ,
         \Data_Mem/n5896 , \Data_Mem/n5895 , \Data_Mem/n5894 ,
         \Data_Mem/n5893 , \Data_Mem/n5892 , \Data_Mem/n5891 ,
         \Data_Mem/n5890 , \Data_Mem/n5889 , \Data_Mem/n5888 ,
         \Data_Mem/n5887 , \Data_Mem/n5886 , \Data_Mem/n5885 ,
         \Data_Mem/n5884 , \Data_Mem/n5883 , \Data_Mem/n5882 ,
         \Data_Mem/n5881 , \Data_Mem/n5880 , \Data_Mem/n5879 ,
         \Data_Mem/n5878 , \Data_Mem/n5877 , \Data_Mem/n5876 ,
         \Data_Mem/n5875 , \Data_Mem/n5874 , \Data_Mem/n5873 ,
         \Data_Mem/n5872 , \Data_Mem/n5871 , \Data_Mem/n5870 ,
         \Data_Mem/n5869 , \Data_Mem/n5868 , \Data_Mem/n5867 ,
         \Data_Mem/n5866 , \Data_Mem/n5865 , \Data_Mem/n5864 ,
         \Data_Mem/n5863 , \Data_Mem/n5862 , \Data_Mem/n5861 ,
         \Data_Mem/n5860 , \Data_Mem/n5859 , \Data_Mem/n5858 ,
         \Data_Mem/n5857 , \Data_Mem/n5856 , \Data_Mem/n5855 ,
         \Data_Mem/n5854 , \Data_Mem/n5853 , \Data_Mem/n5852 ,
         \Data_Mem/n5851 , \Data_Mem/n5850 , \Data_Mem/n5849 ,
         \Data_Mem/n5848 , \Data_Mem/n5847 , \Data_Mem/n5846 ,
         \Data_Mem/n5845 , \Data_Mem/n5844 , \Data_Mem/n5843 ,
         \Data_Mem/n5842 , \Data_Mem/n5841 , \Data_Mem/n5840 ,
         \Data_Mem/n5839 , \Data_Mem/n5838 , \Data_Mem/n5837 ,
         \Data_Mem/n5836 , \Data_Mem/n5835 , \Data_Mem/n5834 ,
         \Data_Mem/n5833 , \Data_Mem/n5832 , \Data_Mem/n5831 ,
         \Data_Mem/n5830 , \Data_Mem/n5829 , \Data_Mem/n5828 ,
         \Data_Mem/n5827 , \Data_Mem/n5826 , \Data_Mem/n5825 ,
         \Data_Mem/n5824 , \Data_Mem/n5823 , \Data_Mem/n5822 ,
         \Data_Mem/n5821 , \Data_Mem/n5820 , \Data_Mem/n5819 ,
         \Data_Mem/n5818 , \Data_Mem/n5817 , \Data_Mem/n5816 ,
         \Data_Mem/n5815 , \Data_Mem/n5814 , \Data_Mem/n5813 ,
         \Data_Mem/n5812 , \Data_Mem/n5811 , \Data_Mem/n5810 ,
         \Data_Mem/n5809 , \Data_Mem/n5808 , \Data_Mem/n5807 ,
         \Data_Mem/n5806 , \Data_Mem/n5805 , \Data_Mem/n5804 ,
         \Data_Mem/n5803 , \Data_Mem/n5802 , \Data_Mem/n5801 ,
         \Data_Mem/n5800 , \Data_Mem/n5799 , \Data_Mem/n5798 ,
         \Data_Mem/n5797 , \Data_Mem/n5796 , \Data_Mem/n5795 ,
         \Data_Mem/n5794 , \Data_Mem/n5793 , \Data_Mem/n5792 ,
         \Data_Mem/n5791 , \Data_Mem/n5790 , \Data_Mem/n5789 ,
         \Data_Mem/n5788 , \Data_Mem/n5787 , \Data_Mem/n5786 ,
         \Data_Mem/n5785 , \Data_Mem/n5784 , \Data_Mem/n5783 ,
         \Data_Mem/n5782 , \Data_Mem/n5781 , \Data_Mem/n5780 ,
         \Data_Mem/n5779 , \Data_Mem/n5778 , \Data_Mem/n5777 ,
         \Data_Mem/n5776 , \Data_Mem/n5775 , \Data_Mem/n5774 ,
         \Data_Mem/n5773 , \Data_Mem/n5772 , \Data_Mem/n5771 ,
         \Data_Mem/n5770 , \Data_Mem/n5769 , \Data_Mem/n5768 ,
         \Data_Mem/n5767 , \Data_Mem/n5766 , \Data_Mem/n5765 ,
         \Data_Mem/n5764 , \Data_Mem/n5763 , \Data_Mem/n5762 ,
         \Data_Mem/n5761 , \Data_Mem/n5760 , \Data_Mem/n5759 ,
         \Data_Mem/n5758 , \Data_Mem/n5757 , \Data_Mem/n5756 ,
         \Data_Mem/n5755 , \Data_Mem/n5754 , \Data_Mem/n5753 ,
         \Data_Mem/n5752 , \Data_Mem/n5751 , \Data_Mem/n5750 ,
         \Data_Mem/n5749 , \Data_Mem/n5748 , \Data_Mem/n5747 ,
         \Data_Mem/n5746 , \Data_Mem/n5745 , \Data_Mem/n5744 ,
         \Data_Mem/n5743 , \Data_Mem/n5742 , \Data_Mem/n5741 ,
         \Data_Mem/n5740 , \Data_Mem/n5739 , \Data_Mem/n5738 ,
         \Data_Mem/n5737 , \Data_Mem/n5736 , \Data_Mem/n5735 ,
         \Data_Mem/n5734 , \Data_Mem/n5733 , \Data_Mem/n5732 ,
         \Data_Mem/n5731 , \Data_Mem/n5730 , \Data_Mem/n5729 ,
         \Data_Mem/n5728 , \Data_Mem/n5727 , \Data_Mem/n5726 ,
         \Data_Mem/n5725 , \Data_Mem/n5724 , \Data_Mem/n5723 ,
         \Data_Mem/n5722 , \Data_Mem/n5721 , \Data_Mem/n5720 ,
         \Data_Mem/n5719 , \Data_Mem/n5718 , \Data_Mem/n5717 ,
         \Data_Mem/n5716 , \Data_Mem/n5715 , \Data_Mem/n5714 ,
         \Data_Mem/n5713 , \Data_Mem/N745 , \Data_Mem/N744 , \Data_Mem/N743 ,
         \Data_Mem/N742 , \Data_Mem/N741 , \Data_Mem/N740 , \Data_Mem/N739 ,
         \Data_Mem/N738 , \Data_Mem/N737 , \Data_Mem/N736 , \Data_Mem/N735 ,
         \Data_Mem/N734 , \Data_Mem/N733 , \Data_Mem/N732 , \Data_Mem/N731 ,
         \Data_Mem/N730 , \Data_Mem/N729 , \Data_Mem/N728 , \Data_Mem/N727 ,
         \Data_Mem/N726 , \Data_Mem/N725 , \Data_Mem/N724 , \Data_Mem/N723 ,
         \Data_Mem/N722 , \Data_Mem/N721 , \Data_Mem/N720 , \Data_Mem/N719 ,
         \Data_Mem/N718 , \Data_Mem/N717 , \Data_Mem/N716 , \Data_Mem/N715 ,
         \Data_Mem/N714 , \Reg_Bank/n5939 , \Reg_Bank/n5938 , \Reg_Bank/n5937 ,
         \Reg_Bank/n5936 , \Reg_Bank/n5935 , \Reg_Bank/n5934 ,
         \Reg_Bank/n5933 , \Reg_Bank/n5932 , \Reg_Bank/n5931 ,
         \Reg_Bank/n5930 , \Reg_Bank/n5929 , \Reg_Bank/n5928 ,
         \Reg_Bank/n5927 , \Reg_Bank/n5926 , \Reg_Bank/n5925 ,
         \Reg_Bank/n5924 , \Reg_Bank/n5923 , \Reg_Bank/n5922 ,
         \Reg_Bank/n5921 , \Reg_Bank/n5920 , \Reg_Bank/n5919 ,
         \Reg_Bank/n5918 , \Reg_Bank/n5917 , \Reg_Bank/n5916 ,
         \Reg_Bank/n5915 , \Reg_Bank/n5914 , \Reg_Bank/n5913 ,
         \Reg_Bank/n5912 , \Reg_Bank/n5911 , \Reg_Bank/n5910 ,
         \Reg_Bank/n5909 , \Reg_Bank/n5908 , \Reg_Bank/n5907 ,
         \Reg_Bank/n5906 , \Reg_Bank/n5905 , \Reg_Bank/n5904 ,
         \Reg_Bank/n5903 , \Reg_Bank/n5902 , \Reg_Bank/n5901 ,
         \Reg_Bank/n5900 , \Reg_Bank/n5899 , \Reg_Bank/n5898 ,
         \Reg_Bank/n5897 , \Reg_Bank/n5896 , \Reg_Bank/n5895 ,
         \Reg_Bank/n5894 , \Reg_Bank/n5893 , \Reg_Bank/n5892 ,
         \Reg_Bank/n5891 , \Reg_Bank/n5890 , \Reg_Bank/n5889 ,
         \Reg_Bank/n5888 , \Reg_Bank/n5887 , \Reg_Bank/n5886 ,
         \Reg_Bank/n5885 , \Reg_Bank/n5884 , \Reg_Bank/n5883 ,
         \Reg_Bank/n5882 , \Reg_Bank/n5881 , \Reg_Bank/n5880 ,
         \Reg_Bank/n5879 , \Reg_Bank/n5878 , \Reg_Bank/n5877 ,
         \Reg_Bank/n5876 , \Reg_Bank/n5875 , \Reg_Bank/n5874 ,
         \Reg_Bank/n5873 , \Reg_Bank/n5872 , \Reg_Bank/n5871 ,
         \Reg_Bank/n5870 , \Reg_Bank/n5869 , \Reg_Bank/n5868 ,
         \Reg_Bank/n5867 , \Reg_Bank/n5866 , \Reg_Bank/n5865 ,
         \Reg_Bank/n5864 , \Reg_Bank/n5863 , \Reg_Bank/n5862 ,
         \Reg_Bank/n5861 , \Reg_Bank/n5860 , \Reg_Bank/n5859 ,
         \Reg_Bank/n5858 , \Reg_Bank/n5857 , \Reg_Bank/n5856 ,
         \Reg_Bank/n5855 , \Reg_Bank/n5854 , \Reg_Bank/n5853 ,
         \Reg_Bank/n5852 , \Reg_Bank/n5851 , \Reg_Bank/n5850 ,
         \Reg_Bank/n5849 , \Reg_Bank/n5848 , \Reg_Bank/n5847 ,
         \Reg_Bank/n5846 , \Reg_Bank/n5845 , \Reg_Bank/n5844 ,
         \Reg_Bank/n5843 , \Reg_Bank/n5842 , \Reg_Bank/n5841 ,
         \Reg_Bank/n5840 , \Reg_Bank/n5839 , \Reg_Bank/n5838 ,
         \Reg_Bank/n5837 , \Reg_Bank/n5836 , \Reg_Bank/n5835 ,
         \Reg_Bank/n5834 , \Reg_Bank/n5833 , \Reg_Bank/n5832 ,
         \Reg_Bank/n5831 , \Reg_Bank/n5830 , \Reg_Bank/n5829 ,
         \Reg_Bank/n5828 , \Reg_Bank/n5827 , \Reg_Bank/n5826 ,
         \Reg_Bank/n5825 , \Reg_Bank/n5824 , \Reg_Bank/n5823 ,
         \Reg_Bank/n5822 , \Reg_Bank/n5821 , \Reg_Bank/n5820 ,
         \Reg_Bank/n5819 , \Reg_Bank/n5818 , \Reg_Bank/n5817 ,
         \Reg_Bank/n5816 , \Reg_Bank/n5815 , \Reg_Bank/n5814 ,
         \Reg_Bank/n5813 , \Reg_Bank/n5812 , \Reg_Bank/n5811 ,
         \Reg_Bank/n5810 , \Reg_Bank/n5809 , \Reg_Bank/n5808 ,
         \Reg_Bank/n5807 , \Reg_Bank/n5806 , \Reg_Bank/n5805 ,
         \Reg_Bank/n5804 , \Reg_Bank/n5803 , \Reg_Bank/n5802 ,
         \Reg_Bank/n5801 , \Reg_Bank/n5800 , \Reg_Bank/n5799 ,
         \Reg_Bank/n5798 , \Reg_Bank/n5797 , \Reg_Bank/n5796 ,
         \Reg_Bank/n5795 , \Reg_Bank/n5794 , \Reg_Bank/n5793 ,
         \Reg_Bank/n5792 , \Reg_Bank/n5791 , \Reg_Bank/n5790 ,
         \Reg_Bank/n5789 , \Reg_Bank/n5788 , \Reg_Bank/n5787 ,
         \Reg_Bank/n5786 , \Reg_Bank/n5785 , \Reg_Bank/n5784 ,
         \Reg_Bank/n5783 , \Reg_Bank/n5782 , \Reg_Bank/n5781 ,
         \Reg_Bank/n5780 , \Reg_Bank/n5779 , \Reg_Bank/n5778 ,
         \Reg_Bank/n5777 , \Reg_Bank/n5776 , \Reg_Bank/n5775 ,
         \Reg_Bank/n5774 , \Reg_Bank/n5773 , \Reg_Bank/n5772 ,
         \Reg_Bank/n5771 , \Reg_Bank/n5770 , \Reg_Bank/n5769 ,
         \Reg_Bank/n5768 , \Reg_Bank/n5767 , \Reg_Bank/n5766 ,
         \Reg_Bank/n5765 , \Reg_Bank/n5764 , \Reg_Bank/n5763 ,
         \Reg_Bank/n5762 , \Reg_Bank/n5761 , \Reg_Bank/n5760 ,
         \Reg_Bank/n5759 , \Reg_Bank/n5758 , \Reg_Bank/n5757 ,
         \Reg_Bank/n5756 , \Reg_Bank/n5755 , \Reg_Bank/n5754 ,
         \Reg_Bank/n5753 , \Reg_Bank/n5752 , \Reg_Bank/n5751 ,
         \Reg_Bank/n5750 , \Reg_Bank/n5749 , \Reg_Bank/n5748 ,
         \Reg_Bank/n5747 , \Reg_Bank/n5746 , \Reg_Bank/n5745 ,
         \Reg_Bank/n5744 , \Reg_Bank/n5743 , \Reg_Bank/n5742 ,
         \Reg_Bank/n5741 , \Reg_Bank/n5740 , \Reg_Bank/n5739 ,
         \Reg_Bank/n5738 , \Reg_Bank/n5737 , \Reg_Bank/n5736 ,
         \Reg_Bank/n5735 , \Reg_Bank/n5734 , \Reg_Bank/n5733 ,
         \Reg_Bank/n5732 , \Reg_Bank/n5731 , \Reg_Bank/n5730 ,
         \Reg_Bank/n5729 , \Reg_Bank/n5728 , \Reg_Bank/n5727 ,
         \Reg_Bank/n5726 , \Reg_Bank/n5725 , \Reg_Bank/n5724 ,
         \Reg_Bank/n5723 , \Reg_Bank/n5722 , \Reg_Bank/n5721 ,
         \Reg_Bank/n5720 , \Reg_Bank/n5719 , \Reg_Bank/n5718 ,
         \Reg_Bank/n5717 , \Reg_Bank/n5716 , \Reg_Bank/n5715 ,
         \Reg_Bank/n5714 , \Reg_Bank/n5713 , \Reg_Bank/n5712 ,
         \Reg_Bank/n5711 , \Reg_Bank/n5710 , \Reg_Bank/n5709 ,
         \Reg_Bank/n5708 , \Reg_Bank/n5707 , \Reg_Bank/n5706 ,
         \Reg_Bank/n5705 , \Reg_Bank/n5704 , \Reg_Bank/n5703 ,
         \Reg_Bank/n5702 , \Reg_Bank/n5701 , \Reg_Bank/n5700 ,
         \Reg_Bank/n5699 , \Reg_Bank/n5698 , \Reg_Bank/n5697 ,
         \Reg_Bank/n5696 , \Reg_Bank/n5695 , \Reg_Bank/n5694 ,
         \Reg_Bank/n5693 , \Reg_Bank/n5692 , \Reg_Bank/n5691 ,
         \Reg_Bank/n5690 , \Reg_Bank/n5689 , \Reg_Bank/n5688 ,
         \Reg_Bank/n5687 , \Reg_Bank/n5686 , \Reg_Bank/n5685 ,
         \Reg_Bank/n5684 , \Reg_Bank/n5683 , \Reg_Bank/n5682 ,
         \Reg_Bank/n5681 , \Reg_Bank/n5680 , \Reg_Bank/n5679 ,
         \Reg_Bank/n5678 , \Reg_Bank/n5677 , \Reg_Bank/n5676 ,
         \Reg_Bank/n5675 , \Reg_Bank/n5674 , \Reg_Bank/n5673 ,
         \Reg_Bank/n5672 , \Reg_Bank/n5671 , \Reg_Bank/n5670 ,
         \Reg_Bank/n5669 , \Reg_Bank/n5668 , \Reg_Bank/n5667 ,
         \Reg_Bank/n5666 , \Reg_Bank/n5665 , \Reg_Bank/n5664 ,
         \Reg_Bank/n5663 , \Reg_Bank/n5662 , \Reg_Bank/n5661 ,
         \Reg_Bank/n5660 , \Reg_Bank/n5659 , \Reg_Bank/n5658 ,
         \Reg_Bank/n5657 , \Reg_Bank/n5656 , \Reg_Bank/n5655 ,
         \Reg_Bank/n5654 , \Reg_Bank/n5653 , \Reg_Bank/n5652 ,
         \Reg_Bank/n5651 , \Reg_Bank/n5650 , \Reg_Bank/n5649 ,
         \Reg_Bank/n5648 , \Reg_Bank/n5647 , \Reg_Bank/n5646 ,
         \Reg_Bank/n5645 , \Reg_Bank/n5644 , \Reg_Bank/n5643 ,
         \Reg_Bank/n5642 , \Reg_Bank/n5641 , \Reg_Bank/n5640 ,
         \Reg_Bank/n5639 , \Reg_Bank/n5638 , \Reg_Bank/n5637 ,
         \Reg_Bank/n5636 , \Reg_Bank/n5635 , \Reg_Bank/n5634 ,
         \Reg_Bank/n5633 , \Reg_Bank/n5632 , \Reg_Bank/n5631 ,
         \Reg_Bank/n5630 , \Reg_Bank/n5629 , \Reg_Bank/n5628 ,
         \Reg_Bank/n5627 , \Reg_Bank/n5626 , \Reg_Bank/n5625 ,
         \Reg_Bank/n5624 , \Reg_Bank/n5623 , \Reg_Bank/n5622 ,
         \Reg_Bank/n5621 , \Reg_Bank/n5620 , \Reg_Bank/n5619 ,
         \Reg_Bank/n5618 , \Reg_Bank/n5617 , \Reg_Bank/n5616 ,
         \Reg_Bank/n5615 , \Reg_Bank/n5614 , \Reg_Bank/n5613 ,
         \Reg_Bank/n5612 , \Reg_Bank/n5611 , \Reg_Bank/n5610 ,
         \Reg_Bank/n5609 , \Reg_Bank/n5608 , \Reg_Bank/n5607 ,
         \Reg_Bank/n5606 , \Reg_Bank/n5605 , \Reg_Bank/n5604 ,
         \Reg_Bank/n5603 , \Reg_Bank/n5602 , \Reg_Bank/n5601 ,
         \Reg_Bank/n5600 , \Reg_Bank/n5599 , \Reg_Bank/n5598 ,
         \Reg_Bank/n5597 , \Reg_Bank/n5596 , \Reg_Bank/n5595 ,
         \Reg_Bank/n5594 , \Reg_Bank/n5593 , \Reg_Bank/n5592 ,
         \Reg_Bank/n5591 , \Reg_Bank/n5590 , \Reg_Bank/n5589 ,
         \Reg_Bank/n5588 , \Reg_Bank/n5587 , \Reg_Bank/n5586 ,
         \Reg_Bank/n5585 , \Reg_Bank/n5584 , \Reg_Bank/n5583 ,
         \Reg_Bank/n5582 , \Reg_Bank/n5581 , \Reg_Bank/n5580 ,
         \Reg_Bank/n5579 , \Reg_Bank/n5578 , \Reg_Bank/n5577 ,
         \Reg_Bank/n5576 , \Reg_Bank/n5575 , \Reg_Bank/n5574 ,
         \Reg_Bank/n5573 , \Reg_Bank/n5572 , \Reg_Bank/n5571 ,
         \Reg_Bank/n5570 , \Reg_Bank/n5569 , \Reg_Bank/n5568 ,
         \Reg_Bank/n5567 , \Reg_Bank/n5566 , \Reg_Bank/n5565 ,
         \Reg_Bank/n5564 , \Reg_Bank/n5563 , \Reg_Bank/n5562 ,
         \Reg_Bank/n5561 , \Reg_Bank/n5560 , \Reg_Bank/n5559 ,
         \Reg_Bank/n5558 , \Reg_Bank/n5557 , \Reg_Bank/n5556 ,
         \Reg_Bank/n5555 , \Reg_Bank/n5554 , \Reg_Bank/n5553 ,
         \Reg_Bank/n5552 , \Reg_Bank/n5551 , \Reg_Bank/n5550 ,
         \Reg_Bank/n5549 , \Reg_Bank/n5548 , \Reg_Bank/n5547 ,
         \Reg_Bank/n5546 , \Reg_Bank/n5545 , \Reg_Bank/n5544 ,
         \Reg_Bank/n5543 , \Reg_Bank/n5542 , \Reg_Bank/n5541 ,
         \Reg_Bank/n5540 , \Reg_Bank/n5539 , \Reg_Bank/n5538 ,
         \Reg_Bank/n5537 , \Reg_Bank/n5536 , \Reg_Bank/n5535 ,
         \Reg_Bank/n5534 , \Reg_Bank/n5533 , \Reg_Bank/n5532 ,
         \Reg_Bank/n5531 , \Reg_Bank/n5530 , \Reg_Bank/n5529 ,
         \Reg_Bank/n5528 , \Reg_Bank/n5527 , \Reg_Bank/n5526 ,
         \Reg_Bank/n5525 , \Reg_Bank/n5524 , \Reg_Bank/n5523 ,
         \Reg_Bank/n5522 , \Reg_Bank/n5521 , \Reg_Bank/n5520 ,
         \Reg_Bank/n5519 , \Reg_Bank/n5518 , \Reg_Bank/n5517 ,
         \Reg_Bank/n5516 , \Reg_Bank/n5515 , \Reg_Bank/n5514 ,
         \Reg_Bank/n5513 , \Reg_Bank/n5512 , \Reg_Bank/n5511 ,
         \Reg_Bank/n5510 , \Reg_Bank/n5509 , \Reg_Bank/n5508 ,
         \Reg_Bank/n5507 , \Reg_Bank/n5506 , \Reg_Bank/n5505 ,
         \Reg_Bank/n5504 , \Reg_Bank/n5503 , \Reg_Bank/n5502 ,
         \Reg_Bank/n5501 , \Reg_Bank/n5500 , \Reg_Bank/n5499 ,
         \Reg_Bank/n5498 , \Reg_Bank/n5497 , \Reg_Bank/n5496 ,
         \Reg_Bank/n5495 , \Reg_Bank/n5494 , \Reg_Bank/n5493 ,
         \Reg_Bank/n5492 , \Reg_Bank/n5491 , \Reg_Bank/n5490 ,
         \Reg_Bank/n5489 , \Reg_Bank/n5488 , \Reg_Bank/n5487 ,
         \Reg_Bank/n5486 , \Reg_Bank/n5485 , \Reg_Bank/n5484 ,
         \Reg_Bank/n5483 , \Reg_Bank/n5482 , \Reg_Bank/n5481 ,
         \Reg_Bank/n5480 , \Reg_Bank/n5479 , \Reg_Bank/n5478 ,
         \Reg_Bank/n5477 , \Reg_Bank/n5476 , \Reg_Bank/n5475 ,
         \Reg_Bank/n5474 , \Reg_Bank/n5473 , \Reg_Bank/n5472 ,
         \Reg_Bank/n5471 , \Reg_Bank/n5470 , \Reg_Bank/n5469 ,
         \Reg_Bank/n5468 , \Reg_Bank/n5467 , \Reg_Bank/n5466 ,
         \Reg_Bank/n5465 , \Reg_Bank/n5464 , \Reg_Bank/n5463 ,
         \Reg_Bank/n5462 , \Reg_Bank/n5461 , \Reg_Bank/n5460 ,
         \Reg_Bank/n5459 , \Reg_Bank/n5458 , \Reg_Bank/n5457 ,
         \Reg_Bank/n5456 , \Reg_Bank/n5455 , \Reg_Bank/n5454 ,
         \Reg_Bank/n5453 , \Reg_Bank/n5452 , \Reg_Bank/n5451 ,
         \Reg_Bank/n5450 , \Reg_Bank/n5449 , \Reg_Bank/n5448 ,
         \Reg_Bank/n5447 , \Reg_Bank/n5446 , \Reg_Bank/n5445 ,
         \Reg_Bank/n5444 , \Reg_Bank/n5443 , \Reg_Bank/n5442 ,
         \Reg_Bank/n5441 , \Reg_Bank/n5440 , \Reg_Bank/n5439 ,
         \Reg_Bank/n5438 , \Reg_Bank/n5437 , \Reg_Bank/n5436 ,
         \Reg_Bank/n5435 , \Reg_Bank/n5434 , \Reg_Bank/n5433 ,
         \Reg_Bank/n5432 , \Reg_Bank/n5431 , \Reg_Bank/n5430 ,
         \Reg_Bank/n5429 , \Reg_Bank/n5428 , \Reg_Bank/n5427 ,
         \Reg_Bank/n5426 , \Reg_Bank/n5425 , \Reg_Bank/n5424 ,
         \Reg_Bank/n5423 , \Reg_Bank/n5422 , \Reg_Bank/n5421 ,
         \Reg_Bank/n5420 , \Reg_Bank/n5419 , \Reg_Bank/n5418 ,
         \Reg_Bank/n5417 , \Reg_Bank/n5416 , \Reg_Bank/n5415 ,
         \Reg_Bank/n5414 , \Reg_Bank/n5413 , \Reg_Bank/n5412 ,
         \Reg_Bank/n5411 , \Reg_Bank/n5410 , \Reg_Bank/n5409 ,
         \Reg_Bank/n5408 , \Reg_Bank/n5407 , \Reg_Bank/n5406 ,
         \Reg_Bank/n5405 , \Reg_Bank/n5404 , \Reg_Bank/n5403 ,
         \Reg_Bank/n5402 , \Reg_Bank/n5401 , \Reg_Bank/n5400 ,
         \Reg_Bank/n5399 , \Reg_Bank/n5398 , \Reg_Bank/n5397 ,
         \Reg_Bank/n5396 , \Reg_Bank/n5395 , \Reg_Bank/n5394 ,
         \Reg_Bank/n5393 , \Reg_Bank/n5392 , \Reg_Bank/n5391 ,
         \Reg_Bank/n5390 , \Reg_Bank/n5389 , \Reg_Bank/n5388 ,
         \Reg_Bank/n5387 , \Reg_Bank/n5386 , \Reg_Bank/n5385 ,
         \Reg_Bank/n5384 , \Reg_Bank/n5383 , \Reg_Bank/n5382 ,
         \Reg_Bank/n5381 , \Reg_Bank/n5380 , \Reg_Bank/n5379 ,
         \Reg_Bank/n5378 , \Reg_Bank/n5377 , \Reg_Bank/n5376 ,
         \Reg_Bank/n5375 , \Reg_Bank/n5374 , \Reg_Bank/n5373 ,
         \Reg_Bank/n5372 , \Reg_Bank/n5371 , \Reg_Bank/n5370 ,
         \Reg_Bank/n5369 , \Reg_Bank/n5368 , \Reg_Bank/n5367 ,
         \Reg_Bank/n5366 , \Reg_Bank/n5365 , \Reg_Bank/n5364 ,
         \Reg_Bank/n5363 , \Reg_Bank/n5362 , \Reg_Bank/n5361 ,
         \Reg_Bank/n5360 , \Reg_Bank/n5359 , \Reg_Bank/n5358 ,
         \Reg_Bank/n5357 , \Reg_Bank/n5356 , \Reg_Bank/n5355 ,
         \Reg_Bank/n5354 , \Reg_Bank/n5353 , \Reg_Bank/n5352 ,
         \Reg_Bank/n5351 , \Reg_Bank/n5350 , \Reg_Bank/n5349 ,
         \Reg_Bank/n5348 , \Reg_Bank/n5347 , \Reg_Bank/n5346 ,
         \Reg_Bank/n5345 , \Reg_Bank/n5344 , \Reg_Bank/n5343 ,
         \Reg_Bank/n5342 , \Reg_Bank/n5341 , \Reg_Bank/n5340 ,
         \Reg_Bank/n5339 , \Reg_Bank/n5338 , \Reg_Bank/n5337 ,
         \Reg_Bank/n5336 , \Reg_Bank/n5335 , \Reg_Bank/n5334 ,
         \Reg_Bank/n5333 , \Reg_Bank/n5332 , \Reg_Bank/n5331 ,
         \Reg_Bank/n5330 , \Reg_Bank/n5329 , \Reg_Bank/n5328 ,
         \Reg_Bank/n5327 , \Reg_Bank/n5326 , \Reg_Bank/n5325 ,
         \Reg_Bank/n5324 , \Reg_Bank/n5323 , \Reg_Bank/n5322 ,
         \Reg_Bank/n5321 , \Reg_Bank/n5320 , \Reg_Bank/n5319 ,
         \Reg_Bank/n5318 , \Reg_Bank/n5317 , \Reg_Bank/n5316 ,
         \Reg_Bank/n5315 , \Reg_Bank/n5314 , \Reg_Bank/n5313 ,
         \Reg_Bank/n5312 , \Reg_Bank/n5311 , \Reg_Bank/n5310 ,
         \Reg_Bank/n5309 , \Reg_Bank/n5308 , \Reg_Bank/n5307 ,
         \Reg_Bank/n5306 , \Reg_Bank/n5305 , \Reg_Bank/n5304 ,
         \Reg_Bank/n5303 , \Reg_Bank/n5302 , \Reg_Bank/n5301 ,
         \Reg_Bank/n5300 , \Reg_Bank/n5299 , \Reg_Bank/n5298 ,
         \Reg_Bank/n5297 , \Reg_Bank/n5296 , \Reg_Bank/n5295 ,
         \Reg_Bank/n5294 , \Reg_Bank/n5293 , \Reg_Bank/n5292 ,
         \Reg_Bank/n5291 , \Reg_Bank/n5290 , \Reg_Bank/n5289 ,
         \Reg_Bank/n5288 , \Reg_Bank/n5287 , \Reg_Bank/n5286 ,
         \Reg_Bank/n5285 , \Reg_Bank/n5284 , \Reg_Bank/n5283 ,
         \Reg_Bank/n5282 , \Reg_Bank/n5281 , \Reg_Bank/n5280 ,
         \Reg_Bank/n5279 , \Reg_Bank/n5278 , \Reg_Bank/n5277 ,
         \Reg_Bank/n5276 , \Reg_Bank/n5275 , \Reg_Bank/n5274 ,
         \Reg_Bank/n5273 , \Reg_Bank/n5272 , \Reg_Bank/n5271 ,
         \Reg_Bank/n5270 , \Reg_Bank/n5269 , \Reg_Bank/n5268 ,
         \Reg_Bank/n5267 , \Reg_Bank/n5266 , \Reg_Bank/n5265 ,
         \Reg_Bank/n5264 , \Reg_Bank/n5263 , \Reg_Bank/n5262 ,
         \Reg_Bank/n5261 , \Reg_Bank/n5260 , \Reg_Bank/n5259 ,
         \Reg_Bank/n5258 , \Reg_Bank/n5257 , \Reg_Bank/n5256 ,
         \Reg_Bank/n5255 , \Reg_Bank/n5254 , \Reg_Bank/n5253 ,
         \Reg_Bank/n5252 , \Reg_Bank/n5251 , \Reg_Bank/n5250 ,
         \Reg_Bank/n5249 , \Reg_Bank/n5248 , \Reg_Bank/n5247 ,
         \Reg_Bank/n5246 , \Reg_Bank/n5245 , \Reg_Bank/n5244 ,
         \Reg_Bank/n5243 , \Reg_Bank/n5242 , \Reg_Bank/n5241 ,
         \Reg_Bank/n5240 , \Reg_Bank/n5239 , \Reg_Bank/n5238 ,
         \Reg_Bank/n5237 , \Reg_Bank/n5236 , \Reg_Bank/n5235 ,
         \Reg_Bank/n5234 , \Reg_Bank/n5233 , \Reg_Bank/n5232 ,
         \Reg_Bank/n5231 , \Reg_Bank/n5230 , \Reg_Bank/n5229 ,
         \Reg_Bank/n5228 , \Reg_Bank/n5227 , \Reg_Bank/n5226 ,
         \Reg_Bank/n5225 , \Reg_Bank/n5224 , \Reg_Bank/n5223 ,
         \Reg_Bank/n5222 , \Reg_Bank/n5221 , \Reg_Bank/n5220 ,
         \Reg_Bank/n5219 , \Reg_Bank/n5218 , \Reg_Bank/n5217 ,
         \Reg_Bank/n5216 , \Reg_Bank/n5215 , \Reg_Bank/n5214 ,
         \Reg_Bank/n5213 , \Reg_Bank/n5212 , \Reg_Bank/n5211 ,
         \Reg_Bank/n5210 , \Reg_Bank/n5209 , \Reg_Bank/n5208 ,
         \Reg_Bank/n5207 , \Reg_Bank/n5206 , \Reg_Bank/n5205 ,
         \Reg_Bank/n5204 , \Reg_Bank/n5203 , \Reg_Bank/n5202 ,
         \Reg_Bank/n5201 , \Reg_Bank/n5200 , \Reg_Bank/n5199 ,
         \Reg_Bank/n5198 , \Reg_Bank/n5197 , \Reg_Bank/n5196 ,
         \Reg_Bank/n5195 , \Reg_Bank/n5194 , \Reg_Bank/n5193 ,
         \Reg_Bank/n5192 , \Reg_Bank/n5191 , \Reg_Bank/n5190 ,
         \Reg_Bank/n5189 , \Reg_Bank/n5188 , \Reg_Bank/n5187 ,
         \Reg_Bank/n5186 , \Reg_Bank/n5185 , \Reg_Bank/n5184 ,
         \Reg_Bank/n5183 , \Reg_Bank/n5182 , \Reg_Bank/n5181 ,
         \Reg_Bank/n5180 , \Reg_Bank/n5179 , \Reg_Bank/n5178 ,
         \Reg_Bank/n5177 , \Reg_Bank/n5176 , \Reg_Bank/n5175 ,
         \Reg_Bank/n5174 , \Reg_Bank/n5173 , \Reg_Bank/n5172 ,
         \Reg_Bank/n5171 , \Reg_Bank/n5170 , \Reg_Bank/n5169 ,
         \Reg_Bank/n5168 , \Reg_Bank/n5167 , \Reg_Bank/n5166 ,
         \Reg_Bank/n5165 , \Reg_Bank/n5164 , \Reg_Bank/n5163 ,
         \Reg_Bank/n5162 , \Reg_Bank/n5161 , \Reg_Bank/n5160 ,
         \Reg_Bank/n5159 , \Reg_Bank/n5158 , \Reg_Bank/n5157 ,
         \Reg_Bank/n5156 , \Reg_Bank/n5155 , \Reg_Bank/n5154 ,
         \Reg_Bank/n5153 , \Reg_Bank/n5152 , \Reg_Bank/n5151 ,
         \Reg_Bank/n5150 , \Reg_Bank/n5149 , \Reg_Bank/n5148 ,
         \Reg_Bank/n5147 , \Reg_Bank/n5146 , \Reg_Bank/n5145 ,
         \Reg_Bank/n5144 , \Reg_Bank/n5143 , \Reg_Bank/n5142 ,
         \Reg_Bank/n5141 , \Reg_Bank/n5140 , \Reg_Bank/n5139 ,
         \Reg_Bank/n5138 , \Reg_Bank/n5137 , \Reg_Bank/n5136 ,
         \Reg_Bank/n5135 , \Reg_Bank/n5134 , \Reg_Bank/n5133 ,
         \Reg_Bank/n5132 , \Reg_Bank/n5131 , \Reg_Bank/n5130 ,
         \Reg_Bank/n5129 , \Reg_Bank/n5128 , \Reg_Bank/n5127 ,
         \Reg_Bank/n5126 , \Reg_Bank/n5125 , \Reg_Bank/n5124 ,
         \Reg_Bank/n5123 , \Reg_Bank/n5122 , \Reg_Bank/n5121 ,
         \Reg_Bank/n5120 , \Reg_Bank/n5119 , \Reg_Bank/n5118 ,
         \Reg_Bank/n5117 , \Reg_Bank/n5116 , \Reg_Bank/n5115 ,
         \Reg_Bank/n5114 , \Reg_Bank/n5113 , \Reg_Bank/n5112 ,
         \Reg_Bank/n5111 , \Reg_Bank/n5110 , \Reg_Bank/n5109 ,
         \Reg_Bank/n5108 , \Reg_Bank/n5107 , \Reg_Bank/n5106 ,
         \Reg_Bank/n5105 , \Reg_Bank/n5104 , \Reg_Bank/n5103 ,
         \Reg_Bank/n5102 , \Reg_Bank/n5101 , \Reg_Bank/n5100 ,
         \Reg_Bank/n5099 , \Reg_Bank/n5098 , \Reg_Bank/n5097 ,
         \Reg_Bank/n5096 , \Reg_Bank/n5095 , \Reg_Bank/n5094 ,
         \Reg_Bank/n5093 , \Reg_Bank/n5092 , \Reg_Bank/n5091 ,
         \Reg_Bank/n5090 , \Reg_Bank/n5089 , \Reg_Bank/n5088 ,
         \Reg_Bank/n5087 , \Reg_Bank/n5086 , \Reg_Bank/n5085 ,
         \Reg_Bank/n5084 , \Reg_Bank/n5083 , \Reg_Bank/n5082 ,
         \Reg_Bank/n5081 , \Reg_Bank/n5080 , \Reg_Bank/n5079 ,
         \Reg_Bank/n5078 , \Reg_Bank/n5077 , \Reg_Bank/n5076 ,
         \Reg_Bank/n5075 , \Reg_Bank/n5074 , \Reg_Bank/n5073 ,
         \Reg_Bank/n5072 , \Reg_Bank/n5071 , \Reg_Bank/n5070 ,
         \Reg_Bank/n5069 , \Reg_Bank/n5068 , \Reg_Bank/n5067 ,
         \Reg_Bank/n5066 , \Reg_Bank/n5065 , \Reg_Bank/n5064 ,
         \Reg_Bank/n5063 , \Reg_Bank/n5062 , \Reg_Bank/n5061 ,
         \Reg_Bank/n5060 , \Reg_Bank/n5059 , \Reg_Bank/n5058 ,
         \Reg_Bank/n5057 , \Reg_Bank/n5056 , \Reg_Bank/n5055 ,
         \Reg_Bank/n5054 , \Reg_Bank/n5053 , \Reg_Bank/n5052 ,
         \Reg_Bank/n5051 , \Reg_Bank/n5050 , \Reg_Bank/n5049 ,
         \Reg_Bank/n5048 , \Reg_Bank/n5047 , \Reg_Bank/n5046 ,
         \Reg_Bank/n5045 , \Reg_Bank/n5044 , \Reg_Bank/n5043 ,
         \Reg_Bank/n5042 , \Reg_Bank/n5041 , \Reg_Bank/n5040 ,
         \Reg_Bank/n5039 , \Reg_Bank/n5038 , \Reg_Bank/n5037 ,
         \Reg_Bank/n5036 , \Reg_Bank/n5035 , \Reg_Bank/n5034 ,
         \Reg_Bank/n5033 , \Reg_Bank/n5032 , \Reg_Bank/n5031 ,
         \Reg_Bank/n5030 , \Reg_Bank/n5029 , \Reg_Bank/n5028 ,
         \Reg_Bank/n5027 , \Reg_Bank/n5026 , \Reg_Bank/n5025 ,
         \Reg_Bank/n5024 , \Reg_Bank/n5023 , \Reg_Bank/n5022 ,
         \Reg_Bank/n5021 , \Reg_Bank/n5020 , \Reg_Bank/n5019 ,
         \Reg_Bank/n5018 , \Reg_Bank/n5017 , \Reg_Bank/n5016 ,
         \Reg_Bank/n5015 , \Reg_Bank/n5014 , \Reg_Bank/n5013 ,
         \Reg_Bank/n5012 , \Reg_Bank/n5011 , \Reg_Bank/n5010 ,
         \Reg_Bank/n5009 , \Reg_Bank/n5008 , \Reg_Bank/n5007 ,
         \Reg_Bank/n5006 , \Reg_Bank/n5005 , \Reg_Bank/n5004 ,
         \Reg_Bank/n5003 , \Reg_Bank/n5002 , \Reg_Bank/n5001 ,
         \Reg_Bank/n5000 , \Reg_Bank/n4999 , \Reg_Bank/n4998 ,
         \Reg_Bank/n4997 , \Reg_Bank/n4996 , \Reg_Bank/n4995 ,
         \Reg_Bank/n4994 , \Reg_Bank/n4993 , \Reg_Bank/n4992 ,
         \Reg_Bank/n4991 , \Reg_Bank/n4990 , \Reg_Bank/n4989 ,
         \Reg_Bank/n4988 , \Reg_Bank/n4987 , \Reg_Bank/n4986 ,
         \Reg_Bank/n4985 , \Reg_Bank/n4984 , \Reg_Bank/n4983 ,
         \Reg_Bank/n4982 , \Reg_Bank/n4981 , \Reg_Bank/n4980 ,
         \Reg_Bank/n4979 , \Reg_Bank/n4978 , \Reg_Bank/n4977 ,
         \Reg_Bank/n4976 , \Reg_Bank/n4975 , \Reg_Bank/n4974 ,
         \Reg_Bank/n4973 , \Reg_Bank/n4972 , \Reg_Bank/n4971 ,
         \Reg_Bank/n4970 , \Reg_Bank/n4969 , \Reg_Bank/n4968 ,
         \Reg_Bank/n4967 , \Reg_Bank/n4966 , \Reg_Bank/n4965 ,
         \Reg_Bank/n4964 , \Reg_Bank/n4963 , \Reg_Bank/n4962 ,
         \Reg_Bank/n4961 , \Reg_Bank/n4960 , \Reg_Bank/n4959 ,
         \Reg_Bank/n4958 , \Reg_Bank/n4957 , \Reg_Bank/n4956 ,
         \Reg_Bank/n4955 , \Reg_Bank/n4954 , \Reg_Bank/n4953 ,
         \Reg_Bank/n4952 , \Reg_Bank/n4951 , \Reg_Bank/n4950 ,
         \Reg_Bank/n4949 , \Reg_Bank/n4948 , \Reg_Bank/n4947 ,
         \Reg_Bank/n4946 , \Reg_Bank/n4945 , \Reg_Bank/n4944 ,
         \Reg_Bank/n4943 , \Reg_Bank/n4942 , \Reg_Bank/n4941 ,
         \Reg_Bank/n4940 , \Reg_Bank/n4939 , \Reg_Bank/n4938 ,
         \Reg_Bank/n4937 , \Reg_Bank/n4936 , \Reg_Bank/n4935 ,
         \Reg_Bank/n4934 , \Reg_Bank/n4933 , \Reg_Bank/n4932 ,
         \Reg_Bank/n4931 , \Reg_Bank/n4930 , \Reg_Bank/n4929 ,
         \Reg_Bank/n4928 , \Reg_Bank/n4927 , \Reg_Bank/n4926 ,
         \Reg_Bank/n4925 , \Reg_Bank/n4924 , \Reg_Bank/n4923 ,
         \Reg_Bank/n4922 , \Reg_Bank/n4921 , \Reg_Bank/n4920 ,
         \Reg_Bank/n4919 , \Reg_Bank/n4918 , \Reg_Bank/n4917 ,
         \Reg_Bank/n4916 , \Reg_Bank/n4915 , \Reg_Bank/n4914 ,
         \Reg_Bank/n4913 , \Reg_Bank/n4912 , \Reg_Bank/n4911 ,
         \Reg_Bank/n4910 , \Reg_Bank/n4909 , \Reg_Bank/n4908 ,
         \Reg_Bank/n4907 , \Reg_Bank/n4906 , \Reg_Bank/n4905 ,
         \Reg_Bank/n4904 , \Reg_Bank/n4903 , \Reg_Bank/n4902 ,
         \Reg_Bank/n4901 , \Reg_Bank/n4900 , \Reg_Bank/n4899 ,
         \Reg_Bank/n4898 , \Reg_Bank/n4897 , \Reg_Bank/n4896 ,
         \Reg_Bank/n4895 , \Reg_Bank/n4894 , \Reg_Bank/n4893 ,
         \Reg_Bank/n4892 , \Reg_Bank/n4891 , \Reg_Bank/n4890 ,
         \Reg_Bank/n4889 , \Reg_Bank/n4888 , \Reg_Bank/n4887 ,
         \Reg_Bank/n4886 , \Reg_Bank/n4885 , \Reg_Bank/n4884 ,
         \Reg_Bank/n4883 , \Reg_Bank/n4882 , \Reg_Bank/n4881 ,
         \Reg_Bank/n4880 , \Reg_Bank/n4879 , \Reg_Bank/n4878 ,
         \Reg_Bank/n4877 , \Reg_Bank/n4876 , \Reg_Bank/n4875 ,
         \Reg_Bank/n4874 , \Reg_Bank/n4873 , \Reg_Bank/n4872 ,
         \Reg_Bank/n4871 , \Reg_Bank/n4870 , \Reg_Bank/n4869 ,
         \Reg_Bank/n4868 , \Reg_Bank/n4867 , \Reg_Bank/n4866 ,
         \Reg_Bank/n4865 , \Reg_Bank/n4864 , \Reg_Bank/n4863 ,
         \Reg_Bank/n4862 , \Reg_Bank/n4861 , \Reg_Bank/n4860 ,
         \Reg_Bank/n4859 , \Reg_Bank/n4858 , \Reg_Bank/n4857 ,
         \Reg_Bank/n4856 , \Reg_Bank/n4855 , \Reg_Bank/n4854 ,
         \Reg_Bank/n4853 , \Reg_Bank/n4852 , \Reg_Bank/n4851 ,
         \Reg_Bank/n4850 , \Reg_Bank/n4849 , \Reg_Bank/n4848 ,
         \Reg_Bank/n4847 , \Reg_Bank/n4846 , \Reg_Bank/n4845 ,
         \Reg_Bank/n4844 , \Reg_Bank/n4843 , \Reg_Bank/n4842 ,
         \Reg_Bank/n4841 , \Reg_Bank/n4840 , \Reg_Bank/n4839 ,
         \Reg_Bank/n4838 , \Reg_Bank/n4837 , \Reg_Bank/n4836 ,
         \Reg_Bank/n4835 , \Reg_Bank/n4834 , \Reg_Bank/n4833 ,
         \Reg_Bank/n4832 , \Reg_Bank/n4831 , \Reg_Bank/n4830 ,
         \Reg_Bank/n4829 , \Reg_Bank/n4828 , \Reg_Bank/n4827 ,
         \Reg_Bank/n4826 , \Reg_Bank/n4825 , \Reg_Bank/n4824 ,
         \Reg_Bank/n4823 , \Reg_Bank/n4822 , \Reg_Bank/n4821 ,
         \Reg_Bank/n4820 , \Reg_Bank/n4819 , \Reg_Bank/n4818 ,
         \Reg_Bank/n4817 , \Reg_Bank/n4816 , \Reg_Bank/n4815 ,
         \Reg_Bank/n4814 , \Reg_Bank/n4813 , \Reg_Bank/n4812 ,
         \Reg_Bank/n4811 , \Reg_Bank/n4810 , \Reg_Bank/n4809 ,
         \Reg_Bank/n4808 , \Reg_Bank/n4807 , \Reg_Bank/n4806 ,
         \Reg_Bank/n4805 , \Reg_Bank/n4804 , \Reg_Bank/n4803 ,
         \Reg_Bank/n4802 , \Reg_Bank/n4801 , \Reg_Bank/n4800 ,
         \Reg_Bank/n4799 , \Reg_Bank/n4798 , \Reg_Bank/n4797 ,
         \Reg_Bank/n4796 , \Reg_Bank/n4795 , \Reg_Bank/n4794 ,
         \Reg_Bank/n4793 , \Reg_Bank/n4792 , \Reg_Bank/n4791 ,
         \Reg_Bank/n4790 , \Reg_Bank/n4789 , \Reg_Bank/n4788 ,
         \Reg_Bank/n4787 , \Reg_Bank/n4786 , \Reg_Bank/n4785 ,
         \Reg_Bank/n4784 , \Reg_Bank/n4783 , \Reg_Bank/n4782 ,
         \Reg_Bank/n4781 , \Reg_Bank/n4780 , \Reg_Bank/n4779 ,
         \Reg_Bank/n4778 , \Reg_Bank/n4777 , \Reg_Bank/n4776 ,
         \Reg_Bank/n4775 , \Reg_Bank/n4774 , \Reg_Bank/n4773 ,
         \Reg_Bank/n4772 , \Reg_Bank/n4771 , \Reg_Bank/n4770 ,
         \Reg_Bank/n4769 , \Reg_Bank/n4768 , \Reg_Bank/n4767 ,
         \Reg_Bank/n4766 , \Reg_Bank/n4765 , \Reg_Bank/n4764 ,
         \Reg_Bank/n4763 , \Reg_Bank/n4762 , \Reg_Bank/n4761 ,
         \Reg_Bank/n4760 , \Reg_Bank/n4759 , \Reg_Bank/n4758 ,
         \Reg_Bank/n4757 , \Reg_Bank/n4756 , \Reg_Bank/n4755 ,
         \Reg_Bank/n4754 , \Reg_Bank/n4753 , \Reg_Bank/n4752 ,
         \Reg_Bank/n4751 , \Reg_Bank/n4750 , \Reg_Bank/n4749 ,
         \Reg_Bank/n4748 , \Reg_Bank/n4747 , \Reg_Bank/n4746 ,
         \Reg_Bank/n4745 , \Reg_Bank/n4744 , \Reg_Bank/n4743 ,
         \Reg_Bank/n4742 , \Reg_Bank/n4741 , \Reg_Bank/n4740 ,
         \Reg_Bank/n4739 , \Reg_Bank/n4738 , \Reg_Bank/n4737 ,
         \Reg_Bank/n4736 , \Reg_Bank/n4735 , \Reg_Bank/n4734 ,
         \Reg_Bank/n4733 , \Reg_Bank/n4732 , \Reg_Bank/n4731 ,
         \Reg_Bank/n4730 , \Reg_Bank/n4729 , \Reg_Bank/n4728 ,
         \Reg_Bank/n4727 , \Reg_Bank/n4726 , \Reg_Bank/n4725 ,
         \Reg_Bank/n4724 , \Reg_Bank/n4723 , \Reg_Bank/n4722 ,
         \Reg_Bank/n4721 , \Reg_Bank/n4720 , \Reg_Bank/n4719 ,
         \Reg_Bank/n4718 , \Reg_Bank/n4717 , \Reg_Bank/n4716 ,
         \Reg_Bank/n4715 , \Reg_Bank/n4714 , \Reg_Bank/n4713 ,
         \Reg_Bank/n4712 , \Reg_Bank/n4711 , \Reg_Bank/n4710 ,
         \Reg_Bank/n4709 , \Reg_Bank/n4708 , \Reg_Bank/n4707 ,
         \Reg_Bank/n4706 , \Reg_Bank/n4705 , \Reg_Bank/n4704 ,
         \Reg_Bank/n4703 , \Reg_Bank/n4702 , \Reg_Bank/n4701 ,
         \Reg_Bank/n4700 , \Reg_Bank/n4699 , \Reg_Bank/n4698 ,
         \Reg_Bank/n4697 , \Reg_Bank/n4696 , \Reg_Bank/n4695 ,
         \Reg_Bank/n4694 , \Reg_Bank/n4693 , \Reg_Bank/n4692 ,
         \Reg_Bank/n4691 , \Reg_Bank/n4690 , \Reg_Bank/n4689 ,
         \Reg_Bank/n4688 , \Reg_Bank/n4687 , \Reg_Bank/n4686 ,
         \Reg_Bank/n4685 , \Reg_Bank/n4684 , \Reg_Bank/n4683 ,
         \Reg_Bank/n4682 , \Reg_Bank/n4681 , \Reg_Bank/n4680 ,
         \Reg_Bank/n4679 , \Reg_Bank/n4678 , \Reg_Bank/n4677 ,
         \Reg_Bank/n4676 , \Reg_Bank/n4675 , \Reg_Bank/n4674 ,
         \Reg_Bank/n4673 , \Reg_Bank/n4672 , \Reg_Bank/n4671 ,
         \Reg_Bank/n4670 , \Reg_Bank/n4669 , \Reg_Bank/n4668 ,
         \Reg_Bank/n4667 , \Reg_Bank/n4666 , \Reg_Bank/n4665 ,
         \Reg_Bank/n4664 , \Reg_Bank/n4663 , \Reg_Bank/n4662 ,
         \Reg_Bank/n4661 , \Reg_Bank/n4660 , \Reg_Bank/n4659 ,
         \Reg_Bank/n4658 , \Reg_Bank/n4657 , \Reg_Bank/n4656 ,
         \Reg_Bank/n4655 , \Reg_Bank/n4654 , \Reg_Bank/n4653 ,
         \Reg_Bank/n4652 , \Reg_Bank/n4651 , \Reg_Bank/n4650 ,
         \Reg_Bank/n4649 , \Reg_Bank/n4648 , \Reg_Bank/n4647 ,
         \Reg_Bank/n4646 , \Reg_Bank/n4645 , \Reg_Bank/n4644 ,
         \Reg_Bank/n4643 , \Reg_Bank/n4642 , \Reg_Bank/n4641 ,
         \Reg_Bank/n4640 , \Reg_Bank/n4639 , \Reg_Bank/n4638 ,
         \Reg_Bank/n4637 , \Reg_Bank/n4636 , \Reg_Bank/n4635 ,
         \Reg_Bank/n4634 , \Reg_Bank/n4633 , \Reg_Bank/n4632 ,
         \Reg_Bank/n4631 , \Reg_Bank/n4630 , \Reg_Bank/n4629 ,
         \Reg_Bank/n4628 , \Reg_Bank/n4627 , \Reg_Bank/n4626 ,
         \Reg_Bank/n4625 , \Reg_Bank/n4624 , \Reg_Bank/n4623 ,
         \Reg_Bank/n4622 , \Reg_Bank/n4621 , \Reg_Bank/n4620 ,
         \Reg_Bank/n4619 , \Reg_Bank/n4618 , \Reg_Bank/n4617 ,
         \Reg_Bank/n4616 , \Reg_Bank/n4615 , \Reg_Bank/n4614 ,
         \Reg_Bank/n4613 , \Reg_Bank/n4612 , \Reg_Bank/n4611 ,
         \Reg_Bank/n4610 , \Reg_Bank/n4609 , \Reg_Bank/n4608 ,
         \Reg_Bank/n4607 , \Reg_Bank/n4606 , \Reg_Bank/n4605 ,
         \Reg_Bank/n4604 , \Reg_Bank/n4603 , \Reg_Bank/n4602 ,
         \Reg_Bank/n4601 , \Reg_Bank/n4600 , \Reg_Bank/n4599 ,
         \Reg_Bank/n4598 , \Reg_Bank/n4597 , \Reg_Bank/n4596 ,
         \Reg_Bank/n4595 , \Reg_Bank/n4594 , \Reg_Bank/n4593 ,
         \Reg_Bank/n4592 , \Reg_Bank/n4591 , \Reg_Bank/n4590 ,
         \Reg_Bank/n4589 , \Reg_Bank/n4588 , \Reg_Bank/n4587 ,
         \Reg_Bank/n4586 , \Reg_Bank/n4585 , \Reg_Bank/n4584 ,
         \Reg_Bank/n4583 , \Reg_Bank/n4582 , \Reg_Bank/n4581 ,
         \Reg_Bank/n4580 , \Reg_Bank/n4579 , \Reg_Bank/n4578 ,
         \Reg_Bank/n4577 , \Reg_Bank/n4576 , \Reg_Bank/n4575 ,
         \Reg_Bank/n4574 , \Reg_Bank/n4573 , \Reg_Bank/n4572 ,
         \Reg_Bank/n4571 , \Reg_Bank/n4570 , \Reg_Bank/n4569 ,
         \Reg_Bank/n4568 , \Reg_Bank/n4567 , \Reg_Bank/n4566 ,
         \Reg_Bank/n4565 , \Reg_Bank/n4564 , \Reg_Bank/n4563 ,
         \Reg_Bank/n4562 , \Reg_Bank/n4561 , \Reg_Bank/n4560 ,
         \Reg_Bank/n4559 , \Reg_Bank/n4558 , \Reg_Bank/n4557 ,
         \Reg_Bank/n4556 , \Reg_Bank/n4555 , \Reg_Bank/n4554 ,
         \Reg_Bank/n4553 , \Reg_Bank/n4552 , \Reg_Bank/n4551 ,
         \Reg_Bank/n4550 , \Reg_Bank/n4549 , \Reg_Bank/n4548 ,
         \Reg_Bank/n4547 , \Reg_Bank/n4546 , \Reg_Bank/n4545 ,
         \Reg_Bank/n4544 , \Reg_Bank/n4543 , \Reg_Bank/n4542 ,
         \Reg_Bank/n4541 , \Reg_Bank/n4540 , \Reg_Bank/n4539 ,
         \Reg_Bank/n4538 , \Reg_Bank/n4537 , \Reg_Bank/n4536 ,
         \Reg_Bank/n4535 , \Reg_Bank/n4534 , \Reg_Bank/n4533 ,
         \Reg_Bank/n4532 , \Reg_Bank/n4531 , \Reg_Bank/n4530 ,
         \Reg_Bank/n4529 , \Reg_Bank/n4528 , \Reg_Bank/n4527 ,
         \Reg_Bank/n4526 , \Reg_Bank/n4525 , \Reg_Bank/n4524 ,
         \Reg_Bank/n4523 , \Reg_Bank/n4522 , \Reg_Bank/n4521 ,
         \Reg_Bank/n4520 , \Reg_Bank/n4519 , \Reg_Bank/n4518 ,
         \Reg_Bank/n4517 , \Reg_Bank/n4516 , \Reg_Bank/n4515 ,
         \Reg_Bank/n4514 , \Reg_Bank/n4513 , \Reg_Bank/n4512 ,
         \Reg_Bank/n4511 , \Reg_Bank/n4510 , \Reg_Bank/n4509 ,
         \Reg_Bank/n4508 , \Reg_Bank/n4507 , \Reg_Bank/n4506 ,
         \Reg_Bank/n4505 , \Reg_Bank/n4504 , \Reg_Bank/n4503 ,
         \Reg_Bank/n4502 , \Reg_Bank/n4501 , \Reg_Bank/n4500 ,
         \Reg_Bank/n4499 , \Reg_Bank/n4498 , \Reg_Bank/n4497 ,
         \Reg_Bank/n4496 , \Reg_Bank/n4495 , \Reg_Bank/n4494 ,
         \Reg_Bank/n4493 , \Reg_Bank/n4492 , \Reg_Bank/n4491 ,
         \Reg_Bank/n4490 , \Reg_Bank/n4489 , \Reg_Bank/n4488 ,
         \Reg_Bank/n4487 , \Reg_Bank/n4486 , \Reg_Bank/n4485 ,
         \Reg_Bank/n4484 , \Reg_Bank/n4483 , \Reg_Bank/n4482 ,
         \Reg_Bank/n4481 , \Reg_Bank/n4480 , \Reg_Bank/n4479 ,
         \Reg_Bank/n4478 , \Reg_Bank/n4477 , \Reg_Bank/n4476 ,
         \Reg_Bank/n4475 , \Reg_Bank/n4474 , \Reg_Bank/n4473 ,
         \Reg_Bank/n4472 , \Reg_Bank/n4471 , \Reg_Bank/n4470 ,
         \Reg_Bank/n4469 , \Reg_Bank/n4468 , \Reg_Bank/n4467 ,
         \Reg_Bank/n4466 , \Reg_Bank/n4465 , \Reg_Bank/n4464 ,
         \Reg_Bank/n4463 , \Reg_Bank/n4462 , \Reg_Bank/n4461 ,
         \Reg_Bank/n4460 , \Reg_Bank/n4459 , \Reg_Bank/n4458 ,
         \Reg_Bank/n4457 , \Reg_Bank/n4456 , \Reg_Bank/n4455 ,
         \Reg_Bank/n4454 , \Reg_Bank/n4453 , \Reg_Bank/n4452 ,
         \Reg_Bank/n4451 , \Reg_Bank/n4450 , \Reg_Bank/n4449 ,
         \Reg_Bank/n4448 , \Reg_Bank/n4447 , \Reg_Bank/n4446 ,
         \Reg_Bank/n4445 , \Reg_Bank/n4444 , \Reg_Bank/n4443 ,
         \Reg_Bank/n4442 , \Reg_Bank/n4441 , \Reg_Bank/n4440 ,
         \Reg_Bank/n4439 , \Reg_Bank/n4438 , \Reg_Bank/n4437 ,
         \Reg_Bank/n4436 , \Reg_Bank/n4435 , \Reg_Bank/n4434 ,
         \Reg_Bank/n4433 , \Reg_Bank/n4432 , \Reg_Bank/n4431 ,
         \Reg_Bank/n4430 , \Reg_Bank/n4429 , \Reg_Bank/n4428 ,
         \Reg_Bank/n4427 , \Reg_Bank/n4426 , \Reg_Bank/n4425 ,
         \Reg_Bank/n4424 , \Reg_Bank/n4423 , \Reg_Bank/n4422 ,
         \Reg_Bank/n4421 , \Reg_Bank/n4420 , \Reg_Bank/n4419 ,
         \Reg_Bank/n4418 , \Reg_Bank/n4417 , \Reg_Bank/n4416 ,
         \Reg_Bank/n4415 , \Reg_Bank/n4414 , \Reg_Bank/n4413 ,
         \Reg_Bank/n4412 , \Reg_Bank/n4411 , \Reg_Bank/n4410 ,
         \Reg_Bank/n4409 , \Reg_Bank/n4408 , \Reg_Bank/n4407 ,
         \Reg_Bank/n4406 , \Reg_Bank/n4405 , \Reg_Bank/n4404 ,
         \Reg_Bank/n4403 , \Reg_Bank/n4402 , \Reg_Bank/n4401 ,
         \Reg_Bank/n4400 , \Reg_Bank/n4399 , \Reg_Bank/n4398 ,
         \Reg_Bank/n4397 , \Reg_Bank/n4396 , \Reg_Bank/n4395 ,
         \Reg_Bank/n4394 , \Reg_Bank/n4393 , \Reg_Bank/n4392 ,
         \Reg_Bank/n4391 , \Reg_Bank/n4390 , \Reg_Bank/n4389 ,
         \Reg_Bank/n4388 , \Reg_Bank/n4387 , \Reg_Bank/n4386 ,
         \Reg_Bank/n4385 , \Reg_Bank/n4384 , \Reg_Bank/n4383 ,
         \Reg_Bank/n4382 , \Reg_Bank/n4381 , \Reg_Bank/n4380 ,
         \Reg_Bank/n4379 , \Reg_Bank/n4378 , \Reg_Bank/n4377 ,
         \Reg_Bank/n4376 , \Reg_Bank/n4375 , \Reg_Bank/n4374 ,
         \Reg_Bank/n4373 , \Reg_Bank/n4372 , \Reg_Bank/n4371 ,
         \Reg_Bank/n4370 , \Reg_Bank/n4369 , \Reg_Bank/n4368 ,
         \Reg_Bank/n4367 , \Reg_Bank/n4366 , \Reg_Bank/n4365 ,
         \Reg_Bank/n4364 , \Reg_Bank/n4363 , \Reg_Bank/n4362 ,
         \Reg_Bank/n4361 , \Reg_Bank/n4360 , \Reg_Bank/n4359 ,
         \Reg_Bank/n4358 , \Reg_Bank/n4357 , \Reg_Bank/n4356 ,
         \Reg_Bank/n4355 , \Reg_Bank/n4354 , \Reg_Bank/n4353 ,
         \Reg_Bank/n4352 , \Reg_Bank/n4351 , \Reg_Bank/n4350 ,
         \Reg_Bank/n4349 , \Reg_Bank/n4348 , \Reg_Bank/n4347 ,
         \Reg_Bank/n4346 , \Reg_Bank/n4345 , \Reg_Bank/n4344 ,
         \Reg_Bank/n4343 , \Reg_Bank/n4342 , \Reg_Bank/n4341 ,
         \Reg_Bank/n4340 , \Reg_Bank/n4339 , \Reg_Bank/n4338 ,
         \Reg_Bank/n4337 , \Reg_Bank/n4336 , \Reg_Bank/n4335 ,
         \Reg_Bank/n4334 , \Reg_Bank/n4333 , \Reg_Bank/n4332 ,
         \Reg_Bank/n4331 , \Reg_Bank/n4330 , \Reg_Bank/n4329 ,
         \Reg_Bank/n4328 , \Reg_Bank/n4327 , \Reg_Bank/n4326 ,
         \Reg_Bank/n4325 , \Reg_Bank/n4324 , \Reg_Bank/n4323 ,
         \Reg_Bank/n4322 , \Reg_Bank/n4321 , \Reg_Bank/n4320 ,
         \Reg_Bank/n4319 , \Reg_Bank/n4318 , \Reg_Bank/n4317 ,
         \Reg_Bank/n4316 , \Reg_Bank/n4315 , \Reg_Bank/n4314 ,
         \Reg_Bank/n4313 , \Reg_Bank/n4312 , \Reg_Bank/n4311 ,
         \Reg_Bank/n4310 , \Reg_Bank/n4309 , \Reg_Bank/n4308 ,
         \Reg_Bank/n4307 , \Reg_Bank/n4306 , \Reg_Bank/n4305 ,
         \Reg_Bank/n4304 , \Reg_Bank/n4303 , \Reg_Bank/n4302 ,
         \Reg_Bank/n4301 , \Reg_Bank/n4300 , \Reg_Bank/n4299 ,
         \Reg_Bank/n4298 , \Reg_Bank/n4297 , \Reg_Bank/n4296 ,
         \Reg_Bank/n4295 , \Reg_Bank/n4294 , \Reg_Bank/n4293 ,
         \Reg_Bank/n4292 , \Reg_Bank/n4291 , \Reg_Bank/n4290 ,
         \Reg_Bank/n4289 , \Reg_Bank/n4288 , \Reg_Bank/n4287 ,
         \Reg_Bank/n4286 , \Reg_Bank/n4285 , \Reg_Bank/n4284 ,
         \Reg_Bank/n4283 , \Reg_Bank/n4282 , \Reg_Bank/n4281 ,
         \Reg_Bank/n4280 , \Reg_Bank/n4279 , \Reg_Bank/n4278 ,
         \Reg_Bank/n4277 , \Reg_Bank/n4276 , \Reg_Bank/n4275 ,
         \Reg_Bank/n4274 , \Reg_Bank/n4273 , \Reg_Bank/n4272 ,
         \Reg_Bank/n4271 , \Reg_Bank/n4270 , \Reg_Bank/n4269 ,
         \Reg_Bank/n4268 , \Reg_Bank/n4267 , \Reg_Bank/n4266 ,
         \Reg_Bank/n4265 , \Reg_Bank/n4264 , \Reg_Bank/n4263 ,
         \Reg_Bank/n4262 , \Reg_Bank/n4261 , \Reg_Bank/n4260 ,
         \Reg_Bank/n4259 , \Reg_Bank/n4258 , \Reg_Bank/n4257 ,
         \Reg_Bank/n4256 , \Reg_Bank/n4255 , \Reg_Bank/n4254 ,
         \Reg_Bank/n4253 , \Reg_Bank/n4252 , \Reg_Bank/n4251 ,
         \Reg_Bank/n4250 , \Reg_Bank/n4249 , \Reg_Bank/n4248 ,
         \Reg_Bank/n4247 , \Reg_Bank/n4246 , \Reg_Bank/n4245 ,
         \Reg_Bank/n4244 , \Reg_Bank/n4243 , \Reg_Bank/n4242 ,
         \Reg_Bank/n4241 , \Reg_Bank/n4240 , \Reg_Bank/n4239 ,
         \Reg_Bank/n4238 , \Reg_Bank/n4237 , \Reg_Bank/n4236 ,
         \Reg_Bank/n4235 , \Reg_Bank/n4234 , \Reg_Bank/n4233 ,
         \Reg_Bank/n4232 , \Reg_Bank/n4231 , \Reg_Bank/n4230 ,
         \Reg_Bank/n4229 , \Reg_Bank/n4228 , \Reg_Bank/n4227 ,
         \Reg_Bank/n4226 , \Reg_Bank/n4225 , \Reg_Bank/n4224 ,
         \Reg_Bank/n4223 , \Reg_Bank/n4222 , \Reg_Bank/n4221 ,
         \Reg_Bank/n4220 , \Reg_Bank/n4219 , \Reg_Bank/n4218 ,
         \Reg_Bank/n4217 , \Reg_Bank/n4216 , \Reg_Bank/n4215 ,
         \Reg_Bank/n4214 , \Reg_Bank/n4213 , \Reg_Bank/n4212 ,
         \Reg_Bank/n4211 , \Reg_Bank/n4210 , \Reg_Bank/n4209 ,
         \Reg_Bank/n4208 , \Reg_Bank/n4207 , \Reg_Bank/n4206 ,
         \Reg_Bank/n4205 , \Reg_Bank/n4204 , \Reg_Bank/n4203 ,
         \Reg_Bank/n4202 , \Reg_Bank/n4201 , \Reg_Bank/n4200 ,
         \Reg_Bank/n4199 , \Reg_Bank/n4198 , \Reg_Bank/n4197 ,
         \Reg_Bank/n4196 , \Reg_Bank/n4195 , \Reg_Bank/n4194 ,
         \Reg_Bank/n4193 , \Reg_Bank/n4192 , \Reg_Bank/n4191 ,
         \Reg_Bank/n4190 , \Reg_Bank/n4189 , \Reg_Bank/n4188 ,
         \Reg_Bank/n4187 , \Reg_Bank/n4186 , \Reg_Bank/n4185 ,
         \Reg_Bank/n4184 , \Reg_Bank/n4183 , \Reg_Bank/n4182 ,
         \Reg_Bank/n4181 , \Reg_Bank/n4180 , \Reg_Bank/n4179 ,
         \Reg_Bank/n4178 , \Reg_Bank/n4177 , \Reg_Bank/n4176 ,
         \Reg_Bank/n4175 , \Reg_Bank/n4174 , \Reg_Bank/n4173 ,
         \Reg_Bank/n4172 , \Reg_Bank/n4171 , \Reg_Bank/n4170 ,
         \Reg_Bank/n4169 , \Reg_Bank/n4168 , \Reg_Bank/n4167 ,
         \Reg_Bank/n4166 , \Reg_Bank/n4165 , \Reg_Bank/n4164 ,
         \Reg_Bank/n4163 , \Reg_Bank/n4162 , \Reg_Bank/n4161 ,
         \Reg_Bank/n4160 , \Reg_Bank/n4159 , \Reg_Bank/n4158 ,
         \Reg_Bank/n4157 , \Reg_Bank/n4156 , \Reg_Bank/n4155 ,
         \Reg_Bank/n4154 , \Reg_Bank/n4153 , \Reg_Bank/n4152 ,
         \Reg_Bank/n4151 , \Reg_Bank/n4150 , \Reg_Bank/n4149 ,
         \Reg_Bank/n4148 , \Reg_Bank/n4147 , \Reg_Bank/n4146 ,
         \Reg_Bank/n4145 , \Reg_Bank/n4144 , \Reg_Bank/n4143 ,
         \Reg_Bank/n4142 , \Reg_Bank/n4141 , \Reg_Bank/n4140 ,
         \Reg_Bank/n4139 , \Reg_Bank/n4138 , \Reg_Bank/n4137 ,
         \Reg_Bank/n4136 , \Reg_Bank/n4135 , \Reg_Bank/n4134 ,
         \Reg_Bank/n4133 , \Reg_Bank/n4132 , \Reg_Bank/n4131 ,
         \Reg_Bank/n4130 , \Reg_Bank/n4129 , \Reg_Bank/n4128 ,
         \Reg_Bank/n4127 , \Reg_Bank/n4126 , \Reg_Bank/n4125 ,
         \Reg_Bank/n4124 , \Reg_Bank/n4123 , \Reg_Bank/n4122 ,
         \Reg_Bank/n4121 , \Reg_Bank/n4120 , \Reg_Bank/n4119 ,
         \Reg_Bank/n4118 , \Reg_Bank/n4117 , \Reg_Bank/n4116 ,
         \Reg_Bank/n4115 , \Reg_Bank/n4114 , \Reg_Bank/n4113 ,
         \Reg_Bank/n4112 , \Reg_Bank/n4111 , \Reg_Bank/n4110 ,
         \Reg_Bank/n4109 , \Reg_Bank/n4108 , \Reg_Bank/n4107 ,
         \Reg_Bank/n4106 , \Reg_Bank/n4105 , \Reg_Bank/n4104 ,
         \Reg_Bank/n4103 , \Reg_Bank/n4102 , \Reg_Bank/n4101 ,
         \Reg_Bank/n4100 , \Reg_Bank/n4099 , \Reg_Bank/n4098 ,
         \Reg_Bank/n4097 , \Reg_Bank/n4096 , \Reg_Bank/n4095 ,
         \Reg_Bank/n4094 , \Reg_Bank/n4093 , \Reg_Bank/n4092 ,
         \Reg_Bank/n4091 , \Reg_Bank/n4090 , \Reg_Bank/n4089 ,
         \Reg_Bank/n4088 , \Reg_Bank/n4087 , \Reg_Bank/n4086 ,
         \Reg_Bank/n4085 , \Reg_Bank/n4084 , \Reg_Bank/n4083 ,
         \Reg_Bank/n4082 , \Reg_Bank/n4081 , \Reg_Bank/n4080 ,
         \Reg_Bank/n4079 , \Reg_Bank/n4078 , \Reg_Bank/n4077 ,
         \Reg_Bank/n4076 , \Reg_Bank/n4075 , \Reg_Bank/n4074 ,
         \Reg_Bank/n4073 , \Reg_Bank/n4072 , \Reg_Bank/n4071 ,
         \Reg_Bank/n4070 , \Reg_Bank/n4069 , \Reg_Bank/n4068 ,
         \Reg_Bank/n4067 , \Reg_Bank/n4066 , \Reg_Bank/n4065 ,
         \Reg_Bank/n4064 , \Reg_Bank/n4063 , \Reg_Bank/n4062 ,
         \Reg_Bank/n4061 , \Reg_Bank/n4060 , \Reg_Bank/n4059 ,
         \Reg_Bank/n4058 , \Reg_Bank/n4057 , \Reg_Bank/n4056 ,
         \Reg_Bank/n4055 , \Reg_Bank/n4054 , \Reg_Bank/n4053 ,
         \Reg_Bank/n4052 , \Reg_Bank/n4051 , \Reg_Bank/n4050 ,
         \Reg_Bank/n4049 , \Reg_Bank/n4048 , \Reg_Bank/n4047 ,
         \Reg_Bank/n4046 , \Reg_Bank/n4045 , \Reg_Bank/n4044 ,
         \Reg_Bank/n4043 , \Reg_Bank/n4042 , \Reg_Bank/n4041 ,
         \Reg_Bank/n4040 , \Reg_Bank/n4039 , \Reg_Bank/n4038 ,
         \Reg_Bank/n4037 , \Reg_Bank/n4036 , \Reg_Bank/n4035 ,
         \Reg_Bank/n4034 , \Reg_Bank/n4033 , \Reg_Bank/n4032 ,
         \Reg_Bank/n4031 , \Reg_Bank/n4030 , \Reg_Bank/n4029 ,
         \Reg_Bank/n4028 , \Reg_Bank/n4027 , \Reg_Bank/n4026 ,
         \Reg_Bank/n4025 , \Reg_Bank/n4024 , \Reg_Bank/n4023 ,
         \Reg_Bank/n4022 , \Reg_Bank/n4021 , \Reg_Bank/n4020 ,
         \Reg_Bank/n4019 , \Reg_Bank/n4018 , \Reg_Bank/n4017 ,
         \Reg_Bank/n4016 , \Reg_Bank/n4015 , \Reg_Bank/n4014 ,
         \Reg_Bank/n4013 , \Reg_Bank/n4012 , \Reg_Bank/n4011 ,
         \Reg_Bank/n4010 , \Reg_Bank/n4009 , \Reg_Bank/n4008 ,
         \Reg_Bank/n4007 , \Reg_Bank/n4006 , \Reg_Bank/n4005 ,
         \Reg_Bank/n4004 , \Reg_Bank/n4003 , \Reg_Bank/n4002 ,
         \Reg_Bank/n4001 , \Reg_Bank/n4000 , \Reg_Bank/n3999 ,
         \Reg_Bank/n3998 , \Reg_Bank/n3997 , \Reg_Bank/n3996 ,
         \Reg_Bank/n3995 , \Reg_Bank/n3994 , \Reg_Bank/n3993 ,
         \Reg_Bank/n3992 , \Reg_Bank/n3991 , \Reg_Bank/n3990 ,
         \Reg_Bank/n3989 , \Reg_Bank/n3988 , \Reg_Bank/n3987 ,
         \Reg_Bank/n3986 , \Reg_Bank/n3985 , \Reg_Bank/n3984 ,
         \Reg_Bank/n3983 , \Reg_Bank/n3982 , \Reg_Bank/n3981 ,
         \Reg_Bank/n3980 , \Reg_Bank/n3979 , \Reg_Bank/n3978 ,
         \Reg_Bank/n3977 , \Reg_Bank/n3976 , \Reg_Bank/n3975 ,
         \Reg_Bank/n3974 , \Reg_Bank/n3973 , \Reg_Bank/n3972 ,
         \Reg_Bank/n3971 , \Reg_Bank/n3970 , \Reg_Bank/n3969 ,
         \Reg_Bank/n3968 , \Reg_Bank/n3967 , \Reg_Bank/n3966 ,
         \Reg_Bank/n3965 , \Reg_Bank/n3964 , \Reg_Bank/n3963 ,
         \Reg_Bank/n3962 , \Reg_Bank/n3961 , \Reg_Bank/n3960 ,
         \Reg_Bank/n3959 , \Reg_Bank/n3958 , \Reg_Bank/n3957 ,
         \Reg_Bank/n3956 , \Reg_Bank/n3955 , \Reg_Bank/n3954 ,
         \Reg_Bank/n3953 , \Reg_Bank/n3952 , \Reg_Bank/n3951 ,
         \Reg_Bank/n3950 , \Reg_Bank/n3949 , \Reg_Bank/n3948 ,
         \Reg_Bank/n3947 , \Reg_Bank/n3946 , \Reg_Bank/n3945 ,
         \Reg_Bank/n3944 , \Reg_Bank/n3943 , \Reg_Bank/n3942 ,
         \Reg_Bank/n3941 , \Reg_Bank/n3940 , \Reg_Bank/n3939 ,
         \Reg_Bank/n3938 , \Reg_Bank/n3937 , \Reg_Bank/n3936 ,
         \Reg_Bank/n3935 , \Reg_Bank/n3934 , \Reg_Bank/n3933 ,
         \Reg_Bank/n3932 , \Reg_Bank/n3931 , \Reg_Bank/n3930 ,
         \Reg_Bank/n3929 , \Reg_Bank/n3928 , \Reg_Bank/n3927 ,
         \Reg_Bank/n3926 , \Reg_Bank/n3925 , \Reg_Bank/n3924 ,
         \Reg_Bank/n3923 , \Reg_Bank/n3922 , \Reg_Bank/n3921 ,
         \Reg_Bank/n3920 , \Reg_Bank/n3919 , \Reg_Bank/n3918 ,
         \Reg_Bank/n3917 , \Reg_Bank/n3916 , \Reg_Bank/n3915 ,
         \Reg_Bank/n3914 , \Reg_Bank/n3913 , \Reg_Bank/n3912 ,
         \Reg_Bank/n3911 , \Reg_Bank/n3910 , \Reg_Bank/n3909 ,
         \Reg_Bank/n3908 , \Reg_Bank/n3907 , \Reg_Bank/n3906 ,
         \Reg_Bank/n3905 , \Reg_Bank/n3904 , \Reg_Bank/n3903 ,
         \Reg_Bank/n3902 , \Reg_Bank/n3901 , \Reg_Bank/n3900 ,
         \Reg_Bank/n3899 , \Reg_Bank/n3898 , \Reg_Bank/n3897 ,
         \Reg_Bank/n3896 , \Reg_Bank/n3895 , \Reg_Bank/n3894 ,
         \Reg_Bank/n3893 , \Reg_Bank/n3892 , \Reg_Bank/n3891 ,
         \Reg_Bank/n3890 , \Reg_Bank/n3889 , \Reg_Bank/n3888 ,
         \Reg_Bank/n3887 , \Reg_Bank/n3886 , \Reg_Bank/n3885 ,
         \Reg_Bank/n3884 , \Reg_Bank/n3883 , \Reg_Bank/n3882 ,
         \Reg_Bank/n3881 , \Reg_Bank/n3880 , \Reg_Bank/n3879 ,
         \Reg_Bank/n3878 , \Reg_Bank/n3877 , \Reg_Bank/n3876 ,
         \Reg_Bank/n3875 , \Reg_Bank/n3874 , \Reg_Bank/n3873 ,
         \Reg_Bank/n3872 , \Reg_Bank/n3871 , \Reg_Bank/n3870 ,
         \Reg_Bank/n3869 , \Reg_Bank/n3868 , \Reg_Bank/n3867 ,
         \Reg_Bank/n3866 , \Reg_Bank/n3865 , \Reg_Bank/n3864 ,
         \Reg_Bank/n3863 , \Reg_Bank/n3862 , \Reg_Bank/n3861 ,
         \Reg_Bank/n3860 , \Reg_Bank/n3859 , \Reg_Bank/n3858 ,
         \Reg_Bank/n3857 , \Reg_Bank/n3856 , \Reg_Bank/n3855 ,
         \Reg_Bank/n3854 , \Reg_Bank/n3853 , \Reg_Bank/n3852 ,
         \Reg_Bank/n3851 , \Reg_Bank/n3850 , \Reg_Bank/n3849 ,
         \Reg_Bank/n3848 , \Reg_Bank/n3847 , \Reg_Bank/n3846 ,
         \Reg_Bank/n3845 , \Reg_Bank/n3844 , \Reg_Bank/n3843 ,
         \Reg_Bank/n3842 , \Reg_Bank/n3841 , \Reg_Bank/n3840 ,
         \Reg_Bank/n3839 , \Reg_Bank/n3838 , \Reg_Bank/n3837 ,
         \Reg_Bank/n3836 , \Reg_Bank/n3835 , \Reg_Bank/n3834 ,
         \Reg_Bank/n3833 , \Reg_Bank/n3832 , \Reg_Bank/n3831 ,
         \Reg_Bank/n3830 , \Reg_Bank/n3829 , \Reg_Bank/n3828 ,
         \Reg_Bank/n3827 , \Reg_Bank/n3826 , \Reg_Bank/n3825 ,
         \Reg_Bank/n3824 , \Reg_Bank/n3823 , \Reg_Bank/n3822 ,
         \Reg_Bank/n3821 , \Reg_Bank/n3820 , \Reg_Bank/n3819 ,
         \Reg_Bank/n3818 , \Reg_Bank/n3817 , \Reg_Bank/n3816 ,
         \Reg_Bank/n3815 , \Reg_Bank/n3814 , \Reg_Bank/n3813 ,
         \Reg_Bank/n3812 , \Reg_Bank/n3811 , \Reg_Bank/n3810 ,
         \Reg_Bank/n3809 , \Reg_Bank/n3808 , \Reg_Bank/n3807 ,
         \Reg_Bank/n3806 , \Reg_Bank/n3805 , \Reg_Bank/n3804 ,
         \Reg_Bank/n3803 , \Reg_Bank/n3802 , \Reg_Bank/n3801 ,
         \Reg_Bank/n3800 , \Reg_Bank/n3799 , \Reg_Bank/n3798 ,
         \Reg_Bank/n3797 , \Reg_Bank/n3796 , \Reg_Bank/n3795 ,
         \Reg_Bank/n3794 , \Reg_Bank/n3793 , \Reg_Bank/n3792 ,
         \Reg_Bank/n3791 , \Reg_Bank/n3790 , \Reg_Bank/n3789 ,
         \Reg_Bank/n3788 , \Reg_Bank/n3787 , \Reg_Bank/n3786 ,
         \Reg_Bank/n3785 , \Reg_Bank/n3784 , \Reg_Bank/n3783 ,
         \Reg_Bank/n3782 , \Reg_Bank/n3781 , \Reg_Bank/n3780 ,
         \Reg_Bank/n3779 , \Reg_Bank/n3778 , \Reg_Bank/n3777 ,
         \Reg_Bank/n3776 , \Reg_Bank/n3775 , \Reg_Bank/n3774 ,
         \Reg_Bank/n3773 , \Reg_Bank/n3772 , \Reg_Bank/n3771 ,
         \Reg_Bank/n3770 , \Reg_Bank/n3769 , \Reg_Bank/n3768 ,
         \Reg_Bank/n3767 , \Reg_Bank/n3766 , \Reg_Bank/n3765 ,
         \Reg_Bank/n3764 , \Reg_Bank/n3763 , \Reg_Bank/n3762 ,
         \Reg_Bank/n3761 , \Reg_Bank/n3760 , \Reg_Bank/n3759 ,
         \Reg_Bank/n3758 , \Reg_Bank/n3757 , \Reg_Bank/n3756 ,
         \Reg_Bank/n3755 , \Reg_Bank/n3754 , \Reg_Bank/n3753 ,
         \Reg_Bank/n3752 , \Reg_Bank/n3751 , \Reg_Bank/n3750 ,
         \Reg_Bank/n3749 , \Reg_Bank/n3748 , \Reg_Bank/n3747 ,
         \Reg_Bank/n3746 , \Reg_Bank/n3745 , \Reg_Bank/n3744 ,
         \Reg_Bank/n3743 , \Reg_Bank/n3742 , \Reg_Bank/n3741 ,
         \Reg_Bank/n3740 , \Reg_Bank/n3739 , \Reg_Bank/n3738 ,
         \Reg_Bank/n3737 , \Reg_Bank/n3736 , \Reg_Bank/n3735 ,
         \Reg_Bank/n3734 , \Reg_Bank/n3733 , \Reg_Bank/n3732 ,
         \Reg_Bank/n3731 , \Reg_Bank/n3730 , \Reg_Bank/n3729 ,
         \Reg_Bank/n3728 , \Reg_Bank/n3727 , \Reg_Bank/n3726 ,
         \Reg_Bank/n3725 , \Reg_Bank/n3724 , \Reg_Bank/n3723 ,
         \Reg_Bank/n3722 , \Reg_Bank/n3721 , \Reg_Bank/n3720 ,
         \Reg_Bank/n3719 , \Reg_Bank/n3718 , \Reg_Bank/n3717 ,
         \Reg_Bank/n3716 , \Reg_Bank/n3715 , \Reg_Bank/n3714 ,
         \Reg_Bank/n3713 , \Reg_Bank/n3712 , \Reg_Bank/n3711 ,
         \Reg_Bank/n3710 , \Reg_Bank/n3709 , \Reg_Bank/n3708 ,
         \Reg_Bank/n3707 , \Reg_Bank/n3706 , \Reg_Bank/n3705 ,
         \Reg_Bank/n3704 , \Reg_Bank/n3703 , \Reg_Bank/n3702 ,
         \Reg_Bank/n3701 , \Reg_Bank/n3700 , \Reg_Bank/n3699 ,
         \Reg_Bank/n3698 , \Reg_Bank/n3697 , \Reg_Bank/n3696 ,
         \Reg_Bank/n3695 , \Reg_Bank/n3694 , \Reg_Bank/n3693 ,
         \Reg_Bank/n3692 , \Reg_Bank/n3691 , \Reg_Bank/n3690 ,
         \Reg_Bank/n3689 , \Reg_Bank/n3688 , \Reg_Bank/n3687 ,
         \Reg_Bank/n3686 , \Reg_Bank/n3685 , \Reg_Bank/n3684 ,
         \Reg_Bank/n3683 , \Reg_Bank/n3682 , \Reg_Bank/n3681 ,
         \Reg_Bank/n3680 , \Reg_Bank/n3679 , \Reg_Bank/n3678 ,
         \Reg_Bank/n3677 , \Reg_Bank/n3676 , \Reg_Bank/n3675 ,
         \Reg_Bank/n3674 , \Reg_Bank/n3673 , \Reg_Bank/n3672 ,
         \Reg_Bank/n3671 , \Reg_Bank/n3670 , \Reg_Bank/n3669 ,
         \Reg_Bank/n3668 , \Reg_Bank/n3667 , \Reg_Bank/n3666 ,
         \Reg_Bank/n3665 , \Reg_Bank/n3664 , \Reg_Bank/n3663 ,
         \Reg_Bank/n3662 , \Reg_Bank/n3661 , \Reg_Bank/n3660 ,
         \Reg_Bank/n3659 , \Reg_Bank/n3658 , \Reg_Bank/n3657 ,
         \Reg_Bank/n3656 , \Reg_Bank/n3655 , \Reg_Bank/n3654 ,
         \Reg_Bank/n3653 , \Reg_Bank/n3652 , \Reg_Bank/n3651 ,
         \Reg_Bank/n3650 , \Reg_Bank/n3649 , \Reg_Bank/n3648 ,
         \Reg_Bank/n3647 , \Reg_Bank/n3646 , \Reg_Bank/n3645 ,
         \Reg_Bank/n3644 , \Reg_Bank/n3643 , \Reg_Bank/n3642 ,
         \Reg_Bank/n3641 , \Reg_Bank/n3640 , \Reg_Bank/n3639 ,
         \Reg_Bank/n3638 , \Reg_Bank/n3637 , \Reg_Bank/n3636 ,
         \Reg_Bank/n3635 , \Reg_Bank/n3634 , \Reg_Bank/n3633 ,
         \Reg_Bank/n3632 , \Reg_Bank/n3631 , \Reg_Bank/n3630 ,
         \Reg_Bank/n3629 , \Reg_Bank/n3628 , \Reg_Bank/n3627 ,
         \Reg_Bank/n3626 , \Reg_Bank/n3625 , \Reg_Bank/n3624 ,
         \Reg_Bank/n3623 , \Reg_Bank/n3622 , \Reg_Bank/n3621 ,
         \Reg_Bank/n3620 , \Reg_Bank/n3619 , \Reg_Bank/n3618 ,
         \Reg_Bank/n3617 , \Reg_Bank/n3616 , \Reg_Bank/n3615 ,
         \Reg_Bank/n3614 , \Reg_Bank/n3613 , \Reg_Bank/n3612 ,
         \Reg_Bank/n3611 , \Reg_Bank/n3610 , \Reg_Bank/n3609 ,
         \Reg_Bank/n3608 , \Reg_Bank/n3607 , \Reg_Bank/n3606 ,
         \Reg_Bank/n3605 , \Reg_Bank/n3604 , \Reg_Bank/n3603 ,
         \Reg_Bank/n3602 , \Reg_Bank/n3601 , \Reg_Bank/n3600 ,
         \Reg_Bank/n3599 , \Reg_Bank/n3598 , \Reg_Bank/n3597 ,
         \Reg_Bank/n3596 , \Reg_Bank/n3595 , \Reg_Bank/n3594 ,
         \Reg_Bank/n3593 , \Reg_Bank/n3592 , \Reg_Bank/n3591 ,
         \Reg_Bank/n3590 , \Reg_Bank/n3589 , \Reg_Bank/n3588 ,
         \Reg_Bank/n3587 , \Reg_Bank/n3586 , \Reg_Bank/n3585 ,
         \Reg_Bank/n3584 , \Reg_Bank/n3583 , \Reg_Bank/n3582 ,
         \Reg_Bank/n3581 , \Reg_Bank/n3580 , \Reg_Bank/n3579 ,
         \Reg_Bank/n3578 , \Reg_Bank/n3577 , \Reg_Bank/n3576 ,
         \Reg_Bank/n3575 , \Reg_Bank/n3574 , \Reg_Bank/n3573 ,
         \Reg_Bank/n3572 , \Reg_Bank/n3571 , \Reg_Bank/n3570 ,
         \Reg_Bank/n3569 , \Reg_Bank/n3568 , \Reg_Bank/n3567 ,
         \Reg_Bank/n3566 , \Reg_Bank/n3565 , \Reg_Bank/n3564 ,
         \Reg_Bank/n3563 , \Reg_Bank/n3562 , \Reg_Bank/n3561 ,
         \Reg_Bank/n3560 , \Reg_Bank/n3559 , \Reg_Bank/n3558 ,
         \Reg_Bank/n3557 , \Reg_Bank/n3556 , \Reg_Bank/n3555 ,
         \Reg_Bank/n3554 , \Reg_Bank/n3553 , \Reg_Bank/n3552 ,
         \Reg_Bank/n3551 , \Reg_Bank/n3550 , \Reg_Bank/n3549 ,
         \Reg_Bank/n3548 , \Reg_Bank/n3547 , \Reg_Bank/n3546 ,
         \Reg_Bank/n3545 , \Reg_Bank/n3544 , \Reg_Bank/n3543 ,
         \Reg_Bank/n3542 , \Reg_Bank/n3541 , \Reg_Bank/n3540 ,
         \Reg_Bank/n3539 , \Reg_Bank/n3538 , \Reg_Bank/n3537 ,
         \Reg_Bank/n3536 , \Reg_Bank/n3535 , \Reg_Bank/n3534 ,
         \Reg_Bank/n3533 , \Reg_Bank/n3532 , \Reg_Bank/n3531 ,
         \Reg_Bank/n3530 , \Reg_Bank/n3529 , \Reg_Bank/n3528 ,
         \Reg_Bank/n3527 , \Reg_Bank/n3526 , \Reg_Bank/n3525 ,
         \Reg_Bank/n3524 , \Reg_Bank/n3523 , \Reg_Bank/n3522 ,
         \Reg_Bank/n3521 , \Reg_Bank/n3520 , \Reg_Bank/n3519 ,
         \Reg_Bank/n3518 , \Reg_Bank/n3517 , \Reg_Bank/n3516 ,
         \Reg_Bank/n3515 , \Reg_Bank/n3514 , \Reg_Bank/n3513 ,
         \Reg_Bank/n3512 , \Reg_Bank/n3511 , \Reg_Bank/n3510 ,
         \Reg_Bank/n3509 , \Reg_Bank/n3508 , \Reg_Bank/n3507 ,
         \Reg_Bank/n3506 , \Reg_Bank/n3505 , \Reg_Bank/n3504 ,
         \Reg_Bank/n3503 , \Reg_Bank/n3502 , \Reg_Bank/n3501 ,
         \Reg_Bank/n3500 , \Reg_Bank/n3499 , \Reg_Bank/n3498 ,
         \Reg_Bank/n3497 , \Reg_Bank/n3496 , \Reg_Bank/n3495 ,
         \Reg_Bank/n3494 , \Reg_Bank/n3493 , \Reg_Bank/n3492 ,
         \Reg_Bank/n3491 , \Reg_Bank/n3490 , \Reg_Bank/n3489 ,
         \Reg_Bank/n3488 , \Reg_Bank/n3487 , \Reg_Bank/n3486 ,
         \Reg_Bank/n3485 , \Reg_Bank/n3484 , \Reg_Bank/n3483 ,
         \Reg_Bank/n3482 , \Reg_Bank/n3481 , \Reg_Bank/n3480 ,
         \Reg_Bank/n3479 , \Reg_Bank/n3478 , \Reg_Bank/n3477 ,
         \Reg_Bank/n3476 , \Reg_Bank/n3475 , \Reg_Bank/n3474 ,
         \Reg_Bank/n3473 , \Reg_Bank/n3472 , \Reg_Bank/n3471 ,
         \Reg_Bank/n3470 , \Reg_Bank/n3469 , \Reg_Bank/n3468 ,
         \Reg_Bank/n3467 , \Reg_Bank/n3466 , \Reg_Bank/n3465 ,
         \Reg_Bank/n3464 , \Reg_Bank/n3463 , \Reg_Bank/n3462 ,
         \Reg_Bank/n3461 , \Reg_Bank/n3460 , \Reg_Bank/n3459 ,
         \Reg_Bank/n3458 , \Reg_Bank/n3457 , \Reg_Bank/n3456 ,
         \Reg_Bank/n3455 , \Reg_Bank/n3454 , \Reg_Bank/n3453 ,
         \Reg_Bank/n3452 , \Reg_Bank/n3451 , \Reg_Bank/n3450 ,
         \Reg_Bank/n3449 , \Reg_Bank/n3448 , \Reg_Bank/n3447 ,
         \Reg_Bank/n3446 , \Reg_Bank/n3445 , \Reg_Bank/n3444 ,
         \Reg_Bank/n3443 , \Reg_Bank/n3442 , \Reg_Bank/n3441 ,
         \Reg_Bank/n3440 , \Reg_Bank/n3439 , \Reg_Bank/n3438 ,
         \Reg_Bank/n3437 , \Reg_Bank/n3436 , \Reg_Bank/n3435 ,
         \Reg_Bank/n3434 , \Reg_Bank/n3433 , \Reg_Bank/n3432 ,
         \Reg_Bank/n3431 , \Reg_Bank/n3430 , \Reg_Bank/n3429 ,
         \Reg_Bank/n3428 , \Reg_Bank/n3427 , \Reg_Bank/n3426 ,
         \Reg_Bank/n3425 , \Reg_Bank/n3424 , \Reg_Bank/n3423 ,
         \Reg_Bank/n3422 , \Reg_Bank/n3421 , \Reg_Bank/n3420 ,
         \Reg_Bank/n3419 , \Reg_Bank/n3418 , \Reg_Bank/n3417 ,
         \Reg_Bank/n3416 , \Reg_Bank/n3415 , \Reg_Bank/n3414 ,
         \Reg_Bank/n3413 , \Reg_Bank/n3412 , \Reg_Bank/n3411 ,
         \Reg_Bank/n3410 , \Reg_Bank/n3409 , \Reg_Bank/n3408 ,
         \Reg_Bank/n3407 , \Reg_Bank/n3406 , \Reg_Bank/n3405 ,
         \Reg_Bank/n3404 , \Reg_Bank/n3403 , \Reg_Bank/n3402 ,
         \Reg_Bank/n3401 , \Reg_Bank/n3400 , \Reg_Bank/n3399 ,
         \Reg_Bank/n3398 , \Reg_Bank/n3397 , \Reg_Bank/n3396 ,
         \Reg_Bank/n3395 , \Reg_Bank/n3394 , \Reg_Bank/n3393 ,
         \Reg_Bank/n3392 , \Reg_Bank/n3391 , \Reg_Bank/n3390 ,
         \Reg_Bank/n3389 , \Reg_Bank/n3388 , \Reg_Bank/n3387 ,
         \Reg_Bank/n3386 , \Reg_Bank/n3385 , \Reg_Bank/n3384 ,
         \Reg_Bank/n3383 , \Reg_Bank/n3382 , \Reg_Bank/n3381 ,
         \Reg_Bank/n3380 , \Reg_Bank/n3379 , \Reg_Bank/n3378 ,
         \Reg_Bank/n3377 , \Reg_Bank/n3376 , \Reg_Bank/n3375 ,
         \Reg_Bank/n3374 , \Reg_Bank/n3373 , \Reg_Bank/n3372 ,
         \Reg_Bank/n3371 , \Reg_Bank/n3370 , \Reg_Bank/n3369 ,
         \Reg_Bank/n3368 , \Reg_Bank/n3367 , \Reg_Bank/n3366 ,
         \Reg_Bank/n3365 , \Reg_Bank/n3364 , \Reg_Bank/n3363 ,
         \Reg_Bank/n3362 , \Reg_Bank/n3361 , \Reg_Bank/n3360 ,
         \Reg_Bank/n3359 , \Reg_Bank/n3358 , \Reg_Bank/n3357 ,
         \Reg_Bank/n3356 , \Reg_Bank/n3355 , \Reg_Bank/n3354 ,
         \Reg_Bank/n3353 , \Reg_Bank/n3352 , \Reg_Bank/n3351 ,
         \Reg_Bank/n3350 , \Reg_Bank/n3349 , \Reg_Bank/n3348 ,
         \Reg_Bank/n3347 , \Reg_Bank/n3346 , \Reg_Bank/n3345 ,
         \Reg_Bank/n3344 , \Reg_Bank/n3343 , \Reg_Bank/n3342 ,
         \Reg_Bank/n3341 , \Reg_Bank/n3340 , \Reg_Bank/n3339 ,
         \Reg_Bank/n3338 , \Reg_Bank/n3337 , \Reg_Bank/n3336 ,
         \Reg_Bank/n3335 , \Reg_Bank/n3334 , \Reg_Bank/n3333 ,
         \Reg_Bank/n3332 , \Reg_Bank/n3331 , \Reg_Bank/n3330 ,
         \Reg_Bank/n3329 , \Reg_Bank/n3328 , \Reg_Bank/n3327 ,
         \Reg_Bank/n3326 , \Reg_Bank/n3325 , \Reg_Bank/n3324 ,
         \Reg_Bank/n3323 , \Reg_Bank/n3322 , \Reg_Bank/n3321 ,
         \Reg_Bank/n3320 , \Reg_Bank/n3319 , \Reg_Bank/n3318 ,
         \Reg_Bank/n3317 , \Reg_Bank/n3316 , \Reg_Bank/n3315 ,
         \Reg_Bank/n3314 , \Reg_Bank/n3313 , \Reg_Bank/n3312 ,
         \Reg_Bank/n3311 , \Reg_Bank/n3310 , \Reg_Bank/n3309 ,
         \Reg_Bank/n3308 , \Reg_Bank/n3307 , \Reg_Bank/n3306 ,
         \Reg_Bank/n3305 , \Reg_Bank/n3304 , \Reg_Bank/n3303 ,
         \Reg_Bank/n3302 , \Reg_Bank/n3301 , \Reg_Bank/n3300 ,
         \Reg_Bank/n3299 , \Reg_Bank/n3298 , \Reg_Bank/n3297 ,
         \Reg_Bank/n3296 , \Reg_Bank/n3295 , \Reg_Bank/n3294 ,
         \Reg_Bank/n3293 , \Reg_Bank/n3292 , \Reg_Bank/n3291 ,
         \Reg_Bank/n3290 , \Reg_Bank/n3289 , \Reg_Bank/n3288 ,
         \Reg_Bank/n3287 , \Reg_Bank/n3286 , \Reg_Bank/n3285 ,
         \Reg_Bank/n3284 , \Reg_Bank/n3283 , \Reg_Bank/n3282 ,
         \Reg_Bank/n3281 , \Reg_Bank/n3280 , \Reg_Bank/n3279 ,
         \Reg_Bank/n3278 , \Reg_Bank/n3277 , \Reg_Bank/n3276 ,
         \Reg_Bank/n3275 , \Reg_Bank/n3274 , \Reg_Bank/n3273 ,
         \Reg_Bank/n3272 , \Reg_Bank/n3271 , \Reg_Bank/n3270 ,
         \Reg_Bank/n3269 , \Reg_Bank/n3268 , \Reg_Bank/n3267 ,
         \Reg_Bank/n3266 , \Reg_Bank/n3265 , \Reg_Bank/n3264 ,
         \Reg_Bank/n3263 , \Reg_Bank/n3262 , \Reg_Bank/n3261 ,
         \Reg_Bank/n3260 , \Reg_Bank/n3259 , \Reg_Bank/n3258 ,
         \Reg_Bank/n3257 , \Reg_Bank/n3256 , \Reg_Bank/n3255 ,
         \Reg_Bank/n3254 , \Reg_Bank/n3253 , \Reg_Bank/n3252 ,
         \Reg_Bank/n3251 , \Reg_Bank/n3250 , \Reg_Bank/n3249 ,
         \Reg_Bank/n3248 , \Reg_Bank/n3247 , \Reg_Bank/n3246 ,
         \Reg_Bank/n3245 , \Reg_Bank/n3244 , \Reg_Bank/n3243 ,
         \Reg_Bank/n3242 , \Reg_Bank/n3241 , \Reg_Bank/n3240 ,
         \Reg_Bank/n3239 , \Reg_Bank/n3238 , \Reg_Bank/n3237 ,
         \Reg_Bank/n3236 , \Reg_Bank/n3235 , \Reg_Bank/n3234 ,
         \Reg_Bank/n3233 , \Reg_Bank/n3232 , \Reg_Bank/n3231 ,
         \Reg_Bank/n3230 , \Reg_Bank/n3229 , \Reg_Bank/n3228 ,
         \Reg_Bank/n3227 , \Reg_Bank/n3226 , \Reg_Bank/n3225 ,
         \Reg_Bank/n3224 , \Reg_Bank/n3223 , \Reg_Bank/n3222 ,
         \Reg_Bank/n3221 , \Reg_Bank/n3220 , \Reg_Bank/n3219 ,
         \Reg_Bank/n3218 , \Reg_Bank/n3217 , \Reg_Bank/n3216 ,
         \Reg_Bank/n3215 , \Reg_Bank/n3214 , \Reg_Bank/n3213 ,
         \Reg_Bank/n3212 , \Reg_Bank/n3211 , \Reg_Bank/n3210 ,
         \Reg_Bank/n3209 , \Reg_Bank/n3208 , \Reg_Bank/n3207 ,
         \Reg_Bank/n3206 , \Reg_Bank/n3205 , \Reg_Bank/n3204 ,
         \Reg_Bank/n3203 , \Reg_Bank/n3202 , \Reg_Bank/n3201 ,
         \Reg_Bank/n3200 , \Reg_Bank/n3199 , \Reg_Bank/n3198 ,
         \Reg_Bank/n3197 , \Reg_Bank/n3196 , \Reg_Bank/n3195 ,
         \Reg_Bank/n3194 , \Reg_Bank/n3193 , \Reg_Bank/n3192 ,
         \Reg_Bank/n3191 , \Reg_Bank/n3190 , \Reg_Bank/n3189 ,
         \Reg_Bank/n3188 , \Reg_Bank/n3187 , \Reg_Bank/n3186 ,
         \Reg_Bank/n3185 , \Reg_Bank/n3184 , \Reg_Bank/n3183 ,
         \Reg_Bank/n3182 , \Reg_Bank/n3181 , \Reg_Bank/n3180 ,
         \Reg_Bank/n3179 , \Reg_Bank/n3178 , \Reg_Bank/n3177 ,
         \Reg_Bank/n3176 , \Reg_Bank/n3175 , \Reg_Bank/n3174 ,
         \Reg_Bank/n3173 , \Reg_Bank/n3172 , \Reg_Bank/n3171 ,
         \Reg_Bank/n3170 , \Reg_Bank/n3169 , \Reg_Bank/n3168 ,
         \Reg_Bank/n3167 , \Reg_Bank/n3166 , \Reg_Bank/n3165 ,
         \Reg_Bank/n3164 , \Reg_Bank/n3163 , \Reg_Bank/n3162 ,
         \Reg_Bank/n3161 , \Reg_Bank/n3160 , \Reg_Bank/n3159 ,
         \Reg_Bank/n3158 , \Reg_Bank/n3157 , \Reg_Bank/n3156 ,
         \Reg_Bank/n3155 , \Reg_Bank/n3154 , \Reg_Bank/n3153 ,
         \Reg_Bank/n3152 , \Reg_Bank/n3151 , \Reg_Bank/n3150 ,
         \Reg_Bank/n3149 , \Reg_Bank/n3148 , \Reg_Bank/n3147 ,
         \Reg_Bank/n3146 , \Reg_Bank/n3145 , \Reg_Bank/n3144 ,
         \Reg_Bank/n3143 , \Reg_Bank/n3142 , \Reg_Bank/n3141 ,
         \Reg_Bank/n3140 , \Reg_Bank/n3139 , \Reg_Bank/n3138 ,
         \Reg_Bank/n3137 , \Reg_Bank/n3136 , \Reg_Bank/n3135 ,
         \Reg_Bank/n3134 , \Reg_Bank/n3133 , \Reg_Bank/n3132 ,
         \Reg_Bank/n3131 , \Reg_Bank/n3130 , \Reg_Bank/n3129 ,
         \Reg_Bank/n3128 , \Reg_Bank/n3127 , \Reg_Bank/n3126 ,
         \Reg_Bank/n3125 , \Reg_Bank/n3124 , \Reg_Bank/n3123 ,
         \Reg_Bank/n3122 , \Reg_Bank/n3121 , \Reg_Bank/n3120 ,
         \Reg_Bank/n3119 , \Reg_Bank/n3118 , \Reg_Bank/n3117 ,
         \Reg_Bank/n3116 , \Reg_Bank/n3115 , \Reg_Bank/n3114 ,
         \Reg_Bank/n3113 , \Reg_Bank/n3112 , \Reg_Bank/n3111 ,
         \Reg_Bank/n3110 , \Reg_Bank/n3109 , \Reg_Bank/n3108 ,
         \Reg_Bank/n3107 , \Reg_Bank/n3106 , \Reg_Bank/n3105 ,
         \Reg_Bank/n3104 , \Reg_Bank/n3103 , \Reg_Bank/n3102 ,
         \Reg_Bank/n3101 , \Reg_Bank/n3100 , \Reg_Bank/n3099 ,
         \Reg_Bank/n3098 , \Reg_Bank/n3097 , \Reg_Bank/n3096 ,
         \Reg_Bank/n3095 , \Reg_Bank/n3094 , \Reg_Bank/n3093 ,
         \Reg_Bank/n3092 , \Reg_Bank/n3091 , \Reg_Bank/n3090 ,
         \Reg_Bank/n3089 , \Reg_Bank/n3088 , \Reg_Bank/n3087 ,
         \Reg_Bank/n3086 , \Reg_Bank/n3085 , \Reg_Bank/n3084 ,
         \Reg_Bank/n3083 , \Reg_Bank/n3082 , \Reg_Bank/n3081 ,
         \Reg_Bank/n3080 , \Reg_Bank/n3079 , \Reg_Bank/n3078 ,
         \Reg_Bank/n3077 , \Reg_Bank/n3076 , \Reg_Bank/n3075 ,
         \Reg_Bank/n3074 , \Reg_Bank/n3073 , \Reg_Bank/n3072 ,
         \Reg_Bank/n3071 , \Reg_Bank/n3070 , \Reg_Bank/n3069 ,
         \Reg_Bank/n3068 , \Reg_Bank/n3067 , \Reg_Bank/n3066 ,
         \Reg_Bank/n3065 , \Reg_Bank/n3064 , \Reg_Bank/n3063 ,
         \Reg_Bank/n3062 , \Reg_Bank/n3061 , \Reg_Bank/n3060 ,
         \Reg_Bank/n3059 , \Reg_Bank/n3058 , \Reg_Bank/n3057 ,
         \Reg_Bank/n3056 , \Reg_Bank/n3055 , \Reg_Bank/n3054 ,
         \Reg_Bank/n3053 , \Reg_Bank/n3052 , \Reg_Bank/n3051 ,
         \Reg_Bank/n3050 , \Reg_Bank/n3049 , \Reg_Bank/n3048 ,
         \Reg_Bank/n3047 , \Reg_Bank/n3046 , \Reg_Bank/n3045 ,
         \Reg_Bank/n3044 , \Reg_Bank/n3043 , \Reg_Bank/n3042 ,
         \Reg_Bank/n3041 , \Reg_Bank/n3040 , \Reg_Bank/n3039 ,
         \Reg_Bank/n3038 , \Reg_Bank/n3037 , \Reg_Bank/n3036 ,
         \Reg_Bank/n3035 , \Reg_Bank/n3034 , \Reg_Bank/n3033 ,
         \Reg_Bank/n3032 , \Reg_Bank/n3031 , \Reg_Bank/n3030 ,
         \Reg_Bank/n3029 , \Reg_Bank/n3028 , \Reg_Bank/registers[1][0] ,
         \Reg_Bank/registers[1][1] , \Reg_Bank/registers[1][2] ,
         \Reg_Bank/registers[1][3] , \Reg_Bank/registers[1][4] ,
         \Reg_Bank/registers[1][5] , \Reg_Bank/registers[1][6] ,
         \Reg_Bank/registers[1][7] , \Reg_Bank/registers[1][8] ,
         \Reg_Bank/registers[1][9] , \Reg_Bank/registers[1][10] ,
         \Reg_Bank/registers[1][11] , \Reg_Bank/registers[1][12] ,
         \Reg_Bank/registers[1][13] , \Reg_Bank/registers[1][14] ,
         \Reg_Bank/registers[1][15] , \Reg_Bank/registers[1][16] ,
         \Reg_Bank/registers[1][17] , \Reg_Bank/registers[1][18] ,
         \Reg_Bank/registers[1][19] , \Reg_Bank/registers[1][20] ,
         \Reg_Bank/registers[1][21] , \Reg_Bank/registers[1][22] ,
         \Reg_Bank/registers[1][23] , \Reg_Bank/registers[1][24] ,
         \Reg_Bank/registers[1][25] , \Reg_Bank/registers[1][26] ,
         \Reg_Bank/registers[1][27] , \Reg_Bank/registers[1][28] ,
         \Reg_Bank/registers[1][29] , \Reg_Bank/registers[1][30] ,
         \Reg_Bank/registers[1][31] , \Reg_Bank/registers[2][0] ,
         \Reg_Bank/registers[2][1] , \Reg_Bank/registers[2][2] ,
         \Reg_Bank/registers[2][3] , \Reg_Bank/registers[2][4] ,
         \Reg_Bank/registers[2][5] , \Reg_Bank/registers[2][6] ,
         \Reg_Bank/registers[2][7] , \Reg_Bank/registers[2][8] ,
         \Reg_Bank/registers[2][9] , \Reg_Bank/registers[2][10] ,
         \Reg_Bank/registers[2][11] , \Reg_Bank/registers[2][12] ,
         \Reg_Bank/registers[2][13] , \Reg_Bank/registers[2][14] ,
         \Reg_Bank/registers[2][15] , \Reg_Bank/registers[2][16] ,
         \Reg_Bank/registers[2][17] , \Reg_Bank/registers[2][18] ,
         \Reg_Bank/registers[2][19] , \Reg_Bank/registers[2][20] ,
         \Reg_Bank/registers[2][21] , \Reg_Bank/registers[2][22] ,
         \Reg_Bank/registers[2][23] , \Reg_Bank/registers[2][24] ,
         \Reg_Bank/registers[2][25] , \Reg_Bank/registers[2][26] ,
         \Reg_Bank/registers[2][27] , \Reg_Bank/registers[2][28] ,
         \Reg_Bank/registers[2][29] , \Reg_Bank/registers[2][30] ,
         \Reg_Bank/registers[2][31] , \Reg_Bank/registers[3][0] ,
         \Reg_Bank/registers[3][1] , \Reg_Bank/registers[3][2] ,
         \Reg_Bank/registers[3][3] , \Reg_Bank/registers[3][4] ,
         \Reg_Bank/registers[3][5] , \Reg_Bank/registers[3][6] ,
         \Reg_Bank/registers[3][7] , \Reg_Bank/registers[3][8] ,
         \Reg_Bank/registers[3][9] , \Reg_Bank/registers[3][10] ,
         \Reg_Bank/registers[3][11] , \Reg_Bank/registers[3][12] ,
         \Reg_Bank/registers[3][13] , \Reg_Bank/registers[3][14] ,
         \Reg_Bank/registers[3][15] , \Reg_Bank/registers[3][16] ,
         \Reg_Bank/registers[3][17] , \Reg_Bank/registers[3][18] ,
         \Reg_Bank/registers[3][19] , \Reg_Bank/registers[3][20] ,
         \Reg_Bank/registers[3][21] , \Reg_Bank/registers[3][22] ,
         \Reg_Bank/registers[3][23] , \Reg_Bank/registers[3][24] ,
         \Reg_Bank/registers[3][25] , \Reg_Bank/registers[3][26] ,
         \Reg_Bank/registers[3][27] , \Reg_Bank/registers[3][28] ,
         \Reg_Bank/registers[3][29] , \Reg_Bank/registers[3][30] ,
         \Reg_Bank/registers[3][31] , \Reg_Bank/registers[4][0] ,
         \Reg_Bank/registers[4][1] , \Reg_Bank/registers[4][2] ,
         \Reg_Bank/registers[4][3] , \Reg_Bank/registers[4][4] ,
         \Reg_Bank/registers[4][5] , \Reg_Bank/registers[4][6] ,
         \Reg_Bank/registers[4][7] , \Reg_Bank/registers[4][8] ,
         \Reg_Bank/registers[4][9] , \Reg_Bank/registers[4][10] ,
         \Reg_Bank/registers[4][11] , \Reg_Bank/registers[4][12] ,
         \Reg_Bank/registers[4][13] , \Reg_Bank/registers[4][14] ,
         \Reg_Bank/registers[4][15] , \Reg_Bank/registers[4][16] ,
         \Reg_Bank/registers[4][17] , \Reg_Bank/registers[4][18] ,
         \Reg_Bank/registers[4][19] , \Reg_Bank/registers[4][20] ,
         \Reg_Bank/registers[4][21] , \Reg_Bank/registers[4][22] ,
         \Reg_Bank/registers[4][23] , \Reg_Bank/registers[4][24] ,
         \Reg_Bank/registers[4][25] , \Reg_Bank/registers[4][26] ,
         \Reg_Bank/registers[4][27] , \Reg_Bank/registers[4][28] ,
         \Reg_Bank/registers[4][29] , \Reg_Bank/registers[4][30] ,
         \Reg_Bank/registers[4][31] , \Reg_Bank/registers[5][0] ,
         \Reg_Bank/registers[5][1] , \Reg_Bank/registers[5][2] ,
         \Reg_Bank/registers[5][3] , \Reg_Bank/registers[5][4] ,
         \Reg_Bank/registers[5][5] , \Reg_Bank/registers[5][6] ,
         \Reg_Bank/registers[5][7] , \Reg_Bank/registers[5][8] ,
         \Reg_Bank/registers[5][9] , \Reg_Bank/registers[5][10] ,
         \Reg_Bank/registers[5][11] , \Reg_Bank/registers[5][12] ,
         \Reg_Bank/registers[5][13] , \Reg_Bank/registers[5][14] ,
         \Reg_Bank/registers[5][15] , \Reg_Bank/registers[5][16] ,
         \Reg_Bank/registers[5][17] , \Reg_Bank/registers[5][18] ,
         \Reg_Bank/registers[5][19] , \Reg_Bank/registers[5][20] ,
         \Reg_Bank/registers[5][21] , \Reg_Bank/registers[5][22] ,
         \Reg_Bank/registers[5][23] , \Reg_Bank/registers[5][24] ,
         \Reg_Bank/registers[5][25] , \Reg_Bank/registers[5][26] ,
         \Reg_Bank/registers[5][27] , \Reg_Bank/registers[5][28] ,
         \Reg_Bank/registers[5][29] , \Reg_Bank/registers[5][30] ,
         \Reg_Bank/registers[5][31] , \Reg_Bank/registers[6][0] ,
         \Reg_Bank/registers[6][1] , \Reg_Bank/registers[6][2] ,
         \Reg_Bank/registers[6][3] , \Reg_Bank/registers[6][4] ,
         \Reg_Bank/registers[6][5] , \Reg_Bank/registers[6][6] ,
         \Reg_Bank/registers[6][7] , \Reg_Bank/registers[6][8] ,
         \Reg_Bank/registers[6][9] , \Reg_Bank/registers[6][10] ,
         \Reg_Bank/registers[6][11] , \Reg_Bank/registers[6][12] ,
         \Reg_Bank/registers[6][13] , \Reg_Bank/registers[6][14] ,
         \Reg_Bank/registers[6][15] , \Reg_Bank/registers[6][16] ,
         \Reg_Bank/registers[6][17] , \Reg_Bank/registers[6][18] ,
         \Reg_Bank/registers[6][19] , \Reg_Bank/registers[6][20] ,
         \Reg_Bank/registers[6][21] , \Reg_Bank/registers[6][22] ,
         \Reg_Bank/registers[6][23] , \Reg_Bank/registers[6][24] ,
         \Reg_Bank/registers[6][25] , \Reg_Bank/registers[6][26] ,
         \Reg_Bank/registers[6][27] , \Reg_Bank/registers[6][28] ,
         \Reg_Bank/registers[6][29] , \Reg_Bank/registers[6][30] ,
         \Reg_Bank/registers[6][31] , \Reg_Bank/registers[7][0] ,
         \Reg_Bank/registers[7][1] , \Reg_Bank/registers[7][2] ,
         \Reg_Bank/registers[7][3] , \Reg_Bank/registers[7][4] ,
         \Reg_Bank/registers[7][5] , \Reg_Bank/registers[7][6] ,
         \Reg_Bank/registers[7][7] , \Reg_Bank/registers[7][8] ,
         \Reg_Bank/registers[7][9] , \Reg_Bank/registers[7][10] ,
         \Reg_Bank/registers[7][11] , \Reg_Bank/registers[7][12] ,
         \Reg_Bank/registers[7][13] , \Reg_Bank/registers[7][14] ,
         \Reg_Bank/registers[7][15] , \Reg_Bank/registers[7][16] ,
         \Reg_Bank/registers[7][17] , \Reg_Bank/registers[7][18] ,
         \Reg_Bank/registers[7][19] , \Reg_Bank/registers[7][20] ,
         \Reg_Bank/registers[7][21] , \Reg_Bank/registers[7][22] ,
         \Reg_Bank/registers[7][23] , \Reg_Bank/registers[7][24] ,
         \Reg_Bank/registers[7][25] , \Reg_Bank/registers[7][26] ,
         \Reg_Bank/registers[7][27] , \Reg_Bank/registers[7][28] ,
         \Reg_Bank/registers[7][29] , \Reg_Bank/registers[7][30] ,
         \Reg_Bank/registers[7][31] , \Reg_Bank/registers[8][0] ,
         \Reg_Bank/registers[8][1] , \Reg_Bank/registers[8][2] ,
         \Reg_Bank/registers[8][3] , \Reg_Bank/registers[8][4] ,
         \Reg_Bank/registers[8][5] , \Reg_Bank/registers[8][6] ,
         \Reg_Bank/registers[8][7] , \Reg_Bank/registers[8][8] ,
         \Reg_Bank/registers[8][9] , \Reg_Bank/registers[8][10] ,
         \Reg_Bank/registers[8][11] , \Reg_Bank/registers[8][12] ,
         \Reg_Bank/registers[8][13] , \Reg_Bank/registers[8][14] ,
         \Reg_Bank/registers[8][15] , \Reg_Bank/registers[8][16] ,
         \Reg_Bank/registers[8][17] , \Reg_Bank/registers[8][18] ,
         \Reg_Bank/registers[8][19] , \Reg_Bank/registers[8][20] ,
         \Reg_Bank/registers[8][21] , \Reg_Bank/registers[8][22] ,
         \Reg_Bank/registers[8][23] , \Reg_Bank/registers[8][24] ,
         \Reg_Bank/registers[8][25] , \Reg_Bank/registers[8][26] ,
         \Reg_Bank/registers[8][27] , \Reg_Bank/registers[8][28] ,
         \Reg_Bank/registers[8][29] , \Reg_Bank/registers[8][30] ,
         \Reg_Bank/registers[8][31] , \Reg_Bank/registers[9][0] ,
         \Reg_Bank/registers[9][1] , \Reg_Bank/registers[9][2] ,
         \Reg_Bank/registers[9][3] , \Reg_Bank/registers[9][4] ,
         \Reg_Bank/registers[9][5] , \Reg_Bank/registers[9][6] ,
         \Reg_Bank/registers[9][7] , \Reg_Bank/registers[9][8] ,
         \Reg_Bank/registers[9][9] , \Reg_Bank/registers[9][10] ,
         \Reg_Bank/registers[9][11] , \Reg_Bank/registers[9][12] ,
         \Reg_Bank/registers[9][13] , \Reg_Bank/registers[9][14] ,
         \Reg_Bank/registers[9][15] , \Reg_Bank/registers[9][16] ,
         \Reg_Bank/registers[9][17] , \Reg_Bank/registers[9][18] ,
         \Reg_Bank/registers[9][19] , \Reg_Bank/registers[9][20] ,
         \Reg_Bank/registers[9][21] , \Reg_Bank/registers[9][22] ,
         \Reg_Bank/registers[9][23] , \Reg_Bank/registers[9][24] ,
         \Reg_Bank/registers[9][25] , \Reg_Bank/registers[9][26] ,
         \Reg_Bank/registers[9][27] , \Reg_Bank/registers[9][28] ,
         \Reg_Bank/registers[9][29] , \Reg_Bank/registers[9][30] ,
         \Reg_Bank/registers[9][31] , \Reg_Bank/registers[10][0] ,
         \Reg_Bank/registers[10][1] , \Reg_Bank/registers[10][2] ,
         \Reg_Bank/registers[10][3] , \Reg_Bank/registers[10][4] ,
         \Reg_Bank/registers[10][5] , \Reg_Bank/registers[10][6] ,
         \Reg_Bank/registers[10][7] , \Reg_Bank/registers[10][8] ,
         \Reg_Bank/registers[10][9] , \Reg_Bank/registers[10][10] ,
         \Reg_Bank/registers[10][11] , \Reg_Bank/registers[10][12] ,
         \Reg_Bank/registers[10][13] , \Reg_Bank/registers[10][14] ,
         \Reg_Bank/registers[10][15] , \Reg_Bank/registers[10][16] ,
         \Reg_Bank/registers[10][17] , \Reg_Bank/registers[10][18] ,
         \Reg_Bank/registers[10][19] , \Reg_Bank/registers[10][20] ,
         \Reg_Bank/registers[10][21] , \Reg_Bank/registers[10][22] ,
         \Reg_Bank/registers[10][23] , \Reg_Bank/registers[10][24] ,
         \Reg_Bank/registers[10][25] , \Reg_Bank/registers[10][26] ,
         \Reg_Bank/registers[10][27] , \Reg_Bank/registers[10][28] ,
         \Reg_Bank/registers[10][29] , \Reg_Bank/registers[10][30] ,
         \Reg_Bank/registers[10][31] , \Reg_Bank/registers[11][0] ,
         \Reg_Bank/registers[11][1] , \Reg_Bank/registers[11][2] ,
         \Reg_Bank/registers[11][3] , \Reg_Bank/registers[11][4] ,
         \Reg_Bank/registers[11][5] , \Reg_Bank/registers[11][6] ,
         \Reg_Bank/registers[11][7] , \Reg_Bank/registers[11][8] ,
         \Reg_Bank/registers[11][9] , \Reg_Bank/registers[11][10] ,
         \Reg_Bank/registers[11][11] , \Reg_Bank/registers[11][12] ,
         \Reg_Bank/registers[11][13] , \Reg_Bank/registers[11][14] ,
         \Reg_Bank/registers[11][15] , \Reg_Bank/registers[11][16] ,
         \Reg_Bank/registers[11][17] , \Reg_Bank/registers[11][18] ,
         \Reg_Bank/registers[11][19] , \Reg_Bank/registers[11][20] ,
         \Reg_Bank/registers[11][21] , \Reg_Bank/registers[11][22] ,
         \Reg_Bank/registers[11][23] , \Reg_Bank/registers[11][24] ,
         \Reg_Bank/registers[11][25] , \Reg_Bank/registers[11][26] ,
         \Reg_Bank/registers[11][27] , \Reg_Bank/registers[11][28] ,
         \Reg_Bank/registers[11][29] , \Reg_Bank/registers[11][30] ,
         \Reg_Bank/registers[11][31] , \Reg_Bank/registers[12][0] ,
         \Reg_Bank/registers[12][1] , \Reg_Bank/registers[12][2] ,
         \Reg_Bank/registers[12][3] , \Reg_Bank/registers[12][4] ,
         \Reg_Bank/registers[12][5] , \Reg_Bank/registers[12][6] ,
         \Reg_Bank/registers[12][7] , \Reg_Bank/registers[12][8] ,
         \Reg_Bank/registers[12][9] , \Reg_Bank/registers[12][10] ,
         \Reg_Bank/registers[12][11] , \Reg_Bank/registers[12][12] ,
         \Reg_Bank/registers[12][13] , \Reg_Bank/registers[12][14] ,
         \Reg_Bank/registers[12][15] , \Reg_Bank/registers[12][16] ,
         \Reg_Bank/registers[12][17] , \Reg_Bank/registers[12][18] ,
         \Reg_Bank/registers[12][19] , \Reg_Bank/registers[12][20] ,
         \Reg_Bank/registers[12][21] , \Reg_Bank/registers[12][22] ,
         \Reg_Bank/registers[12][23] , \Reg_Bank/registers[12][24] ,
         \Reg_Bank/registers[12][25] , \Reg_Bank/registers[12][26] ,
         \Reg_Bank/registers[12][27] , \Reg_Bank/registers[12][28] ,
         \Reg_Bank/registers[12][29] , \Reg_Bank/registers[12][30] ,
         \Reg_Bank/registers[12][31] , \Reg_Bank/registers[13][0] ,
         \Reg_Bank/registers[13][1] , \Reg_Bank/registers[13][2] ,
         \Reg_Bank/registers[13][3] , \Reg_Bank/registers[13][4] ,
         \Reg_Bank/registers[13][5] , \Reg_Bank/registers[13][6] ,
         \Reg_Bank/registers[13][7] , \Reg_Bank/registers[13][8] ,
         \Reg_Bank/registers[13][9] , \Reg_Bank/registers[13][10] ,
         \Reg_Bank/registers[13][11] , \Reg_Bank/registers[13][12] ,
         \Reg_Bank/registers[13][13] , \Reg_Bank/registers[13][14] ,
         \Reg_Bank/registers[13][15] , \Reg_Bank/registers[13][16] ,
         \Reg_Bank/registers[13][17] , \Reg_Bank/registers[13][18] ,
         \Reg_Bank/registers[13][19] , \Reg_Bank/registers[13][20] ,
         \Reg_Bank/registers[13][21] , \Reg_Bank/registers[13][22] ,
         \Reg_Bank/registers[13][23] , \Reg_Bank/registers[13][24] ,
         \Reg_Bank/registers[13][25] , \Reg_Bank/registers[13][26] ,
         \Reg_Bank/registers[13][27] , \Reg_Bank/registers[13][28] ,
         \Reg_Bank/registers[13][29] , \Reg_Bank/registers[13][30] ,
         \Reg_Bank/registers[13][31] , \Reg_Bank/registers[14][0] ,
         \Reg_Bank/registers[14][1] , \Reg_Bank/registers[14][2] ,
         \Reg_Bank/registers[14][3] , \Reg_Bank/registers[14][4] ,
         \Reg_Bank/registers[14][5] , \Reg_Bank/registers[14][6] ,
         \Reg_Bank/registers[14][7] , \Reg_Bank/registers[14][8] ,
         \Reg_Bank/registers[14][9] , \Reg_Bank/registers[14][10] ,
         \Reg_Bank/registers[14][11] , \Reg_Bank/registers[14][12] ,
         \Reg_Bank/registers[14][13] , \Reg_Bank/registers[14][14] ,
         \Reg_Bank/registers[14][15] , \Reg_Bank/registers[14][16] ,
         \Reg_Bank/registers[14][17] , \Reg_Bank/registers[14][18] ,
         \Reg_Bank/registers[14][19] , \Reg_Bank/registers[14][20] ,
         \Reg_Bank/registers[14][21] , \Reg_Bank/registers[14][22] ,
         \Reg_Bank/registers[14][23] , \Reg_Bank/registers[14][24] ,
         \Reg_Bank/registers[14][25] , \Reg_Bank/registers[14][26] ,
         \Reg_Bank/registers[14][27] , \Reg_Bank/registers[14][28] ,
         \Reg_Bank/registers[14][29] , \Reg_Bank/registers[14][30] ,
         \Reg_Bank/registers[14][31] , \Reg_Bank/registers[15][0] ,
         \Reg_Bank/registers[15][1] , \Reg_Bank/registers[15][2] ,
         \Reg_Bank/registers[15][3] , \Reg_Bank/registers[15][4] ,
         \Reg_Bank/registers[15][5] , \Reg_Bank/registers[15][6] ,
         \Reg_Bank/registers[15][7] , \Reg_Bank/registers[15][8] ,
         \Reg_Bank/registers[15][9] , \Reg_Bank/registers[15][10] ,
         \Reg_Bank/registers[15][11] , \Reg_Bank/registers[15][12] ,
         \Reg_Bank/registers[15][13] , \Reg_Bank/registers[15][14] ,
         \Reg_Bank/registers[15][15] , \Reg_Bank/registers[15][16] ,
         \Reg_Bank/registers[15][17] , \Reg_Bank/registers[15][18] ,
         \Reg_Bank/registers[15][19] , \Reg_Bank/registers[15][20] ,
         \Reg_Bank/registers[15][21] , \Reg_Bank/registers[15][22] ,
         \Reg_Bank/registers[15][23] , \Reg_Bank/registers[15][24] ,
         \Reg_Bank/registers[15][25] , \Reg_Bank/registers[15][26] ,
         \Reg_Bank/registers[15][27] , \Reg_Bank/registers[15][28] ,
         \Reg_Bank/registers[15][29] , \Reg_Bank/registers[15][30] ,
         \Reg_Bank/registers[15][31] , \Reg_Bank/registers[16][0] ,
         \Reg_Bank/registers[16][1] , \Reg_Bank/registers[16][2] ,
         \Reg_Bank/registers[16][3] , \Reg_Bank/registers[16][4] ,
         \Reg_Bank/registers[16][5] , \Reg_Bank/registers[16][6] ,
         \Reg_Bank/registers[16][7] , \Reg_Bank/registers[16][8] ,
         \Reg_Bank/registers[16][9] , \Reg_Bank/registers[16][10] ,
         \Reg_Bank/registers[16][11] , \Reg_Bank/registers[16][12] ,
         \Reg_Bank/registers[16][13] , \Reg_Bank/registers[16][14] ,
         \Reg_Bank/registers[16][15] , \Reg_Bank/registers[16][16] ,
         \Reg_Bank/registers[16][17] , \Reg_Bank/registers[16][18] ,
         \Reg_Bank/registers[16][19] , \Reg_Bank/registers[16][20] ,
         \Reg_Bank/registers[16][21] , \Reg_Bank/registers[16][22] ,
         \Reg_Bank/registers[16][23] , \Reg_Bank/registers[16][24] ,
         \Reg_Bank/registers[16][25] , \Reg_Bank/registers[16][26] ,
         \Reg_Bank/registers[16][27] , \Reg_Bank/registers[16][28] ,
         \Reg_Bank/registers[16][29] , \Reg_Bank/registers[16][30] ,
         \Reg_Bank/registers[16][31] , \Reg_Bank/registers[17][0] ,
         \Reg_Bank/registers[17][1] , \Reg_Bank/registers[17][2] ,
         \Reg_Bank/registers[17][3] , \Reg_Bank/registers[17][4] ,
         \Reg_Bank/registers[17][5] , \Reg_Bank/registers[17][6] ,
         \Reg_Bank/registers[17][7] , \Reg_Bank/registers[17][8] ,
         \Reg_Bank/registers[17][9] , \Reg_Bank/registers[17][10] ,
         \Reg_Bank/registers[17][11] , \Reg_Bank/registers[17][12] ,
         \Reg_Bank/registers[17][13] , \Reg_Bank/registers[17][14] ,
         \Reg_Bank/registers[17][15] , \Reg_Bank/registers[17][16] ,
         \Reg_Bank/registers[17][17] , \Reg_Bank/registers[17][18] ,
         \Reg_Bank/registers[17][19] , \Reg_Bank/registers[17][20] ,
         \Reg_Bank/registers[17][21] , \Reg_Bank/registers[17][22] ,
         \Reg_Bank/registers[17][23] , \Reg_Bank/registers[17][24] ,
         \Reg_Bank/registers[17][25] , \Reg_Bank/registers[17][26] ,
         \Reg_Bank/registers[17][27] , \Reg_Bank/registers[17][28] ,
         \Reg_Bank/registers[17][29] , \Reg_Bank/registers[17][30] ,
         \Reg_Bank/registers[17][31] , \Reg_Bank/registers[18][0] ,
         \Reg_Bank/registers[18][1] , \Reg_Bank/registers[18][2] ,
         \Reg_Bank/registers[18][3] , \Reg_Bank/registers[18][4] ,
         \Reg_Bank/registers[18][5] , \Reg_Bank/registers[18][6] ,
         \Reg_Bank/registers[18][7] , \Reg_Bank/registers[18][8] ,
         \Reg_Bank/registers[18][9] , \Reg_Bank/registers[18][10] ,
         \Reg_Bank/registers[18][11] , \Reg_Bank/registers[18][12] ,
         \Reg_Bank/registers[18][13] , \Reg_Bank/registers[18][14] ,
         \Reg_Bank/registers[18][15] , \Reg_Bank/registers[18][16] ,
         \Reg_Bank/registers[18][17] , \Reg_Bank/registers[18][18] ,
         \Reg_Bank/registers[18][19] , \Reg_Bank/registers[18][20] ,
         \Reg_Bank/registers[18][21] , \Reg_Bank/registers[18][22] ,
         \Reg_Bank/registers[18][23] , \Reg_Bank/registers[18][24] ,
         \Reg_Bank/registers[18][25] , \Reg_Bank/registers[18][26] ,
         \Reg_Bank/registers[18][27] , \Reg_Bank/registers[18][28] ,
         \Reg_Bank/registers[18][29] , \Reg_Bank/registers[18][30] ,
         \Reg_Bank/registers[18][31] , \Reg_Bank/registers[19][0] ,
         \Reg_Bank/registers[19][1] , \Reg_Bank/registers[19][2] ,
         \Reg_Bank/registers[19][3] , \Reg_Bank/registers[19][4] ,
         \Reg_Bank/registers[19][5] , \Reg_Bank/registers[19][6] ,
         \Reg_Bank/registers[19][7] , \Reg_Bank/registers[19][8] ,
         \Reg_Bank/registers[19][9] , \Reg_Bank/registers[19][10] ,
         \Reg_Bank/registers[19][11] , \Reg_Bank/registers[19][12] ,
         \Reg_Bank/registers[19][13] , \Reg_Bank/registers[19][14] ,
         \Reg_Bank/registers[19][15] , \Reg_Bank/registers[19][16] ,
         \Reg_Bank/registers[19][17] , \Reg_Bank/registers[19][18] ,
         \Reg_Bank/registers[19][19] , \Reg_Bank/registers[19][20] ,
         \Reg_Bank/registers[19][21] , \Reg_Bank/registers[19][22] ,
         \Reg_Bank/registers[19][23] , \Reg_Bank/registers[19][24] ,
         \Reg_Bank/registers[19][25] , \Reg_Bank/registers[19][26] ,
         \Reg_Bank/registers[19][27] , \Reg_Bank/registers[19][28] ,
         \Reg_Bank/registers[19][29] , \Reg_Bank/registers[19][30] ,
         \Reg_Bank/registers[19][31] , \Reg_Bank/registers[20][0] ,
         \Reg_Bank/registers[20][1] , \Reg_Bank/registers[20][2] ,
         \Reg_Bank/registers[20][3] , \Reg_Bank/registers[20][4] ,
         \Reg_Bank/registers[20][5] , \Reg_Bank/registers[20][6] ,
         \Reg_Bank/registers[20][7] , \Reg_Bank/registers[20][8] ,
         \Reg_Bank/registers[20][9] , \Reg_Bank/registers[20][10] ,
         \Reg_Bank/registers[20][11] , \Reg_Bank/registers[20][12] ,
         \Reg_Bank/registers[20][13] , \Reg_Bank/registers[20][14] ,
         \Reg_Bank/registers[20][15] , \Reg_Bank/registers[20][16] ,
         \Reg_Bank/registers[20][17] , \Reg_Bank/registers[20][18] ,
         \Reg_Bank/registers[20][19] , \Reg_Bank/registers[20][20] ,
         \Reg_Bank/registers[20][21] , \Reg_Bank/registers[20][22] ,
         \Reg_Bank/registers[20][23] , \Reg_Bank/registers[20][24] ,
         \Reg_Bank/registers[20][25] , \Reg_Bank/registers[20][26] ,
         \Reg_Bank/registers[20][27] , \Reg_Bank/registers[20][28] ,
         \Reg_Bank/registers[20][29] , \Reg_Bank/registers[20][30] ,
         \Reg_Bank/registers[20][31] , \Reg_Bank/registers[21][0] ,
         \Reg_Bank/registers[21][1] , \Reg_Bank/registers[21][2] ,
         \Reg_Bank/registers[21][3] , \Reg_Bank/registers[21][4] ,
         \Reg_Bank/registers[21][5] , \Reg_Bank/registers[21][6] ,
         \Reg_Bank/registers[21][7] , \Reg_Bank/registers[21][8] ,
         \Reg_Bank/registers[21][9] , \Reg_Bank/registers[21][10] ,
         \Reg_Bank/registers[21][11] , \Reg_Bank/registers[21][12] ,
         \Reg_Bank/registers[21][13] , \Reg_Bank/registers[21][14] ,
         \Reg_Bank/registers[21][15] , \Reg_Bank/registers[21][16] ,
         \Reg_Bank/registers[21][17] , \Reg_Bank/registers[21][18] ,
         \Reg_Bank/registers[21][19] , \Reg_Bank/registers[21][20] ,
         \Reg_Bank/registers[21][21] , \Reg_Bank/registers[21][22] ,
         \Reg_Bank/registers[21][23] , \Reg_Bank/registers[21][24] ,
         \Reg_Bank/registers[21][25] , \Reg_Bank/registers[21][26] ,
         \Reg_Bank/registers[21][27] , \Reg_Bank/registers[21][28] ,
         \Reg_Bank/registers[21][29] , \Reg_Bank/registers[21][30] ,
         \Reg_Bank/registers[21][31] , \Reg_Bank/registers[22][0] ,
         \Reg_Bank/registers[22][1] , \Reg_Bank/registers[22][2] ,
         \Reg_Bank/registers[22][3] , \Reg_Bank/registers[22][4] ,
         \Reg_Bank/registers[22][5] , \Reg_Bank/registers[22][6] ,
         \Reg_Bank/registers[22][7] , \Reg_Bank/registers[22][8] ,
         \Reg_Bank/registers[22][9] , \Reg_Bank/registers[22][10] ,
         \Reg_Bank/registers[22][11] , \Reg_Bank/registers[22][12] ,
         \Reg_Bank/registers[22][13] , \Reg_Bank/registers[22][14] ,
         \Reg_Bank/registers[22][15] , \Reg_Bank/registers[22][16] ,
         \Reg_Bank/registers[22][17] , \Reg_Bank/registers[22][18] ,
         \Reg_Bank/registers[22][19] , \Reg_Bank/registers[22][20] ,
         \Reg_Bank/registers[22][21] , \Reg_Bank/registers[22][22] ,
         \Reg_Bank/registers[22][23] , \Reg_Bank/registers[22][24] ,
         \Reg_Bank/registers[22][25] , \Reg_Bank/registers[22][26] ,
         \Reg_Bank/registers[22][27] , \Reg_Bank/registers[22][28] ,
         \Reg_Bank/registers[22][29] , \Reg_Bank/registers[22][30] ,
         \Reg_Bank/registers[22][31] , \Reg_Bank/registers[23][0] ,
         \Reg_Bank/registers[23][1] , \Reg_Bank/registers[23][2] ,
         \Reg_Bank/registers[23][3] , \Reg_Bank/registers[23][4] ,
         \Reg_Bank/registers[23][5] , \Reg_Bank/registers[23][6] ,
         \Reg_Bank/registers[23][7] , \Reg_Bank/registers[23][8] ,
         \Reg_Bank/registers[23][9] , \Reg_Bank/registers[23][10] ,
         \Reg_Bank/registers[23][11] , \Reg_Bank/registers[23][12] ,
         \Reg_Bank/registers[23][13] , \Reg_Bank/registers[23][14] ,
         \Reg_Bank/registers[23][15] , \Reg_Bank/registers[23][16] ,
         \Reg_Bank/registers[23][17] , \Reg_Bank/registers[23][18] ,
         \Reg_Bank/registers[23][19] , \Reg_Bank/registers[23][20] ,
         \Reg_Bank/registers[23][21] , \Reg_Bank/registers[23][22] ,
         \Reg_Bank/registers[23][23] , \Reg_Bank/registers[23][24] ,
         \Reg_Bank/registers[23][25] , \Reg_Bank/registers[23][26] ,
         \Reg_Bank/registers[23][27] , \Reg_Bank/registers[23][28] ,
         \Reg_Bank/registers[23][29] , \Reg_Bank/registers[23][30] ,
         \Reg_Bank/registers[23][31] , \Reg_Bank/registers[24][0] ,
         \Reg_Bank/registers[24][1] , \Reg_Bank/registers[24][2] ,
         \Reg_Bank/registers[24][3] , \Reg_Bank/registers[24][4] ,
         \Reg_Bank/registers[24][5] , \Reg_Bank/registers[24][6] ,
         \Reg_Bank/registers[24][7] , \Reg_Bank/registers[24][8] ,
         \Reg_Bank/registers[24][9] , \Reg_Bank/registers[24][10] ,
         \Reg_Bank/registers[24][11] , \Reg_Bank/registers[24][12] ,
         \Reg_Bank/registers[24][13] , \Reg_Bank/registers[24][14] ,
         \Reg_Bank/registers[24][15] , \Reg_Bank/registers[24][16] ,
         \Reg_Bank/registers[24][17] , \Reg_Bank/registers[24][18] ,
         \Reg_Bank/registers[24][19] , \Reg_Bank/registers[24][20] ,
         \Reg_Bank/registers[24][21] , \Reg_Bank/registers[24][22] ,
         \Reg_Bank/registers[24][23] , \Reg_Bank/registers[24][24] ,
         \Reg_Bank/registers[24][25] , \Reg_Bank/registers[24][26] ,
         \Reg_Bank/registers[24][27] , \Reg_Bank/registers[24][28] ,
         \Reg_Bank/registers[24][29] , \Reg_Bank/registers[24][30] ,
         \Reg_Bank/registers[24][31] , \Reg_Bank/registers[25][0] ,
         \Reg_Bank/registers[25][1] , \Reg_Bank/registers[25][2] ,
         \Reg_Bank/registers[25][3] , \Reg_Bank/registers[25][4] ,
         \Reg_Bank/registers[25][5] , \Reg_Bank/registers[25][6] ,
         \Reg_Bank/registers[25][7] , \Reg_Bank/registers[25][8] ,
         \Reg_Bank/registers[25][9] , \Reg_Bank/registers[25][10] ,
         \Reg_Bank/registers[25][11] , \Reg_Bank/registers[25][12] ,
         \Reg_Bank/registers[25][13] , \Reg_Bank/registers[25][14] ,
         \Reg_Bank/registers[25][15] , \Reg_Bank/registers[25][16] ,
         \Reg_Bank/registers[25][17] , \Reg_Bank/registers[25][18] ,
         \Reg_Bank/registers[25][19] , \Reg_Bank/registers[25][20] ,
         \Reg_Bank/registers[25][21] , \Reg_Bank/registers[25][22] ,
         \Reg_Bank/registers[25][23] , \Reg_Bank/registers[25][24] ,
         \Reg_Bank/registers[25][25] , \Reg_Bank/registers[25][26] ,
         \Reg_Bank/registers[25][27] , \Reg_Bank/registers[25][28] ,
         \Reg_Bank/registers[25][29] , \Reg_Bank/registers[25][30] ,
         \Reg_Bank/registers[25][31] , \Reg_Bank/registers[26][0] ,
         \Reg_Bank/registers[26][1] , \Reg_Bank/registers[26][2] ,
         \Reg_Bank/registers[26][3] , \Reg_Bank/registers[26][4] ,
         \Reg_Bank/registers[26][5] , \Reg_Bank/registers[26][6] ,
         \Reg_Bank/registers[26][7] , \Reg_Bank/registers[26][8] ,
         \Reg_Bank/registers[26][9] , \Reg_Bank/registers[26][10] ,
         \Reg_Bank/registers[26][11] , \Reg_Bank/registers[26][12] ,
         \Reg_Bank/registers[26][13] , \Reg_Bank/registers[26][14] ,
         \Reg_Bank/registers[26][15] , \Reg_Bank/registers[26][16] ,
         \Reg_Bank/registers[26][17] , \Reg_Bank/registers[26][18] ,
         \Reg_Bank/registers[26][19] , \Reg_Bank/registers[26][20] ,
         \Reg_Bank/registers[26][21] , \Reg_Bank/registers[26][22] ,
         \Reg_Bank/registers[26][23] , \Reg_Bank/registers[26][24] ,
         \Reg_Bank/registers[26][25] , \Reg_Bank/registers[26][26] ,
         \Reg_Bank/registers[26][27] , \Reg_Bank/registers[26][28] ,
         \Reg_Bank/registers[26][29] , \Reg_Bank/registers[26][30] ,
         \Reg_Bank/registers[26][31] , \Reg_Bank/registers[27][0] ,
         \Reg_Bank/registers[27][1] , \Reg_Bank/registers[27][2] ,
         \Reg_Bank/registers[27][3] , \Reg_Bank/registers[27][4] ,
         \Reg_Bank/registers[27][5] , \Reg_Bank/registers[27][6] ,
         \Reg_Bank/registers[27][7] , \Reg_Bank/registers[27][8] ,
         \Reg_Bank/registers[27][9] , \Reg_Bank/registers[27][10] ,
         \Reg_Bank/registers[27][11] , \Reg_Bank/registers[27][12] ,
         \Reg_Bank/registers[27][13] , \Reg_Bank/registers[27][14] ,
         \Reg_Bank/registers[27][15] , \Reg_Bank/registers[27][16] ,
         \Reg_Bank/registers[27][17] , \Reg_Bank/registers[27][18] ,
         \Reg_Bank/registers[27][19] , \Reg_Bank/registers[27][20] ,
         \Reg_Bank/registers[27][21] , \Reg_Bank/registers[27][22] ,
         \Reg_Bank/registers[27][23] , \Reg_Bank/registers[27][24] ,
         \Reg_Bank/registers[27][25] , \Reg_Bank/registers[27][26] ,
         \Reg_Bank/registers[27][27] , \Reg_Bank/registers[27][28] ,
         \Reg_Bank/registers[27][29] , \Reg_Bank/registers[27][30] ,
         \Reg_Bank/registers[27][31] , \Reg_Bank/registers[28][0] ,
         \Reg_Bank/registers[28][1] , \Reg_Bank/registers[28][2] ,
         \Reg_Bank/registers[28][3] , \Reg_Bank/registers[28][4] ,
         \Reg_Bank/registers[28][5] , \Reg_Bank/registers[28][6] ,
         \Reg_Bank/registers[28][7] , \Reg_Bank/registers[28][8] ,
         \Reg_Bank/registers[28][9] , \Reg_Bank/registers[28][10] ,
         \Reg_Bank/registers[28][11] , \Reg_Bank/registers[28][12] ,
         \Reg_Bank/registers[28][13] , \Reg_Bank/registers[28][14] ,
         \Reg_Bank/registers[28][15] , \Reg_Bank/registers[28][16] ,
         \Reg_Bank/registers[28][17] , \Reg_Bank/registers[28][18] ,
         \Reg_Bank/registers[28][19] , \Reg_Bank/registers[28][20] ,
         \Reg_Bank/registers[28][21] , \Reg_Bank/registers[28][22] ,
         \Reg_Bank/registers[28][23] , \Reg_Bank/registers[28][24] ,
         \Reg_Bank/registers[28][25] , \Reg_Bank/registers[28][26] ,
         \Reg_Bank/registers[28][27] , \Reg_Bank/registers[28][28] ,
         \Reg_Bank/registers[28][29] , \Reg_Bank/registers[28][30] ,
         \Reg_Bank/registers[28][31] , \Reg_Bank/registers[29][0] ,
         \Reg_Bank/registers[29][1] , \Reg_Bank/registers[29][2] ,
         \Reg_Bank/registers[29][3] , \Reg_Bank/registers[29][4] ,
         \Reg_Bank/registers[29][5] , \Reg_Bank/registers[29][6] ,
         \Reg_Bank/registers[29][7] , \Reg_Bank/registers[29][8] ,
         \Reg_Bank/registers[29][9] , \Reg_Bank/registers[29][10] ,
         \Reg_Bank/registers[29][11] , \Reg_Bank/registers[29][12] ,
         \Reg_Bank/registers[29][13] , \Reg_Bank/registers[29][14] ,
         \Reg_Bank/registers[29][15] , \Reg_Bank/registers[29][16] ,
         \Reg_Bank/registers[29][17] , \Reg_Bank/registers[29][18] ,
         \Reg_Bank/registers[29][19] , \Reg_Bank/registers[29][20] ,
         \Reg_Bank/registers[29][21] , \Reg_Bank/registers[29][22] ,
         \Reg_Bank/registers[29][23] , \Reg_Bank/registers[29][24] ,
         \Reg_Bank/registers[29][25] , \Reg_Bank/registers[29][26] ,
         \Reg_Bank/registers[29][27] , \Reg_Bank/registers[29][28] ,
         \Reg_Bank/registers[29][29] , \Reg_Bank/registers[29][30] ,
         \Reg_Bank/registers[29][31] , \Reg_Bank/registers[30][0] ,
         \Reg_Bank/registers[30][1] , \Reg_Bank/registers[30][2] ,
         \Reg_Bank/registers[30][3] , \Reg_Bank/registers[30][4] ,
         \Reg_Bank/registers[30][5] , \Reg_Bank/registers[30][6] ,
         \Reg_Bank/registers[30][7] , \Reg_Bank/registers[30][8] ,
         \Reg_Bank/registers[30][9] , \Reg_Bank/registers[30][10] ,
         \Reg_Bank/registers[30][11] , \Reg_Bank/registers[30][12] ,
         \Reg_Bank/registers[30][13] , \Reg_Bank/registers[30][14] ,
         \Reg_Bank/registers[30][15] , \Reg_Bank/registers[30][16] ,
         \Reg_Bank/registers[30][17] , \Reg_Bank/registers[30][18] ,
         \Reg_Bank/registers[30][19] , \Reg_Bank/registers[30][20] ,
         \Reg_Bank/registers[30][21] , \Reg_Bank/registers[30][22] ,
         \Reg_Bank/registers[30][23] , \Reg_Bank/registers[30][24] ,
         \Reg_Bank/registers[30][25] , \Reg_Bank/registers[30][26] ,
         \Reg_Bank/registers[30][27] , \Reg_Bank/registers[30][28] ,
         \Reg_Bank/registers[30][29] , \Reg_Bank/registers[30][30] ,
         \Reg_Bank/registers[30][31] , \Reg_Bank/registers[31][0] ,
         \Reg_Bank/registers[31][1] , \Reg_Bank/registers[31][2] ,
         \Reg_Bank/registers[31][3] , \Reg_Bank/registers[31][4] ,
         \Reg_Bank/registers[31][5] , \Reg_Bank/registers[31][6] ,
         \Reg_Bank/registers[31][7] , \Reg_Bank/registers[31][8] ,
         \Reg_Bank/registers[31][9] , \Reg_Bank/registers[31][10] ,
         \Reg_Bank/registers[31][11] , \Reg_Bank/registers[31][12] ,
         \Reg_Bank/registers[31][13] , \Reg_Bank/registers[31][14] ,
         \Reg_Bank/registers[31][15] , \Reg_Bank/registers[31][16] ,
         \Reg_Bank/registers[31][17] , \Reg_Bank/registers[31][18] ,
         \Reg_Bank/registers[31][19] , \Reg_Bank/registers[31][20] ,
         \Reg_Bank/registers[31][21] , \Reg_Bank/registers[31][22] ,
         \Reg_Bank/registers[31][23] , \Reg_Bank/registers[31][24] ,
         \Reg_Bank/registers[31][25] , \Reg_Bank/registers[31][26] ,
         \Reg_Bank/registers[31][27] , \Reg_Bank/registers[31][28] ,
         \Reg_Bank/registers[31][29] , \Reg_Bank/registers[31][30] ,
         \Reg_Bank/registers[31][31] , \Shifter/N75 ,
         \Shifter/sll_27/ML_int[5][16] , \Shifter/sll_27/ML_int[5][17] ,
         \Shifter/sll_27/ML_int[5][18] , \Shifter/sll_27/ML_int[5][19] ,
         \Shifter/sll_27/ML_int[5][20] , \Shifter/sll_27/ML_int[5][21] ,
         \Shifter/sll_27/ML_int[5][22] , \Shifter/sll_27/ML_int[5][23] ,
         \Shifter/sll_27/ML_int[5][24] , \Shifter/sll_27/ML_int[5][25] ,
         \Shifter/sll_27/ML_int[5][26] , \Shifter/sll_27/ML_int[5][27] ,
         \Shifter/sll_27/ML_int[5][28] , \Shifter/sll_27/ML_int[5][29] ,
         \Shifter/sll_27/ML_int[5][30] , \Shifter/sll_27/ML_int[5][31] ,
         \Shifter/sll_27/ML_int[4][0] , \Shifter/sll_27/ML_int[4][1] ,
         \Shifter/sll_27/ML_int[4][2] , \Shifter/sll_27/ML_int[4][3] ,
         \Shifter/sll_27/ML_int[4][4] , \Shifter/sll_27/ML_int[4][5] ,
         \Shifter/sll_27/ML_int[4][6] , \Shifter/sll_27/ML_int[4][7] ,
         \Shifter/sll_27/ML_int[4][8] , \Shifter/sll_27/ML_int[4][9] ,
         \Shifter/sll_27/ML_int[4][10] , \Shifter/sll_27/ML_int[4][11] ,
         \Shifter/sll_27/ML_int[4][12] , \Shifter/sll_27/ML_int[4][13] ,
         \Shifter/sll_27/ML_int[4][14] , \Shifter/sll_27/ML_int[4][15] ,
         \Shifter/sll_27/ML_int[4][16] , \Shifter/sll_27/ML_int[4][17] ,
         \Shifter/sll_27/ML_int[4][18] , \Shifter/sll_27/ML_int[4][19] ,
         \Shifter/sll_27/ML_int[4][20] , \Shifter/sll_27/ML_int[4][21] ,
         \Shifter/sll_27/ML_int[4][22] , \Shifter/sll_27/ML_int[4][23] ,
         \Shifter/sll_27/ML_int[4][24] , \Shifter/sll_27/ML_int[4][25] ,
         \Shifter/sll_27/ML_int[4][26] , \Shifter/sll_27/ML_int[4][27] ,
         \Shifter/sll_27/ML_int[4][28] , \Shifter/sll_27/ML_int[4][29] ,
         \Shifter/sll_27/ML_int[4][30] , \Shifter/sll_27/ML_int[4][31] ,
         \Shifter/sll_27/ML_int[3][0] , \Shifter/sll_27/ML_int[3][1] ,
         \Shifter/sll_27/ML_int[3][2] , \Shifter/sll_27/ML_int[3][3] ,
         \Shifter/sll_27/ML_int[3][4] , \Shifter/sll_27/ML_int[3][5] ,
         \Shifter/sll_27/ML_int[3][6] , \Shifter/sll_27/ML_int[3][7] ,
         \Shifter/sll_27/ML_int[3][8] , \Shifter/sll_27/ML_int[3][9] ,
         \Shifter/sll_27/ML_int[3][10] , \Shifter/sll_27/ML_int[3][11] ,
         \Shifter/sll_27/ML_int[3][12] , \Shifter/sll_27/ML_int[3][13] ,
         \Shifter/sll_27/ML_int[3][14] , \Shifter/sll_27/ML_int[3][15] ,
         \Shifter/sll_27/ML_int[3][16] , \Shifter/sll_27/ML_int[3][17] ,
         \Shifter/sll_27/ML_int[3][18] , \Shifter/sll_27/ML_int[3][19] ,
         \Shifter/sll_27/ML_int[3][20] , \Shifter/sll_27/ML_int[3][21] ,
         \Shifter/sll_27/ML_int[3][22] , \Shifter/sll_27/ML_int[3][23] ,
         \Shifter/sll_27/ML_int[3][24] , \Shifter/sll_27/ML_int[3][25] ,
         \Shifter/sll_27/ML_int[3][26] , \Shifter/sll_27/ML_int[3][27] ,
         \Shifter/sll_27/ML_int[3][28] , \Shifter/sll_27/ML_int[3][29] ,
         \Shifter/sll_27/ML_int[3][30] , \Shifter/sll_27/ML_int[3][31] ,
         \Shifter/sll_27/ML_int[2][0] , \Shifter/sll_27/ML_int[2][1] ,
         \Shifter/sll_27/ML_int[2][2] , \Shifter/sll_27/ML_int[2][3] ,
         \Shifter/sll_27/ML_int[2][4] , \Shifter/sll_27/ML_int[2][5] ,
         \Shifter/sll_27/ML_int[2][6] , \Shifter/sll_27/ML_int[2][7] ,
         \Shifter/sll_27/ML_int[2][8] , \Shifter/sll_27/ML_int[2][9] ,
         \Shifter/sll_27/ML_int[2][10] , \Shifter/sll_27/ML_int[2][11] ,
         \Shifter/sll_27/ML_int[2][12] , \Shifter/sll_27/ML_int[2][13] ,
         \Shifter/sll_27/ML_int[2][14] , \Shifter/sll_27/ML_int[2][15] ,
         \Shifter/sll_27/ML_int[2][16] , \Shifter/sll_27/ML_int[2][17] ,
         \Shifter/sll_27/ML_int[2][18] , \Shifter/sll_27/ML_int[2][19] ,
         \Shifter/sll_27/ML_int[2][20] , \Shifter/sll_27/ML_int[2][21] ,
         \Shifter/sll_27/ML_int[2][22] , \Shifter/sll_27/ML_int[2][23] ,
         \Shifter/sll_27/ML_int[2][24] , \Shifter/sll_27/ML_int[2][25] ,
         \Shifter/sll_27/ML_int[2][26] , \Shifter/sll_27/ML_int[2][27] ,
         \Shifter/sll_27/ML_int[2][28] , \Shifter/sll_27/ML_int[2][29] ,
         \Shifter/sll_27/ML_int[2][30] , \Shifter/sll_27/ML_int[2][31] ,
         \Shifter/sll_27/ML_int[1][0] , \Shifter/sll_27/ML_int[1][1] ,
         \Shifter/sll_27/ML_int[1][2] , \Shifter/sll_27/ML_int[1][3] ,
         \Shifter/sll_27/ML_int[1][4] , \Shifter/sll_27/ML_int[1][5] ,
         \Shifter/sll_27/ML_int[1][6] , \Shifter/sll_27/ML_int[1][7] ,
         \Shifter/sll_27/ML_int[1][8] , \Shifter/sll_27/ML_int[1][9] ,
         \Shifter/sll_27/ML_int[1][10] , \Shifter/sll_27/ML_int[1][11] ,
         \Shifter/sll_27/ML_int[1][12] , \Shifter/sll_27/ML_int[1][13] ,
         \Shifter/sll_27/ML_int[1][14] , \Shifter/sll_27/ML_int[1][15] ,
         \Shifter/sll_27/ML_int[1][16] , \Shifter/sll_27/ML_int[1][17] ,
         \Shifter/sll_27/ML_int[1][18] , \Shifter/sll_27/ML_int[1][19] ,
         \Shifter/sll_27/ML_int[1][20] , \Shifter/sll_27/ML_int[1][21] ,
         \Shifter/sll_27/ML_int[1][22] , \Shifter/sll_27/ML_int[1][23] ,
         \Shifter/sll_27/ML_int[1][24] , \Shifter/sll_27/ML_int[1][25] ,
         \Shifter/sll_27/ML_int[1][26] , \Shifter/sll_27/ML_int[1][27] ,
         \Shifter/sll_27/ML_int[1][28] , \Shifter/sll_27/ML_int[1][29] ,
         \Shifter/sll_27/ML_int[1][30] , \Shifter/sll_27/ML_int[1][31] ,
         \PC_Next/add_32/carry[29] , \PC_Next/add_32/carry[28] ,
         \PC_Next/add_32/carry[27] , \PC_Next/add_32/carry[26] ,
         \PC_Next/add_32/carry[25] , \PC_Next/add_32/carry[24] ,
         \PC_Next/add_32/carry[23] , \PC_Next/add_32/carry[22] ,
         \PC_Next/add_32/carry[21] , \PC_Next/add_32/carry[20] ,
         \PC_Next/add_32/carry[19] , \PC_Next/add_32/carry[18] ,
         \PC_Next/add_32/carry[17] , \PC_Next/add_32/carry[16] ,
         \PC_Next/add_32/carry[15] , \PC_Next/add_32/carry[14] ,
         \PC_Next/add_32/carry[13] , \PC_Next/add_32/carry[12] ,
         \PC_Next/add_32/carry[11] , \PC_Next/add_32/carry[10] ,
         \PC_Next/add_32/carry[9] , \PC_Next/add_32/carry[8] ,
         \PC_Next/add_32/carry[7] , \PC_Next/add_32/carry[6] ,
         \PC_Next/add_32/carry[5] , \PC_Next/add_32/carry[4] ,
         \PC_Next/add_32/carry[3] , \PC_Next/add_32/carry[2] ,
         \PC_Next/add_48/carry[29] , \PC_Next/add_48/carry[28] ,
         \PC_Next/add_48/carry[27] , \PC_Next/add_48/carry[26] ,
         \PC_Next/add_48/carry[25] , \PC_Next/add_48/carry[24] ,
         \PC_Next/add_48/carry[23] , \PC_Next/add_48/carry[22] ,
         \PC_Next/add_48/carry[21] , \PC_Next/add_48/carry[20] ,
         \PC_Next/add_48/carry[19] , \PC_Next/add_48/carry[18] ,
         \PC_Next/add_48/carry[17] , \PC_Next/add_48/carry[16] ,
         \PC_Next/add_48/carry[15] , \PC_Next/add_48/carry[14] ,
         \PC_Next/add_48/carry[13] , \PC_Next/add_48/carry[12] ,
         \PC_Next/add_48/carry[11] , \PC_Next/add_48/carry[10] ,
         \PC_Next/add_48/carry[9] , \PC_Next/add_48/carry[8] ,
         \PC_Next/add_48/carry[7] , \PC_Next/add_48/carry[6] ,
         \PC_Next/add_48/carry[5] , \PC_Next/add_48/carry[4] ,
         \PC_Next/add_48/carry[3] , \PC_Next/add_48/carry[2] ,
         \PC_Next/add_48/carry[1] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996;
  wire   [31:0] opcode;
  wire   [31:2] pc_current;
  wire   [31:2] pc_plus4;
  wire   [31:0] reg_target;
  wire   [4:0] rs_index;
  wire   [4:0] rt_index;
  wire   [15:0] imm;
  wire   [31:0] reg_source;
  wire   [31:0] a_bus;
  wire   [31:0] b_bus;

  DFF \PC_Next/pc_reg[30]  ( .D(\PC_Next/n309 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[30]) );
  DFF \PC_Next/pc_reg[29]  ( .D(\PC_Next/n310 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[29]) );
  DFF \PC_Next/pc_reg[28]  ( .D(\PC_Next/n311 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[28]) );
  DFF \PC_Next/pc_reg[27]  ( .D(\PC_Next/pc_future[27] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[27]) );
  DFF \PC_Next/pc_reg[26]  ( .D(\PC_Next/pc_future[26] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[26]) );
  DFF \PC_Next/pc_reg[25]  ( .D(\PC_Next/pc_future[25] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[25]) );
  DFF \PC_Next/pc_reg[24]  ( .D(\PC_Next/pc_future[24] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[24]) );
  DFF \PC_Next/pc_reg[23]  ( .D(\PC_Next/pc_future[23] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[23]) );
  DFF \PC_Next/pc_reg[22]  ( .D(\PC_Next/pc_future[22] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[22]) );
  DFF \PC_Next/pc_reg[21]  ( .D(\PC_Next/pc_future[21] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[21]) );
  DFF \PC_Next/pc_reg[20]  ( .D(\PC_Next/pc_future[20] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[20]) );
  DFF \PC_Next/pc_reg[19]  ( .D(\PC_Next/pc_future[19] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[19]) );
  DFF \PC_Next/pc_reg[18]  ( .D(\PC_Next/pc_future[18] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[18]) );
  DFF \PC_Next/pc_reg[17]  ( .D(\PC_Next/pc_future[17] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[17]) );
  DFF \PC_Next/pc_reg[16]  ( .D(\PC_Next/pc_future[16] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[16]) );
  DFF \PC_Next/pc_reg[15]  ( .D(\PC_Next/pc_future[15] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[15]) );
  DFF \PC_Next/pc_reg[14]  ( .D(\PC_Next/pc_future[14] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[14]) );
  DFF \PC_Next/pc_reg[13]  ( .D(\PC_Next/pc_future[13] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[13]) );
  DFF \PC_Next/pc_reg[12]  ( .D(\PC_Next/pc_future[12] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[12]) );
  DFF \PC_Next/pc_reg[11]  ( .D(\PC_Next/pc_future[11] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[11]) );
  DFF \PC_Next/pc_reg[10]  ( .D(\PC_Next/pc_future[10] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[10]) );
  DFF \PC_Next/pc_reg[9]  ( .D(\PC_Next/pc_future[9] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[9]) );
  DFF \PC_Next/pc_reg[8]  ( .D(\PC_Next/pc_future[8] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[8]) );
  DFF \PC_Next/pc_reg[7]  ( .D(\PC_Next/pc_future[7] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[7]) );
  DFF \PC_Next/pc_reg[6]  ( .D(\PC_Next/pc_future[6] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[6]) );
  DFF \PC_Next/pc_reg[5]  ( .D(\PC_Next/pc_future[5] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[5]) );
  DFF \PC_Next/pc_reg[4]  ( .D(\PC_Next/pc_future[4] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[4]) );
  DFF \PC_Next/pc_reg[3]  ( .D(\PC_Next/pc_future[3] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[3]) );
  DFF \PC_Next/pc_reg[31]  ( .D(\PC_Next/n308 ), .CLK(clk), .RST(rst), .I(1'b0), .Q(pc_current[31]) );
  DFF \PC_Next/pc_reg[2]  ( .D(\PC_Next/pc_future[2] ), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(pc_current[2]) );
  MUX \Inst_Mem/U2019  ( .IN0(\Inst_Mem/n1984 ), .IN1(\Inst_Mem/n1953 ), .SEL(
        pc_current[7]), .F(opcode[31]) );
  MUX \Inst_Mem/U2018  ( .IN0(\Inst_Mem/n1983 ), .IN1(\Inst_Mem/n1968 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1984 ) );
  MUX \Inst_Mem/U2017  ( .IN0(\Inst_Mem/n1982 ), .IN1(\Inst_Mem/n1975 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1983 ) );
  MUX \Inst_Mem/U2016  ( .IN0(\Inst_Mem/n1981 ), .IN1(\Inst_Mem/n1978 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1982 ) );
  MUX \Inst_Mem/U2015  ( .IN0(\Inst_Mem/n1980 ), .IN1(\Inst_Mem/n1979 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1981 ) );
  MUX \Inst_Mem/U2014  ( .IN0(\Inst_Mem/inst_mem_reg[0][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1980 ) );
  MUX \Inst_Mem/U2013  ( .IN0(\Inst_Mem/inst_mem_reg[2][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1979 ) );
  MUX \Inst_Mem/U2012  ( .IN0(\Inst_Mem/n1977 ), .IN1(\Inst_Mem/n1976 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1978 ) );
  MUX \Inst_Mem/U2011  ( .IN0(\Inst_Mem/inst_mem_reg[4][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1977 ) );
  MUX \Inst_Mem/U2010  ( .IN0(\Inst_Mem/inst_mem_reg[6][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1976 ) );
  MUX \Inst_Mem/U2009  ( .IN0(\Inst_Mem/n1974 ), .IN1(\Inst_Mem/n1971 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1975 ) );
  MUX \Inst_Mem/U2008  ( .IN0(\Inst_Mem/n1973 ), .IN1(\Inst_Mem/n1972 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1974 ) );
  MUX \Inst_Mem/U2007  ( .IN0(\Inst_Mem/inst_mem_reg[8][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1973 ) );
  MUX \Inst_Mem/U2006  ( .IN0(\Inst_Mem/inst_mem_reg[10][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1972 ) );
  MUX \Inst_Mem/U2005  ( .IN0(\Inst_Mem/n1970 ), .IN1(\Inst_Mem/n1969 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1971 ) );
  MUX \Inst_Mem/U2004  ( .IN0(\Inst_Mem/inst_mem_reg[12][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1970 ) );
  MUX \Inst_Mem/U2003  ( .IN0(\Inst_Mem/inst_mem_reg[14][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1969 ) );
  MUX \Inst_Mem/U2002  ( .IN0(\Inst_Mem/n1967 ), .IN1(\Inst_Mem/n1960 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1968 ) );
  MUX \Inst_Mem/U2001  ( .IN0(\Inst_Mem/n1966 ), .IN1(\Inst_Mem/n1963 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1967 ) );
  MUX \Inst_Mem/U2000  ( .IN0(\Inst_Mem/n1965 ), .IN1(\Inst_Mem/n1964 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1966 ) );
  MUX \Inst_Mem/U1999  ( .IN0(\Inst_Mem/inst_mem_reg[16][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1965 ) );
  MUX \Inst_Mem/U1998  ( .IN0(\Inst_Mem/inst_mem_reg[18][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1964 ) );
  MUX \Inst_Mem/U1997  ( .IN0(\Inst_Mem/n1962 ), .IN1(\Inst_Mem/n1961 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1963 ) );
  MUX \Inst_Mem/U1996  ( .IN0(\Inst_Mem/inst_mem_reg[20][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1962 ) );
  MUX \Inst_Mem/U1995  ( .IN0(\Inst_Mem/inst_mem_reg[22][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1961 ) );
  MUX \Inst_Mem/U1994  ( .IN0(\Inst_Mem/n1959 ), .IN1(\Inst_Mem/n1956 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1960 ) );
  MUX \Inst_Mem/U1993  ( .IN0(\Inst_Mem/n1958 ), .IN1(\Inst_Mem/n1957 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1959 ) );
  MUX \Inst_Mem/U1992  ( .IN0(\Inst_Mem/inst_mem_reg[24][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1958 ) );
  MUX \Inst_Mem/U1991  ( .IN0(\Inst_Mem/inst_mem_reg[26][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1957 ) );
  MUX \Inst_Mem/U1990  ( .IN0(\Inst_Mem/n1955 ), .IN1(\Inst_Mem/n1954 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1956 ) );
  MUX \Inst_Mem/U1989  ( .IN0(\Inst_Mem/inst_mem_reg[28][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1955 ) );
  MUX \Inst_Mem/U1988  ( .IN0(\Inst_Mem/inst_mem_reg[30][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1954 ) );
  MUX \Inst_Mem/U1987  ( .IN0(\Inst_Mem/n1952 ), .IN1(\Inst_Mem/n1937 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1953 ) );
  MUX \Inst_Mem/U1986  ( .IN0(\Inst_Mem/n1951 ), .IN1(\Inst_Mem/n1944 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1952 ) );
  MUX \Inst_Mem/U1985  ( .IN0(\Inst_Mem/n1950 ), .IN1(\Inst_Mem/n1947 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1951 ) );
  MUX \Inst_Mem/U1984  ( .IN0(\Inst_Mem/n1949 ), .IN1(\Inst_Mem/n1948 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1950 ) );
  MUX \Inst_Mem/U1983  ( .IN0(\Inst_Mem/inst_mem_reg[32][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1949 ) );
  MUX \Inst_Mem/U1982  ( .IN0(\Inst_Mem/inst_mem_reg[34][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1948 ) );
  MUX \Inst_Mem/U1981  ( .IN0(\Inst_Mem/n1946 ), .IN1(\Inst_Mem/n1945 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1947 ) );
  MUX \Inst_Mem/U1980  ( .IN0(\Inst_Mem/inst_mem_reg[36][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1946 ) );
  MUX \Inst_Mem/U1979  ( .IN0(\Inst_Mem/inst_mem_reg[38][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1945 ) );
  MUX \Inst_Mem/U1978  ( .IN0(\Inst_Mem/n1943 ), .IN1(\Inst_Mem/n1940 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1944 ) );
  MUX \Inst_Mem/U1977  ( .IN0(\Inst_Mem/n1942 ), .IN1(\Inst_Mem/n1941 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1943 ) );
  MUX \Inst_Mem/U1976  ( .IN0(\Inst_Mem/inst_mem_reg[40][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1942 ) );
  MUX \Inst_Mem/U1975  ( .IN0(\Inst_Mem/inst_mem_reg[42][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1941 ) );
  MUX \Inst_Mem/U1974  ( .IN0(\Inst_Mem/n1939 ), .IN1(\Inst_Mem/n1938 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1940 ) );
  MUX \Inst_Mem/U1973  ( .IN0(\Inst_Mem/inst_mem_reg[44][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1939 ) );
  MUX \Inst_Mem/U1972  ( .IN0(\Inst_Mem/inst_mem_reg[46][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1938 ) );
  MUX \Inst_Mem/U1971  ( .IN0(\Inst_Mem/n1936 ), .IN1(\Inst_Mem/n1929 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1937 ) );
  MUX \Inst_Mem/U1970  ( .IN0(\Inst_Mem/n1935 ), .IN1(\Inst_Mem/n1932 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1936 ) );
  MUX \Inst_Mem/U1969  ( .IN0(\Inst_Mem/n1934 ), .IN1(\Inst_Mem/n1933 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1935 ) );
  MUX \Inst_Mem/U1968  ( .IN0(\Inst_Mem/inst_mem_reg[48][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1934 ) );
  MUX \Inst_Mem/U1967  ( .IN0(\Inst_Mem/inst_mem_reg[50][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1933 ) );
  MUX \Inst_Mem/U1966  ( .IN0(\Inst_Mem/n1931 ), .IN1(\Inst_Mem/n1930 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1932 ) );
  MUX \Inst_Mem/U1965  ( .IN0(\Inst_Mem/inst_mem_reg[52][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1931 ) );
  MUX \Inst_Mem/U1964  ( .IN0(\Inst_Mem/inst_mem_reg[54][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1930 ) );
  MUX \Inst_Mem/U1963  ( .IN0(\Inst_Mem/n1928 ), .IN1(\Inst_Mem/n1925 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1929 ) );
  MUX \Inst_Mem/U1962  ( .IN0(\Inst_Mem/n1927 ), .IN1(\Inst_Mem/n1926 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1928 ) );
  MUX \Inst_Mem/U1961  ( .IN0(\Inst_Mem/inst_mem_reg[56][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1927 ) );
  MUX \Inst_Mem/U1960  ( .IN0(\Inst_Mem/inst_mem_reg[58][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1926 ) );
  MUX \Inst_Mem/U1959  ( .IN0(\Inst_Mem/n1924 ), .IN1(\Inst_Mem/n1923 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1925 ) );
  MUX \Inst_Mem/U1958  ( .IN0(\Inst_Mem/inst_mem_reg[60][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1924 ) );
  MUX \Inst_Mem/U1957  ( .IN0(\Inst_Mem/inst_mem_reg[62][31] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][31] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1923 ) );
  MUX \Inst_Mem/U1956  ( .IN0(\Inst_Mem/n1922 ), .IN1(\Inst_Mem/n1891 ), .SEL(
        pc_current[7]), .F(opcode[30]) );
  MUX \Inst_Mem/U1955  ( .IN0(\Inst_Mem/n1921 ), .IN1(\Inst_Mem/n1906 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1922 ) );
  MUX \Inst_Mem/U1954  ( .IN0(\Inst_Mem/n1920 ), .IN1(\Inst_Mem/n1913 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1921 ) );
  MUX \Inst_Mem/U1953  ( .IN0(\Inst_Mem/n1919 ), .IN1(\Inst_Mem/n1916 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1920 ) );
  MUX \Inst_Mem/U1952  ( .IN0(\Inst_Mem/n1918 ), .IN1(\Inst_Mem/n1917 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1919 ) );
  MUX \Inst_Mem/U1951  ( .IN0(\Inst_Mem/inst_mem_reg[0][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1918 ) );
  MUX \Inst_Mem/U1950  ( .IN0(\Inst_Mem/inst_mem_reg[2][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1917 ) );
  MUX \Inst_Mem/U1949  ( .IN0(\Inst_Mem/n1915 ), .IN1(\Inst_Mem/n1914 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1916 ) );
  MUX \Inst_Mem/U1948  ( .IN0(\Inst_Mem/inst_mem_reg[4][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1915 ) );
  MUX \Inst_Mem/U1947  ( .IN0(\Inst_Mem/inst_mem_reg[6][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1914 ) );
  MUX \Inst_Mem/U1946  ( .IN0(\Inst_Mem/n1912 ), .IN1(\Inst_Mem/n1909 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1913 ) );
  MUX \Inst_Mem/U1945  ( .IN0(\Inst_Mem/n1911 ), .IN1(\Inst_Mem/n1910 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1912 ) );
  MUX \Inst_Mem/U1944  ( .IN0(\Inst_Mem/inst_mem_reg[8][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1911 ) );
  MUX \Inst_Mem/U1943  ( .IN0(\Inst_Mem/inst_mem_reg[10][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1910 ) );
  MUX \Inst_Mem/U1942  ( .IN0(\Inst_Mem/n1908 ), .IN1(\Inst_Mem/n1907 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1909 ) );
  MUX \Inst_Mem/U1941  ( .IN0(\Inst_Mem/inst_mem_reg[12][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1908 ) );
  MUX \Inst_Mem/U1940  ( .IN0(\Inst_Mem/inst_mem_reg[14][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1907 ) );
  MUX \Inst_Mem/U1939  ( .IN0(\Inst_Mem/n1905 ), .IN1(\Inst_Mem/n1898 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1906 ) );
  MUX \Inst_Mem/U1938  ( .IN0(\Inst_Mem/n1904 ), .IN1(\Inst_Mem/n1901 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1905 ) );
  MUX \Inst_Mem/U1937  ( .IN0(\Inst_Mem/n1903 ), .IN1(\Inst_Mem/n1902 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1904 ) );
  MUX \Inst_Mem/U1936  ( .IN0(\Inst_Mem/inst_mem_reg[16][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1903 ) );
  MUX \Inst_Mem/U1935  ( .IN0(\Inst_Mem/inst_mem_reg[18][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1902 ) );
  MUX \Inst_Mem/U1934  ( .IN0(\Inst_Mem/n1900 ), .IN1(\Inst_Mem/n1899 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1901 ) );
  MUX \Inst_Mem/U1933  ( .IN0(\Inst_Mem/inst_mem_reg[20][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1900 ) );
  MUX \Inst_Mem/U1932  ( .IN0(\Inst_Mem/inst_mem_reg[22][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1899 ) );
  MUX \Inst_Mem/U1931  ( .IN0(\Inst_Mem/n1897 ), .IN1(\Inst_Mem/n1894 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1898 ) );
  MUX \Inst_Mem/U1930  ( .IN0(\Inst_Mem/n1896 ), .IN1(\Inst_Mem/n1895 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1897 ) );
  MUX \Inst_Mem/U1929  ( .IN0(\Inst_Mem/inst_mem_reg[24][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1896 ) );
  MUX \Inst_Mem/U1928  ( .IN0(\Inst_Mem/inst_mem_reg[26][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1895 ) );
  MUX \Inst_Mem/U1927  ( .IN0(\Inst_Mem/n1893 ), .IN1(\Inst_Mem/n1892 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1894 ) );
  MUX \Inst_Mem/U1926  ( .IN0(\Inst_Mem/inst_mem_reg[28][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1893 ) );
  MUX \Inst_Mem/U1925  ( .IN0(\Inst_Mem/inst_mem_reg[30][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1892 ) );
  MUX \Inst_Mem/U1924  ( .IN0(\Inst_Mem/n1890 ), .IN1(\Inst_Mem/n1875 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1891 ) );
  MUX \Inst_Mem/U1923  ( .IN0(\Inst_Mem/n1889 ), .IN1(\Inst_Mem/n1882 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1890 ) );
  MUX \Inst_Mem/U1922  ( .IN0(\Inst_Mem/n1888 ), .IN1(\Inst_Mem/n1885 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1889 ) );
  MUX \Inst_Mem/U1921  ( .IN0(\Inst_Mem/n1887 ), .IN1(\Inst_Mem/n1886 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1888 ) );
  MUX \Inst_Mem/U1920  ( .IN0(\Inst_Mem/inst_mem_reg[32][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1887 ) );
  MUX \Inst_Mem/U1919  ( .IN0(\Inst_Mem/inst_mem_reg[34][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1886 ) );
  MUX \Inst_Mem/U1918  ( .IN0(\Inst_Mem/n1884 ), .IN1(\Inst_Mem/n1883 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1885 ) );
  MUX \Inst_Mem/U1917  ( .IN0(\Inst_Mem/inst_mem_reg[36][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1884 ) );
  MUX \Inst_Mem/U1916  ( .IN0(\Inst_Mem/inst_mem_reg[38][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1883 ) );
  MUX \Inst_Mem/U1915  ( .IN0(\Inst_Mem/n1881 ), .IN1(\Inst_Mem/n1878 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1882 ) );
  MUX \Inst_Mem/U1914  ( .IN0(\Inst_Mem/n1880 ), .IN1(\Inst_Mem/n1879 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1881 ) );
  MUX \Inst_Mem/U1913  ( .IN0(\Inst_Mem/inst_mem_reg[40][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1880 ) );
  MUX \Inst_Mem/U1912  ( .IN0(\Inst_Mem/inst_mem_reg[42][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1879 ) );
  MUX \Inst_Mem/U1911  ( .IN0(\Inst_Mem/n1877 ), .IN1(\Inst_Mem/n1876 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1878 ) );
  MUX \Inst_Mem/U1910  ( .IN0(\Inst_Mem/inst_mem_reg[44][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1877 ) );
  MUX \Inst_Mem/U1909  ( .IN0(\Inst_Mem/inst_mem_reg[46][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1876 ) );
  MUX \Inst_Mem/U1908  ( .IN0(\Inst_Mem/n1874 ), .IN1(\Inst_Mem/n1867 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1875 ) );
  MUX \Inst_Mem/U1907  ( .IN0(\Inst_Mem/n1873 ), .IN1(\Inst_Mem/n1870 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1874 ) );
  MUX \Inst_Mem/U1906  ( .IN0(\Inst_Mem/n1872 ), .IN1(\Inst_Mem/n1871 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1873 ) );
  MUX \Inst_Mem/U1905  ( .IN0(\Inst_Mem/inst_mem_reg[48][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1872 ) );
  MUX \Inst_Mem/U1904  ( .IN0(\Inst_Mem/inst_mem_reg[50][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1871 ) );
  MUX \Inst_Mem/U1903  ( .IN0(\Inst_Mem/n1869 ), .IN1(\Inst_Mem/n1868 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1870 ) );
  MUX \Inst_Mem/U1902  ( .IN0(\Inst_Mem/inst_mem_reg[52][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1869 ) );
  MUX \Inst_Mem/U1901  ( .IN0(\Inst_Mem/inst_mem_reg[54][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1868 ) );
  MUX \Inst_Mem/U1900  ( .IN0(\Inst_Mem/n1866 ), .IN1(\Inst_Mem/n1863 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1867 ) );
  MUX \Inst_Mem/U1899  ( .IN0(\Inst_Mem/n1865 ), .IN1(\Inst_Mem/n1864 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1866 ) );
  MUX \Inst_Mem/U1898  ( .IN0(\Inst_Mem/inst_mem_reg[56][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1865 ) );
  MUX \Inst_Mem/U1897  ( .IN0(\Inst_Mem/inst_mem_reg[58][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1864 ) );
  MUX \Inst_Mem/U1896  ( .IN0(\Inst_Mem/n1862 ), .IN1(\Inst_Mem/n1861 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1863 ) );
  MUX \Inst_Mem/U1895  ( .IN0(\Inst_Mem/inst_mem_reg[60][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1862 ) );
  MUX \Inst_Mem/U1894  ( .IN0(\Inst_Mem/inst_mem_reg[62][30] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][30] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1861 ) );
  MUX \Inst_Mem/U1893  ( .IN0(\Inst_Mem/n1860 ), .IN1(\Inst_Mem/n1829 ), .SEL(
        pc_current[7]), .F(opcode[29]) );
  MUX \Inst_Mem/U1892  ( .IN0(\Inst_Mem/n1859 ), .IN1(\Inst_Mem/n1844 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1860 ) );
  MUX \Inst_Mem/U1891  ( .IN0(\Inst_Mem/n1858 ), .IN1(\Inst_Mem/n1851 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1859 ) );
  MUX \Inst_Mem/U1890  ( .IN0(\Inst_Mem/n1857 ), .IN1(\Inst_Mem/n1854 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1858 ) );
  MUX \Inst_Mem/U1889  ( .IN0(\Inst_Mem/n1856 ), .IN1(\Inst_Mem/n1855 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1857 ) );
  MUX \Inst_Mem/U1888  ( .IN0(\Inst_Mem/inst_mem_reg[0][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1856 ) );
  MUX \Inst_Mem/U1887  ( .IN0(\Inst_Mem/inst_mem_reg[2][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1855 ) );
  MUX \Inst_Mem/U1886  ( .IN0(\Inst_Mem/n1853 ), .IN1(\Inst_Mem/n1852 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1854 ) );
  MUX \Inst_Mem/U1885  ( .IN0(\Inst_Mem/inst_mem_reg[4][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1853 ) );
  MUX \Inst_Mem/U1884  ( .IN0(\Inst_Mem/inst_mem_reg[6][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1852 ) );
  MUX \Inst_Mem/U1883  ( .IN0(\Inst_Mem/n1850 ), .IN1(\Inst_Mem/n1847 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1851 ) );
  MUX \Inst_Mem/U1882  ( .IN0(\Inst_Mem/n1849 ), .IN1(\Inst_Mem/n1848 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1850 ) );
  MUX \Inst_Mem/U1881  ( .IN0(\Inst_Mem/inst_mem_reg[8][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1849 ) );
  MUX \Inst_Mem/U1880  ( .IN0(\Inst_Mem/inst_mem_reg[10][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1848 ) );
  MUX \Inst_Mem/U1879  ( .IN0(\Inst_Mem/n1846 ), .IN1(\Inst_Mem/n1845 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1847 ) );
  MUX \Inst_Mem/U1878  ( .IN0(\Inst_Mem/inst_mem_reg[12][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1846 ) );
  MUX \Inst_Mem/U1877  ( .IN0(\Inst_Mem/inst_mem_reg[14][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1845 ) );
  MUX \Inst_Mem/U1876  ( .IN0(\Inst_Mem/n1843 ), .IN1(\Inst_Mem/n1836 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1844 ) );
  MUX \Inst_Mem/U1875  ( .IN0(\Inst_Mem/n1842 ), .IN1(\Inst_Mem/n1839 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1843 ) );
  MUX \Inst_Mem/U1874  ( .IN0(\Inst_Mem/n1841 ), .IN1(\Inst_Mem/n1840 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1842 ) );
  MUX \Inst_Mem/U1873  ( .IN0(\Inst_Mem/inst_mem_reg[16][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1841 ) );
  MUX \Inst_Mem/U1872  ( .IN0(\Inst_Mem/inst_mem_reg[18][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1840 ) );
  MUX \Inst_Mem/U1871  ( .IN0(\Inst_Mem/n1838 ), .IN1(\Inst_Mem/n1837 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1839 ) );
  MUX \Inst_Mem/U1870  ( .IN0(\Inst_Mem/inst_mem_reg[20][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1838 ) );
  MUX \Inst_Mem/U1869  ( .IN0(\Inst_Mem/inst_mem_reg[22][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1837 ) );
  MUX \Inst_Mem/U1868  ( .IN0(\Inst_Mem/n1835 ), .IN1(\Inst_Mem/n1832 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1836 ) );
  MUX \Inst_Mem/U1867  ( .IN0(\Inst_Mem/n1834 ), .IN1(\Inst_Mem/n1833 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1835 ) );
  MUX \Inst_Mem/U1866  ( .IN0(\Inst_Mem/inst_mem_reg[24][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1834 ) );
  MUX \Inst_Mem/U1865  ( .IN0(\Inst_Mem/inst_mem_reg[26][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1833 ) );
  MUX \Inst_Mem/U1864  ( .IN0(\Inst_Mem/n1831 ), .IN1(\Inst_Mem/n1830 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1832 ) );
  MUX \Inst_Mem/U1863  ( .IN0(\Inst_Mem/inst_mem_reg[28][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1831 ) );
  MUX \Inst_Mem/U1862  ( .IN0(\Inst_Mem/inst_mem_reg[30][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1830 ) );
  MUX \Inst_Mem/U1861  ( .IN0(\Inst_Mem/n1828 ), .IN1(\Inst_Mem/n1813 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1829 ) );
  MUX \Inst_Mem/U1860  ( .IN0(\Inst_Mem/n1827 ), .IN1(\Inst_Mem/n1820 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1828 ) );
  MUX \Inst_Mem/U1859  ( .IN0(\Inst_Mem/n1826 ), .IN1(\Inst_Mem/n1823 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1827 ) );
  MUX \Inst_Mem/U1858  ( .IN0(\Inst_Mem/n1825 ), .IN1(\Inst_Mem/n1824 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1826 ) );
  MUX \Inst_Mem/U1857  ( .IN0(\Inst_Mem/inst_mem_reg[32][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1825 ) );
  MUX \Inst_Mem/U1856  ( .IN0(\Inst_Mem/inst_mem_reg[34][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1824 ) );
  MUX \Inst_Mem/U1855  ( .IN0(\Inst_Mem/n1822 ), .IN1(\Inst_Mem/n1821 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1823 ) );
  MUX \Inst_Mem/U1854  ( .IN0(\Inst_Mem/inst_mem_reg[36][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1822 ) );
  MUX \Inst_Mem/U1853  ( .IN0(\Inst_Mem/inst_mem_reg[38][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1821 ) );
  MUX \Inst_Mem/U1852  ( .IN0(\Inst_Mem/n1819 ), .IN1(\Inst_Mem/n1816 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1820 ) );
  MUX \Inst_Mem/U1851  ( .IN0(\Inst_Mem/n1818 ), .IN1(\Inst_Mem/n1817 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1819 ) );
  MUX \Inst_Mem/U1850  ( .IN0(\Inst_Mem/inst_mem_reg[40][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1818 ) );
  MUX \Inst_Mem/U1849  ( .IN0(\Inst_Mem/inst_mem_reg[42][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1817 ) );
  MUX \Inst_Mem/U1848  ( .IN0(\Inst_Mem/n1815 ), .IN1(\Inst_Mem/n1814 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1816 ) );
  MUX \Inst_Mem/U1847  ( .IN0(\Inst_Mem/inst_mem_reg[44][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1815 ) );
  MUX \Inst_Mem/U1846  ( .IN0(\Inst_Mem/inst_mem_reg[46][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1814 ) );
  MUX \Inst_Mem/U1845  ( .IN0(\Inst_Mem/n1812 ), .IN1(\Inst_Mem/n1805 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1813 ) );
  MUX \Inst_Mem/U1844  ( .IN0(\Inst_Mem/n1811 ), .IN1(\Inst_Mem/n1808 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1812 ) );
  MUX \Inst_Mem/U1843  ( .IN0(\Inst_Mem/n1810 ), .IN1(\Inst_Mem/n1809 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1811 ) );
  MUX \Inst_Mem/U1842  ( .IN0(\Inst_Mem/inst_mem_reg[48][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1810 ) );
  MUX \Inst_Mem/U1841  ( .IN0(\Inst_Mem/inst_mem_reg[50][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1809 ) );
  MUX \Inst_Mem/U1840  ( .IN0(\Inst_Mem/n1807 ), .IN1(\Inst_Mem/n1806 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1808 ) );
  MUX \Inst_Mem/U1839  ( .IN0(\Inst_Mem/inst_mem_reg[52][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1807 ) );
  MUX \Inst_Mem/U1838  ( .IN0(\Inst_Mem/inst_mem_reg[54][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1806 ) );
  MUX \Inst_Mem/U1837  ( .IN0(\Inst_Mem/n1804 ), .IN1(\Inst_Mem/n1801 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1805 ) );
  MUX \Inst_Mem/U1836  ( .IN0(\Inst_Mem/n1803 ), .IN1(\Inst_Mem/n1802 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1804 ) );
  MUX \Inst_Mem/U1835  ( .IN0(\Inst_Mem/inst_mem_reg[56][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1803 ) );
  MUX \Inst_Mem/U1834  ( .IN0(\Inst_Mem/inst_mem_reg[58][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1802 ) );
  MUX \Inst_Mem/U1833  ( .IN0(\Inst_Mem/n1800 ), .IN1(\Inst_Mem/n1799 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1801 ) );
  MUX \Inst_Mem/U1832  ( .IN0(\Inst_Mem/inst_mem_reg[60][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1800 ) );
  MUX \Inst_Mem/U1831  ( .IN0(\Inst_Mem/inst_mem_reg[62][29] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][29] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1799 ) );
  MUX \Inst_Mem/U1830  ( .IN0(\Inst_Mem/n1798 ), .IN1(\Inst_Mem/n1767 ), .SEL(
        pc_current[7]), .F(opcode[28]) );
  MUX \Inst_Mem/U1829  ( .IN0(\Inst_Mem/n1797 ), .IN1(\Inst_Mem/n1782 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1798 ) );
  MUX \Inst_Mem/U1828  ( .IN0(\Inst_Mem/n1796 ), .IN1(\Inst_Mem/n1789 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1797 ) );
  MUX \Inst_Mem/U1827  ( .IN0(\Inst_Mem/n1795 ), .IN1(\Inst_Mem/n1792 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1796 ) );
  MUX \Inst_Mem/U1826  ( .IN0(\Inst_Mem/n1794 ), .IN1(\Inst_Mem/n1793 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1795 ) );
  MUX \Inst_Mem/U1825  ( .IN0(\Inst_Mem/inst_mem_reg[0][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1794 ) );
  MUX \Inst_Mem/U1824  ( .IN0(\Inst_Mem/inst_mem_reg[2][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1793 ) );
  MUX \Inst_Mem/U1823  ( .IN0(\Inst_Mem/n1791 ), .IN1(\Inst_Mem/n1790 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1792 ) );
  MUX \Inst_Mem/U1822  ( .IN0(\Inst_Mem/inst_mem_reg[4][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1791 ) );
  MUX \Inst_Mem/U1821  ( .IN0(\Inst_Mem/inst_mem_reg[6][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1790 ) );
  MUX \Inst_Mem/U1820  ( .IN0(\Inst_Mem/n1788 ), .IN1(\Inst_Mem/n1785 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1789 ) );
  MUX \Inst_Mem/U1819  ( .IN0(\Inst_Mem/n1787 ), .IN1(\Inst_Mem/n1786 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1788 ) );
  MUX \Inst_Mem/U1818  ( .IN0(\Inst_Mem/inst_mem_reg[8][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1787 ) );
  MUX \Inst_Mem/U1817  ( .IN0(\Inst_Mem/inst_mem_reg[10][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1786 ) );
  MUX \Inst_Mem/U1816  ( .IN0(\Inst_Mem/n1784 ), .IN1(\Inst_Mem/n1783 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1785 ) );
  MUX \Inst_Mem/U1815  ( .IN0(\Inst_Mem/inst_mem_reg[12][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1784 ) );
  MUX \Inst_Mem/U1814  ( .IN0(\Inst_Mem/inst_mem_reg[14][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1783 ) );
  MUX \Inst_Mem/U1813  ( .IN0(\Inst_Mem/n1781 ), .IN1(\Inst_Mem/n1774 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1782 ) );
  MUX \Inst_Mem/U1812  ( .IN0(\Inst_Mem/n1780 ), .IN1(\Inst_Mem/n1777 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1781 ) );
  MUX \Inst_Mem/U1811  ( .IN0(\Inst_Mem/n1779 ), .IN1(\Inst_Mem/n1778 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1780 ) );
  MUX \Inst_Mem/U1810  ( .IN0(\Inst_Mem/inst_mem_reg[16][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1779 ) );
  MUX \Inst_Mem/U1809  ( .IN0(\Inst_Mem/inst_mem_reg[18][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1778 ) );
  MUX \Inst_Mem/U1808  ( .IN0(\Inst_Mem/n1776 ), .IN1(\Inst_Mem/n1775 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1777 ) );
  MUX \Inst_Mem/U1807  ( .IN0(\Inst_Mem/inst_mem_reg[20][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1776 ) );
  MUX \Inst_Mem/U1806  ( .IN0(\Inst_Mem/inst_mem_reg[22][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1775 ) );
  MUX \Inst_Mem/U1805  ( .IN0(\Inst_Mem/n1773 ), .IN1(\Inst_Mem/n1770 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1774 ) );
  MUX \Inst_Mem/U1804  ( .IN0(\Inst_Mem/n1772 ), .IN1(\Inst_Mem/n1771 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1773 ) );
  MUX \Inst_Mem/U1803  ( .IN0(\Inst_Mem/inst_mem_reg[24][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1772 ) );
  MUX \Inst_Mem/U1802  ( .IN0(\Inst_Mem/inst_mem_reg[26][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1771 ) );
  MUX \Inst_Mem/U1801  ( .IN0(\Inst_Mem/n1769 ), .IN1(\Inst_Mem/n1768 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1770 ) );
  MUX \Inst_Mem/U1800  ( .IN0(\Inst_Mem/inst_mem_reg[28][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1769 ) );
  MUX \Inst_Mem/U1799  ( .IN0(\Inst_Mem/inst_mem_reg[30][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1768 ) );
  MUX \Inst_Mem/U1798  ( .IN0(\Inst_Mem/n1766 ), .IN1(\Inst_Mem/n1751 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1767 ) );
  MUX \Inst_Mem/U1797  ( .IN0(\Inst_Mem/n1765 ), .IN1(\Inst_Mem/n1758 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1766 ) );
  MUX \Inst_Mem/U1796  ( .IN0(\Inst_Mem/n1764 ), .IN1(\Inst_Mem/n1761 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1765 ) );
  MUX \Inst_Mem/U1795  ( .IN0(\Inst_Mem/n1763 ), .IN1(\Inst_Mem/n1762 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1764 ) );
  MUX \Inst_Mem/U1794  ( .IN0(\Inst_Mem/inst_mem_reg[32][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1763 ) );
  MUX \Inst_Mem/U1793  ( .IN0(\Inst_Mem/inst_mem_reg[34][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1762 ) );
  MUX \Inst_Mem/U1792  ( .IN0(\Inst_Mem/n1760 ), .IN1(\Inst_Mem/n1759 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1761 ) );
  MUX \Inst_Mem/U1791  ( .IN0(\Inst_Mem/inst_mem_reg[36][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1760 ) );
  MUX \Inst_Mem/U1790  ( .IN0(\Inst_Mem/inst_mem_reg[38][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1759 ) );
  MUX \Inst_Mem/U1789  ( .IN0(\Inst_Mem/n1757 ), .IN1(\Inst_Mem/n1754 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1758 ) );
  MUX \Inst_Mem/U1788  ( .IN0(\Inst_Mem/n1756 ), .IN1(\Inst_Mem/n1755 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1757 ) );
  MUX \Inst_Mem/U1787  ( .IN0(\Inst_Mem/inst_mem_reg[40][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1756 ) );
  MUX \Inst_Mem/U1786  ( .IN0(\Inst_Mem/inst_mem_reg[42][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1755 ) );
  MUX \Inst_Mem/U1785  ( .IN0(\Inst_Mem/n1753 ), .IN1(\Inst_Mem/n1752 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1754 ) );
  MUX \Inst_Mem/U1784  ( .IN0(\Inst_Mem/inst_mem_reg[44][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1753 ) );
  MUX \Inst_Mem/U1783  ( .IN0(\Inst_Mem/inst_mem_reg[46][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1752 ) );
  MUX \Inst_Mem/U1782  ( .IN0(\Inst_Mem/n1750 ), .IN1(\Inst_Mem/n1743 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1751 ) );
  MUX \Inst_Mem/U1781  ( .IN0(\Inst_Mem/n1749 ), .IN1(\Inst_Mem/n1746 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1750 ) );
  MUX \Inst_Mem/U1780  ( .IN0(\Inst_Mem/n1748 ), .IN1(\Inst_Mem/n1747 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1749 ) );
  MUX \Inst_Mem/U1779  ( .IN0(\Inst_Mem/inst_mem_reg[48][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1748 ) );
  MUX \Inst_Mem/U1778  ( .IN0(\Inst_Mem/inst_mem_reg[50][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1747 ) );
  MUX \Inst_Mem/U1777  ( .IN0(\Inst_Mem/n1745 ), .IN1(\Inst_Mem/n1744 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1746 ) );
  MUX \Inst_Mem/U1776  ( .IN0(\Inst_Mem/inst_mem_reg[52][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1745 ) );
  MUX \Inst_Mem/U1775  ( .IN0(\Inst_Mem/inst_mem_reg[54][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1744 ) );
  MUX \Inst_Mem/U1774  ( .IN0(\Inst_Mem/n1742 ), .IN1(\Inst_Mem/n1739 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1743 ) );
  MUX \Inst_Mem/U1773  ( .IN0(\Inst_Mem/n1741 ), .IN1(\Inst_Mem/n1740 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1742 ) );
  MUX \Inst_Mem/U1772  ( .IN0(\Inst_Mem/inst_mem_reg[56][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1741 ) );
  MUX \Inst_Mem/U1771  ( .IN0(\Inst_Mem/inst_mem_reg[58][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1740 ) );
  MUX \Inst_Mem/U1770  ( .IN0(\Inst_Mem/n1738 ), .IN1(\Inst_Mem/n1737 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1739 ) );
  MUX \Inst_Mem/U1769  ( .IN0(\Inst_Mem/inst_mem_reg[60][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1738 ) );
  MUX \Inst_Mem/U1768  ( .IN0(\Inst_Mem/inst_mem_reg[62][28] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][28] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1737 ) );
  MUX \Inst_Mem/U1767  ( .IN0(\Inst_Mem/n1736 ), .IN1(\Inst_Mem/n1705 ), .SEL(
        pc_current[7]), .F(opcode[27]) );
  MUX \Inst_Mem/U1766  ( .IN0(\Inst_Mem/n1735 ), .IN1(\Inst_Mem/n1720 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1736 ) );
  MUX \Inst_Mem/U1765  ( .IN0(\Inst_Mem/n1734 ), .IN1(\Inst_Mem/n1727 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1735 ) );
  MUX \Inst_Mem/U1764  ( .IN0(\Inst_Mem/n1733 ), .IN1(\Inst_Mem/n1730 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1734 ) );
  MUX \Inst_Mem/U1763  ( .IN0(\Inst_Mem/n1732 ), .IN1(\Inst_Mem/n1731 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1733 ) );
  MUX \Inst_Mem/U1762  ( .IN0(\Inst_Mem/inst_mem_reg[0][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1732 ) );
  MUX \Inst_Mem/U1761  ( .IN0(\Inst_Mem/inst_mem_reg[2][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1731 ) );
  MUX \Inst_Mem/U1760  ( .IN0(\Inst_Mem/n1729 ), .IN1(\Inst_Mem/n1728 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1730 ) );
  MUX \Inst_Mem/U1759  ( .IN0(\Inst_Mem/inst_mem_reg[4][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1729 ) );
  MUX \Inst_Mem/U1758  ( .IN0(\Inst_Mem/inst_mem_reg[6][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1728 ) );
  MUX \Inst_Mem/U1757  ( .IN0(\Inst_Mem/n1726 ), .IN1(\Inst_Mem/n1723 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1727 ) );
  MUX \Inst_Mem/U1756  ( .IN0(\Inst_Mem/n1725 ), .IN1(\Inst_Mem/n1724 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1726 ) );
  MUX \Inst_Mem/U1755  ( .IN0(\Inst_Mem/inst_mem_reg[8][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1725 ) );
  MUX \Inst_Mem/U1754  ( .IN0(\Inst_Mem/inst_mem_reg[10][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1724 ) );
  MUX \Inst_Mem/U1753  ( .IN0(\Inst_Mem/n1722 ), .IN1(\Inst_Mem/n1721 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1723 ) );
  MUX \Inst_Mem/U1752  ( .IN0(\Inst_Mem/inst_mem_reg[12][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1722 ) );
  MUX \Inst_Mem/U1751  ( .IN0(\Inst_Mem/inst_mem_reg[14][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1721 ) );
  MUX \Inst_Mem/U1750  ( .IN0(\Inst_Mem/n1719 ), .IN1(\Inst_Mem/n1712 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1720 ) );
  MUX \Inst_Mem/U1749  ( .IN0(\Inst_Mem/n1718 ), .IN1(\Inst_Mem/n1715 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1719 ) );
  MUX \Inst_Mem/U1748  ( .IN0(\Inst_Mem/n1717 ), .IN1(\Inst_Mem/n1716 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1718 ) );
  MUX \Inst_Mem/U1747  ( .IN0(\Inst_Mem/inst_mem_reg[16][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1717 ) );
  MUX \Inst_Mem/U1746  ( .IN0(\Inst_Mem/inst_mem_reg[18][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1716 ) );
  MUX \Inst_Mem/U1745  ( .IN0(\Inst_Mem/n1714 ), .IN1(\Inst_Mem/n1713 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1715 ) );
  MUX \Inst_Mem/U1744  ( .IN0(\Inst_Mem/inst_mem_reg[20][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1714 ) );
  MUX \Inst_Mem/U1743  ( .IN0(\Inst_Mem/inst_mem_reg[22][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1713 ) );
  MUX \Inst_Mem/U1742  ( .IN0(\Inst_Mem/n1711 ), .IN1(\Inst_Mem/n1708 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1712 ) );
  MUX \Inst_Mem/U1741  ( .IN0(\Inst_Mem/n1710 ), .IN1(\Inst_Mem/n1709 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1711 ) );
  MUX \Inst_Mem/U1740  ( .IN0(\Inst_Mem/inst_mem_reg[24][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1710 ) );
  MUX \Inst_Mem/U1739  ( .IN0(\Inst_Mem/inst_mem_reg[26][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1709 ) );
  MUX \Inst_Mem/U1738  ( .IN0(\Inst_Mem/n1707 ), .IN1(\Inst_Mem/n1706 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1708 ) );
  MUX \Inst_Mem/U1737  ( .IN0(\Inst_Mem/inst_mem_reg[28][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1707 ) );
  MUX \Inst_Mem/U1736  ( .IN0(\Inst_Mem/inst_mem_reg[30][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1706 ) );
  MUX \Inst_Mem/U1735  ( .IN0(\Inst_Mem/n1704 ), .IN1(\Inst_Mem/n1689 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1705 ) );
  MUX \Inst_Mem/U1734  ( .IN0(\Inst_Mem/n1703 ), .IN1(\Inst_Mem/n1696 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1704 ) );
  MUX \Inst_Mem/U1733  ( .IN0(\Inst_Mem/n1702 ), .IN1(\Inst_Mem/n1699 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1703 ) );
  MUX \Inst_Mem/U1732  ( .IN0(\Inst_Mem/n1701 ), .IN1(\Inst_Mem/n1700 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1702 ) );
  MUX \Inst_Mem/U1731  ( .IN0(\Inst_Mem/inst_mem_reg[32][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1701 ) );
  MUX \Inst_Mem/U1730  ( .IN0(\Inst_Mem/inst_mem_reg[34][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1700 ) );
  MUX \Inst_Mem/U1729  ( .IN0(\Inst_Mem/n1698 ), .IN1(\Inst_Mem/n1697 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1699 ) );
  MUX \Inst_Mem/U1728  ( .IN0(\Inst_Mem/inst_mem_reg[36][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1698 ) );
  MUX \Inst_Mem/U1727  ( .IN0(\Inst_Mem/inst_mem_reg[38][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1697 ) );
  MUX \Inst_Mem/U1726  ( .IN0(\Inst_Mem/n1695 ), .IN1(\Inst_Mem/n1692 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1696 ) );
  MUX \Inst_Mem/U1725  ( .IN0(\Inst_Mem/n1694 ), .IN1(\Inst_Mem/n1693 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1695 ) );
  MUX \Inst_Mem/U1724  ( .IN0(\Inst_Mem/inst_mem_reg[40][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1694 ) );
  MUX \Inst_Mem/U1723  ( .IN0(\Inst_Mem/inst_mem_reg[42][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1693 ) );
  MUX \Inst_Mem/U1722  ( .IN0(\Inst_Mem/n1691 ), .IN1(\Inst_Mem/n1690 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1692 ) );
  MUX \Inst_Mem/U1721  ( .IN0(\Inst_Mem/inst_mem_reg[44][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1691 ) );
  MUX \Inst_Mem/U1720  ( .IN0(\Inst_Mem/inst_mem_reg[46][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1690 ) );
  MUX \Inst_Mem/U1719  ( .IN0(\Inst_Mem/n1688 ), .IN1(\Inst_Mem/n1681 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1689 ) );
  MUX \Inst_Mem/U1718  ( .IN0(\Inst_Mem/n1687 ), .IN1(\Inst_Mem/n1684 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1688 ) );
  MUX \Inst_Mem/U1717  ( .IN0(\Inst_Mem/n1686 ), .IN1(\Inst_Mem/n1685 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1687 ) );
  MUX \Inst_Mem/U1716  ( .IN0(\Inst_Mem/inst_mem_reg[48][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1686 ) );
  MUX \Inst_Mem/U1715  ( .IN0(\Inst_Mem/inst_mem_reg[50][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1685 ) );
  MUX \Inst_Mem/U1714  ( .IN0(\Inst_Mem/n1683 ), .IN1(\Inst_Mem/n1682 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1684 ) );
  MUX \Inst_Mem/U1713  ( .IN0(\Inst_Mem/inst_mem_reg[52][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1683 ) );
  MUX \Inst_Mem/U1712  ( .IN0(\Inst_Mem/inst_mem_reg[54][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1682 ) );
  MUX \Inst_Mem/U1711  ( .IN0(\Inst_Mem/n1680 ), .IN1(\Inst_Mem/n1677 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1681 ) );
  MUX \Inst_Mem/U1710  ( .IN0(\Inst_Mem/n1679 ), .IN1(\Inst_Mem/n1678 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1680 ) );
  MUX \Inst_Mem/U1709  ( .IN0(\Inst_Mem/inst_mem_reg[56][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1679 ) );
  MUX \Inst_Mem/U1708  ( .IN0(\Inst_Mem/inst_mem_reg[58][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1678 ) );
  MUX \Inst_Mem/U1707  ( .IN0(\Inst_Mem/n1676 ), .IN1(\Inst_Mem/n1675 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1677 ) );
  MUX \Inst_Mem/U1706  ( .IN0(\Inst_Mem/inst_mem_reg[60][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1676 ) );
  MUX \Inst_Mem/U1705  ( .IN0(\Inst_Mem/inst_mem_reg[62][27] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][27] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1675 ) );
  MUX \Inst_Mem/U1704  ( .IN0(\Inst_Mem/n1674 ), .IN1(\Inst_Mem/n1643 ), .SEL(
        pc_current[7]), .F(opcode[26]) );
  MUX \Inst_Mem/U1703  ( .IN0(\Inst_Mem/n1673 ), .IN1(\Inst_Mem/n1658 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1674 ) );
  MUX \Inst_Mem/U1702  ( .IN0(\Inst_Mem/n1672 ), .IN1(\Inst_Mem/n1665 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1673 ) );
  MUX \Inst_Mem/U1701  ( .IN0(\Inst_Mem/n1671 ), .IN1(\Inst_Mem/n1668 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1672 ) );
  MUX \Inst_Mem/U1700  ( .IN0(\Inst_Mem/n1670 ), .IN1(\Inst_Mem/n1669 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1671 ) );
  MUX \Inst_Mem/U1699  ( .IN0(\Inst_Mem/inst_mem_reg[0][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1670 ) );
  MUX \Inst_Mem/U1698  ( .IN0(\Inst_Mem/inst_mem_reg[2][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1669 ) );
  MUX \Inst_Mem/U1697  ( .IN0(\Inst_Mem/n1667 ), .IN1(\Inst_Mem/n1666 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1668 ) );
  MUX \Inst_Mem/U1696  ( .IN0(\Inst_Mem/inst_mem_reg[4][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1667 ) );
  MUX \Inst_Mem/U1695  ( .IN0(\Inst_Mem/inst_mem_reg[6][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1666 ) );
  MUX \Inst_Mem/U1694  ( .IN0(\Inst_Mem/n1664 ), .IN1(\Inst_Mem/n1661 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1665 ) );
  MUX \Inst_Mem/U1693  ( .IN0(\Inst_Mem/n1663 ), .IN1(\Inst_Mem/n1662 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1664 ) );
  MUX \Inst_Mem/U1692  ( .IN0(\Inst_Mem/inst_mem_reg[8][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1663 ) );
  MUX \Inst_Mem/U1691  ( .IN0(\Inst_Mem/inst_mem_reg[10][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1662 ) );
  MUX \Inst_Mem/U1690  ( .IN0(\Inst_Mem/n1660 ), .IN1(\Inst_Mem/n1659 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1661 ) );
  MUX \Inst_Mem/U1689  ( .IN0(\Inst_Mem/inst_mem_reg[12][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1660 ) );
  MUX \Inst_Mem/U1688  ( .IN0(\Inst_Mem/inst_mem_reg[14][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1659 ) );
  MUX \Inst_Mem/U1687  ( .IN0(\Inst_Mem/n1657 ), .IN1(\Inst_Mem/n1650 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1658 ) );
  MUX \Inst_Mem/U1686  ( .IN0(\Inst_Mem/n1656 ), .IN1(\Inst_Mem/n1653 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1657 ) );
  MUX \Inst_Mem/U1685  ( .IN0(\Inst_Mem/n1655 ), .IN1(\Inst_Mem/n1654 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1656 ) );
  MUX \Inst_Mem/U1684  ( .IN0(\Inst_Mem/inst_mem_reg[16][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1655 ) );
  MUX \Inst_Mem/U1683  ( .IN0(\Inst_Mem/inst_mem_reg[18][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1654 ) );
  MUX \Inst_Mem/U1682  ( .IN0(\Inst_Mem/n1652 ), .IN1(\Inst_Mem/n1651 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1653 ) );
  MUX \Inst_Mem/U1681  ( .IN0(\Inst_Mem/inst_mem_reg[20][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1652 ) );
  MUX \Inst_Mem/U1680  ( .IN0(\Inst_Mem/inst_mem_reg[22][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1651 ) );
  MUX \Inst_Mem/U1679  ( .IN0(\Inst_Mem/n1649 ), .IN1(\Inst_Mem/n1646 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1650 ) );
  MUX \Inst_Mem/U1678  ( .IN0(\Inst_Mem/n1648 ), .IN1(\Inst_Mem/n1647 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1649 ) );
  MUX \Inst_Mem/U1677  ( .IN0(\Inst_Mem/inst_mem_reg[24][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1648 ) );
  MUX \Inst_Mem/U1676  ( .IN0(\Inst_Mem/inst_mem_reg[26][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1647 ) );
  MUX \Inst_Mem/U1675  ( .IN0(\Inst_Mem/n1645 ), .IN1(\Inst_Mem/n1644 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1646 ) );
  MUX \Inst_Mem/U1674  ( .IN0(\Inst_Mem/inst_mem_reg[28][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1645 ) );
  MUX \Inst_Mem/U1673  ( .IN0(\Inst_Mem/inst_mem_reg[30][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1644 ) );
  MUX \Inst_Mem/U1672  ( .IN0(\Inst_Mem/n1642 ), .IN1(\Inst_Mem/n1627 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1643 ) );
  MUX \Inst_Mem/U1671  ( .IN0(\Inst_Mem/n1641 ), .IN1(\Inst_Mem/n1634 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1642 ) );
  MUX \Inst_Mem/U1670  ( .IN0(\Inst_Mem/n1640 ), .IN1(\Inst_Mem/n1637 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1641 ) );
  MUX \Inst_Mem/U1669  ( .IN0(\Inst_Mem/n1639 ), .IN1(\Inst_Mem/n1638 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1640 ) );
  MUX \Inst_Mem/U1668  ( .IN0(\Inst_Mem/inst_mem_reg[32][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1639 ) );
  MUX \Inst_Mem/U1667  ( .IN0(\Inst_Mem/inst_mem_reg[34][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1638 ) );
  MUX \Inst_Mem/U1666  ( .IN0(\Inst_Mem/n1636 ), .IN1(\Inst_Mem/n1635 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1637 ) );
  MUX \Inst_Mem/U1665  ( .IN0(\Inst_Mem/inst_mem_reg[36][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1636 ) );
  MUX \Inst_Mem/U1664  ( .IN0(\Inst_Mem/inst_mem_reg[38][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1635 ) );
  MUX \Inst_Mem/U1663  ( .IN0(\Inst_Mem/n1633 ), .IN1(\Inst_Mem/n1630 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1634 ) );
  MUX \Inst_Mem/U1662  ( .IN0(\Inst_Mem/n1632 ), .IN1(\Inst_Mem/n1631 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1633 ) );
  MUX \Inst_Mem/U1661  ( .IN0(\Inst_Mem/inst_mem_reg[40][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1632 ) );
  MUX \Inst_Mem/U1660  ( .IN0(\Inst_Mem/inst_mem_reg[42][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1631 ) );
  MUX \Inst_Mem/U1659  ( .IN0(\Inst_Mem/n1629 ), .IN1(\Inst_Mem/n1628 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1630 ) );
  MUX \Inst_Mem/U1658  ( .IN0(\Inst_Mem/inst_mem_reg[44][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1629 ) );
  MUX \Inst_Mem/U1657  ( .IN0(\Inst_Mem/inst_mem_reg[46][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1628 ) );
  MUX \Inst_Mem/U1656  ( .IN0(\Inst_Mem/n1626 ), .IN1(\Inst_Mem/n1619 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1627 ) );
  MUX \Inst_Mem/U1655  ( .IN0(\Inst_Mem/n1625 ), .IN1(\Inst_Mem/n1622 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1626 ) );
  MUX \Inst_Mem/U1654  ( .IN0(\Inst_Mem/n1624 ), .IN1(\Inst_Mem/n1623 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1625 ) );
  MUX \Inst_Mem/U1653  ( .IN0(\Inst_Mem/inst_mem_reg[48][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1624 ) );
  MUX \Inst_Mem/U1652  ( .IN0(\Inst_Mem/inst_mem_reg[50][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1623 ) );
  MUX \Inst_Mem/U1651  ( .IN0(\Inst_Mem/n1621 ), .IN1(\Inst_Mem/n1620 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1622 ) );
  MUX \Inst_Mem/U1650  ( .IN0(\Inst_Mem/inst_mem_reg[52][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1621 ) );
  MUX \Inst_Mem/U1649  ( .IN0(\Inst_Mem/inst_mem_reg[54][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1620 ) );
  MUX \Inst_Mem/U1648  ( .IN0(\Inst_Mem/n1618 ), .IN1(\Inst_Mem/n1615 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1619 ) );
  MUX \Inst_Mem/U1647  ( .IN0(\Inst_Mem/n1617 ), .IN1(\Inst_Mem/n1616 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1618 ) );
  MUX \Inst_Mem/U1646  ( .IN0(\Inst_Mem/inst_mem_reg[56][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1617 ) );
  MUX \Inst_Mem/U1645  ( .IN0(\Inst_Mem/inst_mem_reg[58][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1616 ) );
  MUX \Inst_Mem/U1644  ( .IN0(\Inst_Mem/n1614 ), .IN1(\Inst_Mem/n1613 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1615 ) );
  MUX \Inst_Mem/U1643  ( .IN0(\Inst_Mem/inst_mem_reg[60][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1614 ) );
  MUX \Inst_Mem/U1642  ( .IN0(\Inst_Mem/inst_mem_reg[62][26] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][26] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1613 ) );
  MUX \Inst_Mem/U1641  ( .IN0(\Inst_Mem/n1612 ), .IN1(\Inst_Mem/n1581 ), .SEL(
        pc_current[7]), .F(opcode[25]) );
  MUX \Inst_Mem/U1640  ( .IN0(\Inst_Mem/n1611 ), .IN1(\Inst_Mem/n1596 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1612 ) );
  MUX \Inst_Mem/U1639  ( .IN0(\Inst_Mem/n1610 ), .IN1(\Inst_Mem/n1603 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1611 ) );
  MUX \Inst_Mem/U1638  ( .IN0(\Inst_Mem/n1609 ), .IN1(\Inst_Mem/n1606 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1610 ) );
  MUX \Inst_Mem/U1637  ( .IN0(\Inst_Mem/n1608 ), .IN1(\Inst_Mem/n1607 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1609 ) );
  MUX \Inst_Mem/U1636  ( .IN0(\Inst_Mem/inst_mem_reg[0][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1608 ) );
  MUX \Inst_Mem/U1635  ( .IN0(\Inst_Mem/inst_mem_reg[2][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1607 ) );
  MUX \Inst_Mem/U1634  ( .IN0(\Inst_Mem/n1605 ), .IN1(\Inst_Mem/n1604 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1606 ) );
  MUX \Inst_Mem/U1633  ( .IN0(\Inst_Mem/inst_mem_reg[4][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1605 ) );
  MUX \Inst_Mem/U1632  ( .IN0(\Inst_Mem/inst_mem_reg[6][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1604 ) );
  MUX \Inst_Mem/U1631  ( .IN0(\Inst_Mem/n1602 ), .IN1(\Inst_Mem/n1599 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1603 ) );
  MUX \Inst_Mem/U1630  ( .IN0(\Inst_Mem/n1601 ), .IN1(\Inst_Mem/n1600 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1602 ) );
  MUX \Inst_Mem/U1629  ( .IN0(\Inst_Mem/inst_mem_reg[8][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1601 ) );
  MUX \Inst_Mem/U1628  ( .IN0(\Inst_Mem/inst_mem_reg[10][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1600 ) );
  MUX \Inst_Mem/U1627  ( .IN0(\Inst_Mem/n1598 ), .IN1(\Inst_Mem/n1597 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1599 ) );
  MUX \Inst_Mem/U1626  ( .IN0(\Inst_Mem/inst_mem_reg[12][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1598 ) );
  MUX \Inst_Mem/U1625  ( .IN0(\Inst_Mem/inst_mem_reg[14][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1597 ) );
  MUX \Inst_Mem/U1624  ( .IN0(\Inst_Mem/n1595 ), .IN1(\Inst_Mem/n1588 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1596 ) );
  MUX \Inst_Mem/U1623  ( .IN0(\Inst_Mem/n1594 ), .IN1(\Inst_Mem/n1591 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1595 ) );
  MUX \Inst_Mem/U1622  ( .IN0(\Inst_Mem/n1593 ), .IN1(\Inst_Mem/n1592 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1594 ) );
  MUX \Inst_Mem/U1621  ( .IN0(\Inst_Mem/inst_mem_reg[16][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1593 ) );
  MUX \Inst_Mem/U1620  ( .IN0(\Inst_Mem/inst_mem_reg[18][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1592 ) );
  MUX \Inst_Mem/U1619  ( .IN0(\Inst_Mem/n1590 ), .IN1(\Inst_Mem/n1589 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1591 ) );
  MUX \Inst_Mem/U1618  ( .IN0(\Inst_Mem/inst_mem_reg[20][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1590 ) );
  MUX \Inst_Mem/U1617  ( .IN0(\Inst_Mem/inst_mem_reg[22][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1589 ) );
  MUX \Inst_Mem/U1616  ( .IN0(\Inst_Mem/n1587 ), .IN1(\Inst_Mem/n1584 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1588 ) );
  MUX \Inst_Mem/U1615  ( .IN0(\Inst_Mem/n1586 ), .IN1(\Inst_Mem/n1585 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1587 ) );
  MUX \Inst_Mem/U1614  ( .IN0(\Inst_Mem/inst_mem_reg[24][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1586 ) );
  MUX \Inst_Mem/U1613  ( .IN0(\Inst_Mem/inst_mem_reg[26][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1585 ) );
  MUX \Inst_Mem/U1612  ( .IN0(\Inst_Mem/n1583 ), .IN1(\Inst_Mem/n1582 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1584 ) );
  MUX \Inst_Mem/U1611  ( .IN0(\Inst_Mem/inst_mem_reg[28][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1583 ) );
  MUX \Inst_Mem/U1610  ( .IN0(\Inst_Mem/inst_mem_reg[30][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1582 ) );
  MUX \Inst_Mem/U1609  ( .IN0(\Inst_Mem/n1580 ), .IN1(\Inst_Mem/n1565 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1581 ) );
  MUX \Inst_Mem/U1608  ( .IN0(\Inst_Mem/n1579 ), .IN1(\Inst_Mem/n1572 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1580 ) );
  MUX \Inst_Mem/U1607  ( .IN0(\Inst_Mem/n1578 ), .IN1(\Inst_Mem/n1575 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1579 ) );
  MUX \Inst_Mem/U1606  ( .IN0(\Inst_Mem/n1577 ), .IN1(\Inst_Mem/n1576 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1578 ) );
  MUX \Inst_Mem/U1605  ( .IN0(\Inst_Mem/inst_mem_reg[32][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1577 ) );
  MUX \Inst_Mem/U1604  ( .IN0(\Inst_Mem/inst_mem_reg[34][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1576 ) );
  MUX \Inst_Mem/U1603  ( .IN0(\Inst_Mem/n1574 ), .IN1(\Inst_Mem/n1573 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1575 ) );
  MUX \Inst_Mem/U1602  ( .IN0(\Inst_Mem/inst_mem_reg[36][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1574 ) );
  MUX \Inst_Mem/U1601  ( .IN0(\Inst_Mem/inst_mem_reg[38][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1573 ) );
  MUX \Inst_Mem/U1600  ( .IN0(\Inst_Mem/n1571 ), .IN1(\Inst_Mem/n1568 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1572 ) );
  MUX \Inst_Mem/U1599  ( .IN0(\Inst_Mem/n1570 ), .IN1(\Inst_Mem/n1569 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1571 ) );
  MUX \Inst_Mem/U1598  ( .IN0(\Inst_Mem/inst_mem_reg[40][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1570 ) );
  MUX \Inst_Mem/U1597  ( .IN0(\Inst_Mem/inst_mem_reg[42][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1569 ) );
  MUX \Inst_Mem/U1596  ( .IN0(\Inst_Mem/n1567 ), .IN1(\Inst_Mem/n1566 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1568 ) );
  MUX \Inst_Mem/U1595  ( .IN0(\Inst_Mem/inst_mem_reg[44][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1567 ) );
  MUX \Inst_Mem/U1594  ( .IN0(\Inst_Mem/inst_mem_reg[46][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1566 ) );
  MUX \Inst_Mem/U1593  ( .IN0(\Inst_Mem/n1564 ), .IN1(\Inst_Mem/n1557 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1565 ) );
  MUX \Inst_Mem/U1592  ( .IN0(\Inst_Mem/n1563 ), .IN1(\Inst_Mem/n1560 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1564 ) );
  MUX \Inst_Mem/U1591  ( .IN0(\Inst_Mem/n1562 ), .IN1(\Inst_Mem/n1561 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1563 ) );
  MUX \Inst_Mem/U1590  ( .IN0(\Inst_Mem/inst_mem_reg[48][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1562 ) );
  MUX \Inst_Mem/U1589  ( .IN0(\Inst_Mem/inst_mem_reg[50][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1561 ) );
  MUX \Inst_Mem/U1588  ( .IN0(\Inst_Mem/n1559 ), .IN1(\Inst_Mem/n1558 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1560 ) );
  MUX \Inst_Mem/U1587  ( .IN0(\Inst_Mem/inst_mem_reg[52][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1559 ) );
  MUX \Inst_Mem/U1586  ( .IN0(\Inst_Mem/inst_mem_reg[54][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1558 ) );
  MUX \Inst_Mem/U1585  ( .IN0(\Inst_Mem/n1556 ), .IN1(\Inst_Mem/n1553 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1557 ) );
  MUX \Inst_Mem/U1584  ( .IN0(\Inst_Mem/n1555 ), .IN1(\Inst_Mem/n1554 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1556 ) );
  MUX \Inst_Mem/U1583  ( .IN0(\Inst_Mem/inst_mem_reg[56][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1555 ) );
  MUX \Inst_Mem/U1582  ( .IN0(\Inst_Mem/inst_mem_reg[58][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1554 ) );
  MUX \Inst_Mem/U1581  ( .IN0(\Inst_Mem/n1552 ), .IN1(\Inst_Mem/n1551 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1553 ) );
  MUX \Inst_Mem/U1580  ( .IN0(\Inst_Mem/inst_mem_reg[60][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1552 ) );
  MUX \Inst_Mem/U1579  ( .IN0(\Inst_Mem/inst_mem_reg[62][25] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][25] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1551 ) );
  MUX \Inst_Mem/U1578  ( .IN0(\Inst_Mem/n1550 ), .IN1(\Inst_Mem/n1519 ), .SEL(
        pc_current[7]), .F(opcode[24]) );
  MUX \Inst_Mem/U1577  ( .IN0(\Inst_Mem/n1549 ), .IN1(\Inst_Mem/n1534 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1550 ) );
  MUX \Inst_Mem/U1576  ( .IN0(\Inst_Mem/n1548 ), .IN1(\Inst_Mem/n1541 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1549 ) );
  MUX \Inst_Mem/U1575  ( .IN0(\Inst_Mem/n1547 ), .IN1(\Inst_Mem/n1544 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1548 ) );
  MUX \Inst_Mem/U1574  ( .IN0(\Inst_Mem/n1546 ), .IN1(\Inst_Mem/n1545 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1547 ) );
  MUX \Inst_Mem/U1573  ( .IN0(\Inst_Mem/inst_mem_reg[0][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1546 ) );
  MUX \Inst_Mem/U1572  ( .IN0(\Inst_Mem/inst_mem_reg[2][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1545 ) );
  MUX \Inst_Mem/U1571  ( .IN0(\Inst_Mem/n1543 ), .IN1(\Inst_Mem/n1542 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1544 ) );
  MUX \Inst_Mem/U1570  ( .IN0(\Inst_Mem/inst_mem_reg[4][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1543 ) );
  MUX \Inst_Mem/U1569  ( .IN0(\Inst_Mem/inst_mem_reg[6][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1542 ) );
  MUX \Inst_Mem/U1568  ( .IN0(\Inst_Mem/n1540 ), .IN1(\Inst_Mem/n1537 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1541 ) );
  MUX \Inst_Mem/U1567  ( .IN0(\Inst_Mem/n1539 ), .IN1(\Inst_Mem/n1538 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1540 ) );
  MUX \Inst_Mem/U1566  ( .IN0(\Inst_Mem/inst_mem_reg[8][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1539 ) );
  MUX \Inst_Mem/U1565  ( .IN0(\Inst_Mem/inst_mem_reg[10][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1538 ) );
  MUX \Inst_Mem/U1564  ( .IN0(\Inst_Mem/n1536 ), .IN1(\Inst_Mem/n1535 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1537 ) );
  MUX \Inst_Mem/U1563  ( .IN0(\Inst_Mem/inst_mem_reg[12][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1536 ) );
  MUX \Inst_Mem/U1562  ( .IN0(\Inst_Mem/inst_mem_reg[14][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1535 ) );
  MUX \Inst_Mem/U1561  ( .IN0(\Inst_Mem/n1533 ), .IN1(\Inst_Mem/n1526 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1534 ) );
  MUX \Inst_Mem/U1560  ( .IN0(\Inst_Mem/n1532 ), .IN1(\Inst_Mem/n1529 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1533 ) );
  MUX \Inst_Mem/U1559  ( .IN0(\Inst_Mem/n1531 ), .IN1(\Inst_Mem/n1530 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1532 ) );
  MUX \Inst_Mem/U1558  ( .IN0(\Inst_Mem/inst_mem_reg[16][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1531 ) );
  MUX \Inst_Mem/U1557  ( .IN0(\Inst_Mem/inst_mem_reg[18][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1530 ) );
  MUX \Inst_Mem/U1556  ( .IN0(\Inst_Mem/n1528 ), .IN1(\Inst_Mem/n1527 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1529 ) );
  MUX \Inst_Mem/U1555  ( .IN0(\Inst_Mem/inst_mem_reg[20][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1528 ) );
  MUX \Inst_Mem/U1554  ( .IN0(\Inst_Mem/inst_mem_reg[22][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1527 ) );
  MUX \Inst_Mem/U1553  ( .IN0(\Inst_Mem/n1525 ), .IN1(\Inst_Mem/n1522 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1526 ) );
  MUX \Inst_Mem/U1552  ( .IN0(\Inst_Mem/n1524 ), .IN1(\Inst_Mem/n1523 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1525 ) );
  MUX \Inst_Mem/U1551  ( .IN0(\Inst_Mem/inst_mem_reg[24][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1524 ) );
  MUX \Inst_Mem/U1550  ( .IN0(\Inst_Mem/inst_mem_reg[26][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1523 ) );
  MUX \Inst_Mem/U1549  ( .IN0(\Inst_Mem/n1521 ), .IN1(\Inst_Mem/n1520 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1522 ) );
  MUX \Inst_Mem/U1548  ( .IN0(\Inst_Mem/inst_mem_reg[28][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1521 ) );
  MUX \Inst_Mem/U1547  ( .IN0(\Inst_Mem/inst_mem_reg[30][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1520 ) );
  MUX \Inst_Mem/U1546  ( .IN0(\Inst_Mem/n1518 ), .IN1(\Inst_Mem/n1503 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1519 ) );
  MUX \Inst_Mem/U1545  ( .IN0(\Inst_Mem/n1517 ), .IN1(\Inst_Mem/n1510 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1518 ) );
  MUX \Inst_Mem/U1544  ( .IN0(\Inst_Mem/n1516 ), .IN1(\Inst_Mem/n1513 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1517 ) );
  MUX \Inst_Mem/U1543  ( .IN0(\Inst_Mem/n1515 ), .IN1(\Inst_Mem/n1514 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1516 ) );
  MUX \Inst_Mem/U1542  ( .IN0(\Inst_Mem/inst_mem_reg[32][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1515 ) );
  MUX \Inst_Mem/U1541  ( .IN0(\Inst_Mem/inst_mem_reg[34][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1514 ) );
  MUX \Inst_Mem/U1540  ( .IN0(\Inst_Mem/n1512 ), .IN1(\Inst_Mem/n1511 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1513 ) );
  MUX \Inst_Mem/U1539  ( .IN0(\Inst_Mem/inst_mem_reg[36][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1512 ) );
  MUX \Inst_Mem/U1538  ( .IN0(\Inst_Mem/inst_mem_reg[38][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1511 ) );
  MUX \Inst_Mem/U1537  ( .IN0(\Inst_Mem/n1509 ), .IN1(\Inst_Mem/n1506 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1510 ) );
  MUX \Inst_Mem/U1536  ( .IN0(\Inst_Mem/n1508 ), .IN1(\Inst_Mem/n1507 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1509 ) );
  MUX \Inst_Mem/U1535  ( .IN0(\Inst_Mem/inst_mem_reg[40][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1508 ) );
  MUX \Inst_Mem/U1534  ( .IN0(\Inst_Mem/inst_mem_reg[42][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1507 ) );
  MUX \Inst_Mem/U1533  ( .IN0(\Inst_Mem/n1505 ), .IN1(\Inst_Mem/n1504 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1506 ) );
  MUX \Inst_Mem/U1532  ( .IN0(\Inst_Mem/inst_mem_reg[44][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1505 ) );
  MUX \Inst_Mem/U1531  ( .IN0(\Inst_Mem/inst_mem_reg[46][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1504 ) );
  MUX \Inst_Mem/U1530  ( .IN0(\Inst_Mem/n1502 ), .IN1(\Inst_Mem/n1495 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1503 ) );
  MUX \Inst_Mem/U1529  ( .IN0(\Inst_Mem/n1501 ), .IN1(\Inst_Mem/n1498 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1502 ) );
  MUX \Inst_Mem/U1528  ( .IN0(\Inst_Mem/n1500 ), .IN1(\Inst_Mem/n1499 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1501 ) );
  MUX \Inst_Mem/U1527  ( .IN0(\Inst_Mem/inst_mem_reg[48][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1500 ) );
  MUX \Inst_Mem/U1526  ( .IN0(\Inst_Mem/inst_mem_reg[50][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1499 ) );
  MUX \Inst_Mem/U1525  ( .IN0(\Inst_Mem/n1497 ), .IN1(\Inst_Mem/n1496 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1498 ) );
  MUX \Inst_Mem/U1524  ( .IN0(\Inst_Mem/inst_mem_reg[52][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1497 ) );
  MUX \Inst_Mem/U1523  ( .IN0(\Inst_Mem/inst_mem_reg[54][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1496 ) );
  MUX \Inst_Mem/U1522  ( .IN0(\Inst_Mem/n1494 ), .IN1(\Inst_Mem/n1491 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1495 ) );
  MUX \Inst_Mem/U1521  ( .IN0(\Inst_Mem/n1493 ), .IN1(\Inst_Mem/n1492 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1494 ) );
  MUX \Inst_Mem/U1520  ( .IN0(\Inst_Mem/inst_mem_reg[56][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1493 ) );
  MUX \Inst_Mem/U1519  ( .IN0(\Inst_Mem/inst_mem_reg[58][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1492 ) );
  MUX \Inst_Mem/U1518  ( .IN0(\Inst_Mem/n1490 ), .IN1(\Inst_Mem/n1489 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1491 ) );
  MUX \Inst_Mem/U1517  ( .IN0(\Inst_Mem/inst_mem_reg[60][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1490 ) );
  MUX \Inst_Mem/U1516  ( .IN0(\Inst_Mem/inst_mem_reg[62][24] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][24] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1489 ) );
  MUX \Inst_Mem/U1515  ( .IN0(\Inst_Mem/n1488 ), .IN1(\Inst_Mem/n1457 ), .SEL(
        pc_current[7]), .F(opcode[23]) );
  MUX \Inst_Mem/U1514  ( .IN0(\Inst_Mem/n1487 ), .IN1(\Inst_Mem/n1472 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1488 ) );
  MUX \Inst_Mem/U1513  ( .IN0(\Inst_Mem/n1486 ), .IN1(\Inst_Mem/n1479 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1487 ) );
  MUX \Inst_Mem/U1512  ( .IN0(\Inst_Mem/n1485 ), .IN1(\Inst_Mem/n1482 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1486 ) );
  MUX \Inst_Mem/U1511  ( .IN0(\Inst_Mem/n1484 ), .IN1(\Inst_Mem/n1483 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1485 ) );
  MUX \Inst_Mem/U1510  ( .IN0(\Inst_Mem/inst_mem_reg[0][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1484 ) );
  MUX \Inst_Mem/U1509  ( .IN0(\Inst_Mem/inst_mem_reg[2][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1483 ) );
  MUX \Inst_Mem/U1508  ( .IN0(\Inst_Mem/n1481 ), .IN1(\Inst_Mem/n1480 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1482 ) );
  MUX \Inst_Mem/U1507  ( .IN0(\Inst_Mem/inst_mem_reg[4][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1481 ) );
  MUX \Inst_Mem/U1506  ( .IN0(\Inst_Mem/inst_mem_reg[6][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1480 ) );
  MUX \Inst_Mem/U1505  ( .IN0(\Inst_Mem/n1478 ), .IN1(\Inst_Mem/n1475 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1479 ) );
  MUX \Inst_Mem/U1504  ( .IN0(\Inst_Mem/n1477 ), .IN1(\Inst_Mem/n1476 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1478 ) );
  MUX \Inst_Mem/U1503  ( .IN0(\Inst_Mem/inst_mem_reg[8][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1477 ) );
  MUX \Inst_Mem/U1502  ( .IN0(\Inst_Mem/inst_mem_reg[10][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1476 ) );
  MUX \Inst_Mem/U1501  ( .IN0(\Inst_Mem/n1474 ), .IN1(\Inst_Mem/n1473 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1475 ) );
  MUX \Inst_Mem/U1500  ( .IN0(\Inst_Mem/inst_mem_reg[12][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1474 ) );
  MUX \Inst_Mem/U1499  ( .IN0(\Inst_Mem/inst_mem_reg[14][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1473 ) );
  MUX \Inst_Mem/U1498  ( .IN0(\Inst_Mem/n1471 ), .IN1(\Inst_Mem/n1464 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1472 ) );
  MUX \Inst_Mem/U1497  ( .IN0(\Inst_Mem/n1470 ), .IN1(\Inst_Mem/n1467 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1471 ) );
  MUX \Inst_Mem/U1496  ( .IN0(\Inst_Mem/n1469 ), .IN1(\Inst_Mem/n1468 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1470 ) );
  MUX \Inst_Mem/U1495  ( .IN0(\Inst_Mem/inst_mem_reg[16][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1469 ) );
  MUX \Inst_Mem/U1494  ( .IN0(\Inst_Mem/inst_mem_reg[18][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1468 ) );
  MUX \Inst_Mem/U1493  ( .IN0(\Inst_Mem/n1466 ), .IN1(\Inst_Mem/n1465 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1467 ) );
  MUX \Inst_Mem/U1492  ( .IN0(\Inst_Mem/inst_mem_reg[20][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1466 ) );
  MUX \Inst_Mem/U1491  ( .IN0(\Inst_Mem/inst_mem_reg[22][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1465 ) );
  MUX \Inst_Mem/U1490  ( .IN0(\Inst_Mem/n1463 ), .IN1(\Inst_Mem/n1460 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1464 ) );
  MUX \Inst_Mem/U1489  ( .IN0(\Inst_Mem/n1462 ), .IN1(\Inst_Mem/n1461 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1463 ) );
  MUX \Inst_Mem/U1488  ( .IN0(\Inst_Mem/inst_mem_reg[24][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1462 ) );
  MUX \Inst_Mem/U1487  ( .IN0(\Inst_Mem/inst_mem_reg[26][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1461 ) );
  MUX \Inst_Mem/U1486  ( .IN0(\Inst_Mem/n1459 ), .IN1(\Inst_Mem/n1458 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1460 ) );
  MUX \Inst_Mem/U1485  ( .IN0(\Inst_Mem/inst_mem_reg[28][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1459 ) );
  MUX \Inst_Mem/U1484  ( .IN0(\Inst_Mem/inst_mem_reg[30][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1458 ) );
  MUX \Inst_Mem/U1483  ( .IN0(\Inst_Mem/n1456 ), .IN1(\Inst_Mem/n1441 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1457 ) );
  MUX \Inst_Mem/U1482  ( .IN0(\Inst_Mem/n1455 ), .IN1(\Inst_Mem/n1448 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1456 ) );
  MUX \Inst_Mem/U1481  ( .IN0(\Inst_Mem/n1454 ), .IN1(\Inst_Mem/n1451 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1455 ) );
  MUX \Inst_Mem/U1480  ( .IN0(\Inst_Mem/n1453 ), .IN1(\Inst_Mem/n1452 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1454 ) );
  MUX \Inst_Mem/U1479  ( .IN0(\Inst_Mem/inst_mem_reg[32][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1453 ) );
  MUX \Inst_Mem/U1478  ( .IN0(\Inst_Mem/inst_mem_reg[34][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1452 ) );
  MUX \Inst_Mem/U1477  ( .IN0(\Inst_Mem/n1450 ), .IN1(\Inst_Mem/n1449 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1451 ) );
  MUX \Inst_Mem/U1476  ( .IN0(\Inst_Mem/inst_mem_reg[36][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1450 ) );
  MUX \Inst_Mem/U1475  ( .IN0(\Inst_Mem/inst_mem_reg[38][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1449 ) );
  MUX \Inst_Mem/U1474  ( .IN0(\Inst_Mem/n1447 ), .IN1(\Inst_Mem/n1444 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1448 ) );
  MUX \Inst_Mem/U1473  ( .IN0(\Inst_Mem/n1446 ), .IN1(\Inst_Mem/n1445 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1447 ) );
  MUX \Inst_Mem/U1472  ( .IN0(\Inst_Mem/inst_mem_reg[40][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1446 ) );
  MUX \Inst_Mem/U1471  ( .IN0(\Inst_Mem/inst_mem_reg[42][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1445 ) );
  MUX \Inst_Mem/U1470  ( .IN0(\Inst_Mem/n1443 ), .IN1(\Inst_Mem/n1442 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1444 ) );
  MUX \Inst_Mem/U1469  ( .IN0(\Inst_Mem/inst_mem_reg[44][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1443 ) );
  MUX \Inst_Mem/U1468  ( .IN0(\Inst_Mem/inst_mem_reg[46][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1442 ) );
  MUX \Inst_Mem/U1467  ( .IN0(\Inst_Mem/n1440 ), .IN1(\Inst_Mem/n1433 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1441 ) );
  MUX \Inst_Mem/U1466  ( .IN0(\Inst_Mem/n1439 ), .IN1(\Inst_Mem/n1436 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1440 ) );
  MUX \Inst_Mem/U1465  ( .IN0(\Inst_Mem/n1438 ), .IN1(\Inst_Mem/n1437 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1439 ) );
  MUX \Inst_Mem/U1464  ( .IN0(\Inst_Mem/inst_mem_reg[48][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1438 ) );
  MUX \Inst_Mem/U1463  ( .IN0(\Inst_Mem/inst_mem_reg[50][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1437 ) );
  MUX \Inst_Mem/U1462  ( .IN0(\Inst_Mem/n1435 ), .IN1(\Inst_Mem/n1434 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1436 ) );
  MUX \Inst_Mem/U1461  ( .IN0(\Inst_Mem/inst_mem_reg[52][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1435 ) );
  MUX \Inst_Mem/U1460  ( .IN0(\Inst_Mem/inst_mem_reg[54][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1434 ) );
  MUX \Inst_Mem/U1459  ( .IN0(\Inst_Mem/n1432 ), .IN1(\Inst_Mem/n1429 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1433 ) );
  MUX \Inst_Mem/U1458  ( .IN0(\Inst_Mem/n1431 ), .IN1(\Inst_Mem/n1430 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1432 ) );
  MUX \Inst_Mem/U1457  ( .IN0(\Inst_Mem/inst_mem_reg[56][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1431 ) );
  MUX \Inst_Mem/U1456  ( .IN0(\Inst_Mem/inst_mem_reg[58][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1430 ) );
  MUX \Inst_Mem/U1455  ( .IN0(\Inst_Mem/n1428 ), .IN1(\Inst_Mem/n1427 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1429 ) );
  MUX \Inst_Mem/U1454  ( .IN0(\Inst_Mem/inst_mem_reg[60][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1428 ) );
  MUX \Inst_Mem/U1453  ( .IN0(\Inst_Mem/inst_mem_reg[62][23] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][23] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1427 ) );
  MUX \Inst_Mem/U1452  ( .IN0(\Inst_Mem/n1426 ), .IN1(\Inst_Mem/n1395 ), .SEL(
        pc_current[7]), .F(opcode[22]) );
  MUX \Inst_Mem/U1451  ( .IN0(\Inst_Mem/n1425 ), .IN1(\Inst_Mem/n1410 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1426 ) );
  MUX \Inst_Mem/U1450  ( .IN0(\Inst_Mem/n1424 ), .IN1(\Inst_Mem/n1417 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1425 ) );
  MUX \Inst_Mem/U1449  ( .IN0(\Inst_Mem/n1423 ), .IN1(\Inst_Mem/n1420 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1424 ) );
  MUX \Inst_Mem/U1448  ( .IN0(\Inst_Mem/n1422 ), .IN1(\Inst_Mem/n1421 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1423 ) );
  MUX \Inst_Mem/U1447  ( .IN0(\Inst_Mem/inst_mem_reg[0][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1422 ) );
  MUX \Inst_Mem/U1446  ( .IN0(\Inst_Mem/inst_mem_reg[2][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1421 ) );
  MUX \Inst_Mem/U1445  ( .IN0(\Inst_Mem/n1419 ), .IN1(\Inst_Mem/n1418 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1420 ) );
  MUX \Inst_Mem/U1444  ( .IN0(\Inst_Mem/inst_mem_reg[4][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1419 ) );
  MUX \Inst_Mem/U1443  ( .IN0(\Inst_Mem/inst_mem_reg[6][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1418 ) );
  MUX \Inst_Mem/U1442  ( .IN0(\Inst_Mem/n1416 ), .IN1(\Inst_Mem/n1413 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1417 ) );
  MUX \Inst_Mem/U1441  ( .IN0(\Inst_Mem/n1415 ), .IN1(\Inst_Mem/n1414 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1416 ) );
  MUX \Inst_Mem/U1440  ( .IN0(\Inst_Mem/inst_mem_reg[8][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1415 ) );
  MUX \Inst_Mem/U1439  ( .IN0(\Inst_Mem/inst_mem_reg[10][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1414 ) );
  MUX \Inst_Mem/U1438  ( .IN0(\Inst_Mem/n1412 ), .IN1(\Inst_Mem/n1411 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1413 ) );
  MUX \Inst_Mem/U1437  ( .IN0(\Inst_Mem/inst_mem_reg[12][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1412 ) );
  MUX \Inst_Mem/U1436  ( .IN0(\Inst_Mem/inst_mem_reg[14][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1411 ) );
  MUX \Inst_Mem/U1435  ( .IN0(\Inst_Mem/n1409 ), .IN1(\Inst_Mem/n1402 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1410 ) );
  MUX \Inst_Mem/U1434  ( .IN0(\Inst_Mem/n1408 ), .IN1(\Inst_Mem/n1405 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1409 ) );
  MUX \Inst_Mem/U1433  ( .IN0(\Inst_Mem/n1407 ), .IN1(\Inst_Mem/n1406 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1408 ) );
  MUX \Inst_Mem/U1432  ( .IN0(\Inst_Mem/inst_mem_reg[16][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1407 ) );
  MUX \Inst_Mem/U1431  ( .IN0(\Inst_Mem/inst_mem_reg[18][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1406 ) );
  MUX \Inst_Mem/U1430  ( .IN0(\Inst_Mem/n1404 ), .IN1(\Inst_Mem/n1403 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1405 ) );
  MUX \Inst_Mem/U1429  ( .IN0(\Inst_Mem/inst_mem_reg[20][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1404 ) );
  MUX \Inst_Mem/U1428  ( .IN0(\Inst_Mem/inst_mem_reg[22][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1403 ) );
  MUX \Inst_Mem/U1427  ( .IN0(\Inst_Mem/n1401 ), .IN1(\Inst_Mem/n1398 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1402 ) );
  MUX \Inst_Mem/U1426  ( .IN0(\Inst_Mem/n1400 ), .IN1(\Inst_Mem/n1399 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1401 ) );
  MUX \Inst_Mem/U1425  ( .IN0(\Inst_Mem/inst_mem_reg[24][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1400 ) );
  MUX \Inst_Mem/U1424  ( .IN0(\Inst_Mem/inst_mem_reg[26][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1399 ) );
  MUX \Inst_Mem/U1423  ( .IN0(\Inst_Mem/n1397 ), .IN1(\Inst_Mem/n1396 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1398 ) );
  MUX \Inst_Mem/U1422  ( .IN0(\Inst_Mem/inst_mem_reg[28][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1397 ) );
  MUX \Inst_Mem/U1421  ( .IN0(\Inst_Mem/inst_mem_reg[30][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1396 ) );
  MUX \Inst_Mem/U1420  ( .IN0(\Inst_Mem/n1394 ), .IN1(\Inst_Mem/n1379 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1395 ) );
  MUX \Inst_Mem/U1419  ( .IN0(\Inst_Mem/n1393 ), .IN1(\Inst_Mem/n1386 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1394 ) );
  MUX \Inst_Mem/U1418  ( .IN0(\Inst_Mem/n1392 ), .IN1(\Inst_Mem/n1389 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1393 ) );
  MUX \Inst_Mem/U1417  ( .IN0(\Inst_Mem/n1391 ), .IN1(\Inst_Mem/n1390 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1392 ) );
  MUX \Inst_Mem/U1416  ( .IN0(\Inst_Mem/inst_mem_reg[32][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1391 ) );
  MUX \Inst_Mem/U1415  ( .IN0(\Inst_Mem/inst_mem_reg[34][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1390 ) );
  MUX \Inst_Mem/U1414  ( .IN0(\Inst_Mem/n1388 ), .IN1(\Inst_Mem/n1387 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1389 ) );
  MUX \Inst_Mem/U1413  ( .IN0(\Inst_Mem/inst_mem_reg[36][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1388 ) );
  MUX \Inst_Mem/U1412  ( .IN0(\Inst_Mem/inst_mem_reg[38][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1387 ) );
  MUX \Inst_Mem/U1411  ( .IN0(\Inst_Mem/n1385 ), .IN1(\Inst_Mem/n1382 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1386 ) );
  MUX \Inst_Mem/U1410  ( .IN0(\Inst_Mem/n1384 ), .IN1(\Inst_Mem/n1383 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1385 ) );
  MUX \Inst_Mem/U1409  ( .IN0(\Inst_Mem/inst_mem_reg[40][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1384 ) );
  MUX \Inst_Mem/U1408  ( .IN0(\Inst_Mem/inst_mem_reg[42][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1383 ) );
  MUX \Inst_Mem/U1407  ( .IN0(\Inst_Mem/n1381 ), .IN1(\Inst_Mem/n1380 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1382 ) );
  MUX \Inst_Mem/U1406  ( .IN0(\Inst_Mem/inst_mem_reg[44][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1381 ) );
  MUX \Inst_Mem/U1405  ( .IN0(\Inst_Mem/inst_mem_reg[46][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1380 ) );
  MUX \Inst_Mem/U1404  ( .IN0(\Inst_Mem/n1378 ), .IN1(\Inst_Mem/n1371 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1379 ) );
  MUX \Inst_Mem/U1403  ( .IN0(\Inst_Mem/n1377 ), .IN1(\Inst_Mem/n1374 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1378 ) );
  MUX \Inst_Mem/U1402  ( .IN0(\Inst_Mem/n1376 ), .IN1(\Inst_Mem/n1375 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1377 ) );
  MUX \Inst_Mem/U1401  ( .IN0(\Inst_Mem/inst_mem_reg[48][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1376 ) );
  MUX \Inst_Mem/U1400  ( .IN0(\Inst_Mem/inst_mem_reg[50][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1375 ) );
  MUX \Inst_Mem/U1399  ( .IN0(\Inst_Mem/n1373 ), .IN1(\Inst_Mem/n1372 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1374 ) );
  MUX \Inst_Mem/U1398  ( .IN0(\Inst_Mem/inst_mem_reg[52][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1373 ) );
  MUX \Inst_Mem/U1397  ( .IN0(\Inst_Mem/inst_mem_reg[54][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1372 ) );
  MUX \Inst_Mem/U1396  ( .IN0(\Inst_Mem/n1370 ), .IN1(\Inst_Mem/n1367 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1371 ) );
  MUX \Inst_Mem/U1395  ( .IN0(\Inst_Mem/n1369 ), .IN1(\Inst_Mem/n1368 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1370 ) );
  MUX \Inst_Mem/U1394  ( .IN0(\Inst_Mem/inst_mem_reg[56][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1369 ) );
  MUX \Inst_Mem/U1393  ( .IN0(\Inst_Mem/inst_mem_reg[58][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1368 ) );
  MUX \Inst_Mem/U1392  ( .IN0(\Inst_Mem/n1366 ), .IN1(\Inst_Mem/n1365 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1367 ) );
  MUX \Inst_Mem/U1391  ( .IN0(\Inst_Mem/inst_mem_reg[60][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1366 ) );
  MUX \Inst_Mem/U1390  ( .IN0(\Inst_Mem/inst_mem_reg[62][22] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][22] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1365 ) );
  MUX \Inst_Mem/U1389  ( .IN0(\Inst_Mem/n1364 ), .IN1(\Inst_Mem/n1333 ), .SEL(
        pc_current[7]), .F(opcode[21]) );
  MUX \Inst_Mem/U1388  ( .IN0(\Inst_Mem/n1363 ), .IN1(\Inst_Mem/n1348 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1364 ) );
  MUX \Inst_Mem/U1387  ( .IN0(\Inst_Mem/n1362 ), .IN1(\Inst_Mem/n1355 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1363 ) );
  MUX \Inst_Mem/U1386  ( .IN0(\Inst_Mem/n1361 ), .IN1(\Inst_Mem/n1358 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1362 ) );
  MUX \Inst_Mem/U1385  ( .IN0(\Inst_Mem/n1360 ), .IN1(\Inst_Mem/n1359 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1361 ) );
  MUX \Inst_Mem/U1384  ( .IN0(\Inst_Mem/inst_mem_reg[0][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1360 ) );
  MUX \Inst_Mem/U1383  ( .IN0(\Inst_Mem/inst_mem_reg[2][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1359 ) );
  MUX \Inst_Mem/U1382  ( .IN0(\Inst_Mem/n1357 ), .IN1(\Inst_Mem/n1356 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1358 ) );
  MUX \Inst_Mem/U1381  ( .IN0(\Inst_Mem/inst_mem_reg[4][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1357 ) );
  MUX \Inst_Mem/U1380  ( .IN0(\Inst_Mem/inst_mem_reg[6][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1356 ) );
  MUX \Inst_Mem/U1379  ( .IN0(\Inst_Mem/n1354 ), .IN1(\Inst_Mem/n1351 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1355 ) );
  MUX \Inst_Mem/U1378  ( .IN0(\Inst_Mem/n1353 ), .IN1(\Inst_Mem/n1352 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1354 ) );
  MUX \Inst_Mem/U1377  ( .IN0(\Inst_Mem/inst_mem_reg[8][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1353 ) );
  MUX \Inst_Mem/U1376  ( .IN0(\Inst_Mem/inst_mem_reg[10][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1352 ) );
  MUX \Inst_Mem/U1375  ( .IN0(\Inst_Mem/n1350 ), .IN1(\Inst_Mem/n1349 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1351 ) );
  MUX \Inst_Mem/U1374  ( .IN0(\Inst_Mem/inst_mem_reg[12][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1350 ) );
  MUX \Inst_Mem/U1373  ( .IN0(\Inst_Mem/inst_mem_reg[14][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1349 ) );
  MUX \Inst_Mem/U1372  ( .IN0(\Inst_Mem/n1347 ), .IN1(\Inst_Mem/n1340 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1348 ) );
  MUX \Inst_Mem/U1371  ( .IN0(\Inst_Mem/n1346 ), .IN1(\Inst_Mem/n1343 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1347 ) );
  MUX \Inst_Mem/U1370  ( .IN0(\Inst_Mem/n1345 ), .IN1(\Inst_Mem/n1344 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1346 ) );
  MUX \Inst_Mem/U1369  ( .IN0(\Inst_Mem/inst_mem_reg[16][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1345 ) );
  MUX \Inst_Mem/U1368  ( .IN0(\Inst_Mem/inst_mem_reg[18][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1344 ) );
  MUX \Inst_Mem/U1367  ( .IN0(\Inst_Mem/n1342 ), .IN1(\Inst_Mem/n1341 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1343 ) );
  MUX \Inst_Mem/U1366  ( .IN0(\Inst_Mem/inst_mem_reg[20][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1342 ) );
  MUX \Inst_Mem/U1365  ( .IN0(\Inst_Mem/inst_mem_reg[22][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1341 ) );
  MUX \Inst_Mem/U1364  ( .IN0(\Inst_Mem/n1339 ), .IN1(\Inst_Mem/n1336 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1340 ) );
  MUX \Inst_Mem/U1363  ( .IN0(\Inst_Mem/n1338 ), .IN1(\Inst_Mem/n1337 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1339 ) );
  MUX \Inst_Mem/U1362  ( .IN0(\Inst_Mem/inst_mem_reg[24][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1338 ) );
  MUX \Inst_Mem/U1361  ( .IN0(\Inst_Mem/inst_mem_reg[26][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1337 ) );
  MUX \Inst_Mem/U1360  ( .IN0(\Inst_Mem/n1335 ), .IN1(\Inst_Mem/n1334 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1336 ) );
  MUX \Inst_Mem/U1359  ( .IN0(\Inst_Mem/inst_mem_reg[28][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1335 ) );
  MUX \Inst_Mem/U1358  ( .IN0(\Inst_Mem/inst_mem_reg[30][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1334 ) );
  MUX \Inst_Mem/U1357  ( .IN0(\Inst_Mem/n1332 ), .IN1(\Inst_Mem/n1317 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1333 ) );
  MUX \Inst_Mem/U1356  ( .IN0(\Inst_Mem/n1331 ), .IN1(\Inst_Mem/n1324 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1332 ) );
  MUX \Inst_Mem/U1355  ( .IN0(\Inst_Mem/n1330 ), .IN1(\Inst_Mem/n1327 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1331 ) );
  MUX \Inst_Mem/U1354  ( .IN0(\Inst_Mem/n1329 ), .IN1(\Inst_Mem/n1328 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1330 ) );
  MUX \Inst_Mem/U1353  ( .IN0(\Inst_Mem/inst_mem_reg[32][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1329 ) );
  MUX \Inst_Mem/U1352  ( .IN0(\Inst_Mem/inst_mem_reg[34][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1328 ) );
  MUX \Inst_Mem/U1351  ( .IN0(\Inst_Mem/n1326 ), .IN1(\Inst_Mem/n1325 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1327 ) );
  MUX \Inst_Mem/U1350  ( .IN0(\Inst_Mem/inst_mem_reg[36][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1326 ) );
  MUX \Inst_Mem/U1349  ( .IN0(\Inst_Mem/inst_mem_reg[38][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1325 ) );
  MUX \Inst_Mem/U1348  ( .IN0(\Inst_Mem/n1323 ), .IN1(\Inst_Mem/n1320 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1324 ) );
  MUX \Inst_Mem/U1347  ( .IN0(\Inst_Mem/n1322 ), .IN1(\Inst_Mem/n1321 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1323 ) );
  MUX \Inst_Mem/U1346  ( .IN0(\Inst_Mem/inst_mem_reg[40][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1322 ) );
  MUX \Inst_Mem/U1345  ( .IN0(\Inst_Mem/inst_mem_reg[42][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1321 ) );
  MUX \Inst_Mem/U1344  ( .IN0(\Inst_Mem/n1319 ), .IN1(\Inst_Mem/n1318 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1320 ) );
  MUX \Inst_Mem/U1343  ( .IN0(\Inst_Mem/inst_mem_reg[44][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1319 ) );
  MUX \Inst_Mem/U1342  ( .IN0(\Inst_Mem/inst_mem_reg[46][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1318 ) );
  MUX \Inst_Mem/U1341  ( .IN0(\Inst_Mem/n1316 ), .IN1(\Inst_Mem/n1309 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1317 ) );
  MUX \Inst_Mem/U1340  ( .IN0(\Inst_Mem/n1315 ), .IN1(\Inst_Mem/n1312 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1316 ) );
  MUX \Inst_Mem/U1339  ( .IN0(\Inst_Mem/n1314 ), .IN1(\Inst_Mem/n1313 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1315 ) );
  MUX \Inst_Mem/U1338  ( .IN0(\Inst_Mem/inst_mem_reg[48][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1314 ) );
  MUX \Inst_Mem/U1337  ( .IN0(\Inst_Mem/inst_mem_reg[50][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1313 ) );
  MUX \Inst_Mem/U1336  ( .IN0(\Inst_Mem/n1311 ), .IN1(\Inst_Mem/n1310 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1312 ) );
  MUX \Inst_Mem/U1335  ( .IN0(\Inst_Mem/inst_mem_reg[52][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1311 ) );
  MUX \Inst_Mem/U1334  ( .IN0(\Inst_Mem/inst_mem_reg[54][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1310 ) );
  MUX \Inst_Mem/U1333  ( .IN0(\Inst_Mem/n1308 ), .IN1(\Inst_Mem/n1305 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1309 ) );
  MUX \Inst_Mem/U1332  ( .IN0(\Inst_Mem/n1307 ), .IN1(\Inst_Mem/n1306 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1308 ) );
  MUX \Inst_Mem/U1331  ( .IN0(\Inst_Mem/inst_mem_reg[56][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1307 ) );
  MUX \Inst_Mem/U1330  ( .IN0(\Inst_Mem/inst_mem_reg[58][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1306 ) );
  MUX \Inst_Mem/U1329  ( .IN0(\Inst_Mem/n1304 ), .IN1(\Inst_Mem/n1303 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1305 ) );
  MUX \Inst_Mem/U1328  ( .IN0(\Inst_Mem/inst_mem_reg[60][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1304 ) );
  MUX \Inst_Mem/U1327  ( .IN0(\Inst_Mem/inst_mem_reg[62][21] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][21] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1303 ) );
  MUX \Inst_Mem/U1326  ( .IN0(\Inst_Mem/n1302 ), .IN1(\Inst_Mem/n1271 ), .SEL(
        pc_current[7]), .F(opcode[20]) );
  MUX \Inst_Mem/U1325  ( .IN0(\Inst_Mem/n1301 ), .IN1(\Inst_Mem/n1286 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1302 ) );
  MUX \Inst_Mem/U1324  ( .IN0(\Inst_Mem/n1300 ), .IN1(\Inst_Mem/n1293 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1301 ) );
  MUX \Inst_Mem/U1323  ( .IN0(\Inst_Mem/n1299 ), .IN1(\Inst_Mem/n1296 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1300 ) );
  MUX \Inst_Mem/U1322  ( .IN0(\Inst_Mem/n1298 ), .IN1(\Inst_Mem/n1297 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1299 ) );
  MUX \Inst_Mem/U1321  ( .IN0(\Inst_Mem/inst_mem_reg[0][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1298 ) );
  MUX \Inst_Mem/U1320  ( .IN0(\Inst_Mem/inst_mem_reg[2][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1297 ) );
  MUX \Inst_Mem/U1319  ( .IN0(\Inst_Mem/n1295 ), .IN1(\Inst_Mem/n1294 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1296 ) );
  MUX \Inst_Mem/U1318  ( .IN0(\Inst_Mem/inst_mem_reg[4][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1295 ) );
  MUX \Inst_Mem/U1317  ( .IN0(\Inst_Mem/inst_mem_reg[6][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1294 ) );
  MUX \Inst_Mem/U1316  ( .IN0(\Inst_Mem/n1292 ), .IN1(\Inst_Mem/n1289 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1293 ) );
  MUX \Inst_Mem/U1315  ( .IN0(\Inst_Mem/n1291 ), .IN1(\Inst_Mem/n1290 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1292 ) );
  MUX \Inst_Mem/U1314  ( .IN0(\Inst_Mem/inst_mem_reg[8][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1291 ) );
  MUX \Inst_Mem/U1313  ( .IN0(\Inst_Mem/inst_mem_reg[10][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1290 ) );
  MUX \Inst_Mem/U1312  ( .IN0(\Inst_Mem/n1288 ), .IN1(\Inst_Mem/n1287 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1289 ) );
  MUX \Inst_Mem/U1311  ( .IN0(\Inst_Mem/inst_mem_reg[12][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1288 ) );
  MUX \Inst_Mem/U1310  ( .IN0(\Inst_Mem/inst_mem_reg[14][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1287 ) );
  MUX \Inst_Mem/U1309  ( .IN0(\Inst_Mem/n1285 ), .IN1(\Inst_Mem/n1278 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1286 ) );
  MUX \Inst_Mem/U1308  ( .IN0(\Inst_Mem/n1284 ), .IN1(\Inst_Mem/n1281 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1285 ) );
  MUX \Inst_Mem/U1307  ( .IN0(\Inst_Mem/n1283 ), .IN1(\Inst_Mem/n1282 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1284 ) );
  MUX \Inst_Mem/U1306  ( .IN0(\Inst_Mem/inst_mem_reg[16][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1283 ) );
  MUX \Inst_Mem/U1305  ( .IN0(\Inst_Mem/inst_mem_reg[18][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1282 ) );
  MUX \Inst_Mem/U1304  ( .IN0(\Inst_Mem/n1280 ), .IN1(\Inst_Mem/n1279 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1281 ) );
  MUX \Inst_Mem/U1303  ( .IN0(\Inst_Mem/inst_mem_reg[20][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1280 ) );
  MUX \Inst_Mem/U1302  ( .IN0(\Inst_Mem/inst_mem_reg[22][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1279 ) );
  MUX \Inst_Mem/U1301  ( .IN0(\Inst_Mem/n1277 ), .IN1(\Inst_Mem/n1274 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1278 ) );
  MUX \Inst_Mem/U1300  ( .IN0(\Inst_Mem/n1276 ), .IN1(\Inst_Mem/n1275 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1277 ) );
  MUX \Inst_Mem/U1299  ( .IN0(\Inst_Mem/inst_mem_reg[24][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1276 ) );
  MUX \Inst_Mem/U1298  ( .IN0(\Inst_Mem/inst_mem_reg[26][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1275 ) );
  MUX \Inst_Mem/U1297  ( .IN0(\Inst_Mem/n1273 ), .IN1(\Inst_Mem/n1272 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1274 ) );
  MUX \Inst_Mem/U1296  ( .IN0(\Inst_Mem/inst_mem_reg[28][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1273 ) );
  MUX \Inst_Mem/U1295  ( .IN0(\Inst_Mem/inst_mem_reg[30][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1272 ) );
  MUX \Inst_Mem/U1294  ( .IN0(\Inst_Mem/n1270 ), .IN1(\Inst_Mem/n1255 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1271 ) );
  MUX \Inst_Mem/U1293  ( .IN0(\Inst_Mem/n1269 ), .IN1(\Inst_Mem/n1262 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1270 ) );
  MUX \Inst_Mem/U1292  ( .IN0(\Inst_Mem/n1268 ), .IN1(\Inst_Mem/n1265 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1269 ) );
  MUX \Inst_Mem/U1291  ( .IN0(\Inst_Mem/n1267 ), .IN1(\Inst_Mem/n1266 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1268 ) );
  MUX \Inst_Mem/U1290  ( .IN0(\Inst_Mem/inst_mem_reg[32][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1267 ) );
  MUX \Inst_Mem/U1289  ( .IN0(\Inst_Mem/inst_mem_reg[34][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1266 ) );
  MUX \Inst_Mem/U1288  ( .IN0(\Inst_Mem/n1264 ), .IN1(\Inst_Mem/n1263 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1265 ) );
  MUX \Inst_Mem/U1287  ( .IN0(\Inst_Mem/inst_mem_reg[36][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1264 ) );
  MUX \Inst_Mem/U1286  ( .IN0(\Inst_Mem/inst_mem_reg[38][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1263 ) );
  MUX \Inst_Mem/U1285  ( .IN0(\Inst_Mem/n1261 ), .IN1(\Inst_Mem/n1258 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1262 ) );
  MUX \Inst_Mem/U1284  ( .IN0(\Inst_Mem/n1260 ), .IN1(\Inst_Mem/n1259 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1261 ) );
  MUX \Inst_Mem/U1283  ( .IN0(\Inst_Mem/inst_mem_reg[40][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1260 ) );
  MUX \Inst_Mem/U1282  ( .IN0(\Inst_Mem/inst_mem_reg[42][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1259 ) );
  MUX \Inst_Mem/U1281  ( .IN0(\Inst_Mem/n1257 ), .IN1(\Inst_Mem/n1256 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1258 ) );
  MUX \Inst_Mem/U1280  ( .IN0(\Inst_Mem/inst_mem_reg[44][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1257 ) );
  MUX \Inst_Mem/U1279  ( .IN0(\Inst_Mem/inst_mem_reg[46][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1256 ) );
  MUX \Inst_Mem/U1278  ( .IN0(\Inst_Mem/n1254 ), .IN1(\Inst_Mem/n1247 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1255 ) );
  MUX \Inst_Mem/U1277  ( .IN0(\Inst_Mem/n1253 ), .IN1(\Inst_Mem/n1250 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1254 ) );
  MUX \Inst_Mem/U1276  ( .IN0(\Inst_Mem/n1252 ), .IN1(\Inst_Mem/n1251 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1253 ) );
  MUX \Inst_Mem/U1275  ( .IN0(\Inst_Mem/inst_mem_reg[48][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1252 ) );
  MUX \Inst_Mem/U1274  ( .IN0(\Inst_Mem/inst_mem_reg[50][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1251 ) );
  MUX \Inst_Mem/U1273  ( .IN0(\Inst_Mem/n1249 ), .IN1(\Inst_Mem/n1248 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1250 ) );
  MUX \Inst_Mem/U1272  ( .IN0(\Inst_Mem/inst_mem_reg[52][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1249 ) );
  MUX \Inst_Mem/U1271  ( .IN0(\Inst_Mem/inst_mem_reg[54][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1248 ) );
  MUX \Inst_Mem/U1270  ( .IN0(\Inst_Mem/n1246 ), .IN1(\Inst_Mem/n1243 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1247 ) );
  MUX \Inst_Mem/U1269  ( .IN0(\Inst_Mem/n1245 ), .IN1(\Inst_Mem/n1244 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1246 ) );
  MUX \Inst_Mem/U1268  ( .IN0(\Inst_Mem/inst_mem_reg[56][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1245 ) );
  MUX \Inst_Mem/U1267  ( .IN0(\Inst_Mem/inst_mem_reg[58][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1244 ) );
  MUX \Inst_Mem/U1266  ( .IN0(\Inst_Mem/n1242 ), .IN1(\Inst_Mem/n1241 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1243 ) );
  MUX \Inst_Mem/U1265  ( .IN0(\Inst_Mem/inst_mem_reg[60][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1242 ) );
  MUX \Inst_Mem/U1264  ( .IN0(\Inst_Mem/inst_mem_reg[62][20] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][20] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1241 ) );
  MUX \Inst_Mem/U1263  ( .IN0(\Inst_Mem/n1240 ), .IN1(\Inst_Mem/n1209 ), .SEL(
        pc_current[7]), .F(opcode[19]) );
  MUX \Inst_Mem/U1262  ( .IN0(\Inst_Mem/n1239 ), .IN1(\Inst_Mem/n1224 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1240 ) );
  MUX \Inst_Mem/U1261  ( .IN0(\Inst_Mem/n1238 ), .IN1(\Inst_Mem/n1231 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1239 ) );
  MUX \Inst_Mem/U1260  ( .IN0(\Inst_Mem/n1237 ), .IN1(\Inst_Mem/n1234 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1238 ) );
  MUX \Inst_Mem/U1259  ( .IN0(\Inst_Mem/n1236 ), .IN1(\Inst_Mem/n1235 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1237 ) );
  MUX \Inst_Mem/U1258  ( .IN0(\Inst_Mem/inst_mem_reg[0][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1236 ) );
  MUX \Inst_Mem/U1257  ( .IN0(\Inst_Mem/inst_mem_reg[2][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1235 ) );
  MUX \Inst_Mem/U1256  ( .IN0(\Inst_Mem/n1233 ), .IN1(\Inst_Mem/n1232 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1234 ) );
  MUX \Inst_Mem/U1255  ( .IN0(\Inst_Mem/inst_mem_reg[4][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1233 ) );
  MUX \Inst_Mem/U1254  ( .IN0(\Inst_Mem/inst_mem_reg[6][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1232 ) );
  MUX \Inst_Mem/U1253  ( .IN0(\Inst_Mem/n1230 ), .IN1(\Inst_Mem/n1227 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1231 ) );
  MUX \Inst_Mem/U1252  ( .IN0(\Inst_Mem/n1229 ), .IN1(\Inst_Mem/n1228 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1230 ) );
  MUX \Inst_Mem/U1251  ( .IN0(\Inst_Mem/inst_mem_reg[8][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1229 ) );
  MUX \Inst_Mem/U1250  ( .IN0(\Inst_Mem/inst_mem_reg[10][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1228 ) );
  MUX \Inst_Mem/U1249  ( .IN0(\Inst_Mem/n1226 ), .IN1(\Inst_Mem/n1225 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1227 ) );
  MUX \Inst_Mem/U1248  ( .IN0(\Inst_Mem/inst_mem_reg[12][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1226 ) );
  MUX \Inst_Mem/U1247  ( .IN0(\Inst_Mem/inst_mem_reg[14][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1225 ) );
  MUX \Inst_Mem/U1246  ( .IN0(\Inst_Mem/n1223 ), .IN1(\Inst_Mem/n1216 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1224 ) );
  MUX \Inst_Mem/U1245  ( .IN0(\Inst_Mem/n1222 ), .IN1(\Inst_Mem/n1219 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1223 ) );
  MUX \Inst_Mem/U1244  ( .IN0(\Inst_Mem/n1221 ), .IN1(\Inst_Mem/n1220 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1222 ) );
  MUX \Inst_Mem/U1243  ( .IN0(\Inst_Mem/inst_mem_reg[16][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1221 ) );
  MUX \Inst_Mem/U1242  ( .IN0(\Inst_Mem/inst_mem_reg[18][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1220 ) );
  MUX \Inst_Mem/U1241  ( .IN0(\Inst_Mem/n1218 ), .IN1(\Inst_Mem/n1217 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1219 ) );
  MUX \Inst_Mem/U1240  ( .IN0(\Inst_Mem/inst_mem_reg[20][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1218 ) );
  MUX \Inst_Mem/U1239  ( .IN0(\Inst_Mem/inst_mem_reg[22][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1217 ) );
  MUX \Inst_Mem/U1238  ( .IN0(\Inst_Mem/n1215 ), .IN1(\Inst_Mem/n1212 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1216 ) );
  MUX \Inst_Mem/U1237  ( .IN0(\Inst_Mem/n1214 ), .IN1(\Inst_Mem/n1213 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1215 ) );
  MUX \Inst_Mem/U1236  ( .IN0(\Inst_Mem/inst_mem_reg[24][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1214 ) );
  MUX \Inst_Mem/U1235  ( .IN0(\Inst_Mem/inst_mem_reg[26][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1213 ) );
  MUX \Inst_Mem/U1234  ( .IN0(\Inst_Mem/n1211 ), .IN1(\Inst_Mem/n1210 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1212 ) );
  MUX \Inst_Mem/U1233  ( .IN0(\Inst_Mem/inst_mem_reg[28][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1211 ) );
  MUX \Inst_Mem/U1232  ( .IN0(\Inst_Mem/inst_mem_reg[30][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1210 ) );
  MUX \Inst_Mem/U1231  ( .IN0(\Inst_Mem/n1208 ), .IN1(\Inst_Mem/n1193 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1209 ) );
  MUX \Inst_Mem/U1230  ( .IN0(\Inst_Mem/n1207 ), .IN1(\Inst_Mem/n1200 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1208 ) );
  MUX \Inst_Mem/U1229  ( .IN0(\Inst_Mem/n1206 ), .IN1(\Inst_Mem/n1203 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1207 ) );
  MUX \Inst_Mem/U1228  ( .IN0(\Inst_Mem/n1205 ), .IN1(\Inst_Mem/n1204 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1206 ) );
  MUX \Inst_Mem/U1227  ( .IN0(\Inst_Mem/inst_mem_reg[32][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1205 ) );
  MUX \Inst_Mem/U1226  ( .IN0(\Inst_Mem/inst_mem_reg[34][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1204 ) );
  MUX \Inst_Mem/U1225  ( .IN0(\Inst_Mem/n1202 ), .IN1(\Inst_Mem/n1201 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1203 ) );
  MUX \Inst_Mem/U1224  ( .IN0(\Inst_Mem/inst_mem_reg[36][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1202 ) );
  MUX \Inst_Mem/U1223  ( .IN0(\Inst_Mem/inst_mem_reg[38][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1201 ) );
  MUX \Inst_Mem/U1222  ( .IN0(\Inst_Mem/n1199 ), .IN1(\Inst_Mem/n1196 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1200 ) );
  MUX \Inst_Mem/U1221  ( .IN0(\Inst_Mem/n1198 ), .IN1(\Inst_Mem/n1197 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1199 ) );
  MUX \Inst_Mem/U1220  ( .IN0(\Inst_Mem/inst_mem_reg[40][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1198 ) );
  MUX \Inst_Mem/U1219  ( .IN0(\Inst_Mem/inst_mem_reg[42][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1197 ) );
  MUX \Inst_Mem/U1218  ( .IN0(\Inst_Mem/n1195 ), .IN1(\Inst_Mem/n1194 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1196 ) );
  MUX \Inst_Mem/U1217  ( .IN0(\Inst_Mem/inst_mem_reg[44][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1195 ) );
  MUX \Inst_Mem/U1216  ( .IN0(\Inst_Mem/inst_mem_reg[46][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1194 ) );
  MUX \Inst_Mem/U1215  ( .IN0(\Inst_Mem/n1192 ), .IN1(\Inst_Mem/n1185 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1193 ) );
  MUX \Inst_Mem/U1214  ( .IN0(\Inst_Mem/n1191 ), .IN1(\Inst_Mem/n1188 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1192 ) );
  MUX \Inst_Mem/U1213  ( .IN0(\Inst_Mem/n1190 ), .IN1(\Inst_Mem/n1189 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1191 ) );
  MUX \Inst_Mem/U1212  ( .IN0(\Inst_Mem/inst_mem_reg[48][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1190 ) );
  MUX \Inst_Mem/U1211  ( .IN0(\Inst_Mem/inst_mem_reg[50][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1189 ) );
  MUX \Inst_Mem/U1210  ( .IN0(\Inst_Mem/n1187 ), .IN1(\Inst_Mem/n1186 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1188 ) );
  MUX \Inst_Mem/U1209  ( .IN0(\Inst_Mem/inst_mem_reg[52][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1187 ) );
  MUX \Inst_Mem/U1208  ( .IN0(\Inst_Mem/inst_mem_reg[54][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1186 ) );
  MUX \Inst_Mem/U1207  ( .IN0(\Inst_Mem/n1184 ), .IN1(\Inst_Mem/n1181 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1185 ) );
  MUX \Inst_Mem/U1206  ( .IN0(\Inst_Mem/n1183 ), .IN1(\Inst_Mem/n1182 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1184 ) );
  MUX \Inst_Mem/U1205  ( .IN0(\Inst_Mem/inst_mem_reg[56][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1183 ) );
  MUX \Inst_Mem/U1204  ( .IN0(\Inst_Mem/inst_mem_reg[58][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1182 ) );
  MUX \Inst_Mem/U1203  ( .IN0(\Inst_Mem/n1180 ), .IN1(\Inst_Mem/n1179 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1181 ) );
  MUX \Inst_Mem/U1202  ( .IN0(\Inst_Mem/inst_mem_reg[60][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1180 ) );
  MUX \Inst_Mem/U1201  ( .IN0(\Inst_Mem/inst_mem_reg[62][19] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][19] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1179 ) );
  MUX \Inst_Mem/U1200  ( .IN0(\Inst_Mem/n1178 ), .IN1(\Inst_Mem/n1147 ), .SEL(
        pc_current[7]), .F(opcode[18]) );
  MUX \Inst_Mem/U1199  ( .IN0(\Inst_Mem/n1177 ), .IN1(\Inst_Mem/n1162 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1178 ) );
  MUX \Inst_Mem/U1198  ( .IN0(\Inst_Mem/n1176 ), .IN1(\Inst_Mem/n1169 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1177 ) );
  MUX \Inst_Mem/U1197  ( .IN0(\Inst_Mem/n1175 ), .IN1(\Inst_Mem/n1172 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1176 ) );
  MUX \Inst_Mem/U1196  ( .IN0(\Inst_Mem/n1174 ), .IN1(\Inst_Mem/n1173 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1175 ) );
  MUX \Inst_Mem/U1195  ( .IN0(\Inst_Mem/inst_mem_reg[0][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1174 ) );
  MUX \Inst_Mem/U1194  ( .IN0(\Inst_Mem/inst_mem_reg[2][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1173 ) );
  MUX \Inst_Mem/U1193  ( .IN0(\Inst_Mem/n1171 ), .IN1(\Inst_Mem/n1170 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1172 ) );
  MUX \Inst_Mem/U1192  ( .IN0(\Inst_Mem/inst_mem_reg[4][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1171 ) );
  MUX \Inst_Mem/U1191  ( .IN0(\Inst_Mem/inst_mem_reg[6][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1170 ) );
  MUX \Inst_Mem/U1190  ( .IN0(\Inst_Mem/n1168 ), .IN1(\Inst_Mem/n1165 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1169 ) );
  MUX \Inst_Mem/U1189  ( .IN0(\Inst_Mem/n1167 ), .IN1(\Inst_Mem/n1166 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1168 ) );
  MUX \Inst_Mem/U1188  ( .IN0(\Inst_Mem/inst_mem_reg[8][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1167 ) );
  MUX \Inst_Mem/U1187  ( .IN0(\Inst_Mem/inst_mem_reg[10][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1166 ) );
  MUX \Inst_Mem/U1186  ( .IN0(\Inst_Mem/n1164 ), .IN1(\Inst_Mem/n1163 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1165 ) );
  MUX \Inst_Mem/U1185  ( .IN0(\Inst_Mem/inst_mem_reg[12][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1164 ) );
  MUX \Inst_Mem/U1184  ( .IN0(\Inst_Mem/inst_mem_reg[14][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1163 ) );
  MUX \Inst_Mem/U1183  ( .IN0(\Inst_Mem/n1161 ), .IN1(\Inst_Mem/n1154 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1162 ) );
  MUX \Inst_Mem/U1182  ( .IN0(\Inst_Mem/n1160 ), .IN1(\Inst_Mem/n1157 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1161 ) );
  MUX \Inst_Mem/U1181  ( .IN0(\Inst_Mem/n1159 ), .IN1(\Inst_Mem/n1158 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1160 ) );
  MUX \Inst_Mem/U1180  ( .IN0(\Inst_Mem/inst_mem_reg[16][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1159 ) );
  MUX \Inst_Mem/U1179  ( .IN0(\Inst_Mem/inst_mem_reg[18][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1158 ) );
  MUX \Inst_Mem/U1178  ( .IN0(\Inst_Mem/n1156 ), .IN1(\Inst_Mem/n1155 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1157 ) );
  MUX \Inst_Mem/U1177  ( .IN0(\Inst_Mem/inst_mem_reg[20][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1156 ) );
  MUX \Inst_Mem/U1176  ( .IN0(\Inst_Mem/inst_mem_reg[22][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1155 ) );
  MUX \Inst_Mem/U1175  ( .IN0(\Inst_Mem/n1153 ), .IN1(\Inst_Mem/n1150 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1154 ) );
  MUX \Inst_Mem/U1174  ( .IN0(\Inst_Mem/n1152 ), .IN1(\Inst_Mem/n1151 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1153 ) );
  MUX \Inst_Mem/U1173  ( .IN0(\Inst_Mem/inst_mem_reg[24][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1152 ) );
  MUX \Inst_Mem/U1172  ( .IN0(\Inst_Mem/inst_mem_reg[26][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1151 ) );
  MUX \Inst_Mem/U1171  ( .IN0(\Inst_Mem/n1149 ), .IN1(\Inst_Mem/n1148 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1150 ) );
  MUX \Inst_Mem/U1170  ( .IN0(\Inst_Mem/inst_mem_reg[28][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1149 ) );
  MUX \Inst_Mem/U1169  ( .IN0(\Inst_Mem/inst_mem_reg[30][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1148 ) );
  MUX \Inst_Mem/U1168  ( .IN0(\Inst_Mem/n1146 ), .IN1(\Inst_Mem/n1131 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1147 ) );
  MUX \Inst_Mem/U1167  ( .IN0(\Inst_Mem/n1145 ), .IN1(\Inst_Mem/n1138 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1146 ) );
  MUX \Inst_Mem/U1166  ( .IN0(\Inst_Mem/n1144 ), .IN1(\Inst_Mem/n1141 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1145 ) );
  MUX \Inst_Mem/U1165  ( .IN0(\Inst_Mem/n1143 ), .IN1(\Inst_Mem/n1142 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1144 ) );
  MUX \Inst_Mem/U1164  ( .IN0(\Inst_Mem/inst_mem_reg[32][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1143 ) );
  MUX \Inst_Mem/U1163  ( .IN0(\Inst_Mem/inst_mem_reg[34][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1142 ) );
  MUX \Inst_Mem/U1162  ( .IN0(\Inst_Mem/n1140 ), .IN1(\Inst_Mem/n1139 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1141 ) );
  MUX \Inst_Mem/U1161  ( .IN0(\Inst_Mem/inst_mem_reg[36][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1140 ) );
  MUX \Inst_Mem/U1160  ( .IN0(\Inst_Mem/inst_mem_reg[38][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1139 ) );
  MUX \Inst_Mem/U1159  ( .IN0(\Inst_Mem/n1137 ), .IN1(\Inst_Mem/n1134 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1138 ) );
  MUX \Inst_Mem/U1158  ( .IN0(\Inst_Mem/n1136 ), .IN1(\Inst_Mem/n1135 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1137 ) );
  MUX \Inst_Mem/U1157  ( .IN0(\Inst_Mem/inst_mem_reg[40][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1136 ) );
  MUX \Inst_Mem/U1156  ( .IN0(\Inst_Mem/inst_mem_reg[42][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1135 ) );
  MUX \Inst_Mem/U1155  ( .IN0(\Inst_Mem/n1133 ), .IN1(\Inst_Mem/n1132 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1134 ) );
  MUX \Inst_Mem/U1154  ( .IN0(\Inst_Mem/inst_mem_reg[44][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1133 ) );
  MUX \Inst_Mem/U1153  ( .IN0(\Inst_Mem/inst_mem_reg[46][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1132 ) );
  MUX \Inst_Mem/U1152  ( .IN0(\Inst_Mem/n1130 ), .IN1(\Inst_Mem/n1123 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1131 ) );
  MUX \Inst_Mem/U1151  ( .IN0(\Inst_Mem/n1129 ), .IN1(\Inst_Mem/n1126 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1130 ) );
  MUX \Inst_Mem/U1150  ( .IN0(\Inst_Mem/n1128 ), .IN1(\Inst_Mem/n1127 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1129 ) );
  MUX \Inst_Mem/U1149  ( .IN0(\Inst_Mem/inst_mem_reg[48][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1128 ) );
  MUX \Inst_Mem/U1148  ( .IN0(\Inst_Mem/inst_mem_reg[50][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1127 ) );
  MUX \Inst_Mem/U1147  ( .IN0(\Inst_Mem/n1125 ), .IN1(\Inst_Mem/n1124 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1126 ) );
  MUX \Inst_Mem/U1146  ( .IN0(\Inst_Mem/inst_mem_reg[52][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1125 ) );
  MUX \Inst_Mem/U1145  ( .IN0(\Inst_Mem/inst_mem_reg[54][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1124 ) );
  MUX \Inst_Mem/U1144  ( .IN0(\Inst_Mem/n1122 ), .IN1(\Inst_Mem/n1119 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1123 ) );
  MUX \Inst_Mem/U1143  ( .IN0(\Inst_Mem/n1121 ), .IN1(\Inst_Mem/n1120 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1122 ) );
  MUX \Inst_Mem/U1142  ( .IN0(\Inst_Mem/inst_mem_reg[56][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1121 ) );
  MUX \Inst_Mem/U1141  ( .IN0(\Inst_Mem/inst_mem_reg[58][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1120 ) );
  MUX \Inst_Mem/U1140  ( .IN0(\Inst_Mem/n1118 ), .IN1(\Inst_Mem/n1117 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1119 ) );
  MUX \Inst_Mem/U1139  ( .IN0(\Inst_Mem/inst_mem_reg[60][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1118 ) );
  MUX \Inst_Mem/U1138  ( .IN0(\Inst_Mem/inst_mem_reg[62][18] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][18] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1117 ) );
  MUX \Inst_Mem/U1137  ( .IN0(\Inst_Mem/n1116 ), .IN1(\Inst_Mem/n1085 ), .SEL(
        pc_current[7]), .F(opcode[17]) );
  MUX \Inst_Mem/U1136  ( .IN0(\Inst_Mem/n1115 ), .IN1(\Inst_Mem/n1100 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1116 ) );
  MUX \Inst_Mem/U1135  ( .IN0(\Inst_Mem/n1114 ), .IN1(\Inst_Mem/n1107 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1115 ) );
  MUX \Inst_Mem/U1134  ( .IN0(\Inst_Mem/n1113 ), .IN1(\Inst_Mem/n1110 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1114 ) );
  MUX \Inst_Mem/U1133  ( .IN0(\Inst_Mem/n1112 ), .IN1(\Inst_Mem/n1111 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1113 ) );
  MUX \Inst_Mem/U1132  ( .IN0(\Inst_Mem/inst_mem_reg[0][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1112 ) );
  MUX \Inst_Mem/U1131  ( .IN0(\Inst_Mem/inst_mem_reg[2][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1111 ) );
  MUX \Inst_Mem/U1130  ( .IN0(\Inst_Mem/n1109 ), .IN1(\Inst_Mem/n1108 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1110 ) );
  MUX \Inst_Mem/U1129  ( .IN0(\Inst_Mem/inst_mem_reg[4][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1109 ) );
  MUX \Inst_Mem/U1128  ( .IN0(\Inst_Mem/inst_mem_reg[6][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1108 ) );
  MUX \Inst_Mem/U1127  ( .IN0(\Inst_Mem/n1106 ), .IN1(\Inst_Mem/n1103 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1107 ) );
  MUX \Inst_Mem/U1126  ( .IN0(\Inst_Mem/n1105 ), .IN1(\Inst_Mem/n1104 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1106 ) );
  MUX \Inst_Mem/U1125  ( .IN0(\Inst_Mem/inst_mem_reg[8][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1105 ) );
  MUX \Inst_Mem/U1124  ( .IN0(\Inst_Mem/inst_mem_reg[10][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1104 ) );
  MUX \Inst_Mem/U1123  ( .IN0(\Inst_Mem/n1102 ), .IN1(\Inst_Mem/n1101 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1103 ) );
  MUX \Inst_Mem/U1122  ( .IN0(\Inst_Mem/inst_mem_reg[12][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1102 ) );
  MUX \Inst_Mem/U1121  ( .IN0(\Inst_Mem/inst_mem_reg[14][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1101 ) );
  MUX \Inst_Mem/U1120  ( .IN0(\Inst_Mem/n1099 ), .IN1(\Inst_Mem/n1092 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1100 ) );
  MUX \Inst_Mem/U1119  ( .IN0(\Inst_Mem/n1098 ), .IN1(\Inst_Mem/n1095 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1099 ) );
  MUX \Inst_Mem/U1118  ( .IN0(\Inst_Mem/n1097 ), .IN1(\Inst_Mem/n1096 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1098 ) );
  MUX \Inst_Mem/U1117  ( .IN0(\Inst_Mem/inst_mem_reg[16][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1097 ) );
  MUX \Inst_Mem/U1116  ( .IN0(\Inst_Mem/inst_mem_reg[18][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1096 ) );
  MUX \Inst_Mem/U1115  ( .IN0(\Inst_Mem/n1094 ), .IN1(\Inst_Mem/n1093 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1095 ) );
  MUX \Inst_Mem/U1114  ( .IN0(\Inst_Mem/inst_mem_reg[20][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1094 ) );
  MUX \Inst_Mem/U1113  ( .IN0(\Inst_Mem/inst_mem_reg[22][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1093 ) );
  MUX \Inst_Mem/U1112  ( .IN0(\Inst_Mem/n1091 ), .IN1(\Inst_Mem/n1088 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1092 ) );
  MUX \Inst_Mem/U1111  ( .IN0(\Inst_Mem/n1090 ), .IN1(\Inst_Mem/n1089 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1091 ) );
  MUX \Inst_Mem/U1110  ( .IN0(\Inst_Mem/inst_mem_reg[24][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1090 ) );
  MUX \Inst_Mem/U1109  ( .IN0(\Inst_Mem/inst_mem_reg[26][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1089 ) );
  MUX \Inst_Mem/U1108  ( .IN0(\Inst_Mem/n1087 ), .IN1(\Inst_Mem/n1086 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1088 ) );
  MUX \Inst_Mem/U1107  ( .IN0(\Inst_Mem/inst_mem_reg[28][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1087 ) );
  MUX \Inst_Mem/U1106  ( .IN0(\Inst_Mem/inst_mem_reg[30][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1086 ) );
  MUX \Inst_Mem/U1105  ( .IN0(\Inst_Mem/n1084 ), .IN1(\Inst_Mem/n1069 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1085 ) );
  MUX \Inst_Mem/U1104  ( .IN0(\Inst_Mem/n1083 ), .IN1(\Inst_Mem/n1076 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1084 ) );
  MUX \Inst_Mem/U1103  ( .IN0(\Inst_Mem/n1082 ), .IN1(\Inst_Mem/n1079 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1083 ) );
  MUX \Inst_Mem/U1102  ( .IN0(\Inst_Mem/n1081 ), .IN1(\Inst_Mem/n1080 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1082 ) );
  MUX \Inst_Mem/U1101  ( .IN0(\Inst_Mem/inst_mem_reg[32][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1081 ) );
  MUX \Inst_Mem/U1100  ( .IN0(\Inst_Mem/inst_mem_reg[34][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1080 ) );
  MUX \Inst_Mem/U1099  ( .IN0(\Inst_Mem/n1078 ), .IN1(\Inst_Mem/n1077 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1079 ) );
  MUX \Inst_Mem/U1098  ( .IN0(\Inst_Mem/inst_mem_reg[36][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1078 ) );
  MUX \Inst_Mem/U1097  ( .IN0(\Inst_Mem/inst_mem_reg[38][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1077 ) );
  MUX \Inst_Mem/U1096  ( .IN0(\Inst_Mem/n1075 ), .IN1(\Inst_Mem/n1072 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1076 ) );
  MUX \Inst_Mem/U1095  ( .IN0(\Inst_Mem/n1074 ), .IN1(\Inst_Mem/n1073 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1075 ) );
  MUX \Inst_Mem/U1094  ( .IN0(\Inst_Mem/inst_mem_reg[40][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1074 ) );
  MUX \Inst_Mem/U1093  ( .IN0(\Inst_Mem/inst_mem_reg[42][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1073 ) );
  MUX \Inst_Mem/U1092  ( .IN0(\Inst_Mem/n1071 ), .IN1(\Inst_Mem/n1070 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1072 ) );
  MUX \Inst_Mem/U1091  ( .IN0(\Inst_Mem/inst_mem_reg[44][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1071 ) );
  MUX \Inst_Mem/U1090  ( .IN0(\Inst_Mem/inst_mem_reg[46][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1070 ) );
  MUX \Inst_Mem/U1089  ( .IN0(\Inst_Mem/n1068 ), .IN1(\Inst_Mem/n1061 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1069 ) );
  MUX \Inst_Mem/U1088  ( .IN0(\Inst_Mem/n1067 ), .IN1(\Inst_Mem/n1064 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1068 ) );
  MUX \Inst_Mem/U1087  ( .IN0(\Inst_Mem/n1066 ), .IN1(\Inst_Mem/n1065 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1067 ) );
  MUX \Inst_Mem/U1086  ( .IN0(\Inst_Mem/inst_mem_reg[48][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1066 ) );
  MUX \Inst_Mem/U1085  ( .IN0(\Inst_Mem/inst_mem_reg[50][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1065 ) );
  MUX \Inst_Mem/U1084  ( .IN0(\Inst_Mem/n1063 ), .IN1(\Inst_Mem/n1062 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1064 ) );
  MUX \Inst_Mem/U1083  ( .IN0(\Inst_Mem/inst_mem_reg[52][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1063 ) );
  MUX \Inst_Mem/U1082  ( .IN0(\Inst_Mem/inst_mem_reg[54][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1062 ) );
  MUX \Inst_Mem/U1081  ( .IN0(\Inst_Mem/n1060 ), .IN1(\Inst_Mem/n1057 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1061 ) );
  MUX \Inst_Mem/U1080  ( .IN0(\Inst_Mem/n1059 ), .IN1(\Inst_Mem/n1058 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1060 ) );
  MUX \Inst_Mem/U1079  ( .IN0(\Inst_Mem/inst_mem_reg[56][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1059 ) );
  MUX \Inst_Mem/U1078  ( .IN0(\Inst_Mem/inst_mem_reg[58][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1058 ) );
  MUX \Inst_Mem/U1077  ( .IN0(\Inst_Mem/n1056 ), .IN1(\Inst_Mem/n1055 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1057 ) );
  MUX \Inst_Mem/U1076  ( .IN0(\Inst_Mem/inst_mem_reg[60][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1056 ) );
  MUX \Inst_Mem/U1075  ( .IN0(\Inst_Mem/inst_mem_reg[62][17] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][17] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1055 ) );
  MUX \Inst_Mem/U1074  ( .IN0(\Inst_Mem/n1054 ), .IN1(\Inst_Mem/n1023 ), .SEL(
        pc_current[7]), .F(opcode[16]) );
  MUX \Inst_Mem/U1073  ( .IN0(\Inst_Mem/n1053 ), .IN1(\Inst_Mem/n1038 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1054 ) );
  MUX \Inst_Mem/U1072  ( .IN0(\Inst_Mem/n1052 ), .IN1(\Inst_Mem/n1045 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1053 ) );
  MUX \Inst_Mem/U1071  ( .IN0(\Inst_Mem/n1051 ), .IN1(\Inst_Mem/n1048 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1052 ) );
  MUX \Inst_Mem/U1070  ( .IN0(\Inst_Mem/n1050 ), .IN1(\Inst_Mem/n1049 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1051 ) );
  MUX \Inst_Mem/U1069  ( .IN0(\Inst_Mem/inst_mem_reg[0][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1050 ) );
  MUX \Inst_Mem/U1068  ( .IN0(\Inst_Mem/inst_mem_reg[2][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1049 ) );
  MUX \Inst_Mem/U1067  ( .IN0(\Inst_Mem/n1047 ), .IN1(\Inst_Mem/n1046 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1048 ) );
  MUX \Inst_Mem/U1066  ( .IN0(\Inst_Mem/inst_mem_reg[4][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1047 ) );
  MUX \Inst_Mem/U1065  ( .IN0(\Inst_Mem/inst_mem_reg[6][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1046 ) );
  MUX \Inst_Mem/U1064  ( .IN0(\Inst_Mem/n1044 ), .IN1(\Inst_Mem/n1041 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1045 ) );
  MUX \Inst_Mem/U1063  ( .IN0(\Inst_Mem/n1043 ), .IN1(\Inst_Mem/n1042 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1044 ) );
  MUX \Inst_Mem/U1062  ( .IN0(\Inst_Mem/inst_mem_reg[8][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1043 ) );
  MUX \Inst_Mem/U1061  ( .IN0(\Inst_Mem/inst_mem_reg[10][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1042 ) );
  MUX \Inst_Mem/U1060  ( .IN0(\Inst_Mem/n1040 ), .IN1(\Inst_Mem/n1039 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1041 ) );
  MUX \Inst_Mem/U1059  ( .IN0(\Inst_Mem/inst_mem_reg[12][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1040 ) );
  MUX \Inst_Mem/U1058  ( .IN0(\Inst_Mem/inst_mem_reg[14][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1039 ) );
  MUX \Inst_Mem/U1057  ( .IN0(\Inst_Mem/n1037 ), .IN1(\Inst_Mem/n1030 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1038 ) );
  MUX \Inst_Mem/U1056  ( .IN0(\Inst_Mem/n1036 ), .IN1(\Inst_Mem/n1033 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1037 ) );
  MUX \Inst_Mem/U1055  ( .IN0(\Inst_Mem/n1035 ), .IN1(\Inst_Mem/n1034 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1036 ) );
  MUX \Inst_Mem/U1054  ( .IN0(\Inst_Mem/inst_mem_reg[16][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1035 ) );
  MUX \Inst_Mem/U1053  ( .IN0(\Inst_Mem/inst_mem_reg[18][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1034 ) );
  MUX \Inst_Mem/U1052  ( .IN0(\Inst_Mem/n1032 ), .IN1(\Inst_Mem/n1031 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1033 ) );
  MUX \Inst_Mem/U1051  ( .IN0(\Inst_Mem/inst_mem_reg[20][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1032 ) );
  MUX \Inst_Mem/U1050  ( .IN0(\Inst_Mem/inst_mem_reg[22][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1031 ) );
  MUX \Inst_Mem/U1049  ( .IN0(\Inst_Mem/n1029 ), .IN1(\Inst_Mem/n1026 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1030 ) );
  MUX \Inst_Mem/U1048  ( .IN0(\Inst_Mem/n1028 ), .IN1(\Inst_Mem/n1027 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1029 ) );
  MUX \Inst_Mem/U1047  ( .IN0(\Inst_Mem/inst_mem_reg[24][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1028 ) );
  MUX \Inst_Mem/U1046  ( .IN0(\Inst_Mem/inst_mem_reg[26][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1027 ) );
  MUX \Inst_Mem/U1045  ( .IN0(\Inst_Mem/n1025 ), .IN1(\Inst_Mem/n1024 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1026 ) );
  MUX \Inst_Mem/U1044  ( .IN0(\Inst_Mem/inst_mem_reg[28][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1025 ) );
  MUX \Inst_Mem/U1043  ( .IN0(\Inst_Mem/inst_mem_reg[30][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1024 ) );
  MUX \Inst_Mem/U1042  ( .IN0(\Inst_Mem/n1022 ), .IN1(\Inst_Mem/n1007 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n1023 ) );
  MUX \Inst_Mem/U1041  ( .IN0(\Inst_Mem/n1021 ), .IN1(\Inst_Mem/n1014 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1022 ) );
  MUX \Inst_Mem/U1040  ( .IN0(\Inst_Mem/n1020 ), .IN1(\Inst_Mem/n1017 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1021 ) );
  MUX \Inst_Mem/U1039  ( .IN0(\Inst_Mem/n1019 ), .IN1(\Inst_Mem/n1018 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1020 ) );
  MUX \Inst_Mem/U1038  ( .IN0(\Inst_Mem/inst_mem_reg[32][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1019 ) );
  MUX \Inst_Mem/U1037  ( .IN0(\Inst_Mem/inst_mem_reg[34][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1018 ) );
  MUX \Inst_Mem/U1036  ( .IN0(\Inst_Mem/n1016 ), .IN1(\Inst_Mem/n1015 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1017 ) );
  MUX \Inst_Mem/U1035  ( .IN0(\Inst_Mem/inst_mem_reg[36][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1016 ) );
  MUX \Inst_Mem/U1034  ( .IN0(\Inst_Mem/inst_mem_reg[38][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1015 ) );
  MUX \Inst_Mem/U1033  ( .IN0(\Inst_Mem/n1013 ), .IN1(\Inst_Mem/n1010 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1014 ) );
  MUX \Inst_Mem/U1032  ( .IN0(\Inst_Mem/n1012 ), .IN1(\Inst_Mem/n1011 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1013 ) );
  MUX \Inst_Mem/U1031  ( .IN0(\Inst_Mem/inst_mem_reg[40][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1012 ) );
  MUX \Inst_Mem/U1030  ( .IN0(\Inst_Mem/inst_mem_reg[42][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1011 ) );
  MUX \Inst_Mem/U1029  ( .IN0(\Inst_Mem/n1009 ), .IN1(\Inst_Mem/n1008 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1010 ) );
  MUX \Inst_Mem/U1028  ( .IN0(\Inst_Mem/inst_mem_reg[44][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1009 ) );
  MUX \Inst_Mem/U1027  ( .IN0(\Inst_Mem/inst_mem_reg[46][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1008 ) );
  MUX \Inst_Mem/U1026  ( .IN0(\Inst_Mem/n1006 ), .IN1(\Inst_Mem/n999 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n1007 ) );
  MUX \Inst_Mem/U1025  ( .IN0(\Inst_Mem/n1005 ), .IN1(\Inst_Mem/n1002 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n1006 ) );
  MUX \Inst_Mem/U1024  ( .IN0(\Inst_Mem/n1004 ), .IN1(\Inst_Mem/n1003 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1005 ) );
  MUX \Inst_Mem/U1023  ( .IN0(\Inst_Mem/inst_mem_reg[48][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1004 ) );
  MUX \Inst_Mem/U1022  ( .IN0(\Inst_Mem/inst_mem_reg[50][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1003 ) );
  MUX \Inst_Mem/U1021  ( .IN0(\Inst_Mem/n1001 ), .IN1(\Inst_Mem/n1000 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n1002 ) );
  MUX \Inst_Mem/U1020  ( .IN0(\Inst_Mem/inst_mem_reg[52][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1001 ) );
  MUX \Inst_Mem/U1019  ( .IN0(\Inst_Mem/inst_mem_reg[54][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n1000 ) );
  MUX \Inst_Mem/U1018  ( .IN0(\Inst_Mem/n998 ), .IN1(\Inst_Mem/n995 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n999 ) );
  MUX \Inst_Mem/U1017  ( .IN0(\Inst_Mem/n997 ), .IN1(\Inst_Mem/n996 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n998 ) );
  MUX \Inst_Mem/U1016  ( .IN0(\Inst_Mem/inst_mem_reg[56][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n997 ) );
  MUX \Inst_Mem/U1015  ( .IN0(\Inst_Mem/inst_mem_reg[58][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n996 ) );
  MUX \Inst_Mem/U1014  ( .IN0(\Inst_Mem/n994 ), .IN1(\Inst_Mem/n993 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n995 ) );
  MUX \Inst_Mem/U1013  ( .IN0(\Inst_Mem/inst_mem_reg[60][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n994 ) );
  MUX \Inst_Mem/U1012  ( .IN0(\Inst_Mem/inst_mem_reg[62][16] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][16] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n993 ) );
  MUX \Inst_Mem/U1011  ( .IN0(\Inst_Mem/n992 ), .IN1(\Inst_Mem/n961 ), .SEL(
        pc_current[7]), .F(imm[15]) );
  MUX \Inst_Mem/U1010  ( .IN0(\Inst_Mem/n991 ), .IN1(\Inst_Mem/n976 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n992 ) );
  MUX \Inst_Mem/U1009  ( .IN0(\Inst_Mem/n990 ), .IN1(\Inst_Mem/n983 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n991 ) );
  MUX \Inst_Mem/U1008  ( .IN0(\Inst_Mem/n989 ), .IN1(\Inst_Mem/n986 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n990 ) );
  MUX \Inst_Mem/U1007  ( .IN0(\Inst_Mem/n988 ), .IN1(\Inst_Mem/n987 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n989 ) );
  MUX \Inst_Mem/U1006  ( .IN0(\Inst_Mem/inst_mem_reg[0][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n988 ) );
  MUX \Inst_Mem/U1005  ( .IN0(\Inst_Mem/inst_mem_reg[2][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n987 ) );
  MUX \Inst_Mem/U1004  ( .IN0(\Inst_Mem/n985 ), .IN1(\Inst_Mem/n984 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n986 ) );
  MUX \Inst_Mem/U1003  ( .IN0(\Inst_Mem/inst_mem_reg[4][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n985 ) );
  MUX \Inst_Mem/U1002  ( .IN0(\Inst_Mem/inst_mem_reg[6][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n984 ) );
  MUX \Inst_Mem/U1001  ( .IN0(\Inst_Mem/n982 ), .IN1(\Inst_Mem/n979 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n983 ) );
  MUX \Inst_Mem/U1000  ( .IN0(\Inst_Mem/n981 ), .IN1(\Inst_Mem/n980 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n982 ) );
  MUX \Inst_Mem/U999  ( .IN0(\Inst_Mem/inst_mem_reg[8][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n981 ) );
  MUX \Inst_Mem/U998  ( .IN0(\Inst_Mem/inst_mem_reg[10][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n980 ) );
  MUX \Inst_Mem/U997  ( .IN0(\Inst_Mem/n978 ), .IN1(\Inst_Mem/n977 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n979 ) );
  MUX \Inst_Mem/U996  ( .IN0(\Inst_Mem/inst_mem_reg[12][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n978 ) );
  MUX \Inst_Mem/U995  ( .IN0(\Inst_Mem/inst_mem_reg[14][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n977 ) );
  MUX \Inst_Mem/U994  ( .IN0(\Inst_Mem/n975 ), .IN1(\Inst_Mem/n968 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n976 ) );
  MUX \Inst_Mem/U993  ( .IN0(\Inst_Mem/n974 ), .IN1(\Inst_Mem/n971 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n975 ) );
  MUX \Inst_Mem/U992  ( .IN0(\Inst_Mem/n973 ), .IN1(\Inst_Mem/n972 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n974 ) );
  MUX \Inst_Mem/U991  ( .IN0(\Inst_Mem/inst_mem_reg[16][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n973 ) );
  MUX \Inst_Mem/U990  ( .IN0(\Inst_Mem/inst_mem_reg[18][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n972 ) );
  MUX \Inst_Mem/U989  ( .IN0(\Inst_Mem/n970 ), .IN1(\Inst_Mem/n969 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n971 ) );
  MUX \Inst_Mem/U988  ( .IN0(\Inst_Mem/inst_mem_reg[20][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n970 ) );
  MUX \Inst_Mem/U987  ( .IN0(\Inst_Mem/inst_mem_reg[22][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n969 ) );
  MUX \Inst_Mem/U986  ( .IN0(\Inst_Mem/n967 ), .IN1(\Inst_Mem/n964 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n968 ) );
  MUX \Inst_Mem/U985  ( .IN0(\Inst_Mem/n966 ), .IN1(\Inst_Mem/n965 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n967 ) );
  MUX \Inst_Mem/U984  ( .IN0(\Inst_Mem/inst_mem_reg[24][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n966 ) );
  MUX \Inst_Mem/U983  ( .IN0(\Inst_Mem/inst_mem_reg[26][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n965 ) );
  MUX \Inst_Mem/U982  ( .IN0(\Inst_Mem/n963 ), .IN1(\Inst_Mem/n962 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n964 ) );
  MUX \Inst_Mem/U981  ( .IN0(\Inst_Mem/inst_mem_reg[28][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n963 ) );
  MUX \Inst_Mem/U980  ( .IN0(\Inst_Mem/inst_mem_reg[30][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n962 ) );
  MUX \Inst_Mem/U979  ( .IN0(\Inst_Mem/n960 ), .IN1(\Inst_Mem/n945 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n961 ) );
  MUX \Inst_Mem/U978  ( .IN0(\Inst_Mem/n959 ), .IN1(\Inst_Mem/n952 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n960 ) );
  MUX \Inst_Mem/U977  ( .IN0(\Inst_Mem/n958 ), .IN1(\Inst_Mem/n955 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n959 ) );
  MUX \Inst_Mem/U976  ( .IN0(\Inst_Mem/n957 ), .IN1(\Inst_Mem/n956 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n958 ) );
  MUX \Inst_Mem/U975  ( .IN0(\Inst_Mem/inst_mem_reg[32][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n957 ) );
  MUX \Inst_Mem/U974  ( .IN0(\Inst_Mem/inst_mem_reg[34][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n956 ) );
  MUX \Inst_Mem/U973  ( .IN0(\Inst_Mem/n954 ), .IN1(\Inst_Mem/n953 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n955 ) );
  MUX \Inst_Mem/U972  ( .IN0(\Inst_Mem/inst_mem_reg[36][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n954 ) );
  MUX \Inst_Mem/U971  ( .IN0(\Inst_Mem/inst_mem_reg[38][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n953 ) );
  MUX \Inst_Mem/U970  ( .IN0(\Inst_Mem/n951 ), .IN1(\Inst_Mem/n948 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n952 ) );
  MUX \Inst_Mem/U969  ( .IN0(\Inst_Mem/n950 ), .IN1(\Inst_Mem/n949 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n951 ) );
  MUX \Inst_Mem/U968  ( .IN0(\Inst_Mem/inst_mem_reg[40][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n950 ) );
  MUX \Inst_Mem/U967  ( .IN0(\Inst_Mem/inst_mem_reg[42][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n949 ) );
  MUX \Inst_Mem/U966  ( .IN0(\Inst_Mem/n947 ), .IN1(\Inst_Mem/n946 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n948 ) );
  MUX \Inst_Mem/U965  ( .IN0(\Inst_Mem/inst_mem_reg[44][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n947 ) );
  MUX \Inst_Mem/U964  ( .IN0(\Inst_Mem/inst_mem_reg[46][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n946 ) );
  MUX \Inst_Mem/U963  ( .IN0(\Inst_Mem/n944 ), .IN1(\Inst_Mem/n937 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n945 ) );
  MUX \Inst_Mem/U962  ( .IN0(\Inst_Mem/n943 ), .IN1(\Inst_Mem/n940 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n944 ) );
  MUX \Inst_Mem/U961  ( .IN0(\Inst_Mem/n942 ), .IN1(\Inst_Mem/n941 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n943 ) );
  MUX \Inst_Mem/U960  ( .IN0(\Inst_Mem/inst_mem_reg[48][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n942 ) );
  MUX \Inst_Mem/U959  ( .IN0(\Inst_Mem/inst_mem_reg[50][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n941 ) );
  MUX \Inst_Mem/U958  ( .IN0(\Inst_Mem/n939 ), .IN1(\Inst_Mem/n938 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n940 ) );
  MUX \Inst_Mem/U957  ( .IN0(\Inst_Mem/inst_mem_reg[52][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n939 ) );
  MUX \Inst_Mem/U956  ( .IN0(\Inst_Mem/inst_mem_reg[54][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n938 ) );
  MUX \Inst_Mem/U955  ( .IN0(\Inst_Mem/n936 ), .IN1(\Inst_Mem/n933 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n937 ) );
  MUX \Inst_Mem/U954  ( .IN0(\Inst_Mem/n935 ), .IN1(\Inst_Mem/n934 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n936 ) );
  MUX \Inst_Mem/U953  ( .IN0(\Inst_Mem/inst_mem_reg[56][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n935 ) );
  MUX \Inst_Mem/U952  ( .IN0(\Inst_Mem/inst_mem_reg[58][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n934 ) );
  MUX \Inst_Mem/U951  ( .IN0(\Inst_Mem/n932 ), .IN1(\Inst_Mem/n931 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n933 ) );
  MUX \Inst_Mem/U950  ( .IN0(\Inst_Mem/inst_mem_reg[60][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n932 ) );
  MUX \Inst_Mem/U949  ( .IN0(\Inst_Mem/inst_mem_reg[62][15] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][15] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n931 ) );
  MUX \Inst_Mem/U948  ( .IN0(\Inst_Mem/n930 ), .IN1(\Inst_Mem/n899 ), .SEL(
        pc_current[7]), .F(imm[14]) );
  MUX \Inst_Mem/U947  ( .IN0(\Inst_Mem/n929 ), .IN1(\Inst_Mem/n914 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n930 ) );
  MUX \Inst_Mem/U946  ( .IN0(\Inst_Mem/n928 ), .IN1(\Inst_Mem/n921 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n929 ) );
  MUX \Inst_Mem/U945  ( .IN0(\Inst_Mem/n927 ), .IN1(\Inst_Mem/n924 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n928 ) );
  MUX \Inst_Mem/U944  ( .IN0(\Inst_Mem/n926 ), .IN1(\Inst_Mem/n925 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n927 ) );
  MUX \Inst_Mem/U943  ( .IN0(\Inst_Mem/inst_mem_reg[0][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n926 ) );
  MUX \Inst_Mem/U942  ( .IN0(\Inst_Mem/inst_mem_reg[2][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n925 ) );
  MUX \Inst_Mem/U941  ( .IN0(\Inst_Mem/n923 ), .IN1(\Inst_Mem/n922 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n924 ) );
  MUX \Inst_Mem/U940  ( .IN0(\Inst_Mem/inst_mem_reg[4][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n923 ) );
  MUX \Inst_Mem/U939  ( .IN0(\Inst_Mem/inst_mem_reg[6][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n922 ) );
  MUX \Inst_Mem/U938  ( .IN0(\Inst_Mem/n920 ), .IN1(\Inst_Mem/n917 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n921 ) );
  MUX \Inst_Mem/U937  ( .IN0(\Inst_Mem/n919 ), .IN1(\Inst_Mem/n918 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n920 ) );
  MUX \Inst_Mem/U936  ( .IN0(\Inst_Mem/inst_mem_reg[8][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n919 ) );
  MUX \Inst_Mem/U935  ( .IN0(\Inst_Mem/inst_mem_reg[10][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n918 ) );
  MUX \Inst_Mem/U934  ( .IN0(\Inst_Mem/n916 ), .IN1(\Inst_Mem/n915 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n917 ) );
  MUX \Inst_Mem/U933  ( .IN0(\Inst_Mem/inst_mem_reg[12][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n916 ) );
  MUX \Inst_Mem/U932  ( .IN0(\Inst_Mem/inst_mem_reg[14][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n915 ) );
  MUX \Inst_Mem/U931  ( .IN0(\Inst_Mem/n913 ), .IN1(\Inst_Mem/n906 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n914 ) );
  MUX \Inst_Mem/U930  ( .IN0(\Inst_Mem/n912 ), .IN1(\Inst_Mem/n909 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n913 ) );
  MUX \Inst_Mem/U929  ( .IN0(\Inst_Mem/n911 ), .IN1(\Inst_Mem/n910 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n912 ) );
  MUX \Inst_Mem/U928  ( .IN0(\Inst_Mem/inst_mem_reg[16][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n911 ) );
  MUX \Inst_Mem/U927  ( .IN0(\Inst_Mem/inst_mem_reg[18][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n910 ) );
  MUX \Inst_Mem/U926  ( .IN0(\Inst_Mem/n908 ), .IN1(\Inst_Mem/n907 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n909 ) );
  MUX \Inst_Mem/U925  ( .IN0(\Inst_Mem/inst_mem_reg[20][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n908 ) );
  MUX \Inst_Mem/U924  ( .IN0(\Inst_Mem/inst_mem_reg[22][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n907 ) );
  MUX \Inst_Mem/U923  ( .IN0(\Inst_Mem/n905 ), .IN1(\Inst_Mem/n902 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n906 ) );
  MUX \Inst_Mem/U922  ( .IN0(\Inst_Mem/n904 ), .IN1(\Inst_Mem/n903 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n905 ) );
  MUX \Inst_Mem/U921  ( .IN0(\Inst_Mem/inst_mem_reg[24][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n904 ) );
  MUX \Inst_Mem/U920  ( .IN0(\Inst_Mem/inst_mem_reg[26][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n903 ) );
  MUX \Inst_Mem/U919  ( .IN0(\Inst_Mem/n901 ), .IN1(\Inst_Mem/n900 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n902 ) );
  MUX \Inst_Mem/U918  ( .IN0(\Inst_Mem/inst_mem_reg[28][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n901 ) );
  MUX \Inst_Mem/U917  ( .IN0(\Inst_Mem/inst_mem_reg[30][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n900 ) );
  MUX \Inst_Mem/U916  ( .IN0(\Inst_Mem/n898 ), .IN1(\Inst_Mem/n883 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n899 ) );
  MUX \Inst_Mem/U915  ( .IN0(\Inst_Mem/n897 ), .IN1(\Inst_Mem/n890 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n898 ) );
  MUX \Inst_Mem/U914  ( .IN0(\Inst_Mem/n896 ), .IN1(\Inst_Mem/n893 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n897 ) );
  MUX \Inst_Mem/U913  ( .IN0(\Inst_Mem/n895 ), .IN1(\Inst_Mem/n894 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n896 ) );
  MUX \Inst_Mem/U912  ( .IN0(\Inst_Mem/inst_mem_reg[32][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n895 ) );
  MUX \Inst_Mem/U911  ( .IN0(\Inst_Mem/inst_mem_reg[34][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n894 ) );
  MUX \Inst_Mem/U910  ( .IN0(\Inst_Mem/n892 ), .IN1(\Inst_Mem/n891 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n893 ) );
  MUX \Inst_Mem/U909  ( .IN0(\Inst_Mem/inst_mem_reg[36][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n892 ) );
  MUX \Inst_Mem/U908  ( .IN0(\Inst_Mem/inst_mem_reg[38][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n891 ) );
  MUX \Inst_Mem/U907  ( .IN0(\Inst_Mem/n889 ), .IN1(\Inst_Mem/n886 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n890 ) );
  MUX \Inst_Mem/U906  ( .IN0(\Inst_Mem/n888 ), .IN1(\Inst_Mem/n887 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n889 ) );
  MUX \Inst_Mem/U905  ( .IN0(\Inst_Mem/inst_mem_reg[40][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n888 ) );
  MUX \Inst_Mem/U904  ( .IN0(\Inst_Mem/inst_mem_reg[42][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n887 ) );
  MUX \Inst_Mem/U903  ( .IN0(\Inst_Mem/n885 ), .IN1(\Inst_Mem/n884 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n886 ) );
  MUX \Inst_Mem/U902  ( .IN0(\Inst_Mem/inst_mem_reg[44][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n885 ) );
  MUX \Inst_Mem/U901  ( .IN0(\Inst_Mem/inst_mem_reg[46][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n884 ) );
  MUX \Inst_Mem/U900  ( .IN0(\Inst_Mem/n882 ), .IN1(\Inst_Mem/n875 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n883 ) );
  MUX \Inst_Mem/U899  ( .IN0(\Inst_Mem/n881 ), .IN1(\Inst_Mem/n878 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n882 ) );
  MUX \Inst_Mem/U898  ( .IN0(\Inst_Mem/n880 ), .IN1(\Inst_Mem/n879 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n881 ) );
  MUX \Inst_Mem/U897  ( .IN0(\Inst_Mem/inst_mem_reg[48][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n880 ) );
  MUX \Inst_Mem/U896  ( .IN0(\Inst_Mem/inst_mem_reg[50][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n879 ) );
  MUX \Inst_Mem/U895  ( .IN0(\Inst_Mem/n877 ), .IN1(\Inst_Mem/n876 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n878 ) );
  MUX \Inst_Mem/U894  ( .IN0(\Inst_Mem/inst_mem_reg[52][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n877 ) );
  MUX \Inst_Mem/U893  ( .IN0(\Inst_Mem/inst_mem_reg[54][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n876 ) );
  MUX \Inst_Mem/U892  ( .IN0(\Inst_Mem/n874 ), .IN1(\Inst_Mem/n871 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n875 ) );
  MUX \Inst_Mem/U891  ( .IN0(\Inst_Mem/n873 ), .IN1(\Inst_Mem/n872 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n874 ) );
  MUX \Inst_Mem/U890  ( .IN0(\Inst_Mem/inst_mem_reg[56][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n873 ) );
  MUX \Inst_Mem/U889  ( .IN0(\Inst_Mem/inst_mem_reg[58][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n872 ) );
  MUX \Inst_Mem/U888  ( .IN0(\Inst_Mem/n870 ), .IN1(\Inst_Mem/n869 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n871 ) );
  MUX \Inst_Mem/U887  ( .IN0(\Inst_Mem/inst_mem_reg[60][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n870 ) );
  MUX \Inst_Mem/U886  ( .IN0(\Inst_Mem/inst_mem_reg[62][14] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][14] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n869 ) );
  MUX \Inst_Mem/U885  ( .IN0(\Inst_Mem/n868 ), .IN1(\Inst_Mem/n837 ), .SEL(
        pc_current[7]), .F(imm[13]) );
  MUX \Inst_Mem/U884  ( .IN0(\Inst_Mem/n867 ), .IN1(\Inst_Mem/n852 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n868 ) );
  MUX \Inst_Mem/U883  ( .IN0(\Inst_Mem/n866 ), .IN1(\Inst_Mem/n859 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n867 ) );
  MUX \Inst_Mem/U882  ( .IN0(\Inst_Mem/n865 ), .IN1(\Inst_Mem/n862 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n866 ) );
  MUX \Inst_Mem/U881  ( .IN0(\Inst_Mem/n864 ), .IN1(\Inst_Mem/n863 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n865 ) );
  MUX \Inst_Mem/U880  ( .IN0(\Inst_Mem/inst_mem_reg[0][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n864 ) );
  MUX \Inst_Mem/U879  ( .IN0(\Inst_Mem/inst_mem_reg[2][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n863 ) );
  MUX \Inst_Mem/U878  ( .IN0(\Inst_Mem/n861 ), .IN1(\Inst_Mem/n860 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n862 ) );
  MUX \Inst_Mem/U877  ( .IN0(\Inst_Mem/inst_mem_reg[4][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n861 ) );
  MUX \Inst_Mem/U876  ( .IN0(\Inst_Mem/inst_mem_reg[6][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n860 ) );
  MUX \Inst_Mem/U875  ( .IN0(\Inst_Mem/n858 ), .IN1(\Inst_Mem/n855 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n859 ) );
  MUX \Inst_Mem/U874  ( .IN0(\Inst_Mem/n857 ), .IN1(\Inst_Mem/n856 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n858 ) );
  MUX \Inst_Mem/U873  ( .IN0(\Inst_Mem/inst_mem_reg[8][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n857 ) );
  MUX \Inst_Mem/U872  ( .IN0(\Inst_Mem/inst_mem_reg[10][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n856 ) );
  MUX \Inst_Mem/U871  ( .IN0(\Inst_Mem/n854 ), .IN1(\Inst_Mem/n853 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n855 ) );
  MUX \Inst_Mem/U870  ( .IN0(\Inst_Mem/inst_mem_reg[12][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n854 ) );
  MUX \Inst_Mem/U869  ( .IN0(\Inst_Mem/inst_mem_reg[14][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n853 ) );
  MUX \Inst_Mem/U868  ( .IN0(\Inst_Mem/n851 ), .IN1(\Inst_Mem/n844 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n852 ) );
  MUX \Inst_Mem/U867  ( .IN0(\Inst_Mem/n850 ), .IN1(\Inst_Mem/n847 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n851 ) );
  MUX \Inst_Mem/U866  ( .IN0(\Inst_Mem/n849 ), .IN1(\Inst_Mem/n848 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n850 ) );
  MUX \Inst_Mem/U865  ( .IN0(\Inst_Mem/inst_mem_reg[16][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n849 ) );
  MUX \Inst_Mem/U864  ( .IN0(\Inst_Mem/inst_mem_reg[18][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n848 ) );
  MUX \Inst_Mem/U863  ( .IN0(\Inst_Mem/n846 ), .IN1(\Inst_Mem/n845 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n847 ) );
  MUX \Inst_Mem/U862  ( .IN0(\Inst_Mem/inst_mem_reg[20][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n846 ) );
  MUX \Inst_Mem/U861  ( .IN0(\Inst_Mem/inst_mem_reg[22][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n845 ) );
  MUX \Inst_Mem/U860  ( .IN0(\Inst_Mem/n843 ), .IN1(\Inst_Mem/n840 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n844 ) );
  MUX \Inst_Mem/U859  ( .IN0(\Inst_Mem/n842 ), .IN1(\Inst_Mem/n841 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n843 ) );
  MUX \Inst_Mem/U858  ( .IN0(\Inst_Mem/inst_mem_reg[24][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n842 ) );
  MUX \Inst_Mem/U857  ( .IN0(\Inst_Mem/inst_mem_reg[26][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n841 ) );
  MUX \Inst_Mem/U856  ( .IN0(\Inst_Mem/n839 ), .IN1(\Inst_Mem/n838 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n840 ) );
  MUX \Inst_Mem/U855  ( .IN0(\Inst_Mem/inst_mem_reg[28][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n839 ) );
  MUX \Inst_Mem/U854  ( .IN0(\Inst_Mem/inst_mem_reg[30][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n838 ) );
  MUX \Inst_Mem/U853  ( .IN0(\Inst_Mem/n836 ), .IN1(\Inst_Mem/n821 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n837 ) );
  MUX \Inst_Mem/U852  ( .IN0(\Inst_Mem/n835 ), .IN1(\Inst_Mem/n828 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n836 ) );
  MUX \Inst_Mem/U851  ( .IN0(\Inst_Mem/n834 ), .IN1(\Inst_Mem/n831 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n835 ) );
  MUX \Inst_Mem/U850  ( .IN0(\Inst_Mem/n833 ), .IN1(\Inst_Mem/n832 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n834 ) );
  MUX \Inst_Mem/U849  ( .IN0(\Inst_Mem/inst_mem_reg[32][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n833 ) );
  MUX \Inst_Mem/U848  ( .IN0(\Inst_Mem/inst_mem_reg[34][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n832 ) );
  MUX \Inst_Mem/U847  ( .IN0(\Inst_Mem/n830 ), .IN1(\Inst_Mem/n829 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n831 ) );
  MUX \Inst_Mem/U846  ( .IN0(\Inst_Mem/inst_mem_reg[36][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n830 ) );
  MUX \Inst_Mem/U845  ( .IN0(\Inst_Mem/inst_mem_reg[38][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n829 ) );
  MUX \Inst_Mem/U844  ( .IN0(\Inst_Mem/n827 ), .IN1(\Inst_Mem/n824 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n828 ) );
  MUX \Inst_Mem/U843  ( .IN0(\Inst_Mem/n826 ), .IN1(\Inst_Mem/n825 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n827 ) );
  MUX \Inst_Mem/U842  ( .IN0(\Inst_Mem/inst_mem_reg[40][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n826 ) );
  MUX \Inst_Mem/U841  ( .IN0(\Inst_Mem/inst_mem_reg[42][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n825 ) );
  MUX \Inst_Mem/U840  ( .IN0(\Inst_Mem/n823 ), .IN1(\Inst_Mem/n822 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n824 ) );
  MUX \Inst_Mem/U839  ( .IN0(\Inst_Mem/inst_mem_reg[44][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n823 ) );
  MUX \Inst_Mem/U838  ( .IN0(\Inst_Mem/inst_mem_reg[46][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n822 ) );
  MUX \Inst_Mem/U837  ( .IN0(\Inst_Mem/n820 ), .IN1(\Inst_Mem/n813 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n821 ) );
  MUX \Inst_Mem/U836  ( .IN0(\Inst_Mem/n819 ), .IN1(\Inst_Mem/n816 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n820 ) );
  MUX \Inst_Mem/U835  ( .IN0(\Inst_Mem/n818 ), .IN1(\Inst_Mem/n817 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n819 ) );
  MUX \Inst_Mem/U834  ( .IN0(\Inst_Mem/inst_mem_reg[48][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n818 ) );
  MUX \Inst_Mem/U833  ( .IN0(\Inst_Mem/inst_mem_reg[50][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n817 ) );
  MUX \Inst_Mem/U832  ( .IN0(\Inst_Mem/n815 ), .IN1(\Inst_Mem/n814 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n816 ) );
  MUX \Inst_Mem/U831  ( .IN0(\Inst_Mem/inst_mem_reg[52][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n815 ) );
  MUX \Inst_Mem/U830  ( .IN0(\Inst_Mem/inst_mem_reg[54][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n814 ) );
  MUX \Inst_Mem/U829  ( .IN0(\Inst_Mem/n812 ), .IN1(\Inst_Mem/n809 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n813 ) );
  MUX \Inst_Mem/U828  ( .IN0(\Inst_Mem/n811 ), .IN1(\Inst_Mem/n810 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n812 ) );
  MUX \Inst_Mem/U827  ( .IN0(\Inst_Mem/inst_mem_reg[56][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n811 ) );
  MUX \Inst_Mem/U826  ( .IN0(\Inst_Mem/inst_mem_reg[58][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n810 ) );
  MUX \Inst_Mem/U825  ( .IN0(\Inst_Mem/n808 ), .IN1(\Inst_Mem/n807 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n809 ) );
  MUX \Inst_Mem/U824  ( .IN0(\Inst_Mem/inst_mem_reg[60][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n808 ) );
  MUX \Inst_Mem/U823  ( .IN0(\Inst_Mem/inst_mem_reg[62][13] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][13] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n807 ) );
  MUX \Inst_Mem/U822  ( .IN0(\Inst_Mem/n806 ), .IN1(\Inst_Mem/n775 ), .SEL(
        pc_current[7]), .F(imm[12]) );
  MUX \Inst_Mem/U821  ( .IN0(\Inst_Mem/n805 ), .IN1(\Inst_Mem/n790 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n806 ) );
  MUX \Inst_Mem/U820  ( .IN0(\Inst_Mem/n804 ), .IN1(\Inst_Mem/n797 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n805 ) );
  MUX \Inst_Mem/U819  ( .IN0(\Inst_Mem/n803 ), .IN1(\Inst_Mem/n800 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n804 ) );
  MUX \Inst_Mem/U818  ( .IN0(\Inst_Mem/n802 ), .IN1(\Inst_Mem/n801 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n803 ) );
  MUX \Inst_Mem/U817  ( .IN0(\Inst_Mem/inst_mem_reg[0][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n802 ) );
  MUX \Inst_Mem/U816  ( .IN0(\Inst_Mem/inst_mem_reg[2][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n801 ) );
  MUX \Inst_Mem/U815  ( .IN0(\Inst_Mem/n799 ), .IN1(\Inst_Mem/n798 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n800 ) );
  MUX \Inst_Mem/U814  ( .IN0(\Inst_Mem/inst_mem_reg[4][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n799 ) );
  MUX \Inst_Mem/U813  ( .IN0(\Inst_Mem/inst_mem_reg[6][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n798 ) );
  MUX \Inst_Mem/U812  ( .IN0(\Inst_Mem/n796 ), .IN1(\Inst_Mem/n793 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n797 ) );
  MUX \Inst_Mem/U811  ( .IN0(\Inst_Mem/n795 ), .IN1(\Inst_Mem/n794 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n796 ) );
  MUX \Inst_Mem/U810  ( .IN0(\Inst_Mem/inst_mem_reg[8][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n795 ) );
  MUX \Inst_Mem/U809  ( .IN0(\Inst_Mem/inst_mem_reg[10][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n794 ) );
  MUX \Inst_Mem/U808  ( .IN0(\Inst_Mem/n792 ), .IN1(\Inst_Mem/n791 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n793 ) );
  MUX \Inst_Mem/U807  ( .IN0(\Inst_Mem/inst_mem_reg[12][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n792 ) );
  MUX \Inst_Mem/U806  ( .IN0(\Inst_Mem/inst_mem_reg[14][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n791 ) );
  MUX \Inst_Mem/U805  ( .IN0(\Inst_Mem/n789 ), .IN1(\Inst_Mem/n782 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n790 ) );
  MUX \Inst_Mem/U804  ( .IN0(\Inst_Mem/n788 ), .IN1(\Inst_Mem/n785 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n789 ) );
  MUX \Inst_Mem/U803  ( .IN0(\Inst_Mem/n787 ), .IN1(\Inst_Mem/n786 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n788 ) );
  MUX \Inst_Mem/U802  ( .IN0(\Inst_Mem/inst_mem_reg[16][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n787 ) );
  MUX \Inst_Mem/U801  ( .IN0(\Inst_Mem/inst_mem_reg[18][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n786 ) );
  MUX \Inst_Mem/U800  ( .IN0(\Inst_Mem/n784 ), .IN1(\Inst_Mem/n783 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n785 ) );
  MUX \Inst_Mem/U799  ( .IN0(\Inst_Mem/inst_mem_reg[20][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n784 ) );
  MUX \Inst_Mem/U798  ( .IN0(\Inst_Mem/inst_mem_reg[22][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n783 ) );
  MUX \Inst_Mem/U797  ( .IN0(\Inst_Mem/n781 ), .IN1(\Inst_Mem/n778 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n782 ) );
  MUX \Inst_Mem/U796  ( .IN0(\Inst_Mem/n780 ), .IN1(\Inst_Mem/n779 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n781 ) );
  MUX \Inst_Mem/U795  ( .IN0(\Inst_Mem/inst_mem_reg[24][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n780 ) );
  MUX \Inst_Mem/U794  ( .IN0(\Inst_Mem/inst_mem_reg[26][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n779 ) );
  MUX \Inst_Mem/U793  ( .IN0(\Inst_Mem/n777 ), .IN1(\Inst_Mem/n776 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n778 ) );
  MUX \Inst_Mem/U792  ( .IN0(\Inst_Mem/inst_mem_reg[28][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n777 ) );
  MUX \Inst_Mem/U791  ( .IN0(\Inst_Mem/inst_mem_reg[30][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n776 ) );
  MUX \Inst_Mem/U790  ( .IN0(\Inst_Mem/n774 ), .IN1(\Inst_Mem/n759 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n775 ) );
  MUX \Inst_Mem/U789  ( .IN0(\Inst_Mem/n773 ), .IN1(\Inst_Mem/n766 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n774 ) );
  MUX \Inst_Mem/U788  ( .IN0(\Inst_Mem/n772 ), .IN1(\Inst_Mem/n769 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n773 ) );
  MUX \Inst_Mem/U787  ( .IN0(\Inst_Mem/n771 ), .IN1(\Inst_Mem/n770 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n772 ) );
  MUX \Inst_Mem/U786  ( .IN0(\Inst_Mem/inst_mem_reg[32][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n771 ) );
  MUX \Inst_Mem/U785  ( .IN0(\Inst_Mem/inst_mem_reg[34][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n770 ) );
  MUX \Inst_Mem/U784  ( .IN0(\Inst_Mem/n768 ), .IN1(\Inst_Mem/n767 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n769 ) );
  MUX \Inst_Mem/U783  ( .IN0(\Inst_Mem/inst_mem_reg[36][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n768 ) );
  MUX \Inst_Mem/U782  ( .IN0(\Inst_Mem/inst_mem_reg[38][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n767 ) );
  MUX \Inst_Mem/U781  ( .IN0(\Inst_Mem/n765 ), .IN1(\Inst_Mem/n762 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n766 ) );
  MUX \Inst_Mem/U780  ( .IN0(\Inst_Mem/n764 ), .IN1(\Inst_Mem/n763 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n765 ) );
  MUX \Inst_Mem/U779  ( .IN0(\Inst_Mem/inst_mem_reg[40][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n764 ) );
  MUX \Inst_Mem/U778  ( .IN0(\Inst_Mem/inst_mem_reg[42][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n763 ) );
  MUX \Inst_Mem/U777  ( .IN0(\Inst_Mem/n761 ), .IN1(\Inst_Mem/n760 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n762 ) );
  MUX \Inst_Mem/U776  ( .IN0(\Inst_Mem/inst_mem_reg[44][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n761 ) );
  MUX \Inst_Mem/U775  ( .IN0(\Inst_Mem/inst_mem_reg[46][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n760 ) );
  MUX \Inst_Mem/U774  ( .IN0(\Inst_Mem/n758 ), .IN1(\Inst_Mem/n751 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n759 ) );
  MUX \Inst_Mem/U773  ( .IN0(\Inst_Mem/n757 ), .IN1(\Inst_Mem/n754 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n758 ) );
  MUX \Inst_Mem/U772  ( .IN0(\Inst_Mem/n756 ), .IN1(\Inst_Mem/n755 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n757 ) );
  MUX \Inst_Mem/U771  ( .IN0(\Inst_Mem/inst_mem_reg[48][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n756 ) );
  MUX \Inst_Mem/U770  ( .IN0(\Inst_Mem/inst_mem_reg[50][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n755 ) );
  MUX \Inst_Mem/U769  ( .IN0(\Inst_Mem/n753 ), .IN1(\Inst_Mem/n752 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n754 ) );
  MUX \Inst_Mem/U768  ( .IN0(\Inst_Mem/inst_mem_reg[52][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n753 ) );
  MUX \Inst_Mem/U767  ( .IN0(\Inst_Mem/inst_mem_reg[54][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n752 ) );
  MUX \Inst_Mem/U766  ( .IN0(\Inst_Mem/n750 ), .IN1(\Inst_Mem/n747 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n751 ) );
  MUX \Inst_Mem/U765  ( .IN0(\Inst_Mem/n749 ), .IN1(\Inst_Mem/n748 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n750 ) );
  MUX \Inst_Mem/U764  ( .IN0(\Inst_Mem/inst_mem_reg[56][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n749 ) );
  MUX \Inst_Mem/U763  ( .IN0(\Inst_Mem/inst_mem_reg[58][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n748 ) );
  MUX \Inst_Mem/U762  ( .IN0(\Inst_Mem/n746 ), .IN1(\Inst_Mem/n745 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n747 ) );
  MUX \Inst_Mem/U761  ( .IN0(\Inst_Mem/inst_mem_reg[60][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n746 ) );
  MUX \Inst_Mem/U760  ( .IN0(\Inst_Mem/inst_mem_reg[62][12] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][12] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n745 ) );
  MUX \Inst_Mem/U759  ( .IN0(\Inst_Mem/n744 ), .IN1(\Inst_Mem/n713 ), .SEL(
        pc_current[7]), .F(imm[11]) );
  MUX \Inst_Mem/U758  ( .IN0(\Inst_Mem/n743 ), .IN1(\Inst_Mem/n728 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n744 ) );
  MUX \Inst_Mem/U757  ( .IN0(\Inst_Mem/n742 ), .IN1(\Inst_Mem/n735 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n743 ) );
  MUX \Inst_Mem/U756  ( .IN0(\Inst_Mem/n741 ), .IN1(\Inst_Mem/n738 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n742 ) );
  MUX \Inst_Mem/U755  ( .IN0(\Inst_Mem/n740 ), .IN1(\Inst_Mem/n739 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n741 ) );
  MUX \Inst_Mem/U754  ( .IN0(\Inst_Mem/inst_mem_reg[0][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n740 ) );
  MUX \Inst_Mem/U753  ( .IN0(\Inst_Mem/inst_mem_reg[2][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n739 ) );
  MUX \Inst_Mem/U752  ( .IN0(\Inst_Mem/n737 ), .IN1(\Inst_Mem/n736 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n738 ) );
  MUX \Inst_Mem/U751  ( .IN0(\Inst_Mem/inst_mem_reg[4][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n737 ) );
  MUX \Inst_Mem/U750  ( .IN0(\Inst_Mem/inst_mem_reg[6][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n736 ) );
  MUX \Inst_Mem/U749  ( .IN0(\Inst_Mem/n734 ), .IN1(\Inst_Mem/n731 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n735 ) );
  MUX \Inst_Mem/U748  ( .IN0(\Inst_Mem/n733 ), .IN1(\Inst_Mem/n732 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n734 ) );
  MUX \Inst_Mem/U747  ( .IN0(\Inst_Mem/inst_mem_reg[8][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n733 ) );
  MUX \Inst_Mem/U746  ( .IN0(\Inst_Mem/inst_mem_reg[10][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n732 ) );
  MUX \Inst_Mem/U745  ( .IN0(\Inst_Mem/n730 ), .IN1(\Inst_Mem/n729 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n731 ) );
  MUX \Inst_Mem/U744  ( .IN0(\Inst_Mem/inst_mem_reg[12][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n730 ) );
  MUX \Inst_Mem/U743  ( .IN0(\Inst_Mem/inst_mem_reg[14][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n729 ) );
  MUX \Inst_Mem/U742  ( .IN0(\Inst_Mem/n727 ), .IN1(\Inst_Mem/n720 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n728 ) );
  MUX \Inst_Mem/U741  ( .IN0(\Inst_Mem/n726 ), .IN1(\Inst_Mem/n723 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n727 ) );
  MUX \Inst_Mem/U740  ( .IN0(\Inst_Mem/n725 ), .IN1(\Inst_Mem/n724 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n726 ) );
  MUX \Inst_Mem/U739  ( .IN0(\Inst_Mem/inst_mem_reg[16][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n725 ) );
  MUX \Inst_Mem/U738  ( .IN0(\Inst_Mem/inst_mem_reg[18][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n724 ) );
  MUX \Inst_Mem/U737  ( .IN0(\Inst_Mem/n722 ), .IN1(\Inst_Mem/n721 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n723 ) );
  MUX \Inst_Mem/U736  ( .IN0(\Inst_Mem/inst_mem_reg[20][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n722 ) );
  MUX \Inst_Mem/U735  ( .IN0(\Inst_Mem/inst_mem_reg[22][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n721 ) );
  MUX \Inst_Mem/U734  ( .IN0(\Inst_Mem/n719 ), .IN1(\Inst_Mem/n716 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n720 ) );
  MUX \Inst_Mem/U733  ( .IN0(\Inst_Mem/n718 ), .IN1(\Inst_Mem/n717 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n719 ) );
  MUX \Inst_Mem/U732  ( .IN0(\Inst_Mem/inst_mem_reg[24][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n718 ) );
  MUX \Inst_Mem/U731  ( .IN0(\Inst_Mem/inst_mem_reg[26][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n717 ) );
  MUX \Inst_Mem/U730  ( .IN0(\Inst_Mem/n715 ), .IN1(\Inst_Mem/n714 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n716 ) );
  MUX \Inst_Mem/U729  ( .IN0(\Inst_Mem/inst_mem_reg[28][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n715 ) );
  MUX \Inst_Mem/U728  ( .IN0(\Inst_Mem/inst_mem_reg[30][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n714 ) );
  MUX \Inst_Mem/U727  ( .IN0(\Inst_Mem/n712 ), .IN1(\Inst_Mem/n697 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n713 ) );
  MUX \Inst_Mem/U726  ( .IN0(\Inst_Mem/n711 ), .IN1(\Inst_Mem/n704 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n712 ) );
  MUX \Inst_Mem/U725  ( .IN0(\Inst_Mem/n710 ), .IN1(\Inst_Mem/n707 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n711 ) );
  MUX \Inst_Mem/U724  ( .IN0(\Inst_Mem/n709 ), .IN1(\Inst_Mem/n708 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n710 ) );
  MUX \Inst_Mem/U723  ( .IN0(\Inst_Mem/inst_mem_reg[32][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n709 ) );
  MUX \Inst_Mem/U722  ( .IN0(\Inst_Mem/inst_mem_reg[34][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n708 ) );
  MUX \Inst_Mem/U721  ( .IN0(\Inst_Mem/n706 ), .IN1(\Inst_Mem/n705 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n707 ) );
  MUX \Inst_Mem/U720  ( .IN0(\Inst_Mem/inst_mem_reg[36][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n706 ) );
  MUX \Inst_Mem/U719  ( .IN0(\Inst_Mem/inst_mem_reg[38][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n705 ) );
  MUX \Inst_Mem/U718  ( .IN0(\Inst_Mem/n703 ), .IN1(\Inst_Mem/n700 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n704 ) );
  MUX \Inst_Mem/U717  ( .IN0(\Inst_Mem/n702 ), .IN1(\Inst_Mem/n701 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n703 ) );
  MUX \Inst_Mem/U716  ( .IN0(\Inst_Mem/inst_mem_reg[40][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n702 ) );
  MUX \Inst_Mem/U715  ( .IN0(\Inst_Mem/inst_mem_reg[42][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n701 ) );
  MUX \Inst_Mem/U714  ( .IN0(\Inst_Mem/n699 ), .IN1(\Inst_Mem/n698 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n700 ) );
  MUX \Inst_Mem/U713  ( .IN0(\Inst_Mem/inst_mem_reg[44][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n699 ) );
  MUX \Inst_Mem/U712  ( .IN0(\Inst_Mem/inst_mem_reg[46][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n698 ) );
  MUX \Inst_Mem/U711  ( .IN0(\Inst_Mem/n696 ), .IN1(\Inst_Mem/n689 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n697 ) );
  MUX \Inst_Mem/U710  ( .IN0(\Inst_Mem/n695 ), .IN1(\Inst_Mem/n692 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n696 ) );
  MUX \Inst_Mem/U709  ( .IN0(\Inst_Mem/n694 ), .IN1(\Inst_Mem/n693 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n695 ) );
  MUX \Inst_Mem/U708  ( .IN0(\Inst_Mem/inst_mem_reg[48][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n694 ) );
  MUX \Inst_Mem/U707  ( .IN0(\Inst_Mem/inst_mem_reg[50][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n693 ) );
  MUX \Inst_Mem/U706  ( .IN0(\Inst_Mem/n691 ), .IN1(\Inst_Mem/n690 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n692 ) );
  MUX \Inst_Mem/U705  ( .IN0(\Inst_Mem/inst_mem_reg[52][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n691 ) );
  MUX \Inst_Mem/U704  ( .IN0(\Inst_Mem/inst_mem_reg[54][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n690 ) );
  MUX \Inst_Mem/U703  ( .IN0(\Inst_Mem/n688 ), .IN1(\Inst_Mem/n685 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n689 ) );
  MUX \Inst_Mem/U702  ( .IN0(\Inst_Mem/n687 ), .IN1(\Inst_Mem/n686 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n688 ) );
  MUX \Inst_Mem/U701  ( .IN0(\Inst_Mem/inst_mem_reg[56][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n687 ) );
  MUX \Inst_Mem/U700  ( .IN0(\Inst_Mem/inst_mem_reg[58][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n686 ) );
  MUX \Inst_Mem/U699  ( .IN0(\Inst_Mem/n684 ), .IN1(\Inst_Mem/n683 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n685 ) );
  MUX \Inst_Mem/U698  ( .IN0(\Inst_Mem/inst_mem_reg[60][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n684 ) );
  MUX \Inst_Mem/U697  ( .IN0(\Inst_Mem/inst_mem_reg[62][11] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][11] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n683 ) );
  MUX \Inst_Mem/U696  ( .IN0(\Inst_Mem/n682 ), .IN1(\Inst_Mem/n651 ), .SEL(
        pc_current[7]), .F(imm[10]) );
  MUX \Inst_Mem/U695  ( .IN0(\Inst_Mem/n681 ), .IN1(\Inst_Mem/n666 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n682 ) );
  MUX \Inst_Mem/U694  ( .IN0(\Inst_Mem/n680 ), .IN1(\Inst_Mem/n673 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n681 ) );
  MUX \Inst_Mem/U693  ( .IN0(\Inst_Mem/n679 ), .IN1(\Inst_Mem/n676 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n680 ) );
  MUX \Inst_Mem/U692  ( .IN0(\Inst_Mem/n678 ), .IN1(\Inst_Mem/n677 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n679 ) );
  MUX \Inst_Mem/U691  ( .IN0(\Inst_Mem/inst_mem_reg[0][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n678 ) );
  MUX \Inst_Mem/U690  ( .IN0(\Inst_Mem/inst_mem_reg[2][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n677 ) );
  MUX \Inst_Mem/U689  ( .IN0(\Inst_Mem/n675 ), .IN1(\Inst_Mem/n674 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n676 ) );
  MUX \Inst_Mem/U688  ( .IN0(\Inst_Mem/inst_mem_reg[4][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n675 ) );
  MUX \Inst_Mem/U687  ( .IN0(\Inst_Mem/inst_mem_reg[6][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n674 ) );
  MUX \Inst_Mem/U686  ( .IN0(\Inst_Mem/n672 ), .IN1(\Inst_Mem/n669 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n673 ) );
  MUX \Inst_Mem/U685  ( .IN0(\Inst_Mem/n671 ), .IN1(\Inst_Mem/n670 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n672 ) );
  MUX \Inst_Mem/U684  ( .IN0(\Inst_Mem/inst_mem_reg[8][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n671 ) );
  MUX \Inst_Mem/U683  ( .IN0(\Inst_Mem/inst_mem_reg[10][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n670 ) );
  MUX \Inst_Mem/U682  ( .IN0(\Inst_Mem/n668 ), .IN1(\Inst_Mem/n667 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n669 ) );
  MUX \Inst_Mem/U681  ( .IN0(\Inst_Mem/inst_mem_reg[12][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n668 ) );
  MUX \Inst_Mem/U680  ( .IN0(\Inst_Mem/inst_mem_reg[14][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n667 ) );
  MUX \Inst_Mem/U679  ( .IN0(\Inst_Mem/n665 ), .IN1(\Inst_Mem/n658 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n666 ) );
  MUX \Inst_Mem/U678  ( .IN0(\Inst_Mem/n664 ), .IN1(\Inst_Mem/n661 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n665 ) );
  MUX \Inst_Mem/U677  ( .IN0(\Inst_Mem/n663 ), .IN1(\Inst_Mem/n662 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n664 ) );
  MUX \Inst_Mem/U676  ( .IN0(\Inst_Mem/inst_mem_reg[16][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n663 ) );
  MUX \Inst_Mem/U675  ( .IN0(\Inst_Mem/inst_mem_reg[18][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n662 ) );
  MUX \Inst_Mem/U674  ( .IN0(\Inst_Mem/n660 ), .IN1(\Inst_Mem/n659 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n661 ) );
  MUX \Inst_Mem/U673  ( .IN0(\Inst_Mem/inst_mem_reg[20][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n660 ) );
  MUX \Inst_Mem/U672  ( .IN0(\Inst_Mem/inst_mem_reg[22][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n659 ) );
  MUX \Inst_Mem/U671  ( .IN0(\Inst_Mem/n657 ), .IN1(\Inst_Mem/n654 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n658 ) );
  MUX \Inst_Mem/U670  ( .IN0(\Inst_Mem/n656 ), .IN1(\Inst_Mem/n655 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n657 ) );
  MUX \Inst_Mem/U669  ( .IN0(\Inst_Mem/inst_mem_reg[24][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n656 ) );
  MUX \Inst_Mem/U668  ( .IN0(\Inst_Mem/inst_mem_reg[26][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n655 ) );
  MUX \Inst_Mem/U667  ( .IN0(\Inst_Mem/n653 ), .IN1(\Inst_Mem/n652 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n654 ) );
  MUX \Inst_Mem/U666  ( .IN0(\Inst_Mem/inst_mem_reg[28][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n653 ) );
  MUX \Inst_Mem/U665  ( .IN0(\Inst_Mem/inst_mem_reg[30][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n652 ) );
  MUX \Inst_Mem/U664  ( .IN0(\Inst_Mem/n650 ), .IN1(\Inst_Mem/n635 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n651 ) );
  MUX \Inst_Mem/U663  ( .IN0(\Inst_Mem/n649 ), .IN1(\Inst_Mem/n642 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n650 ) );
  MUX \Inst_Mem/U662  ( .IN0(\Inst_Mem/n648 ), .IN1(\Inst_Mem/n645 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n649 ) );
  MUX \Inst_Mem/U661  ( .IN0(\Inst_Mem/n647 ), .IN1(\Inst_Mem/n646 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n648 ) );
  MUX \Inst_Mem/U660  ( .IN0(\Inst_Mem/inst_mem_reg[32][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n647 ) );
  MUX \Inst_Mem/U659  ( .IN0(\Inst_Mem/inst_mem_reg[34][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n646 ) );
  MUX \Inst_Mem/U658  ( .IN0(\Inst_Mem/n644 ), .IN1(\Inst_Mem/n643 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n645 ) );
  MUX \Inst_Mem/U657  ( .IN0(\Inst_Mem/inst_mem_reg[36][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n644 ) );
  MUX \Inst_Mem/U656  ( .IN0(\Inst_Mem/inst_mem_reg[38][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n643 ) );
  MUX \Inst_Mem/U655  ( .IN0(\Inst_Mem/n641 ), .IN1(\Inst_Mem/n638 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n642 ) );
  MUX \Inst_Mem/U654  ( .IN0(\Inst_Mem/n640 ), .IN1(\Inst_Mem/n639 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n641 ) );
  MUX \Inst_Mem/U653  ( .IN0(\Inst_Mem/inst_mem_reg[40][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n640 ) );
  MUX \Inst_Mem/U652  ( .IN0(\Inst_Mem/inst_mem_reg[42][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n639 ) );
  MUX \Inst_Mem/U651  ( .IN0(\Inst_Mem/n637 ), .IN1(\Inst_Mem/n636 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n638 ) );
  MUX \Inst_Mem/U650  ( .IN0(\Inst_Mem/inst_mem_reg[44][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n637 ) );
  MUX \Inst_Mem/U649  ( .IN0(\Inst_Mem/inst_mem_reg[46][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n636 ) );
  MUX \Inst_Mem/U648  ( .IN0(\Inst_Mem/n634 ), .IN1(\Inst_Mem/n627 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n635 ) );
  MUX \Inst_Mem/U647  ( .IN0(\Inst_Mem/n633 ), .IN1(\Inst_Mem/n630 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n634 ) );
  MUX \Inst_Mem/U646  ( .IN0(\Inst_Mem/n632 ), .IN1(\Inst_Mem/n631 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n633 ) );
  MUX \Inst_Mem/U645  ( .IN0(\Inst_Mem/inst_mem_reg[48][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n632 ) );
  MUX \Inst_Mem/U644  ( .IN0(\Inst_Mem/inst_mem_reg[50][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n631 ) );
  MUX \Inst_Mem/U643  ( .IN0(\Inst_Mem/n629 ), .IN1(\Inst_Mem/n628 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n630 ) );
  MUX \Inst_Mem/U642  ( .IN0(\Inst_Mem/inst_mem_reg[52][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n629 ) );
  MUX \Inst_Mem/U641  ( .IN0(\Inst_Mem/inst_mem_reg[54][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n628 ) );
  MUX \Inst_Mem/U640  ( .IN0(\Inst_Mem/n626 ), .IN1(\Inst_Mem/n623 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n627 ) );
  MUX \Inst_Mem/U639  ( .IN0(\Inst_Mem/n625 ), .IN1(\Inst_Mem/n624 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n626 ) );
  MUX \Inst_Mem/U638  ( .IN0(\Inst_Mem/inst_mem_reg[56][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n625 ) );
  MUX \Inst_Mem/U637  ( .IN0(\Inst_Mem/inst_mem_reg[58][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n624 ) );
  MUX \Inst_Mem/U636  ( .IN0(\Inst_Mem/n622 ), .IN1(\Inst_Mem/n621 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n623 ) );
  MUX \Inst_Mem/U635  ( .IN0(\Inst_Mem/inst_mem_reg[60][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n622 ) );
  MUX \Inst_Mem/U634  ( .IN0(\Inst_Mem/inst_mem_reg[62][10] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][10] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n621 ) );
  MUX \Inst_Mem/U633  ( .IN0(\Inst_Mem/n620 ), .IN1(\Inst_Mem/n589 ), .SEL(
        pc_current[7]), .F(imm[9]) );
  MUX \Inst_Mem/U632  ( .IN0(\Inst_Mem/n619 ), .IN1(\Inst_Mem/n604 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n620 ) );
  MUX \Inst_Mem/U631  ( .IN0(\Inst_Mem/n618 ), .IN1(\Inst_Mem/n611 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n619 ) );
  MUX \Inst_Mem/U630  ( .IN0(\Inst_Mem/n617 ), .IN1(\Inst_Mem/n614 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n618 ) );
  MUX \Inst_Mem/U629  ( .IN0(\Inst_Mem/n616 ), .IN1(\Inst_Mem/n615 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n617 ) );
  MUX \Inst_Mem/U628  ( .IN0(\Inst_Mem/inst_mem_reg[0][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n616 ) );
  MUX \Inst_Mem/U627  ( .IN0(\Inst_Mem/inst_mem_reg[2][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n615 ) );
  MUX \Inst_Mem/U626  ( .IN0(\Inst_Mem/n613 ), .IN1(\Inst_Mem/n612 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n614 ) );
  MUX \Inst_Mem/U625  ( .IN0(\Inst_Mem/inst_mem_reg[4][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n613 ) );
  MUX \Inst_Mem/U624  ( .IN0(\Inst_Mem/inst_mem_reg[6][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n612 ) );
  MUX \Inst_Mem/U623  ( .IN0(\Inst_Mem/n610 ), .IN1(\Inst_Mem/n607 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n611 ) );
  MUX \Inst_Mem/U622  ( .IN0(\Inst_Mem/n609 ), .IN1(\Inst_Mem/n608 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n610 ) );
  MUX \Inst_Mem/U621  ( .IN0(\Inst_Mem/inst_mem_reg[8][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n609 ) );
  MUX \Inst_Mem/U620  ( .IN0(\Inst_Mem/inst_mem_reg[10][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n608 ) );
  MUX \Inst_Mem/U619  ( .IN0(\Inst_Mem/n606 ), .IN1(\Inst_Mem/n605 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n607 ) );
  MUX \Inst_Mem/U618  ( .IN0(\Inst_Mem/inst_mem_reg[12][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n606 ) );
  MUX \Inst_Mem/U617  ( .IN0(\Inst_Mem/inst_mem_reg[14][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n605 ) );
  MUX \Inst_Mem/U616  ( .IN0(\Inst_Mem/n603 ), .IN1(\Inst_Mem/n596 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n604 ) );
  MUX \Inst_Mem/U615  ( .IN0(\Inst_Mem/n602 ), .IN1(\Inst_Mem/n599 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n603 ) );
  MUX \Inst_Mem/U614  ( .IN0(\Inst_Mem/n601 ), .IN1(\Inst_Mem/n600 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n602 ) );
  MUX \Inst_Mem/U613  ( .IN0(\Inst_Mem/inst_mem_reg[16][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n601 ) );
  MUX \Inst_Mem/U612  ( .IN0(\Inst_Mem/inst_mem_reg[18][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n600 ) );
  MUX \Inst_Mem/U611  ( .IN0(\Inst_Mem/n598 ), .IN1(\Inst_Mem/n597 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n599 ) );
  MUX \Inst_Mem/U610  ( .IN0(\Inst_Mem/inst_mem_reg[20][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n598 ) );
  MUX \Inst_Mem/U609  ( .IN0(\Inst_Mem/inst_mem_reg[22][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n597 ) );
  MUX \Inst_Mem/U608  ( .IN0(\Inst_Mem/n595 ), .IN1(\Inst_Mem/n592 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n596 ) );
  MUX \Inst_Mem/U607  ( .IN0(\Inst_Mem/n594 ), .IN1(\Inst_Mem/n593 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n595 ) );
  MUX \Inst_Mem/U606  ( .IN0(\Inst_Mem/inst_mem_reg[24][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n594 ) );
  MUX \Inst_Mem/U605  ( .IN0(\Inst_Mem/inst_mem_reg[26][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n593 ) );
  MUX \Inst_Mem/U604  ( .IN0(\Inst_Mem/n591 ), .IN1(\Inst_Mem/n590 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n592 ) );
  MUX \Inst_Mem/U603  ( .IN0(\Inst_Mem/inst_mem_reg[28][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n591 ) );
  MUX \Inst_Mem/U602  ( .IN0(\Inst_Mem/inst_mem_reg[30][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n590 ) );
  MUX \Inst_Mem/U601  ( .IN0(\Inst_Mem/n588 ), .IN1(\Inst_Mem/n573 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n589 ) );
  MUX \Inst_Mem/U600  ( .IN0(\Inst_Mem/n587 ), .IN1(\Inst_Mem/n580 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n588 ) );
  MUX \Inst_Mem/U599  ( .IN0(\Inst_Mem/n586 ), .IN1(\Inst_Mem/n583 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n587 ) );
  MUX \Inst_Mem/U598  ( .IN0(\Inst_Mem/n585 ), .IN1(\Inst_Mem/n584 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n586 ) );
  MUX \Inst_Mem/U597  ( .IN0(\Inst_Mem/inst_mem_reg[32][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n585 ) );
  MUX \Inst_Mem/U596  ( .IN0(\Inst_Mem/inst_mem_reg[34][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n584 ) );
  MUX \Inst_Mem/U595  ( .IN0(\Inst_Mem/n582 ), .IN1(\Inst_Mem/n581 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n583 ) );
  MUX \Inst_Mem/U594  ( .IN0(\Inst_Mem/inst_mem_reg[36][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n582 ) );
  MUX \Inst_Mem/U593  ( .IN0(\Inst_Mem/inst_mem_reg[38][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n581 ) );
  MUX \Inst_Mem/U592  ( .IN0(\Inst_Mem/n579 ), .IN1(\Inst_Mem/n576 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n580 ) );
  MUX \Inst_Mem/U591  ( .IN0(\Inst_Mem/n578 ), .IN1(\Inst_Mem/n577 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n579 ) );
  MUX \Inst_Mem/U590  ( .IN0(\Inst_Mem/inst_mem_reg[40][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n578 ) );
  MUX \Inst_Mem/U589  ( .IN0(\Inst_Mem/inst_mem_reg[42][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n577 ) );
  MUX \Inst_Mem/U588  ( .IN0(\Inst_Mem/n575 ), .IN1(\Inst_Mem/n574 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n576 ) );
  MUX \Inst_Mem/U587  ( .IN0(\Inst_Mem/inst_mem_reg[44][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n575 ) );
  MUX \Inst_Mem/U586  ( .IN0(\Inst_Mem/inst_mem_reg[46][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n574 ) );
  MUX \Inst_Mem/U585  ( .IN0(\Inst_Mem/n572 ), .IN1(\Inst_Mem/n565 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n573 ) );
  MUX \Inst_Mem/U584  ( .IN0(\Inst_Mem/n571 ), .IN1(\Inst_Mem/n568 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n572 ) );
  MUX \Inst_Mem/U583  ( .IN0(\Inst_Mem/n570 ), .IN1(\Inst_Mem/n569 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n571 ) );
  MUX \Inst_Mem/U582  ( .IN0(\Inst_Mem/inst_mem_reg[48][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n570 ) );
  MUX \Inst_Mem/U581  ( .IN0(\Inst_Mem/inst_mem_reg[50][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n569 ) );
  MUX \Inst_Mem/U580  ( .IN0(\Inst_Mem/n567 ), .IN1(\Inst_Mem/n566 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n568 ) );
  MUX \Inst_Mem/U579  ( .IN0(\Inst_Mem/inst_mem_reg[52][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n567 ) );
  MUX \Inst_Mem/U578  ( .IN0(\Inst_Mem/inst_mem_reg[54][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n566 ) );
  MUX \Inst_Mem/U577  ( .IN0(\Inst_Mem/n564 ), .IN1(\Inst_Mem/n561 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n565 ) );
  MUX \Inst_Mem/U576  ( .IN0(\Inst_Mem/n563 ), .IN1(\Inst_Mem/n562 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n564 ) );
  MUX \Inst_Mem/U575  ( .IN0(\Inst_Mem/inst_mem_reg[56][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n563 ) );
  MUX \Inst_Mem/U574  ( .IN0(\Inst_Mem/inst_mem_reg[58][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n562 ) );
  MUX \Inst_Mem/U573  ( .IN0(\Inst_Mem/n560 ), .IN1(\Inst_Mem/n559 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n561 ) );
  MUX \Inst_Mem/U572  ( .IN0(\Inst_Mem/inst_mem_reg[60][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n560 ) );
  MUX \Inst_Mem/U571  ( .IN0(\Inst_Mem/inst_mem_reg[62][9] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][9] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n559 ) );
  MUX \Inst_Mem/U570  ( .IN0(\Inst_Mem/n558 ), .IN1(\Inst_Mem/n527 ), .SEL(
        pc_current[7]), .F(imm[8]) );
  MUX \Inst_Mem/U569  ( .IN0(\Inst_Mem/n557 ), .IN1(\Inst_Mem/n542 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n558 ) );
  MUX \Inst_Mem/U568  ( .IN0(\Inst_Mem/n556 ), .IN1(\Inst_Mem/n549 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n557 ) );
  MUX \Inst_Mem/U567  ( .IN0(\Inst_Mem/n555 ), .IN1(\Inst_Mem/n552 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n556 ) );
  MUX \Inst_Mem/U566  ( .IN0(\Inst_Mem/n554 ), .IN1(\Inst_Mem/n553 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n555 ) );
  MUX \Inst_Mem/U565  ( .IN0(\Inst_Mem/inst_mem_reg[0][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n554 ) );
  MUX \Inst_Mem/U564  ( .IN0(\Inst_Mem/inst_mem_reg[2][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n553 ) );
  MUX \Inst_Mem/U563  ( .IN0(\Inst_Mem/n551 ), .IN1(\Inst_Mem/n550 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n552 ) );
  MUX \Inst_Mem/U562  ( .IN0(\Inst_Mem/inst_mem_reg[4][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n551 ) );
  MUX \Inst_Mem/U561  ( .IN0(\Inst_Mem/inst_mem_reg[6][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n550 ) );
  MUX \Inst_Mem/U560  ( .IN0(\Inst_Mem/n548 ), .IN1(\Inst_Mem/n545 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n549 ) );
  MUX \Inst_Mem/U559  ( .IN0(\Inst_Mem/n547 ), .IN1(\Inst_Mem/n546 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n548 ) );
  MUX \Inst_Mem/U558  ( .IN0(\Inst_Mem/inst_mem_reg[8][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n547 ) );
  MUX \Inst_Mem/U557  ( .IN0(\Inst_Mem/inst_mem_reg[10][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n546 ) );
  MUX \Inst_Mem/U556  ( .IN0(\Inst_Mem/n544 ), .IN1(\Inst_Mem/n543 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n545 ) );
  MUX \Inst_Mem/U555  ( .IN0(\Inst_Mem/inst_mem_reg[12][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n544 ) );
  MUX \Inst_Mem/U554  ( .IN0(\Inst_Mem/inst_mem_reg[14][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n543 ) );
  MUX \Inst_Mem/U553  ( .IN0(\Inst_Mem/n541 ), .IN1(\Inst_Mem/n534 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n542 ) );
  MUX \Inst_Mem/U552  ( .IN0(\Inst_Mem/n540 ), .IN1(\Inst_Mem/n537 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n541 ) );
  MUX \Inst_Mem/U551  ( .IN0(\Inst_Mem/n539 ), .IN1(\Inst_Mem/n538 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n540 ) );
  MUX \Inst_Mem/U550  ( .IN0(\Inst_Mem/inst_mem_reg[16][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n539 ) );
  MUX \Inst_Mem/U549  ( .IN0(\Inst_Mem/inst_mem_reg[18][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n538 ) );
  MUX \Inst_Mem/U548  ( .IN0(\Inst_Mem/n536 ), .IN1(\Inst_Mem/n535 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n537 ) );
  MUX \Inst_Mem/U547  ( .IN0(\Inst_Mem/inst_mem_reg[20][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n536 ) );
  MUX \Inst_Mem/U546  ( .IN0(\Inst_Mem/inst_mem_reg[22][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n535 ) );
  MUX \Inst_Mem/U545  ( .IN0(\Inst_Mem/n533 ), .IN1(\Inst_Mem/n530 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n534 ) );
  MUX \Inst_Mem/U544  ( .IN0(\Inst_Mem/n532 ), .IN1(\Inst_Mem/n531 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n533 ) );
  MUX \Inst_Mem/U543  ( .IN0(\Inst_Mem/inst_mem_reg[24][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n532 ) );
  MUX \Inst_Mem/U542  ( .IN0(\Inst_Mem/inst_mem_reg[26][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n531 ) );
  MUX \Inst_Mem/U541  ( .IN0(\Inst_Mem/n529 ), .IN1(\Inst_Mem/n528 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n530 ) );
  MUX \Inst_Mem/U540  ( .IN0(\Inst_Mem/inst_mem_reg[28][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n529 ) );
  MUX \Inst_Mem/U539  ( .IN0(\Inst_Mem/inst_mem_reg[30][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n528 ) );
  MUX \Inst_Mem/U538  ( .IN0(\Inst_Mem/n526 ), .IN1(\Inst_Mem/n511 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n527 ) );
  MUX \Inst_Mem/U537  ( .IN0(\Inst_Mem/n525 ), .IN1(\Inst_Mem/n518 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n526 ) );
  MUX \Inst_Mem/U536  ( .IN0(\Inst_Mem/n524 ), .IN1(\Inst_Mem/n521 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n525 ) );
  MUX \Inst_Mem/U535  ( .IN0(\Inst_Mem/n523 ), .IN1(\Inst_Mem/n522 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n524 ) );
  MUX \Inst_Mem/U534  ( .IN0(\Inst_Mem/inst_mem_reg[32][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n523 ) );
  MUX \Inst_Mem/U533  ( .IN0(\Inst_Mem/inst_mem_reg[34][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n522 ) );
  MUX \Inst_Mem/U532  ( .IN0(\Inst_Mem/n520 ), .IN1(\Inst_Mem/n519 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n521 ) );
  MUX \Inst_Mem/U531  ( .IN0(\Inst_Mem/inst_mem_reg[36][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n520 ) );
  MUX \Inst_Mem/U530  ( .IN0(\Inst_Mem/inst_mem_reg[38][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n519 ) );
  MUX \Inst_Mem/U529  ( .IN0(\Inst_Mem/n517 ), .IN1(\Inst_Mem/n514 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n518 ) );
  MUX \Inst_Mem/U528  ( .IN0(\Inst_Mem/n516 ), .IN1(\Inst_Mem/n515 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n517 ) );
  MUX \Inst_Mem/U527  ( .IN0(\Inst_Mem/inst_mem_reg[40][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n516 ) );
  MUX \Inst_Mem/U526  ( .IN0(\Inst_Mem/inst_mem_reg[42][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n515 ) );
  MUX \Inst_Mem/U525  ( .IN0(\Inst_Mem/n513 ), .IN1(\Inst_Mem/n512 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n514 ) );
  MUX \Inst_Mem/U524  ( .IN0(\Inst_Mem/inst_mem_reg[44][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n513 ) );
  MUX \Inst_Mem/U523  ( .IN0(\Inst_Mem/inst_mem_reg[46][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n512 ) );
  MUX \Inst_Mem/U522  ( .IN0(\Inst_Mem/n510 ), .IN1(\Inst_Mem/n503 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n511 ) );
  MUX \Inst_Mem/U521  ( .IN0(\Inst_Mem/n509 ), .IN1(\Inst_Mem/n506 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n510 ) );
  MUX \Inst_Mem/U520  ( .IN0(\Inst_Mem/n508 ), .IN1(\Inst_Mem/n507 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n509 ) );
  MUX \Inst_Mem/U519  ( .IN0(\Inst_Mem/inst_mem_reg[48][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n508 ) );
  MUX \Inst_Mem/U518  ( .IN0(\Inst_Mem/inst_mem_reg[50][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n507 ) );
  MUX \Inst_Mem/U517  ( .IN0(\Inst_Mem/n505 ), .IN1(\Inst_Mem/n504 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n506 ) );
  MUX \Inst_Mem/U516  ( .IN0(\Inst_Mem/inst_mem_reg[52][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n505 ) );
  MUX \Inst_Mem/U515  ( .IN0(\Inst_Mem/inst_mem_reg[54][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n504 ) );
  MUX \Inst_Mem/U514  ( .IN0(\Inst_Mem/n502 ), .IN1(\Inst_Mem/n499 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n503 ) );
  MUX \Inst_Mem/U513  ( .IN0(\Inst_Mem/n501 ), .IN1(\Inst_Mem/n500 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n502 ) );
  MUX \Inst_Mem/U512  ( .IN0(\Inst_Mem/inst_mem_reg[56][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n501 ) );
  MUX \Inst_Mem/U511  ( .IN0(\Inst_Mem/inst_mem_reg[58][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n500 ) );
  MUX \Inst_Mem/U510  ( .IN0(\Inst_Mem/n498 ), .IN1(\Inst_Mem/n497 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n499 ) );
  MUX \Inst_Mem/U509  ( .IN0(\Inst_Mem/inst_mem_reg[60][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n498 ) );
  MUX \Inst_Mem/U508  ( .IN0(\Inst_Mem/inst_mem_reg[62][8] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][8] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n497 ) );
  MUX \Inst_Mem/U507  ( .IN0(\Inst_Mem/n496 ), .IN1(\Inst_Mem/n465 ), .SEL(
        pc_current[7]), .F(imm[7]) );
  MUX \Inst_Mem/U506  ( .IN0(\Inst_Mem/n495 ), .IN1(\Inst_Mem/n480 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n496 ) );
  MUX \Inst_Mem/U505  ( .IN0(\Inst_Mem/n494 ), .IN1(\Inst_Mem/n487 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n495 ) );
  MUX \Inst_Mem/U504  ( .IN0(\Inst_Mem/n493 ), .IN1(\Inst_Mem/n490 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n494 ) );
  MUX \Inst_Mem/U503  ( .IN0(\Inst_Mem/n492 ), .IN1(\Inst_Mem/n491 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n493 ) );
  MUX \Inst_Mem/U502  ( .IN0(\Inst_Mem/inst_mem_reg[0][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n492 ) );
  MUX \Inst_Mem/U501  ( .IN0(\Inst_Mem/inst_mem_reg[2][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n491 ) );
  MUX \Inst_Mem/U500  ( .IN0(\Inst_Mem/n489 ), .IN1(\Inst_Mem/n488 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n490 ) );
  MUX \Inst_Mem/U499  ( .IN0(\Inst_Mem/inst_mem_reg[4][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n489 ) );
  MUX \Inst_Mem/U498  ( .IN0(\Inst_Mem/inst_mem_reg[6][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n488 ) );
  MUX \Inst_Mem/U497  ( .IN0(\Inst_Mem/n486 ), .IN1(\Inst_Mem/n483 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n487 ) );
  MUX \Inst_Mem/U496  ( .IN0(\Inst_Mem/n485 ), .IN1(\Inst_Mem/n484 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n486 ) );
  MUX \Inst_Mem/U495  ( .IN0(\Inst_Mem/inst_mem_reg[8][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n485 ) );
  MUX \Inst_Mem/U494  ( .IN0(\Inst_Mem/inst_mem_reg[10][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n484 ) );
  MUX \Inst_Mem/U493  ( .IN0(\Inst_Mem/n482 ), .IN1(\Inst_Mem/n481 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n483 ) );
  MUX \Inst_Mem/U492  ( .IN0(\Inst_Mem/inst_mem_reg[12][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n482 ) );
  MUX \Inst_Mem/U491  ( .IN0(\Inst_Mem/inst_mem_reg[14][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n481 ) );
  MUX \Inst_Mem/U490  ( .IN0(\Inst_Mem/n479 ), .IN1(\Inst_Mem/n472 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n480 ) );
  MUX \Inst_Mem/U489  ( .IN0(\Inst_Mem/n478 ), .IN1(\Inst_Mem/n475 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n479 ) );
  MUX \Inst_Mem/U488  ( .IN0(\Inst_Mem/n477 ), .IN1(\Inst_Mem/n476 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n478 ) );
  MUX \Inst_Mem/U487  ( .IN0(\Inst_Mem/inst_mem_reg[16][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n477 ) );
  MUX \Inst_Mem/U486  ( .IN0(\Inst_Mem/inst_mem_reg[18][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n476 ) );
  MUX \Inst_Mem/U485  ( .IN0(\Inst_Mem/n474 ), .IN1(\Inst_Mem/n473 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n475 ) );
  MUX \Inst_Mem/U484  ( .IN0(\Inst_Mem/inst_mem_reg[20][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n474 ) );
  MUX \Inst_Mem/U483  ( .IN0(\Inst_Mem/inst_mem_reg[22][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n473 ) );
  MUX \Inst_Mem/U482  ( .IN0(\Inst_Mem/n471 ), .IN1(\Inst_Mem/n468 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n472 ) );
  MUX \Inst_Mem/U481  ( .IN0(\Inst_Mem/n470 ), .IN1(\Inst_Mem/n469 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n471 ) );
  MUX \Inst_Mem/U480  ( .IN0(\Inst_Mem/inst_mem_reg[24][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n470 ) );
  MUX \Inst_Mem/U479  ( .IN0(\Inst_Mem/inst_mem_reg[26][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n469 ) );
  MUX \Inst_Mem/U478  ( .IN0(\Inst_Mem/n467 ), .IN1(\Inst_Mem/n466 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n468 ) );
  MUX \Inst_Mem/U477  ( .IN0(\Inst_Mem/inst_mem_reg[28][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n467 ) );
  MUX \Inst_Mem/U476  ( .IN0(\Inst_Mem/inst_mem_reg[30][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n466 ) );
  MUX \Inst_Mem/U475  ( .IN0(\Inst_Mem/n464 ), .IN1(\Inst_Mem/n449 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n465 ) );
  MUX \Inst_Mem/U474  ( .IN0(\Inst_Mem/n463 ), .IN1(\Inst_Mem/n456 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n464 ) );
  MUX \Inst_Mem/U473  ( .IN0(\Inst_Mem/n462 ), .IN1(\Inst_Mem/n459 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n463 ) );
  MUX \Inst_Mem/U472  ( .IN0(\Inst_Mem/n461 ), .IN1(\Inst_Mem/n460 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n462 ) );
  MUX \Inst_Mem/U471  ( .IN0(\Inst_Mem/inst_mem_reg[32][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n461 ) );
  MUX \Inst_Mem/U470  ( .IN0(\Inst_Mem/inst_mem_reg[34][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n460 ) );
  MUX \Inst_Mem/U469  ( .IN0(\Inst_Mem/n458 ), .IN1(\Inst_Mem/n457 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n459 ) );
  MUX \Inst_Mem/U468  ( .IN0(\Inst_Mem/inst_mem_reg[36][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n458 ) );
  MUX \Inst_Mem/U467  ( .IN0(\Inst_Mem/inst_mem_reg[38][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n457 ) );
  MUX \Inst_Mem/U466  ( .IN0(\Inst_Mem/n455 ), .IN1(\Inst_Mem/n452 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n456 ) );
  MUX \Inst_Mem/U465  ( .IN0(\Inst_Mem/n454 ), .IN1(\Inst_Mem/n453 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n455 ) );
  MUX \Inst_Mem/U464  ( .IN0(\Inst_Mem/inst_mem_reg[40][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n454 ) );
  MUX \Inst_Mem/U463  ( .IN0(\Inst_Mem/inst_mem_reg[42][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n453 ) );
  MUX \Inst_Mem/U462  ( .IN0(\Inst_Mem/n451 ), .IN1(\Inst_Mem/n450 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n452 ) );
  MUX \Inst_Mem/U461  ( .IN0(\Inst_Mem/inst_mem_reg[44][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n451 ) );
  MUX \Inst_Mem/U460  ( .IN0(\Inst_Mem/inst_mem_reg[46][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n450 ) );
  MUX \Inst_Mem/U459  ( .IN0(\Inst_Mem/n448 ), .IN1(\Inst_Mem/n441 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n449 ) );
  MUX \Inst_Mem/U458  ( .IN0(\Inst_Mem/n447 ), .IN1(\Inst_Mem/n444 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n448 ) );
  MUX \Inst_Mem/U457  ( .IN0(\Inst_Mem/n446 ), .IN1(\Inst_Mem/n445 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n447 ) );
  MUX \Inst_Mem/U456  ( .IN0(\Inst_Mem/inst_mem_reg[48][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n446 ) );
  MUX \Inst_Mem/U455  ( .IN0(\Inst_Mem/inst_mem_reg[50][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n445 ) );
  MUX \Inst_Mem/U454  ( .IN0(\Inst_Mem/n443 ), .IN1(\Inst_Mem/n442 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n444 ) );
  MUX \Inst_Mem/U453  ( .IN0(\Inst_Mem/inst_mem_reg[52][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n443 ) );
  MUX \Inst_Mem/U452  ( .IN0(\Inst_Mem/inst_mem_reg[54][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n442 ) );
  MUX \Inst_Mem/U451  ( .IN0(\Inst_Mem/n440 ), .IN1(\Inst_Mem/n437 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n441 ) );
  MUX \Inst_Mem/U450  ( .IN0(\Inst_Mem/n439 ), .IN1(\Inst_Mem/n438 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n440 ) );
  MUX \Inst_Mem/U449  ( .IN0(\Inst_Mem/inst_mem_reg[56][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n439 ) );
  MUX \Inst_Mem/U448  ( .IN0(\Inst_Mem/inst_mem_reg[58][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n438 ) );
  MUX \Inst_Mem/U447  ( .IN0(\Inst_Mem/n436 ), .IN1(\Inst_Mem/n435 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n437 ) );
  MUX \Inst_Mem/U446  ( .IN0(\Inst_Mem/inst_mem_reg[60][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n436 ) );
  MUX \Inst_Mem/U445  ( .IN0(\Inst_Mem/inst_mem_reg[62][7] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][7] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n435 ) );
  MUX \Inst_Mem/U444  ( .IN0(\Inst_Mem/n434 ), .IN1(\Inst_Mem/n403 ), .SEL(
        pc_current[7]), .F(imm[6]) );
  MUX \Inst_Mem/U443  ( .IN0(\Inst_Mem/n433 ), .IN1(\Inst_Mem/n418 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n434 ) );
  MUX \Inst_Mem/U442  ( .IN0(\Inst_Mem/n432 ), .IN1(\Inst_Mem/n425 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n433 ) );
  MUX \Inst_Mem/U441  ( .IN0(\Inst_Mem/n431 ), .IN1(\Inst_Mem/n428 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n432 ) );
  MUX \Inst_Mem/U440  ( .IN0(\Inst_Mem/n430 ), .IN1(\Inst_Mem/n429 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n431 ) );
  MUX \Inst_Mem/U439  ( .IN0(\Inst_Mem/inst_mem_reg[0][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n430 ) );
  MUX \Inst_Mem/U438  ( .IN0(\Inst_Mem/inst_mem_reg[2][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n429 ) );
  MUX \Inst_Mem/U437  ( .IN0(\Inst_Mem/n427 ), .IN1(\Inst_Mem/n426 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n428 ) );
  MUX \Inst_Mem/U436  ( .IN0(\Inst_Mem/inst_mem_reg[4][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n427 ) );
  MUX \Inst_Mem/U435  ( .IN0(\Inst_Mem/inst_mem_reg[6][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n426 ) );
  MUX \Inst_Mem/U434  ( .IN0(\Inst_Mem/n424 ), .IN1(\Inst_Mem/n421 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n425 ) );
  MUX \Inst_Mem/U433  ( .IN0(\Inst_Mem/n423 ), .IN1(\Inst_Mem/n422 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n424 ) );
  MUX \Inst_Mem/U432  ( .IN0(\Inst_Mem/inst_mem_reg[8][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n423 ) );
  MUX \Inst_Mem/U431  ( .IN0(\Inst_Mem/inst_mem_reg[10][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n422 ) );
  MUX \Inst_Mem/U430  ( .IN0(\Inst_Mem/n420 ), .IN1(\Inst_Mem/n419 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n421 ) );
  MUX \Inst_Mem/U429  ( .IN0(\Inst_Mem/inst_mem_reg[12][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n420 ) );
  MUX \Inst_Mem/U428  ( .IN0(\Inst_Mem/inst_mem_reg[14][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n419 ) );
  MUX \Inst_Mem/U427  ( .IN0(\Inst_Mem/n417 ), .IN1(\Inst_Mem/n410 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n418 ) );
  MUX \Inst_Mem/U426  ( .IN0(\Inst_Mem/n416 ), .IN1(\Inst_Mem/n413 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n417 ) );
  MUX \Inst_Mem/U425  ( .IN0(\Inst_Mem/n415 ), .IN1(\Inst_Mem/n414 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n416 ) );
  MUX \Inst_Mem/U424  ( .IN0(\Inst_Mem/inst_mem_reg[16][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n415 ) );
  MUX \Inst_Mem/U423  ( .IN0(\Inst_Mem/inst_mem_reg[18][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n414 ) );
  MUX \Inst_Mem/U422  ( .IN0(\Inst_Mem/n412 ), .IN1(\Inst_Mem/n411 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n413 ) );
  MUX \Inst_Mem/U421  ( .IN0(\Inst_Mem/inst_mem_reg[20][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n412 ) );
  MUX \Inst_Mem/U420  ( .IN0(\Inst_Mem/inst_mem_reg[22][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n411 ) );
  MUX \Inst_Mem/U419  ( .IN0(\Inst_Mem/n409 ), .IN1(\Inst_Mem/n406 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n410 ) );
  MUX \Inst_Mem/U418  ( .IN0(\Inst_Mem/n408 ), .IN1(\Inst_Mem/n407 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n409 ) );
  MUX \Inst_Mem/U417  ( .IN0(\Inst_Mem/inst_mem_reg[24][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n408 ) );
  MUX \Inst_Mem/U416  ( .IN0(\Inst_Mem/inst_mem_reg[26][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n407 ) );
  MUX \Inst_Mem/U415  ( .IN0(\Inst_Mem/n405 ), .IN1(\Inst_Mem/n404 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n406 ) );
  MUX \Inst_Mem/U414  ( .IN0(\Inst_Mem/inst_mem_reg[28][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n405 ) );
  MUX \Inst_Mem/U413  ( .IN0(\Inst_Mem/inst_mem_reg[30][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n404 ) );
  MUX \Inst_Mem/U412  ( .IN0(\Inst_Mem/n402 ), .IN1(\Inst_Mem/n387 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n403 ) );
  MUX \Inst_Mem/U411  ( .IN0(\Inst_Mem/n401 ), .IN1(\Inst_Mem/n394 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n402 ) );
  MUX \Inst_Mem/U410  ( .IN0(\Inst_Mem/n400 ), .IN1(\Inst_Mem/n397 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n401 ) );
  MUX \Inst_Mem/U409  ( .IN0(\Inst_Mem/n399 ), .IN1(\Inst_Mem/n398 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n400 ) );
  MUX \Inst_Mem/U408  ( .IN0(\Inst_Mem/inst_mem_reg[32][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n399 ) );
  MUX \Inst_Mem/U407  ( .IN0(\Inst_Mem/inst_mem_reg[34][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n398 ) );
  MUX \Inst_Mem/U406  ( .IN0(\Inst_Mem/n396 ), .IN1(\Inst_Mem/n395 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n397 ) );
  MUX \Inst_Mem/U405  ( .IN0(\Inst_Mem/inst_mem_reg[36][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n396 ) );
  MUX \Inst_Mem/U404  ( .IN0(\Inst_Mem/inst_mem_reg[38][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n395 ) );
  MUX \Inst_Mem/U403  ( .IN0(\Inst_Mem/n393 ), .IN1(\Inst_Mem/n390 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n394 ) );
  MUX \Inst_Mem/U402  ( .IN0(\Inst_Mem/n392 ), .IN1(\Inst_Mem/n391 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n393 ) );
  MUX \Inst_Mem/U401  ( .IN0(\Inst_Mem/inst_mem_reg[40][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n392 ) );
  MUX \Inst_Mem/U400  ( .IN0(\Inst_Mem/inst_mem_reg[42][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n391 ) );
  MUX \Inst_Mem/U399  ( .IN0(\Inst_Mem/n389 ), .IN1(\Inst_Mem/n388 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n390 ) );
  MUX \Inst_Mem/U398  ( .IN0(\Inst_Mem/inst_mem_reg[44][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n389 ) );
  MUX \Inst_Mem/U397  ( .IN0(\Inst_Mem/inst_mem_reg[46][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n388 ) );
  MUX \Inst_Mem/U396  ( .IN0(\Inst_Mem/n386 ), .IN1(\Inst_Mem/n379 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n387 ) );
  MUX \Inst_Mem/U395  ( .IN0(\Inst_Mem/n385 ), .IN1(\Inst_Mem/n382 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n386 ) );
  MUX \Inst_Mem/U394  ( .IN0(\Inst_Mem/n384 ), .IN1(\Inst_Mem/n383 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n385 ) );
  MUX \Inst_Mem/U393  ( .IN0(\Inst_Mem/inst_mem_reg[48][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n384 ) );
  MUX \Inst_Mem/U392  ( .IN0(\Inst_Mem/inst_mem_reg[50][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n383 ) );
  MUX \Inst_Mem/U391  ( .IN0(\Inst_Mem/n381 ), .IN1(\Inst_Mem/n380 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n382 ) );
  MUX \Inst_Mem/U390  ( .IN0(\Inst_Mem/inst_mem_reg[52][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n381 ) );
  MUX \Inst_Mem/U389  ( .IN0(\Inst_Mem/inst_mem_reg[54][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n380 ) );
  MUX \Inst_Mem/U388  ( .IN0(\Inst_Mem/n378 ), .IN1(\Inst_Mem/n375 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n379 ) );
  MUX \Inst_Mem/U387  ( .IN0(\Inst_Mem/n377 ), .IN1(\Inst_Mem/n376 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n378 ) );
  MUX \Inst_Mem/U386  ( .IN0(\Inst_Mem/inst_mem_reg[56][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n377 ) );
  MUX \Inst_Mem/U385  ( .IN0(\Inst_Mem/inst_mem_reg[58][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n376 ) );
  MUX \Inst_Mem/U384  ( .IN0(\Inst_Mem/n374 ), .IN1(\Inst_Mem/n373 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n375 ) );
  MUX \Inst_Mem/U383  ( .IN0(\Inst_Mem/inst_mem_reg[60][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n374 ) );
  MUX \Inst_Mem/U382  ( .IN0(\Inst_Mem/inst_mem_reg[62][6] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][6] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n373 ) );
  MUX \Inst_Mem/U381  ( .IN0(\Inst_Mem/n372 ), .IN1(\Inst_Mem/n341 ), .SEL(
        pc_current[7]), .F(imm[5]) );
  MUX \Inst_Mem/U380  ( .IN0(\Inst_Mem/n371 ), .IN1(\Inst_Mem/n356 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n372 ) );
  MUX \Inst_Mem/U379  ( .IN0(\Inst_Mem/n370 ), .IN1(\Inst_Mem/n363 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n371 ) );
  MUX \Inst_Mem/U378  ( .IN0(\Inst_Mem/n369 ), .IN1(\Inst_Mem/n366 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n370 ) );
  MUX \Inst_Mem/U377  ( .IN0(\Inst_Mem/n368 ), .IN1(\Inst_Mem/n367 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n369 ) );
  MUX \Inst_Mem/U376  ( .IN0(\Inst_Mem/inst_mem_reg[0][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n368 ) );
  MUX \Inst_Mem/U375  ( .IN0(\Inst_Mem/inst_mem_reg[2][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n367 ) );
  MUX \Inst_Mem/U374  ( .IN0(\Inst_Mem/n365 ), .IN1(\Inst_Mem/n364 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n366 ) );
  MUX \Inst_Mem/U373  ( .IN0(\Inst_Mem/inst_mem_reg[4][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n365 ) );
  MUX \Inst_Mem/U372  ( .IN0(\Inst_Mem/inst_mem_reg[6][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n364 ) );
  MUX \Inst_Mem/U371  ( .IN0(\Inst_Mem/n362 ), .IN1(\Inst_Mem/n359 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n363 ) );
  MUX \Inst_Mem/U370  ( .IN0(\Inst_Mem/n361 ), .IN1(\Inst_Mem/n360 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n362 ) );
  MUX \Inst_Mem/U369  ( .IN0(\Inst_Mem/inst_mem_reg[8][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n361 ) );
  MUX \Inst_Mem/U368  ( .IN0(\Inst_Mem/inst_mem_reg[10][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n360 ) );
  MUX \Inst_Mem/U367  ( .IN0(\Inst_Mem/n358 ), .IN1(\Inst_Mem/n357 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n359 ) );
  MUX \Inst_Mem/U366  ( .IN0(\Inst_Mem/inst_mem_reg[12][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n358 ) );
  MUX \Inst_Mem/U365  ( .IN0(\Inst_Mem/inst_mem_reg[14][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n357 ) );
  MUX \Inst_Mem/U364  ( .IN0(\Inst_Mem/n355 ), .IN1(\Inst_Mem/n348 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n356 ) );
  MUX \Inst_Mem/U363  ( .IN0(\Inst_Mem/n354 ), .IN1(\Inst_Mem/n351 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n355 ) );
  MUX \Inst_Mem/U362  ( .IN0(\Inst_Mem/n353 ), .IN1(\Inst_Mem/n352 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n354 ) );
  MUX \Inst_Mem/U361  ( .IN0(\Inst_Mem/inst_mem_reg[16][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n353 ) );
  MUX \Inst_Mem/U360  ( .IN0(\Inst_Mem/inst_mem_reg[18][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n352 ) );
  MUX \Inst_Mem/U359  ( .IN0(\Inst_Mem/n350 ), .IN1(\Inst_Mem/n349 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n351 ) );
  MUX \Inst_Mem/U358  ( .IN0(\Inst_Mem/inst_mem_reg[20][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n350 ) );
  MUX \Inst_Mem/U357  ( .IN0(\Inst_Mem/inst_mem_reg[22][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n349 ) );
  MUX \Inst_Mem/U356  ( .IN0(\Inst_Mem/n347 ), .IN1(\Inst_Mem/n344 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n348 ) );
  MUX \Inst_Mem/U355  ( .IN0(\Inst_Mem/n346 ), .IN1(\Inst_Mem/n345 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n347 ) );
  MUX \Inst_Mem/U354  ( .IN0(\Inst_Mem/inst_mem_reg[24][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n346 ) );
  MUX \Inst_Mem/U353  ( .IN0(\Inst_Mem/inst_mem_reg[26][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n345 ) );
  MUX \Inst_Mem/U352  ( .IN0(\Inst_Mem/n343 ), .IN1(\Inst_Mem/n342 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n344 ) );
  MUX \Inst_Mem/U351  ( .IN0(\Inst_Mem/inst_mem_reg[28][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n343 ) );
  MUX \Inst_Mem/U350  ( .IN0(\Inst_Mem/inst_mem_reg[30][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n342 ) );
  MUX \Inst_Mem/U349  ( .IN0(\Inst_Mem/n340 ), .IN1(\Inst_Mem/n325 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n341 ) );
  MUX \Inst_Mem/U348  ( .IN0(\Inst_Mem/n339 ), .IN1(\Inst_Mem/n332 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n340 ) );
  MUX \Inst_Mem/U347  ( .IN0(\Inst_Mem/n338 ), .IN1(\Inst_Mem/n335 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n339 ) );
  MUX \Inst_Mem/U346  ( .IN0(\Inst_Mem/n337 ), .IN1(\Inst_Mem/n336 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n338 ) );
  MUX \Inst_Mem/U345  ( .IN0(\Inst_Mem/inst_mem_reg[32][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n337 ) );
  MUX \Inst_Mem/U344  ( .IN0(\Inst_Mem/inst_mem_reg[34][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n336 ) );
  MUX \Inst_Mem/U343  ( .IN0(\Inst_Mem/n334 ), .IN1(\Inst_Mem/n333 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n335 ) );
  MUX \Inst_Mem/U342  ( .IN0(\Inst_Mem/inst_mem_reg[36][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n334 ) );
  MUX \Inst_Mem/U341  ( .IN0(\Inst_Mem/inst_mem_reg[38][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n333 ) );
  MUX \Inst_Mem/U340  ( .IN0(\Inst_Mem/n331 ), .IN1(\Inst_Mem/n328 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n332 ) );
  MUX \Inst_Mem/U339  ( .IN0(\Inst_Mem/n330 ), .IN1(\Inst_Mem/n329 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n331 ) );
  MUX \Inst_Mem/U338  ( .IN0(\Inst_Mem/inst_mem_reg[40][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n330 ) );
  MUX \Inst_Mem/U337  ( .IN0(\Inst_Mem/inst_mem_reg[42][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n329 ) );
  MUX \Inst_Mem/U336  ( .IN0(\Inst_Mem/n327 ), .IN1(\Inst_Mem/n326 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n328 ) );
  MUX \Inst_Mem/U335  ( .IN0(\Inst_Mem/inst_mem_reg[44][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n327 ) );
  MUX \Inst_Mem/U334  ( .IN0(\Inst_Mem/inst_mem_reg[46][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n326 ) );
  MUX \Inst_Mem/U333  ( .IN0(\Inst_Mem/n324 ), .IN1(\Inst_Mem/n317 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n325 ) );
  MUX \Inst_Mem/U332  ( .IN0(\Inst_Mem/n323 ), .IN1(\Inst_Mem/n320 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n324 ) );
  MUX \Inst_Mem/U331  ( .IN0(\Inst_Mem/n322 ), .IN1(\Inst_Mem/n321 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n323 ) );
  MUX \Inst_Mem/U330  ( .IN0(\Inst_Mem/inst_mem_reg[48][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n322 ) );
  MUX \Inst_Mem/U329  ( .IN0(\Inst_Mem/inst_mem_reg[50][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n321 ) );
  MUX \Inst_Mem/U328  ( .IN0(\Inst_Mem/n319 ), .IN1(\Inst_Mem/n318 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n320 ) );
  MUX \Inst_Mem/U327  ( .IN0(\Inst_Mem/inst_mem_reg[52][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n319 ) );
  MUX \Inst_Mem/U326  ( .IN0(\Inst_Mem/inst_mem_reg[54][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n318 ) );
  MUX \Inst_Mem/U325  ( .IN0(\Inst_Mem/n316 ), .IN1(\Inst_Mem/n313 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n317 ) );
  MUX \Inst_Mem/U324  ( .IN0(\Inst_Mem/n315 ), .IN1(\Inst_Mem/n314 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n316 ) );
  MUX \Inst_Mem/U323  ( .IN0(\Inst_Mem/inst_mem_reg[56][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n315 ) );
  MUX \Inst_Mem/U322  ( .IN0(\Inst_Mem/inst_mem_reg[58][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n314 ) );
  MUX \Inst_Mem/U321  ( .IN0(\Inst_Mem/n312 ), .IN1(\Inst_Mem/n311 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n313 ) );
  MUX \Inst_Mem/U320  ( .IN0(\Inst_Mem/inst_mem_reg[60][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n312 ) );
  MUX \Inst_Mem/U319  ( .IN0(\Inst_Mem/inst_mem_reg[62][5] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][5] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n311 ) );
  MUX \Inst_Mem/U318  ( .IN0(\Inst_Mem/n310 ), .IN1(\Inst_Mem/n279 ), .SEL(
        pc_current[7]), .F(imm[4]) );
  MUX \Inst_Mem/U317  ( .IN0(\Inst_Mem/n309 ), .IN1(\Inst_Mem/n294 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n310 ) );
  MUX \Inst_Mem/U316  ( .IN0(\Inst_Mem/n308 ), .IN1(\Inst_Mem/n301 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n309 ) );
  MUX \Inst_Mem/U315  ( .IN0(\Inst_Mem/n307 ), .IN1(\Inst_Mem/n304 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n308 ) );
  MUX \Inst_Mem/U314  ( .IN0(\Inst_Mem/n306 ), .IN1(\Inst_Mem/n305 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n307 ) );
  MUX \Inst_Mem/U313  ( .IN0(\Inst_Mem/inst_mem_reg[0][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n306 ) );
  MUX \Inst_Mem/U312  ( .IN0(\Inst_Mem/inst_mem_reg[2][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n305 ) );
  MUX \Inst_Mem/U311  ( .IN0(\Inst_Mem/n303 ), .IN1(\Inst_Mem/n302 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n304 ) );
  MUX \Inst_Mem/U310  ( .IN0(\Inst_Mem/inst_mem_reg[4][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n303 ) );
  MUX \Inst_Mem/U309  ( .IN0(\Inst_Mem/inst_mem_reg[6][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n302 ) );
  MUX \Inst_Mem/U308  ( .IN0(\Inst_Mem/n300 ), .IN1(\Inst_Mem/n297 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n301 ) );
  MUX \Inst_Mem/U307  ( .IN0(\Inst_Mem/n299 ), .IN1(\Inst_Mem/n298 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n300 ) );
  MUX \Inst_Mem/U306  ( .IN0(\Inst_Mem/inst_mem_reg[8][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n299 ) );
  MUX \Inst_Mem/U305  ( .IN0(\Inst_Mem/inst_mem_reg[10][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n298 ) );
  MUX \Inst_Mem/U304  ( .IN0(\Inst_Mem/n296 ), .IN1(\Inst_Mem/n295 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n297 ) );
  MUX \Inst_Mem/U303  ( .IN0(\Inst_Mem/inst_mem_reg[12][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n296 ) );
  MUX \Inst_Mem/U302  ( .IN0(\Inst_Mem/inst_mem_reg[14][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n295 ) );
  MUX \Inst_Mem/U301  ( .IN0(\Inst_Mem/n293 ), .IN1(\Inst_Mem/n286 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n294 ) );
  MUX \Inst_Mem/U300  ( .IN0(\Inst_Mem/n292 ), .IN1(\Inst_Mem/n289 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n293 ) );
  MUX \Inst_Mem/U299  ( .IN0(\Inst_Mem/n291 ), .IN1(\Inst_Mem/n290 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n292 ) );
  MUX \Inst_Mem/U298  ( .IN0(\Inst_Mem/inst_mem_reg[16][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n291 ) );
  MUX \Inst_Mem/U297  ( .IN0(\Inst_Mem/inst_mem_reg[18][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n290 ) );
  MUX \Inst_Mem/U296  ( .IN0(\Inst_Mem/n288 ), .IN1(\Inst_Mem/n287 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n289 ) );
  MUX \Inst_Mem/U295  ( .IN0(\Inst_Mem/inst_mem_reg[20][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n288 ) );
  MUX \Inst_Mem/U294  ( .IN0(\Inst_Mem/inst_mem_reg[22][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n287 ) );
  MUX \Inst_Mem/U293  ( .IN0(\Inst_Mem/n285 ), .IN1(\Inst_Mem/n282 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n286 ) );
  MUX \Inst_Mem/U292  ( .IN0(\Inst_Mem/n284 ), .IN1(\Inst_Mem/n283 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n285 ) );
  MUX \Inst_Mem/U291  ( .IN0(\Inst_Mem/inst_mem_reg[24][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n284 ) );
  MUX \Inst_Mem/U290  ( .IN0(\Inst_Mem/inst_mem_reg[26][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n283 ) );
  MUX \Inst_Mem/U289  ( .IN0(\Inst_Mem/n281 ), .IN1(\Inst_Mem/n280 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n282 ) );
  MUX \Inst_Mem/U288  ( .IN0(\Inst_Mem/inst_mem_reg[28][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n281 ) );
  MUX \Inst_Mem/U287  ( .IN0(\Inst_Mem/inst_mem_reg[30][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n280 ) );
  MUX \Inst_Mem/U286  ( .IN0(\Inst_Mem/n278 ), .IN1(\Inst_Mem/n263 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n279 ) );
  MUX \Inst_Mem/U285  ( .IN0(\Inst_Mem/n277 ), .IN1(\Inst_Mem/n270 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n278 ) );
  MUX \Inst_Mem/U284  ( .IN0(\Inst_Mem/n276 ), .IN1(\Inst_Mem/n273 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n277 ) );
  MUX \Inst_Mem/U283  ( .IN0(\Inst_Mem/n275 ), .IN1(\Inst_Mem/n274 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n276 ) );
  MUX \Inst_Mem/U282  ( .IN0(\Inst_Mem/inst_mem_reg[32][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n275 ) );
  MUX \Inst_Mem/U281  ( .IN0(\Inst_Mem/inst_mem_reg[34][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n274 ) );
  MUX \Inst_Mem/U280  ( .IN0(\Inst_Mem/n272 ), .IN1(\Inst_Mem/n271 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n273 ) );
  MUX \Inst_Mem/U279  ( .IN0(\Inst_Mem/inst_mem_reg[36][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n272 ) );
  MUX \Inst_Mem/U278  ( .IN0(\Inst_Mem/inst_mem_reg[38][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n271 ) );
  MUX \Inst_Mem/U277  ( .IN0(\Inst_Mem/n269 ), .IN1(\Inst_Mem/n266 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n270 ) );
  MUX \Inst_Mem/U276  ( .IN0(\Inst_Mem/n268 ), .IN1(\Inst_Mem/n267 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n269 ) );
  MUX \Inst_Mem/U275  ( .IN0(\Inst_Mem/inst_mem_reg[40][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n268 ) );
  MUX \Inst_Mem/U274  ( .IN0(\Inst_Mem/inst_mem_reg[42][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n267 ) );
  MUX \Inst_Mem/U273  ( .IN0(\Inst_Mem/n265 ), .IN1(\Inst_Mem/n264 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n266 ) );
  MUX \Inst_Mem/U272  ( .IN0(\Inst_Mem/inst_mem_reg[44][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n265 ) );
  MUX \Inst_Mem/U271  ( .IN0(\Inst_Mem/inst_mem_reg[46][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n264 ) );
  MUX \Inst_Mem/U270  ( .IN0(\Inst_Mem/n262 ), .IN1(\Inst_Mem/n255 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n263 ) );
  MUX \Inst_Mem/U269  ( .IN0(\Inst_Mem/n261 ), .IN1(\Inst_Mem/n258 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n262 ) );
  MUX \Inst_Mem/U268  ( .IN0(\Inst_Mem/n260 ), .IN1(\Inst_Mem/n259 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n261 ) );
  MUX \Inst_Mem/U267  ( .IN0(\Inst_Mem/inst_mem_reg[48][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n260 ) );
  MUX \Inst_Mem/U266  ( .IN0(\Inst_Mem/inst_mem_reg[50][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n259 ) );
  MUX \Inst_Mem/U265  ( .IN0(\Inst_Mem/n257 ), .IN1(\Inst_Mem/n256 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n258 ) );
  MUX \Inst_Mem/U264  ( .IN0(\Inst_Mem/inst_mem_reg[52][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n257 ) );
  MUX \Inst_Mem/U263  ( .IN0(\Inst_Mem/inst_mem_reg[54][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n256 ) );
  MUX \Inst_Mem/U262  ( .IN0(\Inst_Mem/n254 ), .IN1(\Inst_Mem/n251 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n255 ) );
  MUX \Inst_Mem/U261  ( .IN0(\Inst_Mem/n253 ), .IN1(\Inst_Mem/n252 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n254 ) );
  MUX \Inst_Mem/U260  ( .IN0(\Inst_Mem/inst_mem_reg[56][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n253 ) );
  MUX \Inst_Mem/U259  ( .IN0(\Inst_Mem/inst_mem_reg[58][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n252 ) );
  MUX \Inst_Mem/U258  ( .IN0(\Inst_Mem/n250 ), .IN1(\Inst_Mem/n249 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n251 ) );
  MUX \Inst_Mem/U257  ( .IN0(\Inst_Mem/inst_mem_reg[60][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n250 ) );
  MUX \Inst_Mem/U256  ( .IN0(\Inst_Mem/inst_mem_reg[62][4] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][4] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n249 ) );
  MUX \Inst_Mem/U255  ( .IN0(\Inst_Mem/n248 ), .IN1(\Inst_Mem/n217 ), .SEL(
        pc_current[7]), .F(imm[3]) );
  MUX \Inst_Mem/U254  ( .IN0(\Inst_Mem/n247 ), .IN1(\Inst_Mem/n232 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n248 ) );
  MUX \Inst_Mem/U253  ( .IN0(\Inst_Mem/n246 ), .IN1(\Inst_Mem/n239 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n247 ) );
  MUX \Inst_Mem/U252  ( .IN0(\Inst_Mem/n245 ), .IN1(\Inst_Mem/n242 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n246 ) );
  MUX \Inst_Mem/U251  ( .IN0(\Inst_Mem/n244 ), .IN1(\Inst_Mem/n243 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n245 ) );
  MUX \Inst_Mem/U250  ( .IN0(\Inst_Mem/inst_mem_reg[0][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n244 ) );
  MUX \Inst_Mem/U249  ( .IN0(\Inst_Mem/inst_mem_reg[2][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n243 ) );
  MUX \Inst_Mem/U248  ( .IN0(\Inst_Mem/n241 ), .IN1(\Inst_Mem/n240 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n242 ) );
  MUX \Inst_Mem/U247  ( .IN0(\Inst_Mem/inst_mem_reg[4][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n241 ) );
  MUX \Inst_Mem/U246  ( .IN0(\Inst_Mem/inst_mem_reg[6][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n240 ) );
  MUX \Inst_Mem/U245  ( .IN0(\Inst_Mem/n238 ), .IN1(\Inst_Mem/n235 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n239 ) );
  MUX \Inst_Mem/U244  ( .IN0(\Inst_Mem/n237 ), .IN1(\Inst_Mem/n236 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n238 ) );
  MUX \Inst_Mem/U243  ( .IN0(\Inst_Mem/inst_mem_reg[8][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n237 ) );
  MUX \Inst_Mem/U242  ( .IN0(\Inst_Mem/inst_mem_reg[10][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n236 ) );
  MUX \Inst_Mem/U241  ( .IN0(\Inst_Mem/n234 ), .IN1(\Inst_Mem/n233 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n235 ) );
  MUX \Inst_Mem/U240  ( .IN0(\Inst_Mem/inst_mem_reg[12][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n234 ) );
  MUX \Inst_Mem/U239  ( .IN0(\Inst_Mem/inst_mem_reg[14][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n233 ) );
  MUX \Inst_Mem/U238  ( .IN0(\Inst_Mem/n231 ), .IN1(\Inst_Mem/n224 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n232 ) );
  MUX \Inst_Mem/U237  ( .IN0(\Inst_Mem/n230 ), .IN1(\Inst_Mem/n227 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n231 ) );
  MUX \Inst_Mem/U236  ( .IN0(\Inst_Mem/n229 ), .IN1(\Inst_Mem/n228 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n230 ) );
  MUX \Inst_Mem/U235  ( .IN0(\Inst_Mem/inst_mem_reg[16][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n229 ) );
  MUX \Inst_Mem/U234  ( .IN0(\Inst_Mem/inst_mem_reg[18][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n228 ) );
  MUX \Inst_Mem/U233  ( .IN0(\Inst_Mem/n226 ), .IN1(\Inst_Mem/n225 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n227 ) );
  MUX \Inst_Mem/U232  ( .IN0(\Inst_Mem/inst_mem_reg[20][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n226 ) );
  MUX \Inst_Mem/U231  ( .IN0(\Inst_Mem/inst_mem_reg[22][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n225 ) );
  MUX \Inst_Mem/U230  ( .IN0(\Inst_Mem/n223 ), .IN1(\Inst_Mem/n220 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n224 ) );
  MUX \Inst_Mem/U229  ( .IN0(\Inst_Mem/n222 ), .IN1(\Inst_Mem/n221 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n223 ) );
  MUX \Inst_Mem/U228  ( .IN0(\Inst_Mem/inst_mem_reg[24][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n222 ) );
  MUX \Inst_Mem/U227  ( .IN0(\Inst_Mem/inst_mem_reg[26][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n221 ) );
  MUX \Inst_Mem/U226  ( .IN0(\Inst_Mem/n219 ), .IN1(\Inst_Mem/n218 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n220 ) );
  MUX \Inst_Mem/U225  ( .IN0(\Inst_Mem/inst_mem_reg[28][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n219 ) );
  MUX \Inst_Mem/U224  ( .IN0(\Inst_Mem/inst_mem_reg[30][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n218 ) );
  MUX \Inst_Mem/U223  ( .IN0(\Inst_Mem/n216 ), .IN1(\Inst_Mem/n201 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n217 ) );
  MUX \Inst_Mem/U222  ( .IN0(\Inst_Mem/n215 ), .IN1(\Inst_Mem/n208 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n216 ) );
  MUX \Inst_Mem/U221  ( .IN0(\Inst_Mem/n214 ), .IN1(\Inst_Mem/n211 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n215 ) );
  MUX \Inst_Mem/U220  ( .IN0(\Inst_Mem/n213 ), .IN1(\Inst_Mem/n212 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n214 ) );
  MUX \Inst_Mem/U219  ( .IN0(\Inst_Mem/inst_mem_reg[32][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n213 ) );
  MUX \Inst_Mem/U218  ( .IN0(\Inst_Mem/inst_mem_reg[34][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n212 ) );
  MUX \Inst_Mem/U217  ( .IN0(\Inst_Mem/n210 ), .IN1(\Inst_Mem/n209 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n211 ) );
  MUX \Inst_Mem/U216  ( .IN0(\Inst_Mem/inst_mem_reg[36][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n210 ) );
  MUX \Inst_Mem/U215  ( .IN0(\Inst_Mem/inst_mem_reg[38][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n209 ) );
  MUX \Inst_Mem/U214  ( .IN0(\Inst_Mem/n207 ), .IN1(\Inst_Mem/n204 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n208 ) );
  MUX \Inst_Mem/U213  ( .IN0(\Inst_Mem/n206 ), .IN1(\Inst_Mem/n205 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n207 ) );
  MUX \Inst_Mem/U212  ( .IN0(\Inst_Mem/inst_mem_reg[40][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n206 ) );
  MUX \Inst_Mem/U211  ( .IN0(\Inst_Mem/inst_mem_reg[42][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n205 ) );
  MUX \Inst_Mem/U210  ( .IN0(\Inst_Mem/n203 ), .IN1(\Inst_Mem/n202 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n204 ) );
  MUX \Inst_Mem/U209  ( .IN0(\Inst_Mem/inst_mem_reg[44][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n203 ) );
  MUX \Inst_Mem/U208  ( .IN0(\Inst_Mem/inst_mem_reg[46][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n202 ) );
  MUX \Inst_Mem/U207  ( .IN0(\Inst_Mem/n200 ), .IN1(\Inst_Mem/n193 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n201 ) );
  MUX \Inst_Mem/U206  ( .IN0(\Inst_Mem/n199 ), .IN1(\Inst_Mem/n196 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n200 ) );
  MUX \Inst_Mem/U205  ( .IN0(\Inst_Mem/n198 ), .IN1(\Inst_Mem/n197 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n199 ) );
  MUX \Inst_Mem/U204  ( .IN0(\Inst_Mem/inst_mem_reg[48][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n198 ) );
  MUX \Inst_Mem/U203  ( .IN0(\Inst_Mem/inst_mem_reg[50][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n197 ) );
  MUX \Inst_Mem/U202  ( .IN0(\Inst_Mem/n195 ), .IN1(\Inst_Mem/n194 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n196 ) );
  MUX \Inst_Mem/U201  ( .IN0(\Inst_Mem/inst_mem_reg[52][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n195 ) );
  MUX \Inst_Mem/U200  ( .IN0(\Inst_Mem/inst_mem_reg[54][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n194 ) );
  MUX \Inst_Mem/U199  ( .IN0(\Inst_Mem/n192 ), .IN1(\Inst_Mem/n189 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n193 ) );
  MUX \Inst_Mem/U198  ( .IN0(\Inst_Mem/n191 ), .IN1(\Inst_Mem/n190 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n192 ) );
  MUX \Inst_Mem/U197  ( .IN0(\Inst_Mem/inst_mem_reg[56][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n191 ) );
  MUX \Inst_Mem/U196  ( .IN0(\Inst_Mem/inst_mem_reg[58][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n190 ) );
  MUX \Inst_Mem/U195  ( .IN0(\Inst_Mem/n188 ), .IN1(\Inst_Mem/n187 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n189 ) );
  MUX \Inst_Mem/U194  ( .IN0(\Inst_Mem/inst_mem_reg[60][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n188 ) );
  MUX \Inst_Mem/U193  ( .IN0(\Inst_Mem/inst_mem_reg[62][3] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][3] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n187 ) );
  MUX \Inst_Mem/U192  ( .IN0(\Inst_Mem/n186 ), .IN1(\Inst_Mem/n155 ), .SEL(
        pc_current[7]), .F(imm[2]) );
  MUX \Inst_Mem/U191  ( .IN0(\Inst_Mem/n185 ), .IN1(\Inst_Mem/n170 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n186 ) );
  MUX \Inst_Mem/U190  ( .IN0(\Inst_Mem/n184 ), .IN1(\Inst_Mem/n177 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n185 ) );
  MUX \Inst_Mem/U189  ( .IN0(\Inst_Mem/n183 ), .IN1(\Inst_Mem/n180 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n184 ) );
  MUX \Inst_Mem/U188  ( .IN0(\Inst_Mem/n182 ), .IN1(\Inst_Mem/n181 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n183 ) );
  MUX \Inst_Mem/U187  ( .IN0(\Inst_Mem/inst_mem_reg[0][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n182 ) );
  MUX \Inst_Mem/U186  ( .IN0(\Inst_Mem/inst_mem_reg[2][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n181 ) );
  MUX \Inst_Mem/U185  ( .IN0(\Inst_Mem/n179 ), .IN1(\Inst_Mem/n178 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n180 ) );
  MUX \Inst_Mem/U184  ( .IN0(\Inst_Mem/inst_mem_reg[4][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n179 ) );
  MUX \Inst_Mem/U183  ( .IN0(\Inst_Mem/inst_mem_reg[6][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n178 ) );
  MUX \Inst_Mem/U182  ( .IN0(\Inst_Mem/n176 ), .IN1(\Inst_Mem/n173 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n177 ) );
  MUX \Inst_Mem/U181  ( .IN0(\Inst_Mem/n175 ), .IN1(\Inst_Mem/n174 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n176 ) );
  MUX \Inst_Mem/U180  ( .IN0(\Inst_Mem/inst_mem_reg[8][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n175 ) );
  MUX \Inst_Mem/U179  ( .IN0(\Inst_Mem/inst_mem_reg[10][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n174 ) );
  MUX \Inst_Mem/U178  ( .IN0(\Inst_Mem/n172 ), .IN1(\Inst_Mem/n171 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n173 ) );
  MUX \Inst_Mem/U177  ( .IN0(\Inst_Mem/inst_mem_reg[12][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n172 ) );
  MUX \Inst_Mem/U176  ( .IN0(\Inst_Mem/inst_mem_reg[14][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n171 ) );
  MUX \Inst_Mem/U175  ( .IN0(\Inst_Mem/n169 ), .IN1(\Inst_Mem/n162 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n170 ) );
  MUX \Inst_Mem/U174  ( .IN0(\Inst_Mem/n168 ), .IN1(\Inst_Mem/n165 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n169 ) );
  MUX \Inst_Mem/U173  ( .IN0(\Inst_Mem/n167 ), .IN1(\Inst_Mem/n166 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n168 ) );
  MUX \Inst_Mem/U172  ( .IN0(\Inst_Mem/inst_mem_reg[16][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n167 ) );
  MUX \Inst_Mem/U171  ( .IN0(\Inst_Mem/inst_mem_reg[18][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n166 ) );
  MUX \Inst_Mem/U170  ( .IN0(\Inst_Mem/n164 ), .IN1(\Inst_Mem/n163 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n165 ) );
  MUX \Inst_Mem/U169  ( .IN0(\Inst_Mem/inst_mem_reg[20][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n164 ) );
  MUX \Inst_Mem/U168  ( .IN0(\Inst_Mem/inst_mem_reg[22][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n163 ) );
  MUX \Inst_Mem/U167  ( .IN0(\Inst_Mem/n161 ), .IN1(\Inst_Mem/n158 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n162 ) );
  MUX \Inst_Mem/U166  ( .IN0(\Inst_Mem/n160 ), .IN1(\Inst_Mem/n159 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n161 ) );
  MUX \Inst_Mem/U165  ( .IN0(\Inst_Mem/inst_mem_reg[24][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n160 ) );
  MUX \Inst_Mem/U164  ( .IN0(\Inst_Mem/inst_mem_reg[26][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n159 ) );
  MUX \Inst_Mem/U163  ( .IN0(\Inst_Mem/n157 ), .IN1(\Inst_Mem/n156 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n158 ) );
  MUX \Inst_Mem/U162  ( .IN0(\Inst_Mem/inst_mem_reg[28][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n157 ) );
  MUX \Inst_Mem/U161  ( .IN0(\Inst_Mem/inst_mem_reg[30][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n156 ) );
  MUX \Inst_Mem/U160  ( .IN0(\Inst_Mem/n154 ), .IN1(\Inst_Mem/n139 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n155 ) );
  MUX \Inst_Mem/U159  ( .IN0(\Inst_Mem/n153 ), .IN1(\Inst_Mem/n146 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n154 ) );
  MUX \Inst_Mem/U158  ( .IN0(\Inst_Mem/n152 ), .IN1(\Inst_Mem/n149 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n153 ) );
  MUX \Inst_Mem/U157  ( .IN0(\Inst_Mem/n151 ), .IN1(\Inst_Mem/n150 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n152 ) );
  MUX \Inst_Mem/U156  ( .IN0(\Inst_Mem/inst_mem_reg[32][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n151 ) );
  MUX \Inst_Mem/U155  ( .IN0(\Inst_Mem/inst_mem_reg[34][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n150 ) );
  MUX \Inst_Mem/U154  ( .IN0(\Inst_Mem/n148 ), .IN1(\Inst_Mem/n147 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n149 ) );
  MUX \Inst_Mem/U153  ( .IN0(\Inst_Mem/inst_mem_reg[36][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n148 ) );
  MUX \Inst_Mem/U152  ( .IN0(\Inst_Mem/inst_mem_reg[38][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n147 ) );
  MUX \Inst_Mem/U151  ( .IN0(\Inst_Mem/n145 ), .IN1(\Inst_Mem/n142 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n146 ) );
  MUX \Inst_Mem/U150  ( .IN0(\Inst_Mem/n144 ), .IN1(\Inst_Mem/n143 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n145 ) );
  MUX \Inst_Mem/U149  ( .IN0(\Inst_Mem/inst_mem_reg[40][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n144 ) );
  MUX \Inst_Mem/U148  ( .IN0(\Inst_Mem/inst_mem_reg[42][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n143 ) );
  MUX \Inst_Mem/U147  ( .IN0(\Inst_Mem/n141 ), .IN1(\Inst_Mem/n140 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n142 ) );
  MUX \Inst_Mem/U146  ( .IN0(\Inst_Mem/inst_mem_reg[44][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n141 ) );
  MUX \Inst_Mem/U145  ( .IN0(\Inst_Mem/inst_mem_reg[46][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n140 ) );
  MUX \Inst_Mem/U144  ( .IN0(\Inst_Mem/n138 ), .IN1(\Inst_Mem/n131 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n139 ) );
  MUX \Inst_Mem/U143  ( .IN0(\Inst_Mem/n137 ), .IN1(\Inst_Mem/n134 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n138 ) );
  MUX \Inst_Mem/U142  ( .IN0(\Inst_Mem/n136 ), .IN1(\Inst_Mem/n135 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n137 ) );
  MUX \Inst_Mem/U141  ( .IN0(\Inst_Mem/inst_mem_reg[48][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n136 ) );
  MUX \Inst_Mem/U140  ( .IN0(\Inst_Mem/inst_mem_reg[50][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n135 ) );
  MUX \Inst_Mem/U139  ( .IN0(\Inst_Mem/n133 ), .IN1(\Inst_Mem/n132 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n134 ) );
  MUX \Inst_Mem/U138  ( .IN0(\Inst_Mem/inst_mem_reg[52][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n133 ) );
  MUX \Inst_Mem/U137  ( .IN0(\Inst_Mem/inst_mem_reg[54][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n132 ) );
  MUX \Inst_Mem/U136  ( .IN0(\Inst_Mem/n130 ), .IN1(\Inst_Mem/n127 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n131 ) );
  MUX \Inst_Mem/U135  ( .IN0(\Inst_Mem/n129 ), .IN1(\Inst_Mem/n128 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n130 ) );
  MUX \Inst_Mem/U134  ( .IN0(\Inst_Mem/inst_mem_reg[56][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n129 ) );
  MUX \Inst_Mem/U133  ( .IN0(\Inst_Mem/inst_mem_reg[58][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n128 ) );
  MUX \Inst_Mem/U132  ( .IN0(\Inst_Mem/n126 ), .IN1(\Inst_Mem/n125 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n127 ) );
  MUX \Inst_Mem/U131  ( .IN0(\Inst_Mem/inst_mem_reg[60][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n126 ) );
  MUX \Inst_Mem/U130  ( .IN0(\Inst_Mem/inst_mem_reg[62][2] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][2] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n125 ) );
  MUX \Inst_Mem/U129  ( .IN0(\Inst_Mem/n124 ), .IN1(\Inst_Mem/n93 ), .SEL(
        pc_current[7]), .F(imm[1]) );
  MUX \Inst_Mem/U128  ( .IN0(\Inst_Mem/n123 ), .IN1(\Inst_Mem/n108 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n124 ) );
  MUX \Inst_Mem/U127  ( .IN0(\Inst_Mem/n122 ), .IN1(\Inst_Mem/n115 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n123 ) );
  MUX \Inst_Mem/U126  ( .IN0(\Inst_Mem/n121 ), .IN1(\Inst_Mem/n118 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n122 ) );
  MUX \Inst_Mem/U125  ( .IN0(\Inst_Mem/n120 ), .IN1(\Inst_Mem/n119 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n121 ) );
  MUX \Inst_Mem/U124  ( .IN0(\Inst_Mem/inst_mem_reg[0][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n120 ) );
  MUX \Inst_Mem/U123  ( .IN0(\Inst_Mem/inst_mem_reg[2][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n119 ) );
  MUX \Inst_Mem/U122  ( .IN0(\Inst_Mem/n117 ), .IN1(\Inst_Mem/n116 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n118 ) );
  MUX \Inst_Mem/U121  ( .IN0(\Inst_Mem/inst_mem_reg[4][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n117 ) );
  MUX \Inst_Mem/U120  ( .IN0(\Inst_Mem/inst_mem_reg[6][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n116 ) );
  MUX \Inst_Mem/U119  ( .IN0(\Inst_Mem/n114 ), .IN1(\Inst_Mem/n111 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n115 ) );
  MUX \Inst_Mem/U118  ( .IN0(\Inst_Mem/n113 ), .IN1(\Inst_Mem/n112 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n114 ) );
  MUX \Inst_Mem/U117  ( .IN0(\Inst_Mem/inst_mem_reg[8][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n113 ) );
  MUX \Inst_Mem/U116  ( .IN0(\Inst_Mem/inst_mem_reg[10][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n112 ) );
  MUX \Inst_Mem/U115  ( .IN0(\Inst_Mem/n110 ), .IN1(\Inst_Mem/n109 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n111 ) );
  MUX \Inst_Mem/U114  ( .IN0(\Inst_Mem/inst_mem_reg[12][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n110 ) );
  MUX \Inst_Mem/U113  ( .IN0(\Inst_Mem/inst_mem_reg[14][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n109 ) );
  MUX \Inst_Mem/U112  ( .IN0(\Inst_Mem/n107 ), .IN1(\Inst_Mem/n100 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n108 ) );
  MUX \Inst_Mem/U111  ( .IN0(\Inst_Mem/n106 ), .IN1(\Inst_Mem/n103 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n107 ) );
  MUX \Inst_Mem/U110  ( .IN0(\Inst_Mem/n105 ), .IN1(\Inst_Mem/n104 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n106 ) );
  MUX \Inst_Mem/U109  ( .IN0(\Inst_Mem/inst_mem_reg[16][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n105 ) );
  MUX \Inst_Mem/U108  ( .IN0(\Inst_Mem/inst_mem_reg[18][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n104 ) );
  MUX \Inst_Mem/U107  ( .IN0(\Inst_Mem/n102 ), .IN1(\Inst_Mem/n101 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n103 ) );
  MUX \Inst_Mem/U106  ( .IN0(\Inst_Mem/inst_mem_reg[20][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n102 ) );
  MUX \Inst_Mem/U105  ( .IN0(\Inst_Mem/inst_mem_reg[22][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n101 ) );
  MUX \Inst_Mem/U104  ( .IN0(\Inst_Mem/n99 ), .IN1(\Inst_Mem/n96 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n100 ) );
  MUX \Inst_Mem/U103  ( .IN0(\Inst_Mem/n98 ), .IN1(\Inst_Mem/n97 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n99 ) );
  MUX \Inst_Mem/U102  ( .IN0(\Inst_Mem/inst_mem_reg[24][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n98 ) );
  MUX \Inst_Mem/U101  ( .IN0(\Inst_Mem/inst_mem_reg[26][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n97 ) );
  MUX \Inst_Mem/U100  ( .IN0(\Inst_Mem/n95 ), .IN1(\Inst_Mem/n94 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n96 ) );
  MUX \Inst_Mem/U99  ( .IN0(\Inst_Mem/inst_mem_reg[28][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n95 ) );
  MUX \Inst_Mem/U98  ( .IN0(\Inst_Mem/inst_mem_reg[30][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n94 ) );
  MUX \Inst_Mem/U97  ( .IN0(\Inst_Mem/n92 ), .IN1(\Inst_Mem/n77 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n93 ) );
  MUX \Inst_Mem/U96  ( .IN0(\Inst_Mem/n91 ), .IN1(\Inst_Mem/n84 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n92 ) );
  MUX \Inst_Mem/U95  ( .IN0(\Inst_Mem/n90 ), .IN1(\Inst_Mem/n87 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n91 ) );
  MUX \Inst_Mem/U94  ( .IN0(\Inst_Mem/n89 ), .IN1(\Inst_Mem/n88 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n90 ) );
  MUX \Inst_Mem/U93  ( .IN0(\Inst_Mem/inst_mem_reg[32][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n89 ) );
  MUX \Inst_Mem/U92  ( .IN0(\Inst_Mem/inst_mem_reg[34][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n88 ) );
  MUX \Inst_Mem/U91  ( .IN0(\Inst_Mem/n86 ), .IN1(\Inst_Mem/n85 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n87 ) );
  MUX \Inst_Mem/U90  ( .IN0(\Inst_Mem/inst_mem_reg[36][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n86 ) );
  MUX \Inst_Mem/U89  ( .IN0(\Inst_Mem/inst_mem_reg[38][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n85 ) );
  MUX \Inst_Mem/U88  ( .IN0(\Inst_Mem/n83 ), .IN1(\Inst_Mem/n80 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n84 ) );
  MUX \Inst_Mem/U87  ( .IN0(\Inst_Mem/n82 ), .IN1(\Inst_Mem/n81 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n83 ) );
  MUX \Inst_Mem/U86  ( .IN0(\Inst_Mem/inst_mem_reg[40][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n82 ) );
  MUX \Inst_Mem/U85  ( .IN0(\Inst_Mem/inst_mem_reg[42][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n81 ) );
  MUX \Inst_Mem/U84  ( .IN0(\Inst_Mem/n79 ), .IN1(\Inst_Mem/n78 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n80 ) );
  MUX \Inst_Mem/U83  ( .IN0(\Inst_Mem/inst_mem_reg[44][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n79 ) );
  MUX \Inst_Mem/U82  ( .IN0(\Inst_Mem/inst_mem_reg[46][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n78 ) );
  MUX \Inst_Mem/U81  ( .IN0(\Inst_Mem/n76 ), .IN1(\Inst_Mem/n69 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n77 ) );
  MUX \Inst_Mem/U80  ( .IN0(\Inst_Mem/n75 ), .IN1(\Inst_Mem/n72 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n76 ) );
  MUX \Inst_Mem/U79  ( .IN0(\Inst_Mem/n74 ), .IN1(\Inst_Mem/n73 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n75 ) );
  MUX \Inst_Mem/U78  ( .IN0(\Inst_Mem/inst_mem_reg[48][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n74 ) );
  MUX \Inst_Mem/U77  ( .IN0(\Inst_Mem/inst_mem_reg[50][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n73 ) );
  MUX \Inst_Mem/U76  ( .IN0(\Inst_Mem/n71 ), .IN1(\Inst_Mem/n70 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n72 ) );
  MUX \Inst_Mem/U75  ( .IN0(\Inst_Mem/inst_mem_reg[52][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n71 ) );
  MUX \Inst_Mem/U74  ( .IN0(\Inst_Mem/inst_mem_reg[54][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n70 ) );
  MUX \Inst_Mem/U73  ( .IN0(\Inst_Mem/n68 ), .IN1(\Inst_Mem/n65 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n69 ) );
  MUX \Inst_Mem/U72  ( .IN0(\Inst_Mem/n67 ), .IN1(\Inst_Mem/n66 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n68 ) );
  MUX \Inst_Mem/U71  ( .IN0(\Inst_Mem/inst_mem_reg[56][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n67 ) );
  MUX \Inst_Mem/U70  ( .IN0(\Inst_Mem/inst_mem_reg[58][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n66 ) );
  MUX \Inst_Mem/U69  ( .IN0(\Inst_Mem/n64 ), .IN1(\Inst_Mem/n63 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n65 ) );
  MUX \Inst_Mem/U68  ( .IN0(\Inst_Mem/inst_mem_reg[60][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n64 ) );
  MUX \Inst_Mem/U67  ( .IN0(\Inst_Mem/inst_mem_reg[62][1] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][1] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n63 ) );
  MUX \Inst_Mem/U66  ( .IN0(\Inst_Mem/n62 ), .IN1(\Inst_Mem/n31 ), .SEL(
        pc_current[7]), .F(imm[0]) );
  MUX \Inst_Mem/U65  ( .IN0(\Inst_Mem/n61 ), .IN1(\Inst_Mem/n46 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n62 ) );
  MUX \Inst_Mem/U64  ( .IN0(\Inst_Mem/n60 ), .IN1(\Inst_Mem/n53 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n61 ) );
  MUX \Inst_Mem/U63  ( .IN0(\Inst_Mem/n59 ), .IN1(\Inst_Mem/n56 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n60 ) );
  MUX \Inst_Mem/U62  ( .IN0(\Inst_Mem/n58 ), .IN1(\Inst_Mem/n57 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n59 ) );
  MUX \Inst_Mem/U61  ( .IN0(\Inst_Mem/inst_mem_reg[0][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[1][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n58 ) );
  MUX \Inst_Mem/U60  ( .IN0(\Inst_Mem/inst_mem_reg[2][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[3][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n57 ) );
  MUX \Inst_Mem/U59  ( .IN0(\Inst_Mem/n55 ), .IN1(\Inst_Mem/n54 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n56 ) );
  MUX \Inst_Mem/U58  ( .IN0(\Inst_Mem/inst_mem_reg[4][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[5][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n55 ) );
  MUX \Inst_Mem/U57  ( .IN0(\Inst_Mem/inst_mem_reg[6][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[7][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n54 ) );
  MUX \Inst_Mem/U56  ( .IN0(\Inst_Mem/n52 ), .IN1(\Inst_Mem/n49 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n53 ) );
  MUX \Inst_Mem/U55  ( .IN0(\Inst_Mem/n51 ), .IN1(\Inst_Mem/n50 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n52 ) );
  MUX \Inst_Mem/U54  ( .IN0(\Inst_Mem/inst_mem_reg[8][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[9][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n51 ) );
  MUX \Inst_Mem/U53  ( .IN0(\Inst_Mem/inst_mem_reg[10][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[11][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n50 ) );
  MUX \Inst_Mem/U52  ( .IN0(\Inst_Mem/n48 ), .IN1(\Inst_Mem/n47 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n49 ) );
  MUX \Inst_Mem/U51  ( .IN0(\Inst_Mem/inst_mem_reg[12][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[13][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n48 ) );
  MUX \Inst_Mem/U50  ( .IN0(\Inst_Mem/inst_mem_reg[14][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[15][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n47 ) );
  MUX \Inst_Mem/U49  ( .IN0(\Inst_Mem/n45 ), .IN1(\Inst_Mem/n38 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n46 ) );
  MUX \Inst_Mem/U48  ( .IN0(\Inst_Mem/n44 ), .IN1(\Inst_Mem/n41 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n45 ) );
  MUX \Inst_Mem/U47  ( .IN0(\Inst_Mem/n43 ), .IN1(\Inst_Mem/n42 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n44 ) );
  MUX \Inst_Mem/U46  ( .IN0(\Inst_Mem/inst_mem_reg[16][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[17][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n43 ) );
  MUX \Inst_Mem/U45  ( .IN0(\Inst_Mem/inst_mem_reg[18][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[19][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n42 ) );
  MUX \Inst_Mem/U44  ( .IN0(\Inst_Mem/n40 ), .IN1(\Inst_Mem/n39 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n41 ) );
  MUX \Inst_Mem/U43  ( .IN0(\Inst_Mem/inst_mem_reg[20][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[21][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n40 ) );
  MUX \Inst_Mem/U42  ( .IN0(\Inst_Mem/inst_mem_reg[22][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[23][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n39 ) );
  MUX \Inst_Mem/U41  ( .IN0(\Inst_Mem/n37 ), .IN1(\Inst_Mem/n34 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n38 ) );
  MUX \Inst_Mem/U40  ( .IN0(\Inst_Mem/n36 ), .IN1(\Inst_Mem/n35 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n37 ) );
  MUX \Inst_Mem/U39  ( .IN0(\Inst_Mem/inst_mem_reg[24][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[25][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n36 ) );
  MUX \Inst_Mem/U38  ( .IN0(\Inst_Mem/inst_mem_reg[26][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[27][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n35 ) );
  MUX \Inst_Mem/U37  ( .IN0(\Inst_Mem/n33 ), .IN1(\Inst_Mem/n32 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n34 ) );
  MUX \Inst_Mem/U36  ( .IN0(\Inst_Mem/inst_mem_reg[28][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[29][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n33 ) );
  MUX \Inst_Mem/U35  ( .IN0(\Inst_Mem/inst_mem_reg[30][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[31][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n32 ) );
  MUX \Inst_Mem/U34  ( .IN0(\Inst_Mem/n30 ), .IN1(\Inst_Mem/n15 ), .SEL(
        pc_current[6]), .F(\Inst_Mem/n31 ) );
  MUX \Inst_Mem/U33  ( .IN0(\Inst_Mem/n29 ), .IN1(\Inst_Mem/n22 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n30 ) );
  MUX \Inst_Mem/U32  ( .IN0(\Inst_Mem/n28 ), .IN1(\Inst_Mem/n25 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n29 ) );
  MUX \Inst_Mem/U31  ( .IN0(\Inst_Mem/n27 ), .IN1(\Inst_Mem/n26 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n28 ) );
  MUX \Inst_Mem/U30  ( .IN0(\Inst_Mem/inst_mem_reg[32][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[33][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n27 ) );
  MUX \Inst_Mem/U29  ( .IN0(\Inst_Mem/inst_mem_reg[34][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[35][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n26 ) );
  MUX \Inst_Mem/U28  ( .IN0(\Inst_Mem/n24 ), .IN1(\Inst_Mem/n23 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n25 ) );
  MUX \Inst_Mem/U27  ( .IN0(\Inst_Mem/inst_mem_reg[36][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[37][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n24 ) );
  MUX \Inst_Mem/U26  ( .IN0(\Inst_Mem/inst_mem_reg[38][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[39][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n23 ) );
  MUX \Inst_Mem/U25  ( .IN0(\Inst_Mem/n21 ), .IN1(\Inst_Mem/n18 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n22 ) );
  MUX \Inst_Mem/U24  ( .IN0(\Inst_Mem/n20 ), .IN1(\Inst_Mem/n19 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n21 ) );
  MUX \Inst_Mem/U23  ( .IN0(\Inst_Mem/inst_mem_reg[40][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[41][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n20 ) );
  MUX \Inst_Mem/U22  ( .IN0(\Inst_Mem/inst_mem_reg[42][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[43][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n19 ) );
  MUX \Inst_Mem/U21  ( .IN0(\Inst_Mem/n17 ), .IN1(\Inst_Mem/n16 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n18 ) );
  MUX \Inst_Mem/U20  ( .IN0(\Inst_Mem/inst_mem_reg[44][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[45][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n17 ) );
  MUX \Inst_Mem/U19  ( .IN0(\Inst_Mem/inst_mem_reg[46][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[47][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n16 ) );
  MUX \Inst_Mem/U18  ( .IN0(\Inst_Mem/n14 ), .IN1(\Inst_Mem/n7 ), .SEL(
        pc_current[5]), .F(\Inst_Mem/n15 ) );
  MUX \Inst_Mem/U17  ( .IN0(\Inst_Mem/n13 ), .IN1(\Inst_Mem/n10 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n14 ) );
  MUX \Inst_Mem/U16  ( .IN0(\Inst_Mem/n12 ), .IN1(\Inst_Mem/n11 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n13 ) );
  MUX \Inst_Mem/U15  ( .IN0(\Inst_Mem/inst_mem_reg[48][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[49][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n12 ) );
  MUX \Inst_Mem/U14  ( .IN0(\Inst_Mem/inst_mem_reg[50][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[51][0] ), .SEL(pc_current[2]), .F(
        \Inst_Mem/n11 ) );
  MUX \Inst_Mem/U13  ( .IN0(\Inst_Mem/n9 ), .IN1(\Inst_Mem/n8 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n10 ) );
  MUX \Inst_Mem/U12  ( .IN0(\Inst_Mem/inst_mem_reg[52][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[53][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n9 ) );
  MUX \Inst_Mem/U11  ( .IN0(\Inst_Mem/inst_mem_reg[54][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[55][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n8 ) );
  MUX \Inst_Mem/U10  ( .IN0(\Inst_Mem/n6 ), .IN1(\Inst_Mem/n3 ), .SEL(
        pc_current[4]), .F(\Inst_Mem/n7 ) );
  MUX \Inst_Mem/U9  ( .IN0(\Inst_Mem/n5 ), .IN1(\Inst_Mem/n4 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n6 ) );
  MUX \Inst_Mem/U8  ( .IN0(\Inst_Mem/inst_mem_reg[56][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[57][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n5 ) );
  MUX \Inst_Mem/U7  ( .IN0(\Inst_Mem/inst_mem_reg[58][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[59][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n4 ) );
  MUX \Inst_Mem/U6  ( .IN0(\Inst_Mem/n2 ), .IN1(\Inst_Mem/n1 ), .SEL(
        pc_current[3]), .F(\Inst_Mem/n3 ) );
  MUX \Inst_Mem/U5  ( .IN0(\Inst_Mem/inst_mem_reg[60][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[61][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n2 ) );
  MUX \Inst_Mem/U4  ( .IN0(\Inst_Mem/inst_mem_reg[62][0] ), .IN1(
        \Inst_Mem/inst_mem_reg[63][0] ), .SEL(pc_current[2]), .F(\Inst_Mem/n1 ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][0]  ( .D(\Inst_Mem/inst_mem_reg[63][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[2016]), .Q(
        \Inst_Mem/inst_mem_reg[63][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][1]  ( .D(\Inst_Mem/inst_mem_reg[63][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[2017]), .Q(
        \Inst_Mem/inst_mem_reg[63][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][2]  ( .D(\Inst_Mem/inst_mem_reg[63][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[2018]), .Q(
        \Inst_Mem/inst_mem_reg[63][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][3]  ( .D(\Inst_Mem/inst_mem_reg[63][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[2019]), .Q(
        \Inst_Mem/inst_mem_reg[63][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][4]  ( .D(\Inst_Mem/inst_mem_reg[63][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[2020]), .Q(
        \Inst_Mem/inst_mem_reg[63][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][5]  ( .D(\Inst_Mem/inst_mem_reg[63][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[2021]), .Q(
        \Inst_Mem/inst_mem_reg[63][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][6]  ( .D(\Inst_Mem/inst_mem_reg[63][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[2022]), .Q(
        \Inst_Mem/inst_mem_reg[63][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][7]  ( .D(\Inst_Mem/inst_mem_reg[63][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[2023]), .Q(
        \Inst_Mem/inst_mem_reg[63][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][8]  ( .D(\Inst_Mem/inst_mem_reg[63][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[2024]), .Q(
        \Inst_Mem/inst_mem_reg[63][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][9]  ( .D(\Inst_Mem/inst_mem_reg[63][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[2025]), .Q(
        \Inst_Mem/inst_mem_reg[63][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[63][10]  ( .D(\Inst_Mem/inst_mem_reg[63][10] ), .CLK(clk), .RST(rst), .I(g_init[2026]), .Q(\Inst_Mem/inst_mem_reg[63][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][11]  ( .D(\Inst_Mem/inst_mem_reg[63][11] ), .CLK(clk), .RST(rst), .I(g_init[2027]), .Q(\Inst_Mem/inst_mem_reg[63][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][12]  ( .D(\Inst_Mem/inst_mem_reg[63][12] ), .CLK(clk), .RST(rst), .I(g_init[2028]), .Q(\Inst_Mem/inst_mem_reg[63][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][13]  ( .D(\Inst_Mem/inst_mem_reg[63][13] ), .CLK(clk), .RST(rst), .I(g_init[2029]), .Q(\Inst_Mem/inst_mem_reg[63][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][14]  ( .D(\Inst_Mem/inst_mem_reg[63][14] ), .CLK(clk), .RST(rst), .I(g_init[2030]), .Q(\Inst_Mem/inst_mem_reg[63][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][15]  ( .D(\Inst_Mem/inst_mem_reg[63][15] ), .CLK(clk), .RST(rst), .I(g_init[2031]), .Q(\Inst_Mem/inst_mem_reg[63][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][16]  ( .D(\Inst_Mem/inst_mem_reg[63][16] ), .CLK(clk), .RST(rst), .I(g_init[2032]), .Q(\Inst_Mem/inst_mem_reg[63][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][17]  ( .D(\Inst_Mem/inst_mem_reg[63][17] ), .CLK(clk), .RST(rst), .I(g_init[2033]), .Q(\Inst_Mem/inst_mem_reg[63][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][18]  ( .D(\Inst_Mem/inst_mem_reg[63][18] ), .CLK(clk), .RST(rst), .I(g_init[2034]), .Q(\Inst_Mem/inst_mem_reg[63][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][19]  ( .D(\Inst_Mem/inst_mem_reg[63][19] ), .CLK(clk), .RST(rst), .I(g_init[2035]), .Q(\Inst_Mem/inst_mem_reg[63][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][20]  ( .D(\Inst_Mem/inst_mem_reg[63][20] ), .CLK(clk), .RST(rst), .I(g_init[2036]), .Q(\Inst_Mem/inst_mem_reg[63][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][21]  ( .D(\Inst_Mem/inst_mem_reg[63][21] ), .CLK(clk), .RST(rst), .I(g_init[2037]), .Q(\Inst_Mem/inst_mem_reg[63][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][22]  ( .D(\Inst_Mem/inst_mem_reg[63][22] ), .CLK(clk), .RST(rst), .I(g_init[2038]), .Q(\Inst_Mem/inst_mem_reg[63][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][23]  ( .D(\Inst_Mem/inst_mem_reg[63][23] ), .CLK(clk), .RST(rst), .I(g_init[2039]), .Q(\Inst_Mem/inst_mem_reg[63][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][24]  ( .D(\Inst_Mem/inst_mem_reg[63][24] ), .CLK(clk), .RST(rst), .I(g_init[2040]), .Q(\Inst_Mem/inst_mem_reg[63][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][25]  ( .D(\Inst_Mem/inst_mem_reg[63][25] ), .CLK(clk), .RST(rst), .I(g_init[2041]), .Q(\Inst_Mem/inst_mem_reg[63][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][26]  ( .D(\Inst_Mem/inst_mem_reg[63][26] ), .CLK(clk), .RST(rst), .I(g_init[2042]), .Q(\Inst_Mem/inst_mem_reg[63][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][27]  ( .D(\Inst_Mem/inst_mem_reg[63][27] ), .CLK(clk), .RST(rst), .I(g_init[2043]), .Q(\Inst_Mem/inst_mem_reg[63][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][28]  ( .D(\Inst_Mem/inst_mem_reg[63][28] ), .CLK(clk), .RST(rst), .I(g_init[2044]), .Q(\Inst_Mem/inst_mem_reg[63][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][29]  ( .D(\Inst_Mem/inst_mem_reg[63][29] ), .CLK(clk), .RST(rst), .I(g_init[2045]), .Q(\Inst_Mem/inst_mem_reg[63][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][30]  ( .D(\Inst_Mem/inst_mem_reg[63][30] ), .CLK(clk), .RST(rst), .I(g_init[2046]), .Q(\Inst_Mem/inst_mem_reg[63][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[63][31]  ( .D(\Inst_Mem/inst_mem_reg[63][31] ), .CLK(clk), .RST(rst), .I(g_init[2047]), .Q(\Inst_Mem/inst_mem_reg[63][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][0]  ( .D(\Inst_Mem/inst_mem_reg[62][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1984]), .Q(
        \Inst_Mem/inst_mem_reg[62][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][1]  ( .D(\Inst_Mem/inst_mem_reg[62][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1985]), .Q(
        \Inst_Mem/inst_mem_reg[62][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][2]  ( .D(\Inst_Mem/inst_mem_reg[62][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1986]), .Q(
        \Inst_Mem/inst_mem_reg[62][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][3]  ( .D(\Inst_Mem/inst_mem_reg[62][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1987]), .Q(
        \Inst_Mem/inst_mem_reg[62][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][4]  ( .D(\Inst_Mem/inst_mem_reg[62][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1988]), .Q(
        \Inst_Mem/inst_mem_reg[62][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][5]  ( .D(\Inst_Mem/inst_mem_reg[62][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1989]), .Q(
        \Inst_Mem/inst_mem_reg[62][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][6]  ( .D(\Inst_Mem/inst_mem_reg[62][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1990]), .Q(
        \Inst_Mem/inst_mem_reg[62][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][7]  ( .D(\Inst_Mem/inst_mem_reg[62][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1991]), .Q(
        \Inst_Mem/inst_mem_reg[62][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][8]  ( .D(\Inst_Mem/inst_mem_reg[62][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1992]), .Q(
        \Inst_Mem/inst_mem_reg[62][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][9]  ( .D(\Inst_Mem/inst_mem_reg[62][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1993]), .Q(
        \Inst_Mem/inst_mem_reg[62][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[62][10]  ( .D(\Inst_Mem/inst_mem_reg[62][10] ), .CLK(clk), .RST(rst), .I(g_init[1994]), .Q(\Inst_Mem/inst_mem_reg[62][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][11]  ( .D(\Inst_Mem/inst_mem_reg[62][11] ), .CLK(clk), .RST(rst), .I(g_init[1995]), .Q(\Inst_Mem/inst_mem_reg[62][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][12]  ( .D(\Inst_Mem/inst_mem_reg[62][12] ), .CLK(clk), .RST(rst), .I(g_init[1996]), .Q(\Inst_Mem/inst_mem_reg[62][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][13]  ( .D(\Inst_Mem/inst_mem_reg[62][13] ), .CLK(clk), .RST(rst), .I(g_init[1997]), .Q(\Inst_Mem/inst_mem_reg[62][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][14]  ( .D(\Inst_Mem/inst_mem_reg[62][14] ), .CLK(clk), .RST(rst), .I(g_init[1998]), .Q(\Inst_Mem/inst_mem_reg[62][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][15]  ( .D(\Inst_Mem/inst_mem_reg[62][15] ), .CLK(clk), .RST(rst), .I(g_init[1999]), .Q(\Inst_Mem/inst_mem_reg[62][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][16]  ( .D(\Inst_Mem/inst_mem_reg[62][16] ), .CLK(clk), .RST(rst), .I(g_init[2000]), .Q(\Inst_Mem/inst_mem_reg[62][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][17]  ( .D(\Inst_Mem/inst_mem_reg[62][17] ), .CLK(clk), .RST(rst), .I(g_init[2001]), .Q(\Inst_Mem/inst_mem_reg[62][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][18]  ( .D(\Inst_Mem/inst_mem_reg[62][18] ), .CLK(clk), .RST(rst), .I(g_init[2002]), .Q(\Inst_Mem/inst_mem_reg[62][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][19]  ( .D(\Inst_Mem/inst_mem_reg[62][19] ), .CLK(clk), .RST(rst), .I(g_init[2003]), .Q(\Inst_Mem/inst_mem_reg[62][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][20]  ( .D(\Inst_Mem/inst_mem_reg[62][20] ), .CLK(clk), .RST(rst), .I(g_init[2004]), .Q(\Inst_Mem/inst_mem_reg[62][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][21]  ( .D(\Inst_Mem/inst_mem_reg[62][21] ), .CLK(clk), .RST(rst), .I(g_init[2005]), .Q(\Inst_Mem/inst_mem_reg[62][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][22]  ( .D(\Inst_Mem/inst_mem_reg[62][22] ), .CLK(clk), .RST(rst), .I(g_init[2006]), .Q(\Inst_Mem/inst_mem_reg[62][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][23]  ( .D(\Inst_Mem/inst_mem_reg[62][23] ), .CLK(clk), .RST(rst), .I(g_init[2007]), .Q(\Inst_Mem/inst_mem_reg[62][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][24]  ( .D(\Inst_Mem/inst_mem_reg[62][24] ), .CLK(clk), .RST(rst), .I(g_init[2008]), .Q(\Inst_Mem/inst_mem_reg[62][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][25]  ( .D(\Inst_Mem/inst_mem_reg[62][25] ), .CLK(clk), .RST(rst), .I(g_init[2009]), .Q(\Inst_Mem/inst_mem_reg[62][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][26]  ( .D(\Inst_Mem/inst_mem_reg[62][26] ), .CLK(clk), .RST(rst), .I(g_init[2010]), .Q(\Inst_Mem/inst_mem_reg[62][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][27]  ( .D(\Inst_Mem/inst_mem_reg[62][27] ), .CLK(clk), .RST(rst), .I(g_init[2011]), .Q(\Inst_Mem/inst_mem_reg[62][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][28]  ( .D(\Inst_Mem/inst_mem_reg[62][28] ), .CLK(clk), .RST(rst), .I(g_init[2012]), .Q(\Inst_Mem/inst_mem_reg[62][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][29]  ( .D(\Inst_Mem/inst_mem_reg[62][29] ), .CLK(clk), .RST(rst), .I(g_init[2013]), .Q(\Inst_Mem/inst_mem_reg[62][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][30]  ( .D(\Inst_Mem/inst_mem_reg[62][30] ), .CLK(clk), .RST(rst), .I(g_init[2014]), .Q(\Inst_Mem/inst_mem_reg[62][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[62][31]  ( .D(\Inst_Mem/inst_mem_reg[62][31] ), .CLK(clk), .RST(rst), .I(g_init[2015]), .Q(\Inst_Mem/inst_mem_reg[62][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][0]  ( .D(\Inst_Mem/inst_mem_reg[61][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1952]), .Q(
        \Inst_Mem/inst_mem_reg[61][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][1]  ( .D(\Inst_Mem/inst_mem_reg[61][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1953]), .Q(
        \Inst_Mem/inst_mem_reg[61][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][2]  ( .D(\Inst_Mem/inst_mem_reg[61][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1954]), .Q(
        \Inst_Mem/inst_mem_reg[61][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][3]  ( .D(\Inst_Mem/inst_mem_reg[61][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1955]), .Q(
        \Inst_Mem/inst_mem_reg[61][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][4]  ( .D(\Inst_Mem/inst_mem_reg[61][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1956]), .Q(
        \Inst_Mem/inst_mem_reg[61][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][5]  ( .D(\Inst_Mem/inst_mem_reg[61][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1957]), .Q(
        \Inst_Mem/inst_mem_reg[61][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][6]  ( .D(\Inst_Mem/inst_mem_reg[61][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1958]), .Q(
        \Inst_Mem/inst_mem_reg[61][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][7]  ( .D(\Inst_Mem/inst_mem_reg[61][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1959]), .Q(
        \Inst_Mem/inst_mem_reg[61][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][8]  ( .D(\Inst_Mem/inst_mem_reg[61][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1960]), .Q(
        \Inst_Mem/inst_mem_reg[61][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][9]  ( .D(\Inst_Mem/inst_mem_reg[61][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1961]), .Q(
        \Inst_Mem/inst_mem_reg[61][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[61][10]  ( .D(\Inst_Mem/inst_mem_reg[61][10] ), .CLK(clk), .RST(rst), .I(g_init[1962]), .Q(\Inst_Mem/inst_mem_reg[61][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][11]  ( .D(\Inst_Mem/inst_mem_reg[61][11] ), .CLK(clk), .RST(rst), .I(g_init[1963]), .Q(\Inst_Mem/inst_mem_reg[61][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][12]  ( .D(\Inst_Mem/inst_mem_reg[61][12] ), .CLK(clk), .RST(rst), .I(g_init[1964]), .Q(\Inst_Mem/inst_mem_reg[61][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][13]  ( .D(\Inst_Mem/inst_mem_reg[61][13] ), .CLK(clk), .RST(rst), .I(g_init[1965]), .Q(\Inst_Mem/inst_mem_reg[61][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][14]  ( .D(\Inst_Mem/inst_mem_reg[61][14] ), .CLK(clk), .RST(rst), .I(g_init[1966]), .Q(\Inst_Mem/inst_mem_reg[61][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][15]  ( .D(\Inst_Mem/inst_mem_reg[61][15] ), .CLK(clk), .RST(rst), .I(g_init[1967]), .Q(\Inst_Mem/inst_mem_reg[61][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][16]  ( .D(\Inst_Mem/inst_mem_reg[61][16] ), .CLK(clk), .RST(rst), .I(g_init[1968]), .Q(\Inst_Mem/inst_mem_reg[61][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][17]  ( .D(\Inst_Mem/inst_mem_reg[61][17] ), .CLK(clk), .RST(rst), .I(g_init[1969]), .Q(\Inst_Mem/inst_mem_reg[61][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][18]  ( .D(\Inst_Mem/inst_mem_reg[61][18] ), .CLK(clk), .RST(rst), .I(g_init[1970]), .Q(\Inst_Mem/inst_mem_reg[61][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][19]  ( .D(\Inst_Mem/inst_mem_reg[61][19] ), .CLK(clk), .RST(rst), .I(g_init[1971]), .Q(\Inst_Mem/inst_mem_reg[61][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][20]  ( .D(\Inst_Mem/inst_mem_reg[61][20] ), .CLK(clk), .RST(rst), .I(g_init[1972]), .Q(\Inst_Mem/inst_mem_reg[61][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][21]  ( .D(\Inst_Mem/inst_mem_reg[61][21] ), .CLK(clk), .RST(rst), .I(g_init[1973]), .Q(\Inst_Mem/inst_mem_reg[61][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][22]  ( .D(\Inst_Mem/inst_mem_reg[61][22] ), .CLK(clk), .RST(rst), .I(g_init[1974]), .Q(\Inst_Mem/inst_mem_reg[61][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][23]  ( .D(\Inst_Mem/inst_mem_reg[61][23] ), .CLK(clk), .RST(rst), .I(g_init[1975]), .Q(\Inst_Mem/inst_mem_reg[61][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][24]  ( .D(\Inst_Mem/inst_mem_reg[61][24] ), .CLK(clk), .RST(rst), .I(g_init[1976]), .Q(\Inst_Mem/inst_mem_reg[61][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][25]  ( .D(\Inst_Mem/inst_mem_reg[61][25] ), .CLK(clk), .RST(rst), .I(g_init[1977]), .Q(\Inst_Mem/inst_mem_reg[61][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][26]  ( .D(\Inst_Mem/inst_mem_reg[61][26] ), .CLK(clk), .RST(rst), .I(g_init[1978]), .Q(\Inst_Mem/inst_mem_reg[61][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][27]  ( .D(\Inst_Mem/inst_mem_reg[61][27] ), .CLK(clk), .RST(rst), .I(g_init[1979]), .Q(\Inst_Mem/inst_mem_reg[61][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][28]  ( .D(\Inst_Mem/inst_mem_reg[61][28] ), .CLK(clk), .RST(rst), .I(g_init[1980]), .Q(\Inst_Mem/inst_mem_reg[61][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][29]  ( .D(\Inst_Mem/inst_mem_reg[61][29] ), .CLK(clk), .RST(rst), .I(g_init[1981]), .Q(\Inst_Mem/inst_mem_reg[61][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][30]  ( .D(\Inst_Mem/inst_mem_reg[61][30] ), .CLK(clk), .RST(rst), .I(g_init[1982]), .Q(\Inst_Mem/inst_mem_reg[61][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[61][31]  ( .D(\Inst_Mem/inst_mem_reg[61][31] ), .CLK(clk), .RST(rst), .I(g_init[1983]), .Q(\Inst_Mem/inst_mem_reg[61][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][0]  ( .D(\Inst_Mem/inst_mem_reg[60][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1920]), .Q(
        \Inst_Mem/inst_mem_reg[60][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][1]  ( .D(\Inst_Mem/inst_mem_reg[60][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1921]), .Q(
        \Inst_Mem/inst_mem_reg[60][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][2]  ( .D(\Inst_Mem/inst_mem_reg[60][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1922]), .Q(
        \Inst_Mem/inst_mem_reg[60][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][3]  ( .D(\Inst_Mem/inst_mem_reg[60][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1923]), .Q(
        \Inst_Mem/inst_mem_reg[60][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][4]  ( .D(\Inst_Mem/inst_mem_reg[60][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1924]), .Q(
        \Inst_Mem/inst_mem_reg[60][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][5]  ( .D(\Inst_Mem/inst_mem_reg[60][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1925]), .Q(
        \Inst_Mem/inst_mem_reg[60][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][6]  ( .D(\Inst_Mem/inst_mem_reg[60][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1926]), .Q(
        \Inst_Mem/inst_mem_reg[60][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][7]  ( .D(\Inst_Mem/inst_mem_reg[60][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1927]), .Q(
        \Inst_Mem/inst_mem_reg[60][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][8]  ( .D(\Inst_Mem/inst_mem_reg[60][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1928]), .Q(
        \Inst_Mem/inst_mem_reg[60][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][9]  ( .D(\Inst_Mem/inst_mem_reg[60][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1929]), .Q(
        \Inst_Mem/inst_mem_reg[60][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[60][10]  ( .D(\Inst_Mem/inst_mem_reg[60][10] ), .CLK(clk), .RST(rst), .I(g_init[1930]), .Q(\Inst_Mem/inst_mem_reg[60][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][11]  ( .D(\Inst_Mem/inst_mem_reg[60][11] ), .CLK(clk), .RST(rst), .I(g_init[1931]), .Q(\Inst_Mem/inst_mem_reg[60][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][12]  ( .D(\Inst_Mem/inst_mem_reg[60][12] ), .CLK(clk), .RST(rst), .I(g_init[1932]), .Q(\Inst_Mem/inst_mem_reg[60][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][13]  ( .D(\Inst_Mem/inst_mem_reg[60][13] ), .CLK(clk), .RST(rst), .I(g_init[1933]), .Q(\Inst_Mem/inst_mem_reg[60][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][14]  ( .D(\Inst_Mem/inst_mem_reg[60][14] ), .CLK(clk), .RST(rst), .I(g_init[1934]), .Q(\Inst_Mem/inst_mem_reg[60][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][15]  ( .D(\Inst_Mem/inst_mem_reg[60][15] ), .CLK(clk), .RST(rst), .I(g_init[1935]), .Q(\Inst_Mem/inst_mem_reg[60][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][16]  ( .D(\Inst_Mem/inst_mem_reg[60][16] ), .CLK(clk), .RST(rst), .I(g_init[1936]), .Q(\Inst_Mem/inst_mem_reg[60][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][17]  ( .D(\Inst_Mem/inst_mem_reg[60][17] ), .CLK(clk), .RST(rst), .I(g_init[1937]), .Q(\Inst_Mem/inst_mem_reg[60][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][18]  ( .D(\Inst_Mem/inst_mem_reg[60][18] ), .CLK(clk), .RST(rst), .I(g_init[1938]), .Q(\Inst_Mem/inst_mem_reg[60][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][19]  ( .D(\Inst_Mem/inst_mem_reg[60][19] ), .CLK(clk), .RST(rst), .I(g_init[1939]), .Q(\Inst_Mem/inst_mem_reg[60][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][20]  ( .D(\Inst_Mem/inst_mem_reg[60][20] ), .CLK(clk), .RST(rst), .I(g_init[1940]), .Q(\Inst_Mem/inst_mem_reg[60][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][21]  ( .D(\Inst_Mem/inst_mem_reg[60][21] ), .CLK(clk), .RST(rst), .I(g_init[1941]), .Q(\Inst_Mem/inst_mem_reg[60][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][22]  ( .D(\Inst_Mem/inst_mem_reg[60][22] ), .CLK(clk), .RST(rst), .I(g_init[1942]), .Q(\Inst_Mem/inst_mem_reg[60][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][23]  ( .D(\Inst_Mem/inst_mem_reg[60][23] ), .CLK(clk), .RST(rst), .I(g_init[1943]), .Q(\Inst_Mem/inst_mem_reg[60][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][24]  ( .D(\Inst_Mem/inst_mem_reg[60][24] ), .CLK(clk), .RST(rst), .I(g_init[1944]), .Q(\Inst_Mem/inst_mem_reg[60][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][25]  ( .D(\Inst_Mem/inst_mem_reg[60][25] ), .CLK(clk), .RST(rst), .I(g_init[1945]), .Q(\Inst_Mem/inst_mem_reg[60][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][26]  ( .D(\Inst_Mem/inst_mem_reg[60][26] ), .CLK(clk), .RST(rst), .I(g_init[1946]), .Q(\Inst_Mem/inst_mem_reg[60][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][27]  ( .D(\Inst_Mem/inst_mem_reg[60][27] ), .CLK(clk), .RST(rst), .I(g_init[1947]), .Q(\Inst_Mem/inst_mem_reg[60][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][28]  ( .D(\Inst_Mem/inst_mem_reg[60][28] ), .CLK(clk), .RST(rst), .I(g_init[1948]), .Q(\Inst_Mem/inst_mem_reg[60][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][29]  ( .D(\Inst_Mem/inst_mem_reg[60][29] ), .CLK(clk), .RST(rst), .I(g_init[1949]), .Q(\Inst_Mem/inst_mem_reg[60][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][30]  ( .D(\Inst_Mem/inst_mem_reg[60][30] ), .CLK(clk), .RST(rst), .I(g_init[1950]), .Q(\Inst_Mem/inst_mem_reg[60][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[60][31]  ( .D(\Inst_Mem/inst_mem_reg[60][31] ), .CLK(clk), .RST(rst), .I(g_init[1951]), .Q(\Inst_Mem/inst_mem_reg[60][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][0]  ( .D(\Inst_Mem/inst_mem_reg[59][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1888]), .Q(
        \Inst_Mem/inst_mem_reg[59][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][1]  ( .D(\Inst_Mem/inst_mem_reg[59][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1889]), .Q(
        \Inst_Mem/inst_mem_reg[59][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][2]  ( .D(\Inst_Mem/inst_mem_reg[59][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1890]), .Q(
        \Inst_Mem/inst_mem_reg[59][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][3]  ( .D(\Inst_Mem/inst_mem_reg[59][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1891]), .Q(
        \Inst_Mem/inst_mem_reg[59][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][4]  ( .D(\Inst_Mem/inst_mem_reg[59][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1892]), .Q(
        \Inst_Mem/inst_mem_reg[59][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][5]  ( .D(\Inst_Mem/inst_mem_reg[59][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1893]), .Q(
        \Inst_Mem/inst_mem_reg[59][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][6]  ( .D(\Inst_Mem/inst_mem_reg[59][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1894]), .Q(
        \Inst_Mem/inst_mem_reg[59][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][7]  ( .D(\Inst_Mem/inst_mem_reg[59][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1895]), .Q(
        \Inst_Mem/inst_mem_reg[59][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][8]  ( .D(\Inst_Mem/inst_mem_reg[59][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1896]), .Q(
        \Inst_Mem/inst_mem_reg[59][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][9]  ( .D(\Inst_Mem/inst_mem_reg[59][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1897]), .Q(
        \Inst_Mem/inst_mem_reg[59][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[59][10]  ( .D(\Inst_Mem/inst_mem_reg[59][10] ), .CLK(clk), .RST(rst), .I(g_init[1898]), .Q(\Inst_Mem/inst_mem_reg[59][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][11]  ( .D(\Inst_Mem/inst_mem_reg[59][11] ), .CLK(clk), .RST(rst), .I(g_init[1899]), .Q(\Inst_Mem/inst_mem_reg[59][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][12]  ( .D(\Inst_Mem/inst_mem_reg[59][12] ), .CLK(clk), .RST(rst), .I(g_init[1900]), .Q(\Inst_Mem/inst_mem_reg[59][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][13]  ( .D(\Inst_Mem/inst_mem_reg[59][13] ), .CLK(clk), .RST(rst), .I(g_init[1901]), .Q(\Inst_Mem/inst_mem_reg[59][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][14]  ( .D(\Inst_Mem/inst_mem_reg[59][14] ), .CLK(clk), .RST(rst), .I(g_init[1902]), .Q(\Inst_Mem/inst_mem_reg[59][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][15]  ( .D(\Inst_Mem/inst_mem_reg[59][15] ), .CLK(clk), .RST(rst), .I(g_init[1903]), .Q(\Inst_Mem/inst_mem_reg[59][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][16]  ( .D(\Inst_Mem/inst_mem_reg[59][16] ), .CLK(clk), .RST(rst), .I(g_init[1904]), .Q(\Inst_Mem/inst_mem_reg[59][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][17]  ( .D(\Inst_Mem/inst_mem_reg[59][17] ), .CLK(clk), .RST(rst), .I(g_init[1905]), .Q(\Inst_Mem/inst_mem_reg[59][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][18]  ( .D(\Inst_Mem/inst_mem_reg[59][18] ), .CLK(clk), .RST(rst), .I(g_init[1906]), .Q(\Inst_Mem/inst_mem_reg[59][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][19]  ( .D(\Inst_Mem/inst_mem_reg[59][19] ), .CLK(clk), .RST(rst), .I(g_init[1907]), .Q(\Inst_Mem/inst_mem_reg[59][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][20]  ( .D(\Inst_Mem/inst_mem_reg[59][20] ), .CLK(clk), .RST(rst), .I(g_init[1908]), .Q(\Inst_Mem/inst_mem_reg[59][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][21]  ( .D(\Inst_Mem/inst_mem_reg[59][21] ), .CLK(clk), .RST(rst), .I(g_init[1909]), .Q(\Inst_Mem/inst_mem_reg[59][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][22]  ( .D(\Inst_Mem/inst_mem_reg[59][22] ), .CLK(clk), .RST(rst), .I(g_init[1910]), .Q(\Inst_Mem/inst_mem_reg[59][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][23]  ( .D(\Inst_Mem/inst_mem_reg[59][23] ), .CLK(clk), .RST(rst), .I(g_init[1911]), .Q(\Inst_Mem/inst_mem_reg[59][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][24]  ( .D(\Inst_Mem/inst_mem_reg[59][24] ), .CLK(clk), .RST(rst), .I(g_init[1912]), .Q(\Inst_Mem/inst_mem_reg[59][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][25]  ( .D(\Inst_Mem/inst_mem_reg[59][25] ), .CLK(clk), .RST(rst), .I(g_init[1913]), .Q(\Inst_Mem/inst_mem_reg[59][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][26]  ( .D(\Inst_Mem/inst_mem_reg[59][26] ), .CLK(clk), .RST(rst), .I(g_init[1914]), .Q(\Inst_Mem/inst_mem_reg[59][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][27]  ( .D(\Inst_Mem/inst_mem_reg[59][27] ), .CLK(clk), .RST(rst), .I(g_init[1915]), .Q(\Inst_Mem/inst_mem_reg[59][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][28]  ( .D(\Inst_Mem/inst_mem_reg[59][28] ), .CLK(clk), .RST(rst), .I(g_init[1916]), .Q(\Inst_Mem/inst_mem_reg[59][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][29]  ( .D(\Inst_Mem/inst_mem_reg[59][29] ), .CLK(clk), .RST(rst), .I(g_init[1917]), .Q(\Inst_Mem/inst_mem_reg[59][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][30]  ( .D(\Inst_Mem/inst_mem_reg[59][30] ), .CLK(clk), .RST(rst), .I(g_init[1918]), .Q(\Inst_Mem/inst_mem_reg[59][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[59][31]  ( .D(\Inst_Mem/inst_mem_reg[59][31] ), .CLK(clk), .RST(rst), .I(g_init[1919]), .Q(\Inst_Mem/inst_mem_reg[59][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][0]  ( .D(\Inst_Mem/inst_mem_reg[58][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1856]), .Q(
        \Inst_Mem/inst_mem_reg[58][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][1]  ( .D(\Inst_Mem/inst_mem_reg[58][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1857]), .Q(
        \Inst_Mem/inst_mem_reg[58][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][2]  ( .D(\Inst_Mem/inst_mem_reg[58][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1858]), .Q(
        \Inst_Mem/inst_mem_reg[58][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][3]  ( .D(\Inst_Mem/inst_mem_reg[58][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1859]), .Q(
        \Inst_Mem/inst_mem_reg[58][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][4]  ( .D(\Inst_Mem/inst_mem_reg[58][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1860]), .Q(
        \Inst_Mem/inst_mem_reg[58][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][5]  ( .D(\Inst_Mem/inst_mem_reg[58][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1861]), .Q(
        \Inst_Mem/inst_mem_reg[58][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][6]  ( .D(\Inst_Mem/inst_mem_reg[58][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1862]), .Q(
        \Inst_Mem/inst_mem_reg[58][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][7]  ( .D(\Inst_Mem/inst_mem_reg[58][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1863]), .Q(
        \Inst_Mem/inst_mem_reg[58][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][8]  ( .D(\Inst_Mem/inst_mem_reg[58][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1864]), .Q(
        \Inst_Mem/inst_mem_reg[58][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][9]  ( .D(\Inst_Mem/inst_mem_reg[58][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1865]), .Q(
        \Inst_Mem/inst_mem_reg[58][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[58][10]  ( .D(\Inst_Mem/inst_mem_reg[58][10] ), .CLK(clk), .RST(rst), .I(g_init[1866]), .Q(\Inst_Mem/inst_mem_reg[58][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][11]  ( .D(\Inst_Mem/inst_mem_reg[58][11] ), .CLK(clk), .RST(rst), .I(g_init[1867]), .Q(\Inst_Mem/inst_mem_reg[58][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][12]  ( .D(\Inst_Mem/inst_mem_reg[58][12] ), .CLK(clk), .RST(rst), .I(g_init[1868]), .Q(\Inst_Mem/inst_mem_reg[58][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][13]  ( .D(\Inst_Mem/inst_mem_reg[58][13] ), .CLK(clk), .RST(rst), .I(g_init[1869]), .Q(\Inst_Mem/inst_mem_reg[58][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][14]  ( .D(\Inst_Mem/inst_mem_reg[58][14] ), .CLK(clk), .RST(rst), .I(g_init[1870]), .Q(\Inst_Mem/inst_mem_reg[58][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][15]  ( .D(\Inst_Mem/inst_mem_reg[58][15] ), .CLK(clk), .RST(rst), .I(g_init[1871]), .Q(\Inst_Mem/inst_mem_reg[58][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][16]  ( .D(\Inst_Mem/inst_mem_reg[58][16] ), .CLK(clk), .RST(rst), .I(g_init[1872]), .Q(\Inst_Mem/inst_mem_reg[58][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][17]  ( .D(\Inst_Mem/inst_mem_reg[58][17] ), .CLK(clk), .RST(rst), .I(g_init[1873]), .Q(\Inst_Mem/inst_mem_reg[58][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][18]  ( .D(\Inst_Mem/inst_mem_reg[58][18] ), .CLK(clk), .RST(rst), .I(g_init[1874]), .Q(\Inst_Mem/inst_mem_reg[58][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][19]  ( .D(\Inst_Mem/inst_mem_reg[58][19] ), .CLK(clk), .RST(rst), .I(g_init[1875]), .Q(\Inst_Mem/inst_mem_reg[58][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][20]  ( .D(\Inst_Mem/inst_mem_reg[58][20] ), .CLK(clk), .RST(rst), .I(g_init[1876]), .Q(\Inst_Mem/inst_mem_reg[58][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][21]  ( .D(\Inst_Mem/inst_mem_reg[58][21] ), .CLK(clk), .RST(rst), .I(g_init[1877]), .Q(\Inst_Mem/inst_mem_reg[58][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][22]  ( .D(\Inst_Mem/inst_mem_reg[58][22] ), .CLK(clk), .RST(rst), .I(g_init[1878]), .Q(\Inst_Mem/inst_mem_reg[58][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][23]  ( .D(\Inst_Mem/inst_mem_reg[58][23] ), .CLK(clk), .RST(rst), .I(g_init[1879]), .Q(\Inst_Mem/inst_mem_reg[58][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][24]  ( .D(\Inst_Mem/inst_mem_reg[58][24] ), .CLK(clk), .RST(rst), .I(g_init[1880]), .Q(\Inst_Mem/inst_mem_reg[58][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][25]  ( .D(\Inst_Mem/inst_mem_reg[58][25] ), .CLK(clk), .RST(rst), .I(g_init[1881]), .Q(\Inst_Mem/inst_mem_reg[58][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][26]  ( .D(\Inst_Mem/inst_mem_reg[58][26] ), .CLK(clk), .RST(rst), .I(g_init[1882]), .Q(\Inst_Mem/inst_mem_reg[58][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][27]  ( .D(\Inst_Mem/inst_mem_reg[58][27] ), .CLK(clk), .RST(rst), .I(g_init[1883]), .Q(\Inst_Mem/inst_mem_reg[58][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][28]  ( .D(\Inst_Mem/inst_mem_reg[58][28] ), .CLK(clk), .RST(rst), .I(g_init[1884]), .Q(\Inst_Mem/inst_mem_reg[58][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][29]  ( .D(\Inst_Mem/inst_mem_reg[58][29] ), .CLK(clk), .RST(rst), .I(g_init[1885]), .Q(\Inst_Mem/inst_mem_reg[58][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][30]  ( .D(\Inst_Mem/inst_mem_reg[58][30] ), .CLK(clk), .RST(rst), .I(g_init[1886]), .Q(\Inst_Mem/inst_mem_reg[58][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[58][31]  ( .D(\Inst_Mem/inst_mem_reg[58][31] ), .CLK(clk), .RST(rst), .I(g_init[1887]), .Q(\Inst_Mem/inst_mem_reg[58][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][0]  ( .D(\Inst_Mem/inst_mem_reg[57][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1824]), .Q(
        \Inst_Mem/inst_mem_reg[57][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][1]  ( .D(\Inst_Mem/inst_mem_reg[57][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1825]), .Q(
        \Inst_Mem/inst_mem_reg[57][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][2]  ( .D(\Inst_Mem/inst_mem_reg[57][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1826]), .Q(
        \Inst_Mem/inst_mem_reg[57][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][3]  ( .D(\Inst_Mem/inst_mem_reg[57][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1827]), .Q(
        \Inst_Mem/inst_mem_reg[57][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][4]  ( .D(\Inst_Mem/inst_mem_reg[57][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1828]), .Q(
        \Inst_Mem/inst_mem_reg[57][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][5]  ( .D(\Inst_Mem/inst_mem_reg[57][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1829]), .Q(
        \Inst_Mem/inst_mem_reg[57][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][6]  ( .D(\Inst_Mem/inst_mem_reg[57][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1830]), .Q(
        \Inst_Mem/inst_mem_reg[57][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][7]  ( .D(\Inst_Mem/inst_mem_reg[57][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1831]), .Q(
        \Inst_Mem/inst_mem_reg[57][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][8]  ( .D(\Inst_Mem/inst_mem_reg[57][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1832]), .Q(
        \Inst_Mem/inst_mem_reg[57][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][9]  ( .D(\Inst_Mem/inst_mem_reg[57][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1833]), .Q(
        \Inst_Mem/inst_mem_reg[57][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[57][10]  ( .D(\Inst_Mem/inst_mem_reg[57][10] ), .CLK(clk), .RST(rst), .I(g_init[1834]), .Q(\Inst_Mem/inst_mem_reg[57][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][11]  ( .D(\Inst_Mem/inst_mem_reg[57][11] ), .CLK(clk), .RST(rst), .I(g_init[1835]), .Q(\Inst_Mem/inst_mem_reg[57][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][12]  ( .D(\Inst_Mem/inst_mem_reg[57][12] ), .CLK(clk), .RST(rst), .I(g_init[1836]), .Q(\Inst_Mem/inst_mem_reg[57][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][13]  ( .D(\Inst_Mem/inst_mem_reg[57][13] ), .CLK(clk), .RST(rst), .I(g_init[1837]), .Q(\Inst_Mem/inst_mem_reg[57][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][14]  ( .D(\Inst_Mem/inst_mem_reg[57][14] ), .CLK(clk), .RST(rst), .I(g_init[1838]), .Q(\Inst_Mem/inst_mem_reg[57][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][15]  ( .D(\Inst_Mem/inst_mem_reg[57][15] ), .CLK(clk), .RST(rst), .I(g_init[1839]), .Q(\Inst_Mem/inst_mem_reg[57][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][16]  ( .D(\Inst_Mem/inst_mem_reg[57][16] ), .CLK(clk), .RST(rst), .I(g_init[1840]), .Q(\Inst_Mem/inst_mem_reg[57][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][17]  ( .D(\Inst_Mem/inst_mem_reg[57][17] ), .CLK(clk), .RST(rst), .I(g_init[1841]), .Q(\Inst_Mem/inst_mem_reg[57][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][18]  ( .D(\Inst_Mem/inst_mem_reg[57][18] ), .CLK(clk), .RST(rst), .I(g_init[1842]), .Q(\Inst_Mem/inst_mem_reg[57][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][19]  ( .D(\Inst_Mem/inst_mem_reg[57][19] ), .CLK(clk), .RST(rst), .I(g_init[1843]), .Q(\Inst_Mem/inst_mem_reg[57][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][20]  ( .D(\Inst_Mem/inst_mem_reg[57][20] ), .CLK(clk), .RST(rst), .I(g_init[1844]), .Q(\Inst_Mem/inst_mem_reg[57][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][21]  ( .D(\Inst_Mem/inst_mem_reg[57][21] ), .CLK(clk), .RST(rst), .I(g_init[1845]), .Q(\Inst_Mem/inst_mem_reg[57][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][22]  ( .D(\Inst_Mem/inst_mem_reg[57][22] ), .CLK(clk), .RST(rst), .I(g_init[1846]), .Q(\Inst_Mem/inst_mem_reg[57][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][23]  ( .D(\Inst_Mem/inst_mem_reg[57][23] ), .CLK(clk), .RST(rst), .I(g_init[1847]), .Q(\Inst_Mem/inst_mem_reg[57][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][24]  ( .D(\Inst_Mem/inst_mem_reg[57][24] ), .CLK(clk), .RST(rst), .I(g_init[1848]), .Q(\Inst_Mem/inst_mem_reg[57][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][25]  ( .D(\Inst_Mem/inst_mem_reg[57][25] ), .CLK(clk), .RST(rst), .I(g_init[1849]), .Q(\Inst_Mem/inst_mem_reg[57][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][26]  ( .D(\Inst_Mem/inst_mem_reg[57][26] ), .CLK(clk), .RST(rst), .I(g_init[1850]), .Q(\Inst_Mem/inst_mem_reg[57][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][27]  ( .D(\Inst_Mem/inst_mem_reg[57][27] ), .CLK(clk), .RST(rst), .I(g_init[1851]), .Q(\Inst_Mem/inst_mem_reg[57][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][28]  ( .D(\Inst_Mem/inst_mem_reg[57][28] ), .CLK(clk), .RST(rst), .I(g_init[1852]), .Q(\Inst_Mem/inst_mem_reg[57][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][29]  ( .D(\Inst_Mem/inst_mem_reg[57][29] ), .CLK(clk), .RST(rst), .I(g_init[1853]), .Q(\Inst_Mem/inst_mem_reg[57][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][30]  ( .D(\Inst_Mem/inst_mem_reg[57][30] ), .CLK(clk), .RST(rst), .I(g_init[1854]), .Q(\Inst_Mem/inst_mem_reg[57][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[57][31]  ( .D(\Inst_Mem/inst_mem_reg[57][31] ), .CLK(clk), .RST(rst), .I(g_init[1855]), .Q(\Inst_Mem/inst_mem_reg[57][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][0]  ( .D(\Inst_Mem/inst_mem_reg[56][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1792]), .Q(
        \Inst_Mem/inst_mem_reg[56][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][1]  ( .D(\Inst_Mem/inst_mem_reg[56][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1793]), .Q(
        \Inst_Mem/inst_mem_reg[56][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][2]  ( .D(\Inst_Mem/inst_mem_reg[56][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1794]), .Q(
        \Inst_Mem/inst_mem_reg[56][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][3]  ( .D(\Inst_Mem/inst_mem_reg[56][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1795]), .Q(
        \Inst_Mem/inst_mem_reg[56][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][4]  ( .D(\Inst_Mem/inst_mem_reg[56][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1796]), .Q(
        \Inst_Mem/inst_mem_reg[56][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][5]  ( .D(\Inst_Mem/inst_mem_reg[56][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1797]), .Q(
        \Inst_Mem/inst_mem_reg[56][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][6]  ( .D(\Inst_Mem/inst_mem_reg[56][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1798]), .Q(
        \Inst_Mem/inst_mem_reg[56][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][7]  ( .D(\Inst_Mem/inst_mem_reg[56][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1799]), .Q(
        \Inst_Mem/inst_mem_reg[56][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][8]  ( .D(\Inst_Mem/inst_mem_reg[56][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1800]), .Q(
        \Inst_Mem/inst_mem_reg[56][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][9]  ( .D(\Inst_Mem/inst_mem_reg[56][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1801]), .Q(
        \Inst_Mem/inst_mem_reg[56][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[56][10]  ( .D(\Inst_Mem/inst_mem_reg[56][10] ), .CLK(clk), .RST(rst), .I(g_init[1802]), .Q(\Inst_Mem/inst_mem_reg[56][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][11]  ( .D(\Inst_Mem/inst_mem_reg[56][11] ), .CLK(clk), .RST(rst), .I(g_init[1803]), .Q(\Inst_Mem/inst_mem_reg[56][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][12]  ( .D(\Inst_Mem/inst_mem_reg[56][12] ), .CLK(clk), .RST(rst), .I(g_init[1804]), .Q(\Inst_Mem/inst_mem_reg[56][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][13]  ( .D(\Inst_Mem/inst_mem_reg[56][13] ), .CLK(clk), .RST(rst), .I(g_init[1805]), .Q(\Inst_Mem/inst_mem_reg[56][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][14]  ( .D(\Inst_Mem/inst_mem_reg[56][14] ), .CLK(clk), .RST(rst), .I(g_init[1806]), .Q(\Inst_Mem/inst_mem_reg[56][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][15]  ( .D(\Inst_Mem/inst_mem_reg[56][15] ), .CLK(clk), .RST(rst), .I(g_init[1807]), .Q(\Inst_Mem/inst_mem_reg[56][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][16]  ( .D(\Inst_Mem/inst_mem_reg[56][16] ), .CLK(clk), .RST(rst), .I(g_init[1808]), .Q(\Inst_Mem/inst_mem_reg[56][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][17]  ( .D(\Inst_Mem/inst_mem_reg[56][17] ), .CLK(clk), .RST(rst), .I(g_init[1809]), .Q(\Inst_Mem/inst_mem_reg[56][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][18]  ( .D(\Inst_Mem/inst_mem_reg[56][18] ), .CLK(clk), .RST(rst), .I(g_init[1810]), .Q(\Inst_Mem/inst_mem_reg[56][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][19]  ( .D(\Inst_Mem/inst_mem_reg[56][19] ), .CLK(clk), .RST(rst), .I(g_init[1811]), .Q(\Inst_Mem/inst_mem_reg[56][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][20]  ( .D(\Inst_Mem/inst_mem_reg[56][20] ), .CLK(clk), .RST(rst), .I(g_init[1812]), .Q(\Inst_Mem/inst_mem_reg[56][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][21]  ( .D(\Inst_Mem/inst_mem_reg[56][21] ), .CLK(clk), .RST(rst), .I(g_init[1813]), .Q(\Inst_Mem/inst_mem_reg[56][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][22]  ( .D(\Inst_Mem/inst_mem_reg[56][22] ), .CLK(clk), .RST(rst), .I(g_init[1814]), .Q(\Inst_Mem/inst_mem_reg[56][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][23]  ( .D(\Inst_Mem/inst_mem_reg[56][23] ), .CLK(clk), .RST(rst), .I(g_init[1815]), .Q(\Inst_Mem/inst_mem_reg[56][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][24]  ( .D(\Inst_Mem/inst_mem_reg[56][24] ), .CLK(clk), .RST(rst), .I(g_init[1816]), .Q(\Inst_Mem/inst_mem_reg[56][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][25]  ( .D(\Inst_Mem/inst_mem_reg[56][25] ), .CLK(clk), .RST(rst), .I(g_init[1817]), .Q(\Inst_Mem/inst_mem_reg[56][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][26]  ( .D(\Inst_Mem/inst_mem_reg[56][26] ), .CLK(clk), .RST(rst), .I(g_init[1818]), .Q(\Inst_Mem/inst_mem_reg[56][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][27]  ( .D(\Inst_Mem/inst_mem_reg[56][27] ), .CLK(clk), .RST(rst), .I(g_init[1819]), .Q(\Inst_Mem/inst_mem_reg[56][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][28]  ( .D(\Inst_Mem/inst_mem_reg[56][28] ), .CLK(clk), .RST(rst), .I(g_init[1820]), .Q(\Inst_Mem/inst_mem_reg[56][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][29]  ( .D(\Inst_Mem/inst_mem_reg[56][29] ), .CLK(clk), .RST(rst), .I(g_init[1821]), .Q(\Inst_Mem/inst_mem_reg[56][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][30]  ( .D(\Inst_Mem/inst_mem_reg[56][30] ), .CLK(clk), .RST(rst), .I(g_init[1822]), .Q(\Inst_Mem/inst_mem_reg[56][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[56][31]  ( .D(\Inst_Mem/inst_mem_reg[56][31] ), .CLK(clk), .RST(rst), .I(g_init[1823]), .Q(\Inst_Mem/inst_mem_reg[56][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][0]  ( .D(\Inst_Mem/inst_mem_reg[55][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1760]), .Q(
        \Inst_Mem/inst_mem_reg[55][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][1]  ( .D(\Inst_Mem/inst_mem_reg[55][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1761]), .Q(
        \Inst_Mem/inst_mem_reg[55][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][2]  ( .D(\Inst_Mem/inst_mem_reg[55][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1762]), .Q(
        \Inst_Mem/inst_mem_reg[55][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][3]  ( .D(\Inst_Mem/inst_mem_reg[55][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1763]), .Q(
        \Inst_Mem/inst_mem_reg[55][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][4]  ( .D(\Inst_Mem/inst_mem_reg[55][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1764]), .Q(
        \Inst_Mem/inst_mem_reg[55][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][5]  ( .D(\Inst_Mem/inst_mem_reg[55][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1765]), .Q(
        \Inst_Mem/inst_mem_reg[55][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][6]  ( .D(\Inst_Mem/inst_mem_reg[55][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1766]), .Q(
        \Inst_Mem/inst_mem_reg[55][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][7]  ( .D(\Inst_Mem/inst_mem_reg[55][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1767]), .Q(
        \Inst_Mem/inst_mem_reg[55][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][8]  ( .D(\Inst_Mem/inst_mem_reg[55][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1768]), .Q(
        \Inst_Mem/inst_mem_reg[55][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][9]  ( .D(\Inst_Mem/inst_mem_reg[55][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1769]), .Q(
        \Inst_Mem/inst_mem_reg[55][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[55][10]  ( .D(\Inst_Mem/inst_mem_reg[55][10] ), .CLK(clk), .RST(rst), .I(g_init[1770]), .Q(\Inst_Mem/inst_mem_reg[55][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][11]  ( .D(\Inst_Mem/inst_mem_reg[55][11] ), .CLK(clk), .RST(rst), .I(g_init[1771]), .Q(\Inst_Mem/inst_mem_reg[55][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][12]  ( .D(\Inst_Mem/inst_mem_reg[55][12] ), .CLK(clk), .RST(rst), .I(g_init[1772]), .Q(\Inst_Mem/inst_mem_reg[55][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][13]  ( .D(\Inst_Mem/inst_mem_reg[55][13] ), .CLK(clk), .RST(rst), .I(g_init[1773]), .Q(\Inst_Mem/inst_mem_reg[55][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][14]  ( .D(\Inst_Mem/inst_mem_reg[55][14] ), .CLK(clk), .RST(rst), .I(g_init[1774]), .Q(\Inst_Mem/inst_mem_reg[55][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][15]  ( .D(\Inst_Mem/inst_mem_reg[55][15] ), .CLK(clk), .RST(rst), .I(g_init[1775]), .Q(\Inst_Mem/inst_mem_reg[55][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][16]  ( .D(\Inst_Mem/inst_mem_reg[55][16] ), .CLK(clk), .RST(rst), .I(g_init[1776]), .Q(\Inst_Mem/inst_mem_reg[55][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][17]  ( .D(\Inst_Mem/inst_mem_reg[55][17] ), .CLK(clk), .RST(rst), .I(g_init[1777]), .Q(\Inst_Mem/inst_mem_reg[55][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][18]  ( .D(\Inst_Mem/inst_mem_reg[55][18] ), .CLK(clk), .RST(rst), .I(g_init[1778]), .Q(\Inst_Mem/inst_mem_reg[55][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][19]  ( .D(\Inst_Mem/inst_mem_reg[55][19] ), .CLK(clk), .RST(rst), .I(g_init[1779]), .Q(\Inst_Mem/inst_mem_reg[55][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][20]  ( .D(\Inst_Mem/inst_mem_reg[55][20] ), .CLK(clk), .RST(rst), .I(g_init[1780]), .Q(\Inst_Mem/inst_mem_reg[55][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][21]  ( .D(\Inst_Mem/inst_mem_reg[55][21] ), .CLK(clk), .RST(rst), .I(g_init[1781]), .Q(\Inst_Mem/inst_mem_reg[55][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][22]  ( .D(\Inst_Mem/inst_mem_reg[55][22] ), .CLK(clk), .RST(rst), .I(g_init[1782]), .Q(\Inst_Mem/inst_mem_reg[55][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][23]  ( .D(\Inst_Mem/inst_mem_reg[55][23] ), .CLK(clk), .RST(rst), .I(g_init[1783]), .Q(\Inst_Mem/inst_mem_reg[55][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][24]  ( .D(\Inst_Mem/inst_mem_reg[55][24] ), .CLK(clk), .RST(rst), .I(g_init[1784]), .Q(\Inst_Mem/inst_mem_reg[55][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][25]  ( .D(\Inst_Mem/inst_mem_reg[55][25] ), .CLK(clk), .RST(rst), .I(g_init[1785]), .Q(\Inst_Mem/inst_mem_reg[55][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][26]  ( .D(\Inst_Mem/inst_mem_reg[55][26] ), .CLK(clk), .RST(rst), .I(g_init[1786]), .Q(\Inst_Mem/inst_mem_reg[55][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][27]  ( .D(\Inst_Mem/inst_mem_reg[55][27] ), .CLK(clk), .RST(rst), .I(g_init[1787]), .Q(\Inst_Mem/inst_mem_reg[55][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][28]  ( .D(\Inst_Mem/inst_mem_reg[55][28] ), .CLK(clk), .RST(rst), .I(g_init[1788]), .Q(\Inst_Mem/inst_mem_reg[55][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][29]  ( .D(\Inst_Mem/inst_mem_reg[55][29] ), .CLK(clk), .RST(rst), .I(g_init[1789]), .Q(\Inst_Mem/inst_mem_reg[55][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][30]  ( .D(\Inst_Mem/inst_mem_reg[55][30] ), .CLK(clk), .RST(rst), .I(g_init[1790]), .Q(\Inst_Mem/inst_mem_reg[55][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[55][31]  ( .D(\Inst_Mem/inst_mem_reg[55][31] ), .CLK(clk), .RST(rst), .I(g_init[1791]), .Q(\Inst_Mem/inst_mem_reg[55][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][0]  ( .D(\Inst_Mem/inst_mem_reg[54][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1728]), .Q(
        \Inst_Mem/inst_mem_reg[54][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][1]  ( .D(\Inst_Mem/inst_mem_reg[54][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1729]), .Q(
        \Inst_Mem/inst_mem_reg[54][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][2]  ( .D(\Inst_Mem/inst_mem_reg[54][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1730]), .Q(
        \Inst_Mem/inst_mem_reg[54][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][3]  ( .D(\Inst_Mem/inst_mem_reg[54][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1731]), .Q(
        \Inst_Mem/inst_mem_reg[54][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][4]  ( .D(\Inst_Mem/inst_mem_reg[54][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1732]), .Q(
        \Inst_Mem/inst_mem_reg[54][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][5]  ( .D(\Inst_Mem/inst_mem_reg[54][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1733]), .Q(
        \Inst_Mem/inst_mem_reg[54][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][6]  ( .D(\Inst_Mem/inst_mem_reg[54][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1734]), .Q(
        \Inst_Mem/inst_mem_reg[54][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][7]  ( .D(\Inst_Mem/inst_mem_reg[54][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1735]), .Q(
        \Inst_Mem/inst_mem_reg[54][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][8]  ( .D(\Inst_Mem/inst_mem_reg[54][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1736]), .Q(
        \Inst_Mem/inst_mem_reg[54][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][9]  ( .D(\Inst_Mem/inst_mem_reg[54][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1737]), .Q(
        \Inst_Mem/inst_mem_reg[54][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[54][10]  ( .D(\Inst_Mem/inst_mem_reg[54][10] ), .CLK(clk), .RST(rst), .I(g_init[1738]), .Q(\Inst_Mem/inst_mem_reg[54][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][11]  ( .D(\Inst_Mem/inst_mem_reg[54][11] ), .CLK(clk), .RST(rst), .I(g_init[1739]), .Q(\Inst_Mem/inst_mem_reg[54][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][12]  ( .D(\Inst_Mem/inst_mem_reg[54][12] ), .CLK(clk), .RST(rst), .I(g_init[1740]), .Q(\Inst_Mem/inst_mem_reg[54][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][13]  ( .D(\Inst_Mem/inst_mem_reg[54][13] ), .CLK(clk), .RST(rst), .I(g_init[1741]), .Q(\Inst_Mem/inst_mem_reg[54][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][14]  ( .D(\Inst_Mem/inst_mem_reg[54][14] ), .CLK(clk), .RST(rst), .I(g_init[1742]), .Q(\Inst_Mem/inst_mem_reg[54][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][15]  ( .D(\Inst_Mem/inst_mem_reg[54][15] ), .CLK(clk), .RST(rst), .I(g_init[1743]), .Q(\Inst_Mem/inst_mem_reg[54][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][16]  ( .D(\Inst_Mem/inst_mem_reg[54][16] ), .CLK(clk), .RST(rst), .I(g_init[1744]), .Q(\Inst_Mem/inst_mem_reg[54][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][17]  ( .D(\Inst_Mem/inst_mem_reg[54][17] ), .CLK(clk), .RST(rst), .I(g_init[1745]), .Q(\Inst_Mem/inst_mem_reg[54][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][18]  ( .D(\Inst_Mem/inst_mem_reg[54][18] ), .CLK(clk), .RST(rst), .I(g_init[1746]), .Q(\Inst_Mem/inst_mem_reg[54][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][19]  ( .D(\Inst_Mem/inst_mem_reg[54][19] ), .CLK(clk), .RST(rst), .I(g_init[1747]), .Q(\Inst_Mem/inst_mem_reg[54][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][20]  ( .D(\Inst_Mem/inst_mem_reg[54][20] ), .CLK(clk), .RST(rst), .I(g_init[1748]), .Q(\Inst_Mem/inst_mem_reg[54][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][21]  ( .D(\Inst_Mem/inst_mem_reg[54][21] ), .CLK(clk), .RST(rst), .I(g_init[1749]), .Q(\Inst_Mem/inst_mem_reg[54][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][22]  ( .D(\Inst_Mem/inst_mem_reg[54][22] ), .CLK(clk), .RST(rst), .I(g_init[1750]), .Q(\Inst_Mem/inst_mem_reg[54][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][23]  ( .D(\Inst_Mem/inst_mem_reg[54][23] ), .CLK(clk), .RST(rst), .I(g_init[1751]), .Q(\Inst_Mem/inst_mem_reg[54][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][24]  ( .D(\Inst_Mem/inst_mem_reg[54][24] ), .CLK(clk), .RST(rst), .I(g_init[1752]), .Q(\Inst_Mem/inst_mem_reg[54][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][25]  ( .D(\Inst_Mem/inst_mem_reg[54][25] ), .CLK(clk), .RST(rst), .I(g_init[1753]), .Q(\Inst_Mem/inst_mem_reg[54][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][26]  ( .D(\Inst_Mem/inst_mem_reg[54][26] ), .CLK(clk), .RST(rst), .I(g_init[1754]), .Q(\Inst_Mem/inst_mem_reg[54][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][27]  ( .D(\Inst_Mem/inst_mem_reg[54][27] ), .CLK(clk), .RST(rst), .I(g_init[1755]), .Q(\Inst_Mem/inst_mem_reg[54][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][28]  ( .D(\Inst_Mem/inst_mem_reg[54][28] ), .CLK(clk), .RST(rst), .I(g_init[1756]), .Q(\Inst_Mem/inst_mem_reg[54][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][29]  ( .D(\Inst_Mem/inst_mem_reg[54][29] ), .CLK(clk), .RST(rst), .I(g_init[1757]), .Q(\Inst_Mem/inst_mem_reg[54][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][30]  ( .D(\Inst_Mem/inst_mem_reg[54][30] ), .CLK(clk), .RST(rst), .I(g_init[1758]), .Q(\Inst_Mem/inst_mem_reg[54][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[54][31]  ( .D(\Inst_Mem/inst_mem_reg[54][31] ), .CLK(clk), .RST(rst), .I(g_init[1759]), .Q(\Inst_Mem/inst_mem_reg[54][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][0]  ( .D(\Inst_Mem/inst_mem_reg[53][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1696]), .Q(
        \Inst_Mem/inst_mem_reg[53][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][1]  ( .D(\Inst_Mem/inst_mem_reg[53][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1697]), .Q(
        \Inst_Mem/inst_mem_reg[53][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][2]  ( .D(\Inst_Mem/inst_mem_reg[53][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1698]), .Q(
        \Inst_Mem/inst_mem_reg[53][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][3]  ( .D(\Inst_Mem/inst_mem_reg[53][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1699]), .Q(
        \Inst_Mem/inst_mem_reg[53][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][4]  ( .D(\Inst_Mem/inst_mem_reg[53][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1700]), .Q(
        \Inst_Mem/inst_mem_reg[53][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][5]  ( .D(\Inst_Mem/inst_mem_reg[53][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1701]), .Q(
        \Inst_Mem/inst_mem_reg[53][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][6]  ( .D(\Inst_Mem/inst_mem_reg[53][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1702]), .Q(
        \Inst_Mem/inst_mem_reg[53][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][7]  ( .D(\Inst_Mem/inst_mem_reg[53][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1703]), .Q(
        \Inst_Mem/inst_mem_reg[53][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][8]  ( .D(\Inst_Mem/inst_mem_reg[53][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1704]), .Q(
        \Inst_Mem/inst_mem_reg[53][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][9]  ( .D(\Inst_Mem/inst_mem_reg[53][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1705]), .Q(
        \Inst_Mem/inst_mem_reg[53][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[53][10]  ( .D(\Inst_Mem/inst_mem_reg[53][10] ), .CLK(clk), .RST(rst), .I(g_init[1706]), .Q(\Inst_Mem/inst_mem_reg[53][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][11]  ( .D(\Inst_Mem/inst_mem_reg[53][11] ), .CLK(clk), .RST(rst), .I(g_init[1707]), .Q(\Inst_Mem/inst_mem_reg[53][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][12]  ( .D(\Inst_Mem/inst_mem_reg[53][12] ), .CLK(clk), .RST(rst), .I(g_init[1708]), .Q(\Inst_Mem/inst_mem_reg[53][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][13]  ( .D(\Inst_Mem/inst_mem_reg[53][13] ), .CLK(clk), .RST(rst), .I(g_init[1709]), .Q(\Inst_Mem/inst_mem_reg[53][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][14]  ( .D(\Inst_Mem/inst_mem_reg[53][14] ), .CLK(clk), .RST(rst), .I(g_init[1710]), .Q(\Inst_Mem/inst_mem_reg[53][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][15]  ( .D(\Inst_Mem/inst_mem_reg[53][15] ), .CLK(clk), .RST(rst), .I(g_init[1711]), .Q(\Inst_Mem/inst_mem_reg[53][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][16]  ( .D(\Inst_Mem/inst_mem_reg[53][16] ), .CLK(clk), .RST(rst), .I(g_init[1712]), .Q(\Inst_Mem/inst_mem_reg[53][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][17]  ( .D(\Inst_Mem/inst_mem_reg[53][17] ), .CLK(clk), .RST(rst), .I(g_init[1713]), .Q(\Inst_Mem/inst_mem_reg[53][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][18]  ( .D(\Inst_Mem/inst_mem_reg[53][18] ), .CLK(clk), .RST(rst), .I(g_init[1714]), .Q(\Inst_Mem/inst_mem_reg[53][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][19]  ( .D(\Inst_Mem/inst_mem_reg[53][19] ), .CLK(clk), .RST(rst), .I(g_init[1715]), .Q(\Inst_Mem/inst_mem_reg[53][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][20]  ( .D(\Inst_Mem/inst_mem_reg[53][20] ), .CLK(clk), .RST(rst), .I(g_init[1716]), .Q(\Inst_Mem/inst_mem_reg[53][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][21]  ( .D(\Inst_Mem/inst_mem_reg[53][21] ), .CLK(clk), .RST(rst), .I(g_init[1717]), .Q(\Inst_Mem/inst_mem_reg[53][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][22]  ( .D(\Inst_Mem/inst_mem_reg[53][22] ), .CLK(clk), .RST(rst), .I(g_init[1718]), .Q(\Inst_Mem/inst_mem_reg[53][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][23]  ( .D(\Inst_Mem/inst_mem_reg[53][23] ), .CLK(clk), .RST(rst), .I(g_init[1719]), .Q(\Inst_Mem/inst_mem_reg[53][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][24]  ( .D(\Inst_Mem/inst_mem_reg[53][24] ), .CLK(clk), .RST(rst), .I(g_init[1720]), .Q(\Inst_Mem/inst_mem_reg[53][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][25]  ( .D(\Inst_Mem/inst_mem_reg[53][25] ), .CLK(clk), .RST(rst), .I(g_init[1721]), .Q(\Inst_Mem/inst_mem_reg[53][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][26]  ( .D(\Inst_Mem/inst_mem_reg[53][26] ), .CLK(clk), .RST(rst), .I(g_init[1722]), .Q(\Inst_Mem/inst_mem_reg[53][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][27]  ( .D(\Inst_Mem/inst_mem_reg[53][27] ), .CLK(clk), .RST(rst), .I(g_init[1723]), .Q(\Inst_Mem/inst_mem_reg[53][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][28]  ( .D(\Inst_Mem/inst_mem_reg[53][28] ), .CLK(clk), .RST(rst), .I(g_init[1724]), .Q(\Inst_Mem/inst_mem_reg[53][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][29]  ( .D(\Inst_Mem/inst_mem_reg[53][29] ), .CLK(clk), .RST(rst), .I(g_init[1725]), .Q(\Inst_Mem/inst_mem_reg[53][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][30]  ( .D(\Inst_Mem/inst_mem_reg[53][30] ), .CLK(clk), .RST(rst), .I(g_init[1726]), .Q(\Inst_Mem/inst_mem_reg[53][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[53][31]  ( .D(\Inst_Mem/inst_mem_reg[53][31] ), .CLK(clk), .RST(rst), .I(g_init[1727]), .Q(\Inst_Mem/inst_mem_reg[53][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][0]  ( .D(\Inst_Mem/inst_mem_reg[52][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1664]), .Q(
        \Inst_Mem/inst_mem_reg[52][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][1]  ( .D(\Inst_Mem/inst_mem_reg[52][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1665]), .Q(
        \Inst_Mem/inst_mem_reg[52][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][2]  ( .D(\Inst_Mem/inst_mem_reg[52][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1666]), .Q(
        \Inst_Mem/inst_mem_reg[52][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][3]  ( .D(\Inst_Mem/inst_mem_reg[52][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1667]), .Q(
        \Inst_Mem/inst_mem_reg[52][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][4]  ( .D(\Inst_Mem/inst_mem_reg[52][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1668]), .Q(
        \Inst_Mem/inst_mem_reg[52][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][5]  ( .D(\Inst_Mem/inst_mem_reg[52][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1669]), .Q(
        \Inst_Mem/inst_mem_reg[52][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][6]  ( .D(\Inst_Mem/inst_mem_reg[52][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1670]), .Q(
        \Inst_Mem/inst_mem_reg[52][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][7]  ( .D(\Inst_Mem/inst_mem_reg[52][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1671]), .Q(
        \Inst_Mem/inst_mem_reg[52][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][8]  ( .D(\Inst_Mem/inst_mem_reg[52][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1672]), .Q(
        \Inst_Mem/inst_mem_reg[52][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][9]  ( .D(\Inst_Mem/inst_mem_reg[52][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1673]), .Q(
        \Inst_Mem/inst_mem_reg[52][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[52][10]  ( .D(\Inst_Mem/inst_mem_reg[52][10] ), .CLK(clk), .RST(rst), .I(g_init[1674]), .Q(\Inst_Mem/inst_mem_reg[52][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][11]  ( .D(\Inst_Mem/inst_mem_reg[52][11] ), .CLK(clk), .RST(rst), .I(g_init[1675]), .Q(\Inst_Mem/inst_mem_reg[52][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][12]  ( .D(\Inst_Mem/inst_mem_reg[52][12] ), .CLK(clk), .RST(rst), .I(g_init[1676]), .Q(\Inst_Mem/inst_mem_reg[52][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][13]  ( .D(\Inst_Mem/inst_mem_reg[52][13] ), .CLK(clk), .RST(rst), .I(g_init[1677]), .Q(\Inst_Mem/inst_mem_reg[52][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][14]  ( .D(\Inst_Mem/inst_mem_reg[52][14] ), .CLK(clk), .RST(rst), .I(g_init[1678]), .Q(\Inst_Mem/inst_mem_reg[52][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][15]  ( .D(\Inst_Mem/inst_mem_reg[52][15] ), .CLK(clk), .RST(rst), .I(g_init[1679]), .Q(\Inst_Mem/inst_mem_reg[52][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][16]  ( .D(\Inst_Mem/inst_mem_reg[52][16] ), .CLK(clk), .RST(rst), .I(g_init[1680]), .Q(\Inst_Mem/inst_mem_reg[52][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][17]  ( .D(\Inst_Mem/inst_mem_reg[52][17] ), .CLK(clk), .RST(rst), .I(g_init[1681]), .Q(\Inst_Mem/inst_mem_reg[52][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][18]  ( .D(\Inst_Mem/inst_mem_reg[52][18] ), .CLK(clk), .RST(rst), .I(g_init[1682]), .Q(\Inst_Mem/inst_mem_reg[52][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][19]  ( .D(\Inst_Mem/inst_mem_reg[52][19] ), .CLK(clk), .RST(rst), .I(g_init[1683]), .Q(\Inst_Mem/inst_mem_reg[52][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][20]  ( .D(\Inst_Mem/inst_mem_reg[52][20] ), .CLK(clk), .RST(rst), .I(g_init[1684]), .Q(\Inst_Mem/inst_mem_reg[52][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][21]  ( .D(\Inst_Mem/inst_mem_reg[52][21] ), .CLK(clk), .RST(rst), .I(g_init[1685]), .Q(\Inst_Mem/inst_mem_reg[52][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][22]  ( .D(\Inst_Mem/inst_mem_reg[52][22] ), .CLK(clk), .RST(rst), .I(g_init[1686]), .Q(\Inst_Mem/inst_mem_reg[52][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][23]  ( .D(\Inst_Mem/inst_mem_reg[52][23] ), .CLK(clk), .RST(rst), .I(g_init[1687]), .Q(\Inst_Mem/inst_mem_reg[52][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][24]  ( .D(\Inst_Mem/inst_mem_reg[52][24] ), .CLK(clk), .RST(rst), .I(g_init[1688]), .Q(\Inst_Mem/inst_mem_reg[52][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][25]  ( .D(\Inst_Mem/inst_mem_reg[52][25] ), .CLK(clk), .RST(rst), .I(g_init[1689]), .Q(\Inst_Mem/inst_mem_reg[52][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][26]  ( .D(\Inst_Mem/inst_mem_reg[52][26] ), .CLK(clk), .RST(rst), .I(g_init[1690]), .Q(\Inst_Mem/inst_mem_reg[52][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][27]  ( .D(\Inst_Mem/inst_mem_reg[52][27] ), .CLK(clk), .RST(rst), .I(g_init[1691]), .Q(\Inst_Mem/inst_mem_reg[52][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][28]  ( .D(\Inst_Mem/inst_mem_reg[52][28] ), .CLK(clk), .RST(rst), .I(g_init[1692]), .Q(\Inst_Mem/inst_mem_reg[52][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][29]  ( .D(\Inst_Mem/inst_mem_reg[52][29] ), .CLK(clk), .RST(rst), .I(g_init[1693]), .Q(\Inst_Mem/inst_mem_reg[52][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][30]  ( .D(\Inst_Mem/inst_mem_reg[52][30] ), .CLK(clk), .RST(rst), .I(g_init[1694]), .Q(\Inst_Mem/inst_mem_reg[52][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[52][31]  ( .D(\Inst_Mem/inst_mem_reg[52][31] ), .CLK(clk), .RST(rst), .I(g_init[1695]), .Q(\Inst_Mem/inst_mem_reg[52][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][0]  ( .D(\Inst_Mem/inst_mem_reg[51][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1632]), .Q(
        \Inst_Mem/inst_mem_reg[51][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][1]  ( .D(\Inst_Mem/inst_mem_reg[51][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1633]), .Q(
        \Inst_Mem/inst_mem_reg[51][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][2]  ( .D(\Inst_Mem/inst_mem_reg[51][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1634]), .Q(
        \Inst_Mem/inst_mem_reg[51][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][3]  ( .D(\Inst_Mem/inst_mem_reg[51][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1635]), .Q(
        \Inst_Mem/inst_mem_reg[51][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][4]  ( .D(\Inst_Mem/inst_mem_reg[51][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1636]), .Q(
        \Inst_Mem/inst_mem_reg[51][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][5]  ( .D(\Inst_Mem/inst_mem_reg[51][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1637]), .Q(
        \Inst_Mem/inst_mem_reg[51][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][6]  ( .D(\Inst_Mem/inst_mem_reg[51][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1638]), .Q(
        \Inst_Mem/inst_mem_reg[51][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][7]  ( .D(\Inst_Mem/inst_mem_reg[51][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1639]), .Q(
        \Inst_Mem/inst_mem_reg[51][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][8]  ( .D(\Inst_Mem/inst_mem_reg[51][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1640]), .Q(
        \Inst_Mem/inst_mem_reg[51][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][9]  ( .D(\Inst_Mem/inst_mem_reg[51][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1641]), .Q(
        \Inst_Mem/inst_mem_reg[51][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[51][10]  ( .D(\Inst_Mem/inst_mem_reg[51][10] ), .CLK(clk), .RST(rst), .I(g_init[1642]), .Q(\Inst_Mem/inst_mem_reg[51][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][11]  ( .D(\Inst_Mem/inst_mem_reg[51][11] ), .CLK(clk), .RST(rst), .I(g_init[1643]), .Q(\Inst_Mem/inst_mem_reg[51][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][12]  ( .D(\Inst_Mem/inst_mem_reg[51][12] ), .CLK(clk), .RST(rst), .I(g_init[1644]), .Q(\Inst_Mem/inst_mem_reg[51][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][13]  ( .D(\Inst_Mem/inst_mem_reg[51][13] ), .CLK(clk), .RST(rst), .I(g_init[1645]), .Q(\Inst_Mem/inst_mem_reg[51][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][14]  ( .D(\Inst_Mem/inst_mem_reg[51][14] ), .CLK(clk), .RST(rst), .I(g_init[1646]), .Q(\Inst_Mem/inst_mem_reg[51][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][15]  ( .D(\Inst_Mem/inst_mem_reg[51][15] ), .CLK(clk), .RST(rst), .I(g_init[1647]), .Q(\Inst_Mem/inst_mem_reg[51][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][16]  ( .D(\Inst_Mem/inst_mem_reg[51][16] ), .CLK(clk), .RST(rst), .I(g_init[1648]), .Q(\Inst_Mem/inst_mem_reg[51][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][17]  ( .D(\Inst_Mem/inst_mem_reg[51][17] ), .CLK(clk), .RST(rst), .I(g_init[1649]), .Q(\Inst_Mem/inst_mem_reg[51][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][18]  ( .D(\Inst_Mem/inst_mem_reg[51][18] ), .CLK(clk), .RST(rst), .I(g_init[1650]), .Q(\Inst_Mem/inst_mem_reg[51][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][19]  ( .D(\Inst_Mem/inst_mem_reg[51][19] ), .CLK(clk), .RST(rst), .I(g_init[1651]), .Q(\Inst_Mem/inst_mem_reg[51][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][20]  ( .D(\Inst_Mem/inst_mem_reg[51][20] ), .CLK(clk), .RST(rst), .I(g_init[1652]), .Q(\Inst_Mem/inst_mem_reg[51][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][21]  ( .D(\Inst_Mem/inst_mem_reg[51][21] ), .CLK(clk), .RST(rst), .I(g_init[1653]), .Q(\Inst_Mem/inst_mem_reg[51][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][22]  ( .D(\Inst_Mem/inst_mem_reg[51][22] ), .CLK(clk), .RST(rst), .I(g_init[1654]), .Q(\Inst_Mem/inst_mem_reg[51][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][23]  ( .D(\Inst_Mem/inst_mem_reg[51][23] ), .CLK(clk), .RST(rst), .I(g_init[1655]), .Q(\Inst_Mem/inst_mem_reg[51][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][24]  ( .D(\Inst_Mem/inst_mem_reg[51][24] ), .CLK(clk), .RST(rst), .I(g_init[1656]), .Q(\Inst_Mem/inst_mem_reg[51][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][25]  ( .D(\Inst_Mem/inst_mem_reg[51][25] ), .CLK(clk), .RST(rst), .I(g_init[1657]), .Q(\Inst_Mem/inst_mem_reg[51][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][26]  ( .D(\Inst_Mem/inst_mem_reg[51][26] ), .CLK(clk), .RST(rst), .I(g_init[1658]), .Q(\Inst_Mem/inst_mem_reg[51][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][27]  ( .D(\Inst_Mem/inst_mem_reg[51][27] ), .CLK(clk), .RST(rst), .I(g_init[1659]), .Q(\Inst_Mem/inst_mem_reg[51][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][28]  ( .D(\Inst_Mem/inst_mem_reg[51][28] ), .CLK(clk), .RST(rst), .I(g_init[1660]), .Q(\Inst_Mem/inst_mem_reg[51][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][29]  ( .D(\Inst_Mem/inst_mem_reg[51][29] ), .CLK(clk), .RST(rst), .I(g_init[1661]), .Q(\Inst_Mem/inst_mem_reg[51][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][30]  ( .D(\Inst_Mem/inst_mem_reg[51][30] ), .CLK(clk), .RST(rst), .I(g_init[1662]), .Q(\Inst_Mem/inst_mem_reg[51][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[51][31]  ( .D(\Inst_Mem/inst_mem_reg[51][31] ), .CLK(clk), .RST(rst), .I(g_init[1663]), .Q(\Inst_Mem/inst_mem_reg[51][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][0]  ( .D(\Inst_Mem/inst_mem_reg[50][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1600]), .Q(
        \Inst_Mem/inst_mem_reg[50][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][1]  ( .D(\Inst_Mem/inst_mem_reg[50][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1601]), .Q(
        \Inst_Mem/inst_mem_reg[50][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][2]  ( .D(\Inst_Mem/inst_mem_reg[50][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1602]), .Q(
        \Inst_Mem/inst_mem_reg[50][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][3]  ( .D(\Inst_Mem/inst_mem_reg[50][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1603]), .Q(
        \Inst_Mem/inst_mem_reg[50][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][4]  ( .D(\Inst_Mem/inst_mem_reg[50][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1604]), .Q(
        \Inst_Mem/inst_mem_reg[50][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][5]  ( .D(\Inst_Mem/inst_mem_reg[50][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1605]), .Q(
        \Inst_Mem/inst_mem_reg[50][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][6]  ( .D(\Inst_Mem/inst_mem_reg[50][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1606]), .Q(
        \Inst_Mem/inst_mem_reg[50][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][7]  ( .D(\Inst_Mem/inst_mem_reg[50][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1607]), .Q(
        \Inst_Mem/inst_mem_reg[50][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][8]  ( .D(\Inst_Mem/inst_mem_reg[50][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1608]), .Q(
        \Inst_Mem/inst_mem_reg[50][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][9]  ( .D(\Inst_Mem/inst_mem_reg[50][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1609]), .Q(
        \Inst_Mem/inst_mem_reg[50][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[50][10]  ( .D(\Inst_Mem/inst_mem_reg[50][10] ), .CLK(clk), .RST(rst), .I(g_init[1610]), .Q(\Inst_Mem/inst_mem_reg[50][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][11]  ( .D(\Inst_Mem/inst_mem_reg[50][11] ), .CLK(clk), .RST(rst), .I(g_init[1611]), .Q(\Inst_Mem/inst_mem_reg[50][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][12]  ( .D(\Inst_Mem/inst_mem_reg[50][12] ), .CLK(clk), .RST(rst), .I(g_init[1612]), .Q(\Inst_Mem/inst_mem_reg[50][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][13]  ( .D(\Inst_Mem/inst_mem_reg[50][13] ), .CLK(clk), .RST(rst), .I(g_init[1613]), .Q(\Inst_Mem/inst_mem_reg[50][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][14]  ( .D(\Inst_Mem/inst_mem_reg[50][14] ), .CLK(clk), .RST(rst), .I(g_init[1614]), .Q(\Inst_Mem/inst_mem_reg[50][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][15]  ( .D(\Inst_Mem/inst_mem_reg[50][15] ), .CLK(clk), .RST(rst), .I(g_init[1615]), .Q(\Inst_Mem/inst_mem_reg[50][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][16]  ( .D(\Inst_Mem/inst_mem_reg[50][16] ), .CLK(clk), .RST(rst), .I(g_init[1616]), .Q(\Inst_Mem/inst_mem_reg[50][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][17]  ( .D(\Inst_Mem/inst_mem_reg[50][17] ), .CLK(clk), .RST(rst), .I(g_init[1617]), .Q(\Inst_Mem/inst_mem_reg[50][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][18]  ( .D(\Inst_Mem/inst_mem_reg[50][18] ), .CLK(clk), .RST(rst), .I(g_init[1618]), .Q(\Inst_Mem/inst_mem_reg[50][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][19]  ( .D(\Inst_Mem/inst_mem_reg[50][19] ), .CLK(clk), .RST(rst), .I(g_init[1619]), .Q(\Inst_Mem/inst_mem_reg[50][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][20]  ( .D(\Inst_Mem/inst_mem_reg[50][20] ), .CLK(clk), .RST(rst), .I(g_init[1620]), .Q(\Inst_Mem/inst_mem_reg[50][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][21]  ( .D(\Inst_Mem/inst_mem_reg[50][21] ), .CLK(clk), .RST(rst), .I(g_init[1621]), .Q(\Inst_Mem/inst_mem_reg[50][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][22]  ( .D(\Inst_Mem/inst_mem_reg[50][22] ), .CLK(clk), .RST(rst), .I(g_init[1622]), .Q(\Inst_Mem/inst_mem_reg[50][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][23]  ( .D(\Inst_Mem/inst_mem_reg[50][23] ), .CLK(clk), .RST(rst), .I(g_init[1623]), .Q(\Inst_Mem/inst_mem_reg[50][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][24]  ( .D(\Inst_Mem/inst_mem_reg[50][24] ), .CLK(clk), .RST(rst), .I(g_init[1624]), .Q(\Inst_Mem/inst_mem_reg[50][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][25]  ( .D(\Inst_Mem/inst_mem_reg[50][25] ), .CLK(clk), .RST(rst), .I(g_init[1625]), .Q(\Inst_Mem/inst_mem_reg[50][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][26]  ( .D(\Inst_Mem/inst_mem_reg[50][26] ), .CLK(clk), .RST(rst), .I(g_init[1626]), .Q(\Inst_Mem/inst_mem_reg[50][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][27]  ( .D(\Inst_Mem/inst_mem_reg[50][27] ), .CLK(clk), .RST(rst), .I(g_init[1627]), .Q(\Inst_Mem/inst_mem_reg[50][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][28]  ( .D(\Inst_Mem/inst_mem_reg[50][28] ), .CLK(clk), .RST(rst), .I(g_init[1628]), .Q(\Inst_Mem/inst_mem_reg[50][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][29]  ( .D(\Inst_Mem/inst_mem_reg[50][29] ), .CLK(clk), .RST(rst), .I(g_init[1629]), .Q(\Inst_Mem/inst_mem_reg[50][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][30]  ( .D(\Inst_Mem/inst_mem_reg[50][30] ), .CLK(clk), .RST(rst), .I(g_init[1630]), .Q(\Inst_Mem/inst_mem_reg[50][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[50][31]  ( .D(\Inst_Mem/inst_mem_reg[50][31] ), .CLK(clk), .RST(rst), .I(g_init[1631]), .Q(\Inst_Mem/inst_mem_reg[50][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][0]  ( .D(\Inst_Mem/inst_mem_reg[49][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1568]), .Q(
        \Inst_Mem/inst_mem_reg[49][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][1]  ( .D(\Inst_Mem/inst_mem_reg[49][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1569]), .Q(
        \Inst_Mem/inst_mem_reg[49][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][2]  ( .D(\Inst_Mem/inst_mem_reg[49][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1570]), .Q(
        \Inst_Mem/inst_mem_reg[49][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][3]  ( .D(\Inst_Mem/inst_mem_reg[49][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1571]), .Q(
        \Inst_Mem/inst_mem_reg[49][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][4]  ( .D(\Inst_Mem/inst_mem_reg[49][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1572]), .Q(
        \Inst_Mem/inst_mem_reg[49][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][5]  ( .D(\Inst_Mem/inst_mem_reg[49][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1573]), .Q(
        \Inst_Mem/inst_mem_reg[49][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][6]  ( .D(\Inst_Mem/inst_mem_reg[49][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1574]), .Q(
        \Inst_Mem/inst_mem_reg[49][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][7]  ( .D(\Inst_Mem/inst_mem_reg[49][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1575]), .Q(
        \Inst_Mem/inst_mem_reg[49][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][8]  ( .D(\Inst_Mem/inst_mem_reg[49][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1576]), .Q(
        \Inst_Mem/inst_mem_reg[49][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][9]  ( .D(\Inst_Mem/inst_mem_reg[49][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1577]), .Q(
        \Inst_Mem/inst_mem_reg[49][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[49][10]  ( .D(\Inst_Mem/inst_mem_reg[49][10] ), .CLK(clk), .RST(rst), .I(g_init[1578]), .Q(\Inst_Mem/inst_mem_reg[49][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][11]  ( .D(\Inst_Mem/inst_mem_reg[49][11] ), .CLK(clk), .RST(rst), .I(g_init[1579]), .Q(\Inst_Mem/inst_mem_reg[49][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][12]  ( .D(\Inst_Mem/inst_mem_reg[49][12] ), .CLK(clk), .RST(rst), .I(g_init[1580]), .Q(\Inst_Mem/inst_mem_reg[49][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][13]  ( .D(\Inst_Mem/inst_mem_reg[49][13] ), .CLK(clk), .RST(rst), .I(g_init[1581]), .Q(\Inst_Mem/inst_mem_reg[49][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][14]  ( .D(\Inst_Mem/inst_mem_reg[49][14] ), .CLK(clk), .RST(rst), .I(g_init[1582]), .Q(\Inst_Mem/inst_mem_reg[49][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][15]  ( .D(\Inst_Mem/inst_mem_reg[49][15] ), .CLK(clk), .RST(rst), .I(g_init[1583]), .Q(\Inst_Mem/inst_mem_reg[49][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][16]  ( .D(\Inst_Mem/inst_mem_reg[49][16] ), .CLK(clk), .RST(rst), .I(g_init[1584]), .Q(\Inst_Mem/inst_mem_reg[49][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][17]  ( .D(\Inst_Mem/inst_mem_reg[49][17] ), .CLK(clk), .RST(rst), .I(g_init[1585]), .Q(\Inst_Mem/inst_mem_reg[49][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][18]  ( .D(\Inst_Mem/inst_mem_reg[49][18] ), .CLK(clk), .RST(rst), .I(g_init[1586]), .Q(\Inst_Mem/inst_mem_reg[49][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][19]  ( .D(\Inst_Mem/inst_mem_reg[49][19] ), .CLK(clk), .RST(rst), .I(g_init[1587]), .Q(\Inst_Mem/inst_mem_reg[49][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][20]  ( .D(\Inst_Mem/inst_mem_reg[49][20] ), .CLK(clk), .RST(rst), .I(g_init[1588]), .Q(\Inst_Mem/inst_mem_reg[49][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][21]  ( .D(\Inst_Mem/inst_mem_reg[49][21] ), .CLK(clk), .RST(rst), .I(g_init[1589]), .Q(\Inst_Mem/inst_mem_reg[49][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][22]  ( .D(\Inst_Mem/inst_mem_reg[49][22] ), .CLK(clk), .RST(rst), .I(g_init[1590]), .Q(\Inst_Mem/inst_mem_reg[49][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][23]  ( .D(\Inst_Mem/inst_mem_reg[49][23] ), .CLK(clk), .RST(rst), .I(g_init[1591]), .Q(\Inst_Mem/inst_mem_reg[49][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][24]  ( .D(\Inst_Mem/inst_mem_reg[49][24] ), .CLK(clk), .RST(rst), .I(g_init[1592]), .Q(\Inst_Mem/inst_mem_reg[49][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][25]  ( .D(\Inst_Mem/inst_mem_reg[49][25] ), .CLK(clk), .RST(rst), .I(g_init[1593]), .Q(\Inst_Mem/inst_mem_reg[49][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][26]  ( .D(\Inst_Mem/inst_mem_reg[49][26] ), .CLK(clk), .RST(rst), .I(g_init[1594]), .Q(\Inst_Mem/inst_mem_reg[49][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][27]  ( .D(\Inst_Mem/inst_mem_reg[49][27] ), .CLK(clk), .RST(rst), .I(g_init[1595]), .Q(\Inst_Mem/inst_mem_reg[49][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][28]  ( .D(\Inst_Mem/inst_mem_reg[49][28] ), .CLK(clk), .RST(rst), .I(g_init[1596]), .Q(\Inst_Mem/inst_mem_reg[49][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][29]  ( .D(\Inst_Mem/inst_mem_reg[49][29] ), .CLK(clk), .RST(rst), .I(g_init[1597]), .Q(\Inst_Mem/inst_mem_reg[49][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][30]  ( .D(\Inst_Mem/inst_mem_reg[49][30] ), .CLK(clk), .RST(rst), .I(g_init[1598]), .Q(\Inst_Mem/inst_mem_reg[49][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[49][31]  ( .D(\Inst_Mem/inst_mem_reg[49][31] ), .CLK(clk), .RST(rst), .I(g_init[1599]), .Q(\Inst_Mem/inst_mem_reg[49][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][0]  ( .D(\Inst_Mem/inst_mem_reg[48][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1536]), .Q(
        \Inst_Mem/inst_mem_reg[48][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][1]  ( .D(\Inst_Mem/inst_mem_reg[48][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1537]), .Q(
        \Inst_Mem/inst_mem_reg[48][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][2]  ( .D(\Inst_Mem/inst_mem_reg[48][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1538]), .Q(
        \Inst_Mem/inst_mem_reg[48][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][3]  ( .D(\Inst_Mem/inst_mem_reg[48][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1539]), .Q(
        \Inst_Mem/inst_mem_reg[48][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][4]  ( .D(\Inst_Mem/inst_mem_reg[48][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1540]), .Q(
        \Inst_Mem/inst_mem_reg[48][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][5]  ( .D(\Inst_Mem/inst_mem_reg[48][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1541]), .Q(
        \Inst_Mem/inst_mem_reg[48][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][6]  ( .D(\Inst_Mem/inst_mem_reg[48][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1542]), .Q(
        \Inst_Mem/inst_mem_reg[48][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][7]  ( .D(\Inst_Mem/inst_mem_reg[48][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1543]), .Q(
        \Inst_Mem/inst_mem_reg[48][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][8]  ( .D(\Inst_Mem/inst_mem_reg[48][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1544]), .Q(
        \Inst_Mem/inst_mem_reg[48][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][9]  ( .D(\Inst_Mem/inst_mem_reg[48][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1545]), .Q(
        \Inst_Mem/inst_mem_reg[48][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[48][10]  ( .D(\Inst_Mem/inst_mem_reg[48][10] ), .CLK(clk), .RST(rst), .I(g_init[1546]), .Q(\Inst_Mem/inst_mem_reg[48][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][11]  ( .D(\Inst_Mem/inst_mem_reg[48][11] ), .CLK(clk), .RST(rst), .I(g_init[1547]), .Q(\Inst_Mem/inst_mem_reg[48][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][12]  ( .D(\Inst_Mem/inst_mem_reg[48][12] ), .CLK(clk), .RST(rst), .I(g_init[1548]), .Q(\Inst_Mem/inst_mem_reg[48][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][13]  ( .D(\Inst_Mem/inst_mem_reg[48][13] ), .CLK(clk), .RST(rst), .I(g_init[1549]), .Q(\Inst_Mem/inst_mem_reg[48][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][14]  ( .D(\Inst_Mem/inst_mem_reg[48][14] ), .CLK(clk), .RST(rst), .I(g_init[1550]), .Q(\Inst_Mem/inst_mem_reg[48][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][15]  ( .D(\Inst_Mem/inst_mem_reg[48][15] ), .CLK(clk), .RST(rst), .I(g_init[1551]), .Q(\Inst_Mem/inst_mem_reg[48][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][16]  ( .D(\Inst_Mem/inst_mem_reg[48][16] ), .CLK(clk), .RST(rst), .I(g_init[1552]), .Q(\Inst_Mem/inst_mem_reg[48][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][17]  ( .D(\Inst_Mem/inst_mem_reg[48][17] ), .CLK(clk), .RST(rst), .I(g_init[1553]), .Q(\Inst_Mem/inst_mem_reg[48][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][18]  ( .D(\Inst_Mem/inst_mem_reg[48][18] ), .CLK(clk), .RST(rst), .I(g_init[1554]), .Q(\Inst_Mem/inst_mem_reg[48][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][19]  ( .D(\Inst_Mem/inst_mem_reg[48][19] ), .CLK(clk), .RST(rst), .I(g_init[1555]), .Q(\Inst_Mem/inst_mem_reg[48][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][20]  ( .D(\Inst_Mem/inst_mem_reg[48][20] ), .CLK(clk), .RST(rst), .I(g_init[1556]), .Q(\Inst_Mem/inst_mem_reg[48][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][21]  ( .D(\Inst_Mem/inst_mem_reg[48][21] ), .CLK(clk), .RST(rst), .I(g_init[1557]), .Q(\Inst_Mem/inst_mem_reg[48][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][22]  ( .D(\Inst_Mem/inst_mem_reg[48][22] ), .CLK(clk), .RST(rst), .I(g_init[1558]), .Q(\Inst_Mem/inst_mem_reg[48][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][23]  ( .D(\Inst_Mem/inst_mem_reg[48][23] ), .CLK(clk), .RST(rst), .I(g_init[1559]), .Q(\Inst_Mem/inst_mem_reg[48][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][24]  ( .D(\Inst_Mem/inst_mem_reg[48][24] ), .CLK(clk), .RST(rst), .I(g_init[1560]), .Q(\Inst_Mem/inst_mem_reg[48][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][25]  ( .D(\Inst_Mem/inst_mem_reg[48][25] ), .CLK(clk), .RST(rst), .I(g_init[1561]), .Q(\Inst_Mem/inst_mem_reg[48][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][26]  ( .D(\Inst_Mem/inst_mem_reg[48][26] ), .CLK(clk), .RST(rst), .I(g_init[1562]), .Q(\Inst_Mem/inst_mem_reg[48][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][27]  ( .D(\Inst_Mem/inst_mem_reg[48][27] ), .CLK(clk), .RST(rst), .I(g_init[1563]), .Q(\Inst_Mem/inst_mem_reg[48][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][28]  ( .D(\Inst_Mem/inst_mem_reg[48][28] ), .CLK(clk), .RST(rst), .I(g_init[1564]), .Q(\Inst_Mem/inst_mem_reg[48][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][29]  ( .D(\Inst_Mem/inst_mem_reg[48][29] ), .CLK(clk), .RST(rst), .I(g_init[1565]), .Q(\Inst_Mem/inst_mem_reg[48][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][30]  ( .D(\Inst_Mem/inst_mem_reg[48][30] ), .CLK(clk), .RST(rst), .I(g_init[1566]), .Q(\Inst_Mem/inst_mem_reg[48][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[48][31]  ( .D(\Inst_Mem/inst_mem_reg[48][31] ), .CLK(clk), .RST(rst), .I(g_init[1567]), .Q(\Inst_Mem/inst_mem_reg[48][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][0]  ( .D(\Inst_Mem/inst_mem_reg[47][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1504]), .Q(
        \Inst_Mem/inst_mem_reg[47][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][1]  ( .D(\Inst_Mem/inst_mem_reg[47][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1505]), .Q(
        \Inst_Mem/inst_mem_reg[47][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][2]  ( .D(\Inst_Mem/inst_mem_reg[47][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1506]), .Q(
        \Inst_Mem/inst_mem_reg[47][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][3]  ( .D(\Inst_Mem/inst_mem_reg[47][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1507]), .Q(
        \Inst_Mem/inst_mem_reg[47][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][4]  ( .D(\Inst_Mem/inst_mem_reg[47][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1508]), .Q(
        \Inst_Mem/inst_mem_reg[47][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][5]  ( .D(\Inst_Mem/inst_mem_reg[47][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1509]), .Q(
        \Inst_Mem/inst_mem_reg[47][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][6]  ( .D(\Inst_Mem/inst_mem_reg[47][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1510]), .Q(
        \Inst_Mem/inst_mem_reg[47][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][7]  ( .D(\Inst_Mem/inst_mem_reg[47][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1511]), .Q(
        \Inst_Mem/inst_mem_reg[47][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][8]  ( .D(\Inst_Mem/inst_mem_reg[47][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1512]), .Q(
        \Inst_Mem/inst_mem_reg[47][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][9]  ( .D(\Inst_Mem/inst_mem_reg[47][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1513]), .Q(
        \Inst_Mem/inst_mem_reg[47][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[47][10]  ( .D(\Inst_Mem/inst_mem_reg[47][10] ), .CLK(clk), .RST(rst), .I(g_init[1514]), .Q(\Inst_Mem/inst_mem_reg[47][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][11]  ( .D(\Inst_Mem/inst_mem_reg[47][11] ), .CLK(clk), .RST(rst), .I(g_init[1515]), .Q(\Inst_Mem/inst_mem_reg[47][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][12]  ( .D(\Inst_Mem/inst_mem_reg[47][12] ), .CLK(clk), .RST(rst), .I(g_init[1516]), .Q(\Inst_Mem/inst_mem_reg[47][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][13]  ( .D(\Inst_Mem/inst_mem_reg[47][13] ), .CLK(clk), .RST(rst), .I(g_init[1517]), .Q(\Inst_Mem/inst_mem_reg[47][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][14]  ( .D(\Inst_Mem/inst_mem_reg[47][14] ), .CLK(clk), .RST(rst), .I(g_init[1518]), .Q(\Inst_Mem/inst_mem_reg[47][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][15]  ( .D(\Inst_Mem/inst_mem_reg[47][15] ), .CLK(clk), .RST(rst), .I(g_init[1519]), .Q(\Inst_Mem/inst_mem_reg[47][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][16]  ( .D(\Inst_Mem/inst_mem_reg[47][16] ), .CLK(clk), .RST(rst), .I(g_init[1520]), .Q(\Inst_Mem/inst_mem_reg[47][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][17]  ( .D(\Inst_Mem/inst_mem_reg[47][17] ), .CLK(clk), .RST(rst), .I(g_init[1521]), .Q(\Inst_Mem/inst_mem_reg[47][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][18]  ( .D(\Inst_Mem/inst_mem_reg[47][18] ), .CLK(clk), .RST(rst), .I(g_init[1522]), .Q(\Inst_Mem/inst_mem_reg[47][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][19]  ( .D(\Inst_Mem/inst_mem_reg[47][19] ), .CLK(clk), .RST(rst), .I(g_init[1523]), .Q(\Inst_Mem/inst_mem_reg[47][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][20]  ( .D(\Inst_Mem/inst_mem_reg[47][20] ), .CLK(clk), .RST(rst), .I(g_init[1524]), .Q(\Inst_Mem/inst_mem_reg[47][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][21]  ( .D(\Inst_Mem/inst_mem_reg[47][21] ), .CLK(clk), .RST(rst), .I(g_init[1525]), .Q(\Inst_Mem/inst_mem_reg[47][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][22]  ( .D(\Inst_Mem/inst_mem_reg[47][22] ), .CLK(clk), .RST(rst), .I(g_init[1526]), .Q(\Inst_Mem/inst_mem_reg[47][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][23]  ( .D(\Inst_Mem/inst_mem_reg[47][23] ), .CLK(clk), .RST(rst), .I(g_init[1527]), .Q(\Inst_Mem/inst_mem_reg[47][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][24]  ( .D(\Inst_Mem/inst_mem_reg[47][24] ), .CLK(clk), .RST(rst), .I(g_init[1528]), .Q(\Inst_Mem/inst_mem_reg[47][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][25]  ( .D(\Inst_Mem/inst_mem_reg[47][25] ), .CLK(clk), .RST(rst), .I(g_init[1529]), .Q(\Inst_Mem/inst_mem_reg[47][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][26]  ( .D(\Inst_Mem/inst_mem_reg[47][26] ), .CLK(clk), .RST(rst), .I(g_init[1530]), .Q(\Inst_Mem/inst_mem_reg[47][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][27]  ( .D(\Inst_Mem/inst_mem_reg[47][27] ), .CLK(clk), .RST(rst), .I(g_init[1531]), .Q(\Inst_Mem/inst_mem_reg[47][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][28]  ( .D(\Inst_Mem/inst_mem_reg[47][28] ), .CLK(clk), .RST(rst), .I(g_init[1532]), .Q(\Inst_Mem/inst_mem_reg[47][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][29]  ( .D(\Inst_Mem/inst_mem_reg[47][29] ), .CLK(clk), .RST(rst), .I(g_init[1533]), .Q(\Inst_Mem/inst_mem_reg[47][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][30]  ( .D(\Inst_Mem/inst_mem_reg[47][30] ), .CLK(clk), .RST(rst), .I(g_init[1534]), .Q(\Inst_Mem/inst_mem_reg[47][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[47][31]  ( .D(\Inst_Mem/inst_mem_reg[47][31] ), .CLK(clk), .RST(rst), .I(g_init[1535]), .Q(\Inst_Mem/inst_mem_reg[47][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][0]  ( .D(\Inst_Mem/inst_mem_reg[46][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1472]), .Q(
        \Inst_Mem/inst_mem_reg[46][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][1]  ( .D(\Inst_Mem/inst_mem_reg[46][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1473]), .Q(
        \Inst_Mem/inst_mem_reg[46][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][2]  ( .D(\Inst_Mem/inst_mem_reg[46][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1474]), .Q(
        \Inst_Mem/inst_mem_reg[46][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][3]  ( .D(\Inst_Mem/inst_mem_reg[46][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1475]), .Q(
        \Inst_Mem/inst_mem_reg[46][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][4]  ( .D(\Inst_Mem/inst_mem_reg[46][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1476]), .Q(
        \Inst_Mem/inst_mem_reg[46][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][5]  ( .D(\Inst_Mem/inst_mem_reg[46][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1477]), .Q(
        \Inst_Mem/inst_mem_reg[46][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][6]  ( .D(\Inst_Mem/inst_mem_reg[46][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1478]), .Q(
        \Inst_Mem/inst_mem_reg[46][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][7]  ( .D(\Inst_Mem/inst_mem_reg[46][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1479]), .Q(
        \Inst_Mem/inst_mem_reg[46][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][8]  ( .D(\Inst_Mem/inst_mem_reg[46][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1480]), .Q(
        \Inst_Mem/inst_mem_reg[46][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][9]  ( .D(\Inst_Mem/inst_mem_reg[46][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1481]), .Q(
        \Inst_Mem/inst_mem_reg[46][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[46][10]  ( .D(\Inst_Mem/inst_mem_reg[46][10] ), .CLK(clk), .RST(rst), .I(g_init[1482]), .Q(\Inst_Mem/inst_mem_reg[46][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][11]  ( .D(\Inst_Mem/inst_mem_reg[46][11] ), .CLK(clk), .RST(rst), .I(g_init[1483]), .Q(\Inst_Mem/inst_mem_reg[46][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][12]  ( .D(\Inst_Mem/inst_mem_reg[46][12] ), .CLK(clk), .RST(rst), .I(g_init[1484]), .Q(\Inst_Mem/inst_mem_reg[46][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][13]  ( .D(\Inst_Mem/inst_mem_reg[46][13] ), .CLK(clk), .RST(rst), .I(g_init[1485]), .Q(\Inst_Mem/inst_mem_reg[46][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][14]  ( .D(\Inst_Mem/inst_mem_reg[46][14] ), .CLK(clk), .RST(rst), .I(g_init[1486]), .Q(\Inst_Mem/inst_mem_reg[46][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][15]  ( .D(\Inst_Mem/inst_mem_reg[46][15] ), .CLK(clk), .RST(rst), .I(g_init[1487]), .Q(\Inst_Mem/inst_mem_reg[46][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][16]  ( .D(\Inst_Mem/inst_mem_reg[46][16] ), .CLK(clk), .RST(rst), .I(g_init[1488]), .Q(\Inst_Mem/inst_mem_reg[46][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][17]  ( .D(\Inst_Mem/inst_mem_reg[46][17] ), .CLK(clk), .RST(rst), .I(g_init[1489]), .Q(\Inst_Mem/inst_mem_reg[46][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][18]  ( .D(\Inst_Mem/inst_mem_reg[46][18] ), .CLK(clk), .RST(rst), .I(g_init[1490]), .Q(\Inst_Mem/inst_mem_reg[46][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][19]  ( .D(\Inst_Mem/inst_mem_reg[46][19] ), .CLK(clk), .RST(rst), .I(g_init[1491]), .Q(\Inst_Mem/inst_mem_reg[46][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][20]  ( .D(\Inst_Mem/inst_mem_reg[46][20] ), .CLK(clk), .RST(rst), .I(g_init[1492]), .Q(\Inst_Mem/inst_mem_reg[46][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][21]  ( .D(\Inst_Mem/inst_mem_reg[46][21] ), .CLK(clk), .RST(rst), .I(g_init[1493]), .Q(\Inst_Mem/inst_mem_reg[46][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][22]  ( .D(\Inst_Mem/inst_mem_reg[46][22] ), .CLK(clk), .RST(rst), .I(g_init[1494]), .Q(\Inst_Mem/inst_mem_reg[46][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][23]  ( .D(\Inst_Mem/inst_mem_reg[46][23] ), .CLK(clk), .RST(rst), .I(g_init[1495]), .Q(\Inst_Mem/inst_mem_reg[46][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][24]  ( .D(\Inst_Mem/inst_mem_reg[46][24] ), .CLK(clk), .RST(rst), .I(g_init[1496]), .Q(\Inst_Mem/inst_mem_reg[46][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][25]  ( .D(\Inst_Mem/inst_mem_reg[46][25] ), .CLK(clk), .RST(rst), .I(g_init[1497]), .Q(\Inst_Mem/inst_mem_reg[46][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][26]  ( .D(\Inst_Mem/inst_mem_reg[46][26] ), .CLK(clk), .RST(rst), .I(g_init[1498]), .Q(\Inst_Mem/inst_mem_reg[46][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][27]  ( .D(\Inst_Mem/inst_mem_reg[46][27] ), .CLK(clk), .RST(rst), .I(g_init[1499]), .Q(\Inst_Mem/inst_mem_reg[46][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][28]  ( .D(\Inst_Mem/inst_mem_reg[46][28] ), .CLK(clk), .RST(rst), .I(g_init[1500]), .Q(\Inst_Mem/inst_mem_reg[46][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][29]  ( .D(\Inst_Mem/inst_mem_reg[46][29] ), .CLK(clk), .RST(rst), .I(g_init[1501]), .Q(\Inst_Mem/inst_mem_reg[46][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][30]  ( .D(\Inst_Mem/inst_mem_reg[46][30] ), .CLK(clk), .RST(rst), .I(g_init[1502]), .Q(\Inst_Mem/inst_mem_reg[46][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[46][31]  ( .D(\Inst_Mem/inst_mem_reg[46][31] ), .CLK(clk), .RST(rst), .I(g_init[1503]), .Q(\Inst_Mem/inst_mem_reg[46][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][0]  ( .D(\Inst_Mem/inst_mem_reg[45][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1440]), .Q(
        \Inst_Mem/inst_mem_reg[45][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][1]  ( .D(\Inst_Mem/inst_mem_reg[45][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1441]), .Q(
        \Inst_Mem/inst_mem_reg[45][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][2]  ( .D(\Inst_Mem/inst_mem_reg[45][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1442]), .Q(
        \Inst_Mem/inst_mem_reg[45][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][3]  ( .D(\Inst_Mem/inst_mem_reg[45][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1443]), .Q(
        \Inst_Mem/inst_mem_reg[45][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][4]  ( .D(\Inst_Mem/inst_mem_reg[45][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1444]), .Q(
        \Inst_Mem/inst_mem_reg[45][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][5]  ( .D(\Inst_Mem/inst_mem_reg[45][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1445]), .Q(
        \Inst_Mem/inst_mem_reg[45][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][6]  ( .D(\Inst_Mem/inst_mem_reg[45][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1446]), .Q(
        \Inst_Mem/inst_mem_reg[45][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][7]  ( .D(\Inst_Mem/inst_mem_reg[45][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1447]), .Q(
        \Inst_Mem/inst_mem_reg[45][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][8]  ( .D(\Inst_Mem/inst_mem_reg[45][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1448]), .Q(
        \Inst_Mem/inst_mem_reg[45][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][9]  ( .D(\Inst_Mem/inst_mem_reg[45][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1449]), .Q(
        \Inst_Mem/inst_mem_reg[45][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[45][10]  ( .D(\Inst_Mem/inst_mem_reg[45][10] ), .CLK(clk), .RST(rst), .I(g_init[1450]), .Q(\Inst_Mem/inst_mem_reg[45][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][11]  ( .D(\Inst_Mem/inst_mem_reg[45][11] ), .CLK(clk), .RST(rst), .I(g_init[1451]), .Q(\Inst_Mem/inst_mem_reg[45][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][12]  ( .D(\Inst_Mem/inst_mem_reg[45][12] ), .CLK(clk), .RST(rst), .I(g_init[1452]), .Q(\Inst_Mem/inst_mem_reg[45][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][13]  ( .D(\Inst_Mem/inst_mem_reg[45][13] ), .CLK(clk), .RST(rst), .I(g_init[1453]), .Q(\Inst_Mem/inst_mem_reg[45][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][14]  ( .D(\Inst_Mem/inst_mem_reg[45][14] ), .CLK(clk), .RST(rst), .I(g_init[1454]), .Q(\Inst_Mem/inst_mem_reg[45][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][15]  ( .D(\Inst_Mem/inst_mem_reg[45][15] ), .CLK(clk), .RST(rst), .I(g_init[1455]), .Q(\Inst_Mem/inst_mem_reg[45][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][16]  ( .D(\Inst_Mem/inst_mem_reg[45][16] ), .CLK(clk), .RST(rst), .I(g_init[1456]), .Q(\Inst_Mem/inst_mem_reg[45][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][17]  ( .D(\Inst_Mem/inst_mem_reg[45][17] ), .CLK(clk), .RST(rst), .I(g_init[1457]), .Q(\Inst_Mem/inst_mem_reg[45][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][18]  ( .D(\Inst_Mem/inst_mem_reg[45][18] ), .CLK(clk), .RST(rst), .I(g_init[1458]), .Q(\Inst_Mem/inst_mem_reg[45][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][19]  ( .D(\Inst_Mem/inst_mem_reg[45][19] ), .CLK(clk), .RST(rst), .I(g_init[1459]), .Q(\Inst_Mem/inst_mem_reg[45][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][20]  ( .D(\Inst_Mem/inst_mem_reg[45][20] ), .CLK(clk), .RST(rst), .I(g_init[1460]), .Q(\Inst_Mem/inst_mem_reg[45][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][21]  ( .D(\Inst_Mem/inst_mem_reg[45][21] ), .CLK(clk), .RST(rst), .I(g_init[1461]), .Q(\Inst_Mem/inst_mem_reg[45][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][22]  ( .D(\Inst_Mem/inst_mem_reg[45][22] ), .CLK(clk), .RST(rst), .I(g_init[1462]), .Q(\Inst_Mem/inst_mem_reg[45][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][23]  ( .D(\Inst_Mem/inst_mem_reg[45][23] ), .CLK(clk), .RST(rst), .I(g_init[1463]), .Q(\Inst_Mem/inst_mem_reg[45][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][24]  ( .D(\Inst_Mem/inst_mem_reg[45][24] ), .CLK(clk), .RST(rst), .I(g_init[1464]), .Q(\Inst_Mem/inst_mem_reg[45][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][25]  ( .D(\Inst_Mem/inst_mem_reg[45][25] ), .CLK(clk), .RST(rst), .I(g_init[1465]), .Q(\Inst_Mem/inst_mem_reg[45][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][26]  ( .D(\Inst_Mem/inst_mem_reg[45][26] ), .CLK(clk), .RST(rst), .I(g_init[1466]), .Q(\Inst_Mem/inst_mem_reg[45][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][27]  ( .D(\Inst_Mem/inst_mem_reg[45][27] ), .CLK(clk), .RST(rst), .I(g_init[1467]), .Q(\Inst_Mem/inst_mem_reg[45][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][28]  ( .D(\Inst_Mem/inst_mem_reg[45][28] ), .CLK(clk), .RST(rst), .I(g_init[1468]), .Q(\Inst_Mem/inst_mem_reg[45][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][29]  ( .D(\Inst_Mem/inst_mem_reg[45][29] ), .CLK(clk), .RST(rst), .I(g_init[1469]), .Q(\Inst_Mem/inst_mem_reg[45][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][30]  ( .D(\Inst_Mem/inst_mem_reg[45][30] ), .CLK(clk), .RST(rst), .I(g_init[1470]), .Q(\Inst_Mem/inst_mem_reg[45][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[45][31]  ( .D(\Inst_Mem/inst_mem_reg[45][31] ), .CLK(clk), .RST(rst), .I(g_init[1471]), .Q(\Inst_Mem/inst_mem_reg[45][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][0]  ( .D(\Inst_Mem/inst_mem_reg[44][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1408]), .Q(
        \Inst_Mem/inst_mem_reg[44][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][1]  ( .D(\Inst_Mem/inst_mem_reg[44][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1409]), .Q(
        \Inst_Mem/inst_mem_reg[44][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][2]  ( .D(\Inst_Mem/inst_mem_reg[44][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1410]), .Q(
        \Inst_Mem/inst_mem_reg[44][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][3]  ( .D(\Inst_Mem/inst_mem_reg[44][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1411]), .Q(
        \Inst_Mem/inst_mem_reg[44][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][4]  ( .D(\Inst_Mem/inst_mem_reg[44][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1412]), .Q(
        \Inst_Mem/inst_mem_reg[44][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][5]  ( .D(\Inst_Mem/inst_mem_reg[44][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1413]), .Q(
        \Inst_Mem/inst_mem_reg[44][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][6]  ( .D(\Inst_Mem/inst_mem_reg[44][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1414]), .Q(
        \Inst_Mem/inst_mem_reg[44][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][7]  ( .D(\Inst_Mem/inst_mem_reg[44][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1415]), .Q(
        \Inst_Mem/inst_mem_reg[44][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][8]  ( .D(\Inst_Mem/inst_mem_reg[44][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1416]), .Q(
        \Inst_Mem/inst_mem_reg[44][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][9]  ( .D(\Inst_Mem/inst_mem_reg[44][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1417]), .Q(
        \Inst_Mem/inst_mem_reg[44][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[44][10]  ( .D(\Inst_Mem/inst_mem_reg[44][10] ), .CLK(clk), .RST(rst), .I(g_init[1418]), .Q(\Inst_Mem/inst_mem_reg[44][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][11]  ( .D(\Inst_Mem/inst_mem_reg[44][11] ), .CLK(clk), .RST(rst), .I(g_init[1419]), .Q(\Inst_Mem/inst_mem_reg[44][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][12]  ( .D(\Inst_Mem/inst_mem_reg[44][12] ), .CLK(clk), .RST(rst), .I(g_init[1420]), .Q(\Inst_Mem/inst_mem_reg[44][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][13]  ( .D(\Inst_Mem/inst_mem_reg[44][13] ), .CLK(clk), .RST(rst), .I(g_init[1421]), .Q(\Inst_Mem/inst_mem_reg[44][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][14]  ( .D(\Inst_Mem/inst_mem_reg[44][14] ), .CLK(clk), .RST(rst), .I(g_init[1422]), .Q(\Inst_Mem/inst_mem_reg[44][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][15]  ( .D(\Inst_Mem/inst_mem_reg[44][15] ), .CLK(clk), .RST(rst), .I(g_init[1423]), .Q(\Inst_Mem/inst_mem_reg[44][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][16]  ( .D(\Inst_Mem/inst_mem_reg[44][16] ), .CLK(clk), .RST(rst), .I(g_init[1424]), .Q(\Inst_Mem/inst_mem_reg[44][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][17]  ( .D(\Inst_Mem/inst_mem_reg[44][17] ), .CLK(clk), .RST(rst), .I(g_init[1425]), .Q(\Inst_Mem/inst_mem_reg[44][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][18]  ( .D(\Inst_Mem/inst_mem_reg[44][18] ), .CLK(clk), .RST(rst), .I(g_init[1426]), .Q(\Inst_Mem/inst_mem_reg[44][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][19]  ( .D(\Inst_Mem/inst_mem_reg[44][19] ), .CLK(clk), .RST(rst), .I(g_init[1427]), .Q(\Inst_Mem/inst_mem_reg[44][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][20]  ( .D(\Inst_Mem/inst_mem_reg[44][20] ), .CLK(clk), .RST(rst), .I(g_init[1428]), .Q(\Inst_Mem/inst_mem_reg[44][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][21]  ( .D(\Inst_Mem/inst_mem_reg[44][21] ), .CLK(clk), .RST(rst), .I(g_init[1429]), .Q(\Inst_Mem/inst_mem_reg[44][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][22]  ( .D(\Inst_Mem/inst_mem_reg[44][22] ), .CLK(clk), .RST(rst), .I(g_init[1430]), .Q(\Inst_Mem/inst_mem_reg[44][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][23]  ( .D(\Inst_Mem/inst_mem_reg[44][23] ), .CLK(clk), .RST(rst), .I(g_init[1431]), .Q(\Inst_Mem/inst_mem_reg[44][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][24]  ( .D(\Inst_Mem/inst_mem_reg[44][24] ), .CLK(clk), .RST(rst), .I(g_init[1432]), .Q(\Inst_Mem/inst_mem_reg[44][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][25]  ( .D(\Inst_Mem/inst_mem_reg[44][25] ), .CLK(clk), .RST(rst), .I(g_init[1433]), .Q(\Inst_Mem/inst_mem_reg[44][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][26]  ( .D(\Inst_Mem/inst_mem_reg[44][26] ), .CLK(clk), .RST(rst), .I(g_init[1434]), .Q(\Inst_Mem/inst_mem_reg[44][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][27]  ( .D(\Inst_Mem/inst_mem_reg[44][27] ), .CLK(clk), .RST(rst), .I(g_init[1435]), .Q(\Inst_Mem/inst_mem_reg[44][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][28]  ( .D(\Inst_Mem/inst_mem_reg[44][28] ), .CLK(clk), .RST(rst), .I(g_init[1436]), .Q(\Inst_Mem/inst_mem_reg[44][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][29]  ( .D(\Inst_Mem/inst_mem_reg[44][29] ), .CLK(clk), .RST(rst), .I(g_init[1437]), .Q(\Inst_Mem/inst_mem_reg[44][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][30]  ( .D(\Inst_Mem/inst_mem_reg[44][30] ), .CLK(clk), .RST(rst), .I(g_init[1438]), .Q(\Inst_Mem/inst_mem_reg[44][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[44][31]  ( .D(\Inst_Mem/inst_mem_reg[44][31] ), .CLK(clk), .RST(rst), .I(g_init[1439]), .Q(\Inst_Mem/inst_mem_reg[44][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][0]  ( .D(\Inst_Mem/inst_mem_reg[43][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1376]), .Q(
        \Inst_Mem/inst_mem_reg[43][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][1]  ( .D(\Inst_Mem/inst_mem_reg[43][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1377]), .Q(
        \Inst_Mem/inst_mem_reg[43][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][2]  ( .D(\Inst_Mem/inst_mem_reg[43][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1378]), .Q(
        \Inst_Mem/inst_mem_reg[43][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][3]  ( .D(\Inst_Mem/inst_mem_reg[43][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1379]), .Q(
        \Inst_Mem/inst_mem_reg[43][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][4]  ( .D(\Inst_Mem/inst_mem_reg[43][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1380]), .Q(
        \Inst_Mem/inst_mem_reg[43][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][5]  ( .D(\Inst_Mem/inst_mem_reg[43][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1381]), .Q(
        \Inst_Mem/inst_mem_reg[43][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][6]  ( .D(\Inst_Mem/inst_mem_reg[43][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1382]), .Q(
        \Inst_Mem/inst_mem_reg[43][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][7]  ( .D(\Inst_Mem/inst_mem_reg[43][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1383]), .Q(
        \Inst_Mem/inst_mem_reg[43][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][8]  ( .D(\Inst_Mem/inst_mem_reg[43][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1384]), .Q(
        \Inst_Mem/inst_mem_reg[43][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][9]  ( .D(\Inst_Mem/inst_mem_reg[43][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1385]), .Q(
        \Inst_Mem/inst_mem_reg[43][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[43][10]  ( .D(\Inst_Mem/inst_mem_reg[43][10] ), .CLK(clk), .RST(rst), .I(g_init[1386]), .Q(\Inst_Mem/inst_mem_reg[43][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][11]  ( .D(\Inst_Mem/inst_mem_reg[43][11] ), .CLK(clk), .RST(rst), .I(g_init[1387]), .Q(\Inst_Mem/inst_mem_reg[43][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][12]  ( .D(\Inst_Mem/inst_mem_reg[43][12] ), .CLK(clk), .RST(rst), .I(g_init[1388]), .Q(\Inst_Mem/inst_mem_reg[43][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][13]  ( .D(\Inst_Mem/inst_mem_reg[43][13] ), .CLK(clk), .RST(rst), .I(g_init[1389]), .Q(\Inst_Mem/inst_mem_reg[43][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][14]  ( .D(\Inst_Mem/inst_mem_reg[43][14] ), .CLK(clk), .RST(rst), .I(g_init[1390]), .Q(\Inst_Mem/inst_mem_reg[43][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][15]  ( .D(\Inst_Mem/inst_mem_reg[43][15] ), .CLK(clk), .RST(rst), .I(g_init[1391]), .Q(\Inst_Mem/inst_mem_reg[43][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][16]  ( .D(\Inst_Mem/inst_mem_reg[43][16] ), .CLK(clk), .RST(rst), .I(g_init[1392]), .Q(\Inst_Mem/inst_mem_reg[43][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][17]  ( .D(\Inst_Mem/inst_mem_reg[43][17] ), .CLK(clk), .RST(rst), .I(g_init[1393]), .Q(\Inst_Mem/inst_mem_reg[43][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][18]  ( .D(\Inst_Mem/inst_mem_reg[43][18] ), .CLK(clk), .RST(rst), .I(g_init[1394]), .Q(\Inst_Mem/inst_mem_reg[43][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][19]  ( .D(\Inst_Mem/inst_mem_reg[43][19] ), .CLK(clk), .RST(rst), .I(g_init[1395]), .Q(\Inst_Mem/inst_mem_reg[43][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][20]  ( .D(\Inst_Mem/inst_mem_reg[43][20] ), .CLK(clk), .RST(rst), .I(g_init[1396]), .Q(\Inst_Mem/inst_mem_reg[43][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][21]  ( .D(\Inst_Mem/inst_mem_reg[43][21] ), .CLK(clk), .RST(rst), .I(g_init[1397]), .Q(\Inst_Mem/inst_mem_reg[43][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][22]  ( .D(\Inst_Mem/inst_mem_reg[43][22] ), .CLK(clk), .RST(rst), .I(g_init[1398]), .Q(\Inst_Mem/inst_mem_reg[43][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][23]  ( .D(\Inst_Mem/inst_mem_reg[43][23] ), .CLK(clk), .RST(rst), .I(g_init[1399]), .Q(\Inst_Mem/inst_mem_reg[43][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][24]  ( .D(\Inst_Mem/inst_mem_reg[43][24] ), .CLK(clk), .RST(rst), .I(g_init[1400]), .Q(\Inst_Mem/inst_mem_reg[43][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][25]  ( .D(\Inst_Mem/inst_mem_reg[43][25] ), .CLK(clk), .RST(rst), .I(g_init[1401]), .Q(\Inst_Mem/inst_mem_reg[43][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][26]  ( .D(\Inst_Mem/inst_mem_reg[43][26] ), .CLK(clk), .RST(rst), .I(g_init[1402]), .Q(\Inst_Mem/inst_mem_reg[43][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][27]  ( .D(\Inst_Mem/inst_mem_reg[43][27] ), .CLK(clk), .RST(rst), .I(g_init[1403]), .Q(\Inst_Mem/inst_mem_reg[43][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][28]  ( .D(\Inst_Mem/inst_mem_reg[43][28] ), .CLK(clk), .RST(rst), .I(g_init[1404]), .Q(\Inst_Mem/inst_mem_reg[43][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][29]  ( .D(\Inst_Mem/inst_mem_reg[43][29] ), .CLK(clk), .RST(rst), .I(g_init[1405]), .Q(\Inst_Mem/inst_mem_reg[43][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][30]  ( .D(\Inst_Mem/inst_mem_reg[43][30] ), .CLK(clk), .RST(rst), .I(g_init[1406]), .Q(\Inst_Mem/inst_mem_reg[43][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[43][31]  ( .D(\Inst_Mem/inst_mem_reg[43][31] ), .CLK(clk), .RST(rst), .I(g_init[1407]), .Q(\Inst_Mem/inst_mem_reg[43][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][0]  ( .D(\Inst_Mem/inst_mem_reg[42][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1344]), .Q(
        \Inst_Mem/inst_mem_reg[42][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][1]  ( .D(\Inst_Mem/inst_mem_reg[42][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1345]), .Q(
        \Inst_Mem/inst_mem_reg[42][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][2]  ( .D(\Inst_Mem/inst_mem_reg[42][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1346]), .Q(
        \Inst_Mem/inst_mem_reg[42][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][3]  ( .D(\Inst_Mem/inst_mem_reg[42][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1347]), .Q(
        \Inst_Mem/inst_mem_reg[42][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][4]  ( .D(\Inst_Mem/inst_mem_reg[42][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1348]), .Q(
        \Inst_Mem/inst_mem_reg[42][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][5]  ( .D(\Inst_Mem/inst_mem_reg[42][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1349]), .Q(
        \Inst_Mem/inst_mem_reg[42][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][6]  ( .D(\Inst_Mem/inst_mem_reg[42][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1350]), .Q(
        \Inst_Mem/inst_mem_reg[42][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][7]  ( .D(\Inst_Mem/inst_mem_reg[42][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1351]), .Q(
        \Inst_Mem/inst_mem_reg[42][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][8]  ( .D(\Inst_Mem/inst_mem_reg[42][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1352]), .Q(
        \Inst_Mem/inst_mem_reg[42][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][9]  ( .D(\Inst_Mem/inst_mem_reg[42][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1353]), .Q(
        \Inst_Mem/inst_mem_reg[42][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[42][10]  ( .D(\Inst_Mem/inst_mem_reg[42][10] ), .CLK(clk), .RST(rst), .I(g_init[1354]), .Q(\Inst_Mem/inst_mem_reg[42][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][11]  ( .D(\Inst_Mem/inst_mem_reg[42][11] ), .CLK(clk), .RST(rst), .I(g_init[1355]), .Q(\Inst_Mem/inst_mem_reg[42][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][12]  ( .D(\Inst_Mem/inst_mem_reg[42][12] ), .CLK(clk), .RST(rst), .I(g_init[1356]), .Q(\Inst_Mem/inst_mem_reg[42][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][13]  ( .D(\Inst_Mem/inst_mem_reg[42][13] ), .CLK(clk), .RST(rst), .I(g_init[1357]), .Q(\Inst_Mem/inst_mem_reg[42][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][14]  ( .D(\Inst_Mem/inst_mem_reg[42][14] ), .CLK(clk), .RST(rst), .I(g_init[1358]), .Q(\Inst_Mem/inst_mem_reg[42][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][15]  ( .D(\Inst_Mem/inst_mem_reg[42][15] ), .CLK(clk), .RST(rst), .I(g_init[1359]), .Q(\Inst_Mem/inst_mem_reg[42][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][16]  ( .D(\Inst_Mem/inst_mem_reg[42][16] ), .CLK(clk), .RST(rst), .I(g_init[1360]), .Q(\Inst_Mem/inst_mem_reg[42][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][17]  ( .D(\Inst_Mem/inst_mem_reg[42][17] ), .CLK(clk), .RST(rst), .I(g_init[1361]), .Q(\Inst_Mem/inst_mem_reg[42][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][18]  ( .D(\Inst_Mem/inst_mem_reg[42][18] ), .CLK(clk), .RST(rst), .I(g_init[1362]), .Q(\Inst_Mem/inst_mem_reg[42][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][19]  ( .D(\Inst_Mem/inst_mem_reg[42][19] ), .CLK(clk), .RST(rst), .I(g_init[1363]), .Q(\Inst_Mem/inst_mem_reg[42][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][20]  ( .D(\Inst_Mem/inst_mem_reg[42][20] ), .CLK(clk), .RST(rst), .I(g_init[1364]), .Q(\Inst_Mem/inst_mem_reg[42][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][21]  ( .D(\Inst_Mem/inst_mem_reg[42][21] ), .CLK(clk), .RST(rst), .I(g_init[1365]), .Q(\Inst_Mem/inst_mem_reg[42][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][22]  ( .D(\Inst_Mem/inst_mem_reg[42][22] ), .CLK(clk), .RST(rst), .I(g_init[1366]), .Q(\Inst_Mem/inst_mem_reg[42][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][23]  ( .D(\Inst_Mem/inst_mem_reg[42][23] ), .CLK(clk), .RST(rst), .I(g_init[1367]), .Q(\Inst_Mem/inst_mem_reg[42][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][24]  ( .D(\Inst_Mem/inst_mem_reg[42][24] ), .CLK(clk), .RST(rst), .I(g_init[1368]), .Q(\Inst_Mem/inst_mem_reg[42][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][25]  ( .D(\Inst_Mem/inst_mem_reg[42][25] ), .CLK(clk), .RST(rst), .I(g_init[1369]), .Q(\Inst_Mem/inst_mem_reg[42][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][26]  ( .D(\Inst_Mem/inst_mem_reg[42][26] ), .CLK(clk), .RST(rst), .I(g_init[1370]), .Q(\Inst_Mem/inst_mem_reg[42][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][27]  ( .D(\Inst_Mem/inst_mem_reg[42][27] ), .CLK(clk), .RST(rst), .I(g_init[1371]), .Q(\Inst_Mem/inst_mem_reg[42][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][28]  ( .D(\Inst_Mem/inst_mem_reg[42][28] ), .CLK(clk), .RST(rst), .I(g_init[1372]), .Q(\Inst_Mem/inst_mem_reg[42][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][29]  ( .D(\Inst_Mem/inst_mem_reg[42][29] ), .CLK(clk), .RST(rst), .I(g_init[1373]), .Q(\Inst_Mem/inst_mem_reg[42][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][30]  ( .D(\Inst_Mem/inst_mem_reg[42][30] ), .CLK(clk), .RST(rst), .I(g_init[1374]), .Q(\Inst_Mem/inst_mem_reg[42][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[42][31]  ( .D(\Inst_Mem/inst_mem_reg[42][31] ), .CLK(clk), .RST(rst), .I(g_init[1375]), .Q(\Inst_Mem/inst_mem_reg[42][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][0]  ( .D(\Inst_Mem/inst_mem_reg[41][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1312]), .Q(
        \Inst_Mem/inst_mem_reg[41][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][1]  ( .D(\Inst_Mem/inst_mem_reg[41][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1313]), .Q(
        \Inst_Mem/inst_mem_reg[41][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][2]  ( .D(\Inst_Mem/inst_mem_reg[41][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1314]), .Q(
        \Inst_Mem/inst_mem_reg[41][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][3]  ( .D(\Inst_Mem/inst_mem_reg[41][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1315]), .Q(
        \Inst_Mem/inst_mem_reg[41][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][4]  ( .D(\Inst_Mem/inst_mem_reg[41][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1316]), .Q(
        \Inst_Mem/inst_mem_reg[41][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][5]  ( .D(\Inst_Mem/inst_mem_reg[41][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1317]), .Q(
        \Inst_Mem/inst_mem_reg[41][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][6]  ( .D(\Inst_Mem/inst_mem_reg[41][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1318]), .Q(
        \Inst_Mem/inst_mem_reg[41][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][7]  ( .D(\Inst_Mem/inst_mem_reg[41][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1319]), .Q(
        \Inst_Mem/inst_mem_reg[41][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][8]  ( .D(\Inst_Mem/inst_mem_reg[41][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1320]), .Q(
        \Inst_Mem/inst_mem_reg[41][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][9]  ( .D(\Inst_Mem/inst_mem_reg[41][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1321]), .Q(
        \Inst_Mem/inst_mem_reg[41][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[41][10]  ( .D(\Inst_Mem/inst_mem_reg[41][10] ), .CLK(clk), .RST(rst), .I(g_init[1322]), .Q(\Inst_Mem/inst_mem_reg[41][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][11]  ( .D(\Inst_Mem/inst_mem_reg[41][11] ), .CLK(clk), .RST(rst), .I(g_init[1323]), .Q(\Inst_Mem/inst_mem_reg[41][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][12]  ( .D(\Inst_Mem/inst_mem_reg[41][12] ), .CLK(clk), .RST(rst), .I(g_init[1324]), .Q(\Inst_Mem/inst_mem_reg[41][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][13]  ( .D(\Inst_Mem/inst_mem_reg[41][13] ), .CLK(clk), .RST(rst), .I(g_init[1325]), .Q(\Inst_Mem/inst_mem_reg[41][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][14]  ( .D(\Inst_Mem/inst_mem_reg[41][14] ), .CLK(clk), .RST(rst), .I(g_init[1326]), .Q(\Inst_Mem/inst_mem_reg[41][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][15]  ( .D(\Inst_Mem/inst_mem_reg[41][15] ), .CLK(clk), .RST(rst), .I(g_init[1327]), .Q(\Inst_Mem/inst_mem_reg[41][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][16]  ( .D(\Inst_Mem/inst_mem_reg[41][16] ), .CLK(clk), .RST(rst), .I(g_init[1328]), .Q(\Inst_Mem/inst_mem_reg[41][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][17]  ( .D(\Inst_Mem/inst_mem_reg[41][17] ), .CLK(clk), .RST(rst), .I(g_init[1329]), .Q(\Inst_Mem/inst_mem_reg[41][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][18]  ( .D(\Inst_Mem/inst_mem_reg[41][18] ), .CLK(clk), .RST(rst), .I(g_init[1330]), .Q(\Inst_Mem/inst_mem_reg[41][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][19]  ( .D(\Inst_Mem/inst_mem_reg[41][19] ), .CLK(clk), .RST(rst), .I(g_init[1331]), .Q(\Inst_Mem/inst_mem_reg[41][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][20]  ( .D(\Inst_Mem/inst_mem_reg[41][20] ), .CLK(clk), .RST(rst), .I(g_init[1332]), .Q(\Inst_Mem/inst_mem_reg[41][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][21]  ( .D(\Inst_Mem/inst_mem_reg[41][21] ), .CLK(clk), .RST(rst), .I(g_init[1333]), .Q(\Inst_Mem/inst_mem_reg[41][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][22]  ( .D(\Inst_Mem/inst_mem_reg[41][22] ), .CLK(clk), .RST(rst), .I(g_init[1334]), .Q(\Inst_Mem/inst_mem_reg[41][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][23]  ( .D(\Inst_Mem/inst_mem_reg[41][23] ), .CLK(clk), .RST(rst), .I(g_init[1335]), .Q(\Inst_Mem/inst_mem_reg[41][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][24]  ( .D(\Inst_Mem/inst_mem_reg[41][24] ), .CLK(clk), .RST(rst), .I(g_init[1336]), .Q(\Inst_Mem/inst_mem_reg[41][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][25]  ( .D(\Inst_Mem/inst_mem_reg[41][25] ), .CLK(clk), .RST(rst), .I(g_init[1337]), .Q(\Inst_Mem/inst_mem_reg[41][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][26]  ( .D(\Inst_Mem/inst_mem_reg[41][26] ), .CLK(clk), .RST(rst), .I(g_init[1338]), .Q(\Inst_Mem/inst_mem_reg[41][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][27]  ( .D(\Inst_Mem/inst_mem_reg[41][27] ), .CLK(clk), .RST(rst), .I(g_init[1339]), .Q(\Inst_Mem/inst_mem_reg[41][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][28]  ( .D(\Inst_Mem/inst_mem_reg[41][28] ), .CLK(clk), .RST(rst), .I(g_init[1340]), .Q(\Inst_Mem/inst_mem_reg[41][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][29]  ( .D(\Inst_Mem/inst_mem_reg[41][29] ), .CLK(clk), .RST(rst), .I(g_init[1341]), .Q(\Inst_Mem/inst_mem_reg[41][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][30]  ( .D(\Inst_Mem/inst_mem_reg[41][30] ), .CLK(clk), .RST(rst), .I(g_init[1342]), .Q(\Inst_Mem/inst_mem_reg[41][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[41][31]  ( .D(\Inst_Mem/inst_mem_reg[41][31] ), .CLK(clk), .RST(rst), .I(g_init[1343]), .Q(\Inst_Mem/inst_mem_reg[41][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][0]  ( .D(\Inst_Mem/inst_mem_reg[40][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1280]), .Q(
        \Inst_Mem/inst_mem_reg[40][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][1]  ( .D(\Inst_Mem/inst_mem_reg[40][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1281]), .Q(
        \Inst_Mem/inst_mem_reg[40][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][2]  ( .D(\Inst_Mem/inst_mem_reg[40][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1282]), .Q(
        \Inst_Mem/inst_mem_reg[40][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][3]  ( .D(\Inst_Mem/inst_mem_reg[40][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1283]), .Q(
        \Inst_Mem/inst_mem_reg[40][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][4]  ( .D(\Inst_Mem/inst_mem_reg[40][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1284]), .Q(
        \Inst_Mem/inst_mem_reg[40][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][5]  ( .D(\Inst_Mem/inst_mem_reg[40][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1285]), .Q(
        \Inst_Mem/inst_mem_reg[40][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][6]  ( .D(\Inst_Mem/inst_mem_reg[40][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1286]), .Q(
        \Inst_Mem/inst_mem_reg[40][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][7]  ( .D(\Inst_Mem/inst_mem_reg[40][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1287]), .Q(
        \Inst_Mem/inst_mem_reg[40][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][8]  ( .D(\Inst_Mem/inst_mem_reg[40][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1288]), .Q(
        \Inst_Mem/inst_mem_reg[40][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][9]  ( .D(\Inst_Mem/inst_mem_reg[40][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1289]), .Q(
        \Inst_Mem/inst_mem_reg[40][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[40][10]  ( .D(\Inst_Mem/inst_mem_reg[40][10] ), .CLK(clk), .RST(rst), .I(g_init[1290]), .Q(\Inst_Mem/inst_mem_reg[40][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][11]  ( .D(\Inst_Mem/inst_mem_reg[40][11] ), .CLK(clk), .RST(rst), .I(g_init[1291]), .Q(\Inst_Mem/inst_mem_reg[40][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][12]  ( .D(\Inst_Mem/inst_mem_reg[40][12] ), .CLK(clk), .RST(rst), .I(g_init[1292]), .Q(\Inst_Mem/inst_mem_reg[40][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][13]  ( .D(\Inst_Mem/inst_mem_reg[40][13] ), .CLK(clk), .RST(rst), .I(g_init[1293]), .Q(\Inst_Mem/inst_mem_reg[40][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][14]  ( .D(\Inst_Mem/inst_mem_reg[40][14] ), .CLK(clk), .RST(rst), .I(g_init[1294]), .Q(\Inst_Mem/inst_mem_reg[40][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][15]  ( .D(\Inst_Mem/inst_mem_reg[40][15] ), .CLK(clk), .RST(rst), .I(g_init[1295]), .Q(\Inst_Mem/inst_mem_reg[40][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][16]  ( .D(\Inst_Mem/inst_mem_reg[40][16] ), .CLK(clk), .RST(rst), .I(g_init[1296]), .Q(\Inst_Mem/inst_mem_reg[40][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][17]  ( .D(\Inst_Mem/inst_mem_reg[40][17] ), .CLK(clk), .RST(rst), .I(g_init[1297]), .Q(\Inst_Mem/inst_mem_reg[40][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][18]  ( .D(\Inst_Mem/inst_mem_reg[40][18] ), .CLK(clk), .RST(rst), .I(g_init[1298]), .Q(\Inst_Mem/inst_mem_reg[40][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][19]  ( .D(\Inst_Mem/inst_mem_reg[40][19] ), .CLK(clk), .RST(rst), .I(g_init[1299]), .Q(\Inst_Mem/inst_mem_reg[40][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][20]  ( .D(\Inst_Mem/inst_mem_reg[40][20] ), .CLK(clk), .RST(rst), .I(g_init[1300]), .Q(\Inst_Mem/inst_mem_reg[40][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][21]  ( .D(\Inst_Mem/inst_mem_reg[40][21] ), .CLK(clk), .RST(rst), .I(g_init[1301]), .Q(\Inst_Mem/inst_mem_reg[40][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][22]  ( .D(\Inst_Mem/inst_mem_reg[40][22] ), .CLK(clk), .RST(rst), .I(g_init[1302]), .Q(\Inst_Mem/inst_mem_reg[40][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][23]  ( .D(\Inst_Mem/inst_mem_reg[40][23] ), .CLK(clk), .RST(rst), .I(g_init[1303]), .Q(\Inst_Mem/inst_mem_reg[40][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][24]  ( .D(\Inst_Mem/inst_mem_reg[40][24] ), .CLK(clk), .RST(rst), .I(g_init[1304]), .Q(\Inst_Mem/inst_mem_reg[40][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][25]  ( .D(\Inst_Mem/inst_mem_reg[40][25] ), .CLK(clk), .RST(rst), .I(g_init[1305]), .Q(\Inst_Mem/inst_mem_reg[40][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][26]  ( .D(\Inst_Mem/inst_mem_reg[40][26] ), .CLK(clk), .RST(rst), .I(g_init[1306]), .Q(\Inst_Mem/inst_mem_reg[40][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][27]  ( .D(\Inst_Mem/inst_mem_reg[40][27] ), .CLK(clk), .RST(rst), .I(g_init[1307]), .Q(\Inst_Mem/inst_mem_reg[40][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][28]  ( .D(\Inst_Mem/inst_mem_reg[40][28] ), .CLK(clk), .RST(rst), .I(g_init[1308]), .Q(\Inst_Mem/inst_mem_reg[40][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][29]  ( .D(\Inst_Mem/inst_mem_reg[40][29] ), .CLK(clk), .RST(rst), .I(g_init[1309]), .Q(\Inst_Mem/inst_mem_reg[40][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][30]  ( .D(\Inst_Mem/inst_mem_reg[40][30] ), .CLK(clk), .RST(rst), .I(g_init[1310]), .Q(\Inst_Mem/inst_mem_reg[40][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[40][31]  ( .D(\Inst_Mem/inst_mem_reg[40][31] ), .CLK(clk), .RST(rst), .I(g_init[1311]), .Q(\Inst_Mem/inst_mem_reg[40][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][0]  ( .D(\Inst_Mem/inst_mem_reg[39][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1248]), .Q(
        \Inst_Mem/inst_mem_reg[39][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][1]  ( .D(\Inst_Mem/inst_mem_reg[39][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1249]), .Q(
        \Inst_Mem/inst_mem_reg[39][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][2]  ( .D(\Inst_Mem/inst_mem_reg[39][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1250]), .Q(
        \Inst_Mem/inst_mem_reg[39][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][3]  ( .D(\Inst_Mem/inst_mem_reg[39][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1251]), .Q(
        \Inst_Mem/inst_mem_reg[39][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][4]  ( .D(\Inst_Mem/inst_mem_reg[39][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1252]), .Q(
        \Inst_Mem/inst_mem_reg[39][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][5]  ( .D(\Inst_Mem/inst_mem_reg[39][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1253]), .Q(
        \Inst_Mem/inst_mem_reg[39][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][6]  ( .D(\Inst_Mem/inst_mem_reg[39][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1254]), .Q(
        \Inst_Mem/inst_mem_reg[39][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][7]  ( .D(\Inst_Mem/inst_mem_reg[39][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1255]), .Q(
        \Inst_Mem/inst_mem_reg[39][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][8]  ( .D(\Inst_Mem/inst_mem_reg[39][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1256]), .Q(
        \Inst_Mem/inst_mem_reg[39][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][9]  ( .D(\Inst_Mem/inst_mem_reg[39][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1257]), .Q(
        \Inst_Mem/inst_mem_reg[39][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[39][10]  ( .D(\Inst_Mem/inst_mem_reg[39][10] ), .CLK(clk), .RST(rst), .I(g_init[1258]), .Q(\Inst_Mem/inst_mem_reg[39][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][11]  ( .D(\Inst_Mem/inst_mem_reg[39][11] ), .CLK(clk), .RST(rst), .I(g_init[1259]), .Q(\Inst_Mem/inst_mem_reg[39][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][12]  ( .D(\Inst_Mem/inst_mem_reg[39][12] ), .CLK(clk), .RST(rst), .I(g_init[1260]), .Q(\Inst_Mem/inst_mem_reg[39][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][13]  ( .D(\Inst_Mem/inst_mem_reg[39][13] ), .CLK(clk), .RST(rst), .I(g_init[1261]), .Q(\Inst_Mem/inst_mem_reg[39][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][14]  ( .D(\Inst_Mem/inst_mem_reg[39][14] ), .CLK(clk), .RST(rst), .I(g_init[1262]), .Q(\Inst_Mem/inst_mem_reg[39][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][15]  ( .D(\Inst_Mem/inst_mem_reg[39][15] ), .CLK(clk), .RST(rst), .I(g_init[1263]), .Q(\Inst_Mem/inst_mem_reg[39][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][16]  ( .D(\Inst_Mem/inst_mem_reg[39][16] ), .CLK(clk), .RST(rst), .I(g_init[1264]), .Q(\Inst_Mem/inst_mem_reg[39][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][17]  ( .D(\Inst_Mem/inst_mem_reg[39][17] ), .CLK(clk), .RST(rst), .I(g_init[1265]), .Q(\Inst_Mem/inst_mem_reg[39][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][18]  ( .D(\Inst_Mem/inst_mem_reg[39][18] ), .CLK(clk), .RST(rst), .I(g_init[1266]), .Q(\Inst_Mem/inst_mem_reg[39][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][19]  ( .D(\Inst_Mem/inst_mem_reg[39][19] ), .CLK(clk), .RST(rst), .I(g_init[1267]), .Q(\Inst_Mem/inst_mem_reg[39][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][20]  ( .D(\Inst_Mem/inst_mem_reg[39][20] ), .CLK(clk), .RST(rst), .I(g_init[1268]), .Q(\Inst_Mem/inst_mem_reg[39][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][21]  ( .D(\Inst_Mem/inst_mem_reg[39][21] ), .CLK(clk), .RST(rst), .I(g_init[1269]), .Q(\Inst_Mem/inst_mem_reg[39][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][22]  ( .D(\Inst_Mem/inst_mem_reg[39][22] ), .CLK(clk), .RST(rst), .I(g_init[1270]), .Q(\Inst_Mem/inst_mem_reg[39][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][23]  ( .D(\Inst_Mem/inst_mem_reg[39][23] ), .CLK(clk), .RST(rst), .I(g_init[1271]), .Q(\Inst_Mem/inst_mem_reg[39][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][24]  ( .D(\Inst_Mem/inst_mem_reg[39][24] ), .CLK(clk), .RST(rst), .I(g_init[1272]), .Q(\Inst_Mem/inst_mem_reg[39][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][25]  ( .D(\Inst_Mem/inst_mem_reg[39][25] ), .CLK(clk), .RST(rst), .I(g_init[1273]), .Q(\Inst_Mem/inst_mem_reg[39][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][26]  ( .D(\Inst_Mem/inst_mem_reg[39][26] ), .CLK(clk), .RST(rst), .I(g_init[1274]), .Q(\Inst_Mem/inst_mem_reg[39][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][27]  ( .D(\Inst_Mem/inst_mem_reg[39][27] ), .CLK(clk), .RST(rst), .I(g_init[1275]), .Q(\Inst_Mem/inst_mem_reg[39][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][28]  ( .D(\Inst_Mem/inst_mem_reg[39][28] ), .CLK(clk), .RST(rst), .I(g_init[1276]), .Q(\Inst_Mem/inst_mem_reg[39][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][29]  ( .D(\Inst_Mem/inst_mem_reg[39][29] ), .CLK(clk), .RST(rst), .I(g_init[1277]), .Q(\Inst_Mem/inst_mem_reg[39][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][30]  ( .D(\Inst_Mem/inst_mem_reg[39][30] ), .CLK(clk), .RST(rst), .I(g_init[1278]), .Q(\Inst_Mem/inst_mem_reg[39][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[39][31]  ( .D(\Inst_Mem/inst_mem_reg[39][31] ), .CLK(clk), .RST(rst), .I(g_init[1279]), .Q(\Inst_Mem/inst_mem_reg[39][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][0]  ( .D(\Inst_Mem/inst_mem_reg[38][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1216]), .Q(
        \Inst_Mem/inst_mem_reg[38][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][1]  ( .D(\Inst_Mem/inst_mem_reg[38][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1217]), .Q(
        \Inst_Mem/inst_mem_reg[38][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][2]  ( .D(\Inst_Mem/inst_mem_reg[38][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1218]), .Q(
        \Inst_Mem/inst_mem_reg[38][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][3]  ( .D(\Inst_Mem/inst_mem_reg[38][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1219]), .Q(
        \Inst_Mem/inst_mem_reg[38][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][4]  ( .D(\Inst_Mem/inst_mem_reg[38][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1220]), .Q(
        \Inst_Mem/inst_mem_reg[38][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][5]  ( .D(\Inst_Mem/inst_mem_reg[38][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1221]), .Q(
        \Inst_Mem/inst_mem_reg[38][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][6]  ( .D(\Inst_Mem/inst_mem_reg[38][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1222]), .Q(
        \Inst_Mem/inst_mem_reg[38][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][7]  ( .D(\Inst_Mem/inst_mem_reg[38][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1223]), .Q(
        \Inst_Mem/inst_mem_reg[38][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][8]  ( .D(\Inst_Mem/inst_mem_reg[38][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1224]), .Q(
        \Inst_Mem/inst_mem_reg[38][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][9]  ( .D(\Inst_Mem/inst_mem_reg[38][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1225]), .Q(
        \Inst_Mem/inst_mem_reg[38][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[38][10]  ( .D(\Inst_Mem/inst_mem_reg[38][10] ), .CLK(clk), .RST(rst), .I(g_init[1226]), .Q(\Inst_Mem/inst_mem_reg[38][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][11]  ( .D(\Inst_Mem/inst_mem_reg[38][11] ), .CLK(clk), .RST(rst), .I(g_init[1227]), .Q(\Inst_Mem/inst_mem_reg[38][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][12]  ( .D(\Inst_Mem/inst_mem_reg[38][12] ), .CLK(clk), .RST(rst), .I(g_init[1228]), .Q(\Inst_Mem/inst_mem_reg[38][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][13]  ( .D(\Inst_Mem/inst_mem_reg[38][13] ), .CLK(clk), .RST(rst), .I(g_init[1229]), .Q(\Inst_Mem/inst_mem_reg[38][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][14]  ( .D(\Inst_Mem/inst_mem_reg[38][14] ), .CLK(clk), .RST(rst), .I(g_init[1230]), .Q(\Inst_Mem/inst_mem_reg[38][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][15]  ( .D(\Inst_Mem/inst_mem_reg[38][15] ), .CLK(clk), .RST(rst), .I(g_init[1231]), .Q(\Inst_Mem/inst_mem_reg[38][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][16]  ( .D(\Inst_Mem/inst_mem_reg[38][16] ), .CLK(clk), .RST(rst), .I(g_init[1232]), .Q(\Inst_Mem/inst_mem_reg[38][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][17]  ( .D(\Inst_Mem/inst_mem_reg[38][17] ), .CLK(clk), .RST(rst), .I(g_init[1233]), .Q(\Inst_Mem/inst_mem_reg[38][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][18]  ( .D(\Inst_Mem/inst_mem_reg[38][18] ), .CLK(clk), .RST(rst), .I(g_init[1234]), .Q(\Inst_Mem/inst_mem_reg[38][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][19]  ( .D(\Inst_Mem/inst_mem_reg[38][19] ), .CLK(clk), .RST(rst), .I(g_init[1235]), .Q(\Inst_Mem/inst_mem_reg[38][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][20]  ( .D(\Inst_Mem/inst_mem_reg[38][20] ), .CLK(clk), .RST(rst), .I(g_init[1236]), .Q(\Inst_Mem/inst_mem_reg[38][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][21]  ( .D(\Inst_Mem/inst_mem_reg[38][21] ), .CLK(clk), .RST(rst), .I(g_init[1237]), .Q(\Inst_Mem/inst_mem_reg[38][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][22]  ( .D(\Inst_Mem/inst_mem_reg[38][22] ), .CLK(clk), .RST(rst), .I(g_init[1238]), .Q(\Inst_Mem/inst_mem_reg[38][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][23]  ( .D(\Inst_Mem/inst_mem_reg[38][23] ), .CLK(clk), .RST(rst), .I(g_init[1239]), .Q(\Inst_Mem/inst_mem_reg[38][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][24]  ( .D(\Inst_Mem/inst_mem_reg[38][24] ), .CLK(clk), .RST(rst), .I(g_init[1240]), .Q(\Inst_Mem/inst_mem_reg[38][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][25]  ( .D(\Inst_Mem/inst_mem_reg[38][25] ), .CLK(clk), .RST(rst), .I(g_init[1241]), .Q(\Inst_Mem/inst_mem_reg[38][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][26]  ( .D(\Inst_Mem/inst_mem_reg[38][26] ), .CLK(clk), .RST(rst), .I(g_init[1242]), .Q(\Inst_Mem/inst_mem_reg[38][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][27]  ( .D(\Inst_Mem/inst_mem_reg[38][27] ), .CLK(clk), .RST(rst), .I(g_init[1243]), .Q(\Inst_Mem/inst_mem_reg[38][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][28]  ( .D(\Inst_Mem/inst_mem_reg[38][28] ), .CLK(clk), .RST(rst), .I(g_init[1244]), .Q(\Inst_Mem/inst_mem_reg[38][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][29]  ( .D(\Inst_Mem/inst_mem_reg[38][29] ), .CLK(clk), .RST(rst), .I(g_init[1245]), .Q(\Inst_Mem/inst_mem_reg[38][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][30]  ( .D(\Inst_Mem/inst_mem_reg[38][30] ), .CLK(clk), .RST(rst), .I(g_init[1246]), .Q(\Inst_Mem/inst_mem_reg[38][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[38][31]  ( .D(\Inst_Mem/inst_mem_reg[38][31] ), .CLK(clk), .RST(rst), .I(g_init[1247]), .Q(\Inst_Mem/inst_mem_reg[38][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][0]  ( .D(\Inst_Mem/inst_mem_reg[37][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1184]), .Q(
        \Inst_Mem/inst_mem_reg[37][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][1]  ( .D(\Inst_Mem/inst_mem_reg[37][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1185]), .Q(
        \Inst_Mem/inst_mem_reg[37][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][2]  ( .D(\Inst_Mem/inst_mem_reg[37][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1186]), .Q(
        \Inst_Mem/inst_mem_reg[37][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][3]  ( .D(\Inst_Mem/inst_mem_reg[37][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1187]), .Q(
        \Inst_Mem/inst_mem_reg[37][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][4]  ( .D(\Inst_Mem/inst_mem_reg[37][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1188]), .Q(
        \Inst_Mem/inst_mem_reg[37][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][5]  ( .D(\Inst_Mem/inst_mem_reg[37][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1189]), .Q(
        \Inst_Mem/inst_mem_reg[37][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][6]  ( .D(\Inst_Mem/inst_mem_reg[37][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1190]), .Q(
        \Inst_Mem/inst_mem_reg[37][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][7]  ( .D(\Inst_Mem/inst_mem_reg[37][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1191]), .Q(
        \Inst_Mem/inst_mem_reg[37][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][8]  ( .D(\Inst_Mem/inst_mem_reg[37][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1192]), .Q(
        \Inst_Mem/inst_mem_reg[37][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][9]  ( .D(\Inst_Mem/inst_mem_reg[37][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1193]), .Q(
        \Inst_Mem/inst_mem_reg[37][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[37][10]  ( .D(\Inst_Mem/inst_mem_reg[37][10] ), .CLK(clk), .RST(rst), .I(g_init[1194]), .Q(\Inst_Mem/inst_mem_reg[37][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][11]  ( .D(\Inst_Mem/inst_mem_reg[37][11] ), .CLK(clk), .RST(rst), .I(g_init[1195]), .Q(\Inst_Mem/inst_mem_reg[37][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][12]  ( .D(\Inst_Mem/inst_mem_reg[37][12] ), .CLK(clk), .RST(rst), .I(g_init[1196]), .Q(\Inst_Mem/inst_mem_reg[37][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][13]  ( .D(\Inst_Mem/inst_mem_reg[37][13] ), .CLK(clk), .RST(rst), .I(g_init[1197]), .Q(\Inst_Mem/inst_mem_reg[37][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][14]  ( .D(\Inst_Mem/inst_mem_reg[37][14] ), .CLK(clk), .RST(rst), .I(g_init[1198]), .Q(\Inst_Mem/inst_mem_reg[37][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][15]  ( .D(\Inst_Mem/inst_mem_reg[37][15] ), .CLK(clk), .RST(rst), .I(g_init[1199]), .Q(\Inst_Mem/inst_mem_reg[37][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][16]  ( .D(\Inst_Mem/inst_mem_reg[37][16] ), .CLK(clk), .RST(rst), .I(g_init[1200]), .Q(\Inst_Mem/inst_mem_reg[37][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][17]  ( .D(\Inst_Mem/inst_mem_reg[37][17] ), .CLK(clk), .RST(rst), .I(g_init[1201]), .Q(\Inst_Mem/inst_mem_reg[37][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][18]  ( .D(\Inst_Mem/inst_mem_reg[37][18] ), .CLK(clk), .RST(rst), .I(g_init[1202]), .Q(\Inst_Mem/inst_mem_reg[37][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][19]  ( .D(\Inst_Mem/inst_mem_reg[37][19] ), .CLK(clk), .RST(rst), .I(g_init[1203]), .Q(\Inst_Mem/inst_mem_reg[37][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][20]  ( .D(\Inst_Mem/inst_mem_reg[37][20] ), .CLK(clk), .RST(rst), .I(g_init[1204]), .Q(\Inst_Mem/inst_mem_reg[37][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][21]  ( .D(\Inst_Mem/inst_mem_reg[37][21] ), .CLK(clk), .RST(rst), .I(g_init[1205]), .Q(\Inst_Mem/inst_mem_reg[37][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][22]  ( .D(\Inst_Mem/inst_mem_reg[37][22] ), .CLK(clk), .RST(rst), .I(g_init[1206]), .Q(\Inst_Mem/inst_mem_reg[37][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][23]  ( .D(\Inst_Mem/inst_mem_reg[37][23] ), .CLK(clk), .RST(rst), .I(g_init[1207]), .Q(\Inst_Mem/inst_mem_reg[37][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][24]  ( .D(\Inst_Mem/inst_mem_reg[37][24] ), .CLK(clk), .RST(rst), .I(g_init[1208]), .Q(\Inst_Mem/inst_mem_reg[37][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][25]  ( .D(\Inst_Mem/inst_mem_reg[37][25] ), .CLK(clk), .RST(rst), .I(g_init[1209]), .Q(\Inst_Mem/inst_mem_reg[37][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][26]  ( .D(\Inst_Mem/inst_mem_reg[37][26] ), .CLK(clk), .RST(rst), .I(g_init[1210]), .Q(\Inst_Mem/inst_mem_reg[37][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][27]  ( .D(\Inst_Mem/inst_mem_reg[37][27] ), .CLK(clk), .RST(rst), .I(g_init[1211]), .Q(\Inst_Mem/inst_mem_reg[37][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][28]  ( .D(\Inst_Mem/inst_mem_reg[37][28] ), .CLK(clk), .RST(rst), .I(g_init[1212]), .Q(\Inst_Mem/inst_mem_reg[37][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][29]  ( .D(\Inst_Mem/inst_mem_reg[37][29] ), .CLK(clk), .RST(rst), .I(g_init[1213]), .Q(\Inst_Mem/inst_mem_reg[37][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][30]  ( .D(\Inst_Mem/inst_mem_reg[37][30] ), .CLK(clk), .RST(rst), .I(g_init[1214]), .Q(\Inst_Mem/inst_mem_reg[37][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[37][31]  ( .D(\Inst_Mem/inst_mem_reg[37][31] ), .CLK(clk), .RST(rst), .I(g_init[1215]), .Q(\Inst_Mem/inst_mem_reg[37][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][0]  ( .D(\Inst_Mem/inst_mem_reg[36][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1152]), .Q(
        \Inst_Mem/inst_mem_reg[36][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][1]  ( .D(\Inst_Mem/inst_mem_reg[36][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1153]), .Q(
        \Inst_Mem/inst_mem_reg[36][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][2]  ( .D(\Inst_Mem/inst_mem_reg[36][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1154]), .Q(
        \Inst_Mem/inst_mem_reg[36][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][3]  ( .D(\Inst_Mem/inst_mem_reg[36][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1155]), .Q(
        \Inst_Mem/inst_mem_reg[36][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][4]  ( .D(\Inst_Mem/inst_mem_reg[36][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1156]), .Q(
        \Inst_Mem/inst_mem_reg[36][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][5]  ( .D(\Inst_Mem/inst_mem_reg[36][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1157]), .Q(
        \Inst_Mem/inst_mem_reg[36][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][6]  ( .D(\Inst_Mem/inst_mem_reg[36][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1158]), .Q(
        \Inst_Mem/inst_mem_reg[36][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][7]  ( .D(\Inst_Mem/inst_mem_reg[36][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1159]), .Q(
        \Inst_Mem/inst_mem_reg[36][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][8]  ( .D(\Inst_Mem/inst_mem_reg[36][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1160]), .Q(
        \Inst_Mem/inst_mem_reg[36][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][9]  ( .D(\Inst_Mem/inst_mem_reg[36][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1161]), .Q(
        \Inst_Mem/inst_mem_reg[36][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[36][10]  ( .D(\Inst_Mem/inst_mem_reg[36][10] ), .CLK(clk), .RST(rst), .I(g_init[1162]), .Q(\Inst_Mem/inst_mem_reg[36][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][11]  ( .D(\Inst_Mem/inst_mem_reg[36][11] ), .CLK(clk), .RST(rst), .I(g_init[1163]), .Q(\Inst_Mem/inst_mem_reg[36][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][12]  ( .D(\Inst_Mem/inst_mem_reg[36][12] ), .CLK(clk), .RST(rst), .I(g_init[1164]), .Q(\Inst_Mem/inst_mem_reg[36][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][13]  ( .D(\Inst_Mem/inst_mem_reg[36][13] ), .CLK(clk), .RST(rst), .I(g_init[1165]), .Q(\Inst_Mem/inst_mem_reg[36][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][14]  ( .D(\Inst_Mem/inst_mem_reg[36][14] ), .CLK(clk), .RST(rst), .I(g_init[1166]), .Q(\Inst_Mem/inst_mem_reg[36][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][15]  ( .D(\Inst_Mem/inst_mem_reg[36][15] ), .CLK(clk), .RST(rst), .I(g_init[1167]), .Q(\Inst_Mem/inst_mem_reg[36][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][16]  ( .D(\Inst_Mem/inst_mem_reg[36][16] ), .CLK(clk), .RST(rst), .I(g_init[1168]), .Q(\Inst_Mem/inst_mem_reg[36][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][17]  ( .D(\Inst_Mem/inst_mem_reg[36][17] ), .CLK(clk), .RST(rst), .I(g_init[1169]), .Q(\Inst_Mem/inst_mem_reg[36][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][18]  ( .D(\Inst_Mem/inst_mem_reg[36][18] ), .CLK(clk), .RST(rst), .I(g_init[1170]), .Q(\Inst_Mem/inst_mem_reg[36][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][19]  ( .D(\Inst_Mem/inst_mem_reg[36][19] ), .CLK(clk), .RST(rst), .I(g_init[1171]), .Q(\Inst_Mem/inst_mem_reg[36][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][20]  ( .D(\Inst_Mem/inst_mem_reg[36][20] ), .CLK(clk), .RST(rst), .I(g_init[1172]), .Q(\Inst_Mem/inst_mem_reg[36][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][21]  ( .D(\Inst_Mem/inst_mem_reg[36][21] ), .CLK(clk), .RST(rst), .I(g_init[1173]), .Q(\Inst_Mem/inst_mem_reg[36][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][22]  ( .D(\Inst_Mem/inst_mem_reg[36][22] ), .CLK(clk), .RST(rst), .I(g_init[1174]), .Q(\Inst_Mem/inst_mem_reg[36][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][23]  ( .D(\Inst_Mem/inst_mem_reg[36][23] ), .CLK(clk), .RST(rst), .I(g_init[1175]), .Q(\Inst_Mem/inst_mem_reg[36][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][24]  ( .D(\Inst_Mem/inst_mem_reg[36][24] ), .CLK(clk), .RST(rst), .I(g_init[1176]), .Q(\Inst_Mem/inst_mem_reg[36][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][25]  ( .D(\Inst_Mem/inst_mem_reg[36][25] ), .CLK(clk), .RST(rst), .I(g_init[1177]), .Q(\Inst_Mem/inst_mem_reg[36][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][26]  ( .D(\Inst_Mem/inst_mem_reg[36][26] ), .CLK(clk), .RST(rst), .I(g_init[1178]), .Q(\Inst_Mem/inst_mem_reg[36][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][27]  ( .D(\Inst_Mem/inst_mem_reg[36][27] ), .CLK(clk), .RST(rst), .I(g_init[1179]), .Q(\Inst_Mem/inst_mem_reg[36][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][28]  ( .D(\Inst_Mem/inst_mem_reg[36][28] ), .CLK(clk), .RST(rst), .I(g_init[1180]), .Q(\Inst_Mem/inst_mem_reg[36][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][29]  ( .D(\Inst_Mem/inst_mem_reg[36][29] ), .CLK(clk), .RST(rst), .I(g_init[1181]), .Q(\Inst_Mem/inst_mem_reg[36][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][30]  ( .D(\Inst_Mem/inst_mem_reg[36][30] ), .CLK(clk), .RST(rst), .I(g_init[1182]), .Q(\Inst_Mem/inst_mem_reg[36][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[36][31]  ( .D(\Inst_Mem/inst_mem_reg[36][31] ), .CLK(clk), .RST(rst), .I(g_init[1183]), .Q(\Inst_Mem/inst_mem_reg[36][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][0]  ( .D(\Inst_Mem/inst_mem_reg[35][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1120]), .Q(
        \Inst_Mem/inst_mem_reg[35][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][1]  ( .D(\Inst_Mem/inst_mem_reg[35][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1121]), .Q(
        \Inst_Mem/inst_mem_reg[35][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][2]  ( .D(\Inst_Mem/inst_mem_reg[35][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1122]), .Q(
        \Inst_Mem/inst_mem_reg[35][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][3]  ( .D(\Inst_Mem/inst_mem_reg[35][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1123]), .Q(
        \Inst_Mem/inst_mem_reg[35][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][4]  ( .D(\Inst_Mem/inst_mem_reg[35][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1124]), .Q(
        \Inst_Mem/inst_mem_reg[35][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][5]  ( .D(\Inst_Mem/inst_mem_reg[35][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1125]), .Q(
        \Inst_Mem/inst_mem_reg[35][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][6]  ( .D(\Inst_Mem/inst_mem_reg[35][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1126]), .Q(
        \Inst_Mem/inst_mem_reg[35][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][7]  ( .D(\Inst_Mem/inst_mem_reg[35][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1127]), .Q(
        \Inst_Mem/inst_mem_reg[35][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][8]  ( .D(\Inst_Mem/inst_mem_reg[35][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1128]), .Q(
        \Inst_Mem/inst_mem_reg[35][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][9]  ( .D(\Inst_Mem/inst_mem_reg[35][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1129]), .Q(
        \Inst_Mem/inst_mem_reg[35][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[35][10]  ( .D(\Inst_Mem/inst_mem_reg[35][10] ), .CLK(clk), .RST(rst), .I(g_init[1130]), .Q(\Inst_Mem/inst_mem_reg[35][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][11]  ( .D(\Inst_Mem/inst_mem_reg[35][11] ), .CLK(clk), .RST(rst), .I(g_init[1131]), .Q(\Inst_Mem/inst_mem_reg[35][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][12]  ( .D(\Inst_Mem/inst_mem_reg[35][12] ), .CLK(clk), .RST(rst), .I(g_init[1132]), .Q(\Inst_Mem/inst_mem_reg[35][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][13]  ( .D(\Inst_Mem/inst_mem_reg[35][13] ), .CLK(clk), .RST(rst), .I(g_init[1133]), .Q(\Inst_Mem/inst_mem_reg[35][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][14]  ( .D(\Inst_Mem/inst_mem_reg[35][14] ), .CLK(clk), .RST(rst), .I(g_init[1134]), .Q(\Inst_Mem/inst_mem_reg[35][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][15]  ( .D(\Inst_Mem/inst_mem_reg[35][15] ), .CLK(clk), .RST(rst), .I(g_init[1135]), .Q(\Inst_Mem/inst_mem_reg[35][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][16]  ( .D(\Inst_Mem/inst_mem_reg[35][16] ), .CLK(clk), .RST(rst), .I(g_init[1136]), .Q(\Inst_Mem/inst_mem_reg[35][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][17]  ( .D(\Inst_Mem/inst_mem_reg[35][17] ), .CLK(clk), .RST(rst), .I(g_init[1137]), .Q(\Inst_Mem/inst_mem_reg[35][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][18]  ( .D(\Inst_Mem/inst_mem_reg[35][18] ), .CLK(clk), .RST(rst), .I(g_init[1138]), .Q(\Inst_Mem/inst_mem_reg[35][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][19]  ( .D(\Inst_Mem/inst_mem_reg[35][19] ), .CLK(clk), .RST(rst), .I(g_init[1139]), .Q(\Inst_Mem/inst_mem_reg[35][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][20]  ( .D(\Inst_Mem/inst_mem_reg[35][20] ), .CLK(clk), .RST(rst), .I(g_init[1140]), .Q(\Inst_Mem/inst_mem_reg[35][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][21]  ( .D(\Inst_Mem/inst_mem_reg[35][21] ), .CLK(clk), .RST(rst), .I(g_init[1141]), .Q(\Inst_Mem/inst_mem_reg[35][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][22]  ( .D(\Inst_Mem/inst_mem_reg[35][22] ), .CLK(clk), .RST(rst), .I(g_init[1142]), .Q(\Inst_Mem/inst_mem_reg[35][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][23]  ( .D(\Inst_Mem/inst_mem_reg[35][23] ), .CLK(clk), .RST(rst), .I(g_init[1143]), .Q(\Inst_Mem/inst_mem_reg[35][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][24]  ( .D(\Inst_Mem/inst_mem_reg[35][24] ), .CLK(clk), .RST(rst), .I(g_init[1144]), .Q(\Inst_Mem/inst_mem_reg[35][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][25]  ( .D(\Inst_Mem/inst_mem_reg[35][25] ), .CLK(clk), .RST(rst), .I(g_init[1145]), .Q(\Inst_Mem/inst_mem_reg[35][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][26]  ( .D(\Inst_Mem/inst_mem_reg[35][26] ), .CLK(clk), .RST(rst), .I(g_init[1146]), .Q(\Inst_Mem/inst_mem_reg[35][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][27]  ( .D(\Inst_Mem/inst_mem_reg[35][27] ), .CLK(clk), .RST(rst), .I(g_init[1147]), .Q(\Inst_Mem/inst_mem_reg[35][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][28]  ( .D(\Inst_Mem/inst_mem_reg[35][28] ), .CLK(clk), .RST(rst), .I(g_init[1148]), .Q(\Inst_Mem/inst_mem_reg[35][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][29]  ( .D(\Inst_Mem/inst_mem_reg[35][29] ), .CLK(clk), .RST(rst), .I(g_init[1149]), .Q(\Inst_Mem/inst_mem_reg[35][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][30]  ( .D(\Inst_Mem/inst_mem_reg[35][30] ), .CLK(clk), .RST(rst), .I(g_init[1150]), .Q(\Inst_Mem/inst_mem_reg[35][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[35][31]  ( .D(\Inst_Mem/inst_mem_reg[35][31] ), .CLK(clk), .RST(rst), .I(g_init[1151]), .Q(\Inst_Mem/inst_mem_reg[35][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][0]  ( .D(\Inst_Mem/inst_mem_reg[34][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1088]), .Q(
        \Inst_Mem/inst_mem_reg[34][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][1]  ( .D(\Inst_Mem/inst_mem_reg[34][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1089]), .Q(
        \Inst_Mem/inst_mem_reg[34][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][2]  ( .D(\Inst_Mem/inst_mem_reg[34][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1090]), .Q(
        \Inst_Mem/inst_mem_reg[34][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][3]  ( .D(\Inst_Mem/inst_mem_reg[34][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1091]), .Q(
        \Inst_Mem/inst_mem_reg[34][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][4]  ( .D(\Inst_Mem/inst_mem_reg[34][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1092]), .Q(
        \Inst_Mem/inst_mem_reg[34][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][5]  ( .D(\Inst_Mem/inst_mem_reg[34][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1093]), .Q(
        \Inst_Mem/inst_mem_reg[34][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][6]  ( .D(\Inst_Mem/inst_mem_reg[34][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1094]), .Q(
        \Inst_Mem/inst_mem_reg[34][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][7]  ( .D(\Inst_Mem/inst_mem_reg[34][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1095]), .Q(
        \Inst_Mem/inst_mem_reg[34][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][8]  ( .D(\Inst_Mem/inst_mem_reg[34][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1096]), .Q(
        \Inst_Mem/inst_mem_reg[34][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][9]  ( .D(\Inst_Mem/inst_mem_reg[34][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1097]), .Q(
        \Inst_Mem/inst_mem_reg[34][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[34][10]  ( .D(\Inst_Mem/inst_mem_reg[34][10] ), .CLK(clk), .RST(rst), .I(g_init[1098]), .Q(\Inst_Mem/inst_mem_reg[34][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][11]  ( .D(\Inst_Mem/inst_mem_reg[34][11] ), .CLK(clk), .RST(rst), .I(g_init[1099]), .Q(\Inst_Mem/inst_mem_reg[34][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][12]  ( .D(\Inst_Mem/inst_mem_reg[34][12] ), .CLK(clk), .RST(rst), .I(g_init[1100]), .Q(\Inst_Mem/inst_mem_reg[34][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][13]  ( .D(\Inst_Mem/inst_mem_reg[34][13] ), .CLK(clk), .RST(rst), .I(g_init[1101]), .Q(\Inst_Mem/inst_mem_reg[34][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][14]  ( .D(\Inst_Mem/inst_mem_reg[34][14] ), .CLK(clk), .RST(rst), .I(g_init[1102]), .Q(\Inst_Mem/inst_mem_reg[34][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][15]  ( .D(\Inst_Mem/inst_mem_reg[34][15] ), .CLK(clk), .RST(rst), .I(g_init[1103]), .Q(\Inst_Mem/inst_mem_reg[34][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][16]  ( .D(\Inst_Mem/inst_mem_reg[34][16] ), .CLK(clk), .RST(rst), .I(g_init[1104]), .Q(\Inst_Mem/inst_mem_reg[34][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][17]  ( .D(\Inst_Mem/inst_mem_reg[34][17] ), .CLK(clk), .RST(rst), .I(g_init[1105]), .Q(\Inst_Mem/inst_mem_reg[34][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][18]  ( .D(\Inst_Mem/inst_mem_reg[34][18] ), .CLK(clk), .RST(rst), .I(g_init[1106]), .Q(\Inst_Mem/inst_mem_reg[34][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][19]  ( .D(\Inst_Mem/inst_mem_reg[34][19] ), .CLK(clk), .RST(rst), .I(g_init[1107]), .Q(\Inst_Mem/inst_mem_reg[34][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][20]  ( .D(\Inst_Mem/inst_mem_reg[34][20] ), .CLK(clk), .RST(rst), .I(g_init[1108]), .Q(\Inst_Mem/inst_mem_reg[34][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][21]  ( .D(\Inst_Mem/inst_mem_reg[34][21] ), .CLK(clk), .RST(rst), .I(g_init[1109]), .Q(\Inst_Mem/inst_mem_reg[34][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][22]  ( .D(\Inst_Mem/inst_mem_reg[34][22] ), .CLK(clk), .RST(rst), .I(g_init[1110]), .Q(\Inst_Mem/inst_mem_reg[34][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][23]  ( .D(\Inst_Mem/inst_mem_reg[34][23] ), .CLK(clk), .RST(rst), .I(g_init[1111]), .Q(\Inst_Mem/inst_mem_reg[34][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][24]  ( .D(\Inst_Mem/inst_mem_reg[34][24] ), .CLK(clk), .RST(rst), .I(g_init[1112]), .Q(\Inst_Mem/inst_mem_reg[34][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][25]  ( .D(\Inst_Mem/inst_mem_reg[34][25] ), .CLK(clk), .RST(rst), .I(g_init[1113]), .Q(\Inst_Mem/inst_mem_reg[34][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][26]  ( .D(\Inst_Mem/inst_mem_reg[34][26] ), .CLK(clk), .RST(rst), .I(g_init[1114]), .Q(\Inst_Mem/inst_mem_reg[34][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][27]  ( .D(\Inst_Mem/inst_mem_reg[34][27] ), .CLK(clk), .RST(rst), .I(g_init[1115]), .Q(\Inst_Mem/inst_mem_reg[34][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][28]  ( .D(\Inst_Mem/inst_mem_reg[34][28] ), .CLK(clk), .RST(rst), .I(g_init[1116]), .Q(\Inst_Mem/inst_mem_reg[34][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][29]  ( .D(\Inst_Mem/inst_mem_reg[34][29] ), .CLK(clk), .RST(rst), .I(g_init[1117]), .Q(\Inst_Mem/inst_mem_reg[34][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][30]  ( .D(\Inst_Mem/inst_mem_reg[34][30] ), .CLK(clk), .RST(rst), .I(g_init[1118]), .Q(\Inst_Mem/inst_mem_reg[34][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[34][31]  ( .D(\Inst_Mem/inst_mem_reg[34][31] ), .CLK(clk), .RST(rst), .I(g_init[1119]), .Q(\Inst_Mem/inst_mem_reg[34][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][0]  ( .D(\Inst_Mem/inst_mem_reg[33][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1056]), .Q(
        \Inst_Mem/inst_mem_reg[33][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][1]  ( .D(\Inst_Mem/inst_mem_reg[33][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1057]), .Q(
        \Inst_Mem/inst_mem_reg[33][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][2]  ( .D(\Inst_Mem/inst_mem_reg[33][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1058]), .Q(
        \Inst_Mem/inst_mem_reg[33][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][3]  ( .D(\Inst_Mem/inst_mem_reg[33][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1059]), .Q(
        \Inst_Mem/inst_mem_reg[33][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][4]  ( .D(\Inst_Mem/inst_mem_reg[33][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1060]), .Q(
        \Inst_Mem/inst_mem_reg[33][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][5]  ( .D(\Inst_Mem/inst_mem_reg[33][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1061]), .Q(
        \Inst_Mem/inst_mem_reg[33][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][6]  ( .D(\Inst_Mem/inst_mem_reg[33][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1062]), .Q(
        \Inst_Mem/inst_mem_reg[33][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][7]  ( .D(\Inst_Mem/inst_mem_reg[33][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1063]), .Q(
        \Inst_Mem/inst_mem_reg[33][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][8]  ( .D(\Inst_Mem/inst_mem_reg[33][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1064]), .Q(
        \Inst_Mem/inst_mem_reg[33][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][9]  ( .D(\Inst_Mem/inst_mem_reg[33][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1065]), .Q(
        \Inst_Mem/inst_mem_reg[33][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[33][10]  ( .D(\Inst_Mem/inst_mem_reg[33][10] ), .CLK(clk), .RST(rst), .I(g_init[1066]), .Q(\Inst_Mem/inst_mem_reg[33][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][11]  ( .D(\Inst_Mem/inst_mem_reg[33][11] ), .CLK(clk), .RST(rst), .I(g_init[1067]), .Q(\Inst_Mem/inst_mem_reg[33][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][12]  ( .D(\Inst_Mem/inst_mem_reg[33][12] ), .CLK(clk), .RST(rst), .I(g_init[1068]), .Q(\Inst_Mem/inst_mem_reg[33][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][13]  ( .D(\Inst_Mem/inst_mem_reg[33][13] ), .CLK(clk), .RST(rst), .I(g_init[1069]), .Q(\Inst_Mem/inst_mem_reg[33][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][14]  ( .D(\Inst_Mem/inst_mem_reg[33][14] ), .CLK(clk), .RST(rst), .I(g_init[1070]), .Q(\Inst_Mem/inst_mem_reg[33][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][15]  ( .D(\Inst_Mem/inst_mem_reg[33][15] ), .CLK(clk), .RST(rst), .I(g_init[1071]), .Q(\Inst_Mem/inst_mem_reg[33][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][16]  ( .D(\Inst_Mem/inst_mem_reg[33][16] ), .CLK(clk), .RST(rst), .I(g_init[1072]), .Q(\Inst_Mem/inst_mem_reg[33][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][17]  ( .D(\Inst_Mem/inst_mem_reg[33][17] ), .CLK(clk), .RST(rst), .I(g_init[1073]), .Q(\Inst_Mem/inst_mem_reg[33][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][18]  ( .D(\Inst_Mem/inst_mem_reg[33][18] ), .CLK(clk), .RST(rst), .I(g_init[1074]), .Q(\Inst_Mem/inst_mem_reg[33][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][19]  ( .D(\Inst_Mem/inst_mem_reg[33][19] ), .CLK(clk), .RST(rst), .I(g_init[1075]), .Q(\Inst_Mem/inst_mem_reg[33][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][20]  ( .D(\Inst_Mem/inst_mem_reg[33][20] ), .CLK(clk), .RST(rst), .I(g_init[1076]), .Q(\Inst_Mem/inst_mem_reg[33][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][21]  ( .D(\Inst_Mem/inst_mem_reg[33][21] ), .CLK(clk), .RST(rst), .I(g_init[1077]), .Q(\Inst_Mem/inst_mem_reg[33][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][22]  ( .D(\Inst_Mem/inst_mem_reg[33][22] ), .CLK(clk), .RST(rst), .I(g_init[1078]), .Q(\Inst_Mem/inst_mem_reg[33][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][23]  ( .D(\Inst_Mem/inst_mem_reg[33][23] ), .CLK(clk), .RST(rst), .I(g_init[1079]), .Q(\Inst_Mem/inst_mem_reg[33][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][24]  ( .D(\Inst_Mem/inst_mem_reg[33][24] ), .CLK(clk), .RST(rst), .I(g_init[1080]), .Q(\Inst_Mem/inst_mem_reg[33][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][25]  ( .D(\Inst_Mem/inst_mem_reg[33][25] ), .CLK(clk), .RST(rst), .I(g_init[1081]), .Q(\Inst_Mem/inst_mem_reg[33][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][26]  ( .D(\Inst_Mem/inst_mem_reg[33][26] ), .CLK(clk), .RST(rst), .I(g_init[1082]), .Q(\Inst_Mem/inst_mem_reg[33][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][27]  ( .D(\Inst_Mem/inst_mem_reg[33][27] ), .CLK(clk), .RST(rst), .I(g_init[1083]), .Q(\Inst_Mem/inst_mem_reg[33][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][28]  ( .D(\Inst_Mem/inst_mem_reg[33][28] ), .CLK(clk), .RST(rst), .I(g_init[1084]), .Q(\Inst_Mem/inst_mem_reg[33][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][29]  ( .D(\Inst_Mem/inst_mem_reg[33][29] ), .CLK(clk), .RST(rst), .I(g_init[1085]), .Q(\Inst_Mem/inst_mem_reg[33][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][30]  ( .D(\Inst_Mem/inst_mem_reg[33][30] ), .CLK(clk), .RST(rst), .I(g_init[1086]), .Q(\Inst_Mem/inst_mem_reg[33][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[33][31]  ( .D(\Inst_Mem/inst_mem_reg[33][31] ), .CLK(clk), .RST(rst), .I(g_init[1087]), .Q(\Inst_Mem/inst_mem_reg[33][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][0]  ( .D(\Inst_Mem/inst_mem_reg[32][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[1024]), .Q(
        \Inst_Mem/inst_mem_reg[32][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][1]  ( .D(\Inst_Mem/inst_mem_reg[32][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1025]), .Q(
        \Inst_Mem/inst_mem_reg[32][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][2]  ( .D(\Inst_Mem/inst_mem_reg[32][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[1026]), .Q(
        \Inst_Mem/inst_mem_reg[32][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][3]  ( .D(\Inst_Mem/inst_mem_reg[32][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[1027]), .Q(
        \Inst_Mem/inst_mem_reg[32][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][4]  ( .D(\Inst_Mem/inst_mem_reg[32][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[1028]), .Q(
        \Inst_Mem/inst_mem_reg[32][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][5]  ( .D(\Inst_Mem/inst_mem_reg[32][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[1029]), .Q(
        \Inst_Mem/inst_mem_reg[32][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][6]  ( .D(\Inst_Mem/inst_mem_reg[32][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[1030]), .Q(
        \Inst_Mem/inst_mem_reg[32][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][7]  ( .D(\Inst_Mem/inst_mem_reg[32][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[1031]), .Q(
        \Inst_Mem/inst_mem_reg[32][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][8]  ( .D(\Inst_Mem/inst_mem_reg[32][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1032]), .Q(
        \Inst_Mem/inst_mem_reg[32][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][9]  ( .D(\Inst_Mem/inst_mem_reg[32][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1033]), .Q(
        \Inst_Mem/inst_mem_reg[32][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[32][10]  ( .D(\Inst_Mem/inst_mem_reg[32][10] ), .CLK(clk), .RST(rst), .I(g_init[1034]), .Q(\Inst_Mem/inst_mem_reg[32][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][11]  ( .D(\Inst_Mem/inst_mem_reg[32][11] ), .CLK(clk), .RST(rst), .I(g_init[1035]), .Q(\Inst_Mem/inst_mem_reg[32][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][12]  ( .D(\Inst_Mem/inst_mem_reg[32][12] ), .CLK(clk), .RST(rst), .I(g_init[1036]), .Q(\Inst_Mem/inst_mem_reg[32][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][13]  ( .D(\Inst_Mem/inst_mem_reg[32][13] ), .CLK(clk), .RST(rst), .I(g_init[1037]), .Q(\Inst_Mem/inst_mem_reg[32][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][14]  ( .D(\Inst_Mem/inst_mem_reg[32][14] ), .CLK(clk), .RST(rst), .I(g_init[1038]), .Q(\Inst_Mem/inst_mem_reg[32][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][15]  ( .D(\Inst_Mem/inst_mem_reg[32][15] ), .CLK(clk), .RST(rst), .I(g_init[1039]), .Q(\Inst_Mem/inst_mem_reg[32][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][16]  ( .D(\Inst_Mem/inst_mem_reg[32][16] ), .CLK(clk), .RST(rst), .I(g_init[1040]), .Q(\Inst_Mem/inst_mem_reg[32][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][17]  ( .D(\Inst_Mem/inst_mem_reg[32][17] ), .CLK(clk), .RST(rst), .I(g_init[1041]), .Q(\Inst_Mem/inst_mem_reg[32][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][18]  ( .D(\Inst_Mem/inst_mem_reg[32][18] ), .CLK(clk), .RST(rst), .I(g_init[1042]), .Q(\Inst_Mem/inst_mem_reg[32][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][19]  ( .D(\Inst_Mem/inst_mem_reg[32][19] ), .CLK(clk), .RST(rst), .I(g_init[1043]), .Q(\Inst_Mem/inst_mem_reg[32][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][20]  ( .D(\Inst_Mem/inst_mem_reg[32][20] ), .CLK(clk), .RST(rst), .I(g_init[1044]), .Q(\Inst_Mem/inst_mem_reg[32][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][21]  ( .D(\Inst_Mem/inst_mem_reg[32][21] ), .CLK(clk), .RST(rst), .I(g_init[1045]), .Q(\Inst_Mem/inst_mem_reg[32][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][22]  ( .D(\Inst_Mem/inst_mem_reg[32][22] ), .CLK(clk), .RST(rst), .I(g_init[1046]), .Q(\Inst_Mem/inst_mem_reg[32][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][23]  ( .D(\Inst_Mem/inst_mem_reg[32][23] ), .CLK(clk), .RST(rst), .I(g_init[1047]), .Q(\Inst_Mem/inst_mem_reg[32][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][24]  ( .D(\Inst_Mem/inst_mem_reg[32][24] ), .CLK(clk), .RST(rst), .I(g_init[1048]), .Q(\Inst_Mem/inst_mem_reg[32][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][25]  ( .D(\Inst_Mem/inst_mem_reg[32][25] ), .CLK(clk), .RST(rst), .I(g_init[1049]), .Q(\Inst_Mem/inst_mem_reg[32][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][26]  ( .D(\Inst_Mem/inst_mem_reg[32][26] ), .CLK(clk), .RST(rst), .I(g_init[1050]), .Q(\Inst_Mem/inst_mem_reg[32][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][27]  ( .D(\Inst_Mem/inst_mem_reg[32][27] ), .CLK(clk), .RST(rst), .I(g_init[1051]), .Q(\Inst_Mem/inst_mem_reg[32][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][28]  ( .D(\Inst_Mem/inst_mem_reg[32][28] ), .CLK(clk), .RST(rst), .I(g_init[1052]), .Q(\Inst_Mem/inst_mem_reg[32][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][29]  ( .D(\Inst_Mem/inst_mem_reg[32][29] ), .CLK(clk), .RST(rst), .I(g_init[1053]), .Q(\Inst_Mem/inst_mem_reg[32][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][30]  ( .D(\Inst_Mem/inst_mem_reg[32][30] ), .CLK(clk), .RST(rst), .I(g_init[1054]), .Q(\Inst_Mem/inst_mem_reg[32][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[32][31]  ( .D(\Inst_Mem/inst_mem_reg[32][31] ), .CLK(clk), .RST(rst), .I(g_init[1055]), .Q(\Inst_Mem/inst_mem_reg[32][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][0]  ( .D(\Inst_Mem/inst_mem_reg[31][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[992]), .Q(
        \Inst_Mem/inst_mem_reg[31][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][1]  ( .D(\Inst_Mem/inst_mem_reg[31][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[993]), .Q(
        \Inst_Mem/inst_mem_reg[31][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][2]  ( .D(\Inst_Mem/inst_mem_reg[31][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[994]), .Q(
        \Inst_Mem/inst_mem_reg[31][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][3]  ( .D(\Inst_Mem/inst_mem_reg[31][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[995]), .Q(
        \Inst_Mem/inst_mem_reg[31][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][4]  ( .D(\Inst_Mem/inst_mem_reg[31][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[996]), .Q(
        \Inst_Mem/inst_mem_reg[31][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][5]  ( .D(\Inst_Mem/inst_mem_reg[31][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[997]), .Q(
        \Inst_Mem/inst_mem_reg[31][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][6]  ( .D(\Inst_Mem/inst_mem_reg[31][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[998]), .Q(
        \Inst_Mem/inst_mem_reg[31][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][7]  ( .D(\Inst_Mem/inst_mem_reg[31][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[999]), .Q(
        \Inst_Mem/inst_mem_reg[31][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][8]  ( .D(\Inst_Mem/inst_mem_reg[31][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[1000]), .Q(
        \Inst_Mem/inst_mem_reg[31][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][9]  ( .D(\Inst_Mem/inst_mem_reg[31][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[1001]), .Q(
        \Inst_Mem/inst_mem_reg[31][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[31][10]  ( .D(\Inst_Mem/inst_mem_reg[31][10] ), .CLK(clk), .RST(rst), .I(g_init[1002]), .Q(\Inst_Mem/inst_mem_reg[31][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][11]  ( .D(\Inst_Mem/inst_mem_reg[31][11] ), .CLK(clk), .RST(rst), .I(g_init[1003]), .Q(\Inst_Mem/inst_mem_reg[31][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][12]  ( .D(\Inst_Mem/inst_mem_reg[31][12] ), .CLK(clk), .RST(rst), .I(g_init[1004]), .Q(\Inst_Mem/inst_mem_reg[31][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][13]  ( .D(\Inst_Mem/inst_mem_reg[31][13] ), .CLK(clk), .RST(rst), .I(g_init[1005]), .Q(\Inst_Mem/inst_mem_reg[31][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][14]  ( .D(\Inst_Mem/inst_mem_reg[31][14] ), .CLK(clk), .RST(rst), .I(g_init[1006]), .Q(\Inst_Mem/inst_mem_reg[31][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][15]  ( .D(\Inst_Mem/inst_mem_reg[31][15] ), .CLK(clk), .RST(rst), .I(g_init[1007]), .Q(\Inst_Mem/inst_mem_reg[31][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][16]  ( .D(\Inst_Mem/inst_mem_reg[31][16] ), .CLK(clk), .RST(rst), .I(g_init[1008]), .Q(\Inst_Mem/inst_mem_reg[31][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][17]  ( .D(\Inst_Mem/inst_mem_reg[31][17] ), .CLK(clk), .RST(rst), .I(g_init[1009]), .Q(\Inst_Mem/inst_mem_reg[31][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][18]  ( .D(\Inst_Mem/inst_mem_reg[31][18] ), .CLK(clk), .RST(rst), .I(g_init[1010]), .Q(\Inst_Mem/inst_mem_reg[31][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][19]  ( .D(\Inst_Mem/inst_mem_reg[31][19] ), .CLK(clk), .RST(rst), .I(g_init[1011]), .Q(\Inst_Mem/inst_mem_reg[31][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][20]  ( .D(\Inst_Mem/inst_mem_reg[31][20] ), .CLK(clk), .RST(rst), .I(g_init[1012]), .Q(\Inst_Mem/inst_mem_reg[31][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][21]  ( .D(\Inst_Mem/inst_mem_reg[31][21] ), .CLK(clk), .RST(rst), .I(g_init[1013]), .Q(\Inst_Mem/inst_mem_reg[31][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][22]  ( .D(\Inst_Mem/inst_mem_reg[31][22] ), .CLK(clk), .RST(rst), .I(g_init[1014]), .Q(\Inst_Mem/inst_mem_reg[31][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][23]  ( .D(\Inst_Mem/inst_mem_reg[31][23] ), .CLK(clk), .RST(rst), .I(g_init[1015]), .Q(\Inst_Mem/inst_mem_reg[31][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][24]  ( .D(\Inst_Mem/inst_mem_reg[31][24] ), .CLK(clk), .RST(rst), .I(g_init[1016]), .Q(\Inst_Mem/inst_mem_reg[31][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][25]  ( .D(\Inst_Mem/inst_mem_reg[31][25] ), .CLK(clk), .RST(rst), .I(g_init[1017]), .Q(\Inst_Mem/inst_mem_reg[31][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][26]  ( .D(\Inst_Mem/inst_mem_reg[31][26] ), .CLK(clk), .RST(rst), .I(g_init[1018]), .Q(\Inst_Mem/inst_mem_reg[31][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][27]  ( .D(\Inst_Mem/inst_mem_reg[31][27] ), .CLK(clk), .RST(rst), .I(g_init[1019]), .Q(\Inst_Mem/inst_mem_reg[31][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][28]  ( .D(\Inst_Mem/inst_mem_reg[31][28] ), .CLK(clk), .RST(rst), .I(g_init[1020]), .Q(\Inst_Mem/inst_mem_reg[31][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][29]  ( .D(\Inst_Mem/inst_mem_reg[31][29] ), .CLK(clk), .RST(rst), .I(g_init[1021]), .Q(\Inst_Mem/inst_mem_reg[31][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][30]  ( .D(\Inst_Mem/inst_mem_reg[31][30] ), .CLK(clk), .RST(rst), .I(g_init[1022]), .Q(\Inst_Mem/inst_mem_reg[31][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[31][31]  ( .D(\Inst_Mem/inst_mem_reg[31][31] ), .CLK(clk), .RST(rst), .I(g_init[1023]), .Q(\Inst_Mem/inst_mem_reg[31][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][0]  ( .D(\Inst_Mem/inst_mem_reg[30][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[960]), .Q(
        \Inst_Mem/inst_mem_reg[30][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][1]  ( .D(\Inst_Mem/inst_mem_reg[30][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[961]), .Q(
        \Inst_Mem/inst_mem_reg[30][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][2]  ( .D(\Inst_Mem/inst_mem_reg[30][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[962]), .Q(
        \Inst_Mem/inst_mem_reg[30][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][3]  ( .D(\Inst_Mem/inst_mem_reg[30][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[963]), .Q(
        \Inst_Mem/inst_mem_reg[30][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][4]  ( .D(\Inst_Mem/inst_mem_reg[30][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[964]), .Q(
        \Inst_Mem/inst_mem_reg[30][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][5]  ( .D(\Inst_Mem/inst_mem_reg[30][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[965]), .Q(
        \Inst_Mem/inst_mem_reg[30][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][6]  ( .D(\Inst_Mem/inst_mem_reg[30][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[966]), .Q(
        \Inst_Mem/inst_mem_reg[30][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][7]  ( .D(\Inst_Mem/inst_mem_reg[30][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[967]), .Q(
        \Inst_Mem/inst_mem_reg[30][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][8]  ( .D(\Inst_Mem/inst_mem_reg[30][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[968]), .Q(
        \Inst_Mem/inst_mem_reg[30][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][9]  ( .D(\Inst_Mem/inst_mem_reg[30][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[969]), .Q(
        \Inst_Mem/inst_mem_reg[30][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[30][10]  ( .D(\Inst_Mem/inst_mem_reg[30][10] ), .CLK(clk), .RST(rst), .I(g_init[970]), .Q(\Inst_Mem/inst_mem_reg[30][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][11]  ( .D(\Inst_Mem/inst_mem_reg[30][11] ), .CLK(clk), .RST(rst), .I(g_init[971]), .Q(\Inst_Mem/inst_mem_reg[30][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][12]  ( .D(\Inst_Mem/inst_mem_reg[30][12] ), .CLK(clk), .RST(rst), .I(g_init[972]), .Q(\Inst_Mem/inst_mem_reg[30][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][13]  ( .D(\Inst_Mem/inst_mem_reg[30][13] ), .CLK(clk), .RST(rst), .I(g_init[973]), .Q(\Inst_Mem/inst_mem_reg[30][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][14]  ( .D(\Inst_Mem/inst_mem_reg[30][14] ), .CLK(clk), .RST(rst), .I(g_init[974]), .Q(\Inst_Mem/inst_mem_reg[30][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][15]  ( .D(\Inst_Mem/inst_mem_reg[30][15] ), .CLK(clk), .RST(rst), .I(g_init[975]), .Q(\Inst_Mem/inst_mem_reg[30][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][16]  ( .D(\Inst_Mem/inst_mem_reg[30][16] ), .CLK(clk), .RST(rst), .I(g_init[976]), .Q(\Inst_Mem/inst_mem_reg[30][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][17]  ( .D(\Inst_Mem/inst_mem_reg[30][17] ), .CLK(clk), .RST(rst), .I(g_init[977]), .Q(\Inst_Mem/inst_mem_reg[30][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][18]  ( .D(\Inst_Mem/inst_mem_reg[30][18] ), .CLK(clk), .RST(rst), .I(g_init[978]), .Q(\Inst_Mem/inst_mem_reg[30][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][19]  ( .D(\Inst_Mem/inst_mem_reg[30][19] ), .CLK(clk), .RST(rst), .I(g_init[979]), .Q(\Inst_Mem/inst_mem_reg[30][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][20]  ( .D(\Inst_Mem/inst_mem_reg[30][20] ), .CLK(clk), .RST(rst), .I(g_init[980]), .Q(\Inst_Mem/inst_mem_reg[30][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][21]  ( .D(\Inst_Mem/inst_mem_reg[30][21] ), .CLK(clk), .RST(rst), .I(g_init[981]), .Q(\Inst_Mem/inst_mem_reg[30][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][22]  ( .D(\Inst_Mem/inst_mem_reg[30][22] ), .CLK(clk), .RST(rst), .I(g_init[982]), .Q(\Inst_Mem/inst_mem_reg[30][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][23]  ( .D(\Inst_Mem/inst_mem_reg[30][23] ), .CLK(clk), .RST(rst), .I(g_init[983]), .Q(\Inst_Mem/inst_mem_reg[30][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][24]  ( .D(\Inst_Mem/inst_mem_reg[30][24] ), .CLK(clk), .RST(rst), .I(g_init[984]), .Q(\Inst_Mem/inst_mem_reg[30][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][25]  ( .D(\Inst_Mem/inst_mem_reg[30][25] ), .CLK(clk), .RST(rst), .I(g_init[985]), .Q(\Inst_Mem/inst_mem_reg[30][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][26]  ( .D(\Inst_Mem/inst_mem_reg[30][26] ), .CLK(clk), .RST(rst), .I(g_init[986]), .Q(\Inst_Mem/inst_mem_reg[30][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][27]  ( .D(\Inst_Mem/inst_mem_reg[30][27] ), .CLK(clk), .RST(rst), .I(g_init[987]), .Q(\Inst_Mem/inst_mem_reg[30][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][28]  ( .D(\Inst_Mem/inst_mem_reg[30][28] ), .CLK(clk), .RST(rst), .I(g_init[988]), .Q(\Inst_Mem/inst_mem_reg[30][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][29]  ( .D(\Inst_Mem/inst_mem_reg[30][29] ), .CLK(clk), .RST(rst), .I(g_init[989]), .Q(\Inst_Mem/inst_mem_reg[30][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][30]  ( .D(\Inst_Mem/inst_mem_reg[30][30] ), .CLK(clk), .RST(rst), .I(g_init[990]), .Q(\Inst_Mem/inst_mem_reg[30][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[30][31]  ( .D(\Inst_Mem/inst_mem_reg[30][31] ), .CLK(clk), .RST(rst), .I(g_init[991]), .Q(\Inst_Mem/inst_mem_reg[30][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][0]  ( .D(\Inst_Mem/inst_mem_reg[29][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[928]), .Q(
        \Inst_Mem/inst_mem_reg[29][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][1]  ( .D(\Inst_Mem/inst_mem_reg[29][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[929]), .Q(
        \Inst_Mem/inst_mem_reg[29][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][2]  ( .D(\Inst_Mem/inst_mem_reg[29][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[930]), .Q(
        \Inst_Mem/inst_mem_reg[29][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][3]  ( .D(\Inst_Mem/inst_mem_reg[29][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[931]), .Q(
        \Inst_Mem/inst_mem_reg[29][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][4]  ( .D(\Inst_Mem/inst_mem_reg[29][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[932]), .Q(
        \Inst_Mem/inst_mem_reg[29][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][5]  ( .D(\Inst_Mem/inst_mem_reg[29][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[933]), .Q(
        \Inst_Mem/inst_mem_reg[29][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][6]  ( .D(\Inst_Mem/inst_mem_reg[29][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[934]), .Q(
        \Inst_Mem/inst_mem_reg[29][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][7]  ( .D(\Inst_Mem/inst_mem_reg[29][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[935]), .Q(
        \Inst_Mem/inst_mem_reg[29][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][8]  ( .D(\Inst_Mem/inst_mem_reg[29][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[936]), .Q(
        \Inst_Mem/inst_mem_reg[29][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][9]  ( .D(\Inst_Mem/inst_mem_reg[29][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[937]), .Q(
        \Inst_Mem/inst_mem_reg[29][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[29][10]  ( .D(\Inst_Mem/inst_mem_reg[29][10] ), .CLK(clk), .RST(rst), .I(g_init[938]), .Q(\Inst_Mem/inst_mem_reg[29][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][11]  ( .D(\Inst_Mem/inst_mem_reg[29][11] ), .CLK(clk), .RST(rst), .I(g_init[939]), .Q(\Inst_Mem/inst_mem_reg[29][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][12]  ( .D(\Inst_Mem/inst_mem_reg[29][12] ), .CLK(clk), .RST(rst), .I(g_init[940]), .Q(\Inst_Mem/inst_mem_reg[29][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][13]  ( .D(\Inst_Mem/inst_mem_reg[29][13] ), .CLK(clk), .RST(rst), .I(g_init[941]), .Q(\Inst_Mem/inst_mem_reg[29][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][14]  ( .D(\Inst_Mem/inst_mem_reg[29][14] ), .CLK(clk), .RST(rst), .I(g_init[942]), .Q(\Inst_Mem/inst_mem_reg[29][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][15]  ( .D(\Inst_Mem/inst_mem_reg[29][15] ), .CLK(clk), .RST(rst), .I(g_init[943]), .Q(\Inst_Mem/inst_mem_reg[29][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][16]  ( .D(\Inst_Mem/inst_mem_reg[29][16] ), .CLK(clk), .RST(rst), .I(g_init[944]), .Q(\Inst_Mem/inst_mem_reg[29][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][17]  ( .D(\Inst_Mem/inst_mem_reg[29][17] ), .CLK(clk), .RST(rst), .I(g_init[945]), .Q(\Inst_Mem/inst_mem_reg[29][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][18]  ( .D(\Inst_Mem/inst_mem_reg[29][18] ), .CLK(clk), .RST(rst), .I(g_init[946]), .Q(\Inst_Mem/inst_mem_reg[29][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][19]  ( .D(\Inst_Mem/inst_mem_reg[29][19] ), .CLK(clk), .RST(rst), .I(g_init[947]), .Q(\Inst_Mem/inst_mem_reg[29][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][20]  ( .D(\Inst_Mem/inst_mem_reg[29][20] ), .CLK(clk), .RST(rst), .I(g_init[948]), .Q(\Inst_Mem/inst_mem_reg[29][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][21]  ( .D(\Inst_Mem/inst_mem_reg[29][21] ), .CLK(clk), .RST(rst), .I(g_init[949]), .Q(\Inst_Mem/inst_mem_reg[29][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][22]  ( .D(\Inst_Mem/inst_mem_reg[29][22] ), .CLK(clk), .RST(rst), .I(g_init[950]), .Q(\Inst_Mem/inst_mem_reg[29][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][23]  ( .D(\Inst_Mem/inst_mem_reg[29][23] ), .CLK(clk), .RST(rst), .I(g_init[951]), .Q(\Inst_Mem/inst_mem_reg[29][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][24]  ( .D(\Inst_Mem/inst_mem_reg[29][24] ), .CLK(clk), .RST(rst), .I(g_init[952]), .Q(\Inst_Mem/inst_mem_reg[29][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][25]  ( .D(\Inst_Mem/inst_mem_reg[29][25] ), .CLK(clk), .RST(rst), .I(g_init[953]), .Q(\Inst_Mem/inst_mem_reg[29][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][26]  ( .D(\Inst_Mem/inst_mem_reg[29][26] ), .CLK(clk), .RST(rst), .I(g_init[954]), .Q(\Inst_Mem/inst_mem_reg[29][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][27]  ( .D(\Inst_Mem/inst_mem_reg[29][27] ), .CLK(clk), .RST(rst), .I(g_init[955]), .Q(\Inst_Mem/inst_mem_reg[29][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][28]  ( .D(\Inst_Mem/inst_mem_reg[29][28] ), .CLK(clk), .RST(rst), .I(g_init[956]), .Q(\Inst_Mem/inst_mem_reg[29][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][29]  ( .D(\Inst_Mem/inst_mem_reg[29][29] ), .CLK(clk), .RST(rst), .I(g_init[957]), .Q(\Inst_Mem/inst_mem_reg[29][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][30]  ( .D(\Inst_Mem/inst_mem_reg[29][30] ), .CLK(clk), .RST(rst), .I(g_init[958]), .Q(\Inst_Mem/inst_mem_reg[29][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[29][31]  ( .D(\Inst_Mem/inst_mem_reg[29][31] ), .CLK(clk), .RST(rst), .I(g_init[959]), .Q(\Inst_Mem/inst_mem_reg[29][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][0]  ( .D(\Inst_Mem/inst_mem_reg[28][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[896]), .Q(
        \Inst_Mem/inst_mem_reg[28][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][1]  ( .D(\Inst_Mem/inst_mem_reg[28][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[897]), .Q(
        \Inst_Mem/inst_mem_reg[28][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][2]  ( .D(\Inst_Mem/inst_mem_reg[28][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[898]), .Q(
        \Inst_Mem/inst_mem_reg[28][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][3]  ( .D(\Inst_Mem/inst_mem_reg[28][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[899]), .Q(
        \Inst_Mem/inst_mem_reg[28][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][4]  ( .D(\Inst_Mem/inst_mem_reg[28][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[900]), .Q(
        \Inst_Mem/inst_mem_reg[28][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][5]  ( .D(\Inst_Mem/inst_mem_reg[28][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[901]), .Q(
        \Inst_Mem/inst_mem_reg[28][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][6]  ( .D(\Inst_Mem/inst_mem_reg[28][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[902]), .Q(
        \Inst_Mem/inst_mem_reg[28][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][7]  ( .D(\Inst_Mem/inst_mem_reg[28][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[903]), .Q(
        \Inst_Mem/inst_mem_reg[28][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][8]  ( .D(\Inst_Mem/inst_mem_reg[28][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[904]), .Q(
        \Inst_Mem/inst_mem_reg[28][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][9]  ( .D(\Inst_Mem/inst_mem_reg[28][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[905]), .Q(
        \Inst_Mem/inst_mem_reg[28][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[28][10]  ( .D(\Inst_Mem/inst_mem_reg[28][10] ), .CLK(clk), .RST(rst), .I(g_init[906]), .Q(\Inst_Mem/inst_mem_reg[28][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][11]  ( .D(\Inst_Mem/inst_mem_reg[28][11] ), .CLK(clk), .RST(rst), .I(g_init[907]), .Q(\Inst_Mem/inst_mem_reg[28][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][12]  ( .D(\Inst_Mem/inst_mem_reg[28][12] ), .CLK(clk), .RST(rst), .I(g_init[908]), .Q(\Inst_Mem/inst_mem_reg[28][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][13]  ( .D(\Inst_Mem/inst_mem_reg[28][13] ), .CLK(clk), .RST(rst), .I(g_init[909]), .Q(\Inst_Mem/inst_mem_reg[28][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][14]  ( .D(\Inst_Mem/inst_mem_reg[28][14] ), .CLK(clk), .RST(rst), .I(g_init[910]), .Q(\Inst_Mem/inst_mem_reg[28][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][15]  ( .D(\Inst_Mem/inst_mem_reg[28][15] ), .CLK(clk), .RST(rst), .I(g_init[911]), .Q(\Inst_Mem/inst_mem_reg[28][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][16]  ( .D(\Inst_Mem/inst_mem_reg[28][16] ), .CLK(clk), .RST(rst), .I(g_init[912]), .Q(\Inst_Mem/inst_mem_reg[28][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][17]  ( .D(\Inst_Mem/inst_mem_reg[28][17] ), .CLK(clk), .RST(rst), .I(g_init[913]), .Q(\Inst_Mem/inst_mem_reg[28][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][18]  ( .D(\Inst_Mem/inst_mem_reg[28][18] ), .CLK(clk), .RST(rst), .I(g_init[914]), .Q(\Inst_Mem/inst_mem_reg[28][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][19]  ( .D(\Inst_Mem/inst_mem_reg[28][19] ), .CLK(clk), .RST(rst), .I(g_init[915]), .Q(\Inst_Mem/inst_mem_reg[28][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][20]  ( .D(\Inst_Mem/inst_mem_reg[28][20] ), .CLK(clk), .RST(rst), .I(g_init[916]), .Q(\Inst_Mem/inst_mem_reg[28][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][21]  ( .D(\Inst_Mem/inst_mem_reg[28][21] ), .CLK(clk), .RST(rst), .I(g_init[917]), .Q(\Inst_Mem/inst_mem_reg[28][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][22]  ( .D(\Inst_Mem/inst_mem_reg[28][22] ), .CLK(clk), .RST(rst), .I(g_init[918]), .Q(\Inst_Mem/inst_mem_reg[28][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][23]  ( .D(\Inst_Mem/inst_mem_reg[28][23] ), .CLK(clk), .RST(rst), .I(g_init[919]), .Q(\Inst_Mem/inst_mem_reg[28][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][24]  ( .D(\Inst_Mem/inst_mem_reg[28][24] ), .CLK(clk), .RST(rst), .I(g_init[920]), .Q(\Inst_Mem/inst_mem_reg[28][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][25]  ( .D(\Inst_Mem/inst_mem_reg[28][25] ), .CLK(clk), .RST(rst), .I(g_init[921]), .Q(\Inst_Mem/inst_mem_reg[28][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][26]  ( .D(\Inst_Mem/inst_mem_reg[28][26] ), .CLK(clk), .RST(rst), .I(g_init[922]), .Q(\Inst_Mem/inst_mem_reg[28][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][27]  ( .D(\Inst_Mem/inst_mem_reg[28][27] ), .CLK(clk), .RST(rst), .I(g_init[923]), .Q(\Inst_Mem/inst_mem_reg[28][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][28]  ( .D(\Inst_Mem/inst_mem_reg[28][28] ), .CLK(clk), .RST(rst), .I(g_init[924]), .Q(\Inst_Mem/inst_mem_reg[28][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][29]  ( .D(\Inst_Mem/inst_mem_reg[28][29] ), .CLK(clk), .RST(rst), .I(g_init[925]), .Q(\Inst_Mem/inst_mem_reg[28][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][30]  ( .D(\Inst_Mem/inst_mem_reg[28][30] ), .CLK(clk), .RST(rst), .I(g_init[926]), .Q(\Inst_Mem/inst_mem_reg[28][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[28][31]  ( .D(\Inst_Mem/inst_mem_reg[28][31] ), .CLK(clk), .RST(rst), .I(g_init[927]), .Q(\Inst_Mem/inst_mem_reg[28][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][0]  ( .D(\Inst_Mem/inst_mem_reg[27][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[864]), .Q(
        \Inst_Mem/inst_mem_reg[27][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][1]  ( .D(\Inst_Mem/inst_mem_reg[27][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[865]), .Q(
        \Inst_Mem/inst_mem_reg[27][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][2]  ( .D(\Inst_Mem/inst_mem_reg[27][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[866]), .Q(
        \Inst_Mem/inst_mem_reg[27][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][3]  ( .D(\Inst_Mem/inst_mem_reg[27][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[867]), .Q(
        \Inst_Mem/inst_mem_reg[27][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][4]  ( .D(\Inst_Mem/inst_mem_reg[27][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[868]), .Q(
        \Inst_Mem/inst_mem_reg[27][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][5]  ( .D(\Inst_Mem/inst_mem_reg[27][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[869]), .Q(
        \Inst_Mem/inst_mem_reg[27][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][6]  ( .D(\Inst_Mem/inst_mem_reg[27][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[870]), .Q(
        \Inst_Mem/inst_mem_reg[27][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][7]  ( .D(\Inst_Mem/inst_mem_reg[27][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[871]), .Q(
        \Inst_Mem/inst_mem_reg[27][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][8]  ( .D(\Inst_Mem/inst_mem_reg[27][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[872]), .Q(
        \Inst_Mem/inst_mem_reg[27][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][9]  ( .D(\Inst_Mem/inst_mem_reg[27][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[873]), .Q(
        \Inst_Mem/inst_mem_reg[27][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[27][10]  ( .D(\Inst_Mem/inst_mem_reg[27][10] ), .CLK(clk), .RST(rst), .I(g_init[874]), .Q(\Inst_Mem/inst_mem_reg[27][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][11]  ( .D(\Inst_Mem/inst_mem_reg[27][11] ), .CLK(clk), .RST(rst), .I(g_init[875]), .Q(\Inst_Mem/inst_mem_reg[27][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][12]  ( .D(\Inst_Mem/inst_mem_reg[27][12] ), .CLK(clk), .RST(rst), .I(g_init[876]), .Q(\Inst_Mem/inst_mem_reg[27][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][13]  ( .D(\Inst_Mem/inst_mem_reg[27][13] ), .CLK(clk), .RST(rst), .I(g_init[877]), .Q(\Inst_Mem/inst_mem_reg[27][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][14]  ( .D(\Inst_Mem/inst_mem_reg[27][14] ), .CLK(clk), .RST(rst), .I(g_init[878]), .Q(\Inst_Mem/inst_mem_reg[27][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][15]  ( .D(\Inst_Mem/inst_mem_reg[27][15] ), .CLK(clk), .RST(rst), .I(g_init[879]), .Q(\Inst_Mem/inst_mem_reg[27][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][16]  ( .D(\Inst_Mem/inst_mem_reg[27][16] ), .CLK(clk), .RST(rst), .I(g_init[880]), .Q(\Inst_Mem/inst_mem_reg[27][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][17]  ( .D(\Inst_Mem/inst_mem_reg[27][17] ), .CLK(clk), .RST(rst), .I(g_init[881]), .Q(\Inst_Mem/inst_mem_reg[27][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][18]  ( .D(\Inst_Mem/inst_mem_reg[27][18] ), .CLK(clk), .RST(rst), .I(g_init[882]), .Q(\Inst_Mem/inst_mem_reg[27][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][19]  ( .D(\Inst_Mem/inst_mem_reg[27][19] ), .CLK(clk), .RST(rst), .I(g_init[883]), .Q(\Inst_Mem/inst_mem_reg[27][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][20]  ( .D(\Inst_Mem/inst_mem_reg[27][20] ), .CLK(clk), .RST(rst), .I(g_init[884]), .Q(\Inst_Mem/inst_mem_reg[27][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][21]  ( .D(\Inst_Mem/inst_mem_reg[27][21] ), .CLK(clk), .RST(rst), .I(g_init[885]), .Q(\Inst_Mem/inst_mem_reg[27][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][22]  ( .D(\Inst_Mem/inst_mem_reg[27][22] ), .CLK(clk), .RST(rst), .I(g_init[886]), .Q(\Inst_Mem/inst_mem_reg[27][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][23]  ( .D(\Inst_Mem/inst_mem_reg[27][23] ), .CLK(clk), .RST(rst), .I(g_init[887]), .Q(\Inst_Mem/inst_mem_reg[27][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][24]  ( .D(\Inst_Mem/inst_mem_reg[27][24] ), .CLK(clk), .RST(rst), .I(g_init[888]), .Q(\Inst_Mem/inst_mem_reg[27][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][25]  ( .D(\Inst_Mem/inst_mem_reg[27][25] ), .CLK(clk), .RST(rst), .I(g_init[889]), .Q(\Inst_Mem/inst_mem_reg[27][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][26]  ( .D(\Inst_Mem/inst_mem_reg[27][26] ), .CLK(clk), .RST(rst), .I(g_init[890]), .Q(\Inst_Mem/inst_mem_reg[27][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][27]  ( .D(\Inst_Mem/inst_mem_reg[27][27] ), .CLK(clk), .RST(rst), .I(g_init[891]), .Q(\Inst_Mem/inst_mem_reg[27][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][28]  ( .D(\Inst_Mem/inst_mem_reg[27][28] ), .CLK(clk), .RST(rst), .I(g_init[892]), .Q(\Inst_Mem/inst_mem_reg[27][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][29]  ( .D(\Inst_Mem/inst_mem_reg[27][29] ), .CLK(clk), .RST(rst), .I(g_init[893]), .Q(\Inst_Mem/inst_mem_reg[27][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][30]  ( .D(\Inst_Mem/inst_mem_reg[27][30] ), .CLK(clk), .RST(rst), .I(g_init[894]), .Q(\Inst_Mem/inst_mem_reg[27][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[27][31]  ( .D(\Inst_Mem/inst_mem_reg[27][31] ), .CLK(clk), .RST(rst), .I(g_init[895]), .Q(\Inst_Mem/inst_mem_reg[27][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][0]  ( .D(\Inst_Mem/inst_mem_reg[26][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[832]), .Q(
        \Inst_Mem/inst_mem_reg[26][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][1]  ( .D(\Inst_Mem/inst_mem_reg[26][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[833]), .Q(
        \Inst_Mem/inst_mem_reg[26][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][2]  ( .D(\Inst_Mem/inst_mem_reg[26][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[834]), .Q(
        \Inst_Mem/inst_mem_reg[26][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][3]  ( .D(\Inst_Mem/inst_mem_reg[26][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[835]), .Q(
        \Inst_Mem/inst_mem_reg[26][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][4]  ( .D(\Inst_Mem/inst_mem_reg[26][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[836]), .Q(
        \Inst_Mem/inst_mem_reg[26][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][5]  ( .D(\Inst_Mem/inst_mem_reg[26][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[837]), .Q(
        \Inst_Mem/inst_mem_reg[26][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][6]  ( .D(\Inst_Mem/inst_mem_reg[26][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[838]), .Q(
        \Inst_Mem/inst_mem_reg[26][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][7]  ( .D(\Inst_Mem/inst_mem_reg[26][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[839]), .Q(
        \Inst_Mem/inst_mem_reg[26][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][8]  ( .D(\Inst_Mem/inst_mem_reg[26][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[840]), .Q(
        \Inst_Mem/inst_mem_reg[26][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][9]  ( .D(\Inst_Mem/inst_mem_reg[26][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[841]), .Q(
        \Inst_Mem/inst_mem_reg[26][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[26][10]  ( .D(\Inst_Mem/inst_mem_reg[26][10] ), .CLK(clk), .RST(rst), .I(g_init[842]), .Q(\Inst_Mem/inst_mem_reg[26][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][11]  ( .D(\Inst_Mem/inst_mem_reg[26][11] ), .CLK(clk), .RST(rst), .I(g_init[843]), .Q(\Inst_Mem/inst_mem_reg[26][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][12]  ( .D(\Inst_Mem/inst_mem_reg[26][12] ), .CLK(clk), .RST(rst), .I(g_init[844]), .Q(\Inst_Mem/inst_mem_reg[26][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][13]  ( .D(\Inst_Mem/inst_mem_reg[26][13] ), .CLK(clk), .RST(rst), .I(g_init[845]), .Q(\Inst_Mem/inst_mem_reg[26][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][14]  ( .D(\Inst_Mem/inst_mem_reg[26][14] ), .CLK(clk), .RST(rst), .I(g_init[846]), .Q(\Inst_Mem/inst_mem_reg[26][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][15]  ( .D(\Inst_Mem/inst_mem_reg[26][15] ), .CLK(clk), .RST(rst), .I(g_init[847]), .Q(\Inst_Mem/inst_mem_reg[26][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][16]  ( .D(\Inst_Mem/inst_mem_reg[26][16] ), .CLK(clk), .RST(rst), .I(g_init[848]), .Q(\Inst_Mem/inst_mem_reg[26][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][17]  ( .D(\Inst_Mem/inst_mem_reg[26][17] ), .CLK(clk), .RST(rst), .I(g_init[849]), .Q(\Inst_Mem/inst_mem_reg[26][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][18]  ( .D(\Inst_Mem/inst_mem_reg[26][18] ), .CLK(clk), .RST(rst), .I(g_init[850]), .Q(\Inst_Mem/inst_mem_reg[26][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][19]  ( .D(\Inst_Mem/inst_mem_reg[26][19] ), .CLK(clk), .RST(rst), .I(g_init[851]), .Q(\Inst_Mem/inst_mem_reg[26][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][20]  ( .D(\Inst_Mem/inst_mem_reg[26][20] ), .CLK(clk), .RST(rst), .I(g_init[852]), .Q(\Inst_Mem/inst_mem_reg[26][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][21]  ( .D(\Inst_Mem/inst_mem_reg[26][21] ), .CLK(clk), .RST(rst), .I(g_init[853]), .Q(\Inst_Mem/inst_mem_reg[26][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][22]  ( .D(\Inst_Mem/inst_mem_reg[26][22] ), .CLK(clk), .RST(rst), .I(g_init[854]), .Q(\Inst_Mem/inst_mem_reg[26][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][23]  ( .D(\Inst_Mem/inst_mem_reg[26][23] ), .CLK(clk), .RST(rst), .I(g_init[855]), .Q(\Inst_Mem/inst_mem_reg[26][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][24]  ( .D(\Inst_Mem/inst_mem_reg[26][24] ), .CLK(clk), .RST(rst), .I(g_init[856]), .Q(\Inst_Mem/inst_mem_reg[26][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][25]  ( .D(\Inst_Mem/inst_mem_reg[26][25] ), .CLK(clk), .RST(rst), .I(g_init[857]), .Q(\Inst_Mem/inst_mem_reg[26][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][26]  ( .D(\Inst_Mem/inst_mem_reg[26][26] ), .CLK(clk), .RST(rst), .I(g_init[858]), .Q(\Inst_Mem/inst_mem_reg[26][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][27]  ( .D(\Inst_Mem/inst_mem_reg[26][27] ), .CLK(clk), .RST(rst), .I(g_init[859]), .Q(\Inst_Mem/inst_mem_reg[26][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][28]  ( .D(\Inst_Mem/inst_mem_reg[26][28] ), .CLK(clk), .RST(rst), .I(g_init[860]), .Q(\Inst_Mem/inst_mem_reg[26][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][29]  ( .D(\Inst_Mem/inst_mem_reg[26][29] ), .CLK(clk), .RST(rst), .I(g_init[861]), .Q(\Inst_Mem/inst_mem_reg[26][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][30]  ( .D(\Inst_Mem/inst_mem_reg[26][30] ), .CLK(clk), .RST(rst), .I(g_init[862]), .Q(\Inst_Mem/inst_mem_reg[26][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[26][31]  ( .D(\Inst_Mem/inst_mem_reg[26][31] ), .CLK(clk), .RST(rst), .I(g_init[863]), .Q(\Inst_Mem/inst_mem_reg[26][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][0]  ( .D(\Inst_Mem/inst_mem_reg[25][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[800]), .Q(
        \Inst_Mem/inst_mem_reg[25][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][1]  ( .D(\Inst_Mem/inst_mem_reg[25][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[801]), .Q(
        \Inst_Mem/inst_mem_reg[25][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][2]  ( .D(\Inst_Mem/inst_mem_reg[25][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[802]), .Q(
        \Inst_Mem/inst_mem_reg[25][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][3]  ( .D(\Inst_Mem/inst_mem_reg[25][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[803]), .Q(
        \Inst_Mem/inst_mem_reg[25][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][4]  ( .D(\Inst_Mem/inst_mem_reg[25][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[804]), .Q(
        \Inst_Mem/inst_mem_reg[25][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][5]  ( .D(\Inst_Mem/inst_mem_reg[25][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[805]), .Q(
        \Inst_Mem/inst_mem_reg[25][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][6]  ( .D(\Inst_Mem/inst_mem_reg[25][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[806]), .Q(
        \Inst_Mem/inst_mem_reg[25][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][7]  ( .D(\Inst_Mem/inst_mem_reg[25][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[807]), .Q(
        \Inst_Mem/inst_mem_reg[25][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][8]  ( .D(\Inst_Mem/inst_mem_reg[25][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[808]), .Q(
        \Inst_Mem/inst_mem_reg[25][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][9]  ( .D(\Inst_Mem/inst_mem_reg[25][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[809]), .Q(
        \Inst_Mem/inst_mem_reg[25][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[25][10]  ( .D(\Inst_Mem/inst_mem_reg[25][10] ), .CLK(clk), .RST(rst), .I(g_init[810]), .Q(\Inst_Mem/inst_mem_reg[25][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][11]  ( .D(\Inst_Mem/inst_mem_reg[25][11] ), .CLK(clk), .RST(rst), .I(g_init[811]), .Q(\Inst_Mem/inst_mem_reg[25][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][12]  ( .D(\Inst_Mem/inst_mem_reg[25][12] ), .CLK(clk), .RST(rst), .I(g_init[812]), .Q(\Inst_Mem/inst_mem_reg[25][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][13]  ( .D(\Inst_Mem/inst_mem_reg[25][13] ), .CLK(clk), .RST(rst), .I(g_init[813]), .Q(\Inst_Mem/inst_mem_reg[25][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][14]  ( .D(\Inst_Mem/inst_mem_reg[25][14] ), .CLK(clk), .RST(rst), .I(g_init[814]), .Q(\Inst_Mem/inst_mem_reg[25][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][15]  ( .D(\Inst_Mem/inst_mem_reg[25][15] ), .CLK(clk), .RST(rst), .I(g_init[815]), .Q(\Inst_Mem/inst_mem_reg[25][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][16]  ( .D(\Inst_Mem/inst_mem_reg[25][16] ), .CLK(clk), .RST(rst), .I(g_init[816]), .Q(\Inst_Mem/inst_mem_reg[25][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][17]  ( .D(\Inst_Mem/inst_mem_reg[25][17] ), .CLK(clk), .RST(rst), .I(g_init[817]), .Q(\Inst_Mem/inst_mem_reg[25][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][18]  ( .D(\Inst_Mem/inst_mem_reg[25][18] ), .CLK(clk), .RST(rst), .I(g_init[818]), .Q(\Inst_Mem/inst_mem_reg[25][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][19]  ( .D(\Inst_Mem/inst_mem_reg[25][19] ), .CLK(clk), .RST(rst), .I(g_init[819]), .Q(\Inst_Mem/inst_mem_reg[25][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][20]  ( .D(\Inst_Mem/inst_mem_reg[25][20] ), .CLK(clk), .RST(rst), .I(g_init[820]), .Q(\Inst_Mem/inst_mem_reg[25][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][21]  ( .D(\Inst_Mem/inst_mem_reg[25][21] ), .CLK(clk), .RST(rst), .I(g_init[821]), .Q(\Inst_Mem/inst_mem_reg[25][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][22]  ( .D(\Inst_Mem/inst_mem_reg[25][22] ), .CLK(clk), .RST(rst), .I(g_init[822]), .Q(\Inst_Mem/inst_mem_reg[25][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][23]  ( .D(\Inst_Mem/inst_mem_reg[25][23] ), .CLK(clk), .RST(rst), .I(g_init[823]), .Q(\Inst_Mem/inst_mem_reg[25][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][24]  ( .D(\Inst_Mem/inst_mem_reg[25][24] ), .CLK(clk), .RST(rst), .I(g_init[824]), .Q(\Inst_Mem/inst_mem_reg[25][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][25]  ( .D(\Inst_Mem/inst_mem_reg[25][25] ), .CLK(clk), .RST(rst), .I(g_init[825]), .Q(\Inst_Mem/inst_mem_reg[25][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][26]  ( .D(\Inst_Mem/inst_mem_reg[25][26] ), .CLK(clk), .RST(rst), .I(g_init[826]), .Q(\Inst_Mem/inst_mem_reg[25][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][27]  ( .D(\Inst_Mem/inst_mem_reg[25][27] ), .CLK(clk), .RST(rst), .I(g_init[827]), .Q(\Inst_Mem/inst_mem_reg[25][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][28]  ( .D(\Inst_Mem/inst_mem_reg[25][28] ), .CLK(clk), .RST(rst), .I(g_init[828]), .Q(\Inst_Mem/inst_mem_reg[25][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][29]  ( .D(\Inst_Mem/inst_mem_reg[25][29] ), .CLK(clk), .RST(rst), .I(g_init[829]), .Q(\Inst_Mem/inst_mem_reg[25][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][30]  ( .D(\Inst_Mem/inst_mem_reg[25][30] ), .CLK(clk), .RST(rst), .I(g_init[830]), .Q(\Inst_Mem/inst_mem_reg[25][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[25][31]  ( .D(\Inst_Mem/inst_mem_reg[25][31] ), .CLK(clk), .RST(rst), .I(g_init[831]), .Q(\Inst_Mem/inst_mem_reg[25][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][0]  ( .D(\Inst_Mem/inst_mem_reg[24][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[768]), .Q(
        \Inst_Mem/inst_mem_reg[24][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][1]  ( .D(\Inst_Mem/inst_mem_reg[24][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[769]), .Q(
        \Inst_Mem/inst_mem_reg[24][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][2]  ( .D(\Inst_Mem/inst_mem_reg[24][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[770]), .Q(
        \Inst_Mem/inst_mem_reg[24][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][3]  ( .D(\Inst_Mem/inst_mem_reg[24][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[771]), .Q(
        \Inst_Mem/inst_mem_reg[24][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][4]  ( .D(\Inst_Mem/inst_mem_reg[24][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[772]), .Q(
        \Inst_Mem/inst_mem_reg[24][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][5]  ( .D(\Inst_Mem/inst_mem_reg[24][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[773]), .Q(
        \Inst_Mem/inst_mem_reg[24][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][6]  ( .D(\Inst_Mem/inst_mem_reg[24][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[774]), .Q(
        \Inst_Mem/inst_mem_reg[24][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][7]  ( .D(\Inst_Mem/inst_mem_reg[24][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[775]), .Q(
        \Inst_Mem/inst_mem_reg[24][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][8]  ( .D(\Inst_Mem/inst_mem_reg[24][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[776]), .Q(
        \Inst_Mem/inst_mem_reg[24][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][9]  ( .D(\Inst_Mem/inst_mem_reg[24][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[777]), .Q(
        \Inst_Mem/inst_mem_reg[24][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[24][10]  ( .D(\Inst_Mem/inst_mem_reg[24][10] ), .CLK(clk), .RST(rst), .I(g_init[778]), .Q(\Inst_Mem/inst_mem_reg[24][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][11]  ( .D(\Inst_Mem/inst_mem_reg[24][11] ), .CLK(clk), .RST(rst), .I(g_init[779]), .Q(\Inst_Mem/inst_mem_reg[24][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][12]  ( .D(\Inst_Mem/inst_mem_reg[24][12] ), .CLK(clk), .RST(rst), .I(g_init[780]), .Q(\Inst_Mem/inst_mem_reg[24][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][13]  ( .D(\Inst_Mem/inst_mem_reg[24][13] ), .CLK(clk), .RST(rst), .I(g_init[781]), .Q(\Inst_Mem/inst_mem_reg[24][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][14]  ( .D(\Inst_Mem/inst_mem_reg[24][14] ), .CLK(clk), .RST(rst), .I(g_init[782]), .Q(\Inst_Mem/inst_mem_reg[24][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][15]  ( .D(\Inst_Mem/inst_mem_reg[24][15] ), .CLK(clk), .RST(rst), .I(g_init[783]), .Q(\Inst_Mem/inst_mem_reg[24][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][16]  ( .D(\Inst_Mem/inst_mem_reg[24][16] ), .CLK(clk), .RST(rst), .I(g_init[784]), .Q(\Inst_Mem/inst_mem_reg[24][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][17]  ( .D(\Inst_Mem/inst_mem_reg[24][17] ), .CLK(clk), .RST(rst), .I(g_init[785]), .Q(\Inst_Mem/inst_mem_reg[24][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][18]  ( .D(\Inst_Mem/inst_mem_reg[24][18] ), .CLK(clk), .RST(rst), .I(g_init[786]), .Q(\Inst_Mem/inst_mem_reg[24][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][19]  ( .D(\Inst_Mem/inst_mem_reg[24][19] ), .CLK(clk), .RST(rst), .I(g_init[787]), .Q(\Inst_Mem/inst_mem_reg[24][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][20]  ( .D(\Inst_Mem/inst_mem_reg[24][20] ), .CLK(clk), .RST(rst), .I(g_init[788]), .Q(\Inst_Mem/inst_mem_reg[24][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][21]  ( .D(\Inst_Mem/inst_mem_reg[24][21] ), .CLK(clk), .RST(rst), .I(g_init[789]), .Q(\Inst_Mem/inst_mem_reg[24][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][22]  ( .D(\Inst_Mem/inst_mem_reg[24][22] ), .CLK(clk), .RST(rst), .I(g_init[790]), .Q(\Inst_Mem/inst_mem_reg[24][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][23]  ( .D(\Inst_Mem/inst_mem_reg[24][23] ), .CLK(clk), .RST(rst), .I(g_init[791]), .Q(\Inst_Mem/inst_mem_reg[24][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][24]  ( .D(\Inst_Mem/inst_mem_reg[24][24] ), .CLK(clk), .RST(rst), .I(g_init[792]), .Q(\Inst_Mem/inst_mem_reg[24][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][25]  ( .D(\Inst_Mem/inst_mem_reg[24][25] ), .CLK(clk), .RST(rst), .I(g_init[793]), .Q(\Inst_Mem/inst_mem_reg[24][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][26]  ( .D(\Inst_Mem/inst_mem_reg[24][26] ), .CLK(clk), .RST(rst), .I(g_init[794]), .Q(\Inst_Mem/inst_mem_reg[24][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][27]  ( .D(\Inst_Mem/inst_mem_reg[24][27] ), .CLK(clk), .RST(rst), .I(g_init[795]), .Q(\Inst_Mem/inst_mem_reg[24][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][28]  ( .D(\Inst_Mem/inst_mem_reg[24][28] ), .CLK(clk), .RST(rst), .I(g_init[796]), .Q(\Inst_Mem/inst_mem_reg[24][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][29]  ( .D(\Inst_Mem/inst_mem_reg[24][29] ), .CLK(clk), .RST(rst), .I(g_init[797]), .Q(\Inst_Mem/inst_mem_reg[24][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][30]  ( .D(\Inst_Mem/inst_mem_reg[24][30] ), .CLK(clk), .RST(rst), .I(g_init[798]), .Q(\Inst_Mem/inst_mem_reg[24][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[24][31]  ( .D(\Inst_Mem/inst_mem_reg[24][31] ), .CLK(clk), .RST(rst), .I(g_init[799]), .Q(\Inst_Mem/inst_mem_reg[24][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][0]  ( .D(\Inst_Mem/inst_mem_reg[23][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[736]), .Q(
        \Inst_Mem/inst_mem_reg[23][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][1]  ( .D(\Inst_Mem/inst_mem_reg[23][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[737]), .Q(
        \Inst_Mem/inst_mem_reg[23][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][2]  ( .D(\Inst_Mem/inst_mem_reg[23][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[738]), .Q(
        \Inst_Mem/inst_mem_reg[23][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][3]  ( .D(\Inst_Mem/inst_mem_reg[23][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[739]), .Q(
        \Inst_Mem/inst_mem_reg[23][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][4]  ( .D(\Inst_Mem/inst_mem_reg[23][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[740]), .Q(
        \Inst_Mem/inst_mem_reg[23][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][5]  ( .D(\Inst_Mem/inst_mem_reg[23][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[741]), .Q(
        \Inst_Mem/inst_mem_reg[23][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][6]  ( .D(\Inst_Mem/inst_mem_reg[23][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[742]), .Q(
        \Inst_Mem/inst_mem_reg[23][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][7]  ( .D(\Inst_Mem/inst_mem_reg[23][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[743]), .Q(
        \Inst_Mem/inst_mem_reg[23][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][8]  ( .D(\Inst_Mem/inst_mem_reg[23][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[744]), .Q(
        \Inst_Mem/inst_mem_reg[23][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][9]  ( .D(\Inst_Mem/inst_mem_reg[23][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[745]), .Q(
        \Inst_Mem/inst_mem_reg[23][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[23][10]  ( .D(\Inst_Mem/inst_mem_reg[23][10] ), .CLK(clk), .RST(rst), .I(g_init[746]), .Q(\Inst_Mem/inst_mem_reg[23][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][11]  ( .D(\Inst_Mem/inst_mem_reg[23][11] ), .CLK(clk), .RST(rst), .I(g_init[747]), .Q(\Inst_Mem/inst_mem_reg[23][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][12]  ( .D(\Inst_Mem/inst_mem_reg[23][12] ), .CLK(clk), .RST(rst), .I(g_init[748]), .Q(\Inst_Mem/inst_mem_reg[23][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][13]  ( .D(\Inst_Mem/inst_mem_reg[23][13] ), .CLK(clk), .RST(rst), .I(g_init[749]), .Q(\Inst_Mem/inst_mem_reg[23][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][14]  ( .D(\Inst_Mem/inst_mem_reg[23][14] ), .CLK(clk), .RST(rst), .I(g_init[750]), .Q(\Inst_Mem/inst_mem_reg[23][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][15]  ( .D(\Inst_Mem/inst_mem_reg[23][15] ), .CLK(clk), .RST(rst), .I(g_init[751]), .Q(\Inst_Mem/inst_mem_reg[23][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][16]  ( .D(\Inst_Mem/inst_mem_reg[23][16] ), .CLK(clk), .RST(rst), .I(g_init[752]), .Q(\Inst_Mem/inst_mem_reg[23][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][17]  ( .D(\Inst_Mem/inst_mem_reg[23][17] ), .CLK(clk), .RST(rst), .I(g_init[753]), .Q(\Inst_Mem/inst_mem_reg[23][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][18]  ( .D(\Inst_Mem/inst_mem_reg[23][18] ), .CLK(clk), .RST(rst), .I(g_init[754]), .Q(\Inst_Mem/inst_mem_reg[23][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][19]  ( .D(\Inst_Mem/inst_mem_reg[23][19] ), .CLK(clk), .RST(rst), .I(g_init[755]), .Q(\Inst_Mem/inst_mem_reg[23][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][20]  ( .D(\Inst_Mem/inst_mem_reg[23][20] ), .CLK(clk), .RST(rst), .I(g_init[756]), .Q(\Inst_Mem/inst_mem_reg[23][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][21]  ( .D(\Inst_Mem/inst_mem_reg[23][21] ), .CLK(clk), .RST(rst), .I(g_init[757]), .Q(\Inst_Mem/inst_mem_reg[23][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][22]  ( .D(\Inst_Mem/inst_mem_reg[23][22] ), .CLK(clk), .RST(rst), .I(g_init[758]), .Q(\Inst_Mem/inst_mem_reg[23][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][23]  ( .D(\Inst_Mem/inst_mem_reg[23][23] ), .CLK(clk), .RST(rst), .I(g_init[759]), .Q(\Inst_Mem/inst_mem_reg[23][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][24]  ( .D(\Inst_Mem/inst_mem_reg[23][24] ), .CLK(clk), .RST(rst), .I(g_init[760]), .Q(\Inst_Mem/inst_mem_reg[23][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][25]  ( .D(\Inst_Mem/inst_mem_reg[23][25] ), .CLK(clk), .RST(rst), .I(g_init[761]), .Q(\Inst_Mem/inst_mem_reg[23][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][26]  ( .D(\Inst_Mem/inst_mem_reg[23][26] ), .CLK(clk), .RST(rst), .I(g_init[762]), .Q(\Inst_Mem/inst_mem_reg[23][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][27]  ( .D(\Inst_Mem/inst_mem_reg[23][27] ), .CLK(clk), .RST(rst), .I(g_init[763]), .Q(\Inst_Mem/inst_mem_reg[23][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][28]  ( .D(\Inst_Mem/inst_mem_reg[23][28] ), .CLK(clk), .RST(rst), .I(g_init[764]), .Q(\Inst_Mem/inst_mem_reg[23][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][29]  ( .D(\Inst_Mem/inst_mem_reg[23][29] ), .CLK(clk), .RST(rst), .I(g_init[765]), .Q(\Inst_Mem/inst_mem_reg[23][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][30]  ( .D(\Inst_Mem/inst_mem_reg[23][30] ), .CLK(clk), .RST(rst), .I(g_init[766]), .Q(\Inst_Mem/inst_mem_reg[23][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[23][31]  ( .D(\Inst_Mem/inst_mem_reg[23][31] ), .CLK(clk), .RST(rst), .I(g_init[767]), .Q(\Inst_Mem/inst_mem_reg[23][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][0]  ( .D(\Inst_Mem/inst_mem_reg[22][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[704]), .Q(
        \Inst_Mem/inst_mem_reg[22][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][1]  ( .D(\Inst_Mem/inst_mem_reg[22][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[705]), .Q(
        \Inst_Mem/inst_mem_reg[22][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][2]  ( .D(\Inst_Mem/inst_mem_reg[22][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[706]), .Q(
        \Inst_Mem/inst_mem_reg[22][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][3]  ( .D(\Inst_Mem/inst_mem_reg[22][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[707]), .Q(
        \Inst_Mem/inst_mem_reg[22][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][4]  ( .D(\Inst_Mem/inst_mem_reg[22][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[708]), .Q(
        \Inst_Mem/inst_mem_reg[22][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][5]  ( .D(\Inst_Mem/inst_mem_reg[22][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[709]), .Q(
        \Inst_Mem/inst_mem_reg[22][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][6]  ( .D(\Inst_Mem/inst_mem_reg[22][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[710]), .Q(
        \Inst_Mem/inst_mem_reg[22][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][7]  ( .D(\Inst_Mem/inst_mem_reg[22][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[711]), .Q(
        \Inst_Mem/inst_mem_reg[22][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][8]  ( .D(\Inst_Mem/inst_mem_reg[22][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[712]), .Q(
        \Inst_Mem/inst_mem_reg[22][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][9]  ( .D(\Inst_Mem/inst_mem_reg[22][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[713]), .Q(
        \Inst_Mem/inst_mem_reg[22][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[22][10]  ( .D(\Inst_Mem/inst_mem_reg[22][10] ), .CLK(clk), .RST(rst), .I(g_init[714]), .Q(\Inst_Mem/inst_mem_reg[22][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][11]  ( .D(\Inst_Mem/inst_mem_reg[22][11] ), .CLK(clk), .RST(rst), .I(g_init[715]), .Q(\Inst_Mem/inst_mem_reg[22][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][12]  ( .D(\Inst_Mem/inst_mem_reg[22][12] ), .CLK(clk), .RST(rst), .I(g_init[716]), .Q(\Inst_Mem/inst_mem_reg[22][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][13]  ( .D(\Inst_Mem/inst_mem_reg[22][13] ), .CLK(clk), .RST(rst), .I(g_init[717]), .Q(\Inst_Mem/inst_mem_reg[22][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][14]  ( .D(\Inst_Mem/inst_mem_reg[22][14] ), .CLK(clk), .RST(rst), .I(g_init[718]), .Q(\Inst_Mem/inst_mem_reg[22][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][15]  ( .D(\Inst_Mem/inst_mem_reg[22][15] ), .CLK(clk), .RST(rst), .I(g_init[719]), .Q(\Inst_Mem/inst_mem_reg[22][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][16]  ( .D(\Inst_Mem/inst_mem_reg[22][16] ), .CLK(clk), .RST(rst), .I(g_init[720]), .Q(\Inst_Mem/inst_mem_reg[22][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][17]  ( .D(\Inst_Mem/inst_mem_reg[22][17] ), .CLK(clk), .RST(rst), .I(g_init[721]), .Q(\Inst_Mem/inst_mem_reg[22][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][18]  ( .D(\Inst_Mem/inst_mem_reg[22][18] ), .CLK(clk), .RST(rst), .I(g_init[722]), .Q(\Inst_Mem/inst_mem_reg[22][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][19]  ( .D(\Inst_Mem/inst_mem_reg[22][19] ), .CLK(clk), .RST(rst), .I(g_init[723]), .Q(\Inst_Mem/inst_mem_reg[22][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][20]  ( .D(\Inst_Mem/inst_mem_reg[22][20] ), .CLK(clk), .RST(rst), .I(g_init[724]), .Q(\Inst_Mem/inst_mem_reg[22][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][21]  ( .D(\Inst_Mem/inst_mem_reg[22][21] ), .CLK(clk), .RST(rst), .I(g_init[725]), .Q(\Inst_Mem/inst_mem_reg[22][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][22]  ( .D(\Inst_Mem/inst_mem_reg[22][22] ), .CLK(clk), .RST(rst), .I(g_init[726]), .Q(\Inst_Mem/inst_mem_reg[22][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][23]  ( .D(\Inst_Mem/inst_mem_reg[22][23] ), .CLK(clk), .RST(rst), .I(g_init[727]), .Q(\Inst_Mem/inst_mem_reg[22][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][24]  ( .D(\Inst_Mem/inst_mem_reg[22][24] ), .CLK(clk), .RST(rst), .I(g_init[728]), .Q(\Inst_Mem/inst_mem_reg[22][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][25]  ( .D(\Inst_Mem/inst_mem_reg[22][25] ), .CLK(clk), .RST(rst), .I(g_init[729]), .Q(\Inst_Mem/inst_mem_reg[22][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][26]  ( .D(\Inst_Mem/inst_mem_reg[22][26] ), .CLK(clk), .RST(rst), .I(g_init[730]), .Q(\Inst_Mem/inst_mem_reg[22][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][27]  ( .D(\Inst_Mem/inst_mem_reg[22][27] ), .CLK(clk), .RST(rst), .I(g_init[731]), .Q(\Inst_Mem/inst_mem_reg[22][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][28]  ( .D(\Inst_Mem/inst_mem_reg[22][28] ), .CLK(clk), .RST(rst), .I(g_init[732]), .Q(\Inst_Mem/inst_mem_reg[22][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][29]  ( .D(\Inst_Mem/inst_mem_reg[22][29] ), .CLK(clk), .RST(rst), .I(g_init[733]), .Q(\Inst_Mem/inst_mem_reg[22][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][30]  ( .D(\Inst_Mem/inst_mem_reg[22][30] ), .CLK(clk), .RST(rst), .I(g_init[734]), .Q(\Inst_Mem/inst_mem_reg[22][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[22][31]  ( .D(\Inst_Mem/inst_mem_reg[22][31] ), .CLK(clk), .RST(rst), .I(g_init[735]), .Q(\Inst_Mem/inst_mem_reg[22][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][0]  ( .D(\Inst_Mem/inst_mem_reg[21][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[672]), .Q(
        \Inst_Mem/inst_mem_reg[21][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][1]  ( .D(\Inst_Mem/inst_mem_reg[21][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[673]), .Q(
        \Inst_Mem/inst_mem_reg[21][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][2]  ( .D(\Inst_Mem/inst_mem_reg[21][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[674]), .Q(
        \Inst_Mem/inst_mem_reg[21][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][3]  ( .D(\Inst_Mem/inst_mem_reg[21][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[675]), .Q(
        \Inst_Mem/inst_mem_reg[21][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][4]  ( .D(\Inst_Mem/inst_mem_reg[21][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[676]), .Q(
        \Inst_Mem/inst_mem_reg[21][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][5]  ( .D(\Inst_Mem/inst_mem_reg[21][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[677]), .Q(
        \Inst_Mem/inst_mem_reg[21][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][6]  ( .D(\Inst_Mem/inst_mem_reg[21][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[678]), .Q(
        \Inst_Mem/inst_mem_reg[21][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][7]  ( .D(\Inst_Mem/inst_mem_reg[21][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[679]), .Q(
        \Inst_Mem/inst_mem_reg[21][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][8]  ( .D(\Inst_Mem/inst_mem_reg[21][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[680]), .Q(
        \Inst_Mem/inst_mem_reg[21][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][9]  ( .D(\Inst_Mem/inst_mem_reg[21][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[681]), .Q(
        \Inst_Mem/inst_mem_reg[21][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[21][10]  ( .D(\Inst_Mem/inst_mem_reg[21][10] ), .CLK(clk), .RST(rst), .I(g_init[682]), .Q(\Inst_Mem/inst_mem_reg[21][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][11]  ( .D(\Inst_Mem/inst_mem_reg[21][11] ), .CLK(clk), .RST(rst), .I(g_init[683]), .Q(\Inst_Mem/inst_mem_reg[21][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][12]  ( .D(\Inst_Mem/inst_mem_reg[21][12] ), .CLK(clk), .RST(rst), .I(g_init[684]), .Q(\Inst_Mem/inst_mem_reg[21][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][13]  ( .D(\Inst_Mem/inst_mem_reg[21][13] ), .CLK(clk), .RST(rst), .I(g_init[685]), .Q(\Inst_Mem/inst_mem_reg[21][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][14]  ( .D(\Inst_Mem/inst_mem_reg[21][14] ), .CLK(clk), .RST(rst), .I(g_init[686]), .Q(\Inst_Mem/inst_mem_reg[21][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][15]  ( .D(\Inst_Mem/inst_mem_reg[21][15] ), .CLK(clk), .RST(rst), .I(g_init[687]), .Q(\Inst_Mem/inst_mem_reg[21][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][16]  ( .D(\Inst_Mem/inst_mem_reg[21][16] ), .CLK(clk), .RST(rst), .I(g_init[688]), .Q(\Inst_Mem/inst_mem_reg[21][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][17]  ( .D(\Inst_Mem/inst_mem_reg[21][17] ), .CLK(clk), .RST(rst), .I(g_init[689]), .Q(\Inst_Mem/inst_mem_reg[21][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][18]  ( .D(\Inst_Mem/inst_mem_reg[21][18] ), .CLK(clk), .RST(rst), .I(g_init[690]), .Q(\Inst_Mem/inst_mem_reg[21][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][19]  ( .D(\Inst_Mem/inst_mem_reg[21][19] ), .CLK(clk), .RST(rst), .I(g_init[691]), .Q(\Inst_Mem/inst_mem_reg[21][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][20]  ( .D(\Inst_Mem/inst_mem_reg[21][20] ), .CLK(clk), .RST(rst), .I(g_init[692]), .Q(\Inst_Mem/inst_mem_reg[21][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][21]  ( .D(\Inst_Mem/inst_mem_reg[21][21] ), .CLK(clk), .RST(rst), .I(g_init[693]), .Q(\Inst_Mem/inst_mem_reg[21][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][22]  ( .D(\Inst_Mem/inst_mem_reg[21][22] ), .CLK(clk), .RST(rst), .I(g_init[694]), .Q(\Inst_Mem/inst_mem_reg[21][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][23]  ( .D(\Inst_Mem/inst_mem_reg[21][23] ), .CLK(clk), .RST(rst), .I(g_init[695]), .Q(\Inst_Mem/inst_mem_reg[21][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][24]  ( .D(\Inst_Mem/inst_mem_reg[21][24] ), .CLK(clk), .RST(rst), .I(g_init[696]), .Q(\Inst_Mem/inst_mem_reg[21][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][25]  ( .D(\Inst_Mem/inst_mem_reg[21][25] ), .CLK(clk), .RST(rst), .I(g_init[697]), .Q(\Inst_Mem/inst_mem_reg[21][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][26]  ( .D(\Inst_Mem/inst_mem_reg[21][26] ), .CLK(clk), .RST(rst), .I(g_init[698]), .Q(\Inst_Mem/inst_mem_reg[21][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][27]  ( .D(\Inst_Mem/inst_mem_reg[21][27] ), .CLK(clk), .RST(rst), .I(g_init[699]), .Q(\Inst_Mem/inst_mem_reg[21][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][28]  ( .D(\Inst_Mem/inst_mem_reg[21][28] ), .CLK(clk), .RST(rst), .I(g_init[700]), .Q(\Inst_Mem/inst_mem_reg[21][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][29]  ( .D(\Inst_Mem/inst_mem_reg[21][29] ), .CLK(clk), .RST(rst), .I(g_init[701]), .Q(\Inst_Mem/inst_mem_reg[21][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][30]  ( .D(\Inst_Mem/inst_mem_reg[21][30] ), .CLK(clk), .RST(rst), .I(g_init[702]), .Q(\Inst_Mem/inst_mem_reg[21][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[21][31]  ( .D(\Inst_Mem/inst_mem_reg[21][31] ), .CLK(clk), .RST(rst), .I(g_init[703]), .Q(\Inst_Mem/inst_mem_reg[21][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][0]  ( .D(\Inst_Mem/inst_mem_reg[20][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[640]), .Q(
        \Inst_Mem/inst_mem_reg[20][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][1]  ( .D(\Inst_Mem/inst_mem_reg[20][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[641]), .Q(
        \Inst_Mem/inst_mem_reg[20][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][2]  ( .D(\Inst_Mem/inst_mem_reg[20][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[642]), .Q(
        \Inst_Mem/inst_mem_reg[20][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][3]  ( .D(\Inst_Mem/inst_mem_reg[20][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[643]), .Q(
        \Inst_Mem/inst_mem_reg[20][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][4]  ( .D(\Inst_Mem/inst_mem_reg[20][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[644]), .Q(
        \Inst_Mem/inst_mem_reg[20][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][5]  ( .D(\Inst_Mem/inst_mem_reg[20][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[645]), .Q(
        \Inst_Mem/inst_mem_reg[20][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][6]  ( .D(\Inst_Mem/inst_mem_reg[20][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[646]), .Q(
        \Inst_Mem/inst_mem_reg[20][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][7]  ( .D(\Inst_Mem/inst_mem_reg[20][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[647]), .Q(
        \Inst_Mem/inst_mem_reg[20][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][8]  ( .D(\Inst_Mem/inst_mem_reg[20][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[648]), .Q(
        \Inst_Mem/inst_mem_reg[20][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][9]  ( .D(\Inst_Mem/inst_mem_reg[20][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[649]), .Q(
        \Inst_Mem/inst_mem_reg[20][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[20][10]  ( .D(\Inst_Mem/inst_mem_reg[20][10] ), .CLK(clk), .RST(rst), .I(g_init[650]), .Q(\Inst_Mem/inst_mem_reg[20][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][11]  ( .D(\Inst_Mem/inst_mem_reg[20][11] ), .CLK(clk), .RST(rst), .I(g_init[651]), .Q(\Inst_Mem/inst_mem_reg[20][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][12]  ( .D(\Inst_Mem/inst_mem_reg[20][12] ), .CLK(clk), .RST(rst), .I(g_init[652]), .Q(\Inst_Mem/inst_mem_reg[20][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][13]  ( .D(\Inst_Mem/inst_mem_reg[20][13] ), .CLK(clk), .RST(rst), .I(g_init[653]), .Q(\Inst_Mem/inst_mem_reg[20][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][14]  ( .D(\Inst_Mem/inst_mem_reg[20][14] ), .CLK(clk), .RST(rst), .I(g_init[654]), .Q(\Inst_Mem/inst_mem_reg[20][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][15]  ( .D(\Inst_Mem/inst_mem_reg[20][15] ), .CLK(clk), .RST(rst), .I(g_init[655]), .Q(\Inst_Mem/inst_mem_reg[20][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][16]  ( .D(\Inst_Mem/inst_mem_reg[20][16] ), .CLK(clk), .RST(rst), .I(g_init[656]), .Q(\Inst_Mem/inst_mem_reg[20][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][17]  ( .D(\Inst_Mem/inst_mem_reg[20][17] ), .CLK(clk), .RST(rst), .I(g_init[657]), .Q(\Inst_Mem/inst_mem_reg[20][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][18]  ( .D(\Inst_Mem/inst_mem_reg[20][18] ), .CLK(clk), .RST(rst), .I(g_init[658]), .Q(\Inst_Mem/inst_mem_reg[20][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][19]  ( .D(\Inst_Mem/inst_mem_reg[20][19] ), .CLK(clk), .RST(rst), .I(g_init[659]), .Q(\Inst_Mem/inst_mem_reg[20][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][20]  ( .D(\Inst_Mem/inst_mem_reg[20][20] ), .CLK(clk), .RST(rst), .I(g_init[660]), .Q(\Inst_Mem/inst_mem_reg[20][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][21]  ( .D(\Inst_Mem/inst_mem_reg[20][21] ), .CLK(clk), .RST(rst), .I(g_init[661]), .Q(\Inst_Mem/inst_mem_reg[20][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][22]  ( .D(\Inst_Mem/inst_mem_reg[20][22] ), .CLK(clk), .RST(rst), .I(g_init[662]), .Q(\Inst_Mem/inst_mem_reg[20][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][23]  ( .D(\Inst_Mem/inst_mem_reg[20][23] ), .CLK(clk), .RST(rst), .I(g_init[663]), .Q(\Inst_Mem/inst_mem_reg[20][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][24]  ( .D(\Inst_Mem/inst_mem_reg[20][24] ), .CLK(clk), .RST(rst), .I(g_init[664]), .Q(\Inst_Mem/inst_mem_reg[20][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][25]  ( .D(\Inst_Mem/inst_mem_reg[20][25] ), .CLK(clk), .RST(rst), .I(g_init[665]), .Q(\Inst_Mem/inst_mem_reg[20][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][26]  ( .D(\Inst_Mem/inst_mem_reg[20][26] ), .CLK(clk), .RST(rst), .I(g_init[666]), .Q(\Inst_Mem/inst_mem_reg[20][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][27]  ( .D(\Inst_Mem/inst_mem_reg[20][27] ), .CLK(clk), .RST(rst), .I(g_init[667]), .Q(\Inst_Mem/inst_mem_reg[20][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][28]  ( .D(\Inst_Mem/inst_mem_reg[20][28] ), .CLK(clk), .RST(rst), .I(g_init[668]), .Q(\Inst_Mem/inst_mem_reg[20][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][29]  ( .D(\Inst_Mem/inst_mem_reg[20][29] ), .CLK(clk), .RST(rst), .I(g_init[669]), .Q(\Inst_Mem/inst_mem_reg[20][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][30]  ( .D(\Inst_Mem/inst_mem_reg[20][30] ), .CLK(clk), .RST(rst), .I(g_init[670]), .Q(\Inst_Mem/inst_mem_reg[20][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[20][31]  ( .D(\Inst_Mem/inst_mem_reg[20][31] ), .CLK(clk), .RST(rst), .I(g_init[671]), .Q(\Inst_Mem/inst_mem_reg[20][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][0]  ( .D(\Inst_Mem/inst_mem_reg[19][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[608]), .Q(
        \Inst_Mem/inst_mem_reg[19][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][1]  ( .D(\Inst_Mem/inst_mem_reg[19][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[609]), .Q(
        \Inst_Mem/inst_mem_reg[19][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][2]  ( .D(\Inst_Mem/inst_mem_reg[19][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[610]), .Q(
        \Inst_Mem/inst_mem_reg[19][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][3]  ( .D(\Inst_Mem/inst_mem_reg[19][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[611]), .Q(
        \Inst_Mem/inst_mem_reg[19][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][4]  ( .D(\Inst_Mem/inst_mem_reg[19][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[612]), .Q(
        \Inst_Mem/inst_mem_reg[19][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][5]  ( .D(\Inst_Mem/inst_mem_reg[19][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[613]), .Q(
        \Inst_Mem/inst_mem_reg[19][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][6]  ( .D(\Inst_Mem/inst_mem_reg[19][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[614]), .Q(
        \Inst_Mem/inst_mem_reg[19][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][7]  ( .D(\Inst_Mem/inst_mem_reg[19][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[615]), .Q(
        \Inst_Mem/inst_mem_reg[19][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][8]  ( .D(\Inst_Mem/inst_mem_reg[19][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[616]), .Q(
        \Inst_Mem/inst_mem_reg[19][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][9]  ( .D(\Inst_Mem/inst_mem_reg[19][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[617]), .Q(
        \Inst_Mem/inst_mem_reg[19][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[19][10]  ( .D(\Inst_Mem/inst_mem_reg[19][10] ), .CLK(clk), .RST(rst), .I(g_init[618]), .Q(\Inst_Mem/inst_mem_reg[19][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][11]  ( .D(\Inst_Mem/inst_mem_reg[19][11] ), .CLK(clk), .RST(rst), .I(g_init[619]), .Q(\Inst_Mem/inst_mem_reg[19][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][12]  ( .D(\Inst_Mem/inst_mem_reg[19][12] ), .CLK(clk), .RST(rst), .I(g_init[620]), .Q(\Inst_Mem/inst_mem_reg[19][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][13]  ( .D(\Inst_Mem/inst_mem_reg[19][13] ), .CLK(clk), .RST(rst), .I(g_init[621]), .Q(\Inst_Mem/inst_mem_reg[19][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][14]  ( .D(\Inst_Mem/inst_mem_reg[19][14] ), .CLK(clk), .RST(rst), .I(g_init[622]), .Q(\Inst_Mem/inst_mem_reg[19][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][15]  ( .D(\Inst_Mem/inst_mem_reg[19][15] ), .CLK(clk), .RST(rst), .I(g_init[623]), .Q(\Inst_Mem/inst_mem_reg[19][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][16]  ( .D(\Inst_Mem/inst_mem_reg[19][16] ), .CLK(clk), .RST(rst), .I(g_init[624]), .Q(\Inst_Mem/inst_mem_reg[19][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][17]  ( .D(\Inst_Mem/inst_mem_reg[19][17] ), .CLK(clk), .RST(rst), .I(g_init[625]), .Q(\Inst_Mem/inst_mem_reg[19][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][18]  ( .D(\Inst_Mem/inst_mem_reg[19][18] ), .CLK(clk), .RST(rst), .I(g_init[626]), .Q(\Inst_Mem/inst_mem_reg[19][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][19]  ( .D(\Inst_Mem/inst_mem_reg[19][19] ), .CLK(clk), .RST(rst), .I(g_init[627]), .Q(\Inst_Mem/inst_mem_reg[19][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][20]  ( .D(\Inst_Mem/inst_mem_reg[19][20] ), .CLK(clk), .RST(rst), .I(g_init[628]), .Q(\Inst_Mem/inst_mem_reg[19][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][21]  ( .D(\Inst_Mem/inst_mem_reg[19][21] ), .CLK(clk), .RST(rst), .I(g_init[629]), .Q(\Inst_Mem/inst_mem_reg[19][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][22]  ( .D(\Inst_Mem/inst_mem_reg[19][22] ), .CLK(clk), .RST(rst), .I(g_init[630]), .Q(\Inst_Mem/inst_mem_reg[19][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][23]  ( .D(\Inst_Mem/inst_mem_reg[19][23] ), .CLK(clk), .RST(rst), .I(g_init[631]), .Q(\Inst_Mem/inst_mem_reg[19][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][24]  ( .D(\Inst_Mem/inst_mem_reg[19][24] ), .CLK(clk), .RST(rst), .I(g_init[632]), .Q(\Inst_Mem/inst_mem_reg[19][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][25]  ( .D(\Inst_Mem/inst_mem_reg[19][25] ), .CLK(clk), .RST(rst), .I(g_init[633]), .Q(\Inst_Mem/inst_mem_reg[19][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][26]  ( .D(\Inst_Mem/inst_mem_reg[19][26] ), .CLK(clk), .RST(rst), .I(g_init[634]), .Q(\Inst_Mem/inst_mem_reg[19][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][27]  ( .D(\Inst_Mem/inst_mem_reg[19][27] ), .CLK(clk), .RST(rst), .I(g_init[635]), .Q(\Inst_Mem/inst_mem_reg[19][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][28]  ( .D(\Inst_Mem/inst_mem_reg[19][28] ), .CLK(clk), .RST(rst), .I(g_init[636]), .Q(\Inst_Mem/inst_mem_reg[19][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][29]  ( .D(\Inst_Mem/inst_mem_reg[19][29] ), .CLK(clk), .RST(rst), .I(g_init[637]), .Q(\Inst_Mem/inst_mem_reg[19][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][30]  ( .D(\Inst_Mem/inst_mem_reg[19][30] ), .CLK(clk), .RST(rst), .I(g_init[638]), .Q(\Inst_Mem/inst_mem_reg[19][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[19][31]  ( .D(\Inst_Mem/inst_mem_reg[19][31] ), .CLK(clk), .RST(rst), .I(g_init[639]), .Q(\Inst_Mem/inst_mem_reg[19][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][0]  ( .D(\Inst_Mem/inst_mem_reg[18][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[576]), .Q(
        \Inst_Mem/inst_mem_reg[18][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][1]  ( .D(\Inst_Mem/inst_mem_reg[18][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[577]), .Q(
        \Inst_Mem/inst_mem_reg[18][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][2]  ( .D(\Inst_Mem/inst_mem_reg[18][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[578]), .Q(
        \Inst_Mem/inst_mem_reg[18][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][3]  ( .D(\Inst_Mem/inst_mem_reg[18][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[579]), .Q(
        \Inst_Mem/inst_mem_reg[18][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][4]  ( .D(\Inst_Mem/inst_mem_reg[18][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[580]), .Q(
        \Inst_Mem/inst_mem_reg[18][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][5]  ( .D(\Inst_Mem/inst_mem_reg[18][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[581]), .Q(
        \Inst_Mem/inst_mem_reg[18][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][6]  ( .D(\Inst_Mem/inst_mem_reg[18][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[582]), .Q(
        \Inst_Mem/inst_mem_reg[18][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][7]  ( .D(\Inst_Mem/inst_mem_reg[18][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[583]), .Q(
        \Inst_Mem/inst_mem_reg[18][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][8]  ( .D(\Inst_Mem/inst_mem_reg[18][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[584]), .Q(
        \Inst_Mem/inst_mem_reg[18][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][9]  ( .D(\Inst_Mem/inst_mem_reg[18][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[585]), .Q(
        \Inst_Mem/inst_mem_reg[18][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[18][10]  ( .D(\Inst_Mem/inst_mem_reg[18][10] ), .CLK(clk), .RST(rst), .I(g_init[586]), .Q(\Inst_Mem/inst_mem_reg[18][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][11]  ( .D(\Inst_Mem/inst_mem_reg[18][11] ), .CLK(clk), .RST(rst), .I(g_init[587]), .Q(\Inst_Mem/inst_mem_reg[18][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][12]  ( .D(\Inst_Mem/inst_mem_reg[18][12] ), .CLK(clk), .RST(rst), .I(g_init[588]), .Q(\Inst_Mem/inst_mem_reg[18][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][13]  ( .D(\Inst_Mem/inst_mem_reg[18][13] ), .CLK(clk), .RST(rst), .I(g_init[589]), .Q(\Inst_Mem/inst_mem_reg[18][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][14]  ( .D(\Inst_Mem/inst_mem_reg[18][14] ), .CLK(clk), .RST(rst), .I(g_init[590]), .Q(\Inst_Mem/inst_mem_reg[18][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][15]  ( .D(\Inst_Mem/inst_mem_reg[18][15] ), .CLK(clk), .RST(rst), .I(g_init[591]), .Q(\Inst_Mem/inst_mem_reg[18][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][16]  ( .D(\Inst_Mem/inst_mem_reg[18][16] ), .CLK(clk), .RST(rst), .I(g_init[592]), .Q(\Inst_Mem/inst_mem_reg[18][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][17]  ( .D(\Inst_Mem/inst_mem_reg[18][17] ), .CLK(clk), .RST(rst), .I(g_init[593]), .Q(\Inst_Mem/inst_mem_reg[18][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][18]  ( .D(\Inst_Mem/inst_mem_reg[18][18] ), .CLK(clk), .RST(rst), .I(g_init[594]), .Q(\Inst_Mem/inst_mem_reg[18][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][19]  ( .D(\Inst_Mem/inst_mem_reg[18][19] ), .CLK(clk), .RST(rst), .I(g_init[595]), .Q(\Inst_Mem/inst_mem_reg[18][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][20]  ( .D(\Inst_Mem/inst_mem_reg[18][20] ), .CLK(clk), .RST(rst), .I(g_init[596]), .Q(\Inst_Mem/inst_mem_reg[18][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][21]  ( .D(\Inst_Mem/inst_mem_reg[18][21] ), .CLK(clk), .RST(rst), .I(g_init[597]), .Q(\Inst_Mem/inst_mem_reg[18][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][22]  ( .D(\Inst_Mem/inst_mem_reg[18][22] ), .CLK(clk), .RST(rst), .I(g_init[598]), .Q(\Inst_Mem/inst_mem_reg[18][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][23]  ( .D(\Inst_Mem/inst_mem_reg[18][23] ), .CLK(clk), .RST(rst), .I(g_init[599]), .Q(\Inst_Mem/inst_mem_reg[18][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][24]  ( .D(\Inst_Mem/inst_mem_reg[18][24] ), .CLK(clk), .RST(rst), .I(g_init[600]), .Q(\Inst_Mem/inst_mem_reg[18][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][25]  ( .D(\Inst_Mem/inst_mem_reg[18][25] ), .CLK(clk), .RST(rst), .I(g_init[601]), .Q(\Inst_Mem/inst_mem_reg[18][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][26]  ( .D(\Inst_Mem/inst_mem_reg[18][26] ), .CLK(clk), .RST(rst), .I(g_init[602]), .Q(\Inst_Mem/inst_mem_reg[18][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][27]  ( .D(\Inst_Mem/inst_mem_reg[18][27] ), .CLK(clk), .RST(rst), .I(g_init[603]), .Q(\Inst_Mem/inst_mem_reg[18][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][28]  ( .D(\Inst_Mem/inst_mem_reg[18][28] ), .CLK(clk), .RST(rst), .I(g_init[604]), .Q(\Inst_Mem/inst_mem_reg[18][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][29]  ( .D(\Inst_Mem/inst_mem_reg[18][29] ), .CLK(clk), .RST(rst), .I(g_init[605]), .Q(\Inst_Mem/inst_mem_reg[18][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][30]  ( .D(\Inst_Mem/inst_mem_reg[18][30] ), .CLK(clk), .RST(rst), .I(g_init[606]), .Q(\Inst_Mem/inst_mem_reg[18][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[18][31]  ( .D(\Inst_Mem/inst_mem_reg[18][31] ), .CLK(clk), .RST(rst), .I(g_init[607]), .Q(\Inst_Mem/inst_mem_reg[18][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][0]  ( .D(\Inst_Mem/inst_mem_reg[17][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[544]), .Q(
        \Inst_Mem/inst_mem_reg[17][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][1]  ( .D(\Inst_Mem/inst_mem_reg[17][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[545]), .Q(
        \Inst_Mem/inst_mem_reg[17][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][2]  ( .D(\Inst_Mem/inst_mem_reg[17][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[546]), .Q(
        \Inst_Mem/inst_mem_reg[17][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][3]  ( .D(\Inst_Mem/inst_mem_reg[17][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[547]), .Q(
        \Inst_Mem/inst_mem_reg[17][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][4]  ( .D(\Inst_Mem/inst_mem_reg[17][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[548]), .Q(
        \Inst_Mem/inst_mem_reg[17][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][5]  ( .D(\Inst_Mem/inst_mem_reg[17][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[549]), .Q(
        \Inst_Mem/inst_mem_reg[17][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][6]  ( .D(\Inst_Mem/inst_mem_reg[17][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[550]), .Q(
        \Inst_Mem/inst_mem_reg[17][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][7]  ( .D(\Inst_Mem/inst_mem_reg[17][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[551]), .Q(
        \Inst_Mem/inst_mem_reg[17][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][8]  ( .D(\Inst_Mem/inst_mem_reg[17][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[552]), .Q(
        \Inst_Mem/inst_mem_reg[17][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][9]  ( .D(\Inst_Mem/inst_mem_reg[17][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[553]), .Q(
        \Inst_Mem/inst_mem_reg[17][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[17][10]  ( .D(\Inst_Mem/inst_mem_reg[17][10] ), .CLK(clk), .RST(rst), .I(g_init[554]), .Q(\Inst_Mem/inst_mem_reg[17][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][11]  ( .D(\Inst_Mem/inst_mem_reg[17][11] ), .CLK(clk), .RST(rst), .I(g_init[555]), .Q(\Inst_Mem/inst_mem_reg[17][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][12]  ( .D(\Inst_Mem/inst_mem_reg[17][12] ), .CLK(clk), .RST(rst), .I(g_init[556]), .Q(\Inst_Mem/inst_mem_reg[17][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][13]  ( .D(\Inst_Mem/inst_mem_reg[17][13] ), .CLK(clk), .RST(rst), .I(g_init[557]), .Q(\Inst_Mem/inst_mem_reg[17][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][14]  ( .D(\Inst_Mem/inst_mem_reg[17][14] ), .CLK(clk), .RST(rst), .I(g_init[558]), .Q(\Inst_Mem/inst_mem_reg[17][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][15]  ( .D(\Inst_Mem/inst_mem_reg[17][15] ), .CLK(clk), .RST(rst), .I(g_init[559]), .Q(\Inst_Mem/inst_mem_reg[17][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][16]  ( .D(\Inst_Mem/inst_mem_reg[17][16] ), .CLK(clk), .RST(rst), .I(g_init[560]), .Q(\Inst_Mem/inst_mem_reg[17][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][17]  ( .D(\Inst_Mem/inst_mem_reg[17][17] ), .CLK(clk), .RST(rst), .I(g_init[561]), .Q(\Inst_Mem/inst_mem_reg[17][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][18]  ( .D(\Inst_Mem/inst_mem_reg[17][18] ), .CLK(clk), .RST(rst), .I(g_init[562]), .Q(\Inst_Mem/inst_mem_reg[17][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][19]  ( .D(\Inst_Mem/inst_mem_reg[17][19] ), .CLK(clk), .RST(rst), .I(g_init[563]), .Q(\Inst_Mem/inst_mem_reg[17][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][20]  ( .D(\Inst_Mem/inst_mem_reg[17][20] ), .CLK(clk), .RST(rst), .I(g_init[564]), .Q(\Inst_Mem/inst_mem_reg[17][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][21]  ( .D(\Inst_Mem/inst_mem_reg[17][21] ), .CLK(clk), .RST(rst), .I(g_init[565]), .Q(\Inst_Mem/inst_mem_reg[17][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][22]  ( .D(\Inst_Mem/inst_mem_reg[17][22] ), .CLK(clk), .RST(rst), .I(g_init[566]), .Q(\Inst_Mem/inst_mem_reg[17][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][23]  ( .D(\Inst_Mem/inst_mem_reg[17][23] ), .CLK(clk), .RST(rst), .I(g_init[567]), .Q(\Inst_Mem/inst_mem_reg[17][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][24]  ( .D(\Inst_Mem/inst_mem_reg[17][24] ), .CLK(clk), .RST(rst), .I(g_init[568]), .Q(\Inst_Mem/inst_mem_reg[17][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][25]  ( .D(\Inst_Mem/inst_mem_reg[17][25] ), .CLK(clk), .RST(rst), .I(g_init[569]), .Q(\Inst_Mem/inst_mem_reg[17][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][26]  ( .D(\Inst_Mem/inst_mem_reg[17][26] ), .CLK(clk), .RST(rst), .I(g_init[570]), .Q(\Inst_Mem/inst_mem_reg[17][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][27]  ( .D(\Inst_Mem/inst_mem_reg[17][27] ), .CLK(clk), .RST(rst), .I(g_init[571]), .Q(\Inst_Mem/inst_mem_reg[17][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][28]  ( .D(\Inst_Mem/inst_mem_reg[17][28] ), .CLK(clk), .RST(rst), .I(g_init[572]), .Q(\Inst_Mem/inst_mem_reg[17][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][29]  ( .D(\Inst_Mem/inst_mem_reg[17][29] ), .CLK(clk), .RST(rst), .I(g_init[573]), .Q(\Inst_Mem/inst_mem_reg[17][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][30]  ( .D(\Inst_Mem/inst_mem_reg[17][30] ), .CLK(clk), .RST(rst), .I(g_init[574]), .Q(\Inst_Mem/inst_mem_reg[17][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[17][31]  ( .D(\Inst_Mem/inst_mem_reg[17][31] ), .CLK(clk), .RST(rst), .I(g_init[575]), .Q(\Inst_Mem/inst_mem_reg[17][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][0]  ( .D(\Inst_Mem/inst_mem_reg[16][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[512]), .Q(
        \Inst_Mem/inst_mem_reg[16][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][1]  ( .D(\Inst_Mem/inst_mem_reg[16][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[513]), .Q(
        \Inst_Mem/inst_mem_reg[16][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][2]  ( .D(\Inst_Mem/inst_mem_reg[16][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[514]), .Q(
        \Inst_Mem/inst_mem_reg[16][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][3]  ( .D(\Inst_Mem/inst_mem_reg[16][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[515]), .Q(
        \Inst_Mem/inst_mem_reg[16][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][4]  ( .D(\Inst_Mem/inst_mem_reg[16][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[516]), .Q(
        \Inst_Mem/inst_mem_reg[16][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][5]  ( .D(\Inst_Mem/inst_mem_reg[16][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[517]), .Q(
        \Inst_Mem/inst_mem_reg[16][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][6]  ( .D(\Inst_Mem/inst_mem_reg[16][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[518]), .Q(
        \Inst_Mem/inst_mem_reg[16][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][7]  ( .D(\Inst_Mem/inst_mem_reg[16][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[519]), .Q(
        \Inst_Mem/inst_mem_reg[16][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][8]  ( .D(\Inst_Mem/inst_mem_reg[16][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[520]), .Q(
        \Inst_Mem/inst_mem_reg[16][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][9]  ( .D(\Inst_Mem/inst_mem_reg[16][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[521]), .Q(
        \Inst_Mem/inst_mem_reg[16][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[16][10]  ( .D(\Inst_Mem/inst_mem_reg[16][10] ), .CLK(clk), .RST(rst), .I(g_init[522]), .Q(\Inst_Mem/inst_mem_reg[16][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][11]  ( .D(\Inst_Mem/inst_mem_reg[16][11] ), .CLK(clk), .RST(rst), .I(g_init[523]), .Q(\Inst_Mem/inst_mem_reg[16][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][12]  ( .D(\Inst_Mem/inst_mem_reg[16][12] ), .CLK(clk), .RST(rst), .I(g_init[524]), .Q(\Inst_Mem/inst_mem_reg[16][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][13]  ( .D(\Inst_Mem/inst_mem_reg[16][13] ), .CLK(clk), .RST(rst), .I(g_init[525]), .Q(\Inst_Mem/inst_mem_reg[16][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][14]  ( .D(\Inst_Mem/inst_mem_reg[16][14] ), .CLK(clk), .RST(rst), .I(g_init[526]), .Q(\Inst_Mem/inst_mem_reg[16][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][15]  ( .D(\Inst_Mem/inst_mem_reg[16][15] ), .CLK(clk), .RST(rst), .I(g_init[527]), .Q(\Inst_Mem/inst_mem_reg[16][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][16]  ( .D(\Inst_Mem/inst_mem_reg[16][16] ), .CLK(clk), .RST(rst), .I(g_init[528]), .Q(\Inst_Mem/inst_mem_reg[16][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][17]  ( .D(\Inst_Mem/inst_mem_reg[16][17] ), .CLK(clk), .RST(rst), .I(g_init[529]), .Q(\Inst_Mem/inst_mem_reg[16][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][18]  ( .D(\Inst_Mem/inst_mem_reg[16][18] ), .CLK(clk), .RST(rst), .I(g_init[530]), .Q(\Inst_Mem/inst_mem_reg[16][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][19]  ( .D(\Inst_Mem/inst_mem_reg[16][19] ), .CLK(clk), .RST(rst), .I(g_init[531]), .Q(\Inst_Mem/inst_mem_reg[16][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][20]  ( .D(\Inst_Mem/inst_mem_reg[16][20] ), .CLK(clk), .RST(rst), .I(g_init[532]), .Q(\Inst_Mem/inst_mem_reg[16][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][21]  ( .D(\Inst_Mem/inst_mem_reg[16][21] ), .CLK(clk), .RST(rst), .I(g_init[533]), .Q(\Inst_Mem/inst_mem_reg[16][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][22]  ( .D(\Inst_Mem/inst_mem_reg[16][22] ), .CLK(clk), .RST(rst), .I(g_init[534]), .Q(\Inst_Mem/inst_mem_reg[16][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][23]  ( .D(\Inst_Mem/inst_mem_reg[16][23] ), .CLK(clk), .RST(rst), .I(g_init[535]), .Q(\Inst_Mem/inst_mem_reg[16][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][24]  ( .D(\Inst_Mem/inst_mem_reg[16][24] ), .CLK(clk), .RST(rst), .I(g_init[536]), .Q(\Inst_Mem/inst_mem_reg[16][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][25]  ( .D(\Inst_Mem/inst_mem_reg[16][25] ), .CLK(clk), .RST(rst), .I(g_init[537]), .Q(\Inst_Mem/inst_mem_reg[16][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][26]  ( .D(\Inst_Mem/inst_mem_reg[16][26] ), .CLK(clk), .RST(rst), .I(g_init[538]), .Q(\Inst_Mem/inst_mem_reg[16][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][27]  ( .D(\Inst_Mem/inst_mem_reg[16][27] ), .CLK(clk), .RST(rst), .I(g_init[539]), .Q(\Inst_Mem/inst_mem_reg[16][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][28]  ( .D(\Inst_Mem/inst_mem_reg[16][28] ), .CLK(clk), .RST(rst), .I(g_init[540]), .Q(\Inst_Mem/inst_mem_reg[16][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][29]  ( .D(\Inst_Mem/inst_mem_reg[16][29] ), .CLK(clk), .RST(rst), .I(g_init[541]), .Q(\Inst_Mem/inst_mem_reg[16][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][30]  ( .D(\Inst_Mem/inst_mem_reg[16][30] ), .CLK(clk), .RST(rst), .I(g_init[542]), .Q(\Inst_Mem/inst_mem_reg[16][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[16][31]  ( .D(\Inst_Mem/inst_mem_reg[16][31] ), .CLK(clk), .RST(rst), .I(g_init[543]), .Q(\Inst_Mem/inst_mem_reg[16][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][0]  ( .D(\Inst_Mem/inst_mem_reg[15][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[480]), .Q(
        \Inst_Mem/inst_mem_reg[15][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][1]  ( .D(\Inst_Mem/inst_mem_reg[15][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[481]), .Q(
        \Inst_Mem/inst_mem_reg[15][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][2]  ( .D(\Inst_Mem/inst_mem_reg[15][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[482]), .Q(
        \Inst_Mem/inst_mem_reg[15][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][3]  ( .D(\Inst_Mem/inst_mem_reg[15][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[483]), .Q(
        \Inst_Mem/inst_mem_reg[15][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][4]  ( .D(\Inst_Mem/inst_mem_reg[15][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[484]), .Q(
        \Inst_Mem/inst_mem_reg[15][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][5]  ( .D(\Inst_Mem/inst_mem_reg[15][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[485]), .Q(
        \Inst_Mem/inst_mem_reg[15][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][6]  ( .D(\Inst_Mem/inst_mem_reg[15][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[486]), .Q(
        \Inst_Mem/inst_mem_reg[15][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][7]  ( .D(\Inst_Mem/inst_mem_reg[15][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[487]), .Q(
        \Inst_Mem/inst_mem_reg[15][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][8]  ( .D(\Inst_Mem/inst_mem_reg[15][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[488]), .Q(
        \Inst_Mem/inst_mem_reg[15][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][9]  ( .D(\Inst_Mem/inst_mem_reg[15][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[489]), .Q(
        \Inst_Mem/inst_mem_reg[15][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[15][10]  ( .D(\Inst_Mem/inst_mem_reg[15][10] ), .CLK(clk), .RST(rst), .I(g_init[490]), .Q(\Inst_Mem/inst_mem_reg[15][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][11]  ( .D(\Inst_Mem/inst_mem_reg[15][11] ), .CLK(clk), .RST(rst), .I(g_init[491]), .Q(\Inst_Mem/inst_mem_reg[15][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][12]  ( .D(\Inst_Mem/inst_mem_reg[15][12] ), .CLK(clk), .RST(rst), .I(g_init[492]), .Q(\Inst_Mem/inst_mem_reg[15][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][13]  ( .D(\Inst_Mem/inst_mem_reg[15][13] ), .CLK(clk), .RST(rst), .I(g_init[493]), .Q(\Inst_Mem/inst_mem_reg[15][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][14]  ( .D(\Inst_Mem/inst_mem_reg[15][14] ), .CLK(clk), .RST(rst), .I(g_init[494]), .Q(\Inst_Mem/inst_mem_reg[15][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][15]  ( .D(\Inst_Mem/inst_mem_reg[15][15] ), .CLK(clk), .RST(rst), .I(g_init[495]), .Q(\Inst_Mem/inst_mem_reg[15][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][16]  ( .D(\Inst_Mem/inst_mem_reg[15][16] ), .CLK(clk), .RST(rst), .I(g_init[496]), .Q(\Inst_Mem/inst_mem_reg[15][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][17]  ( .D(\Inst_Mem/inst_mem_reg[15][17] ), .CLK(clk), .RST(rst), .I(g_init[497]), .Q(\Inst_Mem/inst_mem_reg[15][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][18]  ( .D(\Inst_Mem/inst_mem_reg[15][18] ), .CLK(clk), .RST(rst), .I(g_init[498]), .Q(\Inst_Mem/inst_mem_reg[15][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][19]  ( .D(\Inst_Mem/inst_mem_reg[15][19] ), .CLK(clk), .RST(rst), .I(g_init[499]), .Q(\Inst_Mem/inst_mem_reg[15][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][20]  ( .D(\Inst_Mem/inst_mem_reg[15][20] ), .CLK(clk), .RST(rst), .I(g_init[500]), .Q(\Inst_Mem/inst_mem_reg[15][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][21]  ( .D(\Inst_Mem/inst_mem_reg[15][21] ), .CLK(clk), .RST(rst), .I(g_init[501]), .Q(\Inst_Mem/inst_mem_reg[15][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][22]  ( .D(\Inst_Mem/inst_mem_reg[15][22] ), .CLK(clk), .RST(rst), .I(g_init[502]), .Q(\Inst_Mem/inst_mem_reg[15][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][23]  ( .D(\Inst_Mem/inst_mem_reg[15][23] ), .CLK(clk), .RST(rst), .I(g_init[503]), .Q(\Inst_Mem/inst_mem_reg[15][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][24]  ( .D(\Inst_Mem/inst_mem_reg[15][24] ), .CLK(clk), .RST(rst), .I(g_init[504]), .Q(\Inst_Mem/inst_mem_reg[15][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][25]  ( .D(\Inst_Mem/inst_mem_reg[15][25] ), .CLK(clk), .RST(rst), .I(g_init[505]), .Q(\Inst_Mem/inst_mem_reg[15][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][26]  ( .D(\Inst_Mem/inst_mem_reg[15][26] ), .CLK(clk), .RST(rst), .I(g_init[506]), .Q(\Inst_Mem/inst_mem_reg[15][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][27]  ( .D(\Inst_Mem/inst_mem_reg[15][27] ), .CLK(clk), .RST(rst), .I(g_init[507]), .Q(\Inst_Mem/inst_mem_reg[15][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][28]  ( .D(\Inst_Mem/inst_mem_reg[15][28] ), .CLK(clk), .RST(rst), .I(g_init[508]), .Q(\Inst_Mem/inst_mem_reg[15][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][29]  ( .D(\Inst_Mem/inst_mem_reg[15][29] ), .CLK(clk), .RST(rst), .I(g_init[509]), .Q(\Inst_Mem/inst_mem_reg[15][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][30]  ( .D(\Inst_Mem/inst_mem_reg[15][30] ), .CLK(clk), .RST(rst), .I(g_init[510]), .Q(\Inst_Mem/inst_mem_reg[15][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[15][31]  ( .D(\Inst_Mem/inst_mem_reg[15][31] ), .CLK(clk), .RST(rst), .I(g_init[511]), .Q(\Inst_Mem/inst_mem_reg[15][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][0]  ( .D(\Inst_Mem/inst_mem_reg[14][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[448]), .Q(
        \Inst_Mem/inst_mem_reg[14][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][1]  ( .D(\Inst_Mem/inst_mem_reg[14][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[449]), .Q(
        \Inst_Mem/inst_mem_reg[14][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][2]  ( .D(\Inst_Mem/inst_mem_reg[14][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[450]), .Q(
        \Inst_Mem/inst_mem_reg[14][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][3]  ( .D(\Inst_Mem/inst_mem_reg[14][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[451]), .Q(
        \Inst_Mem/inst_mem_reg[14][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][4]  ( .D(\Inst_Mem/inst_mem_reg[14][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[452]), .Q(
        \Inst_Mem/inst_mem_reg[14][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][5]  ( .D(\Inst_Mem/inst_mem_reg[14][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[453]), .Q(
        \Inst_Mem/inst_mem_reg[14][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][6]  ( .D(\Inst_Mem/inst_mem_reg[14][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[454]), .Q(
        \Inst_Mem/inst_mem_reg[14][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][7]  ( .D(\Inst_Mem/inst_mem_reg[14][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[455]), .Q(
        \Inst_Mem/inst_mem_reg[14][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][8]  ( .D(\Inst_Mem/inst_mem_reg[14][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[456]), .Q(
        \Inst_Mem/inst_mem_reg[14][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][9]  ( .D(\Inst_Mem/inst_mem_reg[14][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[457]), .Q(
        \Inst_Mem/inst_mem_reg[14][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[14][10]  ( .D(\Inst_Mem/inst_mem_reg[14][10] ), .CLK(clk), .RST(rst), .I(g_init[458]), .Q(\Inst_Mem/inst_mem_reg[14][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][11]  ( .D(\Inst_Mem/inst_mem_reg[14][11] ), .CLK(clk), .RST(rst), .I(g_init[459]), .Q(\Inst_Mem/inst_mem_reg[14][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][12]  ( .D(\Inst_Mem/inst_mem_reg[14][12] ), .CLK(clk), .RST(rst), .I(g_init[460]), .Q(\Inst_Mem/inst_mem_reg[14][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][13]  ( .D(\Inst_Mem/inst_mem_reg[14][13] ), .CLK(clk), .RST(rst), .I(g_init[461]), .Q(\Inst_Mem/inst_mem_reg[14][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][14]  ( .D(\Inst_Mem/inst_mem_reg[14][14] ), .CLK(clk), .RST(rst), .I(g_init[462]), .Q(\Inst_Mem/inst_mem_reg[14][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][15]  ( .D(\Inst_Mem/inst_mem_reg[14][15] ), .CLK(clk), .RST(rst), .I(g_init[463]), .Q(\Inst_Mem/inst_mem_reg[14][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][16]  ( .D(\Inst_Mem/inst_mem_reg[14][16] ), .CLK(clk), .RST(rst), .I(g_init[464]), .Q(\Inst_Mem/inst_mem_reg[14][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][17]  ( .D(\Inst_Mem/inst_mem_reg[14][17] ), .CLK(clk), .RST(rst), .I(g_init[465]), .Q(\Inst_Mem/inst_mem_reg[14][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][18]  ( .D(\Inst_Mem/inst_mem_reg[14][18] ), .CLK(clk), .RST(rst), .I(g_init[466]), .Q(\Inst_Mem/inst_mem_reg[14][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][19]  ( .D(\Inst_Mem/inst_mem_reg[14][19] ), .CLK(clk), .RST(rst), .I(g_init[467]), .Q(\Inst_Mem/inst_mem_reg[14][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][20]  ( .D(\Inst_Mem/inst_mem_reg[14][20] ), .CLK(clk), .RST(rst), .I(g_init[468]), .Q(\Inst_Mem/inst_mem_reg[14][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][21]  ( .D(\Inst_Mem/inst_mem_reg[14][21] ), .CLK(clk), .RST(rst), .I(g_init[469]), .Q(\Inst_Mem/inst_mem_reg[14][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][22]  ( .D(\Inst_Mem/inst_mem_reg[14][22] ), .CLK(clk), .RST(rst), .I(g_init[470]), .Q(\Inst_Mem/inst_mem_reg[14][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][23]  ( .D(\Inst_Mem/inst_mem_reg[14][23] ), .CLK(clk), .RST(rst), .I(g_init[471]), .Q(\Inst_Mem/inst_mem_reg[14][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][24]  ( .D(\Inst_Mem/inst_mem_reg[14][24] ), .CLK(clk), .RST(rst), .I(g_init[472]), .Q(\Inst_Mem/inst_mem_reg[14][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][25]  ( .D(\Inst_Mem/inst_mem_reg[14][25] ), .CLK(clk), .RST(rst), .I(g_init[473]), .Q(\Inst_Mem/inst_mem_reg[14][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][26]  ( .D(\Inst_Mem/inst_mem_reg[14][26] ), .CLK(clk), .RST(rst), .I(g_init[474]), .Q(\Inst_Mem/inst_mem_reg[14][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][27]  ( .D(\Inst_Mem/inst_mem_reg[14][27] ), .CLK(clk), .RST(rst), .I(g_init[475]), .Q(\Inst_Mem/inst_mem_reg[14][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][28]  ( .D(\Inst_Mem/inst_mem_reg[14][28] ), .CLK(clk), .RST(rst), .I(g_init[476]), .Q(\Inst_Mem/inst_mem_reg[14][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][29]  ( .D(\Inst_Mem/inst_mem_reg[14][29] ), .CLK(clk), .RST(rst), .I(g_init[477]), .Q(\Inst_Mem/inst_mem_reg[14][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][30]  ( .D(\Inst_Mem/inst_mem_reg[14][30] ), .CLK(clk), .RST(rst), .I(g_init[478]), .Q(\Inst_Mem/inst_mem_reg[14][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[14][31]  ( .D(\Inst_Mem/inst_mem_reg[14][31] ), .CLK(clk), .RST(rst), .I(g_init[479]), .Q(\Inst_Mem/inst_mem_reg[14][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][0]  ( .D(\Inst_Mem/inst_mem_reg[13][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[416]), .Q(
        \Inst_Mem/inst_mem_reg[13][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][1]  ( .D(\Inst_Mem/inst_mem_reg[13][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[417]), .Q(
        \Inst_Mem/inst_mem_reg[13][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][2]  ( .D(\Inst_Mem/inst_mem_reg[13][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[418]), .Q(
        \Inst_Mem/inst_mem_reg[13][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][3]  ( .D(\Inst_Mem/inst_mem_reg[13][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[419]), .Q(
        \Inst_Mem/inst_mem_reg[13][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][4]  ( .D(\Inst_Mem/inst_mem_reg[13][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[420]), .Q(
        \Inst_Mem/inst_mem_reg[13][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][5]  ( .D(\Inst_Mem/inst_mem_reg[13][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[421]), .Q(
        \Inst_Mem/inst_mem_reg[13][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][6]  ( .D(\Inst_Mem/inst_mem_reg[13][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[422]), .Q(
        \Inst_Mem/inst_mem_reg[13][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][7]  ( .D(\Inst_Mem/inst_mem_reg[13][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[423]), .Q(
        \Inst_Mem/inst_mem_reg[13][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][8]  ( .D(\Inst_Mem/inst_mem_reg[13][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[424]), .Q(
        \Inst_Mem/inst_mem_reg[13][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][9]  ( .D(\Inst_Mem/inst_mem_reg[13][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[425]), .Q(
        \Inst_Mem/inst_mem_reg[13][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[13][10]  ( .D(\Inst_Mem/inst_mem_reg[13][10] ), .CLK(clk), .RST(rst), .I(g_init[426]), .Q(\Inst_Mem/inst_mem_reg[13][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][11]  ( .D(\Inst_Mem/inst_mem_reg[13][11] ), .CLK(clk), .RST(rst), .I(g_init[427]), .Q(\Inst_Mem/inst_mem_reg[13][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][12]  ( .D(\Inst_Mem/inst_mem_reg[13][12] ), .CLK(clk), .RST(rst), .I(g_init[428]), .Q(\Inst_Mem/inst_mem_reg[13][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][13]  ( .D(\Inst_Mem/inst_mem_reg[13][13] ), .CLK(clk), .RST(rst), .I(g_init[429]), .Q(\Inst_Mem/inst_mem_reg[13][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][14]  ( .D(\Inst_Mem/inst_mem_reg[13][14] ), .CLK(clk), .RST(rst), .I(g_init[430]), .Q(\Inst_Mem/inst_mem_reg[13][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][15]  ( .D(\Inst_Mem/inst_mem_reg[13][15] ), .CLK(clk), .RST(rst), .I(g_init[431]), .Q(\Inst_Mem/inst_mem_reg[13][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][16]  ( .D(\Inst_Mem/inst_mem_reg[13][16] ), .CLK(clk), .RST(rst), .I(g_init[432]), .Q(\Inst_Mem/inst_mem_reg[13][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][17]  ( .D(\Inst_Mem/inst_mem_reg[13][17] ), .CLK(clk), .RST(rst), .I(g_init[433]), .Q(\Inst_Mem/inst_mem_reg[13][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][18]  ( .D(\Inst_Mem/inst_mem_reg[13][18] ), .CLK(clk), .RST(rst), .I(g_init[434]), .Q(\Inst_Mem/inst_mem_reg[13][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][19]  ( .D(\Inst_Mem/inst_mem_reg[13][19] ), .CLK(clk), .RST(rst), .I(g_init[435]), .Q(\Inst_Mem/inst_mem_reg[13][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][20]  ( .D(\Inst_Mem/inst_mem_reg[13][20] ), .CLK(clk), .RST(rst), .I(g_init[436]), .Q(\Inst_Mem/inst_mem_reg[13][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][21]  ( .D(\Inst_Mem/inst_mem_reg[13][21] ), .CLK(clk), .RST(rst), .I(g_init[437]), .Q(\Inst_Mem/inst_mem_reg[13][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][22]  ( .D(\Inst_Mem/inst_mem_reg[13][22] ), .CLK(clk), .RST(rst), .I(g_init[438]), .Q(\Inst_Mem/inst_mem_reg[13][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][23]  ( .D(\Inst_Mem/inst_mem_reg[13][23] ), .CLK(clk), .RST(rst), .I(g_init[439]), .Q(\Inst_Mem/inst_mem_reg[13][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][24]  ( .D(\Inst_Mem/inst_mem_reg[13][24] ), .CLK(clk), .RST(rst), .I(g_init[440]), .Q(\Inst_Mem/inst_mem_reg[13][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][25]  ( .D(\Inst_Mem/inst_mem_reg[13][25] ), .CLK(clk), .RST(rst), .I(g_init[441]), .Q(\Inst_Mem/inst_mem_reg[13][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][26]  ( .D(\Inst_Mem/inst_mem_reg[13][26] ), .CLK(clk), .RST(rst), .I(g_init[442]), .Q(\Inst_Mem/inst_mem_reg[13][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][27]  ( .D(\Inst_Mem/inst_mem_reg[13][27] ), .CLK(clk), .RST(rst), .I(g_init[443]), .Q(\Inst_Mem/inst_mem_reg[13][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][28]  ( .D(\Inst_Mem/inst_mem_reg[13][28] ), .CLK(clk), .RST(rst), .I(g_init[444]), .Q(\Inst_Mem/inst_mem_reg[13][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][29]  ( .D(\Inst_Mem/inst_mem_reg[13][29] ), .CLK(clk), .RST(rst), .I(g_init[445]), .Q(\Inst_Mem/inst_mem_reg[13][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][30]  ( .D(\Inst_Mem/inst_mem_reg[13][30] ), .CLK(clk), .RST(rst), .I(g_init[446]), .Q(\Inst_Mem/inst_mem_reg[13][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[13][31]  ( .D(\Inst_Mem/inst_mem_reg[13][31] ), .CLK(clk), .RST(rst), .I(g_init[447]), .Q(\Inst_Mem/inst_mem_reg[13][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][0]  ( .D(\Inst_Mem/inst_mem_reg[12][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[384]), .Q(
        \Inst_Mem/inst_mem_reg[12][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][1]  ( .D(\Inst_Mem/inst_mem_reg[12][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[385]), .Q(
        \Inst_Mem/inst_mem_reg[12][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][2]  ( .D(\Inst_Mem/inst_mem_reg[12][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[386]), .Q(
        \Inst_Mem/inst_mem_reg[12][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][3]  ( .D(\Inst_Mem/inst_mem_reg[12][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[387]), .Q(
        \Inst_Mem/inst_mem_reg[12][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][4]  ( .D(\Inst_Mem/inst_mem_reg[12][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[388]), .Q(
        \Inst_Mem/inst_mem_reg[12][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][5]  ( .D(\Inst_Mem/inst_mem_reg[12][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[389]), .Q(
        \Inst_Mem/inst_mem_reg[12][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][6]  ( .D(\Inst_Mem/inst_mem_reg[12][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[390]), .Q(
        \Inst_Mem/inst_mem_reg[12][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][7]  ( .D(\Inst_Mem/inst_mem_reg[12][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[391]), .Q(
        \Inst_Mem/inst_mem_reg[12][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][8]  ( .D(\Inst_Mem/inst_mem_reg[12][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[392]), .Q(
        \Inst_Mem/inst_mem_reg[12][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][9]  ( .D(\Inst_Mem/inst_mem_reg[12][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[393]), .Q(
        \Inst_Mem/inst_mem_reg[12][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[12][10]  ( .D(\Inst_Mem/inst_mem_reg[12][10] ), .CLK(clk), .RST(rst), .I(g_init[394]), .Q(\Inst_Mem/inst_mem_reg[12][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][11]  ( .D(\Inst_Mem/inst_mem_reg[12][11] ), .CLK(clk), .RST(rst), .I(g_init[395]), .Q(\Inst_Mem/inst_mem_reg[12][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][12]  ( .D(\Inst_Mem/inst_mem_reg[12][12] ), .CLK(clk), .RST(rst), .I(g_init[396]), .Q(\Inst_Mem/inst_mem_reg[12][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][13]  ( .D(\Inst_Mem/inst_mem_reg[12][13] ), .CLK(clk), .RST(rst), .I(g_init[397]), .Q(\Inst_Mem/inst_mem_reg[12][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][14]  ( .D(\Inst_Mem/inst_mem_reg[12][14] ), .CLK(clk), .RST(rst), .I(g_init[398]), .Q(\Inst_Mem/inst_mem_reg[12][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][15]  ( .D(\Inst_Mem/inst_mem_reg[12][15] ), .CLK(clk), .RST(rst), .I(g_init[399]), .Q(\Inst_Mem/inst_mem_reg[12][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][16]  ( .D(\Inst_Mem/inst_mem_reg[12][16] ), .CLK(clk), .RST(rst), .I(g_init[400]), .Q(\Inst_Mem/inst_mem_reg[12][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][17]  ( .D(\Inst_Mem/inst_mem_reg[12][17] ), .CLK(clk), .RST(rst), .I(g_init[401]), .Q(\Inst_Mem/inst_mem_reg[12][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][18]  ( .D(\Inst_Mem/inst_mem_reg[12][18] ), .CLK(clk), .RST(rst), .I(g_init[402]), .Q(\Inst_Mem/inst_mem_reg[12][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][19]  ( .D(\Inst_Mem/inst_mem_reg[12][19] ), .CLK(clk), .RST(rst), .I(g_init[403]), .Q(\Inst_Mem/inst_mem_reg[12][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][20]  ( .D(\Inst_Mem/inst_mem_reg[12][20] ), .CLK(clk), .RST(rst), .I(g_init[404]), .Q(\Inst_Mem/inst_mem_reg[12][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][21]  ( .D(\Inst_Mem/inst_mem_reg[12][21] ), .CLK(clk), .RST(rst), .I(g_init[405]), .Q(\Inst_Mem/inst_mem_reg[12][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][22]  ( .D(\Inst_Mem/inst_mem_reg[12][22] ), .CLK(clk), .RST(rst), .I(g_init[406]), .Q(\Inst_Mem/inst_mem_reg[12][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][23]  ( .D(\Inst_Mem/inst_mem_reg[12][23] ), .CLK(clk), .RST(rst), .I(g_init[407]), .Q(\Inst_Mem/inst_mem_reg[12][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][24]  ( .D(\Inst_Mem/inst_mem_reg[12][24] ), .CLK(clk), .RST(rst), .I(g_init[408]), .Q(\Inst_Mem/inst_mem_reg[12][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][25]  ( .D(\Inst_Mem/inst_mem_reg[12][25] ), .CLK(clk), .RST(rst), .I(g_init[409]), .Q(\Inst_Mem/inst_mem_reg[12][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][26]  ( .D(\Inst_Mem/inst_mem_reg[12][26] ), .CLK(clk), .RST(rst), .I(g_init[410]), .Q(\Inst_Mem/inst_mem_reg[12][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][27]  ( .D(\Inst_Mem/inst_mem_reg[12][27] ), .CLK(clk), .RST(rst), .I(g_init[411]), .Q(\Inst_Mem/inst_mem_reg[12][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][28]  ( .D(\Inst_Mem/inst_mem_reg[12][28] ), .CLK(clk), .RST(rst), .I(g_init[412]), .Q(\Inst_Mem/inst_mem_reg[12][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][29]  ( .D(\Inst_Mem/inst_mem_reg[12][29] ), .CLK(clk), .RST(rst), .I(g_init[413]), .Q(\Inst_Mem/inst_mem_reg[12][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][30]  ( .D(\Inst_Mem/inst_mem_reg[12][30] ), .CLK(clk), .RST(rst), .I(g_init[414]), .Q(\Inst_Mem/inst_mem_reg[12][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[12][31]  ( .D(\Inst_Mem/inst_mem_reg[12][31] ), .CLK(clk), .RST(rst), .I(g_init[415]), .Q(\Inst_Mem/inst_mem_reg[12][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][0]  ( .D(\Inst_Mem/inst_mem_reg[11][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[352]), .Q(
        \Inst_Mem/inst_mem_reg[11][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][1]  ( .D(\Inst_Mem/inst_mem_reg[11][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[353]), .Q(
        \Inst_Mem/inst_mem_reg[11][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][2]  ( .D(\Inst_Mem/inst_mem_reg[11][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[354]), .Q(
        \Inst_Mem/inst_mem_reg[11][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][3]  ( .D(\Inst_Mem/inst_mem_reg[11][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[355]), .Q(
        \Inst_Mem/inst_mem_reg[11][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][4]  ( .D(\Inst_Mem/inst_mem_reg[11][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[356]), .Q(
        \Inst_Mem/inst_mem_reg[11][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][5]  ( .D(\Inst_Mem/inst_mem_reg[11][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[357]), .Q(
        \Inst_Mem/inst_mem_reg[11][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][6]  ( .D(\Inst_Mem/inst_mem_reg[11][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[358]), .Q(
        \Inst_Mem/inst_mem_reg[11][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][7]  ( .D(\Inst_Mem/inst_mem_reg[11][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[359]), .Q(
        \Inst_Mem/inst_mem_reg[11][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][8]  ( .D(\Inst_Mem/inst_mem_reg[11][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[360]), .Q(
        \Inst_Mem/inst_mem_reg[11][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][9]  ( .D(\Inst_Mem/inst_mem_reg[11][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[361]), .Q(
        \Inst_Mem/inst_mem_reg[11][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[11][10]  ( .D(\Inst_Mem/inst_mem_reg[11][10] ), .CLK(clk), .RST(rst), .I(g_init[362]), .Q(\Inst_Mem/inst_mem_reg[11][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][11]  ( .D(\Inst_Mem/inst_mem_reg[11][11] ), .CLK(clk), .RST(rst), .I(g_init[363]), .Q(\Inst_Mem/inst_mem_reg[11][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][12]  ( .D(\Inst_Mem/inst_mem_reg[11][12] ), .CLK(clk), .RST(rst), .I(g_init[364]), .Q(\Inst_Mem/inst_mem_reg[11][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][13]  ( .D(\Inst_Mem/inst_mem_reg[11][13] ), .CLK(clk), .RST(rst), .I(g_init[365]), .Q(\Inst_Mem/inst_mem_reg[11][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][14]  ( .D(\Inst_Mem/inst_mem_reg[11][14] ), .CLK(clk), .RST(rst), .I(g_init[366]), .Q(\Inst_Mem/inst_mem_reg[11][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][15]  ( .D(\Inst_Mem/inst_mem_reg[11][15] ), .CLK(clk), .RST(rst), .I(g_init[367]), .Q(\Inst_Mem/inst_mem_reg[11][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][16]  ( .D(\Inst_Mem/inst_mem_reg[11][16] ), .CLK(clk), .RST(rst), .I(g_init[368]), .Q(\Inst_Mem/inst_mem_reg[11][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][17]  ( .D(\Inst_Mem/inst_mem_reg[11][17] ), .CLK(clk), .RST(rst), .I(g_init[369]), .Q(\Inst_Mem/inst_mem_reg[11][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][18]  ( .D(\Inst_Mem/inst_mem_reg[11][18] ), .CLK(clk), .RST(rst), .I(g_init[370]), .Q(\Inst_Mem/inst_mem_reg[11][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][19]  ( .D(\Inst_Mem/inst_mem_reg[11][19] ), .CLK(clk), .RST(rst), .I(g_init[371]), .Q(\Inst_Mem/inst_mem_reg[11][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][20]  ( .D(\Inst_Mem/inst_mem_reg[11][20] ), .CLK(clk), .RST(rst), .I(g_init[372]), .Q(\Inst_Mem/inst_mem_reg[11][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][21]  ( .D(\Inst_Mem/inst_mem_reg[11][21] ), .CLK(clk), .RST(rst), .I(g_init[373]), .Q(\Inst_Mem/inst_mem_reg[11][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][22]  ( .D(\Inst_Mem/inst_mem_reg[11][22] ), .CLK(clk), .RST(rst), .I(g_init[374]), .Q(\Inst_Mem/inst_mem_reg[11][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][23]  ( .D(\Inst_Mem/inst_mem_reg[11][23] ), .CLK(clk), .RST(rst), .I(g_init[375]), .Q(\Inst_Mem/inst_mem_reg[11][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][24]  ( .D(\Inst_Mem/inst_mem_reg[11][24] ), .CLK(clk), .RST(rst), .I(g_init[376]), .Q(\Inst_Mem/inst_mem_reg[11][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][25]  ( .D(\Inst_Mem/inst_mem_reg[11][25] ), .CLK(clk), .RST(rst), .I(g_init[377]), .Q(\Inst_Mem/inst_mem_reg[11][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][26]  ( .D(\Inst_Mem/inst_mem_reg[11][26] ), .CLK(clk), .RST(rst), .I(g_init[378]), .Q(\Inst_Mem/inst_mem_reg[11][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][27]  ( .D(\Inst_Mem/inst_mem_reg[11][27] ), .CLK(clk), .RST(rst), .I(g_init[379]), .Q(\Inst_Mem/inst_mem_reg[11][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][28]  ( .D(\Inst_Mem/inst_mem_reg[11][28] ), .CLK(clk), .RST(rst), .I(g_init[380]), .Q(\Inst_Mem/inst_mem_reg[11][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][29]  ( .D(\Inst_Mem/inst_mem_reg[11][29] ), .CLK(clk), .RST(rst), .I(g_init[381]), .Q(\Inst_Mem/inst_mem_reg[11][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][30]  ( .D(\Inst_Mem/inst_mem_reg[11][30] ), .CLK(clk), .RST(rst), .I(g_init[382]), .Q(\Inst_Mem/inst_mem_reg[11][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[11][31]  ( .D(\Inst_Mem/inst_mem_reg[11][31] ), .CLK(clk), .RST(rst), .I(g_init[383]), .Q(\Inst_Mem/inst_mem_reg[11][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][0]  ( .D(\Inst_Mem/inst_mem_reg[10][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[320]), .Q(
        \Inst_Mem/inst_mem_reg[10][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][1]  ( .D(\Inst_Mem/inst_mem_reg[10][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[321]), .Q(
        \Inst_Mem/inst_mem_reg[10][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][2]  ( .D(\Inst_Mem/inst_mem_reg[10][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[322]), .Q(
        \Inst_Mem/inst_mem_reg[10][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][3]  ( .D(\Inst_Mem/inst_mem_reg[10][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[323]), .Q(
        \Inst_Mem/inst_mem_reg[10][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][4]  ( .D(\Inst_Mem/inst_mem_reg[10][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[324]), .Q(
        \Inst_Mem/inst_mem_reg[10][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][5]  ( .D(\Inst_Mem/inst_mem_reg[10][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[325]), .Q(
        \Inst_Mem/inst_mem_reg[10][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][6]  ( .D(\Inst_Mem/inst_mem_reg[10][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[326]), .Q(
        \Inst_Mem/inst_mem_reg[10][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][7]  ( .D(\Inst_Mem/inst_mem_reg[10][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[327]), .Q(
        \Inst_Mem/inst_mem_reg[10][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][8]  ( .D(\Inst_Mem/inst_mem_reg[10][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[328]), .Q(
        \Inst_Mem/inst_mem_reg[10][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][9]  ( .D(\Inst_Mem/inst_mem_reg[10][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[329]), .Q(
        \Inst_Mem/inst_mem_reg[10][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[10][10]  ( .D(\Inst_Mem/inst_mem_reg[10][10] ), .CLK(clk), .RST(rst), .I(g_init[330]), .Q(\Inst_Mem/inst_mem_reg[10][10] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][11]  ( .D(\Inst_Mem/inst_mem_reg[10][11] ), .CLK(clk), .RST(rst), .I(g_init[331]), .Q(\Inst_Mem/inst_mem_reg[10][11] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][12]  ( .D(\Inst_Mem/inst_mem_reg[10][12] ), .CLK(clk), .RST(rst), .I(g_init[332]), .Q(\Inst_Mem/inst_mem_reg[10][12] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][13]  ( .D(\Inst_Mem/inst_mem_reg[10][13] ), .CLK(clk), .RST(rst), .I(g_init[333]), .Q(\Inst_Mem/inst_mem_reg[10][13] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][14]  ( .D(\Inst_Mem/inst_mem_reg[10][14] ), .CLK(clk), .RST(rst), .I(g_init[334]), .Q(\Inst_Mem/inst_mem_reg[10][14] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][15]  ( .D(\Inst_Mem/inst_mem_reg[10][15] ), .CLK(clk), .RST(rst), .I(g_init[335]), .Q(\Inst_Mem/inst_mem_reg[10][15] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][16]  ( .D(\Inst_Mem/inst_mem_reg[10][16] ), .CLK(clk), .RST(rst), .I(g_init[336]), .Q(\Inst_Mem/inst_mem_reg[10][16] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][17]  ( .D(\Inst_Mem/inst_mem_reg[10][17] ), .CLK(clk), .RST(rst), .I(g_init[337]), .Q(\Inst_Mem/inst_mem_reg[10][17] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][18]  ( .D(\Inst_Mem/inst_mem_reg[10][18] ), .CLK(clk), .RST(rst), .I(g_init[338]), .Q(\Inst_Mem/inst_mem_reg[10][18] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][19]  ( .D(\Inst_Mem/inst_mem_reg[10][19] ), .CLK(clk), .RST(rst), .I(g_init[339]), .Q(\Inst_Mem/inst_mem_reg[10][19] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][20]  ( .D(\Inst_Mem/inst_mem_reg[10][20] ), .CLK(clk), .RST(rst), .I(g_init[340]), .Q(\Inst_Mem/inst_mem_reg[10][20] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][21]  ( .D(\Inst_Mem/inst_mem_reg[10][21] ), .CLK(clk), .RST(rst), .I(g_init[341]), .Q(\Inst_Mem/inst_mem_reg[10][21] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][22]  ( .D(\Inst_Mem/inst_mem_reg[10][22] ), .CLK(clk), .RST(rst), .I(g_init[342]), .Q(\Inst_Mem/inst_mem_reg[10][22] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][23]  ( .D(\Inst_Mem/inst_mem_reg[10][23] ), .CLK(clk), .RST(rst), .I(g_init[343]), .Q(\Inst_Mem/inst_mem_reg[10][23] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][24]  ( .D(\Inst_Mem/inst_mem_reg[10][24] ), .CLK(clk), .RST(rst), .I(g_init[344]), .Q(\Inst_Mem/inst_mem_reg[10][24] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][25]  ( .D(\Inst_Mem/inst_mem_reg[10][25] ), .CLK(clk), .RST(rst), .I(g_init[345]), .Q(\Inst_Mem/inst_mem_reg[10][25] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][26]  ( .D(\Inst_Mem/inst_mem_reg[10][26] ), .CLK(clk), .RST(rst), .I(g_init[346]), .Q(\Inst_Mem/inst_mem_reg[10][26] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][27]  ( .D(\Inst_Mem/inst_mem_reg[10][27] ), .CLK(clk), .RST(rst), .I(g_init[347]), .Q(\Inst_Mem/inst_mem_reg[10][27] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][28]  ( .D(\Inst_Mem/inst_mem_reg[10][28] ), .CLK(clk), .RST(rst), .I(g_init[348]), .Q(\Inst_Mem/inst_mem_reg[10][28] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][29]  ( .D(\Inst_Mem/inst_mem_reg[10][29] ), .CLK(clk), .RST(rst), .I(g_init[349]), .Q(\Inst_Mem/inst_mem_reg[10][29] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][30]  ( .D(\Inst_Mem/inst_mem_reg[10][30] ), .CLK(clk), .RST(rst), .I(g_init[350]), .Q(\Inst_Mem/inst_mem_reg[10][30] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[10][31]  ( .D(\Inst_Mem/inst_mem_reg[10][31] ), .CLK(clk), .RST(rst), .I(g_init[351]), .Q(\Inst_Mem/inst_mem_reg[10][31] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[9][0]  ( .D(\Inst_Mem/inst_mem_reg[9][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[288]), .Q(
        \Inst_Mem/inst_mem_reg[9][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][1]  ( .D(\Inst_Mem/inst_mem_reg[9][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[289]), .Q(
        \Inst_Mem/inst_mem_reg[9][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][2]  ( .D(\Inst_Mem/inst_mem_reg[9][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[290]), .Q(
        \Inst_Mem/inst_mem_reg[9][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][3]  ( .D(\Inst_Mem/inst_mem_reg[9][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[291]), .Q(
        \Inst_Mem/inst_mem_reg[9][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][4]  ( .D(\Inst_Mem/inst_mem_reg[9][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[292]), .Q(
        \Inst_Mem/inst_mem_reg[9][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][5]  ( .D(\Inst_Mem/inst_mem_reg[9][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[293]), .Q(
        \Inst_Mem/inst_mem_reg[9][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][6]  ( .D(\Inst_Mem/inst_mem_reg[9][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[294]), .Q(
        \Inst_Mem/inst_mem_reg[9][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][7]  ( .D(\Inst_Mem/inst_mem_reg[9][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[295]), .Q(
        \Inst_Mem/inst_mem_reg[9][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][8]  ( .D(\Inst_Mem/inst_mem_reg[9][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[296]), .Q(
        \Inst_Mem/inst_mem_reg[9][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][9]  ( .D(\Inst_Mem/inst_mem_reg[9][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[297]), .Q(
        \Inst_Mem/inst_mem_reg[9][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][10]  ( .D(\Inst_Mem/inst_mem_reg[9][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[298]), .Q(
        \Inst_Mem/inst_mem_reg[9][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][11]  ( .D(\Inst_Mem/inst_mem_reg[9][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[299]), .Q(
        \Inst_Mem/inst_mem_reg[9][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][12]  ( .D(\Inst_Mem/inst_mem_reg[9][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[300]), .Q(
        \Inst_Mem/inst_mem_reg[9][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][13]  ( .D(\Inst_Mem/inst_mem_reg[9][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[301]), .Q(
        \Inst_Mem/inst_mem_reg[9][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][14]  ( .D(\Inst_Mem/inst_mem_reg[9][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[302]), .Q(
        \Inst_Mem/inst_mem_reg[9][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][15]  ( .D(\Inst_Mem/inst_mem_reg[9][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[303]), .Q(
        \Inst_Mem/inst_mem_reg[9][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][16]  ( .D(\Inst_Mem/inst_mem_reg[9][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[304]), .Q(
        \Inst_Mem/inst_mem_reg[9][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][17]  ( .D(\Inst_Mem/inst_mem_reg[9][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[305]), .Q(
        \Inst_Mem/inst_mem_reg[9][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][18]  ( .D(\Inst_Mem/inst_mem_reg[9][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[306]), .Q(
        \Inst_Mem/inst_mem_reg[9][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][19]  ( .D(\Inst_Mem/inst_mem_reg[9][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[307]), .Q(
        \Inst_Mem/inst_mem_reg[9][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][20]  ( .D(\Inst_Mem/inst_mem_reg[9][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[308]), .Q(
        \Inst_Mem/inst_mem_reg[9][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][21]  ( .D(\Inst_Mem/inst_mem_reg[9][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[309]), .Q(
        \Inst_Mem/inst_mem_reg[9][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][22]  ( .D(\Inst_Mem/inst_mem_reg[9][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[310]), .Q(
        \Inst_Mem/inst_mem_reg[9][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][23]  ( .D(\Inst_Mem/inst_mem_reg[9][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[311]), .Q(
        \Inst_Mem/inst_mem_reg[9][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][24]  ( .D(\Inst_Mem/inst_mem_reg[9][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[312]), .Q(
        \Inst_Mem/inst_mem_reg[9][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][25]  ( .D(\Inst_Mem/inst_mem_reg[9][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[313]), .Q(
        \Inst_Mem/inst_mem_reg[9][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][26]  ( .D(\Inst_Mem/inst_mem_reg[9][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[314]), .Q(
        \Inst_Mem/inst_mem_reg[9][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][27]  ( .D(\Inst_Mem/inst_mem_reg[9][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[315]), .Q(
        \Inst_Mem/inst_mem_reg[9][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][28]  ( .D(\Inst_Mem/inst_mem_reg[9][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[316]), .Q(
        \Inst_Mem/inst_mem_reg[9][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][29]  ( .D(\Inst_Mem/inst_mem_reg[9][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[317]), .Q(
        \Inst_Mem/inst_mem_reg[9][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][30]  ( .D(\Inst_Mem/inst_mem_reg[9][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[318]), .Q(
        \Inst_Mem/inst_mem_reg[9][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[9][31]  ( .D(\Inst_Mem/inst_mem_reg[9][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[319]), .Q(
        \Inst_Mem/inst_mem_reg[9][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][0]  ( .D(\Inst_Mem/inst_mem_reg[8][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[256]), .Q(
        \Inst_Mem/inst_mem_reg[8][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][1]  ( .D(\Inst_Mem/inst_mem_reg[8][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[257]), .Q(
        \Inst_Mem/inst_mem_reg[8][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][2]  ( .D(\Inst_Mem/inst_mem_reg[8][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[258]), .Q(
        \Inst_Mem/inst_mem_reg[8][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][3]  ( .D(\Inst_Mem/inst_mem_reg[8][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[259]), .Q(
        \Inst_Mem/inst_mem_reg[8][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][4]  ( .D(\Inst_Mem/inst_mem_reg[8][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[260]), .Q(
        \Inst_Mem/inst_mem_reg[8][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][5]  ( .D(\Inst_Mem/inst_mem_reg[8][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[261]), .Q(
        \Inst_Mem/inst_mem_reg[8][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][6]  ( .D(\Inst_Mem/inst_mem_reg[8][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[262]), .Q(
        \Inst_Mem/inst_mem_reg[8][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][7]  ( .D(\Inst_Mem/inst_mem_reg[8][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[263]), .Q(
        \Inst_Mem/inst_mem_reg[8][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][8]  ( .D(\Inst_Mem/inst_mem_reg[8][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[264]), .Q(
        \Inst_Mem/inst_mem_reg[8][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][9]  ( .D(\Inst_Mem/inst_mem_reg[8][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[265]), .Q(
        \Inst_Mem/inst_mem_reg[8][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][10]  ( .D(\Inst_Mem/inst_mem_reg[8][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[266]), .Q(
        \Inst_Mem/inst_mem_reg[8][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][11]  ( .D(\Inst_Mem/inst_mem_reg[8][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[267]), .Q(
        \Inst_Mem/inst_mem_reg[8][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][12]  ( .D(\Inst_Mem/inst_mem_reg[8][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[268]), .Q(
        \Inst_Mem/inst_mem_reg[8][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][13]  ( .D(\Inst_Mem/inst_mem_reg[8][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[269]), .Q(
        \Inst_Mem/inst_mem_reg[8][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][14]  ( .D(\Inst_Mem/inst_mem_reg[8][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[270]), .Q(
        \Inst_Mem/inst_mem_reg[8][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][15]  ( .D(\Inst_Mem/inst_mem_reg[8][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[271]), .Q(
        \Inst_Mem/inst_mem_reg[8][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][16]  ( .D(\Inst_Mem/inst_mem_reg[8][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[272]), .Q(
        \Inst_Mem/inst_mem_reg[8][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][17]  ( .D(\Inst_Mem/inst_mem_reg[8][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[273]), .Q(
        \Inst_Mem/inst_mem_reg[8][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][18]  ( .D(\Inst_Mem/inst_mem_reg[8][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[274]), .Q(
        \Inst_Mem/inst_mem_reg[8][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][19]  ( .D(\Inst_Mem/inst_mem_reg[8][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[275]), .Q(
        \Inst_Mem/inst_mem_reg[8][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][20]  ( .D(\Inst_Mem/inst_mem_reg[8][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[276]), .Q(
        \Inst_Mem/inst_mem_reg[8][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][21]  ( .D(\Inst_Mem/inst_mem_reg[8][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[277]), .Q(
        \Inst_Mem/inst_mem_reg[8][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][22]  ( .D(\Inst_Mem/inst_mem_reg[8][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[278]), .Q(
        \Inst_Mem/inst_mem_reg[8][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][23]  ( .D(\Inst_Mem/inst_mem_reg[8][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[279]), .Q(
        \Inst_Mem/inst_mem_reg[8][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][24]  ( .D(\Inst_Mem/inst_mem_reg[8][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[280]), .Q(
        \Inst_Mem/inst_mem_reg[8][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][25]  ( .D(\Inst_Mem/inst_mem_reg[8][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[281]), .Q(
        \Inst_Mem/inst_mem_reg[8][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][26]  ( .D(\Inst_Mem/inst_mem_reg[8][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[282]), .Q(
        \Inst_Mem/inst_mem_reg[8][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][27]  ( .D(\Inst_Mem/inst_mem_reg[8][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[283]), .Q(
        \Inst_Mem/inst_mem_reg[8][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][28]  ( .D(\Inst_Mem/inst_mem_reg[8][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[284]), .Q(
        \Inst_Mem/inst_mem_reg[8][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][29]  ( .D(\Inst_Mem/inst_mem_reg[8][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[285]), .Q(
        \Inst_Mem/inst_mem_reg[8][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][30]  ( .D(\Inst_Mem/inst_mem_reg[8][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[286]), .Q(
        \Inst_Mem/inst_mem_reg[8][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[8][31]  ( .D(\Inst_Mem/inst_mem_reg[8][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[287]), .Q(
        \Inst_Mem/inst_mem_reg[8][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][0]  ( .D(\Inst_Mem/inst_mem_reg[7][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[224]), .Q(
        \Inst_Mem/inst_mem_reg[7][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][1]  ( .D(\Inst_Mem/inst_mem_reg[7][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[225]), .Q(
        \Inst_Mem/inst_mem_reg[7][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][2]  ( .D(\Inst_Mem/inst_mem_reg[7][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[226]), .Q(
        \Inst_Mem/inst_mem_reg[7][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][3]  ( .D(\Inst_Mem/inst_mem_reg[7][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[227]), .Q(
        \Inst_Mem/inst_mem_reg[7][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][4]  ( .D(\Inst_Mem/inst_mem_reg[7][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[228]), .Q(
        \Inst_Mem/inst_mem_reg[7][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][5]  ( .D(\Inst_Mem/inst_mem_reg[7][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[229]), .Q(
        \Inst_Mem/inst_mem_reg[7][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][6]  ( .D(\Inst_Mem/inst_mem_reg[7][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[230]), .Q(
        \Inst_Mem/inst_mem_reg[7][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][7]  ( .D(\Inst_Mem/inst_mem_reg[7][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[231]), .Q(
        \Inst_Mem/inst_mem_reg[7][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][8]  ( .D(\Inst_Mem/inst_mem_reg[7][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[232]), .Q(
        \Inst_Mem/inst_mem_reg[7][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][9]  ( .D(\Inst_Mem/inst_mem_reg[7][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[233]), .Q(
        \Inst_Mem/inst_mem_reg[7][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][10]  ( .D(\Inst_Mem/inst_mem_reg[7][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[234]), .Q(
        \Inst_Mem/inst_mem_reg[7][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][11]  ( .D(\Inst_Mem/inst_mem_reg[7][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[235]), .Q(
        \Inst_Mem/inst_mem_reg[7][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][12]  ( .D(\Inst_Mem/inst_mem_reg[7][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[236]), .Q(
        \Inst_Mem/inst_mem_reg[7][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][13]  ( .D(\Inst_Mem/inst_mem_reg[7][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[237]), .Q(
        \Inst_Mem/inst_mem_reg[7][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][14]  ( .D(\Inst_Mem/inst_mem_reg[7][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[238]), .Q(
        \Inst_Mem/inst_mem_reg[7][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][15]  ( .D(\Inst_Mem/inst_mem_reg[7][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[239]), .Q(
        \Inst_Mem/inst_mem_reg[7][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][16]  ( .D(\Inst_Mem/inst_mem_reg[7][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[240]), .Q(
        \Inst_Mem/inst_mem_reg[7][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][17]  ( .D(\Inst_Mem/inst_mem_reg[7][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[241]), .Q(
        \Inst_Mem/inst_mem_reg[7][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][18]  ( .D(\Inst_Mem/inst_mem_reg[7][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[242]), .Q(
        \Inst_Mem/inst_mem_reg[7][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][19]  ( .D(\Inst_Mem/inst_mem_reg[7][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[243]), .Q(
        \Inst_Mem/inst_mem_reg[7][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][20]  ( .D(\Inst_Mem/inst_mem_reg[7][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[244]), .Q(
        \Inst_Mem/inst_mem_reg[7][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][21]  ( .D(\Inst_Mem/inst_mem_reg[7][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[245]), .Q(
        \Inst_Mem/inst_mem_reg[7][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][22]  ( .D(\Inst_Mem/inst_mem_reg[7][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[246]), .Q(
        \Inst_Mem/inst_mem_reg[7][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][23]  ( .D(\Inst_Mem/inst_mem_reg[7][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[247]), .Q(
        \Inst_Mem/inst_mem_reg[7][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][24]  ( .D(\Inst_Mem/inst_mem_reg[7][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[248]), .Q(
        \Inst_Mem/inst_mem_reg[7][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][25]  ( .D(\Inst_Mem/inst_mem_reg[7][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[249]), .Q(
        \Inst_Mem/inst_mem_reg[7][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][26]  ( .D(\Inst_Mem/inst_mem_reg[7][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[250]), .Q(
        \Inst_Mem/inst_mem_reg[7][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][27]  ( .D(\Inst_Mem/inst_mem_reg[7][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[251]), .Q(
        \Inst_Mem/inst_mem_reg[7][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][28]  ( .D(\Inst_Mem/inst_mem_reg[7][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[252]), .Q(
        \Inst_Mem/inst_mem_reg[7][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][29]  ( .D(\Inst_Mem/inst_mem_reg[7][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[253]), .Q(
        \Inst_Mem/inst_mem_reg[7][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][30]  ( .D(\Inst_Mem/inst_mem_reg[7][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[254]), .Q(
        \Inst_Mem/inst_mem_reg[7][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[7][31]  ( .D(\Inst_Mem/inst_mem_reg[7][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[255]), .Q(
        \Inst_Mem/inst_mem_reg[7][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][0]  ( .D(\Inst_Mem/inst_mem_reg[6][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[192]), .Q(
        \Inst_Mem/inst_mem_reg[6][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][1]  ( .D(\Inst_Mem/inst_mem_reg[6][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[193]), .Q(
        \Inst_Mem/inst_mem_reg[6][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][2]  ( .D(\Inst_Mem/inst_mem_reg[6][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[194]), .Q(
        \Inst_Mem/inst_mem_reg[6][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][3]  ( .D(\Inst_Mem/inst_mem_reg[6][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[195]), .Q(
        \Inst_Mem/inst_mem_reg[6][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][4]  ( .D(\Inst_Mem/inst_mem_reg[6][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[196]), .Q(
        \Inst_Mem/inst_mem_reg[6][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][5]  ( .D(\Inst_Mem/inst_mem_reg[6][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[197]), .Q(
        \Inst_Mem/inst_mem_reg[6][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][6]  ( .D(\Inst_Mem/inst_mem_reg[6][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[198]), .Q(
        \Inst_Mem/inst_mem_reg[6][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][7]  ( .D(\Inst_Mem/inst_mem_reg[6][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[199]), .Q(
        \Inst_Mem/inst_mem_reg[6][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][8]  ( .D(\Inst_Mem/inst_mem_reg[6][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[200]), .Q(
        \Inst_Mem/inst_mem_reg[6][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][9]  ( .D(\Inst_Mem/inst_mem_reg[6][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[201]), .Q(
        \Inst_Mem/inst_mem_reg[6][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][10]  ( .D(\Inst_Mem/inst_mem_reg[6][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[202]), .Q(
        \Inst_Mem/inst_mem_reg[6][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][11]  ( .D(\Inst_Mem/inst_mem_reg[6][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[203]), .Q(
        \Inst_Mem/inst_mem_reg[6][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][12]  ( .D(\Inst_Mem/inst_mem_reg[6][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[204]), .Q(
        \Inst_Mem/inst_mem_reg[6][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][13]  ( .D(\Inst_Mem/inst_mem_reg[6][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[205]), .Q(
        \Inst_Mem/inst_mem_reg[6][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][14]  ( .D(\Inst_Mem/inst_mem_reg[6][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[206]), .Q(
        \Inst_Mem/inst_mem_reg[6][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][15]  ( .D(\Inst_Mem/inst_mem_reg[6][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[207]), .Q(
        \Inst_Mem/inst_mem_reg[6][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][16]  ( .D(\Inst_Mem/inst_mem_reg[6][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[208]), .Q(
        \Inst_Mem/inst_mem_reg[6][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][17]  ( .D(\Inst_Mem/inst_mem_reg[6][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[209]), .Q(
        \Inst_Mem/inst_mem_reg[6][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][18]  ( .D(\Inst_Mem/inst_mem_reg[6][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[210]), .Q(
        \Inst_Mem/inst_mem_reg[6][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][19]  ( .D(\Inst_Mem/inst_mem_reg[6][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[211]), .Q(
        \Inst_Mem/inst_mem_reg[6][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][20]  ( .D(\Inst_Mem/inst_mem_reg[6][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[212]), .Q(
        \Inst_Mem/inst_mem_reg[6][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][21]  ( .D(\Inst_Mem/inst_mem_reg[6][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[213]), .Q(
        \Inst_Mem/inst_mem_reg[6][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][22]  ( .D(\Inst_Mem/inst_mem_reg[6][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[214]), .Q(
        \Inst_Mem/inst_mem_reg[6][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][23]  ( .D(\Inst_Mem/inst_mem_reg[6][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[215]), .Q(
        \Inst_Mem/inst_mem_reg[6][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][24]  ( .D(\Inst_Mem/inst_mem_reg[6][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[216]), .Q(
        \Inst_Mem/inst_mem_reg[6][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][25]  ( .D(\Inst_Mem/inst_mem_reg[6][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[217]), .Q(
        \Inst_Mem/inst_mem_reg[6][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][26]  ( .D(\Inst_Mem/inst_mem_reg[6][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[218]), .Q(
        \Inst_Mem/inst_mem_reg[6][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][27]  ( .D(\Inst_Mem/inst_mem_reg[6][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[219]), .Q(
        \Inst_Mem/inst_mem_reg[6][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][28]  ( .D(\Inst_Mem/inst_mem_reg[6][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[220]), .Q(
        \Inst_Mem/inst_mem_reg[6][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][29]  ( .D(\Inst_Mem/inst_mem_reg[6][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[221]), .Q(
        \Inst_Mem/inst_mem_reg[6][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][30]  ( .D(\Inst_Mem/inst_mem_reg[6][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[222]), .Q(
        \Inst_Mem/inst_mem_reg[6][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[6][31]  ( .D(\Inst_Mem/inst_mem_reg[6][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[223]), .Q(
        \Inst_Mem/inst_mem_reg[6][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][0]  ( .D(\Inst_Mem/inst_mem_reg[5][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[160]), .Q(
        \Inst_Mem/inst_mem_reg[5][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][1]  ( .D(\Inst_Mem/inst_mem_reg[5][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[161]), .Q(
        \Inst_Mem/inst_mem_reg[5][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][2]  ( .D(\Inst_Mem/inst_mem_reg[5][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[162]), .Q(
        \Inst_Mem/inst_mem_reg[5][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][3]  ( .D(\Inst_Mem/inst_mem_reg[5][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[163]), .Q(
        \Inst_Mem/inst_mem_reg[5][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][4]  ( .D(\Inst_Mem/inst_mem_reg[5][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[164]), .Q(
        \Inst_Mem/inst_mem_reg[5][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][5]  ( .D(\Inst_Mem/inst_mem_reg[5][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[165]), .Q(
        \Inst_Mem/inst_mem_reg[5][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][6]  ( .D(\Inst_Mem/inst_mem_reg[5][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[166]), .Q(
        \Inst_Mem/inst_mem_reg[5][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][7]  ( .D(\Inst_Mem/inst_mem_reg[5][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[167]), .Q(
        \Inst_Mem/inst_mem_reg[5][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][8]  ( .D(\Inst_Mem/inst_mem_reg[5][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[168]), .Q(
        \Inst_Mem/inst_mem_reg[5][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][9]  ( .D(\Inst_Mem/inst_mem_reg[5][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[169]), .Q(
        \Inst_Mem/inst_mem_reg[5][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][10]  ( .D(\Inst_Mem/inst_mem_reg[5][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[170]), .Q(
        \Inst_Mem/inst_mem_reg[5][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][11]  ( .D(\Inst_Mem/inst_mem_reg[5][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[171]), .Q(
        \Inst_Mem/inst_mem_reg[5][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][12]  ( .D(\Inst_Mem/inst_mem_reg[5][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[172]), .Q(
        \Inst_Mem/inst_mem_reg[5][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][13]  ( .D(\Inst_Mem/inst_mem_reg[5][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[173]), .Q(
        \Inst_Mem/inst_mem_reg[5][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][14]  ( .D(\Inst_Mem/inst_mem_reg[5][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[174]), .Q(
        \Inst_Mem/inst_mem_reg[5][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][15]  ( .D(\Inst_Mem/inst_mem_reg[5][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[175]), .Q(
        \Inst_Mem/inst_mem_reg[5][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][16]  ( .D(\Inst_Mem/inst_mem_reg[5][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[176]), .Q(
        \Inst_Mem/inst_mem_reg[5][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][17]  ( .D(\Inst_Mem/inst_mem_reg[5][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[177]), .Q(
        \Inst_Mem/inst_mem_reg[5][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][18]  ( .D(\Inst_Mem/inst_mem_reg[5][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[178]), .Q(
        \Inst_Mem/inst_mem_reg[5][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][19]  ( .D(\Inst_Mem/inst_mem_reg[5][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[179]), .Q(
        \Inst_Mem/inst_mem_reg[5][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][20]  ( .D(\Inst_Mem/inst_mem_reg[5][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[180]), .Q(
        \Inst_Mem/inst_mem_reg[5][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][21]  ( .D(\Inst_Mem/inst_mem_reg[5][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[181]), .Q(
        \Inst_Mem/inst_mem_reg[5][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][22]  ( .D(\Inst_Mem/inst_mem_reg[5][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[182]), .Q(
        \Inst_Mem/inst_mem_reg[5][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][23]  ( .D(\Inst_Mem/inst_mem_reg[5][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[183]), .Q(
        \Inst_Mem/inst_mem_reg[5][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][24]  ( .D(\Inst_Mem/inst_mem_reg[5][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[184]), .Q(
        \Inst_Mem/inst_mem_reg[5][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][25]  ( .D(\Inst_Mem/inst_mem_reg[5][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[185]), .Q(
        \Inst_Mem/inst_mem_reg[5][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][26]  ( .D(\Inst_Mem/inst_mem_reg[5][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[186]), .Q(
        \Inst_Mem/inst_mem_reg[5][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][27]  ( .D(\Inst_Mem/inst_mem_reg[5][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[187]), .Q(
        \Inst_Mem/inst_mem_reg[5][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][28]  ( .D(\Inst_Mem/inst_mem_reg[5][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[188]), .Q(
        \Inst_Mem/inst_mem_reg[5][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][29]  ( .D(\Inst_Mem/inst_mem_reg[5][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[189]), .Q(
        \Inst_Mem/inst_mem_reg[5][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][30]  ( .D(\Inst_Mem/inst_mem_reg[5][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[190]), .Q(
        \Inst_Mem/inst_mem_reg[5][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[5][31]  ( .D(\Inst_Mem/inst_mem_reg[5][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[191]), .Q(
        \Inst_Mem/inst_mem_reg[5][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][0]  ( .D(\Inst_Mem/inst_mem_reg[4][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[128]), .Q(
        \Inst_Mem/inst_mem_reg[4][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][1]  ( .D(\Inst_Mem/inst_mem_reg[4][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[129]), .Q(
        \Inst_Mem/inst_mem_reg[4][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][2]  ( .D(\Inst_Mem/inst_mem_reg[4][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[130]), .Q(
        \Inst_Mem/inst_mem_reg[4][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][3]  ( .D(\Inst_Mem/inst_mem_reg[4][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[131]), .Q(
        \Inst_Mem/inst_mem_reg[4][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][4]  ( .D(\Inst_Mem/inst_mem_reg[4][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[132]), .Q(
        \Inst_Mem/inst_mem_reg[4][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][5]  ( .D(\Inst_Mem/inst_mem_reg[4][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[133]), .Q(
        \Inst_Mem/inst_mem_reg[4][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][6]  ( .D(\Inst_Mem/inst_mem_reg[4][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[134]), .Q(
        \Inst_Mem/inst_mem_reg[4][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][7]  ( .D(\Inst_Mem/inst_mem_reg[4][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[135]), .Q(
        \Inst_Mem/inst_mem_reg[4][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][8]  ( .D(\Inst_Mem/inst_mem_reg[4][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[136]), .Q(
        \Inst_Mem/inst_mem_reg[4][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][9]  ( .D(\Inst_Mem/inst_mem_reg[4][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[137]), .Q(
        \Inst_Mem/inst_mem_reg[4][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][10]  ( .D(\Inst_Mem/inst_mem_reg[4][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[138]), .Q(
        \Inst_Mem/inst_mem_reg[4][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][11]  ( .D(\Inst_Mem/inst_mem_reg[4][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[139]), .Q(
        \Inst_Mem/inst_mem_reg[4][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][12]  ( .D(\Inst_Mem/inst_mem_reg[4][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[140]), .Q(
        \Inst_Mem/inst_mem_reg[4][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][13]  ( .D(\Inst_Mem/inst_mem_reg[4][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[141]), .Q(
        \Inst_Mem/inst_mem_reg[4][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][14]  ( .D(\Inst_Mem/inst_mem_reg[4][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[142]), .Q(
        \Inst_Mem/inst_mem_reg[4][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][15]  ( .D(\Inst_Mem/inst_mem_reg[4][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[143]), .Q(
        \Inst_Mem/inst_mem_reg[4][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][16]  ( .D(\Inst_Mem/inst_mem_reg[4][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[144]), .Q(
        \Inst_Mem/inst_mem_reg[4][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][17]  ( .D(\Inst_Mem/inst_mem_reg[4][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[145]), .Q(
        \Inst_Mem/inst_mem_reg[4][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][18]  ( .D(\Inst_Mem/inst_mem_reg[4][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[146]), .Q(
        \Inst_Mem/inst_mem_reg[4][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][19]  ( .D(\Inst_Mem/inst_mem_reg[4][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[147]), .Q(
        \Inst_Mem/inst_mem_reg[4][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][20]  ( .D(\Inst_Mem/inst_mem_reg[4][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[148]), .Q(
        \Inst_Mem/inst_mem_reg[4][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][21]  ( .D(\Inst_Mem/inst_mem_reg[4][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[149]), .Q(
        \Inst_Mem/inst_mem_reg[4][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][22]  ( .D(\Inst_Mem/inst_mem_reg[4][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[150]), .Q(
        \Inst_Mem/inst_mem_reg[4][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][23]  ( .D(\Inst_Mem/inst_mem_reg[4][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[151]), .Q(
        \Inst_Mem/inst_mem_reg[4][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][24]  ( .D(\Inst_Mem/inst_mem_reg[4][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[152]), .Q(
        \Inst_Mem/inst_mem_reg[4][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][25]  ( .D(\Inst_Mem/inst_mem_reg[4][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[153]), .Q(
        \Inst_Mem/inst_mem_reg[4][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][26]  ( .D(\Inst_Mem/inst_mem_reg[4][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[154]), .Q(
        \Inst_Mem/inst_mem_reg[4][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][27]  ( .D(\Inst_Mem/inst_mem_reg[4][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[155]), .Q(
        \Inst_Mem/inst_mem_reg[4][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][28]  ( .D(\Inst_Mem/inst_mem_reg[4][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[156]), .Q(
        \Inst_Mem/inst_mem_reg[4][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][29]  ( .D(\Inst_Mem/inst_mem_reg[4][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[157]), .Q(
        \Inst_Mem/inst_mem_reg[4][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][30]  ( .D(\Inst_Mem/inst_mem_reg[4][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[158]), .Q(
        \Inst_Mem/inst_mem_reg[4][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[4][31]  ( .D(\Inst_Mem/inst_mem_reg[4][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[159]), .Q(
        \Inst_Mem/inst_mem_reg[4][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][0]  ( .D(\Inst_Mem/inst_mem_reg[3][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[96]), .Q(\Inst_Mem/inst_mem_reg[3][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][1]  ( .D(\Inst_Mem/inst_mem_reg[3][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[97]), .Q(\Inst_Mem/inst_mem_reg[3][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][2]  ( .D(\Inst_Mem/inst_mem_reg[3][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[98]), .Q(\Inst_Mem/inst_mem_reg[3][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][3]  ( .D(\Inst_Mem/inst_mem_reg[3][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[99]), .Q(\Inst_Mem/inst_mem_reg[3][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][4]  ( .D(\Inst_Mem/inst_mem_reg[3][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[100]), .Q(
        \Inst_Mem/inst_mem_reg[3][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][5]  ( .D(\Inst_Mem/inst_mem_reg[3][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[101]), .Q(
        \Inst_Mem/inst_mem_reg[3][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][6]  ( .D(\Inst_Mem/inst_mem_reg[3][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[102]), .Q(
        \Inst_Mem/inst_mem_reg[3][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][7]  ( .D(\Inst_Mem/inst_mem_reg[3][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[103]), .Q(
        \Inst_Mem/inst_mem_reg[3][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][8]  ( .D(\Inst_Mem/inst_mem_reg[3][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[104]), .Q(
        \Inst_Mem/inst_mem_reg[3][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][9]  ( .D(\Inst_Mem/inst_mem_reg[3][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[105]), .Q(
        \Inst_Mem/inst_mem_reg[3][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][10]  ( .D(\Inst_Mem/inst_mem_reg[3][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[106]), .Q(
        \Inst_Mem/inst_mem_reg[3][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][11]  ( .D(\Inst_Mem/inst_mem_reg[3][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[107]), .Q(
        \Inst_Mem/inst_mem_reg[3][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][12]  ( .D(\Inst_Mem/inst_mem_reg[3][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[108]), .Q(
        \Inst_Mem/inst_mem_reg[3][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][13]  ( .D(\Inst_Mem/inst_mem_reg[3][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[109]), .Q(
        \Inst_Mem/inst_mem_reg[3][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][14]  ( .D(\Inst_Mem/inst_mem_reg[3][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[110]), .Q(
        \Inst_Mem/inst_mem_reg[3][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][15]  ( .D(\Inst_Mem/inst_mem_reg[3][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[111]), .Q(
        \Inst_Mem/inst_mem_reg[3][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][16]  ( .D(\Inst_Mem/inst_mem_reg[3][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[112]), .Q(
        \Inst_Mem/inst_mem_reg[3][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][17]  ( .D(\Inst_Mem/inst_mem_reg[3][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[113]), .Q(
        \Inst_Mem/inst_mem_reg[3][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][18]  ( .D(\Inst_Mem/inst_mem_reg[3][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[114]), .Q(
        \Inst_Mem/inst_mem_reg[3][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][19]  ( .D(\Inst_Mem/inst_mem_reg[3][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[115]), .Q(
        \Inst_Mem/inst_mem_reg[3][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][20]  ( .D(\Inst_Mem/inst_mem_reg[3][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[116]), .Q(
        \Inst_Mem/inst_mem_reg[3][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][21]  ( .D(\Inst_Mem/inst_mem_reg[3][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[117]), .Q(
        \Inst_Mem/inst_mem_reg[3][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][22]  ( .D(\Inst_Mem/inst_mem_reg[3][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[118]), .Q(
        \Inst_Mem/inst_mem_reg[3][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][23]  ( .D(\Inst_Mem/inst_mem_reg[3][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[119]), .Q(
        \Inst_Mem/inst_mem_reg[3][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][24]  ( .D(\Inst_Mem/inst_mem_reg[3][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[120]), .Q(
        \Inst_Mem/inst_mem_reg[3][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][25]  ( .D(\Inst_Mem/inst_mem_reg[3][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[121]), .Q(
        \Inst_Mem/inst_mem_reg[3][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][26]  ( .D(\Inst_Mem/inst_mem_reg[3][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[122]), .Q(
        \Inst_Mem/inst_mem_reg[3][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][27]  ( .D(\Inst_Mem/inst_mem_reg[3][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[123]), .Q(
        \Inst_Mem/inst_mem_reg[3][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][28]  ( .D(\Inst_Mem/inst_mem_reg[3][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[124]), .Q(
        \Inst_Mem/inst_mem_reg[3][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][29]  ( .D(\Inst_Mem/inst_mem_reg[3][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[125]), .Q(
        \Inst_Mem/inst_mem_reg[3][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][30]  ( .D(\Inst_Mem/inst_mem_reg[3][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[126]), .Q(
        \Inst_Mem/inst_mem_reg[3][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[3][31]  ( .D(\Inst_Mem/inst_mem_reg[3][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[127]), .Q(
        \Inst_Mem/inst_mem_reg[3][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][0]  ( .D(\Inst_Mem/inst_mem_reg[2][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[64]), .Q(\Inst_Mem/inst_mem_reg[2][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][1]  ( .D(\Inst_Mem/inst_mem_reg[2][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[65]), .Q(\Inst_Mem/inst_mem_reg[2][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][2]  ( .D(\Inst_Mem/inst_mem_reg[2][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[66]), .Q(\Inst_Mem/inst_mem_reg[2][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][3]  ( .D(\Inst_Mem/inst_mem_reg[2][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[67]), .Q(\Inst_Mem/inst_mem_reg[2][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][4]  ( .D(\Inst_Mem/inst_mem_reg[2][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[68]), .Q(\Inst_Mem/inst_mem_reg[2][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][5]  ( .D(\Inst_Mem/inst_mem_reg[2][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[69]), .Q(\Inst_Mem/inst_mem_reg[2][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][6]  ( .D(\Inst_Mem/inst_mem_reg[2][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[70]), .Q(\Inst_Mem/inst_mem_reg[2][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][7]  ( .D(\Inst_Mem/inst_mem_reg[2][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[71]), .Q(\Inst_Mem/inst_mem_reg[2][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][8]  ( .D(\Inst_Mem/inst_mem_reg[2][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[72]), .Q(\Inst_Mem/inst_mem_reg[2][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][9]  ( .D(\Inst_Mem/inst_mem_reg[2][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[73]), .Q(\Inst_Mem/inst_mem_reg[2][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][10]  ( .D(\Inst_Mem/inst_mem_reg[2][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[74]), .Q(
        \Inst_Mem/inst_mem_reg[2][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][11]  ( .D(\Inst_Mem/inst_mem_reg[2][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[75]), .Q(
        \Inst_Mem/inst_mem_reg[2][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][12]  ( .D(\Inst_Mem/inst_mem_reg[2][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[76]), .Q(
        \Inst_Mem/inst_mem_reg[2][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][13]  ( .D(\Inst_Mem/inst_mem_reg[2][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[77]), .Q(
        \Inst_Mem/inst_mem_reg[2][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][14]  ( .D(\Inst_Mem/inst_mem_reg[2][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[78]), .Q(
        \Inst_Mem/inst_mem_reg[2][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][15]  ( .D(\Inst_Mem/inst_mem_reg[2][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[79]), .Q(
        \Inst_Mem/inst_mem_reg[2][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][16]  ( .D(\Inst_Mem/inst_mem_reg[2][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[80]), .Q(
        \Inst_Mem/inst_mem_reg[2][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][17]  ( .D(\Inst_Mem/inst_mem_reg[2][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[81]), .Q(
        \Inst_Mem/inst_mem_reg[2][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][18]  ( .D(\Inst_Mem/inst_mem_reg[2][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[82]), .Q(
        \Inst_Mem/inst_mem_reg[2][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][19]  ( .D(\Inst_Mem/inst_mem_reg[2][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[83]), .Q(
        \Inst_Mem/inst_mem_reg[2][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][20]  ( .D(\Inst_Mem/inst_mem_reg[2][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[84]), .Q(
        \Inst_Mem/inst_mem_reg[2][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][21]  ( .D(\Inst_Mem/inst_mem_reg[2][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[85]), .Q(
        \Inst_Mem/inst_mem_reg[2][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][22]  ( .D(\Inst_Mem/inst_mem_reg[2][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[86]), .Q(
        \Inst_Mem/inst_mem_reg[2][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][23]  ( .D(\Inst_Mem/inst_mem_reg[2][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[87]), .Q(
        \Inst_Mem/inst_mem_reg[2][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][24]  ( .D(\Inst_Mem/inst_mem_reg[2][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[88]), .Q(
        \Inst_Mem/inst_mem_reg[2][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][25]  ( .D(\Inst_Mem/inst_mem_reg[2][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[89]), .Q(
        \Inst_Mem/inst_mem_reg[2][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][26]  ( .D(\Inst_Mem/inst_mem_reg[2][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[90]), .Q(
        \Inst_Mem/inst_mem_reg[2][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][27]  ( .D(\Inst_Mem/inst_mem_reg[2][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[91]), .Q(
        \Inst_Mem/inst_mem_reg[2][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][28]  ( .D(\Inst_Mem/inst_mem_reg[2][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[92]), .Q(
        \Inst_Mem/inst_mem_reg[2][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][29]  ( .D(\Inst_Mem/inst_mem_reg[2][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[93]), .Q(
        \Inst_Mem/inst_mem_reg[2][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][30]  ( .D(\Inst_Mem/inst_mem_reg[2][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[94]), .Q(
        \Inst_Mem/inst_mem_reg[2][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[2][31]  ( .D(\Inst_Mem/inst_mem_reg[2][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[95]), .Q(
        \Inst_Mem/inst_mem_reg[2][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][0]  ( .D(\Inst_Mem/inst_mem_reg[1][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[32]), .Q(\Inst_Mem/inst_mem_reg[1][0] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][1]  ( .D(\Inst_Mem/inst_mem_reg[1][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[33]), .Q(\Inst_Mem/inst_mem_reg[1][1] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][2]  ( .D(\Inst_Mem/inst_mem_reg[1][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[34]), .Q(\Inst_Mem/inst_mem_reg[1][2] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][3]  ( .D(\Inst_Mem/inst_mem_reg[1][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[35]), .Q(\Inst_Mem/inst_mem_reg[1][3] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][4]  ( .D(\Inst_Mem/inst_mem_reg[1][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[36]), .Q(\Inst_Mem/inst_mem_reg[1][4] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][5]  ( .D(\Inst_Mem/inst_mem_reg[1][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[37]), .Q(\Inst_Mem/inst_mem_reg[1][5] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][6]  ( .D(\Inst_Mem/inst_mem_reg[1][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[38]), .Q(\Inst_Mem/inst_mem_reg[1][6] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][7]  ( .D(\Inst_Mem/inst_mem_reg[1][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[39]), .Q(\Inst_Mem/inst_mem_reg[1][7] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][8]  ( .D(\Inst_Mem/inst_mem_reg[1][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[40]), .Q(\Inst_Mem/inst_mem_reg[1][8] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][9]  ( .D(\Inst_Mem/inst_mem_reg[1][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[41]), .Q(\Inst_Mem/inst_mem_reg[1][9] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][10]  ( .D(\Inst_Mem/inst_mem_reg[1][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[42]), .Q(
        \Inst_Mem/inst_mem_reg[1][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][11]  ( .D(\Inst_Mem/inst_mem_reg[1][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[43]), .Q(
        \Inst_Mem/inst_mem_reg[1][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][12]  ( .D(\Inst_Mem/inst_mem_reg[1][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[44]), .Q(
        \Inst_Mem/inst_mem_reg[1][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][13]  ( .D(\Inst_Mem/inst_mem_reg[1][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[45]), .Q(
        \Inst_Mem/inst_mem_reg[1][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][14]  ( .D(\Inst_Mem/inst_mem_reg[1][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[46]), .Q(
        \Inst_Mem/inst_mem_reg[1][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][15]  ( .D(\Inst_Mem/inst_mem_reg[1][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[47]), .Q(
        \Inst_Mem/inst_mem_reg[1][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][16]  ( .D(\Inst_Mem/inst_mem_reg[1][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[48]), .Q(
        \Inst_Mem/inst_mem_reg[1][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][17]  ( .D(\Inst_Mem/inst_mem_reg[1][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[49]), .Q(
        \Inst_Mem/inst_mem_reg[1][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][18]  ( .D(\Inst_Mem/inst_mem_reg[1][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[50]), .Q(
        \Inst_Mem/inst_mem_reg[1][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][19]  ( .D(\Inst_Mem/inst_mem_reg[1][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[51]), .Q(
        \Inst_Mem/inst_mem_reg[1][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][20]  ( .D(\Inst_Mem/inst_mem_reg[1][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[52]), .Q(
        \Inst_Mem/inst_mem_reg[1][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][21]  ( .D(\Inst_Mem/inst_mem_reg[1][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[53]), .Q(
        \Inst_Mem/inst_mem_reg[1][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][22]  ( .D(\Inst_Mem/inst_mem_reg[1][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[54]), .Q(
        \Inst_Mem/inst_mem_reg[1][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][23]  ( .D(\Inst_Mem/inst_mem_reg[1][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[55]), .Q(
        \Inst_Mem/inst_mem_reg[1][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][24]  ( .D(\Inst_Mem/inst_mem_reg[1][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[56]), .Q(
        \Inst_Mem/inst_mem_reg[1][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][25]  ( .D(\Inst_Mem/inst_mem_reg[1][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[57]), .Q(
        \Inst_Mem/inst_mem_reg[1][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][26]  ( .D(\Inst_Mem/inst_mem_reg[1][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[58]), .Q(
        \Inst_Mem/inst_mem_reg[1][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][27]  ( .D(\Inst_Mem/inst_mem_reg[1][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[59]), .Q(
        \Inst_Mem/inst_mem_reg[1][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][28]  ( .D(\Inst_Mem/inst_mem_reg[1][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[60]), .Q(
        \Inst_Mem/inst_mem_reg[1][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][29]  ( .D(\Inst_Mem/inst_mem_reg[1][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[61]), .Q(
        \Inst_Mem/inst_mem_reg[1][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][30]  ( .D(\Inst_Mem/inst_mem_reg[1][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[62]), .Q(
        \Inst_Mem/inst_mem_reg[1][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[1][31]  ( .D(\Inst_Mem/inst_mem_reg[1][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[63]), .Q(
        \Inst_Mem/inst_mem_reg[1][31] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][0]  ( .D(\Inst_Mem/inst_mem_reg[0][0] ), 
        .CLK(clk), .RST(rst), .I(g_init[0]), .Q(\Inst_Mem/inst_mem_reg[0][0] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][1]  ( .D(\Inst_Mem/inst_mem_reg[0][1] ), 
        .CLK(clk), .RST(rst), .I(g_init[1]), .Q(\Inst_Mem/inst_mem_reg[0][1] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][2]  ( .D(\Inst_Mem/inst_mem_reg[0][2] ), 
        .CLK(clk), .RST(rst), .I(g_init[2]), .Q(\Inst_Mem/inst_mem_reg[0][2] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][3]  ( .D(\Inst_Mem/inst_mem_reg[0][3] ), 
        .CLK(clk), .RST(rst), .I(g_init[3]), .Q(\Inst_Mem/inst_mem_reg[0][3] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][4]  ( .D(\Inst_Mem/inst_mem_reg[0][4] ), 
        .CLK(clk), .RST(rst), .I(g_init[4]), .Q(\Inst_Mem/inst_mem_reg[0][4] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][5]  ( .D(\Inst_Mem/inst_mem_reg[0][5] ), 
        .CLK(clk), .RST(rst), .I(g_init[5]), .Q(\Inst_Mem/inst_mem_reg[0][5] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][6]  ( .D(\Inst_Mem/inst_mem_reg[0][6] ), 
        .CLK(clk), .RST(rst), .I(g_init[6]), .Q(\Inst_Mem/inst_mem_reg[0][6] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][7]  ( .D(\Inst_Mem/inst_mem_reg[0][7] ), 
        .CLK(clk), .RST(rst), .I(g_init[7]), .Q(\Inst_Mem/inst_mem_reg[0][7] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][8]  ( .D(\Inst_Mem/inst_mem_reg[0][8] ), 
        .CLK(clk), .RST(rst), .I(g_init[8]), .Q(\Inst_Mem/inst_mem_reg[0][8] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][9]  ( .D(\Inst_Mem/inst_mem_reg[0][9] ), 
        .CLK(clk), .RST(rst), .I(g_init[9]), .Q(\Inst_Mem/inst_mem_reg[0][9] )
         );
  DFF \Inst_Mem/inst_mem_reg_reg[0][10]  ( .D(\Inst_Mem/inst_mem_reg[0][10] ), 
        .CLK(clk), .RST(rst), .I(g_init[10]), .Q(
        \Inst_Mem/inst_mem_reg[0][10] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][11]  ( .D(\Inst_Mem/inst_mem_reg[0][11] ), 
        .CLK(clk), .RST(rst), .I(g_init[11]), .Q(
        \Inst_Mem/inst_mem_reg[0][11] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][12]  ( .D(\Inst_Mem/inst_mem_reg[0][12] ), 
        .CLK(clk), .RST(rst), .I(g_init[12]), .Q(
        \Inst_Mem/inst_mem_reg[0][12] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][13]  ( .D(\Inst_Mem/inst_mem_reg[0][13] ), 
        .CLK(clk), .RST(rst), .I(g_init[13]), .Q(
        \Inst_Mem/inst_mem_reg[0][13] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][14]  ( .D(\Inst_Mem/inst_mem_reg[0][14] ), 
        .CLK(clk), .RST(rst), .I(g_init[14]), .Q(
        \Inst_Mem/inst_mem_reg[0][14] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][15]  ( .D(\Inst_Mem/inst_mem_reg[0][15] ), 
        .CLK(clk), .RST(rst), .I(g_init[15]), .Q(
        \Inst_Mem/inst_mem_reg[0][15] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][16]  ( .D(\Inst_Mem/inst_mem_reg[0][16] ), 
        .CLK(clk), .RST(rst), .I(g_init[16]), .Q(
        \Inst_Mem/inst_mem_reg[0][16] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][17]  ( .D(\Inst_Mem/inst_mem_reg[0][17] ), 
        .CLK(clk), .RST(rst), .I(g_init[17]), .Q(
        \Inst_Mem/inst_mem_reg[0][17] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][18]  ( .D(\Inst_Mem/inst_mem_reg[0][18] ), 
        .CLK(clk), .RST(rst), .I(g_init[18]), .Q(
        \Inst_Mem/inst_mem_reg[0][18] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][19]  ( .D(\Inst_Mem/inst_mem_reg[0][19] ), 
        .CLK(clk), .RST(rst), .I(g_init[19]), .Q(
        \Inst_Mem/inst_mem_reg[0][19] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][20]  ( .D(\Inst_Mem/inst_mem_reg[0][20] ), 
        .CLK(clk), .RST(rst), .I(g_init[20]), .Q(
        \Inst_Mem/inst_mem_reg[0][20] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][21]  ( .D(\Inst_Mem/inst_mem_reg[0][21] ), 
        .CLK(clk), .RST(rst), .I(g_init[21]), .Q(
        \Inst_Mem/inst_mem_reg[0][21] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][22]  ( .D(\Inst_Mem/inst_mem_reg[0][22] ), 
        .CLK(clk), .RST(rst), .I(g_init[22]), .Q(
        \Inst_Mem/inst_mem_reg[0][22] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][23]  ( .D(\Inst_Mem/inst_mem_reg[0][23] ), 
        .CLK(clk), .RST(rst), .I(g_init[23]), .Q(
        \Inst_Mem/inst_mem_reg[0][23] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][24]  ( .D(\Inst_Mem/inst_mem_reg[0][24] ), 
        .CLK(clk), .RST(rst), .I(g_init[24]), .Q(
        \Inst_Mem/inst_mem_reg[0][24] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][25]  ( .D(\Inst_Mem/inst_mem_reg[0][25] ), 
        .CLK(clk), .RST(rst), .I(g_init[25]), .Q(
        \Inst_Mem/inst_mem_reg[0][25] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][26]  ( .D(\Inst_Mem/inst_mem_reg[0][26] ), 
        .CLK(clk), .RST(rst), .I(g_init[26]), .Q(
        \Inst_Mem/inst_mem_reg[0][26] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][27]  ( .D(\Inst_Mem/inst_mem_reg[0][27] ), 
        .CLK(clk), .RST(rst), .I(g_init[27]), .Q(
        \Inst_Mem/inst_mem_reg[0][27] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][28]  ( .D(\Inst_Mem/inst_mem_reg[0][28] ), 
        .CLK(clk), .RST(rst), .I(g_init[28]), .Q(
        \Inst_Mem/inst_mem_reg[0][28] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][29]  ( .D(\Inst_Mem/inst_mem_reg[0][29] ), 
        .CLK(clk), .RST(rst), .I(g_init[29]), .Q(
        \Inst_Mem/inst_mem_reg[0][29] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][30]  ( .D(\Inst_Mem/inst_mem_reg[0][30] ), 
        .CLK(clk), .RST(rst), .I(g_init[30]), .Q(
        \Inst_Mem/inst_mem_reg[0][30] ) );
  DFF \Inst_Mem/inst_mem_reg_reg[0][31]  ( .D(\Inst_Mem/inst_mem_reg[0][31] ), 
        .CLK(clk), .RST(rst), .I(g_init[31]), .Q(
        \Inst_Mem/inst_mem_reg[0][31] ) );
  MUX \Data_Mem/U9809  ( .IN0(\Data_Mem/n9744 ), .IN1(\Data_Mem/n9713 ), .SEL(
        N24), .F(\Data_Mem/N714 ) );
  MUX \Data_Mem/U9808  ( .IN0(\Data_Mem/n9743 ), .IN1(\Data_Mem/n9728 ), .SEL(
        N25), .F(\Data_Mem/n9744 ) );
  MUX \Data_Mem/U9807  ( .IN0(\Data_Mem/n9742 ), .IN1(\Data_Mem/n9735 ), .SEL(
        N26), .F(\Data_Mem/n9743 ) );
  MUX \Data_Mem/U9806  ( .IN0(\Data_Mem/n9741 ), .IN1(\Data_Mem/n9738 ), .SEL(
        N27), .F(\Data_Mem/n9742 ) );
  MUX \Data_Mem/U9805  ( .IN0(\Data_Mem/n9740 ), .IN1(\Data_Mem/n9739 ), .SEL(
        N28), .F(\Data_Mem/n9741 ) );
  MUX \Data_Mem/U9804  ( .IN0(o[31]), .IN1(o[63]), .SEL(N29), .F(
        \Data_Mem/n9740 ) );
  MUX \Data_Mem/U9803  ( .IN0(o[95]), .IN1(o[127]), .SEL(N29), .F(
        \Data_Mem/n9739 ) );
  MUX \Data_Mem/U9802  ( .IN0(\Data_Mem/n9737 ), .IN1(\Data_Mem/n9736 ), .SEL(
        N28), .F(\Data_Mem/n9738 ) );
  MUX \Data_Mem/U9801  ( .IN0(o[159]), .IN1(o[191]), .SEL(N29), .F(
        \Data_Mem/n9737 ) );
  MUX \Data_Mem/U9800  ( .IN0(o[223]), .IN1(o[255]), .SEL(N29), .F(
        \Data_Mem/n9736 ) );
  MUX \Data_Mem/U9799  ( .IN0(\Data_Mem/n9734 ), .IN1(\Data_Mem/n9731 ), .SEL(
        N27), .F(\Data_Mem/n9735 ) );
  MUX \Data_Mem/U9798  ( .IN0(\Data_Mem/n9733 ), .IN1(\Data_Mem/n9732 ), .SEL(
        N28), .F(\Data_Mem/n9734 ) );
  MUX \Data_Mem/U9797  ( .IN0(o[287]), .IN1(o[319]), .SEL(N29), .F(
        \Data_Mem/n9733 ) );
  MUX \Data_Mem/U9796  ( .IN0(o[351]), .IN1(o[383]), .SEL(N29), .F(
        \Data_Mem/n9732 ) );
  MUX \Data_Mem/U9795  ( .IN0(\Data_Mem/n9730 ), .IN1(\Data_Mem/n9729 ), .SEL(
        N28), .F(\Data_Mem/n9731 ) );
  MUX \Data_Mem/U9794  ( .IN0(o[415]), .IN1(o[447]), .SEL(N29), .F(
        \Data_Mem/n9730 ) );
  MUX \Data_Mem/U9793  ( .IN0(o[479]), .IN1(o[511]), .SEL(N29), .F(
        \Data_Mem/n9729 ) );
  MUX \Data_Mem/U9792  ( .IN0(\Data_Mem/n9727 ), .IN1(\Data_Mem/n9720 ), .SEL(
        N26), .F(\Data_Mem/n9728 ) );
  MUX \Data_Mem/U9791  ( .IN0(\Data_Mem/n9726 ), .IN1(\Data_Mem/n9723 ), .SEL(
        N27), .F(\Data_Mem/n9727 ) );
  MUX \Data_Mem/U9790  ( .IN0(\Data_Mem/n9725 ), .IN1(\Data_Mem/n9724 ), .SEL(
        N28), .F(\Data_Mem/n9726 ) );
  MUX \Data_Mem/U9789  ( .IN0(o[543]), .IN1(o[575]), .SEL(N29), .F(
        \Data_Mem/n9725 ) );
  MUX \Data_Mem/U9788  ( .IN0(o[607]), .IN1(o[639]), .SEL(N29), .F(
        \Data_Mem/n9724 ) );
  MUX \Data_Mem/U9787  ( .IN0(\Data_Mem/n9722 ), .IN1(\Data_Mem/n9721 ), .SEL(
        N28), .F(\Data_Mem/n9723 ) );
  MUX \Data_Mem/U9786  ( .IN0(o[671]), .IN1(o[703]), .SEL(N29), .F(
        \Data_Mem/n9722 ) );
  MUX \Data_Mem/U9785  ( .IN0(o[735]), .IN1(o[767]), .SEL(N29), .F(
        \Data_Mem/n9721 ) );
  MUX \Data_Mem/U9784  ( .IN0(\Data_Mem/n9719 ), .IN1(\Data_Mem/n9716 ), .SEL(
        N27), .F(\Data_Mem/n9720 ) );
  MUX \Data_Mem/U9783  ( .IN0(\Data_Mem/n9718 ), .IN1(\Data_Mem/n9717 ), .SEL(
        N28), .F(\Data_Mem/n9719 ) );
  MUX \Data_Mem/U9782  ( .IN0(o[799]), .IN1(o[831]), .SEL(N29), .F(
        \Data_Mem/n9718 ) );
  MUX \Data_Mem/U9781  ( .IN0(o[863]), .IN1(o[895]), .SEL(N29), .F(
        \Data_Mem/n9717 ) );
  MUX \Data_Mem/U9780  ( .IN0(\Data_Mem/n9715 ), .IN1(\Data_Mem/n9714 ), .SEL(
        N28), .F(\Data_Mem/n9716 ) );
  MUX \Data_Mem/U9779  ( .IN0(o[927]), .IN1(o[959]), .SEL(N29), .F(
        \Data_Mem/n9715 ) );
  MUX \Data_Mem/U9778  ( .IN0(o[991]), .IN1(o[1023]), .SEL(N29), .F(
        \Data_Mem/n9714 ) );
  MUX \Data_Mem/U9777  ( .IN0(\Data_Mem/n9712 ), .IN1(\Data_Mem/n9697 ), .SEL(
        N25), .F(\Data_Mem/n9713 ) );
  MUX \Data_Mem/U9776  ( .IN0(\Data_Mem/n9711 ), .IN1(\Data_Mem/n9704 ), .SEL(
        N26), .F(\Data_Mem/n9712 ) );
  MUX \Data_Mem/U9775  ( .IN0(\Data_Mem/n9710 ), .IN1(\Data_Mem/n9707 ), .SEL(
        N27), .F(\Data_Mem/n9711 ) );
  MUX \Data_Mem/U9774  ( .IN0(\Data_Mem/n9709 ), .IN1(\Data_Mem/n9708 ), .SEL(
        N28), .F(\Data_Mem/n9710 ) );
  MUX \Data_Mem/U9773  ( .IN0(o[1055]), .IN1(o[1087]), .SEL(N29), .F(
        \Data_Mem/n9709 ) );
  MUX \Data_Mem/U9772  ( .IN0(o[1119]), .IN1(o[1151]), .SEL(N29), .F(
        \Data_Mem/n9708 ) );
  MUX \Data_Mem/U9771  ( .IN0(\Data_Mem/n9706 ), .IN1(\Data_Mem/n9705 ), .SEL(
        N28), .F(\Data_Mem/n9707 ) );
  MUX \Data_Mem/U9770  ( .IN0(o[1183]), .IN1(o[1215]), .SEL(N29), .F(
        \Data_Mem/n9706 ) );
  MUX \Data_Mem/U9769  ( .IN0(o[1247]), .IN1(o[1279]), .SEL(N29), .F(
        \Data_Mem/n9705 ) );
  MUX \Data_Mem/U9768  ( .IN0(\Data_Mem/n9703 ), .IN1(\Data_Mem/n9700 ), .SEL(
        N27), .F(\Data_Mem/n9704 ) );
  MUX \Data_Mem/U9767  ( .IN0(\Data_Mem/n9702 ), .IN1(\Data_Mem/n9701 ), .SEL(
        N28), .F(\Data_Mem/n9703 ) );
  MUX \Data_Mem/U9766  ( .IN0(o[1311]), .IN1(o[1343]), .SEL(N29), .F(
        \Data_Mem/n9702 ) );
  MUX \Data_Mem/U9765  ( .IN0(o[1375]), .IN1(o[1407]), .SEL(N29), .F(
        \Data_Mem/n9701 ) );
  MUX \Data_Mem/U9764  ( .IN0(\Data_Mem/n9699 ), .IN1(\Data_Mem/n9698 ), .SEL(
        N28), .F(\Data_Mem/n9700 ) );
  MUX \Data_Mem/U9763  ( .IN0(o[1439]), .IN1(o[1471]), .SEL(N29), .F(
        \Data_Mem/n9699 ) );
  MUX \Data_Mem/U9762  ( .IN0(o[1503]), .IN1(o[1535]), .SEL(N29), .F(
        \Data_Mem/n9698 ) );
  MUX \Data_Mem/U9761  ( .IN0(\Data_Mem/n9696 ), .IN1(\Data_Mem/n9689 ), .SEL(
        N26), .F(\Data_Mem/n9697 ) );
  MUX \Data_Mem/U9760  ( .IN0(\Data_Mem/n9695 ), .IN1(\Data_Mem/n9692 ), .SEL(
        N27), .F(\Data_Mem/n9696 ) );
  MUX \Data_Mem/U9759  ( .IN0(\Data_Mem/n9694 ), .IN1(\Data_Mem/n9693 ), .SEL(
        N28), .F(\Data_Mem/n9695 ) );
  MUX \Data_Mem/U9758  ( .IN0(o[1567]), .IN1(o[1599]), .SEL(N29), .F(
        \Data_Mem/n9694 ) );
  MUX \Data_Mem/U9757  ( .IN0(o[1631]), .IN1(o[1663]), .SEL(N29), .F(
        \Data_Mem/n9693 ) );
  MUX \Data_Mem/U9756  ( .IN0(\Data_Mem/n9691 ), .IN1(\Data_Mem/n9690 ), .SEL(
        N28), .F(\Data_Mem/n9692 ) );
  MUX \Data_Mem/U9755  ( .IN0(o[1695]), .IN1(o[1727]), .SEL(N29), .F(
        \Data_Mem/n9691 ) );
  MUX \Data_Mem/U9754  ( .IN0(o[1759]), .IN1(o[1791]), .SEL(N29), .F(
        \Data_Mem/n9690 ) );
  MUX \Data_Mem/U9753  ( .IN0(\Data_Mem/n9688 ), .IN1(\Data_Mem/n9685 ), .SEL(
        N27), .F(\Data_Mem/n9689 ) );
  MUX \Data_Mem/U9752  ( .IN0(\Data_Mem/n9687 ), .IN1(\Data_Mem/n9686 ), .SEL(
        N28), .F(\Data_Mem/n9688 ) );
  MUX \Data_Mem/U9751  ( .IN0(o[1823]), .IN1(o[1855]), .SEL(N29), .F(
        \Data_Mem/n9687 ) );
  MUX \Data_Mem/U9750  ( .IN0(o[1887]), .IN1(o[1919]), .SEL(N29), .F(
        \Data_Mem/n9686 ) );
  MUX \Data_Mem/U9749  ( .IN0(\Data_Mem/n9684 ), .IN1(\Data_Mem/n9683 ), .SEL(
        N28), .F(\Data_Mem/n9685 ) );
  MUX \Data_Mem/U9748  ( .IN0(o[1951]), .IN1(o[1983]), .SEL(N29), .F(
        \Data_Mem/n9684 ) );
  MUX \Data_Mem/U9747  ( .IN0(o[2015]), .IN1(o[2047]), .SEL(N29), .F(
        \Data_Mem/n9683 ) );
  MUX \Data_Mem/U9746  ( .IN0(\Data_Mem/n9682 ), .IN1(\Data_Mem/n9651 ), .SEL(
        N24), .F(\Data_Mem/N715 ) );
  MUX \Data_Mem/U9745  ( .IN0(\Data_Mem/n9681 ), .IN1(\Data_Mem/n9666 ), .SEL(
        N25), .F(\Data_Mem/n9682 ) );
  MUX \Data_Mem/U9744  ( .IN0(\Data_Mem/n9680 ), .IN1(\Data_Mem/n9673 ), .SEL(
        N26), .F(\Data_Mem/n9681 ) );
  MUX \Data_Mem/U9743  ( .IN0(\Data_Mem/n9679 ), .IN1(\Data_Mem/n9676 ), .SEL(
        N27), .F(\Data_Mem/n9680 ) );
  MUX \Data_Mem/U9742  ( .IN0(\Data_Mem/n9678 ), .IN1(\Data_Mem/n9677 ), .SEL(
        N28), .F(\Data_Mem/n9679 ) );
  MUX \Data_Mem/U9741  ( .IN0(o[30]), .IN1(o[62]), .SEL(N29), .F(
        \Data_Mem/n9678 ) );
  MUX \Data_Mem/U9740  ( .IN0(o[94]), .IN1(o[126]), .SEL(N29), .F(
        \Data_Mem/n9677 ) );
  MUX \Data_Mem/U9739  ( .IN0(\Data_Mem/n9675 ), .IN1(\Data_Mem/n9674 ), .SEL(
        N28), .F(\Data_Mem/n9676 ) );
  MUX \Data_Mem/U9738  ( .IN0(o[158]), .IN1(o[190]), .SEL(N29), .F(
        \Data_Mem/n9675 ) );
  MUX \Data_Mem/U9737  ( .IN0(o[222]), .IN1(o[254]), .SEL(N29), .F(
        \Data_Mem/n9674 ) );
  MUX \Data_Mem/U9736  ( .IN0(\Data_Mem/n9672 ), .IN1(\Data_Mem/n9669 ), .SEL(
        N27), .F(\Data_Mem/n9673 ) );
  MUX \Data_Mem/U9735  ( .IN0(\Data_Mem/n9671 ), .IN1(\Data_Mem/n9670 ), .SEL(
        N28), .F(\Data_Mem/n9672 ) );
  MUX \Data_Mem/U9734  ( .IN0(o[286]), .IN1(o[318]), .SEL(N29), .F(
        \Data_Mem/n9671 ) );
  MUX \Data_Mem/U9733  ( .IN0(o[350]), .IN1(o[382]), .SEL(N29), .F(
        \Data_Mem/n9670 ) );
  MUX \Data_Mem/U9732  ( .IN0(\Data_Mem/n9668 ), .IN1(\Data_Mem/n9667 ), .SEL(
        N28), .F(\Data_Mem/n9669 ) );
  MUX \Data_Mem/U9731  ( .IN0(o[414]), .IN1(o[446]), .SEL(N29), .F(
        \Data_Mem/n9668 ) );
  MUX \Data_Mem/U9730  ( .IN0(o[478]), .IN1(o[510]), .SEL(N29), .F(
        \Data_Mem/n9667 ) );
  MUX \Data_Mem/U9729  ( .IN0(\Data_Mem/n9665 ), .IN1(\Data_Mem/n9658 ), .SEL(
        N26), .F(\Data_Mem/n9666 ) );
  MUX \Data_Mem/U9728  ( .IN0(\Data_Mem/n9664 ), .IN1(\Data_Mem/n9661 ), .SEL(
        N27), .F(\Data_Mem/n9665 ) );
  MUX \Data_Mem/U9727  ( .IN0(\Data_Mem/n9663 ), .IN1(\Data_Mem/n9662 ), .SEL(
        N28), .F(\Data_Mem/n9664 ) );
  MUX \Data_Mem/U9726  ( .IN0(o[542]), .IN1(o[574]), .SEL(N29), .F(
        \Data_Mem/n9663 ) );
  MUX \Data_Mem/U9725  ( .IN0(o[606]), .IN1(o[638]), .SEL(N29), .F(
        \Data_Mem/n9662 ) );
  MUX \Data_Mem/U9724  ( .IN0(\Data_Mem/n9660 ), .IN1(\Data_Mem/n9659 ), .SEL(
        N28), .F(\Data_Mem/n9661 ) );
  MUX \Data_Mem/U9723  ( .IN0(o[670]), .IN1(o[702]), .SEL(N29), .F(
        \Data_Mem/n9660 ) );
  MUX \Data_Mem/U9722  ( .IN0(o[734]), .IN1(o[766]), .SEL(N29), .F(
        \Data_Mem/n9659 ) );
  MUX \Data_Mem/U9721  ( .IN0(\Data_Mem/n9657 ), .IN1(\Data_Mem/n9654 ), .SEL(
        N27), .F(\Data_Mem/n9658 ) );
  MUX \Data_Mem/U9720  ( .IN0(\Data_Mem/n9656 ), .IN1(\Data_Mem/n9655 ), .SEL(
        N28), .F(\Data_Mem/n9657 ) );
  MUX \Data_Mem/U9719  ( .IN0(o[798]), .IN1(o[830]), .SEL(N29), .F(
        \Data_Mem/n9656 ) );
  MUX \Data_Mem/U9718  ( .IN0(o[862]), .IN1(o[894]), .SEL(N29), .F(
        \Data_Mem/n9655 ) );
  MUX \Data_Mem/U9717  ( .IN0(\Data_Mem/n9653 ), .IN1(\Data_Mem/n9652 ), .SEL(
        N28), .F(\Data_Mem/n9654 ) );
  MUX \Data_Mem/U9716  ( .IN0(o[926]), .IN1(o[958]), .SEL(N29), .F(
        \Data_Mem/n9653 ) );
  MUX \Data_Mem/U9715  ( .IN0(o[990]), .IN1(o[1022]), .SEL(N29), .F(
        \Data_Mem/n9652 ) );
  MUX \Data_Mem/U9714  ( .IN0(\Data_Mem/n9650 ), .IN1(\Data_Mem/n9635 ), .SEL(
        N25), .F(\Data_Mem/n9651 ) );
  MUX \Data_Mem/U9713  ( .IN0(\Data_Mem/n9649 ), .IN1(\Data_Mem/n9642 ), .SEL(
        N26), .F(\Data_Mem/n9650 ) );
  MUX \Data_Mem/U9712  ( .IN0(\Data_Mem/n9648 ), .IN1(\Data_Mem/n9645 ), .SEL(
        N27), .F(\Data_Mem/n9649 ) );
  MUX \Data_Mem/U9711  ( .IN0(\Data_Mem/n9647 ), .IN1(\Data_Mem/n9646 ), .SEL(
        N28), .F(\Data_Mem/n9648 ) );
  MUX \Data_Mem/U9710  ( .IN0(o[1054]), .IN1(o[1086]), .SEL(N29), .F(
        \Data_Mem/n9647 ) );
  MUX \Data_Mem/U9709  ( .IN0(o[1118]), .IN1(o[1150]), .SEL(N29), .F(
        \Data_Mem/n9646 ) );
  MUX \Data_Mem/U9708  ( .IN0(\Data_Mem/n9644 ), .IN1(\Data_Mem/n9643 ), .SEL(
        N28), .F(\Data_Mem/n9645 ) );
  MUX \Data_Mem/U9707  ( .IN0(o[1182]), .IN1(o[1214]), .SEL(N29), .F(
        \Data_Mem/n9644 ) );
  MUX \Data_Mem/U9706  ( .IN0(o[1246]), .IN1(o[1278]), .SEL(N29), .F(
        \Data_Mem/n9643 ) );
  MUX \Data_Mem/U9705  ( .IN0(\Data_Mem/n9641 ), .IN1(\Data_Mem/n9638 ), .SEL(
        N27), .F(\Data_Mem/n9642 ) );
  MUX \Data_Mem/U9704  ( .IN0(\Data_Mem/n9640 ), .IN1(\Data_Mem/n9639 ), .SEL(
        N28), .F(\Data_Mem/n9641 ) );
  MUX \Data_Mem/U9703  ( .IN0(o[1310]), .IN1(o[1342]), .SEL(N29), .F(
        \Data_Mem/n9640 ) );
  MUX \Data_Mem/U9702  ( .IN0(o[1374]), .IN1(o[1406]), .SEL(N29), .F(
        \Data_Mem/n9639 ) );
  MUX \Data_Mem/U9701  ( .IN0(\Data_Mem/n9637 ), .IN1(\Data_Mem/n9636 ), .SEL(
        N28), .F(\Data_Mem/n9638 ) );
  MUX \Data_Mem/U9700  ( .IN0(o[1438]), .IN1(o[1470]), .SEL(N29), .F(
        \Data_Mem/n9637 ) );
  MUX \Data_Mem/U9699  ( .IN0(o[1502]), .IN1(o[1534]), .SEL(N29), .F(
        \Data_Mem/n9636 ) );
  MUX \Data_Mem/U9698  ( .IN0(\Data_Mem/n9634 ), .IN1(\Data_Mem/n9627 ), .SEL(
        N26), .F(\Data_Mem/n9635 ) );
  MUX \Data_Mem/U9697  ( .IN0(\Data_Mem/n9633 ), .IN1(\Data_Mem/n9630 ), .SEL(
        N27), .F(\Data_Mem/n9634 ) );
  MUX \Data_Mem/U9696  ( .IN0(\Data_Mem/n9632 ), .IN1(\Data_Mem/n9631 ), .SEL(
        N28), .F(\Data_Mem/n9633 ) );
  MUX \Data_Mem/U9695  ( .IN0(o[1566]), .IN1(o[1598]), .SEL(N29), .F(
        \Data_Mem/n9632 ) );
  MUX \Data_Mem/U9694  ( .IN0(o[1630]), .IN1(o[1662]), .SEL(N29), .F(
        \Data_Mem/n9631 ) );
  MUX \Data_Mem/U9693  ( .IN0(\Data_Mem/n9629 ), .IN1(\Data_Mem/n9628 ), .SEL(
        N28), .F(\Data_Mem/n9630 ) );
  MUX \Data_Mem/U9692  ( .IN0(o[1694]), .IN1(o[1726]), .SEL(N29), .F(
        \Data_Mem/n9629 ) );
  MUX \Data_Mem/U9691  ( .IN0(o[1758]), .IN1(o[1790]), .SEL(N29), .F(
        \Data_Mem/n9628 ) );
  MUX \Data_Mem/U9690  ( .IN0(\Data_Mem/n9626 ), .IN1(\Data_Mem/n9623 ), .SEL(
        N27), .F(\Data_Mem/n9627 ) );
  MUX \Data_Mem/U9689  ( .IN0(\Data_Mem/n9625 ), .IN1(\Data_Mem/n9624 ), .SEL(
        N28), .F(\Data_Mem/n9626 ) );
  MUX \Data_Mem/U9688  ( .IN0(o[1822]), .IN1(o[1854]), .SEL(N29), .F(
        \Data_Mem/n9625 ) );
  MUX \Data_Mem/U9687  ( .IN0(o[1886]), .IN1(o[1918]), .SEL(N29), .F(
        \Data_Mem/n9624 ) );
  MUX \Data_Mem/U9686  ( .IN0(\Data_Mem/n9622 ), .IN1(\Data_Mem/n9621 ), .SEL(
        N28), .F(\Data_Mem/n9623 ) );
  MUX \Data_Mem/U9685  ( .IN0(o[1950]), .IN1(o[1982]), .SEL(N29), .F(
        \Data_Mem/n9622 ) );
  MUX \Data_Mem/U9684  ( .IN0(o[2014]), .IN1(o[2046]), .SEL(N29), .F(
        \Data_Mem/n9621 ) );
  MUX \Data_Mem/U9683  ( .IN0(\Data_Mem/n9620 ), .IN1(\Data_Mem/n9589 ), .SEL(
        N24), .F(\Data_Mem/N716 ) );
  MUX \Data_Mem/U9682  ( .IN0(\Data_Mem/n9619 ), .IN1(\Data_Mem/n9604 ), .SEL(
        N25), .F(\Data_Mem/n9620 ) );
  MUX \Data_Mem/U9681  ( .IN0(\Data_Mem/n9618 ), .IN1(\Data_Mem/n9611 ), .SEL(
        N26), .F(\Data_Mem/n9619 ) );
  MUX \Data_Mem/U9680  ( .IN0(\Data_Mem/n9617 ), .IN1(\Data_Mem/n9614 ), .SEL(
        N27), .F(\Data_Mem/n9618 ) );
  MUX \Data_Mem/U9679  ( .IN0(\Data_Mem/n9616 ), .IN1(\Data_Mem/n9615 ), .SEL(
        N28), .F(\Data_Mem/n9617 ) );
  MUX \Data_Mem/U9678  ( .IN0(o[29]), .IN1(o[61]), .SEL(N29), .F(
        \Data_Mem/n9616 ) );
  MUX \Data_Mem/U9677  ( .IN0(o[93]), .IN1(o[125]), .SEL(N29), .F(
        \Data_Mem/n9615 ) );
  MUX \Data_Mem/U9676  ( .IN0(\Data_Mem/n9613 ), .IN1(\Data_Mem/n9612 ), .SEL(
        N28), .F(\Data_Mem/n9614 ) );
  MUX \Data_Mem/U9675  ( .IN0(o[157]), .IN1(o[189]), .SEL(N29), .F(
        \Data_Mem/n9613 ) );
  MUX \Data_Mem/U9674  ( .IN0(o[221]), .IN1(o[253]), .SEL(N29), .F(
        \Data_Mem/n9612 ) );
  MUX \Data_Mem/U9673  ( .IN0(\Data_Mem/n9610 ), .IN1(\Data_Mem/n9607 ), .SEL(
        N27), .F(\Data_Mem/n9611 ) );
  MUX \Data_Mem/U9672  ( .IN0(\Data_Mem/n9609 ), .IN1(\Data_Mem/n9608 ), .SEL(
        N28), .F(\Data_Mem/n9610 ) );
  MUX \Data_Mem/U9671  ( .IN0(o[285]), .IN1(o[317]), .SEL(N29), .F(
        \Data_Mem/n9609 ) );
  MUX \Data_Mem/U9670  ( .IN0(o[349]), .IN1(o[381]), .SEL(N29), .F(
        \Data_Mem/n9608 ) );
  MUX \Data_Mem/U9669  ( .IN0(\Data_Mem/n9606 ), .IN1(\Data_Mem/n9605 ), .SEL(
        N28), .F(\Data_Mem/n9607 ) );
  MUX \Data_Mem/U9668  ( .IN0(o[413]), .IN1(o[445]), .SEL(N29), .F(
        \Data_Mem/n9606 ) );
  MUX \Data_Mem/U9667  ( .IN0(o[477]), .IN1(o[509]), .SEL(N29), .F(
        \Data_Mem/n9605 ) );
  MUX \Data_Mem/U9666  ( .IN0(\Data_Mem/n9603 ), .IN1(\Data_Mem/n9596 ), .SEL(
        N26), .F(\Data_Mem/n9604 ) );
  MUX \Data_Mem/U9665  ( .IN0(\Data_Mem/n9602 ), .IN1(\Data_Mem/n9599 ), .SEL(
        N27), .F(\Data_Mem/n9603 ) );
  MUX \Data_Mem/U9664  ( .IN0(\Data_Mem/n9601 ), .IN1(\Data_Mem/n9600 ), .SEL(
        N28), .F(\Data_Mem/n9602 ) );
  MUX \Data_Mem/U9663  ( .IN0(o[541]), .IN1(o[573]), .SEL(N29), .F(
        \Data_Mem/n9601 ) );
  MUX \Data_Mem/U9662  ( .IN0(o[605]), .IN1(o[637]), .SEL(N29), .F(
        \Data_Mem/n9600 ) );
  MUX \Data_Mem/U9661  ( .IN0(\Data_Mem/n9598 ), .IN1(\Data_Mem/n9597 ), .SEL(
        N28), .F(\Data_Mem/n9599 ) );
  MUX \Data_Mem/U9660  ( .IN0(o[669]), .IN1(o[701]), .SEL(N29), .F(
        \Data_Mem/n9598 ) );
  MUX \Data_Mem/U9659  ( .IN0(o[733]), .IN1(o[765]), .SEL(N29), .F(
        \Data_Mem/n9597 ) );
  MUX \Data_Mem/U9658  ( .IN0(\Data_Mem/n9595 ), .IN1(\Data_Mem/n9592 ), .SEL(
        N27), .F(\Data_Mem/n9596 ) );
  MUX \Data_Mem/U9657  ( .IN0(\Data_Mem/n9594 ), .IN1(\Data_Mem/n9593 ), .SEL(
        N28), .F(\Data_Mem/n9595 ) );
  MUX \Data_Mem/U9656  ( .IN0(o[797]), .IN1(o[829]), .SEL(N29), .F(
        \Data_Mem/n9594 ) );
  MUX \Data_Mem/U9655  ( .IN0(o[861]), .IN1(o[893]), .SEL(N29), .F(
        \Data_Mem/n9593 ) );
  MUX \Data_Mem/U9654  ( .IN0(\Data_Mem/n9591 ), .IN1(\Data_Mem/n9590 ), .SEL(
        N28), .F(\Data_Mem/n9592 ) );
  MUX \Data_Mem/U9653  ( .IN0(o[925]), .IN1(o[957]), .SEL(N29), .F(
        \Data_Mem/n9591 ) );
  MUX \Data_Mem/U9652  ( .IN0(o[989]), .IN1(o[1021]), .SEL(N29), .F(
        \Data_Mem/n9590 ) );
  MUX \Data_Mem/U9651  ( .IN0(\Data_Mem/n9588 ), .IN1(\Data_Mem/n9573 ), .SEL(
        N25), .F(\Data_Mem/n9589 ) );
  MUX \Data_Mem/U9650  ( .IN0(\Data_Mem/n9587 ), .IN1(\Data_Mem/n9580 ), .SEL(
        N26), .F(\Data_Mem/n9588 ) );
  MUX \Data_Mem/U9649  ( .IN0(\Data_Mem/n9586 ), .IN1(\Data_Mem/n9583 ), .SEL(
        N27), .F(\Data_Mem/n9587 ) );
  MUX \Data_Mem/U9648  ( .IN0(\Data_Mem/n9585 ), .IN1(\Data_Mem/n9584 ), .SEL(
        N28), .F(\Data_Mem/n9586 ) );
  MUX \Data_Mem/U9647  ( .IN0(o[1053]), .IN1(o[1085]), .SEL(N29), .F(
        \Data_Mem/n9585 ) );
  MUX \Data_Mem/U9646  ( .IN0(o[1117]), .IN1(o[1149]), .SEL(N29), .F(
        \Data_Mem/n9584 ) );
  MUX \Data_Mem/U9645  ( .IN0(\Data_Mem/n9582 ), .IN1(\Data_Mem/n9581 ), .SEL(
        N28), .F(\Data_Mem/n9583 ) );
  MUX \Data_Mem/U9644  ( .IN0(o[1181]), .IN1(o[1213]), .SEL(N29), .F(
        \Data_Mem/n9582 ) );
  MUX \Data_Mem/U9643  ( .IN0(o[1245]), .IN1(o[1277]), .SEL(N29), .F(
        \Data_Mem/n9581 ) );
  MUX \Data_Mem/U9642  ( .IN0(\Data_Mem/n9579 ), .IN1(\Data_Mem/n9576 ), .SEL(
        N27), .F(\Data_Mem/n9580 ) );
  MUX \Data_Mem/U9641  ( .IN0(\Data_Mem/n9578 ), .IN1(\Data_Mem/n9577 ), .SEL(
        N28), .F(\Data_Mem/n9579 ) );
  MUX \Data_Mem/U9640  ( .IN0(o[1309]), .IN1(o[1341]), .SEL(N29), .F(
        \Data_Mem/n9578 ) );
  MUX \Data_Mem/U9639  ( .IN0(o[1373]), .IN1(o[1405]), .SEL(N29), .F(
        \Data_Mem/n9577 ) );
  MUX \Data_Mem/U9638  ( .IN0(\Data_Mem/n9575 ), .IN1(\Data_Mem/n9574 ), .SEL(
        N28), .F(\Data_Mem/n9576 ) );
  MUX \Data_Mem/U9637  ( .IN0(o[1437]), .IN1(o[1469]), .SEL(N29), .F(
        \Data_Mem/n9575 ) );
  MUX \Data_Mem/U9636  ( .IN0(o[1501]), .IN1(o[1533]), .SEL(N29), .F(
        \Data_Mem/n9574 ) );
  MUX \Data_Mem/U9635  ( .IN0(\Data_Mem/n9572 ), .IN1(\Data_Mem/n9565 ), .SEL(
        N26), .F(\Data_Mem/n9573 ) );
  MUX \Data_Mem/U9634  ( .IN0(\Data_Mem/n9571 ), .IN1(\Data_Mem/n9568 ), .SEL(
        N27), .F(\Data_Mem/n9572 ) );
  MUX \Data_Mem/U9633  ( .IN0(\Data_Mem/n9570 ), .IN1(\Data_Mem/n9569 ), .SEL(
        N28), .F(\Data_Mem/n9571 ) );
  MUX \Data_Mem/U9632  ( .IN0(o[1565]), .IN1(o[1597]), .SEL(N29), .F(
        \Data_Mem/n9570 ) );
  MUX \Data_Mem/U9631  ( .IN0(o[1629]), .IN1(o[1661]), .SEL(N29), .F(
        \Data_Mem/n9569 ) );
  MUX \Data_Mem/U9630  ( .IN0(\Data_Mem/n9567 ), .IN1(\Data_Mem/n9566 ), .SEL(
        N28), .F(\Data_Mem/n9568 ) );
  MUX \Data_Mem/U9629  ( .IN0(o[1693]), .IN1(o[1725]), .SEL(N29), .F(
        \Data_Mem/n9567 ) );
  MUX \Data_Mem/U9628  ( .IN0(o[1757]), .IN1(o[1789]), .SEL(N29), .F(
        \Data_Mem/n9566 ) );
  MUX \Data_Mem/U9627  ( .IN0(\Data_Mem/n9564 ), .IN1(\Data_Mem/n9561 ), .SEL(
        N27), .F(\Data_Mem/n9565 ) );
  MUX \Data_Mem/U9626  ( .IN0(\Data_Mem/n9563 ), .IN1(\Data_Mem/n9562 ), .SEL(
        N28), .F(\Data_Mem/n9564 ) );
  MUX \Data_Mem/U9625  ( .IN0(o[1821]), .IN1(o[1853]), .SEL(N29), .F(
        \Data_Mem/n9563 ) );
  MUX \Data_Mem/U9624  ( .IN0(o[1885]), .IN1(o[1917]), .SEL(N29), .F(
        \Data_Mem/n9562 ) );
  MUX \Data_Mem/U9623  ( .IN0(\Data_Mem/n9560 ), .IN1(\Data_Mem/n9559 ), .SEL(
        N28), .F(\Data_Mem/n9561 ) );
  MUX \Data_Mem/U9622  ( .IN0(o[1949]), .IN1(o[1981]), .SEL(N29), .F(
        \Data_Mem/n9560 ) );
  MUX \Data_Mem/U9621  ( .IN0(o[2013]), .IN1(o[2045]), .SEL(N29), .F(
        \Data_Mem/n9559 ) );
  MUX \Data_Mem/U9620  ( .IN0(\Data_Mem/n9558 ), .IN1(\Data_Mem/n9527 ), .SEL(
        N24), .F(\Data_Mem/N717 ) );
  MUX \Data_Mem/U9619  ( .IN0(\Data_Mem/n9557 ), .IN1(\Data_Mem/n9542 ), .SEL(
        N25), .F(\Data_Mem/n9558 ) );
  MUX \Data_Mem/U9618  ( .IN0(\Data_Mem/n9556 ), .IN1(\Data_Mem/n9549 ), .SEL(
        N26), .F(\Data_Mem/n9557 ) );
  MUX \Data_Mem/U9617  ( .IN0(\Data_Mem/n9555 ), .IN1(\Data_Mem/n9552 ), .SEL(
        N27), .F(\Data_Mem/n9556 ) );
  MUX \Data_Mem/U9616  ( .IN0(\Data_Mem/n9554 ), .IN1(\Data_Mem/n9553 ), .SEL(
        N28), .F(\Data_Mem/n9555 ) );
  MUX \Data_Mem/U9615  ( .IN0(o[28]), .IN1(o[60]), .SEL(N29), .F(
        \Data_Mem/n9554 ) );
  MUX \Data_Mem/U9614  ( .IN0(o[92]), .IN1(o[124]), .SEL(N29), .F(
        \Data_Mem/n9553 ) );
  MUX \Data_Mem/U9613  ( .IN0(\Data_Mem/n9551 ), .IN1(\Data_Mem/n9550 ), .SEL(
        N28), .F(\Data_Mem/n9552 ) );
  MUX \Data_Mem/U9612  ( .IN0(o[156]), .IN1(o[188]), .SEL(N29), .F(
        \Data_Mem/n9551 ) );
  MUX \Data_Mem/U9611  ( .IN0(o[220]), .IN1(o[252]), .SEL(N29), .F(
        \Data_Mem/n9550 ) );
  MUX \Data_Mem/U9610  ( .IN0(\Data_Mem/n9548 ), .IN1(\Data_Mem/n9545 ), .SEL(
        N27), .F(\Data_Mem/n9549 ) );
  MUX \Data_Mem/U9609  ( .IN0(\Data_Mem/n9547 ), .IN1(\Data_Mem/n9546 ), .SEL(
        N28), .F(\Data_Mem/n9548 ) );
  MUX \Data_Mem/U9608  ( .IN0(o[284]), .IN1(o[316]), .SEL(N29), .F(
        \Data_Mem/n9547 ) );
  MUX \Data_Mem/U9607  ( .IN0(o[348]), .IN1(o[380]), .SEL(N29), .F(
        \Data_Mem/n9546 ) );
  MUX \Data_Mem/U9606  ( .IN0(\Data_Mem/n9544 ), .IN1(\Data_Mem/n9543 ), .SEL(
        N28), .F(\Data_Mem/n9545 ) );
  MUX \Data_Mem/U9605  ( .IN0(o[412]), .IN1(o[444]), .SEL(N29), .F(
        \Data_Mem/n9544 ) );
  MUX \Data_Mem/U9604  ( .IN0(o[476]), .IN1(o[508]), .SEL(N29), .F(
        \Data_Mem/n9543 ) );
  MUX \Data_Mem/U9603  ( .IN0(\Data_Mem/n9541 ), .IN1(\Data_Mem/n9534 ), .SEL(
        N26), .F(\Data_Mem/n9542 ) );
  MUX \Data_Mem/U9602  ( .IN0(\Data_Mem/n9540 ), .IN1(\Data_Mem/n9537 ), .SEL(
        N27), .F(\Data_Mem/n9541 ) );
  MUX \Data_Mem/U9601  ( .IN0(\Data_Mem/n9539 ), .IN1(\Data_Mem/n9538 ), .SEL(
        N28), .F(\Data_Mem/n9540 ) );
  MUX \Data_Mem/U9600  ( .IN0(o[540]), .IN1(o[572]), .SEL(N29), .F(
        \Data_Mem/n9539 ) );
  MUX \Data_Mem/U9599  ( .IN0(o[604]), .IN1(o[636]), .SEL(N29), .F(
        \Data_Mem/n9538 ) );
  MUX \Data_Mem/U9598  ( .IN0(\Data_Mem/n9536 ), .IN1(\Data_Mem/n9535 ), .SEL(
        N28), .F(\Data_Mem/n9537 ) );
  MUX \Data_Mem/U9597  ( .IN0(o[668]), .IN1(o[700]), .SEL(N29), .F(
        \Data_Mem/n9536 ) );
  MUX \Data_Mem/U9596  ( .IN0(o[732]), .IN1(o[764]), .SEL(N29), .F(
        \Data_Mem/n9535 ) );
  MUX \Data_Mem/U9595  ( .IN0(\Data_Mem/n9533 ), .IN1(\Data_Mem/n9530 ), .SEL(
        N27), .F(\Data_Mem/n9534 ) );
  MUX \Data_Mem/U9594  ( .IN0(\Data_Mem/n9532 ), .IN1(\Data_Mem/n9531 ), .SEL(
        N28), .F(\Data_Mem/n9533 ) );
  MUX \Data_Mem/U9593  ( .IN0(o[796]), .IN1(o[828]), .SEL(N29), .F(
        \Data_Mem/n9532 ) );
  MUX \Data_Mem/U9592  ( .IN0(o[860]), .IN1(o[892]), .SEL(N29), .F(
        \Data_Mem/n9531 ) );
  MUX \Data_Mem/U9591  ( .IN0(\Data_Mem/n9529 ), .IN1(\Data_Mem/n9528 ), .SEL(
        N28), .F(\Data_Mem/n9530 ) );
  MUX \Data_Mem/U9590  ( .IN0(o[924]), .IN1(o[956]), .SEL(N29), .F(
        \Data_Mem/n9529 ) );
  MUX \Data_Mem/U9589  ( .IN0(o[988]), .IN1(o[1020]), .SEL(N29), .F(
        \Data_Mem/n9528 ) );
  MUX \Data_Mem/U9588  ( .IN0(\Data_Mem/n9526 ), .IN1(\Data_Mem/n9511 ), .SEL(
        N25), .F(\Data_Mem/n9527 ) );
  MUX \Data_Mem/U9587  ( .IN0(\Data_Mem/n9525 ), .IN1(\Data_Mem/n9518 ), .SEL(
        N26), .F(\Data_Mem/n9526 ) );
  MUX \Data_Mem/U9586  ( .IN0(\Data_Mem/n9524 ), .IN1(\Data_Mem/n9521 ), .SEL(
        N27), .F(\Data_Mem/n9525 ) );
  MUX \Data_Mem/U9585  ( .IN0(\Data_Mem/n9523 ), .IN1(\Data_Mem/n9522 ), .SEL(
        N28), .F(\Data_Mem/n9524 ) );
  MUX \Data_Mem/U9584  ( .IN0(o[1052]), .IN1(o[1084]), .SEL(N29), .F(
        \Data_Mem/n9523 ) );
  MUX \Data_Mem/U9583  ( .IN0(o[1116]), .IN1(o[1148]), .SEL(N29), .F(
        \Data_Mem/n9522 ) );
  MUX \Data_Mem/U9582  ( .IN0(\Data_Mem/n9520 ), .IN1(\Data_Mem/n9519 ), .SEL(
        N28), .F(\Data_Mem/n9521 ) );
  MUX \Data_Mem/U9581  ( .IN0(o[1180]), .IN1(o[1212]), .SEL(N29), .F(
        \Data_Mem/n9520 ) );
  MUX \Data_Mem/U9580  ( .IN0(o[1244]), .IN1(o[1276]), .SEL(N29), .F(
        \Data_Mem/n9519 ) );
  MUX \Data_Mem/U9579  ( .IN0(\Data_Mem/n9517 ), .IN1(\Data_Mem/n9514 ), .SEL(
        N27), .F(\Data_Mem/n9518 ) );
  MUX \Data_Mem/U9578  ( .IN0(\Data_Mem/n9516 ), .IN1(\Data_Mem/n9515 ), .SEL(
        N28), .F(\Data_Mem/n9517 ) );
  MUX \Data_Mem/U9577  ( .IN0(o[1308]), .IN1(o[1340]), .SEL(N29), .F(
        \Data_Mem/n9516 ) );
  MUX \Data_Mem/U9576  ( .IN0(o[1372]), .IN1(o[1404]), .SEL(N29), .F(
        \Data_Mem/n9515 ) );
  MUX \Data_Mem/U9575  ( .IN0(\Data_Mem/n9513 ), .IN1(\Data_Mem/n9512 ), .SEL(
        N28), .F(\Data_Mem/n9514 ) );
  MUX \Data_Mem/U9574  ( .IN0(o[1436]), .IN1(o[1468]), .SEL(N29), .F(
        \Data_Mem/n9513 ) );
  MUX \Data_Mem/U9573  ( .IN0(o[1500]), .IN1(o[1532]), .SEL(N29), .F(
        \Data_Mem/n9512 ) );
  MUX \Data_Mem/U9572  ( .IN0(\Data_Mem/n9510 ), .IN1(\Data_Mem/n9503 ), .SEL(
        N26), .F(\Data_Mem/n9511 ) );
  MUX \Data_Mem/U9571  ( .IN0(\Data_Mem/n9509 ), .IN1(\Data_Mem/n9506 ), .SEL(
        N27), .F(\Data_Mem/n9510 ) );
  MUX \Data_Mem/U9570  ( .IN0(\Data_Mem/n9508 ), .IN1(\Data_Mem/n9507 ), .SEL(
        N28), .F(\Data_Mem/n9509 ) );
  MUX \Data_Mem/U9569  ( .IN0(o[1564]), .IN1(o[1596]), .SEL(N29), .F(
        \Data_Mem/n9508 ) );
  MUX \Data_Mem/U9568  ( .IN0(o[1628]), .IN1(o[1660]), .SEL(N29), .F(
        \Data_Mem/n9507 ) );
  MUX \Data_Mem/U9567  ( .IN0(\Data_Mem/n9505 ), .IN1(\Data_Mem/n9504 ), .SEL(
        N28), .F(\Data_Mem/n9506 ) );
  MUX \Data_Mem/U9566  ( .IN0(o[1692]), .IN1(o[1724]), .SEL(N29), .F(
        \Data_Mem/n9505 ) );
  MUX \Data_Mem/U9565  ( .IN0(o[1756]), .IN1(o[1788]), .SEL(N29), .F(
        \Data_Mem/n9504 ) );
  MUX \Data_Mem/U9564  ( .IN0(\Data_Mem/n9502 ), .IN1(\Data_Mem/n9499 ), .SEL(
        N27), .F(\Data_Mem/n9503 ) );
  MUX \Data_Mem/U9563  ( .IN0(\Data_Mem/n9501 ), .IN1(\Data_Mem/n9500 ), .SEL(
        N28), .F(\Data_Mem/n9502 ) );
  MUX \Data_Mem/U9562  ( .IN0(o[1820]), .IN1(o[1852]), .SEL(N29), .F(
        \Data_Mem/n9501 ) );
  MUX \Data_Mem/U9561  ( .IN0(o[1884]), .IN1(o[1916]), .SEL(N29), .F(
        \Data_Mem/n9500 ) );
  MUX \Data_Mem/U9560  ( .IN0(\Data_Mem/n9498 ), .IN1(\Data_Mem/n9497 ), .SEL(
        N28), .F(\Data_Mem/n9499 ) );
  MUX \Data_Mem/U9559  ( .IN0(o[1948]), .IN1(o[1980]), .SEL(N29), .F(
        \Data_Mem/n9498 ) );
  MUX \Data_Mem/U9558  ( .IN0(o[2012]), .IN1(o[2044]), .SEL(N29), .F(
        \Data_Mem/n9497 ) );
  MUX \Data_Mem/U9557  ( .IN0(\Data_Mem/n9496 ), .IN1(\Data_Mem/n9465 ), .SEL(
        N24), .F(\Data_Mem/N718 ) );
  MUX \Data_Mem/U9556  ( .IN0(\Data_Mem/n9495 ), .IN1(\Data_Mem/n9480 ), .SEL(
        N25), .F(\Data_Mem/n9496 ) );
  MUX \Data_Mem/U9555  ( .IN0(\Data_Mem/n9494 ), .IN1(\Data_Mem/n9487 ), .SEL(
        N26), .F(\Data_Mem/n9495 ) );
  MUX \Data_Mem/U9554  ( .IN0(\Data_Mem/n9493 ), .IN1(\Data_Mem/n9490 ), .SEL(
        N27), .F(\Data_Mem/n9494 ) );
  MUX \Data_Mem/U9553  ( .IN0(\Data_Mem/n9492 ), .IN1(\Data_Mem/n9491 ), .SEL(
        N28), .F(\Data_Mem/n9493 ) );
  MUX \Data_Mem/U9552  ( .IN0(o[27]), .IN1(o[59]), .SEL(N29), .F(
        \Data_Mem/n9492 ) );
  MUX \Data_Mem/U9551  ( .IN0(o[91]), .IN1(o[123]), .SEL(N29), .F(
        \Data_Mem/n9491 ) );
  MUX \Data_Mem/U9550  ( .IN0(\Data_Mem/n9489 ), .IN1(\Data_Mem/n9488 ), .SEL(
        N28), .F(\Data_Mem/n9490 ) );
  MUX \Data_Mem/U9549  ( .IN0(o[155]), .IN1(o[187]), .SEL(N29), .F(
        \Data_Mem/n9489 ) );
  MUX \Data_Mem/U9548  ( .IN0(o[219]), .IN1(o[251]), .SEL(N29), .F(
        \Data_Mem/n9488 ) );
  MUX \Data_Mem/U9547  ( .IN0(\Data_Mem/n9486 ), .IN1(\Data_Mem/n9483 ), .SEL(
        N27), .F(\Data_Mem/n9487 ) );
  MUX \Data_Mem/U9546  ( .IN0(\Data_Mem/n9485 ), .IN1(\Data_Mem/n9484 ), .SEL(
        N28), .F(\Data_Mem/n9486 ) );
  MUX \Data_Mem/U9545  ( .IN0(o[283]), .IN1(o[315]), .SEL(N29), .F(
        \Data_Mem/n9485 ) );
  MUX \Data_Mem/U9544  ( .IN0(o[347]), .IN1(o[379]), .SEL(N29), .F(
        \Data_Mem/n9484 ) );
  MUX \Data_Mem/U9543  ( .IN0(\Data_Mem/n9482 ), .IN1(\Data_Mem/n9481 ), .SEL(
        N28), .F(\Data_Mem/n9483 ) );
  MUX \Data_Mem/U9542  ( .IN0(o[411]), .IN1(o[443]), .SEL(N29), .F(
        \Data_Mem/n9482 ) );
  MUX \Data_Mem/U9541  ( .IN0(o[475]), .IN1(o[507]), .SEL(N29), .F(
        \Data_Mem/n9481 ) );
  MUX \Data_Mem/U9540  ( .IN0(\Data_Mem/n9479 ), .IN1(\Data_Mem/n9472 ), .SEL(
        N26), .F(\Data_Mem/n9480 ) );
  MUX \Data_Mem/U9539  ( .IN0(\Data_Mem/n9478 ), .IN1(\Data_Mem/n9475 ), .SEL(
        N27), .F(\Data_Mem/n9479 ) );
  MUX \Data_Mem/U9538  ( .IN0(\Data_Mem/n9477 ), .IN1(\Data_Mem/n9476 ), .SEL(
        N28), .F(\Data_Mem/n9478 ) );
  MUX \Data_Mem/U9537  ( .IN0(o[539]), .IN1(o[571]), .SEL(N29), .F(
        \Data_Mem/n9477 ) );
  MUX \Data_Mem/U9536  ( .IN0(o[603]), .IN1(o[635]), .SEL(N29), .F(
        \Data_Mem/n9476 ) );
  MUX \Data_Mem/U9535  ( .IN0(\Data_Mem/n9474 ), .IN1(\Data_Mem/n9473 ), .SEL(
        N28), .F(\Data_Mem/n9475 ) );
  MUX \Data_Mem/U9534  ( .IN0(o[667]), .IN1(o[699]), .SEL(N29), .F(
        \Data_Mem/n9474 ) );
  MUX \Data_Mem/U9533  ( .IN0(o[731]), .IN1(o[763]), .SEL(N29), .F(
        \Data_Mem/n9473 ) );
  MUX \Data_Mem/U9532  ( .IN0(\Data_Mem/n9471 ), .IN1(\Data_Mem/n9468 ), .SEL(
        N27), .F(\Data_Mem/n9472 ) );
  MUX \Data_Mem/U9531  ( .IN0(\Data_Mem/n9470 ), .IN1(\Data_Mem/n9469 ), .SEL(
        N28), .F(\Data_Mem/n9471 ) );
  MUX \Data_Mem/U9530  ( .IN0(o[795]), .IN1(o[827]), .SEL(N29), .F(
        \Data_Mem/n9470 ) );
  MUX \Data_Mem/U9529  ( .IN0(o[859]), .IN1(o[891]), .SEL(N29), .F(
        \Data_Mem/n9469 ) );
  MUX \Data_Mem/U9528  ( .IN0(\Data_Mem/n9467 ), .IN1(\Data_Mem/n9466 ), .SEL(
        N28), .F(\Data_Mem/n9468 ) );
  MUX \Data_Mem/U9527  ( .IN0(o[923]), .IN1(o[955]), .SEL(N29), .F(
        \Data_Mem/n9467 ) );
  MUX \Data_Mem/U9526  ( .IN0(o[987]), .IN1(o[1019]), .SEL(N29), .F(
        \Data_Mem/n9466 ) );
  MUX \Data_Mem/U9525  ( .IN0(\Data_Mem/n9464 ), .IN1(\Data_Mem/n9449 ), .SEL(
        N25), .F(\Data_Mem/n9465 ) );
  MUX \Data_Mem/U9524  ( .IN0(\Data_Mem/n9463 ), .IN1(\Data_Mem/n9456 ), .SEL(
        N26), .F(\Data_Mem/n9464 ) );
  MUX \Data_Mem/U9523  ( .IN0(\Data_Mem/n9462 ), .IN1(\Data_Mem/n9459 ), .SEL(
        N27), .F(\Data_Mem/n9463 ) );
  MUX \Data_Mem/U9522  ( .IN0(\Data_Mem/n9461 ), .IN1(\Data_Mem/n9460 ), .SEL(
        N28), .F(\Data_Mem/n9462 ) );
  MUX \Data_Mem/U9521  ( .IN0(o[1051]), .IN1(o[1083]), .SEL(N29), .F(
        \Data_Mem/n9461 ) );
  MUX \Data_Mem/U9520  ( .IN0(o[1115]), .IN1(o[1147]), .SEL(N29), .F(
        \Data_Mem/n9460 ) );
  MUX \Data_Mem/U9519  ( .IN0(\Data_Mem/n9458 ), .IN1(\Data_Mem/n9457 ), .SEL(
        N28), .F(\Data_Mem/n9459 ) );
  MUX \Data_Mem/U9518  ( .IN0(o[1179]), .IN1(o[1211]), .SEL(N29), .F(
        \Data_Mem/n9458 ) );
  MUX \Data_Mem/U9517  ( .IN0(o[1243]), .IN1(o[1275]), .SEL(N29), .F(
        \Data_Mem/n9457 ) );
  MUX \Data_Mem/U9516  ( .IN0(\Data_Mem/n9455 ), .IN1(\Data_Mem/n9452 ), .SEL(
        N27), .F(\Data_Mem/n9456 ) );
  MUX \Data_Mem/U9515  ( .IN0(\Data_Mem/n9454 ), .IN1(\Data_Mem/n9453 ), .SEL(
        N28), .F(\Data_Mem/n9455 ) );
  MUX \Data_Mem/U9514  ( .IN0(o[1307]), .IN1(o[1339]), .SEL(N29), .F(
        \Data_Mem/n9454 ) );
  MUX \Data_Mem/U9513  ( .IN0(o[1371]), .IN1(o[1403]), .SEL(N29), .F(
        \Data_Mem/n9453 ) );
  MUX \Data_Mem/U9512  ( .IN0(\Data_Mem/n9451 ), .IN1(\Data_Mem/n9450 ), .SEL(
        N28), .F(\Data_Mem/n9452 ) );
  MUX \Data_Mem/U9511  ( .IN0(o[1435]), .IN1(o[1467]), .SEL(N29), .F(
        \Data_Mem/n9451 ) );
  MUX \Data_Mem/U9510  ( .IN0(o[1499]), .IN1(o[1531]), .SEL(N29), .F(
        \Data_Mem/n9450 ) );
  MUX \Data_Mem/U9509  ( .IN0(\Data_Mem/n9448 ), .IN1(\Data_Mem/n9441 ), .SEL(
        N26), .F(\Data_Mem/n9449 ) );
  MUX \Data_Mem/U9508  ( .IN0(\Data_Mem/n9447 ), .IN1(\Data_Mem/n9444 ), .SEL(
        N27), .F(\Data_Mem/n9448 ) );
  MUX \Data_Mem/U9507  ( .IN0(\Data_Mem/n9446 ), .IN1(\Data_Mem/n9445 ), .SEL(
        N28), .F(\Data_Mem/n9447 ) );
  MUX \Data_Mem/U9506  ( .IN0(o[1563]), .IN1(o[1595]), .SEL(N29), .F(
        \Data_Mem/n9446 ) );
  MUX \Data_Mem/U9505  ( .IN0(o[1627]), .IN1(o[1659]), .SEL(N29), .F(
        \Data_Mem/n9445 ) );
  MUX \Data_Mem/U9504  ( .IN0(\Data_Mem/n9443 ), .IN1(\Data_Mem/n9442 ), .SEL(
        N28), .F(\Data_Mem/n9444 ) );
  MUX \Data_Mem/U9503  ( .IN0(o[1691]), .IN1(o[1723]), .SEL(N29), .F(
        \Data_Mem/n9443 ) );
  MUX \Data_Mem/U9502  ( .IN0(o[1755]), .IN1(o[1787]), .SEL(N29), .F(
        \Data_Mem/n9442 ) );
  MUX \Data_Mem/U9501  ( .IN0(\Data_Mem/n9440 ), .IN1(\Data_Mem/n9437 ), .SEL(
        N27), .F(\Data_Mem/n9441 ) );
  MUX \Data_Mem/U9500  ( .IN0(\Data_Mem/n9439 ), .IN1(\Data_Mem/n9438 ), .SEL(
        N28), .F(\Data_Mem/n9440 ) );
  MUX \Data_Mem/U9499  ( .IN0(o[1819]), .IN1(o[1851]), .SEL(N29), .F(
        \Data_Mem/n9439 ) );
  MUX \Data_Mem/U9498  ( .IN0(o[1883]), .IN1(o[1915]), .SEL(N29), .F(
        \Data_Mem/n9438 ) );
  MUX \Data_Mem/U9497  ( .IN0(\Data_Mem/n9436 ), .IN1(\Data_Mem/n9435 ), .SEL(
        N28), .F(\Data_Mem/n9437 ) );
  MUX \Data_Mem/U9496  ( .IN0(o[1947]), .IN1(o[1979]), .SEL(N29), .F(
        \Data_Mem/n9436 ) );
  MUX \Data_Mem/U9495  ( .IN0(o[2011]), .IN1(o[2043]), .SEL(N29), .F(
        \Data_Mem/n9435 ) );
  MUX \Data_Mem/U9494  ( .IN0(\Data_Mem/n9434 ), .IN1(\Data_Mem/n9403 ), .SEL(
        N24), .F(\Data_Mem/N719 ) );
  MUX \Data_Mem/U9493  ( .IN0(\Data_Mem/n9433 ), .IN1(\Data_Mem/n9418 ), .SEL(
        N25), .F(\Data_Mem/n9434 ) );
  MUX \Data_Mem/U9492  ( .IN0(\Data_Mem/n9432 ), .IN1(\Data_Mem/n9425 ), .SEL(
        N26), .F(\Data_Mem/n9433 ) );
  MUX \Data_Mem/U9491  ( .IN0(\Data_Mem/n9431 ), .IN1(\Data_Mem/n9428 ), .SEL(
        N27), .F(\Data_Mem/n9432 ) );
  MUX \Data_Mem/U9490  ( .IN0(\Data_Mem/n9430 ), .IN1(\Data_Mem/n9429 ), .SEL(
        N28), .F(\Data_Mem/n9431 ) );
  MUX \Data_Mem/U9489  ( .IN0(o[26]), .IN1(o[58]), .SEL(N29), .F(
        \Data_Mem/n9430 ) );
  MUX \Data_Mem/U9488  ( .IN0(o[90]), .IN1(o[122]), .SEL(N29), .F(
        \Data_Mem/n9429 ) );
  MUX \Data_Mem/U9487  ( .IN0(\Data_Mem/n9427 ), .IN1(\Data_Mem/n9426 ), .SEL(
        N28), .F(\Data_Mem/n9428 ) );
  MUX \Data_Mem/U9486  ( .IN0(o[154]), .IN1(o[186]), .SEL(N29), .F(
        \Data_Mem/n9427 ) );
  MUX \Data_Mem/U9485  ( .IN0(o[218]), .IN1(o[250]), .SEL(N29), .F(
        \Data_Mem/n9426 ) );
  MUX \Data_Mem/U9484  ( .IN0(\Data_Mem/n9424 ), .IN1(\Data_Mem/n9421 ), .SEL(
        N27), .F(\Data_Mem/n9425 ) );
  MUX \Data_Mem/U9483  ( .IN0(\Data_Mem/n9423 ), .IN1(\Data_Mem/n9422 ), .SEL(
        N28), .F(\Data_Mem/n9424 ) );
  MUX \Data_Mem/U9482  ( .IN0(o[282]), .IN1(o[314]), .SEL(N29), .F(
        \Data_Mem/n9423 ) );
  MUX \Data_Mem/U9481  ( .IN0(o[346]), .IN1(o[378]), .SEL(N29), .F(
        \Data_Mem/n9422 ) );
  MUX \Data_Mem/U9480  ( .IN0(\Data_Mem/n9420 ), .IN1(\Data_Mem/n9419 ), .SEL(
        N28), .F(\Data_Mem/n9421 ) );
  MUX \Data_Mem/U9479  ( .IN0(o[410]), .IN1(o[442]), .SEL(N29), .F(
        \Data_Mem/n9420 ) );
  MUX \Data_Mem/U9478  ( .IN0(o[474]), .IN1(o[506]), .SEL(N29), .F(
        \Data_Mem/n9419 ) );
  MUX \Data_Mem/U9477  ( .IN0(\Data_Mem/n9417 ), .IN1(\Data_Mem/n9410 ), .SEL(
        N26), .F(\Data_Mem/n9418 ) );
  MUX \Data_Mem/U9476  ( .IN0(\Data_Mem/n9416 ), .IN1(\Data_Mem/n9413 ), .SEL(
        N27), .F(\Data_Mem/n9417 ) );
  MUX \Data_Mem/U9475  ( .IN0(\Data_Mem/n9415 ), .IN1(\Data_Mem/n9414 ), .SEL(
        N28), .F(\Data_Mem/n9416 ) );
  MUX \Data_Mem/U9474  ( .IN0(o[538]), .IN1(o[570]), .SEL(N29), .F(
        \Data_Mem/n9415 ) );
  MUX \Data_Mem/U9473  ( .IN0(o[602]), .IN1(o[634]), .SEL(N29), .F(
        \Data_Mem/n9414 ) );
  MUX \Data_Mem/U9472  ( .IN0(\Data_Mem/n9412 ), .IN1(\Data_Mem/n9411 ), .SEL(
        N28), .F(\Data_Mem/n9413 ) );
  MUX \Data_Mem/U9471  ( .IN0(o[666]), .IN1(o[698]), .SEL(N29), .F(
        \Data_Mem/n9412 ) );
  MUX \Data_Mem/U9470  ( .IN0(o[730]), .IN1(o[762]), .SEL(N29), .F(
        \Data_Mem/n9411 ) );
  MUX \Data_Mem/U9469  ( .IN0(\Data_Mem/n9409 ), .IN1(\Data_Mem/n9406 ), .SEL(
        N27), .F(\Data_Mem/n9410 ) );
  MUX \Data_Mem/U9468  ( .IN0(\Data_Mem/n9408 ), .IN1(\Data_Mem/n9407 ), .SEL(
        N28), .F(\Data_Mem/n9409 ) );
  MUX \Data_Mem/U9467  ( .IN0(o[794]), .IN1(o[826]), .SEL(N29), .F(
        \Data_Mem/n9408 ) );
  MUX \Data_Mem/U9466  ( .IN0(o[858]), .IN1(o[890]), .SEL(N29), .F(
        \Data_Mem/n9407 ) );
  MUX \Data_Mem/U9465  ( .IN0(\Data_Mem/n9405 ), .IN1(\Data_Mem/n9404 ), .SEL(
        N28), .F(\Data_Mem/n9406 ) );
  MUX \Data_Mem/U9464  ( .IN0(o[922]), .IN1(o[954]), .SEL(N29), .F(
        \Data_Mem/n9405 ) );
  MUX \Data_Mem/U9463  ( .IN0(o[986]), .IN1(o[1018]), .SEL(N29), .F(
        \Data_Mem/n9404 ) );
  MUX \Data_Mem/U9462  ( .IN0(\Data_Mem/n9402 ), .IN1(\Data_Mem/n9387 ), .SEL(
        N25), .F(\Data_Mem/n9403 ) );
  MUX \Data_Mem/U9461  ( .IN0(\Data_Mem/n9401 ), .IN1(\Data_Mem/n9394 ), .SEL(
        N26), .F(\Data_Mem/n9402 ) );
  MUX \Data_Mem/U9460  ( .IN0(\Data_Mem/n9400 ), .IN1(\Data_Mem/n9397 ), .SEL(
        N27), .F(\Data_Mem/n9401 ) );
  MUX \Data_Mem/U9459  ( .IN0(\Data_Mem/n9399 ), .IN1(\Data_Mem/n9398 ), .SEL(
        N28), .F(\Data_Mem/n9400 ) );
  MUX \Data_Mem/U9458  ( .IN0(o[1050]), .IN1(o[1082]), .SEL(N29), .F(
        \Data_Mem/n9399 ) );
  MUX \Data_Mem/U9457  ( .IN0(o[1114]), .IN1(o[1146]), .SEL(N29), .F(
        \Data_Mem/n9398 ) );
  MUX \Data_Mem/U9456  ( .IN0(\Data_Mem/n9396 ), .IN1(\Data_Mem/n9395 ), .SEL(
        N28), .F(\Data_Mem/n9397 ) );
  MUX \Data_Mem/U9455  ( .IN0(o[1178]), .IN1(o[1210]), .SEL(N29), .F(
        \Data_Mem/n9396 ) );
  MUX \Data_Mem/U9454  ( .IN0(o[1242]), .IN1(o[1274]), .SEL(N29), .F(
        \Data_Mem/n9395 ) );
  MUX \Data_Mem/U9453  ( .IN0(\Data_Mem/n9393 ), .IN1(\Data_Mem/n9390 ), .SEL(
        N27), .F(\Data_Mem/n9394 ) );
  MUX \Data_Mem/U9452  ( .IN0(\Data_Mem/n9392 ), .IN1(\Data_Mem/n9391 ), .SEL(
        N28), .F(\Data_Mem/n9393 ) );
  MUX \Data_Mem/U9451  ( .IN0(o[1306]), .IN1(o[1338]), .SEL(N29), .F(
        \Data_Mem/n9392 ) );
  MUX \Data_Mem/U9450  ( .IN0(o[1370]), .IN1(o[1402]), .SEL(N29), .F(
        \Data_Mem/n9391 ) );
  MUX \Data_Mem/U9449  ( .IN0(\Data_Mem/n9389 ), .IN1(\Data_Mem/n9388 ), .SEL(
        N28), .F(\Data_Mem/n9390 ) );
  MUX \Data_Mem/U9448  ( .IN0(o[1434]), .IN1(o[1466]), .SEL(N29), .F(
        \Data_Mem/n9389 ) );
  MUX \Data_Mem/U9447  ( .IN0(o[1498]), .IN1(o[1530]), .SEL(N29), .F(
        \Data_Mem/n9388 ) );
  MUX \Data_Mem/U9446  ( .IN0(\Data_Mem/n9386 ), .IN1(\Data_Mem/n9379 ), .SEL(
        N26), .F(\Data_Mem/n9387 ) );
  MUX \Data_Mem/U9445  ( .IN0(\Data_Mem/n9385 ), .IN1(\Data_Mem/n9382 ), .SEL(
        N27), .F(\Data_Mem/n9386 ) );
  MUX \Data_Mem/U9444  ( .IN0(\Data_Mem/n9384 ), .IN1(\Data_Mem/n9383 ), .SEL(
        N28), .F(\Data_Mem/n9385 ) );
  MUX \Data_Mem/U9443  ( .IN0(o[1562]), .IN1(o[1594]), .SEL(N29), .F(
        \Data_Mem/n9384 ) );
  MUX \Data_Mem/U9442  ( .IN0(o[1626]), .IN1(o[1658]), .SEL(N29), .F(
        \Data_Mem/n9383 ) );
  MUX \Data_Mem/U9441  ( .IN0(\Data_Mem/n9381 ), .IN1(\Data_Mem/n9380 ), .SEL(
        N28), .F(\Data_Mem/n9382 ) );
  MUX \Data_Mem/U9440  ( .IN0(o[1690]), .IN1(o[1722]), .SEL(N29), .F(
        \Data_Mem/n9381 ) );
  MUX \Data_Mem/U9439  ( .IN0(o[1754]), .IN1(o[1786]), .SEL(N29), .F(
        \Data_Mem/n9380 ) );
  MUX \Data_Mem/U9438  ( .IN0(\Data_Mem/n9378 ), .IN1(\Data_Mem/n9375 ), .SEL(
        N27), .F(\Data_Mem/n9379 ) );
  MUX \Data_Mem/U9437  ( .IN0(\Data_Mem/n9377 ), .IN1(\Data_Mem/n9376 ), .SEL(
        N28), .F(\Data_Mem/n9378 ) );
  MUX \Data_Mem/U9436  ( .IN0(o[1818]), .IN1(o[1850]), .SEL(N29), .F(
        \Data_Mem/n9377 ) );
  MUX \Data_Mem/U9435  ( .IN0(o[1882]), .IN1(o[1914]), .SEL(N29), .F(
        \Data_Mem/n9376 ) );
  MUX \Data_Mem/U9434  ( .IN0(\Data_Mem/n9374 ), .IN1(\Data_Mem/n9373 ), .SEL(
        N28), .F(\Data_Mem/n9375 ) );
  MUX \Data_Mem/U9433  ( .IN0(o[1946]), .IN1(o[1978]), .SEL(N29), .F(
        \Data_Mem/n9374 ) );
  MUX \Data_Mem/U9432  ( .IN0(o[2010]), .IN1(o[2042]), .SEL(N29), .F(
        \Data_Mem/n9373 ) );
  MUX \Data_Mem/U9431  ( .IN0(\Data_Mem/n9372 ), .IN1(\Data_Mem/n9341 ), .SEL(
        N24), .F(\Data_Mem/N720 ) );
  MUX \Data_Mem/U9430  ( .IN0(\Data_Mem/n9371 ), .IN1(\Data_Mem/n9356 ), .SEL(
        N25), .F(\Data_Mem/n9372 ) );
  MUX \Data_Mem/U9429  ( .IN0(\Data_Mem/n9370 ), .IN1(\Data_Mem/n9363 ), .SEL(
        N26), .F(\Data_Mem/n9371 ) );
  MUX \Data_Mem/U9428  ( .IN0(\Data_Mem/n9369 ), .IN1(\Data_Mem/n9366 ), .SEL(
        N27), .F(\Data_Mem/n9370 ) );
  MUX \Data_Mem/U9427  ( .IN0(\Data_Mem/n9368 ), .IN1(\Data_Mem/n9367 ), .SEL(
        N28), .F(\Data_Mem/n9369 ) );
  MUX \Data_Mem/U9426  ( .IN0(o[25]), .IN1(o[57]), .SEL(N29), .F(
        \Data_Mem/n9368 ) );
  MUX \Data_Mem/U9425  ( .IN0(o[89]), .IN1(o[121]), .SEL(N29), .F(
        \Data_Mem/n9367 ) );
  MUX \Data_Mem/U9424  ( .IN0(\Data_Mem/n9365 ), .IN1(\Data_Mem/n9364 ), .SEL(
        N28), .F(\Data_Mem/n9366 ) );
  MUX \Data_Mem/U9423  ( .IN0(o[153]), .IN1(o[185]), .SEL(N29), .F(
        \Data_Mem/n9365 ) );
  MUX \Data_Mem/U9422  ( .IN0(o[217]), .IN1(o[249]), .SEL(N29), .F(
        \Data_Mem/n9364 ) );
  MUX \Data_Mem/U9421  ( .IN0(\Data_Mem/n9362 ), .IN1(\Data_Mem/n9359 ), .SEL(
        N27), .F(\Data_Mem/n9363 ) );
  MUX \Data_Mem/U9420  ( .IN0(\Data_Mem/n9361 ), .IN1(\Data_Mem/n9360 ), .SEL(
        N28), .F(\Data_Mem/n9362 ) );
  MUX \Data_Mem/U9419  ( .IN0(o[281]), .IN1(o[313]), .SEL(N29), .F(
        \Data_Mem/n9361 ) );
  MUX \Data_Mem/U9418  ( .IN0(o[345]), .IN1(o[377]), .SEL(N29), .F(
        \Data_Mem/n9360 ) );
  MUX \Data_Mem/U9417  ( .IN0(\Data_Mem/n9358 ), .IN1(\Data_Mem/n9357 ), .SEL(
        N28), .F(\Data_Mem/n9359 ) );
  MUX \Data_Mem/U9416  ( .IN0(o[409]), .IN1(o[441]), .SEL(N29), .F(
        \Data_Mem/n9358 ) );
  MUX \Data_Mem/U9415  ( .IN0(o[473]), .IN1(o[505]), .SEL(N29), .F(
        \Data_Mem/n9357 ) );
  MUX \Data_Mem/U9414  ( .IN0(\Data_Mem/n9355 ), .IN1(\Data_Mem/n9348 ), .SEL(
        N26), .F(\Data_Mem/n9356 ) );
  MUX \Data_Mem/U9413  ( .IN0(\Data_Mem/n9354 ), .IN1(\Data_Mem/n9351 ), .SEL(
        N27), .F(\Data_Mem/n9355 ) );
  MUX \Data_Mem/U9412  ( .IN0(\Data_Mem/n9353 ), .IN1(\Data_Mem/n9352 ), .SEL(
        N28), .F(\Data_Mem/n9354 ) );
  MUX \Data_Mem/U9411  ( .IN0(o[537]), .IN1(o[569]), .SEL(N29), .F(
        \Data_Mem/n9353 ) );
  MUX \Data_Mem/U9410  ( .IN0(o[601]), .IN1(o[633]), .SEL(N29), .F(
        \Data_Mem/n9352 ) );
  MUX \Data_Mem/U9409  ( .IN0(\Data_Mem/n9350 ), .IN1(\Data_Mem/n9349 ), .SEL(
        N28), .F(\Data_Mem/n9351 ) );
  MUX \Data_Mem/U9408  ( .IN0(o[665]), .IN1(o[697]), .SEL(N29), .F(
        \Data_Mem/n9350 ) );
  MUX \Data_Mem/U9407  ( .IN0(o[729]), .IN1(o[761]), .SEL(N29), .F(
        \Data_Mem/n9349 ) );
  MUX \Data_Mem/U9406  ( .IN0(\Data_Mem/n9347 ), .IN1(\Data_Mem/n9344 ), .SEL(
        N27), .F(\Data_Mem/n9348 ) );
  MUX \Data_Mem/U9405  ( .IN0(\Data_Mem/n9346 ), .IN1(\Data_Mem/n9345 ), .SEL(
        N28), .F(\Data_Mem/n9347 ) );
  MUX \Data_Mem/U9404  ( .IN0(o[793]), .IN1(o[825]), .SEL(N29), .F(
        \Data_Mem/n9346 ) );
  MUX \Data_Mem/U9403  ( .IN0(o[857]), .IN1(o[889]), .SEL(N29), .F(
        \Data_Mem/n9345 ) );
  MUX \Data_Mem/U9402  ( .IN0(\Data_Mem/n9343 ), .IN1(\Data_Mem/n9342 ), .SEL(
        N28), .F(\Data_Mem/n9344 ) );
  MUX \Data_Mem/U9401  ( .IN0(o[921]), .IN1(o[953]), .SEL(N29), .F(
        \Data_Mem/n9343 ) );
  MUX \Data_Mem/U9400  ( .IN0(o[985]), .IN1(o[1017]), .SEL(N29), .F(
        \Data_Mem/n9342 ) );
  MUX \Data_Mem/U9399  ( .IN0(\Data_Mem/n9340 ), .IN1(\Data_Mem/n9325 ), .SEL(
        N25), .F(\Data_Mem/n9341 ) );
  MUX \Data_Mem/U9398  ( .IN0(\Data_Mem/n9339 ), .IN1(\Data_Mem/n9332 ), .SEL(
        N26), .F(\Data_Mem/n9340 ) );
  MUX \Data_Mem/U9397  ( .IN0(\Data_Mem/n9338 ), .IN1(\Data_Mem/n9335 ), .SEL(
        N27), .F(\Data_Mem/n9339 ) );
  MUX \Data_Mem/U9396  ( .IN0(\Data_Mem/n9337 ), .IN1(\Data_Mem/n9336 ), .SEL(
        N28), .F(\Data_Mem/n9338 ) );
  MUX \Data_Mem/U9395  ( .IN0(o[1049]), .IN1(o[1081]), .SEL(N29), .F(
        \Data_Mem/n9337 ) );
  MUX \Data_Mem/U9394  ( .IN0(o[1113]), .IN1(o[1145]), .SEL(N29), .F(
        \Data_Mem/n9336 ) );
  MUX \Data_Mem/U9393  ( .IN0(\Data_Mem/n9334 ), .IN1(\Data_Mem/n9333 ), .SEL(
        N28), .F(\Data_Mem/n9335 ) );
  MUX \Data_Mem/U9392  ( .IN0(o[1177]), .IN1(o[1209]), .SEL(N29), .F(
        \Data_Mem/n9334 ) );
  MUX \Data_Mem/U9391  ( .IN0(o[1241]), .IN1(o[1273]), .SEL(N29), .F(
        \Data_Mem/n9333 ) );
  MUX \Data_Mem/U9390  ( .IN0(\Data_Mem/n9331 ), .IN1(\Data_Mem/n9328 ), .SEL(
        N27), .F(\Data_Mem/n9332 ) );
  MUX \Data_Mem/U9389  ( .IN0(\Data_Mem/n9330 ), .IN1(\Data_Mem/n9329 ), .SEL(
        N28), .F(\Data_Mem/n9331 ) );
  MUX \Data_Mem/U9388  ( .IN0(o[1305]), .IN1(o[1337]), .SEL(N29), .F(
        \Data_Mem/n9330 ) );
  MUX \Data_Mem/U9387  ( .IN0(o[1369]), .IN1(o[1401]), .SEL(N29), .F(
        \Data_Mem/n9329 ) );
  MUX \Data_Mem/U9386  ( .IN0(\Data_Mem/n9327 ), .IN1(\Data_Mem/n9326 ), .SEL(
        N28), .F(\Data_Mem/n9328 ) );
  MUX \Data_Mem/U9385  ( .IN0(o[1433]), .IN1(o[1465]), .SEL(N29), .F(
        \Data_Mem/n9327 ) );
  MUX \Data_Mem/U9384  ( .IN0(o[1497]), .IN1(o[1529]), .SEL(N29), .F(
        \Data_Mem/n9326 ) );
  MUX \Data_Mem/U9383  ( .IN0(\Data_Mem/n9324 ), .IN1(\Data_Mem/n9317 ), .SEL(
        N26), .F(\Data_Mem/n9325 ) );
  MUX \Data_Mem/U9382  ( .IN0(\Data_Mem/n9323 ), .IN1(\Data_Mem/n9320 ), .SEL(
        N27), .F(\Data_Mem/n9324 ) );
  MUX \Data_Mem/U9381  ( .IN0(\Data_Mem/n9322 ), .IN1(\Data_Mem/n9321 ), .SEL(
        N28), .F(\Data_Mem/n9323 ) );
  MUX \Data_Mem/U9380  ( .IN0(o[1561]), .IN1(o[1593]), .SEL(N29), .F(
        \Data_Mem/n9322 ) );
  MUX \Data_Mem/U9379  ( .IN0(o[1625]), .IN1(o[1657]), .SEL(N29), .F(
        \Data_Mem/n9321 ) );
  MUX \Data_Mem/U9378  ( .IN0(\Data_Mem/n9319 ), .IN1(\Data_Mem/n9318 ), .SEL(
        N28), .F(\Data_Mem/n9320 ) );
  MUX \Data_Mem/U9377  ( .IN0(o[1689]), .IN1(o[1721]), .SEL(N29), .F(
        \Data_Mem/n9319 ) );
  MUX \Data_Mem/U9376  ( .IN0(o[1753]), .IN1(o[1785]), .SEL(N29), .F(
        \Data_Mem/n9318 ) );
  MUX \Data_Mem/U9375  ( .IN0(\Data_Mem/n9316 ), .IN1(\Data_Mem/n9313 ), .SEL(
        N27), .F(\Data_Mem/n9317 ) );
  MUX \Data_Mem/U9374  ( .IN0(\Data_Mem/n9315 ), .IN1(\Data_Mem/n9314 ), .SEL(
        N28), .F(\Data_Mem/n9316 ) );
  MUX \Data_Mem/U9373  ( .IN0(o[1817]), .IN1(o[1849]), .SEL(N29), .F(
        \Data_Mem/n9315 ) );
  MUX \Data_Mem/U9372  ( .IN0(o[1881]), .IN1(o[1913]), .SEL(N29), .F(
        \Data_Mem/n9314 ) );
  MUX \Data_Mem/U9371  ( .IN0(\Data_Mem/n9312 ), .IN1(\Data_Mem/n9311 ), .SEL(
        N28), .F(\Data_Mem/n9313 ) );
  MUX \Data_Mem/U9370  ( .IN0(o[1945]), .IN1(o[1977]), .SEL(N29), .F(
        \Data_Mem/n9312 ) );
  MUX \Data_Mem/U9369  ( .IN0(o[2009]), .IN1(o[2041]), .SEL(N29), .F(
        \Data_Mem/n9311 ) );
  MUX \Data_Mem/U9368  ( .IN0(\Data_Mem/n9310 ), .IN1(\Data_Mem/n9279 ), .SEL(
        N24), .F(\Data_Mem/N721 ) );
  MUX \Data_Mem/U9367  ( .IN0(\Data_Mem/n9309 ), .IN1(\Data_Mem/n9294 ), .SEL(
        N25), .F(\Data_Mem/n9310 ) );
  MUX \Data_Mem/U9366  ( .IN0(\Data_Mem/n9308 ), .IN1(\Data_Mem/n9301 ), .SEL(
        N26), .F(\Data_Mem/n9309 ) );
  MUX \Data_Mem/U9365  ( .IN0(\Data_Mem/n9307 ), .IN1(\Data_Mem/n9304 ), .SEL(
        N27), .F(\Data_Mem/n9308 ) );
  MUX \Data_Mem/U9364  ( .IN0(\Data_Mem/n9306 ), .IN1(\Data_Mem/n9305 ), .SEL(
        N28), .F(\Data_Mem/n9307 ) );
  MUX \Data_Mem/U9363  ( .IN0(o[24]), .IN1(o[56]), .SEL(N29), .F(
        \Data_Mem/n9306 ) );
  MUX \Data_Mem/U9362  ( .IN0(o[88]), .IN1(o[120]), .SEL(N29), .F(
        \Data_Mem/n9305 ) );
  MUX \Data_Mem/U9361  ( .IN0(\Data_Mem/n9303 ), .IN1(\Data_Mem/n9302 ), .SEL(
        N28), .F(\Data_Mem/n9304 ) );
  MUX \Data_Mem/U9360  ( .IN0(o[152]), .IN1(o[184]), .SEL(N29), .F(
        \Data_Mem/n9303 ) );
  MUX \Data_Mem/U9359  ( .IN0(o[216]), .IN1(o[248]), .SEL(N29), .F(
        \Data_Mem/n9302 ) );
  MUX \Data_Mem/U9358  ( .IN0(\Data_Mem/n9300 ), .IN1(\Data_Mem/n9297 ), .SEL(
        N27), .F(\Data_Mem/n9301 ) );
  MUX \Data_Mem/U9357  ( .IN0(\Data_Mem/n9299 ), .IN1(\Data_Mem/n9298 ), .SEL(
        N28), .F(\Data_Mem/n9300 ) );
  MUX \Data_Mem/U9356  ( .IN0(o[280]), .IN1(o[312]), .SEL(N29), .F(
        \Data_Mem/n9299 ) );
  MUX \Data_Mem/U9355  ( .IN0(o[344]), .IN1(o[376]), .SEL(N29), .F(
        \Data_Mem/n9298 ) );
  MUX \Data_Mem/U9354  ( .IN0(\Data_Mem/n9296 ), .IN1(\Data_Mem/n9295 ), .SEL(
        N28), .F(\Data_Mem/n9297 ) );
  MUX \Data_Mem/U9353  ( .IN0(o[408]), .IN1(o[440]), .SEL(N29), .F(
        \Data_Mem/n9296 ) );
  MUX \Data_Mem/U9352  ( .IN0(o[472]), .IN1(o[504]), .SEL(N29), .F(
        \Data_Mem/n9295 ) );
  MUX \Data_Mem/U9351  ( .IN0(\Data_Mem/n9293 ), .IN1(\Data_Mem/n9286 ), .SEL(
        N26), .F(\Data_Mem/n9294 ) );
  MUX \Data_Mem/U9350  ( .IN0(\Data_Mem/n9292 ), .IN1(\Data_Mem/n9289 ), .SEL(
        N27), .F(\Data_Mem/n9293 ) );
  MUX \Data_Mem/U9349  ( .IN0(\Data_Mem/n9291 ), .IN1(\Data_Mem/n9290 ), .SEL(
        N28), .F(\Data_Mem/n9292 ) );
  MUX \Data_Mem/U9348  ( .IN0(o[536]), .IN1(o[568]), .SEL(N29), .F(
        \Data_Mem/n9291 ) );
  MUX \Data_Mem/U9347  ( .IN0(o[600]), .IN1(o[632]), .SEL(N29), .F(
        \Data_Mem/n9290 ) );
  MUX \Data_Mem/U9346  ( .IN0(\Data_Mem/n9288 ), .IN1(\Data_Mem/n9287 ), .SEL(
        N28), .F(\Data_Mem/n9289 ) );
  MUX \Data_Mem/U9345  ( .IN0(o[664]), .IN1(o[696]), .SEL(N29), .F(
        \Data_Mem/n9288 ) );
  MUX \Data_Mem/U9344  ( .IN0(o[728]), .IN1(o[760]), .SEL(N29), .F(
        \Data_Mem/n9287 ) );
  MUX \Data_Mem/U9343  ( .IN0(\Data_Mem/n9285 ), .IN1(\Data_Mem/n9282 ), .SEL(
        N27), .F(\Data_Mem/n9286 ) );
  MUX \Data_Mem/U9342  ( .IN0(\Data_Mem/n9284 ), .IN1(\Data_Mem/n9283 ), .SEL(
        N28), .F(\Data_Mem/n9285 ) );
  MUX \Data_Mem/U9341  ( .IN0(o[792]), .IN1(o[824]), .SEL(N29), .F(
        \Data_Mem/n9284 ) );
  MUX \Data_Mem/U9340  ( .IN0(o[856]), .IN1(o[888]), .SEL(N29), .F(
        \Data_Mem/n9283 ) );
  MUX \Data_Mem/U9339  ( .IN0(\Data_Mem/n9281 ), .IN1(\Data_Mem/n9280 ), .SEL(
        N28), .F(\Data_Mem/n9282 ) );
  MUX \Data_Mem/U9338  ( .IN0(o[920]), .IN1(o[952]), .SEL(N29), .F(
        \Data_Mem/n9281 ) );
  MUX \Data_Mem/U9337  ( .IN0(o[984]), .IN1(o[1016]), .SEL(N29), .F(
        \Data_Mem/n9280 ) );
  MUX \Data_Mem/U9336  ( .IN0(\Data_Mem/n9278 ), .IN1(\Data_Mem/n9263 ), .SEL(
        N25), .F(\Data_Mem/n9279 ) );
  MUX \Data_Mem/U9335  ( .IN0(\Data_Mem/n9277 ), .IN1(\Data_Mem/n9270 ), .SEL(
        N26), .F(\Data_Mem/n9278 ) );
  MUX \Data_Mem/U9334  ( .IN0(\Data_Mem/n9276 ), .IN1(\Data_Mem/n9273 ), .SEL(
        N27), .F(\Data_Mem/n9277 ) );
  MUX \Data_Mem/U9333  ( .IN0(\Data_Mem/n9275 ), .IN1(\Data_Mem/n9274 ), .SEL(
        N28), .F(\Data_Mem/n9276 ) );
  MUX \Data_Mem/U9332  ( .IN0(o[1048]), .IN1(o[1080]), .SEL(N29), .F(
        \Data_Mem/n9275 ) );
  MUX \Data_Mem/U9331  ( .IN0(o[1112]), .IN1(o[1144]), .SEL(N29), .F(
        \Data_Mem/n9274 ) );
  MUX \Data_Mem/U9330  ( .IN0(\Data_Mem/n9272 ), .IN1(\Data_Mem/n9271 ), .SEL(
        N28), .F(\Data_Mem/n9273 ) );
  MUX \Data_Mem/U9329  ( .IN0(o[1176]), .IN1(o[1208]), .SEL(N29), .F(
        \Data_Mem/n9272 ) );
  MUX \Data_Mem/U9328  ( .IN0(o[1240]), .IN1(o[1272]), .SEL(N29), .F(
        \Data_Mem/n9271 ) );
  MUX \Data_Mem/U9327  ( .IN0(\Data_Mem/n9269 ), .IN1(\Data_Mem/n9266 ), .SEL(
        N27), .F(\Data_Mem/n9270 ) );
  MUX \Data_Mem/U9326  ( .IN0(\Data_Mem/n9268 ), .IN1(\Data_Mem/n9267 ), .SEL(
        N28), .F(\Data_Mem/n9269 ) );
  MUX \Data_Mem/U9325  ( .IN0(o[1304]), .IN1(o[1336]), .SEL(N29), .F(
        \Data_Mem/n9268 ) );
  MUX \Data_Mem/U9324  ( .IN0(o[1368]), .IN1(o[1400]), .SEL(N29), .F(
        \Data_Mem/n9267 ) );
  MUX \Data_Mem/U9323  ( .IN0(\Data_Mem/n9265 ), .IN1(\Data_Mem/n9264 ), .SEL(
        N28), .F(\Data_Mem/n9266 ) );
  MUX \Data_Mem/U9322  ( .IN0(o[1432]), .IN1(o[1464]), .SEL(N29), .F(
        \Data_Mem/n9265 ) );
  MUX \Data_Mem/U9321  ( .IN0(o[1496]), .IN1(o[1528]), .SEL(N29), .F(
        \Data_Mem/n9264 ) );
  MUX \Data_Mem/U9320  ( .IN0(\Data_Mem/n9262 ), .IN1(\Data_Mem/n9255 ), .SEL(
        N26), .F(\Data_Mem/n9263 ) );
  MUX \Data_Mem/U9319  ( .IN0(\Data_Mem/n9261 ), .IN1(\Data_Mem/n9258 ), .SEL(
        N27), .F(\Data_Mem/n9262 ) );
  MUX \Data_Mem/U9318  ( .IN0(\Data_Mem/n9260 ), .IN1(\Data_Mem/n9259 ), .SEL(
        N28), .F(\Data_Mem/n9261 ) );
  MUX \Data_Mem/U9317  ( .IN0(o[1560]), .IN1(o[1592]), .SEL(N29), .F(
        \Data_Mem/n9260 ) );
  MUX \Data_Mem/U9316  ( .IN0(o[1624]), .IN1(o[1656]), .SEL(N29), .F(
        \Data_Mem/n9259 ) );
  MUX \Data_Mem/U9315  ( .IN0(\Data_Mem/n9257 ), .IN1(\Data_Mem/n9256 ), .SEL(
        N28), .F(\Data_Mem/n9258 ) );
  MUX \Data_Mem/U9314  ( .IN0(o[1688]), .IN1(o[1720]), .SEL(N29), .F(
        \Data_Mem/n9257 ) );
  MUX \Data_Mem/U9313  ( .IN0(o[1752]), .IN1(o[1784]), .SEL(N29), .F(
        \Data_Mem/n9256 ) );
  MUX \Data_Mem/U9312  ( .IN0(\Data_Mem/n9254 ), .IN1(\Data_Mem/n9251 ), .SEL(
        N27), .F(\Data_Mem/n9255 ) );
  MUX \Data_Mem/U9311  ( .IN0(\Data_Mem/n9253 ), .IN1(\Data_Mem/n9252 ), .SEL(
        N28), .F(\Data_Mem/n9254 ) );
  MUX \Data_Mem/U9310  ( .IN0(o[1816]), .IN1(o[1848]), .SEL(N29), .F(
        \Data_Mem/n9253 ) );
  MUX \Data_Mem/U9309  ( .IN0(o[1880]), .IN1(o[1912]), .SEL(N29), .F(
        \Data_Mem/n9252 ) );
  MUX \Data_Mem/U9308  ( .IN0(\Data_Mem/n9250 ), .IN1(\Data_Mem/n9249 ), .SEL(
        N28), .F(\Data_Mem/n9251 ) );
  MUX \Data_Mem/U9307  ( .IN0(o[1944]), .IN1(o[1976]), .SEL(N29), .F(
        \Data_Mem/n9250 ) );
  MUX \Data_Mem/U9306  ( .IN0(o[2008]), .IN1(o[2040]), .SEL(N29), .F(
        \Data_Mem/n9249 ) );
  MUX \Data_Mem/U9305  ( .IN0(\Data_Mem/n9248 ), .IN1(\Data_Mem/n9217 ), .SEL(
        N24), .F(\Data_Mem/N722 ) );
  MUX \Data_Mem/U9304  ( .IN0(\Data_Mem/n9247 ), .IN1(\Data_Mem/n9232 ), .SEL(
        N25), .F(\Data_Mem/n9248 ) );
  MUX \Data_Mem/U9303  ( .IN0(\Data_Mem/n9246 ), .IN1(\Data_Mem/n9239 ), .SEL(
        N26), .F(\Data_Mem/n9247 ) );
  MUX \Data_Mem/U9302  ( .IN0(\Data_Mem/n9245 ), .IN1(\Data_Mem/n9242 ), .SEL(
        N27), .F(\Data_Mem/n9246 ) );
  MUX \Data_Mem/U9301  ( .IN0(\Data_Mem/n9244 ), .IN1(\Data_Mem/n9243 ), .SEL(
        N28), .F(\Data_Mem/n9245 ) );
  MUX \Data_Mem/U9300  ( .IN0(o[23]), .IN1(o[55]), .SEL(N29), .F(
        \Data_Mem/n9244 ) );
  MUX \Data_Mem/U9299  ( .IN0(o[87]), .IN1(o[119]), .SEL(N29), .F(
        \Data_Mem/n9243 ) );
  MUX \Data_Mem/U9298  ( .IN0(\Data_Mem/n9241 ), .IN1(\Data_Mem/n9240 ), .SEL(
        N28), .F(\Data_Mem/n9242 ) );
  MUX \Data_Mem/U9297  ( .IN0(o[151]), .IN1(o[183]), .SEL(N29), .F(
        \Data_Mem/n9241 ) );
  MUX \Data_Mem/U9296  ( .IN0(o[215]), .IN1(o[247]), .SEL(N29), .F(
        \Data_Mem/n9240 ) );
  MUX \Data_Mem/U9295  ( .IN0(\Data_Mem/n9238 ), .IN1(\Data_Mem/n9235 ), .SEL(
        N27), .F(\Data_Mem/n9239 ) );
  MUX \Data_Mem/U9294  ( .IN0(\Data_Mem/n9237 ), .IN1(\Data_Mem/n9236 ), .SEL(
        N28), .F(\Data_Mem/n9238 ) );
  MUX \Data_Mem/U9293  ( .IN0(o[279]), .IN1(o[311]), .SEL(N29), .F(
        \Data_Mem/n9237 ) );
  MUX \Data_Mem/U9292  ( .IN0(o[343]), .IN1(o[375]), .SEL(N29), .F(
        \Data_Mem/n9236 ) );
  MUX \Data_Mem/U9291  ( .IN0(\Data_Mem/n9234 ), .IN1(\Data_Mem/n9233 ), .SEL(
        N28), .F(\Data_Mem/n9235 ) );
  MUX \Data_Mem/U9290  ( .IN0(o[407]), .IN1(o[439]), .SEL(N29), .F(
        \Data_Mem/n9234 ) );
  MUX \Data_Mem/U9289  ( .IN0(o[471]), .IN1(o[503]), .SEL(N29), .F(
        \Data_Mem/n9233 ) );
  MUX \Data_Mem/U9288  ( .IN0(\Data_Mem/n9231 ), .IN1(\Data_Mem/n9224 ), .SEL(
        N26), .F(\Data_Mem/n9232 ) );
  MUX \Data_Mem/U9287  ( .IN0(\Data_Mem/n9230 ), .IN1(\Data_Mem/n9227 ), .SEL(
        N27), .F(\Data_Mem/n9231 ) );
  MUX \Data_Mem/U9286  ( .IN0(\Data_Mem/n9229 ), .IN1(\Data_Mem/n9228 ), .SEL(
        N28), .F(\Data_Mem/n9230 ) );
  MUX \Data_Mem/U9285  ( .IN0(o[535]), .IN1(o[567]), .SEL(N29), .F(
        \Data_Mem/n9229 ) );
  MUX \Data_Mem/U9284  ( .IN0(o[599]), .IN1(o[631]), .SEL(N29), .F(
        \Data_Mem/n9228 ) );
  MUX \Data_Mem/U9283  ( .IN0(\Data_Mem/n9226 ), .IN1(\Data_Mem/n9225 ), .SEL(
        N28), .F(\Data_Mem/n9227 ) );
  MUX \Data_Mem/U9282  ( .IN0(o[663]), .IN1(o[695]), .SEL(N29), .F(
        \Data_Mem/n9226 ) );
  MUX \Data_Mem/U9281  ( .IN0(o[727]), .IN1(o[759]), .SEL(N29), .F(
        \Data_Mem/n9225 ) );
  MUX \Data_Mem/U9280  ( .IN0(\Data_Mem/n9223 ), .IN1(\Data_Mem/n9220 ), .SEL(
        N27), .F(\Data_Mem/n9224 ) );
  MUX \Data_Mem/U9279  ( .IN0(\Data_Mem/n9222 ), .IN1(\Data_Mem/n9221 ), .SEL(
        N28), .F(\Data_Mem/n9223 ) );
  MUX \Data_Mem/U9278  ( .IN0(o[791]), .IN1(o[823]), .SEL(N29), .F(
        \Data_Mem/n9222 ) );
  MUX \Data_Mem/U9277  ( .IN0(o[855]), .IN1(o[887]), .SEL(N29), .F(
        \Data_Mem/n9221 ) );
  MUX \Data_Mem/U9276  ( .IN0(\Data_Mem/n9219 ), .IN1(\Data_Mem/n9218 ), .SEL(
        N28), .F(\Data_Mem/n9220 ) );
  MUX \Data_Mem/U9275  ( .IN0(o[919]), .IN1(o[951]), .SEL(N29), .F(
        \Data_Mem/n9219 ) );
  MUX \Data_Mem/U9274  ( .IN0(o[983]), .IN1(o[1015]), .SEL(N29), .F(
        \Data_Mem/n9218 ) );
  MUX \Data_Mem/U9273  ( .IN0(\Data_Mem/n9216 ), .IN1(\Data_Mem/n9201 ), .SEL(
        N25), .F(\Data_Mem/n9217 ) );
  MUX \Data_Mem/U9272  ( .IN0(\Data_Mem/n9215 ), .IN1(\Data_Mem/n9208 ), .SEL(
        N26), .F(\Data_Mem/n9216 ) );
  MUX \Data_Mem/U9271  ( .IN0(\Data_Mem/n9214 ), .IN1(\Data_Mem/n9211 ), .SEL(
        N27), .F(\Data_Mem/n9215 ) );
  MUX \Data_Mem/U9270  ( .IN0(\Data_Mem/n9213 ), .IN1(\Data_Mem/n9212 ), .SEL(
        N28), .F(\Data_Mem/n9214 ) );
  MUX \Data_Mem/U9269  ( .IN0(o[1047]), .IN1(o[1079]), .SEL(N29), .F(
        \Data_Mem/n9213 ) );
  MUX \Data_Mem/U9268  ( .IN0(o[1111]), .IN1(o[1143]), .SEL(N29), .F(
        \Data_Mem/n9212 ) );
  MUX \Data_Mem/U9267  ( .IN0(\Data_Mem/n9210 ), .IN1(\Data_Mem/n9209 ), .SEL(
        N28), .F(\Data_Mem/n9211 ) );
  MUX \Data_Mem/U9266  ( .IN0(o[1175]), .IN1(o[1207]), .SEL(N29), .F(
        \Data_Mem/n9210 ) );
  MUX \Data_Mem/U9265  ( .IN0(o[1239]), .IN1(o[1271]), .SEL(N29), .F(
        \Data_Mem/n9209 ) );
  MUX \Data_Mem/U9264  ( .IN0(\Data_Mem/n9207 ), .IN1(\Data_Mem/n9204 ), .SEL(
        N27), .F(\Data_Mem/n9208 ) );
  MUX \Data_Mem/U9263  ( .IN0(\Data_Mem/n9206 ), .IN1(\Data_Mem/n9205 ), .SEL(
        N28), .F(\Data_Mem/n9207 ) );
  MUX \Data_Mem/U9262  ( .IN0(o[1303]), .IN1(o[1335]), .SEL(N29), .F(
        \Data_Mem/n9206 ) );
  MUX \Data_Mem/U9261  ( .IN0(o[1367]), .IN1(o[1399]), .SEL(N29), .F(
        \Data_Mem/n9205 ) );
  MUX \Data_Mem/U9260  ( .IN0(\Data_Mem/n9203 ), .IN1(\Data_Mem/n9202 ), .SEL(
        N28), .F(\Data_Mem/n9204 ) );
  MUX \Data_Mem/U9259  ( .IN0(o[1431]), .IN1(o[1463]), .SEL(N29), .F(
        \Data_Mem/n9203 ) );
  MUX \Data_Mem/U9258  ( .IN0(o[1495]), .IN1(o[1527]), .SEL(N29), .F(
        \Data_Mem/n9202 ) );
  MUX \Data_Mem/U9257  ( .IN0(\Data_Mem/n9200 ), .IN1(\Data_Mem/n9193 ), .SEL(
        N26), .F(\Data_Mem/n9201 ) );
  MUX \Data_Mem/U9256  ( .IN0(\Data_Mem/n9199 ), .IN1(\Data_Mem/n9196 ), .SEL(
        N27), .F(\Data_Mem/n9200 ) );
  MUX \Data_Mem/U9255  ( .IN0(\Data_Mem/n9198 ), .IN1(\Data_Mem/n9197 ), .SEL(
        N28), .F(\Data_Mem/n9199 ) );
  MUX \Data_Mem/U9254  ( .IN0(o[1559]), .IN1(o[1591]), .SEL(N29), .F(
        \Data_Mem/n9198 ) );
  MUX \Data_Mem/U9253  ( .IN0(o[1623]), .IN1(o[1655]), .SEL(N29), .F(
        \Data_Mem/n9197 ) );
  MUX \Data_Mem/U9252  ( .IN0(\Data_Mem/n9195 ), .IN1(\Data_Mem/n9194 ), .SEL(
        N28), .F(\Data_Mem/n9196 ) );
  MUX \Data_Mem/U9251  ( .IN0(o[1687]), .IN1(o[1719]), .SEL(N29), .F(
        \Data_Mem/n9195 ) );
  MUX \Data_Mem/U9250  ( .IN0(o[1751]), .IN1(o[1783]), .SEL(N29), .F(
        \Data_Mem/n9194 ) );
  MUX \Data_Mem/U9249  ( .IN0(\Data_Mem/n9192 ), .IN1(\Data_Mem/n9189 ), .SEL(
        N27), .F(\Data_Mem/n9193 ) );
  MUX \Data_Mem/U9248  ( .IN0(\Data_Mem/n9191 ), .IN1(\Data_Mem/n9190 ), .SEL(
        N28), .F(\Data_Mem/n9192 ) );
  MUX \Data_Mem/U9247  ( .IN0(o[1815]), .IN1(o[1847]), .SEL(N29), .F(
        \Data_Mem/n9191 ) );
  MUX \Data_Mem/U9246  ( .IN0(o[1879]), .IN1(o[1911]), .SEL(N29), .F(
        \Data_Mem/n9190 ) );
  MUX \Data_Mem/U9245  ( .IN0(\Data_Mem/n9188 ), .IN1(\Data_Mem/n9187 ), .SEL(
        N28), .F(\Data_Mem/n9189 ) );
  MUX \Data_Mem/U9244  ( .IN0(o[1943]), .IN1(o[1975]), .SEL(N29), .F(
        \Data_Mem/n9188 ) );
  MUX \Data_Mem/U9243  ( .IN0(o[2007]), .IN1(o[2039]), .SEL(N29), .F(
        \Data_Mem/n9187 ) );
  MUX \Data_Mem/U9242  ( .IN0(\Data_Mem/n9186 ), .IN1(\Data_Mem/n9155 ), .SEL(
        N24), .F(\Data_Mem/N723 ) );
  MUX \Data_Mem/U9241  ( .IN0(\Data_Mem/n9185 ), .IN1(\Data_Mem/n9170 ), .SEL(
        N25), .F(\Data_Mem/n9186 ) );
  MUX \Data_Mem/U9240  ( .IN0(\Data_Mem/n9184 ), .IN1(\Data_Mem/n9177 ), .SEL(
        N26), .F(\Data_Mem/n9185 ) );
  MUX \Data_Mem/U9239  ( .IN0(\Data_Mem/n9183 ), .IN1(\Data_Mem/n9180 ), .SEL(
        N27), .F(\Data_Mem/n9184 ) );
  MUX \Data_Mem/U9238  ( .IN0(\Data_Mem/n9182 ), .IN1(\Data_Mem/n9181 ), .SEL(
        N28), .F(\Data_Mem/n9183 ) );
  MUX \Data_Mem/U9237  ( .IN0(o[22]), .IN1(o[54]), .SEL(N29), .F(
        \Data_Mem/n9182 ) );
  MUX \Data_Mem/U9236  ( .IN0(o[86]), .IN1(o[118]), .SEL(N29), .F(
        \Data_Mem/n9181 ) );
  MUX \Data_Mem/U9235  ( .IN0(\Data_Mem/n9179 ), .IN1(\Data_Mem/n9178 ), .SEL(
        N28), .F(\Data_Mem/n9180 ) );
  MUX \Data_Mem/U9234  ( .IN0(o[150]), .IN1(o[182]), .SEL(N29), .F(
        \Data_Mem/n9179 ) );
  MUX \Data_Mem/U9233  ( .IN0(o[214]), .IN1(o[246]), .SEL(N29), .F(
        \Data_Mem/n9178 ) );
  MUX \Data_Mem/U9232  ( .IN0(\Data_Mem/n9176 ), .IN1(\Data_Mem/n9173 ), .SEL(
        N27), .F(\Data_Mem/n9177 ) );
  MUX \Data_Mem/U9231  ( .IN0(\Data_Mem/n9175 ), .IN1(\Data_Mem/n9174 ), .SEL(
        N28), .F(\Data_Mem/n9176 ) );
  MUX \Data_Mem/U9230  ( .IN0(o[278]), .IN1(o[310]), .SEL(N29), .F(
        \Data_Mem/n9175 ) );
  MUX \Data_Mem/U9229  ( .IN0(o[342]), .IN1(o[374]), .SEL(N29), .F(
        \Data_Mem/n9174 ) );
  MUX \Data_Mem/U9228  ( .IN0(\Data_Mem/n9172 ), .IN1(\Data_Mem/n9171 ), .SEL(
        N28), .F(\Data_Mem/n9173 ) );
  MUX \Data_Mem/U9227  ( .IN0(o[406]), .IN1(o[438]), .SEL(N29), .F(
        \Data_Mem/n9172 ) );
  MUX \Data_Mem/U9226  ( .IN0(o[470]), .IN1(o[502]), .SEL(N29), .F(
        \Data_Mem/n9171 ) );
  MUX \Data_Mem/U9225  ( .IN0(\Data_Mem/n9169 ), .IN1(\Data_Mem/n9162 ), .SEL(
        N26), .F(\Data_Mem/n9170 ) );
  MUX \Data_Mem/U9224  ( .IN0(\Data_Mem/n9168 ), .IN1(\Data_Mem/n9165 ), .SEL(
        N27), .F(\Data_Mem/n9169 ) );
  MUX \Data_Mem/U9223  ( .IN0(\Data_Mem/n9167 ), .IN1(\Data_Mem/n9166 ), .SEL(
        N28), .F(\Data_Mem/n9168 ) );
  MUX \Data_Mem/U9222  ( .IN0(o[534]), .IN1(o[566]), .SEL(N29), .F(
        \Data_Mem/n9167 ) );
  MUX \Data_Mem/U9221  ( .IN0(o[598]), .IN1(o[630]), .SEL(N29), .F(
        \Data_Mem/n9166 ) );
  MUX \Data_Mem/U9220  ( .IN0(\Data_Mem/n9164 ), .IN1(\Data_Mem/n9163 ), .SEL(
        N28), .F(\Data_Mem/n9165 ) );
  MUX \Data_Mem/U9219  ( .IN0(o[662]), .IN1(o[694]), .SEL(N29), .F(
        \Data_Mem/n9164 ) );
  MUX \Data_Mem/U9218  ( .IN0(o[726]), .IN1(o[758]), .SEL(N29), .F(
        \Data_Mem/n9163 ) );
  MUX \Data_Mem/U9217  ( .IN0(\Data_Mem/n9161 ), .IN1(\Data_Mem/n9158 ), .SEL(
        N27), .F(\Data_Mem/n9162 ) );
  MUX \Data_Mem/U9216  ( .IN0(\Data_Mem/n9160 ), .IN1(\Data_Mem/n9159 ), .SEL(
        N28), .F(\Data_Mem/n9161 ) );
  MUX \Data_Mem/U9215  ( .IN0(o[790]), .IN1(o[822]), .SEL(N29), .F(
        \Data_Mem/n9160 ) );
  MUX \Data_Mem/U9214  ( .IN0(o[854]), .IN1(o[886]), .SEL(N29), .F(
        \Data_Mem/n9159 ) );
  MUX \Data_Mem/U9213  ( .IN0(\Data_Mem/n9157 ), .IN1(\Data_Mem/n9156 ), .SEL(
        N28), .F(\Data_Mem/n9158 ) );
  MUX \Data_Mem/U9212  ( .IN0(o[918]), .IN1(o[950]), .SEL(N29), .F(
        \Data_Mem/n9157 ) );
  MUX \Data_Mem/U9211  ( .IN0(o[982]), .IN1(o[1014]), .SEL(N29), .F(
        \Data_Mem/n9156 ) );
  MUX \Data_Mem/U9210  ( .IN0(\Data_Mem/n9154 ), .IN1(\Data_Mem/n9139 ), .SEL(
        N25), .F(\Data_Mem/n9155 ) );
  MUX \Data_Mem/U9209  ( .IN0(\Data_Mem/n9153 ), .IN1(\Data_Mem/n9146 ), .SEL(
        N26), .F(\Data_Mem/n9154 ) );
  MUX \Data_Mem/U9208  ( .IN0(\Data_Mem/n9152 ), .IN1(\Data_Mem/n9149 ), .SEL(
        N27), .F(\Data_Mem/n9153 ) );
  MUX \Data_Mem/U9207  ( .IN0(\Data_Mem/n9151 ), .IN1(\Data_Mem/n9150 ), .SEL(
        N28), .F(\Data_Mem/n9152 ) );
  MUX \Data_Mem/U9206  ( .IN0(o[1046]), .IN1(o[1078]), .SEL(N29), .F(
        \Data_Mem/n9151 ) );
  MUX \Data_Mem/U9205  ( .IN0(o[1110]), .IN1(o[1142]), .SEL(N29), .F(
        \Data_Mem/n9150 ) );
  MUX \Data_Mem/U9204  ( .IN0(\Data_Mem/n9148 ), .IN1(\Data_Mem/n9147 ), .SEL(
        N28), .F(\Data_Mem/n9149 ) );
  MUX \Data_Mem/U9203  ( .IN0(o[1174]), .IN1(o[1206]), .SEL(N29), .F(
        \Data_Mem/n9148 ) );
  MUX \Data_Mem/U9202  ( .IN0(o[1238]), .IN1(o[1270]), .SEL(N29), .F(
        \Data_Mem/n9147 ) );
  MUX \Data_Mem/U9201  ( .IN0(\Data_Mem/n9145 ), .IN1(\Data_Mem/n9142 ), .SEL(
        N27), .F(\Data_Mem/n9146 ) );
  MUX \Data_Mem/U9200  ( .IN0(\Data_Mem/n9144 ), .IN1(\Data_Mem/n9143 ), .SEL(
        N28), .F(\Data_Mem/n9145 ) );
  MUX \Data_Mem/U9199  ( .IN0(o[1302]), .IN1(o[1334]), .SEL(N29), .F(
        \Data_Mem/n9144 ) );
  MUX \Data_Mem/U9198  ( .IN0(o[1366]), .IN1(o[1398]), .SEL(N29), .F(
        \Data_Mem/n9143 ) );
  MUX \Data_Mem/U9197  ( .IN0(\Data_Mem/n9141 ), .IN1(\Data_Mem/n9140 ), .SEL(
        N28), .F(\Data_Mem/n9142 ) );
  MUX \Data_Mem/U9196  ( .IN0(o[1430]), .IN1(o[1462]), .SEL(N29), .F(
        \Data_Mem/n9141 ) );
  MUX \Data_Mem/U9195  ( .IN0(o[1494]), .IN1(o[1526]), .SEL(N29), .F(
        \Data_Mem/n9140 ) );
  MUX \Data_Mem/U9194  ( .IN0(\Data_Mem/n9138 ), .IN1(\Data_Mem/n9131 ), .SEL(
        N26), .F(\Data_Mem/n9139 ) );
  MUX \Data_Mem/U9193  ( .IN0(\Data_Mem/n9137 ), .IN1(\Data_Mem/n9134 ), .SEL(
        N27), .F(\Data_Mem/n9138 ) );
  MUX \Data_Mem/U9192  ( .IN0(\Data_Mem/n9136 ), .IN1(\Data_Mem/n9135 ), .SEL(
        N28), .F(\Data_Mem/n9137 ) );
  MUX \Data_Mem/U9191  ( .IN0(o[1558]), .IN1(o[1590]), .SEL(N29), .F(
        \Data_Mem/n9136 ) );
  MUX \Data_Mem/U9190  ( .IN0(o[1622]), .IN1(o[1654]), .SEL(N29), .F(
        \Data_Mem/n9135 ) );
  MUX \Data_Mem/U9189  ( .IN0(\Data_Mem/n9133 ), .IN1(\Data_Mem/n9132 ), .SEL(
        N28), .F(\Data_Mem/n9134 ) );
  MUX \Data_Mem/U9188  ( .IN0(o[1686]), .IN1(o[1718]), .SEL(N29), .F(
        \Data_Mem/n9133 ) );
  MUX \Data_Mem/U9187  ( .IN0(o[1750]), .IN1(o[1782]), .SEL(N29), .F(
        \Data_Mem/n9132 ) );
  MUX \Data_Mem/U9186  ( .IN0(\Data_Mem/n9130 ), .IN1(\Data_Mem/n9127 ), .SEL(
        N27), .F(\Data_Mem/n9131 ) );
  MUX \Data_Mem/U9185  ( .IN0(\Data_Mem/n9129 ), .IN1(\Data_Mem/n9128 ), .SEL(
        N28), .F(\Data_Mem/n9130 ) );
  MUX \Data_Mem/U9184  ( .IN0(o[1814]), .IN1(o[1846]), .SEL(N29), .F(
        \Data_Mem/n9129 ) );
  MUX \Data_Mem/U9183  ( .IN0(o[1878]), .IN1(o[1910]), .SEL(N29), .F(
        \Data_Mem/n9128 ) );
  MUX \Data_Mem/U9182  ( .IN0(\Data_Mem/n9126 ), .IN1(\Data_Mem/n9125 ), .SEL(
        N28), .F(\Data_Mem/n9127 ) );
  MUX \Data_Mem/U9181  ( .IN0(o[1942]), .IN1(o[1974]), .SEL(N29), .F(
        \Data_Mem/n9126 ) );
  MUX \Data_Mem/U9180  ( .IN0(o[2006]), .IN1(o[2038]), .SEL(N29), .F(
        \Data_Mem/n9125 ) );
  MUX \Data_Mem/U9179  ( .IN0(\Data_Mem/n9124 ), .IN1(\Data_Mem/n9093 ), .SEL(
        N24), .F(\Data_Mem/N724 ) );
  MUX \Data_Mem/U9178  ( .IN0(\Data_Mem/n9123 ), .IN1(\Data_Mem/n9108 ), .SEL(
        N25), .F(\Data_Mem/n9124 ) );
  MUX \Data_Mem/U9177  ( .IN0(\Data_Mem/n9122 ), .IN1(\Data_Mem/n9115 ), .SEL(
        N26), .F(\Data_Mem/n9123 ) );
  MUX \Data_Mem/U9176  ( .IN0(\Data_Mem/n9121 ), .IN1(\Data_Mem/n9118 ), .SEL(
        N27), .F(\Data_Mem/n9122 ) );
  MUX \Data_Mem/U9175  ( .IN0(\Data_Mem/n9120 ), .IN1(\Data_Mem/n9119 ), .SEL(
        N28), .F(\Data_Mem/n9121 ) );
  MUX \Data_Mem/U9174  ( .IN0(o[21]), .IN1(o[53]), .SEL(N29), .F(
        \Data_Mem/n9120 ) );
  MUX \Data_Mem/U9173  ( .IN0(o[85]), .IN1(o[117]), .SEL(N29), .F(
        \Data_Mem/n9119 ) );
  MUX \Data_Mem/U9172  ( .IN0(\Data_Mem/n9117 ), .IN1(\Data_Mem/n9116 ), .SEL(
        N28), .F(\Data_Mem/n9118 ) );
  MUX \Data_Mem/U9171  ( .IN0(o[149]), .IN1(o[181]), .SEL(N29), .F(
        \Data_Mem/n9117 ) );
  MUX \Data_Mem/U9170  ( .IN0(o[213]), .IN1(o[245]), .SEL(N29), .F(
        \Data_Mem/n9116 ) );
  MUX \Data_Mem/U9169  ( .IN0(\Data_Mem/n9114 ), .IN1(\Data_Mem/n9111 ), .SEL(
        N27), .F(\Data_Mem/n9115 ) );
  MUX \Data_Mem/U9168  ( .IN0(\Data_Mem/n9113 ), .IN1(\Data_Mem/n9112 ), .SEL(
        N28), .F(\Data_Mem/n9114 ) );
  MUX \Data_Mem/U9167  ( .IN0(o[277]), .IN1(o[309]), .SEL(N29), .F(
        \Data_Mem/n9113 ) );
  MUX \Data_Mem/U9166  ( .IN0(o[341]), .IN1(o[373]), .SEL(N29), .F(
        \Data_Mem/n9112 ) );
  MUX \Data_Mem/U9165  ( .IN0(\Data_Mem/n9110 ), .IN1(\Data_Mem/n9109 ), .SEL(
        N28), .F(\Data_Mem/n9111 ) );
  MUX \Data_Mem/U9164  ( .IN0(o[405]), .IN1(o[437]), .SEL(N29), .F(
        \Data_Mem/n9110 ) );
  MUX \Data_Mem/U9163  ( .IN0(o[469]), .IN1(o[501]), .SEL(N29), .F(
        \Data_Mem/n9109 ) );
  MUX \Data_Mem/U9162  ( .IN0(\Data_Mem/n9107 ), .IN1(\Data_Mem/n9100 ), .SEL(
        N26), .F(\Data_Mem/n9108 ) );
  MUX \Data_Mem/U9161  ( .IN0(\Data_Mem/n9106 ), .IN1(\Data_Mem/n9103 ), .SEL(
        N27), .F(\Data_Mem/n9107 ) );
  MUX \Data_Mem/U9160  ( .IN0(\Data_Mem/n9105 ), .IN1(\Data_Mem/n9104 ), .SEL(
        N28), .F(\Data_Mem/n9106 ) );
  MUX \Data_Mem/U9159  ( .IN0(o[533]), .IN1(o[565]), .SEL(N29), .F(
        \Data_Mem/n9105 ) );
  MUX \Data_Mem/U9158  ( .IN0(o[597]), .IN1(o[629]), .SEL(N29), .F(
        \Data_Mem/n9104 ) );
  MUX \Data_Mem/U9157  ( .IN0(\Data_Mem/n9102 ), .IN1(\Data_Mem/n9101 ), .SEL(
        N28), .F(\Data_Mem/n9103 ) );
  MUX \Data_Mem/U9156  ( .IN0(o[661]), .IN1(o[693]), .SEL(N29), .F(
        \Data_Mem/n9102 ) );
  MUX \Data_Mem/U9155  ( .IN0(o[725]), .IN1(o[757]), .SEL(N29), .F(
        \Data_Mem/n9101 ) );
  MUX \Data_Mem/U9154  ( .IN0(\Data_Mem/n9099 ), .IN1(\Data_Mem/n9096 ), .SEL(
        N27), .F(\Data_Mem/n9100 ) );
  MUX \Data_Mem/U9153  ( .IN0(\Data_Mem/n9098 ), .IN1(\Data_Mem/n9097 ), .SEL(
        N28), .F(\Data_Mem/n9099 ) );
  MUX \Data_Mem/U9152  ( .IN0(o[789]), .IN1(o[821]), .SEL(N29), .F(
        \Data_Mem/n9098 ) );
  MUX \Data_Mem/U9151  ( .IN0(o[853]), .IN1(o[885]), .SEL(N29), .F(
        \Data_Mem/n9097 ) );
  MUX \Data_Mem/U9150  ( .IN0(\Data_Mem/n9095 ), .IN1(\Data_Mem/n9094 ), .SEL(
        N28), .F(\Data_Mem/n9096 ) );
  MUX \Data_Mem/U9149  ( .IN0(o[917]), .IN1(o[949]), .SEL(N29), .F(
        \Data_Mem/n9095 ) );
  MUX \Data_Mem/U9148  ( .IN0(o[981]), .IN1(o[1013]), .SEL(N29), .F(
        \Data_Mem/n9094 ) );
  MUX \Data_Mem/U9147  ( .IN0(\Data_Mem/n9092 ), .IN1(\Data_Mem/n9077 ), .SEL(
        N25), .F(\Data_Mem/n9093 ) );
  MUX \Data_Mem/U9146  ( .IN0(\Data_Mem/n9091 ), .IN1(\Data_Mem/n9084 ), .SEL(
        N26), .F(\Data_Mem/n9092 ) );
  MUX \Data_Mem/U9145  ( .IN0(\Data_Mem/n9090 ), .IN1(\Data_Mem/n9087 ), .SEL(
        N27), .F(\Data_Mem/n9091 ) );
  MUX \Data_Mem/U9144  ( .IN0(\Data_Mem/n9089 ), .IN1(\Data_Mem/n9088 ), .SEL(
        N28), .F(\Data_Mem/n9090 ) );
  MUX \Data_Mem/U9143  ( .IN0(o[1045]), .IN1(o[1077]), .SEL(N29), .F(
        \Data_Mem/n9089 ) );
  MUX \Data_Mem/U9142  ( .IN0(o[1109]), .IN1(o[1141]), .SEL(N29), .F(
        \Data_Mem/n9088 ) );
  MUX \Data_Mem/U9141  ( .IN0(\Data_Mem/n9086 ), .IN1(\Data_Mem/n9085 ), .SEL(
        N28), .F(\Data_Mem/n9087 ) );
  MUX \Data_Mem/U9140  ( .IN0(o[1173]), .IN1(o[1205]), .SEL(N29), .F(
        \Data_Mem/n9086 ) );
  MUX \Data_Mem/U9139  ( .IN0(o[1237]), .IN1(o[1269]), .SEL(N29), .F(
        \Data_Mem/n9085 ) );
  MUX \Data_Mem/U9138  ( .IN0(\Data_Mem/n9083 ), .IN1(\Data_Mem/n9080 ), .SEL(
        N27), .F(\Data_Mem/n9084 ) );
  MUX \Data_Mem/U9137  ( .IN0(\Data_Mem/n9082 ), .IN1(\Data_Mem/n9081 ), .SEL(
        N28), .F(\Data_Mem/n9083 ) );
  MUX \Data_Mem/U9136  ( .IN0(o[1301]), .IN1(o[1333]), .SEL(N29), .F(
        \Data_Mem/n9082 ) );
  MUX \Data_Mem/U9135  ( .IN0(o[1365]), .IN1(o[1397]), .SEL(N29), .F(
        \Data_Mem/n9081 ) );
  MUX \Data_Mem/U9134  ( .IN0(\Data_Mem/n9079 ), .IN1(\Data_Mem/n9078 ), .SEL(
        N28), .F(\Data_Mem/n9080 ) );
  MUX \Data_Mem/U9133  ( .IN0(o[1429]), .IN1(o[1461]), .SEL(N29), .F(
        \Data_Mem/n9079 ) );
  MUX \Data_Mem/U9132  ( .IN0(o[1493]), .IN1(o[1525]), .SEL(N29), .F(
        \Data_Mem/n9078 ) );
  MUX \Data_Mem/U9131  ( .IN0(\Data_Mem/n9076 ), .IN1(\Data_Mem/n9069 ), .SEL(
        N26), .F(\Data_Mem/n9077 ) );
  MUX \Data_Mem/U9130  ( .IN0(\Data_Mem/n9075 ), .IN1(\Data_Mem/n9072 ), .SEL(
        N27), .F(\Data_Mem/n9076 ) );
  MUX \Data_Mem/U9129  ( .IN0(\Data_Mem/n9074 ), .IN1(\Data_Mem/n9073 ), .SEL(
        N28), .F(\Data_Mem/n9075 ) );
  MUX \Data_Mem/U9128  ( .IN0(o[1557]), .IN1(o[1589]), .SEL(N29), .F(
        \Data_Mem/n9074 ) );
  MUX \Data_Mem/U9127  ( .IN0(o[1621]), .IN1(o[1653]), .SEL(N29), .F(
        \Data_Mem/n9073 ) );
  MUX \Data_Mem/U9126  ( .IN0(\Data_Mem/n9071 ), .IN1(\Data_Mem/n9070 ), .SEL(
        N28), .F(\Data_Mem/n9072 ) );
  MUX \Data_Mem/U9125  ( .IN0(o[1685]), .IN1(o[1717]), .SEL(N29), .F(
        \Data_Mem/n9071 ) );
  MUX \Data_Mem/U9124  ( .IN0(o[1749]), .IN1(o[1781]), .SEL(N29), .F(
        \Data_Mem/n9070 ) );
  MUX \Data_Mem/U9123  ( .IN0(\Data_Mem/n9068 ), .IN1(\Data_Mem/n9065 ), .SEL(
        N27), .F(\Data_Mem/n9069 ) );
  MUX \Data_Mem/U9122  ( .IN0(\Data_Mem/n9067 ), .IN1(\Data_Mem/n9066 ), .SEL(
        N28), .F(\Data_Mem/n9068 ) );
  MUX \Data_Mem/U9121  ( .IN0(o[1813]), .IN1(o[1845]), .SEL(N29), .F(
        \Data_Mem/n9067 ) );
  MUX \Data_Mem/U9120  ( .IN0(o[1877]), .IN1(o[1909]), .SEL(N29), .F(
        \Data_Mem/n9066 ) );
  MUX \Data_Mem/U9119  ( .IN0(\Data_Mem/n9064 ), .IN1(\Data_Mem/n9063 ), .SEL(
        N28), .F(\Data_Mem/n9065 ) );
  MUX \Data_Mem/U9118  ( .IN0(o[1941]), .IN1(o[1973]), .SEL(N29), .F(
        \Data_Mem/n9064 ) );
  MUX \Data_Mem/U9117  ( .IN0(o[2005]), .IN1(o[2037]), .SEL(N29), .F(
        \Data_Mem/n9063 ) );
  MUX \Data_Mem/U9116  ( .IN0(\Data_Mem/n9062 ), .IN1(\Data_Mem/n9031 ), .SEL(
        N24), .F(\Data_Mem/N725 ) );
  MUX \Data_Mem/U9115  ( .IN0(\Data_Mem/n9061 ), .IN1(\Data_Mem/n9046 ), .SEL(
        N25), .F(\Data_Mem/n9062 ) );
  MUX \Data_Mem/U9114  ( .IN0(\Data_Mem/n9060 ), .IN1(\Data_Mem/n9053 ), .SEL(
        N26), .F(\Data_Mem/n9061 ) );
  MUX \Data_Mem/U9113  ( .IN0(\Data_Mem/n9059 ), .IN1(\Data_Mem/n9056 ), .SEL(
        N27), .F(\Data_Mem/n9060 ) );
  MUX \Data_Mem/U9112  ( .IN0(\Data_Mem/n9058 ), .IN1(\Data_Mem/n9057 ), .SEL(
        N28), .F(\Data_Mem/n9059 ) );
  MUX \Data_Mem/U9111  ( .IN0(o[20]), .IN1(o[52]), .SEL(N29), .F(
        \Data_Mem/n9058 ) );
  MUX \Data_Mem/U9110  ( .IN0(o[84]), .IN1(o[116]), .SEL(N29), .F(
        \Data_Mem/n9057 ) );
  MUX \Data_Mem/U9109  ( .IN0(\Data_Mem/n9055 ), .IN1(\Data_Mem/n9054 ), .SEL(
        N28), .F(\Data_Mem/n9056 ) );
  MUX \Data_Mem/U9108  ( .IN0(o[148]), .IN1(o[180]), .SEL(N29), .F(
        \Data_Mem/n9055 ) );
  MUX \Data_Mem/U9107  ( .IN0(o[212]), .IN1(o[244]), .SEL(N29), .F(
        \Data_Mem/n9054 ) );
  MUX \Data_Mem/U9106  ( .IN0(\Data_Mem/n9052 ), .IN1(\Data_Mem/n9049 ), .SEL(
        N27), .F(\Data_Mem/n9053 ) );
  MUX \Data_Mem/U9105  ( .IN0(\Data_Mem/n9051 ), .IN1(\Data_Mem/n9050 ), .SEL(
        N28), .F(\Data_Mem/n9052 ) );
  MUX \Data_Mem/U9104  ( .IN0(o[276]), .IN1(o[308]), .SEL(N29), .F(
        \Data_Mem/n9051 ) );
  MUX \Data_Mem/U9103  ( .IN0(o[340]), .IN1(o[372]), .SEL(N29), .F(
        \Data_Mem/n9050 ) );
  MUX \Data_Mem/U9102  ( .IN0(\Data_Mem/n9048 ), .IN1(\Data_Mem/n9047 ), .SEL(
        N28), .F(\Data_Mem/n9049 ) );
  MUX \Data_Mem/U9101  ( .IN0(o[404]), .IN1(o[436]), .SEL(N29), .F(
        \Data_Mem/n9048 ) );
  MUX \Data_Mem/U9100  ( .IN0(o[468]), .IN1(o[500]), .SEL(N29), .F(
        \Data_Mem/n9047 ) );
  MUX \Data_Mem/U9099  ( .IN0(\Data_Mem/n9045 ), .IN1(\Data_Mem/n9038 ), .SEL(
        N26), .F(\Data_Mem/n9046 ) );
  MUX \Data_Mem/U9098  ( .IN0(\Data_Mem/n9044 ), .IN1(\Data_Mem/n9041 ), .SEL(
        N27), .F(\Data_Mem/n9045 ) );
  MUX \Data_Mem/U9097  ( .IN0(\Data_Mem/n9043 ), .IN1(\Data_Mem/n9042 ), .SEL(
        N28), .F(\Data_Mem/n9044 ) );
  MUX \Data_Mem/U9096  ( .IN0(o[532]), .IN1(o[564]), .SEL(N29), .F(
        \Data_Mem/n9043 ) );
  MUX \Data_Mem/U9095  ( .IN0(o[596]), .IN1(o[628]), .SEL(N29), .F(
        \Data_Mem/n9042 ) );
  MUX \Data_Mem/U9094  ( .IN0(\Data_Mem/n9040 ), .IN1(\Data_Mem/n9039 ), .SEL(
        N28), .F(\Data_Mem/n9041 ) );
  MUX \Data_Mem/U9093  ( .IN0(o[660]), .IN1(o[692]), .SEL(N29), .F(
        \Data_Mem/n9040 ) );
  MUX \Data_Mem/U9092  ( .IN0(o[724]), .IN1(o[756]), .SEL(N29), .F(
        \Data_Mem/n9039 ) );
  MUX \Data_Mem/U9091  ( .IN0(\Data_Mem/n9037 ), .IN1(\Data_Mem/n9034 ), .SEL(
        N27), .F(\Data_Mem/n9038 ) );
  MUX \Data_Mem/U9090  ( .IN0(\Data_Mem/n9036 ), .IN1(\Data_Mem/n9035 ), .SEL(
        N28), .F(\Data_Mem/n9037 ) );
  MUX \Data_Mem/U9089  ( .IN0(o[788]), .IN1(o[820]), .SEL(N29), .F(
        \Data_Mem/n9036 ) );
  MUX \Data_Mem/U9088  ( .IN0(o[852]), .IN1(o[884]), .SEL(N29), .F(
        \Data_Mem/n9035 ) );
  MUX \Data_Mem/U9087  ( .IN0(\Data_Mem/n9033 ), .IN1(\Data_Mem/n9032 ), .SEL(
        N28), .F(\Data_Mem/n9034 ) );
  MUX \Data_Mem/U9086  ( .IN0(o[916]), .IN1(o[948]), .SEL(N29), .F(
        \Data_Mem/n9033 ) );
  MUX \Data_Mem/U9085  ( .IN0(o[980]), .IN1(o[1012]), .SEL(N29), .F(
        \Data_Mem/n9032 ) );
  MUX \Data_Mem/U9084  ( .IN0(\Data_Mem/n9030 ), .IN1(\Data_Mem/n9015 ), .SEL(
        N25), .F(\Data_Mem/n9031 ) );
  MUX \Data_Mem/U9083  ( .IN0(\Data_Mem/n9029 ), .IN1(\Data_Mem/n9022 ), .SEL(
        N26), .F(\Data_Mem/n9030 ) );
  MUX \Data_Mem/U9082  ( .IN0(\Data_Mem/n9028 ), .IN1(\Data_Mem/n9025 ), .SEL(
        N27), .F(\Data_Mem/n9029 ) );
  MUX \Data_Mem/U9081  ( .IN0(\Data_Mem/n9027 ), .IN1(\Data_Mem/n9026 ), .SEL(
        N28), .F(\Data_Mem/n9028 ) );
  MUX \Data_Mem/U9080  ( .IN0(o[1044]), .IN1(o[1076]), .SEL(N29), .F(
        \Data_Mem/n9027 ) );
  MUX \Data_Mem/U9079  ( .IN0(o[1108]), .IN1(o[1140]), .SEL(N29), .F(
        \Data_Mem/n9026 ) );
  MUX \Data_Mem/U9078  ( .IN0(\Data_Mem/n9024 ), .IN1(\Data_Mem/n9023 ), .SEL(
        N28), .F(\Data_Mem/n9025 ) );
  MUX \Data_Mem/U9077  ( .IN0(o[1172]), .IN1(o[1204]), .SEL(N29), .F(
        \Data_Mem/n9024 ) );
  MUX \Data_Mem/U9076  ( .IN0(o[1236]), .IN1(o[1268]), .SEL(N29), .F(
        \Data_Mem/n9023 ) );
  MUX \Data_Mem/U9075  ( .IN0(\Data_Mem/n9021 ), .IN1(\Data_Mem/n9018 ), .SEL(
        N27), .F(\Data_Mem/n9022 ) );
  MUX \Data_Mem/U9074  ( .IN0(\Data_Mem/n9020 ), .IN1(\Data_Mem/n9019 ), .SEL(
        N28), .F(\Data_Mem/n9021 ) );
  MUX \Data_Mem/U9073  ( .IN0(o[1300]), .IN1(o[1332]), .SEL(N29), .F(
        \Data_Mem/n9020 ) );
  MUX \Data_Mem/U9072  ( .IN0(o[1364]), .IN1(o[1396]), .SEL(N29), .F(
        \Data_Mem/n9019 ) );
  MUX \Data_Mem/U9071  ( .IN0(\Data_Mem/n9017 ), .IN1(\Data_Mem/n9016 ), .SEL(
        N28), .F(\Data_Mem/n9018 ) );
  MUX \Data_Mem/U9070  ( .IN0(o[1428]), .IN1(o[1460]), .SEL(N29), .F(
        \Data_Mem/n9017 ) );
  MUX \Data_Mem/U9069  ( .IN0(o[1492]), .IN1(o[1524]), .SEL(N29), .F(
        \Data_Mem/n9016 ) );
  MUX \Data_Mem/U9068  ( .IN0(\Data_Mem/n9014 ), .IN1(\Data_Mem/n9007 ), .SEL(
        N26), .F(\Data_Mem/n9015 ) );
  MUX \Data_Mem/U9067  ( .IN0(\Data_Mem/n9013 ), .IN1(\Data_Mem/n9010 ), .SEL(
        N27), .F(\Data_Mem/n9014 ) );
  MUX \Data_Mem/U9066  ( .IN0(\Data_Mem/n9012 ), .IN1(\Data_Mem/n9011 ), .SEL(
        N28), .F(\Data_Mem/n9013 ) );
  MUX \Data_Mem/U9065  ( .IN0(o[1556]), .IN1(o[1588]), .SEL(N29), .F(
        \Data_Mem/n9012 ) );
  MUX \Data_Mem/U9064  ( .IN0(o[1620]), .IN1(o[1652]), .SEL(N29), .F(
        \Data_Mem/n9011 ) );
  MUX \Data_Mem/U9063  ( .IN0(\Data_Mem/n9009 ), .IN1(\Data_Mem/n9008 ), .SEL(
        N28), .F(\Data_Mem/n9010 ) );
  MUX \Data_Mem/U9062  ( .IN0(o[1684]), .IN1(o[1716]), .SEL(N29), .F(
        \Data_Mem/n9009 ) );
  MUX \Data_Mem/U9061  ( .IN0(o[1748]), .IN1(o[1780]), .SEL(N29), .F(
        \Data_Mem/n9008 ) );
  MUX \Data_Mem/U9060  ( .IN0(\Data_Mem/n9006 ), .IN1(\Data_Mem/n9003 ), .SEL(
        N27), .F(\Data_Mem/n9007 ) );
  MUX \Data_Mem/U9059  ( .IN0(\Data_Mem/n9005 ), .IN1(\Data_Mem/n9004 ), .SEL(
        N28), .F(\Data_Mem/n9006 ) );
  MUX \Data_Mem/U9058  ( .IN0(o[1812]), .IN1(o[1844]), .SEL(N29), .F(
        \Data_Mem/n9005 ) );
  MUX \Data_Mem/U9057  ( .IN0(o[1876]), .IN1(o[1908]), .SEL(N29), .F(
        \Data_Mem/n9004 ) );
  MUX \Data_Mem/U9056  ( .IN0(\Data_Mem/n9002 ), .IN1(\Data_Mem/n9001 ), .SEL(
        N28), .F(\Data_Mem/n9003 ) );
  MUX \Data_Mem/U9055  ( .IN0(o[1940]), .IN1(o[1972]), .SEL(N29), .F(
        \Data_Mem/n9002 ) );
  MUX \Data_Mem/U9054  ( .IN0(o[2004]), .IN1(o[2036]), .SEL(N29), .F(
        \Data_Mem/n9001 ) );
  MUX \Data_Mem/U9053  ( .IN0(\Data_Mem/n9000 ), .IN1(\Data_Mem/n8969 ), .SEL(
        N24), .F(\Data_Mem/N726 ) );
  MUX \Data_Mem/U9052  ( .IN0(\Data_Mem/n8999 ), .IN1(\Data_Mem/n8984 ), .SEL(
        N25), .F(\Data_Mem/n9000 ) );
  MUX \Data_Mem/U9051  ( .IN0(\Data_Mem/n8998 ), .IN1(\Data_Mem/n8991 ), .SEL(
        N26), .F(\Data_Mem/n8999 ) );
  MUX \Data_Mem/U9050  ( .IN0(\Data_Mem/n8997 ), .IN1(\Data_Mem/n8994 ), .SEL(
        N27), .F(\Data_Mem/n8998 ) );
  MUX \Data_Mem/U9049  ( .IN0(\Data_Mem/n8996 ), .IN1(\Data_Mem/n8995 ), .SEL(
        N28), .F(\Data_Mem/n8997 ) );
  MUX \Data_Mem/U9048  ( .IN0(o[19]), .IN1(o[51]), .SEL(N29), .F(
        \Data_Mem/n8996 ) );
  MUX \Data_Mem/U9047  ( .IN0(o[83]), .IN1(o[115]), .SEL(N29), .F(
        \Data_Mem/n8995 ) );
  MUX \Data_Mem/U9046  ( .IN0(\Data_Mem/n8993 ), .IN1(\Data_Mem/n8992 ), .SEL(
        N28), .F(\Data_Mem/n8994 ) );
  MUX \Data_Mem/U9045  ( .IN0(o[147]), .IN1(o[179]), .SEL(N29), .F(
        \Data_Mem/n8993 ) );
  MUX \Data_Mem/U9044  ( .IN0(o[211]), .IN1(o[243]), .SEL(N29), .F(
        \Data_Mem/n8992 ) );
  MUX \Data_Mem/U9043  ( .IN0(\Data_Mem/n8990 ), .IN1(\Data_Mem/n8987 ), .SEL(
        N27), .F(\Data_Mem/n8991 ) );
  MUX \Data_Mem/U9042  ( .IN0(\Data_Mem/n8989 ), .IN1(\Data_Mem/n8988 ), .SEL(
        N28), .F(\Data_Mem/n8990 ) );
  MUX \Data_Mem/U9041  ( .IN0(o[275]), .IN1(o[307]), .SEL(N29), .F(
        \Data_Mem/n8989 ) );
  MUX \Data_Mem/U9040  ( .IN0(o[339]), .IN1(o[371]), .SEL(N29), .F(
        \Data_Mem/n8988 ) );
  MUX \Data_Mem/U9039  ( .IN0(\Data_Mem/n8986 ), .IN1(\Data_Mem/n8985 ), .SEL(
        N28), .F(\Data_Mem/n8987 ) );
  MUX \Data_Mem/U9038  ( .IN0(o[403]), .IN1(o[435]), .SEL(N29), .F(
        \Data_Mem/n8986 ) );
  MUX \Data_Mem/U9037  ( .IN0(o[467]), .IN1(o[499]), .SEL(N29), .F(
        \Data_Mem/n8985 ) );
  MUX \Data_Mem/U9036  ( .IN0(\Data_Mem/n8983 ), .IN1(\Data_Mem/n8976 ), .SEL(
        N26), .F(\Data_Mem/n8984 ) );
  MUX \Data_Mem/U9035  ( .IN0(\Data_Mem/n8982 ), .IN1(\Data_Mem/n8979 ), .SEL(
        N27), .F(\Data_Mem/n8983 ) );
  MUX \Data_Mem/U9034  ( .IN0(\Data_Mem/n8981 ), .IN1(\Data_Mem/n8980 ), .SEL(
        N28), .F(\Data_Mem/n8982 ) );
  MUX \Data_Mem/U9033  ( .IN0(o[531]), .IN1(o[563]), .SEL(N29), .F(
        \Data_Mem/n8981 ) );
  MUX \Data_Mem/U9032  ( .IN0(o[595]), .IN1(o[627]), .SEL(N29), .F(
        \Data_Mem/n8980 ) );
  MUX \Data_Mem/U9031  ( .IN0(\Data_Mem/n8978 ), .IN1(\Data_Mem/n8977 ), .SEL(
        N28), .F(\Data_Mem/n8979 ) );
  MUX \Data_Mem/U9030  ( .IN0(o[659]), .IN1(o[691]), .SEL(N29), .F(
        \Data_Mem/n8978 ) );
  MUX \Data_Mem/U9029  ( .IN0(o[723]), .IN1(o[755]), .SEL(N29), .F(
        \Data_Mem/n8977 ) );
  MUX \Data_Mem/U9028  ( .IN0(\Data_Mem/n8975 ), .IN1(\Data_Mem/n8972 ), .SEL(
        N27), .F(\Data_Mem/n8976 ) );
  MUX \Data_Mem/U9027  ( .IN0(\Data_Mem/n8974 ), .IN1(\Data_Mem/n8973 ), .SEL(
        N28), .F(\Data_Mem/n8975 ) );
  MUX \Data_Mem/U9026  ( .IN0(o[787]), .IN1(o[819]), .SEL(N29), .F(
        \Data_Mem/n8974 ) );
  MUX \Data_Mem/U9025  ( .IN0(o[851]), .IN1(o[883]), .SEL(N29), .F(
        \Data_Mem/n8973 ) );
  MUX \Data_Mem/U9024  ( .IN0(\Data_Mem/n8971 ), .IN1(\Data_Mem/n8970 ), .SEL(
        N28), .F(\Data_Mem/n8972 ) );
  MUX \Data_Mem/U9023  ( .IN0(o[915]), .IN1(o[947]), .SEL(N29), .F(
        \Data_Mem/n8971 ) );
  MUX \Data_Mem/U9022  ( .IN0(o[979]), .IN1(o[1011]), .SEL(N29), .F(
        \Data_Mem/n8970 ) );
  MUX \Data_Mem/U9021  ( .IN0(\Data_Mem/n8968 ), .IN1(\Data_Mem/n8953 ), .SEL(
        N25), .F(\Data_Mem/n8969 ) );
  MUX \Data_Mem/U9020  ( .IN0(\Data_Mem/n8967 ), .IN1(\Data_Mem/n8960 ), .SEL(
        N26), .F(\Data_Mem/n8968 ) );
  MUX \Data_Mem/U9019  ( .IN0(\Data_Mem/n8966 ), .IN1(\Data_Mem/n8963 ), .SEL(
        N27), .F(\Data_Mem/n8967 ) );
  MUX \Data_Mem/U9018  ( .IN0(\Data_Mem/n8965 ), .IN1(\Data_Mem/n8964 ), .SEL(
        N28), .F(\Data_Mem/n8966 ) );
  MUX \Data_Mem/U9017  ( .IN0(o[1043]), .IN1(o[1075]), .SEL(N29), .F(
        \Data_Mem/n8965 ) );
  MUX \Data_Mem/U9016  ( .IN0(o[1107]), .IN1(o[1139]), .SEL(N29), .F(
        \Data_Mem/n8964 ) );
  MUX \Data_Mem/U9015  ( .IN0(\Data_Mem/n8962 ), .IN1(\Data_Mem/n8961 ), .SEL(
        N28), .F(\Data_Mem/n8963 ) );
  MUX \Data_Mem/U9014  ( .IN0(o[1171]), .IN1(o[1203]), .SEL(N29), .F(
        \Data_Mem/n8962 ) );
  MUX \Data_Mem/U9013  ( .IN0(o[1235]), .IN1(o[1267]), .SEL(N29), .F(
        \Data_Mem/n8961 ) );
  MUX \Data_Mem/U9012  ( .IN0(\Data_Mem/n8959 ), .IN1(\Data_Mem/n8956 ), .SEL(
        N27), .F(\Data_Mem/n8960 ) );
  MUX \Data_Mem/U9011  ( .IN0(\Data_Mem/n8958 ), .IN1(\Data_Mem/n8957 ), .SEL(
        N28), .F(\Data_Mem/n8959 ) );
  MUX \Data_Mem/U9010  ( .IN0(o[1299]), .IN1(o[1331]), .SEL(N29), .F(
        \Data_Mem/n8958 ) );
  MUX \Data_Mem/U9009  ( .IN0(o[1363]), .IN1(o[1395]), .SEL(N29), .F(
        \Data_Mem/n8957 ) );
  MUX \Data_Mem/U9008  ( .IN0(\Data_Mem/n8955 ), .IN1(\Data_Mem/n8954 ), .SEL(
        N28), .F(\Data_Mem/n8956 ) );
  MUX \Data_Mem/U9007  ( .IN0(o[1427]), .IN1(o[1459]), .SEL(N29), .F(
        \Data_Mem/n8955 ) );
  MUX \Data_Mem/U9006  ( .IN0(o[1491]), .IN1(o[1523]), .SEL(N29), .F(
        \Data_Mem/n8954 ) );
  MUX \Data_Mem/U9005  ( .IN0(\Data_Mem/n8952 ), .IN1(\Data_Mem/n8945 ), .SEL(
        N26), .F(\Data_Mem/n8953 ) );
  MUX \Data_Mem/U9004  ( .IN0(\Data_Mem/n8951 ), .IN1(\Data_Mem/n8948 ), .SEL(
        N27), .F(\Data_Mem/n8952 ) );
  MUX \Data_Mem/U9003  ( .IN0(\Data_Mem/n8950 ), .IN1(\Data_Mem/n8949 ), .SEL(
        N28), .F(\Data_Mem/n8951 ) );
  MUX \Data_Mem/U9002  ( .IN0(o[1555]), .IN1(o[1587]), .SEL(N29), .F(
        \Data_Mem/n8950 ) );
  MUX \Data_Mem/U9001  ( .IN0(o[1619]), .IN1(o[1651]), .SEL(N29), .F(
        \Data_Mem/n8949 ) );
  MUX \Data_Mem/U9000  ( .IN0(\Data_Mem/n8947 ), .IN1(\Data_Mem/n8946 ), .SEL(
        N28), .F(\Data_Mem/n8948 ) );
  MUX \Data_Mem/U8999  ( .IN0(o[1683]), .IN1(o[1715]), .SEL(N29), .F(
        \Data_Mem/n8947 ) );
  MUX \Data_Mem/U8998  ( .IN0(o[1747]), .IN1(o[1779]), .SEL(N29), .F(
        \Data_Mem/n8946 ) );
  MUX \Data_Mem/U8997  ( .IN0(\Data_Mem/n8944 ), .IN1(\Data_Mem/n8941 ), .SEL(
        N27), .F(\Data_Mem/n8945 ) );
  MUX \Data_Mem/U8996  ( .IN0(\Data_Mem/n8943 ), .IN1(\Data_Mem/n8942 ), .SEL(
        N28), .F(\Data_Mem/n8944 ) );
  MUX \Data_Mem/U8995  ( .IN0(o[1811]), .IN1(o[1843]), .SEL(N29), .F(
        \Data_Mem/n8943 ) );
  MUX \Data_Mem/U8994  ( .IN0(o[1875]), .IN1(o[1907]), .SEL(N29), .F(
        \Data_Mem/n8942 ) );
  MUX \Data_Mem/U8993  ( .IN0(\Data_Mem/n8940 ), .IN1(\Data_Mem/n8939 ), .SEL(
        N28), .F(\Data_Mem/n8941 ) );
  MUX \Data_Mem/U8992  ( .IN0(o[1939]), .IN1(o[1971]), .SEL(N29), .F(
        \Data_Mem/n8940 ) );
  MUX \Data_Mem/U8991  ( .IN0(o[2003]), .IN1(o[2035]), .SEL(N29), .F(
        \Data_Mem/n8939 ) );
  MUX \Data_Mem/U8990  ( .IN0(\Data_Mem/n8938 ), .IN1(\Data_Mem/n8907 ), .SEL(
        N24), .F(\Data_Mem/N727 ) );
  MUX \Data_Mem/U8989  ( .IN0(\Data_Mem/n8937 ), .IN1(\Data_Mem/n8922 ), .SEL(
        N25), .F(\Data_Mem/n8938 ) );
  MUX \Data_Mem/U8988  ( .IN0(\Data_Mem/n8936 ), .IN1(\Data_Mem/n8929 ), .SEL(
        N26), .F(\Data_Mem/n8937 ) );
  MUX \Data_Mem/U8987  ( .IN0(\Data_Mem/n8935 ), .IN1(\Data_Mem/n8932 ), .SEL(
        N27), .F(\Data_Mem/n8936 ) );
  MUX \Data_Mem/U8986  ( .IN0(\Data_Mem/n8934 ), .IN1(\Data_Mem/n8933 ), .SEL(
        N28), .F(\Data_Mem/n8935 ) );
  MUX \Data_Mem/U8985  ( .IN0(o[18]), .IN1(o[50]), .SEL(N29), .F(
        \Data_Mem/n8934 ) );
  MUX \Data_Mem/U8984  ( .IN0(o[82]), .IN1(o[114]), .SEL(N29), .F(
        \Data_Mem/n8933 ) );
  MUX \Data_Mem/U8983  ( .IN0(\Data_Mem/n8931 ), .IN1(\Data_Mem/n8930 ), .SEL(
        N28), .F(\Data_Mem/n8932 ) );
  MUX \Data_Mem/U8982  ( .IN0(o[146]), .IN1(o[178]), .SEL(N29), .F(
        \Data_Mem/n8931 ) );
  MUX \Data_Mem/U8981  ( .IN0(o[210]), .IN1(o[242]), .SEL(N29), .F(
        \Data_Mem/n8930 ) );
  MUX \Data_Mem/U8980  ( .IN0(\Data_Mem/n8928 ), .IN1(\Data_Mem/n8925 ), .SEL(
        N27), .F(\Data_Mem/n8929 ) );
  MUX \Data_Mem/U8979  ( .IN0(\Data_Mem/n8927 ), .IN1(\Data_Mem/n8926 ), .SEL(
        N28), .F(\Data_Mem/n8928 ) );
  MUX \Data_Mem/U8978  ( .IN0(o[274]), .IN1(o[306]), .SEL(N29), .F(
        \Data_Mem/n8927 ) );
  MUX \Data_Mem/U8977  ( .IN0(o[338]), .IN1(o[370]), .SEL(N29), .F(
        \Data_Mem/n8926 ) );
  MUX \Data_Mem/U8976  ( .IN0(\Data_Mem/n8924 ), .IN1(\Data_Mem/n8923 ), .SEL(
        N28), .F(\Data_Mem/n8925 ) );
  MUX \Data_Mem/U8975  ( .IN0(o[402]), .IN1(o[434]), .SEL(N29), .F(
        \Data_Mem/n8924 ) );
  MUX \Data_Mem/U8974  ( .IN0(o[466]), .IN1(o[498]), .SEL(N29), .F(
        \Data_Mem/n8923 ) );
  MUX \Data_Mem/U8973  ( .IN0(\Data_Mem/n8921 ), .IN1(\Data_Mem/n8914 ), .SEL(
        N26), .F(\Data_Mem/n8922 ) );
  MUX \Data_Mem/U8972  ( .IN0(\Data_Mem/n8920 ), .IN1(\Data_Mem/n8917 ), .SEL(
        N27), .F(\Data_Mem/n8921 ) );
  MUX \Data_Mem/U8971  ( .IN0(\Data_Mem/n8919 ), .IN1(\Data_Mem/n8918 ), .SEL(
        N28), .F(\Data_Mem/n8920 ) );
  MUX \Data_Mem/U8970  ( .IN0(o[530]), .IN1(o[562]), .SEL(N29), .F(
        \Data_Mem/n8919 ) );
  MUX \Data_Mem/U8969  ( .IN0(o[594]), .IN1(o[626]), .SEL(N29), .F(
        \Data_Mem/n8918 ) );
  MUX \Data_Mem/U8968  ( .IN0(\Data_Mem/n8916 ), .IN1(\Data_Mem/n8915 ), .SEL(
        N28), .F(\Data_Mem/n8917 ) );
  MUX \Data_Mem/U8967  ( .IN0(o[658]), .IN1(o[690]), .SEL(N29), .F(
        \Data_Mem/n8916 ) );
  MUX \Data_Mem/U8966  ( .IN0(o[722]), .IN1(o[754]), .SEL(N29), .F(
        \Data_Mem/n8915 ) );
  MUX \Data_Mem/U8965  ( .IN0(\Data_Mem/n8913 ), .IN1(\Data_Mem/n8910 ), .SEL(
        N27), .F(\Data_Mem/n8914 ) );
  MUX \Data_Mem/U8964  ( .IN0(\Data_Mem/n8912 ), .IN1(\Data_Mem/n8911 ), .SEL(
        N28), .F(\Data_Mem/n8913 ) );
  MUX \Data_Mem/U8963  ( .IN0(o[786]), .IN1(o[818]), .SEL(N29), .F(
        \Data_Mem/n8912 ) );
  MUX \Data_Mem/U8962  ( .IN0(o[850]), .IN1(o[882]), .SEL(N29), .F(
        \Data_Mem/n8911 ) );
  MUX \Data_Mem/U8961  ( .IN0(\Data_Mem/n8909 ), .IN1(\Data_Mem/n8908 ), .SEL(
        N28), .F(\Data_Mem/n8910 ) );
  MUX \Data_Mem/U8960  ( .IN0(o[914]), .IN1(o[946]), .SEL(N29), .F(
        \Data_Mem/n8909 ) );
  MUX \Data_Mem/U8959  ( .IN0(o[978]), .IN1(o[1010]), .SEL(N29), .F(
        \Data_Mem/n8908 ) );
  MUX \Data_Mem/U8958  ( .IN0(\Data_Mem/n8906 ), .IN1(\Data_Mem/n8891 ), .SEL(
        N25), .F(\Data_Mem/n8907 ) );
  MUX \Data_Mem/U8957  ( .IN0(\Data_Mem/n8905 ), .IN1(\Data_Mem/n8898 ), .SEL(
        N26), .F(\Data_Mem/n8906 ) );
  MUX \Data_Mem/U8956  ( .IN0(\Data_Mem/n8904 ), .IN1(\Data_Mem/n8901 ), .SEL(
        N27), .F(\Data_Mem/n8905 ) );
  MUX \Data_Mem/U8955  ( .IN0(\Data_Mem/n8903 ), .IN1(\Data_Mem/n8902 ), .SEL(
        N28), .F(\Data_Mem/n8904 ) );
  MUX \Data_Mem/U8954  ( .IN0(o[1042]), .IN1(o[1074]), .SEL(N29), .F(
        \Data_Mem/n8903 ) );
  MUX \Data_Mem/U8953  ( .IN0(o[1106]), .IN1(o[1138]), .SEL(N29), .F(
        \Data_Mem/n8902 ) );
  MUX \Data_Mem/U8952  ( .IN0(\Data_Mem/n8900 ), .IN1(\Data_Mem/n8899 ), .SEL(
        N28), .F(\Data_Mem/n8901 ) );
  MUX \Data_Mem/U8951  ( .IN0(o[1170]), .IN1(o[1202]), .SEL(N29), .F(
        \Data_Mem/n8900 ) );
  MUX \Data_Mem/U8950  ( .IN0(o[1234]), .IN1(o[1266]), .SEL(N29), .F(
        \Data_Mem/n8899 ) );
  MUX \Data_Mem/U8949  ( .IN0(\Data_Mem/n8897 ), .IN1(\Data_Mem/n8894 ), .SEL(
        N27), .F(\Data_Mem/n8898 ) );
  MUX \Data_Mem/U8948  ( .IN0(\Data_Mem/n8896 ), .IN1(\Data_Mem/n8895 ), .SEL(
        N28), .F(\Data_Mem/n8897 ) );
  MUX \Data_Mem/U8947  ( .IN0(o[1298]), .IN1(o[1330]), .SEL(N29), .F(
        \Data_Mem/n8896 ) );
  MUX \Data_Mem/U8946  ( .IN0(o[1362]), .IN1(o[1394]), .SEL(N29), .F(
        \Data_Mem/n8895 ) );
  MUX \Data_Mem/U8945  ( .IN0(\Data_Mem/n8893 ), .IN1(\Data_Mem/n8892 ), .SEL(
        N28), .F(\Data_Mem/n8894 ) );
  MUX \Data_Mem/U8944  ( .IN0(o[1426]), .IN1(o[1458]), .SEL(N29), .F(
        \Data_Mem/n8893 ) );
  MUX \Data_Mem/U8943  ( .IN0(o[1490]), .IN1(o[1522]), .SEL(N29), .F(
        \Data_Mem/n8892 ) );
  MUX \Data_Mem/U8942  ( .IN0(\Data_Mem/n8890 ), .IN1(\Data_Mem/n8883 ), .SEL(
        N26), .F(\Data_Mem/n8891 ) );
  MUX \Data_Mem/U8941  ( .IN0(\Data_Mem/n8889 ), .IN1(\Data_Mem/n8886 ), .SEL(
        N27), .F(\Data_Mem/n8890 ) );
  MUX \Data_Mem/U8940  ( .IN0(\Data_Mem/n8888 ), .IN1(\Data_Mem/n8887 ), .SEL(
        N28), .F(\Data_Mem/n8889 ) );
  MUX \Data_Mem/U8939  ( .IN0(o[1554]), .IN1(o[1586]), .SEL(N29), .F(
        \Data_Mem/n8888 ) );
  MUX \Data_Mem/U8938  ( .IN0(o[1618]), .IN1(o[1650]), .SEL(N29), .F(
        \Data_Mem/n8887 ) );
  MUX \Data_Mem/U8937  ( .IN0(\Data_Mem/n8885 ), .IN1(\Data_Mem/n8884 ), .SEL(
        N28), .F(\Data_Mem/n8886 ) );
  MUX \Data_Mem/U8936  ( .IN0(o[1682]), .IN1(o[1714]), .SEL(N29), .F(
        \Data_Mem/n8885 ) );
  MUX \Data_Mem/U8935  ( .IN0(o[1746]), .IN1(o[1778]), .SEL(N29), .F(
        \Data_Mem/n8884 ) );
  MUX \Data_Mem/U8934  ( .IN0(\Data_Mem/n8882 ), .IN1(\Data_Mem/n8879 ), .SEL(
        N27), .F(\Data_Mem/n8883 ) );
  MUX \Data_Mem/U8933  ( .IN0(\Data_Mem/n8881 ), .IN1(\Data_Mem/n8880 ), .SEL(
        N28), .F(\Data_Mem/n8882 ) );
  MUX \Data_Mem/U8932  ( .IN0(o[1810]), .IN1(o[1842]), .SEL(N29), .F(
        \Data_Mem/n8881 ) );
  MUX \Data_Mem/U8931  ( .IN0(o[1874]), .IN1(o[1906]), .SEL(N29), .F(
        \Data_Mem/n8880 ) );
  MUX \Data_Mem/U8930  ( .IN0(\Data_Mem/n8878 ), .IN1(\Data_Mem/n8877 ), .SEL(
        N28), .F(\Data_Mem/n8879 ) );
  MUX \Data_Mem/U8929  ( .IN0(o[1938]), .IN1(o[1970]), .SEL(N29), .F(
        \Data_Mem/n8878 ) );
  MUX \Data_Mem/U8928  ( .IN0(o[2002]), .IN1(o[2034]), .SEL(N29), .F(
        \Data_Mem/n8877 ) );
  MUX \Data_Mem/U8927  ( .IN0(\Data_Mem/n8876 ), .IN1(\Data_Mem/n8845 ), .SEL(
        N24), .F(\Data_Mem/N728 ) );
  MUX \Data_Mem/U8926  ( .IN0(\Data_Mem/n8875 ), .IN1(\Data_Mem/n8860 ), .SEL(
        N25), .F(\Data_Mem/n8876 ) );
  MUX \Data_Mem/U8925  ( .IN0(\Data_Mem/n8874 ), .IN1(\Data_Mem/n8867 ), .SEL(
        N26), .F(\Data_Mem/n8875 ) );
  MUX \Data_Mem/U8924  ( .IN0(\Data_Mem/n8873 ), .IN1(\Data_Mem/n8870 ), .SEL(
        N27), .F(\Data_Mem/n8874 ) );
  MUX \Data_Mem/U8923  ( .IN0(\Data_Mem/n8872 ), .IN1(\Data_Mem/n8871 ), .SEL(
        N28), .F(\Data_Mem/n8873 ) );
  MUX \Data_Mem/U8922  ( .IN0(o[17]), .IN1(o[49]), .SEL(N29), .F(
        \Data_Mem/n8872 ) );
  MUX \Data_Mem/U8921  ( .IN0(o[81]), .IN1(o[113]), .SEL(N29), .F(
        \Data_Mem/n8871 ) );
  MUX \Data_Mem/U8920  ( .IN0(\Data_Mem/n8869 ), .IN1(\Data_Mem/n8868 ), .SEL(
        N28), .F(\Data_Mem/n8870 ) );
  MUX \Data_Mem/U8919  ( .IN0(o[145]), .IN1(o[177]), .SEL(N29), .F(
        \Data_Mem/n8869 ) );
  MUX \Data_Mem/U8918  ( .IN0(o[209]), .IN1(o[241]), .SEL(N29), .F(
        \Data_Mem/n8868 ) );
  MUX \Data_Mem/U8917  ( .IN0(\Data_Mem/n8866 ), .IN1(\Data_Mem/n8863 ), .SEL(
        N27), .F(\Data_Mem/n8867 ) );
  MUX \Data_Mem/U8916  ( .IN0(\Data_Mem/n8865 ), .IN1(\Data_Mem/n8864 ), .SEL(
        N28), .F(\Data_Mem/n8866 ) );
  MUX \Data_Mem/U8915  ( .IN0(o[273]), .IN1(o[305]), .SEL(N29), .F(
        \Data_Mem/n8865 ) );
  MUX \Data_Mem/U8914  ( .IN0(o[337]), .IN1(o[369]), .SEL(N29), .F(
        \Data_Mem/n8864 ) );
  MUX \Data_Mem/U8913  ( .IN0(\Data_Mem/n8862 ), .IN1(\Data_Mem/n8861 ), .SEL(
        N28), .F(\Data_Mem/n8863 ) );
  MUX \Data_Mem/U8912  ( .IN0(o[401]), .IN1(o[433]), .SEL(N29), .F(
        \Data_Mem/n8862 ) );
  MUX \Data_Mem/U8911  ( .IN0(o[465]), .IN1(o[497]), .SEL(N29), .F(
        \Data_Mem/n8861 ) );
  MUX \Data_Mem/U8910  ( .IN0(\Data_Mem/n8859 ), .IN1(\Data_Mem/n8852 ), .SEL(
        N26), .F(\Data_Mem/n8860 ) );
  MUX \Data_Mem/U8909  ( .IN0(\Data_Mem/n8858 ), .IN1(\Data_Mem/n8855 ), .SEL(
        N27), .F(\Data_Mem/n8859 ) );
  MUX \Data_Mem/U8908  ( .IN0(\Data_Mem/n8857 ), .IN1(\Data_Mem/n8856 ), .SEL(
        N28), .F(\Data_Mem/n8858 ) );
  MUX \Data_Mem/U8907  ( .IN0(o[529]), .IN1(o[561]), .SEL(N29), .F(
        \Data_Mem/n8857 ) );
  MUX \Data_Mem/U8906  ( .IN0(o[593]), .IN1(o[625]), .SEL(N29), .F(
        \Data_Mem/n8856 ) );
  MUX \Data_Mem/U8905  ( .IN0(\Data_Mem/n8854 ), .IN1(\Data_Mem/n8853 ), .SEL(
        N28), .F(\Data_Mem/n8855 ) );
  MUX \Data_Mem/U8904  ( .IN0(o[657]), .IN1(o[689]), .SEL(N29), .F(
        \Data_Mem/n8854 ) );
  MUX \Data_Mem/U8903  ( .IN0(o[721]), .IN1(o[753]), .SEL(N29), .F(
        \Data_Mem/n8853 ) );
  MUX \Data_Mem/U8902  ( .IN0(\Data_Mem/n8851 ), .IN1(\Data_Mem/n8848 ), .SEL(
        N27), .F(\Data_Mem/n8852 ) );
  MUX \Data_Mem/U8901  ( .IN0(\Data_Mem/n8850 ), .IN1(\Data_Mem/n8849 ), .SEL(
        N28), .F(\Data_Mem/n8851 ) );
  MUX \Data_Mem/U8900  ( .IN0(o[785]), .IN1(o[817]), .SEL(N29), .F(
        \Data_Mem/n8850 ) );
  MUX \Data_Mem/U8899  ( .IN0(o[849]), .IN1(o[881]), .SEL(N29), .F(
        \Data_Mem/n8849 ) );
  MUX \Data_Mem/U8898  ( .IN0(\Data_Mem/n8847 ), .IN1(\Data_Mem/n8846 ), .SEL(
        N28), .F(\Data_Mem/n8848 ) );
  MUX \Data_Mem/U8897  ( .IN0(o[913]), .IN1(o[945]), .SEL(N29), .F(
        \Data_Mem/n8847 ) );
  MUX \Data_Mem/U8896  ( .IN0(o[977]), .IN1(o[1009]), .SEL(N29), .F(
        \Data_Mem/n8846 ) );
  MUX \Data_Mem/U8895  ( .IN0(\Data_Mem/n8844 ), .IN1(\Data_Mem/n8829 ), .SEL(
        N25), .F(\Data_Mem/n8845 ) );
  MUX \Data_Mem/U8894  ( .IN0(\Data_Mem/n8843 ), .IN1(\Data_Mem/n8836 ), .SEL(
        N26), .F(\Data_Mem/n8844 ) );
  MUX \Data_Mem/U8893  ( .IN0(\Data_Mem/n8842 ), .IN1(\Data_Mem/n8839 ), .SEL(
        N27), .F(\Data_Mem/n8843 ) );
  MUX \Data_Mem/U8892  ( .IN0(\Data_Mem/n8841 ), .IN1(\Data_Mem/n8840 ), .SEL(
        N28), .F(\Data_Mem/n8842 ) );
  MUX \Data_Mem/U8891  ( .IN0(o[1041]), .IN1(o[1073]), .SEL(N29), .F(
        \Data_Mem/n8841 ) );
  MUX \Data_Mem/U8890  ( .IN0(o[1105]), .IN1(o[1137]), .SEL(N29), .F(
        \Data_Mem/n8840 ) );
  MUX \Data_Mem/U8889  ( .IN0(\Data_Mem/n8838 ), .IN1(\Data_Mem/n8837 ), .SEL(
        N28), .F(\Data_Mem/n8839 ) );
  MUX \Data_Mem/U8888  ( .IN0(o[1169]), .IN1(o[1201]), .SEL(N29), .F(
        \Data_Mem/n8838 ) );
  MUX \Data_Mem/U8887  ( .IN0(o[1233]), .IN1(o[1265]), .SEL(N29), .F(
        \Data_Mem/n8837 ) );
  MUX \Data_Mem/U8886  ( .IN0(\Data_Mem/n8835 ), .IN1(\Data_Mem/n8832 ), .SEL(
        N27), .F(\Data_Mem/n8836 ) );
  MUX \Data_Mem/U8885  ( .IN0(\Data_Mem/n8834 ), .IN1(\Data_Mem/n8833 ), .SEL(
        N28), .F(\Data_Mem/n8835 ) );
  MUX \Data_Mem/U8884  ( .IN0(o[1297]), .IN1(o[1329]), .SEL(N29), .F(
        \Data_Mem/n8834 ) );
  MUX \Data_Mem/U8883  ( .IN0(o[1361]), .IN1(o[1393]), .SEL(N29), .F(
        \Data_Mem/n8833 ) );
  MUX \Data_Mem/U8882  ( .IN0(\Data_Mem/n8831 ), .IN1(\Data_Mem/n8830 ), .SEL(
        N28), .F(\Data_Mem/n8832 ) );
  MUX \Data_Mem/U8881  ( .IN0(o[1425]), .IN1(o[1457]), .SEL(N29), .F(
        \Data_Mem/n8831 ) );
  MUX \Data_Mem/U8880  ( .IN0(o[1489]), .IN1(o[1521]), .SEL(N29), .F(
        \Data_Mem/n8830 ) );
  MUX \Data_Mem/U8879  ( .IN0(\Data_Mem/n8828 ), .IN1(\Data_Mem/n8821 ), .SEL(
        N26), .F(\Data_Mem/n8829 ) );
  MUX \Data_Mem/U8878  ( .IN0(\Data_Mem/n8827 ), .IN1(\Data_Mem/n8824 ), .SEL(
        N27), .F(\Data_Mem/n8828 ) );
  MUX \Data_Mem/U8877  ( .IN0(\Data_Mem/n8826 ), .IN1(\Data_Mem/n8825 ), .SEL(
        N28), .F(\Data_Mem/n8827 ) );
  MUX \Data_Mem/U8876  ( .IN0(o[1553]), .IN1(o[1585]), .SEL(N29), .F(
        \Data_Mem/n8826 ) );
  MUX \Data_Mem/U8875  ( .IN0(o[1617]), .IN1(o[1649]), .SEL(N29), .F(
        \Data_Mem/n8825 ) );
  MUX \Data_Mem/U8874  ( .IN0(\Data_Mem/n8823 ), .IN1(\Data_Mem/n8822 ), .SEL(
        N28), .F(\Data_Mem/n8824 ) );
  MUX \Data_Mem/U8873  ( .IN0(o[1681]), .IN1(o[1713]), .SEL(N29), .F(
        \Data_Mem/n8823 ) );
  MUX \Data_Mem/U8872  ( .IN0(o[1745]), .IN1(o[1777]), .SEL(N29), .F(
        \Data_Mem/n8822 ) );
  MUX \Data_Mem/U8871  ( .IN0(\Data_Mem/n8820 ), .IN1(\Data_Mem/n8817 ), .SEL(
        N27), .F(\Data_Mem/n8821 ) );
  MUX \Data_Mem/U8870  ( .IN0(\Data_Mem/n8819 ), .IN1(\Data_Mem/n8818 ), .SEL(
        N28), .F(\Data_Mem/n8820 ) );
  MUX \Data_Mem/U8869  ( .IN0(o[1809]), .IN1(o[1841]), .SEL(N29), .F(
        \Data_Mem/n8819 ) );
  MUX \Data_Mem/U8868  ( .IN0(o[1873]), .IN1(o[1905]), .SEL(N29), .F(
        \Data_Mem/n8818 ) );
  MUX \Data_Mem/U8867  ( .IN0(\Data_Mem/n8816 ), .IN1(\Data_Mem/n8815 ), .SEL(
        N28), .F(\Data_Mem/n8817 ) );
  MUX \Data_Mem/U8866  ( .IN0(o[1937]), .IN1(o[1969]), .SEL(N29), .F(
        \Data_Mem/n8816 ) );
  MUX \Data_Mem/U8865  ( .IN0(o[2001]), .IN1(o[2033]), .SEL(N29), .F(
        \Data_Mem/n8815 ) );
  MUX \Data_Mem/U8864  ( .IN0(\Data_Mem/n8814 ), .IN1(\Data_Mem/n8783 ), .SEL(
        N24), .F(\Data_Mem/N729 ) );
  MUX \Data_Mem/U8863  ( .IN0(\Data_Mem/n8813 ), .IN1(\Data_Mem/n8798 ), .SEL(
        N25), .F(\Data_Mem/n8814 ) );
  MUX \Data_Mem/U8862  ( .IN0(\Data_Mem/n8812 ), .IN1(\Data_Mem/n8805 ), .SEL(
        N26), .F(\Data_Mem/n8813 ) );
  MUX \Data_Mem/U8861  ( .IN0(\Data_Mem/n8811 ), .IN1(\Data_Mem/n8808 ), .SEL(
        N27), .F(\Data_Mem/n8812 ) );
  MUX \Data_Mem/U8860  ( .IN0(\Data_Mem/n8810 ), .IN1(\Data_Mem/n8809 ), .SEL(
        N28), .F(\Data_Mem/n8811 ) );
  MUX \Data_Mem/U8859  ( .IN0(o[16]), .IN1(o[48]), .SEL(N29), .F(
        \Data_Mem/n8810 ) );
  MUX \Data_Mem/U8858  ( .IN0(o[80]), .IN1(o[112]), .SEL(N29), .F(
        \Data_Mem/n8809 ) );
  MUX \Data_Mem/U8857  ( .IN0(\Data_Mem/n8807 ), .IN1(\Data_Mem/n8806 ), .SEL(
        N28), .F(\Data_Mem/n8808 ) );
  MUX \Data_Mem/U8856  ( .IN0(o[144]), .IN1(o[176]), .SEL(N29), .F(
        \Data_Mem/n8807 ) );
  MUX \Data_Mem/U8855  ( .IN0(o[208]), .IN1(o[240]), .SEL(N29), .F(
        \Data_Mem/n8806 ) );
  MUX \Data_Mem/U8854  ( .IN0(\Data_Mem/n8804 ), .IN1(\Data_Mem/n8801 ), .SEL(
        N27), .F(\Data_Mem/n8805 ) );
  MUX \Data_Mem/U8853  ( .IN0(\Data_Mem/n8803 ), .IN1(\Data_Mem/n8802 ), .SEL(
        N28), .F(\Data_Mem/n8804 ) );
  MUX \Data_Mem/U8852  ( .IN0(o[272]), .IN1(o[304]), .SEL(N29), .F(
        \Data_Mem/n8803 ) );
  MUX \Data_Mem/U8851  ( .IN0(o[336]), .IN1(o[368]), .SEL(N29), .F(
        \Data_Mem/n8802 ) );
  MUX \Data_Mem/U8850  ( .IN0(\Data_Mem/n8800 ), .IN1(\Data_Mem/n8799 ), .SEL(
        N28), .F(\Data_Mem/n8801 ) );
  MUX \Data_Mem/U8849  ( .IN0(o[400]), .IN1(o[432]), .SEL(N29), .F(
        \Data_Mem/n8800 ) );
  MUX \Data_Mem/U8848  ( .IN0(o[464]), .IN1(o[496]), .SEL(N29), .F(
        \Data_Mem/n8799 ) );
  MUX \Data_Mem/U8847  ( .IN0(\Data_Mem/n8797 ), .IN1(\Data_Mem/n8790 ), .SEL(
        N26), .F(\Data_Mem/n8798 ) );
  MUX \Data_Mem/U8846  ( .IN0(\Data_Mem/n8796 ), .IN1(\Data_Mem/n8793 ), .SEL(
        N27), .F(\Data_Mem/n8797 ) );
  MUX \Data_Mem/U8845  ( .IN0(\Data_Mem/n8795 ), .IN1(\Data_Mem/n8794 ), .SEL(
        N28), .F(\Data_Mem/n8796 ) );
  MUX \Data_Mem/U8844  ( .IN0(o[528]), .IN1(o[560]), .SEL(N29), .F(
        \Data_Mem/n8795 ) );
  MUX \Data_Mem/U8843  ( .IN0(o[592]), .IN1(o[624]), .SEL(N29), .F(
        \Data_Mem/n8794 ) );
  MUX \Data_Mem/U8842  ( .IN0(\Data_Mem/n8792 ), .IN1(\Data_Mem/n8791 ), .SEL(
        N28), .F(\Data_Mem/n8793 ) );
  MUX \Data_Mem/U8841  ( .IN0(o[656]), .IN1(o[688]), .SEL(N29), .F(
        \Data_Mem/n8792 ) );
  MUX \Data_Mem/U8840  ( .IN0(o[720]), .IN1(o[752]), .SEL(N29), .F(
        \Data_Mem/n8791 ) );
  MUX \Data_Mem/U8839  ( .IN0(\Data_Mem/n8789 ), .IN1(\Data_Mem/n8786 ), .SEL(
        N27), .F(\Data_Mem/n8790 ) );
  MUX \Data_Mem/U8838  ( .IN0(\Data_Mem/n8788 ), .IN1(\Data_Mem/n8787 ), .SEL(
        N28), .F(\Data_Mem/n8789 ) );
  MUX \Data_Mem/U8837  ( .IN0(o[784]), .IN1(o[816]), .SEL(N29), .F(
        \Data_Mem/n8788 ) );
  MUX \Data_Mem/U8836  ( .IN0(o[848]), .IN1(o[880]), .SEL(N29), .F(
        \Data_Mem/n8787 ) );
  MUX \Data_Mem/U8835  ( .IN0(\Data_Mem/n8785 ), .IN1(\Data_Mem/n8784 ), .SEL(
        N28), .F(\Data_Mem/n8786 ) );
  MUX \Data_Mem/U8834  ( .IN0(o[912]), .IN1(o[944]), .SEL(N29), .F(
        \Data_Mem/n8785 ) );
  MUX \Data_Mem/U8833  ( .IN0(o[976]), .IN1(o[1008]), .SEL(N29), .F(
        \Data_Mem/n8784 ) );
  MUX \Data_Mem/U8832  ( .IN0(\Data_Mem/n8782 ), .IN1(\Data_Mem/n8767 ), .SEL(
        N25), .F(\Data_Mem/n8783 ) );
  MUX \Data_Mem/U8831  ( .IN0(\Data_Mem/n8781 ), .IN1(\Data_Mem/n8774 ), .SEL(
        N26), .F(\Data_Mem/n8782 ) );
  MUX \Data_Mem/U8830  ( .IN0(\Data_Mem/n8780 ), .IN1(\Data_Mem/n8777 ), .SEL(
        N27), .F(\Data_Mem/n8781 ) );
  MUX \Data_Mem/U8829  ( .IN0(\Data_Mem/n8779 ), .IN1(\Data_Mem/n8778 ), .SEL(
        N28), .F(\Data_Mem/n8780 ) );
  MUX \Data_Mem/U8828  ( .IN0(o[1040]), .IN1(o[1072]), .SEL(N29), .F(
        \Data_Mem/n8779 ) );
  MUX \Data_Mem/U8827  ( .IN0(o[1104]), .IN1(o[1136]), .SEL(N29), .F(
        \Data_Mem/n8778 ) );
  MUX \Data_Mem/U8826  ( .IN0(\Data_Mem/n8776 ), .IN1(\Data_Mem/n8775 ), .SEL(
        N28), .F(\Data_Mem/n8777 ) );
  MUX \Data_Mem/U8825  ( .IN0(o[1168]), .IN1(o[1200]), .SEL(N29), .F(
        \Data_Mem/n8776 ) );
  MUX \Data_Mem/U8824  ( .IN0(o[1232]), .IN1(o[1264]), .SEL(N29), .F(
        \Data_Mem/n8775 ) );
  MUX \Data_Mem/U8823  ( .IN0(\Data_Mem/n8773 ), .IN1(\Data_Mem/n8770 ), .SEL(
        N27), .F(\Data_Mem/n8774 ) );
  MUX \Data_Mem/U8822  ( .IN0(\Data_Mem/n8772 ), .IN1(\Data_Mem/n8771 ), .SEL(
        N28), .F(\Data_Mem/n8773 ) );
  MUX \Data_Mem/U8821  ( .IN0(o[1296]), .IN1(o[1328]), .SEL(N29), .F(
        \Data_Mem/n8772 ) );
  MUX \Data_Mem/U8820  ( .IN0(o[1360]), .IN1(o[1392]), .SEL(N29), .F(
        \Data_Mem/n8771 ) );
  MUX \Data_Mem/U8819  ( .IN0(\Data_Mem/n8769 ), .IN1(\Data_Mem/n8768 ), .SEL(
        N28), .F(\Data_Mem/n8770 ) );
  MUX \Data_Mem/U8818  ( .IN0(o[1424]), .IN1(o[1456]), .SEL(N29), .F(
        \Data_Mem/n8769 ) );
  MUX \Data_Mem/U8817  ( .IN0(o[1488]), .IN1(o[1520]), .SEL(N29), .F(
        \Data_Mem/n8768 ) );
  MUX \Data_Mem/U8816  ( .IN0(\Data_Mem/n8766 ), .IN1(\Data_Mem/n8759 ), .SEL(
        N26), .F(\Data_Mem/n8767 ) );
  MUX \Data_Mem/U8815  ( .IN0(\Data_Mem/n8765 ), .IN1(\Data_Mem/n8762 ), .SEL(
        N27), .F(\Data_Mem/n8766 ) );
  MUX \Data_Mem/U8814  ( .IN0(\Data_Mem/n8764 ), .IN1(\Data_Mem/n8763 ), .SEL(
        N28), .F(\Data_Mem/n8765 ) );
  MUX \Data_Mem/U8813  ( .IN0(o[1552]), .IN1(o[1584]), .SEL(N29), .F(
        \Data_Mem/n8764 ) );
  MUX \Data_Mem/U8812  ( .IN0(o[1616]), .IN1(o[1648]), .SEL(N29), .F(
        \Data_Mem/n8763 ) );
  MUX \Data_Mem/U8811  ( .IN0(\Data_Mem/n8761 ), .IN1(\Data_Mem/n8760 ), .SEL(
        N28), .F(\Data_Mem/n8762 ) );
  MUX \Data_Mem/U8810  ( .IN0(o[1680]), .IN1(o[1712]), .SEL(N29), .F(
        \Data_Mem/n8761 ) );
  MUX \Data_Mem/U8809  ( .IN0(o[1744]), .IN1(o[1776]), .SEL(N29), .F(
        \Data_Mem/n8760 ) );
  MUX \Data_Mem/U8808  ( .IN0(\Data_Mem/n8758 ), .IN1(\Data_Mem/n8755 ), .SEL(
        N27), .F(\Data_Mem/n8759 ) );
  MUX \Data_Mem/U8807  ( .IN0(\Data_Mem/n8757 ), .IN1(\Data_Mem/n8756 ), .SEL(
        N28), .F(\Data_Mem/n8758 ) );
  MUX \Data_Mem/U8806  ( .IN0(o[1808]), .IN1(o[1840]), .SEL(N29), .F(
        \Data_Mem/n8757 ) );
  MUX \Data_Mem/U8805  ( .IN0(o[1872]), .IN1(o[1904]), .SEL(N29), .F(
        \Data_Mem/n8756 ) );
  MUX \Data_Mem/U8804  ( .IN0(\Data_Mem/n8754 ), .IN1(\Data_Mem/n8753 ), .SEL(
        N28), .F(\Data_Mem/n8755 ) );
  MUX \Data_Mem/U8803  ( .IN0(o[1936]), .IN1(o[1968]), .SEL(N29), .F(
        \Data_Mem/n8754 ) );
  MUX \Data_Mem/U8802  ( .IN0(o[2000]), .IN1(o[2032]), .SEL(N29), .F(
        \Data_Mem/n8753 ) );
  MUX \Data_Mem/U8801  ( .IN0(\Data_Mem/n8752 ), .IN1(\Data_Mem/n8721 ), .SEL(
        N24), .F(\Data_Mem/N730 ) );
  MUX \Data_Mem/U8800  ( .IN0(\Data_Mem/n8751 ), .IN1(\Data_Mem/n8736 ), .SEL(
        N25), .F(\Data_Mem/n8752 ) );
  MUX \Data_Mem/U8799  ( .IN0(\Data_Mem/n8750 ), .IN1(\Data_Mem/n8743 ), .SEL(
        N26), .F(\Data_Mem/n8751 ) );
  MUX \Data_Mem/U8798  ( .IN0(\Data_Mem/n8749 ), .IN1(\Data_Mem/n8746 ), .SEL(
        N27), .F(\Data_Mem/n8750 ) );
  MUX \Data_Mem/U8797  ( .IN0(\Data_Mem/n8748 ), .IN1(\Data_Mem/n8747 ), .SEL(
        N28), .F(\Data_Mem/n8749 ) );
  MUX \Data_Mem/U8796  ( .IN0(o[15]), .IN1(o[47]), .SEL(N29), .F(
        \Data_Mem/n8748 ) );
  MUX \Data_Mem/U8795  ( .IN0(o[79]), .IN1(o[111]), .SEL(N29), .F(
        \Data_Mem/n8747 ) );
  MUX \Data_Mem/U8794  ( .IN0(\Data_Mem/n8745 ), .IN1(\Data_Mem/n8744 ), .SEL(
        N28), .F(\Data_Mem/n8746 ) );
  MUX \Data_Mem/U8793  ( .IN0(o[143]), .IN1(o[175]), .SEL(N29), .F(
        \Data_Mem/n8745 ) );
  MUX \Data_Mem/U8792  ( .IN0(o[207]), .IN1(o[239]), .SEL(N29), .F(
        \Data_Mem/n8744 ) );
  MUX \Data_Mem/U8791  ( .IN0(\Data_Mem/n8742 ), .IN1(\Data_Mem/n8739 ), .SEL(
        N27), .F(\Data_Mem/n8743 ) );
  MUX \Data_Mem/U8790  ( .IN0(\Data_Mem/n8741 ), .IN1(\Data_Mem/n8740 ), .SEL(
        N28), .F(\Data_Mem/n8742 ) );
  MUX \Data_Mem/U8789  ( .IN0(o[271]), .IN1(o[303]), .SEL(N29), .F(
        \Data_Mem/n8741 ) );
  MUX \Data_Mem/U8788  ( .IN0(o[335]), .IN1(o[367]), .SEL(N29), .F(
        \Data_Mem/n8740 ) );
  MUX \Data_Mem/U8787  ( .IN0(\Data_Mem/n8738 ), .IN1(\Data_Mem/n8737 ), .SEL(
        N28), .F(\Data_Mem/n8739 ) );
  MUX \Data_Mem/U8786  ( .IN0(o[399]), .IN1(o[431]), .SEL(N29), .F(
        \Data_Mem/n8738 ) );
  MUX \Data_Mem/U8785  ( .IN0(o[463]), .IN1(o[495]), .SEL(N29), .F(
        \Data_Mem/n8737 ) );
  MUX \Data_Mem/U8784  ( .IN0(\Data_Mem/n8735 ), .IN1(\Data_Mem/n8728 ), .SEL(
        N26), .F(\Data_Mem/n8736 ) );
  MUX \Data_Mem/U8783  ( .IN0(\Data_Mem/n8734 ), .IN1(\Data_Mem/n8731 ), .SEL(
        N27), .F(\Data_Mem/n8735 ) );
  MUX \Data_Mem/U8782  ( .IN0(\Data_Mem/n8733 ), .IN1(\Data_Mem/n8732 ), .SEL(
        N28), .F(\Data_Mem/n8734 ) );
  MUX \Data_Mem/U8781  ( .IN0(o[527]), .IN1(o[559]), .SEL(N29), .F(
        \Data_Mem/n8733 ) );
  MUX \Data_Mem/U8780  ( .IN0(o[591]), .IN1(o[623]), .SEL(N29), .F(
        \Data_Mem/n8732 ) );
  MUX \Data_Mem/U8779  ( .IN0(\Data_Mem/n8730 ), .IN1(\Data_Mem/n8729 ), .SEL(
        N28), .F(\Data_Mem/n8731 ) );
  MUX \Data_Mem/U8778  ( .IN0(o[655]), .IN1(o[687]), .SEL(N29), .F(
        \Data_Mem/n8730 ) );
  MUX \Data_Mem/U8777  ( .IN0(o[719]), .IN1(o[751]), .SEL(N29), .F(
        \Data_Mem/n8729 ) );
  MUX \Data_Mem/U8776  ( .IN0(\Data_Mem/n8727 ), .IN1(\Data_Mem/n8724 ), .SEL(
        N27), .F(\Data_Mem/n8728 ) );
  MUX \Data_Mem/U8775  ( .IN0(\Data_Mem/n8726 ), .IN1(\Data_Mem/n8725 ), .SEL(
        N28), .F(\Data_Mem/n8727 ) );
  MUX \Data_Mem/U8774  ( .IN0(o[783]), .IN1(o[815]), .SEL(N29), .F(
        \Data_Mem/n8726 ) );
  MUX \Data_Mem/U8773  ( .IN0(o[847]), .IN1(o[879]), .SEL(N29), .F(
        \Data_Mem/n8725 ) );
  MUX \Data_Mem/U8772  ( .IN0(\Data_Mem/n8723 ), .IN1(\Data_Mem/n8722 ), .SEL(
        N28), .F(\Data_Mem/n8724 ) );
  MUX \Data_Mem/U8771  ( .IN0(o[911]), .IN1(o[943]), .SEL(N29), .F(
        \Data_Mem/n8723 ) );
  MUX \Data_Mem/U8770  ( .IN0(o[975]), .IN1(o[1007]), .SEL(N29), .F(
        \Data_Mem/n8722 ) );
  MUX \Data_Mem/U8769  ( .IN0(\Data_Mem/n8720 ), .IN1(\Data_Mem/n8705 ), .SEL(
        N25), .F(\Data_Mem/n8721 ) );
  MUX \Data_Mem/U8768  ( .IN0(\Data_Mem/n8719 ), .IN1(\Data_Mem/n8712 ), .SEL(
        N26), .F(\Data_Mem/n8720 ) );
  MUX \Data_Mem/U8767  ( .IN0(\Data_Mem/n8718 ), .IN1(\Data_Mem/n8715 ), .SEL(
        N27), .F(\Data_Mem/n8719 ) );
  MUX \Data_Mem/U8766  ( .IN0(\Data_Mem/n8717 ), .IN1(\Data_Mem/n8716 ), .SEL(
        N28), .F(\Data_Mem/n8718 ) );
  MUX \Data_Mem/U8765  ( .IN0(o[1039]), .IN1(o[1071]), .SEL(N29), .F(
        \Data_Mem/n8717 ) );
  MUX \Data_Mem/U8764  ( .IN0(o[1103]), .IN1(o[1135]), .SEL(N29), .F(
        \Data_Mem/n8716 ) );
  MUX \Data_Mem/U8763  ( .IN0(\Data_Mem/n8714 ), .IN1(\Data_Mem/n8713 ), .SEL(
        N28), .F(\Data_Mem/n8715 ) );
  MUX \Data_Mem/U8762  ( .IN0(o[1167]), .IN1(o[1199]), .SEL(N29), .F(
        \Data_Mem/n8714 ) );
  MUX \Data_Mem/U8761  ( .IN0(o[1231]), .IN1(o[1263]), .SEL(N29), .F(
        \Data_Mem/n8713 ) );
  MUX \Data_Mem/U8760  ( .IN0(\Data_Mem/n8711 ), .IN1(\Data_Mem/n8708 ), .SEL(
        N27), .F(\Data_Mem/n8712 ) );
  MUX \Data_Mem/U8759  ( .IN0(\Data_Mem/n8710 ), .IN1(\Data_Mem/n8709 ), .SEL(
        N28), .F(\Data_Mem/n8711 ) );
  MUX \Data_Mem/U8758  ( .IN0(o[1295]), .IN1(o[1327]), .SEL(N29), .F(
        \Data_Mem/n8710 ) );
  MUX \Data_Mem/U8757  ( .IN0(o[1359]), .IN1(o[1391]), .SEL(N29), .F(
        \Data_Mem/n8709 ) );
  MUX \Data_Mem/U8756  ( .IN0(\Data_Mem/n8707 ), .IN1(\Data_Mem/n8706 ), .SEL(
        N28), .F(\Data_Mem/n8708 ) );
  MUX \Data_Mem/U8755  ( .IN0(o[1423]), .IN1(o[1455]), .SEL(N29), .F(
        \Data_Mem/n8707 ) );
  MUX \Data_Mem/U8754  ( .IN0(o[1487]), .IN1(o[1519]), .SEL(N29), .F(
        \Data_Mem/n8706 ) );
  MUX \Data_Mem/U8753  ( .IN0(\Data_Mem/n8704 ), .IN1(\Data_Mem/n8697 ), .SEL(
        N26), .F(\Data_Mem/n8705 ) );
  MUX \Data_Mem/U8752  ( .IN0(\Data_Mem/n8703 ), .IN1(\Data_Mem/n8700 ), .SEL(
        N27), .F(\Data_Mem/n8704 ) );
  MUX \Data_Mem/U8751  ( .IN0(\Data_Mem/n8702 ), .IN1(\Data_Mem/n8701 ), .SEL(
        N28), .F(\Data_Mem/n8703 ) );
  MUX \Data_Mem/U8750  ( .IN0(o[1551]), .IN1(o[1583]), .SEL(N29), .F(
        \Data_Mem/n8702 ) );
  MUX \Data_Mem/U8749  ( .IN0(o[1615]), .IN1(o[1647]), .SEL(N29), .F(
        \Data_Mem/n8701 ) );
  MUX \Data_Mem/U8748  ( .IN0(\Data_Mem/n8699 ), .IN1(\Data_Mem/n8698 ), .SEL(
        N28), .F(\Data_Mem/n8700 ) );
  MUX \Data_Mem/U8747  ( .IN0(o[1679]), .IN1(o[1711]), .SEL(N29), .F(
        \Data_Mem/n8699 ) );
  MUX \Data_Mem/U8746  ( .IN0(o[1743]), .IN1(o[1775]), .SEL(N29), .F(
        \Data_Mem/n8698 ) );
  MUX \Data_Mem/U8745  ( .IN0(\Data_Mem/n8696 ), .IN1(\Data_Mem/n8693 ), .SEL(
        N27), .F(\Data_Mem/n8697 ) );
  MUX \Data_Mem/U8744  ( .IN0(\Data_Mem/n8695 ), .IN1(\Data_Mem/n8694 ), .SEL(
        N28), .F(\Data_Mem/n8696 ) );
  MUX \Data_Mem/U8743  ( .IN0(o[1807]), .IN1(o[1839]), .SEL(N29), .F(
        \Data_Mem/n8695 ) );
  MUX \Data_Mem/U8742  ( .IN0(o[1871]), .IN1(o[1903]), .SEL(N29), .F(
        \Data_Mem/n8694 ) );
  MUX \Data_Mem/U8741  ( .IN0(\Data_Mem/n8692 ), .IN1(\Data_Mem/n8691 ), .SEL(
        N28), .F(\Data_Mem/n8693 ) );
  MUX \Data_Mem/U8740  ( .IN0(o[1935]), .IN1(o[1967]), .SEL(N29), .F(
        \Data_Mem/n8692 ) );
  MUX \Data_Mem/U8739  ( .IN0(o[1999]), .IN1(o[2031]), .SEL(N29), .F(
        \Data_Mem/n8691 ) );
  MUX \Data_Mem/U8738  ( .IN0(\Data_Mem/n8690 ), .IN1(\Data_Mem/n8659 ), .SEL(
        N24), .F(\Data_Mem/N731 ) );
  MUX \Data_Mem/U8737  ( .IN0(\Data_Mem/n8689 ), .IN1(\Data_Mem/n8674 ), .SEL(
        N25), .F(\Data_Mem/n8690 ) );
  MUX \Data_Mem/U8736  ( .IN0(\Data_Mem/n8688 ), .IN1(\Data_Mem/n8681 ), .SEL(
        N26), .F(\Data_Mem/n8689 ) );
  MUX \Data_Mem/U8735  ( .IN0(\Data_Mem/n8687 ), .IN1(\Data_Mem/n8684 ), .SEL(
        N27), .F(\Data_Mem/n8688 ) );
  MUX \Data_Mem/U8734  ( .IN0(\Data_Mem/n8686 ), .IN1(\Data_Mem/n8685 ), .SEL(
        N28), .F(\Data_Mem/n8687 ) );
  MUX \Data_Mem/U8733  ( .IN0(o[14]), .IN1(o[46]), .SEL(N29), .F(
        \Data_Mem/n8686 ) );
  MUX \Data_Mem/U8732  ( .IN0(o[78]), .IN1(o[110]), .SEL(N29), .F(
        \Data_Mem/n8685 ) );
  MUX \Data_Mem/U8731  ( .IN0(\Data_Mem/n8683 ), .IN1(\Data_Mem/n8682 ), .SEL(
        N28), .F(\Data_Mem/n8684 ) );
  MUX \Data_Mem/U8730  ( .IN0(o[142]), .IN1(o[174]), .SEL(N29), .F(
        \Data_Mem/n8683 ) );
  MUX \Data_Mem/U8729  ( .IN0(o[206]), .IN1(o[238]), .SEL(N29), .F(
        \Data_Mem/n8682 ) );
  MUX \Data_Mem/U8728  ( .IN0(\Data_Mem/n8680 ), .IN1(\Data_Mem/n8677 ), .SEL(
        N27), .F(\Data_Mem/n8681 ) );
  MUX \Data_Mem/U8727  ( .IN0(\Data_Mem/n8679 ), .IN1(\Data_Mem/n8678 ), .SEL(
        N28), .F(\Data_Mem/n8680 ) );
  MUX \Data_Mem/U8726  ( .IN0(o[270]), .IN1(o[302]), .SEL(N29), .F(
        \Data_Mem/n8679 ) );
  MUX \Data_Mem/U8725  ( .IN0(o[334]), .IN1(o[366]), .SEL(N29), .F(
        \Data_Mem/n8678 ) );
  MUX \Data_Mem/U8724  ( .IN0(\Data_Mem/n8676 ), .IN1(\Data_Mem/n8675 ), .SEL(
        N28), .F(\Data_Mem/n8677 ) );
  MUX \Data_Mem/U8723  ( .IN0(o[398]), .IN1(o[430]), .SEL(N29), .F(
        \Data_Mem/n8676 ) );
  MUX \Data_Mem/U8722  ( .IN0(o[462]), .IN1(o[494]), .SEL(N29), .F(
        \Data_Mem/n8675 ) );
  MUX \Data_Mem/U8721  ( .IN0(\Data_Mem/n8673 ), .IN1(\Data_Mem/n8666 ), .SEL(
        N26), .F(\Data_Mem/n8674 ) );
  MUX \Data_Mem/U8720  ( .IN0(\Data_Mem/n8672 ), .IN1(\Data_Mem/n8669 ), .SEL(
        N27), .F(\Data_Mem/n8673 ) );
  MUX \Data_Mem/U8719  ( .IN0(\Data_Mem/n8671 ), .IN1(\Data_Mem/n8670 ), .SEL(
        N28), .F(\Data_Mem/n8672 ) );
  MUX \Data_Mem/U8718  ( .IN0(o[526]), .IN1(o[558]), .SEL(N29), .F(
        \Data_Mem/n8671 ) );
  MUX \Data_Mem/U8717  ( .IN0(o[590]), .IN1(o[622]), .SEL(N29), .F(
        \Data_Mem/n8670 ) );
  MUX \Data_Mem/U8716  ( .IN0(\Data_Mem/n8668 ), .IN1(\Data_Mem/n8667 ), .SEL(
        N28), .F(\Data_Mem/n8669 ) );
  MUX \Data_Mem/U8715  ( .IN0(o[654]), .IN1(o[686]), .SEL(N29), .F(
        \Data_Mem/n8668 ) );
  MUX \Data_Mem/U8714  ( .IN0(o[718]), .IN1(o[750]), .SEL(N29), .F(
        \Data_Mem/n8667 ) );
  MUX \Data_Mem/U8713  ( .IN0(\Data_Mem/n8665 ), .IN1(\Data_Mem/n8662 ), .SEL(
        N27), .F(\Data_Mem/n8666 ) );
  MUX \Data_Mem/U8712  ( .IN0(\Data_Mem/n8664 ), .IN1(\Data_Mem/n8663 ), .SEL(
        N28), .F(\Data_Mem/n8665 ) );
  MUX \Data_Mem/U8711  ( .IN0(o[782]), .IN1(o[814]), .SEL(N29), .F(
        \Data_Mem/n8664 ) );
  MUX \Data_Mem/U8710  ( .IN0(o[846]), .IN1(o[878]), .SEL(N29), .F(
        \Data_Mem/n8663 ) );
  MUX \Data_Mem/U8709  ( .IN0(\Data_Mem/n8661 ), .IN1(\Data_Mem/n8660 ), .SEL(
        N28), .F(\Data_Mem/n8662 ) );
  MUX \Data_Mem/U8708  ( .IN0(o[910]), .IN1(o[942]), .SEL(N29), .F(
        \Data_Mem/n8661 ) );
  MUX \Data_Mem/U8707  ( .IN0(o[974]), .IN1(o[1006]), .SEL(N29), .F(
        \Data_Mem/n8660 ) );
  MUX \Data_Mem/U8706  ( .IN0(\Data_Mem/n8658 ), .IN1(\Data_Mem/n8643 ), .SEL(
        N25), .F(\Data_Mem/n8659 ) );
  MUX \Data_Mem/U8705  ( .IN0(\Data_Mem/n8657 ), .IN1(\Data_Mem/n8650 ), .SEL(
        N26), .F(\Data_Mem/n8658 ) );
  MUX \Data_Mem/U8704  ( .IN0(\Data_Mem/n8656 ), .IN1(\Data_Mem/n8653 ), .SEL(
        N27), .F(\Data_Mem/n8657 ) );
  MUX \Data_Mem/U8703  ( .IN0(\Data_Mem/n8655 ), .IN1(\Data_Mem/n8654 ), .SEL(
        N28), .F(\Data_Mem/n8656 ) );
  MUX \Data_Mem/U8702  ( .IN0(o[1038]), .IN1(o[1070]), .SEL(N29), .F(
        \Data_Mem/n8655 ) );
  MUX \Data_Mem/U8701  ( .IN0(o[1102]), .IN1(o[1134]), .SEL(N29), .F(
        \Data_Mem/n8654 ) );
  MUX \Data_Mem/U8700  ( .IN0(\Data_Mem/n8652 ), .IN1(\Data_Mem/n8651 ), .SEL(
        N28), .F(\Data_Mem/n8653 ) );
  MUX \Data_Mem/U8699  ( .IN0(o[1166]), .IN1(o[1198]), .SEL(N29), .F(
        \Data_Mem/n8652 ) );
  MUX \Data_Mem/U8698  ( .IN0(o[1230]), .IN1(o[1262]), .SEL(N29), .F(
        \Data_Mem/n8651 ) );
  MUX \Data_Mem/U8697  ( .IN0(\Data_Mem/n8649 ), .IN1(\Data_Mem/n8646 ), .SEL(
        N27), .F(\Data_Mem/n8650 ) );
  MUX \Data_Mem/U8696  ( .IN0(\Data_Mem/n8648 ), .IN1(\Data_Mem/n8647 ), .SEL(
        N28), .F(\Data_Mem/n8649 ) );
  MUX \Data_Mem/U8695  ( .IN0(o[1294]), .IN1(o[1326]), .SEL(N29), .F(
        \Data_Mem/n8648 ) );
  MUX \Data_Mem/U8694  ( .IN0(o[1358]), .IN1(o[1390]), .SEL(N29), .F(
        \Data_Mem/n8647 ) );
  MUX \Data_Mem/U8693  ( .IN0(\Data_Mem/n8645 ), .IN1(\Data_Mem/n8644 ), .SEL(
        N28), .F(\Data_Mem/n8646 ) );
  MUX \Data_Mem/U8692  ( .IN0(o[1422]), .IN1(o[1454]), .SEL(N29), .F(
        \Data_Mem/n8645 ) );
  MUX \Data_Mem/U8691  ( .IN0(o[1486]), .IN1(o[1518]), .SEL(N29), .F(
        \Data_Mem/n8644 ) );
  MUX \Data_Mem/U8690  ( .IN0(\Data_Mem/n8642 ), .IN1(\Data_Mem/n8635 ), .SEL(
        N26), .F(\Data_Mem/n8643 ) );
  MUX \Data_Mem/U8689  ( .IN0(\Data_Mem/n8641 ), .IN1(\Data_Mem/n8638 ), .SEL(
        N27), .F(\Data_Mem/n8642 ) );
  MUX \Data_Mem/U8688  ( .IN0(\Data_Mem/n8640 ), .IN1(\Data_Mem/n8639 ), .SEL(
        N28), .F(\Data_Mem/n8641 ) );
  MUX \Data_Mem/U8687  ( .IN0(o[1550]), .IN1(o[1582]), .SEL(N29), .F(
        \Data_Mem/n8640 ) );
  MUX \Data_Mem/U8686  ( .IN0(o[1614]), .IN1(o[1646]), .SEL(N29), .F(
        \Data_Mem/n8639 ) );
  MUX \Data_Mem/U8685  ( .IN0(\Data_Mem/n8637 ), .IN1(\Data_Mem/n8636 ), .SEL(
        N28), .F(\Data_Mem/n8638 ) );
  MUX \Data_Mem/U8684  ( .IN0(o[1678]), .IN1(o[1710]), .SEL(N29), .F(
        \Data_Mem/n8637 ) );
  MUX \Data_Mem/U8683  ( .IN0(o[1742]), .IN1(o[1774]), .SEL(N29), .F(
        \Data_Mem/n8636 ) );
  MUX \Data_Mem/U8682  ( .IN0(\Data_Mem/n8634 ), .IN1(\Data_Mem/n8631 ), .SEL(
        N27), .F(\Data_Mem/n8635 ) );
  MUX \Data_Mem/U8681  ( .IN0(\Data_Mem/n8633 ), .IN1(\Data_Mem/n8632 ), .SEL(
        N28), .F(\Data_Mem/n8634 ) );
  MUX \Data_Mem/U8680  ( .IN0(o[1806]), .IN1(o[1838]), .SEL(N29), .F(
        \Data_Mem/n8633 ) );
  MUX \Data_Mem/U8679  ( .IN0(o[1870]), .IN1(o[1902]), .SEL(N29), .F(
        \Data_Mem/n8632 ) );
  MUX \Data_Mem/U8678  ( .IN0(\Data_Mem/n8630 ), .IN1(\Data_Mem/n8629 ), .SEL(
        N28), .F(\Data_Mem/n8631 ) );
  MUX \Data_Mem/U8677  ( .IN0(o[1934]), .IN1(o[1966]), .SEL(N29), .F(
        \Data_Mem/n8630 ) );
  MUX \Data_Mem/U8676  ( .IN0(o[1998]), .IN1(o[2030]), .SEL(N29), .F(
        \Data_Mem/n8629 ) );
  MUX \Data_Mem/U8675  ( .IN0(\Data_Mem/n8628 ), .IN1(\Data_Mem/n8597 ), .SEL(
        N24), .F(\Data_Mem/N732 ) );
  MUX \Data_Mem/U8674  ( .IN0(\Data_Mem/n8627 ), .IN1(\Data_Mem/n8612 ), .SEL(
        N25), .F(\Data_Mem/n8628 ) );
  MUX \Data_Mem/U8673  ( .IN0(\Data_Mem/n8626 ), .IN1(\Data_Mem/n8619 ), .SEL(
        N26), .F(\Data_Mem/n8627 ) );
  MUX \Data_Mem/U8672  ( .IN0(\Data_Mem/n8625 ), .IN1(\Data_Mem/n8622 ), .SEL(
        N27), .F(\Data_Mem/n8626 ) );
  MUX \Data_Mem/U8671  ( .IN0(\Data_Mem/n8624 ), .IN1(\Data_Mem/n8623 ), .SEL(
        N28), .F(\Data_Mem/n8625 ) );
  MUX \Data_Mem/U8670  ( .IN0(o[13]), .IN1(o[45]), .SEL(N29), .F(
        \Data_Mem/n8624 ) );
  MUX \Data_Mem/U8669  ( .IN0(o[77]), .IN1(o[109]), .SEL(N29), .F(
        \Data_Mem/n8623 ) );
  MUX \Data_Mem/U8668  ( .IN0(\Data_Mem/n8621 ), .IN1(\Data_Mem/n8620 ), .SEL(
        N28), .F(\Data_Mem/n8622 ) );
  MUX \Data_Mem/U8667  ( .IN0(o[141]), .IN1(o[173]), .SEL(N29), .F(
        \Data_Mem/n8621 ) );
  MUX \Data_Mem/U8666  ( .IN0(o[205]), .IN1(o[237]), .SEL(N29), .F(
        \Data_Mem/n8620 ) );
  MUX \Data_Mem/U8665  ( .IN0(\Data_Mem/n8618 ), .IN1(\Data_Mem/n8615 ), .SEL(
        N27), .F(\Data_Mem/n8619 ) );
  MUX \Data_Mem/U8664  ( .IN0(\Data_Mem/n8617 ), .IN1(\Data_Mem/n8616 ), .SEL(
        N28), .F(\Data_Mem/n8618 ) );
  MUX \Data_Mem/U8663  ( .IN0(o[269]), .IN1(o[301]), .SEL(N29), .F(
        \Data_Mem/n8617 ) );
  MUX \Data_Mem/U8662  ( .IN0(o[333]), .IN1(o[365]), .SEL(N29), .F(
        \Data_Mem/n8616 ) );
  MUX \Data_Mem/U8661  ( .IN0(\Data_Mem/n8614 ), .IN1(\Data_Mem/n8613 ), .SEL(
        N28), .F(\Data_Mem/n8615 ) );
  MUX \Data_Mem/U8660  ( .IN0(o[397]), .IN1(o[429]), .SEL(N29), .F(
        \Data_Mem/n8614 ) );
  MUX \Data_Mem/U8659  ( .IN0(o[461]), .IN1(o[493]), .SEL(N29), .F(
        \Data_Mem/n8613 ) );
  MUX \Data_Mem/U8658  ( .IN0(\Data_Mem/n8611 ), .IN1(\Data_Mem/n8604 ), .SEL(
        N26), .F(\Data_Mem/n8612 ) );
  MUX \Data_Mem/U8657  ( .IN0(\Data_Mem/n8610 ), .IN1(\Data_Mem/n8607 ), .SEL(
        N27), .F(\Data_Mem/n8611 ) );
  MUX \Data_Mem/U8656  ( .IN0(\Data_Mem/n8609 ), .IN1(\Data_Mem/n8608 ), .SEL(
        N28), .F(\Data_Mem/n8610 ) );
  MUX \Data_Mem/U8655  ( .IN0(o[525]), .IN1(o[557]), .SEL(N29), .F(
        \Data_Mem/n8609 ) );
  MUX \Data_Mem/U8654  ( .IN0(o[589]), .IN1(o[621]), .SEL(N29), .F(
        \Data_Mem/n8608 ) );
  MUX \Data_Mem/U8653  ( .IN0(\Data_Mem/n8606 ), .IN1(\Data_Mem/n8605 ), .SEL(
        N28), .F(\Data_Mem/n8607 ) );
  MUX \Data_Mem/U8652  ( .IN0(o[653]), .IN1(o[685]), .SEL(N29), .F(
        \Data_Mem/n8606 ) );
  MUX \Data_Mem/U8651  ( .IN0(o[717]), .IN1(o[749]), .SEL(N29), .F(
        \Data_Mem/n8605 ) );
  MUX \Data_Mem/U8650  ( .IN0(\Data_Mem/n8603 ), .IN1(\Data_Mem/n8600 ), .SEL(
        N27), .F(\Data_Mem/n8604 ) );
  MUX \Data_Mem/U8649  ( .IN0(\Data_Mem/n8602 ), .IN1(\Data_Mem/n8601 ), .SEL(
        N28), .F(\Data_Mem/n8603 ) );
  MUX \Data_Mem/U8648  ( .IN0(o[781]), .IN1(o[813]), .SEL(N29), .F(
        \Data_Mem/n8602 ) );
  MUX \Data_Mem/U8647  ( .IN0(o[845]), .IN1(o[877]), .SEL(N29), .F(
        \Data_Mem/n8601 ) );
  MUX \Data_Mem/U8646  ( .IN0(\Data_Mem/n8599 ), .IN1(\Data_Mem/n8598 ), .SEL(
        N28), .F(\Data_Mem/n8600 ) );
  MUX \Data_Mem/U8645  ( .IN0(o[909]), .IN1(o[941]), .SEL(N29), .F(
        \Data_Mem/n8599 ) );
  MUX \Data_Mem/U8644  ( .IN0(o[973]), .IN1(o[1005]), .SEL(N29), .F(
        \Data_Mem/n8598 ) );
  MUX \Data_Mem/U8643  ( .IN0(\Data_Mem/n8596 ), .IN1(\Data_Mem/n8581 ), .SEL(
        N25), .F(\Data_Mem/n8597 ) );
  MUX \Data_Mem/U8642  ( .IN0(\Data_Mem/n8595 ), .IN1(\Data_Mem/n8588 ), .SEL(
        N26), .F(\Data_Mem/n8596 ) );
  MUX \Data_Mem/U8641  ( .IN0(\Data_Mem/n8594 ), .IN1(\Data_Mem/n8591 ), .SEL(
        N27), .F(\Data_Mem/n8595 ) );
  MUX \Data_Mem/U8640  ( .IN0(\Data_Mem/n8593 ), .IN1(\Data_Mem/n8592 ), .SEL(
        N28), .F(\Data_Mem/n8594 ) );
  MUX \Data_Mem/U8639  ( .IN0(o[1037]), .IN1(o[1069]), .SEL(N29), .F(
        \Data_Mem/n8593 ) );
  MUX \Data_Mem/U8638  ( .IN0(o[1101]), .IN1(o[1133]), .SEL(N29), .F(
        \Data_Mem/n8592 ) );
  MUX \Data_Mem/U8637  ( .IN0(\Data_Mem/n8590 ), .IN1(\Data_Mem/n8589 ), .SEL(
        N28), .F(\Data_Mem/n8591 ) );
  MUX \Data_Mem/U8636  ( .IN0(o[1165]), .IN1(o[1197]), .SEL(N29), .F(
        \Data_Mem/n8590 ) );
  MUX \Data_Mem/U8635  ( .IN0(o[1229]), .IN1(o[1261]), .SEL(N29), .F(
        \Data_Mem/n8589 ) );
  MUX \Data_Mem/U8634  ( .IN0(\Data_Mem/n8587 ), .IN1(\Data_Mem/n8584 ), .SEL(
        N27), .F(\Data_Mem/n8588 ) );
  MUX \Data_Mem/U8633  ( .IN0(\Data_Mem/n8586 ), .IN1(\Data_Mem/n8585 ), .SEL(
        N28), .F(\Data_Mem/n8587 ) );
  MUX \Data_Mem/U8632  ( .IN0(o[1293]), .IN1(o[1325]), .SEL(N29), .F(
        \Data_Mem/n8586 ) );
  MUX \Data_Mem/U8631  ( .IN0(o[1357]), .IN1(o[1389]), .SEL(N29), .F(
        \Data_Mem/n8585 ) );
  MUX \Data_Mem/U8630  ( .IN0(\Data_Mem/n8583 ), .IN1(\Data_Mem/n8582 ), .SEL(
        N28), .F(\Data_Mem/n8584 ) );
  MUX \Data_Mem/U8629  ( .IN0(o[1421]), .IN1(o[1453]), .SEL(N29), .F(
        \Data_Mem/n8583 ) );
  MUX \Data_Mem/U8628  ( .IN0(o[1485]), .IN1(o[1517]), .SEL(N29), .F(
        \Data_Mem/n8582 ) );
  MUX \Data_Mem/U8627  ( .IN0(\Data_Mem/n8580 ), .IN1(\Data_Mem/n8573 ), .SEL(
        N26), .F(\Data_Mem/n8581 ) );
  MUX \Data_Mem/U8626  ( .IN0(\Data_Mem/n8579 ), .IN1(\Data_Mem/n8576 ), .SEL(
        N27), .F(\Data_Mem/n8580 ) );
  MUX \Data_Mem/U8625  ( .IN0(\Data_Mem/n8578 ), .IN1(\Data_Mem/n8577 ), .SEL(
        N28), .F(\Data_Mem/n8579 ) );
  MUX \Data_Mem/U8624  ( .IN0(o[1549]), .IN1(o[1581]), .SEL(N29), .F(
        \Data_Mem/n8578 ) );
  MUX \Data_Mem/U8623  ( .IN0(o[1613]), .IN1(o[1645]), .SEL(N29), .F(
        \Data_Mem/n8577 ) );
  MUX \Data_Mem/U8622  ( .IN0(\Data_Mem/n8575 ), .IN1(\Data_Mem/n8574 ), .SEL(
        N28), .F(\Data_Mem/n8576 ) );
  MUX \Data_Mem/U8621  ( .IN0(o[1677]), .IN1(o[1709]), .SEL(N29), .F(
        \Data_Mem/n8575 ) );
  MUX \Data_Mem/U8620  ( .IN0(o[1741]), .IN1(o[1773]), .SEL(N29), .F(
        \Data_Mem/n8574 ) );
  MUX \Data_Mem/U8619  ( .IN0(\Data_Mem/n8572 ), .IN1(\Data_Mem/n8569 ), .SEL(
        N27), .F(\Data_Mem/n8573 ) );
  MUX \Data_Mem/U8618  ( .IN0(\Data_Mem/n8571 ), .IN1(\Data_Mem/n8570 ), .SEL(
        N28), .F(\Data_Mem/n8572 ) );
  MUX \Data_Mem/U8617  ( .IN0(o[1805]), .IN1(o[1837]), .SEL(N29), .F(
        \Data_Mem/n8571 ) );
  MUX \Data_Mem/U8616  ( .IN0(o[1869]), .IN1(o[1901]), .SEL(N29), .F(
        \Data_Mem/n8570 ) );
  MUX \Data_Mem/U8615  ( .IN0(\Data_Mem/n8568 ), .IN1(\Data_Mem/n8567 ), .SEL(
        N28), .F(\Data_Mem/n8569 ) );
  MUX \Data_Mem/U8614  ( .IN0(o[1933]), .IN1(o[1965]), .SEL(N29), .F(
        \Data_Mem/n8568 ) );
  MUX \Data_Mem/U8613  ( .IN0(o[1997]), .IN1(o[2029]), .SEL(N29), .F(
        \Data_Mem/n8567 ) );
  MUX \Data_Mem/U8612  ( .IN0(\Data_Mem/n8566 ), .IN1(\Data_Mem/n8535 ), .SEL(
        N24), .F(\Data_Mem/N733 ) );
  MUX \Data_Mem/U8611  ( .IN0(\Data_Mem/n8565 ), .IN1(\Data_Mem/n8550 ), .SEL(
        N25), .F(\Data_Mem/n8566 ) );
  MUX \Data_Mem/U8610  ( .IN0(\Data_Mem/n8564 ), .IN1(\Data_Mem/n8557 ), .SEL(
        N26), .F(\Data_Mem/n8565 ) );
  MUX \Data_Mem/U8609  ( .IN0(\Data_Mem/n8563 ), .IN1(\Data_Mem/n8560 ), .SEL(
        N27), .F(\Data_Mem/n8564 ) );
  MUX \Data_Mem/U8608  ( .IN0(\Data_Mem/n8562 ), .IN1(\Data_Mem/n8561 ), .SEL(
        N28), .F(\Data_Mem/n8563 ) );
  MUX \Data_Mem/U8607  ( .IN0(o[12]), .IN1(o[44]), .SEL(N29), .F(
        \Data_Mem/n8562 ) );
  MUX \Data_Mem/U8606  ( .IN0(o[76]), .IN1(o[108]), .SEL(N29), .F(
        \Data_Mem/n8561 ) );
  MUX \Data_Mem/U8605  ( .IN0(\Data_Mem/n8559 ), .IN1(\Data_Mem/n8558 ), .SEL(
        N28), .F(\Data_Mem/n8560 ) );
  MUX \Data_Mem/U8604  ( .IN0(o[140]), .IN1(o[172]), .SEL(N29), .F(
        \Data_Mem/n8559 ) );
  MUX \Data_Mem/U8603  ( .IN0(o[204]), .IN1(o[236]), .SEL(N29), .F(
        \Data_Mem/n8558 ) );
  MUX \Data_Mem/U8602  ( .IN0(\Data_Mem/n8556 ), .IN1(\Data_Mem/n8553 ), .SEL(
        N27), .F(\Data_Mem/n8557 ) );
  MUX \Data_Mem/U8601  ( .IN0(\Data_Mem/n8555 ), .IN1(\Data_Mem/n8554 ), .SEL(
        N28), .F(\Data_Mem/n8556 ) );
  MUX \Data_Mem/U8600  ( .IN0(o[268]), .IN1(o[300]), .SEL(N29), .F(
        \Data_Mem/n8555 ) );
  MUX \Data_Mem/U8599  ( .IN0(o[332]), .IN1(o[364]), .SEL(N29), .F(
        \Data_Mem/n8554 ) );
  MUX \Data_Mem/U8598  ( .IN0(\Data_Mem/n8552 ), .IN1(\Data_Mem/n8551 ), .SEL(
        N28), .F(\Data_Mem/n8553 ) );
  MUX \Data_Mem/U8597  ( .IN0(o[396]), .IN1(o[428]), .SEL(N29), .F(
        \Data_Mem/n8552 ) );
  MUX \Data_Mem/U8596  ( .IN0(o[460]), .IN1(o[492]), .SEL(N29), .F(
        \Data_Mem/n8551 ) );
  MUX \Data_Mem/U8595  ( .IN0(\Data_Mem/n8549 ), .IN1(\Data_Mem/n8542 ), .SEL(
        N26), .F(\Data_Mem/n8550 ) );
  MUX \Data_Mem/U8594  ( .IN0(\Data_Mem/n8548 ), .IN1(\Data_Mem/n8545 ), .SEL(
        N27), .F(\Data_Mem/n8549 ) );
  MUX \Data_Mem/U8593  ( .IN0(\Data_Mem/n8547 ), .IN1(\Data_Mem/n8546 ), .SEL(
        N28), .F(\Data_Mem/n8548 ) );
  MUX \Data_Mem/U8592  ( .IN0(o[524]), .IN1(o[556]), .SEL(N29), .F(
        \Data_Mem/n8547 ) );
  MUX \Data_Mem/U8591  ( .IN0(o[588]), .IN1(o[620]), .SEL(N29), .F(
        \Data_Mem/n8546 ) );
  MUX \Data_Mem/U8590  ( .IN0(\Data_Mem/n8544 ), .IN1(\Data_Mem/n8543 ), .SEL(
        N28), .F(\Data_Mem/n8545 ) );
  MUX \Data_Mem/U8589  ( .IN0(o[652]), .IN1(o[684]), .SEL(N29), .F(
        \Data_Mem/n8544 ) );
  MUX \Data_Mem/U8588  ( .IN0(o[716]), .IN1(o[748]), .SEL(N29), .F(
        \Data_Mem/n8543 ) );
  MUX \Data_Mem/U8587  ( .IN0(\Data_Mem/n8541 ), .IN1(\Data_Mem/n8538 ), .SEL(
        N27), .F(\Data_Mem/n8542 ) );
  MUX \Data_Mem/U8586  ( .IN0(\Data_Mem/n8540 ), .IN1(\Data_Mem/n8539 ), .SEL(
        N28), .F(\Data_Mem/n8541 ) );
  MUX \Data_Mem/U8585  ( .IN0(o[780]), .IN1(o[812]), .SEL(N29), .F(
        \Data_Mem/n8540 ) );
  MUX \Data_Mem/U8584  ( .IN0(o[844]), .IN1(o[876]), .SEL(N29), .F(
        \Data_Mem/n8539 ) );
  MUX \Data_Mem/U8583  ( .IN0(\Data_Mem/n8537 ), .IN1(\Data_Mem/n8536 ), .SEL(
        N28), .F(\Data_Mem/n8538 ) );
  MUX \Data_Mem/U8582  ( .IN0(o[908]), .IN1(o[940]), .SEL(N29), .F(
        \Data_Mem/n8537 ) );
  MUX \Data_Mem/U8581  ( .IN0(o[972]), .IN1(o[1004]), .SEL(N29), .F(
        \Data_Mem/n8536 ) );
  MUX \Data_Mem/U8580  ( .IN0(\Data_Mem/n8534 ), .IN1(\Data_Mem/n8519 ), .SEL(
        N25), .F(\Data_Mem/n8535 ) );
  MUX \Data_Mem/U8579  ( .IN0(\Data_Mem/n8533 ), .IN1(\Data_Mem/n8526 ), .SEL(
        N26), .F(\Data_Mem/n8534 ) );
  MUX \Data_Mem/U8578  ( .IN0(\Data_Mem/n8532 ), .IN1(\Data_Mem/n8529 ), .SEL(
        N27), .F(\Data_Mem/n8533 ) );
  MUX \Data_Mem/U8577  ( .IN0(\Data_Mem/n8531 ), .IN1(\Data_Mem/n8530 ), .SEL(
        N28), .F(\Data_Mem/n8532 ) );
  MUX \Data_Mem/U8576  ( .IN0(o[1036]), .IN1(o[1068]), .SEL(N29), .F(
        \Data_Mem/n8531 ) );
  MUX \Data_Mem/U8575  ( .IN0(o[1100]), .IN1(o[1132]), .SEL(N29), .F(
        \Data_Mem/n8530 ) );
  MUX \Data_Mem/U8574  ( .IN0(\Data_Mem/n8528 ), .IN1(\Data_Mem/n8527 ), .SEL(
        N28), .F(\Data_Mem/n8529 ) );
  MUX \Data_Mem/U8573  ( .IN0(o[1164]), .IN1(o[1196]), .SEL(N29), .F(
        \Data_Mem/n8528 ) );
  MUX \Data_Mem/U8572  ( .IN0(o[1228]), .IN1(o[1260]), .SEL(N29), .F(
        \Data_Mem/n8527 ) );
  MUX \Data_Mem/U8571  ( .IN0(\Data_Mem/n8525 ), .IN1(\Data_Mem/n8522 ), .SEL(
        N27), .F(\Data_Mem/n8526 ) );
  MUX \Data_Mem/U8570  ( .IN0(\Data_Mem/n8524 ), .IN1(\Data_Mem/n8523 ), .SEL(
        N28), .F(\Data_Mem/n8525 ) );
  MUX \Data_Mem/U8569  ( .IN0(o[1292]), .IN1(o[1324]), .SEL(N29), .F(
        \Data_Mem/n8524 ) );
  MUX \Data_Mem/U8568  ( .IN0(o[1356]), .IN1(o[1388]), .SEL(N29), .F(
        \Data_Mem/n8523 ) );
  MUX \Data_Mem/U8567  ( .IN0(\Data_Mem/n8521 ), .IN1(\Data_Mem/n8520 ), .SEL(
        N28), .F(\Data_Mem/n8522 ) );
  MUX \Data_Mem/U8566  ( .IN0(o[1420]), .IN1(o[1452]), .SEL(N29), .F(
        \Data_Mem/n8521 ) );
  MUX \Data_Mem/U8565  ( .IN0(o[1484]), .IN1(o[1516]), .SEL(N29), .F(
        \Data_Mem/n8520 ) );
  MUX \Data_Mem/U8564  ( .IN0(\Data_Mem/n8518 ), .IN1(\Data_Mem/n8511 ), .SEL(
        N26), .F(\Data_Mem/n8519 ) );
  MUX \Data_Mem/U8563  ( .IN0(\Data_Mem/n8517 ), .IN1(\Data_Mem/n8514 ), .SEL(
        N27), .F(\Data_Mem/n8518 ) );
  MUX \Data_Mem/U8562  ( .IN0(\Data_Mem/n8516 ), .IN1(\Data_Mem/n8515 ), .SEL(
        N28), .F(\Data_Mem/n8517 ) );
  MUX \Data_Mem/U8561  ( .IN0(o[1548]), .IN1(o[1580]), .SEL(N29), .F(
        \Data_Mem/n8516 ) );
  MUX \Data_Mem/U8560  ( .IN0(o[1612]), .IN1(o[1644]), .SEL(N29), .F(
        \Data_Mem/n8515 ) );
  MUX \Data_Mem/U8559  ( .IN0(\Data_Mem/n8513 ), .IN1(\Data_Mem/n8512 ), .SEL(
        N28), .F(\Data_Mem/n8514 ) );
  MUX \Data_Mem/U8558  ( .IN0(o[1676]), .IN1(o[1708]), .SEL(N29), .F(
        \Data_Mem/n8513 ) );
  MUX \Data_Mem/U8557  ( .IN0(o[1740]), .IN1(o[1772]), .SEL(N29), .F(
        \Data_Mem/n8512 ) );
  MUX \Data_Mem/U8556  ( .IN0(\Data_Mem/n8510 ), .IN1(\Data_Mem/n8507 ), .SEL(
        N27), .F(\Data_Mem/n8511 ) );
  MUX \Data_Mem/U8555  ( .IN0(\Data_Mem/n8509 ), .IN1(\Data_Mem/n8508 ), .SEL(
        N28), .F(\Data_Mem/n8510 ) );
  MUX \Data_Mem/U8554  ( .IN0(o[1804]), .IN1(o[1836]), .SEL(N29), .F(
        \Data_Mem/n8509 ) );
  MUX \Data_Mem/U8553  ( .IN0(o[1868]), .IN1(o[1900]), .SEL(N29), .F(
        \Data_Mem/n8508 ) );
  MUX \Data_Mem/U8552  ( .IN0(\Data_Mem/n8506 ), .IN1(\Data_Mem/n8505 ), .SEL(
        N28), .F(\Data_Mem/n8507 ) );
  MUX \Data_Mem/U8551  ( .IN0(o[1932]), .IN1(o[1964]), .SEL(N29), .F(
        \Data_Mem/n8506 ) );
  MUX \Data_Mem/U8550  ( .IN0(o[1996]), .IN1(o[2028]), .SEL(N29), .F(
        \Data_Mem/n8505 ) );
  MUX \Data_Mem/U8549  ( .IN0(\Data_Mem/n8504 ), .IN1(\Data_Mem/n8473 ), .SEL(
        N24), .F(\Data_Mem/N734 ) );
  MUX \Data_Mem/U8548  ( .IN0(\Data_Mem/n8503 ), .IN1(\Data_Mem/n8488 ), .SEL(
        N25), .F(\Data_Mem/n8504 ) );
  MUX \Data_Mem/U8547  ( .IN0(\Data_Mem/n8502 ), .IN1(\Data_Mem/n8495 ), .SEL(
        N26), .F(\Data_Mem/n8503 ) );
  MUX \Data_Mem/U8546  ( .IN0(\Data_Mem/n8501 ), .IN1(\Data_Mem/n8498 ), .SEL(
        N27), .F(\Data_Mem/n8502 ) );
  MUX \Data_Mem/U8545  ( .IN0(\Data_Mem/n8500 ), .IN1(\Data_Mem/n8499 ), .SEL(
        N28), .F(\Data_Mem/n8501 ) );
  MUX \Data_Mem/U8544  ( .IN0(o[11]), .IN1(o[43]), .SEL(N29), .F(
        \Data_Mem/n8500 ) );
  MUX \Data_Mem/U8543  ( .IN0(o[75]), .IN1(o[107]), .SEL(N29), .F(
        \Data_Mem/n8499 ) );
  MUX \Data_Mem/U8542  ( .IN0(\Data_Mem/n8497 ), .IN1(\Data_Mem/n8496 ), .SEL(
        N28), .F(\Data_Mem/n8498 ) );
  MUX \Data_Mem/U8541  ( .IN0(o[139]), .IN1(o[171]), .SEL(N29), .F(
        \Data_Mem/n8497 ) );
  MUX \Data_Mem/U8540  ( .IN0(o[203]), .IN1(o[235]), .SEL(N29), .F(
        \Data_Mem/n8496 ) );
  MUX \Data_Mem/U8539  ( .IN0(\Data_Mem/n8494 ), .IN1(\Data_Mem/n8491 ), .SEL(
        N27), .F(\Data_Mem/n8495 ) );
  MUX \Data_Mem/U8538  ( .IN0(\Data_Mem/n8493 ), .IN1(\Data_Mem/n8492 ), .SEL(
        N28), .F(\Data_Mem/n8494 ) );
  MUX \Data_Mem/U8537  ( .IN0(o[267]), .IN1(o[299]), .SEL(N29), .F(
        \Data_Mem/n8493 ) );
  MUX \Data_Mem/U8536  ( .IN0(o[331]), .IN1(o[363]), .SEL(N29), .F(
        \Data_Mem/n8492 ) );
  MUX \Data_Mem/U8535  ( .IN0(\Data_Mem/n8490 ), .IN1(\Data_Mem/n8489 ), .SEL(
        N28), .F(\Data_Mem/n8491 ) );
  MUX \Data_Mem/U8534  ( .IN0(o[395]), .IN1(o[427]), .SEL(N29), .F(
        \Data_Mem/n8490 ) );
  MUX \Data_Mem/U8533  ( .IN0(o[459]), .IN1(o[491]), .SEL(N29), .F(
        \Data_Mem/n8489 ) );
  MUX \Data_Mem/U8532  ( .IN0(\Data_Mem/n8487 ), .IN1(\Data_Mem/n8480 ), .SEL(
        N26), .F(\Data_Mem/n8488 ) );
  MUX \Data_Mem/U8531  ( .IN0(\Data_Mem/n8486 ), .IN1(\Data_Mem/n8483 ), .SEL(
        N27), .F(\Data_Mem/n8487 ) );
  MUX \Data_Mem/U8530  ( .IN0(\Data_Mem/n8485 ), .IN1(\Data_Mem/n8484 ), .SEL(
        N28), .F(\Data_Mem/n8486 ) );
  MUX \Data_Mem/U8529  ( .IN0(o[523]), .IN1(o[555]), .SEL(N29), .F(
        \Data_Mem/n8485 ) );
  MUX \Data_Mem/U8528  ( .IN0(o[587]), .IN1(o[619]), .SEL(N29), .F(
        \Data_Mem/n8484 ) );
  MUX \Data_Mem/U8527  ( .IN0(\Data_Mem/n8482 ), .IN1(\Data_Mem/n8481 ), .SEL(
        N28), .F(\Data_Mem/n8483 ) );
  MUX \Data_Mem/U8526  ( .IN0(o[651]), .IN1(o[683]), .SEL(N29), .F(
        \Data_Mem/n8482 ) );
  MUX \Data_Mem/U8525  ( .IN0(o[715]), .IN1(o[747]), .SEL(N29), .F(
        \Data_Mem/n8481 ) );
  MUX \Data_Mem/U8524  ( .IN0(\Data_Mem/n8479 ), .IN1(\Data_Mem/n8476 ), .SEL(
        N27), .F(\Data_Mem/n8480 ) );
  MUX \Data_Mem/U8523  ( .IN0(\Data_Mem/n8478 ), .IN1(\Data_Mem/n8477 ), .SEL(
        N28), .F(\Data_Mem/n8479 ) );
  MUX \Data_Mem/U8522  ( .IN0(o[779]), .IN1(o[811]), .SEL(N29), .F(
        \Data_Mem/n8478 ) );
  MUX \Data_Mem/U8521  ( .IN0(o[843]), .IN1(o[875]), .SEL(N29), .F(
        \Data_Mem/n8477 ) );
  MUX \Data_Mem/U8520  ( .IN0(\Data_Mem/n8475 ), .IN1(\Data_Mem/n8474 ), .SEL(
        N28), .F(\Data_Mem/n8476 ) );
  MUX \Data_Mem/U8519  ( .IN0(o[907]), .IN1(o[939]), .SEL(N29), .F(
        \Data_Mem/n8475 ) );
  MUX \Data_Mem/U8518  ( .IN0(o[971]), .IN1(o[1003]), .SEL(N29), .F(
        \Data_Mem/n8474 ) );
  MUX \Data_Mem/U8517  ( .IN0(\Data_Mem/n8472 ), .IN1(\Data_Mem/n8457 ), .SEL(
        N25), .F(\Data_Mem/n8473 ) );
  MUX \Data_Mem/U8516  ( .IN0(\Data_Mem/n8471 ), .IN1(\Data_Mem/n8464 ), .SEL(
        N26), .F(\Data_Mem/n8472 ) );
  MUX \Data_Mem/U8515  ( .IN0(\Data_Mem/n8470 ), .IN1(\Data_Mem/n8467 ), .SEL(
        N27), .F(\Data_Mem/n8471 ) );
  MUX \Data_Mem/U8514  ( .IN0(\Data_Mem/n8469 ), .IN1(\Data_Mem/n8468 ), .SEL(
        N28), .F(\Data_Mem/n8470 ) );
  MUX \Data_Mem/U8513  ( .IN0(o[1035]), .IN1(o[1067]), .SEL(N29), .F(
        \Data_Mem/n8469 ) );
  MUX \Data_Mem/U8512  ( .IN0(o[1099]), .IN1(o[1131]), .SEL(N29), .F(
        \Data_Mem/n8468 ) );
  MUX \Data_Mem/U8511  ( .IN0(\Data_Mem/n8466 ), .IN1(\Data_Mem/n8465 ), .SEL(
        N28), .F(\Data_Mem/n8467 ) );
  MUX \Data_Mem/U8510  ( .IN0(o[1163]), .IN1(o[1195]), .SEL(N29), .F(
        \Data_Mem/n8466 ) );
  MUX \Data_Mem/U8509  ( .IN0(o[1227]), .IN1(o[1259]), .SEL(N29), .F(
        \Data_Mem/n8465 ) );
  MUX \Data_Mem/U8508  ( .IN0(\Data_Mem/n8463 ), .IN1(\Data_Mem/n8460 ), .SEL(
        N27), .F(\Data_Mem/n8464 ) );
  MUX \Data_Mem/U8507  ( .IN0(\Data_Mem/n8462 ), .IN1(\Data_Mem/n8461 ), .SEL(
        N28), .F(\Data_Mem/n8463 ) );
  MUX \Data_Mem/U8506  ( .IN0(o[1291]), .IN1(o[1323]), .SEL(N29), .F(
        \Data_Mem/n8462 ) );
  MUX \Data_Mem/U8505  ( .IN0(o[1355]), .IN1(o[1387]), .SEL(N29), .F(
        \Data_Mem/n8461 ) );
  MUX \Data_Mem/U8504  ( .IN0(\Data_Mem/n8459 ), .IN1(\Data_Mem/n8458 ), .SEL(
        N28), .F(\Data_Mem/n8460 ) );
  MUX \Data_Mem/U8503  ( .IN0(o[1419]), .IN1(o[1451]), .SEL(N29), .F(
        \Data_Mem/n8459 ) );
  MUX \Data_Mem/U8502  ( .IN0(o[1483]), .IN1(o[1515]), .SEL(N29), .F(
        \Data_Mem/n8458 ) );
  MUX \Data_Mem/U8501  ( .IN0(\Data_Mem/n8456 ), .IN1(\Data_Mem/n8449 ), .SEL(
        N26), .F(\Data_Mem/n8457 ) );
  MUX \Data_Mem/U8500  ( .IN0(\Data_Mem/n8455 ), .IN1(\Data_Mem/n8452 ), .SEL(
        N27), .F(\Data_Mem/n8456 ) );
  MUX \Data_Mem/U8499  ( .IN0(\Data_Mem/n8454 ), .IN1(\Data_Mem/n8453 ), .SEL(
        N28), .F(\Data_Mem/n8455 ) );
  MUX \Data_Mem/U8498  ( .IN0(o[1547]), .IN1(o[1579]), .SEL(N29), .F(
        \Data_Mem/n8454 ) );
  MUX \Data_Mem/U8497  ( .IN0(o[1611]), .IN1(o[1643]), .SEL(N29), .F(
        \Data_Mem/n8453 ) );
  MUX \Data_Mem/U8496  ( .IN0(\Data_Mem/n8451 ), .IN1(\Data_Mem/n8450 ), .SEL(
        N28), .F(\Data_Mem/n8452 ) );
  MUX \Data_Mem/U8495  ( .IN0(o[1675]), .IN1(o[1707]), .SEL(N29), .F(
        \Data_Mem/n8451 ) );
  MUX \Data_Mem/U8494  ( .IN0(o[1739]), .IN1(o[1771]), .SEL(N29), .F(
        \Data_Mem/n8450 ) );
  MUX \Data_Mem/U8493  ( .IN0(\Data_Mem/n8448 ), .IN1(\Data_Mem/n8445 ), .SEL(
        N27), .F(\Data_Mem/n8449 ) );
  MUX \Data_Mem/U8492  ( .IN0(\Data_Mem/n8447 ), .IN1(\Data_Mem/n8446 ), .SEL(
        N28), .F(\Data_Mem/n8448 ) );
  MUX \Data_Mem/U8491  ( .IN0(o[1803]), .IN1(o[1835]), .SEL(N29), .F(
        \Data_Mem/n8447 ) );
  MUX \Data_Mem/U8490  ( .IN0(o[1867]), .IN1(o[1899]), .SEL(N29), .F(
        \Data_Mem/n8446 ) );
  MUX \Data_Mem/U8489  ( .IN0(\Data_Mem/n8444 ), .IN1(\Data_Mem/n8443 ), .SEL(
        N28), .F(\Data_Mem/n8445 ) );
  MUX \Data_Mem/U8488  ( .IN0(o[1931]), .IN1(o[1963]), .SEL(N29), .F(
        \Data_Mem/n8444 ) );
  MUX \Data_Mem/U8487  ( .IN0(o[1995]), .IN1(o[2027]), .SEL(N29), .F(
        \Data_Mem/n8443 ) );
  MUX \Data_Mem/U8486  ( .IN0(\Data_Mem/n8442 ), .IN1(\Data_Mem/n8411 ), .SEL(
        N24), .F(\Data_Mem/N735 ) );
  MUX \Data_Mem/U8485  ( .IN0(\Data_Mem/n8441 ), .IN1(\Data_Mem/n8426 ), .SEL(
        N25), .F(\Data_Mem/n8442 ) );
  MUX \Data_Mem/U8484  ( .IN0(\Data_Mem/n8440 ), .IN1(\Data_Mem/n8433 ), .SEL(
        N26), .F(\Data_Mem/n8441 ) );
  MUX \Data_Mem/U8483  ( .IN0(\Data_Mem/n8439 ), .IN1(\Data_Mem/n8436 ), .SEL(
        N27), .F(\Data_Mem/n8440 ) );
  MUX \Data_Mem/U8482  ( .IN0(\Data_Mem/n8438 ), .IN1(\Data_Mem/n8437 ), .SEL(
        N28), .F(\Data_Mem/n8439 ) );
  MUX \Data_Mem/U8481  ( .IN0(o[10]), .IN1(o[42]), .SEL(N29), .F(
        \Data_Mem/n8438 ) );
  MUX \Data_Mem/U8480  ( .IN0(o[74]), .IN1(o[106]), .SEL(N29), .F(
        \Data_Mem/n8437 ) );
  MUX \Data_Mem/U8479  ( .IN0(\Data_Mem/n8435 ), .IN1(\Data_Mem/n8434 ), .SEL(
        N28), .F(\Data_Mem/n8436 ) );
  MUX \Data_Mem/U8478  ( .IN0(o[138]), .IN1(o[170]), .SEL(N29), .F(
        \Data_Mem/n8435 ) );
  MUX \Data_Mem/U8477  ( .IN0(o[202]), .IN1(o[234]), .SEL(N29), .F(
        \Data_Mem/n8434 ) );
  MUX \Data_Mem/U8476  ( .IN0(\Data_Mem/n8432 ), .IN1(\Data_Mem/n8429 ), .SEL(
        N27), .F(\Data_Mem/n8433 ) );
  MUX \Data_Mem/U8475  ( .IN0(\Data_Mem/n8431 ), .IN1(\Data_Mem/n8430 ), .SEL(
        N28), .F(\Data_Mem/n8432 ) );
  MUX \Data_Mem/U8474  ( .IN0(o[266]), .IN1(o[298]), .SEL(N29), .F(
        \Data_Mem/n8431 ) );
  MUX \Data_Mem/U8473  ( .IN0(o[330]), .IN1(o[362]), .SEL(N29), .F(
        \Data_Mem/n8430 ) );
  MUX \Data_Mem/U8472  ( .IN0(\Data_Mem/n8428 ), .IN1(\Data_Mem/n8427 ), .SEL(
        N28), .F(\Data_Mem/n8429 ) );
  MUX \Data_Mem/U8471  ( .IN0(o[394]), .IN1(o[426]), .SEL(N29), .F(
        \Data_Mem/n8428 ) );
  MUX \Data_Mem/U8470  ( .IN0(o[458]), .IN1(o[490]), .SEL(N29), .F(
        \Data_Mem/n8427 ) );
  MUX \Data_Mem/U8469  ( .IN0(\Data_Mem/n8425 ), .IN1(\Data_Mem/n8418 ), .SEL(
        N26), .F(\Data_Mem/n8426 ) );
  MUX \Data_Mem/U8468  ( .IN0(\Data_Mem/n8424 ), .IN1(\Data_Mem/n8421 ), .SEL(
        N27), .F(\Data_Mem/n8425 ) );
  MUX \Data_Mem/U8467  ( .IN0(\Data_Mem/n8423 ), .IN1(\Data_Mem/n8422 ), .SEL(
        N28), .F(\Data_Mem/n8424 ) );
  MUX \Data_Mem/U8466  ( .IN0(o[522]), .IN1(o[554]), .SEL(N29), .F(
        \Data_Mem/n8423 ) );
  MUX \Data_Mem/U8465  ( .IN0(o[586]), .IN1(o[618]), .SEL(N29), .F(
        \Data_Mem/n8422 ) );
  MUX \Data_Mem/U8464  ( .IN0(\Data_Mem/n8420 ), .IN1(\Data_Mem/n8419 ), .SEL(
        N28), .F(\Data_Mem/n8421 ) );
  MUX \Data_Mem/U8463  ( .IN0(o[650]), .IN1(o[682]), .SEL(N29), .F(
        \Data_Mem/n8420 ) );
  MUX \Data_Mem/U8462  ( .IN0(o[714]), .IN1(o[746]), .SEL(N29), .F(
        \Data_Mem/n8419 ) );
  MUX \Data_Mem/U8461  ( .IN0(\Data_Mem/n8417 ), .IN1(\Data_Mem/n8414 ), .SEL(
        N27), .F(\Data_Mem/n8418 ) );
  MUX \Data_Mem/U8460  ( .IN0(\Data_Mem/n8416 ), .IN1(\Data_Mem/n8415 ), .SEL(
        N28), .F(\Data_Mem/n8417 ) );
  MUX \Data_Mem/U8459  ( .IN0(o[778]), .IN1(o[810]), .SEL(N29), .F(
        \Data_Mem/n8416 ) );
  MUX \Data_Mem/U8458  ( .IN0(o[842]), .IN1(o[874]), .SEL(N29), .F(
        \Data_Mem/n8415 ) );
  MUX \Data_Mem/U8457  ( .IN0(\Data_Mem/n8413 ), .IN1(\Data_Mem/n8412 ), .SEL(
        N28), .F(\Data_Mem/n8414 ) );
  MUX \Data_Mem/U8456  ( .IN0(o[906]), .IN1(o[938]), .SEL(N29), .F(
        \Data_Mem/n8413 ) );
  MUX \Data_Mem/U8455  ( .IN0(o[970]), .IN1(o[1002]), .SEL(N29), .F(
        \Data_Mem/n8412 ) );
  MUX \Data_Mem/U8454  ( .IN0(\Data_Mem/n8410 ), .IN1(\Data_Mem/n8395 ), .SEL(
        N25), .F(\Data_Mem/n8411 ) );
  MUX \Data_Mem/U8453  ( .IN0(\Data_Mem/n8409 ), .IN1(\Data_Mem/n8402 ), .SEL(
        N26), .F(\Data_Mem/n8410 ) );
  MUX \Data_Mem/U8452  ( .IN0(\Data_Mem/n8408 ), .IN1(\Data_Mem/n8405 ), .SEL(
        N27), .F(\Data_Mem/n8409 ) );
  MUX \Data_Mem/U8451  ( .IN0(\Data_Mem/n8407 ), .IN1(\Data_Mem/n8406 ), .SEL(
        N28), .F(\Data_Mem/n8408 ) );
  MUX \Data_Mem/U8450  ( .IN0(o[1034]), .IN1(o[1066]), .SEL(N29), .F(
        \Data_Mem/n8407 ) );
  MUX \Data_Mem/U8449  ( .IN0(o[1098]), .IN1(o[1130]), .SEL(N29), .F(
        \Data_Mem/n8406 ) );
  MUX \Data_Mem/U8448  ( .IN0(\Data_Mem/n8404 ), .IN1(\Data_Mem/n8403 ), .SEL(
        N28), .F(\Data_Mem/n8405 ) );
  MUX \Data_Mem/U8447  ( .IN0(o[1162]), .IN1(o[1194]), .SEL(N29), .F(
        \Data_Mem/n8404 ) );
  MUX \Data_Mem/U8446  ( .IN0(o[1226]), .IN1(o[1258]), .SEL(N29), .F(
        \Data_Mem/n8403 ) );
  MUX \Data_Mem/U8445  ( .IN0(\Data_Mem/n8401 ), .IN1(\Data_Mem/n8398 ), .SEL(
        N27), .F(\Data_Mem/n8402 ) );
  MUX \Data_Mem/U8444  ( .IN0(\Data_Mem/n8400 ), .IN1(\Data_Mem/n8399 ), .SEL(
        N28), .F(\Data_Mem/n8401 ) );
  MUX \Data_Mem/U8443  ( .IN0(o[1290]), .IN1(o[1322]), .SEL(N29), .F(
        \Data_Mem/n8400 ) );
  MUX \Data_Mem/U8442  ( .IN0(o[1354]), .IN1(o[1386]), .SEL(N29), .F(
        \Data_Mem/n8399 ) );
  MUX \Data_Mem/U8441  ( .IN0(\Data_Mem/n8397 ), .IN1(\Data_Mem/n8396 ), .SEL(
        N28), .F(\Data_Mem/n8398 ) );
  MUX \Data_Mem/U8440  ( .IN0(o[1418]), .IN1(o[1450]), .SEL(N29), .F(
        \Data_Mem/n8397 ) );
  MUX \Data_Mem/U8439  ( .IN0(o[1482]), .IN1(o[1514]), .SEL(N29), .F(
        \Data_Mem/n8396 ) );
  MUX \Data_Mem/U8438  ( .IN0(\Data_Mem/n8394 ), .IN1(\Data_Mem/n8387 ), .SEL(
        N26), .F(\Data_Mem/n8395 ) );
  MUX \Data_Mem/U8437  ( .IN0(\Data_Mem/n8393 ), .IN1(\Data_Mem/n8390 ), .SEL(
        N27), .F(\Data_Mem/n8394 ) );
  MUX \Data_Mem/U8436  ( .IN0(\Data_Mem/n8392 ), .IN1(\Data_Mem/n8391 ), .SEL(
        N28), .F(\Data_Mem/n8393 ) );
  MUX \Data_Mem/U8435  ( .IN0(o[1546]), .IN1(o[1578]), .SEL(N29), .F(
        \Data_Mem/n8392 ) );
  MUX \Data_Mem/U8434  ( .IN0(o[1610]), .IN1(o[1642]), .SEL(N29), .F(
        \Data_Mem/n8391 ) );
  MUX \Data_Mem/U8433  ( .IN0(\Data_Mem/n8389 ), .IN1(\Data_Mem/n8388 ), .SEL(
        N28), .F(\Data_Mem/n8390 ) );
  MUX \Data_Mem/U8432  ( .IN0(o[1674]), .IN1(o[1706]), .SEL(N29), .F(
        \Data_Mem/n8389 ) );
  MUX \Data_Mem/U8431  ( .IN0(o[1738]), .IN1(o[1770]), .SEL(N29), .F(
        \Data_Mem/n8388 ) );
  MUX \Data_Mem/U8430  ( .IN0(\Data_Mem/n8386 ), .IN1(\Data_Mem/n8383 ), .SEL(
        N27), .F(\Data_Mem/n8387 ) );
  MUX \Data_Mem/U8429  ( .IN0(\Data_Mem/n8385 ), .IN1(\Data_Mem/n8384 ), .SEL(
        N28), .F(\Data_Mem/n8386 ) );
  MUX \Data_Mem/U8428  ( .IN0(o[1802]), .IN1(o[1834]), .SEL(N29), .F(
        \Data_Mem/n8385 ) );
  MUX \Data_Mem/U8427  ( .IN0(o[1866]), .IN1(o[1898]), .SEL(N29), .F(
        \Data_Mem/n8384 ) );
  MUX \Data_Mem/U8426  ( .IN0(\Data_Mem/n8382 ), .IN1(\Data_Mem/n8381 ), .SEL(
        N28), .F(\Data_Mem/n8383 ) );
  MUX \Data_Mem/U8425  ( .IN0(o[1930]), .IN1(o[1962]), .SEL(N29), .F(
        \Data_Mem/n8382 ) );
  MUX \Data_Mem/U8424  ( .IN0(o[1994]), .IN1(o[2026]), .SEL(N29), .F(
        \Data_Mem/n8381 ) );
  MUX \Data_Mem/U8423  ( .IN0(\Data_Mem/n8380 ), .IN1(\Data_Mem/n8349 ), .SEL(
        N24), .F(\Data_Mem/N736 ) );
  MUX \Data_Mem/U8422  ( .IN0(\Data_Mem/n8379 ), .IN1(\Data_Mem/n8364 ), .SEL(
        N25), .F(\Data_Mem/n8380 ) );
  MUX \Data_Mem/U8421  ( .IN0(\Data_Mem/n8378 ), .IN1(\Data_Mem/n8371 ), .SEL(
        N26), .F(\Data_Mem/n8379 ) );
  MUX \Data_Mem/U8420  ( .IN0(\Data_Mem/n8377 ), .IN1(\Data_Mem/n8374 ), .SEL(
        N27), .F(\Data_Mem/n8378 ) );
  MUX \Data_Mem/U8419  ( .IN0(\Data_Mem/n8376 ), .IN1(\Data_Mem/n8375 ), .SEL(
        N28), .F(\Data_Mem/n8377 ) );
  MUX \Data_Mem/U8418  ( .IN0(o[9]), .IN1(o[41]), .SEL(N29), .F(
        \Data_Mem/n8376 ) );
  MUX \Data_Mem/U8417  ( .IN0(o[73]), .IN1(o[105]), .SEL(N29), .F(
        \Data_Mem/n8375 ) );
  MUX \Data_Mem/U8416  ( .IN0(\Data_Mem/n8373 ), .IN1(\Data_Mem/n8372 ), .SEL(
        N28), .F(\Data_Mem/n8374 ) );
  MUX \Data_Mem/U8415  ( .IN0(o[137]), .IN1(o[169]), .SEL(N29), .F(
        \Data_Mem/n8373 ) );
  MUX \Data_Mem/U8414  ( .IN0(o[201]), .IN1(o[233]), .SEL(N29), .F(
        \Data_Mem/n8372 ) );
  MUX \Data_Mem/U8413  ( .IN0(\Data_Mem/n8370 ), .IN1(\Data_Mem/n8367 ), .SEL(
        N27), .F(\Data_Mem/n8371 ) );
  MUX \Data_Mem/U8412  ( .IN0(\Data_Mem/n8369 ), .IN1(\Data_Mem/n8368 ), .SEL(
        N28), .F(\Data_Mem/n8370 ) );
  MUX \Data_Mem/U8411  ( .IN0(o[265]), .IN1(o[297]), .SEL(N29), .F(
        \Data_Mem/n8369 ) );
  MUX \Data_Mem/U8410  ( .IN0(o[329]), .IN1(o[361]), .SEL(N29), .F(
        \Data_Mem/n8368 ) );
  MUX \Data_Mem/U8409  ( .IN0(\Data_Mem/n8366 ), .IN1(\Data_Mem/n8365 ), .SEL(
        N28), .F(\Data_Mem/n8367 ) );
  MUX \Data_Mem/U8408  ( .IN0(o[393]), .IN1(o[425]), .SEL(N29), .F(
        \Data_Mem/n8366 ) );
  MUX \Data_Mem/U8407  ( .IN0(o[457]), .IN1(o[489]), .SEL(N29), .F(
        \Data_Mem/n8365 ) );
  MUX \Data_Mem/U8406  ( .IN0(\Data_Mem/n8363 ), .IN1(\Data_Mem/n8356 ), .SEL(
        N26), .F(\Data_Mem/n8364 ) );
  MUX \Data_Mem/U8405  ( .IN0(\Data_Mem/n8362 ), .IN1(\Data_Mem/n8359 ), .SEL(
        N27), .F(\Data_Mem/n8363 ) );
  MUX \Data_Mem/U8404  ( .IN0(\Data_Mem/n8361 ), .IN1(\Data_Mem/n8360 ), .SEL(
        N28), .F(\Data_Mem/n8362 ) );
  MUX \Data_Mem/U8403  ( .IN0(o[521]), .IN1(o[553]), .SEL(N29), .F(
        \Data_Mem/n8361 ) );
  MUX \Data_Mem/U8402  ( .IN0(o[585]), .IN1(o[617]), .SEL(N29), .F(
        \Data_Mem/n8360 ) );
  MUX \Data_Mem/U8401  ( .IN0(\Data_Mem/n8358 ), .IN1(\Data_Mem/n8357 ), .SEL(
        N28), .F(\Data_Mem/n8359 ) );
  MUX \Data_Mem/U8400  ( .IN0(o[649]), .IN1(o[681]), .SEL(N29), .F(
        \Data_Mem/n8358 ) );
  MUX \Data_Mem/U8399  ( .IN0(o[713]), .IN1(o[745]), .SEL(N29), .F(
        \Data_Mem/n8357 ) );
  MUX \Data_Mem/U8398  ( .IN0(\Data_Mem/n8355 ), .IN1(\Data_Mem/n8352 ), .SEL(
        N27), .F(\Data_Mem/n8356 ) );
  MUX \Data_Mem/U8397  ( .IN0(\Data_Mem/n8354 ), .IN1(\Data_Mem/n8353 ), .SEL(
        N28), .F(\Data_Mem/n8355 ) );
  MUX \Data_Mem/U8396  ( .IN0(o[777]), .IN1(o[809]), .SEL(N29), .F(
        \Data_Mem/n8354 ) );
  MUX \Data_Mem/U8395  ( .IN0(o[841]), .IN1(o[873]), .SEL(N29), .F(
        \Data_Mem/n8353 ) );
  MUX \Data_Mem/U8394  ( .IN0(\Data_Mem/n8351 ), .IN1(\Data_Mem/n8350 ), .SEL(
        N28), .F(\Data_Mem/n8352 ) );
  MUX \Data_Mem/U8393  ( .IN0(o[905]), .IN1(o[937]), .SEL(N29), .F(
        \Data_Mem/n8351 ) );
  MUX \Data_Mem/U8392  ( .IN0(o[969]), .IN1(o[1001]), .SEL(N29), .F(
        \Data_Mem/n8350 ) );
  MUX \Data_Mem/U8391  ( .IN0(\Data_Mem/n8348 ), .IN1(\Data_Mem/n8333 ), .SEL(
        N25), .F(\Data_Mem/n8349 ) );
  MUX \Data_Mem/U8390  ( .IN0(\Data_Mem/n8347 ), .IN1(\Data_Mem/n8340 ), .SEL(
        N26), .F(\Data_Mem/n8348 ) );
  MUX \Data_Mem/U8389  ( .IN0(\Data_Mem/n8346 ), .IN1(\Data_Mem/n8343 ), .SEL(
        N27), .F(\Data_Mem/n8347 ) );
  MUX \Data_Mem/U8388  ( .IN0(\Data_Mem/n8345 ), .IN1(\Data_Mem/n8344 ), .SEL(
        N28), .F(\Data_Mem/n8346 ) );
  MUX \Data_Mem/U8387  ( .IN0(o[1033]), .IN1(o[1065]), .SEL(N29), .F(
        \Data_Mem/n8345 ) );
  MUX \Data_Mem/U8386  ( .IN0(o[1097]), .IN1(o[1129]), .SEL(N29), .F(
        \Data_Mem/n8344 ) );
  MUX \Data_Mem/U8385  ( .IN0(\Data_Mem/n8342 ), .IN1(\Data_Mem/n8341 ), .SEL(
        N28), .F(\Data_Mem/n8343 ) );
  MUX \Data_Mem/U8384  ( .IN0(o[1161]), .IN1(o[1193]), .SEL(N29), .F(
        \Data_Mem/n8342 ) );
  MUX \Data_Mem/U8383  ( .IN0(o[1225]), .IN1(o[1257]), .SEL(N29), .F(
        \Data_Mem/n8341 ) );
  MUX \Data_Mem/U8382  ( .IN0(\Data_Mem/n8339 ), .IN1(\Data_Mem/n8336 ), .SEL(
        N27), .F(\Data_Mem/n8340 ) );
  MUX \Data_Mem/U8381  ( .IN0(\Data_Mem/n8338 ), .IN1(\Data_Mem/n8337 ), .SEL(
        N28), .F(\Data_Mem/n8339 ) );
  MUX \Data_Mem/U8380  ( .IN0(o[1289]), .IN1(o[1321]), .SEL(N29), .F(
        \Data_Mem/n8338 ) );
  MUX \Data_Mem/U8379  ( .IN0(o[1353]), .IN1(o[1385]), .SEL(N29), .F(
        \Data_Mem/n8337 ) );
  MUX \Data_Mem/U8378  ( .IN0(\Data_Mem/n8335 ), .IN1(\Data_Mem/n8334 ), .SEL(
        N28), .F(\Data_Mem/n8336 ) );
  MUX \Data_Mem/U8377  ( .IN0(o[1417]), .IN1(o[1449]), .SEL(N29), .F(
        \Data_Mem/n8335 ) );
  MUX \Data_Mem/U8376  ( .IN0(o[1481]), .IN1(o[1513]), .SEL(N29), .F(
        \Data_Mem/n8334 ) );
  MUX \Data_Mem/U8375  ( .IN0(\Data_Mem/n8332 ), .IN1(\Data_Mem/n8325 ), .SEL(
        N26), .F(\Data_Mem/n8333 ) );
  MUX \Data_Mem/U8374  ( .IN0(\Data_Mem/n8331 ), .IN1(\Data_Mem/n8328 ), .SEL(
        N27), .F(\Data_Mem/n8332 ) );
  MUX \Data_Mem/U8373  ( .IN0(\Data_Mem/n8330 ), .IN1(\Data_Mem/n8329 ), .SEL(
        N28), .F(\Data_Mem/n8331 ) );
  MUX \Data_Mem/U8372  ( .IN0(o[1545]), .IN1(o[1577]), .SEL(N29), .F(
        \Data_Mem/n8330 ) );
  MUX \Data_Mem/U8371  ( .IN0(o[1609]), .IN1(o[1641]), .SEL(N29), .F(
        \Data_Mem/n8329 ) );
  MUX \Data_Mem/U8370  ( .IN0(\Data_Mem/n8327 ), .IN1(\Data_Mem/n8326 ), .SEL(
        N28), .F(\Data_Mem/n8328 ) );
  MUX \Data_Mem/U8369  ( .IN0(o[1673]), .IN1(o[1705]), .SEL(N29), .F(
        \Data_Mem/n8327 ) );
  MUX \Data_Mem/U8368  ( .IN0(o[1737]), .IN1(o[1769]), .SEL(N29), .F(
        \Data_Mem/n8326 ) );
  MUX \Data_Mem/U8367  ( .IN0(\Data_Mem/n8324 ), .IN1(\Data_Mem/n8321 ), .SEL(
        N27), .F(\Data_Mem/n8325 ) );
  MUX \Data_Mem/U8366  ( .IN0(\Data_Mem/n8323 ), .IN1(\Data_Mem/n8322 ), .SEL(
        N28), .F(\Data_Mem/n8324 ) );
  MUX \Data_Mem/U8365  ( .IN0(o[1801]), .IN1(o[1833]), .SEL(N29), .F(
        \Data_Mem/n8323 ) );
  MUX \Data_Mem/U8364  ( .IN0(o[1865]), .IN1(o[1897]), .SEL(N29), .F(
        \Data_Mem/n8322 ) );
  MUX \Data_Mem/U8363  ( .IN0(\Data_Mem/n8320 ), .IN1(\Data_Mem/n8319 ), .SEL(
        N28), .F(\Data_Mem/n8321 ) );
  MUX \Data_Mem/U8362  ( .IN0(o[1929]), .IN1(o[1961]), .SEL(N29), .F(
        \Data_Mem/n8320 ) );
  MUX \Data_Mem/U8361  ( .IN0(o[1993]), .IN1(o[2025]), .SEL(N29), .F(
        \Data_Mem/n8319 ) );
  MUX \Data_Mem/U8360  ( .IN0(\Data_Mem/n8318 ), .IN1(\Data_Mem/n8287 ), .SEL(
        N24), .F(\Data_Mem/N737 ) );
  MUX \Data_Mem/U8359  ( .IN0(\Data_Mem/n8317 ), .IN1(\Data_Mem/n8302 ), .SEL(
        N25), .F(\Data_Mem/n8318 ) );
  MUX \Data_Mem/U8358  ( .IN0(\Data_Mem/n8316 ), .IN1(\Data_Mem/n8309 ), .SEL(
        N26), .F(\Data_Mem/n8317 ) );
  MUX \Data_Mem/U8357  ( .IN0(\Data_Mem/n8315 ), .IN1(\Data_Mem/n8312 ), .SEL(
        N27), .F(\Data_Mem/n8316 ) );
  MUX \Data_Mem/U8356  ( .IN0(\Data_Mem/n8314 ), .IN1(\Data_Mem/n8313 ), .SEL(
        N28), .F(\Data_Mem/n8315 ) );
  MUX \Data_Mem/U8355  ( .IN0(o[8]), .IN1(o[40]), .SEL(N29), .F(
        \Data_Mem/n8314 ) );
  MUX \Data_Mem/U8354  ( .IN0(o[72]), .IN1(o[104]), .SEL(N29), .F(
        \Data_Mem/n8313 ) );
  MUX \Data_Mem/U8353  ( .IN0(\Data_Mem/n8311 ), .IN1(\Data_Mem/n8310 ), .SEL(
        N28), .F(\Data_Mem/n8312 ) );
  MUX \Data_Mem/U8352  ( .IN0(o[136]), .IN1(o[168]), .SEL(N29), .F(
        \Data_Mem/n8311 ) );
  MUX \Data_Mem/U8351  ( .IN0(o[200]), .IN1(o[232]), .SEL(N29), .F(
        \Data_Mem/n8310 ) );
  MUX \Data_Mem/U8350  ( .IN0(\Data_Mem/n8308 ), .IN1(\Data_Mem/n8305 ), .SEL(
        N27), .F(\Data_Mem/n8309 ) );
  MUX \Data_Mem/U8349  ( .IN0(\Data_Mem/n8307 ), .IN1(\Data_Mem/n8306 ), .SEL(
        N28), .F(\Data_Mem/n8308 ) );
  MUX \Data_Mem/U8348  ( .IN0(o[264]), .IN1(o[296]), .SEL(N29), .F(
        \Data_Mem/n8307 ) );
  MUX \Data_Mem/U8347  ( .IN0(o[328]), .IN1(o[360]), .SEL(N29), .F(
        \Data_Mem/n8306 ) );
  MUX \Data_Mem/U8346  ( .IN0(\Data_Mem/n8304 ), .IN1(\Data_Mem/n8303 ), .SEL(
        N28), .F(\Data_Mem/n8305 ) );
  MUX \Data_Mem/U8345  ( .IN0(o[392]), .IN1(o[424]), .SEL(N29), .F(
        \Data_Mem/n8304 ) );
  MUX \Data_Mem/U8344  ( .IN0(o[456]), .IN1(o[488]), .SEL(N29), .F(
        \Data_Mem/n8303 ) );
  MUX \Data_Mem/U8343  ( .IN0(\Data_Mem/n8301 ), .IN1(\Data_Mem/n8294 ), .SEL(
        N26), .F(\Data_Mem/n8302 ) );
  MUX \Data_Mem/U8342  ( .IN0(\Data_Mem/n8300 ), .IN1(\Data_Mem/n8297 ), .SEL(
        N27), .F(\Data_Mem/n8301 ) );
  MUX \Data_Mem/U8341  ( .IN0(\Data_Mem/n8299 ), .IN1(\Data_Mem/n8298 ), .SEL(
        N28), .F(\Data_Mem/n8300 ) );
  MUX \Data_Mem/U8340  ( .IN0(o[520]), .IN1(o[552]), .SEL(N29), .F(
        \Data_Mem/n8299 ) );
  MUX \Data_Mem/U8339  ( .IN0(o[584]), .IN1(o[616]), .SEL(N29), .F(
        \Data_Mem/n8298 ) );
  MUX \Data_Mem/U8338  ( .IN0(\Data_Mem/n8296 ), .IN1(\Data_Mem/n8295 ), .SEL(
        N28), .F(\Data_Mem/n8297 ) );
  MUX \Data_Mem/U8337  ( .IN0(o[648]), .IN1(o[680]), .SEL(N29), .F(
        \Data_Mem/n8296 ) );
  MUX \Data_Mem/U8336  ( .IN0(o[712]), .IN1(o[744]), .SEL(N29), .F(
        \Data_Mem/n8295 ) );
  MUX \Data_Mem/U8335  ( .IN0(\Data_Mem/n8293 ), .IN1(\Data_Mem/n8290 ), .SEL(
        N27), .F(\Data_Mem/n8294 ) );
  MUX \Data_Mem/U8334  ( .IN0(\Data_Mem/n8292 ), .IN1(\Data_Mem/n8291 ), .SEL(
        N28), .F(\Data_Mem/n8293 ) );
  MUX \Data_Mem/U8333  ( .IN0(o[776]), .IN1(o[808]), .SEL(N29), .F(
        \Data_Mem/n8292 ) );
  MUX \Data_Mem/U8332  ( .IN0(o[840]), .IN1(o[872]), .SEL(N29), .F(
        \Data_Mem/n8291 ) );
  MUX \Data_Mem/U8331  ( .IN0(\Data_Mem/n8289 ), .IN1(\Data_Mem/n8288 ), .SEL(
        N28), .F(\Data_Mem/n8290 ) );
  MUX \Data_Mem/U8330  ( .IN0(o[904]), .IN1(o[936]), .SEL(N29), .F(
        \Data_Mem/n8289 ) );
  MUX \Data_Mem/U8329  ( .IN0(o[968]), .IN1(o[1000]), .SEL(N29), .F(
        \Data_Mem/n8288 ) );
  MUX \Data_Mem/U8328  ( .IN0(\Data_Mem/n8286 ), .IN1(\Data_Mem/n8271 ), .SEL(
        N25), .F(\Data_Mem/n8287 ) );
  MUX \Data_Mem/U8327  ( .IN0(\Data_Mem/n8285 ), .IN1(\Data_Mem/n8278 ), .SEL(
        N26), .F(\Data_Mem/n8286 ) );
  MUX \Data_Mem/U8326  ( .IN0(\Data_Mem/n8284 ), .IN1(\Data_Mem/n8281 ), .SEL(
        N27), .F(\Data_Mem/n8285 ) );
  MUX \Data_Mem/U8325  ( .IN0(\Data_Mem/n8283 ), .IN1(\Data_Mem/n8282 ), .SEL(
        N28), .F(\Data_Mem/n8284 ) );
  MUX \Data_Mem/U8324  ( .IN0(o[1032]), .IN1(o[1064]), .SEL(N29), .F(
        \Data_Mem/n8283 ) );
  MUX \Data_Mem/U8323  ( .IN0(o[1096]), .IN1(o[1128]), .SEL(N29), .F(
        \Data_Mem/n8282 ) );
  MUX \Data_Mem/U8322  ( .IN0(\Data_Mem/n8280 ), .IN1(\Data_Mem/n8279 ), .SEL(
        N28), .F(\Data_Mem/n8281 ) );
  MUX \Data_Mem/U8321  ( .IN0(o[1160]), .IN1(o[1192]), .SEL(N29), .F(
        \Data_Mem/n8280 ) );
  MUX \Data_Mem/U8320  ( .IN0(o[1224]), .IN1(o[1256]), .SEL(N29), .F(
        \Data_Mem/n8279 ) );
  MUX \Data_Mem/U8319  ( .IN0(\Data_Mem/n8277 ), .IN1(\Data_Mem/n8274 ), .SEL(
        N27), .F(\Data_Mem/n8278 ) );
  MUX \Data_Mem/U8318  ( .IN0(\Data_Mem/n8276 ), .IN1(\Data_Mem/n8275 ), .SEL(
        N28), .F(\Data_Mem/n8277 ) );
  MUX \Data_Mem/U8317  ( .IN0(o[1288]), .IN1(o[1320]), .SEL(N29), .F(
        \Data_Mem/n8276 ) );
  MUX \Data_Mem/U8316  ( .IN0(o[1352]), .IN1(o[1384]), .SEL(N29), .F(
        \Data_Mem/n8275 ) );
  MUX \Data_Mem/U8315  ( .IN0(\Data_Mem/n8273 ), .IN1(\Data_Mem/n8272 ), .SEL(
        N28), .F(\Data_Mem/n8274 ) );
  MUX \Data_Mem/U8314  ( .IN0(o[1416]), .IN1(o[1448]), .SEL(N29), .F(
        \Data_Mem/n8273 ) );
  MUX \Data_Mem/U8313  ( .IN0(o[1480]), .IN1(o[1512]), .SEL(N29), .F(
        \Data_Mem/n8272 ) );
  MUX \Data_Mem/U8312  ( .IN0(\Data_Mem/n8270 ), .IN1(\Data_Mem/n8263 ), .SEL(
        N26), .F(\Data_Mem/n8271 ) );
  MUX \Data_Mem/U8311  ( .IN0(\Data_Mem/n8269 ), .IN1(\Data_Mem/n8266 ), .SEL(
        N27), .F(\Data_Mem/n8270 ) );
  MUX \Data_Mem/U8310  ( .IN0(\Data_Mem/n8268 ), .IN1(\Data_Mem/n8267 ), .SEL(
        N28), .F(\Data_Mem/n8269 ) );
  MUX \Data_Mem/U8309  ( .IN0(o[1544]), .IN1(o[1576]), .SEL(N29), .F(
        \Data_Mem/n8268 ) );
  MUX \Data_Mem/U8308  ( .IN0(o[1608]), .IN1(o[1640]), .SEL(N29), .F(
        \Data_Mem/n8267 ) );
  MUX \Data_Mem/U8307  ( .IN0(\Data_Mem/n8265 ), .IN1(\Data_Mem/n8264 ), .SEL(
        N28), .F(\Data_Mem/n8266 ) );
  MUX \Data_Mem/U8306  ( .IN0(o[1672]), .IN1(o[1704]), .SEL(N29), .F(
        \Data_Mem/n8265 ) );
  MUX \Data_Mem/U8305  ( .IN0(o[1736]), .IN1(o[1768]), .SEL(N29), .F(
        \Data_Mem/n8264 ) );
  MUX \Data_Mem/U8304  ( .IN0(\Data_Mem/n8262 ), .IN1(\Data_Mem/n8259 ), .SEL(
        N27), .F(\Data_Mem/n8263 ) );
  MUX \Data_Mem/U8303  ( .IN0(\Data_Mem/n8261 ), .IN1(\Data_Mem/n8260 ), .SEL(
        N28), .F(\Data_Mem/n8262 ) );
  MUX \Data_Mem/U8302  ( .IN0(o[1800]), .IN1(o[1832]), .SEL(N29), .F(
        \Data_Mem/n8261 ) );
  MUX \Data_Mem/U8301  ( .IN0(o[1864]), .IN1(o[1896]), .SEL(N29), .F(
        \Data_Mem/n8260 ) );
  MUX \Data_Mem/U8300  ( .IN0(\Data_Mem/n8258 ), .IN1(\Data_Mem/n8257 ), .SEL(
        N28), .F(\Data_Mem/n8259 ) );
  MUX \Data_Mem/U8299  ( .IN0(o[1928]), .IN1(o[1960]), .SEL(N29), .F(
        \Data_Mem/n8258 ) );
  MUX \Data_Mem/U8298  ( .IN0(o[1992]), .IN1(o[2024]), .SEL(N29), .F(
        \Data_Mem/n8257 ) );
  MUX \Data_Mem/U8297  ( .IN0(\Data_Mem/n8256 ), .IN1(\Data_Mem/n8225 ), .SEL(
        N24), .F(\Data_Mem/N738 ) );
  MUX \Data_Mem/U8296  ( .IN0(\Data_Mem/n8255 ), .IN1(\Data_Mem/n8240 ), .SEL(
        N25), .F(\Data_Mem/n8256 ) );
  MUX \Data_Mem/U8295  ( .IN0(\Data_Mem/n8254 ), .IN1(\Data_Mem/n8247 ), .SEL(
        N26), .F(\Data_Mem/n8255 ) );
  MUX \Data_Mem/U8294  ( .IN0(\Data_Mem/n8253 ), .IN1(\Data_Mem/n8250 ), .SEL(
        N27), .F(\Data_Mem/n8254 ) );
  MUX \Data_Mem/U8293  ( .IN0(\Data_Mem/n8252 ), .IN1(\Data_Mem/n8251 ), .SEL(
        N28), .F(\Data_Mem/n8253 ) );
  MUX \Data_Mem/U8292  ( .IN0(o[7]), .IN1(o[39]), .SEL(N29), .F(
        \Data_Mem/n8252 ) );
  MUX \Data_Mem/U8291  ( .IN0(o[71]), .IN1(o[103]), .SEL(N29), .F(
        \Data_Mem/n8251 ) );
  MUX \Data_Mem/U8290  ( .IN0(\Data_Mem/n8249 ), .IN1(\Data_Mem/n8248 ), .SEL(
        N28), .F(\Data_Mem/n8250 ) );
  MUX \Data_Mem/U8289  ( .IN0(o[135]), .IN1(o[167]), .SEL(N29), .F(
        \Data_Mem/n8249 ) );
  MUX \Data_Mem/U8288  ( .IN0(o[199]), .IN1(o[231]), .SEL(N29), .F(
        \Data_Mem/n8248 ) );
  MUX \Data_Mem/U8287  ( .IN0(\Data_Mem/n8246 ), .IN1(\Data_Mem/n8243 ), .SEL(
        N27), .F(\Data_Mem/n8247 ) );
  MUX \Data_Mem/U8286  ( .IN0(\Data_Mem/n8245 ), .IN1(\Data_Mem/n8244 ), .SEL(
        N28), .F(\Data_Mem/n8246 ) );
  MUX \Data_Mem/U8285  ( .IN0(o[263]), .IN1(o[295]), .SEL(N29), .F(
        \Data_Mem/n8245 ) );
  MUX \Data_Mem/U8284  ( .IN0(o[327]), .IN1(o[359]), .SEL(N29), .F(
        \Data_Mem/n8244 ) );
  MUX \Data_Mem/U8283  ( .IN0(\Data_Mem/n8242 ), .IN1(\Data_Mem/n8241 ), .SEL(
        N28), .F(\Data_Mem/n8243 ) );
  MUX \Data_Mem/U8282  ( .IN0(o[391]), .IN1(o[423]), .SEL(N29), .F(
        \Data_Mem/n8242 ) );
  MUX \Data_Mem/U8281  ( .IN0(o[455]), .IN1(o[487]), .SEL(N29), .F(
        \Data_Mem/n8241 ) );
  MUX \Data_Mem/U8280  ( .IN0(\Data_Mem/n8239 ), .IN1(\Data_Mem/n8232 ), .SEL(
        N26), .F(\Data_Mem/n8240 ) );
  MUX \Data_Mem/U8279  ( .IN0(\Data_Mem/n8238 ), .IN1(\Data_Mem/n8235 ), .SEL(
        N27), .F(\Data_Mem/n8239 ) );
  MUX \Data_Mem/U8278  ( .IN0(\Data_Mem/n8237 ), .IN1(\Data_Mem/n8236 ), .SEL(
        N28), .F(\Data_Mem/n8238 ) );
  MUX \Data_Mem/U8277  ( .IN0(o[519]), .IN1(o[551]), .SEL(N29), .F(
        \Data_Mem/n8237 ) );
  MUX \Data_Mem/U8276  ( .IN0(o[583]), .IN1(o[615]), .SEL(N29), .F(
        \Data_Mem/n8236 ) );
  MUX \Data_Mem/U8275  ( .IN0(\Data_Mem/n8234 ), .IN1(\Data_Mem/n8233 ), .SEL(
        N28), .F(\Data_Mem/n8235 ) );
  MUX \Data_Mem/U8274  ( .IN0(o[647]), .IN1(o[679]), .SEL(N29), .F(
        \Data_Mem/n8234 ) );
  MUX \Data_Mem/U8273  ( .IN0(o[711]), .IN1(o[743]), .SEL(N29), .F(
        \Data_Mem/n8233 ) );
  MUX \Data_Mem/U8272  ( .IN0(\Data_Mem/n8231 ), .IN1(\Data_Mem/n8228 ), .SEL(
        N27), .F(\Data_Mem/n8232 ) );
  MUX \Data_Mem/U8271  ( .IN0(\Data_Mem/n8230 ), .IN1(\Data_Mem/n8229 ), .SEL(
        N28), .F(\Data_Mem/n8231 ) );
  MUX \Data_Mem/U8270  ( .IN0(o[775]), .IN1(o[807]), .SEL(N29), .F(
        \Data_Mem/n8230 ) );
  MUX \Data_Mem/U8269  ( .IN0(o[839]), .IN1(o[871]), .SEL(N29), .F(
        \Data_Mem/n8229 ) );
  MUX \Data_Mem/U8268  ( .IN0(\Data_Mem/n8227 ), .IN1(\Data_Mem/n8226 ), .SEL(
        N28), .F(\Data_Mem/n8228 ) );
  MUX \Data_Mem/U8267  ( .IN0(o[903]), .IN1(o[935]), .SEL(N29), .F(
        \Data_Mem/n8227 ) );
  MUX \Data_Mem/U8266  ( .IN0(o[967]), .IN1(o[999]), .SEL(N29), .F(
        \Data_Mem/n8226 ) );
  MUX \Data_Mem/U8265  ( .IN0(\Data_Mem/n8224 ), .IN1(\Data_Mem/n8209 ), .SEL(
        N25), .F(\Data_Mem/n8225 ) );
  MUX \Data_Mem/U8264  ( .IN0(\Data_Mem/n8223 ), .IN1(\Data_Mem/n8216 ), .SEL(
        N26), .F(\Data_Mem/n8224 ) );
  MUX \Data_Mem/U8263  ( .IN0(\Data_Mem/n8222 ), .IN1(\Data_Mem/n8219 ), .SEL(
        N27), .F(\Data_Mem/n8223 ) );
  MUX \Data_Mem/U8262  ( .IN0(\Data_Mem/n8221 ), .IN1(\Data_Mem/n8220 ), .SEL(
        N28), .F(\Data_Mem/n8222 ) );
  MUX \Data_Mem/U8261  ( .IN0(o[1031]), .IN1(o[1063]), .SEL(N29), .F(
        \Data_Mem/n8221 ) );
  MUX \Data_Mem/U8260  ( .IN0(o[1095]), .IN1(o[1127]), .SEL(N29), .F(
        \Data_Mem/n8220 ) );
  MUX \Data_Mem/U8259  ( .IN0(\Data_Mem/n8218 ), .IN1(\Data_Mem/n8217 ), .SEL(
        N28), .F(\Data_Mem/n8219 ) );
  MUX \Data_Mem/U8258  ( .IN0(o[1159]), .IN1(o[1191]), .SEL(N29), .F(
        \Data_Mem/n8218 ) );
  MUX \Data_Mem/U8257  ( .IN0(o[1223]), .IN1(o[1255]), .SEL(N29), .F(
        \Data_Mem/n8217 ) );
  MUX \Data_Mem/U8256  ( .IN0(\Data_Mem/n8215 ), .IN1(\Data_Mem/n8212 ), .SEL(
        N27), .F(\Data_Mem/n8216 ) );
  MUX \Data_Mem/U8255  ( .IN0(\Data_Mem/n8214 ), .IN1(\Data_Mem/n8213 ), .SEL(
        N28), .F(\Data_Mem/n8215 ) );
  MUX \Data_Mem/U8254  ( .IN0(o[1287]), .IN1(o[1319]), .SEL(N29), .F(
        \Data_Mem/n8214 ) );
  MUX \Data_Mem/U8253  ( .IN0(o[1351]), .IN1(o[1383]), .SEL(N29), .F(
        \Data_Mem/n8213 ) );
  MUX \Data_Mem/U8252  ( .IN0(\Data_Mem/n8211 ), .IN1(\Data_Mem/n8210 ), .SEL(
        N28), .F(\Data_Mem/n8212 ) );
  MUX \Data_Mem/U8251  ( .IN0(o[1415]), .IN1(o[1447]), .SEL(N29), .F(
        \Data_Mem/n8211 ) );
  MUX \Data_Mem/U8250  ( .IN0(o[1479]), .IN1(o[1511]), .SEL(N29), .F(
        \Data_Mem/n8210 ) );
  MUX \Data_Mem/U8249  ( .IN0(\Data_Mem/n8208 ), .IN1(\Data_Mem/n8201 ), .SEL(
        N26), .F(\Data_Mem/n8209 ) );
  MUX \Data_Mem/U8248  ( .IN0(\Data_Mem/n8207 ), .IN1(\Data_Mem/n8204 ), .SEL(
        N27), .F(\Data_Mem/n8208 ) );
  MUX \Data_Mem/U8247  ( .IN0(\Data_Mem/n8206 ), .IN1(\Data_Mem/n8205 ), .SEL(
        N28), .F(\Data_Mem/n8207 ) );
  MUX \Data_Mem/U8246  ( .IN0(o[1543]), .IN1(o[1575]), .SEL(N29), .F(
        \Data_Mem/n8206 ) );
  MUX \Data_Mem/U8245  ( .IN0(o[1607]), .IN1(o[1639]), .SEL(N29), .F(
        \Data_Mem/n8205 ) );
  MUX \Data_Mem/U8244  ( .IN0(\Data_Mem/n8203 ), .IN1(\Data_Mem/n8202 ), .SEL(
        N28), .F(\Data_Mem/n8204 ) );
  MUX \Data_Mem/U8243  ( .IN0(o[1671]), .IN1(o[1703]), .SEL(N29), .F(
        \Data_Mem/n8203 ) );
  MUX \Data_Mem/U8242  ( .IN0(o[1735]), .IN1(o[1767]), .SEL(N29), .F(
        \Data_Mem/n8202 ) );
  MUX \Data_Mem/U8241  ( .IN0(\Data_Mem/n8200 ), .IN1(\Data_Mem/n8197 ), .SEL(
        N27), .F(\Data_Mem/n8201 ) );
  MUX \Data_Mem/U8240  ( .IN0(\Data_Mem/n8199 ), .IN1(\Data_Mem/n8198 ), .SEL(
        N28), .F(\Data_Mem/n8200 ) );
  MUX \Data_Mem/U8239  ( .IN0(o[1799]), .IN1(o[1831]), .SEL(N29), .F(
        \Data_Mem/n8199 ) );
  MUX \Data_Mem/U8238  ( .IN0(o[1863]), .IN1(o[1895]), .SEL(N29), .F(
        \Data_Mem/n8198 ) );
  MUX \Data_Mem/U8237  ( .IN0(\Data_Mem/n8196 ), .IN1(\Data_Mem/n8195 ), .SEL(
        N28), .F(\Data_Mem/n8197 ) );
  MUX \Data_Mem/U8236  ( .IN0(o[1927]), .IN1(o[1959]), .SEL(N29), .F(
        \Data_Mem/n8196 ) );
  MUX \Data_Mem/U8235  ( .IN0(o[1991]), .IN1(o[2023]), .SEL(N29), .F(
        \Data_Mem/n8195 ) );
  MUX \Data_Mem/U8234  ( .IN0(\Data_Mem/n8194 ), .IN1(\Data_Mem/n8163 ), .SEL(
        N24), .F(\Data_Mem/N739 ) );
  MUX \Data_Mem/U8233  ( .IN0(\Data_Mem/n8193 ), .IN1(\Data_Mem/n8178 ), .SEL(
        N25), .F(\Data_Mem/n8194 ) );
  MUX \Data_Mem/U8232  ( .IN0(\Data_Mem/n8192 ), .IN1(\Data_Mem/n8185 ), .SEL(
        N26), .F(\Data_Mem/n8193 ) );
  MUX \Data_Mem/U8231  ( .IN0(\Data_Mem/n8191 ), .IN1(\Data_Mem/n8188 ), .SEL(
        N27), .F(\Data_Mem/n8192 ) );
  MUX \Data_Mem/U8230  ( .IN0(\Data_Mem/n8190 ), .IN1(\Data_Mem/n8189 ), .SEL(
        N28), .F(\Data_Mem/n8191 ) );
  MUX \Data_Mem/U8229  ( .IN0(o[6]), .IN1(o[38]), .SEL(N29), .F(
        \Data_Mem/n8190 ) );
  MUX \Data_Mem/U8228  ( .IN0(o[70]), .IN1(o[102]), .SEL(N29), .F(
        \Data_Mem/n8189 ) );
  MUX \Data_Mem/U8227  ( .IN0(\Data_Mem/n8187 ), .IN1(\Data_Mem/n8186 ), .SEL(
        N28), .F(\Data_Mem/n8188 ) );
  MUX \Data_Mem/U8226  ( .IN0(o[134]), .IN1(o[166]), .SEL(N29), .F(
        \Data_Mem/n8187 ) );
  MUX \Data_Mem/U8225  ( .IN0(o[198]), .IN1(o[230]), .SEL(N29), .F(
        \Data_Mem/n8186 ) );
  MUX \Data_Mem/U8224  ( .IN0(\Data_Mem/n8184 ), .IN1(\Data_Mem/n8181 ), .SEL(
        N27), .F(\Data_Mem/n8185 ) );
  MUX \Data_Mem/U8223  ( .IN0(\Data_Mem/n8183 ), .IN1(\Data_Mem/n8182 ), .SEL(
        N28), .F(\Data_Mem/n8184 ) );
  MUX \Data_Mem/U8222  ( .IN0(o[262]), .IN1(o[294]), .SEL(N29), .F(
        \Data_Mem/n8183 ) );
  MUX \Data_Mem/U8221  ( .IN0(o[326]), .IN1(o[358]), .SEL(N29), .F(
        \Data_Mem/n8182 ) );
  MUX \Data_Mem/U8220  ( .IN0(\Data_Mem/n8180 ), .IN1(\Data_Mem/n8179 ), .SEL(
        N28), .F(\Data_Mem/n8181 ) );
  MUX \Data_Mem/U8219  ( .IN0(o[390]), .IN1(o[422]), .SEL(N29), .F(
        \Data_Mem/n8180 ) );
  MUX \Data_Mem/U8218  ( .IN0(o[454]), .IN1(o[486]), .SEL(N29), .F(
        \Data_Mem/n8179 ) );
  MUX \Data_Mem/U8217  ( .IN0(\Data_Mem/n8177 ), .IN1(\Data_Mem/n8170 ), .SEL(
        N26), .F(\Data_Mem/n8178 ) );
  MUX \Data_Mem/U8216  ( .IN0(\Data_Mem/n8176 ), .IN1(\Data_Mem/n8173 ), .SEL(
        N27), .F(\Data_Mem/n8177 ) );
  MUX \Data_Mem/U8215  ( .IN0(\Data_Mem/n8175 ), .IN1(\Data_Mem/n8174 ), .SEL(
        N28), .F(\Data_Mem/n8176 ) );
  MUX \Data_Mem/U8214  ( .IN0(o[518]), .IN1(o[550]), .SEL(N29), .F(
        \Data_Mem/n8175 ) );
  MUX \Data_Mem/U8213  ( .IN0(o[582]), .IN1(o[614]), .SEL(N29), .F(
        \Data_Mem/n8174 ) );
  MUX \Data_Mem/U8212  ( .IN0(\Data_Mem/n8172 ), .IN1(\Data_Mem/n8171 ), .SEL(
        N28), .F(\Data_Mem/n8173 ) );
  MUX \Data_Mem/U8211  ( .IN0(o[646]), .IN1(o[678]), .SEL(N29), .F(
        \Data_Mem/n8172 ) );
  MUX \Data_Mem/U8210  ( .IN0(o[710]), .IN1(o[742]), .SEL(N29), .F(
        \Data_Mem/n8171 ) );
  MUX \Data_Mem/U8209  ( .IN0(\Data_Mem/n8169 ), .IN1(\Data_Mem/n8166 ), .SEL(
        N27), .F(\Data_Mem/n8170 ) );
  MUX \Data_Mem/U8208  ( .IN0(\Data_Mem/n8168 ), .IN1(\Data_Mem/n8167 ), .SEL(
        N28), .F(\Data_Mem/n8169 ) );
  MUX \Data_Mem/U8207  ( .IN0(o[774]), .IN1(o[806]), .SEL(N29), .F(
        \Data_Mem/n8168 ) );
  MUX \Data_Mem/U8206  ( .IN0(o[838]), .IN1(o[870]), .SEL(N29), .F(
        \Data_Mem/n8167 ) );
  MUX \Data_Mem/U8205  ( .IN0(\Data_Mem/n8165 ), .IN1(\Data_Mem/n8164 ), .SEL(
        N28), .F(\Data_Mem/n8166 ) );
  MUX \Data_Mem/U8204  ( .IN0(o[902]), .IN1(o[934]), .SEL(N29), .F(
        \Data_Mem/n8165 ) );
  MUX \Data_Mem/U8203  ( .IN0(o[966]), .IN1(o[998]), .SEL(N29), .F(
        \Data_Mem/n8164 ) );
  MUX \Data_Mem/U8202  ( .IN0(\Data_Mem/n8162 ), .IN1(\Data_Mem/n8147 ), .SEL(
        N25), .F(\Data_Mem/n8163 ) );
  MUX \Data_Mem/U8201  ( .IN0(\Data_Mem/n8161 ), .IN1(\Data_Mem/n8154 ), .SEL(
        N26), .F(\Data_Mem/n8162 ) );
  MUX \Data_Mem/U8200  ( .IN0(\Data_Mem/n8160 ), .IN1(\Data_Mem/n8157 ), .SEL(
        N27), .F(\Data_Mem/n8161 ) );
  MUX \Data_Mem/U8199  ( .IN0(\Data_Mem/n8159 ), .IN1(\Data_Mem/n8158 ), .SEL(
        N28), .F(\Data_Mem/n8160 ) );
  MUX \Data_Mem/U8198  ( .IN0(o[1030]), .IN1(o[1062]), .SEL(N29), .F(
        \Data_Mem/n8159 ) );
  MUX \Data_Mem/U8197  ( .IN0(o[1094]), .IN1(o[1126]), .SEL(N29), .F(
        \Data_Mem/n8158 ) );
  MUX \Data_Mem/U8196  ( .IN0(\Data_Mem/n8156 ), .IN1(\Data_Mem/n8155 ), .SEL(
        N28), .F(\Data_Mem/n8157 ) );
  MUX \Data_Mem/U8195  ( .IN0(o[1158]), .IN1(o[1190]), .SEL(N29), .F(
        \Data_Mem/n8156 ) );
  MUX \Data_Mem/U8194  ( .IN0(o[1222]), .IN1(o[1254]), .SEL(N29), .F(
        \Data_Mem/n8155 ) );
  MUX \Data_Mem/U8193  ( .IN0(\Data_Mem/n8153 ), .IN1(\Data_Mem/n8150 ), .SEL(
        N27), .F(\Data_Mem/n8154 ) );
  MUX \Data_Mem/U8192  ( .IN0(\Data_Mem/n8152 ), .IN1(\Data_Mem/n8151 ), .SEL(
        N28), .F(\Data_Mem/n8153 ) );
  MUX \Data_Mem/U8191  ( .IN0(o[1286]), .IN1(o[1318]), .SEL(N29), .F(
        \Data_Mem/n8152 ) );
  MUX \Data_Mem/U8190  ( .IN0(o[1350]), .IN1(o[1382]), .SEL(N29), .F(
        \Data_Mem/n8151 ) );
  MUX \Data_Mem/U8189  ( .IN0(\Data_Mem/n8149 ), .IN1(\Data_Mem/n8148 ), .SEL(
        N28), .F(\Data_Mem/n8150 ) );
  MUX \Data_Mem/U8188  ( .IN0(o[1414]), .IN1(o[1446]), .SEL(N29), .F(
        \Data_Mem/n8149 ) );
  MUX \Data_Mem/U8187  ( .IN0(o[1478]), .IN1(o[1510]), .SEL(N29), .F(
        \Data_Mem/n8148 ) );
  MUX \Data_Mem/U8186  ( .IN0(\Data_Mem/n8146 ), .IN1(\Data_Mem/n8139 ), .SEL(
        N26), .F(\Data_Mem/n8147 ) );
  MUX \Data_Mem/U8185  ( .IN0(\Data_Mem/n8145 ), .IN1(\Data_Mem/n8142 ), .SEL(
        N27), .F(\Data_Mem/n8146 ) );
  MUX \Data_Mem/U8184  ( .IN0(\Data_Mem/n8144 ), .IN1(\Data_Mem/n8143 ), .SEL(
        N28), .F(\Data_Mem/n8145 ) );
  MUX \Data_Mem/U8183  ( .IN0(o[1542]), .IN1(o[1574]), .SEL(N29), .F(
        \Data_Mem/n8144 ) );
  MUX \Data_Mem/U8182  ( .IN0(o[1606]), .IN1(o[1638]), .SEL(N29), .F(
        \Data_Mem/n8143 ) );
  MUX \Data_Mem/U8181  ( .IN0(\Data_Mem/n8141 ), .IN1(\Data_Mem/n8140 ), .SEL(
        N28), .F(\Data_Mem/n8142 ) );
  MUX \Data_Mem/U8180  ( .IN0(o[1670]), .IN1(o[1702]), .SEL(N29), .F(
        \Data_Mem/n8141 ) );
  MUX \Data_Mem/U8179  ( .IN0(o[1734]), .IN1(o[1766]), .SEL(N29), .F(
        \Data_Mem/n8140 ) );
  MUX \Data_Mem/U8178  ( .IN0(\Data_Mem/n8138 ), .IN1(\Data_Mem/n8135 ), .SEL(
        N27), .F(\Data_Mem/n8139 ) );
  MUX \Data_Mem/U8177  ( .IN0(\Data_Mem/n8137 ), .IN1(\Data_Mem/n8136 ), .SEL(
        N28), .F(\Data_Mem/n8138 ) );
  MUX \Data_Mem/U8176  ( .IN0(o[1798]), .IN1(o[1830]), .SEL(N29), .F(
        \Data_Mem/n8137 ) );
  MUX \Data_Mem/U8175  ( .IN0(o[1862]), .IN1(o[1894]), .SEL(N29), .F(
        \Data_Mem/n8136 ) );
  MUX \Data_Mem/U8174  ( .IN0(\Data_Mem/n8134 ), .IN1(\Data_Mem/n8133 ), .SEL(
        N28), .F(\Data_Mem/n8135 ) );
  MUX \Data_Mem/U8173  ( .IN0(o[1926]), .IN1(o[1958]), .SEL(N29), .F(
        \Data_Mem/n8134 ) );
  MUX \Data_Mem/U8172  ( .IN0(o[1990]), .IN1(o[2022]), .SEL(N29), .F(
        \Data_Mem/n8133 ) );
  MUX \Data_Mem/U8171  ( .IN0(\Data_Mem/n8132 ), .IN1(\Data_Mem/n8101 ), .SEL(
        N24), .F(\Data_Mem/N740 ) );
  MUX \Data_Mem/U8170  ( .IN0(\Data_Mem/n8131 ), .IN1(\Data_Mem/n8116 ), .SEL(
        N25), .F(\Data_Mem/n8132 ) );
  MUX \Data_Mem/U8169  ( .IN0(\Data_Mem/n8130 ), .IN1(\Data_Mem/n8123 ), .SEL(
        N26), .F(\Data_Mem/n8131 ) );
  MUX \Data_Mem/U8168  ( .IN0(\Data_Mem/n8129 ), .IN1(\Data_Mem/n8126 ), .SEL(
        N27), .F(\Data_Mem/n8130 ) );
  MUX \Data_Mem/U8167  ( .IN0(\Data_Mem/n8128 ), .IN1(\Data_Mem/n8127 ), .SEL(
        N28), .F(\Data_Mem/n8129 ) );
  MUX \Data_Mem/U8166  ( .IN0(o[5]), .IN1(o[37]), .SEL(N29), .F(
        \Data_Mem/n8128 ) );
  MUX \Data_Mem/U8165  ( .IN0(o[69]), .IN1(o[101]), .SEL(N29), .F(
        \Data_Mem/n8127 ) );
  MUX \Data_Mem/U8164  ( .IN0(\Data_Mem/n8125 ), .IN1(\Data_Mem/n8124 ), .SEL(
        N28), .F(\Data_Mem/n8126 ) );
  MUX \Data_Mem/U8163  ( .IN0(o[133]), .IN1(o[165]), .SEL(N29), .F(
        \Data_Mem/n8125 ) );
  MUX \Data_Mem/U8162  ( .IN0(o[197]), .IN1(o[229]), .SEL(N29), .F(
        \Data_Mem/n8124 ) );
  MUX \Data_Mem/U8161  ( .IN0(\Data_Mem/n8122 ), .IN1(\Data_Mem/n8119 ), .SEL(
        N27), .F(\Data_Mem/n8123 ) );
  MUX \Data_Mem/U8160  ( .IN0(\Data_Mem/n8121 ), .IN1(\Data_Mem/n8120 ), .SEL(
        N28), .F(\Data_Mem/n8122 ) );
  MUX \Data_Mem/U8159  ( .IN0(o[261]), .IN1(o[293]), .SEL(N29), .F(
        \Data_Mem/n8121 ) );
  MUX \Data_Mem/U8158  ( .IN0(o[325]), .IN1(o[357]), .SEL(N29), .F(
        \Data_Mem/n8120 ) );
  MUX \Data_Mem/U8157  ( .IN0(\Data_Mem/n8118 ), .IN1(\Data_Mem/n8117 ), .SEL(
        N28), .F(\Data_Mem/n8119 ) );
  MUX \Data_Mem/U8156  ( .IN0(o[389]), .IN1(o[421]), .SEL(N29), .F(
        \Data_Mem/n8118 ) );
  MUX \Data_Mem/U8155  ( .IN0(o[453]), .IN1(o[485]), .SEL(N29), .F(
        \Data_Mem/n8117 ) );
  MUX \Data_Mem/U8154  ( .IN0(\Data_Mem/n8115 ), .IN1(\Data_Mem/n8108 ), .SEL(
        N26), .F(\Data_Mem/n8116 ) );
  MUX \Data_Mem/U8153  ( .IN0(\Data_Mem/n8114 ), .IN1(\Data_Mem/n8111 ), .SEL(
        N27), .F(\Data_Mem/n8115 ) );
  MUX \Data_Mem/U8152  ( .IN0(\Data_Mem/n8113 ), .IN1(\Data_Mem/n8112 ), .SEL(
        N28), .F(\Data_Mem/n8114 ) );
  MUX \Data_Mem/U8151  ( .IN0(o[517]), .IN1(o[549]), .SEL(N29), .F(
        \Data_Mem/n8113 ) );
  MUX \Data_Mem/U8150  ( .IN0(o[581]), .IN1(o[613]), .SEL(N29), .F(
        \Data_Mem/n8112 ) );
  MUX \Data_Mem/U8149  ( .IN0(\Data_Mem/n8110 ), .IN1(\Data_Mem/n8109 ), .SEL(
        N28), .F(\Data_Mem/n8111 ) );
  MUX \Data_Mem/U8148  ( .IN0(o[645]), .IN1(o[677]), .SEL(N29), .F(
        \Data_Mem/n8110 ) );
  MUX \Data_Mem/U8147  ( .IN0(o[709]), .IN1(o[741]), .SEL(N29), .F(
        \Data_Mem/n8109 ) );
  MUX \Data_Mem/U8146  ( .IN0(\Data_Mem/n8107 ), .IN1(\Data_Mem/n8104 ), .SEL(
        N27), .F(\Data_Mem/n8108 ) );
  MUX \Data_Mem/U8145  ( .IN0(\Data_Mem/n8106 ), .IN1(\Data_Mem/n8105 ), .SEL(
        N28), .F(\Data_Mem/n8107 ) );
  MUX \Data_Mem/U8144  ( .IN0(o[773]), .IN1(o[805]), .SEL(N29), .F(
        \Data_Mem/n8106 ) );
  MUX \Data_Mem/U8143  ( .IN0(o[837]), .IN1(o[869]), .SEL(N29), .F(
        \Data_Mem/n8105 ) );
  MUX \Data_Mem/U8142  ( .IN0(\Data_Mem/n8103 ), .IN1(\Data_Mem/n8102 ), .SEL(
        N28), .F(\Data_Mem/n8104 ) );
  MUX \Data_Mem/U8141  ( .IN0(o[901]), .IN1(o[933]), .SEL(N29), .F(
        \Data_Mem/n8103 ) );
  MUX \Data_Mem/U8140  ( .IN0(o[965]), .IN1(o[997]), .SEL(N29), .F(
        \Data_Mem/n8102 ) );
  MUX \Data_Mem/U8139  ( .IN0(\Data_Mem/n8100 ), .IN1(\Data_Mem/n8085 ), .SEL(
        N25), .F(\Data_Mem/n8101 ) );
  MUX \Data_Mem/U8138  ( .IN0(\Data_Mem/n8099 ), .IN1(\Data_Mem/n8092 ), .SEL(
        N26), .F(\Data_Mem/n8100 ) );
  MUX \Data_Mem/U8137  ( .IN0(\Data_Mem/n8098 ), .IN1(\Data_Mem/n8095 ), .SEL(
        N27), .F(\Data_Mem/n8099 ) );
  MUX \Data_Mem/U8136  ( .IN0(\Data_Mem/n8097 ), .IN1(\Data_Mem/n8096 ), .SEL(
        N28), .F(\Data_Mem/n8098 ) );
  MUX \Data_Mem/U8135  ( .IN0(o[1029]), .IN1(o[1061]), .SEL(N29), .F(
        \Data_Mem/n8097 ) );
  MUX \Data_Mem/U8134  ( .IN0(o[1093]), .IN1(o[1125]), .SEL(N29), .F(
        \Data_Mem/n8096 ) );
  MUX \Data_Mem/U8133  ( .IN0(\Data_Mem/n8094 ), .IN1(\Data_Mem/n8093 ), .SEL(
        N28), .F(\Data_Mem/n8095 ) );
  MUX \Data_Mem/U8132  ( .IN0(o[1157]), .IN1(o[1189]), .SEL(N29), .F(
        \Data_Mem/n8094 ) );
  MUX \Data_Mem/U8131  ( .IN0(o[1221]), .IN1(o[1253]), .SEL(N29), .F(
        \Data_Mem/n8093 ) );
  MUX \Data_Mem/U8130  ( .IN0(\Data_Mem/n8091 ), .IN1(\Data_Mem/n8088 ), .SEL(
        N27), .F(\Data_Mem/n8092 ) );
  MUX \Data_Mem/U8129  ( .IN0(\Data_Mem/n8090 ), .IN1(\Data_Mem/n8089 ), .SEL(
        N28), .F(\Data_Mem/n8091 ) );
  MUX \Data_Mem/U8128  ( .IN0(o[1285]), .IN1(o[1317]), .SEL(N29), .F(
        \Data_Mem/n8090 ) );
  MUX \Data_Mem/U8127  ( .IN0(o[1349]), .IN1(o[1381]), .SEL(N29), .F(
        \Data_Mem/n8089 ) );
  MUX \Data_Mem/U8126  ( .IN0(\Data_Mem/n8087 ), .IN1(\Data_Mem/n8086 ), .SEL(
        N28), .F(\Data_Mem/n8088 ) );
  MUX \Data_Mem/U8125  ( .IN0(o[1413]), .IN1(o[1445]), .SEL(N29), .F(
        \Data_Mem/n8087 ) );
  MUX \Data_Mem/U8124  ( .IN0(o[1477]), .IN1(o[1509]), .SEL(N29), .F(
        \Data_Mem/n8086 ) );
  MUX \Data_Mem/U8123  ( .IN0(\Data_Mem/n8084 ), .IN1(\Data_Mem/n8077 ), .SEL(
        N26), .F(\Data_Mem/n8085 ) );
  MUX \Data_Mem/U8122  ( .IN0(\Data_Mem/n8083 ), .IN1(\Data_Mem/n8080 ), .SEL(
        N27), .F(\Data_Mem/n8084 ) );
  MUX \Data_Mem/U8121  ( .IN0(\Data_Mem/n8082 ), .IN1(\Data_Mem/n8081 ), .SEL(
        N28), .F(\Data_Mem/n8083 ) );
  MUX \Data_Mem/U8120  ( .IN0(o[1541]), .IN1(o[1573]), .SEL(N29), .F(
        \Data_Mem/n8082 ) );
  MUX \Data_Mem/U8119  ( .IN0(o[1605]), .IN1(o[1637]), .SEL(N29), .F(
        \Data_Mem/n8081 ) );
  MUX \Data_Mem/U8118  ( .IN0(\Data_Mem/n8079 ), .IN1(\Data_Mem/n8078 ), .SEL(
        N28), .F(\Data_Mem/n8080 ) );
  MUX \Data_Mem/U8117  ( .IN0(o[1669]), .IN1(o[1701]), .SEL(N29), .F(
        \Data_Mem/n8079 ) );
  MUX \Data_Mem/U8116  ( .IN0(o[1733]), .IN1(o[1765]), .SEL(N29), .F(
        \Data_Mem/n8078 ) );
  MUX \Data_Mem/U8115  ( .IN0(\Data_Mem/n8076 ), .IN1(\Data_Mem/n8073 ), .SEL(
        N27), .F(\Data_Mem/n8077 ) );
  MUX \Data_Mem/U8114  ( .IN0(\Data_Mem/n8075 ), .IN1(\Data_Mem/n8074 ), .SEL(
        N28), .F(\Data_Mem/n8076 ) );
  MUX \Data_Mem/U8113  ( .IN0(o[1797]), .IN1(o[1829]), .SEL(N29), .F(
        \Data_Mem/n8075 ) );
  MUX \Data_Mem/U8112  ( .IN0(o[1861]), .IN1(o[1893]), .SEL(N29), .F(
        \Data_Mem/n8074 ) );
  MUX \Data_Mem/U8111  ( .IN0(\Data_Mem/n8072 ), .IN1(\Data_Mem/n8071 ), .SEL(
        N28), .F(\Data_Mem/n8073 ) );
  MUX \Data_Mem/U8110  ( .IN0(o[1925]), .IN1(o[1957]), .SEL(N29), .F(
        \Data_Mem/n8072 ) );
  MUX \Data_Mem/U8109  ( .IN0(o[1989]), .IN1(o[2021]), .SEL(N29), .F(
        \Data_Mem/n8071 ) );
  MUX \Data_Mem/U8108  ( .IN0(\Data_Mem/n8070 ), .IN1(\Data_Mem/n8039 ), .SEL(
        N24), .F(\Data_Mem/N741 ) );
  MUX \Data_Mem/U8107  ( .IN0(\Data_Mem/n8069 ), .IN1(\Data_Mem/n8054 ), .SEL(
        N25), .F(\Data_Mem/n8070 ) );
  MUX \Data_Mem/U8106  ( .IN0(\Data_Mem/n8068 ), .IN1(\Data_Mem/n8061 ), .SEL(
        N26), .F(\Data_Mem/n8069 ) );
  MUX \Data_Mem/U8105  ( .IN0(\Data_Mem/n8067 ), .IN1(\Data_Mem/n8064 ), .SEL(
        N27), .F(\Data_Mem/n8068 ) );
  MUX \Data_Mem/U8104  ( .IN0(\Data_Mem/n8066 ), .IN1(\Data_Mem/n8065 ), .SEL(
        N28), .F(\Data_Mem/n8067 ) );
  MUX \Data_Mem/U8103  ( .IN0(o[4]), .IN1(o[36]), .SEL(N29), .F(
        \Data_Mem/n8066 ) );
  MUX \Data_Mem/U8102  ( .IN0(o[68]), .IN1(o[100]), .SEL(N29), .F(
        \Data_Mem/n8065 ) );
  MUX \Data_Mem/U8101  ( .IN0(\Data_Mem/n8063 ), .IN1(\Data_Mem/n8062 ), .SEL(
        N28), .F(\Data_Mem/n8064 ) );
  MUX \Data_Mem/U8100  ( .IN0(o[132]), .IN1(o[164]), .SEL(N29), .F(
        \Data_Mem/n8063 ) );
  MUX \Data_Mem/U8099  ( .IN0(o[196]), .IN1(o[228]), .SEL(N29), .F(
        \Data_Mem/n8062 ) );
  MUX \Data_Mem/U8098  ( .IN0(\Data_Mem/n8060 ), .IN1(\Data_Mem/n8057 ), .SEL(
        N27), .F(\Data_Mem/n8061 ) );
  MUX \Data_Mem/U8097  ( .IN0(\Data_Mem/n8059 ), .IN1(\Data_Mem/n8058 ), .SEL(
        N28), .F(\Data_Mem/n8060 ) );
  MUX \Data_Mem/U8096  ( .IN0(o[260]), .IN1(o[292]), .SEL(N29), .F(
        \Data_Mem/n8059 ) );
  MUX \Data_Mem/U8095  ( .IN0(o[324]), .IN1(o[356]), .SEL(N29), .F(
        \Data_Mem/n8058 ) );
  MUX \Data_Mem/U8094  ( .IN0(\Data_Mem/n8056 ), .IN1(\Data_Mem/n8055 ), .SEL(
        N28), .F(\Data_Mem/n8057 ) );
  MUX \Data_Mem/U8093  ( .IN0(o[388]), .IN1(o[420]), .SEL(N29), .F(
        \Data_Mem/n8056 ) );
  MUX \Data_Mem/U8092  ( .IN0(o[452]), .IN1(o[484]), .SEL(N29), .F(
        \Data_Mem/n8055 ) );
  MUX \Data_Mem/U8091  ( .IN0(\Data_Mem/n8053 ), .IN1(\Data_Mem/n8046 ), .SEL(
        N26), .F(\Data_Mem/n8054 ) );
  MUX \Data_Mem/U8090  ( .IN0(\Data_Mem/n8052 ), .IN1(\Data_Mem/n8049 ), .SEL(
        N27), .F(\Data_Mem/n8053 ) );
  MUX \Data_Mem/U8089  ( .IN0(\Data_Mem/n8051 ), .IN1(\Data_Mem/n8050 ), .SEL(
        N28), .F(\Data_Mem/n8052 ) );
  MUX \Data_Mem/U8088  ( .IN0(o[516]), .IN1(o[548]), .SEL(N29), .F(
        \Data_Mem/n8051 ) );
  MUX \Data_Mem/U8087  ( .IN0(o[580]), .IN1(o[612]), .SEL(N29), .F(
        \Data_Mem/n8050 ) );
  MUX \Data_Mem/U8086  ( .IN0(\Data_Mem/n8048 ), .IN1(\Data_Mem/n8047 ), .SEL(
        N28), .F(\Data_Mem/n8049 ) );
  MUX \Data_Mem/U8085  ( .IN0(o[644]), .IN1(o[676]), .SEL(N29), .F(
        \Data_Mem/n8048 ) );
  MUX \Data_Mem/U8084  ( .IN0(o[708]), .IN1(o[740]), .SEL(N29), .F(
        \Data_Mem/n8047 ) );
  MUX \Data_Mem/U8083  ( .IN0(\Data_Mem/n8045 ), .IN1(\Data_Mem/n8042 ), .SEL(
        N27), .F(\Data_Mem/n8046 ) );
  MUX \Data_Mem/U8082  ( .IN0(\Data_Mem/n8044 ), .IN1(\Data_Mem/n8043 ), .SEL(
        N28), .F(\Data_Mem/n8045 ) );
  MUX \Data_Mem/U8081  ( .IN0(o[772]), .IN1(o[804]), .SEL(N29), .F(
        \Data_Mem/n8044 ) );
  MUX \Data_Mem/U8080  ( .IN0(o[836]), .IN1(o[868]), .SEL(N29), .F(
        \Data_Mem/n8043 ) );
  MUX \Data_Mem/U8079  ( .IN0(\Data_Mem/n8041 ), .IN1(\Data_Mem/n8040 ), .SEL(
        N28), .F(\Data_Mem/n8042 ) );
  MUX \Data_Mem/U8078  ( .IN0(o[900]), .IN1(o[932]), .SEL(N29), .F(
        \Data_Mem/n8041 ) );
  MUX \Data_Mem/U8077  ( .IN0(o[964]), .IN1(o[996]), .SEL(N29), .F(
        \Data_Mem/n8040 ) );
  MUX \Data_Mem/U8076  ( .IN0(\Data_Mem/n8038 ), .IN1(\Data_Mem/n8023 ), .SEL(
        N25), .F(\Data_Mem/n8039 ) );
  MUX \Data_Mem/U8075  ( .IN0(\Data_Mem/n8037 ), .IN1(\Data_Mem/n8030 ), .SEL(
        N26), .F(\Data_Mem/n8038 ) );
  MUX \Data_Mem/U8074  ( .IN0(\Data_Mem/n8036 ), .IN1(\Data_Mem/n8033 ), .SEL(
        N27), .F(\Data_Mem/n8037 ) );
  MUX \Data_Mem/U8073  ( .IN0(\Data_Mem/n8035 ), .IN1(\Data_Mem/n8034 ), .SEL(
        N28), .F(\Data_Mem/n8036 ) );
  MUX \Data_Mem/U8072  ( .IN0(o[1028]), .IN1(o[1060]), .SEL(N29), .F(
        \Data_Mem/n8035 ) );
  MUX \Data_Mem/U8071  ( .IN0(o[1092]), .IN1(o[1124]), .SEL(N29), .F(
        \Data_Mem/n8034 ) );
  MUX \Data_Mem/U8070  ( .IN0(\Data_Mem/n8032 ), .IN1(\Data_Mem/n8031 ), .SEL(
        N28), .F(\Data_Mem/n8033 ) );
  MUX \Data_Mem/U8069  ( .IN0(o[1156]), .IN1(o[1188]), .SEL(N29), .F(
        \Data_Mem/n8032 ) );
  MUX \Data_Mem/U8068  ( .IN0(o[1220]), .IN1(o[1252]), .SEL(N29), .F(
        \Data_Mem/n8031 ) );
  MUX \Data_Mem/U8067  ( .IN0(\Data_Mem/n8029 ), .IN1(\Data_Mem/n8026 ), .SEL(
        N27), .F(\Data_Mem/n8030 ) );
  MUX \Data_Mem/U8066  ( .IN0(\Data_Mem/n8028 ), .IN1(\Data_Mem/n8027 ), .SEL(
        N28), .F(\Data_Mem/n8029 ) );
  MUX \Data_Mem/U8065  ( .IN0(o[1284]), .IN1(o[1316]), .SEL(N29), .F(
        \Data_Mem/n8028 ) );
  MUX \Data_Mem/U8064  ( .IN0(o[1348]), .IN1(o[1380]), .SEL(N29), .F(
        \Data_Mem/n8027 ) );
  MUX \Data_Mem/U8063  ( .IN0(\Data_Mem/n8025 ), .IN1(\Data_Mem/n8024 ), .SEL(
        N28), .F(\Data_Mem/n8026 ) );
  MUX \Data_Mem/U8062  ( .IN0(o[1412]), .IN1(o[1444]), .SEL(N29), .F(
        \Data_Mem/n8025 ) );
  MUX \Data_Mem/U8061  ( .IN0(o[1476]), .IN1(o[1508]), .SEL(N29), .F(
        \Data_Mem/n8024 ) );
  MUX \Data_Mem/U8060  ( .IN0(\Data_Mem/n8022 ), .IN1(\Data_Mem/n8015 ), .SEL(
        N26), .F(\Data_Mem/n8023 ) );
  MUX \Data_Mem/U8059  ( .IN0(\Data_Mem/n8021 ), .IN1(\Data_Mem/n8018 ), .SEL(
        N27), .F(\Data_Mem/n8022 ) );
  MUX \Data_Mem/U8058  ( .IN0(\Data_Mem/n8020 ), .IN1(\Data_Mem/n8019 ), .SEL(
        N28), .F(\Data_Mem/n8021 ) );
  MUX \Data_Mem/U8057  ( .IN0(o[1540]), .IN1(o[1572]), .SEL(N29), .F(
        \Data_Mem/n8020 ) );
  MUX \Data_Mem/U8056  ( .IN0(o[1604]), .IN1(o[1636]), .SEL(N29), .F(
        \Data_Mem/n8019 ) );
  MUX \Data_Mem/U8055  ( .IN0(\Data_Mem/n8017 ), .IN1(\Data_Mem/n8016 ), .SEL(
        N28), .F(\Data_Mem/n8018 ) );
  MUX \Data_Mem/U8054  ( .IN0(o[1668]), .IN1(o[1700]), .SEL(N29), .F(
        \Data_Mem/n8017 ) );
  MUX \Data_Mem/U8053  ( .IN0(o[1732]), .IN1(o[1764]), .SEL(N29), .F(
        \Data_Mem/n8016 ) );
  MUX \Data_Mem/U8052  ( .IN0(\Data_Mem/n8014 ), .IN1(\Data_Mem/n8011 ), .SEL(
        N27), .F(\Data_Mem/n8015 ) );
  MUX \Data_Mem/U8051  ( .IN0(\Data_Mem/n8013 ), .IN1(\Data_Mem/n8012 ), .SEL(
        N28), .F(\Data_Mem/n8014 ) );
  MUX \Data_Mem/U8050  ( .IN0(o[1796]), .IN1(o[1828]), .SEL(N29), .F(
        \Data_Mem/n8013 ) );
  MUX \Data_Mem/U8049  ( .IN0(o[1860]), .IN1(o[1892]), .SEL(N29), .F(
        \Data_Mem/n8012 ) );
  MUX \Data_Mem/U8048  ( .IN0(\Data_Mem/n8010 ), .IN1(\Data_Mem/n8009 ), .SEL(
        N28), .F(\Data_Mem/n8011 ) );
  MUX \Data_Mem/U8047  ( .IN0(o[1924]), .IN1(o[1956]), .SEL(N29), .F(
        \Data_Mem/n8010 ) );
  MUX \Data_Mem/U8046  ( .IN0(o[1988]), .IN1(o[2020]), .SEL(N29), .F(
        \Data_Mem/n8009 ) );
  MUX \Data_Mem/U8045  ( .IN0(\Data_Mem/n8008 ), .IN1(\Data_Mem/n7977 ), .SEL(
        N24), .F(\Data_Mem/N742 ) );
  MUX \Data_Mem/U8044  ( .IN0(\Data_Mem/n8007 ), .IN1(\Data_Mem/n7992 ), .SEL(
        N25), .F(\Data_Mem/n8008 ) );
  MUX \Data_Mem/U8043  ( .IN0(\Data_Mem/n8006 ), .IN1(\Data_Mem/n7999 ), .SEL(
        N26), .F(\Data_Mem/n8007 ) );
  MUX \Data_Mem/U8042  ( .IN0(\Data_Mem/n8005 ), .IN1(\Data_Mem/n8002 ), .SEL(
        N27), .F(\Data_Mem/n8006 ) );
  MUX \Data_Mem/U8041  ( .IN0(\Data_Mem/n8004 ), .IN1(\Data_Mem/n8003 ), .SEL(
        N28), .F(\Data_Mem/n8005 ) );
  MUX \Data_Mem/U8040  ( .IN0(o[3]), .IN1(o[35]), .SEL(N29), .F(
        \Data_Mem/n8004 ) );
  MUX \Data_Mem/U8039  ( .IN0(o[67]), .IN1(o[99]), .SEL(N29), .F(
        \Data_Mem/n8003 ) );
  MUX \Data_Mem/U8038  ( .IN0(\Data_Mem/n8001 ), .IN1(\Data_Mem/n8000 ), .SEL(
        N28), .F(\Data_Mem/n8002 ) );
  MUX \Data_Mem/U8037  ( .IN0(o[131]), .IN1(o[163]), .SEL(N29), .F(
        \Data_Mem/n8001 ) );
  MUX \Data_Mem/U8036  ( .IN0(o[195]), .IN1(o[227]), .SEL(N29), .F(
        \Data_Mem/n8000 ) );
  MUX \Data_Mem/U8035  ( .IN0(\Data_Mem/n7998 ), .IN1(\Data_Mem/n7995 ), .SEL(
        N27), .F(\Data_Mem/n7999 ) );
  MUX \Data_Mem/U8034  ( .IN0(\Data_Mem/n7997 ), .IN1(\Data_Mem/n7996 ), .SEL(
        N28), .F(\Data_Mem/n7998 ) );
  MUX \Data_Mem/U8033  ( .IN0(o[259]), .IN1(o[291]), .SEL(N29), .F(
        \Data_Mem/n7997 ) );
  MUX \Data_Mem/U8032  ( .IN0(o[323]), .IN1(o[355]), .SEL(N29), .F(
        \Data_Mem/n7996 ) );
  MUX \Data_Mem/U8031  ( .IN0(\Data_Mem/n7994 ), .IN1(\Data_Mem/n7993 ), .SEL(
        N28), .F(\Data_Mem/n7995 ) );
  MUX \Data_Mem/U8030  ( .IN0(o[387]), .IN1(o[419]), .SEL(N29), .F(
        \Data_Mem/n7994 ) );
  MUX \Data_Mem/U8029  ( .IN0(o[451]), .IN1(o[483]), .SEL(N29), .F(
        \Data_Mem/n7993 ) );
  MUX \Data_Mem/U8028  ( .IN0(\Data_Mem/n7991 ), .IN1(\Data_Mem/n7984 ), .SEL(
        N26), .F(\Data_Mem/n7992 ) );
  MUX \Data_Mem/U8027  ( .IN0(\Data_Mem/n7990 ), .IN1(\Data_Mem/n7987 ), .SEL(
        N27), .F(\Data_Mem/n7991 ) );
  MUX \Data_Mem/U8026  ( .IN0(\Data_Mem/n7989 ), .IN1(\Data_Mem/n7988 ), .SEL(
        N28), .F(\Data_Mem/n7990 ) );
  MUX \Data_Mem/U8025  ( .IN0(o[515]), .IN1(o[547]), .SEL(N29), .F(
        \Data_Mem/n7989 ) );
  MUX \Data_Mem/U8024  ( .IN0(o[579]), .IN1(o[611]), .SEL(N29), .F(
        \Data_Mem/n7988 ) );
  MUX \Data_Mem/U8023  ( .IN0(\Data_Mem/n7986 ), .IN1(\Data_Mem/n7985 ), .SEL(
        N28), .F(\Data_Mem/n7987 ) );
  MUX \Data_Mem/U8022  ( .IN0(o[643]), .IN1(o[675]), .SEL(N29), .F(
        \Data_Mem/n7986 ) );
  MUX \Data_Mem/U8021  ( .IN0(o[707]), .IN1(o[739]), .SEL(N29), .F(
        \Data_Mem/n7985 ) );
  MUX \Data_Mem/U8020  ( .IN0(\Data_Mem/n7983 ), .IN1(\Data_Mem/n7980 ), .SEL(
        N27), .F(\Data_Mem/n7984 ) );
  MUX \Data_Mem/U8019  ( .IN0(\Data_Mem/n7982 ), .IN1(\Data_Mem/n7981 ), .SEL(
        N28), .F(\Data_Mem/n7983 ) );
  MUX \Data_Mem/U8018  ( .IN0(o[771]), .IN1(o[803]), .SEL(N29), .F(
        \Data_Mem/n7982 ) );
  MUX \Data_Mem/U8017  ( .IN0(o[835]), .IN1(o[867]), .SEL(N29), .F(
        \Data_Mem/n7981 ) );
  MUX \Data_Mem/U8016  ( .IN0(\Data_Mem/n7979 ), .IN1(\Data_Mem/n7978 ), .SEL(
        N28), .F(\Data_Mem/n7980 ) );
  MUX \Data_Mem/U8015  ( .IN0(o[899]), .IN1(o[931]), .SEL(N29), .F(
        \Data_Mem/n7979 ) );
  MUX \Data_Mem/U8014  ( .IN0(o[963]), .IN1(o[995]), .SEL(N29), .F(
        \Data_Mem/n7978 ) );
  MUX \Data_Mem/U8013  ( .IN0(\Data_Mem/n7976 ), .IN1(\Data_Mem/n7961 ), .SEL(
        N25), .F(\Data_Mem/n7977 ) );
  MUX \Data_Mem/U8012  ( .IN0(\Data_Mem/n7975 ), .IN1(\Data_Mem/n7968 ), .SEL(
        N26), .F(\Data_Mem/n7976 ) );
  MUX \Data_Mem/U8011  ( .IN0(\Data_Mem/n7974 ), .IN1(\Data_Mem/n7971 ), .SEL(
        N27), .F(\Data_Mem/n7975 ) );
  MUX \Data_Mem/U8010  ( .IN0(\Data_Mem/n7973 ), .IN1(\Data_Mem/n7972 ), .SEL(
        N28), .F(\Data_Mem/n7974 ) );
  MUX \Data_Mem/U8009  ( .IN0(o[1027]), .IN1(o[1059]), .SEL(N29), .F(
        \Data_Mem/n7973 ) );
  MUX \Data_Mem/U8008  ( .IN0(o[1091]), .IN1(o[1123]), .SEL(N29), .F(
        \Data_Mem/n7972 ) );
  MUX \Data_Mem/U8007  ( .IN0(\Data_Mem/n7970 ), .IN1(\Data_Mem/n7969 ), .SEL(
        N28), .F(\Data_Mem/n7971 ) );
  MUX \Data_Mem/U8006  ( .IN0(o[1155]), .IN1(o[1187]), .SEL(N29), .F(
        \Data_Mem/n7970 ) );
  MUX \Data_Mem/U8005  ( .IN0(o[1219]), .IN1(o[1251]), .SEL(N29), .F(
        \Data_Mem/n7969 ) );
  MUX \Data_Mem/U8004  ( .IN0(\Data_Mem/n7967 ), .IN1(\Data_Mem/n7964 ), .SEL(
        N27), .F(\Data_Mem/n7968 ) );
  MUX \Data_Mem/U8003  ( .IN0(\Data_Mem/n7966 ), .IN1(\Data_Mem/n7965 ), .SEL(
        N28), .F(\Data_Mem/n7967 ) );
  MUX \Data_Mem/U8002  ( .IN0(o[1283]), .IN1(o[1315]), .SEL(N29), .F(
        \Data_Mem/n7966 ) );
  MUX \Data_Mem/U8001  ( .IN0(o[1347]), .IN1(o[1379]), .SEL(N29), .F(
        \Data_Mem/n7965 ) );
  MUX \Data_Mem/U8000  ( .IN0(\Data_Mem/n7963 ), .IN1(\Data_Mem/n7962 ), .SEL(
        N28), .F(\Data_Mem/n7964 ) );
  MUX \Data_Mem/U7999  ( .IN0(o[1411]), .IN1(o[1443]), .SEL(N29), .F(
        \Data_Mem/n7963 ) );
  MUX \Data_Mem/U7998  ( .IN0(o[1475]), .IN1(o[1507]), .SEL(N29), .F(
        \Data_Mem/n7962 ) );
  MUX \Data_Mem/U7997  ( .IN0(\Data_Mem/n7960 ), .IN1(\Data_Mem/n7953 ), .SEL(
        N26), .F(\Data_Mem/n7961 ) );
  MUX \Data_Mem/U7996  ( .IN0(\Data_Mem/n7959 ), .IN1(\Data_Mem/n7956 ), .SEL(
        N27), .F(\Data_Mem/n7960 ) );
  MUX \Data_Mem/U7995  ( .IN0(\Data_Mem/n7958 ), .IN1(\Data_Mem/n7957 ), .SEL(
        N28), .F(\Data_Mem/n7959 ) );
  MUX \Data_Mem/U7994  ( .IN0(o[1539]), .IN1(o[1571]), .SEL(N29), .F(
        \Data_Mem/n7958 ) );
  MUX \Data_Mem/U7993  ( .IN0(o[1603]), .IN1(o[1635]), .SEL(N29), .F(
        \Data_Mem/n7957 ) );
  MUX \Data_Mem/U7992  ( .IN0(\Data_Mem/n7955 ), .IN1(\Data_Mem/n7954 ), .SEL(
        N28), .F(\Data_Mem/n7956 ) );
  MUX \Data_Mem/U7991  ( .IN0(o[1667]), .IN1(o[1699]), .SEL(N29), .F(
        \Data_Mem/n7955 ) );
  MUX \Data_Mem/U7990  ( .IN0(o[1731]), .IN1(o[1763]), .SEL(N29), .F(
        \Data_Mem/n7954 ) );
  MUX \Data_Mem/U7989  ( .IN0(\Data_Mem/n7952 ), .IN1(\Data_Mem/n7949 ), .SEL(
        N27), .F(\Data_Mem/n7953 ) );
  MUX \Data_Mem/U7988  ( .IN0(\Data_Mem/n7951 ), .IN1(\Data_Mem/n7950 ), .SEL(
        N28), .F(\Data_Mem/n7952 ) );
  MUX \Data_Mem/U7987  ( .IN0(o[1795]), .IN1(o[1827]), .SEL(N29), .F(
        \Data_Mem/n7951 ) );
  MUX \Data_Mem/U7986  ( .IN0(o[1859]), .IN1(o[1891]), .SEL(N29), .F(
        \Data_Mem/n7950 ) );
  MUX \Data_Mem/U7985  ( .IN0(\Data_Mem/n7948 ), .IN1(\Data_Mem/n7947 ), .SEL(
        N28), .F(\Data_Mem/n7949 ) );
  MUX \Data_Mem/U7984  ( .IN0(o[1923]), .IN1(o[1955]), .SEL(N29), .F(
        \Data_Mem/n7948 ) );
  MUX \Data_Mem/U7983  ( .IN0(o[1987]), .IN1(o[2019]), .SEL(N29), .F(
        \Data_Mem/n7947 ) );
  MUX \Data_Mem/U7982  ( .IN0(\Data_Mem/n7946 ), .IN1(\Data_Mem/n7915 ), .SEL(
        N24), .F(\Data_Mem/N743 ) );
  MUX \Data_Mem/U7981  ( .IN0(\Data_Mem/n7945 ), .IN1(\Data_Mem/n7930 ), .SEL(
        N25), .F(\Data_Mem/n7946 ) );
  MUX \Data_Mem/U7980  ( .IN0(\Data_Mem/n7944 ), .IN1(\Data_Mem/n7937 ), .SEL(
        N26), .F(\Data_Mem/n7945 ) );
  MUX \Data_Mem/U7979  ( .IN0(\Data_Mem/n7943 ), .IN1(\Data_Mem/n7940 ), .SEL(
        N27), .F(\Data_Mem/n7944 ) );
  MUX \Data_Mem/U7978  ( .IN0(\Data_Mem/n7942 ), .IN1(\Data_Mem/n7941 ), .SEL(
        N28), .F(\Data_Mem/n7943 ) );
  MUX \Data_Mem/U7977  ( .IN0(o[2]), .IN1(o[34]), .SEL(N29), .F(
        \Data_Mem/n7942 ) );
  MUX \Data_Mem/U7976  ( .IN0(o[66]), .IN1(o[98]), .SEL(N29), .F(
        \Data_Mem/n7941 ) );
  MUX \Data_Mem/U7975  ( .IN0(\Data_Mem/n7939 ), .IN1(\Data_Mem/n7938 ), .SEL(
        N28), .F(\Data_Mem/n7940 ) );
  MUX \Data_Mem/U7974  ( .IN0(o[130]), .IN1(o[162]), .SEL(N29), .F(
        \Data_Mem/n7939 ) );
  MUX \Data_Mem/U7973  ( .IN0(o[194]), .IN1(o[226]), .SEL(N29), .F(
        \Data_Mem/n7938 ) );
  MUX \Data_Mem/U7972  ( .IN0(\Data_Mem/n7936 ), .IN1(\Data_Mem/n7933 ), .SEL(
        N27), .F(\Data_Mem/n7937 ) );
  MUX \Data_Mem/U7971  ( .IN0(\Data_Mem/n7935 ), .IN1(\Data_Mem/n7934 ), .SEL(
        N28), .F(\Data_Mem/n7936 ) );
  MUX \Data_Mem/U7970  ( .IN0(o[258]), .IN1(o[290]), .SEL(N29), .F(
        \Data_Mem/n7935 ) );
  MUX \Data_Mem/U7969  ( .IN0(o[322]), .IN1(o[354]), .SEL(N29), .F(
        \Data_Mem/n7934 ) );
  MUX \Data_Mem/U7968  ( .IN0(\Data_Mem/n7932 ), .IN1(\Data_Mem/n7931 ), .SEL(
        N28), .F(\Data_Mem/n7933 ) );
  MUX \Data_Mem/U7967  ( .IN0(o[386]), .IN1(o[418]), .SEL(N29), .F(
        \Data_Mem/n7932 ) );
  MUX \Data_Mem/U7966  ( .IN0(o[450]), .IN1(o[482]), .SEL(N29), .F(
        \Data_Mem/n7931 ) );
  MUX \Data_Mem/U7965  ( .IN0(\Data_Mem/n7929 ), .IN1(\Data_Mem/n7922 ), .SEL(
        N26), .F(\Data_Mem/n7930 ) );
  MUX \Data_Mem/U7964  ( .IN0(\Data_Mem/n7928 ), .IN1(\Data_Mem/n7925 ), .SEL(
        N27), .F(\Data_Mem/n7929 ) );
  MUX \Data_Mem/U7963  ( .IN0(\Data_Mem/n7927 ), .IN1(\Data_Mem/n7926 ), .SEL(
        N28), .F(\Data_Mem/n7928 ) );
  MUX \Data_Mem/U7962  ( .IN0(o[514]), .IN1(o[546]), .SEL(N29), .F(
        \Data_Mem/n7927 ) );
  MUX \Data_Mem/U7961  ( .IN0(o[578]), .IN1(o[610]), .SEL(N29), .F(
        \Data_Mem/n7926 ) );
  MUX \Data_Mem/U7960  ( .IN0(\Data_Mem/n7924 ), .IN1(\Data_Mem/n7923 ), .SEL(
        N28), .F(\Data_Mem/n7925 ) );
  MUX \Data_Mem/U7959  ( .IN0(o[642]), .IN1(o[674]), .SEL(N29), .F(
        \Data_Mem/n7924 ) );
  MUX \Data_Mem/U7958  ( .IN0(o[706]), .IN1(o[738]), .SEL(N29), .F(
        \Data_Mem/n7923 ) );
  MUX \Data_Mem/U7957  ( .IN0(\Data_Mem/n7921 ), .IN1(\Data_Mem/n7918 ), .SEL(
        N27), .F(\Data_Mem/n7922 ) );
  MUX \Data_Mem/U7956  ( .IN0(\Data_Mem/n7920 ), .IN1(\Data_Mem/n7919 ), .SEL(
        N28), .F(\Data_Mem/n7921 ) );
  MUX \Data_Mem/U7955  ( .IN0(o[770]), .IN1(o[802]), .SEL(N29), .F(
        \Data_Mem/n7920 ) );
  MUX \Data_Mem/U7954  ( .IN0(o[834]), .IN1(o[866]), .SEL(N29), .F(
        \Data_Mem/n7919 ) );
  MUX \Data_Mem/U7953  ( .IN0(\Data_Mem/n7917 ), .IN1(\Data_Mem/n7916 ), .SEL(
        N28), .F(\Data_Mem/n7918 ) );
  MUX \Data_Mem/U7952  ( .IN0(o[898]), .IN1(o[930]), .SEL(N29), .F(
        \Data_Mem/n7917 ) );
  MUX \Data_Mem/U7951  ( .IN0(o[962]), .IN1(o[994]), .SEL(N29), .F(
        \Data_Mem/n7916 ) );
  MUX \Data_Mem/U7950  ( .IN0(\Data_Mem/n7914 ), .IN1(\Data_Mem/n7899 ), .SEL(
        N25), .F(\Data_Mem/n7915 ) );
  MUX \Data_Mem/U7949  ( .IN0(\Data_Mem/n7913 ), .IN1(\Data_Mem/n7906 ), .SEL(
        N26), .F(\Data_Mem/n7914 ) );
  MUX \Data_Mem/U7948  ( .IN0(\Data_Mem/n7912 ), .IN1(\Data_Mem/n7909 ), .SEL(
        N27), .F(\Data_Mem/n7913 ) );
  MUX \Data_Mem/U7947  ( .IN0(\Data_Mem/n7911 ), .IN1(\Data_Mem/n7910 ), .SEL(
        N28), .F(\Data_Mem/n7912 ) );
  MUX \Data_Mem/U7946  ( .IN0(o[1026]), .IN1(o[1058]), .SEL(N29), .F(
        \Data_Mem/n7911 ) );
  MUX \Data_Mem/U7945  ( .IN0(o[1090]), .IN1(o[1122]), .SEL(N29), .F(
        \Data_Mem/n7910 ) );
  MUX \Data_Mem/U7944  ( .IN0(\Data_Mem/n7908 ), .IN1(\Data_Mem/n7907 ), .SEL(
        N28), .F(\Data_Mem/n7909 ) );
  MUX \Data_Mem/U7943  ( .IN0(o[1154]), .IN1(o[1186]), .SEL(N29), .F(
        \Data_Mem/n7908 ) );
  MUX \Data_Mem/U7942  ( .IN0(o[1218]), .IN1(o[1250]), .SEL(N29), .F(
        \Data_Mem/n7907 ) );
  MUX \Data_Mem/U7941  ( .IN0(\Data_Mem/n7905 ), .IN1(\Data_Mem/n7902 ), .SEL(
        N27), .F(\Data_Mem/n7906 ) );
  MUX \Data_Mem/U7940  ( .IN0(\Data_Mem/n7904 ), .IN1(\Data_Mem/n7903 ), .SEL(
        N28), .F(\Data_Mem/n7905 ) );
  MUX \Data_Mem/U7939  ( .IN0(o[1282]), .IN1(o[1314]), .SEL(N29), .F(
        \Data_Mem/n7904 ) );
  MUX \Data_Mem/U7938  ( .IN0(o[1346]), .IN1(o[1378]), .SEL(N29), .F(
        \Data_Mem/n7903 ) );
  MUX \Data_Mem/U7937  ( .IN0(\Data_Mem/n7901 ), .IN1(\Data_Mem/n7900 ), .SEL(
        N28), .F(\Data_Mem/n7902 ) );
  MUX \Data_Mem/U7936  ( .IN0(o[1410]), .IN1(o[1442]), .SEL(N29), .F(
        \Data_Mem/n7901 ) );
  MUX \Data_Mem/U7935  ( .IN0(o[1474]), .IN1(o[1506]), .SEL(N29), .F(
        \Data_Mem/n7900 ) );
  MUX \Data_Mem/U7934  ( .IN0(\Data_Mem/n7898 ), .IN1(\Data_Mem/n7891 ), .SEL(
        N26), .F(\Data_Mem/n7899 ) );
  MUX \Data_Mem/U7933  ( .IN0(\Data_Mem/n7897 ), .IN1(\Data_Mem/n7894 ), .SEL(
        N27), .F(\Data_Mem/n7898 ) );
  MUX \Data_Mem/U7932  ( .IN0(\Data_Mem/n7896 ), .IN1(\Data_Mem/n7895 ), .SEL(
        N28), .F(\Data_Mem/n7897 ) );
  MUX \Data_Mem/U7931  ( .IN0(o[1538]), .IN1(o[1570]), .SEL(N29), .F(
        \Data_Mem/n7896 ) );
  MUX \Data_Mem/U7930  ( .IN0(o[1602]), .IN1(o[1634]), .SEL(N29), .F(
        \Data_Mem/n7895 ) );
  MUX \Data_Mem/U7929  ( .IN0(\Data_Mem/n7893 ), .IN1(\Data_Mem/n7892 ), .SEL(
        N28), .F(\Data_Mem/n7894 ) );
  MUX \Data_Mem/U7928  ( .IN0(o[1666]), .IN1(o[1698]), .SEL(N29), .F(
        \Data_Mem/n7893 ) );
  MUX \Data_Mem/U7927  ( .IN0(o[1730]), .IN1(o[1762]), .SEL(N29), .F(
        \Data_Mem/n7892 ) );
  MUX \Data_Mem/U7926  ( .IN0(\Data_Mem/n7890 ), .IN1(\Data_Mem/n7887 ), .SEL(
        N27), .F(\Data_Mem/n7891 ) );
  MUX \Data_Mem/U7925  ( .IN0(\Data_Mem/n7889 ), .IN1(\Data_Mem/n7888 ), .SEL(
        N28), .F(\Data_Mem/n7890 ) );
  MUX \Data_Mem/U7924  ( .IN0(o[1794]), .IN1(o[1826]), .SEL(N29), .F(
        \Data_Mem/n7889 ) );
  MUX \Data_Mem/U7923  ( .IN0(o[1858]), .IN1(o[1890]), .SEL(N29), .F(
        \Data_Mem/n7888 ) );
  MUX \Data_Mem/U7922  ( .IN0(\Data_Mem/n7886 ), .IN1(\Data_Mem/n7885 ), .SEL(
        N28), .F(\Data_Mem/n7887 ) );
  MUX \Data_Mem/U7921  ( .IN0(o[1922]), .IN1(o[1954]), .SEL(N29), .F(
        \Data_Mem/n7886 ) );
  MUX \Data_Mem/U7920  ( .IN0(o[1986]), .IN1(o[2018]), .SEL(N29), .F(
        \Data_Mem/n7885 ) );
  MUX \Data_Mem/U7919  ( .IN0(\Data_Mem/n7884 ), .IN1(\Data_Mem/n7853 ), .SEL(
        N24), .F(\Data_Mem/N744 ) );
  MUX \Data_Mem/U7918  ( .IN0(\Data_Mem/n7883 ), .IN1(\Data_Mem/n7868 ), .SEL(
        N25), .F(\Data_Mem/n7884 ) );
  MUX \Data_Mem/U7917  ( .IN0(\Data_Mem/n7882 ), .IN1(\Data_Mem/n7875 ), .SEL(
        N26), .F(\Data_Mem/n7883 ) );
  MUX \Data_Mem/U7916  ( .IN0(\Data_Mem/n7881 ), .IN1(\Data_Mem/n7878 ), .SEL(
        N27), .F(\Data_Mem/n7882 ) );
  MUX \Data_Mem/U7915  ( .IN0(\Data_Mem/n7880 ), .IN1(\Data_Mem/n7879 ), .SEL(
        N28), .F(\Data_Mem/n7881 ) );
  MUX \Data_Mem/U7914  ( .IN0(o[1]), .IN1(o[33]), .SEL(N29), .F(
        \Data_Mem/n7880 ) );
  MUX \Data_Mem/U7913  ( .IN0(o[65]), .IN1(o[97]), .SEL(N29), .F(
        \Data_Mem/n7879 ) );
  MUX \Data_Mem/U7912  ( .IN0(\Data_Mem/n7877 ), .IN1(\Data_Mem/n7876 ), .SEL(
        N28), .F(\Data_Mem/n7878 ) );
  MUX \Data_Mem/U7911  ( .IN0(o[129]), .IN1(o[161]), .SEL(N29), .F(
        \Data_Mem/n7877 ) );
  MUX \Data_Mem/U7910  ( .IN0(o[193]), .IN1(o[225]), .SEL(N29), .F(
        \Data_Mem/n7876 ) );
  MUX \Data_Mem/U7909  ( .IN0(\Data_Mem/n7874 ), .IN1(\Data_Mem/n7871 ), .SEL(
        N27), .F(\Data_Mem/n7875 ) );
  MUX \Data_Mem/U7908  ( .IN0(\Data_Mem/n7873 ), .IN1(\Data_Mem/n7872 ), .SEL(
        N28), .F(\Data_Mem/n7874 ) );
  MUX \Data_Mem/U7907  ( .IN0(o[257]), .IN1(o[289]), .SEL(N29), .F(
        \Data_Mem/n7873 ) );
  MUX \Data_Mem/U7906  ( .IN0(o[321]), .IN1(o[353]), .SEL(N29), .F(
        \Data_Mem/n7872 ) );
  MUX \Data_Mem/U7905  ( .IN0(\Data_Mem/n7870 ), .IN1(\Data_Mem/n7869 ), .SEL(
        N28), .F(\Data_Mem/n7871 ) );
  MUX \Data_Mem/U7904  ( .IN0(o[385]), .IN1(o[417]), .SEL(N29), .F(
        \Data_Mem/n7870 ) );
  MUX \Data_Mem/U7903  ( .IN0(o[449]), .IN1(o[481]), .SEL(N29), .F(
        \Data_Mem/n7869 ) );
  MUX \Data_Mem/U7902  ( .IN0(\Data_Mem/n7867 ), .IN1(\Data_Mem/n7860 ), .SEL(
        N26), .F(\Data_Mem/n7868 ) );
  MUX \Data_Mem/U7901  ( .IN0(\Data_Mem/n7866 ), .IN1(\Data_Mem/n7863 ), .SEL(
        N27), .F(\Data_Mem/n7867 ) );
  MUX \Data_Mem/U7900  ( .IN0(\Data_Mem/n7865 ), .IN1(\Data_Mem/n7864 ), .SEL(
        N28), .F(\Data_Mem/n7866 ) );
  MUX \Data_Mem/U7899  ( .IN0(o[513]), .IN1(o[545]), .SEL(N29), .F(
        \Data_Mem/n7865 ) );
  MUX \Data_Mem/U7898  ( .IN0(o[577]), .IN1(o[609]), .SEL(N29), .F(
        \Data_Mem/n7864 ) );
  MUX \Data_Mem/U7897  ( .IN0(\Data_Mem/n7862 ), .IN1(\Data_Mem/n7861 ), .SEL(
        N28), .F(\Data_Mem/n7863 ) );
  MUX \Data_Mem/U7896  ( .IN0(o[641]), .IN1(o[673]), .SEL(N29), .F(
        \Data_Mem/n7862 ) );
  MUX \Data_Mem/U7895  ( .IN0(o[705]), .IN1(o[737]), .SEL(N29), .F(
        \Data_Mem/n7861 ) );
  MUX \Data_Mem/U7894  ( .IN0(\Data_Mem/n7859 ), .IN1(\Data_Mem/n7856 ), .SEL(
        N27), .F(\Data_Mem/n7860 ) );
  MUX \Data_Mem/U7893  ( .IN0(\Data_Mem/n7858 ), .IN1(\Data_Mem/n7857 ), .SEL(
        N28), .F(\Data_Mem/n7859 ) );
  MUX \Data_Mem/U7892  ( .IN0(o[769]), .IN1(o[801]), .SEL(N29), .F(
        \Data_Mem/n7858 ) );
  MUX \Data_Mem/U7891  ( .IN0(o[833]), .IN1(o[865]), .SEL(N29), .F(
        \Data_Mem/n7857 ) );
  MUX \Data_Mem/U7890  ( .IN0(\Data_Mem/n7855 ), .IN1(\Data_Mem/n7854 ), .SEL(
        N28), .F(\Data_Mem/n7856 ) );
  MUX \Data_Mem/U7889  ( .IN0(o[897]), .IN1(o[929]), .SEL(N29), .F(
        \Data_Mem/n7855 ) );
  MUX \Data_Mem/U7888  ( .IN0(o[961]), .IN1(o[993]), .SEL(N29), .F(
        \Data_Mem/n7854 ) );
  MUX \Data_Mem/U7887  ( .IN0(\Data_Mem/n7852 ), .IN1(\Data_Mem/n7837 ), .SEL(
        N25), .F(\Data_Mem/n7853 ) );
  MUX \Data_Mem/U7886  ( .IN0(\Data_Mem/n7851 ), .IN1(\Data_Mem/n7844 ), .SEL(
        N26), .F(\Data_Mem/n7852 ) );
  MUX \Data_Mem/U7885  ( .IN0(\Data_Mem/n7850 ), .IN1(\Data_Mem/n7847 ), .SEL(
        N27), .F(\Data_Mem/n7851 ) );
  MUX \Data_Mem/U7884  ( .IN0(\Data_Mem/n7849 ), .IN1(\Data_Mem/n7848 ), .SEL(
        N28), .F(\Data_Mem/n7850 ) );
  MUX \Data_Mem/U7883  ( .IN0(o[1025]), .IN1(o[1057]), .SEL(N29), .F(
        \Data_Mem/n7849 ) );
  MUX \Data_Mem/U7882  ( .IN0(o[1089]), .IN1(o[1121]), .SEL(N29), .F(
        \Data_Mem/n7848 ) );
  MUX \Data_Mem/U7881  ( .IN0(\Data_Mem/n7846 ), .IN1(\Data_Mem/n7845 ), .SEL(
        N28), .F(\Data_Mem/n7847 ) );
  MUX \Data_Mem/U7880  ( .IN0(o[1153]), .IN1(o[1185]), .SEL(N29), .F(
        \Data_Mem/n7846 ) );
  MUX \Data_Mem/U7879  ( .IN0(o[1217]), .IN1(o[1249]), .SEL(N29), .F(
        \Data_Mem/n7845 ) );
  MUX \Data_Mem/U7878  ( .IN0(\Data_Mem/n7843 ), .IN1(\Data_Mem/n7840 ), .SEL(
        N27), .F(\Data_Mem/n7844 ) );
  MUX \Data_Mem/U7877  ( .IN0(\Data_Mem/n7842 ), .IN1(\Data_Mem/n7841 ), .SEL(
        N28), .F(\Data_Mem/n7843 ) );
  MUX \Data_Mem/U7876  ( .IN0(o[1281]), .IN1(o[1313]), .SEL(N29), .F(
        \Data_Mem/n7842 ) );
  MUX \Data_Mem/U7875  ( .IN0(o[1345]), .IN1(o[1377]), .SEL(N29), .F(
        \Data_Mem/n7841 ) );
  MUX \Data_Mem/U7874  ( .IN0(\Data_Mem/n7839 ), .IN1(\Data_Mem/n7838 ), .SEL(
        N28), .F(\Data_Mem/n7840 ) );
  MUX \Data_Mem/U7873  ( .IN0(o[1409]), .IN1(o[1441]), .SEL(N29), .F(
        \Data_Mem/n7839 ) );
  MUX \Data_Mem/U7872  ( .IN0(o[1473]), .IN1(o[1505]), .SEL(N29), .F(
        \Data_Mem/n7838 ) );
  MUX \Data_Mem/U7871  ( .IN0(\Data_Mem/n7836 ), .IN1(\Data_Mem/n7829 ), .SEL(
        N26), .F(\Data_Mem/n7837 ) );
  MUX \Data_Mem/U7870  ( .IN0(\Data_Mem/n7835 ), .IN1(\Data_Mem/n7832 ), .SEL(
        N27), .F(\Data_Mem/n7836 ) );
  MUX \Data_Mem/U7869  ( .IN0(\Data_Mem/n7834 ), .IN1(\Data_Mem/n7833 ), .SEL(
        N28), .F(\Data_Mem/n7835 ) );
  MUX \Data_Mem/U7868  ( .IN0(o[1537]), .IN1(o[1569]), .SEL(N29), .F(
        \Data_Mem/n7834 ) );
  MUX \Data_Mem/U7867  ( .IN0(o[1601]), .IN1(o[1633]), .SEL(N29), .F(
        \Data_Mem/n7833 ) );
  MUX \Data_Mem/U7866  ( .IN0(\Data_Mem/n7831 ), .IN1(\Data_Mem/n7830 ), .SEL(
        N28), .F(\Data_Mem/n7832 ) );
  MUX \Data_Mem/U7865  ( .IN0(o[1665]), .IN1(o[1697]), .SEL(N29), .F(
        \Data_Mem/n7831 ) );
  MUX \Data_Mem/U7864  ( .IN0(o[1729]), .IN1(o[1761]), .SEL(N29), .F(
        \Data_Mem/n7830 ) );
  MUX \Data_Mem/U7863  ( .IN0(\Data_Mem/n7828 ), .IN1(\Data_Mem/n7825 ), .SEL(
        N27), .F(\Data_Mem/n7829 ) );
  MUX \Data_Mem/U7862  ( .IN0(\Data_Mem/n7827 ), .IN1(\Data_Mem/n7826 ), .SEL(
        N28), .F(\Data_Mem/n7828 ) );
  MUX \Data_Mem/U7861  ( .IN0(o[1793]), .IN1(o[1825]), .SEL(N29), .F(
        \Data_Mem/n7827 ) );
  MUX \Data_Mem/U7860  ( .IN0(o[1857]), .IN1(o[1889]), .SEL(N29), .F(
        \Data_Mem/n7826 ) );
  MUX \Data_Mem/U7859  ( .IN0(\Data_Mem/n7824 ), .IN1(\Data_Mem/n7823 ), .SEL(
        N28), .F(\Data_Mem/n7825 ) );
  MUX \Data_Mem/U7858  ( .IN0(o[1921]), .IN1(o[1953]), .SEL(N29), .F(
        \Data_Mem/n7824 ) );
  MUX \Data_Mem/U7857  ( .IN0(o[1985]), .IN1(o[2017]), .SEL(N29), .F(
        \Data_Mem/n7823 ) );
  MUX \Data_Mem/U7856  ( .IN0(\Data_Mem/n7822 ), .IN1(\Data_Mem/n7791 ), .SEL(
        N24), .F(\Data_Mem/N745 ) );
  MUX \Data_Mem/U7855  ( .IN0(\Data_Mem/n7821 ), .IN1(\Data_Mem/n7806 ), .SEL(
        N25), .F(\Data_Mem/n7822 ) );
  MUX \Data_Mem/U7854  ( .IN0(\Data_Mem/n7820 ), .IN1(\Data_Mem/n7813 ), .SEL(
        N26), .F(\Data_Mem/n7821 ) );
  MUX \Data_Mem/U7853  ( .IN0(\Data_Mem/n7819 ), .IN1(\Data_Mem/n7816 ), .SEL(
        N27), .F(\Data_Mem/n7820 ) );
  MUX \Data_Mem/U7852  ( .IN0(\Data_Mem/n7818 ), .IN1(\Data_Mem/n7817 ), .SEL(
        N28), .F(\Data_Mem/n7819 ) );
  MUX \Data_Mem/U7851  ( .IN0(o[0]), .IN1(o[32]), .SEL(N29), .F(
        \Data_Mem/n7818 ) );
  MUX \Data_Mem/U7850  ( .IN0(o[64]), .IN1(o[96]), .SEL(N29), .F(
        \Data_Mem/n7817 ) );
  MUX \Data_Mem/U7849  ( .IN0(\Data_Mem/n7815 ), .IN1(\Data_Mem/n7814 ), .SEL(
        N28), .F(\Data_Mem/n7816 ) );
  MUX \Data_Mem/U7848  ( .IN0(o[128]), .IN1(o[160]), .SEL(N29), .F(
        \Data_Mem/n7815 ) );
  MUX \Data_Mem/U7847  ( .IN0(o[192]), .IN1(o[224]), .SEL(N29), .F(
        \Data_Mem/n7814 ) );
  MUX \Data_Mem/U7846  ( .IN0(\Data_Mem/n7812 ), .IN1(\Data_Mem/n7809 ), .SEL(
        N27), .F(\Data_Mem/n7813 ) );
  MUX \Data_Mem/U7845  ( .IN0(\Data_Mem/n7811 ), .IN1(\Data_Mem/n7810 ), .SEL(
        N28), .F(\Data_Mem/n7812 ) );
  MUX \Data_Mem/U7844  ( .IN0(o[256]), .IN1(o[288]), .SEL(N29), .F(
        \Data_Mem/n7811 ) );
  MUX \Data_Mem/U7843  ( .IN0(o[320]), .IN1(o[352]), .SEL(N29), .F(
        \Data_Mem/n7810 ) );
  MUX \Data_Mem/U7842  ( .IN0(\Data_Mem/n7808 ), .IN1(\Data_Mem/n7807 ), .SEL(
        N28), .F(\Data_Mem/n7809 ) );
  MUX \Data_Mem/U7841  ( .IN0(o[384]), .IN1(o[416]), .SEL(N29), .F(
        \Data_Mem/n7808 ) );
  MUX \Data_Mem/U7840  ( .IN0(o[448]), .IN1(o[480]), .SEL(N29), .F(
        \Data_Mem/n7807 ) );
  MUX \Data_Mem/U7839  ( .IN0(\Data_Mem/n7805 ), .IN1(\Data_Mem/n7798 ), .SEL(
        N26), .F(\Data_Mem/n7806 ) );
  MUX \Data_Mem/U7838  ( .IN0(\Data_Mem/n7804 ), .IN1(\Data_Mem/n7801 ), .SEL(
        N27), .F(\Data_Mem/n7805 ) );
  MUX \Data_Mem/U7837  ( .IN0(\Data_Mem/n7803 ), .IN1(\Data_Mem/n7802 ), .SEL(
        N28), .F(\Data_Mem/n7804 ) );
  MUX \Data_Mem/U7836  ( .IN0(o[512]), .IN1(o[544]), .SEL(N29), .F(
        \Data_Mem/n7803 ) );
  MUX \Data_Mem/U7835  ( .IN0(o[576]), .IN1(o[608]), .SEL(N29), .F(
        \Data_Mem/n7802 ) );
  MUX \Data_Mem/U7834  ( .IN0(\Data_Mem/n7800 ), .IN1(\Data_Mem/n7799 ), .SEL(
        N28), .F(\Data_Mem/n7801 ) );
  MUX \Data_Mem/U7833  ( .IN0(o[640]), .IN1(o[672]), .SEL(N29), .F(
        \Data_Mem/n7800 ) );
  MUX \Data_Mem/U7832  ( .IN0(o[704]), .IN1(o[736]), .SEL(N29), .F(
        \Data_Mem/n7799 ) );
  MUX \Data_Mem/U7831  ( .IN0(\Data_Mem/n7797 ), .IN1(\Data_Mem/n7794 ), .SEL(
        N27), .F(\Data_Mem/n7798 ) );
  MUX \Data_Mem/U7830  ( .IN0(\Data_Mem/n7796 ), .IN1(\Data_Mem/n7795 ), .SEL(
        N28), .F(\Data_Mem/n7797 ) );
  MUX \Data_Mem/U7829  ( .IN0(o[768]), .IN1(o[800]), .SEL(N29), .F(
        \Data_Mem/n7796 ) );
  MUX \Data_Mem/U7828  ( .IN0(o[832]), .IN1(o[864]), .SEL(N29), .F(
        \Data_Mem/n7795 ) );
  MUX \Data_Mem/U7827  ( .IN0(\Data_Mem/n7793 ), .IN1(\Data_Mem/n7792 ), .SEL(
        N28), .F(\Data_Mem/n7794 ) );
  MUX \Data_Mem/U7826  ( .IN0(o[896]), .IN1(o[928]), .SEL(N29), .F(
        \Data_Mem/n7793 ) );
  MUX \Data_Mem/U7825  ( .IN0(o[960]), .IN1(o[992]), .SEL(N29), .F(
        \Data_Mem/n7792 ) );
  MUX \Data_Mem/U7824  ( .IN0(\Data_Mem/n7790 ), .IN1(\Data_Mem/n7775 ), .SEL(
        N25), .F(\Data_Mem/n7791 ) );
  MUX \Data_Mem/U7823  ( .IN0(\Data_Mem/n7789 ), .IN1(\Data_Mem/n7782 ), .SEL(
        N26), .F(\Data_Mem/n7790 ) );
  MUX \Data_Mem/U7822  ( .IN0(\Data_Mem/n7788 ), .IN1(\Data_Mem/n7785 ), .SEL(
        N27), .F(\Data_Mem/n7789 ) );
  MUX \Data_Mem/U7821  ( .IN0(\Data_Mem/n7787 ), .IN1(\Data_Mem/n7786 ), .SEL(
        N28), .F(\Data_Mem/n7788 ) );
  MUX \Data_Mem/U7820  ( .IN0(o[1024]), .IN1(o[1056]), .SEL(N29), .F(
        \Data_Mem/n7787 ) );
  MUX \Data_Mem/U7819  ( .IN0(o[1088]), .IN1(o[1120]), .SEL(N29), .F(
        \Data_Mem/n7786 ) );
  MUX \Data_Mem/U7818  ( .IN0(\Data_Mem/n7784 ), .IN1(\Data_Mem/n7783 ), .SEL(
        N28), .F(\Data_Mem/n7785 ) );
  MUX \Data_Mem/U7817  ( .IN0(o[1152]), .IN1(o[1184]), .SEL(N29), .F(
        \Data_Mem/n7784 ) );
  MUX \Data_Mem/U7816  ( .IN0(o[1216]), .IN1(o[1248]), .SEL(N29), .F(
        \Data_Mem/n7783 ) );
  MUX \Data_Mem/U7815  ( .IN0(\Data_Mem/n7781 ), .IN1(\Data_Mem/n7778 ), .SEL(
        N27), .F(\Data_Mem/n7782 ) );
  MUX \Data_Mem/U7814  ( .IN0(\Data_Mem/n7780 ), .IN1(\Data_Mem/n7779 ), .SEL(
        N28), .F(\Data_Mem/n7781 ) );
  MUX \Data_Mem/U7813  ( .IN0(o[1280]), .IN1(o[1312]), .SEL(N29), .F(
        \Data_Mem/n7780 ) );
  MUX \Data_Mem/U7812  ( .IN0(o[1344]), .IN1(o[1376]), .SEL(N29), .F(
        \Data_Mem/n7779 ) );
  MUX \Data_Mem/U7811  ( .IN0(\Data_Mem/n7777 ), .IN1(\Data_Mem/n7776 ), .SEL(
        N28), .F(\Data_Mem/n7778 ) );
  MUX \Data_Mem/U7810  ( .IN0(o[1408]), .IN1(o[1440]), .SEL(N29), .F(
        \Data_Mem/n7777 ) );
  MUX \Data_Mem/U7809  ( .IN0(o[1472]), .IN1(o[1504]), .SEL(N29), .F(
        \Data_Mem/n7776 ) );
  MUX \Data_Mem/U7808  ( .IN0(\Data_Mem/n7774 ), .IN1(\Data_Mem/n7767 ), .SEL(
        N26), .F(\Data_Mem/n7775 ) );
  MUX \Data_Mem/U7807  ( .IN0(\Data_Mem/n7773 ), .IN1(\Data_Mem/n7770 ), .SEL(
        N27), .F(\Data_Mem/n7774 ) );
  MUX \Data_Mem/U7806  ( .IN0(\Data_Mem/n7772 ), .IN1(\Data_Mem/n7771 ), .SEL(
        N28), .F(\Data_Mem/n7773 ) );
  MUX \Data_Mem/U7805  ( .IN0(o[1536]), .IN1(o[1568]), .SEL(N29), .F(
        \Data_Mem/n7772 ) );
  MUX \Data_Mem/U7804  ( .IN0(o[1600]), .IN1(o[1632]), .SEL(N29), .F(
        \Data_Mem/n7771 ) );
  MUX \Data_Mem/U7803  ( .IN0(\Data_Mem/n7769 ), .IN1(\Data_Mem/n7768 ), .SEL(
        N28), .F(\Data_Mem/n7770 ) );
  MUX \Data_Mem/U7802  ( .IN0(o[1664]), .IN1(o[1696]), .SEL(N29), .F(
        \Data_Mem/n7769 ) );
  MUX \Data_Mem/U7801  ( .IN0(o[1728]), .IN1(o[1760]), .SEL(N29), .F(
        \Data_Mem/n7768 ) );
  MUX \Data_Mem/U7800  ( .IN0(\Data_Mem/n7766 ), .IN1(\Data_Mem/n7763 ), .SEL(
        N27), .F(\Data_Mem/n7767 ) );
  MUX \Data_Mem/U7799  ( .IN0(\Data_Mem/n7765 ), .IN1(\Data_Mem/n7764 ), .SEL(
        N28), .F(\Data_Mem/n7766 ) );
  MUX \Data_Mem/U7798  ( .IN0(o[1792]), .IN1(o[1824]), .SEL(N29), .F(
        \Data_Mem/n7765 ) );
  MUX \Data_Mem/U7797  ( .IN0(o[1856]), .IN1(o[1888]), .SEL(N29), .F(
        \Data_Mem/n7764 ) );
  MUX \Data_Mem/U7796  ( .IN0(\Data_Mem/n7762 ), .IN1(\Data_Mem/n7761 ), .SEL(
        N28), .F(\Data_Mem/n7763 ) );
  MUX \Data_Mem/U7795  ( .IN0(o[1920]), .IN1(o[1952]), .SEL(N29), .F(
        \Data_Mem/n7762 ) );
  MUX \Data_Mem/U7794  ( .IN0(o[1984]), .IN1(o[2016]), .SEL(N29), .F(
        \Data_Mem/n7761 ) );
  DFF \Data_Mem/memory_reg[63][0]  ( .D(\Data_Mem/n5713 ), .CLK(clk), .RST(rst), .I(e_init[2016]), .Q(o[2016]) );
  DFF \Data_Mem/memory_reg[63][1]  ( .D(\Data_Mem/n5714 ), .CLK(clk), .RST(rst), .I(e_init[2017]), .Q(o[2017]) );
  DFF \Data_Mem/memory_reg[63][2]  ( .D(\Data_Mem/n5715 ), .CLK(clk), .RST(rst), .I(e_init[2018]), .Q(o[2018]) );
  DFF \Data_Mem/memory_reg[63][3]  ( .D(\Data_Mem/n5716 ), .CLK(clk), .RST(rst), .I(e_init[2019]), .Q(o[2019]) );
  DFF \Data_Mem/memory_reg[63][4]  ( .D(\Data_Mem/n5717 ), .CLK(clk), .RST(rst), .I(e_init[2020]), .Q(o[2020]) );
  DFF \Data_Mem/memory_reg[63][5]  ( .D(\Data_Mem/n5718 ), .CLK(clk), .RST(rst), .I(e_init[2021]), .Q(o[2021]) );
  DFF \Data_Mem/memory_reg[63][6]  ( .D(\Data_Mem/n5719 ), .CLK(clk), .RST(rst), .I(e_init[2022]), .Q(o[2022]) );
  DFF \Data_Mem/memory_reg[63][7]  ( .D(\Data_Mem/n5720 ), .CLK(clk), .RST(rst), .I(e_init[2023]), .Q(o[2023]) );
  DFF \Data_Mem/memory_reg[63][8]  ( .D(\Data_Mem/n5721 ), .CLK(clk), .RST(rst), .I(e_init[2024]), .Q(o[2024]) );
  DFF \Data_Mem/memory_reg[63][9]  ( .D(\Data_Mem/n5722 ), .CLK(clk), .RST(rst), .I(e_init[2025]), .Q(o[2025]) );
  DFF \Data_Mem/memory_reg[63][10]  ( .D(\Data_Mem/n5723 ), .CLK(clk), .RST(
        rst), .I(e_init[2026]), .Q(o[2026]) );
  DFF \Data_Mem/memory_reg[63][11]  ( .D(\Data_Mem/n5724 ), .CLK(clk), .RST(
        rst), .I(e_init[2027]), .Q(o[2027]) );
  DFF \Data_Mem/memory_reg[63][12]  ( .D(\Data_Mem/n5725 ), .CLK(clk), .RST(
        rst), .I(e_init[2028]), .Q(o[2028]) );
  DFF \Data_Mem/memory_reg[63][13]  ( .D(\Data_Mem/n5726 ), .CLK(clk), .RST(
        rst), .I(e_init[2029]), .Q(o[2029]) );
  DFF \Data_Mem/memory_reg[63][14]  ( .D(\Data_Mem/n5727 ), .CLK(clk), .RST(
        rst), .I(e_init[2030]), .Q(o[2030]) );
  DFF \Data_Mem/memory_reg[63][15]  ( .D(\Data_Mem/n5728 ), .CLK(clk), .RST(
        rst), .I(e_init[2031]), .Q(o[2031]) );
  DFF \Data_Mem/memory_reg[63][16]  ( .D(\Data_Mem/n5729 ), .CLK(clk), .RST(
        rst), .I(e_init[2032]), .Q(o[2032]) );
  DFF \Data_Mem/memory_reg[63][17]  ( .D(\Data_Mem/n5730 ), .CLK(clk), .RST(
        rst), .I(e_init[2033]), .Q(o[2033]) );
  DFF \Data_Mem/memory_reg[63][18]  ( .D(\Data_Mem/n5731 ), .CLK(clk), .RST(
        rst), .I(e_init[2034]), .Q(o[2034]) );
  DFF \Data_Mem/memory_reg[63][19]  ( .D(\Data_Mem/n5732 ), .CLK(clk), .RST(
        rst), .I(e_init[2035]), .Q(o[2035]) );
  DFF \Data_Mem/memory_reg[63][20]  ( .D(\Data_Mem/n5733 ), .CLK(clk), .RST(
        rst), .I(e_init[2036]), .Q(o[2036]) );
  DFF \Data_Mem/memory_reg[63][21]  ( .D(\Data_Mem/n5734 ), .CLK(clk), .RST(
        rst), .I(e_init[2037]), .Q(o[2037]) );
  DFF \Data_Mem/memory_reg[63][22]  ( .D(\Data_Mem/n5735 ), .CLK(clk), .RST(
        rst), .I(e_init[2038]), .Q(o[2038]) );
  DFF \Data_Mem/memory_reg[63][23]  ( .D(\Data_Mem/n5736 ), .CLK(clk), .RST(
        rst), .I(e_init[2039]), .Q(o[2039]) );
  DFF \Data_Mem/memory_reg[63][24]  ( .D(\Data_Mem/n5737 ), .CLK(clk), .RST(
        rst), .I(e_init[2040]), .Q(o[2040]) );
  DFF \Data_Mem/memory_reg[63][25]  ( .D(\Data_Mem/n5738 ), .CLK(clk), .RST(
        rst), .I(e_init[2041]), .Q(o[2041]) );
  DFF \Data_Mem/memory_reg[63][26]  ( .D(\Data_Mem/n5739 ), .CLK(clk), .RST(
        rst), .I(e_init[2042]), .Q(o[2042]) );
  DFF \Data_Mem/memory_reg[63][27]  ( .D(\Data_Mem/n5740 ), .CLK(clk), .RST(
        rst), .I(e_init[2043]), .Q(o[2043]) );
  DFF \Data_Mem/memory_reg[63][28]  ( .D(\Data_Mem/n5741 ), .CLK(clk), .RST(
        rst), .I(e_init[2044]), .Q(o[2044]) );
  DFF \Data_Mem/memory_reg[63][29]  ( .D(\Data_Mem/n5742 ), .CLK(clk), .RST(
        rst), .I(e_init[2045]), .Q(o[2045]) );
  DFF \Data_Mem/memory_reg[63][30]  ( .D(\Data_Mem/n5743 ), .CLK(clk), .RST(
        rst), .I(e_init[2046]), .Q(o[2046]) );
  DFF \Data_Mem/memory_reg[63][31]  ( .D(\Data_Mem/n5744 ), .CLK(clk), .RST(
        rst), .I(e_init[2047]), .Q(o[2047]) );
  DFF \Data_Mem/memory_reg[62][0]  ( .D(\Data_Mem/n5745 ), .CLK(clk), .RST(rst), .I(e_init[1984]), .Q(o[1984]) );
  DFF \Data_Mem/memory_reg[62][1]  ( .D(\Data_Mem/n5746 ), .CLK(clk), .RST(rst), .I(e_init[1985]), .Q(o[1985]) );
  DFF \Data_Mem/memory_reg[62][2]  ( .D(\Data_Mem/n5747 ), .CLK(clk), .RST(rst), .I(e_init[1986]), .Q(o[1986]) );
  DFF \Data_Mem/memory_reg[62][3]  ( .D(\Data_Mem/n5748 ), .CLK(clk), .RST(rst), .I(e_init[1987]), .Q(o[1987]) );
  DFF \Data_Mem/memory_reg[62][4]  ( .D(\Data_Mem/n5749 ), .CLK(clk), .RST(rst), .I(e_init[1988]), .Q(o[1988]) );
  DFF \Data_Mem/memory_reg[62][5]  ( .D(\Data_Mem/n5750 ), .CLK(clk), .RST(rst), .I(e_init[1989]), .Q(o[1989]) );
  DFF \Data_Mem/memory_reg[62][6]  ( .D(\Data_Mem/n5751 ), .CLK(clk), .RST(rst), .I(e_init[1990]), .Q(o[1990]) );
  DFF \Data_Mem/memory_reg[62][7]  ( .D(\Data_Mem/n5752 ), .CLK(clk), .RST(rst), .I(e_init[1991]), .Q(o[1991]) );
  DFF \Data_Mem/memory_reg[62][8]  ( .D(\Data_Mem/n5753 ), .CLK(clk), .RST(rst), .I(e_init[1992]), .Q(o[1992]) );
  DFF \Data_Mem/memory_reg[62][9]  ( .D(\Data_Mem/n5754 ), .CLK(clk), .RST(rst), .I(e_init[1993]), .Q(o[1993]) );
  DFF \Data_Mem/memory_reg[62][10]  ( .D(\Data_Mem/n5755 ), .CLK(clk), .RST(
        rst), .I(e_init[1994]), .Q(o[1994]) );
  DFF \Data_Mem/memory_reg[62][11]  ( .D(\Data_Mem/n5756 ), .CLK(clk), .RST(
        rst), .I(e_init[1995]), .Q(o[1995]) );
  DFF \Data_Mem/memory_reg[62][12]  ( .D(\Data_Mem/n5757 ), .CLK(clk), .RST(
        rst), .I(e_init[1996]), .Q(o[1996]) );
  DFF \Data_Mem/memory_reg[62][13]  ( .D(\Data_Mem/n5758 ), .CLK(clk), .RST(
        rst), .I(e_init[1997]), .Q(o[1997]) );
  DFF \Data_Mem/memory_reg[62][14]  ( .D(\Data_Mem/n5759 ), .CLK(clk), .RST(
        rst), .I(e_init[1998]), .Q(o[1998]) );
  DFF \Data_Mem/memory_reg[62][15]  ( .D(\Data_Mem/n5760 ), .CLK(clk), .RST(
        rst), .I(e_init[1999]), .Q(o[1999]) );
  DFF \Data_Mem/memory_reg[62][16]  ( .D(\Data_Mem/n5761 ), .CLK(clk), .RST(
        rst), .I(e_init[2000]), .Q(o[2000]) );
  DFF \Data_Mem/memory_reg[62][17]  ( .D(\Data_Mem/n5762 ), .CLK(clk), .RST(
        rst), .I(e_init[2001]), .Q(o[2001]) );
  DFF \Data_Mem/memory_reg[62][18]  ( .D(\Data_Mem/n5763 ), .CLK(clk), .RST(
        rst), .I(e_init[2002]), .Q(o[2002]) );
  DFF \Data_Mem/memory_reg[62][19]  ( .D(\Data_Mem/n5764 ), .CLK(clk), .RST(
        rst), .I(e_init[2003]), .Q(o[2003]) );
  DFF \Data_Mem/memory_reg[62][20]  ( .D(\Data_Mem/n5765 ), .CLK(clk), .RST(
        rst), .I(e_init[2004]), .Q(o[2004]) );
  DFF \Data_Mem/memory_reg[62][21]  ( .D(\Data_Mem/n5766 ), .CLK(clk), .RST(
        rst), .I(e_init[2005]), .Q(o[2005]) );
  DFF \Data_Mem/memory_reg[62][22]  ( .D(\Data_Mem/n5767 ), .CLK(clk), .RST(
        rst), .I(e_init[2006]), .Q(o[2006]) );
  DFF \Data_Mem/memory_reg[62][23]  ( .D(\Data_Mem/n5768 ), .CLK(clk), .RST(
        rst), .I(e_init[2007]), .Q(o[2007]) );
  DFF \Data_Mem/memory_reg[62][24]  ( .D(\Data_Mem/n5769 ), .CLK(clk), .RST(
        rst), .I(e_init[2008]), .Q(o[2008]) );
  DFF \Data_Mem/memory_reg[62][25]  ( .D(\Data_Mem/n5770 ), .CLK(clk), .RST(
        rst), .I(e_init[2009]), .Q(o[2009]) );
  DFF \Data_Mem/memory_reg[62][26]  ( .D(\Data_Mem/n5771 ), .CLK(clk), .RST(
        rst), .I(e_init[2010]), .Q(o[2010]) );
  DFF \Data_Mem/memory_reg[62][27]  ( .D(\Data_Mem/n5772 ), .CLK(clk), .RST(
        rst), .I(e_init[2011]), .Q(o[2011]) );
  DFF \Data_Mem/memory_reg[62][28]  ( .D(\Data_Mem/n5773 ), .CLK(clk), .RST(
        rst), .I(e_init[2012]), .Q(o[2012]) );
  DFF \Data_Mem/memory_reg[62][29]  ( .D(\Data_Mem/n5774 ), .CLK(clk), .RST(
        rst), .I(e_init[2013]), .Q(o[2013]) );
  DFF \Data_Mem/memory_reg[62][30]  ( .D(\Data_Mem/n5775 ), .CLK(clk), .RST(
        rst), .I(e_init[2014]), .Q(o[2014]) );
  DFF \Data_Mem/memory_reg[62][31]  ( .D(\Data_Mem/n5776 ), .CLK(clk), .RST(
        rst), .I(e_init[2015]), .Q(o[2015]) );
  DFF \Data_Mem/memory_reg[61][0]  ( .D(\Data_Mem/n5777 ), .CLK(clk), .RST(rst), .I(e_init[1952]), .Q(o[1952]) );
  DFF \Data_Mem/memory_reg[61][1]  ( .D(\Data_Mem/n5778 ), .CLK(clk), .RST(rst), .I(e_init[1953]), .Q(o[1953]) );
  DFF \Data_Mem/memory_reg[61][2]  ( .D(\Data_Mem/n5779 ), .CLK(clk), .RST(rst), .I(e_init[1954]), .Q(o[1954]) );
  DFF \Data_Mem/memory_reg[61][3]  ( .D(\Data_Mem/n5780 ), .CLK(clk), .RST(rst), .I(e_init[1955]), .Q(o[1955]) );
  DFF \Data_Mem/memory_reg[61][4]  ( .D(\Data_Mem/n5781 ), .CLK(clk), .RST(rst), .I(e_init[1956]), .Q(o[1956]) );
  DFF \Data_Mem/memory_reg[61][5]  ( .D(\Data_Mem/n5782 ), .CLK(clk), .RST(rst), .I(e_init[1957]), .Q(o[1957]) );
  DFF \Data_Mem/memory_reg[61][6]  ( .D(\Data_Mem/n5783 ), .CLK(clk), .RST(rst), .I(e_init[1958]), .Q(o[1958]) );
  DFF \Data_Mem/memory_reg[61][7]  ( .D(\Data_Mem/n5784 ), .CLK(clk), .RST(rst), .I(e_init[1959]), .Q(o[1959]) );
  DFF \Data_Mem/memory_reg[61][8]  ( .D(\Data_Mem/n5785 ), .CLK(clk), .RST(rst), .I(e_init[1960]), .Q(o[1960]) );
  DFF \Data_Mem/memory_reg[61][9]  ( .D(\Data_Mem/n5786 ), .CLK(clk), .RST(rst), .I(e_init[1961]), .Q(o[1961]) );
  DFF \Data_Mem/memory_reg[61][10]  ( .D(\Data_Mem/n5787 ), .CLK(clk), .RST(
        rst), .I(e_init[1962]), .Q(o[1962]) );
  DFF \Data_Mem/memory_reg[61][11]  ( .D(\Data_Mem/n5788 ), .CLK(clk), .RST(
        rst), .I(e_init[1963]), .Q(o[1963]) );
  DFF \Data_Mem/memory_reg[61][12]  ( .D(\Data_Mem/n5789 ), .CLK(clk), .RST(
        rst), .I(e_init[1964]), .Q(o[1964]) );
  DFF \Data_Mem/memory_reg[61][13]  ( .D(\Data_Mem/n5790 ), .CLK(clk), .RST(
        rst), .I(e_init[1965]), .Q(o[1965]) );
  DFF \Data_Mem/memory_reg[61][14]  ( .D(\Data_Mem/n5791 ), .CLK(clk), .RST(
        rst), .I(e_init[1966]), .Q(o[1966]) );
  DFF \Data_Mem/memory_reg[61][15]  ( .D(\Data_Mem/n5792 ), .CLK(clk), .RST(
        rst), .I(e_init[1967]), .Q(o[1967]) );
  DFF \Data_Mem/memory_reg[61][16]  ( .D(\Data_Mem/n5793 ), .CLK(clk), .RST(
        rst), .I(e_init[1968]), .Q(o[1968]) );
  DFF \Data_Mem/memory_reg[61][17]  ( .D(\Data_Mem/n5794 ), .CLK(clk), .RST(
        rst), .I(e_init[1969]), .Q(o[1969]) );
  DFF \Data_Mem/memory_reg[61][18]  ( .D(\Data_Mem/n5795 ), .CLK(clk), .RST(
        rst), .I(e_init[1970]), .Q(o[1970]) );
  DFF \Data_Mem/memory_reg[61][19]  ( .D(\Data_Mem/n5796 ), .CLK(clk), .RST(
        rst), .I(e_init[1971]), .Q(o[1971]) );
  DFF \Data_Mem/memory_reg[61][20]  ( .D(\Data_Mem/n5797 ), .CLK(clk), .RST(
        rst), .I(e_init[1972]), .Q(o[1972]) );
  DFF \Data_Mem/memory_reg[61][21]  ( .D(\Data_Mem/n5798 ), .CLK(clk), .RST(
        rst), .I(e_init[1973]), .Q(o[1973]) );
  DFF \Data_Mem/memory_reg[61][22]  ( .D(\Data_Mem/n5799 ), .CLK(clk), .RST(
        rst), .I(e_init[1974]), .Q(o[1974]) );
  DFF \Data_Mem/memory_reg[61][23]  ( .D(\Data_Mem/n5800 ), .CLK(clk), .RST(
        rst), .I(e_init[1975]), .Q(o[1975]) );
  DFF \Data_Mem/memory_reg[61][24]  ( .D(\Data_Mem/n5801 ), .CLK(clk), .RST(
        rst), .I(e_init[1976]), .Q(o[1976]) );
  DFF \Data_Mem/memory_reg[61][25]  ( .D(\Data_Mem/n5802 ), .CLK(clk), .RST(
        rst), .I(e_init[1977]), .Q(o[1977]) );
  DFF \Data_Mem/memory_reg[61][26]  ( .D(\Data_Mem/n5803 ), .CLK(clk), .RST(
        rst), .I(e_init[1978]), .Q(o[1978]) );
  DFF \Data_Mem/memory_reg[61][27]  ( .D(\Data_Mem/n5804 ), .CLK(clk), .RST(
        rst), .I(e_init[1979]), .Q(o[1979]) );
  DFF \Data_Mem/memory_reg[61][28]  ( .D(\Data_Mem/n5805 ), .CLK(clk), .RST(
        rst), .I(e_init[1980]), .Q(o[1980]) );
  DFF \Data_Mem/memory_reg[61][29]  ( .D(\Data_Mem/n5806 ), .CLK(clk), .RST(
        rst), .I(e_init[1981]), .Q(o[1981]) );
  DFF \Data_Mem/memory_reg[61][30]  ( .D(\Data_Mem/n5807 ), .CLK(clk), .RST(
        rst), .I(e_init[1982]), .Q(o[1982]) );
  DFF \Data_Mem/memory_reg[61][31]  ( .D(\Data_Mem/n5808 ), .CLK(clk), .RST(
        rst), .I(e_init[1983]), .Q(o[1983]) );
  DFF \Data_Mem/memory_reg[60][0]  ( .D(\Data_Mem/n5809 ), .CLK(clk), .RST(rst), .I(e_init[1920]), .Q(o[1920]) );
  DFF \Data_Mem/memory_reg[60][1]  ( .D(\Data_Mem/n5810 ), .CLK(clk), .RST(rst), .I(e_init[1921]), .Q(o[1921]) );
  DFF \Data_Mem/memory_reg[60][2]  ( .D(\Data_Mem/n5811 ), .CLK(clk), .RST(rst), .I(e_init[1922]), .Q(o[1922]) );
  DFF \Data_Mem/memory_reg[60][3]  ( .D(\Data_Mem/n5812 ), .CLK(clk), .RST(rst), .I(e_init[1923]), .Q(o[1923]) );
  DFF \Data_Mem/memory_reg[60][4]  ( .D(\Data_Mem/n5813 ), .CLK(clk), .RST(rst), .I(e_init[1924]), .Q(o[1924]) );
  DFF \Data_Mem/memory_reg[60][5]  ( .D(\Data_Mem/n5814 ), .CLK(clk), .RST(rst), .I(e_init[1925]), .Q(o[1925]) );
  DFF \Data_Mem/memory_reg[60][6]  ( .D(\Data_Mem/n5815 ), .CLK(clk), .RST(rst), .I(e_init[1926]), .Q(o[1926]) );
  DFF \Data_Mem/memory_reg[60][7]  ( .D(\Data_Mem/n5816 ), .CLK(clk), .RST(rst), .I(e_init[1927]), .Q(o[1927]) );
  DFF \Data_Mem/memory_reg[60][8]  ( .D(\Data_Mem/n5817 ), .CLK(clk), .RST(rst), .I(e_init[1928]), .Q(o[1928]) );
  DFF \Data_Mem/memory_reg[60][9]  ( .D(\Data_Mem/n5818 ), .CLK(clk), .RST(rst), .I(e_init[1929]), .Q(o[1929]) );
  DFF \Data_Mem/memory_reg[60][10]  ( .D(\Data_Mem/n5819 ), .CLK(clk), .RST(
        rst), .I(e_init[1930]), .Q(o[1930]) );
  DFF \Data_Mem/memory_reg[60][11]  ( .D(\Data_Mem/n5820 ), .CLK(clk), .RST(
        rst), .I(e_init[1931]), .Q(o[1931]) );
  DFF \Data_Mem/memory_reg[60][12]  ( .D(\Data_Mem/n5821 ), .CLK(clk), .RST(
        rst), .I(e_init[1932]), .Q(o[1932]) );
  DFF \Data_Mem/memory_reg[60][13]  ( .D(\Data_Mem/n5822 ), .CLK(clk), .RST(
        rst), .I(e_init[1933]), .Q(o[1933]) );
  DFF \Data_Mem/memory_reg[60][14]  ( .D(\Data_Mem/n5823 ), .CLK(clk), .RST(
        rst), .I(e_init[1934]), .Q(o[1934]) );
  DFF \Data_Mem/memory_reg[60][15]  ( .D(\Data_Mem/n5824 ), .CLK(clk), .RST(
        rst), .I(e_init[1935]), .Q(o[1935]) );
  DFF \Data_Mem/memory_reg[60][16]  ( .D(\Data_Mem/n5825 ), .CLK(clk), .RST(
        rst), .I(e_init[1936]), .Q(o[1936]) );
  DFF \Data_Mem/memory_reg[60][17]  ( .D(\Data_Mem/n5826 ), .CLK(clk), .RST(
        rst), .I(e_init[1937]), .Q(o[1937]) );
  DFF \Data_Mem/memory_reg[60][18]  ( .D(\Data_Mem/n5827 ), .CLK(clk), .RST(
        rst), .I(e_init[1938]), .Q(o[1938]) );
  DFF \Data_Mem/memory_reg[60][19]  ( .D(\Data_Mem/n5828 ), .CLK(clk), .RST(
        rst), .I(e_init[1939]), .Q(o[1939]) );
  DFF \Data_Mem/memory_reg[60][20]  ( .D(\Data_Mem/n5829 ), .CLK(clk), .RST(
        rst), .I(e_init[1940]), .Q(o[1940]) );
  DFF \Data_Mem/memory_reg[60][21]  ( .D(\Data_Mem/n5830 ), .CLK(clk), .RST(
        rst), .I(e_init[1941]), .Q(o[1941]) );
  DFF \Data_Mem/memory_reg[60][22]  ( .D(\Data_Mem/n5831 ), .CLK(clk), .RST(
        rst), .I(e_init[1942]), .Q(o[1942]) );
  DFF \Data_Mem/memory_reg[60][23]  ( .D(\Data_Mem/n5832 ), .CLK(clk), .RST(
        rst), .I(e_init[1943]), .Q(o[1943]) );
  DFF \Data_Mem/memory_reg[60][24]  ( .D(\Data_Mem/n5833 ), .CLK(clk), .RST(
        rst), .I(e_init[1944]), .Q(o[1944]) );
  DFF \Data_Mem/memory_reg[60][25]  ( .D(\Data_Mem/n5834 ), .CLK(clk), .RST(
        rst), .I(e_init[1945]), .Q(o[1945]) );
  DFF \Data_Mem/memory_reg[60][26]  ( .D(\Data_Mem/n5835 ), .CLK(clk), .RST(
        rst), .I(e_init[1946]), .Q(o[1946]) );
  DFF \Data_Mem/memory_reg[60][27]  ( .D(\Data_Mem/n5836 ), .CLK(clk), .RST(
        rst), .I(e_init[1947]), .Q(o[1947]) );
  DFF \Data_Mem/memory_reg[60][28]  ( .D(\Data_Mem/n5837 ), .CLK(clk), .RST(
        rst), .I(e_init[1948]), .Q(o[1948]) );
  DFF \Data_Mem/memory_reg[60][29]  ( .D(\Data_Mem/n5838 ), .CLK(clk), .RST(
        rst), .I(e_init[1949]), .Q(o[1949]) );
  DFF \Data_Mem/memory_reg[60][30]  ( .D(\Data_Mem/n5839 ), .CLK(clk), .RST(
        rst), .I(e_init[1950]), .Q(o[1950]) );
  DFF \Data_Mem/memory_reg[60][31]  ( .D(\Data_Mem/n5840 ), .CLK(clk), .RST(
        rst), .I(e_init[1951]), .Q(o[1951]) );
  DFF \Data_Mem/memory_reg[59][0]  ( .D(\Data_Mem/n5841 ), .CLK(clk), .RST(rst), .I(e_init[1888]), .Q(o[1888]) );
  DFF \Data_Mem/memory_reg[59][1]  ( .D(\Data_Mem/n5842 ), .CLK(clk), .RST(rst), .I(e_init[1889]), .Q(o[1889]) );
  DFF \Data_Mem/memory_reg[59][2]  ( .D(\Data_Mem/n5843 ), .CLK(clk), .RST(rst), .I(e_init[1890]), .Q(o[1890]) );
  DFF \Data_Mem/memory_reg[59][3]  ( .D(\Data_Mem/n5844 ), .CLK(clk), .RST(rst), .I(e_init[1891]), .Q(o[1891]) );
  DFF \Data_Mem/memory_reg[59][4]  ( .D(\Data_Mem/n5845 ), .CLK(clk), .RST(rst), .I(e_init[1892]), .Q(o[1892]) );
  DFF \Data_Mem/memory_reg[59][5]  ( .D(\Data_Mem/n5846 ), .CLK(clk), .RST(rst), .I(e_init[1893]), .Q(o[1893]) );
  DFF \Data_Mem/memory_reg[59][6]  ( .D(\Data_Mem/n5847 ), .CLK(clk), .RST(rst), .I(e_init[1894]), .Q(o[1894]) );
  DFF \Data_Mem/memory_reg[59][7]  ( .D(\Data_Mem/n5848 ), .CLK(clk), .RST(rst), .I(e_init[1895]), .Q(o[1895]) );
  DFF \Data_Mem/memory_reg[59][8]  ( .D(\Data_Mem/n5849 ), .CLK(clk), .RST(rst), .I(e_init[1896]), .Q(o[1896]) );
  DFF \Data_Mem/memory_reg[59][9]  ( .D(\Data_Mem/n5850 ), .CLK(clk), .RST(rst), .I(e_init[1897]), .Q(o[1897]) );
  DFF \Data_Mem/memory_reg[59][10]  ( .D(\Data_Mem/n5851 ), .CLK(clk), .RST(
        rst), .I(e_init[1898]), .Q(o[1898]) );
  DFF \Data_Mem/memory_reg[59][11]  ( .D(\Data_Mem/n5852 ), .CLK(clk), .RST(
        rst), .I(e_init[1899]), .Q(o[1899]) );
  DFF \Data_Mem/memory_reg[59][12]  ( .D(\Data_Mem/n5853 ), .CLK(clk), .RST(
        rst), .I(e_init[1900]), .Q(o[1900]) );
  DFF \Data_Mem/memory_reg[59][13]  ( .D(\Data_Mem/n5854 ), .CLK(clk), .RST(
        rst), .I(e_init[1901]), .Q(o[1901]) );
  DFF \Data_Mem/memory_reg[59][14]  ( .D(\Data_Mem/n5855 ), .CLK(clk), .RST(
        rst), .I(e_init[1902]), .Q(o[1902]) );
  DFF \Data_Mem/memory_reg[59][15]  ( .D(\Data_Mem/n5856 ), .CLK(clk), .RST(
        rst), .I(e_init[1903]), .Q(o[1903]) );
  DFF \Data_Mem/memory_reg[59][16]  ( .D(\Data_Mem/n5857 ), .CLK(clk), .RST(
        rst), .I(e_init[1904]), .Q(o[1904]) );
  DFF \Data_Mem/memory_reg[59][17]  ( .D(\Data_Mem/n5858 ), .CLK(clk), .RST(
        rst), .I(e_init[1905]), .Q(o[1905]) );
  DFF \Data_Mem/memory_reg[59][18]  ( .D(\Data_Mem/n5859 ), .CLK(clk), .RST(
        rst), .I(e_init[1906]), .Q(o[1906]) );
  DFF \Data_Mem/memory_reg[59][19]  ( .D(\Data_Mem/n5860 ), .CLK(clk), .RST(
        rst), .I(e_init[1907]), .Q(o[1907]) );
  DFF \Data_Mem/memory_reg[59][20]  ( .D(\Data_Mem/n5861 ), .CLK(clk), .RST(
        rst), .I(e_init[1908]), .Q(o[1908]) );
  DFF \Data_Mem/memory_reg[59][21]  ( .D(\Data_Mem/n5862 ), .CLK(clk), .RST(
        rst), .I(e_init[1909]), .Q(o[1909]) );
  DFF \Data_Mem/memory_reg[59][22]  ( .D(\Data_Mem/n5863 ), .CLK(clk), .RST(
        rst), .I(e_init[1910]), .Q(o[1910]) );
  DFF \Data_Mem/memory_reg[59][23]  ( .D(\Data_Mem/n5864 ), .CLK(clk), .RST(
        rst), .I(e_init[1911]), .Q(o[1911]) );
  DFF \Data_Mem/memory_reg[59][24]  ( .D(\Data_Mem/n5865 ), .CLK(clk), .RST(
        rst), .I(e_init[1912]), .Q(o[1912]) );
  DFF \Data_Mem/memory_reg[59][25]  ( .D(\Data_Mem/n5866 ), .CLK(clk), .RST(
        rst), .I(e_init[1913]), .Q(o[1913]) );
  DFF \Data_Mem/memory_reg[59][26]  ( .D(\Data_Mem/n5867 ), .CLK(clk), .RST(
        rst), .I(e_init[1914]), .Q(o[1914]) );
  DFF \Data_Mem/memory_reg[59][27]  ( .D(\Data_Mem/n5868 ), .CLK(clk), .RST(
        rst), .I(e_init[1915]), .Q(o[1915]) );
  DFF \Data_Mem/memory_reg[59][28]  ( .D(\Data_Mem/n5869 ), .CLK(clk), .RST(
        rst), .I(e_init[1916]), .Q(o[1916]) );
  DFF \Data_Mem/memory_reg[59][29]  ( .D(\Data_Mem/n5870 ), .CLK(clk), .RST(
        rst), .I(e_init[1917]), .Q(o[1917]) );
  DFF \Data_Mem/memory_reg[59][30]  ( .D(\Data_Mem/n5871 ), .CLK(clk), .RST(
        rst), .I(e_init[1918]), .Q(o[1918]) );
  DFF \Data_Mem/memory_reg[59][31]  ( .D(\Data_Mem/n5872 ), .CLK(clk), .RST(
        rst), .I(e_init[1919]), .Q(o[1919]) );
  DFF \Data_Mem/memory_reg[58][0]  ( .D(\Data_Mem/n5873 ), .CLK(clk), .RST(rst), .I(e_init[1856]), .Q(o[1856]) );
  DFF \Data_Mem/memory_reg[58][1]  ( .D(\Data_Mem/n5874 ), .CLK(clk), .RST(rst), .I(e_init[1857]), .Q(o[1857]) );
  DFF \Data_Mem/memory_reg[58][2]  ( .D(\Data_Mem/n5875 ), .CLK(clk), .RST(rst), .I(e_init[1858]), .Q(o[1858]) );
  DFF \Data_Mem/memory_reg[58][3]  ( .D(\Data_Mem/n5876 ), .CLK(clk), .RST(rst), .I(e_init[1859]), .Q(o[1859]) );
  DFF \Data_Mem/memory_reg[58][4]  ( .D(\Data_Mem/n5877 ), .CLK(clk), .RST(rst), .I(e_init[1860]), .Q(o[1860]) );
  DFF \Data_Mem/memory_reg[58][5]  ( .D(\Data_Mem/n5878 ), .CLK(clk), .RST(rst), .I(e_init[1861]), .Q(o[1861]) );
  DFF \Data_Mem/memory_reg[58][6]  ( .D(\Data_Mem/n5879 ), .CLK(clk), .RST(rst), .I(e_init[1862]), .Q(o[1862]) );
  DFF \Data_Mem/memory_reg[58][7]  ( .D(\Data_Mem/n5880 ), .CLK(clk), .RST(rst), .I(e_init[1863]), .Q(o[1863]) );
  DFF \Data_Mem/memory_reg[58][8]  ( .D(\Data_Mem/n5881 ), .CLK(clk), .RST(rst), .I(e_init[1864]), .Q(o[1864]) );
  DFF \Data_Mem/memory_reg[58][9]  ( .D(\Data_Mem/n5882 ), .CLK(clk), .RST(rst), .I(e_init[1865]), .Q(o[1865]) );
  DFF \Data_Mem/memory_reg[58][10]  ( .D(\Data_Mem/n5883 ), .CLK(clk), .RST(
        rst), .I(e_init[1866]), .Q(o[1866]) );
  DFF \Data_Mem/memory_reg[58][11]  ( .D(\Data_Mem/n5884 ), .CLK(clk), .RST(
        rst), .I(e_init[1867]), .Q(o[1867]) );
  DFF \Data_Mem/memory_reg[58][12]  ( .D(\Data_Mem/n5885 ), .CLK(clk), .RST(
        rst), .I(e_init[1868]), .Q(o[1868]) );
  DFF \Data_Mem/memory_reg[58][13]  ( .D(\Data_Mem/n5886 ), .CLK(clk), .RST(
        rst), .I(e_init[1869]), .Q(o[1869]) );
  DFF \Data_Mem/memory_reg[58][14]  ( .D(\Data_Mem/n5887 ), .CLK(clk), .RST(
        rst), .I(e_init[1870]), .Q(o[1870]) );
  DFF \Data_Mem/memory_reg[58][15]  ( .D(\Data_Mem/n5888 ), .CLK(clk), .RST(
        rst), .I(e_init[1871]), .Q(o[1871]) );
  DFF \Data_Mem/memory_reg[58][16]  ( .D(\Data_Mem/n5889 ), .CLK(clk), .RST(
        rst), .I(e_init[1872]), .Q(o[1872]) );
  DFF \Data_Mem/memory_reg[58][17]  ( .D(\Data_Mem/n5890 ), .CLK(clk), .RST(
        rst), .I(e_init[1873]), .Q(o[1873]) );
  DFF \Data_Mem/memory_reg[58][18]  ( .D(\Data_Mem/n5891 ), .CLK(clk), .RST(
        rst), .I(e_init[1874]), .Q(o[1874]) );
  DFF \Data_Mem/memory_reg[58][19]  ( .D(\Data_Mem/n5892 ), .CLK(clk), .RST(
        rst), .I(e_init[1875]), .Q(o[1875]) );
  DFF \Data_Mem/memory_reg[58][20]  ( .D(\Data_Mem/n5893 ), .CLK(clk), .RST(
        rst), .I(e_init[1876]), .Q(o[1876]) );
  DFF \Data_Mem/memory_reg[58][21]  ( .D(\Data_Mem/n5894 ), .CLK(clk), .RST(
        rst), .I(e_init[1877]), .Q(o[1877]) );
  DFF \Data_Mem/memory_reg[58][22]  ( .D(\Data_Mem/n5895 ), .CLK(clk), .RST(
        rst), .I(e_init[1878]), .Q(o[1878]) );
  DFF \Data_Mem/memory_reg[58][23]  ( .D(\Data_Mem/n5896 ), .CLK(clk), .RST(
        rst), .I(e_init[1879]), .Q(o[1879]) );
  DFF \Data_Mem/memory_reg[58][24]  ( .D(\Data_Mem/n5897 ), .CLK(clk), .RST(
        rst), .I(e_init[1880]), .Q(o[1880]) );
  DFF \Data_Mem/memory_reg[58][25]  ( .D(\Data_Mem/n5898 ), .CLK(clk), .RST(
        rst), .I(e_init[1881]), .Q(o[1881]) );
  DFF \Data_Mem/memory_reg[58][26]  ( .D(\Data_Mem/n5899 ), .CLK(clk), .RST(
        rst), .I(e_init[1882]), .Q(o[1882]) );
  DFF \Data_Mem/memory_reg[58][27]  ( .D(\Data_Mem/n5900 ), .CLK(clk), .RST(
        rst), .I(e_init[1883]), .Q(o[1883]) );
  DFF \Data_Mem/memory_reg[58][28]  ( .D(\Data_Mem/n5901 ), .CLK(clk), .RST(
        rst), .I(e_init[1884]), .Q(o[1884]) );
  DFF \Data_Mem/memory_reg[58][29]  ( .D(\Data_Mem/n5902 ), .CLK(clk), .RST(
        rst), .I(e_init[1885]), .Q(o[1885]) );
  DFF \Data_Mem/memory_reg[58][30]  ( .D(\Data_Mem/n5903 ), .CLK(clk), .RST(
        rst), .I(e_init[1886]), .Q(o[1886]) );
  DFF \Data_Mem/memory_reg[58][31]  ( .D(\Data_Mem/n5904 ), .CLK(clk), .RST(
        rst), .I(e_init[1887]), .Q(o[1887]) );
  DFF \Data_Mem/memory_reg[57][0]  ( .D(\Data_Mem/n5905 ), .CLK(clk), .RST(rst), .I(e_init[1824]), .Q(o[1824]) );
  DFF \Data_Mem/memory_reg[57][1]  ( .D(\Data_Mem/n5906 ), .CLK(clk), .RST(rst), .I(e_init[1825]), .Q(o[1825]) );
  DFF \Data_Mem/memory_reg[57][2]  ( .D(\Data_Mem/n5907 ), .CLK(clk), .RST(rst), .I(e_init[1826]), .Q(o[1826]) );
  DFF \Data_Mem/memory_reg[57][3]  ( .D(\Data_Mem/n5908 ), .CLK(clk), .RST(rst), .I(e_init[1827]), .Q(o[1827]) );
  DFF \Data_Mem/memory_reg[57][4]  ( .D(\Data_Mem/n5909 ), .CLK(clk), .RST(rst), .I(e_init[1828]), .Q(o[1828]) );
  DFF \Data_Mem/memory_reg[57][5]  ( .D(\Data_Mem/n5910 ), .CLK(clk), .RST(rst), .I(e_init[1829]), .Q(o[1829]) );
  DFF \Data_Mem/memory_reg[57][6]  ( .D(\Data_Mem/n5911 ), .CLK(clk), .RST(rst), .I(e_init[1830]), .Q(o[1830]) );
  DFF \Data_Mem/memory_reg[57][7]  ( .D(\Data_Mem/n5912 ), .CLK(clk), .RST(rst), .I(e_init[1831]), .Q(o[1831]) );
  DFF \Data_Mem/memory_reg[57][8]  ( .D(\Data_Mem/n5913 ), .CLK(clk), .RST(rst), .I(e_init[1832]), .Q(o[1832]) );
  DFF \Data_Mem/memory_reg[57][9]  ( .D(\Data_Mem/n5914 ), .CLK(clk), .RST(rst), .I(e_init[1833]), .Q(o[1833]) );
  DFF \Data_Mem/memory_reg[57][10]  ( .D(\Data_Mem/n5915 ), .CLK(clk), .RST(
        rst), .I(e_init[1834]), .Q(o[1834]) );
  DFF \Data_Mem/memory_reg[57][11]  ( .D(\Data_Mem/n5916 ), .CLK(clk), .RST(
        rst), .I(e_init[1835]), .Q(o[1835]) );
  DFF \Data_Mem/memory_reg[57][12]  ( .D(\Data_Mem/n5917 ), .CLK(clk), .RST(
        rst), .I(e_init[1836]), .Q(o[1836]) );
  DFF \Data_Mem/memory_reg[57][13]  ( .D(\Data_Mem/n5918 ), .CLK(clk), .RST(
        rst), .I(e_init[1837]), .Q(o[1837]) );
  DFF \Data_Mem/memory_reg[57][14]  ( .D(\Data_Mem/n5919 ), .CLK(clk), .RST(
        rst), .I(e_init[1838]), .Q(o[1838]) );
  DFF \Data_Mem/memory_reg[57][15]  ( .D(\Data_Mem/n5920 ), .CLK(clk), .RST(
        rst), .I(e_init[1839]), .Q(o[1839]) );
  DFF \Data_Mem/memory_reg[57][16]  ( .D(\Data_Mem/n5921 ), .CLK(clk), .RST(
        rst), .I(e_init[1840]), .Q(o[1840]) );
  DFF \Data_Mem/memory_reg[57][17]  ( .D(\Data_Mem/n5922 ), .CLK(clk), .RST(
        rst), .I(e_init[1841]), .Q(o[1841]) );
  DFF \Data_Mem/memory_reg[57][18]  ( .D(\Data_Mem/n5923 ), .CLK(clk), .RST(
        rst), .I(e_init[1842]), .Q(o[1842]) );
  DFF \Data_Mem/memory_reg[57][19]  ( .D(\Data_Mem/n5924 ), .CLK(clk), .RST(
        rst), .I(e_init[1843]), .Q(o[1843]) );
  DFF \Data_Mem/memory_reg[57][20]  ( .D(\Data_Mem/n5925 ), .CLK(clk), .RST(
        rst), .I(e_init[1844]), .Q(o[1844]) );
  DFF \Data_Mem/memory_reg[57][21]  ( .D(\Data_Mem/n5926 ), .CLK(clk), .RST(
        rst), .I(e_init[1845]), .Q(o[1845]) );
  DFF \Data_Mem/memory_reg[57][22]  ( .D(\Data_Mem/n5927 ), .CLK(clk), .RST(
        rst), .I(e_init[1846]), .Q(o[1846]) );
  DFF \Data_Mem/memory_reg[57][23]  ( .D(\Data_Mem/n5928 ), .CLK(clk), .RST(
        rst), .I(e_init[1847]), .Q(o[1847]) );
  DFF \Data_Mem/memory_reg[57][24]  ( .D(\Data_Mem/n5929 ), .CLK(clk), .RST(
        rst), .I(e_init[1848]), .Q(o[1848]) );
  DFF \Data_Mem/memory_reg[57][25]  ( .D(\Data_Mem/n5930 ), .CLK(clk), .RST(
        rst), .I(e_init[1849]), .Q(o[1849]) );
  DFF \Data_Mem/memory_reg[57][26]  ( .D(\Data_Mem/n5931 ), .CLK(clk), .RST(
        rst), .I(e_init[1850]), .Q(o[1850]) );
  DFF \Data_Mem/memory_reg[57][27]  ( .D(\Data_Mem/n5932 ), .CLK(clk), .RST(
        rst), .I(e_init[1851]), .Q(o[1851]) );
  DFF \Data_Mem/memory_reg[57][28]  ( .D(\Data_Mem/n5933 ), .CLK(clk), .RST(
        rst), .I(e_init[1852]), .Q(o[1852]) );
  DFF \Data_Mem/memory_reg[57][29]  ( .D(\Data_Mem/n5934 ), .CLK(clk), .RST(
        rst), .I(e_init[1853]), .Q(o[1853]) );
  DFF \Data_Mem/memory_reg[57][30]  ( .D(\Data_Mem/n5935 ), .CLK(clk), .RST(
        rst), .I(e_init[1854]), .Q(o[1854]) );
  DFF \Data_Mem/memory_reg[57][31]  ( .D(\Data_Mem/n5936 ), .CLK(clk), .RST(
        rst), .I(e_init[1855]), .Q(o[1855]) );
  DFF \Data_Mem/memory_reg[56][0]  ( .D(\Data_Mem/n5937 ), .CLK(clk), .RST(rst), .I(e_init[1792]), .Q(o[1792]) );
  DFF \Data_Mem/memory_reg[56][1]  ( .D(\Data_Mem/n5938 ), .CLK(clk), .RST(rst), .I(e_init[1793]), .Q(o[1793]) );
  DFF \Data_Mem/memory_reg[56][2]  ( .D(\Data_Mem/n5939 ), .CLK(clk), .RST(rst), .I(e_init[1794]), .Q(o[1794]) );
  DFF \Data_Mem/memory_reg[56][3]  ( .D(\Data_Mem/n5940 ), .CLK(clk), .RST(rst), .I(e_init[1795]), .Q(o[1795]) );
  DFF \Data_Mem/memory_reg[56][4]  ( .D(\Data_Mem/n5941 ), .CLK(clk), .RST(rst), .I(e_init[1796]), .Q(o[1796]) );
  DFF \Data_Mem/memory_reg[56][5]  ( .D(\Data_Mem/n5942 ), .CLK(clk), .RST(rst), .I(e_init[1797]), .Q(o[1797]) );
  DFF \Data_Mem/memory_reg[56][6]  ( .D(\Data_Mem/n5943 ), .CLK(clk), .RST(rst), .I(e_init[1798]), .Q(o[1798]) );
  DFF \Data_Mem/memory_reg[56][7]  ( .D(\Data_Mem/n5944 ), .CLK(clk), .RST(rst), .I(e_init[1799]), .Q(o[1799]) );
  DFF \Data_Mem/memory_reg[56][8]  ( .D(\Data_Mem/n5945 ), .CLK(clk), .RST(rst), .I(e_init[1800]), .Q(o[1800]) );
  DFF \Data_Mem/memory_reg[56][9]  ( .D(\Data_Mem/n5946 ), .CLK(clk), .RST(rst), .I(e_init[1801]), .Q(o[1801]) );
  DFF \Data_Mem/memory_reg[56][10]  ( .D(\Data_Mem/n5947 ), .CLK(clk), .RST(
        rst), .I(e_init[1802]), .Q(o[1802]) );
  DFF \Data_Mem/memory_reg[56][11]  ( .D(\Data_Mem/n5948 ), .CLK(clk), .RST(
        rst), .I(e_init[1803]), .Q(o[1803]) );
  DFF \Data_Mem/memory_reg[56][12]  ( .D(\Data_Mem/n5949 ), .CLK(clk), .RST(
        rst), .I(e_init[1804]), .Q(o[1804]) );
  DFF \Data_Mem/memory_reg[56][13]  ( .D(\Data_Mem/n5950 ), .CLK(clk), .RST(
        rst), .I(e_init[1805]), .Q(o[1805]) );
  DFF \Data_Mem/memory_reg[56][14]  ( .D(\Data_Mem/n5951 ), .CLK(clk), .RST(
        rst), .I(e_init[1806]), .Q(o[1806]) );
  DFF \Data_Mem/memory_reg[56][15]  ( .D(\Data_Mem/n5952 ), .CLK(clk), .RST(
        rst), .I(e_init[1807]), .Q(o[1807]) );
  DFF \Data_Mem/memory_reg[56][16]  ( .D(\Data_Mem/n5953 ), .CLK(clk), .RST(
        rst), .I(e_init[1808]), .Q(o[1808]) );
  DFF \Data_Mem/memory_reg[56][17]  ( .D(\Data_Mem/n5954 ), .CLK(clk), .RST(
        rst), .I(e_init[1809]), .Q(o[1809]) );
  DFF \Data_Mem/memory_reg[56][18]  ( .D(\Data_Mem/n5955 ), .CLK(clk), .RST(
        rst), .I(e_init[1810]), .Q(o[1810]) );
  DFF \Data_Mem/memory_reg[56][19]  ( .D(\Data_Mem/n5956 ), .CLK(clk), .RST(
        rst), .I(e_init[1811]), .Q(o[1811]) );
  DFF \Data_Mem/memory_reg[56][20]  ( .D(\Data_Mem/n5957 ), .CLK(clk), .RST(
        rst), .I(e_init[1812]), .Q(o[1812]) );
  DFF \Data_Mem/memory_reg[56][21]  ( .D(\Data_Mem/n5958 ), .CLK(clk), .RST(
        rst), .I(e_init[1813]), .Q(o[1813]) );
  DFF \Data_Mem/memory_reg[56][22]  ( .D(\Data_Mem/n5959 ), .CLK(clk), .RST(
        rst), .I(e_init[1814]), .Q(o[1814]) );
  DFF \Data_Mem/memory_reg[56][23]  ( .D(\Data_Mem/n5960 ), .CLK(clk), .RST(
        rst), .I(e_init[1815]), .Q(o[1815]) );
  DFF \Data_Mem/memory_reg[56][24]  ( .D(\Data_Mem/n5961 ), .CLK(clk), .RST(
        rst), .I(e_init[1816]), .Q(o[1816]) );
  DFF \Data_Mem/memory_reg[56][25]  ( .D(\Data_Mem/n5962 ), .CLK(clk), .RST(
        rst), .I(e_init[1817]), .Q(o[1817]) );
  DFF \Data_Mem/memory_reg[56][26]  ( .D(\Data_Mem/n5963 ), .CLK(clk), .RST(
        rst), .I(e_init[1818]), .Q(o[1818]) );
  DFF \Data_Mem/memory_reg[56][27]  ( .D(\Data_Mem/n5964 ), .CLK(clk), .RST(
        rst), .I(e_init[1819]), .Q(o[1819]) );
  DFF \Data_Mem/memory_reg[56][28]  ( .D(\Data_Mem/n5965 ), .CLK(clk), .RST(
        rst), .I(e_init[1820]), .Q(o[1820]) );
  DFF \Data_Mem/memory_reg[56][29]  ( .D(\Data_Mem/n5966 ), .CLK(clk), .RST(
        rst), .I(e_init[1821]), .Q(o[1821]) );
  DFF \Data_Mem/memory_reg[56][30]  ( .D(\Data_Mem/n5967 ), .CLK(clk), .RST(
        rst), .I(e_init[1822]), .Q(o[1822]) );
  DFF \Data_Mem/memory_reg[56][31]  ( .D(\Data_Mem/n5968 ), .CLK(clk), .RST(
        rst), .I(e_init[1823]), .Q(o[1823]) );
  DFF \Data_Mem/memory_reg[55][0]  ( .D(\Data_Mem/n5969 ), .CLK(clk), .RST(rst), .I(e_init[1760]), .Q(o[1760]) );
  DFF \Data_Mem/memory_reg[55][1]  ( .D(\Data_Mem/n5970 ), .CLK(clk), .RST(rst), .I(e_init[1761]), .Q(o[1761]) );
  DFF \Data_Mem/memory_reg[55][2]  ( .D(\Data_Mem/n5971 ), .CLK(clk), .RST(rst), .I(e_init[1762]), .Q(o[1762]) );
  DFF \Data_Mem/memory_reg[55][3]  ( .D(\Data_Mem/n5972 ), .CLK(clk), .RST(rst), .I(e_init[1763]), .Q(o[1763]) );
  DFF \Data_Mem/memory_reg[55][4]  ( .D(\Data_Mem/n5973 ), .CLK(clk), .RST(rst), .I(e_init[1764]), .Q(o[1764]) );
  DFF \Data_Mem/memory_reg[55][5]  ( .D(\Data_Mem/n5974 ), .CLK(clk), .RST(rst), .I(e_init[1765]), .Q(o[1765]) );
  DFF \Data_Mem/memory_reg[55][6]  ( .D(\Data_Mem/n5975 ), .CLK(clk), .RST(rst), .I(e_init[1766]), .Q(o[1766]) );
  DFF \Data_Mem/memory_reg[55][7]  ( .D(\Data_Mem/n5976 ), .CLK(clk), .RST(rst), .I(e_init[1767]), .Q(o[1767]) );
  DFF \Data_Mem/memory_reg[55][8]  ( .D(\Data_Mem/n5977 ), .CLK(clk), .RST(rst), .I(e_init[1768]), .Q(o[1768]) );
  DFF \Data_Mem/memory_reg[55][9]  ( .D(\Data_Mem/n5978 ), .CLK(clk), .RST(rst), .I(e_init[1769]), .Q(o[1769]) );
  DFF \Data_Mem/memory_reg[55][10]  ( .D(\Data_Mem/n5979 ), .CLK(clk), .RST(
        rst), .I(e_init[1770]), .Q(o[1770]) );
  DFF \Data_Mem/memory_reg[55][11]  ( .D(\Data_Mem/n5980 ), .CLK(clk), .RST(
        rst), .I(e_init[1771]), .Q(o[1771]) );
  DFF \Data_Mem/memory_reg[55][12]  ( .D(\Data_Mem/n5981 ), .CLK(clk), .RST(
        rst), .I(e_init[1772]), .Q(o[1772]) );
  DFF \Data_Mem/memory_reg[55][13]  ( .D(\Data_Mem/n5982 ), .CLK(clk), .RST(
        rst), .I(e_init[1773]), .Q(o[1773]) );
  DFF \Data_Mem/memory_reg[55][14]  ( .D(\Data_Mem/n5983 ), .CLK(clk), .RST(
        rst), .I(e_init[1774]), .Q(o[1774]) );
  DFF \Data_Mem/memory_reg[55][15]  ( .D(\Data_Mem/n5984 ), .CLK(clk), .RST(
        rst), .I(e_init[1775]), .Q(o[1775]) );
  DFF \Data_Mem/memory_reg[55][16]  ( .D(\Data_Mem/n5985 ), .CLK(clk), .RST(
        rst), .I(e_init[1776]), .Q(o[1776]) );
  DFF \Data_Mem/memory_reg[55][17]  ( .D(\Data_Mem/n5986 ), .CLK(clk), .RST(
        rst), .I(e_init[1777]), .Q(o[1777]) );
  DFF \Data_Mem/memory_reg[55][18]  ( .D(\Data_Mem/n5987 ), .CLK(clk), .RST(
        rst), .I(e_init[1778]), .Q(o[1778]) );
  DFF \Data_Mem/memory_reg[55][19]  ( .D(\Data_Mem/n5988 ), .CLK(clk), .RST(
        rst), .I(e_init[1779]), .Q(o[1779]) );
  DFF \Data_Mem/memory_reg[55][20]  ( .D(\Data_Mem/n5989 ), .CLK(clk), .RST(
        rst), .I(e_init[1780]), .Q(o[1780]) );
  DFF \Data_Mem/memory_reg[55][21]  ( .D(\Data_Mem/n5990 ), .CLK(clk), .RST(
        rst), .I(e_init[1781]), .Q(o[1781]) );
  DFF \Data_Mem/memory_reg[55][22]  ( .D(\Data_Mem/n5991 ), .CLK(clk), .RST(
        rst), .I(e_init[1782]), .Q(o[1782]) );
  DFF \Data_Mem/memory_reg[55][23]  ( .D(\Data_Mem/n5992 ), .CLK(clk), .RST(
        rst), .I(e_init[1783]), .Q(o[1783]) );
  DFF \Data_Mem/memory_reg[55][24]  ( .D(\Data_Mem/n5993 ), .CLK(clk), .RST(
        rst), .I(e_init[1784]), .Q(o[1784]) );
  DFF \Data_Mem/memory_reg[55][25]  ( .D(\Data_Mem/n5994 ), .CLK(clk), .RST(
        rst), .I(e_init[1785]), .Q(o[1785]) );
  DFF \Data_Mem/memory_reg[55][26]  ( .D(\Data_Mem/n5995 ), .CLK(clk), .RST(
        rst), .I(e_init[1786]), .Q(o[1786]) );
  DFF \Data_Mem/memory_reg[55][27]  ( .D(\Data_Mem/n5996 ), .CLK(clk), .RST(
        rst), .I(e_init[1787]), .Q(o[1787]) );
  DFF \Data_Mem/memory_reg[55][28]  ( .D(\Data_Mem/n5997 ), .CLK(clk), .RST(
        rst), .I(e_init[1788]), .Q(o[1788]) );
  DFF \Data_Mem/memory_reg[55][29]  ( .D(\Data_Mem/n5998 ), .CLK(clk), .RST(
        rst), .I(e_init[1789]), .Q(o[1789]) );
  DFF \Data_Mem/memory_reg[55][30]  ( .D(\Data_Mem/n5999 ), .CLK(clk), .RST(
        rst), .I(e_init[1790]), .Q(o[1790]) );
  DFF \Data_Mem/memory_reg[55][31]  ( .D(\Data_Mem/n6000 ), .CLK(clk), .RST(
        rst), .I(e_init[1791]), .Q(o[1791]) );
  DFF \Data_Mem/memory_reg[54][0]  ( .D(\Data_Mem/n6001 ), .CLK(clk), .RST(rst), .I(e_init[1728]), .Q(o[1728]) );
  DFF \Data_Mem/memory_reg[54][1]  ( .D(\Data_Mem/n6002 ), .CLK(clk), .RST(rst), .I(e_init[1729]), .Q(o[1729]) );
  DFF \Data_Mem/memory_reg[54][2]  ( .D(\Data_Mem/n6003 ), .CLK(clk), .RST(rst), .I(e_init[1730]), .Q(o[1730]) );
  DFF \Data_Mem/memory_reg[54][3]  ( .D(\Data_Mem/n6004 ), .CLK(clk), .RST(rst), .I(e_init[1731]), .Q(o[1731]) );
  DFF \Data_Mem/memory_reg[54][4]  ( .D(\Data_Mem/n6005 ), .CLK(clk), .RST(rst), .I(e_init[1732]), .Q(o[1732]) );
  DFF \Data_Mem/memory_reg[54][5]  ( .D(\Data_Mem/n6006 ), .CLK(clk), .RST(rst), .I(e_init[1733]), .Q(o[1733]) );
  DFF \Data_Mem/memory_reg[54][6]  ( .D(\Data_Mem/n6007 ), .CLK(clk), .RST(rst), .I(e_init[1734]), .Q(o[1734]) );
  DFF \Data_Mem/memory_reg[54][7]  ( .D(\Data_Mem/n6008 ), .CLK(clk), .RST(rst), .I(e_init[1735]), .Q(o[1735]) );
  DFF \Data_Mem/memory_reg[54][8]  ( .D(\Data_Mem/n6009 ), .CLK(clk), .RST(rst), .I(e_init[1736]), .Q(o[1736]) );
  DFF \Data_Mem/memory_reg[54][9]  ( .D(\Data_Mem/n6010 ), .CLK(clk), .RST(rst), .I(e_init[1737]), .Q(o[1737]) );
  DFF \Data_Mem/memory_reg[54][10]  ( .D(\Data_Mem/n6011 ), .CLK(clk), .RST(
        rst), .I(e_init[1738]), .Q(o[1738]) );
  DFF \Data_Mem/memory_reg[54][11]  ( .D(\Data_Mem/n6012 ), .CLK(clk), .RST(
        rst), .I(e_init[1739]), .Q(o[1739]) );
  DFF \Data_Mem/memory_reg[54][12]  ( .D(\Data_Mem/n6013 ), .CLK(clk), .RST(
        rst), .I(e_init[1740]), .Q(o[1740]) );
  DFF \Data_Mem/memory_reg[54][13]  ( .D(\Data_Mem/n6014 ), .CLK(clk), .RST(
        rst), .I(e_init[1741]), .Q(o[1741]) );
  DFF \Data_Mem/memory_reg[54][14]  ( .D(\Data_Mem/n6015 ), .CLK(clk), .RST(
        rst), .I(e_init[1742]), .Q(o[1742]) );
  DFF \Data_Mem/memory_reg[54][15]  ( .D(\Data_Mem/n6016 ), .CLK(clk), .RST(
        rst), .I(e_init[1743]), .Q(o[1743]) );
  DFF \Data_Mem/memory_reg[54][16]  ( .D(\Data_Mem/n6017 ), .CLK(clk), .RST(
        rst), .I(e_init[1744]), .Q(o[1744]) );
  DFF \Data_Mem/memory_reg[54][17]  ( .D(\Data_Mem/n6018 ), .CLK(clk), .RST(
        rst), .I(e_init[1745]), .Q(o[1745]) );
  DFF \Data_Mem/memory_reg[54][18]  ( .D(\Data_Mem/n6019 ), .CLK(clk), .RST(
        rst), .I(e_init[1746]), .Q(o[1746]) );
  DFF \Data_Mem/memory_reg[54][19]  ( .D(\Data_Mem/n6020 ), .CLK(clk), .RST(
        rst), .I(e_init[1747]), .Q(o[1747]) );
  DFF \Data_Mem/memory_reg[54][20]  ( .D(\Data_Mem/n6021 ), .CLK(clk), .RST(
        rst), .I(e_init[1748]), .Q(o[1748]) );
  DFF \Data_Mem/memory_reg[54][21]  ( .D(\Data_Mem/n6022 ), .CLK(clk), .RST(
        rst), .I(e_init[1749]), .Q(o[1749]) );
  DFF \Data_Mem/memory_reg[54][22]  ( .D(\Data_Mem/n6023 ), .CLK(clk), .RST(
        rst), .I(e_init[1750]), .Q(o[1750]) );
  DFF \Data_Mem/memory_reg[54][23]  ( .D(\Data_Mem/n6024 ), .CLK(clk), .RST(
        rst), .I(e_init[1751]), .Q(o[1751]) );
  DFF \Data_Mem/memory_reg[54][24]  ( .D(\Data_Mem/n6025 ), .CLK(clk), .RST(
        rst), .I(e_init[1752]), .Q(o[1752]) );
  DFF \Data_Mem/memory_reg[54][25]  ( .D(\Data_Mem/n6026 ), .CLK(clk), .RST(
        rst), .I(e_init[1753]), .Q(o[1753]) );
  DFF \Data_Mem/memory_reg[54][26]  ( .D(\Data_Mem/n6027 ), .CLK(clk), .RST(
        rst), .I(e_init[1754]), .Q(o[1754]) );
  DFF \Data_Mem/memory_reg[54][27]  ( .D(\Data_Mem/n6028 ), .CLK(clk), .RST(
        rst), .I(e_init[1755]), .Q(o[1755]) );
  DFF \Data_Mem/memory_reg[54][28]  ( .D(\Data_Mem/n6029 ), .CLK(clk), .RST(
        rst), .I(e_init[1756]), .Q(o[1756]) );
  DFF \Data_Mem/memory_reg[54][29]  ( .D(\Data_Mem/n6030 ), .CLK(clk), .RST(
        rst), .I(e_init[1757]), .Q(o[1757]) );
  DFF \Data_Mem/memory_reg[54][30]  ( .D(\Data_Mem/n6031 ), .CLK(clk), .RST(
        rst), .I(e_init[1758]), .Q(o[1758]) );
  DFF \Data_Mem/memory_reg[54][31]  ( .D(\Data_Mem/n6032 ), .CLK(clk), .RST(
        rst), .I(e_init[1759]), .Q(o[1759]) );
  DFF \Data_Mem/memory_reg[53][0]  ( .D(\Data_Mem/n6033 ), .CLK(clk), .RST(rst), .I(e_init[1696]), .Q(o[1696]) );
  DFF \Data_Mem/memory_reg[53][1]  ( .D(\Data_Mem/n6034 ), .CLK(clk), .RST(rst), .I(e_init[1697]), .Q(o[1697]) );
  DFF \Data_Mem/memory_reg[53][2]  ( .D(\Data_Mem/n6035 ), .CLK(clk), .RST(rst), .I(e_init[1698]), .Q(o[1698]) );
  DFF \Data_Mem/memory_reg[53][3]  ( .D(\Data_Mem/n6036 ), .CLK(clk), .RST(rst), .I(e_init[1699]), .Q(o[1699]) );
  DFF \Data_Mem/memory_reg[53][4]  ( .D(\Data_Mem/n6037 ), .CLK(clk), .RST(rst), .I(e_init[1700]), .Q(o[1700]) );
  DFF \Data_Mem/memory_reg[53][5]  ( .D(\Data_Mem/n6038 ), .CLK(clk), .RST(rst), .I(e_init[1701]), .Q(o[1701]) );
  DFF \Data_Mem/memory_reg[53][6]  ( .D(\Data_Mem/n6039 ), .CLK(clk), .RST(rst), .I(e_init[1702]), .Q(o[1702]) );
  DFF \Data_Mem/memory_reg[53][7]  ( .D(\Data_Mem/n6040 ), .CLK(clk), .RST(rst), .I(e_init[1703]), .Q(o[1703]) );
  DFF \Data_Mem/memory_reg[53][8]  ( .D(\Data_Mem/n6041 ), .CLK(clk), .RST(rst), .I(e_init[1704]), .Q(o[1704]) );
  DFF \Data_Mem/memory_reg[53][9]  ( .D(\Data_Mem/n6042 ), .CLK(clk), .RST(rst), .I(e_init[1705]), .Q(o[1705]) );
  DFF \Data_Mem/memory_reg[53][10]  ( .D(\Data_Mem/n6043 ), .CLK(clk), .RST(
        rst), .I(e_init[1706]), .Q(o[1706]) );
  DFF \Data_Mem/memory_reg[53][11]  ( .D(\Data_Mem/n6044 ), .CLK(clk), .RST(
        rst), .I(e_init[1707]), .Q(o[1707]) );
  DFF \Data_Mem/memory_reg[53][12]  ( .D(\Data_Mem/n6045 ), .CLK(clk), .RST(
        rst), .I(e_init[1708]), .Q(o[1708]) );
  DFF \Data_Mem/memory_reg[53][13]  ( .D(\Data_Mem/n6046 ), .CLK(clk), .RST(
        rst), .I(e_init[1709]), .Q(o[1709]) );
  DFF \Data_Mem/memory_reg[53][14]  ( .D(\Data_Mem/n6047 ), .CLK(clk), .RST(
        rst), .I(e_init[1710]), .Q(o[1710]) );
  DFF \Data_Mem/memory_reg[53][15]  ( .D(\Data_Mem/n6048 ), .CLK(clk), .RST(
        rst), .I(e_init[1711]), .Q(o[1711]) );
  DFF \Data_Mem/memory_reg[53][16]  ( .D(\Data_Mem/n6049 ), .CLK(clk), .RST(
        rst), .I(e_init[1712]), .Q(o[1712]) );
  DFF \Data_Mem/memory_reg[53][17]  ( .D(\Data_Mem/n6050 ), .CLK(clk), .RST(
        rst), .I(e_init[1713]), .Q(o[1713]) );
  DFF \Data_Mem/memory_reg[53][18]  ( .D(\Data_Mem/n6051 ), .CLK(clk), .RST(
        rst), .I(e_init[1714]), .Q(o[1714]) );
  DFF \Data_Mem/memory_reg[53][19]  ( .D(\Data_Mem/n6052 ), .CLK(clk), .RST(
        rst), .I(e_init[1715]), .Q(o[1715]) );
  DFF \Data_Mem/memory_reg[53][20]  ( .D(\Data_Mem/n6053 ), .CLK(clk), .RST(
        rst), .I(e_init[1716]), .Q(o[1716]) );
  DFF \Data_Mem/memory_reg[53][21]  ( .D(\Data_Mem/n6054 ), .CLK(clk), .RST(
        rst), .I(e_init[1717]), .Q(o[1717]) );
  DFF \Data_Mem/memory_reg[53][22]  ( .D(\Data_Mem/n6055 ), .CLK(clk), .RST(
        rst), .I(e_init[1718]), .Q(o[1718]) );
  DFF \Data_Mem/memory_reg[53][23]  ( .D(\Data_Mem/n6056 ), .CLK(clk), .RST(
        rst), .I(e_init[1719]), .Q(o[1719]) );
  DFF \Data_Mem/memory_reg[53][24]  ( .D(\Data_Mem/n6057 ), .CLK(clk), .RST(
        rst), .I(e_init[1720]), .Q(o[1720]) );
  DFF \Data_Mem/memory_reg[53][25]  ( .D(\Data_Mem/n6058 ), .CLK(clk), .RST(
        rst), .I(e_init[1721]), .Q(o[1721]) );
  DFF \Data_Mem/memory_reg[53][26]  ( .D(\Data_Mem/n6059 ), .CLK(clk), .RST(
        rst), .I(e_init[1722]), .Q(o[1722]) );
  DFF \Data_Mem/memory_reg[53][27]  ( .D(\Data_Mem/n6060 ), .CLK(clk), .RST(
        rst), .I(e_init[1723]), .Q(o[1723]) );
  DFF \Data_Mem/memory_reg[53][28]  ( .D(\Data_Mem/n6061 ), .CLK(clk), .RST(
        rst), .I(e_init[1724]), .Q(o[1724]) );
  DFF \Data_Mem/memory_reg[53][29]  ( .D(\Data_Mem/n6062 ), .CLK(clk), .RST(
        rst), .I(e_init[1725]), .Q(o[1725]) );
  DFF \Data_Mem/memory_reg[53][30]  ( .D(\Data_Mem/n6063 ), .CLK(clk), .RST(
        rst), .I(e_init[1726]), .Q(o[1726]) );
  DFF \Data_Mem/memory_reg[53][31]  ( .D(\Data_Mem/n6064 ), .CLK(clk), .RST(
        rst), .I(e_init[1727]), .Q(o[1727]) );
  DFF \Data_Mem/memory_reg[52][0]  ( .D(\Data_Mem/n6065 ), .CLK(clk), .RST(rst), .I(e_init[1664]), .Q(o[1664]) );
  DFF \Data_Mem/memory_reg[52][1]  ( .D(\Data_Mem/n6066 ), .CLK(clk), .RST(rst), .I(e_init[1665]), .Q(o[1665]) );
  DFF \Data_Mem/memory_reg[52][2]  ( .D(\Data_Mem/n6067 ), .CLK(clk), .RST(rst), .I(e_init[1666]), .Q(o[1666]) );
  DFF \Data_Mem/memory_reg[52][3]  ( .D(\Data_Mem/n6068 ), .CLK(clk), .RST(rst), .I(e_init[1667]), .Q(o[1667]) );
  DFF \Data_Mem/memory_reg[52][4]  ( .D(\Data_Mem/n6069 ), .CLK(clk), .RST(rst), .I(e_init[1668]), .Q(o[1668]) );
  DFF \Data_Mem/memory_reg[52][5]  ( .D(\Data_Mem/n6070 ), .CLK(clk), .RST(rst), .I(e_init[1669]), .Q(o[1669]) );
  DFF \Data_Mem/memory_reg[52][6]  ( .D(\Data_Mem/n6071 ), .CLK(clk), .RST(rst), .I(e_init[1670]), .Q(o[1670]) );
  DFF \Data_Mem/memory_reg[52][7]  ( .D(\Data_Mem/n6072 ), .CLK(clk), .RST(rst), .I(e_init[1671]), .Q(o[1671]) );
  DFF \Data_Mem/memory_reg[52][8]  ( .D(\Data_Mem/n6073 ), .CLK(clk), .RST(rst), .I(e_init[1672]), .Q(o[1672]) );
  DFF \Data_Mem/memory_reg[52][9]  ( .D(\Data_Mem/n6074 ), .CLK(clk), .RST(rst), .I(e_init[1673]), .Q(o[1673]) );
  DFF \Data_Mem/memory_reg[52][10]  ( .D(\Data_Mem/n6075 ), .CLK(clk), .RST(
        rst), .I(e_init[1674]), .Q(o[1674]) );
  DFF \Data_Mem/memory_reg[52][11]  ( .D(\Data_Mem/n6076 ), .CLK(clk), .RST(
        rst), .I(e_init[1675]), .Q(o[1675]) );
  DFF \Data_Mem/memory_reg[52][12]  ( .D(\Data_Mem/n6077 ), .CLK(clk), .RST(
        rst), .I(e_init[1676]), .Q(o[1676]) );
  DFF \Data_Mem/memory_reg[52][13]  ( .D(\Data_Mem/n6078 ), .CLK(clk), .RST(
        rst), .I(e_init[1677]), .Q(o[1677]) );
  DFF \Data_Mem/memory_reg[52][14]  ( .D(\Data_Mem/n6079 ), .CLK(clk), .RST(
        rst), .I(e_init[1678]), .Q(o[1678]) );
  DFF \Data_Mem/memory_reg[52][15]  ( .D(\Data_Mem/n6080 ), .CLK(clk), .RST(
        rst), .I(e_init[1679]), .Q(o[1679]) );
  DFF \Data_Mem/memory_reg[52][16]  ( .D(\Data_Mem/n6081 ), .CLK(clk), .RST(
        rst), .I(e_init[1680]), .Q(o[1680]) );
  DFF \Data_Mem/memory_reg[52][17]  ( .D(\Data_Mem/n6082 ), .CLK(clk), .RST(
        rst), .I(e_init[1681]), .Q(o[1681]) );
  DFF \Data_Mem/memory_reg[52][18]  ( .D(\Data_Mem/n6083 ), .CLK(clk), .RST(
        rst), .I(e_init[1682]), .Q(o[1682]) );
  DFF \Data_Mem/memory_reg[52][19]  ( .D(\Data_Mem/n6084 ), .CLK(clk), .RST(
        rst), .I(e_init[1683]), .Q(o[1683]) );
  DFF \Data_Mem/memory_reg[52][20]  ( .D(\Data_Mem/n6085 ), .CLK(clk), .RST(
        rst), .I(e_init[1684]), .Q(o[1684]) );
  DFF \Data_Mem/memory_reg[52][21]  ( .D(\Data_Mem/n6086 ), .CLK(clk), .RST(
        rst), .I(e_init[1685]), .Q(o[1685]) );
  DFF \Data_Mem/memory_reg[52][22]  ( .D(\Data_Mem/n6087 ), .CLK(clk), .RST(
        rst), .I(e_init[1686]), .Q(o[1686]) );
  DFF \Data_Mem/memory_reg[52][23]  ( .D(\Data_Mem/n6088 ), .CLK(clk), .RST(
        rst), .I(e_init[1687]), .Q(o[1687]) );
  DFF \Data_Mem/memory_reg[52][24]  ( .D(\Data_Mem/n6089 ), .CLK(clk), .RST(
        rst), .I(e_init[1688]), .Q(o[1688]) );
  DFF \Data_Mem/memory_reg[52][25]  ( .D(\Data_Mem/n6090 ), .CLK(clk), .RST(
        rst), .I(e_init[1689]), .Q(o[1689]) );
  DFF \Data_Mem/memory_reg[52][26]  ( .D(\Data_Mem/n6091 ), .CLK(clk), .RST(
        rst), .I(e_init[1690]), .Q(o[1690]) );
  DFF \Data_Mem/memory_reg[52][27]  ( .D(\Data_Mem/n6092 ), .CLK(clk), .RST(
        rst), .I(e_init[1691]), .Q(o[1691]) );
  DFF \Data_Mem/memory_reg[52][28]  ( .D(\Data_Mem/n6093 ), .CLK(clk), .RST(
        rst), .I(e_init[1692]), .Q(o[1692]) );
  DFF \Data_Mem/memory_reg[52][29]  ( .D(\Data_Mem/n6094 ), .CLK(clk), .RST(
        rst), .I(e_init[1693]), .Q(o[1693]) );
  DFF \Data_Mem/memory_reg[52][30]  ( .D(\Data_Mem/n6095 ), .CLK(clk), .RST(
        rst), .I(e_init[1694]), .Q(o[1694]) );
  DFF \Data_Mem/memory_reg[52][31]  ( .D(\Data_Mem/n6096 ), .CLK(clk), .RST(
        rst), .I(e_init[1695]), .Q(o[1695]) );
  DFF \Data_Mem/memory_reg[51][0]  ( .D(\Data_Mem/n6097 ), .CLK(clk), .RST(rst), .I(e_init[1632]), .Q(o[1632]) );
  DFF \Data_Mem/memory_reg[51][1]  ( .D(\Data_Mem/n6098 ), .CLK(clk), .RST(rst), .I(e_init[1633]), .Q(o[1633]) );
  DFF \Data_Mem/memory_reg[51][2]  ( .D(\Data_Mem/n6099 ), .CLK(clk), .RST(rst), .I(e_init[1634]), .Q(o[1634]) );
  DFF \Data_Mem/memory_reg[51][3]  ( .D(\Data_Mem/n6100 ), .CLK(clk), .RST(rst), .I(e_init[1635]), .Q(o[1635]) );
  DFF \Data_Mem/memory_reg[51][4]  ( .D(\Data_Mem/n6101 ), .CLK(clk), .RST(rst), .I(e_init[1636]), .Q(o[1636]) );
  DFF \Data_Mem/memory_reg[51][5]  ( .D(\Data_Mem/n6102 ), .CLK(clk), .RST(rst), .I(e_init[1637]), .Q(o[1637]) );
  DFF \Data_Mem/memory_reg[51][6]  ( .D(\Data_Mem/n6103 ), .CLK(clk), .RST(rst), .I(e_init[1638]), .Q(o[1638]) );
  DFF \Data_Mem/memory_reg[51][7]  ( .D(\Data_Mem/n6104 ), .CLK(clk), .RST(rst), .I(e_init[1639]), .Q(o[1639]) );
  DFF \Data_Mem/memory_reg[51][8]  ( .D(\Data_Mem/n6105 ), .CLK(clk), .RST(rst), .I(e_init[1640]), .Q(o[1640]) );
  DFF \Data_Mem/memory_reg[51][9]  ( .D(\Data_Mem/n6106 ), .CLK(clk), .RST(rst), .I(e_init[1641]), .Q(o[1641]) );
  DFF \Data_Mem/memory_reg[51][10]  ( .D(\Data_Mem/n6107 ), .CLK(clk), .RST(
        rst), .I(e_init[1642]), .Q(o[1642]) );
  DFF \Data_Mem/memory_reg[51][11]  ( .D(\Data_Mem/n6108 ), .CLK(clk), .RST(
        rst), .I(e_init[1643]), .Q(o[1643]) );
  DFF \Data_Mem/memory_reg[51][12]  ( .D(\Data_Mem/n6109 ), .CLK(clk), .RST(
        rst), .I(e_init[1644]), .Q(o[1644]) );
  DFF \Data_Mem/memory_reg[51][13]  ( .D(\Data_Mem/n6110 ), .CLK(clk), .RST(
        rst), .I(e_init[1645]), .Q(o[1645]) );
  DFF \Data_Mem/memory_reg[51][14]  ( .D(\Data_Mem/n6111 ), .CLK(clk), .RST(
        rst), .I(e_init[1646]), .Q(o[1646]) );
  DFF \Data_Mem/memory_reg[51][15]  ( .D(\Data_Mem/n6112 ), .CLK(clk), .RST(
        rst), .I(e_init[1647]), .Q(o[1647]) );
  DFF \Data_Mem/memory_reg[51][16]  ( .D(\Data_Mem/n6113 ), .CLK(clk), .RST(
        rst), .I(e_init[1648]), .Q(o[1648]) );
  DFF \Data_Mem/memory_reg[51][17]  ( .D(\Data_Mem/n6114 ), .CLK(clk), .RST(
        rst), .I(e_init[1649]), .Q(o[1649]) );
  DFF \Data_Mem/memory_reg[51][18]  ( .D(\Data_Mem/n6115 ), .CLK(clk), .RST(
        rst), .I(e_init[1650]), .Q(o[1650]) );
  DFF \Data_Mem/memory_reg[51][19]  ( .D(\Data_Mem/n6116 ), .CLK(clk), .RST(
        rst), .I(e_init[1651]), .Q(o[1651]) );
  DFF \Data_Mem/memory_reg[51][20]  ( .D(\Data_Mem/n6117 ), .CLK(clk), .RST(
        rst), .I(e_init[1652]), .Q(o[1652]) );
  DFF \Data_Mem/memory_reg[51][21]  ( .D(\Data_Mem/n6118 ), .CLK(clk), .RST(
        rst), .I(e_init[1653]), .Q(o[1653]) );
  DFF \Data_Mem/memory_reg[51][22]  ( .D(\Data_Mem/n6119 ), .CLK(clk), .RST(
        rst), .I(e_init[1654]), .Q(o[1654]) );
  DFF \Data_Mem/memory_reg[51][23]  ( .D(\Data_Mem/n6120 ), .CLK(clk), .RST(
        rst), .I(e_init[1655]), .Q(o[1655]) );
  DFF \Data_Mem/memory_reg[51][24]  ( .D(\Data_Mem/n6121 ), .CLK(clk), .RST(
        rst), .I(e_init[1656]), .Q(o[1656]) );
  DFF \Data_Mem/memory_reg[51][25]  ( .D(\Data_Mem/n6122 ), .CLK(clk), .RST(
        rst), .I(e_init[1657]), .Q(o[1657]) );
  DFF \Data_Mem/memory_reg[51][26]  ( .D(\Data_Mem/n6123 ), .CLK(clk), .RST(
        rst), .I(e_init[1658]), .Q(o[1658]) );
  DFF \Data_Mem/memory_reg[51][27]  ( .D(\Data_Mem/n6124 ), .CLK(clk), .RST(
        rst), .I(e_init[1659]), .Q(o[1659]) );
  DFF \Data_Mem/memory_reg[51][28]  ( .D(\Data_Mem/n6125 ), .CLK(clk), .RST(
        rst), .I(e_init[1660]), .Q(o[1660]) );
  DFF \Data_Mem/memory_reg[51][29]  ( .D(\Data_Mem/n6126 ), .CLK(clk), .RST(
        rst), .I(e_init[1661]), .Q(o[1661]) );
  DFF \Data_Mem/memory_reg[51][30]  ( .D(\Data_Mem/n6127 ), .CLK(clk), .RST(
        rst), .I(e_init[1662]), .Q(o[1662]) );
  DFF \Data_Mem/memory_reg[51][31]  ( .D(\Data_Mem/n6128 ), .CLK(clk), .RST(
        rst), .I(e_init[1663]), .Q(o[1663]) );
  DFF \Data_Mem/memory_reg[50][0]  ( .D(\Data_Mem/n6129 ), .CLK(clk), .RST(rst), .I(e_init[1600]), .Q(o[1600]) );
  DFF \Data_Mem/memory_reg[50][1]  ( .D(\Data_Mem/n6130 ), .CLK(clk), .RST(rst), .I(e_init[1601]), .Q(o[1601]) );
  DFF \Data_Mem/memory_reg[50][2]  ( .D(\Data_Mem/n6131 ), .CLK(clk), .RST(rst), .I(e_init[1602]), .Q(o[1602]) );
  DFF \Data_Mem/memory_reg[50][3]  ( .D(\Data_Mem/n6132 ), .CLK(clk), .RST(rst), .I(e_init[1603]), .Q(o[1603]) );
  DFF \Data_Mem/memory_reg[50][4]  ( .D(\Data_Mem/n6133 ), .CLK(clk), .RST(rst), .I(e_init[1604]), .Q(o[1604]) );
  DFF \Data_Mem/memory_reg[50][5]  ( .D(\Data_Mem/n6134 ), .CLK(clk), .RST(rst), .I(e_init[1605]), .Q(o[1605]) );
  DFF \Data_Mem/memory_reg[50][6]  ( .D(\Data_Mem/n6135 ), .CLK(clk), .RST(rst), .I(e_init[1606]), .Q(o[1606]) );
  DFF \Data_Mem/memory_reg[50][7]  ( .D(\Data_Mem/n6136 ), .CLK(clk), .RST(rst), .I(e_init[1607]), .Q(o[1607]) );
  DFF \Data_Mem/memory_reg[50][8]  ( .D(\Data_Mem/n6137 ), .CLK(clk), .RST(rst), .I(e_init[1608]), .Q(o[1608]) );
  DFF \Data_Mem/memory_reg[50][9]  ( .D(\Data_Mem/n6138 ), .CLK(clk), .RST(rst), .I(e_init[1609]), .Q(o[1609]) );
  DFF \Data_Mem/memory_reg[50][10]  ( .D(\Data_Mem/n6139 ), .CLK(clk), .RST(
        rst), .I(e_init[1610]), .Q(o[1610]) );
  DFF \Data_Mem/memory_reg[50][11]  ( .D(\Data_Mem/n6140 ), .CLK(clk), .RST(
        rst), .I(e_init[1611]), .Q(o[1611]) );
  DFF \Data_Mem/memory_reg[50][12]  ( .D(\Data_Mem/n6141 ), .CLK(clk), .RST(
        rst), .I(e_init[1612]), .Q(o[1612]) );
  DFF \Data_Mem/memory_reg[50][13]  ( .D(\Data_Mem/n6142 ), .CLK(clk), .RST(
        rst), .I(e_init[1613]), .Q(o[1613]) );
  DFF \Data_Mem/memory_reg[50][14]  ( .D(\Data_Mem/n6143 ), .CLK(clk), .RST(
        rst), .I(e_init[1614]), .Q(o[1614]) );
  DFF \Data_Mem/memory_reg[50][15]  ( .D(\Data_Mem/n6144 ), .CLK(clk), .RST(
        rst), .I(e_init[1615]), .Q(o[1615]) );
  DFF \Data_Mem/memory_reg[50][16]  ( .D(\Data_Mem/n6145 ), .CLK(clk), .RST(
        rst), .I(e_init[1616]), .Q(o[1616]) );
  DFF \Data_Mem/memory_reg[50][17]  ( .D(\Data_Mem/n6146 ), .CLK(clk), .RST(
        rst), .I(e_init[1617]), .Q(o[1617]) );
  DFF \Data_Mem/memory_reg[50][18]  ( .D(\Data_Mem/n6147 ), .CLK(clk), .RST(
        rst), .I(e_init[1618]), .Q(o[1618]) );
  DFF \Data_Mem/memory_reg[50][19]  ( .D(\Data_Mem/n6148 ), .CLK(clk), .RST(
        rst), .I(e_init[1619]), .Q(o[1619]) );
  DFF \Data_Mem/memory_reg[50][20]  ( .D(\Data_Mem/n6149 ), .CLK(clk), .RST(
        rst), .I(e_init[1620]), .Q(o[1620]) );
  DFF \Data_Mem/memory_reg[50][21]  ( .D(\Data_Mem/n6150 ), .CLK(clk), .RST(
        rst), .I(e_init[1621]), .Q(o[1621]) );
  DFF \Data_Mem/memory_reg[50][22]  ( .D(\Data_Mem/n6151 ), .CLK(clk), .RST(
        rst), .I(e_init[1622]), .Q(o[1622]) );
  DFF \Data_Mem/memory_reg[50][23]  ( .D(\Data_Mem/n6152 ), .CLK(clk), .RST(
        rst), .I(e_init[1623]), .Q(o[1623]) );
  DFF \Data_Mem/memory_reg[50][24]  ( .D(\Data_Mem/n6153 ), .CLK(clk), .RST(
        rst), .I(e_init[1624]), .Q(o[1624]) );
  DFF \Data_Mem/memory_reg[50][25]  ( .D(\Data_Mem/n6154 ), .CLK(clk), .RST(
        rst), .I(e_init[1625]), .Q(o[1625]) );
  DFF \Data_Mem/memory_reg[50][26]  ( .D(\Data_Mem/n6155 ), .CLK(clk), .RST(
        rst), .I(e_init[1626]), .Q(o[1626]) );
  DFF \Data_Mem/memory_reg[50][27]  ( .D(\Data_Mem/n6156 ), .CLK(clk), .RST(
        rst), .I(e_init[1627]), .Q(o[1627]) );
  DFF \Data_Mem/memory_reg[50][28]  ( .D(\Data_Mem/n6157 ), .CLK(clk), .RST(
        rst), .I(e_init[1628]), .Q(o[1628]) );
  DFF \Data_Mem/memory_reg[50][29]  ( .D(\Data_Mem/n6158 ), .CLK(clk), .RST(
        rst), .I(e_init[1629]), .Q(o[1629]) );
  DFF \Data_Mem/memory_reg[50][30]  ( .D(\Data_Mem/n6159 ), .CLK(clk), .RST(
        rst), .I(e_init[1630]), .Q(o[1630]) );
  DFF \Data_Mem/memory_reg[50][31]  ( .D(\Data_Mem/n6160 ), .CLK(clk), .RST(
        rst), .I(e_init[1631]), .Q(o[1631]) );
  DFF \Data_Mem/memory_reg[49][0]  ( .D(\Data_Mem/n6161 ), .CLK(clk), .RST(rst), .I(e_init[1568]), .Q(o[1568]) );
  DFF \Data_Mem/memory_reg[49][1]  ( .D(\Data_Mem/n6162 ), .CLK(clk), .RST(rst), .I(e_init[1569]), .Q(o[1569]) );
  DFF \Data_Mem/memory_reg[49][2]  ( .D(\Data_Mem/n6163 ), .CLK(clk), .RST(rst), .I(e_init[1570]), .Q(o[1570]) );
  DFF \Data_Mem/memory_reg[49][3]  ( .D(\Data_Mem/n6164 ), .CLK(clk), .RST(rst), .I(e_init[1571]), .Q(o[1571]) );
  DFF \Data_Mem/memory_reg[49][4]  ( .D(\Data_Mem/n6165 ), .CLK(clk), .RST(rst), .I(e_init[1572]), .Q(o[1572]) );
  DFF \Data_Mem/memory_reg[49][5]  ( .D(\Data_Mem/n6166 ), .CLK(clk), .RST(rst), .I(e_init[1573]), .Q(o[1573]) );
  DFF \Data_Mem/memory_reg[49][6]  ( .D(\Data_Mem/n6167 ), .CLK(clk), .RST(rst), .I(e_init[1574]), .Q(o[1574]) );
  DFF \Data_Mem/memory_reg[49][7]  ( .D(\Data_Mem/n6168 ), .CLK(clk), .RST(rst), .I(e_init[1575]), .Q(o[1575]) );
  DFF \Data_Mem/memory_reg[49][8]  ( .D(\Data_Mem/n6169 ), .CLK(clk), .RST(rst), .I(e_init[1576]), .Q(o[1576]) );
  DFF \Data_Mem/memory_reg[49][9]  ( .D(\Data_Mem/n6170 ), .CLK(clk), .RST(rst), .I(e_init[1577]), .Q(o[1577]) );
  DFF \Data_Mem/memory_reg[49][10]  ( .D(\Data_Mem/n6171 ), .CLK(clk), .RST(
        rst), .I(e_init[1578]), .Q(o[1578]) );
  DFF \Data_Mem/memory_reg[49][11]  ( .D(\Data_Mem/n6172 ), .CLK(clk), .RST(
        rst), .I(e_init[1579]), .Q(o[1579]) );
  DFF \Data_Mem/memory_reg[49][12]  ( .D(\Data_Mem/n6173 ), .CLK(clk), .RST(
        rst), .I(e_init[1580]), .Q(o[1580]) );
  DFF \Data_Mem/memory_reg[49][13]  ( .D(\Data_Mem/n6174 ), .CLK(clk), .RST(
        rst), .I(e_init[1581]), .Q(o[1581]) );
  DFF \Data_Mem/memory_reg[49][14]  ( .D(\Data_Mem/n6175 ), .CLK(clk), .RST(
        rst), .I(e_init[1582]), .Q(o[1582]) );
  DFF \Data_Mem/memory_reg[49][15]  ( .D(\Data_Mem/n6176 ), .CLK(clk), .RST(
        rst), .I(e_init[1583]), .Q(o[1583]) );
  DFF \Data_Mem/memory_reg[49][16]  ( .D(\Data_Mem/n6177 ), .CLK(clk), .RST(
        rst), .I(e_init[1584]), .Q(o[1584]) );
  DFF \Data_Mem/memory_reg[49][17]  ( .D(\Data_Mem/n6178 ), .CLK(clk), .RST(
        rst), .I(e_init[1585]), .Q(o[1585]) );
  DFF \Data_Mem/memory_reg[49][18]  ( .D(\Data_Mem/n6179 ), .CLK(clk), .RST(
        rst), .I(e_init[1586]), .Q(o[1586]) );
  DFF \Data_Mem/memory_reg[49][19]  ( .D(\Data_Mem/n6180 ), .CLK(clk), .RST(
        rst), .I(e_init[1587]), .Q(o[1587]) );
  DFF \Data_Mem/memory_reg[49][20]  ( .D(\Data_Mem/n6181 ), .CLK(clk), .RST(
        rst), .I(e_init[1588]), .Q(o[1588]) );
  DFF \Data_Mem/memory_reg[49][21]  ( .D(\Data_Mem/n6182 ), .CLK(clk), .RST(
        rst), .I(e_init[1589]), .Q(o[1589]) );
  DFF \Data_Mem/memory_reg[49][22]  ( .D(\Data_Mem/n6183 ), .CLK(clk), .RST(
        rst), .I(e_init[1590]), .Q(o[1590]) );
  DFF \Data_Mem/memory_reg[49][23]  ( .D(\Data_Mem/n6184 ), .CLK(clk), .RST(
        rst), .I(e_init[1591]), .Q(o[1591]) );
  DFF \Data_Mem/memory_reg[49][24]  ( .D(\Data_Mem/n6185 ), .CLK(clk), .RST(
        rst), .I(e_init[1592]), .Q(o[1592]) );
  DFF \Data_Mem/memory_reg[49][25]  ( .D(\Data_Mem/n6186 ), .CLK(clk), .RST(
        rst), .I(e_init[1593]), .Q(o[1593]) );
  DFF \Data_Mem/memory_reg[49][26]  ( .D(\Data_Mem/n6187 ), .CLK(clk), .RST(
        rst), .I(e_init[1594]), .Q(o[1594]) );
  DFF \Data_Mem/memory_reg[49][27]  ( .D(\Data_Mem/n6188 ), .CLK(clk), .RST(
        rst), .I(e_init[1595]), .Q(o[1595]) );
  DFF \Data_Mem/memory_reg[49][28]  ( .D(\Data_Mem/n6189 ), .CLK(clk), .RST(
        rst), .I(e_init[1596]), .Q(o[1596]) );
  DFF \Data_Mem/memory_reg[49][29]  ( .D(\Data_Mem/n6190 ), .CLK(clk), .RST(
        rst), .I(e_init[1597]), .Q(o[1597]) );
  DFF \Data_Mem/memory_reg[49][30]  ( .D(\Data_Mem/n6191 ), .CLK(clk), .RST(
        rst), .I(e_init[1598]), .Q(o[1598]) );
  DFF \Data_Mem/memory_reg[49][31]  ( .D(\Data_Mem/n6192 ), .CLK(clk), .RST(
        rst), .I(e_init[1599]), .Q(o[1599]) );
  DFF \Data_Mem/memory_reg[48][0]  ( .D(\Data_Mem/n6193 ), .CLK(clk), .RST(rst), .I(e_init[1536]), .Q(o[1536]) );
  DFF \Data_Mem/memory_reg[48][1]  ( .D(\Data_Mem/n6194 ), .CLK(clk), .RST(rst), .I(e_init[1537]), .Q(o[1537]) );
  DFF \Data_Mem/memory_reg[48][2]  ( .D(\Data_Mem/n6195 ), .CLK(clk), .RST(rst), .I(e_init[1538]), .Q(o[1538]) );
  DFF \Data_Mem/memory_reg[48][3]  ( .D(\Data_Mem/n6196 ), .CLK(clk), .RST(rst), .I(e_init[1539]), .Q(o[1539]) );
  DFF \Data_Mem/memory_reg[48][4]  ( .D(\Data_Mem/n6197 ), .CLK(clk), .RST(rst), .I(e_init[1540]), .Q(o[1540]) );
  DFF \Data_Mem/memory_reg[48][5]  ( .D(\Data_Mem/n6198 ), .CLK(clk), .RST(rst), .I(e_init[1541]), .Q(o[1541]) );
  DFF \Data_Mem/memory_reg[48][6]  ( .D(\Data_Mem/n6199 ), .CLK(clk), .RST(rst), .I(e_init[1542]), .Q(o[1542]) );
  DFF \Data_Mem/memory_reg[48][7]  ( .D(\Data_Mem/n6200 ), .CLK(clk), .RST(rst), .I(e_init[1543]), .Q(o[1543]) );
  DFF \Data_Mem/memory_reg[48][8]  ( .D(\Data_Mem/n6201 ), .CLK(clk), .RST(rst), .I(e_init[1544]), .Q(o[1544]) );
  DFF \Data_Mem/memory_reg[48][9]  ( .D(\Data_Mem/n6202 ), .CLK(clk), .RST(rst), .I(e_init[1545]), .Q(o[1545]) );
  DFF \Data_Mem/memory_reg[48][10]  ( .D(\Data_Mem/n6203 ), .CLK(clk), .RST(
        rst), .I(e_init[1546]), .Q(o[1546]) );
  DFF \Data_Mem/memory_reg[48][11]  ( .D(\Data_Mem/n6204 ), .CLK(clk), .RST(
        rst), .I(e_init[1547]), .Q(o[1547]) );
  DFF \Data_Mem/memory_reg[48][12]  ( .D(\Data_Mem/n6205 ), .CLK(clk), .RST(
        rst), .I(e_init[1548]), .Q(o[1548]) );
  DFF \Data_Mem/memory_reg[48][13]  ( .D(\Data_Mem/n6206 ), .CLK(clk), .RST(
        rst), .I(e_init[1549]), .Q(o[1549]) );
  DFF \Data_Mem/memory_reg[48][14]  ( .D(\Data_Mem/n6207 ), .CLK(clk), .RST(
        rst), .I(e_init[1550]), .Q(o[1550]) );
  DFF \Data_Mem/memory_reg[48][15]  ( .D(\Data_Mem/n6208 ), .CLK(clk), .RST(
        rst), .I(e_init[1551]), .Q(o[1551]) );
  DFF \Data_Mem/memory_reg[48][16]  ( .D(\Data_Mem/n6209 ), .CLK(clk), .RST(
        rst), .I(e_init[1552]), .Q(o[1552]) );
  DFF \Data_Mem/memory_reg[48][17]  ( .D(\Data_Mem/n6210 ), .CLK(clk), .RST(
        rst), .I(e_init[1553]), .Q(o[1553]) );
  DFF \Data_Mem/memory_reg[48][18]  ( .D(\Data_Mem/n6211 ), .CLK(clk), .RST(
        rst), .I(e_init[1554]), .Q(o[1554]) );
  DFF \Data_Mem/memory_reg[48][19]  ( .D(\Data_Mem/n6212 ), .CLK(clk), .RST(
        rst), .I(e_init[1555]), .Q(o[1555]) );
  DFF \Data_Mem/memory_reg[48][20]  ( .D(\Data_Mem/n6213 ), .CLK(clk), .RST(
        rst), .I(e_init[1556]), .Q(o[1556]) );
  DFF \Data_Mem/memory_reg[48][21]  ( .D(\Data_Mem/n6214 ), .CLK(clk), .RST(
        rst), .I(e_init[1557]), .Q(o[1557]) );
  DFF \Data_Mem/memory_reg[48][22]  ( .D(\Data_Mem/n6215 ), .CLK(clk), .RST(
        rst), .I(e_init[1558]), .Q(o[1558]) );
  DFF \Data_Mem/memory_reg[48][23]  ( .D(\Data_Mem/n6216 ), .CLK(clk), .RST(
        rst), .I(e_init[1559]), .Q(o[1559]) );
  DFF \Data_Mem/memory_reg[48][24]  ( .D(\Data_Mem/n6217 ), .CLK(clk), .RST(
        rst), .I(e_init[1560]), .Q(o[1560]) );
  DFF \Data_Mem/memory_reg[48][25]  ( .D(\Data_Mem/n6218 ), .CLK(clk), .RST(
        rst), .I(e_init[1561]), .Q(o[1561]) );
  DFF \Data_Mem/memory_reg[48][26]  ( .D(\Data_Mem/n6219 ), .CLK(clk), .RST(
        rst), .I(e_init[1562]), .Q(o[1562]) );
  DFF \Data_Mem/memory_reg[48][27]  ( .D(\Data_Mem/n6220 ), .CLK(clk), .RST(
        rst), .I(e_init[1563]), .Q(o[1563]) );
  DFF \Data_Mem/memory_reg[48][28]  ( .D(\Data_Mem/n6221 ), .CLK(clk), .RST(
        rst), .I(e_init[1564]), .Q(o[1564]) );
  DFF \Data_Mem/memory_reg[48][29]  ( .D(\Data_Mem/n6222 ), .CLK(clk), .RST(
        rst), .I(e_init[1565]), .Q(o[1565]) );
  DFF \Data_Mem/memory_reg[48][30]  ( .D(\Data_Mem/n6223 ), .CLK(clk), .RST(
        rst), .I(e_init[1566]), .Q(o[1566]) );
  DFF \Data_Mem/memory_reg[48][31]  ( .D(\Data_Mem/n6224 ), .CLK(clk), .RST(
        rst), .I(e_init[1567]), .Q(o[1567]) );
  DFF \Data_Mem/memory_reg[47][0]  ( .D(\Data_Mem/n6225 ), .CLK(clk), .RST(rst), .I(e_init[1504]), .Q(o[1504]) );
  DFF \Data_Mem/memory_reg[47][1]  ( .D(\Data_Mem/n6226 ), .CLK(clk), .RST(rst), .I(e_init[1505]), .Q(o[1505]) );
  DFF \Data_Mem/memory_reg[47][2]  ( .D(\Data_Mem/n6227 ), .CLK(clk), .RST(rst), .I(e_init[1506]), .Q(o[1506]) );
  DFF \Data_Mem/memory_reg[47][3]  ( .D(\Data_Mem/n6228 ), .CLK(clk), .RST(rst), .I(e_init[1507]), .Q(o[1507]) );
  DFF \Data_Mem/memory_reg[47][4]  ( .D(\Data_Mem/n6229 ), .CLK(clk), .RST(rst), .I(e_init[1508]), .Q(o[1508]) );
  DFF \Data_Mem/memory_reg[47][5]  ( .D(\Data_Mem/n6230 ), .CLK(clk), .RST(rst), .I(e_init[1509]), .Q(o[1509]) );
  DFF \Data_Mem/memory_reg[47][6]  ( .D(\Data_Mem/n6231 ), .CLK(clk), .RST(rst), .I(e_init[1510]), .Q(o[1510]) );
  DFF \Data_Mem/memory_reg[47][7]  ( .D(\Data_Mem/n6232 ), .CLK(clk), .RST(rst), .I(e_init[1511]), .Q(o[1511]) );
  DFF \Data_Mem/memory_reg[47][8]  ( .D(\Data_Mem/n6233 ), .CLK(clk), .RST(rst), .I(e_init[1512]), .Q(o[1512]) );
  DFF \Data_Mem/memory_reg[47][9]  ( .D(\Data_Mem/n6234 ), .CLK(clk), .RST(rst), .I(e_init[1513]), .Q(o[1513]) );
  DFF \Data_Mem/memory_reg[47][10]  ( .D(\Data_Mem/n6235 ), .CLK(clk), .RST(
        rst), .I(e_init[1514]), .Q(o[1514]) );
  DFF \Data_Mem/memory_reg[47][11]  ( .D(\Data_Mem/n6236 ), .CLK(clk), .RST(
        rst), .I(e_init[1515]), .Q(o[1515]) );
  DFF \Data_Mem/memory_reg[47][12]  ( .D(\Data_Mem/n6237 ), .CLK(clk), .RST(
        rst), .I(e_init[1516]), .Q(o[1516]) );
  DFF \Data_Mem/memory_reg[47][13]  ( .D(\Data_Mem/n6238 ), .CLK(clk), .RST(
        rst), .I(e_init[1517]), .Q(o[1517]) );
  DFF \Data_Mem/memory_reg[47][14]  ( .D(\Data_Mem/n6239 ), .CLK(clk), .RST(
        rst), .I(e_init[1518]), .Q(o[1518]) );
  DFF \Data_Mem/memory_reg[47][15]  ( .D(\Data_Mem/n6240 ), .CLK(clk), .RST(
        rst), .I(e_init[1519]), .Q(o[1519]) );
  DFF \Data_Mem/memory_reg[47][16]  ( .D(\Data_Mem/n6241 ), .CLK(clk), .RST(
        rst), .I(e_init[1520]), .Q(o[1520]) );
  DFF \Data_Mem/memory_reg[47][17]  ( .D(\Data_Mem/n6242 ), .CLK(clk), .RST(
        rst), .I(e_init[1521]), .Q(o[1521]) );
  DFF \Data_Mem/memory_reg[47][18]  ( .D(\Data_Mem/n6243 ), .CLK(clk), .RST(
        rst), .I(e_init[1522]), .Q(o[1522]) );
  DFF \Data_Mem/memory_reg[47][19]  ( .D(\Data_Mem/n6244 ), .CLK(clk), .RST(
        rst), .I(e_init[1523]), .Q(o[1523]) );
  DFF \Data_Mem/memory_reg[47][20]  ( .D(\Data_Mem/n6245 ), .CLK(clk), .RST(
        rst), .I(e_init[1524]), .Q(o[1524]) );
  DFF \Data_Mem/memory_reg[47][21]  ( .D(\Data_Mem/n6246 ), .CLK(clk), .RST(
        rst), .I(e_init[1525]), .Q(o[1525]) );
  DFF \Data_Mem/memory_reg[47][22]  ( .D(\Data_Mem/n6247 ), .CLK(clk), .RST(
        rst), .I(e_init[1526]), .Q(o[1526]) );
  DFF \Data_Mem/memory_reg[47][23]  ( .D(\Data_Mem/n6248 ), .CLK(clk), .RST(
        rst), .I(e_init[1527]), .Q(o[1527]) );
  DFF \Data_Mem/memory_reg[47][24]  ( .D(\Data_Mem/n6249 ), .CLK(clk), .RST(
        rst), .I(e_init[1528]), .Q(o[1528]) );
  DFF \Data_Mem/memory_reg[47][25]  ( .D(\Data_Mem/n6250 ), .CLK(clk), .RST(
        rst), .I(e_init[1529]), .Q(o[1529]) );
  DFF \Data_Mem/memory_reg[47][26]  ( .D(\Data_Mem/n6251 ), .CLK(clk), .RST(
        rst), .I(e_init[1530]), .Q(o[1530]) );
  DFF \Data_Mem/memory_reg[47][27]  ( .D(\Data_Mem/n6252 ), .CLK(clk), .RST(
        rst), .I(e_init[1531]), .Q(o[1531]) );
  DFF \Data_Mem/memory_reg[47][28]  ( .D(\Data_Mem/n6253 ), .CLK(clk), .RST(
        rst), .I(e_init[1532]), .Q(o[1532]) );
  DFF \Data_Mem/memory_reg[47][29]  ( .D(\Data_Mem/n6254 ), .CLK(clk), .RST(
        rst), .I(e_init[1533]), .Q(o[1533]) );
  DFF \Data_Mem/memory_reg[47][30]  ( .D(\Data_Mem/n6255 ), .CLK(clk), .RST(
        rst), .I(e_init[1534]), .Q(o[1534]) );
  DFF \Data_Mem/memory_reg[47][31]  ( .D(\Data_Mem/n6256 ), .CLK(clk), .RST(
        rst), .I(e_init[1535]), .Q(o[1535]) );
  DFF \Data_Mem/memory_reg[46][0]  ( .D(\Data_Mem/n6257 ), .CLK(clk), .RST(rst), .I(e_init[1472]), .Q(o[1472]) );
  DFF \Data_Mem/memory_reg[46][1]  ( .D(\Data_Mem/n6258 ), .CLK(clk), .RST(rst), .I(e_init[1473]), .Q(o[1473]) );
  DFF \Data_Mem/memory_reg[46][2]  ( .D(\Data_Mem/n6259 ), .CLK(clk), .RST(rst), .I(e_init[1474]), .Q(o[1474]) );
  DFF \Data_Mem/memory_reg[46][3]  ( .D(\Data_Mem/n6260 ), .CLK(clk), .RST(rst), .I(e_init[1475]), .Q(o[1475]) );
  DFF \Data_Mem/memory_reg[46][4]  ( .D(\Data_Mem/n6261 ), .CLK(clk), .RST(rst), .I(e_init[1476]), .Q(o[1476]) );
  DFF \Data_Mem/memory_reg[46][5]  ( .D(\Data_Mem/n6262 ), .CLK(clk), .RST(rst), .I(e_init[1477]), .Q(o[1477]) );
  DFF \Data_Mem/memory_reg[46][6]  ( .D(\Data_Mem/n6263 ), .CLK(clk), .RST(rst), .I(e_init[1478]), .Q(o[1478]) );
  DFF \Data_Mem/memory_reg[46][7]  ( .D(\Data_Mem/n6264 ), .CLK(clk), .RST(rst), .I(e_init[1479]), .Q(o[1479]) );
  DFF \Data_Mem/memory_reg[46][8]  ( .D(\Data_Mem/n6265 ), .CLK(clk), .RST(rst), .I(e_init[1480]), .Q(o[1480]) );
  DFF \Data_Mem/memory_reg[46][9]  ( .D(\Data_Mem/n6266 ), .CLK(clk), .RST(rst), .I(e_init[1481]), .Q(o[1481]) );
  DFF \Data_Mem/memory_reg[46][10]  ( .D(\Data_Mem/n6267 ), .CLK(clk), .RST(
        rst), .I(e_init[1482]), .Q(o[1482]) );
  DFF \Data_Mem/memory_reg[46][11]  ( .D(\Data_Mem/n6268 ), .CLK(clk), .RST(
        rst), .I(e_init[1483]), .Q(o[1483]) );
  DFF \Data_Mem/memory_reg[46][12]  ( .D(\Data_Mem/n6269 ), .CLK(clk), .RST(
        rst), .I(e_init[1484]), .Q(o[1484]) );
  DFF \Data_Mem/memory_reg[46][13]  ( .D(\Data_Mem/n6270 ), .CLK(clk), .RST(
        rst), .I(e_init[1485]), .Q(o[1485]) );
  DFF \Data_Mem/memory_reg[46][14]  ( .D(\Data_Mem/n6271 ), .CLK(clk), .RST(
        rst), .I(e_init[1486]), .Q(o[1486]) );
  DFF \Data_Mem/memory_reg[46][15]  ( .D(\Data_Mem/n6272 ), .CLK(clk), .RST(
        rst), .I(e_init[1487]), .Q(o[1487]) );
  DFF \Data_Mem/memory_reg[46][16]  ( .D(\Data_Mem/n6273 ), .CLK(clk), .RST(
        rst), .I(e_init[1488]), .Q(o[1488]) );
  DFF \Data_Mem/memory_reg[46][17]  ( .D(\Data_Mem/n6274 ), .CLK(clk), .RST(
        rst), .I(e_init[1489]), .Q(o[1489]) );
  DFF \Data_Mem/memory_reg[46][18]  ( .D(\Data_Mem/n6275 ), .CLK(clk), .RST(
        rst), .I(e_init[1490]), .Q(o[1490]) );
  DFF \Data_Mem/memory_reg[46][19]  ( .D(\Data_Mem/n6276 ), .CLK(clk), .RST(
        rst), .I(e_init[1491]), .Q(o[1491]) );
  DFF \Data_Mem/memory_reg[46][20]  ( .D(\Data_Mem/n6277 ), .CLK(clk), .RST(
        rst), .I(e_init[1492]), .Q(o[1492]) );
  DFF \Data_Mem/memory_reg[46][21]  ( .D(\Data_Mem/n6278 ), .CLK(clk), .RST(
        rst), .I(e_init[1493]), .Q(o[1493]) );
  DFF \Data_Mem/memory_reg[46][22]  ( .D(\Data_Mem/n6279 ), .CLK(clk), .RST(
        rst), .I(e_init[1494]), .Q(o[1494]) );
  DFF \Data_Mem/memory_reg[46][23]  ( .D(\Data_Mem/n6280 ), .CLK(clk), .RST(
        rst), .I(e_init[1495]), .Q(o[1495]) );
  DFF \Data_Mem/memory_reg[46][24]  ( .D(\Data_Mem/n6281 ), .CLK(clk), .RST(
        rst), .I(e_init[1496]), .Q(o[1496]) );
  DFF \Data_Mem/memory_reg[46][25]  ( .D(\Data_Mem/n6282 ), .CLK(clk), .RST(
        rst), .I(e_init[1497]), .Q(o[1497]) );
  DFF \Data_Mem/memory_reg[46][26]  ( .D(\Data_Mem/n6283 ), .CLK(clk), .RST(
        rst), .I(e_init[1498]), .Q(o[1498]) );
  DFF \Data_Mem/memory_reg[46][27]  ( .D(\Data_Mem/n6284 ), .CLK(clk), .RST(
        rst), .I(e_init[1499]), .Q(o[1499]) );
  DFF \Data_Mem/memory_reg[46][28]  ( .D(\Data_Mem/n6285 ), .CLK(clk), .RST(
        rst), .I(e_init[1500]), .Q(o[1500]) );
  DFF \Data_Mem/memory_reg[46][29]  ( .D(\Data_Mem/n6286 ), .CLK(clk), .RST(
        rst), .I(e_init[1501]), .Q(o[1501]) );
  DFF \Data_Mem/memory_reg[46][30]  ( .D(\Data_Mem/n6287 ), .CLK(clk), .RST(
        rst), .I(e_init[1502]), .Q(o[1502]) );
  DFF \Data_Mem/memory_reg[46][31]  ( .D(\Data_Mem/n6288 ), .CLK(clk), .RST(
        rst), .I(e_init[1503]), .Q(o[1503]) );
  DFF \Data_Mem/memory_reg[45][0]  ( .D(\Data_Mem/n6289 ), .CLK(clk), .RST(rst), .I(e_init[1440]), .Q(o[1440]) );
  DFF \Data_Mem/memory_reg[45][1]  ( .D(\Data_Mem/n6290 ), .CLK(clk), .RST(rst), .I(e_init[1441]), .Q(o[1441]) );
  DFF \Data_Mem/memory_reg[45][2]  ( .D(\Data_Mem/n6291 ), .CLK(clk), .RST(rst), .I(e_init[1442]), .Q(o[1442]) );
  DFF \Data_Mem/memory_reg[45][3]  ( .D(\Data_Mem/n6292 ), .CLK(clk), .RST(rst), .I(e_init[1443]), .Q(o[1443]) );
  DFF \Data_Mem/memory_reg[45][4]  ( .D(\Data_Mem/n6293 ), .CLK(clk), .RST(rst), .I(e_init[1444]), .Q(o[1444]) );
  DFF \Data_Mem/memory_reg[45][5]  ( .D(\Data_Mem/n6294 ), .CLK(clk), .RST(rst), .I(e_init[1445]), .Q(o[1445]) );
  DFF \Data_Mem/memory_reg[45][6]  ( .D(\Data_Mem/n6295 ), .CLK(clk), .RST(rst), .I(e_init[1446]), .Q(o[1446]) );
  DFF \Data_Mem/memory_reg[45][7]  ( .D(\Data_Mem/n6296 ), .CLK(clk), .RST(rst), .I(e_init[1447]), .Q(o[1447]) );
  DFF \Data_Mem/memory_reg[45][8]  ( .D(\Data_Mem/n6297 ), .CLK(clk), .RST(rst), .I(e_init[1448]), .Q(o[1448]) );
  DFF \Data_Mem/memory_reg[45][9]  ( .D(\Data_Mem/n6298 ), .CLK(clk), .RST(rst), .I(e_init[1449]), .Q(o[1449]) );
  DFF \Data_Mem/memory_reg[45][10]  ( .D(\Data_Mem/n6299 ), .CLK(clk), .RST(
        rst), .I(e_init[1450]), .Q(o[1450]) );
  DFF \Data_Mem/memory_reg[45][11]  ( .D(\Data_Mem/n6300 ), .CLK(clk), .RST(
        rst), .I(e_init[1451]), .Q(o[1451]) );
  DFF \Data_Mem/memory_reg[45][12]  ( .D(\Data_Mem/n6301 ), .CLK(clk), .RST(
        rst), .I(e_init[1452]), .Q(o[1452]) );
  DFF \Data_Mem/memory_reg[45][13]  ( .D(\Data_Mem/n6302 ), .CLK(clk), .RST(
        rst), .I(e_init[1453]), .Q(o[1453]) );
  DFF \Data_Mem/memory_reg[45][14]  ( .D(\Data_Mem/n6303 ), .CLK(clk), .RST(
        rst), .I(e_init[1454]), .Q(o[1454]) );
  DFF \Data_Mem/memory_reg[45][15]  ( .D(\Data_Mem/n6304 ), .CLK(clk), .RST(
        rst), .I(e_init[1455]), .Q(o[1455]) );
  DFF \Data_Mem/memory_reg[45][16]  ( .D(\Data_Mem/n6305 ), .CLK(clk), .RST(
        rst), .I(e_init[1456]), .Q(o[1456]) );
  DFF \Data_Mem/memory_reg[45][17]  ( .D(\Data_Mem/n6306 ), .CLK(clk), .RST(
        rst), .I(e_init[1457]), .Q(o[1457]) );
  DFF \Data_Mem/memory_reg[45][18]  ( .D(\Data_Mem/n6307 ), .CLK(clk), .RST(
        rst), .I(e_init[1458]), .Q(o[1458]) );
  DFF \Data_Mem/memory_reg[45][19]  ( .D(\Data_Mem/n6308 ), .CLK(clk), .RST(
        rst), .I(e_init[1459]), .Q(o[1459]) );
  DFF \Data_Mem/memory_reg[45][20]  ( .D(\Data_Mem/n6309 ), .CLK(clk), .RST(
        rst), .I(e_init[1460]), .Q(o[1460]) );
  DFF \Data_Mem/memory_reg[45][21]  ( .D(\Data_Mem/n6310 ), .CLK(clk), .RST(
        rst), .I(e_init[1461]), .Q(o[1461]) );
  DFF \Data_Mem/memory_reg[45][22]  ( .D(\Data_Mem/n6311 ), .CLK(clk), .RST(
        rst), .I(e_init[1462]), .Q(o[1462]) );
  DFF \Data_Mem/memory_reg[45][23]  ( .D(\Data_Mem/n6312 ), .CLK(clk), .RST(
        rst), .I(e_init[1463]), .Q(o[1463]) );
  DFF \Data_Mem/memory_reg[45][24]  ( .D(\Data_Mem/n6313 ), .CLK(clk), .RST(
        rst), .I(e_init[1464]), .Q(o[1464]) );
  DFF \Data_Mem/memory_reg[45][25]  ( .D(\Data_Mem/n6314 ), .CLK(clk), .RST(
        rst), .I(e_init[1465]), .Q(o[1465]) );
  DFF \Data_Mem/memory_reg[45][26]  ( .D(\Data_Mem/n6315 ), .CLK(clk), .RST(
        rst), .I(e_init[1466]), .Q(o[1466]) );
  DFF \Data_Mem/memory_reg[45][27]  ( .D(\Data_Mem/n6316 ), .CLK(clk), .RST(
        rst), .I(e_init[1467]), .Q(o[1467]) );
  DFF \Data_Mem/memory_reg[45][28]  ( .D(\Data_Mem/n6317 ), .CLK(clk), .RST(
        rst), .I(e_init[1468]), .Q(o[1468]) );
  DFF \Data_Mem/memory_reg[45][29]  ( .D(\Data_Mem/n6318 ), .CLK(clk), .RST(
        rst), .I(e_init[1469]), .Q(o[1469]) );
  DFF \Data_Mem/memory_reg[45][30]  ( .D(\Data_Mem/n6319 ), .CLK(clk), .RST(
        rst), .I(e_init[1470]), .Q(o[1470]) );
  DFF \Data_Mem/memory_reg[45][31]  ( .D(\Data_Mem/n6320 ), .CLK(clk), .RST(
        rst), .I(e_init[1471]), .Q(o[1471]) );
  DFF \Data_Mem/memory_reg[44][0]  ( .D(\Data_Mem/n6321 ), .CLK(clk), .RST(rst), .I(e_init[1408]), .Q(o[1408]) );
  DFF \Data_Mem/memory_reg[44][1]  ( .D(\Data_Mem/n6322 ), .CLK(clk), .RST(rst), .I(e_init[1409]), .Q(o[1409]) );
  DFF \Data_Mem/memory_reg[44][2]  ( .D(\Data_Mem/n6323 ), .CLK(clk), .RST(rst), .I(e_init[1410]), .Q(o[1410]) );
  DFF \Data_Mem/memory_reg[44][3]  ( .D(\Data_Mem/n6324 ), .CLK(clk), .RST(rst), .I(e_init[1411]), .Q(o[1411]) );
  DFF \Data_Mem/memory_reg[44][4]  ( .D(\Data_Mem/n6325 ), .CLK(clk), .RST(rst), .I(e_init[1412]), .Q(o[1412]) );
  DFF \Data_Mem/memory_reg[44][5]  ( .D(\Data_Mem/n6326 ), .CLK(clk), .RST(rst), .I(e_init[1413]), .Q(o[1413]) );
  DFF \Data_Mem/memory_reg[44][6]  ( .D(\Data_Mem/n6327 ), .CLK(clk), .RST(rst), .I(e_init[1414]), .Q(o[1414]) );
  DFF \Data_Mem/memory_reg[44][7]  ( .D(\Data_Mem/n6328 ), .CLK(clk), .RST(rst), .I(e_init[1415]), .Q(o[1415]) );
  DFF \Data_Mem/memory_reg[44][8]  ( .D(\Data_Mem/n6329 ), .CLK(clk), .RST(rst), .I(e_init[1416]), .Q(o[1416]) );
  DFF \Data_Mem/memory_reg[44][9]  ( .D(\Data_Mem/n6330 ), .CLK(clk), .RST(rst), .I(e_init[1417]), .Q(o[1417]) );
  DFF \Data_Mem/memory_reg[44][10]  ( .D(\Data_Mem/n6331 ), .CLK(clk), .RST(
        rst), .I(e_init[1418]), .Q(o[1418]) );
  DFF \Data_Mem/memory_reg[44][11]  ( .D(\Data_Mem/n6332 ), .CLK(clk), .RST(
        rst), .I(e_init[1419]), .Q(o[1419]) );
  DFF \Data_Mem/memory_reg[44][12]  ( .D(\Data_Mem/n6333 ), .CLK(clk), .RST(
        rst), .I(e_init[1420]), .Q(o[1420]) );
  DFF \Data_Mem/memory_reg[44][13]  ( .D(\Data_Mem/n6334 ), .CLK(clk), .RST(
        rst), .I(e_init[1421]), .Q(o[1421]) );
  DFF \Data_Mem/memory_reg[44][14]  ( .D(\Data_Mem/n6335 ), .CLK(clk), .RST(
        rst), .I(e_init[1422]), .Q(o[1422]) );
  DFF \Data_Mem/memory_reg[44][15]  ( .D(\Data_Mem/n6336 ), .CLK(clk), .RST(
        rst), .I(e_init[1423]), .Q(o[1423]) );
  DFF \Data_Mem/memory_reg[44][16]  ( .D(\Data_Mem/n6337 ), .CLK(clk), .RST(
        rst), .I(e_init[1424]), .Q(o[1424]) );
  DFF \Data_Mem/memory_reg[44][17]  ( .D(\Data_Mem/n6338 ), .CLK(clk), .RST(
        rst), .I(e_init[1425]), .Q(o[1425]) );
  DFF \Data_Mem/memory_reg[44][18]  ( .D(\Data_Mem/n6339 ), .CLK(clk), .RST(
        rst), .I(e_init[1426]), .Q(o[1426]) );
  DFF \Data_Mem/memory_reg[44][19]  ( .D(\Data_Mem/n6340 ), .CLK(clk), .RST(
        rst), .I(e_init[1427]), .Q(o[1427]) );
  DFF \Data_Mem/memory_reg[44][20]  ( .D(\Data_Mem/n6341 ), .CLK(clk), .RST(
        rst), .I(e_init[1428]), .Q(o[1428]) );
  DFF \Data_Mem/memory_reg[44][21]  ( .D(\Data_Mem/n6342 ), .CLK(clk), .RST(
        rst), .I(e_init[1429]), .Q(o[1429]) );
  DFF \Data_Mem/memory_reg[44][22]  ( .D(\Data_Mem/n6343 ), .CLK(clk), .RST(
        rst), .I(e_init[1430]), .Q(o[1430]) );
  DFF \Data_Mem/memory_reg[44][23]  ( .D(\Data_Mem/n6344 ), .CLK(clk), .RST(
        rst), .I(e_init[1431]), .Q(o[1431]) );
  DFF \Data_Mem/memory_reg[44][24]  ( .D(\Data_Mem/n6345 ), .CLK(clk), .RST(
        rst), .I(e_init[1432]), .Q(o[1432]) );
  DFF \Data_Mem/memory_reg[44][25]  ( .D(\Data_Mem/n6346 ), .CLK(clk), .RST(
        rst), .I(e_init[1433]), .Q(o[1433]) );
  DFF \Data_Mem/memory_reg[44][26]  ( .D(\Data_Mem/n6347 ), .CLK(clk), .RST(
        rst), .I(e_init[1434]), .Q(o[1434]) );
  DFF \Data_Mem/memory_reg[44][27]  ( .D(\Data_Mem/n6348 ), .CLK(clk), .RST(
        rst), .I(e_init[1435]), .Q(o[1435]) );
  DFF \Data_Mem/memory_reg[44][28]  ( .D(\Data_Mem/n6349 ), .CLK(clk), .RST(
        rst), .I(e_init[1436]), .Q(o[1436]) );
  DFF \Data_Mem/memory_reg[44][29]  ( .D(\Data_Mem/n6350 ), .CLK(clk), .RST(
        rst), .I(e_init[1437]), .Q(o[1437]) );
  DFF \Data_Mem/memory_reg[44][30]  ( .D(\Data_Mem/n6351 ), .CLK(clk), .RST(
        rst), .I(e_init[1438]), .Q(o[1438]) );
  DFF \Data_Mem/memory_reg[44][31]  ( .D(\Data_Mem/n6352 ), .CLK(clk), .RST(
        rst), .I(e_init[1439]), .Q(o[1439]) );
  DFF \Data_Mem/memory_reg[43][0]  ( .D(\Data_Mem/n6353 ), .CLK(clk), .RST(rst), .I(e_init[1376]), .Q(o[1376]) );
  DFF \Data_Mem/memory_reg[43][1]  ( .D(\Data_Mem/n6354 ), .CLK(clk), .RST(rst), .I(e_init[1377]), .Q(o[1377]) );
  DFF \Data_Mem/memory_reg[43][2]  ( .D(\Data_Mem/n6355 ), .CLK(clk), .RST(rst), .I(e_init[1378]), .Q(o[1378]) );
  DFF \Data_Mem/memory_reg[43][3]  ( .D(\Data_Mem/n6356 ), .CLK(clk), .RST(rst), .I(e_init[1379]), .Q(o[1379]) );
  DFF \Data_Mem/memory_reg[43][4]  ( .D(\Data_Mem/n6357 ), .CLK(clk), .RST(rst), .I(e_init[1380]), .Q(o[1380]) );
  DFF \Data_Mem/memory_reg[43][5]  ( .D(\Data_Mem/n6358 ), .CLK(clk), .RST(rst), .I(e_init[1381]), .Q(o[1381]) );
  DFF \Data_Mem/memory_reg[43][6]  ( .D(\Data_Mem/n6359 ), .CLK(clk), .RST(rst), .I(e_init[1382]), .Q(o[1382]) );
  DFF \Data_Mem/memory_reg[43][7]  ( .D(\Data_Mem/n6360 ), .CLK(clk), .RST(rst), .I(e_init[1383]), .Q(o[1383]) );
  DFF \Data_Mem/memory_reg[43][8]  ( .D(\Data_Mem/n6361 ), .CLK(clk), .RST(rst), .I(e_init[1384]), .Q(o[1384]) );
  DFF \Data_Mem/memory_reg[43][9]  ( .D(\Data_Mem/n6362 ), .CLK(clk), .RST(rst), .I(e_init[1385]), .Q(o[1385]) );
  DFF \Data_Mem/memory_reg[43][10]  ( .D(\Data_Mem/n6363 ), .CLK(clk), .RST(
        rst), .I(e_init[1386]), .Q(o[1386]) );
  DFF \Data_Mem/memory_reg[43][11]  ( .D(\Data_Mem/n6364 ), .CLK(clk), .RST(
        rst), .I(e_init[1387]), .Q(o[1387]) );
  DFF \Data_Mem/memory_reg[43][12]  ( .D(\Data_Mem/n6365 ), .CLK(clk), .RST(
        rst), .I(e_init[1388]), .Q(o[1388]) );
  DFF \Data_Mem/memory_reg[43][13]  ( .D(\Data_Mem/n6366 ), .CLK(clk), .RST(
        rst), .I(e_init[1389]), .Q(o[1389]) );
  DFF \Data_Mem/memory_reg[43][14]  ( .D(\Data_Mem/n6367 ), .CLK(clk), .RST(
        rst), .I(e_init[1390]), .Q(o[1390]) );
  DFF \Data_Mem/memory_reg[43][15]  ( .D(\Data_Mem/n6368 ), .CLK(clk), .RST(
        rst), .I(e_init[1391]), .Q(o[1391]) );
  DFF \Data_Mem/memory_reg[43][16]  ( .D(\Data_Mem/n6369 ), .CLK(clk), .RST(
        rst), .I(e_init[1392]), .Q(o[1392]) );
  DFF \Data_Mem/memory_reg[43][17]  ( .D(\Data_Mem/n6370 ), .CLK(clk), .RST(
        rst), .I(e_init[1393]), .Q(o[1393]) );
  DFF \Data_Mem/memory_reg[43][18]  ( .D(\Data_Mem/n6371 ), .CLK(clk), .RST(
        rst), .I(e_init[1394]), .Q(o[1394]) );
  DFF \Data_Mem/memory_reg[43][19]  ( .D(\Data_Mem/n6372 ), .CLK(clk), .RST(
        rst), .I(e_init[1395]), .Q(o[1395]) );
  DFF \Data_Mem/memory_reg[43][20]  ( .D(\Data_Mem/n6373 ), .CLK(clk), .RST(
        rst), .I(e_init[1396]), .Q(o[1396]) );
  DFF \Data_Mem/memory_reg[43][21]  ( .D(\Data_Mem/n6374 ), .CLK(clk), .RST(
        rst), .I(e_init[1397]), .Q(o[1397]) );
  DFF \Data_Mem/memory_reg[43][22]  ( .D(\Data_Mem/n6375 ), .CLK(clk), .RST(
        rst), .I(e_init[1398]), .Q(o[1398]) );
  DFF \Data_Mem/memory_reg[43][23]  ( .D(\Data_Mem/n6376 ), .CLK(clk), .RST(
        rst), .I(e_init[1399]), .Q(o[1399]) );
  DFF \Data_Mem/memory_reg[43][24]  ( .D(\Data_Mem/n6377 ), .CLK(clk), .RST(
        rst), .I(e_init[1400]), .Q(o[1400]) );
  DFF \Data_Mem/memory_reg[43][25]  ( .D(\Data_Mem/n6378 ), .CLK(clk), .RST(
        rst), .I(e_init[1401]), .Q(o[1401]) );
  DFF \Data_Mem/memory_reg[43][26]  ( .D(\Data_Mem/n6379 ), .CLK(clk), .RST(
        rst), .I(e_init[1402]), .Q(o[1402]) );
  DFF \Data_Mem/memory_reg[43][27]  ( .D(\Data_Mem/n6380 ), .CLK(clk), .RST(
        rst), .I(e_init[1403]), .Q(o[1403]) );
  DFF \Data_Mem/memory_reg[43][28]  ( .D(\Data_Mem/n6381 ), .CLK(clk), .RST(
        rst), .I(e_init[1404]), .Q(o[1404]) );
  DFF \Data_Mem/memory_reg[43][29]  ( .D(\Data_Mem/n6382 ), .CLK(clk), .RST(
        rst), .I(e_init[1405]), .Q(o[1405]) );
  DFF \Data_Mem/memory_reg[43][30]  ( .D(\Data_Mem/n6383 ), .CLK(clk), .RST(
        rst), .I(e_init[1406]), .Q(o[1406]) );
  DFF \Data_Mem/memory_reg[43][31]  ( .D(\Data_Mem/n6384 ), .CLK(clk), .RST(
        rst), .I(e_init[1407]), .Q(o[1407]) );
  DFF \Data_Mem/memory_reg[42][0]  ( .D(\Data_Mem/n6385 ), .CLK(clk), .RST(rst), .I(e_init[1344]), .Q(o[1344]) );
  DFF \Data_Mem/memory_reg[42][1]  ( .D(\Data_Mem/n6386 ), .CLK(clk), .RST(rst), .I(e_init[1345]), .Q(o[1345]) );
  DFF \Data_Mem/memory_reg[42][2]  ( .D(\Data_Mem/n6387 ), .CLK(clk), .RST(rst), .I(e_init[1346]), .Q(o[1346]) );
  DFF \Data_Mem/memory_reg[42][3]  ( .D(\Data_Mem/n6388 ), .CLK(clk), .RST(rst), .I(e_init[1347]), .Q(o[1347]) );
  DFF \Data_Mem/memory_reg[42][4]  ( .D(\Data_Mem/n6389 ), .CLK(clk), .RST(rst), .I(e_init[1348]), .Q(o[1348]) );
  DFF \Data_Mem/memory_reg[42][5]  ( .D(\Data_Mem/n6390 ), .CLK(clk), .RST(rst), .I(e_init[1349]), .Q(o[1349]) );
  DFF \Data_Mem/memory_reg[42][6]  ( .D(\Data_Mem/n6391 ), .CLK(clk), .RST(rst), .I(e_init[1350]), .Q(o[1350]) );
  DFF \Data_Mem/memory_reg[42][7]  ( .D(\Data_Mem/n6392 ), .CLK(clk), .RST(rst), .I(e_init[1351]), .Q(o[1351]) );
  DFF \Data_Mem/memory_reg[42][8]  ( .D(\Data_Mem/n6393 ), .CLK(clk), .RST(rst), .I(e_init[1352]), .Q(o[1352]) );
  DFF \Data_Mem/memory_reg[42][9]  ( .D(\Data_Mem/n6394 ), .CLK(clk), .RST(rst), .I(e_init[1353]), .Q(o[1353]) );
  DFF \Data_Mem/memory_reg[42][10]  ( .D(\Data_Mem/n6395 ), .CLK(clk), .RST(
        rst), .I(e_init[1354]), .Q(o[1354]) );
  DFF \Data_Mem/memory_reg[42][11]  ( .D(\Data_Mem/n6396 ), .CLK(clk), .RST(
        rst), .I(e_init[1355]), .Q(o[1355]) );
  DFF \Data_Mem/memory_reg[42][12]  ( .D(\Data_Mem/n6397 ), .CLK(clk), .RST(
        rst), .I(e_init[1356]), .Q(o[1356]) );
  DFF \Data_Mem/memory_reg[42][13]  ( .D(\Data_Mem/n6398 ), .CLK(clk), .RST(
        rst), .I(e_init[1357]), .Q(o[1357]) );
  DFF \Data_Mem/memory_reg[42][14]  ( .D(\Data_Mem/n6399 ), .CLK(clk), .RST(
        rst), .I(e_init[1358]), .Q(o[1358]) );
  DFF \Data_Mem/memory_reg[42][15]  ( .D(\Data_Mem/n6400 ), .CLK(clk), .RST(
        rst), .I(e_init[1359]), .Q(o[1359]) );
  DFF \Data_Mem/memory_reg[42][16]  ( .D(\Data_Mem/n6401 ), .CLK(clk), .RST(
        rst), .I(e_init[1360]), .Q(o[1360]) );
  DFF \Data_Mem/memory_reg[42][17]  ( .D(\Data_Mem/n6402 ), .CLK(clk), .RST(
        rst), .I(e_init[1361]), .Q(o[1361]) );
  DFF \Data_Mem/memory_reg[42][18]  ( .D(\Data_Mem/n6403 ), .CLK(clk), .RST(
        rst), .I(e_init[1362]), .Q(o[1362]) );
  DFF \Data_Mem/memory_reg[42][19]  ( .D(\Data_Mem/n6404 ), .CLK(clk), .RST(
        rst), .I(e_init[1363]), .Q(o[1363]) );
  DFF \Data_Mem/memory_reg[42][20]  ( .D(\Data_Mem/n6405 ), .CLK(clk), .RST(
        rst), .I(e_init[1364]), .Q(o[1364]) );
  DFF \Data_Mem/memory_reg[42][21]  ( .D(\Data_Mem/n6406 ), .CLK(clk), .RST(
        rst), .I(e_init[1365]), .Q(o[1365]) );
  DFF \Data_Mem/memory_reg[42][22]  ( .D(\Data_Mem/n6407 ), .CLK(clk), .RST(
        rst), .I(e_init[1366]), .Q(o[1366]) );
  DFF \Data_Mem/memory_reg[42][23]  ( .D(\Data_Mem/n6408 ), .CLK(clk), .RST(
        rst), .I(e_init[1367]), .Q(o[1367]) );
  DFF \Data_Mem/memory_reg[42][24]  ( .D(\Data_Mem/n6409 ), .CLK(clk), .RST(
        rst), .I(e_init[1368]), .Q(o[1368]) );
  DFF \Data_Mem/memory_reg[42][25]  ( .D(\Data_Mem/n6410 ), .CLK(clk), .RST(
        rst), .I(e_init[1369]), .Q(o[1369]) );
  DFF \Data_Mem/memory_reg[42][26]  ( .D(\Data_Mem/n6411 ), .CLK(clk), .RST(
        rst), .I(e_init[1370]), .Q(o[1370]) );
  DFF \Data_Mem/memory_reg[42][27]  ( .D(\Data_Mem/n6412 ), .CLK(clk), .RST(
        rst), .I(e_init[1371]), .Q(o[1371]) );
  DFF \Data_Mem/memory_reg[42][28]  ( .D(\Data_Mem/n6413 ), .CLK(clk), .RST(
        rst), .I(e_init[1372]), .Q(o[1372]) );
  DFF \Data_Mem/memory_reg[42][29]  ( .D(\Data_Mem/n6414 ), .CLK(clk), .RST(
        rst), .I(e_init[1373]), .Q(o[1373]) );
  DFF \Data_Mem/memory_reg[42][30]  ( .D(\Data_Mem/n6415 ), .CLK(clk), .RST(
        rst), .I(e_init[1374]), .Q(o[1374]) );
  DFF \Data_Mem/memory_reg[42][31]  ( .D(\Data_Mem/n6416 ), .CLK(clk), .RST(
        rst), .I(e_init[1375]), .Q(o[1375]) );
  DFF \Data_Mem/memory_reg[41][0]  ( .D(\Data_Mem/n6417 ), .CLK(clk), .RST(rst), .I(e_init[1312]), .Q(o[1312]) );
  DFF \Data_Mem/memory_reg[41][1]  ( .D(\Data_Mem/n6418 ), .CLK(clk), .RST(rst), .I(e_init[1313]), .Q(o[1313]) );
  DFF \Data_Mem/memory_reg[41][2]  ( .D(\Data_Mem/n6419 ), .CLK(clk), .RST(rst), .I(e_init[1314]), .Q(o[1314]) );
  DFF \Data_Mem/memory_reg[41][3]  ( .D(\Data_Mem/n6420 ), .CLK(clk), .RST(rst), .I(e_init[1315]), .Q(o[1315]) );
  DFF \Data_Mem/memory_reg[41][4]  ( .D(\Data_Mem/n6421 ), .CLK(clk), .RST(rst), .I(e_init[1316]), .Q(o[1316]) );
  DFF \Data_Mem/memory_reg[41][5]  ( .D(\Data_Mem/n6422 ), .CLK(clk), .RST(rst), .I(e_init[1317]), .Q(o[1317]) );
  DFF \Data_Mem/memory_reg[41][6]  ( .D(\Data_Mem/n6423 ), .CLK(clk), .RST(rst), .I(e_init[1318]), .Q(o[1318]) );
  DFF \Data_Mem/memory_reg[41][7]  ( .D(\Data_Mem/n6424 ), .CLK(clk), .RST(rst), .I(e_init[1319]), .Q(o[1319]) );
  DFF \Data_Mem/memory_reg[41][8]  ( .D(\Data_Mem/n6425 ), .CLK(clk), .RST(rst), .I(e_init[1320]), .Q(o[1320]) );
  DFF \Data_Mem/memory_reg[41][9]  ( .D(\Data_Mem/n6426 ), .CLK(clk), .RST(rst), .I(e_init[1321]), .Q(o[1321]) );
  DFF \Data_Mem/memory_reg[41][10]  ( .D(\Data_Mem/n6427 ), .CLK(clk), .RST(
        rst), .I(e_init[1322]), .Q(o[1322]) );
  DFF \Data_Mem/memory_reg[41][11]  ( .D(\Data_Mem/n6428 ), .CLK(clk), .RST(
        rst), .I(e_init[1323]), .Q(o[1323]) );
  DFF \Data_Mem/memory_reg[41][12]  ( .D(\Data_Mem/n6429 ), .CLK(clk), .RST(
        rst), .I(e_init[1324]), .Q(o[1324]) );
  DFF \Data_Mem/memory_reg[41][13]  ( .D(\Data_Mem/n6430 ), .CLK(clk), .RST(
        rst), .I(e_init[1325]), .Q(o[1325]) );
  DFF \Data_Mem/memory_reg[41][14]  ( .D(\Data_Mem/n6431 ), .CLK(clk), .RST(
        rst), .I(e_init[1326]), .Q(o[1326]) );
  DFF \Data_Mem/memory_reg[41][15]  ( .D(\Data_Mem/n6432 ), .CLK(clk), .RST(
        rst), .I(e_init[1327]), .Q(o[1327]) );
  DFF \Data_Mem/memory_reg[41][16]  ( .D(\Data_Mem/n6433 ), .CLK(clk), .RST(
        rst), .I(e_init[1328]), .Q(o[1328]) );
  DFF \Data_Mem/memory_reg[41][17]  ( .D(\Data_Mem/n6434 ), .CLK(clk), .RST(
        rst), .I(e_init[1329]), .Q(o[1329]) );
  DFF \Data_Mem/memory_reg[41][18]  ( .D(\Data_Mem/n6435 ), .CLK(clk), .RST(
        rst), .I(e_init[1330]), .Q(o[1330]) );
  DFF \Data_Mem/memory_reg[41][19]  ( .D(\Data_Mem/n6436 ), .CLK(clk), .RST(
        rst), .I(e_init[1331]), .Q(o[1331]) );
  DFF \Data_Mem/memory_reg[41][20]  ( .D(\Data_Mem/n6437 ), .CLK(clk), .RST(
        rst), .I(e_init[1332]), .Q(o[1332]) );
  DFF \Data_Mem/memory_reg[41][21]  ( .D(\Data_Mem/n6438 ), .CLK(clk), .RST(
        rst), .I(e_init[1333]), .Q(o[1333]) );
  DFF \Data_Mem/memory_reg[41][22]  ( .D(\Data_Mem/n6439 ), .CLK(clk), .RST(
        rst), .I(e_init[1334]), .Q(o[1334]) );
  DFF \Data_Mem/memory_reg[41][23]  ( .D(\Data_Mem/n6440 ), .CLK(clk), .RST(
        rst), .I(e_init[1335]), .Q(o[1335]) );
  DFF \Data_Mem/memory_reg[41][24]  ( .D(\Data_Mem/n6441 ), .CLK(clk), .RST(
        rst), .I(e_init[1336]), .Q(o[1336]) );
  DFF \Data_Mem/memory_reg[41][25]  ( .D(\Data_Mem/n6442 ), .CLK(clk), .RST(
        rst), .I(e_init[1337]), .Q(o[1337]) );
  DFF \Data_Mem/memory_reg[41][26]  ( .D(\Data_Mem/n6443 ), .CLK(clk), .RST(
        rst), .I(e_init[1338]), .Q(o[1338]) );
  DFF \Data_Mem/memory_reg[41][27]  ( .D(\Data_Mem/n6444 ), .CLK(clk), .RST(
        rst), .I(e_init[1339]), .Q(o[1339]) );
  DFF \Data_Mem/memory_reg[41][28]  ( .D(\Data_Mem/n6445 ), .CLK(clk), .RST(
        rst), .I(e_init[1340]), .Q(o[1340]) );
  DFF \Data_Mem/memory_reg[41][29]  ( .D(\Data_Mem/n6446 ), .CLK(clk), .RST(
        rst), .I(e_init[1341]), .Q(o[1341]) );
  DFF \Data_Mem/memory_reg[41][30]  ( .D(\Data_Mem/n6447 ), .CLK(clk), .RST(
        rst), .I(e_init[1342]), .Q(o[1342]) );
  DFF \Data_Mem/memory_reg[41][31]  ( .D(\Data_Mem/n6448 ), .CLK(clk), .RST(
        rst), .I(e_init[1343]), .Q(o[1343]) );
  DFF \Data_Mem/memory_reg[40][0]  ( .D(\Data_Mem/n6449 ), .CLK(clk), .RST(rst), .I(e_init[1280]), .Q(o[1280]) );
  DFF \Data_Mem/memory_reg[40][1]  ( .D(\Data_Mem/n6450 ), .CLK(clk), .RST(rst), .I(e_init[1281]), .Q(o[1281]) );
  DFF \Data_Mem/memory_reg[40][2]  ( .D(\Data_Mem/n6451 ), .CLK(clk), .RST(rst), .I(e_init[1282]), .Q(o[1282]) );
  DFF \Data_Mem/memory_reg[40][3]  ( .D(\Data_Mem/n6452 ), .CLK(clk), .RST(rst), .I(e_init[1283]), .Q(o[1283]) );
  DFF \Data_Mem/memory_reg[40][4]  ( .D(\Data_Mem/n6453 ), .CLK(clk), .RST(rst), .I(e_init[1284]), .Q(o[1284]) );
  DFF \Data_Mem/memory_reg[40][5]  ( .D(\Data_Mem/n6454 ), .CLK(clk), .RST(rst), .I(e_init[1285]), .Q(o[1285]) );
  DFF \Data_Mem/memory_reg[40][6]  ( .D(\Data_Mem/n6455 ), .CLK(clk), .RST(rst), .I(e_init[1286]), .Q(o[1286]) );
  DFF \Data_Mem/memory_reg[40][7]  ( .D(\Data_Mem/n6456 ), .CLK(clk), .RST(rst), .I(e_init[1287]), .Q(o[1287]) );
  DFF \Data_Mem/memory_reg[40][8]  ( .D(\Data_Mem/n6457 ), .CLK(clk), .RST(rst), .I(e_init[1288]), .Q(o[1288]) );
  DFF \Data_Mem/memory_reg[40][9]  ( .D(\Data_Mem/n6458 ), .CLK(clk), .RST(rst), .I(e_init[1289]), .Q(o[1289]) );
  DFF \Data_Mem/memory_reg[40][10]  ( .D(\Data_Mem/n6459 ), .CLK(clk), .RST(
        rst), .I(e_init[1290]), .Q(o[1290]) );
  DFF \Data_Mem/memory_reg[40][11]  ( .D(\Data_Mem/n6460 ), .CLK(clk), .RST(
        rst), .I(e_init[1291]), .Q(o[1291]) );
  DFF \Data_Mem/memory_reg[40][12]  ( .D(\Data_Mem/n6461 ), .CLK(clk), .RST(
        rst), .I(e_init[1292]), .Q(o[1292]) );
  DFF \Data_Mem/memory_reg[40][13]  ( .D(\Data_Mem/n6462 ), .CLK(clk), .RST(
        rst), .I(e_init[1293]), .Q(o[1293]) );
  DFF \Data_Mem/memory_reg[40][14]  ( .D(\Data_Mem/n6463 ), .CLK(clk), .RST(
        rst), .I(e_init[1294]), .Q(o[1294]) );
  DFF \Data_Mem/memory_reg[40][15]  ( .D(\Data_Mem/n6464 ), .CLK(clk), .RST(
        rst), .I(e_init[1295]), .Q(o[1295]) );
  DFF \Data_Mem/memory_reg[40][16]  ( .D(\Data_Mem/n6465 ), .CLK(clk), .RST(
        rst), .I(e_init[1296]), .Q(o[1296]) );
  DFF \Data_Mem/memory_reg[40][17]  ( .D(\Data_Mem/n6466 ), .CLK(clk), .RST(
        rst), .I(e_init[1297]), .Q(o[1297]) );
  DFF \Data_Mem/memory_reg[40][18]  ( .D(\Data_Mem/n6467 ), .CLK(clk), .RST(
        rst), .I(e_init[1298]), .Q(o[1298]) );
  DFF \Data_Mem/memory_reg[40][19]  ( .D(\Data_Mem/n6468 ), .CLK(clk), .RST(
        rst), .I(e_init[1299]), .Q(o[1299]) );
  DFF \Data_Mem/memory_reg[40][20]  ( .D(\Data_Mem/n6469 ), .CLK(clk), .RST(
        rst), .I(e_init[1300]), .Q(o[1300]) );
  DFF \Data_Mem/memory_reg[40][21]  ( .D(\Data_Mem/n6470 ), .CLK(clk), .RST(
        rst), .I(e_init[1301]), .Q(o[1301]) );
  DFF \Data_Mem/memory_reg[40][22]  ( .D(\Data_Mem/n6471 ), .CLK(clk), .RST(
        rst), .I(e_init[1302]), .Q(o[1302]) );
  DFF \Data_Mem/memory_reg[40][23]  ( .D(\Data_Mem/n6472 ), .CLK(clk), .RST(
        rst), .I(e_init[1303]), .Q(o[1303]) );
  DFF \Data_Mem/memory_reg[40][24]  ( .D(\Data_Mem/n6473 ), .CLK(clk), .RST(
        rst), .I(e_init[1304]), .Q(o[1304]) );
  DFF \Data_Mem/memory_reg[40][25]  ( .D(\Data_Mem/n6474 ), .CLK(clk), .RST(
        rst), .I(e_init[1305]), .Q(o[1305]) );
  DFF \Data_Mem/memory_reg[40][26]  ( .D(\Data_Mem/n6475 ), .CLK(clk), .RST(
        rst), .I(e_init[1306]), .Q(o[1306]) );
  DFF \Data_Mem/memory_reg[40][27]  ( .D(\Data_Mem/n6476 ), .CLK(clk), .RST(
        rst), .I(e_init[1307]), .Q(o[1307]) );
  DFF \Data_Mem/memory_reg[40][28]  ( .D(\Data_Mem/n6477 ), .CLK(clk), .RST(
        rst), .I(e_init[1308]), .Q(o[1308]) );
  DFF \Data_Mem/memory_reg[40][29]  ( .D(\Data_Mem/n6478 ), .CLK(clk), .RST(
        rst), .I(e_init[1309]), .Q(o[1309]) );
  DFF \Data_Mem/memory_reg[40][30]  ( .D(\Data_Mem/n6479 ), .CLK(clk), .RST(
        rst), .I(e_init[1310]), .Q(o[1310]) );
  DFF \Data_Mem/memory_reg[40][31]  ( .D(\Data_Mem/n6480 ), .CLK(clk), .RST(
        rst), .I(e_init[1311]), .Q(o[1311]) );
  DFF \Data_Mem/memory_reg[39][0]  ( .D(\Data_Mem/n6481 ), .CLK(clk), .RST(rst), .I(e_init[1248]), .Q(o[1248]) );
  DFF \Data_Mem/memory_reg[39][1]  ( .D(\Data_Mem/n6482 ), .CLK(clk), .RST(rst), .I(e_init[1249]), .Q(o[1249]) );
  DFF \Data_Mem/memory_reg[39][2]  ( .D(\Data_Mem/n6483 ), .CLK(clk), .RST(rst), .I(e_init[1250]), .Q(o[1250]) );
  DFF \Data_Mem/memory_reg[39][3]  ( .D(\Data_Mem/n6484 ), .CLK(clk), .RST(rst), .I(e_init[1251]), .Q(o[1251]) );
  DFF \Data_Mem/memory_reg[39][4]  ( .D(\Data_Mem/n6485 ), .CLK(clk), .RST(rst), .I(e_init[1252]), .Q(o[1252]) );
  DFF \Data_Mem/memory_reg[39][5]  ( .D(\Data_Mem/n6486 ), .CLK(clk), .RST(rst), .I(e_init[1253]), .Q(o[1253]) );
  DFF \Data_Mem/memory_reg[39][6]  ( .D(\Data_Mem/n6487 ), .CLK(clk), .RST(rst), .I(e_init[1254]), .Q(o[1254]) );
  DFF \Data_Mem/memory_reg[39][7]  ( .D(\Data_Mem/n6488 ), .CLK(clk), .RST(rst), .I(e_init[1255]), .Q(o[1255]) );
  DFF \Data_Mem/memory_reg[39][8]  ( .D(\Data_Mem/n6489 ), .CLK(clk), .RST(rst), .I(e_init[1256]), .Q(o[1256]) );
  DFF \Data_Mem/memory_reg[39][9]  ( .D(\Data_Mem/n6490 ), .CLK(clk), .RST(rst), .I(e_init[1257]), .Q(o[1257]) );
  DFF \Data_Mem/memory_reg[39][10]  ( .D(\Data_Mem/n6491 ), .CLK(clk), .RST(
        rst), .I(e_init[1258]), .Q(o[1258]) );
  DFF \Data_Mem/memory_reg[39][11]  ( .D(\Data_Mem/n6492 ), .CLK(clk), .RST(
        rst), .I(e_init[1259]), .Q(o[1259]) );
  DFF \Data_Mem/memory_reg[39][12]  ( .D(\Data_Mem/n6493 ), .CLK(clk), .RST(
        rst), .I(e_init[1260]), .Q(o[1260]) );
  DFF \Data_Mem/memory_reg[39][13]  ( .D(\Data_Mem/n6494 ), .CLK(clk), .RST(
        rst), .I(e_init[1261]), .Q(o[1261]) );
  DFF \Data_Mem/memory_reg[39][14]  ( .D(\Data_Mem/n6495 ), .CLK(clk), .RST(
        rst), .I(e_init[1262]), .Q(o[1262]) );
  DFF \Data_Mem/memory_reg[39][15]  ( .D(\Data_Mem/n6496 ), .CLK(clk), .RST(
        rst), .I(e_init[1263]), .Q(o[1263]) );
  DFF \Data_Mem/memory_reg[39][16]  ( .D(\Data_Mem/n6497 ), .CLK(clk), .RST(
        rst), .I(e_init[1264]), .Q(o[1264]) );
  DFF \Data_Mem/memory_reg[39][17]  ( .D(\Data_Mem/n6498 ), .CLK(clk), .RST(
        rst), .I(e_init[1265]), .Q(o[1265]) );
  DFF \Data_Mem/memory_reg[39][18]  ( .D(\Data_Mem/n6499 ), .CLK(clk), .RST(
        rst), .I(e_init[1266]), .Q(o[1266]) );
  DFF \Data_Mem/memory_reg[39][19]  ( .D(\Data_Mem/n6500 ), .CLK(clk), .RST(
        rst), .I(e_init[1267]), .Q(o[1267]) );
  DFF \Data_Mem/memory_reg[39][20]  ( .D(\Data_Mem/n6501 ), .CLK(clk), .RST(
        rst), .I(e_init[1268]), .Q(o[1268]) );
  DFF \Data_Mem/memory_reg[39][21]  ( .D(\Data_Mem/n6502 ), .CLK(clk), .RST(
        rst), .I(e_init[1269]), .Q(o[1269]) );
  DFF \Data_Mem/memory_reg[39][22]  ( .D(\Data_Mem/n6503 ), .CLK(clk), .RST(
        rst), .I(e_init[1270]), .Q(o[1270]) );
  DFF \Data_Mem/memory_reg[39][23]  ( .D(\Data_Mem/n6504 ), .CLK(clk), .RST(
        rst), .I(e_init[1271]), .Q(o[1271]) );
  DFF \Data_Mem/memory_reg[39][24]  ( .D(\Data_Mem/n6505 ), .CLK(clk), .RST(
        rst), .I(e_init[1272]), .Q(o[1272]) );
  DFF \Data_Mem/memory_reg[39][25]  ( .D(\Data_Mem/n6506 ), .CLK(clk), .RST(
        rst), .I(e_init[1273]), .Q(o[1273]) );
  DFF \Data_Mem/memory_reg[39][26]  ( .D(\Data_Mem/n6507 ), .CLK(clk), .RST(
        rst), .I(e_init[1274]), .Q(o[1274]) );
  DFF \Data_Mem/memory_reg[39][27]  ( .D(\Data_Mem/n6508 ), .CLK(clk), .RST(
        rst), .I(e_init[1275]), .Q(o[1275]) );
  DFF \Data_Mem/memory_reg[39][28]  ( .D(\Data_Mem/n6509 ), .CLK(clk), .RST(
        rst), .I(e_init[1276]), .Q(o[1276]) );
  DFF \Data_Mem/memory_reg[39][29]  ( .D(\Data_Mem/n6510 ), .CLK(clk), .RST(
        rst), .I(e_init[1277]), .Q(o[1277]) );
  DFF \Data_Mem/memory_reg[39][30]  ( .D(\Data_Mem/n6511 ), .CLK(clk), .RST(
        rst), .I(e_init[1278]), .Q(o[1278]) );
  DFF \Data_Mem/memory_reg[39][31]  ( .D(\Data_Mem/n6512 ), .CLK(clk), .RST(
        rst), .I(e_init[1279]), .Q(o[1279]) );
  DFF \Data_Mem/memory_reg[38][0]  ( .D(\Data_Mem/n6513 ), .CLK(clk), .RST(rst), .I(e_init[1216]), .Q(o[1216]) );
  DFF \Data_Mem/memory_reg[38][1]  ( .D(\Data_Mem/n6514 ), .CLK(clk), .RST(rst), .I(e_init[1217]), .Q(o[1217]) );
  DFF \Data_Mem/memory_reg[38][2]  ( .D(\Data_Mem/n6515 ), .CLK(clk), .RST(rst), .I(e_init[1218]), .Q(o[1218]) );
  DFF \Data_Mem/memory_reg[38][3]  ( .D(\Data_Mem/n6516 ), .CLK(clk), .RST(rst), .I(e_init[1219]), .Q(o[1219]) );
  DFF \Data_Mem/memory_reg[38][4]  ( .D(\Data_Mem/n6517 ), .CLK(clk), .RST(rst), .I(e_init[1220]), .Q(o[1220]) );
  DFF \Data_Mem/memory_reg[38][5]  ( .D(\Data_Mem/n6518 ), .CLK(clk), .RST(rst), .I(e_init[1221]), .Q(o[1221]) );
  DFF \Data_Mem/memory_reg[38][6]  ( .D(\Data_Mem/n6519 ), .CLK(clk), .RST(rst), .I(e_init[1222]), .Q(o[1222]) );
  DFF \Data_Mem/memory_reg[38][7]  ( .D(\Data_Mem/n6520 ), .CLK(clk), .RST(rst), .I(e_init[1223]), .Q(o[1223]) );
  DFF \Data_Mem/memory_reg[38][8]  ( .D(\Data_Mem/n6521 ), .CLK(clk), .RST(rst), .I(e_init[1224]), .Q(o[1224]) );
  DFF \Data_Mem/memory_reg[38][9]  ( .D(\Data_Mem/n6522 ), .CLK(clk), .RST(rst), .I(e_init[1225]), .Q(o[1225]) );
  DFF \Data_Mem/memory_reg[38][10]  ( .D(\Data_Mem/n6523 ), .CLK(clk), .RST(
        rst), .I(e_init[1226]), .Q(o[1226]) );
  DFF \Data_Mem/memory_reg[38][11]  ( .D(\Data_Mem/n6524 ), .CLK(clk), .RST(
        rst), .I(e_init[1227]), .Q(o[1227]) );
  DFF \Data_Mem/memory_reg[38][12]  ( .D(\Data_Mem/n6525 ), .CLK(clk), .RST(
        rst), .I(e_init[1228]), .Q(o[1228]) );
  DFF \Data_Mem/memory_reg[38][13]  ( .D(\Data_Mem/n6526 ), .CLK(clk), .RST(
        rst), .I(e_init[1229]), .Q(o[1229]) );
  DFF \Data_Mem/memory_reg[38][14]  ( .D(\Data_Mem/n6527 ), .CLK(clk), .RST(
        rst), .I(e_init[1230]), .Q(o[1230]) );
  DFF \Data_Mem/memory_reg[38][15]  ( .D(\Data_Mem/n6528 ), .CLK(clk), .RST(
        rst), .I(e_init[1231]), .Q(o[1231]) );
  DFF \Data_Mem/memory_reg[38][16]  ( .D(\Data_Mem/n6529 ), .CLK(clk), .RST(
        rst), .I(e_init[1232]), .Q(o[1232]) );
  DFF \Data_Mem/memory_reg[38][17]  ( .D(\Data_Mem/n6530 ), .CLK(clk), .RST(
        rst), .I(e_init[1233]), .Q(o[1233]) );
  DFF \Data_Mem/memory_reg[38][18]  ( .D(\Data_Mem/n6531 ), .CLK(clk), .RST(
        rst), .I(e_init[1234]), .Q(o[1234]) );
  DFF \Data_Mem/memory_reg[38][19]  ( .D(\Data_Mem/n6532 ), .CLK(clk), .RST(
        rst), .I(e_init[1235]), .Q(o[1235]) );
  DFF \Data_Mem/memory_reg[38][20]  ( .D(\Data_Mem/n6533 ), .CLK(clk), .RST(
        rst), .I(e_init[1236]), .Q(o[1236]) );
  DFF \Data_Mem/memory_reg[38][21]  ( .D(\Data_Mem/n6534 ), .CLK(clk), .RST(
        rst), .I(e_init[1237]), .Q(o[1237]) );
  DFF \Data_Mem/memory_reg[38][22]  ( .D(\Data_Mem/n6535 ), .CLK(clk), .RST(
        rst), .I(e_init[1238]), .Q(o[1238]) );
  DFF \Data_Mem/memory_reg[38][23]  ( .D(\Data_Mem/n6536 ), .CLK(clk), .RST(
        rst), .I(e_init[1239]), .Q(o[1239]) );
  DFF \Data_Mem/memory_reg[38][24]  ( .D(\Data_Mem/n6537 ), .CLK(clk), .RST(
        rst), .I(e_init[1240]), .Q(o[1240]) );
  DFF \Data_Mem/memory_reg[38][25]  ( .D(\Data_Mem/n6538 ), .CLK(clk), .RST(
        rst), .I(e_init[1241]), .Q(o[1241]) );
  DFF \Data_Mem/memory_reg[38][26]  ( .D(\Data_Mem/n6539 ), .CLK(clk), .RST(
        rst), .I(e_init[1242]), .Q(o[1242]) );
  DFF \Data_Mem/memory_reg[38][27]  ( .D(\Data_Mem/n6540 ), .CLK(clk), .RST(
        rst), .I(e_init[1243]), .Q(o[1243]) );
  DFF \Data_Mem/memory_reg[38][28]  ( .D(\Data_Mem/n6541 ), .CLK(clk), .RST(
        rst), .I(e_init[1244]), .Q(o[1244]) );
  DFF \Data_Mem/memory_reg[38][29]  ( .D(\Data_Mem/n6542 ), .CLK(clk), .RST(
        rst), .I(e_init[1245]), .Q(o[1245]) );
  DFF \Data_Mem/memory_reg[38][30]  ( .D(\Data_Mem/n6543 ), .CLK(clk), .RST(
        rst), .I(e_init[1246]), .Q(o[1246]) );
  DFF \Data_Mem/memory_reg[38][31]  ( .D(\Data_Mem/n6544 ), .CLK(clk), .RST(
        rst), .I(e_init[1247]), .Q(o[1247]) );
  DFF \Data_Mem/memory_reg[37][0]  ( .D(\Data_Mem/n6545 ), .CLK(clk), .RST(rst), .I(e_init[1184]), .Q(o[1184]) );
  DFF \Data_Mem/memory_reg[37][1]  ( .D(\Data_Mem/n6546 ), .CLK(clk), .RST(rst), .I(e_init[1185]), .Q(o[1185]) );
  DFF \Data_Mem/memory_reg[37][2]  ( .D(\Data_Mem/n6547 ), .CLK(clk), .RST(rst), .I(e_init[1186]), .Q(o[1186]) );
  DFF \Data_Mem/memory_reg[37][3]  ( .D(\Data_Mem/n6548 ), .CLK(clk), .RST(rst), .I(e_init[1187]), .Q(o[1187]) );
  DFF \Data_Mem/memory_reg[37][4]  ( .D(\Data_Mem/n6549 ), .CLK(clk), .RST(rst), .I(e_init[1188]), .Q(o[1188]) );
  DFF \Data_Mem/memory_reg[37][5]  ( .D(\Data_Mem/n6550 ), .CLK(clk), .RST(rst), .I(e_init[1189]), .Q(o[1189]) );
  DFF \Data_Mem/memory_reg[37][6]  ( .D(\Data_Mem/n6551 ), .CLK(clk), .RST(rst), .I(e_init[1190]), .Q(o[1190]) );
  DFF \Data_Mem/memory_reg[37][7]  ( .D(\Data_Mem/n6552 ), .CLK(clk), .RST(rst), .I(e_init[1191]), .Q(o[1191]) );
  DFF \Data_Mem/memory_reg[37][8]  ( .D(\Data_Mem/n6553 ), .CLK(clk), .RST(rst), .I(e_init[1192]), .Q(o[1192]) );
  DFF \Data_Mem/memory_reg[37][9]  ( .D(\Data_Mem/n6554 ), .CLK(clk), .RST(rst), .I(e_init[1193]), .Q(o[1193]) );
  DFF \Data_Mem/memory_reg[37][10]  ( .D(\Data_Mem/n6555 ), .CLK(clk), .RST(
        rst), .I(e_init[1194]), .Q(o[1194]) );
  DFF \Data_Mem/memory_reg[37][11]  ( .D(\Data_Mem/n6556 ), .CLK(clk), .RST(
        rst), .I(e_init[1195]), .Q(o[1195]) );
  DFF \Data_Mem/memory_reg[37][12]  ( .D(\Data_Mem/n6557 ), .CLK(clk), .RST(
        rst), .I(e_init[1196]), .Q(o[1196]) );
  DFF \Data_Mem/memory_reg[37][13]  ( .D(\Data_Mem/n6558 ), .CLK(clk), .RST(
        rst), .I(e_init[1197]), .Q(o[1197]) );
  DFF \Data_Mem/memory_reg[37][14]  ( .D(\Data_Mem/n6559 ), .CLK(clk), .RST(
        rst), .I(e_init[1198]), .Q(o[1198]) );
  DFF \Data_Mem/memory_reg[37][15]  ( .D(\Data_Mem/n6560 ), .CLK(clk), .RST(
        rst), .I(e_init[1199]), .Q(o[1199]) );
  DFF \Data_Mem/memory_reg[37][16]  ( .D(\Data_Mem/n6561 ), .CLK(clk), .RST(
        rst), .I(e_init[1200]), .Q(o[1200]) );
  DFF \Data_Mem/memory_reg[37][17]  ( .D(\Data_Mem/n6562 ), .CLK(clk), .RST(
        rst), .I(e_init[1201]), .Q(o[1201]) );
  DFF \Data_Mem/memory_reg[37][18]  ( .D(\Data_Mem/n6563 ), .CLK(clk), .RST(
        rst), .I(e_init[1202]), .Q(o[1202]) );
  DFF \Data_Mem/memory_reg[37][19]  ( .D(\Data_Mem/n6564 ), .CLK(clk), .RST(
        rst), .I(e_init[1203]), .Q(o[1203]) );
  DFF \Data_Mem/memory_reg[37][20]  ( .D(\Data_Mem/n6565 ), .CLK(clk), .RST(
        rst), .I(e_init[1204]), .Q(o[1204]) );
  DFF \Data_Mem/memory_reg[37][21]  ( .D(\Data_Mem/n6566 ), .CLK(clk), .RST(
        rst), .I(e_init[1205]), .Q(o[1205]) );
  DFF \Data_Mem/memory_reg[37][22]  ( .D(\Data_Mem/n6567 ), .CLK(clk), .RST(
        rst), .I(e_init[1206]), .Q(o[1206]) );
  DFF \Data_Mem/memory_reg[37][23]  ( .D(\Data_Mem/n6568 ), .CLK(clk), .RST(
        rst), .I(e_init[1207]), .Q(o[1207]) );
  DFF \Data_Mem/memory_reg[37][24]  ( .D(\Data_Mem/n6569 ), .CLK(clk), .RST(
        rst), .I(e_init[1208]), .Q(o[1208]) );
  DFF \Data_Mem/memory_reg[37][25]  ( .D(\Data_Mem/n6570 ), .CLK(clk), .RST(
        rst), .I(e_init[1209]), .Q(o[1209]) );
  DFF \Data_Mem/memory_reg[37][26]  ( .D(\Data_Mem/n6571 ), .CLK(clk), .RST(
        rst), .I(e_init[1210]), .Q(o[1210]) );
  DFF \Data_Mem/memory_reg[37][27]  ( .D(\Data_Mem/n6572 ), .CLK(clk), .RST(
        rst), .I(e_init[1211]), .Q(o[1211]) );
  DFF \Data_Mem/memory_reg[37][28]  ( .D(\Data_Mem/n6573 ), .CLK(clk), .RST(
        rst), .I(e_init[1212]), .Q(o[1212]) );
  DFF \Data_Mem/memory_reg[37][29]  ( .D(\Data_Mem/n6574 ), .CLK(clk), .RST(
        rst), .I(e_init[1213]), .Q(o[1213]) );
  DFF \Data_Mem/memory_reg[37][30]  ( .D(\Data_Mem/n6575 ), .CLK(clk), .RST(
        rst), .I(e_init[1214]), .Q(o[1214]) );
  DFF \Data_Mem/memory_reg[37][31]  ( .D(\Data_Mem/n6576 ), .CLK(clk), .RST(
        rst), .I(e_init[1215]), .Q(o[1215]) );
  DFF \Data_Mem/memory_reg[36][0]  ( .D(\Data_Mem/n6577 ), .CLK(clk), .RST(rst), .I(e_init[1152]), .Q(o[1152]) );
  DFF \Data_Mem/memory_reg[36][1]  ( .D(\Data_Mem/n6578 ), .CLK(clk), .RST(rst), .I(e_init[1153]), .Q(o[1153]) );
  DFF \Data_Mem/memory_reg[36][2]  ( .D(\Data_Mem/n6579 ), .CLK(clk), .RST(rst), .I(e_init[1154]), .Q(o[1154]) );
  DFF \Data_Mem/memory_reg[36][3]  ( .D(\Data_Mem/n6580 ), .CLK(clk), .RST(rst), .I(e_init[1155]), .Q(o[1155]) );
  DFF \Data_Mem/memory_reg[36][4]  ( .D(\Data_Mem/n6581 ), .CLK(clk), .RST(rst), .I(e_init[1156]), .Q(o[1156]) );
  DFF \Data_Mem/memory_reg[36][5]  ( .D(\Data_Mem/n6582 ), .CLK(clk), .RST(rst), .I(e_init[1157]), .Q(o[1157]) );
  DFF \Data_Mem/memory_reg[36][6]  ( .D(\Data_Mem/n6583 ), .CLK(clk), .RST(rst), .I(e_init[1158]), .Q(o[1158]) );
  DFF \Data_Mem/memory_reg[36][7]  ( .D(\Data_Mem/n6584 ), .CLK(clk), .RST(rst), .I(e_init[1159]), .Q(o[1159]) );
  DFF \Data_Mem/memory_reg[36][8]  ( .D(\Data_Mem/n6585 ), .CLK(clk), .RST(rst), .I(e_init[1160]), .Q(o[1160]) );
  DFF \Data_Mem/memory_reg[36][9]  ( .D(\Data_Mem/n6586 ), .CLK(clk), .RST(rst), .I(e_init[1161]), .Q(o[1161]) );
  DFF \Data_Mem/memory_reg[36][10]  ( .D(\Data_Mem/n6587 ), .CLK(clk), .RST(
        rst), .I(e_init[1162]), .Q(o[1162]) );
  DFF \Data_Mem/memory_reg[36][11]  ( .D(\Data_Mem/n6588 ), .CLK(clk), .RST(
        rst), .I(e_init[1163]), .Q(o[1163]) );
  DFF \Data_Mem/memory_reg[36][12]  ( .D(\Data_Mem/n6589 ), .CLK(clk), .RST(
        rst), .I(e_init[1164]), .Q(o[1164]) );
  DFF \Data_Mem/memory_reg[36][13]  ( .D(\Data_Mem/n6590 ), .CLK(clk), .RST(
        rst), .I(e_init[1165]), .Q(o[1165]) );
  DFF \Data_Mem/memory_reg[36][14]  ( .D(\Data_Mem/n6591 ), .CLK(clk), .RST(
        rst), .I(e_init[1166]), .Q(o[1166]) );
  DFF \Data_Mem/memory_reg[36][15]  ( .D(\Data_Mem/n6592 ), .CLK(clk), .RST(
        rst), .I(e_init[1167]), .Q(o[1167]) );
  DFF \Data_Mem/memory_reg[36][16]  ( .D(\Data_Mem/n6593 ), .CLK(clk), .RST(
        rst), .I(e_init[1168]), .Q(o[1168]) );
  DFF \Data_Mem/memory_reg[36][17]  ( .D(\Data_Mem/n6594 ), .CLK(clk), .RST(
        rst), .I(e_init[1169]), .Q(o[1169]) );
  DFF \Data_Mem/memory_reg[36][18]  ( .D(\Data_Mem/n6595 ), .CLK(clk), .RST(
        rst), .I(e_init[1170]), .Q(o[1170]) );
  DFF \Data_Mem/memory_reg[36][19]  ( .D(\Data_Mem/n6596 ), .CLK(clk), .RST(
        rst), .I(e_init[1171]), .Q(o[1171]) );
  DFF \Data_Mem/memory_reg[36][20]  ( .D(\Data_Mem/n6597 ), .CLK(clk), .RST(
        rst), .I(e_init[1172]), .Q(o[1172]) );
  DFF \Data_Mem/memory_reg[36][21]  ( .D(\Data_Mem/n6598 ), .CLK(clk), .RST(
        rst), .I(e_init[1173]), .Q(o[1173]) );
  DFF \Data_Mem/memory_reg[36][22]  ( .D(\Data_Mem/n6599 ), .CLK(clk), .RST(
        rst), .I(e_init[1174]), .Q(o[1174]) );
  DFF \Data_Mem/memory_reg[36][23]  ( .D(\Data_Mem/n6600 ), .CLK(clk), .RST(
        rst), .I(e_init[1175]), .Q(o[1175]) );
  DFF \Data_Mem/memory_reg[36][24]  ( .D(\Data_Mem/n6601 ), .CLK(clk), .RST(
        rst), .I(e_init[1176]), .Q(o[1176]) );
  DFF \Data_Mem/memory_reg[36][25]  ( .D(\Data_Mem/n6602 ), .CLK(clk), .RST(
        rst), .I(e_init[1177]), .Q(o[1177]) );
  DFF \Data_Mem/memory_reg[36][26]  ( .D(\Data_Mem/n6603 ), .CLK(clk), .RST(
        rst), .I(e_init[1178]), .Q(o[1178]) );
  DFF \Data_Mem/memory_reg[36][27]  ( .D(\Data_Mem/n6604 ), .CLK(clk), .RST(
        rst), .I(e_init[1179]), .Q(o[1179]) );
  DFF \Data_Mem/memory_reg[36][28]  ( .D(\Data_Mem/n6605 ), .CLK(clk), .RST(
        rst), .I(e_init[1180]), .Q(o[1180]) );
  DFF \Data_Mem/memory_reg[36][29]  ( .D(\Data_Mem/n6606 ), .CLK(clk), .RST(
        rst), .I(e_init[1181]), .Q(o[1181]) );
  DFF \Data_Mem/memory_reg[36][30]  ( .D(\Data_Mem/n6607 ), .CLK(clk), .RST(
        rst), .I(e_init[1182]), .Q(o[1182]) );
  DFF \Data_Mem/memory_reg[36][31]  ( .D(\Data_Mem/n6608 ), .CLK(clk), .RST(
        rst), .I(e_init[1183]), .Q(o[1183]) );
  DFF \Data_Mem/memory_reg[35][0]  ( .D(\Data_Mem/n6609 ), .CLK(clk), .RST(rst), .I(e_init[1120]), .Q(o[1120]) );
  DFF \Data_Mem/memory_reg[35][1]  ( .D(\Data_Mem/n6610 ), .CLK(clk), .RST(rst), .I(e_init[1121]), .Q(o[1121]) );
  DFF \Data_Mem/memory_reg[35][2]  ( .D(\Data_Mem/n6611 ), .CLK(clk), .RST(rst), .I(e_init[1122]), .Q(o[1122]) );
  DFF \Data_Mem/memory_reg[35][3]  ( .D(\Data_Mem/n6612 ), .CLK(clk), .RST(rst), .I(e_init[1123]), .Q(o[1123]) );
  DFF \Data_Mem/memory_reg[35][4]  ( .D(\Data_Mem/n6613 ), .CLK(clk), .RST(rst), .I(e_init[1124]), .Q(o[1124]) );
  DFF \Data_Mem/memory_reg[35][5]  ( .D(\Data_Mem/n6614 ), .CLK(clk), .RST(rst), .I(e_init[1125]), .Q(o[1125]) );
  DFF \Data_Mem/memory_reg[35][6]  ( .D(\Data_Mem/n6615 ), .CLK(clk), .RST(rst), .I(e_init[1126]), .Q(o[1126]) );
  DFF \Data_Mem/memory_reg[35][7]  ( .D(\Data_Mem/n6616 ), .CLK(clk), .RST(rst), .I(e_init[1127]), .Q(o[1127]) );
  DFF \Data_Mem/memory_reg[35][8]  ( .D(\Data_Mem/n6617 ), .CLK(clk), .RST(rst), .I(e_init[1128]), .Q(o[1128]) );
  DFF \Data_Mem/memory_reg[35][9]  ( .D(\Data_Mem/n6618 ), .CLK(clk), .RST(rst), .I(e_init[1129]), .Q(o[1129]) );
  DFF \Data_Mem/memory_reg[35][10]  ( .D(\Data_Mem/n6619 ), .CLK(clk), .RST(
        rst), .I(e_init[1130]), .Q(o[1130]) );
  DFF \Data_Mem/memory_reg[35][11]  ( .D(\Data_Mem/n6620 ), .CLK(clk), .RST(
        rst), .I(e_init[1131]), .Q(o[1131]) );
  DFF \Data_Mem/memory_reg[35][12]  ( .D(\Data_Mem/n6621 ), .CLK(clk), .RST(
        rst), .I(e_init[1132]), .Q(o[1132]) );
  DFF \Data_Mem/memory_reg[35][13]  ( .D(\Data_Mem/n6622 ), .CLK(clk), .RST(
        rst), .I(e_init[1133]), .Q(o[1133]) );
  DFF \Data_Mem/memory_reg[35][14]  ( .D(\Data_Mem/n6623 ), .CLK(clk), .RST(
        rst), .I(e_init[1134]), .Q(o[1134]) );
  DFF \Data_Mem/memory_reg[35][15]  ( .D(\Data_Mem/n6624 ), .CLK(clk), .RST(
        rst), .I(e_init[1135]), .Q(o[1135]) );
  DFF \Data_Mem/memory_reg[35][16]  ( .D(\Data_Mem/n6625 ), .CLK(clk), .RST(
        rst), .I(e_init[1136]), .Q(o[1136]) );
  DFF \Data_Mem/memory_reg[35][17]  ( .D(\Data_Mem/n6626 ), .CLK(clk), .RST(
        rst), .I(e_init[1137]), .Q(o[1137]) );
  DFF \Data_Mem/memory_reg[35][18]  ( .D(\Data_Mem/n6627 ), .CLK(clk), .RST(
        rst), .I(e_init[1138]), .Q(o[1138]) );
  DFF \Data_Mem/memory_reg[35][19]  ( .D(\Data_Mem/n6628 ), .CLK(clk), .RST(
        rst), .I(e_init[1139]), .Q(o[1139]) );
  DFF \Data_Mem/memory_reg[35][20]  ( .D(\Data_Mem/n6629 ), .CLK(clk), .RST(
        rst), .I(e_init[1140]), .Q(o[1140]) );
  DFF \Data_Mem/memory_reg[35][21]  ( .D(\Data_Mem/n6630 ), .CLK(clk), .RST(
        rst), .I(e_init[1141]), .Q(o[1141]) );
  DFF \Data_Mem/memory_reg[35][22]  ( .D(\Data_Mem/n6631 ), .CLK(clk), .RST(
        rst), .I(e_init[1142]), .Q(o[1142]) );
  DFF \Data_Mem/memory_reg[35][23]  ( .D(\Data_Mem/n6632 ), .CLK(clk), .RST(
        rst), .I(e_init[1143]), .Q(o[1143]) );
  DFF \Data_Mem/memory_reg[35][24]  ( .D(\Data_Mem/n6633 ), .CLK(clk), .RST(
        rst), .I(e_init[1144]), .Q(o[1144]) );
  DFF \Data_Mem/memory_reg[35][25]  ( .D(\Data_Mem/n6634 ), .CLK(clk), .RST(
        rst), .I(e_init[1145]), .Q(o[1145]) );
  DFF \Data_Mem/memory_reg[35][26]  ( .D(\Data_Mem/n6635 ), .CLK(clk), .RST(
        rst), .I(e_init[1146]), .Q(o[1146]) );
  DFF \Data_Mem/memory_reg[35][27]  ( .D(\Data_Mem/n6636 ), .CLK(clk), .RST(
        rst), .I(e_init[1147]), .Q(o[1147]) );
  DFF \Data_Mem/memory_reg[35][28]  ( .D(\Data_Mem/n6637 ), .CLK(clk), .RST(
        rst), .I(e_init[1148]), .Q(o[1148]) );
  DFF \Data_Mem/memory_reg[35][29]  ( .D(\Data_Mem/n6638 ), .CLK(clk), .RST(
        rst), .I(e_init[1149]), .Q(o[1149]) );
  DFF \Data_Mem/memory_reg[35][30]  ( .D(\Data_Mem/n6639 ), .CLK(clk), .RST(
        rst), .I(e_init[1150]), .Q(o[1150]) );
  DFF \Data_Mem/memory_reg[35][31]  ( .D(\Data_Mem/n6640 ), .CLK(clk), .RST(
        rst), .I(e_init[1151]), .Q(o[1151]) );
  DFF \Data_Mem/memory_reg[34][0]  ( .D(\Data_Mem/n6641 ), .CLK(clk), .RST(rst), .I(e_init[1088]), .Q(o[1088]) );
  DFF \Data_Mem/memory_reg[34][1]  ( .D(\Data_Mem/n6642 ), .CLK(clk), .RST(rst), .I(e_init[1089]), .Q(o[1089]) );
  DFF \Data_Mem/memory_reg[34][2]  ( .D(\Data_Mem/n6643 ), .CLK(clk), .RST(rst), .I(e_init[1090]), .Q(o[1090]) );
  DFF \Data_Mem/memory_reg[34][3]  ( .D(\Data_Mem/n6644 ), .CLK(clk), .RST(rst), .I(e_init[1091]), .Q(o[1091]) );
  DFF \Data_Mem/memory_reg[34][4]  ( .D(\Data_Mem/n6645 ), .CLK(clk), .RST(rst), .I(e_init[1092]), .Q(o[1092]) );
  DFF \Data_Mem/memory_reg[34][5]  ( .D(\Data_Mem/n6646 ), .CLK(clk), .RST(rst), .I(e_init[1093]), .Q(o[1093]) );
  DFF \Data_Mem/memory_reg[34][6]  ( .D(\Data_Mem/n6647 ), .CLK(clk), .RST(rst), .I(e_init[1094]), .Q(o[1094]) );
  DFF \Data_Mem/memory_reg[34][7]  ( .D(\Data_Mem/n6648 ), .CLK(clk), .RST(rst), .I(e_init[1095]), .Q(o[1095]) );
  DFF \Data_Mem/memory_reg[34][8]  ( .D(\Data_Mem/n6649 ), .CLK(clk), .RST(rst), .I(e_init[1096]), .Q(o[1096]) );
  DFF \Data_Mem/memory_reg[34][9]  ( .D(\Data_Mem/n6650 ), .CLK(clk), .RST(rst), .I(e_init[1097]), .Q(o[1097]) );
  DFF \Data_Mem/memory_reg[34][10]  ( .D(\Data_Mem/n6651 ), .CLK(clk), .RST(
        rst), .I(e_init[1098]), .Q(o[1098]) );
  DFF \Data_Mem/memory_reg[34][11]  ( .D(\Data_Mem/n6652 ), .CLK(clk), .RST(
        rst), .I(e_init[1099]), .Q(o[1099]) );
  DFF \Data_Mem/memory_reg[34][12]  ( .D(\Data_Mem/n6653 ), .CLK(clk), .RST(
        rst), .I(e_init[1100]), .Q(o[1100]) );
  DFF \Data_Mem/memory_reg[34][13]  ( .D(\Data_Mem/n6654 ), .CLK(clk), .RST(
        rst), .I(e_init[1101]), .Q(o[1101]) );
  DFF \Data_Mem/memory_reg[34][14]  ( .D(\Data_Mem/n6655 ), .CLK(clk), .RST(
        rst), .I(e_init[1102]), .Q(o[1102]) );
  DFF \Data_Mem/memory_reg[34][15]  ( .D(\Data_Mem/n6656 ), .CLK(clk), .RST(
        rst), .I(e_init[1103]), .Q(o[1103]) );
  DFF \Data_Mem/memory_reg[34][16]  ( .D(\Data_Mem/n6657 ), .CLK(clk), .RST(
        rst), .I(e_init[1104]), .Q(o[1104]) );
  DFF \Data_Mem/memory_reg[34][17]  ( .D(\Data_Mem/n6658 ), .CLK(clk), .RST(
        rst), .I(e_init[1105]), .Q(o[1105]) );
  DFF \Data_Mem/memory_reg[34][18]  ( .D(\Data_Mem/n6659 ), .CLK(clk), .RST(
        rst), .I(e_init[1106]), .Q(o[1106]) );
  DFF \Data_Mem/memory_reg[34][19]  ( .D(\Data_Mem/n6660 ), .CLK(clk), .RST(
        rst), .I(e_init[1107]), .Q(o[1107]) );
  DFF \Data_Mem/memory_reg[34][20]  ( .D(\Data_Mem/n6661 ), .CLK(clk), .RST(
        rst), .I(e_init[1108]), .Q(o[1108]) );
  DFF \Data_Mem/memory_reg[34][21]  ( .D(\Data_Mem/n6662 ), .CLK(clk), .RST(
        rst), .I(e_init[1109]), .Q(o[1109]) );
  DFF \Data_Mem/memory_reg[34][22]  ( .D(\Data_Mem/n6663 ), .CLK(clk), .RST(
        rst), .I(e_init[1110]), .Q(o[1110]) );
  DFF \Data_Mem/memory_reg[34][23]  ( .D(\Data_Mem/n6664 ), .CLK(clk), .RST(
        rst), .I(e_init[1111]), .Q(o[1111]) );
  DFF \Data_Mem/memory_reg[34][24]  ( .D(\Data_Mem/n6665 ), .CLK(clk), .RST(
        rst), .I(e_init[1112]), .Q(o[1112]) );
  DFF \Data_Mem/memory_reg[34][25]  ( .D(\Data_Mem/n6666 ), .CLK(clk), .RST(
        rst), .I(e_init[1113]), .Q(o[1113]) );
  DFF \Data_Mem/memory_reg[34][26]  ( .D(\Data_Mem/n6667 ), .CLK(clk), .RST(
        rst), .I(e_init[1114]), .Q(o[1114]) );
  DFF \Data_Mem/memory_reg[34][27]  ( .D(\Data_Mem/n6668 ), .CLK(clk), .RST(
        rst), .I(e_init[1115]), .Q(o[1115]) );
  DFF \Data_Mem/memory_reg[34][28]  ( .D(\Data_Mem/n6669 ), .CLK(clk), .RST(
        rst), .I(e_init[1116]), .Q(o[1116]) );
  DFF \Data_Mem/memory_reg[34][29]  ( .D(\Data_Mem/n6670 ), .CLK(clk), .RST(
        rst), .I(e_init[1117]), .Q(o[1117]) );
  DFF \Data_Mem/memory_reg[34][30]  ( .D(\Data_Mem/n6671 ), .CLK(clk), .RST(
        rst), .I(e_init[1118]), .Q(o[1118]) );
  DFF \Data_Mem/memory_reg[34][31]  ( .D(\Data_Mem/n6672 ), .CLK(clk), .RST(
        rst), .I(e_init[1119]), .Q(o[1119]) );
  DFF \Data_Mem/memory_reg[33][0]  ( .D(\Data_Mem/n6673 ), .CLK(clk), .RST(rst), .I(e_init[1056]), .Q(o[1056]) );
  DFF \Data_Mem/memory_reg[33][1]  ( .D(\Data_Mem/n6674 ), .CLK(clk), .RST(rst), .I(e_init[1057]), .Q(o[1057]) );
  DFF \Data_Mem/memory_reg[33][2]  ( .D(\Data_Mem/n6675 ), .CLK(clk), .RST(rst), .I(e_init[1058]), .Q(o[1058]) );
  DFF \Data_Mem/memory_reg[33][3]  ( .D(\Data_Mem/n6676 ), .CLK(clk), .RST(rst), .I(e_init[1059]), .Q(o[1059]) );
  DFF \Data_Mem/memory_reg[33][4]  ( .D(\Data_Mem/n6677 ), .CLK(clk), .RST(rst), .I(e_init[1060]), .Q(o[1060]) );
  DFF \Data_Mem/memory_reg[33][5]  ( .D(\Data_Mem/n6678 ), .CLK(clk), .RST(rst), .I(e_init[1061]), .Q(o[1061]) );
  DFF \Data_Mem/memory_reg[33][6]  ( .D(\Data_Mem/n6679 ), .CLK(clk), .RST(rst), .I(e_init[1062]), .Q(o[1062]) );
  DFF \Data_Mem/memory_reg[33][7]  ( .D(\Data_Mem/n6680 ), .CLK(clk), .RST(rst), .I(e_init[1063]), .Q(o[1063]) );
  DFF \Data_Mem/memory_reg[33][8]  ( .D(\Data_Mem/n6681 ), .CLK(clk), .RST(rst), .I(e_init[1064]), .Q(o[1064]) );
  DFF \Data_Mem/memory_reg[33][9]  ( .D(\Data_Mem/n6682 ), .CLK(clk), .RST(rst), .I(e_init[1065]), .Q(o[1065]) );
  DFF \Data_Mem/memory_reg[33][10]  ( .D(\Data_Mem/n6683 ), .CLK(clk), .RST(
        rst), .I(e_init[1066]), .Q(o[1066]) );
  DFF \Data_Mem/memory_reg[33][11]  ( .D(\Data_Mem/n6684 ), .CLK(clk), .RST(
        rst), .I(e_init[1067]), .Q(o[1067]) );
  DFF \Data_Mem/memory_reg[33][12]  ( .D(\Data_Mem/n6685 ), .CLK(clk), .RST(
        rst), .I(e_init[1068]), .Q(o[1068]) );
  DFF \Data_Mem/memory_reg[33][13]  ( .D(\Data_Mem/n6686 ), .CLK(clk), .RST(
        rst), .I(e_init[1069]), .Q(o[1069]) );
  DFF \Data_Mem/memory_reg[33][14]  ( .D(\Data_Mem/n6687 ), .CLK(clk), .RST(
        rst), .I(e_init[1070]), .Q(o[1070]) );
  DFF \Data_Mem/memory_reg[33][15]  ( .D(\Data_Mem/n6688 ), .CLK(clk), .RST(
        rst), .I(e_init[1071]), .Q(o[1071]) );
  DFF \Data_Mem/memory_reg[33][16]  ( .D(\Data_Mem/n6689 ), .CLK(clk), .RST(
        rst), .I(e_init[1072]), .Q(o[1072]) );
  DFF \Data_Mem/memory_reg[33][17]  ( .D(\Data_Mem/n6690 ), .CLK(clk), .RST(
        rst), .I(e_init[1073]), .Q(o[1073]) );
  DFF \Data_Mem/memory_reg[33][18]  ( .D(\Data_Mem/n6691 ), .CLK(clk), .RST(
        rst), .I(e_init[1074]), .Q(o[1074]) );
  DFF \Data_Mem/memory_reg[33][19]  ( .D(\Data_Mem/n6692 ), .CLK(clk), .RST(
        rst), .I(e_init[1075]), .Q(o[1075]) );
  DFF \Data_Mem/memory_reg[33][20]  ( .D(\Data_Mem/n6693 ), .CLK(clk), .RST(
        rst), .I(e_init[1076]), .Q(o[1076]) );
  DFF \Data_Mem/memory_reg[33][21]  ( .D(\Data_Mem/n6694 ), .CLK(clk), .RST(
        rst), .I(e_init[1077]), .Q(o[1077]) );
  DFF \Data_Mem/memory_reg[33][22]  ( .D(\Data_Mem/n6695 ), .CLK(clk), .RST(
        rst), .I(e_init[1078]), .Q(o[1078]) );
  DFF \Data_Mem/memory_reg[33][23]  ( .D(\Data_Mem/n6696 ), .CLK(clk), .RST(
        rst), .I(e_init[1079]), .Q(o[1079]) );
  DFF \Data_Mem/memory_reg[33][24]  ( .D(\Data_Mem/n6697 ), .CLK(clk), .RST(
        rst), .I(e_init[1080]), .Q(o[1080]) );
  DFF \Data_Mem/memory_reg[33][25]  ( .D(\Data_Mem/n6698 ), .CLK(clk), .RST(
        rst), .I(e_init[1081]), .Q(o[1081]) );
  DFF \Data_Mem/memory_reg[33][26]  ( .D(\Data_Mem/n6699 ), .CLK(clk), .RST(
        rst), .I(e_init[1082]), .Q(o[1082]) );
  DFF \Data_Mem/memory_reg[33][27]  ( .D(\Data_Mem/n6700 ), .CLK(clk), .RST(
        rst), .I(e_init[1083]), .Q(o[1083]) );
  DFF \Data_Mem/memory_reg[33][28]  ( .D(\Data_Mem/n6701 ), .CLK(clk), .RST(
        rst), .I(e_init[1084]), .Q(o[1084]) );
  DFF \Data_Mem/memory_reg[33][29]  ( .D(\Data_Mem/n6702 ), .CLK(clk), .RST(
        rst), .I(e_init[1085]), .Q(o[1085]) );
  DFF \Data_Mem/memory_reg[33][30]  ( .D(\Data_Mem/n6703 ), .CLK(clk), .RST(
        rst), .I(e_init[1086]), .Q(o[1086]) );
  DFF \Data_Mem/memory_reg[33][31]  ( .D(\Data_Mem/n6704 ), .CLK(clk), .RST(
        rst), .I(e_init[1087]), .Q(o[1087]) );
  DFF \Data_Mem/memory_reg[32][0]  ( .D(\Data_Mem/n6705 ), .CLK(clk), .RST(rst), .I(e_init[1024]), .Q(o[1024]) );
  DFF \Data_Mem/memory_reg[32][1]  ( .D(\Data_Mem/n6706 ), .CLK(clk), .RST(rst), .I(e_init[1025]), .Q(o[1025]) );
  DFF \Data_Mem/memory_reg[32][2]  ( .D(\Data_Mem/n6707 ), .CLK(clk), .RST(rst), .I(e_init[1026]), .Q(o[1026]) );
  DFF \Data_Mem/memory_reg[32][3]  ( .D(\Data_Mem/n6708 ), .CLK(clk), .RST(rst), .I(e_init[1027]), .Q(o[1027]) );
  DFF \Data_Mem/memory_reg[32][4]  ( .D(\Data_Mem/n6709 ), .CLK(clk), .RST(rst), .I(e_init[1028]), .Q(o[1028]) );
  DFF \Data_Mem/memory_reg[32][5]  ( .D(\Data_Mem/n6710 ), .CLK(clk), .RST(rst), .I(e_init[1029]), .Q(o[1029]) );
  DFF \Data_Mem/memory_reg[32][6]  ( .D(\Data_Mem/n6711 ), .CLK(clk), .RST(rst), .I(e_init[1030]), .Q(o[1030]) );
  DFF \Data_Mem/memory_reg[32][7]  ( .D(\Data_Mem/n6712 ), .CLK(clk), .RST(rst), .I(e_init[1031]), .Q(o[1031]) );
  DFF \Data_Mem/memory_reg[32][8]  ( .D(\Data_Mem/n6713 ), .CLK(clk), .RST(rst), .I(e_init[1032]), .Q(o[1032]) );
  DFF \Data_Mem/memory_reg[32][9]  ( .D(\Data_Mem/n6714 ), .CLK(clk), .RST(rst), .I(e_init[1033]), .Q(o[1033]) );
  DFF \Data_Mem/memory_reg[32][10]  ( .D(\Data_Mem/n6715 ), .CLK(clk), .RST(
        rst), .I(e_init[1034]), .Q(o[1034]) );
  DFF \Data_Mem/memory_reg[32][11]  ( .D(\Data_Mem/n6716 ), .CLK(clk), .RST(
        rst), .I(e_init[1035]), .Q(o[1035]) );
  DFF \Data_Mem/memory_reg[32][12]  ( .D(\Data_Mem/n6717 ), .CLK(clk), .RST(
        rst), .I(e_init[1036]), .Q(o[1036]) );
  DFF \Data_Mem/memory_reg[32][13]  ( .D(\Data_Mem/n6718 ), .CLK(clk), .RST(
        rst), .I(e_init[1037]), .Q(o[1037]) );
  DFF \Data_Mem/memory_reg[32][14]  ( .D(\Data_Mem/n6719 ), .CLK(clk), .RST(
        rst), .I(e_init[1038]), .Q(o[1038]) );
  DFF \Data_Mem/memory_reg[32][15]  ( .D(\Data_Mem/n6720 ), .CLK(clk), .RST(
        rst), .I(e_init[1039]), .Q(o[1039]) );
  DFF \Data_Mem/memory_reg[32][16]  ( .D(\Data_Mem/n6721 ), .CLK(clk), .RST(
        rst), .I(e_init[1040]), .Q(o[1040]) );
  DFF \Data_Mem/memory_reg[32][17]  ( .D(\Data_Mem/n6722 ), .CLK(clk), .RST(
        rst), .I(e_init[1041]), .Q(o[1041]) );
  DFF \Data_Mem/memory_reg[32][18]  ( .D(\Data_Mem/n6723 ), .CLK(clk), .RST(
        rst), .I(e_init[1042]), .Q(o[1042]) );
  DFF \Data_Mem/memory_reg[32][19]  ( .D(\Data_Mem/n6724 ), .CLK(clk), .RST(
        rst), .I(e_init[1043]), .Q(o[1043]) );
  DFF \Data_Mem/memory_reg[32][20]  ( .D(\Data_Mem/n6725 ), .CLK(clk), .RST(
        rst), .I(e_init[1044]), .Q(o[1044]) );
  DFF \Data_Mem/memory_reg[32][21]  ( .D(\Data_Mem/n6726 ), .CLK(clk), .RST(
        rst), .I(e_init[1045]), .Q(o[1045]) );
  DFF \Data_Mem/memory_reg[32][22]  ( .D(\Data_Mem/n6727 ), .CLK(clk), .RST(
        rst), .I(e_init[1046]), .Q(o[1046]) );
  DFF \Data_Mem/memory_reg[32][23]  ( .D(\Data_Mem/n6728 ), .CLK(clk), .RST(
        rst), .I(e_init[1047]), .Q(o[1047]) );
  DFF \Data_Mem/memory_reg[32][24]  ( .D(\Data_Mem/n6729 ), .CLK(clk), .RST(
        rst), .I(e_init[1048]), .Q(o[1048]) );
  DFF \Data_Mem/memory_reg[32][25]  ( .D(\Data_Mem/n6730 ), .CLK(clk), .RST(
        rst), .I(e_init[1049]), .Q(o[1049]) );
  DFF \Data_Mem/memory_reg[32][26]  ( .D(\Data_Mem/n6731 ), .CLK(clk), .RST(
        rst), .I(e_init[1050]), .Q(o[1050]) );
  DFF \Data_Mem/memory_reg[32][27]  ( .D(\Data_Mem/n6732 ), .CLK(clk), .RST(
        rst), .I(e_init[1051]), .Q(o[1051]) );
  DFF \Data_Mem/memory_reg[32][28]  ( .D(\Data_Mem/n6733 ), .CLK(clk), .RST(
        rst), .I(e_init[1052]), .Q(o[1052]) );
  DFF \Data_Mem/memory_reg[32][29]  ( .D(\Data_Mem/n6734 ), .CLK(clk), .RST(
        rst), .I(e_init[1053]), .Q(o[1053]) );
  DFF \Data_Mem/memory_reg[32][30]  ( .D(\Data_Mem/n6735 ), .CLK(clk), .RST(
        rst), .I(e_init[1054]), .Q(o[1054]) );
  DFF \Data_Mem/memory_reg[32][31]  ( .D(\Data_Mem/n6736 ), .CLK(clk), .RST(
        rst), .I(e_init[1055]), .Q(o[1055]) );
  DFF \Data_Mem/memory_reg[31][0]  ( .D(\Data_Mem/n6737 ), .CLK(clk), .RST(rst), .I(e_init[992]), .Q(o[992]) );
  DFF \Data_Mem/memory_reg[31][1]  ( .D(\Data_Mem/n6738 ), .CLK(clk), .RST(rst), .I(e_init[993]), .Q(o[993]) );
  DFF \Data_Mem/memory_reg[31][2]  ( .D(\Data_Mem/n6739 ), .CLK(clk), .RST(rst), .I(e_init[994]), .Q(o[994]) );
  DFF \Data_Mem/memory_reg[31][3]  ( .D(\Data_Mem/n6740 ), .CLK(clk), .RST(rst), .I(e_init[995]), .Q(o[995]) );
  DFF \Data_Mem/memory_reg[31][4]  ( .D(\Data_Mem/n6741 ), .CLK(clk), .RST(rst), .I(e_init[996]), .Q(o[996]) );
  DFF \Data_Mem/memory_reg[31][5]  ( .D(\Data_Mem/n6742 ), .CLK(clk), .RST(rst), .I(e_init[997]), .Q(o[997]) );
  DFF \Data_Mem/memory_reg[31][6]  ( .D(\Data_Mem/n6743 ), .CLK(clk), .RST(rst), .I(e_init[998]), .Q(o[998]) );
  DFF \Data_Mem/memory_reg[31][7]  ( .D(\Data_Mem/n6744 ), .CLK(clk), .RST(rst), .I(e_init[999]), .Q(o[999]) );
  DFF \Data_Mem/memory_reg[31][8]  ( .D(\Data_Mem/n6745 ), .CLK(clk), .RST(rst), .I(e_init[1000]), .Q(o[1000]) );
  DFF \Data_Mem/memory_reg[31][9]  ( .D(\Data_Mem/n6746 ), .CLK(clk), .RST(rst), .I(e_init[1001]), .Q(o[1001]) );
  DFF \Data_Mem/memory_reg[31][10]  ( .D(\Data_Mem/n6747 ), .CLK(clk), .RST(
        rst), .I(e_init[1002]), .Q(o[1002]) );
  DFF \Data_Mem/memory_reg[31][11]  ( .D(\Data_Mem/n6748 ), .CLK(clk), .RST(
        rst), .I(e_init[1003]), .Q(o[1003]) );
  DFF \Data_Mem/memory_reg[31][12]  ( .D(\Data_Mem/n6749 ), .CLK(clk), .RST(
        rst), .I(e_init[1004]), .Q(o[1004]) );
  DFF \Data_Mem/memory_reg[31][13]  ( .D(\Data_Mem/n6750 ), .CLK(clk), .RST(
        rst), .I(e_init[1005]), .Q(o[1005]) );
  DFF \Data_Mem/memory_reg[31][14]  ( .D(\Data_Mem/n6751 ), .CLK(clk), .RST(
        rst), .I(e_init[1006]), .Q(o[1006]) );
  DFF \Data_Mem/memory_reg[31][15]  ( .D(\Data_Mem/n6752 ), .CLK(clk), .RST(
        rst), .I(e_init[1007]), .Q(o[1007]) );
  DFF \Data_Mem/memory_reg[31][16]  ( .D(\Data_Mem/n6753 ), .CLK(clk), .RST(
        rst), .I(e_init[1008]), .Q(o[1008]) );
  DFF \Data_Mem/memory_reg[31][17]  ( .D(\Data_Mem/n6754 ), .CLK(clk), .RST(
        rst), .I(e_init[1009]), .Q(o[1009]) );
  DFF \Data_Mem/memory_reg[31][18]  ( .D(\Data_Mem/n6755 ), .CLK(clk), .RST(
        rst), .I(e_init[1010]), .Q(o[1010]) );
  DFF \Data_Mem/memory_reg[31][19]  ( .D(\Data_Mem/n6756 ), .CLK(clk), .RST(
        rst), .I(e_init[1011]), .Q(o[1011]) );
  DFF \Data_Mem/memory_reg[31][20]  ( .D(\Data_Mem/n6757 ), .CLK(clk), .RST(
        rst), .I(e_init[1012]), .Q(o[1012]) );
  DFF \Data_Mem/memory_reg[31][21]  ( .D(\Data_Mem/n6758 ), .CLK(clk), .RST(
        rst), .I(e_init[1013]), .Q(o[1013]) );
  DFF \Data_Mem/memory_reg[31][22]  ( .D(\Data_Mem/n6759 ), .CLK(clk), .RST(
        rst), .I(e_init[1014]), .Q(o[1014]) );
  DFF \Data_Mem/memory_reg[31][23]  ( .D(\Data_Mem/n6760 ), .CLK(clk), .RST(
        rst), .I(e_init[1015]), .Q(o[1015]) );
  DFF \Data_Mem/memory_reg[31][24]  ( .D(\Data_Mem/n6761 ), .CLK(clk), .RST(
        rst), .I(e_init[1016]), .Q(o[1016]) );
  DFF \Data_Mem/memory_reg[31][25]  ( .D(\Data_Mem/n6762 ), .CLK(clk), .RST(
        rst), .I(e_init[1017]), .Q(o[1017]) );
  DFF \Data_Mem/memory_reg[31][26]  ( .D(\Data_Mem/n6763 ), .CLK(clk), .RST(
        rst), .I(e_init[1018]), .Q(o[1018]) );
  DFF \Data_Mem/memory_reg[31][27]  ( .D(\Data_Mem/n6764 ), .CLK(clk), .RST(
        rst), .I(e_init[1019]), .Q(o[1019]) );
  DFF \Data_Mem/memory_reg[31][28]  ( .D(\Data_Mem/n6765 ), .CLK(clk), .RST(
        rst), .I(e_init[1020]), .Q(o[1020]) );
  DFF \Data_Mem/memory_reg[31][29]  ( .D(\Data_Mem/n6766 ), .CLK(clk), .RST(
        rst), .I(e_init[1021]), .Q(o[1021]) );
  DFF \Data_Mem/memory_reg[31][30]  ( .D(\Data_Mem/n6767 ), .CLK(clk), .RST(
        rst), .I(e_init[1022]), .Q(o[1022]) );
  DFF \Data_Mem/memory_reg[31][31]  ( .D(\Data_Mem/n6768 ), .CLK(clk), .RST(
        rst), .I(e_init[1023]), .Q(o[1023]) );
  DFF \Data_Mem/memory_reg[30][0]  ( .D(\Data_Mem/n6769 ), .CLK(clk), .RST(rst), .I(e_init[960]), .Q(o[960]) );
  DFF \Data_Mem/memory_reg[30][1]  ( .D(\Data_Mem/n6770 ), .CLK(clk), .RST(rst), .I(e_init[961]), .Q(o[961]) );
  DFF \Data_Mem/memory_reg[30][2]  ( .D(\Data_Mem/n6771 ), .CLK(clk), .RST(rst), .I(e_init[962]), .Q(o[962]) );
  DFF \Data_Mem/memory_reg[30][3]  ( .D(\Data_Mem/n6772 ), .CLK(clk), .RST(rst), .I(e_init[963]), .Q(o[963]) );
  DFF \Data_Mem/memory_reg[30][4]  ( .D(\Data_Mem/n6773 ), .CLK(clk), .RST(rst), .I(e_init[964]), .Q(o[964]) );
  DFF \Data_Mem/memory_reg[30][5]  ( .D(\Data_Mem/n6774 ), .CLK(clk), .RST(rst), .I(e_init[965]), .Q(o[965]) );
  DFF \Data_Mem/memory_reg[30][6]  ( .D(\Data_Mem/n6775 ), .CLK(clk), .RST(rst), .I(e_init[966]), .Q(o[966]) );
  DFF \Data_Mem/memory_reg[30][7]  ( .D(\Data_Mem/n6776 ), .CLK(clk), .RST(rst), .I(e_init[967]), .Q(o[967]) );
  DFF \Data_Mem/memory_reg[30][8]  ( .D(\Data_Mem/n6777 ), .CLK(clk), .RST(rst), .I(e_init[968]), .Q(o[968]) );
  DFF \Data_Mem/memory_reg[30][9]  ( .D(\Data_Mem/n6778 ), .CLK(clk), .RST(rst), .I(e_init[969]), .Q(o[969]) );
  DFF \Data_Mem/memory_reg[30][10]  ( .D(\Data_Mem/n6779 ), .CLK(clk), .RST(
        rst), .I(e_init[970]), .Q(o[970]) );
  DFF \Data_Mem/memory_reg[30][11]  ( .D(\Data_Mem/n6780 ), .CLK(clk), .RST(
        rst), .I(e_init[971]), .Q(o[971]) );
  DFF \Data_Mem/memory_reg[30][12]  ( .D(\Data_Mem/n6781 ), .CLK(clk), .RST(
        rst), .I(e_init[972]), .Q(o[972]) );
  DFF \Data_Mem/memory_reg[30][13]  ( .D(\Data_Mem/n6782 ), .CLK(clk), .RST(
        rst), .I(e_init[973]), .Q(o[973]) );
  DFF \Data_Mem/memory_reg[30][14]  ( .D(\Data_Mem/n6783 ), .CLK(clk), .RST(
        rst), .I(e_init[974]), .Q(o[974]) );
  DFF \Data_Mem/memory_reg[30][15]  ( .D(\Data_Mem/n6784 ), .CLK(clk), .RST(
        rst), .I(e_init[975]), .Q(o[975]) );
  DFF \Data_Mem/memory_reg[30][16]  ( .D(\Data_Mem/n6785 ), .CLK(clk), .RST(
        rst), .I(e_init[976]), .Q(o[976]) );
  DFF \Data_Mem/memory_reg[30][17]  ( .D(\Data_Mem/n6786 ), .CLK(clk), .RST(
        rst), .I(e_init[977]), .Q(o[977]) );
  DFF \Data_Mem/memory_reg[30][18]  ( .D(\Data_Mem/n6787 ), .CLK(clk), .RST(
        rst), .I(e_init[978]), .Q(o[978]) );
  DFF \Data_Mem/memory_reg[30][19]  ( .D(\Data_Mem/n6788 ), .CLK(clk), .RST(
        rst), .I(e_init[979]), .Q(o[979]) );
  DFF \Data_Mem/memory_reg[30][20]  ( .D(\Data_Mem/n6789 ), .CLK(clk), .RST(
        rst), .I(e_init[980]), .Q(o[980]) );
  DFF \Data_Mem/memory_reg[30][21]  ( .D(\Data_Mem/n6790 ), .CLK(clk), .RST(
        rst), .I(e_init[981]), .Q(o[981]) );
  DFF \Data_Mem/memory_reg[30][22]  ( .D(\Data_Mem/n6791 ), .CLK(clk), .RST(
        rst), .I(e_init[982]), .Q(o[982]) );
  DFF \Data_Mem/memory_reg[30][23]  ( .D(\Data_Mem/n6792 ), .CLK(clk), .RST(
        rst), .I(e_init[983]), .Q(o[983]) );
  DFF \Data_Mem/memory_reg[30][24]  ( .D(\Data_Mem/n6793 ), .CLK(clk), .RST(
        rst), .I(e_init[984]), .Q(o[984]) );
  DFF \Data_Mem/memory_reg[30][25]  ( .D(\Data_Mem/n6794 ), .CLK(clk), .RST(
        rst), .I(e_init[985]), .Q(o[985]) );
  DFF \Data_Mem/memory_reg[30][26]  ( .D(\Data_Mem/n6795 ), .CLK(clk), .RST(
        rst), .I(e_init[986]), .Q(o[986]) );
  DFF \Data_Mem/memory_reg[30][27]  ( .D(\Data_Mem/n6796 ), .CLK(clk), .RST(
        rst), .I(e_init[987]), .Q(o[987]) );
  DFF \Data_Mem/memory_reg[30][28]  ( .D(\Data_Mem/n6797 ), .CLK(clk), .RST(
        rst), .I(e_init[988]), .Q(o[988]) );
  DFF \Data_Mem/memory_reg[30][29]  ( .D(\Data_Mem/n6798 ), .CLK(clk), .RST(
        rst), .I(e_init[989]), .Q(o[989]) );
  DFF \Data_Mem/memory_reg[30][30]  ( .D(\Data_Mem/n6799 ), .CLK(clk), .RST(
        rst), .I(e_init[990]), .Q(o[990]) );
  DFF \Data_Mem/memory_reg[30][31]  ( .D(\Data_Mem/n6800 ), .CLK(clk), .RST(
        rst), .I(e_init[991]), .Q(o[991]) );
  DFF \Data_Mem/memory_reg[29][0]  ( .D(\Data_Mem/n6801 ), .CLK(clk), .RST(rst), .I(e_init[928]), .Q(o[928]) );
  DFF \Data_Mem/memory_reg[29][1]  ( .D(\Data_Mem/n6802 ), .CLK(clk), .RST(rst), .I(e_init[929]), .Q(o[929]) );
  DFF \Data_Mem/memory_reg[29][2]  ( .D(\Data_Mem/n6803 ), .CLK(clk), .RST(rst), .I(e_init[930]), .Q(o[930]) );
  DFF \Data_Mem/memory_reg[29][3]  ( .D(\Data_Mem/n6804 ), .CLK(clk), .RST(rst), .I(e_init[931]), .Q(o[931]) );
  DFF \Data_Mem/memory_reg[29][4]  ( .D(\Data_Mem/n6805 ), .CLK(clk), .RST(rst), .I(e_init[932]), .Q(o[932]) );
  DFF \Data_Mem/memory_reg[29][5]  ( .D(\Data_Mem/n6806 ), .CLK(clk), .RST(rst), .I(e_init[933]), .Q(o[933]) );
  DFF \Data_Mem/memory_reg[29][6]  ( .D(\Data_Mem/n6807 ), .CLK(clk), .RST(rst), .I(e_init[934]), .Q(o[934]) );
  DFF \Data_Mem/memory_reg[29][7]  ( .D(\Data_Mem/n6808 ), .CLK(clk), .RST(rst), .I(e_init[935]), .Q(o[935]) );
  DFF \Data_Mem/memory_reg[29][8]  ( .D(\Data_Mem/n6809 ), .CLK(clk), .RST(rst), .I(e_init[936]), .Q(o[936]) );
  DFF \Data_Mem/memory_reg[29][9]  ( .D(\Data_Mem/n6810 ), .CLK(clk), .RST(rst), .I(e_init[937]), .Q(o[937]) );
  DFF \Data_Mem/memory_reg[29][10]  ( .D(\Data_Mem/n6811 ), .CLK(clk), .RST(
        rst), .I(e_init[938]), .Q(o[938]) );
  DFF \Data_Mem/memory_reg[29][11]  ( .D(\Data_Mem/n6812 ), .CLK(clk), .RST(
        rst), .I(e_init[939]), .Q(o[939]) );
  DFF \Data_Mem/memory_reg[29][12]  ( .D(\Data_Mem/n6813 ), .CLK(clk), .RST(
        rst), .I(e_init[940]), .Q(o[940]) );
  DFF \Data_Mem/memory_reg[29][13]  ( .D(\Data_Mem/n6814 ), .CLK(clk), .RST(
        rst), .I(e_init[941]), .Q(o[941]) );
  DFF \Data_Mem/memory_reg[29][14]  ( .D(\Data_Mem/n6815 ), .CLK(clk), .RST(
        rst), .I(e_init[942]), .Q(o[942]) );
  DFF \Data_Mem/memory_reg[29][15]  ( .D(\Data_Mem/n6816 ), .CLK(clk), .RST(
        rst), .I(e_init[943]), .Q(o[943]) );
  DFF \Data_Mem/memory_reg[29][16]  ( .D(\Data_Mem/n6817 ), .CLK(clk), .RST(
        rst), .I(e_init[944]), .Q(o[944]) );
  DFF \Data_Mem/memory_reg[29][17]  ( .D(\Data_Mem/n6818 ), .CLK(clk), .RST(
        rst), .I(e_init[945]), .Q(o[945]) );
  DFF \Data_Mem/memory_reg[29][18]  ( .D(\Data_Mem/n6819 ), .CLK(clk), .RST(
        rst), .I(e_init[946]), .Q(o[946]) );
  DFF \Data_Mem/memory_reg[29][19]  ( .D(\Data_Mem/n6820 ), .CLK(clk), .RST(
        rst), .I(e_init[947]), .Q(o[947]) );
  DFF \Data_Mem/memory_reg[29][20]  ( .D(\Data_Mem/n6821 ), .CLK(clk), .RST(
        rst), .I(e_init[948]), .Q(o[948]) );
  DFF \Data_Mem/memory_reg[29][21]  ( .D(\Data_Mem/n6822 ), .CLK(clk), .RST(
        rst), .I(e_init[949]), .Q(o[949]) );
  DFF \Data_Mem/memory_reg[29][22]  ( .D(\Data_Mem/n6823 ), .CLK(clk), .RST(
        rst), .I(e_init[950]), .Q(o[950]) );
  DFF \Data_Mem/memory_reg[29][23]  ( .D(\Data_Mem/n6824 ), .CLK(clk), .RST(
        rst), .I(e_init[951]), .Q(o[951]) );
  DFF \Data_Mem/memory_reg[29][24]  ( .D(\Data_Mem/n6825 ), .CLK(clk), .RST(
        rst), .I(e_init[952]), .Q(o[952]) );
  DFF \Data_Mem/memory_reg[29][25]  ( .D(\Data_Mem/n6826 ), .CLK(clk), .RST(
        rst), .I(e_init[953]), .Q(o[953]) );
  DFF \Data_Mem/memory_reg[29][26]  ( .D(\Data_Mem/n6827 ), .CLK(clk), .RST(
        rst), .I(e_init[954]), .Q(o[954]) );
  DFF \Data_Mem/memory_reg[29][27]  ( .D(\Data_Mem/n6828 ), .CLK(clk), .RST(
        rst), .I(e_init[955]), .Q(o[955]) );
  DFF \Data_Mem/memory_reg[29][28]  ( .D(\Data_Mem/n6829 ), .CLK(clk), .RST(
        rst), .I(e_init[956]), .Q(o[956]) );
  DFF \Data_Mem/memory_reg[29][29]  ( .D(\Data_Mem/n6830 ), .CLK(clk), .RST(
        rst), .I(e_init[957]), .Q(o[957]) );
  DFF \Data_Mem/memory_reg[29][30]  ( .D(\Data_Mem/n6831 ), .CLK(clk), .RST(
        rst), .I(e_init[958]), .Q(o[958]) );
  DFF \Data_Mem/memory_reg[29][31]  ( .D(\Data_Mem/n6832 ), .CLK(clk), .RST(
        rst), .I(e_init[959]), .Q(o[959]) );
  DFF \Data_Mem/memory_reg[28][0]  ( .D(\Data_Mem/n6833 ), .CLK(clk), .RST(rst), .I(e_init[896]), .Q(o[896]) );
  DFF \Data_Mem/memory_reg[28][1]  ( .D(\Data_Mem/n6834 ), .CLK(clk), .RST(rst), .I(e_init[897]), .Q(o[897]) );
  DFF \Data_Mem/memory_reg[28][2]  ( .D(\Data_Mem/n6835 ), .CLK(clk), .RST(rst), .I(e_init[898]), .Q(o[898]) );
  DFF \Data_Mem/memory_reg[28][3]  ( .D(\Data_Mem/n6836 ), .CLK(clk), .RST(rst), .I(e_init[899]), .Q(o[899]) );
  DFF \Data_Mem/memory_reg[28][4]  ( .D(\Data_Mem/n6837 ), .CLK(clk), .RST(rst), .I(e_init[900]), .Q(o[900]) );
  DFF \Data_Mem/memory_reg[28][5]  ( .D(\Data_Mem/n6838 ), .CLK(clk), .RST(rst), .I(e_init[901]), .Q(o[901]) );
  DFF \Data_Mem/memory_reg[28][6]  ( .D(\Data_Mem/n6839 ), .CLK(clk), .RST(rst), .I(e_init[902]), .Q(o[902]) );
  DFF \Data_Mem/memory_reg[28][7]  ( .D(\Data_Mem/n6840 ), .CLK(clk), .RST(rst), .I(e_init[903]), .Q(o[903]) );
  DFF \Data_Mem/memory_reg[28][8]  ( .D(\Data_Mem/n6841 ), .CLK(clk), .RST(rst), .I(e_init[904]), .Q(o[904]) );
  DFF \Data_Mem/memory_reg[28][9]  ( .D(\Data_Mem/n6842 ), .CLK(clk), .RST(rst), .I(e_init[905]), .Q(o[905]) );
  DFF \Data_Mem/memory_reg[28][10]  ( .D(\Data_Mem/n6843 ), .CLK(clk), .RST(
        rst), .I(e_init[906]), .Q(o[906]) );
  DFF \Data_Mem/memory_reg[28][11]  ( .D(\Data_Mem/n6844 ), .CLK(clk), .RST(
        rst), .I(e_init[907]), .Q(o[907]) );
  DFF \Data_Mem/memory_reg[28][12]  ( .D(\Data_Mem/n6845 ), .CLK(clk), .RST(
        rst), .I(e_init[908]), .Q(o[908]) );
  DFF \Data_Mem/memory_reg[28][13]  ( .D(\Data_Mem/n6846 ), .CLK(clk), .RST(
        rst), .I(e_init[909]), .Q(o[909]) );
  DFF \Data_Mem/memory_reg[28][14]  ( .D(\Data_Mem/n6847 ), .CLK(clk), .RST(
        rst), .I(e_init[910]), .Q(o[910]) );
  DFF \Data_Mem/memory_reg[28][15]  ( .D(\Data_Mem/n6848 ), .CLK(clk), .RST(
        rst), .I(e_init[911]), .Q(o[911]) );
  DFF \Data_Mem/memory_reg[28][16]  ( .D(\Data_Mem/n6849 ), .CLK(clk), .RST(
        rst), .I(e_init[912]), .Q(o[912]) );
  DFF \Data_Mem/memory_reg[28][17]  ( .D(\Data_Mem/n6850 ), .CLK(clk), .RST(
        rst), .I(e_init[913]), .Q(o[913]) );
  DFF \Data_Mem/memory_reg[28][18]  ( .D(\Data_Mem/n6851 ), .CLK(clk), .RST(
        rst), .I(e_init[914]), .Q(o[914]) );
  DFF \Data_Mem/memory_reg[28][19]  ( .D(\Data_Mem/n6852 ), .CLK(clk), .RST(
        rst), .I(e_init[915]), .Q(o[915]) );
  DFF \Data_Mem/memory_reg[28][20]  ( .D(\Data_Mem/n6853 ), .CLK(clk), .RST(
        rst), .I(e_init[916]), .Q(o[916]) );
  DFF \Data_Mem/memory_reg[28][21]  ( .D(\Data_Mem/n6854 ), .CLK(clk), .RST(
        rst), .I(e_init[917]), .Q(o[917]) );
  DFF \Data_Mem/memory_reg[28][22]  ( .D(\Data_Mem/n6855 ), .CLK(clk), .RST(
        rst), .I(e_init[918]), .Q(o[918]) );
  DFF \Data_Mem/memory_reg[28][23]  ( .D(\Data_Mem/n6856 ), .CLK(clk), .RST(
        rst), .I(e_init[919]), .Q(o[919]) );
  DFF \Data_Mem/memory_reg[28][24]  ( .D(\Data_Mem/n6857 ), .CLK(clk), .RST(
        rst), .I(e_init[920]), .Q(o[920]) );
  DFF \Data_Mem/memory_reg[28][25]  ( .D(\Data_Mem/n6858 ), .CLK(clk), .RST(
        rst), .I(e_init[921]), .Q(o[921]) );
  DFF \Data_Mem/memory_reg[28][26]  ( .D(\Data_Mem/n6859 ), .CLK(clk), .RST(
        rst), .I(e_init[922]), .Q(o[922]) );
  DFF \Data_Mem/memory_reg[28][27]  ( .D(\Data_Mem/n6860 ), .CLK(clk), .RST(
        rst), .I(e_init[923]), .Q(o[923]) );
  DFF \Data_Mem/memory_reg[28][28]  ( .D(\Data_Mem/n6861 ), .CLK(clk), .RST(
        rst), .I(e_init[924]), .Q(o[924]) );
  DFF \Data_Mem/memory_reg[28][29]  ( .D(\Data_Mem/n6862 ), .CLK(clk), .RST(
        rst), .I(e_init[925]), .Q(o[925]) );
  DFF \Data_Mem/memory_reg[28][30]  ( .D(\Data_Mem/n6863 ), .CLK(clk), .RST(
        rst), .I(e_init[926]), .Q(o[926]) );
  DFF \Data_Mem/memory_reg[28][31]  ( .D(\Data_Mem/n6864 ), .CLK(clk), .RST(
        rst), .I(e_init[927]), .Q(o[927]) );
  DFF \Data_Mem/memory_reg[27][0]  ( .D(\Data_Mem/n6865 ), .CLK(clk), .RST(rst), .I(e_init[864]), .Q(o[864]) );
  DFF \Data_Mem/memory_reg[27][1]  ( .D(\Data_Mem/n6866 ), .CLK(clk), .RST(rst), .I(e_init[865]), .Q(o[865]) );
  DFF \Data_Mem/memory_reg[27][2]  ( .D(\Data_Mem/n6867 ), .CLK(clk), .RST(rst), .I(e_init[866]), .Q(o[866]) );
  DFF \Data_Mem/memory_reg[27][3]  ( .D(\Data_Mem/n6868 ), .CLK(clk), .RST(rst), .I(e_init[867]), .Q(o[867]) );
  DFF \Data_Mem/memory_reg[27][4]  ( .D(\Data_Mem/n6869 ), .CLK(clk), .RST(rst), .I(e_init[868]), .Q(o[868]) );
  DFF \Data_Mem/memory_reg[27][5]  ( .D(\Data_Mem/n6870 ), .CLK(clk), .RST(rst), .I(e_init[869]), .Q(o[869]) );
  DFF \Data_Mem/memory_reg[27][6]  ( .D(\Data_Mem/n6871 ), .CLK(clk), .RST(rst), .I(e_init[870]), .Q(o[870]) );
  DFF \Data_Mem/memory_reg[27][7]  ( .D(\Data_Mem/n6872 ), .CLK(clk), .RST(rst), .I(e_init[871]), .Q(o[871]) );
  DFF \Data_Mem/memory_reg[27][8]  ( .D(\Data_Mem/n6873 ), .CLK(clk), .RST(rst), .I(e_init[872]), .Q(o[872]) );
  DFF \Data_Mem/memory_reg[27][9]  ( .D(\Data_Mem/n6874 ), .CLK(clk), .RST(rst), .I(e_init[873]), .Q(o[873]) );
  DFF \Data_Mem/memory_reg[27][10]  ( .D(\Data_Mem/n6875 ), .CLK(clk), .RST(
        rst), .I(e_init[874]), .Q(o[874]) );
  DFF \Data_Mem/memory_reg[27][11]  ( .D(\Data_Mem/n6876 ), .CLK(clk), .RST(
        rst), .I(e_init[875]), .Q(o[875]) );
  DFF \Data_Mem/memory_reg[27][12]  ( .D(\Data_Mem/n6877 ), .CLK(clk), .RST(
        rst), .I(e_init[876]), .Q(o[876]) );
  DFF \Data_Mem/memory_reg[27][13]  ( .D(\Data_Mem/n6878 ), .CLK(clk), .RST(
        rst), .I(e_init[877]), .Q(o[877]) );
  DFF \Data_Mem/memory_reg[27][14]  ( .D(\Data_Mem/n6879 ), .CLK(clk), .RST(
        rst), .I(e_init[878]), .Q(o[878]) );
  DFF \Data_Mem/memory_reg[27][15]  ( .D(\Data_Mem/n6880 ), .CLK(clk), .RST(
        rst), .I(e_init[879]), .Q(o[879]) );
  DFF \Data_Mem/memory_reg[27][16]  ( .D(\Data_Mem/n6881 ), .CLK(clk), .RST(
        rst), .I(e_init[880]), .Q(o[880]) );
  DFF \Data_Mem/memory_reg[27][17]  ( .D(\Data_Mem/n6882 ), .CLK(clk), .RST(
        rst), .I(e_init[881]), .Q(o[881]) );
  DFF \Data_Mem/memory_reg[27][18]  ( .D(\Data_Mem/n6883 ), .CLK(clk), .RST(
        rst), .I(e_init[882]), .Q(o[882]) );
  DFF \Data_Mem/memory_reg[27][19]  ( .D(\Data_Mem/n6884 ), .CLK(clk), .RST(
        rst), .I(e_init[883]), .Q(o[883]) );
  DFF \Data_Mem/memory_reg[27][20]  ( .D(\Data_Mem/n6885 ), .CLK(clk), .RST(
        rst), .I(e_init[884]), .Q(o[884]) );
  DFF \Data_Mem/memory_reg[27][21]  ( .D(\Data_Mem/n6886 ), .CLK(clk), .RST(
        rst), .I(e_init[885]), .Q(o[885]) );
  DFF \Data_Mem/memory_reg[27][22]  ( .D(\Data_Mem/n6887 ), .CLK(clk), .RST(
        rst), .I(e_init[886]), .Q(o[886]) );
  DFF \Data_Mem/memory_reg[27][23]  ( .D(\Data_Mem/n6888 ), .CLK(clk), .RST(
        rst), .I(e_init[887]), .Q(o[887]) );
  DFF \Data_Mem/memory_reg[27][24]  ( .D(\Data_Mem/n6889 ), .CLK(clk), .RST(
        rst), .I(e_init[888]), .Q(o[888]) );
  DFF \Data_Mem/memory_reg[27][25]  ( .D(\Data_Mem/n6890 ), .CLK(clk), .RST(
        rst), .I(e_init[889]), .Q(o[889]) );
  DFF \Data_Mem/memory_reg[27][26]  ( .D(\Data_Mem/n6891 ), .CLK(clk), .RST(
        rst), .I(e_init[890]), .Q(o[890]) );
  DFF \Data_Mem/memory_reg[27][27]  ( .D(\Data_Mem/n6892 ), .CLK(clk), .RST(
        rst), .I(e_init[891]), .Q(o[891]) );
  DFF \Data_Mem/memory_reg[27][28]  ( .D(\Data_Mem/n6893 ), .CLK(clk), .RST(
        rst), .I(e_init[892]), .Q(o[892]) );
  DFF \Data_Mem/memory_reg[27][29]  ( .D(\Data_Mem/n6894 ), .CLK(clk), .RST(
        rst), .I(e_init[893]), .Q(o[893]) );
  DFF \Data_Mem/memory_reg[27][30]  ( .D(\Data_Mem/n6895 ), .CLK(clk), .RST(
        rst), .I(e_init[894]), .Q(o[894]) );
  DFF \Data_Mem/memory_reg[27][31]  ( .D(\Data_Mem/n6896 ), .CLK(clk), .RST(
        rst), .I(e_init[895]), .Q(o[895]) );
  DFF \Data_Mem/memory_reg[26][0]  ( .D(\Data_Mem/n6897 ), .CLK(clk), .RST(rst), .I(e_init[832]), .Q(o[832]) );
  DFF \Data_Mem/memory_reg[26][1]  ( .D(\Data_Mem/n6898 ), .CLK(clk), .RST(rst), .I(e_init[833]), .Q(o[833]) );
  DFF \Data_Mem/memory_reg[26][2]  ( .D(\Data_Mem/n6899 ), .CLK(clk), .RST(rst), .I(e_init[834]), .Q(o[834]) );
  DFF \Data_Mem/memory_reg[26][3]  ( .D(\Data_Mem/n6900 ), .CLK(clk), .RST(rst), .I(e_init[835]), .Q(o[835]) );
  DFF \Data_Mem/memory_reg[26][4]  ( .D(\Data_Mem/n6901 ), .CLK(clk), .RST(rst), .I(e_init[836]), .Q(o[836]) );
  DFF \Data_Mem/memory_reg[26][5]  ( .D(\Data_Mem/n6902 ), .CLK(clk), .RST(rst), .I(e_init[837]), .Q(o[837]) );
  DFF \Data_Mem/memory_reg[26][6]  ( .D(\Data_Mem/n6903 ), .CLK(clk), .RST(rst), .I(e_init[838]), .Q(o[838]) );
  DFF \Data_Mem/memory_reg[26][7]  ( .D(\Data_Mem/n6904 ), .CLK(clk), .RST(rst), .I(e_init[839]), .Q(o[839]) );
  DFF \Data_Mem/memory_reg[26][8]  ( .D(\Data_Mem/n6905 ), .CLK(clk), .RST(rst), .I(e_init[840]), .Q(o[840]) );
  DFF \Data_Mem/memory_reg[26][9]  ( .D(\Data_Mem/n6906 ), .CLK(clk), .RST(rst), .I(e_init[841]), .Q(o[841]) );
  DFF \Data_Mem/memory_reg[26][10]  ( .D(\Data_Mem/n6907 ), .CLK(clk), .RST(
        rst), .I(e_init[842]), .Q(o[842]) );
  DFF \Data_Mem/memory_reg[26][11]  ( .D(\Data_Mem/n6908 ), .CLK(clk), .RST(
        rst), .I(e_init[843]), .Q(o[843]) );
  DFF \Data_Mem/memory_reg[26][12]  ( .D(\Data_Mem/n6909 ), .CLK(clk), .RST(
        rst), .I(e_init[844]), .Q(o[844]) );
  DFF \Data_Mem/memory_reg[26][13]  ( .D(\Data_Mem/n6910 ), .CLK(clk), .RST(
        rst), .I(e_init[845]), .Q(o[845]) );
  DFF \Data_Mem/memory_reg[26][14]  ( .D(\Data_Mem/n6911 ), .CLK(clk), .RST(
        rst), .I(e_init[846]), .Q(o[846]) );
  DFF \Data_Mem/memory_reg[26][15]  ( .D(\Data_Mem/n6912 ), .CLK(clk), .RST(
        rst), .I(e_init[847]), .Q(o[847]) );
  DFF \Data_Mem/memory_reg[26][16]  ( .D(\Data_Mem/n6913 ), .CLK(clk), .RST(
        rst), .I(e_init[848]), .Q(o[848]) );
  DFF \Data_Mem/memory_reg[26][17]  ( .D(\Data_Mem/n6914 ), .CLK(clk), .RST(
        rst), .I(e_init[849]), .Q(o[849]) );
  DFF \Data_Mem/memory_reg[26][18]  ( .D(\Data_Mem/n6915 ), .CLK(clk), .RST(
        rst), .I(e_init[850]), .Q(o[850]) );
  DFF \Data_Mem/memory_reg[26][19]  ( .D(\Data_Mem/n6916 ), .CLK(clk), .RST(
        rst), .I(e_init[851]), .Q(o[851]) );
  DFF \Data_Mem/memory_reg[26][20]  ( .D(\Data_Mem/n6917 ), .CLK(clk), .RST(
        rst), .I(e_init[852]), .Q(o[852]) );
  DFF \Data_Mem/memory_reg[26][21]  ( .D(\Data_Mem/n6918 ), .CLK(clk), .RST(
        rst), .I(e_init[853]), .Q(o[853]) );
  DFF \Data_Mem/memory_reg[26][22]  ( .D(\Data_Mem/n6919 ), .CLK(clk), .RST(
        rst), .I(e_init[854]), .Q(o[854]) );
  DFF \Data_Mem/memory_reg[26][23]  ( .D(\Data_Mem/n6920 ), .CLK(clk), .RST(
        rst), .I(e_init[855]), .Q(o[855]) );
  DFF \Data_Mem/memory_reg[26][24]  ( .D(\Data_Mem/n6921 ), .CLK(clk), .RST(
        rst), .I(e_init[856]), .Q(o[856]) );
  DFF \Data_Mem/memory_reg[26][25]  ( .D(\Data_Mem/n6922 ), .CLK(clk), .RST(
        rst), .I(e_init[857]), .Q(o[857]) );
  DFF \Data_Mem/memory_reg[26][26]  ( .D(\Data_Mem/n6923 ), .CLK(clk), .RST(
        rst), .I(e_init[858]), .Q(o[858]) );
  DFF \Data_Mem/memory_reg[26][27]  ( .D(\Data_Mem/n6924 ), .CLK(clk), .RST(
        rst), .I(e_init[859]), .Q(o[859]) );
  DFF \Data_Mem/memory_reg[26][28]  ( .D(\Data_Mem/n6925 ), .CLK(clk), .RST(
        rst), .I(e_init[860]), .Q(o[860]) );
  DFF \Data_Mem/memory_reg[26][29]  ( .D(\Data_Mem/n6926 ), .CLK(clk), .RST(
        rst), .I(e_init[861]), .Q(o[861]) );
  DFF \Data_Mem/memory_reg[26][30]  ( .D(\Data_Mem/n6927 ), .CLK(clk), .RST(
        rst), .I(e_init[862]), .Q(o[862]) );
  DFF \Data_Mem/memory_reg[26][31]  ( .D(\Data_Mem/n6928 ), .CLK(clk), .RST(
        rst), .I(e_init[863]), .Q(o[863]) );
  DFF \Data_Mem/memory_reg[25][0]  ( .D(\Data_Mem/n6929 ), .CLK(clk), .RST(rst), .I(e_init[800]), .Q(o[800]) );
  DFF \Data_Mem/memory_reg[25][1]  ( .D(\Data_Mem/n6930 ), .CLK(clk), .RST(rst), .I(e_init[801]), .Q(o[801]) );
  DFF \Data_Mem/memory_reg[25][2]  ( .D(\Data_Mem/n6931 ), .CLK(clk), .RST(rst), .I(e_init[802]), .Q(o[802]) );
  DFF \Data_Mem/memory_reg[25][3]  ( .D(\Data_Mem/n6932 ), .CLK(clk), .RST(rst), .I(e_init[803]), .Q(o[803]) );
  DFF \Data_Mem/memory_reg[25][4]  ( .D(\Data_Mem/n6933 ), .CLK(clk), .RST(rst), .I(e_init[804]), .Q(o[804]) );
  DFF \Data_Mem/memory_reg[25][5]  ( .D(\Data_Mem/n6934 ), .CLK(clk), .RST(rst), .I(e_init[805]), .Q(o[805]) );
  DFF \Data_Mem/memory_reg[25][6]  ( .D(\Data_Mem/n6935 ), .CLK(clk), .RST(rst), .I(e_init[806]), .Q(o[806]) );
  DFF \Data_Mem/memory_reg[25][7]  ( .D(\Data_Mem/n6936 ), .CLK(clk), .RST(rst), .I(e_init[807]), .Q(o[807]) );
  DFF \Data_Mem/memory_reg[25][8]  ( .D(\Data_Mem/n6937 ), .CLK(clk), .RST(rst), .I(e_init[808]), .Q(o[808]) );
  DFF \Data_Mem/memory_reg[25][9]  ( .D(\Data_Mem/n6938 ), .CLK(clk), .RST(rst), .I(e_init[809]), .Q(o[809]) );
  DFF \Data_Mem/memory_reg[25][10]  ( .D(\Data_Mem/n6939 ), .CLK(clk), .RST(
        rst), .I(e_init[810]), .Q(o[810]) );
  DFF \Data_Mem/memory_reg[25][11]  ( .D(\Data_Mem/n6940 ), .CLK(clk), .RST(
        rst), .I(e_init[811]), .Q(o[811]) );
  DFF \Data_Mem/memory_reg[25][12]  ( .D(\Data_Mem/n6941 ), .CLK(clk), .RST(
        rst), .I(e_init[812]), .Q(o[812]) );
  DFF \Data_Mem/memory_reg[25][13]  ( .D(\Data_Mem/n6942 ), .CLK(clk), .RST(
        rst), .I(e_init[813]), .Q(o[813]) );
  DFF \Data_Mem/memory_reg[25][14]  ( .D(\Data_Mem/n6943 ), .CLK(clk), .RST(
        rst), .I(e_init[814]), .Q(o[814]) );
  DFF \Data_Mem/memory_reg[25][15]  ( .D(\Data_Mem/n6944 ), .CLK(clk), .RST(
        rst), .I(e_init[815]), .Q(o[815]) );
  DFF \Data_Mem/memory_reg[25][16]  ( .D(\Data_Mem/n6945 ), .CLK(clk), .RST(
        rst), .I(e_init[816]), .Q(o[816]) );
  DFF \Data_Mem/memory_reg[25][17]  ( .D(\Data_Mem/n6946 ), .CLK(clk), .RST(
        rst), .I(e_init[817]), .Q(o[817]) );
  DFF \Data_Mem/memory_reg[25][18]  ( .D(\Data_Mem/n6947 ), .CLK(clk), .RST(
        rst), .I(e_init[818]), .Q(o[818]) );
  DFF \Data_Mem/memory_reg[25][19]  ( .D(\Data_Mem/n6948 ), .CLK(clk), .RST(
        rst), .I(e_init[819]), .Q(o[819]) );
  DFF \Data_Mem/memory_reg[25][20]  ( .D(\Data_Mem/n6949 ), .CLK(clk), .RST(
        rst), .I(e_init[820]), .Q(o[820]) );
  DFF \Data_Mem/memory_reg[25][21]  ( .D(\Data_Mem/n6950 ), .CLK(clk), .RST(
        rst), .I(e_init[821]), .Q(o[821]) );
  DFF \Data_Mem/memory_reg[25][22]  ( .D(\Data_Mem/n6951 ), .CLK(clk), .RST(
        rst), .I(e_init[822]), .Q(o[822]) );
  DFF \Data_Mem/memory_reg[25][23]  ( .D(\Data_Mem/n6952 ), .CLK(clk), .RST(
        rst), .I(e_init[823]), .Q(o[823]) );
  DFF \Data_Mem/memory_reg[25][24]  ( .D(\Data_Mem/n6953 ), .CLK(clk), .RST(
        rst), .I(e_init[824]), .Q(o[824]) );
  DFF \Data_Mem/memory_reg[25][25]  ( .D(\Data_Mem/n6954 ), .CLK(clk), .RST(
        rst), .I(e_init[825]), .Q(o[825]) );
  DFF \Data_Mem/memory_reg[25][26]  ( .D(\Data_Mem/n6955 ), .CLK(clk), .RST(
        rst), .I(e_init[826]), .Q(o[826]) );
  DFF \Data_Mem/memory_reg[25][27]  ( .D(\Data_Mem/n6956 ), .CLK(clk), .RST(
        rst), .I(e_init[827]), .Q(o[827]) );
  DFF \Data_Mem/memory_reg[25][28]  ( .D(\Data_Mem/n6957 ), .CLK(clk), .RST(
        rst), .I(e_init[828]), .Q(o[828]) );
  DFF \Data_Mem/memory_reg[25][29]  ( .D(\Data_Mem/n6958 ), .CLK(clk), .RST(
        rst), .I(e_init[829]), .Q(o[829]) );
  DFF \Data_Mem/memory_reg[25][30]  ( .D(\Data_Mem/n6959 ), .CLK(clk), .RST(
        rst), .I(e_init[830]), .Q(o[830]) );
  DFF \Data_Mem/memory_reg[25][31]  ( .D(\Data_Mem/n6960 ), .CLK(clk), .RST(
        rst), .I(e_init[831]), .Q(o[831]) );
  DFF \Data_Mem/memory_reg[24][0]  ( .D(\Data_Mem/n6961 ), .CLK(clk), .RST(rst), .I(e_init[768]), .Q(o[768]) );
  DFF \Data_Mem/memory_reg[24][1]  ( .D(\Data_Mem/n6962 ), .CLK(clk), .RST(rst), .I(e_init[769]), .Q(o[769]) );
  DFF \Data_Mem/memory_reg[24][2]  ( .D(\Data_Mem/n6963 ), .CLK(clk), .RST(rst), .I(e_init[770]), .Q(o[770]) );
  DFF \Data_Mem/memory_reg[24][3]  ( .D(\Data_Mem/n6964 ), .CLK(clk), .RST(rst), .I(e_init[771]), .Q(o[771]) );
  DFF \Data_Mem/memory_reg[24][4]  ( .D(\Data_Mem/n6965 ), .CLK(clk), .RST(rst), .I(e_init[772]), .Q(o[772]) );
  DFF \Data_Mem/memory_reg[24][5]  ( .D(\Data_Mem/n6966 ), .CLK(clk), .RST(rst), .I(e_init[773]), .Q(o[773]) );
  DFF \Data_Mem/memory_reg[24][6]  ( .D(\Data_Mem/n6967 ), .CLK(clk), .RST(rst), .I(e_init[774]), .Q(o[774]) );
  DFF \Data_Mem/memory_reg[24][7]  ( .D(\Data_Mem/n6968 ), .CLK(clk), .RST(rst), .I(e_init[775]), .Q(o[775]) );
  DFF \Data_Mem/memory_reg[24][8]  ( .D(\Data_Mem/n6969 ), .CLK(clk), .RST(rst), .I(e_init[776]), .Q(o[776]) );
  DFF \Data_Mem/memory_reg[24][9]  ( .D(\Data_Mem/n6970 ), .CLK(clk), .RST(rst), .I(e_init[777]), .Q(o[777]) );
  DFF \Data_Mem/memory_reg[24][10]  ( .D(\Data_Mem/n6971 ), .CLK(clk), .RST(
        rst), .I(e_init[778]), .Q(o[778]) );
  DFF \Data_Mem/memory_reg[24][11]  ( .D(\Data_Mem/n6972 ), .CLK(clk), .RST(
        rst), .I(e_init[779]), .Q(o[779]) );
  DFF \Data_Mem/memory_reg[24][12]  ( .D(\Data_Mem/n6973 ), .CLK(clk), .RST(
        rst), .I(e_init[780]), .Q(o[780]) );
  DFF \Data_Mem/memory_reg[24][13]  ( .D(\Data_Mem/n6974 ), .CLK(clk), .RST(
        rst), .I(e_init[781]), .Q(o[781]) );
  DFF \Data_Mem/memory_reg[24][14]  ( .D(\Data_Mem/n6975 ), .CLK(clk), .RST(
        rst), .I(e_init[782]), .Q(o[782]) );
  DFF \Data_Mem/memory_reg[24][15]  ( .D(\Data_Mem/n6976 ), .CLK(clk), .RST(
        rst), .I(e_init[783]), .Q(o[783]) );
  DFF \Data_Mem/memory_reg[24][16]  ( .D(\Data_Mem/n6977 ), .CLK(clk), .RST(
        rst), .I(e_init[784]), .Q(o[784]) );
  DFF \Data_Mem/memory_reg[24][17]  ( .D(\Data_Mem/n6978 ), .CLK(clk), .RST(
        rst), .I(e_init[785]), .Q(o[785]) );
  DFF \Data_Mem/memory_reg[24][18]  ( .D(\Data_Mem/n6979 ), .CLK(clk), .RST(
        rst), .I(e_init[786]), .Q(o[786]) );
  DFF \Data_Mem/memory_reg[24][19]  ( .D(\Data_Mem/n6980 ), .CLK(clk), .RST(
        rst), .I(e_init[787]), .Q(o[787]) );
  DFF \Data_Mem/memory_reg[24][20]  ( .D(\Data_Mem/n6981 ), .CLK(clk), .RST(
        rst), .I(e_init[788]), .Q(o[788]) );
  DFF \Data_Mem/memory_reg[24][21]  ( .D(\Data_Mem/n6982 ), .CLK(clk), .RST(
        rst), .I(e_init[789]), .Q(o[789]) );
  DFF \Data_Mem/memory_reg[24][22]  ( .D(\Data_Mem/n6983 ), .CLK(clk), .RST(
        rst), .I(e_init[790]), .Q(o[790]) );
  DFF \Data_Mem/memory_reg[24][23]  ( .D(\Data_Mem/n6984 ), .CLK(clk), .RST(
        rst), .I(e_init[791]), .Q(o[791]) );
  DFF \Data_Mem/memory_reg[24][24]  ( .D(\Data_Mem/n6985 ), .CLK(clk), .RST(
        rst), .I(e_init[792]), .Q(o[792]) );
  DFF \Data_Mem/memory_reg[24][25]  ( .D(\Data_Mem/n6986 ), .CLK(clk), .RST(
        rst), .I(e_init[793]), .Q(o[793]) );
  DFF \Data_Mem/memory_reg[24][26]  ( .D(\Data_Mem/n6987 ), .CLK(clk), .RST(
        rst), .I(e_init[794]), .Q(o[794]) );
  DFF \Data_Mem/memory_reg[24][27]  ( .D(\Data_Mem/n6988 ), .CLK(clk), .RST(
        rst), .I(e_init[795]), .Q(o[795]) );
  DFF \Data_Mem/memory_reg[24][28]  ( .D(\Data_Mem/n6989 ), .CLK(clk), .RST(
        rst), .I(e_init[796]), .Q(o[796]) );
  DFF \Data_Mem/memory_reg[24][29]  ( .D(\Data_Mem/n6990 ), .CLK(clk), .RST(
        rst), .I(e_init[797]), .Q(o[797]) );
  DFF \Data_Mem/memory_reg[24][30]  ( .D(\Data_Mem/n6991 ), .CLK(clk), .RST(
        rst), .I(e_init[798]), .Q(o[798]) );
  DFF \Data_Mem/memory_reg[24][31]  ( .D(\Data_Mem/n6992 ), .CLK(clk), .RST(
        rst), .I(e_init[799]), .Q(o[799]) );
  DFF \Data_Mem/memory_reg[23][0]  ( .D(\Data_Mem/n6993 ), .CLK(clk), .RST(rst), .I(e_init[736]), .Q(o[736]) );
  DFF \Data_Mem/memory_reg[23][1]  ( .D(\Data_Mem/n6994 ), .CLK(clk), .RST(rst), .I(e_init[737]), .Q(o[737]) );
  DFF \Data_Mem/memory_reg[23][2]  ( .D(\Data_Mem/n6995 ), .CLK(clk), .RST(rst), .I(e_init[738]), .Q(o[738]) );
  DFF \Data_Mem/memory_reg[23][3]  ( .D(\Data_Mem/n6996 ), .CLK(clk), .RST(rst), .I(e_init[739]), .Q(o[739]) );
  DFF \Data_Mem/memory_reg[23][4]  ( .D(\Data_Mem/n6997 ), .CLK(clk), .RST(rst), .I(e_init[740]), .Q(o[740]) );
  DFF \Data_Mem/memory_reg[23][5]  ( .D(\Data_Mem/n6998 ), .CLK(clk), .RST(rst), .I(e_init[741]), .Q(o[741]) );
  DFF \Data_Mem/memory_reg[23][6]  ( .D(\Data_Mem/n6999 ), .CLK(clk), .RST(rst), .I(e_init[742]), .Q(o[742]) );
  DFF \Data_Mem/memory_reg[23][7]  ( .D(\Data_Mem/n7000 ), .CLK(clk), .RST(rst), .I(e_init[743]), .Q(o[743]) );
  DFF \Data_Mem/memory_reg[23][8]  ( .D(\Data_Mem/n7001 ), .CLK(clk), .RST(rst), .I(e_init[744]), .Q(o[744]) );
  DFF \Data_Mem/memory_reg[23][9]  ( .D(\Data_Mem/n7002 ), .CLK(clk), .RST(rst), .I(e_init[745]), .Q(o[745]) );
  DFF \Data_Mem/memory_reg[23][10]  ( .D(\Data_Mem/n7003 ), .CLK(clk), .RST(
        rst), .I(e_init[746]), .Q(o[746]) );
  DFF \Data_Mem/memory_reg[23][11]  ( .D(\Data_Mem/n7004 ), .CLK(clk), .RST(
        rst), .I(e_init[747]), .Q(o[747]) );
  DFF \Data_Mem/memory_reg[23][12]  ( .D(\Data_Mem/n7005 ), .CLK(clk), .RST(
        rst), .I(e_init[748]), .Q(o[748]) );
  DFF \Data_Mem/memory_reg[23][13]  ( .D(\Data_Mem/n7006 ), .CLK(clk), .RST(
        rst), .I(e_init[749]), .Q(o[749]) );
  DFF \Data_Mem/memory_reg[23][14]  ( .D(\Data_Mem/n7007 ), .CLK(clk), .RST(
        rst), .I(e_init[750]), .Q(o[750]) );
  DFF \Data_Mem/memory_reg[23][15]  ( .D(\Data_Mem/n7008 ), .CLK(clk), .RST(
        rst), .I(e_init[751]), .Q(o[751]) );
  DFF \Data_Mem/memory_reg[23][16]  ( .D(\Data_Mem/n7009 ), .CLK(clk), .RST(
        rst), .I(e_init[752]), .Q(o[752]) );
  DFF \Data_Mem/memory_reg[23][17]  ( .D(\Data_Mem/n7010 ), .CLK(clk), .RST(
        rst), .I(e_init[753]), .Q(o[753]) );
  DFF \Data_Mem/memory_reg[23][18]  ( .D(\Data_Mem/n7011 ), .CLK(clk), .RST(
        rst), .I(e_init[754]), .Q(o[754]) );
  DFF \Data_Mem/memory_reg[23][19]  ( .D(\Data_Mem/n7012 ), .CLK(clk), .RST(
        rst), .I(e_init[755]), .Q(o[755]) );
  DFF \Data_Mem/memory_reg[23][20]  ( .D(\Data_Mem/n7013 ), .CLK(clk), .RST(
        rst), .I(e_init[756]), .Q(o[756]) );
  DFF \Data_Mem/memory_reg[23][21]  ( .D(\Data_Mem/n7014 ), .CLK(clk), .RST(
        rst), .I(e_init[757]), .Q(o[757]) );
  DFF \Data_Mem/memory_reg[23][22]  ( .D(\Data_Mem/n7015 ), .CLK(clk), .RST(
        rst), .I(e_init[758]), .Q(o[758]) );
  DFF \Data_Mem/memory_reg[23][23]  ( .D(\Data_Mem/n7016 ), .CLK(clk), .RST(
        rst), .I(e_init[759]), .Q(o[759]) );
  DFF \Data_Mem/memory_reg[23][24]  ( .D(\Data_Mem/n7017 ), .CLK(clk), .RST(
        rst), .I(e_init[760]), .Q(o[760]) );
  DFF \Data_Mem/memory_reg[23][25]  ( .D(\Data_Mem/n7018 ), .CLK(clk), .RST(
        rst), .I(e_init[761]), .Q(o[761]) );
  DFF \Data_Mem/memory_reg[23][26]  ( .D(\Data_Mem/n7019 ), .CLK(clk), .RST(
        rst), .I(e_init[762]), .Q(o[762]) );
  DFF \Data_Mem/memory_reg[23][27]  ( .D(\Data_Mem/n7020 ), .CLK(clk), .RST(
        rst), .I(e_init[763]), .Q(o[763]) );
  DFF \Data_Mem/memory_reg[23][28]  ( .D(\Data_Mem/n7021 ), .CLK(clk), .RST(
        rst), .I(e_init[764]), .Q(o[764]) );
  DFF \Data_Mem/memory_reg[23][29]  ( .D(\Data_Mem/n7022 ), .CLK(clk), .RST(
        rst), .I(e_init[765]), .Q(o[765]) );
  DFF \Data_Mem/memory_reg[23][30]  ( .D(\Data_Mem/n7023 ), .CLK(clk), .RST(
        rst), .I(e_init[766]), .Q(o[766]) );
  DFF \Data_Mem/memory_reg[23][31]  ( .D(\Data_Mem/n7024 ), .CLK(clk), .RST(
        rst), .I(e_init[767]), .Q(o[767]) );
  DFF \Data_Mem/memory_reg[22][0]  ( .D(\Data_Mem/n7025 ), .CLK(clk), .RST(rst), .I(e_init[704]), .Q(o[704]) );
  DFF \Data_Mem/memory_reg[22][1]  ( .D(\Data_Mem/n7026 ), .CLK(clk), .RST(rst), .I(e_init[705]), .Q(o[705]) );
  DFF \Data_Mem/memory_reg[22][2]  ( .D(\Data_Mem/n7027 ), .CLK(clk), .RST(rst), .I(e_init[706]), .Q(o[706]) );
  DFF \Data_Mem/memory_reg[22][3]  ( .D(\Data_Mem/n7028 ), .CLK(clk), .RST(rst), .I(e_init[707]), .Q(o[707]) );
  DFF \Data_Mem/memory_reg[22][4]  ( .D(\Data_Mem/n7029 ), .CLK(clk), .RST(rst), .I(e_init[708]), .Q(o[708]) );
  DFF \Data_Mem/memory_reg[22][5]  ( .D(\Data_Mem/n7030 ), .CLK(clk), .RST(rst), .I(e_init[709]), .Q(o[709]) );
  DFF \Data_Mem/memory_reg[22][6]  ( .D(\Data_Mem/n7031 ), .CLK(clk), .RST(rst), .I(e_init[710]), .Q(o[710]) );
  DFF \Data_Mem/memory_reg[22][7]  ( .D(\Data_Mem/n7032 ), .CLK(clk), .RST(rst), .I(e_init[711]), .Q(o[711]) );
  DFF \Data_Mem/memory_reg[22][8]  ( .D(\Data_Mem/n7033 ), .CLK(clk), .RST(rst), .I(e_init[712]), .Q(o[712]) );
  DFF \Data_Mem/memory_reg[22][9]  ( .D(\Data_Mem/n7034 ), .CLK(clk), .RST(rst), .I(e_init[713]), .Q(o[713]) );
  DFF \Data_Mem/memory_reg[22][10]  ( .D(\Data_Mem/n7035 ), .CLK(clk), .RST(
        rst), .I(e_init[714]), .Q(o[714]) );
  DFF \Data_Mem/memory_reg[22][11]  ( .D(\Data_Mem/n7036 ), .CLK(clk), .RST(
        rst), .I(e_init[715]), .Q(o[715]) );
  DFF \Data_Mem/memory_reg[22][12]  ( .D(\Data_Mem/n7037 ), .CLK(clk), .RST(
        rst), .I(e_init[716]), .Q(o[716]) );
  DFF \Data_Mem/memory_reg[22][13]  ( .D(\Data_Mem/n7038 ), .CLK(clk), .RST(
        rst), .I(e_init[717]), .Q(o[717]) );
  DFF \Data_Mem/memory_reg[22][14]  ( .D(\Data_Mem/n7039 ), .CLK(clk), .RST(
        rst), .I(e_init[718]), .Q(o[718]) );
  DFF \Data_Mem/memory_reg[22][15]  ( .D(\Data_Mem/n7040 ), .CLK(clk), .RST(
        rst), .I(e_init[719]), .Q(o[719]) );
  DFF \Data_Mem/memory_reg[22][16]  ( .D(\Data_Mem/n7041 ), .CLK(clk), .RST(
        rst), .I(e_init[720]), .Q(o[720]) );
  DFF \Data_Mem/memory_reg[22][17]  ( .D(\Data_Mem/n7042 ), .CLK(clk), .RST(
        rst), .I(e_init[721]), .Q(o[721]) );
  DFF \Data_Mem/memory_reg[22][18]  ( .D(\Data_Mem/n7043 ), .CLK(clk), .RST(
        rst), .I(e_init[722]), .Q(o[722]) );
  DFF \Data_Mem/memory_reg[22][19]  ( .D(\Data_Mem/n7044 ), .CLK(clk), .RST(
        rst), .I(e_init[723]), .Q(o[723]) );
  DFF \Data_Mem/memory_reg[22][20]  ( .D(\Data_Mem/n7045 ), .CLK(clk), .RST(
        rst), .I(e_init[724]), .Q(o[724]) );
  DFF \Data_Mem/memory_reg[22][21]  ( .D(\Data_Mem/n7046 ), .CLK(clk), .RST(
        rst), .I(e_init[725]), .Q(o[725]) );
  DFF \Data_Mem/memory_reg[22][22]  ( .D(\Data_Mem/n7047 ), .CLK(clk), .RST(
        rst), .I(e_init[726]), .Q(o[726]) );
  DFF \Data_Mem/memory_reg[22][23]  ( .D(\Data_Mem/n7048 ), .CLK(clk), .RST(
        rst), .I(e_init[727]), .Q(o[727]) );
  DFF \Data_Mem/memory_reg[22][24]  ( .D(\Data_Mem/n7049 ), .CLK(clk), .RST(
        rst), .I(e_init[728]), .Q(o[728]) );
  DFF \Data_Mem/memory_reg[22][25]  ( .D(\Data_Mem/n7050 ), .CLK(clk), .RST(
        rst), .I(e_init[729]), .Q(o[729]) );
  DFF \Data_Mem/memory_reg[22][26]  ( .D(\Data_Mem/n7051 ), .CLK(clk), .RST(
        rst), .I(e_init[730]), .Q(o[730]) );
  DFF \Data_Mem/memory_reg[22][27]  ( .D(\Data_Mem/n7052 ), .CLK(clk), .RST(
        rst), .I(e_init[731]), .Q(o[731]) );
  DFF \Data_Mem/memory_reg[22][28]  ( .D(\Data_Mem/n7053 ), .CLK(clk), .RST(
        rst), .I(e_init[732]), .Q(o[732]) );
  DFF \Data_Mem/memory_reg[22][29]  ( .D(\Data_Mem/n7054 ), .CLK(clk), .RST(
        rst), .I(e_init[733]), .Q(o[733]) );
  DFF \Data_Mem/memory_reg[22][30]  ( .D(\Data_Mem/n7055 ), .CLK(clk), .RST(
        rst), .I(e_init[734]), .Q(o[734]) );
  DFF \Data_Mem/memory_reg[22][31]  ( .D(\Data_Mem/n7056 ), .CLK(clk), .RST(
        rst), .I(e_init[735]), .Q(o[735]) );
  DFF \Data_Mem/memory_reg[21][0]  ( .D(\Data_Mem/n7057 ), .CLK(clk), .RST(rst), .I(e_init[672]), .Q(o[672]) );
  DFF \Data_Mem/memory_reg[21][1]  ( .D(\Data_Mem/n7058 ), .CLK(clk), .RST(rst), .I(e_init[673]), .Q(o[673]) );
  DFF \Data_Mem/memory_reg[21][2]  ( .D(\Data_Mem/n7059 ), .CLK(clk), .RST(rst), .I(e_init[674]), .Q(o[674]) );
  DFF \Data_Mem/memory_reg[21][3]  ( .D(\Data_Mem/n7060 ), .CLK(clk), .RST(rst), .I(e_init[675]), .Q(o[675]) );
  DFF \Data_Mem/memory_reg[21][4]  ( .D(\Data_Mem/n7061 ), .CLK(clk), .RST(rst), .I(e_init[676]), .Q(o[676]) );
  DFF \Data_Mem/memory_reg[21][5]  ( .D(\Data_Mem/n7062 ), .CLK(clk), .RST(rst), .I(e_init[677]), .Q(o[677]) );
  DFF \Data_Mem/memory_reg[21][6]  ( .D(\Data_Mem/n7063 ), .CLK(clk), .RST(rst), .I(e_init[678]), .Q(o[678]) );
  DFF \Data_Mem/memory_reg[21][7]  ( .D(\Data_Mem/n7064 ), .CLK(clk), .RST(rst), .I(e_init[679]), .Q(o[679]) );
  DFF \Data_Mem/memory_reg[21][8]  ( .D(\Data_Mem/n7065 ), .CLK(clk), .RST(rst), .I(e_init[680]), .Q(o[680]) );
  DFF \Data_Mem/memory_reg[21][9]  ( .D(\Data_Mem/n7066 ), .CLK(clk), .RST(rst), .I(e_init[681]), .Q(o[681]) );
  DFF \Data_Mem/memory_reg[21][10]  ( .D(\Data_Mem/n7067 ), .CLK(clk), .RST(
        rst), .I(e_init[682]), .Q(o[682]) );
  DFF \Data_Mem/memory_reg[21][11]  ( .D(\Data_Mem/n7068 ), .CLK(clk), .RST(
        rst), .I(e_init[683]), .Q(o[683]) );
  DFF \Data_Mem/memory_reg[21][12]  ( .D(\Data_Mem/n7069 ), .CLK(clk), .RST(
        rst), .I(e_init[684]), .Q(o[684]) );
  DFF \Data_Mem/memory_reg[21][13]  ( .D(\Data_Mem/n7070 ), .CLK(clk), .RST(
        rst), .I(e_init[685]), .Q(o[685]) );
  DFF \Data_Mem/memory_reg[21][14]  ( .D(\Data_Mem/n7071 ), .CLK(clk), .RST(
        rst), .I(e_init[686]), .Q(o[686]) );
  DFF \Data_Mem/memory_reg[21][15]  ( .D(\Data_Mem/n7072 ), .CLK(clk), .RST(
        rst), .I(e_init[687]), .Q(o[687]) );
  DFF \Data_Mem/memory_reg[21][16]  ( .D(\Data_Mem/n7073 ), .CLK(clk), .RST(
        rst), .I(e_init[688]), .Q(o[688]) );
  DFF \Data_Mem/memory_reg[21][17]  ( .D(\Data_Mem/n7074 ), .CLK(clk), .RST(
        rst), .I(e_init[689]), .Q(o[689]) );
  DFF \Data_Mem/memory_reg[21][18]  ( .D(\Data_Mem/n7075 ), .CLK(clk), .RST(
        rst), .I(e_init[690]), .Q(o[690]) );
  DFF \Data_Mem/memory_reg[21][19]  ( .D(\Data_Mem/n7076 ), .CLK(clk), .RST(
        rst), .I(e_init[691]), .Q(o[691]) );
  DFF \Data_Mem/memory_reg[21][20]  ( .D(\Data_Mem/n7077 ), .CLK(clk), .RST(
        rst), .I(e_init[692]), .Q(o[692]) );
  DFF \Data_Mem/memory_reg[21][21]  ( .D(\Data_Mem/n7078 ), .CLK(clk), .RST(
        rst), .I(e_init[693]), .Q(o[693]) );
  DFF \Data_Mem/memory_reg[21][22]  ( .D(\Data_Mem/n7079 ), .CLK(clk), .RST(
        rst), .I(e_init[694]), .Q(o[694]) );
  DFF \Data_Mem/memory_reg[21][23]  ( .D(\Data_Mem/n7080 ), .CLK(clk), .RST(
        rst), .I(e_init[695]), .Q(o[695]) );
  DFF \Data_Mem/memory_reg[21][24]  ( .D(\Data_Mem/n7081 ), .CLK(clk), .RST(
        rst), .I(e_init[696]), .Q(o[696]) );
  DFF \Data_Mem/memory_reg[21][25]  ( .D(\Data_Mem/n7082 ), .CLK(clk), .RST(
        rst), .I(e_init[697]), .Q(o[697]) );
  DFF \Data_Mem/memory_reg[21][26]  ( .D(\Data_Mem/n7083 ), .CLK(clk), .RST(
        rst), .I(e_init[698]), .Q(o[698]) );
  DFF \Data_Mem/memory_reg[21][27]  ( .D(\Data_Mem/n7084 ), .CLK(clk), .RST(
        rst), .I(e_init[699]), .Q(o[699]) );
  DFF \Data_Mem/memory_reg[21][28]  ( .D(\Data_Mem/n7085 ), .CLK(clk), .RST(
        rst), .I(e_init[700]), .Q(o[700]) );
  DFF \Data_Mem/memory_reg[21][29]  ( .D(\Data_Mem/n7086 ), .CLK(clk), .RST(
        rst), .I(e_init[701]), .Q(o[701]) );
  DFF \Data_Mem/memory_reg[21][30]  ( .D(\Data_Mem/n7087 ), .CLK(clk), .RST(
        rst), .I(e_init[702]), .Q(o[702]) );
  DFF \Data_Mem/memory_reg[21][31]  ( .D(\Data_Mem/n7088 ), .CLK(clk), .RST(
        rst), .I(e_init[703]), .Q(o[703]) );
  DFF \Data_Mem/memory_reg[20][0]  ( .D(\Data_Mem/n7089 ), .CLK(clk), .RST(rst), .I(e_init[640]), .Q(o[640]) );
  DFF \Data_Mem/memory_reg[20][1]  ( .D(\Data_Mem/n7090 ), .CLK(clk), .RST(rst), .I(e_init[641]), .Q(o[641]) );
  DFF \Data_Mem/memory_reg[20][2]  ( .D(\Data_Mem/n7091 ), .CLK(clk), .RST(rst), .I(e_init[642]), .Q(o[642]) );
  DFF \Data_Mem/memory_reg[20][3]  ( .D(\Data_Mem/n7092 ), .CLK(clk), .RST(rst), .I(e_init[643]), .Q(o[643]) );
  DFF \Data_Mem/memory_reg[20][4]  ( .D(\Data_Mem/n7093 ), .CLK(clk), .RST(rst), .I(e_init[644]), .Q(o[644]) );
  DFF \Data_Mem/memory_reg[20][5]  ( .D(\Data_Mem/n7094 ), .CLK(clk), .RST(rst), .I(e_init[645]), .Q(o[645]) );
  DFF \Data_Mem/memory_reg[20][6]  ( .D(\Data_Mem/n7095 ), .CLK(clk), .RST(rst), .I(e_init[646]), .Q(o[646]) );
  DFF \Data_Mem/memory_reg[20][7]  ( .D(\Data_Mem/n7096 ), .CLK(clk), .RST(rst), .I(e_init[647]), .Q(o[647]) );
  DFF \Data_Mem/memory_reg[20][8]  ( .D(\Data_Mem/n7097 ), .CLK(clk), .RST(rst), .I(e_init[648]), .Q(o[648]) );
  DFF \Data_Mem/memory_reg[20][9]  ( .D(\Data_Mem/n7098 ), .CLK(clk), .RST(rst), .I(e_init[649]), .Q(o[649]) );
  DFF \Data_Mem/memory_reg[20][10]  ( .D(\Data_Mem/n7099 ), .CLK(clk), .RST(
        rst), .I(e_init[650]), .Q(o[650]) );
  DFF \Data_Mem/memory_reg[20][11]  ( .D(\Data_Mem/n7100 ), .CLK(clk), .RST(
        rst), .I(e_init[651]), .Q(o[651]) );
  DFF \Data_Mem/memory_reg[20][12]  ( .D(\Data_Mem/n7101 ), .CLK(clk), .RST(
        rst), .I(e_init[652]), .Q(o[652]) );
  DFF \Data_Mem/memory_reg[20][13]  ( .D(\Data_Mem/n7102 ), .CLK(clk), .RST(
        rst), .I(e_init[653]), .Q(o[653]) );
  DFF \Data_Mem/memory_reg[20][14]  ( .D(\Data_Mem/n7103 ), .CLK(clk), .RST(
        rst), .I(e_init[654]), .Q(o[654]) );
  DFF \Data_Mem/memory_reg[20][15]  ( .D(\Data_Mem/n7104 ), .CLK(clk), .RST(
        rst), .I(e_init[655]), .Q(o[655]) );
  DFF \Data_Mem/memory_reg[20][16]  ( .D(\Data_Mem/n7105 ), .CLK(clk), .RST(
        rst), .I(e_init[656]), .Q(o[656]) );
  DFF \Data_Mem/memory_reg[20][17]  ( .D(\Data_Mem/n7106 ), .CLK(clk), .RST(
        rst), .I(e_init[657]), .Q(o[657]) );
  DFF \Data_Mem/memory_reg[20][18]  ( .D(\Data_Mem/n7107 ), .CLK(clk), .RST(
        rst), .I(e_init[658]), .Q(o[658]) );
  DFF \Data_Mem/memory_reg[20][19]  ( .D(\Data_Mem/n7108 ), .CLK(clk), .RST(
        rst), .I(e_init[659]), .Q(o[659]) );
  DFF \Data_Mem/memory_reg[20][20]  ( .D(\Data_Mem/n7109 ), .CLK(clk), .RST(
        rst), .I(e_init[660]), .Q(o[660]) );
  DFF \Data_Mem/memory_reg[20][21]  ( .D(\Data_Mem/n7110 ), .CLK(clk), .RST(
        rst), .I(e_init[661]), .Q(o[661]) );
  DFF \Data_Mem/memory_reg[20][22]  ( .D(\Data_Mem/n7111 ), .CLK(clk), .RST(
        rst), .I(e_init[662]), .Q(o[662]) );
  DFF \Data_Mem/memory_reg[20][23]  ( .D(\Data_Mem/n7112 ), .CLK(clk), .RST(
        rst), .I(e_init[663]), .Q(o[663]) );
  DFF \Data_Mem/memory_reg[20][24]  ( .D(\Data_Mem/n7113 ), .CLK(clk), .RST(
        rst), .I(e_init[664]), .Q(o[664]) );
  DFF \Data_Mem/memory_reg[20][25]  ( .D(\Data_Mem/n7114 ), .CLK(clk), .RST(
        rst), .I(e_init[665]), .Q(o[665]) );
  DFF \Data_Mem/memory_reg[20][26]  ( .D(\Data_Mem/n7115 ), .CLK(clk), .RST(
        rst), .I(e_init[666]), .Q(o[666]) );
  DFF \Data_Mem/memory_reg[20][27]  ( .D(\Data_Mem/n7116 ), .CLK(clk), .RST(
        rst), .I(e_init[667]), .Q(o[667]) );
  DFF \Data_Mem/memory_reg[20][28]  ( .D(\Data_Mem/n7117 ), .CLK(clk), .RST(
        rst), .I(e_init[668]), .Q(o[668]) );
  DFF \Data_Mem/memory_reg[20][29]  ( .D(\Data_Mem/n7118 ), .CLK(clk), .RST(
        rst), .I(e_init[669]), .Q(o[669]) );
  DFF \Data_Mem/memory_reg[20][30]  ( .D(\Data_Mem/n7119 ), .CLK(clk), .RST(
        rst), .I(e_init[670]), .Q(o[670]) );
  DFF \Data_Mem/memory_reg[20][31]  ( .D(\Data_Mem/n7120 ), .CLK(clk), .RST(
        rst), .I(e_init[671]), .Q(o[671]) );
  DFF \Data_Mem/memory_reg[19][0]  ( .D(\Data_Mem/n7121 ), .CLK(clk), .RST(rst), .I(e_init[608]), .Q(o[608]) );
  DFF \Data_Mem/memory_reg[19][1]  ( .D(\Data_Mem/n7122 ), .CLK(clk), .RST(rst), .I(e_init[609]), .Q(o[609]) );
  DFF \Data_Mem/memory_reg[19][2]  ( .D(\Data_Mem/n7123 ), .CLK(clk), .RST(rst), .I(e_init[610]), .Q(o[610]) );
  DFF \Data_Mem/memory_reg[19][3]  ( .D(\Data_Mem/n7124 ), .CLK(clk), .RST(rst), .I(e_init[611]), .Q(o[611]) );
  DFF \Data_Mem/memory_reg[19][4]  ( .D(\Data_Mem/n7125 ), .CLK(clk), .RST(rst), .I(e_init[612]), .Q(o[612]) );
  DFF \Data_Mem/memory_reg[19][5]  ( .D(\Data_Mem/n7126 ), .CLK(clk), .RST(rst), .I(e_init[613]), .Q(o[613]) );
  DFF \Data_Mem/memory_reg[19][6]  ( .D(\Data_Mem/n7127 ), .CLK(clk), .RST(rst), .I(e_init[614]), .Q(o[614]) );
  DFF \Data_Mem/memory_reg[19][7]  ( .D(\Data_Mem/n7128 ), .CLK(clk), .RST(rst), .I(e_init[615]), .Q(o[615]) );
  DFF \Data_Mem/memory_reg[19][8]  ( .D(\Data_Mem/n7129 ), .CLK(clk), .RST(rst), .I(e_init[616]), .Q(o[616]) );
  DFF \Data_Mem/memory_reg[19][9]  ( .D(\Data_Mem/n7130 ), .CLK(clk), .RST(rst), .I(e_init[617]), .Q(o[617]) );
  DFF \Data_Mem/memory_reg[19][10]  ( .D(\Data_Mem/n7131 ), .CLK(clk), .RST(
        rst), .I(e_init[618]), .Q(o[618]) );
  DFF \Data_Mem/memory_reg[19][11]  ( .D(\Data_Mem/n7132 ), .CLK(clk), .RST(
        rst), .I(e_init[619]), .Q(o[619]) );
  DFF \Data_Mem/memory_reg[19][12]  ( .D(\Data_Mem/n7133 ), .CLK(clk), .RST(
        rst), .I(e_init[620]), .Q(o[620]) );
  DFF \Data_Mem/memory_reg[19][13]  ( .D(\Data_Mem/n7134 ), .CLK(clk), .RST(
        rst), .I(e_init[621]), .Q(o[621]) );
  DFF \Data_Mem/memory_reg[19][14]  ( .D(\Data_Mem/n7135 ), .CLK(clk), .RST(
        rst), .I(e_init[622]), .Q(o[622]) );
  DFF \Data_Mem/memory_reg[19][15]  ( .D(\Data_Mem/n7136 ), .CLK(clk), .RST(
        rst), .I(e_init[623]), .Q(o[623]) );
  DFF \Data_Mem/memory_reg[19][16]  ( .D(\Data_Mem/n7137 ), .CLK(clk), .RST(
        rst), .I(e_init[624]), .Q(o[624]) );
  DFF \Data_Mem/memory_reg[19][17]  ( .D(\Data_Mem/n7138 ), .CLK(clk), .RST(
        rst), .I(e_init[625]), .Q(o[625]) );
  DFF \Data_Mem/memory_reg[19][18]  ( .D(\Data_Mem/n7139 ), .CLK(clk), .RST(
        rst), .I(e_init[626]), .Q(o[626]) );
  DFF \Data_Mem/memory_reg[19][19]  ( .D(\Data_Mem/n7140 ), .CLK(clk), .RST(
        rst), .I(e_init[627]), .Q(o[627]) );
  DFF \Data_Mem/memory_reg[19][20]  ( .D(\Data_Mem/n7141 ), .CLK(clk), .RST(
        rst), .I(e_init[628]), .Q(o[628]) );
  DFF \Data_Mem/memory_reg[19][21]  ( .D(\Data_Mem/n7142 ), .CLK(clk), .RST(
        rst), .I(e_init[629]), .Q(o[629]) );
  DFF \Data_Mem/memory_reg[19][22]  ( .D(\Data_Mem/n7143 ), .CLK(clk), .RST(
        rst), .I(e_init[630]), .Q(o[630]) );
  DFF \Data_Mem/memory_reg[19][23]  ( .D(\Data_Mem/n7144 ), .CLK(clk), .RST(
        rst), .I(e_init[631]), .Q(o[631]) );
  DFF \Data_Mem/memory_reg[19][24]  ( .D(\Data_Mem/n7145 ), .CLK(clk), .RST(
        rst), .I(e_init[632]), .Q(o[632]) );
  DFF \Data_Mem/memory_reg[19][25]  ( .D(\Data_Mem/n7146 ), .CLK(clk), .RST(
        rst), .I(e_init[633]), .Q(o[633]) );
  DFF \Data_Mem/memory_reg[19][26]  ( .D(\Data_Mem/n7147 ), .CLK(clk), .RST(
        rst), .I(e_init[634]), .Q(o[634]) );
  DFF \Data_Mem/memory_reg[19][27]  ( .D(\Data_Mem/n7148 ), .CLK(clk), .RST(
        rst), .I(e_init[635]), .Q(o[635]) );
  DFF \Data_Mem/memory_reg[19][28]  ( .D(\Data_Mem/n7149 ), .CLK(clk), .RST(
        rst), .I(e_init[636]), .Q(o[636]) );
  DFF \Data_Mem/memory_reg[19][29]  ( .D(\Data_Mem/n7150 ), .CLK(clk), .RST(
        rst), .I(e_init[637]), .Q(o[637]) );
  DFF \Data_Mem/memory_reg[19][30]  ( .D(\Data_Mem/n7151 ), .CLK(clk), .RST(
        rst), .I(e_init[638]), .Q(o[638]) );
  DFF \Data_Mem/memory_reg[19][31]  ( .D(\Data_Mem/n7152 ), .CLK(clk), .RST(
        rst), .I(e_init[639]), .Q(o[639]) );
  DFF \Data_Mem/memory_reg[18][0]  ( .D(\Data_Mem/n7153 ), .CLK(clk), .RST(rst), .I(e_init[576]), .Q(o[576]) );
  DFF \Data_Mem/memory_reg[18][1]  ( .D(\Data_Mem/n7154 ), .CLK(clk), .RST(rst), .I(e_init[577]), .Q(o[577]) );
  DFF \Data_Mem/memory_reg[18][2]  ( .D(\Data_Mem/n7155 ), .CLK(clk), .RST(rst), .I(e_init[578]), .Q(o[578]) );
  DFF \Data_Mem/memory_reg[18][3]  ( .D(\Data_Mem/n7156 ), .CLK(clk), .RST(rst), .I(e_init[579]), .Q(o[579]) );
  DFF \Data_Mem/memory_reg[18][4]  ( .D(\Data_Mem/n7157 ), .CLK(clk), .RST(rst), .I(e_init[580]), .Q(o[580]) );
  DFF \Data_Mem/memory_reg[18][5]  ( .D(\Data_Mem/n7158 ), .CLK(clk), .RST(rst), .I(e_init[581]), .Q(o[581]) );
  DFF \Data_Mem/memory_reg[18][6]  ( .D(\Data_Mem/n7159 ), .CLK(clk), .RST(rst), .I(e_init[582]), .Q(o[582]) );
  DFF \Data_Mem/memory_reg[18][7]  ( .D(\Data_Mem/n7160 ), .CLK(clk), .RST(rst), .I(e_init[583]), .Q(o[583]) );
  DFF \Data_Mem/memory_reg[18][8]  ( .D(\Data_Mem/n7161 ), .CLK(clk), .RST(rst), .I(e_init[584]), .Q(o[584]) );
  DFF \Data_Mem/memory_reg[18][9]  ( .D(\Data_Mem/n7162 ), .CLK(clk), .RST(rst), .I(e_init[585]), .Q(o[585]) );
  DFF \Data_Mem/memory_reg[18][10]  ( .D(\Data_Mem/n7163 ), .CLK(clk), .RST(
        rst), .I(e_init[586]), .Q(o[586]) );
  DFF \Data_Mem/memory_reg[18][11]  ( .D(\Data_Mem/n7164 ), .CLK(clk), .RST(
        rst), .I(e_init[587]), .Q(o[587]) );
  DFF \Data_Mem/memory_reg[18][12]  ( .D(\Data_Mem/n7165 ), .CLK(clk), .RST(
        rst), .I(e_init[588]), .Q(o[588]) );
  DFF \Data_Mem/memory_reg[18][13]  ( .D(\Data_Mem/n7166 ), .CLK(clk), .RST(
        rst), .I(e_init[589]), .Q(o[589]) );
  DFF \Data_Mem/memory_reg[18][14]  ( .D(\Data_Mem/n7167 ), .CLK(clk), .RST(
        rst), .I(e_init[590]), .Q(o[590]) );
  DFF \Data_Mem/memory_reg[18][15]  ( .D(\Data_Mem/n7168 ), .CLK(clk), .RST(
        rst), .I(e_init[591]), .Q(o[591]) );
  DFF \Data_Mem/memory_reg[18][16]  ( .D(\Data_Mem/n7169 ), .CLK(clk), .RST(
        rst), .I(e_init[592]), .Q(o[592]) );
  DFF \Data_Mem/memory_reg[18][17]  ( .D(\Data_Mem/n7170 ), .CLK(clk), .RST(
        rst), .I(e_init[593]), .Q(o[593]) );
  DFF \Data_Mem/memory_reg[18][18]  ( .D(\Data_Mem/n7171 ), .CLK(clk), .RST(
        rst), .I(e_init[594]), .Q(o[594]) );
  DFF \Data_Mem/memory_reg[18][19]  ( .D(\Data_Mem/n7172 ), .CLK(clk), .RST(
        rst), .I(e_init[595]), .Q(o[595]) );
  DFF \Data_Mem/memory_reg[18][20]  ( .D(\Data_Mem/n7173 ), .CLK(clk), .RST(
        rst), .I(e_init[596]), .Q(o[596]) );
  DFF \Data_Mem/memory_reg[18][21]  ( .D(\Data_Mem/n7174 ), .CLK(clk), .RST(
        rst), .I(e_init[597]), .Q(o[597]) );
  DFF \Data_Mem/memory_reg[18][22]  ( .D(\Data_Mem/n7175 ), .CLK(clk), .RST(
        rst), .I(e_init[598]), .Q(o[598]) );
  DFF \Data_Mem/memory_reg[18][23]  ( .D(\Data_Mem/n7176 ), .CLK(clk), .RST(
        rst), .I(e_init[599]), .Q(o[599]) );
  DFF \Data_Mem/memory_reg[18][24]  ( .D(\Data_Mem/n7177 ), .CLK(clk), .RST(
        rst), .I(e_init[600]), .Q(o[600]) );
  DFF \Data_Mem/memory_reg[18][25]  ( .D(\Data_Mem/n7178 ), .CLK(clk), .RST(
        rst), .I(e_init[601]), .Q(o[601]) );
  DFF \Data_Mem/memory_reg[18][26]  ( .D(\Data_Mem/n7179 ), .CLK(clk), .RST(
        rst), .I(e_init[602]), .Q(o[602]) );
  DFF \Data_Mem/memory_reg[18][27]  ( .D(\Data_Mem/n7180 ), .CLK(clk), .RST(
        rst), .I(e_init[603]), .Q(o[603]) );
  DFF \Data_Mem/memory_reg[18][28]  ( .D(\Data_Mem/n7181 ), .CLK(clk), .RST(
        rst), .I(e_init[604]), .Q(o[604]) );
  DFF \Data_Mem/memory_reg[18][29]  ( .D(\Data_Mem/n7182 ), .CLK(clk), .RST(
        rst), .I(e_init[605]), .Q(o[605]) );
  DFF \Data_Mem/memory_reg[18][30]  ( .D(\Data_Mem/n7183 ), .CLK(clk), .RST(
        rst), .I(e_init[606]), .Q(o[606]) );
  DFF \Data_Mem/memory_reg[18][31]  ( .D(\Data_Mem/n7184 ), .CLK(clk), .RST(
        rst), .I(e_init[607]), .Q(o[607]) );
  DFF \Data_Mem/memory_reg[17][0]  ( .D(\Data_Mem/n7185 ), .CLK(clk), .RST(rst), .I(e_init[544]), .Q(o[544]) );
  DFF \Data_Mem/memory_reg[17][1]  ( .D(\Data_Mem/n7186 ), .CLK(clk), .RST(rst), .I(e_init[545]), .Q(o[545]) );
  DFF \Data_Mem/memory_reg[17][2]  ( .D(\Data_Mem/n7187 ), .CLK(clk), .RST(rst), .I(e_init[546]), .Q(o[546]) );
  DFF \Data_Mem/memory_reg[17][3]  ( .D(\Data_Mem/n7188 ), .CLK(clk), .RST(rst), .I(e_init[547]), .Q(o[547]) );
  DFF \Data_Mem/memory_reg[17][4]  ( .D(\Data_Mem/n7189 ), .CLK(clk), .RST(rst), .I(e_init[548]), .Q(o[548]) );
  DFF \Data_Mem/memory_reg[17][5]  ( .D(\Data_Mem/n7190 ), .CLK(clk), .RST(rst), .I(e_init[549]), .Q(o[549]) );
  DFF \Data_Mem/memory_reg[17][6]  ( .D(\Data_Mem/n7191 ), .CLK(clk), .RST(rst), .I(e_init[550]), .Q(o[550]) );
  DFF \Data_Mem/memory_reg[17][7]  ( .D(\Data_Mem/n7192 ), .CLK(clk), .RST(rst), .I(e_init[551]), .Q(o[551]) );
  DFF \Data_Mem/memory_reg[17][8]  ( .D(\Data_Mem/n7193 ), .CLK(clk), .RST(rst), .I(e_init[552]), .Q(o[552]) );
  DFF \Data_Mem/memory_reg[17][9]  ( .D(\Data_Mem/n7194 ), .CLK(clk), .RST(rst), .I(e_init[553]), .Q(o[553]) );
  DFF \Data_Mem/memory_reg[17][10]  ( .D(\Data_Mem/n7195 ), .CLK(clk), .RST(
        rst), .I(e_init[554]), .Q(o[554]) );
  DFF \Data_Mem/memory_reg[17][11]  ( .D(\Data_Mem/n7196 ), .CLK(clk), .RST(
        rst), .I(e_init[555]), .Q(o[555]) );
  DFF \Data_Mem/memory_reg[17][12]  ( .D(\Data_Mem/n7197 ), .CLK(clk), .RST(
        rst), .I(e_init[556]), .Q(o[556]) );
  DFF \Data_Mem/memory_reg[17][13]  ( .D(\Data_Mem/n7198 ), .CLK(clk), .RST(
        rst), .I(e_init[557]), .Q(o[557]) );
  DFF \Data_Mem/memory_reg[17][14]  ( .D(\Data_Mem/n7199 ), .CLK(clk), .RST(
        rst), .I(e_init[558]), .Q(o[558]) );
  DFF \Data_Mem/memory_reg[17][15]  ( .D(\Data_Mem/n7200 ), .CLK(clk), .RST(
        rst), .I(e_init[559]), .Q(o[559]) );
  DFF \Data_Mem/memory_reg[17][16]  ( .D(\Data_Mem/n7201 ), .CLK(clk), .RST(
        rst), .I(e_init[560]), .Q(o[560]) );
  DFF \Data_Mem/memory_reg[17][17]  ( .D(\Data_Mem/n7202 ), .CLK(clk), .RST(
        rst), .I(e_init[561]), .Q(o[561]) );
  DFF \Data_Mem/memory_reg[17][18]  ( .D(\Data_Mem/n7203 ), .CLK(clk), .RST(
        rst), .I(e_init[562]), .Q(o[562]) );
  DFF \Data_Mem/memory_reg[17][19]  ( .D(\Data_Mem/n7204 ), .CLK(clk), .RST(
        rst), .I(e_init[563]), .Q(o[563]) );
  DFF \Data_Mem/memory_reg[17][20]  ( .D(\Data_Mem/n7205 ), .CLK(clk), .RST(
        rst), .I(e_init[564]), .Q(o[564]) );
  DFF \Data_Mem/memory_reg[17][21]  ( .D(\Data_Mem/n7206 ), .CLK(clk), .RST(
        rst), .I(e_init[565]), .Q(o[565]) );
  DFF \Data_Mem/memory_reg[17][22]  ( .D(\Data_Mem/n7207 ), .CLK(clk), .RST(
        rst), .I(e_init[566]), .Q(o[566]) );
  DFF \Data_Mem/memory_reg[17][23]  ( .D(\Data_Mem/n7208 ), .CLK(clk), .RST(
        rst), .I(e_init[567]), .Q(o[567]) );
  DFF \Data_Mem/memory_reg[17][24]  ( .D(\Data_Mem/n7209 ), .CLK(clk), .RST(
        rst), .I(e_init[568]), .Q(o[568]) );
  DFF \Data_Mem/memory_reg[17][25]  ( .D(\Data_Mem/n7210 ), .CLK(clk), .RST(
        rst), .I(e_init[569]), .Q(o[569]) );
  DFF \Data_Mem/memory_reg[17][26]  ( .D(\Data_Mem/n7211 ), .CLK(clk), .RST(
        rst), .I(e_init[570]), .Q(o[570]) );
  DFF \Data_Mem/memory_reg[17][27]  ( .D(\Data_Mem/n7212 ), .CLK(clk), .RST(
        rst), .I(e_init[571]), .Q(o[571]) );
  DFF \Data_Mem/memory_reg[17][28]  ( .D(\Data_Mem/n7213 ), .CLK(clk), .RST(
        rst), .I(e_init[572]), .Q(o[572]) );
  DFF \Data_Mem/memory_reg[17][29]  ( .D(\Data_Mem/n7214 ), .CLK(clk), .RST(
        rst), .I(e_init[573]), .Q(o[573]) );
  DFF \Data_Mem/memory_reg[17][30]  ( .D(\Data_Mem/n7215 ), .CLK(clk), .RST(
        rst), .I(e_init[574]), .Q(o[574]) );
  DFF \Data_Mem/memory_reg[17][31]  ( .D(\Data_Mem/n7216 ), .CLK(clk), .RST(
        rst), .I(e_init[575]), .Q(o[575]) );
  DFF \Data_Mem/memory_reg[16][0]  ( .D(\Data_Mem/n7217 ), .CLK(clk), .RST(rst), .I(e_init[512]), .Q(o[512]) );
  DFF \Data_Mem/memory_reg[16][1]  ( .D(\Data_Mem/n7218 ), .CLK(clk), .RST(rst), .I(e_init[513]), .Q(o[513]) );
  DFF \Data_Mem/memory_reg[16][2]  ( .D(\Data_Mem/n7219 ), .CLK(clk), .RST(rst), .I(e_init[514]), .Q(o[514]) );
  DFF \Data_Mem/memory_reg[16][3]  ( .D(\Data_Mem/n7220 ), .CLK(clk), .RST(rst), .I(e_init[515]), .Q(o[515]) );
  DFF \Data_Mem/memory_reg[16][4]  ( .D(\Data_Mem/n7221 ), .CLK(clk), .RST(rst), .I(e_init[516]), .Q(o[516]) );
  DFF \Data_Mem/memory_reg[16][5]  ( .D(\Data_Mem/n7222 ), .CLK(clk), .RST(rst), .I(e_init[517]), .Q(o[517]) );
  DFF \Data_Mem/memory_reg[16][6]  ( .D(\Data_Mem/n7223 ), .CLK(clk), .RST(rst), .I(e_init[518]), .Q(o[518]) );
  DFF \Data_Mem/memory_reg[16][7]  ( .D(\Data_Mem/n7224 ), .CLK(clk), .RST(rst), .I(e_init[519]), .Q(o[519]) );
  DFF \Data_Mem/memory_reg[16][8]  ( .D(\Data_Mem/n7225 ), .CLK(clk), .RST(rst), .I(e_init[520]), .Q(o[520]) );
  DFF \Data_Mem/memory_reg[16][9]  ( .D(\Data_Mem/n7226 ), .CLK(clk), .RST(rst), .I(e_init[521]), .Q(o[521]) );
  DFF \Data_Mem/memory_reg[16][10]  ( .D(\Data_Mem/n7227 ), .CLK(clk), .RST(
        rst), .I(e_init[522]), .Q(o[522]) );
  DFF \Data_Mem/memory_reg[16][11]  ( .D(\Data_Mem/n7228 ), .CLK(clk), .RST(
        rst), .I(e_init[523]), .Q(o[523]) );
  DFF \Data_Mem/memory_reg[16][12]  ( .D(\Data_Mem/n7229 ), .CLK(clk), .RST(
        rst), .I(e_init[524]), .Q(o[524]) );
  DFF \Data_Mem/memory_reg[16][13]  ( .D(\Data_Mem/n7230 ), .CLK(clk), .RST(
        rst), .I(e_init[525]), .Q(o[525]) );
  DFF \Data_Mem/memory_reg[16][14]  ( .D(\Data_Mem/n7231 ), .CLK(clk), .RST(
        rst), .I(e_init[526]), .Q(o[526]) );
  DFF \Data_Mem/memory_reg[16][15]  ( .D(\Data_Mem/n7232 ), .CLK(clk), .RST(
        rst), .I(e_init[527]), .Q(o[527]) );
  DFF \Data_Mem/memory_reg[16][16]  ( .D(\Data_Mem/n7233 ), .CLK(clk), .RST(
        rst), .I(e_init[528]), .Q(o[528]) );
  DFF \Data_Mem/memory_reg[16][17]  ( .D(\Data_Mem/n7234 ), .CLK(clk), .RST(
        rst), .I(e_init[529]), .Q(o[529]) );
  DFF \Data_Mem/memory_reg[16][18]  ( .D(\Data_Mem/n7235 ), .CLK(clk), .RST(
        rst), .I(e_init[530]), .Q(o[530]) );
  DFF \Data_Mem/memory_reg[16][19]  ( .D(\Data_Mem/n7236 ), .CLK(clk), .RST(
        rst), .I(e_init[531]), .Q(o[531]) );
  DFF \Data_Mem/memory_reg[16][20]  ( .D(\Data_Mem/n7237 ), .CLK(clk), .RST(
        rst), .I(e_init[532]), .Q(o[532]) );
  DFF \Data_Mem/memory_reg[16][21]  ( .D(\Data_Mem/n7238 ), .CLK(clk), .RST(
        rst), .I(e_init[533]), .Q(o[533]) );
  DFF \Data_Mem/memory_reg[16][22]  ( .D(\Data_Mem/n7239 ), .CLK(clk), .RST(
        rst), .I(e_init[534]), .Q(o[534]) );
  DFF \Data_Mem/memory_reg[16][23]  ( .D(\Data_Mem/n7240 ), .CLK(clk), .RST(
        rst), .I(e_init[535]), .Q(o[535]) );
  DFF \Data_Mem/memory_reg[16][24]  ( .D(\Data_Mem/n7241 ), .CLK(clk), .RST(
        rst), .I(e_init[536]), .Q(o[536]) );
  DFF \Data_Mem/memory_reg[16][25]  ( .D(\Data_Mem/n7242 ), .CLK(clk), .RST(
        rst), .I(e_init[537]), .Q(o[537]) );
  DFF \Data_Mem/memory_reg[16][26]  ( .D(\Data_Mem/n7243 ), .CLK(clk), .RST(
        rst), .I(e_init[538]), .Q(o[538]) );
  DFF \Data_Mem/memory_reg[16][27]  ( .D(\Data_Mem/n7244 ), .CLK(clk), .RST(
        rst), .I(e_init[539]), .Q(o[539]) );
  DFF \Data_Mem/memory_reg[16][28]  ( .D(\Data_Mem/n7245 ), .CLK(clk), .RST(
        rst), .I(e_init[540]), .Q(o[540]) );
  DFF \Data_Mem/memory_reg[16][29]  ( .D(\Data_Mem/n7246 ), .CLK(clk), .RST(
        rst), .I(e_init[541]), .Q(o[541]) );
  DFF \Data_Mem/memory_reg[16][30]  ( .D(\Data_Mem/n7247 ), .CLK(clk), .RST(
        rst), .I(e_init[542]), .Q(o[542]) );
  DFF \Data_Mem/memory_reg[16][31]  ( .D(\Data_Mem/n7248 ), .CLK(clk), .RST(
        rst), .I(e_init[543]), .Q(o[543]) );
  DFF \Data_Mem/memory_reg[15][0]  ( .D(\Data_Mem/n7249 ), .CLK(clk), .RST(rst), .I(e_init[480]), .Q(o[480]) );
  DFF \Data_Mem/memory_reg[15][1]  ( .D(\Data_Mem/n7250 ), .CLK(clk), .RST(rst), .I(e_init[481]), .Q(o[481]) );
  DFF \Data_Mem/memory_reg[15][2]  ( .D(\Data_Mem/n7251 ), .CLK(clk), .RST(rst), .I(e_init[482]), .Q(o[482]) );
  DFF \Data_Mem/memory_reg[15][3]  ( .D(\Data_Mem/n7252 ), .CLK(clk), .RST(rst), .I(e_init[483]), .Q(o[483]) );
  DFF \Data_Mem/memory_reg[15][4]  ( .D(\Data_Mem/n7253 ), .CLK(clk), .RST(rst), .I(e_init[484]), .Q(o[484]) );
  DFF \Data_Mem/memory_reg[15][5]  ( .D(\Data_Mem/n7254 ), .CLK(clk), .RST(rst), .I(e_init[485]), .Q(o[485]) );
  DFF \Data_Mem/memory_reg[15][6]  ( .D(\Data_Mem/n7255 ), .CLK(clk), .RST(rst), .I(e_init[486]), .Q(o[486]) );
  DFF \Data_Mem/memory_reg[15][7]  ( .D(\Data_Mem/n7256 ), .CLK(clk), .RST(rst), .I(e_init[487]), .Q(o[487]) );
  DFF \Data_Mem/memory_reg[15][8]  ( .D(\Data_Mem/n7257 ), .CLK(clk), .RST(rst), .I(e_init[488]), .Q(o[488]) );
  DFF \Data_Mem/memory_reg[15][9]  ( .D(\Data_Mem/n7258 ), .CLK(clk), .RST(rst), .I(e_init[489]), .Q(o[489]) );
  DFF \Data_Mem/memory_reg[15][10]  ( .D(\Data_Mem/n7259 ), .CLK(clk), .RST(
        rst), .I(e_init[490]), .Q(o[490]) );
  DFF \Data_Mem/memory_reg[15][11]  ( .D(\Data_Mem/n7260 ), .CLK(clk), .RST(
        rst), .I(e_init[491]), .Q(o[491]) );
  DFF \Data_Mem/memory_reg[15][12]  ( .D(\Data_Mem/n7261 ), .CLK(clk), .RST(
        rst), .I(e_init[492]), .Q(o[492]) );
  DFF \Data_Mem/memory_reg[15][13]  ( .D(\Data_Mem/n7262 ), .CLK(clk), .RST(
        rst), .I(e_init[493]), .Q(o[493]) );
  DFF \Data_Mem/memory_reg[15][14]  ( .D(\Data_Mem/n7263 ), .CLK(clk), .RST(
        rst), .I(e_init[494]), .Q(o[494]) );
  DFF \Data_Mem/memory_reg[15][15]  ( .D(\Data_Mem/n7264 ), .CLK(clk), .RST(
        rst), .I(e_init[495]), .Q(o[495]) );
  DFF \Data_Mem/memory_reg[15][16]  ( .D(\Data_Mem/n7265 ), .CLK(clk), .RST(
        rst), .I(e_init[496]), .Q(o[496]) );
  DFF \Data_Mem/memory_reg[15][17]  ( .D(\Data_Mem/n7266 ), .CLK(clk), .RST(
        rst), .I(e_init[497]), .Q(o[497]) );
  DFF \Data_Mem/memory_reg[15][18]  ( .D(\Data_Mem/n7267 ), .CLK(clk), .RST(
        rst), .I(e_init[498]), .Q(o[498]) );
  DFF \Data_Mem/memory_reg[15][19]  ( .D(\Data_Mem/n7268 ), .CLK(clk), .RST(
        rst), .I(e_init[499]), .Q(o[499]) );
  DFF \Data_Mem/memory_reg[15][20]  ( .D(\Data_Mem/n7269 ), .CLK(clk), .RST(
        rst), .I(e_init[500]), .Q(o[500]) );
  DFF \Data_Mem/memory_reg[15][21]  ( .D(\Data_Mem/n7270 ), .CLK(clk), .RST(
        rst), .I(e_init[501]), .Q(o[501]) );
  DFF \Data_Mem/memory_reg[15][22]  ( .D(\Data_Mem/n7271 ), .CLK(clk), .RST(
        rst), .I(e_init[502]), .Q(o[502]) );
  DFF \Data_Mem/memory_reg[15][23]  ( .D(\Data_Mem/n7272 ), .CLK(clk), .RST(
        rst), .I(e_init[503]), .Q(o[503]) );
  DFF \Data_Mem/memory_reg[15][24]  ( .D(\Data_Mem/n7273 ), .CLK(clk), .RST(
        rst), .I(e_init[504]), .Q(o[504]) );
  DFF \Data_Mem/memory_reg[15][25]  ( .D(\Data_Mem/n7274 ), .CLK(clk), .RST(
        rst), .I(e_init[505]), .Q(o[505]) );
  DFF \Data_Mem/memory_reg[15][26]  ( .D(\Data_Mem/n7275 ), .CLK(clk), .RST(
        rst), .I(e_init[506]), .Q(o[506]) );
  DFF \Data_Mem/memory_reg[15][27]  ( .D(\Data_Mem/n7276 ), .CLK(clk), .RST(
        rst), .I(e_init[507]), .Q(o[507]) );
  DFF \Data_Mem/memory_reg[15][28]  ( .D(\Data_Mem/n7277 ), .CLK(clk), .RST(
        rst), .I(e_init[508]), .Q(o[508]) );
  DFF \Data_Mem/memory_reg[15][29]  ( .D(\Data_Mem/n7278 ), .CLK(clk), .RST(
        rst), .I(e_init[509]), .Q(o[509]) );
  DFF \Data_Mem/memory_reg[15][30]  ( .D(\Data_Mem/n7279 ), .CLK(clk), .RST(
        rst), .I(e_init[510]), .Q(o[510]) );
  DFF \Data_Mem/memory_reg[15][31]  ( .D(\Data_Mem/n7280 ), .CLK(clk), .RST(
        rst), .I(e_init[511]), .Q(o[511]) );
  DFF \Data_Mem/memory_reg[14][0]  ( .D(\Data_Mem/n7281 ), .CLK(clk), .RST(rst), .I(e_init[448]), .Q(o[448]) );
  DFF \Data_Mem/memory_reg[14][1]  ( .D(\Data_Mem/n7282 ), .CLK(clk), .RST(rst), .I(e_init[449]), .Q(o[449]) );
  DFF \Data_Mem/memory_reg[14][2]  ( .D(\Data_Mem/n7283 ), .CLK(clk), .RST(rst), .I(e_init[450]), .Q(o[450]) );
  DFF \Data_Mem/memory_reg[14][3]  ( .D(\Data_Mem/n7284 ), .CLK(clk), .RST(rst), .I(e_init[451]), .Q(o[451]) );
  DFF \Data_Mem/memory_reg[14][4]  ( .D(\Data_Mem/n7285 ), .CLK(clk), .RST(rst), .I(e_init[452]), .Q(o[452]) );
  DFF \Data_Mem/memory_reg[14][5]  ( .D(\Data_Mem/n7286 ), .CLK(clk), .RST(rst), .I(e_init[453]), .Q(o[453]) );
  DFF \Data_Mem/memory_reg[14][6]  ( .D(\Data_Mem/n7287 ), .CLK(clk), .RST(rst), .I(e_init[454]), .Q(o[454]) );
  DFF \Data_Mem/memory_reg[14][7]  ( .D(\Data_Mem/n7288 ), .CLK(clk), .RST(rst), .I(e_init[455]), .Q(o[455]) );
  DFF \Data_Mem/memory_reg[14][8]  ( .D(\Data_Mem/n7289 ), .CLK(clk), .RST(rst), .I(e_init[456]), .Q(o[456]) );
  DFF \Data_Mem/memory_reg[14][9]  ( .D(\Data_Mem/n7290 ), .CLK(clk), .RST(rst), .I(e_init[457]), .Q(o[457]) );
  DFF \Data_Mem/memory_reg[14][10]  ( .D(\Data_Mem/n7291 ), .CLK(clk), .RST(
        rst), .I(e_init[458]), .Q(o[458]) );
  DFF \Data_Mem/memory_reg[14][11]  ( .D(\Data_Mem/n7292 ), .CLK(clk), .RST(
        rst), .I(e_init[459]), .Q(o[459]) );
  DFF \Data_Mem/memory_reg[14][12]  ( .D(\Data_Mem/n7293 ), .CLK(clk), .RST(
        rst), .I(e_init[460]), .Q(o[460]) );
  DFF \Data_Mem/memory_reg[14][13]  ( .D(\Data_Mem/n7294 ), .CLK(clk), .RST(
        rst), .I(e_init[461]), .Q(o[461]) );
  DFF \Data_Mem/memory_reg[14][14]  ( .D(\Data_Mem/n7295 ), .CLK(clk), .RST(
        rst), .I(e_init[462]), .Q(o[462]) );
  DFF \Data_Mem/memory_reg[14][15]  ( .D(\Data_Mem/n7296 ), .CLK(clk), .RST(
        rst), .I(e_init[463]), .Q(o[463]) );
  DFF \Data_Mem/memory_reg[14][16]  ( .D(\Data_Mem/n7297 ), .CLK(clk), .RST(
        rst), .I(e_init[464]), .Q(o[464]) );
  DFF \Data_Mem/memory_reg[14][17]  ( .D(\Data_Mem/n7298 ), .CLK(clk), .RST(
        rst), .I(e_init[465]), .Q(o[465]) );
  DFF \Data_Mem/memory_reg[14][18]  ( .D(\Data_Mem/n7299 ), .CLK(clk), .RST(
        rst), .I(e_init[466]), .Q(o[466]) );
  DFF \Data_Mem/memory_reg[14][19]  ( .D(\Data_Mem/n7300 ), .CLK(clk), .RST(
        rst), .I(e_init[467]), .Q(o[467]) );
  DFF \Data_Mem/memory_reg[14][20]  ( .D(\Data_Mem/n7301 ), .CLK(clk), .RST(
        rst), .I(e_init[468]), .Q(o[468]) );
  DFF \Data_Mem/memory_reg[14][21]  ( .D(\Data_Mem/n7302 ), .CLK(clk), .RST(
        rst), .I(e_init[469]), .Q(o[469]) );
  DFF \Data_Mem/memory_reg[14][22]  ( .D(\Data_Mem/n7303 ), .CLK(clk), .RST(
        rst), .I(e_init[470]), .Q(o[470]) );
  DFF \Data_Mem/memory_reg[14][23]  ( .D(\Data_Mem/n7304 ), .CLK(clk), .RST(
        rst), .I(e_init[471]), .Q(o[471]) );
  DFF \Data_Mem/memory_reg[14][24]  ( .D(\Data_Mem/n7305 ), .CLK(clk), .RST(
        rst), .I(e_init[472]), .Q(o[472]) );
  DFF \Data_Mem/memory_reg[14][25]  ( .D(\Data_Mem/n7306 ), .CLK(clk), .RST(
        rst), .I(e_init[473]), .Q(o[473]) );
  DFF \Data_Mem/memory_reg[14][26]  ( .D(\Data_Mem/n7307 ), .CLK(clk), .RST(
        rst), .I(e_init[474]), .Q(o[474]) );
  DFF \Data_Mem/memory_reg[14][27]  ( .D(\Data_Mem/n7308 ), .CLK(clk), .RST(
        rst), .I(e_init[475]), .Q(o[475]) );
  DFF \Data_Mem/memory_reg[14][28]  ( .D(\Data_Mem/n7309 ), .CLK(clk), .RST(
        rst), .I(e_init[476]), .Q(o[476]) );
  DFF \Data_Mem/memory_reg[14][29]  ( .D(\Data_Mem/n7310 ), .CLK(clk), .RST(
        rst), .I(e_init[477]), .Q(o[477]) );
  DFF \Data_Mem/memory_reg[14][30]  ( .D(\Data_Mem/n7311 ), .CLK(clk), .RST(
        rst), .I(e_init[478]), .Q(o[478]) );
  DFF \Data_Mem/memory_reg[14][31]  ( .D(\Data_Mem/n7312 ), .CLK(clk), .RST(
        rst), .I(e_init[479]), .Q(o[479]) );
  DFF \Data_Mem/memory_reg[13][0]  ( .D(\Data_Mem/n7313 ), .CLK(clk), .RST(rst), .I(e_init[416]), .Q(o[416]) );
  DFF \Data_Mem/memory_reg[13][1]  ( .D(\Data_Mem/n7314 ), .CLK(clk), .RST(rst), .I(e_init[417]), .Q(o[417]) );
  DFF \Data_Mem/memory_reg[13][2]  ( .D(\Data_Mem/n7315 ), .CLK(clk), .RST(rst), .I(e_init[418]), .Q(o[418]) );
  DFF \Data_Mem/memory_reg[13][3]  ( .D(\Data_Mem/n7316 ), .CLK(clk), .RST(rst), .I(e_init[419]), .Q(o[419]) );
  DFF \Data_Mem/memory_reg[13][4]  ( .D(\Data_Mem/n7317 ), .CLK(clk), .RST(rst), .I(e_init[420]), .Q(o[420]) );
  DFF \Data_Mem/memory_reg[13][5]  ( .D(\Data_Mem/n7318 ), .CLK(clk), .RST(rst), .I(e_init[421]), .Q(o[421]) );
  DFF \Data_Mem/memory_reg[13][6]  ( .D(\Data_Mem/n7319 ), .CLK(clk), .RST(rst), .I(e_init[422]), .Q(o[422]) );
  DFF \Data_Mem/memory_reg[13][7]  ( .D(\Data_Mem/n7320 ), .CLK(clk), .RST(rst), .I(e_init[423]), .Q(o[423]) );
  DFF \Data_Mem/memory_reg[13][8]  ( .D(\Data_Mem/n7321 ), .CLK(clk), .RST(rst), .I(e_init[424]), .Q(o[424]) );
  DFF \Data_Mem/memory_reg[13][9]  ( .D(\Data_Mem/n7322 ), .CLK(clk), .RST(rst), .I(e_init[425]), .Q(o[425]) );
  DFF \Data_Mem/memory_reg[13][10]  ( .D(\Data_Mem/n7323 ), .CLK(clk), .RST(
        rst), .I(e_init[426]), .Q(o[426]) );
  DFF \Data_Mem/memory_reg[13][11]  ( .D(\Data_Mem/n7324 ), .CLK(clk), .RST(
        rst), .I(e_init[427]), .Q(o[427]) );
  DFF \Data_Mem/memory_reg[13][12]  ( .D(\Data_Mem/n7325 ), .CLK(clk), .RST(
        rst), .I(e_init[428]), .Q(o[428]) );
  DFF \Data_Mem/memory_reg[13][13]  ( .D(\Data_Mem/n7326 ), .CLK(clk), .RST(
        rst), .I(e_init[429]), .Q(o[429]) );
  DFF \Data_Mem/memory_reg[13][14]  ( .D(\Data_Mem/n7327 ), .CLK(clk), .RST(
        rst), .I(e_init[430]), .Q(o[430]) );
  DFF \Data_Mem/memory_reg[13][15]  ( .D(\Data_Mem/n7328 ), .CLK(clk), .RST(
        rst), .I(e_init[431]), .Q(o[431]) );
  DFF \Data_Mem/memory_reg[13][16]  ( .D(\Data_Mem/n7329 ), .CLK(clk), .RST(
        rst), .I(e_init[432]), .Q(o[432]) );
  DFF \Data_Mem/memory_reg[13][17]  ( .D(\Data_Mem/n7330 ), .CLK(clk), .RST(
        rst), .I(e_init[433]), .Q(o[433]) );
  DFF \Data_Mem/memory_reg[13][18]  ( .D(\Data_Mem/n7331 ), .CLK(clk), .RST(
        rst), .I(e_init[434]), .Q(o[434]) );
  DFF \Data_Mem/memory_reg[13][19]  ( .D(\Data_Mem/n7332 ), .CLK(clk), .RST(
        rst), .I(e_init[435]), .Q(o[435]) );
  DFF \Data_Mem/memory_reg[13][20]  ( .D(\Data_Mem/n7333 ), .CLK(clk), .RST(
        rst), .I(e_init[436]), .Q(o[436]) );
  DFF \Data_Mem/memory_reg[13][21]  ( .D(\Data_Mem/n7334 ), .CLK(clk), .RST(
        rst), .I(e_init[437]), .Q(o[437]) );
  DFF \Data_Mem/memory_reg[13][22]  ( .D(\Data_Mem/n7335 ), .CLK(clk), .RST(
        rst), .I(e_init[438]), .Q(o[438]) );
  DFF \Data_Mem/memory_reg[13][23]  ( .D(\Data_Mem/n7336 ), .CLK(clk), .RST(
        rst), .I(e_init[439]), .Q(o[439]) );
  DFF \Data_Mem/memory_reg[13][24]  ( .D(\Data_Mem/n7337 ), .CLK(clk), .RST(
        rst), .I(e_init[440]), .Q(o[440]) );
  DFF \Data_Mem/memory_reg[13][25]  ( .D(\Data_Mem/n7338 ), .CLK(clk), .RST(
        rst), .I(e_init[441]), .Q(o[441]) );
  DFF \Data_Mem/memory_reg[13][26]  ( .D(\Data_Mem/n7339 ), .CLK(clk), .RST(
        rst), .I(e_init[442]), .Q(o[442]) );
  DFF \Data_Mem/memory_reg[13][27]  ( .D(\Data_Mem/n7340 ), .CLK(clk), .RST(
        rst), .I(e_init[443]), .Q(o[443]) );
  DFF \Data_Mem/memory_reg[13][28]  ( .D(\Data_Mem/n7341 ), .CLK(clk), .RST(
        rst), .I(e_init[444]), .Q(o[444]) );
  DFF \Data_Mem/memory_reg[13][29]  ( .D(\Data_Mem/n7342 ), .CLK(clk), .RST(
        rst), .I(e_init[445]), .Q(o[445]) );
  DFF \Data_Mem/memory_reg[13][30]  ( .D(\Data_Mem/n7343 ), .CLK(clk), .RST(
        rst), .I(e_init[446]), .Q(o[446]) );
  DFF \Data_Mem/memory_reg[13][31]  ( .D(\Data_Mem/n7344 ), .CLK(clk), .RST(
        rst), .I(e_init[447]), .Q(o[447]) );
  DFF \Data_Mem/memory_reg[12][0]  ( .D(\Data_Mem/n7345 ), .CLK(clk), .RST(rst), .I(e_init[384]), .Q(o[384]) );
  DFF \Data_Mem/memory_reg[12][1]  ( .D(\Data_Mem/n7346 ), .CLK(clk), .RST(rst), .I(e_init[385]), .Q(o[385]) );
  DFF \Data_Mem/memory_reg[12][2]  ( .D(\Data_Mem/n7347 ), .CLK(clk), .RST(rst), .I(e_init[386]), .Q(o[386]) );
  DFF \Data_Mem/memory_reg[12][3]  ( .D(\Data_Mem/n7348 ), .CLK(clk), .RST(rst), .I(e_init[387]), .Q(o[387]) );
  DFF \Data_Mem/memory_reg[12][4]  ( .D(\Data_Mem/n7349 ), .CLK(clk), .RST(rst), .I(e_init[388]), .Q(o[388]) );
  DFF \Data_Mem/memory_reg[12][5]  ( .D(\Data_Mem/n7350 ), .CLK(clk), .RST(rst), .I(e_init[389]), .Q(o[389]) );
  DFF \Data_Mem/memory_reg[12][6]  ( .D(\Data_Mem/n7351 ), .CLK(clk), .RST(rst), .I(e_init[390]), .Q(o[390]) );
  DFF \Data_Mem/memory_reg[12][7]  ( .D(\Data_Mem/n7352 ), .CLK(clk), .RST(rst), .I(e_init[391]), .Q(o[391]) );
  DFF \Data_Mem/memory_reg[12][8]  ( .D(\Data_Mem/n7353 ), .CLK(clk), .RST(rst), .I(e_init[392]), .Q(o[392]) );
  DFF \Data_Mem/memory_reg[12][9]  ( .D(\Data_Mem/n7354 ), .CLK(clk), .RST(rst), .I(e_init[393]), .Q(o[393]) );
  DFF \Data_Mem/memory_reg[12][10]  ( .D(\Data_Mem/n7355 ), .CLK(clk), .RST(
        rst), .I(e_init[394]), .Q(o[394]) );
  DFF \Data_Mem/memory_reg[12][11]  ( .D(\Data_Mem/n7356 ), .CLK(clk), .RST(
        rst), .I(e_init[395]), .Q(o[395]) );
  DFF \Data_Mem/memory_reg[12][12]  ( .D(\Data_Mem/n7357 ), .CLK(clk), .RST(
        rst), .I(e_init[396]), .Q(o[396]) );
  DFF \Data_Mem/memory_reg[12][13]  ( .D(\Data_Mem/n7358 ), .CLK(clk), .RST(
        rst), .I(e_init[397]), .Q(o[397]) );
  DFF \Data_Mem/memory_reg[12][14]  ( .D(\Data_Mem/n7359 ), .CLK(clk), .RST(
        rst), .I(e_init[398]), .Q(o[398]) );
  DFF \Data_Mem/memory_reg[12][15]  ( .D(\Data_Mem/n7360 ), .CLK(clk), .RST(
        rst), .I(e_init[399]), .Q(o[399]) );
  DFF \Data_Mem/memory_reg[12][16]  ( .D(\Data_Mem/n7361 ), .CLK(clk), .RST(
        rst), .I(e_init[400]), .Q(o[400]) );
  DFF \Data_Mem/memory_reg[12][17]  ( .D(\Data_Mem/n7362 ), .CLK(clk), .RST(
        rst), .I(e_init[401]), .Q(o[401]) );
  DFF \Data_Mem/memory_reg[12][18]  ( .D(\Data_Mem/n7363 ), .CLK(clk), .RST(
        rst), .I(e_init[402]), .Q(o[402]) );
  DFF \Data_Mem/memory_reg[12][19]  ( .D(\Data_Mem/n7364 ), .CLK(clk), .RST(
        rst), .I(e_init[403]), .Q(o[403]) );
  DFF \Data_Mem/memory_reg[12][20]  ( .D(\Data_Mem/n7365 ), .CLK(clk), .RST(
        rst), .I(e_init[404]), .Q(o[404]) );
  DFF \Data_Mem/memory_reg[12][21]  ( .D(\Data_Mem/n7366 ), .CLK(clk), .RST(
        rst), .I(e_init[405]), .Q(o[405]) );
  DFF \Data_Mem/memory_reg[12][22]  ( .D(\Data_Mem/n7367 ), .CLK(clk), .RST(
        rst), .I(e_init[406]), .Q(o[406]) );
  DFF \Data_Mem/memory_reg[12][23]  ( .D(\Data_Mem/n7368 ), .CLK(clk), .RST(
        rst), .I(e_init[407]), .Q(o[407]) );
  DFF \Data_Mem/memory_reg[12][24]  ( .D(\Data_Mem/n7369 ), .CLK(clk), .RST(
        rst), .I(e_init[408]), .Q(o[408]) );
  DFF \Data_Mem/memory_reg[12][25]  ( .D(\Data_Mem/n7370 ), .CLK(clk), .RST(
        rst), .I(e_init[409]), .Q(o[409]) );
  DFF \Data_Mem/memory_reg[12][26]  ( .D(\Data_Mem/n7371 ), .CLK(clk), .RST(
        rst), .I(e_init[410]), .Q(o[410]) );
  DFF \Data_Mem/memory_reg[12][27]  ( .D(\Data_Mem/n7372 ), .CLK(clk), .RST(
        rst), .I(e_init[411]), .Q(o[411]) );
  DFF \Data_Mem/memory_reg[12][28]  ( .D(\Data_Mem/n7373 ), .CLK(clk), .RST(
        rst), .I(e_init[412]), .Q(o[412]) );
  DFF \Data_Mem/memory_reg[12][29]  ( .D(\Data_Mem/n7374 ), .CLK(clk), .RST(
        rst), .I(e_init[413]), .Q(o[413]) );
  DFF \Data_Mem/memory_reg[12][30]  ( .D(\Data_Mem/n7375 ), .CLK(clk), .RST(
        rst), .I(e_init[414]), .Q(o[414]) );
  DFF \Data_Mem/memory_reg[12][31]  ( .D(\Data_Mem/n7376 ), .CLK(clk), .RST(
        rst), .I(e_init[415]), .Q(o[415]) );
  DFF \Data_Mem/memory_reg[11][0]  ( .D(\Data_Mem/n7377 ), .CLK(clk), .RST(rst), .I(e_init[352]), .Q(o[352]) );
  DFF \Data_Mem/memory_reg[11][1]  ( .D(\Data_Mem/n7378 ), .CLK(clk), .RST(rst), .I(e_init[353]), .Q(o[353]) );
  DFF \Data_Mem/memory_reg[11][2]  ( .D(\Data_Mem/n7379 ), .CLK(clk), .RST(rst), .I(e_init[354]), .Q(o[354]) );
  DFF \Data_Mem/memory_reg[11][3]  ( .D(\Data_Mem/n7380 ), .CLK(clk), .RST(rst), .I(e_init[355]), .Q(o[355]) );
  DFF \Data_Mem/memory_reg[11][4]  ( .D(\Data_Mem/n7381 ), .CLK(clk), .RST(rst), .I(e_init[356]), .Q(o[356]) );
  DFF \Data_Mem/memory_reg[11][5]  ( .D(\Data_Mem/n7382 ), .CLK(clk), .RST(rst), .I(e_init[357]), .Q(o[357]) );
  DFF \Data_Mem/memory_reg[11][6]  ( .D(\Data_Mem/n7383 ), .CLK(clk), .RST(rst), .I(e_init[358]), .Q(o[358]) );
  DFF \Data_Mem/memory_reg[11][7]  ( .D(\Data_Mem/n7384 ), .CLK(clk), .RST(rst), .I(e_init[359]), .Q(o[359]) );
  DFF \Data_Mem/memory_reg[11][8]  ( .D(\Data_Mem/n7385 ), .CLK(clk), .RST(rst), .I(e_init[360]), .Q(o[360]) );
  DFF \Data_Mem/memory_reg[11][9]  ( .D(\Data_Mem/n7386 ), .CLK(clk), .RST(rst), .I(e_init[361]), .Q(o[361]) );
  DFF \Data_Mem/memory_reg[11][10]  ( .D(\Data_Mem/n7387 ), .CLK(clk), .RST(
        rst), .I(e_init[362]), .Q(o[362]) );
  DFF \Data_Mem/memory_reg[11][11]  ( .D(\Data_Mem/n7388 ), .CLK(clk), .RST(
        rst), .I(e_init[363]), .Q(o[363]) );
  DFF \Data_Mem/memory_reg[11][12]  ( .D(\Data_Mem/n7389 ), .CLK(clk), .RST(
        rst), .I(e_init[364]), .Q(o[364]) );
  DFF \Data_Mem/memory_reg[11][13]  ( .D(\Data_Mem/n7390 ), .CLK(clk), .RST(
        rst), .I(e_init[365]), .Q(o[365]) );
  DFF \Data_Mem/memory_reg[11][14]  ( .D(\Data_Mem/n7391 ), .CLK(clk), .RST(
        rst), .I(e_init[366]), .Q(o[366]) );
  DFF \Data_Mem/memory_reg[11][15]  ( .D(\Data_Mem/n7392 ), .CLK(clk), .RST(
        rst), .I(e_init[367]), .Q(o[367]) );
  DFF \Data_Mem/memory_reg[11][16]  ( .D(\Data_Mem/n7393 ), .CLK(clk), .RST(
        rst), .I(e_init[368]), .Q(o[368]) );
  DFF \Data_Mem/memory_reg[11][17]  ( .D(\Data_Mem/n7394 ), .CLK(clk), .RST(
        rst), .I(e_init[369]), .Q(o[369]) );
  DFF \Data_Mem/memory_reg[11][18]  ( .D(\Data_Mem/n7395 ), .CLK(clk), .RST(
        rst), .I(e_init[370]), .Q(o[370]) );
  DFF \Data_Mem/memory_reg[11][19]  ( .D(\Data_Mem/n7396 ), .CLK(clk), .RST(
        rst), .I(e_init[371]), .Q(o[371]) );
  DFF \Data_Mem/memory_reg[11][20]  ( .D(\Data_Mem/n7397 ), .CLK(clk), .RST(
        rst), .I(e_init[372]), .Q(o[372]) );
  DFF \Data_Mem/memory_reg[11][21]  ( .D(\Data_Mem/n7398 ), .CLK(clk), .RST(
        rst), .I(e_init[373]), .Q(o[373]) );
  DFF \Data_Mem/memory_reg[11][22]  ( .D(\Data_Mem/n7399 ), .CLK(clk), .RST(
        rst), .I(e_init[374]), .Q(o[374]) );
  DFF \Data_Mem/memory_reg[11][23]  ( .D(\Data_Mem/n7400 ), .CLK(clk), .RST(
        rst), .I(e_init[375]), .Q(o[375]) );
  DFF \Data_Mem/memory_reg[11][24]  ( .D(\Data_Mem/n7401 ), .CLK(clk), .RST(
        rst), .I(e_init[376]), .Q(o[376]) );
  DFF \Data_Mem/memory_reg[11][25]  ( .D(\Data_Mem/n7402 ), .CLK(clk), .RST(
        rst), .I(e_init[377]), .Q(o[377]) );
  DFF \Data_Mem/memory_reg[11][26]  ( .D(\Data_Mem/n7403 ), .CLK(clk), .RST(
        rst), .I(e_init[378]), .Q(o[378]) );
  DFF \Data_Mem/memory_reg[11][27]  ( .D(\Data_Mem/n7404 ), .CLK(clk), .RST(
        rst), .I(e_init[379]), .Q(o[379]) );
  DFF \Data_Mem/memory_reg[11][28]  ( .D(\Data_Mem/n7405 ), .CLK(clk), .RST(
        rst), .I(e_init[380]), .Q(o[380]) );
  DFF \Data_Mem/memory_reg[11][29]  ( .D(\Data_Mem/n7406 ), .CLK(clk), .RST(
        rst), .I(e_init[381]), .Q(o[381]) );
  DFF \Data_Mem/memory_reg[11][30]  ( .D(\Data_Mem/n7407 ), .CLK(clk), .RST(
        rst), .I(e_init[382]), .Q(o[382]) );
  DFF \Data_Mem/memory_reg[11][31]  ( .D(\Data_Mem/n7408 ), .CLK(clk), .RST(
        rst), .I(e_init[383]), .Q(o[383]) );
  DFF \Data_Mem/memory_reg[10][0]  ( .D(\Data_Mem/n7409 ), .CLK(clk), .RST(rst), .I(e_init[320]), .Q(o[320]) );
  DFF \Data_Mem/memory_reg[10][1]  ( .D(\Data_Mem/n7410 ), .CLK(clk), .RST(rst), .I(e_init[321]), .Q(o[321]) );
  DFF \Data_Mem/memory_reg[10][2]  ( .D(\Data_Mem/n7411 ), .CLK(clk), .RST(rst), .I(e_init[322]), .Q(o[322]) );
  DFF \Data_Mem/memory_reg[10][3]  ( .D(\Data_Mem/n7412 ), .CLK(clk), .RST(rst), .I(e_init[323]), .Q(o[323]) );
  DFF \Data_Mem/memory_reg[10][4]  ( .D(\Data_Mem/n7413 ), .CLK(clk), .RST(rst), .I(e_init[324]), .Q(o[324]) );
  DFF \Data_Mem/memory_reg[10][5]  ( .D(\Data_Mem/n7414 ), .CLK(clk), .RST(rst), .I(e_init[325]), .Q(o[325]) );
  DFF \Data_Mem/memory_reg[10][6]  ( .D(\Data_Mem/n7415 ), .CLK(clk), .RST(rst), .I(e_init[326]), .Q(o[326]) );
  DFF \Data_Mem/memory_reg[10][7]  ( .D(\Data_Mem/n7416 ), .CLK(clk), .RST(rst), .I(e_init[327]), .Q(o[327]) );
  DFF \Data_Mem/memory_reg[10][8]  ( .D(\Data_Mem/n7417 ), .CLK(clk), .RST(rst), .I(e_init[328]), .Q(o[328]) );
  DFF \Data_Mem/memory_reg[10][9]  ( .D(\Data_Mem/n7418 ), .CLK(clk), .RST(rst), .I(e_init[329]), .Q(o[329]) );
  DFF \Data_Mem/memory_reg[10][10]  ( .D(\Data_Mem/n7419 ), .CLK(clk), .RST(
        rst), .I(e_init[330]), .Q(o[330]) );
  DFF \Data_Mem/memory_reg[10][11]  ( .D(\Data_Mem/n7420 ), .CLK(clk), .RST(
        rst), .I(e_init[331]), .Q(o[331]) );
  DFF \Data_Mem/memory_reg[10][12]  ( .D(\Data_Mem/n7421 ), .CLK(clk), .RST(
        rst), .I(e_init[332]), .Q(o[332]) );
  DFF \Data_Mem/memory_reg[10][13]  ( .D(\Data_Mem/n7422 ), .CLK(clk), .RST(
        rst), .I(e_init[333]), .Q(o[333]) );
  DFF \Data_Mem/memory_reg[10][14]  ( .D(\Data_Mem/n7423 ), .CLK(clk), .RST(
        rst), .I(e_init[334]), .Q(o[334]) );
  DFF \Data_Mem/memory_reg[10][15]  ( .D(\Data_Mem/n7424 ), .CLK(clk), .RST(
        rst), .I(e_init[335]), .Q(o[335]) );
  DFF \Data_Mem/memory_reg[10][16]  ( .D(\Data_Mem/n7425 ), .CLK(clk), .RST(
        rst), .I(e_init[336]), .Q(o[336]) );
  DFF \Data_Mem/memory_reg[10][17]  ( .D(\Data_Mem/n7426 ), .CLK(clk), .RST(
        rst), .I(e_init[337]), .Q(o[337]) );
  DFF \Data_Mem/memory_reg[10][18]  ( .D(\Data_Mem/n7427 ), .CLK(clk), .RST(
        rst), .I(e_init[338]), .Q(o[338]) );
  DFF \Data_Mem/memory_reg[10][19]  ( .D(\Data_Mem/n7428 ), .CLK(clk), .RST(
        rst), .I(e_init[339]), .Q(o[339]) );
  DFF \Data_Mem/memory_reg[10][20]  ( .D(\Data_Mem/n7429 ), .CLK(clk), .RST(
        rst), .I(e_init[340]), .Q(o[340]) );
  DFF \Data_Mem/memory_reg[10][21]  ( .D(\Data_Mem/n7430 ), .CLK(clk), .RST(
        rst), .I(e_init[341]), .Q(o[341]) );
  DFF \Data_Mem/memory_reg[10][22]  ( .D(\Data_Mem/n7431 ), .CLK(clk), .RST(
        rst), .I(e_init[342]), .Q(o[342]) );
  DFF \Data_Mem/memory_reg[10][23]  ( .D(\Data_Mem/n7432 ), .CLK(clk), .RST(
        rst), .I(e_init[343]), .Q(o[343]) );
  DFF \Data_Mem/memory_reg[10][24]  ( .D(\Data_Mem/n7433 ), .CLK(clk), .RST(
        rst), .I(e_init[344]), .Q(o[344]) );
  DFF \Data_Mem/memory_reg[10][25]  ( .D(\Data_Mem/n7434 ), .CLK(clk), .RST(
        rst), .I(e_init[345]), .Q(o[345]) );
  DFF \Data_Mem/memory_reg[10][26]  ( .D(\Data_Mem/n7435 ), .CLK(clk), .RST(
        rst), .I(e_init[346]), .Q(o[346]) );
  DFF \Data_Mem/memory_reg[10][27]  ( .D(\Data_Mem/n7436 ), .CLK(clk), .RST(
        rst), .I(e_init[347]), .Q(o[347]) );
  DFF \Data_Mem/memory_reg[10][28]  ( .D(\Data_Mem/n7437 ), .CLK(clk), .RST(
        rst), .I(e_init[348]), .Q(o[348]) );
  DFF \Data_Mem/memory_reg[10][29]  ( .D(\Data_Mem/n7438 ), .CLK(clk), .RST(
        rst), .I(e_init[349]), .Q(o[349]) );
  DFF \Data_Mem/memory_reg[10][30]  ( .D(\Data_Mem/n7439 ), .CLK(clk), .RST(
        rst), .I(e_init[350]), .Q(o[350]) );
  DFF \Data_Mem/memory_reg[10][31]  ( .D(\Data_Mem/n7440 ), .CLK(clk), .RST(
        rst), .I(e_init[351]), .Q(o[351]) );
  DFF \Data_Mem/memory_reg[9][0]  ( .D(\Data_Mem/n7441 ), .CLK(clk), .RST(rst), 
        .I(e_init[288]), .Q(o[288]) );
  DFF \Data_Mem/memory_reg[9][1]  ( .D(\Data_Mem/n7442 ), .CLK(clk), .RST(rst), 
        .I(e_init[289]), .Q(o[289]) );
  DFF \Data_Mem/memory_reg[9][2]  ( .D(\Data_Mem/n7443 ), .CLK(clk), .RST(rst), 
        .I(e_init[290]), .Q(o[290]) );
  DFF \Data_Mem/memory_reg[9][3]  ( .D(\Data_Mem/n7444 ), .CLK(clk), .RST(rst), 
        .I(e_init[291]), .Q(o[291]) );
  DFF \Data_Mem/memory_reg[9][4]  ( .D(\Data_Mem/n7445 ), .CLK(clk), .RST(rst), 
        .I(e_init[292]), .Q(o[292]) );
  DFF \Data_Mem/memory_reg[9][5]  ( .D(\Data_Mem/n7446 ), .CLK(clk), .RST(rst), 
        .I(e_init[293]), .Q(o[293]) );
  DFF \Data_Mem/memory_reg[9][6]  ( .D(\Data_Mem/n7447 ), .CLK(clk), .RST(rst), 
        .I(e_init[294]), .Q(o[294]) );
  DFF \Data_Mem/memory_reg[9][7]  ( .D(\Data_Mem/n7448 ), .CLK(clk), .RST(rst), 
        .I(e_init[295]), .Q(o[295]) );
  DFF \Data_Mem/memory_reg[9][8]  ( .D(\Data_Mem/n7449 ), .CLK(clk), .RST(rst), 
        .I(e_init[296]), .Q(o[296]) );
  DFF \Data_Mem/memory_reg[9][9]  ( .D(\Data_Mem/n7450 ), .CLK(clk), .RST(rst), 
        .I(e_init[297]), .Q(o[297]) );
  DFF \Data_Mem/memory_reg[9][10]  ( .D(\Data_Mem/n7451 ), .CLK(clk), .RST(rst), .I(e_init[298]), .Q(o[298]) );
  DFF \Data_Mem/memory_reg[9][11]  ( .D(\Data_Mem/n7452 ), .CLK(clk), .RST(rst), .I(e_init[299]), .Q(o[299]) );
  DFF \Data_Mem/memory_reg[9][12]  ( .D(\Data_Mem/n7453 ), .CLK(clk), .RST(rst), .I(e_init[300]), .Q(o[300]) );
  DFF \Data_Mem/memory_reg[9][13]  ( .D(\Data_Mem/n7454 ), .CLK(clk), .RST(rst), .I(e_init[301]), .Q(o[301]) );
  DFF \Data_Mem/memory_reg[9][14]  ( .D(\Data_Mem/n7455 ), .CLK(clk), .RST(rst), .I(e_init[302]), .Q(o[302]) );
  DFF \Data_Mem/memory_reg[9][15]  ( .D(\Data_Mem/n7456 ), .CLK(clk), .RST(rst), .I(e_init[303]), .Q(o[303]) );
  DFF \Data_Mem/memory_reg[9][16]  ( .D(\Data_Mem/n7457 ), .CLK(clk), .RST(rst), .I(e_init[304]), .Q(o[304]) );
  DFF \Data_Mem/memory_reg[9][17]  ( .D(\Data_Mem/n7458 ), .CLK(clk), .RST(rst), .I(e_init[305]), .Q(o[305]) );
  DFF \Data_Mem/memory_reg[9][18]  ( .D(\Data_Mem/n7459 ), .CLK(clk), .RST(rst), .I(e_init[306]), .Q(o[306]) );
  DFF \Data_Mem/memory_reg[9][19]  ( .D(\Data_Mem/n7460 ), .CLK(clk), .RST(rst), .I(e_init[307]), .Q(o[307]) );
  DFF \Data_Mem/memory_reg[9][20]  ( .D(\Data_Mem/n7461 ), .CLK(clk), .RST(rst), .I(e_init[308]), .Q(o[308]) );
  DFF \Data_Mem/memory_reg[9][21]  ( .D(\Data_Mem/n7462 ), .CLK(clk), .RST(rst), .I(e_init[309]), .Q(o[309]) );
  DFF \Data_Mem/memory_reg[9][22]  ( .D(\Data_Mem/n7463 ), .CLK(clk), .RST(rst), .I(e_init[310]), .Q(o[310]) );
  DFF \Data_Mem/memory_reg[9][23]  ( .D(\Data_Mem/n7464 ), .CLK(clk), .RST(rst), .I(e_init[311]), .Q(o[311]) );
  DFF \Data_Mem/memory_reg[9][24]  ( .D(\Data_Mem/n7465 ), .CLK(clk), .RST(rst), .I(e_init[312]), .Q(o[312]) );
  DFF \Data_Mem/memory_reg[9][25]  ( .D(\Data_Mem/n7466 ), .CLK(clk), .RST(rst), .I(e_init[313]), .Q(o[313]) );
  DFF \Data_Mem/memory_reg[9][26]  ( .D(\Data_Mem/n7467 ), .CLK(clk), .RST(rst), .I(e_init[314]), .Q(o[314]) );
  DFF \Data_Mem/memory_reg[9][27]  ( .D(\Data_Mem/n7468 ), .CLK(clk), .RST(rst), .I(e_init[315]), .Q(o[315]) );
  DFF \Data_Mem/memory_reg[9][28]  ( .D(\Data_Mem/n7469 ), .CLK(clk), .RST(rst), .I(e_init[316]), .Q(o[316]) );
  DFF \Data_Mem/memory_reg[9][29]  ( .D(\Data_Mem/n7470 ), .CLK(clk), .RST(rst), .I(e_init[317]), .Q(o[317]) );
  DFF \Data_Mem/memory_reg[9][30]  ( .D(\Data_Mem/n7471 ), .CLK(clk), .RST(rst), .I(e_init[318]), .Q(o[318]) );
  DFF \Data_Mem/memory_reg[9][31]  ( .D(\Data_Mem/n7472 ), .CLK(clk), .RST(rst), .I(e_init[319]), .Q(o[319]) );
  DFF \Data_Mem/memory_reg[8][0]  ( .D(\Data_Mem/n7473 ), .CLK(clk), .RST(rst), 
        .I(e_init[256]), .Q(o[256]) );
  DFF \Data_Mem/memory_reg[8][1]  ( .D(\Data_Mem/n7474 ), .CLK(clk), .RST(rst), 
        .I(e_init[257]), .Q(o[257]) );
  DFF \Data_Mem/memory_reg[8][2]  ( .D(\Data_Mem/n7475 ), .CLK(clk), .RST(rst), 
        .I(e_init[258]), .Q(o[258]) );
  DFF \Data_Mem/memory_reg[8][3]  ( .D(\Data_Mem/n7476 ), .CLK(clk), .RST(rst), 
        .I(e_init[259]), .Q(o[259]) );
  DFF \Data_Mem/memory_reg[8][4]  ( .D(\Data_Mem/n7477 ), .CLK(clk), .RST(rst), 
        .I(e_init[260]), .Q(o[260]) );
  DFF \Data_Mem/memory_reg[8][5]  ( .D(\Data_Mem/n7478 ), .CLK(clk), .RST(rst), 
        .I(e_init[261]), .Q(o[261]) );
  DFF \Data_Mem/memory_reg[8][6]  ( .D(\Data_Mem/n7479 ), .CLK(clk), .RST(rst), 
        .I(e_init[262]), .Q(o[262]) );
  DFF \Data_Mem/memory_reg[8][7]  ( .D(\Data_Mem/n7480 ), .CLK(clk), .RST(rst), 
        .I(e_init[263]), .Q(o[263]) );
  DFF \Data_Mem/memory_reg[8][8]  ( .D(\Data_Mem/n7481 ), .CLK(clk), .RST(rst), 
        .I(e_init[264]), .Q(o[264]) );
  DFF \Data_Mem/memory_reg[8][9]  ( .D(\Data_Mem/n7482 ), .CLK(clk), .RST(rst), 
        .I(e_init[265]), .Q(o[265]) );
  DFF \Data_Mem/memory_reg[8][10]  ( .D(\Data_Mem/n7483 ), .CLK(clk), .RST(rst), .I(e_init[266]), .Q(o[266]) );
  DFF \Data_Mem/memory_reg[8][11]  ( .D(\Data_Mem/n7484 ), .CLK(clk), .RST(rst), .I(e_init[267]), .Q(o[267]) );
  DFF \Data_Mem/memory_reg[8][12]  ( .D(\Data_Mem/n7485 ), .CLK(clk), .RST(rst), .I(e_init[268]), .Q(o[268]) );
  DFF \Data_Mem/memory_reg[8][13]  ( .D(\Data_Mem/n7486 ), .CLK(clk), .RST(rst), .I(e_init[269]), .Q(o[269]) );
  DFF \Data_Mem/memory_reg[8][14]  ( .D(\Data_Mem/n7487 ), .CLK(clk), .RST(rst), .I(e_init[270]), .Q(o[270]) );
  DFF \Data_Mem/memory_reg[8][15]  ( .D(\Data_Mem/n7488 ), .CLK(clk), .RST(rst), .I(e_init[271]), .Q(o[271]) );
  DFF \Data_Mem/memory_reg[8][16]  ( .D(\Data_Mem/n7489 ), .CLK(clk), .RST(rst), .I(e_init[272]), .Q(o[272]) );
  DFF \Data_Mem/memory_reg[8][17]  ( .D(\Data_Mem/n7490 ), .CLK(clk), .RST(rst), .I(e_init[273]), .Q(o[273]) );
  DFF \Data_Mem/memory_reg[8][18]  ( .D(\Data_Mem/n7491 ), .CLK(clk), .RST(rst), .I(e_init[274]), .Q(o[274]) );
  DFF \Data_Mem/memory_reg[8][19]  ( .D(\Data_Mem/n7492 ), .CLK(clk), .RST(rst), .I(e_init[275]), .Q(o[275]) );
  DFF \Data_Mem/memory_reg[8][20]  ( .D(\Data_Mem/n7493 ), .CLK(clk), .RST(rst), .I(e_init[276]), .Q(o[276]) );
  DFF \Data_Mem/memory_reg[8][21]  ( .D(\Data_Mem/n7494 ), .CLK(clk), .RST(rst), .I(e_init[277]), .Q(o[277]) );
  DFF \Data_Mem/memory_reg[8][22]  ( .D(\Data_Mem/n7495 ), .CLK(clk), .RST(rst), .I(e_init[278]), .Q(o[278]) );
  DFF \Data_Mem/memory_reg[8][23]  ( .D(\Data_Mem/n7496 ), .CLK(clk), .RST(rst), .I(e_init[279]), .Q(o[279]) );
  DFF \Data_Mem/memory_reg[8][24]  ( .D(\Data_Mem/n7497 ), .CLK(clk), .RST(rst), .I(e_init[280]), .Q(o[280]) );
  DFF \Data_Mem/memory_reg[8][25]  ( .D(\Data_Mem/n7498 ), .CLK(clk), .RST(rst), .I(e_init[281]), .Q(o[281]) );
  DFF \Data_Mem/memory_reg[8][26]  ( .D(\Data_Mem/n7499 ), .CLK(clk), .RST(rst), .I(e_init[282]), .Q(o[282]) );
  DFF \Data_Mem/memory_reg[8][27]  ( .D(\Data_Mem/n7500 ), .CLK(clk), .RST(rst), .I(e_init[283]), .Q(o[283]) );
  DFF \Data_Mem/memory_reg[8][28]  ( .D(\Data_Mem/n7501 ), .CLK(clk), .RST(rst), .I(e_init[284]), .Q(o[284]) );
  DFF \Data_Mem/memory_reg[8][29]  ( .D(\Data_Mem/n7502 ), .CLK(clk), .RST(rst), .I(e_init[285]), .Q(o[285]) );
  DFF \Data_Mem/memory_reg[8][30]  ( .D(\Data_Mem/n7503 ), .CLK(clk), .RST(rst), .I(e_init[286]), .Q(o[286]) );
  DFF \Data_Mem/memory_reg[8][31]  ( .D(\Data_Mem/n7504 ), .CLK(clk), .RST(rst), .I(e_init[287]), .Q(o[287]) );
  DFF \Data_Mem/memory_reg[7][0]  ( .D(\Data_Mem/n7505 ), .CLK(clk), .RST(rst), 
        .I(e_init[224]), .Q(o[224]) );
  DFF \Data_Mem/memory_reg[7][1]  ( .D(\Data_Mem/n7506 ), .CLK(clk), .RST(rst), 
        .I(e_init[225]), .Q(o[225]) );
  DFF \Data_Mem/memory_reg[7][2]  ( .D(\Data_Mem/n7507 ), .CLK(clk), .RST(rst), 
        .I(e_init[226]), .Q(o[226]) );
  DFF \Data_Mem/memory_reg[7][3]  ( .D(\Data_Mem/n7508 ), .CLK(clk), .RST(rst), 
        .I(e_init[227]), .Q(o[227]) );
  DFF \Data_Mem/memory_reg[7][4]  ( .D(\Data_Mem/n7509 ), .CLK(clk), .RST(rst), 
        .I(e_init[228]), .Q(o[228]) );
  DFF \Data_Mem/memory_reg[7][5]  ( .D(\Data_Mem/n7510 ), .CLK(clk), .RST(rst), 
        .I(e_init[229]), .Q(o[229]) );
  DFF \Data_Mem/memory_reg[7][6]  ( .D(\Data_Mem/n7511 ), .CLK(clk), .RST(rst), 
        .I(e_init[230]), .Q(o[230]) );
  DFF \Data_Mem/memory_reg[7][7]  ( .D(\Data_Mem/n7512 ), .CLK(clk), .RST(rst), 
        .I(e_init[231]), .Q(o[231]) );
  DFF \Data_Mem/memory_reg[7][8]  ( .D(\Data_Mem/n7513 ), .CLK(clk), .RST(rst), 
        .I(e_init[232]), .Q(o[232]) );
  DFF \Data_Mem/memory_reg[7][9]  ( .D(\Data_Mem/n7514 ), .CLK(clk), .RST(rst), 
        .I(e_init[233]), .Q(o[233]) );
  DFF \Data_Mem/memory_reg[7][10]  ( .D(\Data_Mem/n7515 ), .CLK(clk), .RST(rst), .I(e_init[234]), .Q(o[234]) );
  DFF \Data_Mem/memory_reg[7][11]  ( .D(\Data_Mem/n7516 ), .CLK(clk), .RST(rst), .I(e_init[235]), .Q(o[235]) );
  DFF \Data_Mem/memory_reg[7][12]  ( .D(\Data_Mem/n7517 ), .CLK(clk), .RST(rst), .I(e_init[236]), .Q(o[236]) );
  DFF \Data_Mem/memory_reg[7][13]  ( .D(\Data_Mem/n7518 ), .CLK(clk), .RST(rst), .I(e_init[237]), .Q(o[237]) );
  DFF \Data_Mem/memory_reg[7][14]  ( .D(\Data_Mem/n7519 ), .CLK(clk), .RST(rst), .I(e_init[238]), .Q(o[238]) );
  DFF \Data_Mem/memory_reg[7][15]  ( .D(\Data_Mem/n7520 ), .CLK(clk), .RST(rst), .I(e_init[239]), .Q(o[239]) );
  DFF \Data_Mem/memory_reg[7][16]  ( .D(\Data_Mem/n7521 ), .CLK(clk), .RST(rst), .I(e_init[240]), .Q(o[240]) );
  DFF \Data_Mem/memory_reg[7][17]  ( .D(\Data_Mem/n7522 ), .CLK(clk), .RST(rst), .I(e_init[241]), .Q(o[241]) );
  DFF \Data_Mem/memory_reg[7][18]  ( .D(\Data_Mem/n7523 ), .CLK(clk), .RST(rst), .I(e_init[242]), .Q(o[242]) );
  DFF \Data_Mem/memory_reg[7][19]  ( .D(\Data_Mem/n7524 ), .CLK(clk), .RST(rst), .I(e_init[243]), .Q(o[243]) );
  DFF \Data_Mem/memory_reg[7][20]  ( .D(\Data_Mem/n7525 ), .CLK(clk), .RST(rst), .I(e_init[244]), .Q(o[244]) );
  DFF \Data_Mem/memory_reg[7][21]  ( .D(\Data_Mem/n7526 ), .CLK(clk), .RST(rst), .I(e_init[245]), .Q(o[245]) );
  DFF \Data_Mem/memory_reg[7][22]  ( .D(\Data_Mem/n7527 ), .CLK(clk), .RST(rst), .I(e_init[246]), .Q(o[246]) );
  DFF \Data_Mem/memory_reg[7][23]  ( .D(\Data_Mem/n7528 ), .CLK(clk), .RST(rst), .I(e_init[247]), .Q(o[247]) );
  DFF \Data_Mem/memory_reg[7][24]  ( .D(\Data_Mem/n7529 ), .CLK(clk), .RST(rst), .I(e_init[248]), .Q(o[248]) );
  DFF \Data_Mem/memory_reg[7][25]  ( .D(\Data_Mem/n7530 ), .CLK(clk), .RST(rst), .I(e_init[249]), .Q(o[249]) );
  DFF \Data_Mem/memory_reg[7][26]  ( .D(\Data_Mem/n7531 ), .CLK(clk), .RST(rst), .I(e_init[250]), .Q(o[250]) );
  DFF \Data_Mem/memory_reg[7][27]  ( .D(\Data_Mem/n7532 ), .CLK(clk), .RST(rst), .I(e_init[251]), .Q(o[251]) );
  DFF \Data_Mem/memory_reg[7][28]  ( .D(\Data_Mem/n7533 ), .CLK(clk), .RST(rst), .I(e_init[252]), .Q(o[252]) );
  DFF \Data_Mem/memory_reg[7][29]  ( .D(\Data_Mem/n7534 ), .CLK(clk), .RST(rst), .I(e_init[253]), .Q(o[253]) );
  DFF \Data_Mem/memory_reg[7][30]  ( .D(\Data_Mem/n7535 ), .CLK(clk), .RST(rst), .I(e_init[254]), .Q(o[254]) );
  DFF \Data_Mem/memory_reg[7][31]  ( .D(\Data_Mem/n7536 ), .CLK(clk), .RST(rst), .I(e_init[255]), .Q(o[255]) );
  DFF \Data_Mem/memory_reg[6][0]  ( .D(\Data_Mem/n7537 ), .CLK(clk), .RST(rst), 
        .I(e_init[192]), .Q(o[192]) );
  DFF \Data_Mem/memory_reg[6][1]  ( .D(\Data_Mem/n7538 ), .CLK(clk), .RST(rst), 
        .I(e_init[193]), .Q(o[193]) );
  DFF \Data_Mem/memory_reg[6][2]  ( .D(\Data_Mem/n7539 ), .CLK(clk), .RST(rst), 
        .I(e_init[194]), .Q(o[194]) );
  DFF \Data_Mem/memory_reg[6][3]  ( .D(\Data_Mem/n7540 ), .CLK(clk), .RST(rst), 
        .I(e_init[195]), .Q(o[195]) );
  DFF \Data_Mem/memory_reg[6][4]  ( .D(\Data_Mem/n7541 ), .CLK(clk), .RST(rst), 
        .I(e_init[196]), .Q(o[196]) );
  DFF \Data_Mem/memory_reg[6][5]  ( .D(\Data_Mem/n7542 ), .CLK(clk), .RST(rst), 
        .I(e_init[197]), .Q(o[197]) );
  DFF \Data_Mem/memory_reg[6][6]  ( .D(\Data_Mem/n7543 ), .CLK(clk), .RST(rst), 
        .I(e_init[198]), .Q(o[198]) );
  DFF \Data_Mem/memory_reg[6][7]  ( .D(\Data_Mem/n7544 ), .CLK(clk), .RST(rst), 
        .I(e_init[199]), .Q(o[199]) );
  DFF \Data_Mem/memory_reg[6][8]  ( .D(\Data_Mem/n7545 ), .CLK(clk), .RST(rst), 
        .I(e_init[200]), .Q(o[200]) );
  DFF \Data_Mem/memory_reg[6][9]  ( .D(\Data_Mem/n7546 ), .CLK(clk), .RST(rst), 
        .I(e_init[201]), .Q(o[201]) );
  DFF \Data_Mem/memory_reg[6][10]  ( .D(\Data_Mem/n7547 ), .CLK(clk), .RST(rst), .I(e_init[202]), .Q(o[202]) );
  DFF \Data_Mem/memory_reg[6][11]  ( .D(\Data_Mem/n7548 ), .CLK(clk), .RST(rst), .I(e_init[203]), .Q(o[203]) );
  DFF \Data_Mem/memory_reg[6][12]  ( .D(\Data_Mem/n7549 ), .CLK(clk), .RST(rst), .I(e_init[204]), .Q(o[204]) );
  DFF \Data_Mem/memory_reg[6][13]  ( .D(\Data_Mem/n7550 ), .CLK(clk), .RST(rst), .I(e_init[205]), .Q(o[205]) );
  DFF \Data_Mem/memory_reg[6][14]  ( .D(\Data_Mem/n7551 ), .CLK(clk), .RST(rst), .I(e_init[206]), .Q(o[206]) );
  DFF \Data_Mem/memory_reg[6][15]  ( .D(\Data_Mem/n7552 ), .CLK(clk), .RST(rst), .I(e_init[207]), .Q(o[207]) );
  DFF \Data_Mem/memory_reg[6][16]  ( .D(\Data_Mem/n7553 ), .CLK(clk), .RST(rst), .I(e_init[208]), .Q(o[208]) );
  DFF \Data_Mem/memory_reg[6][17]  ( .D(\Data_Mem/n7554 ), .CLK(clk), .RST(rst), .I(e_init[209]), .Q(o[209]) );
  DFF \Data_Mem/memory_reg[6][18]  ( .D(\Data_Mem/n7555 ), .CLK(clk), .RST(rst), .I(e_init[210]), .Q(o[210]) );
  DFF \Data_Mem/memory_reg[6][19]  ( .D(\Data_Mem/n7556 ), .CLK(clk), .RST(rst), .I(e_init[211]), .Q(o[211]) );
  DFF \Data_Mem/memory_reg[6][20]  ( .D(\Data_Mem/n7557 ), .CLK(clk), .RST(rst), .I(e_init[212]), .Q(o[212]) );
  DFF \Data_Mem/memory_reg[6][21]  ( .D(\Data_Mem/n7558 ), .CLK(clk), .RST(rst), .I(e_init[213]), .Q(o[213]) );
  DFF \Data_Mem/memory_reg[6][22]  ( .D(\Data_Mem/n7559 ), .CLK(clk), .RST(rst), .I(e_init[214]), .Q(o[214]) );
  DFF \Data_Mem/memory_reg[6][23]  ( .D(\Data_Mem/n7560 ), .CLK(clk), .RST(rst), .I(e_init[215]), .Q(o[215]) );
  DFF \Data_Mem/memory_reg[6][24]  ( .D(\Data_Mem/n7561 ), .CLK(clk), .RST(rst), .I(e_init[216]), .Q(o[216]) );
  DFF \Data_Mem/memory_reg[6][25]  ( .D(\Data_Mem/n7562 ), .CLK(clk), .RST(rst), .I(e_init[217]), .Q(o[217]) );
  DFF \Data_Mem/memory_reg[6][26]  ( .D(\Data_Mem/n7563 ), .CLK(clk), .RST(rst), .I(e_init[218]), .Q(o[218]) );
  DFF \Data_Mem/memory_reg[6][27]  ( .D(\Data_Mem/n7564 ), .CLK(clk), .RST(rst), .I(e_init[219]), .Q(o[219]) );
  DFF \Data_Mem/memory_reg[6][28]  ( .D(\Data_Mem/n7565 ), .CLK(clk), .RST(rst), .I(e_init[220]), .Q(o[220]) );
  DFF \Data_Mem/memory_reg[6][29]  ( .D(\Data_Mem/n7566 ), .CLK(clk), .RST(rst), .I(e_init[221]), .Q(o[221]) );
  DFF \Data_Mem/memory_reg[6][30]  ( .D(\Data_Mem/n7567 ), .CLK(clk), .RST(rst), .I(e_init[222]), .Q(o[222]) );
  DFF \Data_Mem/memory_reg[6][31]  ( .D(\Data_Mem/n7568 ), .CLK(clk), .RST(rst), .I(e_init[223]), .Q(o[223]) );
  DFF \Data_Mem/memory_reg[5][0]  ( .D(\Data_Mem/n7569 ), .CLK(clk), .RST(rst), 
        .I(e_init[160]), .Q(o[160]) );
  DFF \Data_Mem/memory_reg[5][1]  ( .D(\Data_Mem/n7570 ), .CLK(clk), .RST(rst), 
        .I(e_init[161]), .Q(o[161]) );
  DFF \Data_Mem/memory_reg[5][2]  ( .D(\Data_Mem/n7571 ), .CLK(clk), .RST(rst), 
        .I(e_init[162]), .Q(o[162]) );
  DFF \Data_Mem/memory_reg[5][3]  ( .D(\Data_Mem/n7572 ), .CLK(clk), .RST(rst), 
        .I(e_init[163]), .Q(o[163]) );
  DFF \Data_Mem/memory_reg[5][4]  ( .D(\Data_Mem/n7573 ), .CLK(clk), .RST(rst), 
        .I(e_init[164]), .Q(o[164]) );
  DFF \Data_Mem/memory_reg[5][5]  ( .D(\Data_Mem/n7574 ), .CLK(clk), .RST(rst), 
        .I(e_init[165]), .Q(o[165]) );
  DFF \Data_Mem/memory_reg[5][6]  ( .D(\Data_Mem/n7575 ), .CLK(clk), .RST(rst), 
        .I(e_init[166]), .Q(o[166]) );
  DFF \Data_Mem/memory_reg[5][7]  ( .D(\Data_Mem/n7576 ), .CLK(clk), .RST(rst), 
        .I(e_init[167]), .Q(o[167]) );
  DFF \Data_Mem/memory_reg[5][8]  ( .D(\Data_Mem/n7577 ), .CLK(clk), .RST(rst), 
        .I(e_init[168]), .Q(o[168]) );
  DFF \Data_Mem/memory_reg[5][9]  ( .D(\Data_Mem/n7578 ), .CLK(clk), .RST(rst), 
        .I(e_init[169]), .Q(o[169]) );
  DFF \Data_Mem/memory_reg[5][10]  ( .D(\Data_Mem/n7579 ), .CLK(clk), .RST(rst), .I(e_init[170]), .Q(o[170]) );
  DFF \Data_Mem/memory_reg[5][11]  ( .D(\Data_Mem/n7580 ), .CLK(clk), .RST(rst), .I(e_init[171]), .Q(o[171]) );
  DFF \Data_Mem/memory_reg[5][12]  ( .D(\Data_Mem/n7581 ), .CLK(clk), .RST(rst), .I(e_init[172]), .Q(o[172]) );
  DFF \Data_Mem/memory_reg[5][13]  ( .D(\Data_Mem/n7582 ), .CLK(clk), .RST(rst), .I(e_init[173]), .Q(o[173]) );
  DFF \Data_Mem/memory_reg[5][14]  ( .D(\Data_Mem/n7583 ), .CLK(clk), .RST(rst), .I(e_init[174]), .Q(o[174]) );
  DFF \Data_Mem/memory_reg[5][15]  ( .D(\Data_Mem/n7584 ), .CLK(clk), .RST(rst), .I(e_init[175]), .Q(o[175]) );
  DFF \Data_Mem/memory_reg[5][16]  ( .D(\Data_Mem/n7585 ), .CLK(clk), .RST(rst), .I(e_init[176]), .Q(o[176]) );
  DFF \Data_Mem/memory_reg[5][17]  ( .D(\Data_Mem/n7586 ), .CLK(clk), .RST(rst), .I(e_init[177]), .Q(o[177]) );
  DFF \Data_Mem/memory_reg[5][18]  ( .D(\Data_Mem/n7587 ), .CLK(clk), .RST(rst), .I(e_init[178]), .Q(o[178]) );
  DFF \Data_Mem/memory_reg[5][19]  ( .D(\Data_Mem/n7588 ), .CLK(clk), .RST(rst), .I(e_init[179]), .Q(o[179]) );
  DFF \Data_Mem/memory_reg[5][20]  ( .D(\Data_Mem/n7589 ), .CLK(clk), .RST(rst), .I(e_init[180]), .Q(o[180]) );
  DFF \Data_Mem/memory_reg[5][21]  ( .D(\Data_Mem/n7590 ), .CLK(clk), .RST(rst), .I(e_init[181]), .Q(o[181]) );
  DFF \Data_Mem/memory_reg[5][22]  ( .D(\Data_Mem/n7591 ), .CLK(clk), .RST(rst), .I(e_init[182]), .Q(o[182]) );
  DFF \Data_Mem/memory_reg[5][23]  ( .D(\Data_Mem/n7592 ), .CLK(clk), .RST(rst), .I(e_init[183]), .Q(o[183]) );
  DFF \Data_Mem/memory_reg[5][24]  ( .D(\Data_Mem/n7593 ), .CLK(clk), .RST(rst), .I(e_init[184]), .Q(o[184]) );
  DFF \Data_Mem/memory_reg[5][25]  ( .D(\Data_Mem/n7594 ), .CLK(clk), .RST(rst), .I(e_init[185]), .Q(o[185]) );
  DFF \Data_Mem/memory_reg[5][26]  ( .D(\Data_Mem/n7595 ), .CLK(clk), .RST(rst), .I(e_init[186]), .Q(o[186]) );
  DFF \Data_Mem/memory_reg[5][27]  ( .D(\Data_Mem/n7596 ), .CLK(clk), .RST(rst), .I(e_init[187]), .Q(o[187]) );
  DFF \Data_Mem/memory_reg[5][28]  ( .D(\Data_Mem/n7597 ), .CLK(clk), .RST(rst), .I(e_init[188]), .Q(o[188]) );
  DFF \Data_Mem/memory_reg[5][29]  ( .D(\Data_Mem/n7598 ), .CLK(clk), .RST(rst), .I(e_init[189]), .Q(o[189]) );
  DFF \Data_Mem/memory_reg[5][30]  ( .D(\Data_Mem/n7599 ), .CLK(clk), .RST(rst), .I(e_init[190]), .Q(o[190]) );
  DFF \Data_Mem/memory_reg[5][31]  ( .D(\Data_Mem/n7600 ), .CLK(clk), .RST(rst), .I(e_init[191]), .Q(o[191]) );
  DFF \Data_Mem/memory_reg[4][0]  ( .D(\Data_Mem/n7601 ), .CLK(clk), .RST(rst), 
        .I(e_init[128]), .Q(o[128]) );
  DFF \Data_Mem/memory_reg[4][1]  ( .D(\Data_Mem/n7602 ), .CLK(clk), .RST(rst), 
        .I(e_init[129]), .Q(o[129]) );
  DFF \Data_Mem/memory_reg[4][2]  ( .D(\Data_Mem/n7603 ), .CLK(clk), .RST(rst), 
        .I(e_init[130]), .Q(o[130]) );
  DFF \Data_Mem/memory_reg[4][3]  ( .D(\Data_Mem/n7604 ), .CLK(clk), .RST(rst), 
        .I(e_init[131]), .Q(o[131]) );
  DFF \Data_Mem/memory_reg[4][4]  ( .D(\Data_Mem/n7605 ), .CLK(clk), .RST(rst), 
        .I(e_init[132]), .Q(o[132]) );
  DFF \Data_Mem/memory_reg[4][5]  ( .D(\Data_Mem/n7606 ), .CLK(clk), .RST(rst), 
        .I(e_init[133]), .Q(o[133]) );
  DFF \Data_Mem/memory_reg[4][6]  ( .D(\Data_Mem/n7607 ), .CLK(clk), .RST(rst), 
        .I(e_init[134]), .Q(o[134]) );
  DFF \Data_Mem/memory_reg[4][7]  ( .D(\Data_Mem/n7608 ), .CLK(clk), .RST(rst), 
        .I(e_init[135]), .Q(o[135]) );
  DFF \Data_Mem/memory_reg[4][8]  ( .D(\Data_Mem/n7609 ), .CLK(clk), .RST(rst), 
        .I(e_init[136]), .Q(o[136]) );
  DFF \Data_Mem/memory_reg[4][9]  ( .D(\Data_Mem/n7610 ), .CLK(clk), .RST(rst), 
        .I(e_init[137]), .Q(o[137]) );
  DFF \Data_Mem/memory_reg[4][10]  ( .D(\Data_Mem/n7611 ), .CLK(clk), .RST(rst), .I(e_init[138]), .Q(o[138]) );
  DFF \Data_Mem/memory_reg[4][11]  ( .D(\Data_Mem/n7612 ), .CLK(clk), .RST(rst), .I(e_init[139]), .Q(o[139]) );
  DFF \Data_Mem/memory_reg[4][12]  ( .D(\Data_Mem/n7613 ), .CLK(clk), .RST(rst), .I(e_init[140]), .Q(o[140]) );
  DFF \Data_Mem/memory_reg[4][13]  ( .D(\Data_Mem/n7614 ), .CLK(clk), .RST(rst), .I(e_init[141]), .Q(o[141]) );
  DFF \Data_Mem/memory_reg[4][14]  ( .D(\Data_Mem/n7615 ), .CLK(clk), .RST(rst), .I(e_init[142]), .Q(o[142]) );
  DFF \Data_Mem/memory_reg[4][15]  ( .D(\Data_Mem/n7616 ), .CLK(clk), .RST(rst), .I(e_init[143]), .Q(o[143]) );
  DFF \Data_Mem/memory_reg[4][16]  ( .D(\Data_Mem/n7617 ), .CLK(clk), .RST(rst), .I(e_init[144]), .Q(o[144]) );
  DFF \Data_Mem/memory_reg[4][17]  ( .D(\Data_Mem/n7618 ), .CLK(clk), .RST(rst), .I(e_init[145]), .Q(o[145]) );
  DFF \Data_Mem/memory_reg[4][18]  ( .D(\Data_Mem/n7619 ), .CLK(clk), .RST(rst), .I(e_init[146]), .Q(o[146]) );
  DFF \Data_Mem/memory_reg[4][19]  ( .D(\Data_Mem/n7620 ), .CLK(clk), .RST(rst), .I(e_init[147]), .Q(o[147]) );
  DFF \Data_Mem/memory_reg[4][20]  ( .D(\Data_Mem/n7621 ), .CLK(clk), .RST(rst), .I(e_init[148]), .Q(o[148]) );
  DFF \Data_Mem/memory_reg[4][21]  ( .D(\Data_Mem/n7622 ), .CLK(clk), .RST(rst), .I(e_init[149]), .Q(o[149]) );
  DFF \Data_Mem/memory_reg[4][22]  ( .D(\Data_Mem/n7623 ), .CLK(clk), .RST(rst), .I(e_init[150]), .Q(o[150]) );
  DFF \Data_Mem/memory_reg[4][23]  ( .D(\Data_Mem/n7624 ), .CLK(clk), .RST(rst), .I(e_init[151]), .Q(o[151]) );
  DFF \Data_Mem/memory_reg[4][24]  ( .D(\Data_Mem/n7625 ), .CLK(clk), .RST(rst), .I(e_init[152]), .Q(o[152]) );
  DFF \Data_Mem/memory_reg[4][25]  ( .D(\Data_Mem/n7626 ), .CLK(clk), .RST(rst), .I(e_init[153]), .Q(o[153]) );
  DFF \Data_Mem/memory_reg[4][26]  ( .D(\Data_Mem/n7627 ), .CLK(clk), .RST(rst), .I(e_init[154]), .Q(o[154]) );
  DFF \Data_Mem/memory_reg[4][27]  ( .D(\Data_Mem/n7628 ), .CLK(clk), .RST(rst), .I(e_init[155]), .Q(o[155]) );
  DFF \Data_Mem/memory_reg[4][28]  ( .D(\Data_Mem/n7629 ), .CLK(clk), .RST(rst), .I(e_init[156]), .Q(o[156]) );
  DFF \Data_Mem/memory_reg[4][29]  ( .D(\Data_Mem/n7630 ), .CLK(clk), .RST(rst), .I(e_init[157]), .Q(o[157]) );
  DFF \Data_Mem/memory_reg[4][30]  ( .D(\Data_Mem/n7631 ), .CLK(clk), .RST(rst), .I(e_init[158]), .Q(o[158]) );
  DFF \Data_Mem/memory_reg[4][31]  ( .D(\Data_Mem/n7632 ), .CLK(clk), .RST(rst), .I(e_init[159]), .Q(o[159]) );
  DFF \Data_Mem/memory_reg[3][0]  ( .D(\Data_Mem/n7633 ), .CLK(clk), .RST(rst), 
        .I(e_init[96]), .Q(o[96]) );
  DFF \Data_Mem/memory_reg[3][1]  ( .D(\Data_Mem/n7634 ), .CLK(clk), .RST(rst), 
        .I(e_init[97]), .Q(o[97]) );
  DFF \Data_Mem/memory_reg[3][2]  ( .D(\Data_Mem/n7635 ), .CLK(clk), .RST(rst), 
        .I(e_init[98]), .Q(o[98]) );
  DFF \Data_Mem/memory_reg[3][3]  ( .D(\Data_Mem/n7636 ), .CLK(clk), .RST(rst), 
        .I(e_init[99]), .Q(o[99]) );
  DFF \Data_Mem/memory_reg[3][4]  ( .D(\Data_Mem/n7637 ), .CLK(clk), .RST(rst), 
        .I(e_init[100]), .Q(o[100]) );
  DFF \Data_Mem/memory_reg[3][5]  ( .D(\Data_Mem/n7638 ), .CLK(clk), .RST(rst), 
        .I(e_init[101]), .Q(o[101]) );
  DFF \Data_Mem/memory_reg[3][6]  ( .D(\Data_Mem/n7639 ), .CLK(clk), .RST(rst), 
        .I(e_init[102]), .Q(o[102]) );
  DFF \Data_Mem/memory_reg[3][7]  ( .D(\Data_Mem/n7640 ), .CLK(clk), .RST(rst), 
        .I(e_init[103]), .Q(o[103]) );
  DFF \Data_Mem/memory_reg[3][8]  ( .D(\Data_Mem/n7641 ), .CLK(clk), .RST(rst), 
        .I(e_init[104]), .Q(o[104]) );
  DFF \Data_Mem/memory_reg[3][9]  ( .D(\Data_Mem/n7642 ), .CLK(clk), .RST(rst), 
        .I(e_init[105]), .Q(o[105]) );
  DFF \Data_Mem/memory_reg[3][10]  ( .D(\Data_Mem/n7643 ), .CLK(clk), .RST(rst), .I(e_init[106]), .Q(o[106]) );
  DFF \Data_Mem/memory_reg[3][11]  ( .D(\Data_Mem/n7644 ), .CLK(clk), .RST(rst), .I(e_init[107]), .Q(o[107]) );
  DFF \Data_Mem/memory_reg[3][12]  ( .D(\Data_Mem/n7645 ), .CLK(clk), .RST(rst), .I(e_init[108]), .Q(o[108]) );
  DFF \Data_Mem/memory_reg[3][13]  ( .D(\Data_Mem/n7646 ), .CLK(clk), .RST(rst), .I(e_init[109]), .Q(o[109]) );
  DFF \Data_Mem/memory_reg[3][14]  ( .D(\Data_Mem/n7647 ), .CLK(clk), .RST(rst), .I(e_init[110]), .Q(o[110]) );
  DFF \Data_Mem/memory_reg[3][15]  ( .D(\Data_Mem/n7648 ), .CLK(clk), .RST(rst), .I(e_init[111]), .Q(o[111]) );
  DFF \Data_Mem/memory_reg[3][16]  ( .D(\Data_Mem/n7649 ), .CLK(clk), .RST(rst), .I(e_init[112]), .Q(o[112]) );
  DFF \Data_Mem/memory_reg[3][17]  ( .D(\Data_Mem/n7650 ), .CLK(clk), .RST(rst), .I(e_init[113]), .Q(o[113]) );
  DFF \Data_Mem/memory_reg[3][18]  ( .D(\Data_Mem/n7651 ), .CLK(clk), .RST(rst), .I(e_init[114]), .Q(o[114]) );
  DFF \Data_Mem/memory_reg[3][19]  ( .D(\Data_Mem/n7652 ), .CLK(clk), .RST(rst), .I(e_init[115]), .Q(o[115]) );
  DFF \Data_Mem/memory_reg[3][20]  ( .D(\Data_Mem/n7653 ), .CLK(clk), .RST(rst), .I(e_init[116]), .Q(o[116]) );
  DFF \Data_Mem/memory_reg[3][21]  ( .D(\Data_Mem/n7654 ), .CLK(clk), .RST(rst), .I(e_init[117]), .Q(o[117]) );
  DFF \Data_Mem/memory_reg[3][22]  ( .D(\Data_Mem/n7655 ), .CLK(clk), .RST(rst), .I(e_init[118]), .Q(o[118]) );
  DFF \Data_Mem/memory_reg[3][23]  ( .D(\Data_Mem/n7656 ), .CLK(clk), .RST(rst), .I(e_init[119]), .Q(o[119]) );
  DFF \Data_Mem/memory_reg[3][24]  ( .D(\Data_Mem/n7657 ), .CLK(clk), .RST(rst), .I(e_init[120]), .Q(o[120]) );
  DFF \Data_Mem/memory_reg[3][25]  ( .D(\Data_Mem/n7658 ), .CLK(clk), .RST(rst), .I(e_init[121]), .Q(o[121]) );
  DFF \Data_Mem/memory_reg[3][26]  ( .D(\Data_Mem/n7659 ), .CLK(clk), .RST(rst), .I(e_init[122]), .Q(o[122]) );
  DFF \Data_Mem/memory_reg[3][27]  ( .D(\Data_Mem/n7660 ), .CLK(clk), .RST(rst), .I(e_init[123]), .Q(o[123]) );
  DFF \Data_Mem/memory_reg[3][28]  ( .D(\Data_Mem/n7661 ), .CLK(clk), .RST(rst), .I(e_init[124]), .Q(o[124]) );
  DFF \Data_Mem/memory_reg[3][29]  ( .D(\Data_Mem/n7662 ), .CLK(clk), .RST(rst), .I(e_init[125]), .Q(o[125]) );
  DFF \Data_Mem/memory_reg[3][30]  ( .D(\Data_Mem/n7663 ), .CLK(clk), .RST(rst), .I(e_init[126]), .Q(o[126]) );
  DFF \Data_Mem/memory_reg[3][31]  ( .D(\Data_Mem/n7664 ), .CLK(clk), .RST(rst), .I(e_init[127]), .Q(o[127]) );
  DFF \Data_Mem/memory_reg[2][0]  ( .D(\Data_Mem/n7665 ), .CLK(clk), .RST(rst), 
        .I(e_init[64]), .Q(o[64]) );
  DFF \Data_Mem/memory_reg[2][1]  ( .D(\Data_Mem/n7666 ), .CLK(clk), .RST(rst), 
        .I(e_init[65]), .Q(o[65]) );
  DFF \Data_Mem/memory_reg[2][2]  ( .D(\Data_Mem/n7667 ), .CLK(clk), .RST(rst), 
        .I(e_init[66]), .Q(o[66]) );
  DFF \Data_Mem/memory_reg[2][3]  ( .D(\Data_Mem/n7668 ), .CLK(clk), .RST(rst), 
        .I(e_init[67]), .Q(o[67]) );
  DFF \Data_Mem/memory_reg[2][4]  ( .D(\Data_Mem/n7669 ), .CLK(clk), .RST(rst), 
        .I(e_init[68]), .Q(o[68]) );
  DFF \Data_Mem/memory_reg[2][5]  ( .D(\Data_Mem/n7670 ), .CLK(clk), .RST(rst), 
        .I(e_init[69]), .Q(o[69]) );
  DFF \Data_Mem/memory_reg[2][6]  ( .D(\Data_Mem/n7671 ), .CLK(clk), .RST(rst), 
        .I(e_init[70]), .Q(o[70]) );
  DFF \Data_Mem/memory_reg[2][7]  ( .D(\Data_Mem/n7672 ), .CLK(clk), .RST(rst), 
        .I(e_init[71]), .Q(o[71]) );
  DFF \Data_Mem/memory_reg[2][8]  ( .D(\Data_Mem/n7673 ), .CLK(clk), .RST(rst), 
        .I(e_init[72]), .Q(o[72]) );
  DFF \Data_Mem/memory_reg[2][9]  ( .D(\Data_Mem/n7674 ), .CLK(clk), .RST(rst), 
        .I(e_init[73]), .Q(o[73]) );
  DFF \Data_Mem/memory_reg[2][10]  ( .D(\Data_Mem/n7675 ), .CLK(clk), .RST(rst), .I(e_init[74]), .Q(o[74]) );
  DFF \Data_Mem/memory_reg[2][11]  ( .D(\Data_Mem/n7676 ), .CLK(clk), .RST(rst), .I(e_init[75]), .Q(o[75]) );
  DFF \Data_Mem/memory_reg[2][12]  ( .D(\Data_Mem/n7677 ), .CLK(clk), .RST(rst), .I(e_init[76]), .Q(o[76]) );
  DFF \Data_Mem/memory_reg[2][13]  ( .D(\Data_Mem/n7678 ), .CLK(clk), .RST(rst), .I(e_init[77]), .Q(o[77]) );
  DFF \Data_Mem/memory_reg[2][14]  ( .D(\Data_Mem/n7679 ), .CLK(clk), .RST(rst), .I(e_init[78]), .Q(o[78]) );
  DFF \Data_Mem/memory_reg[2][15]  ( .D(\Data_Mem/n7680 ), .CLK(clk), .RST(rst), .I(e_init[79]), .Q(o[79]) );
  DFF \Data_Mem/memory_reg[2][16]  ( .D(\Data_Mem/n7681 ), .CLK(clk), .RST(rst), .I(e_init[80]), .Q(o[80]) );
  DFF \Data_Mem/memory_reg[2][17]  ( .D(\Data_Mem/n7682 ), .CLK(clk), .RST(rst), .I(e_init[81]), .Q(o[81]) );
  DFF \Data_Mem/memory_reg[2][18]  ( .D(\Data_Mem/n7683 ), .CLK(clk), .RST(rst), .I(e_init[82]), .Q(o[82]) );
  DFF \Data_Mem/memory_reg[2][19]  ( .D(\Data_Mem/n7684 ), .CLK(clk), .RST(rst), .I(e_init[83]), .Q(o[83]) );
  DFF \Data_Mem/memory_reg[2][20]  ( .D(\Data_Mem/n7685 ), .CLK(clk), .RST(rst), .I(e_init[84]), .Q(o[84]) );
  DFF \Data_Mem/memory_reg[2][21]  ( .D(\Data_Mem/n7686 ), .CLK(clk), .RST(rst), .I(e_init[85]), .Q(o[85]) );
  DFF \Data_Mem/memory_reg[2][22]  ( .D(\Data_Mem/n7687 ), .CLK(clk), .RST(rst), .I(e_init[86]), .Q(o[86]) );
  DFF \Data_Mem/memory_reg[2][23]  ( .D(\Data_Mem/n7688 ), .CLK(clk), .RST(rst), .I(e_init[87]), .Q(o[87]) );
  DFF \Data_Mem/memory_reg[2][24]  ( .D(\Data_Mem/n7689 ), .CLK(clk), .RST(rst), .I(e_init[88]), .Q(o[88]) );
  DFF \Data_Mem/memory_reg[2][25]  ( .D(\Data_Mem/n7690 ), .CLK(clk), .RST(rst), .I(e_init[89]), .Q(o[89]) );
  DFF \Data_Mem/memory_reg[2][26]  ( .D(\Data_Mem/n7691 ), .CLK(clk), .RST(rst), .I(e_init[90]), .Q(o[90]) );
  DFF \Data_Mem/memory_reg[2][27]  ( .D(\Data_Mem/n7692 ), .CLK(clk), .RST(rst), .I(e_init[91]), .Q(o[91]) );
  DFF \Data_Mem/memory_reg[2][28]  ( .D(\Data_Mem/n7693 ), .CLK(clk), .RST(rst), .I(e_init[92]), .Q(o[92]) );
  DFF \Data_Mem/memory_reg[2][29]  ( .D(\Data_Mem/n7694 ), .CLK(clk), .RST(rst), .I(e_init[93]), .Q(o[93]) );
  DFF \Data_Mem/memory_reg[2][30]  ( .D(\Data_Mem/n7695 ), .CLK(clk), .RST(rst), .I(e_init[94]), .Q(o[94]) );
  DFF \Data_Mem/memory_reg[2][31]  ( .D(\Data_Mem/n7696 ), .CLK(clk), .RST(rst), .I(e_init[95]), .Q(o[95]) );
  DFF \Data_Mem/memory_reg[1][0]  ( .D(\Data_Mem/n7697 ), .CLK(clk), .RST(rst), 
        .I(e_init[32]), .Q(o[32]) );
  DFF \Data_Mem/memory_reg[1][1]  ( .D(\Data_Mem/n7698 ), .CLK(clk), .RST(rst), 
        .I(e_init[33]), .Q(o[33]) );
  DFF \Data_Mem/memory_reg[1][2]  ( .D(\Data_Mem/n7699 ), .CLK(clk), .RST(rst), 
        .I(e_init[34]), .Q(o[34]) );
  DFF \Data_Mem/memory_reg[1][3]  ( .D(\Data_Mem/n7700 ), .CLK(clk), .RST(rst), 
        .I(e_init[35]), .Q(o[35]) );
  DFF \Data_Mem/memory_reg[1][4]  ( .D(\Data_Mem/n7701 ), .CLK(clk), .RST(rst), 
        .I(e_init[36]), .Q(o[36]) );
  DFF \Data_Mem/memory_reg[1][5]  ( .D(\Data_Mem/n7702 ), .CLK(clk), .RST(rst), 
        .I(e_init[37]), .Q(o[37]) );
  DFF \Data_Mem/memory_reg[1][6]  ( .D(\Data_Mem/n7703 ), .CLK(clk), .RST(rst), 
        .I(e_init[38]), .Q(o[38]) );
  DFF \Data_Mem/memory_reg[1][7]  ( .D(\Data_Mem/n7704 ), .CLK(clk), .RST(rst), 
        .I(e_init[39]), .Q(o[39]) );
  DFF \Data_Mem/memory_reg[1][8]  ( .D(\Data_Mem/n7705 ), .CLK(clk), .RST(rst), 
        .I(e_init[40]), .Q(o[40]) );
  DFF \Data_Mem/memory_reg[1][9]  ( .D(\Data_Mem/n7706 ), .CLK(clk), .RST(rst), 
        .I(e_init[41]), .Q(o[41]) );
  DFF \Data_Mem/memory_reg[1][10]  ( .D(\Data_Mem/n7707 ), .CLK(clk), .RST(rst), .I(e_init[42]), .Q(o[42]) );
  DFF \Data_Mem/memory_reg[1][11]  ( .D(\Data_Mem/n7708 ), .CLK(clk), .RST(rst), .I(e_init[43]), .Q(o[43]) );
  DFF \Data_Mem/memory_reg[1][12]  ( .D(\Data_Mem/n7709 ), .CLK(clk), .RST(rst), .I(e_init[44]), .Q(o[44]) );
  DFF \Data_Mem/memory_reg[1][13]  ( .D(\Data_Mem/n7710 ), .CLK(clk), .RST(rst), .I(e_init[45]), .Q(o[45]) );
  DFF \Data_Mem/memory_reg[1][14]  ( .D(\Data_Mem/n7711 ), .CLK(clk), .RST(rst), .I(e_init[46]), .Q(o[46]) );
  DFF \Data_Mem/memory_reg[1][15]  ( .D(\Data_Mem/n7712 ), .CLK(clk), .RST(rst), .I(e_init[47]), .Q(o[47]) );
  DFF \Data_Mem/memory_reg[1][16]  ( .D(\Data_Mem/n7713 ), .CLK(clk), .RST(rst), .I(e_init[48]), .Q(o[48]) );
  DFF \Data_Mem/memory_reg[1][17]  ( .D(\Data_Mem/n7714 ), .CLK(clk), .RST(rst), .I(e_init[49]), .Q(o[49]) );
  DFF \Data_Mem/memory_reg[1][18]  ( .D(\Data_Mem/n7715 ), .CLK(clk), .RST(rst), .I(e_init[50]), .Q(o[50]) );
  DFF \Data_Mem/memory_reg[1][19]  ( .D(\Data_Mem/n7716 ), .CLK(clk), .RST(rst), .I(e_init[51]), .Q(o[51]) );
  DFF \Data_Mem/memory_reg[1][20]  ( .D(\Data_Mem/n7717 ), .CLK(clk), .RST(rst), .I(e_init[52]), .Q(o[52]) );
  DFF \Data_Mem/memory_reg[1][21]  ( .D(\Data_Mem/n7718 ), .CLK(clk), .RST(rst), .I(e_init[53]), .Q(o[53]) );
  DFF \Data_Mem/memory_reg[1][22]  ( .D(\Data_Mem/n7719 ), .CLK(clk), .RST(rst), .I(e_init[54]), .Q(o[54]) );
  DFF \Data_Mem/memory_reg[1][23]  ( .D(\Data_Mem/n7720 ), .CLK(clk), .RST(rst), .I(e_init[55]), .Q(o[55]) );
  DFF \Data_Mem/memory_reg[1][24]  ( .D(\Data_Mem/n7721 ), .CLK(clk), .RST(rst), .I(e_init[56]), .Q(o[56]) );
  DFF \Data_Mem/memory_reg[1][25]  ( .D(\Data_Mem/n7722 ), .CLK(clk), .RST(rst), .I(e_init[57]), .Q(o[57]) );
  DFF \Data_Mem/memory_reg[1][26]  ( .D(\Data_Mem/n7723 ), .CLK(clk), .RST(rst), .I(e_init[58]), .Q(o[58]) );
  DFF \Data_Mem/memory_reg[1][27]  ( .D(\Data_Mem/n7724 ), .CLK(clk), .RST(rst), .I(e_init[59]), .Q(o[59]) );
  DFF \Data_Mem/memory_reg[1][28]  ( .D(\Data_Mem/n7725 ), .CLK(clk), .RST(rst), .I(e_init[60]), .Q(o[60]) );
  DFF \Data_Mem/memory_reg[1][29]  ( .D(\Data_Mem/n7726 ), .CLK(clk), .RST(rst), .I(e_init[61]), .Q(o[61]) );
  DFF \Data_Mem/memory_reg[1][30]  ( .D(\Data_Mem/n7727 ), .CLK(clk), .RST(rst), .I(e_init[62]), .Q(o[62]) );
  DFF \Data_Mem/memory_reg[1][31]  ( .D(\Data_Mem/n7728 ), .CLK(clk), .RST(rst), .I(e_init[63]), .Q(o[63]) );
  DFF \Data_Mem/memory_reg[0][0]  ( .D(\Data_Mem/n7729 ), .CLK(clk), .RST(rst), 
        .I(e_init[0]), .Q(o[0]) );
  DFF \Data_Mem/memory_reg[0][1]  ( .D(\Data_Mem/n7730 ), .CLK(clk), .RST(rst), 
        .I(e_init[1]), .Q(o[1]) );
  DFF \Data_Mem/memory_reg[0][2]  ( .D(\Data_Mem/n7731 ), .CLK(clk), .RST(rst), 
        .I(e_init[2]), .Q(o[2]) );
  DFF \Data_Mem/memory_reg[0][3]  ( .D(\Data_Mem/n7732 ), .CLK(clk), .RST(rst), 
        .I(e_init[3]), .Q(o[3]) );
  DFF \Data_Mem/memory_reg[0][4]  ( .D(\Data_Mem/n7733 ), .CLK(clk), .RST(rst), 
        .I(e_init[4]), .Q(o[4]) );
  DFF \Data_Mem/memory_reg[0][5]  ( .D(\Data_Mem/n7734 ), .CLK(clk), .RST(rst), 
        .I(e_init[5]), .Q(o[5]) );
  DFF \Data_Mem/memory_reg[0][6]  ( .D(\Data_Mem/n7735 ), .CLK(clk), .RST(rst), 
        .I(e_init[6]), .Q(o[6]) );
  DFF \Data_Mem/memory_reg[0][7]  ( .D(\Data_Mem/n7736 ), .CLK(clk), .RST(rst), 
        .I(e_init[7]), .Q(o[7]) );
  DFF \Data_Mem/memory_reg[0][8]  ( .D(\Data_Mem/n7737 ), .CLK(clk), .RST(rst), 
        .I(e_init[8]), .Q(o[8]) );
  DFF \Data_Mem/memory_reg[0][9]  ( .D(\Data_Mem/n7738 ), .CLK(clk), .RST(rst), 
        .I(e_init[9]), .Q(o[9]) );
  DFF \Data_Mem/memory_reg[0][10]  ( .D(\Data_Mem/n7739 ), .CLK(clk), .RST(rst), .I(e_init[10]), .Q(o[10]) );
  DFF \Data_Mem/memory_reg[0][11]  ( .D(\Data_Mem/n7740 ), .CLK(clk), .RST(rst), .I(e_init[11]), .Q(o[11]) );
  DFF \Data_Mem/memory_reg[0][12]  ( .D(\Data_Mem/n7741 ), .CLK(clk), .RST(rst), .I(e_init[12]), .Q(o[12]) );
  DFF \Data_Mem/memory_reg[0][13]  ( .D(\Data_Mem/n7742 ), .CLK(clk), .RST(rst), .I(e_init[13]), .Q(o[13]) );
  DFF \Data_Mem/memory_reg[0][14]  ( .D(\Data_Mem/n7743 ), .CLK(clk), .RST(rst), .I(e_init[14]), .Q(o[14]) );
  DFF \Data_Mem/memory_reg[0][15]  ( .D(\Data_Mem/n7744 ), .CLK(clk), .RST(rst), .I(e_init[15]), .Q(o[15]) );
  DFF \Data_Mem/memory_reg[0][16]  ( .D(\Data_Mem/n7745 ), .CLK(clk), .RST(rst), .I(e_init[16]), .Q(o[16]) );
  DFF \Data_Mem/memory_reg[0][17]  ( .D(\Data_Mem/n7746 ), .CLK(clk), .RST(rst), .I(e_init[17]), .Q(o[17]) );
  DFF \Data_Mem/memory_reg[0][18]  ( .D(\Data_Mem/n7747 ), .CLK(clk), .RST(rst), .I(e_init[18]), .Q(o[18]) );
  DFF \Data_Mem/memory_reg[0][19]  ( .D(\Data_Mem/n7748 ), .CLK(clk), .RST(rst), .I(e_init[19]), .Q(o[19]) );
  DFF \Data_Mem/memory_reg[0][20]  ( .D(\Data_Mem/n7749 ), .CLK(clk), .RST(rst), .I(e_init[20]), .Q(o[20]) );
  DFF \Data_Mem/memory_reg[0][21]  ( .D(\Data_Mem/n7750 ), .CLK(clk), .RST(rst), .I(e_init[21]), .Q(o[21]) );
  DFF \Data_Mem/memory_reg[0][22]  ( .D(\Data_Mem/n7751 ), .CLK(clk), .RST(rst), .I(e_init[22]), .Q(o[22]) );
  DFF \Data_Mem/memory_reg[0][23]  ( .D(\Data_Mem/n7752 ), .CLK(clk), .RST(rst), .I(e_init[23]), .Q(o[23]) );
  DFF \Data_Mem/memory_reg[0][24]  ( .D(\Data_Mem/n7753 ), .CLK(clk), .RST(rst), .I(e_init[24]), .Q(o[24]) );
  DFF \Data_Mem/memory_reg[0][25]  ( .D(\Data_Mem/n7754 ), .CLK(clk), .RST(rst), .I(e_init[25]), .Q(o[25]) );
  DFF \Data_Mem/memory_reg[0][26]  ( .D(\Data_Mem/n7755 ), .CLK(clk), .RST(rst), .I(e_init[26]), .Q(o[26]) );
  DFF \Data_Mem/memory_reg[0][27]  ( .D(\Data_Mem/n7756 ), .CLK(clk), .RST(rst), .I(e_init[27]), .Q(o[27]) );
  DFF \Data_Mem/memory_reg[0][28]  ( .D(\Data_Mem/n7757 ), .CLK(clk), .RST(rst), .I(e_init[28]), .Q(o[28]) );
  DFF \Data_Mem/memory_reg[0][29]  ( .D(\Data_Mem/n7758 ), .CLK(clk), .RST(rst), .I(e_init[29]), .Q(o[29]) );
  DFF \Data_Mem/memory_reg[0][30]  ( .D(\Data_Mem/n7759 ), .CLK(clk), .RST(rst), .I(e_init[30]), .Q(o[30]) );
  DFF \Data_Mem/memory_reg[0][31]  ( .D(\Data_Mem/n7760 ), .CLK(clk), .RST(rst), .I(e_init[31]), .Q(o[31]) );
  MUX \Reg_Bank/U6036  ( .IN0(\Reg_Bank/n5939 ), .IN1(\Reg_Bank/n5924 ), .SEL(
        rt_index[4]), .F(reg_target[31]) );
  MUX \Reg_Bank/U6035  ( .IN0(\Reg_Bank/n5938 ), .IN1(\Reg_Bank/n5931 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5939 ) );
  MUX \Reg_Bank/U6034  ( .IN0(\Reg_Bank/n5937 ), .IN1(\Reg_Bank/n5934 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5938 ) );
  MUX \Reg_Bank/U6033  ( .IN0(\Reg_Bank/n5936 ), .IN1(\Reg_Bank/n5935 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5937 ) );
  MUX \Reg_Bank/U6031  ( .IN0(\Reg_Bank/registers[2][31] ), .IN1(
        \Reg_Bank/registers[3][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5935 )
         );
  MUX \Reg_Bank/U6030  ( .IN0(\Reg_Bank/n5933 ), .IN1(\Reg_Bank/n5932 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5934 ) );
  MUX \Reg_Bank/U6029  ( .IN0(\Reg_Bank/registers[4][31] ), .IN1(
        \Reg_Bank/registers[5][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5933 )
         );
  MUX \Reg_Bank/U6028  ( .IN0(\Reg_Bank/registers[6][31] ), .IN1(
        \Reg_Bank/registers[7][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5932 )
         );
  MUX \Reg_Bank/U6027  ( .IN0(\Reg_Bank/n5930 ), .IN1(\Reg_Bank/n5927 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5931 ) );
  MUX \Reg_Bank/U6026  ( .IN0(\Reg_Bank/n5929 ), .IN1(\Reg_Bank/n5928 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5930 ) );
  MUX \Reg_Bank/U6025  ( .IN0(\Reg_Bank/registers[8][31] ), .IN1(
        \Reg_Bank/registers[9][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5929 )
         );
  MUX \Reg_Bank/U6024  ( .IN0(\Reg_Bank/registers[10][31] ), .IN1(
        \Reg_Bank/registers[11][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5928 )
         );
  MUX \Reg_Bank/U6023  ( .IN0(\Reg_Bank/n5926 ), .IN1(\Reg_Bank/n5925 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5927 ) );
  MUX \Reg_Bank/U6022  ( .IN0(\Reg_Bank/registers[12][31] ), .IN1(
        \Reg_Bank/registers[13][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5926 )
         );
  MUX \Reg_Bank/U6021  ( .IN0(\Reg_Bank/registers[14][31] ), .IN1(
        \Reg_Bank/registers[15][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5925 )
         );
  MUX \Reg_Bank/U6020  ( .IN0(\Reg_Bank/n5923 ), .IN1(\Reg_Bank/n5916 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5924 ) );
  MUX \Reg_Bank/U6019  ( .IN0(\Reg_Bank/n5922 ), .IN1(\Reg_Bank/n5919 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5923 ) );
  MUX \Reg_Bank/U6018  ( .IN0(\Reg_Bank/n5921 ), .IN1(\Reg_Bank/n5920 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5922 ) );
  MUX \Reg_Bank/U6017  ( .IN0(\Reg_Bank/registers[16][31] ), .IN1(
        \Reg_Bank/registers[17][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5921 )
         );
  MUX \Reg_Bank/U6016  ( .IN0(\Reg_Bank/registers[18][31] ), .IN1(
        \Reg_Bank/registers[19][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5920 )
         );
  MUX \Reg_Bank/U6015  ( .IN0(\Reg_Bank/n5918 ), .IN1(\Reg_Bank/n5917 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5919 ) );
  MUX \Reg_Bank/U6014  ( .IN0(\Reg_Bank/registers[20][31] ), .IN1(
        \Reg_Bank/registers[21][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5918 )
         );
  MUX \Reg_Bank/U6013  ( .IN0(\Reg_Bank/registers[22][31] ), .IN1(
        \Reg_Bank/registers[23][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5917 )
         );
  MUX \Reg_Bank/U6012  ( .IN0(\Reg_Bank/n5915 ), .IN1(\Reg_Bank/n5912 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5916 ) );
  MUX \Reg_Bank/U6011  ( .IN0(\Reg_Bank/n5914 ), .IN1(\Reg_Bank/n5913 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5915 ) );
  MUX \Reg_Bank/U6010  ( .IN0(\Reg_Bank/registers[24][31] ), .IN1(
        \Reg_Bank/registers[25][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5914 )
         );
  MUX \Reg_Bank/U6009  ( .IN0(\Reg_Bank/registers[26][31] ), .IN1(
        \Reg_Bank/registers[27][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5913 )
         );
  MUX \Reg_Bank/U6008  ( .IN0(\Reg_Bank/n5911 ), .IN1(\Reg_Bank/n5910 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5912 ) );
  MUX \Reg_Bank/U6007  ( .IN0(\Reg_Bank/registers[28][31] ), .IN1(
        \Reg_Bank/registers[29][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5911 )
         );
  MUX \Reg_Bank/U6006  ( .IN0(\Reg_Bank/registers[30][31] ), .IN1(
        \Reg_Bank/registers[31][31] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5910 )
         );
  MUX \Reg_Bank/U6005  ( .IN0(\Reg_Bank/n5909 ), .IN1(\Reg_Bank/n5894 ), .SEL(
        rt_index[4]), .F(reg_target[30]) );
  MUX \Reg_Bank/U6004  ( .IN0(\Reg_Bank/n5908 ), .IN1(\Reg_Bank/n5901 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5909 ) );
  MUX \Reg_Bank/U6003  ( .IN0(\Reg_Bank/n5907 ), .IN1(\Reg_Bank/n5904 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5908 ) );
  MUX \Reg_Bank/U6002  ( .IN0(\Reg_Bank/n5906 ), .IN1(\Reg_Bank/n5905 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5907 ) );
  MUX \Reg_Bank/U6000  ( .IN0(\Reg_Bank/registers[2][30] ), .IN1(
        \Reg_Bank/registers[3][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5905 )
         );
  MUX \Reg_Bank/U5999  ( .IN0(\Reg_Bank/n5903 ), .IN1(\Reg_Bank/n5902 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5904 ) );
  MUX \Reg_Bank/U5998  ( .IN0(\Reg_Bank/registers[4][30] ), .IN1(
        \Reg_Bank/registers[5][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5903 )
         );
  MUX \Reg_Bank/U5997  ( .IN0(\Reg_Bank/registers[6][30] ), .IN1(
        \Reg_Bank/registers[7][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5902 )
         );
  MUX \Reg_Bank/U5996  ( .IN0(\Reg_Bank/n5900 ), .IN1(\Reg_Bank/n5897 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5901 ) );
  MUX \Reg_Bank/U5995  ( .IN0(\Reg_Bank/n5899 ), .IN1(\Reg_Bank/n5898 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5900 ) );
  MUX \Reg_Bank/U5994  ( .IN0(\Reg_Bank/registers[8][30] ), .IN1(
        \Reg_Bank/registers[9][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5899 )
         );
  MUX \Reg_Bank/U5993  ( .IN0(\Reg_Bank/registers[10][30] ), .IN1(
        \Reg_Bank/registers[11][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5898 )
         );
  MUX \Reg_Bank/U5992  ( .IN0(\Reg_Bank/n5896 ), .IN1(\Reg_Bank/n5895 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5897 ) );
  MUX \Reg_Bank/U5991  ( .IN0(\Reg_Bank/registers[12][30] ), .IN1(
        \Reg_Bank/registers[13][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5896 )
         );
  MUX \Reg_Bank/U5990  ( .IN0(\Reg_Bank/registers[14][30] ), .IN1(
        \Reg_Bank/registers[15][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5895 )
         );
  MUX \Reg_Bank/U5989  ( .IN0(\Reg_Bank/n5893 ), .IN1(\Reg_Bank/n5886 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5894 ) );
  MUX \Reg_Bank/U5988  ( .IN0(\Reg_Bank/n5892 ), .IN1(\Reg_Bank/n5889 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5893 ) );
  MUX \Reg_Bank/U5987  ( .IN0(\Reg_Bank/n5891 ), .IN1(\Reg_Bank/n5890 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5892 ) );
  MUX \Reg_Bank/U5986  ( .IN0(\Reg_Bank/registers[16][30] ), .IN1(
        \Reg_Bank/registers[17][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5891 )
         );
  MUX \Reg_Bank/U5985  ( .IN0(\Reg_Bank/registers[18][30] ), .IN1(
        \Reg_Bank/registers[19][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5890 )
         );
  MUX \Reg_Bank/U5984  ( .IN0(\Reg_Bank/n5888 ), .IN1(\Reg_Bank/n5887 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5889 ) );
  MUX \Reg_Bank/U5983  ( .IN0(\Reg_Bank/registers[20][30] ), .IN1(
        \Reg_Bank/registers[21][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5888 )
         );
  MUX \Reg_Bank/U5982  ( .IN0(\Reg_Bank/registers[22][30] ), .IN1(
        \Reg_Bank/registers[23][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5887 )
         );
  MUX \Reg_Bank/U5981  ( .IN0(\Reg_Bank/n5885 ), .IN1(\Reg_Bank/n5882 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5886 ) );
  MUX \Reg_Bank/U5980  ( .IN0(\Reg_Bank/n5884 ), .IN1(\Reg_Bank/n5883 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5885 ) );
  MUX \Reg_Bank/U5979  ( .IN0(\Reg_Bank/registers[24][30] ), .IN1(
        \Reg_Bank/registers[25][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5884 )
         );
  MUX \Reg_Bank/U5978  ( .IN0(\Reg_Bank/registers[26][30] ), .IN1(
        \Reg_Bank/registers[27][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5883 )
         );
  MUX \Reg_Bank/U5977  ( .IN0(\Reg_Bank/n5881 ), .IN1(\Reg_Bank/n5880 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5882 ) );
  MUX \Reg_Bank/U5976  ( .IN0(\Reg_Bank/registers[28][30] ), .IN1(
        \Reg_Bank/registers[29][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5881 )
         );
  MUX \Reg_Bank/U5975  ( .IN0(\Reg_Bank/registers[30][30] ), .IN1(
        \Reg_Bank/registers[31][30] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5880 )
         );
  MUX \Reg_Bank/U5974  ( .IN0(\Reg_Bank/n5879 ), .IN1(\Reg_Bank/n5864 ), .SEL(
        rt_index[4]), .F(reg_target[29]) );
  MUX \Reg_Bank/U5973  ( .IN0(\Reg_Bank/n5878 ), .IN1(\Reg_Bank/n5871 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5879 ) );
  MUX \Reg_Bank/U5972  ( .IN0(\Reg_Bank/n5877 ), .IN1(\Reg_Bank/n5874 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5878 ) );
  MUX \Reg_Bank/U5971  ( .IN0(\Reg_Bank/n5876 ), .IN1(\Reg_Bank/n5875 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5877 ) );
  MUX \Reg_Bank/U5969  ( .IN0(\Reg_Bank/registers[2][29] ), .IN1(
        \Reg_Bank/registers[3][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5875 )
         );
  MUX \Reg_Bank/U5968  ( .IN0(\Reg_Bank/n5873 ), .IN1(\Reg_Bank/n5872 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5874 ) );
  MUX \Reg_Bank/U5967  ( .IN0(\Reg_Bank/registers[4][29] ), .IN1(
        \Reg_Bank/registers[5][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5873 )
         );
  MUX \Reg_Bank/U5966  ( .IN0(\Reg_Bank/registers[6][29] ), .IN1(
        \Reg_Bank/registers[7][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5872 )
         );
  MUX \Reg_Bank/U5965  ( .IN0(\Reg_Bank/n5870 ), .IN1(\Reg_Bank/n5867 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5871 ) );
  MUX \Reg_Bank/U5964  ( .IN0(\Reg_Bank/n5869 ), .IN1(\Reg_Bank/n5868 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5870 ) );
  MUX \Reg_Bank/U5963  ( .IN0(\Reg_Bank/registers[8][29] ), .IN1(
        \Reg_Bank/registers[9][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5869 )
         );
  MUX \Reg_Bank/U5962  ( .IN0(\Reg_Bank/registers[10][29] ), .IN1(
        \Reg_Bank/registers[11][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5868 )
         );
  MUX \Reg_Bank/U5961  ( .IN0(\Reg_Bank/n5866 ), .IN1(\Reg_Bank/n5865 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5867 ) );
  MUX \Reg_Bank/U5960  ( .IN0(\Reg_Bank/registers[12][29] ), .IN1(
        \Reg_Bank/registers[13][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5866 )
         );
  MUX \Reg_Bank/U5959  ( .IN0(\Reg_Bank/registers[14][29] ), .IN1(
        \Reg_Bank/registers[15][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5865 )
         );
  MUX \Reg_Bank/U5958  ( .IN0(\Reg_Bank/n5863 ), .IN1(\Reg_Bank/n5856 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5864 ) );
  MUX \Reg_Bank/U5957  ( .IN0(\Reg_Bank/n5862 ), .IN1(\Reg_Bank/n5859 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5863 ) );
  MUX \Reg_Bank/U5956  ( .IN0(\Reg_Bank/n5861 ), .IN1(\Reg_Bank/n5860 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5862 ) );
  MUX \Reg_Bank/U5955  ( .IN0(\Reg_Bank/registers[16][29] ), .IN1(
        \Reg_Bank/registers[17][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5861 )
         );
  MUX \Reg_Bank/U5954  ( .IN0(\Reg_Bank/registers[18][29] ), .IN1(
        \Reg_Bank/registers[19][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5860 )
         );
  MUX \Reg_Bank/U5953  ( .IN0(\Reg_Bank/n5858 ), .IN1(\Reg_Bank/n5857 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5859 ) );
  MUX \Reg_Bank/U5952  ( .IN0(\Reg_Bank/registers[20][29] ), .IN1(
        \Reg_Bank/registers[21][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5858 )
         );
  MUX \Reg_Bank/U5951  ( .IN0(\Reg_Bank/registers[22][29] ), .IN1(
        \Reg_Bank/registers[23][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5857 )
         );
  MUX \Reg_Bank/U5950  ( .IN0(\Reg_Bank/n5855 ), .IN1(\Reg_Bank/n5852 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5856 ) );
  MUX \Reg_Bank/U5949  ( .IN0(\Reg_Bank/n5854 ), .IN1(\Reg_Bank/n5853 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5855 ) );
  MUX \Reg_Bank/U5948  ( .IN0(\Reg_Bank/registers[24][29] ), .IN1(
        \Reg_Bank/registers[25][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5854 )
         );
  MUX \Reg_Bank/U5947  ( .IN0(\Reg_Bank/registers[26][29] ), .IN1(
        \Reg_Bank/registers[27][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5853 )
         );
  MUX \Reg_Bank/U5946  ( .IN0(\Reg_Bank/n5851 ), .IN1(\Reg_Bank/n5850 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5852 ) );
  MUX \Reg_Bank/U5945  ( .IN0(\Reg_Bank/registers[28][29] ), .IN1(
        \Reg_Bank/registers[29][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5851 )
         );
  MUX \Reg_Bank/U5944  ( .IN0(\Reg_Bank/registers[30][29] ), .IN1(
        \Reg_Bank/registers[31][29] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5850 )
         );
  MUX \Reg_Bank/U5943  ( .IN0(\Reg_Bank/n5849 ), .IN1(\Reg_Bank/n5834 ), .SEL(
        rt_index[4]), .F(reg_target[28]) );
  MUX \Reg_Bank/U5942  ( .IN0(\Reg_Bank/n5848 ), .IN1(\Reg_Bank/n5841 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5849 ) );
  MUX \Reg_Bank/U5941  ( .IN0(\Reg_Bank/n5847 ), .IN1(\Reg_Bank/n5844 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5848 ) );
  MUX \Reg_Bank/U5940  ( .IN0(\Reg_Bank/n5846 ), .IN1(\Reg_Bank/n5845 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5847 ) );
  MUX \Reg_Bank/U5938  ( .IN0(\Reg_Bank/registers[2][28] ), .IN1(
        \Reg_Bank/registers[3][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5845 )
         );
  MUX \Reg_Bank/U5937  ( .IN0(\Reg_Bank/n5843 ), .IN1(\Reg_Bank/n5842 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5844 ) );
  MUX \Reg_Bank/U5936  ( .IN0(\Reg_Bank/registers[4][28] ), .IN1(
        \Reg_Bank/registers[5][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5843 )
         );
  MUX \Reg_Bank/U5935  ( .IN0(\Reg_Bank/registers[6][28] ), .IN1(
        \Reg_Bank/registers[7][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5842 )
         );
  MUX \Reg_Bank/U5934  ( .IN0(\Reg_Bank/n5840 ), .IN1(\Reg_Bank/n5837 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5841 ) );
  MUX \Reg_Bank/U5933  ( .IN0(\Reg_Bank/n5839 ), .IN1(\Reg_Bank/n5838 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5840 ) );
  MUX \Reg_Bank/U5932  ( .IN0(\Reg_Bank/registers[8][28] ), .IN1(
        \Reg_Bank/registers[9][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5839 )
         );
  MUX \Reg_Bank/U5931  ( .IN0(\Reg_Bank/registers[10][28] ), .IN1(
        \Reg_Bank/registers[11][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5838 )
         );
  MUX \Reg_Bank/U5930  ( .IN0(\Reg_Bank/n5836 ), .IN1(\Reg_Bank/n5835 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5837 ) );
  MUX \Reg_Bank/U5929  ( .IN0(\Reg_Bank/registers[12][28] ), .IN1(
        \Reg_Bank/registers[13][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5836 )
         );
  MUX \Reg_Bank/U5928  ( .IN0(\Reg_Bank/registers[14][28] ), .IN1(
        \Reg_Bank/registers[15][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5835 )
         );
  MUX \Reg_Bank/U5927  ( .IN0(\Reg_Bank/n5833 ), .IN1(\Reg_Bank/n5826 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5834 ) );
  MUX \Reg_Bank/U5926  ( .IN0(\Reg_Bank/n5832 ), .IN1(\Reg_Bank/n5829 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5833 ) );
  MUX \Reg_Bank/U5925  ( .IN0(\Reg_Bank/n5831 ), .IN1(\Reg_Bank/n5830 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5832 ) );
  MUX \Reg_Bank/U5924  ( .IN0(\Reg_Bank/registers[16][28] ), .IN1(
        \Reg_Bank/registers[17][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5831 )
         );
  MUX \Reg_Bank/U5923  ( .IN0(\Reg_Bank/registers[18][28] ), .IN1(
        \Reg_Bank/registers[19][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5830 )
         );
  MUX \Reg_Bank/U5922  ( .IN0(\Reg_Bank/n5828 ), .IN1(\Reg_Bank/n5827 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5829 ) );
  MUX \Reg_Bank/U5921  ( .IN0(\Reg_Bank/registers[20][28] ), .IN1(
        \Reg_Bank/registers[21][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5828 )
         );
  MUX \Reg_Bank/U5920  ( .IN0(\Reg_Bank/registers[22][28] ), .IN1(
        \Reg_Bank/registers[23][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5827 )
         );
  MUX \Reg_Bank/U5919  ( .IN0(\Reg_Bank/n5825 ), .IN1(\Reg_Bank/n5822 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5826 ) );
  MUX \Reg_Bank/U5918  ( .IN0(\Reg_Bank/n5824 ), .IN1(\Reg_Bank/n5823 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5825 ) );
  MUX \Reg_Bank/U5917  ( .IN0(\Reg_Bank/registers[24][28] ), .IN1(
        \Reg_Bank/registers[25][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5824 )
         );
  MUX \Reg_Bank/U5916  ( .IN0(\Reg_Bank/registers[26][28] ), .IN1(
        \Reg_Bank/registers[27][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5823 )
         );
  MUX \Reg_Bank/U5915  ( .IN0(\Reg_Bank/n5821 ), .IN1(\Reg_Bank/n5820 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5822 ) );
  MUX \Reg_Bank/U5914  ( .IN0(\Reg_Bank/registers[28][28] ), .IN1(
        \Reg_Bank/registers[29][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5821 )
         );
  MUX \Reg_Bank/U5913  ( .IN0(\Reg_Bank/registers[30][28] ), .IN1(
        \Reg_Bank/registers[31][28] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5820 )
         );
  MUX \Reg_Bank/U5912  ( .IN0(\Reg_Bank/n5819 ), .IN1(\Reg_Bank/n5804 ), .SEL(
        rt_index[4]), .F(reg_target[27]) );
  MUX \Reg_Bank/U5911  ( .IN0(\Reg_Bank/n5818 ), .IN1(\Reg_Bank/n5811 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5819 ) );
  MUX \Reg_Bank/U5910  ( .IN0(\Reg_Bank/n5817 ), .IN1(\Reg_Bank/n5814 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5818 ) );
  MUX \Reg_Bank/U5909  ( .IN0(\Reg_Bank/n5816 ), .IN1(\Reg_Bank/n5815 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5817 ) );
  MUX \Reg_Bank/U5907  ( .IN0(\Reg_Bank/registers[2][27] ), .IN1(
        \Reg_Bank/registers[3][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5815 )
         );
  MUX \Reg_Bank/U5906  ( .IN0(\Reg_Bank/n5813 ), .IN1(\Reg_Bank/n5812 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5814 ) );
  MUX \Reg_Bank/U5905  ( .IN0(\Reg_Bank/registers[4][27] ), .IN1(
        \Reg_Bank/registers[5][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5813 )
         );
  MUX \Reg_Bank/U5904  ( .IN0(\Reg_Bank/registers[6][27] ), .IN1(
        \Reg_Bank/registers[7][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5812 )
         );
  MUX \Reg_Bank/U5903  ( .IN0(\Reg_Bank/n5810 ), .IN1(\Reg_Bank/n5807 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5811 ) );
  MUX \Reg_Bank/U5902  ( .IN0(\Reg_Bank/n5809 ), .IN1(\Reg_Bank/n5808 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5810 ) );
  MUX \Reg_Bank/U5901  ( .IN0(\Reg_Bank/registers[8][27] ), .IN1(
        \Reg_Bank/registers[9][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5809 )
         );
  MUX \Reg_Bank/U5900  ( .IN0(\Reg_Bank/registers[10][27] ), .IN1(
        \Reg_Bank/registers[11][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5808 )
         );
  MUX \Reg_Bank/U5899  ( .IN0(\Reg_Bank/n5806 ), .IN1(\Reg_Bank/n5805 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5807 ) );
  MUX \Reg_Bank/U5898  ( .IN0(\Reg_Bank/registers[12][27] ), .IN1(
        \Reg_Bank/registers[13][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5806 )
         );
  MUX \Reg_Bank/U5897  ( .IN0(\Reg_Bank/registers[14][27] ), .IN1(
        \Reg_Bank/registers[15][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5805 )
         );
  MUX \Reg_Bank/U5896  ( .IN0(\Reg_Bank/n5803 ), .IN1(\Reg_Bank/n5796 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5804 ) );
  MUX \Reg_Bank/U5895  ( .IN0(\Reg_Bank/n5802 ), .IN1(\Reg_Bank/n5799 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5803 ) );
  MUX \Reg_Bank/U5894  ( .IN0(\Reg_Bank/n5801 ), .IN1(\Reg_Bank/n5800 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5802 ) );
  MUX \Reg_Bank/U5893  ( .IN0(\Reg_Bank/registers[16][27] ), .IN1(
        \Reg_Bank/registers[17][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5801 )
         );
  MUX \Reg_Bank/U5892  ( .IN0(\Reg_Bank/registers[18][27] ), .IN1(
        \Reg_Bank/registers[19][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5800 )
         );
  MUX \Reg_Bank/U5891  ( .IN0(\Reg_Bank/n5798 ), .IN1(\Reg_Bank/n5797 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5799 ) );
  MUX \Reg_Bank/U5890  ( .IN0(\Reg_Bank/registers[20][27] ), .IN1(
        \Reg_Bank/registers[21][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5798 )
         );
  MUX \Reg_Bank/U5889  ( .IN0(\Reg_Bank/registers[22][27] ), .IN1(
        \Reg_Bank/registers[23][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5797 )
         );
  MUX \Reg_Bank/U5888  ( .IN0(\Reg_Bank/n5795 ), .IN1(\Reg_Bank/n5792 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5796 ) );
  MUX \Reg_Bank/U5887  ( .IN0(\Reg_Bank/n5794 ), .IN1(\Reg_Bank/n5793 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5795 ) );
  MUX \Reg_Bank/U5886  ( .IN0(\Reg_Bank/registers[24][27] ), .IN1(
        \Reg_Bank/registers[25][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5794 )
         );
  MUX \Reg_Bank/U5885  ( .IN0(\Reg_Bank/registers[26][27] ), .IN1(
        \Reg_Bank/registers[27][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5793 )
         );
  MUX \Reg_Bank/U5884  ( .IN0(\Reg_Bank/n5791 ), .IN1(\Reg_Bank/n5790 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5792 ) );
  MUX \Reg_Bank/U5883  ( .IN0(\Reg_Bank/registers[28][27] ), .IN1(
        \Reg_Bank/registers[29][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5791 )
         );
  MUX \Reg_Bank/U5882  ( .IN0(\Reg_Bank/registers[30][27] ), .IN1(
        \Reg_Bank/registers[31][27] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5790 )
         );
  MUX \Reg_Bank/U5881  ( .IN0(\Reg_Bank/n5789 ), .IN1(\Reg_Bank/n5774 ), .SEL(
        rt_index[4]), .F(reg_target[26]) );
  MUX \Reg_Bank/U5880  ( .IN0(\Reg_Bank/n5788 ), .IN1(\Reg_Bank/n5781 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5789 ) );
  MUX \Reg_Bank/U5879  ( .IN0(\Reg_Bank/n5787 ), .IN1(\Reg_Bank/n5784 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5788 ) );
  MUX \Reg_Bank/U5878  ( .IN0(\Reg_Bank/n5786 ), .IN1(\Reg_Bank/n5785 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5787 ) );
  MUX \Reg_Bank/U5876  ( .IN0(\Reg_Bank/registers[2][26] ), .IN1(
        \Reg_Bank/registers[3][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5785 )
         );
  MUX \Reg_Bank/U5875  ( .IN0(\Reg_Bank/n5783 ), .IN1(\Reg_Bank/n5782 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5784 ) );
  MUX \Reg_Bank/U5874  ( .IN0(\Reg_Bank/registers[4][26] ), .IN1(
        \Reg_Bank/registers[5][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5783 )
         );
  MUX \Reg_Bank/U5873  ( .IN0(\Reg_Bank/registers[6][26] ), .IN1(
        \Reg_Bank/registers[7][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5782 )
         );
  MUX \Reg_Bank/U5872  ( .IN0(\Reg_Bank/n5780 ), .IN1(\Reg_Bank/n5777 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5781 ) );
  MUX \Reg_Bank/U5871  ( .IN0(\Reg_Bank/n5779 ), .IN1(\Reg_Bank/n5778 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5780 ) );
  MUX \Reg_Bank/U5870  ( .IN0(\Reg_Bank/registers[8][26] ), .IN1(
        \Reg_Bank/registers[9][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5779 )
         );
  MUX \Reg_Bank/U5869  ( .IN0(\Reg_Bank/registers[10][26] ), .IN1(
        \Reg_Bank/registers[11][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5778 )
         );
  MUX \Reg_Bank/U5868  ( .IN0(\Reg_Bank/n5776 ), .IN1(\Reg_Bank/n5775 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5777 ) );
  MUX \Reg_Bank/U5867  ( .IN0(\Reg_Bank/registers[12][26] ), .IN1(
        \Reg_Bank/registers[13][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5776 )
         );
  MUX \Reg_Bank/U5866  ( .IN0(\Reg_Bank/registers[14][26] ), .IN1(
        \Reg_Bank/registers[15][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5775 )
         );
  MUX \Reg_Bank/U5865  ( .IN0(\Reg_Bank/n5773 ), .IN1(\Reg_Bank/n5766 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5774 ) );
  MUX \Reg_Bank/U5864  ( .IN0(\Reg_Bank/n5772 ), .IN1(\Reg_Bank/n5769 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5773 ) );
  MUX \Reg_Bank/U5863  ( .IN0(\Reg_Bank/n5771 ), .IN1(\Reg_Bank/n5770 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5772 ) );
  MUX \Reg_Bank/U5862  ( .IN0(\Reg_Bank/registers[16][26] ), .IN1(
        \Reg_Bank/registers[17][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5771 )
         );
  MUX \Reg_Bank/U5861  ( .IN0(\Reg_Bank/registers[18][26] ), .IN1(
        \Reg_Bank/registers[19][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5770 )
         );
  MUX \Reg_Bank/U5860  ( .IN0(\Reg_Bank/n5768 ), .IN1(\Reg_Bank/n5767 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5769 ) );
  MUX \Reg_Bank/U5859  ( .IN0(\Reg_Bank/registers[20][26] ), .IN1(
        \Reg_Bank/registers[21][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5768 )
         );
  MUX \Reg_Bank/U5858  ( .IN0(\Reg_Bank/registers[22][26] ), .IN1(
        \Reg_Bank/registers[23][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5767 )
         );
  MUX \Reg_Bank/U5857  ( .IN0(\Reg_Bank/n5765 ), .IN1(\Reg_Bank/n5762 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5766 ) );
  MUX \Reg_Bank/U5856  ( .IN0(\Reg_Bank/n5764 ), .IN1(\Reg_Bank/n5763 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5765 ) );
  MUX \Reg_Bank/U5855  ( .IN0(\Reg_Bank/registers[24][26] ), .IN1(
        \Reg_Bank/registers[25][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5764 )
         );
  MUX \Reg_Bank/U5854  ( .IN0(\Reg_Bank/registers[26][26] ), .IN1(
        \Reg_Bank/registers[27][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5763 )
         );
  MUX \Reg_Bank/U5853  ( .IN0(\Reg_Bank/n5761 ), .IN1(\Reg_Bank/n5760 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5762 ) );
  MUX \Reg_Bank/U5852  ( .IN0(\Reg_Bank/registers[28][26] ), .IN1(
        \Reg_Bank/registers[29][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5761 )
         );
  MUX \Reg_Bank/U5851  ( .IN0(\Reg_Bank/registers[30][26] ), .IN1(
        \Reg_Bank/registers[31][26] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5760 )
         );
  MUX \Reg_Bank/U5850  ( .IN0(\Reg_Bank/n5759 ), .IN1(\Reg_Bank/n5744 ), .SEL(
        rt_index[4]), .F(reg_target[25]) );
  MUX \Reg_Bank/U5849  ( .IN0(\Reg_Bank/n5758 ), .IN1(\Reg_Bank/n5751 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5759 ) );
  MUX \Reg_Bank/U5848  ( .IN0(\Reg_Bank/n5757 ), .IN1(\Reg_Bank/n5754 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5758 ) );
  MUX \Reg_Bank/U5847  ( .IN0(\Reg_Bank/n5756 ), .IN1(\Reg_Bank/n5755 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5757 ) );
  MUX \Reg_Bank/U5845  ( .IN0(\Reg_Bank/registers[2][25] ), .IN1(
        \Reg_Bank/registers[3][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5755 )
         );
  MUX \Reg_Bank/U5844  ( .IN0(\Reg_Bank/n5753 ), .IN1(\Reg_Bank/n5752 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5754 ) );
  MUX \Reg_Bank/U5843  ( .IN0(\Reg_Bank/registers[4][25] ), .IN1(
        \Reg_Bank/registers[5][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5753 )
         );
  MUX \Reg_Bank/U5842  ( .IN0(\Reg_Bank/registers[6][25] ), .IN1(
        \Reg_Bank/registers[7][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5752 )
         );
  MUX \Reg_Bank/U5841  ( .IN0(\Reg_Bank/n5750 ), .IN1(\Reg_Bank/n5747 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5751 ) );
  MUX \Reg_Bank/U5840  ( .IN0(\Reg_Bank/n5749 ), .IN1(\Reg_Bank/n5748 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5750 ) );
  MUX \Reg_Bank/U5839  ( .IN0(\Reg_Bank/registers[8][25] ), .IN1(
        \Reg_Bank/registers[9][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5749 )
         );
  MUX \Reg_Bank/U5838  ( .IN0(\Reg_Bank/registers[10][25] ), .IN1(
        \Reg_Bank/registers[11][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5748 )
         );
  MUX \Reg_Bank/U5837  ( .IN0(\Reg_Bank/n5746 ), .IN1(\Reg_Bank/n5745 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5747 ) );
  MUX \Reg_Bank/U5836  ( .IN0(\Reg_Bank/registers[12][25] ), .IN1(
        \Reg_Bank/registers[13][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5746 )
         );
  MUX \Reg_Bank/U5835  ( .IN0(\Reg_Bank/registers[14][25] ), .IN1(
        \Reg_Bank/registers[15][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5745 )
         );
  MUX \Reg_Bank/U5834  ( .IN0(\Reg_Bank/n5743 ), .IN1(\Reg_Bank/n5736 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5744 ) );
  MUX \Reg_Bank/U5833  ( .IN0(\Reg_Bank/n5742 ), .IN1(\Reg_Bank/n5739 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5743 ) );
  MUX \Reg_Bank/U5832  ( .IN0(\Reg_Bank/n5741 ), .IN1(\Reg_Bank/n5740 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5742 ) );
  MUX \Reg_Bank/U5831  ( .IN0(\Reg_Bank/registers[16][25] ), .IN1(
        \Reg_Bank/registers[17][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5741 )
         );
  MUX \Reg_Bank/U5830  ( .IN0(\Reg_Bank/registers[18][25] ), .IN1(
        \Reg_Bank/registers[19][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5740 )
         );
  MUX \Reg_Bank/U5829  ( .IN0(\Reg_Bank/n5738 ), .IN1(\Reg_Bank/n5737 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5739 ) );
  MUX \Reg_Bank/U5828  ( .IN0(\Reg_Bank/registers[20][25] ), .IN1(
        \Reg_Bank/registers[21][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5738 )
         );
  MUX \Reg_Bank/U5827  ( .IN0(\Reg_Bank/registers[22][25] ), .IN1(
        \Reg_Bank/registers[23][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5737 )
         );
  MUX \Reg_Bank/U5826  ( .IN0(\Reg_Bank/n5735 ), .IN1(\Reg_Bank/n5732 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5736 ) );
  MUX \Reg_Bank/U5825  ( .IN0(\Reg_Bank/n5734 ), .IN1(\Reg_Bank/n5733 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5735 ) );
  MUX \Reg_Bank/U5824  ( .IN0(\Reg_Bank/registers[24][25] ), .IN1(
        \Reg_Bank/registers[25][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5734 )
         );
  MUX \Reg_Bank/U5823  ( .IN0(\Reg_Bank/registers[26][25] ), .IN1(
        \Reg_Bank/registers[27][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5733 )
         );
  MUX \Reg_Bank/U5822  ( .IN0(\Reg_Bank/n5731 ), .IN1(\Reg_Bank/n5730 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5732 ) );
  MUX \Reg_Bank/U5821  ( .IN0(\Reg_Bank/registers[28][25] ), .IN1(
        \Reg_Bank/registers[29][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5731 )
         );
  MUX \Reg_Bank/U5820  ( .IN0(\Reg_Bank/registers[30][25] ), .IN1(
        \Reg_Bank/registers[31][25] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5730 )
         );
  MUX \Reg_Bank/U5819  ( .IN0(\Reg_Bank/n5729 ), .IN1(\Reg_Bank/n5714 ), .SEL(
        rt_index[4]), .F(reg_target[24]) );
  MUX \Reg_Bank/U5818  ( .IN0(\Reg_Bank/n5728 ), .IN1(\Reg_Bank/n5721 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5729 ) );
  MUX \Reg_Bank/U5817  ( .IN0(\Reg_Bank/n5727 ), .IN1(\Reg_Bank/n5724 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5728 ) );
  MUX \Reg_Bank/U5816  ( .IN0(\Reg_Bank/n5726 ), .IN1(\Reg_Bank/n5725 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5727 ) );
  MUX \Reg_Bank/U5814  ( .IN0(\Reg_Bank/registers[2][24] ), .IN1(
        \Reg_Bank/registers[3][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5725 )
         );
  MUX \Reg_Bank/U5813  ( .IN0(\Reg_Bank/n5723 ), .IN1(\Reg_Bank/n5722 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5724 ) );
  MUX \Reg_Bank/U5812  ( .IN0(\Reg_Bank/registers[4][24] ), .IN1(
        \Reg_Bank/registers[5][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5723 )
         );
  MUX \Reg_Bank/U5811  ( .IN0(\Reg_Bank/registers[6][24] ), .IN1(
        \Reg_Bank/registers[7][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5722 )
         );
  MUX \Reg_Bank/U5810  ( .IN0(\Reg_Bank/n5720 ), .IN1(\Reg_Bank/n5717 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5721 ) );
  MUX \Reg_Bank/U5809  ( .IN0(\Reg_Bank/n5719 ), .IN1(\Reg_Bank/n5718 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5720 ) );
  MUX \Reg_Bank/U5808  ( .IN0(\Reg_Bank/registers[8][24] ), .IN1(
        \Reg_Bank/registers[9][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5719 )
         );
  MUX \Reg_Bank/U5807  ( .IN0(\Reg_Bank/registers[10][24] ), .IN1(
        \Reg_Bank/registers[11][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5718 )
         );
  MUX \Reg_Bank/U5806  ( .IN0(\Reg_Bank/n5716 ), .IN1(\Reg_Bank/n5715 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5717 ) );
  MUX \Reg_Bank/U5805  ( .IN0(\Reg_Bank/registers[12][24] ), .IN1(
        \Reg_Bank/registers[13][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5716 )
         );
  MUX \Reg_Bank/U5804  ( .IN0(\Reg_Bank/registers[14][24] ), .IN1(
        \Reg_Bank/registers[15][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5715 )
         );
  MUX \Reg_Bank/U5803  ( .IN0(\Reg_Bank/n5713 ), .IN1(\Reg_Bank/n5706 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5714 ) );
  MUX \Reg_Bank/U5802  ( .IN0(\Reg_Bank/n5712 ), .IN1(\Reg_Bank/n5709 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5713 ) );
  MUX \Reg_Bank/U5801  ( .IN0(\Reg_Bank/n5711 ), .IN1(\Reg_Bank/n5710 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5712 ) );
  MUX \Reg_Bank/U5800  ( .IN0(\Reg_Bank/registers[16][24] ), .IN1(
        \Reg_Bank/registers[17][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5711 )
         );
  MUX \Reg_Bank/U5799  ( .IN0(\Reg_Bank/registers[18][24] ), .IN1(
        \Reg_Bank/registers[19][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5710 )
         );
  MUX \Reg_Bank/U5798  ( .IN0(\Reg_Bank/n5708 ), .IN1(\Reg_Bank/n5707 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5709 ) );
  MUX \Reg_Bank/U5797  ( .IN0(\Reg_Bank/registers[20][24] ), .IN1(
        \Reg_Bank/registers[21][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5708 )
         );
  MUX \Reg_Bank/U5796  ( .IN0(\Reg_Bank/registers[22][24] ), .IN1(
        \Reg_Bank/registers[23][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5707 )
         );
  MUX \Reg_Bank/U5795  ( .IN0(\Reg_Bank/n5705 ), .IN1(\Reg_Bank/n5702 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5706 ) );
  MUX \Reg_Bank/U5794  ( .IN0(\Reg_Bank/n5704 ), .IN1(\Reg_Bank/n5703 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5705 ) );
  MUX \Reg_Bank/U5793  ( .IN0(\Reg_Bank/registers[24][24] ), .IN1(
        \Reg_Bank/registers[25][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5704 )
         );
  MUX \Reg_Bank/U5792  ( .IN0(\Reg_Bank/registers[26][24] ), .IN1(
        \Reg_Bank/registers[27][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5703 )
         );
  MUX \Reg_Bank/U5791  ( .IN0(\Reg_Bank/n5701 ), .IN1(\Reg_Bank/n5700 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5702 ) );
  MUX \Reg_Bank/U5790  ( .IN0(\Reg_Bank/registers[28][24] ), .IN1(
        \Reg_Bank/registers[29][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5701 )
         );
  MUX \Reg_Bank/U5789  ( .IN0(\Reg_Bank/registers[30][24] ), .IN1(
        \Reg_Bank/registers[31][24] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5700 )
         );
  MUX \Reg_Bank/U5788  ( .IN0(\Reg_Bank/n5699 ), .IN1(\Reg_Bank/n5684 ), .SEL(
        rt_index[4]), .F(reg_target[23]) );
  MUX \Reg_Bank/U5787  ( .IN0(\Reg_Bank/n5698 ), .IN1(\Reg_Bank/n5691 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5699 ) );
  MUX \Reg_Bank/U5786  ( .IN0(\Reg_Bank/n5697 ), .IN1(\Reg_Bank/n5694 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5698 ) );
  MUX \Reg_Bank/U5785  ( .IN0(\Reg_Bank/n5696 ), .IN1(\Reg_Bank/n5695 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5697 ) );
  MUX \Reg_Bank/U5783  ( .IN0(\Reg_Bank/registers[2][23] ), .IN1(
        \Reg_Bank/registers[3][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5695 )
         );
  MUX \Reg_Bank/U5782  ( .IN0(\Reg_Bank/n5693 ), .IN1(\Reg_Bank/n5692 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5694 ) );
  MUX \Reg_Bank/U5781  ( .IN0(\Reg_Bank/registers[4][23] ), .IN1(
        \Reg_Bank/registers[5][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5693 )
         );
  MUX \Reg_Bank/U5780  ( .IN0(\Reg_Bank/registers[6][23] ), .IN1(
        \Reg_Bank/registers[7][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5692 )
         );
  MUX \Reg_Bank/U5779  ( .IN0(\Reg_Bank/n5690 ), .IN1(\Reg_Bank/n5687 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5691 ) );
  MUX \Reg_Bank/U5778  ( .IN0(\Reg_Bank/n5689 ), .IN1(\Reg_Bank/n5688 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5690 ) );
  MUX \Reg_Bank/U5777  ( .IN0(\Reg_Bank/registers[8][23] ), .IN1(
        \Reg_Bank/registers[9][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5689 )
         );
  MUX \Reg_Bank/U5776  ( .IN0(\Reg_Bank/registers[10][23] ), .IN1(
        \Reg_Bank/registers[11][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5688 )
         );
  MUX \Reg_Bank/U5775  ( .IN0(\Reg_Bank/n5686 ), .IN1(\Reg_Bank/n5685 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5687 ) );
  MUX \Reg_Bank/U5774  ( .IN0(\Reg_Bank/registers[12][23] ), .IN1(
        \Reg_Bank/registers[13][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5686 )
         );
  MUX \Reg_Bank/U5773  ( .IN0(\Reg_Bank/registers[14][23] ), .IN1(
        \Reg_Bank/registers[15][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5685 )
         );
  MUX \Reg_Bank/U5772  ( .IN0(\Reg_Bank/n5683 ), .IN1(\Reg_Bank/n5676 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5684 ) );
  MUX \Reg_Bank/U5771  ( .IN0(\Reg_Bank/n5682 ), .IN1(\Reg_Bank/n5679 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5683 ) );
  MUX \Reg_Bank/U5770  ( .IN0(\Reg_Bank/n5681 ), .IN1(\Reg_Bank/n5680 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5682 ) );
  MUX \Reg_Bank/U5769  ( .IN0(\Reg_Bank/registers[16][23] ), .IN1(
        \Reg_Bank/registers[17][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5681 )
         );
  MUX \Reg_Bank/U5768  ( .IN0(\Reg_Bank/registers[18][23] ), .IN1(
        \Reg_Bank/registers[19][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5680 )
         );
  MUX \Reg_Bank/U5767  ( .IN0(\Reg_Bank/n5678 ), .IN1(\Reg_Bank/n5677 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5679 ) );
  MUX \Reg_Bank/U5766  ( .IN0(\Reg_Bank/registers[20][23] ), .IN1(
        \Reg_Bank/registers[21][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5678 )
         );
  MUX \Reg_Bank/U5765  ( .IN0(\Reg_Bank/registers[22][23] ), .IN1(
        \Reg_Bank/registers[23][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5677 )
         );
  MUX \Reg_Bank/U5764  ( .IN0(\Reg_Bank/n5675 ), .IN1(\Reg_Bank/n5672 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5676 ) );
  MUX \Reg_Bank/U5763  ( .IN0(\Reg_Bank/n5674 ), .IN1(\Reg_Bank/n5673 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5675 ) );
  MUX \Reg_Bank/U5762  ( .IN0(\Reg_Bank/registers[24][23] ), .IN1(
        \Reg_Bank/registers[25][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5674 )
         );
  MUX \Reg_Bank/U5761  ( .IN0(\Reg_Bank/registers[26][23] ), .IN1(
        \Reg_Bank/registers[27][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5673 )
         );
  MUX \Reg_Bank/U5760  ( .IN0(\Reg_Bank/n5671 ), .IN1(\Reg_Bank/n5670 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5672 ) );
  MUX \Reg_Bank/U5759  ( .IN0(\Reg_Bank/registers[28][23] ), .IN1(
        \Reg_Bank/registers[29][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5671 )
         );
  MUX \Reg_Bank/U5758  ( .IN0(\Reg_Bank/registers[30][23] ), .IN1(
        \Reg_Bank/registers[31][23] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5670 )
         );
  MUX \Reg_Bank/U5757  ( .IN0(\Reg_Bank/n5669 ), .IN1(\Reg_Bank/n5654 ), .SEL(
        rt_index[4]), .F(reg_target[22]) );
  MUX \Reg_Bank/U5756  ( .IN0(\Reg_Bank/n5668 ), .IN1(\Reg_Bank/n5661 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5669 ) );
  MUX \Reg_Bank/U5755  ( .IN0(\Reg_Bank/n5667 ), .IN1(\Reg_Bank/n5664 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5668 ) );
  MUX \Reg_Bank/U5754  ( .IN0(\Reg_Bank/n5666 ), .IN1(\Reg_Bank/n5665 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5667 ) );
  MUX \Reg_Bank/U5752  ( .IN0(\Reg_Bank/registers[2][22] ), .IN1(
        \Reg_Bank/registers[3][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5665 )
         );
  MUX \Reg_Bank/U5751  ( .IN0(\Reg_Bank/n5663 ), .IN1(\Reg_Bank/n5662 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5664 ) );
  MUX \Reg_Bank/U5750  ( .IN0(\Reg_Bank/registers[4][22] ), .IN1(
        \Reg_Bank/registers[5][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5663 )
         );
  MUX \Reg_Bank/U5749  ( .IN0(\Reg_Bank/registers[6][22] ), .IN1(
        \Reg_Bank/registers[7][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5662 )
         );
  MUX \Reg_Bank/U5748  ( .IN0(\Reg_Bank/n5660 ), .IN1(\Reg_Bank/n5657 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5661 ) );
  MUX \Reg_Bank/U5747  ( .IN0(\Reg_Bank/n5659 ), .IN1(\Reg_Bank/n5658 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5660 ) );
  MUX \Reg_Bank/U5746  ( .IN0(\Reg_Bank/registers[8][22] ), .IN1(
        \Reg_Bank/registers[9][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5659 )
         );
  MUX \Reg_Bank/U5745  ( .IN0(\Reg_Bank/registers[10][22] ), .IN1(
        \Reg_Bank/registers[11][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5658 )
         );
  MUX \Reg_Bank/U5744  ( .IN0(\Reg_Bank/n5656 ), .IN1(\Reg_Bank/n5655 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5657 ) );
  MUX \Reg_Bank/U5743  ( .IN0(\Reg_Bank/registers[12][22] ), .IN1(
        \Reg_Bank/registers[13][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5656 )
         );
  MUX \Reg_Bank/U5742  ( .IN0(\Reg_Bank/registers[14][22] ), .IN1(
        \Reg_Bank/registers[15][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5655 )
         );
  MUX \Reg_Bank/U5741  ( .IN0(\Reg_Bank/n5653 ), .IN1(\Reg_Bank/n5646 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5654 ) );
  MUX \Reg_Bank/U5740  ( .IN0(\Reg_Bank/n5652 ), .IN1(\Reg_Bank/n5649 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5653 ) );
  MUX \Reg_Bank/U5739  ( .IN0(\Reg_Bank/n5651 ), .IN1(\Reg_Bank/n5650 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5652 ) );
  MUX \Reg_Bank/U5738  ( .IN0(\Reg_Bank/registers[16][22] ), .IN1(
        \Reg_Bank/registers[17][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5651 )
         );
  MUX \Reg_Bank/U5737  ( .IN0(\Reg_Bank/registers[18][22] ), .IN1(
        \Reg_Bank/registers[19][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5650 )
         );
  MUX \Reg_Bank/U5736  ( .IN0(\Reg_Bank/n5648 ), .IN1(\Reg_Bank/n5647 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5649 ) );
  MUX \Reg_Bank/U5735  ( .IN0(\Reg_Bank/registers[20][22] ), .IN1(
        \Reg_Bank/registers[21][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5648 )
         );
  MUX \Reg_Bank/U5734  ( .IN0(\Reg_Bank/registers[22][22] ), .IN1(
        \Reg_Bank/registers[23][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5647 )
         );
  MUX \Reg_Bank/U5733  ( .IN0(\Reg_Bank/n5645 ), .IN1(\Reg_Bank/n5642 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5646 ) );
  MUX \Reg_Bank/U5732  ( .IN0(\Reg_Bank/n5644 ), .IN1(\Reg_Bank/n5643 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5645 ) );
  MUX \Reg_Bank/U5731  ( .IN0(\Reg_Bank/registers[24][22] ), .IN1(
        \Reg_Bank/registers[25][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5644 )
         );
  MUX \Reg_Bank/U5730  ( .IN0(\Reg_Bank/registers[26][22] ), .IN1(
        \Reg_Bank/registers[27][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5643 )
         );
  MUX \Reg_Bank/U5729  ( .IN0(\Reg_Bank/n5641 ), .IN1(\Reg_Bank/n5640 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5642 ) );
  MUX \Reg_Bank/U5728  ( .IN0(\Reg_Bank/registers[28][22] ), .IN1(
        \Reg_Bank/registers[29][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5641 )
         );
  MUX \Reg_Bank/U5727  ( .IN0(\Reg_Bank/registers[30][22] ), .IN1(
        \Reg_Bank/registers[31][22] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5640 )
         );
  MUX \Reg_Bank/U5726  ( .IN0(\Reg_Bank/n5639 ), .IN1(\Reg_Bank/n5624 ), .SEL(
        rt_index[4]), .F(reg_target[21]) );
  MUX \Reg_Bank/U5725  ( .IN0(\Reg_Bank/n5638 ), .IN1(\Reg_Bank/n5631 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5639 ) );
  MUX \Reg_Bank/U5724  ( .IN0(\Reg_Bank/n5637 ), .IN1(\Reg_Bank/n5634 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5638 ) );
  MUX \Reg_Bank/U5723  ( .IN0(\Reg_Bank/n5636 ), .IN1(\Reg_Bank/n5635 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5637 ) );
  MUX \Reg_Bank/U5721  ( .IN0(\Reg_Bank/registers[2][21] ), .IN1(
        \Reg_Bank/registers[3][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5635 )
         );
  MUX \Reg_Bank/U5720  ( .IN0(\Reg_Bank/n5633 ), .IN1(\Reg_Bank/n5632 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5634 ) );
  MUX \Reg_Bank/U5719  ( .IN0(\Reg_Bank/registers[4][21] ), .IN1(
        \Reg_Bank/registers[5][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5633 )
         );
  MUX \Reg_Bank/U5718  ( .IN0(\Reg_Bank/registers[6][21] ), .IN1(
        \Reg_Bank/registers[7][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5632 )
         );
  MUX \Reg_Bank/U5717  ( .IN0(\Reg_Bank/n5630 ), .IN1(\Reg_Bank/n5627 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5631 ) );
  MUX \Reg_Bank/U5716  ( .IN0(\Reg_Bank/n5629 ), .IN1(\Reg_Bank/n5628 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5630 ) );
  MUX \Reg_Bank/U5715  ( .IN0(\Reg_Bank/registers[8][21] ), .IN1(
        \Reg_Bank/registers[9][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5629 )
         );
  MUX \Reg_Bank/U5714  ( .IN0(\Reg_Bank/registers[10][21] ), .IN1(
        \Reg_Bank/registers[11][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5628 )
         );
  MUX \Reg_Bank/U5713  ( .IN0(\Reg_Bank/n5626 ), .IN1(\Reg_Bank/n5625 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5627 ) );
  MUX \Reg_Bank/U5712  ( .IN0(\Reg_Bank/registers[12][21] ), .IN1(
        \Reg_Bank/registers[13][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5626 )
         );
  MUX \Reg_Bank/U5711  ( .IN0(\Reg_Bank/registers[14][21] ), .IN1(
        \Reg_Bank/registers[15][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5625 )
         );
  MUX \Reg_Bank/U5710  ( .IN0(\Reg_Bank/n5623 ), .IN1(\Reg_Bank/n5616 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5624 ) );
  MUX \Reg_Bank/U5709  ( .IN0(\Reg_Bank/n5622 ), .IN1(\Reg_Bank/n5619 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5623 ) );
  MUX \Reg_Bank/U5708  ( .IN0(\Reg_Bank/n5621 ), .IN1(\Reg_Bank/n5620 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5622 ) );
  MUX \Reg_Bank/U5707  ( .IN0(\Reg_Bank/registers[16][21] ), .IN1(
        \Reg_Bank/registers[17][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5621 )
         );
  MUX \Reg_Bank/U5706  ( .IN0(\Reg_Bank/registers[18][21] ), .IN1(
        \Reg_Bank/registers[19][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5620 )
         );
  MUX \Reg_Bank/U5705  ( .IN0(\Reg_Bank/n5618 ), .IN1(\Reg_Bank/n5617 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5619 ) );
  MUX \Reg_Bank/U5704  ( .IN0(\Reg_Bank/registers[20][21] ), .IN1(
        \Reg_Bank/registers[21][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5618 )
         );
  MUX \Reg_Bank/U5703  ( .IN0(\Reg_Bank/registers[22][21] ), .IN1(
        \Reg_Bank/registers[23][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5617 )
         );
  MUX \Reg_Bank/U5702  ( .IN0(\Reg_Bank/n5615 ), .IN1(\Reg_Bank/n5612 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5616 ) );
  MUX \Reg_Bank/U5701  ( .IN0(\Reg_Bank/n5614 ), .IN1(\Reg_Bank/n5613 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5615 ) );
  MUX \Reg_Bank/U5700  ( .IN0(\Reg_Bank/registers[24][21] ), .IN1(
        \Reg_Bank/registers[25][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5614 )
         );
  MUX \Reg_Bank/U5699  ( .IN0(\Reg_Bank/registers[26][21] ), .IN1(
        \Reg_Bank/registers[27][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5613 )
         );
  MUX \Reg_Bank/U5698  ( .IN0(\Reg_Bank/n5611 ), .IN1(\Reg_Bank/n5610 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5612 ) );
  MUX \Reg_Bank/U5697  ( .IN0(\Reg_Bank/registers[28][21] ), .IN1(
        \Reg_Bank/registers[29][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5611 )
         );
  MUX \Reg_Bank/U5696  ( .IN0(\Reg_Bank/registers[30][21] ), .IN1(
        \Reg_Bank/registers[31][21] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5610 )
         );
  MUX \Reg_Bank/U5695  ( .IN0(\Reg_Bank/n5609 ), .IN1(\Reg_Bank/n5594 ), .SEL(
        rt_index[4]), .F(reg_target[20]) );
  MUX \Reg_Bank/U5694  ( .IN0(\Reg_Bank/n5608 ), .IN1(\Reg_Bank/n5601 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5609 ) );
  MUX \Reg_Bank/U5693  ( .IN0(\Reg_Bank/n5607 ), .IN1(\Reg_Bank/n5604 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5608 ) );
  MUX \Reg_Bank/U5692  ( .IN0(\Reg_Bank/n5606 ), .IN1(\Reg_Bank/n5605 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5607 ) );
  MUX \Reg_Bank/U5690  ( .IN0(\Reg_Bank/registers[2][20] ), .IN1(
        \Reg_Bank/registers[3][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5605 )
         );
  MUX \Reg_Bank/U5689  ( .IN0(\Reg_Bank/n5603 ), .IN1(\Reg_Bank/n5602 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5604 ) );
  MUX \Reg_Bank/U5688  ( .IN0(\Reg_Bank/registers[4][20] ), .IN1(
        \Reg_Bank/registers[5][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5603 )
         );
  MUX \Reg_Bank/U5687  ( .IN0(\Reg_Bank/registers[6][20] ), .IN1(
        \Reg_Bank/registers[7][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5602 )
         );
  MUX \Reg_Bank/U5686  ( .IN0(\Reg_Bank/n5600 ), .IN1(\Reg_Bank/n5597 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5601 ) );
  MUX \Reg_Bank/U5685  ( .IN0(\Reg_Bank/n5599 ), .IN1(\Reg_Bank/n5598 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5600 ) );
  MUX \Reg_Bank/U5684  ( .IN0(\Reg_Bank/registers[8][20] ), .IN1(
        \Reg_Bank/registers[9][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5599 )
         );
  MUX \Reg_Bank/U5683  ( .IN0(\Reg_Bank/registers[10][20] ), .IN1(
        \Reg_Bank/registers[11][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5598 )
         );
  MUX \Reg_Bank/U5682  ( .IN0(\Reg_Bank/n5596 ), .IN1(\Reg_Bank/n5595 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5597 ) );
  MUX \Reg_Bank/U5681  ( .IN0(\Reg_Bank/registers[12][20] ), .IN1(
        \Reg_Bank/registers[13][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5596 )
         );
  MUX \Reg_Bank/U5680  ( .IN0(\Reg_Bank/registers[14][20] ), .IN1(
        \Reg_Bank/registers[15][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5595 )
         );
  MUX \Reg_Bank/U5679  ( .IN0(\Reg_Bank/n5593 ), .IN1(\Reg_Bank/n5586 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5594 ) );
  MUX \Reg_Bank/U5678  ( .IN0(\Reg_Bank/n5592 ), .IN1(\Reg_Bank/n5589 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5593 ) );
  MUX \Reg_Bank/U5677  ( .IN0(\Reg_Bank/n5591 ), .IN1(\Reg_Bank/n5590 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5592 ) );
  MUX \Reg_Bank/U5676  ( .IN0(\Reg_Bank/registers[16][20] ), .IN1(
        \Reg_Bank/registers[17][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5591 )
         );
  MUX \Reg_Bank/U5675  ( .IN0(\Reg_Bank/registers[18][20] ), .IN1(
        \Reg_Bank/registers[19][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5590 )
         );
  MUX \Reg_Bank/U5674  ( .IN0(\Reg_Bank/n5588 ), .IN1(\Reg_Bank/n5587 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5589 ) );
  MUX \Reg_Bank/U5673  ( .IN0(\Reg_Bank/registers[20][20] ), .IN1(
        \Reg_Bank/registers[21][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5588 )
         );
  MUX \Reg_Bank/U5672  ( .IN0(\Reg_Bank/registers[22][20] ), .IN1(
        \Reg_Bank/registers[23][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5587 )
         );
  MUX \Reg_Bank/U5671  ( .IN0(\Reg_Bank/n5585 ), .IN1(\Reg_Bank/n5582 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5586 ) );
  MUX \Reg_Bank/U5670  ( .IN0(\Reg_Bank/n5584 ), .IN1(\Reg_Bank/n5583 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5585 ) );
  MUX \Reg_Bank/U5669  ( .IN0(\Reg_Bank/registers[24][20] ), .IN1(
        \Reg_Bank/registers[25][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5584 )
         );
  MUX \Reg_Bank/U5668  ( .IN0(\Reg_Bank/registers[26][20] ), .IN1(
        \Reg_Bank/registers[27][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5583 )
         );
  MUX \Reg_Bank/U5667  ( .IN0(\Reg_Bank/n5581 ), .IN1(\Reg_Bank/n5580 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5582 ) );
  MUX \Reg_Bank/U5666  ( .IN0(\Reg_Bank/registers[28][20] ), .IN1(
        \Reg_Bank/registers[29][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5581 )
         );
  MUX \Reg_Bank/U5665  ( .IN0(\Reg_Bank/registers[30][20] ), .IN1(
        \Reg_Bank/registers[31][20] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5580 )
         );
  MUX \Reg_Bank/U5664  ( .IN0(\Reg_Bank/n5579 ), .IN1(\Reg_Bank/n5564 ), .SEL(
        rt_index[4]), .F(reg_target[19]) );
  MUX \Reg_Bank/U5663  ( .IN0(\Reg_Bank/n5578 ), .IN1(\Reg_Bank/n5571 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5579 ) );
  MUX \Reg_Bank/U5662  ( .IN0(\Reg_Bank/n5577 ), .IN1(\Reg_Bank/n5574 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5578 ) );
  MUX \Reg_Bank/U5661  ( .IN0(\Reg_Bank/n5576 ), .IN1(\Reg_Bank/n5575 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5577 ) );
  MUX \Reg_Bank/U5659  ( .IN0(\Reg_Bank/registers[2][19] ), .IN1(
        \Reg_Bank/registers[3][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5575 )
         );
  MUX \Reg_Bank/U5658  ( .IN0(\Reg_Bank/n5573 ), .IN1(\Reg_Bank/n5572 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5574 ) );
  MUX \Reg_Bank/U5657  ( .IN0(\Reg_Bank/registers[4][19] ), .IN1(
        \Reg_Bank/registers[5][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5573 )
         );
  MUX \Reg_Bank/U5656  ( .IN0(\Reg_Bank/registers[6][19] ), .IN1(
        \Reg_Bank/registers[7][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5572 )
         );
  MUX \Reg_Bank/U5655  ( .IN0(\Reg_Bank/n5570 ), .IN1(\Reg_Bank/n5567 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5571 ) );
  MUX \Reg_Bank/U5654  ( .IN0(\Reg_Bank/n5569 ), .IN1(\Reg_Bank/n5568 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5570 ) );
  MUX \Reg_Bank/U5653  ( .IN0(\Reg_Bank/registers[8][19] ), .IN1(
        \Reg_Bank/registers[9][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5569 )
         );
  MUX \Reg_Bank/U5652  ( .IN0(\Reg_Bank/registers[10][19] ), .IN1(
        \Reg_Bank/registers[11][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5568 )
         );
  MUX \Reg_Bank/U5651  ( .IN0(\Reg_Bank/n5566 ), .IN1(\Reg_Bank/n5565 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5567 ) );
  MUX \Reg_Bank/U5650  ( .IN0(\Reg_Bank/registers[12][19] ), .IN1(
        \Reg_Bank/registers[13][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5566 )
         );
  MUX \Reg_Bank/U5649  ( .IN0(\Reg_Bank/registers[14][19] ), .IN1(
        \Reg_Bank/registers[15][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5565 )
         );
  MUX \Reg_Bank/U5648  ( .IN0(\Reg_Bank/n5563 ), .IN1(\Reg_Bank/n5556 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5564 ) );
  MUX \Reg_Bank/U5647  ( .IN0(\Reg_Bank/n5562 ), .IN1(\Reg_Bank/n5559 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5563 ) );
  MUX \Reg_Bank/U5646  ( .IN0(\Reg_Bank/n5561 ), .IN1(\Reg_Bank/n5560 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5562 ) );
  MUX \Reg_Bank/U5645  ( .IN0(\Reg_Bank/registers[16][19] ), .IN1(
        \Reg_Bank/registers[17][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5561 )
         );
  MUX \Reg_Bank/U5644  ( .IN0(\Reg_Bank/registers[18][19] ), .IN1(
        \Reg_Bank/registers[19][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5560 )
         );
  MUX \Reg_Bank/U5643  ( .IN0(\Reg_Bank/n5558 ), .IN1(\Reg_Bank/n5557 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5559 ) );
  MUX \Reg_Bank/U5642  ( .IN0(\Reg_Bank/registers[20][19] ), .IN1(
        \Reg_Bank/registers[21][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5558 )
         );
  MUX \Reg_Bank/U5641  ( .IN0(\Reg_Bank/registers[22][19] ), .IN1(
        \Reg_Bank/registers[23][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5557 )
         );
  MUX \Reg_Bank/U5640  ( .IN0(\Reg_Bank/n5555 ), .IN1(\Reg_Bank/n5552 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5556 ) );
  MUX \Reg_Bank/U5639  ( .IN0(\Reg_Bank/n5554 ), .IN1(\Reg_Bank/n5553 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5555 ) );
  MUX \Reg_Bank/U5638  ( .IN0(\Reg_Bank/registers[24][19] ), .IN1(
        \Reg_Bank/registers[25][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5554 )
         );
  MUX \Reg_Bank/U5637  ( .IN0(\Reg_Bank/registers[26][19] ), .IN1(
        \Reg_Bank/registers[27][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5553 )
         );
  MUX \Reg_Bank/U5636  ( .IN0(\Reg_Bank/n5551 ), .IN1(\Reg_Bank/n5550 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5552 ) );
  MUX \Reg_Bank/U5635  ( .IN0(\Reg_Bank/registers[28][19] ), .IN1(
        \Reg_Bank/registers[29][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5551 )
         );
  MUX \Reg_Bank/U5634  ( .IN0(\Reg_Bank/registers[30][19] ), .IN1(
        \Reg_Bank/registers[31][19] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5550 )
         );
  MUX \Reg_Bank/U5633  ( .IN0(\Reg_Bank/n5549 ), .IN1(\Reg_Bank/n5534 ), .SEL(
        rt_index[4]), .F(reg_target[18]) );
  MUX \Reg_Bank/U5632  ( .IN0(\Reg_Bank/n5548 ), .IN1(\Reg_Bank/n5541 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5549 ) );
  MUX \Reg_Bank/U5631  ( .IN0(\Reg_Bank/n5547 ), .IN1(\Reg_Bank/n5544 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5548 ) );
  MUX \Reg_Bank/U5630  ( .IN0(\Reg_Bank/n5546 ), .IN1(\Reg_Bank/n5545 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5547 ) );
  MUX \Reg_Bank/U5628  ( .IN0(\Reg_Bank/registers[2][18] ), .IN1(
        \Reg_Bank/registers[3][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5545 )
         );
  MUX \Reg_Bank/U5627  ( .IN0(\Reg_Bank/n5543 ), .IN1(\Reg_Bank/n5542 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5544 ) );
  MUX \Reg_Bank/U5626  ( .IN0(\Reg_Bank/registers[4][18] ), .IN1(
        \Reg_Bank/registers[5][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5543 )
         );
  MUX \Reg_Bank/U5625  ( .IN0(\Reg_Bank/registers[6][18] ), .IN1(
        \Reg_Bank/registers[7][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5542 )
         );
  MUX \Reg_Bank/U5624  ( .IN0(\Reg_Bank/n5540 ), .IN1(\Reg_Bank/n5537 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5541 ) );
  MUX \Reg_Bank/U5623  ( .IN0(\Reg_Bank/n5539 ), .IN1(\Reg_Bank/n5538 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5540 ) );
  MUX \Reg_Bank/U5622  ( .IN0(\Reg_Bank/registers[8][18] ), .IN1(
        \Reg_Bank/registers[9][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5539 )
         );
  MUX \Reg_Bank/U5621  ( .IN0(\Reg_Bank/registers[10][18] ), .IN1(
        \Reg_Bank/registers[11][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5538 )
         );
  MUX \Reg_Bank/U5620  ( .IN0(\Reg_Bank/n5536 ), .IN1(\Reg_Bank/n5535 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5537 ) );
  MUX \Reg_Bank/U5619  ( .IN0(\Reg_Bank/registers[12][18] ), .IN1(
        \Reg_Bank/registers[13][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5536 )
         );
  MUX \Reg_Bank/U5618  ( .IN0(\Reg_Bank/registers[14][18] ), .IN1(
        \Reg_Bank/registers[15][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5535 )
         );
  MUX \Reg_Bank/U5617  ( .IN0(\Reg_Bank/n5533 ), .IN1(\Reg_Bank/n5526 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5534 ) );
  MUX \Reg_Bank/U5616  ( .IN0(\Reg_Bank/n5532 ), .IN1(\Reg_Bank/n5529 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5533 ) );
  MUX \Reg_Bank/U5615  ( .IN0(\Reg_Bank/n5531 ), .IN1(\Reg_Bank/n5530 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5532 ) );
  MUX \Reg_Bank/U5614  ( .IN0(\Reg_Bank/registers[16][18] ), .IN1(
        \Reg_Bank/registers[17][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5531 )
         );
  MUX \Reg_Bank/U5613  ( .IN0(\Reg_Bank/registers[18][18] ), .IN1(
        \Reg_Bank/registers[19][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5530 )
         );
  MUX \Reg_Bank/U5612  ( .IN0(\Reg_Bank/n5528 ), .IN1(\Reg_Bank/n5527 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5529 ) );
  MUX \Reg_Bank/U5611  ( .IN0(\Reg_Bank/registers[20][18] ), .IN1(
        \Reg_Bank/registers[21][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5528 )
         );
  MUX \Reg_Bank/U5610  ( .IN0(\Reg_Bank/registers[22][18] ), .IN1(
        \Reg_Bank/registers[23][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5527 )
         );
  MUX \Reg_Bank/U5609  ( .IN0(\Reg_Bank/n5525 ), .IN1(\Reg_Bank/n5522 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5526 ) );
  MUX \Reg_Bank/U5608  ( .IN0(\Reg_Bank/n5524 ), .IN1(\Reg_Bank/n5523 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5525 ) );
  MUX \Reg_Bank/U5607  ( .IN0(\Reg_Bank/registers[24][18] ), .IN1(
        \Reg_Bank/registers[25][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5524 )
         );
  MUX \Reg_Bank/U5606  ( .IN0(\Reg_Bank/registers[26][18] ), .IN1(
        \Reg_Bank/registers[27][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5523 )
         );
  MUX \Reg_Bank/U5605  ( .IN0(\Reg_Bank/n5521 ), .IN1(\Reg_Bank/n5520 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5522 ) );
  MUX \Reg_Bank/U5604  ( .IN0(\Reg_Bank/registers[28][18] ), .IN1(
        \Reg_Bank/registers[29][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5521 )
         );
  MUX \Reg_Bank/U5603  ( .IN0(\Reg_Bank/registers[30][18] ), .IN1(
        \Reg_Bank/registers[31][18] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5520 )
         );
  MUX \Reg_Bank/U5602  ( .IN0(\Reg_Bank/n5519 ), .IN1(\Reg_Bank/n5504 ), .SEL(
        rt_index[4]), .F(reg_target[17]) );
  MUX \Reg_Bank/U5601  ( .IN0(\Reg_Bank/n5518 ), .IN1(\Reg_Bank/n5511 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5519 ) );
  MUX \Reg_Bank/U5600  ( .IN0(\Reg_Bank/n5517 ), .IN1(\Reg_Bank/n5514 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5518 ) );
  MUX \Reg_Bank/U5599  ( .IN0(\Reg_Bank/n5516 ), .IN1(\Reg_Bank/n5515 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5517 ) );
  MUX \Reg_Bank/U5597  ( .IN0(\Reg_Bank/registers[2][17] ), .IN1(
        \Reg_Bank/registers[3][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5515 )
         );
  MUX \Reg_Bank/U5596  ( .IN0(\Reg_Bank/n5513 ), .IN1(\Reg_Bank/n5512 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5514 ) );
  MUX \Reg_Bank/U5595  ( .IN0(\Reg_Bank/registers[4][17] ), .IN1(
        \Reg_Bank/registers[5][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5513 )
         );
  MUX \Reg_Bank/U5594  ( .IN0(\Reg_Bank/registers[6][17] ), .IN1(
        \Reg_Bank/registers[7][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5512 )
         );
  MUX \Reg_Bank/U5593  ( .IN0(\Reg_Bank/n5510 ), .IN1(\Reg_Bank/n5507 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5511 ) );
  MUX \Reg_Bank/U5592  ( .IN0(\Reg_Bank/n5509 ), .IN1(\Reg_Bank/n5508 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5510 ) );
  MUX \Reg_Bank/U5591  ( .IN0(\Reg_Bank/registers[8][17] ), .IN1(
        \Reg_Bank/registers[9][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5509 )
         );
  MUX \Reg_Bank/U5590  ( .IN0(\Reg_Bank/registers[10][17] ), .IN1(
        \Reg_Bank/registers[11][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5508 )
         );
  MUX \Reg_Bank/U5589  ( .IN0(\Reg_Bank/n5506 ), .IN1(\Reg_Bank/n5505 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5507 ) );
  MUX \Reg_Bank/U5588  ( .IN0(\Reg_Bank/registers[12][17] ), .IN1(
        \Reg_Bank/registers[13][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5506 )
         );
  MUX \Reg_Bank/U5587  ( .IN0(\Reg_Bank/registers[14][17] ), .IN1(
        \Reg_Bank/registers[15][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5505 )
         );
  MUX \Reg_Bank/U5586  ( .IN0(\Reg_Bank/n5503 ), .IN1(\Reg_Bank/n5496 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5504 ) );
  MUX \Reg_Bank/U5585  ( .IN0(\Reg_Bank/n5502 ), .IN1(\Reg_Bank/n5499 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5503 ) );
  MUX \Reg_Bank/U5584  ( .IN0(\Reg_Bank/n5501 ), .IN1(\Reg_Bank/n5500 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5502 ) );
  MUX \Reg_Bank/U5583  ( .IN0(\Reg_Bank/registers[16][17] ), .IN1(
        \Reg_Bank/registers[17][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5501 )
         );
  MUX \Reg_Bank/U5582  ( .IN0(\Reg_Bank/registers[18][17] ), .IN1(
        \Reg_Bank/registers[19][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5500 )
         );
  MUX \Reg_Bank/U5581  ( .IN0(\Reg_Bank/n5498 ), .IN1(\Reg_Bank/n5497 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5499 ) );
  MUX \Reg_Bank/U5580  ( .IN0(\Reg_Bank/registers[20][17] ), .IN1(
        \Reg_Bank/registers[21][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5498 )
         );
  MUX \Reg_Bank/U5579  ( .IN0(\Reg_Bank/registers[22][17] ), .IN1(
        \Reg_Bank/registers[23][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5497 )
         );
  MUX \Reg_Bank/U5578  ( .IN0(\Reg_Bank/n5495 ), .IN1(\Reg_Bank/n5492 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5496 ) );
  MUX \Reg_Bank/U5577  ( .IN0(\Reg_Bank/n5494 ), .IN1(\Reg_Bank/n5493 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5495 ) );
  MUX \Reg_Bank/U5576  ( .IN0(\Reg_Bank/registers[24][17] ), .IN1(
        \Reg_Bank/registers[25][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5494 )
         );
  MUX \Reg_Bank/U5575  ( .IN0(\Reg_Bank/registers[26][17] ), .IN1(
        \Reg_Bank/registers[27][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5493 )
         );
  MUX \Reg_Bank/U5574  ( .IN0(\Reg_Bank/n5491 ), .IN1(\Reg_Bank/n5490 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5492 ) );
  MUX \Reg_Bank/U5573  ( .IN0(\Reg_Bank/registers[28][17] ), .IN1(
        \Reg_Bank/registers[29][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5491 )
         );
  MUX \Reg_Bank/U5572  ( .IN0(\Reg_Bank/registers[30][17] ), .IN1(
        \Reg_Bank/registers[31][17] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5490 )
         );
  MUX \Reg_Bank/U5571  ( .IN0(\Reg_Bank/n5489 ), .IN1(\Reg_Bank/n5474 ), .SEL(
        rt_index[4]), .F(reg_target[16]) );
  MUX \Reg_Bank/U5570  ( .IN0(\Reg_Bank/n5488 ), .IN1(\Reg_Bank/n5481 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5489 ) );
  MUX \Reg_Bank/U5569  ( .IN0(\Reg_Bank/n5487 ), .IN1(\Reg_Bank/n5484 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5488 ) );
  MUX \Reg_Bank/U5568  ( .IN0(\Reg_Bank/n5486 ), .IN1(\Reg_Bank/n5485 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5487 ) );
  MUX \Reg_Bank/U5566  ( .IN0(\Reg_Bank/registers[2][16] ), .IN1(
        \Reg_Bank/registers[3][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5485 )
         );
  MUX \Reg_Bank/U5565  ( .IN0(\Reg_Bank/n5483 ), .IN1(\Reg_Bank/n5482 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5484 ) );
  MUX \Reg_Bank/U5564  ( .IN0(\Reg_Bank/registers[4][16] ), .IN1(
        \Reg_Bank/registers[5][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5483 )
         );
  MUX \Reg_Bank/U5563  ( .IN0(\Reg_Bank/registers[6][16] ), .IN1(
        \Reg_Bank/registers[7][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5482 )
         );
  MUX \Reg_Bank/U5562  ( .IN0(\Reg_Bank/n5480 ), .IN1(\Reg_Bank/n5477 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5481 ) );
  MUX \Reg_Bank/U5561  ( .IN0(\Reg_Bank/n5479 ), .IN1(\Reg_Bank/n5478 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5480 ) );
  MUX \Reg_Bank/U5560  ( .IN0(\Reg_Bank/registers[8][16] ), .IN1(
        \Reg_Bank/registers[9][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5479 )
         );
  MUX \Reg_Bank/U5559  ( .IN0(\Reg_Bank/registers[10][16] ), .IN1(
        \Reg_Bank/registers[11][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5478 )
         );
  MUX \Reg_Bank/U5558  ( .IN0(\Reg_Bank/n5476 ), .IN1(\Reg_Bank/n5475 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5477 ) );
  MUX \Reg_Bank/U5557  ( .IN0(\Reg_Bank/registers[12][16] ), .IN1(
        \Reg_Bank/registers[13][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5476 )
         );
  MUX \Reg_Bank/U5556  ( .IN0(\Reg_Bank/registers[14][16] ), .IN1(
        \Reg_Bank/registers[15][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5475 )
         );
  MUX \Reg_Bank/U5555  ( .IN0(\Reg_Bank/n5473 ), .IN1(\Reg_Bank/n5466 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5474 ) );
  MUX \Reg_Bank/U5554  ( .IN0(\Reg_Bank/n5472 ), .IN1(\Reg_Bank/n5469 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5473 ) );
  MUX \Reg_Bank/U5553  ( .IN0(\Reg_Bank/n5471 ), .IN1(\Reg_Bank/n5470 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5472 ) );
  MUX \Reg_Bank/U5552  ( .IN0(\Reg_Bank/registers[16][16] ), .IN1(
        \Reg_Bank/registers[17][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5471 )
         );
  MUX \Reg_Bank/U5551  ( .IN0(\Reg_Bank/registers[18][16] ), .IN1(
        \Reg_Bank/registers[19][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5470 )
         );
  MUX \Reg_Bank/U5550  ( .IN0(\Reg_Bank/n5468 ), .IN1(\Reg_Bank/n5467 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5469 ) );
  MUX \Reg_Bank/U5549  ( .IN0(\Reg_Bank/registers[20][16] ), .IN1(
        \Reg_Bank/registers[21][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5468 )
         );
  MUX \Reg_Bank/U5548  ( .IN0(\Reg_Bank/registers[22][16] ), .IN1(
        \Reg_Bank/registers[23][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5467 )
         );
  MUX \Reg_Bank/U5547  ( .IN0(\Reg_Bank/n5465 ), .IN1(\Reg_Bank/n5462 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5466 ) );
  MUX \Reg_Bank/U5546  ( .IN0(\Reg_Bank/n5464 ), .IN1(\Reg_Bank/n5463 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5465 ) );
  MUX \Reg_Bank/U5545  ( .IN0(\Reg_Bank/registers[24][16] ), .IN1(
        \Reg_Bank/registers[25][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5464 )
         );
  MUX \Reg_Bank/U5544  ( .IN0(\Reg_Bank/registers[26][16] ), .IN1(
        \Reg_Bank/registers[27][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5463 )
         );
  MUX \Reg_Bank/U5543  ( .IN0(\Reg_Bank/n5461 ), .IN1(\Reg_Bank/n5460 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5462 ) );
  MUX \Reg_Bank/U5542  ( .IN0(\Reg_Bank/registers[28][16] ), .IN1(
        \Reg_Bank/registers[29][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5461 )
         );
  MUX \Reg_Bank/U5541  ( .IN0(\Reg_Bank/registers[30][16] ), .IN1(
        \Reg_Bank/registers[31][16] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5460 )
         );
  MUX \Reg_Bank/U5540  ( .IN0(\Reg_Bank/n5459 ), .IN1(\Reg_Bank/n5444 ), .SEL(
        rt_index[4]), .F(reg_target[15]) );
  MUX \Reg_Bank/U5539  ( .IN0(\Reg_Bank/n5458 ), .IN1(\Reg_Bank/n5451 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5459 ) );
  MUX \Reg_Bank/U5538  ( .IN0(\Reg_Bank/n5457 ), .IN1(\Reg_Bank/n5454 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5458 ) );
  MUX \Reg_Bank/U5537  ( .IN0(\Reg_Bank/n5456 ), .IN1(\Reg_Bank/n5455 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5457 ) );
  MUX \Reg_Bank/U5535  ( .IN0(\Reg_Bank/registers[2][15] ), .IN1(
        \Reg_Bank/registers[3][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5455 )
         );
  MUX \Reg_Bank/U5534  ( .IN0(\Reg_Bank/n5453 ), .IN1(\Reg_Bank/n5452 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5454 ) );
  MUX \Reg_Bank/U5533  ( .IN0(\Reg_Bank/registers[4][15] ), .IN1(
        \Reg_Bank/registers[5][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5453 )
         );
  MUX \Reg_Bank/U5532  ( .IN0(\Reg_Bank/registers[6][15] ), .IN1(
        \Reg_Bank/registers[7][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5452 )
         );
  MUX \Reg_Bank/U5531  ( .IN0(\Reg_Bank/n5450 ), .IN1(\Reg_Bank/n5447 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5451 ) );
  MUX \Reg_Bank/U5530  ( .IN0(\Reg_Bank/n5449 ), .IN1(\Reg_Bank/n5448 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5450 ) );
  MUX \Reg_Bank/U5529  ( .IN0(\Reg_Bank/registers[8][15] ), .IN1(
        \Reg_Bank/registers[9][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5449 )
         );
  MUX \Reg_Bank/U5528  ( .IN0(\Reg_Bank/registers[10][15] ), .IN1(
        \Reg_Bank/registers[11][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5448 )
         );
  MUX \Reg_Bank/U5527  ( .IN0(\Reg_Bank/n5446 ), .IN1(\Reg_Bank/n5445 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5447 ) );
  MUX \Reg_Bank/U5526  ( .IN0(\Reg_Bank/registers[12][15] ), .IN1(
        \Reg_Bank/registers[13][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5446 )
         );
  MUX \Reg_Bank/U5525  ( .IN0(\Reg_Bank/registers[14][15] ), .IN1(
        \Reg_Bank/registers[15][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5445 )
         );
  MUX \Reg_Bank/U5524  ( .IN0(\Reg_Bank/n5443 ), .IN1(\Reg_Bank/n5436 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5444 ) );
  MUX \Reg_Bank/U5523  ( .IN0(\Reg_Bank/n5442 ), .IN1(\Reg_Bank/n5439 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5443 ) );
  MUX \Reg_Bank/U5522  ( .IN0(\Reg_Bank/n5441 ), .IN1(\Reg_Bank/n5440 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5442 ) );
  MUX \Reg_Bank/U5521  ( .IN0(\Reg_Bank/registers[16][15] ), .IN1(
        \Reg_Bank/registers[17][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5441 )
         );
  MUX \Reg_Bank/U5520  ( .IN0(\Reg_Bank/registers[18][15] ), .IN1(
        \Reg_Bank/registers[19][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5440 )
         );
  MUX \Reg_Bank/U5519  ( .IN0(\Reg_Bank/n5438 ), .IN1(\Reg_Bank/n5437 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5439 ) );
  MUX \Reg_Bank/U5518  ( .IN0(\Reg_Bank/registers[20][15] ), .IN1(
        \Reg_Bank/registers[21][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5438 )
         );
  MUX \Reg_Bank/U5517  ( .IN0(\Reg_Bank/registers[22][15] ), .IN1(
        \Reg_Bank/registers[23][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5437 )
         );
  MUX \Reg_Bank/U5516  ( .IN0(\Reg_Bank/n5435 ), .IN1(\Reg_Bank/n5432 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5436 ) );
  MUX \Reg_Bank/U5515  ( .IN0(\Reg_Bank/n5434 ), .IN1(\Reg_Bank/n5433 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5435 ) );
  MUX \Reg_Bank/U5514  ( .IN0(\Reg_Bank/registers[24][15] ), .IN1(
        \Reg_Bank/registers[25][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5434 )
         );
  MUX \Reg_Bank/U5513  ( .IN0(\Reg_Bank/registers[26][15] ), .IN1(
        \Reg_Bank/registers[27][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5433 )
         );
  MUX \Reg_Bank/U5512  ( .IN0(\Reg_Bank/n5431 ), .IN1(\Reg_Bank/n5430 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5432 ) );
  MUX \Reg_Bank/U5511  ( .IN0(\Reg_Bank/registers[28][15] ), .IN1(
        \Reg_Bank/registers[29][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5431 )
         );
  MUX \Reg_Bank/U5510  ( .IN0(\Reg_Bank/registers[30][15] ), .IN1(
        \Reg_Bank/registers[31][15] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5430 )
         );
  MUX \Reg_Bank/U5509  ( .IN0(\Reg_Bank/n5429 ), .IN1(\Reg_Bank/n5414 ), .SEL(
        rt_index[4]), .F(reg_target[14]) );
  MUX \Reg_Bank/U5508  ( .IN0(\Reg_Bank/n5428 ), .IN1(\Reg_Bank/n5421 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5429 ) );
  MUX \Reg_Bank/U5507  ( .IN0(\Reg_Bank/n5427 ), .IN1(\Reg_Bank/n5424 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5428 ) );
  MUX \Reg_Bank/U5506  ( .IN0(\Reg_Bank/n5426 ), .IN1(\Reg_Bank/n5425 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5427 ) );
  MUX \Reg_Bank/U5504  ( .IN0(\Reg_Bank/registers[2][14] ), .IN1(
        \Reg_Bank/registers[3][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5425 )
         );
  MUX \Reg_Bank/U5503  ( .IN0(\Reg_Bank/n5423 ), .IN1(\Reg_Bank/n5422 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5424 ) );
  MUX \Reg_Bank/U5502  ( .IN0(\Reg_Bank/registers[4][14] ), .IN1(
        \Reg_Bank/registers[5][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5423 )
         );
  MUX \Reg_Bank/U5501  ( .IN0(\Reg_Bank/registers[6][14] ), .IN1(
        \Reg_Bank/registers[7][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5422 )
         );
  MUX \Reg_Bank/U5500  ( .IN0(\Reg_Bank/n5420 ), .IN1(\Reg_Bank/n5417 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5421 ) );
  MUX \Reg_Bank/U5499  ( .IN0(\Reg_Bank/n5419 ), .IN1(\Reg_Bank/n5418 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5420 ) );
  MUX \Reg_Bank/U5498  ( .IN0(\Reg_Bank/registers[8][14] ), .IN1(
        \Reg_Bank/registers[9][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5419 )
         );
  MUX \Reg_Bank/U5497  ( .IN0(\Reg_Bank/registers[10][14] ), .IN1(
        \Reg_Bank/registers[11][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5418 )
         );
  MUX \Reg_Bank/U5496  ( .IN0(\Reg_Bank/n5416 ), .IN1(\Reg_Bank/n5415 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5417 ) );
  MUX \Reg_Bank/U5495  ( .IN0(\Reg_Bank/registers[12][14] ), .IN1(
        \Reg_Bank/registers[13][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5416 )
         );
  MUX \Reg_Bank/U5494  ( .IN0(\Reg_Bank/registers[14][14] ), .IN1(
        \Reg_Bank/registers[15][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5415 )
         );
  MUX \Reg_Bank/U5493  ( .IN0(\Reg_Bank/n5413 ), .IN1(\Reg_Bank/n5406 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5414 ) );
  MUX \Reg_Bank/U5492  ( .IN0(\Reg_Bank/n5412 ), .IN1(\Reg_Bank/n5409 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5413 ) );
  MUX \Reg_Bank/U5491  ( .IN0(\Reg_Bank/n5411 ), .IN1(\Reg_Bank/n5410 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5412 ) );
  MUX \Reg_Bank/U5490  ( .IN0(\Reg_Bank/registers[16][14] ), .IN1(
        \Reg_Bank/registers[17][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5411 )
         );
  MUX \Reg_Bank/U5489  ( .IN0(\Reg_Bank/registers[18][14] ), .IN1(
        \Reg_Bank/registers[19][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5410 )
         );
  MUX \Reg_Bank/U5488  ( .IN0(\Reg_Bank/n5408 ), .IN1(\Reg_Bank/n5407 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5409 ) );
  MUX \Reg_Bank/U5487  ( .IN0(\Reg_Bank/registers[20][14] ), .IN1(
        \Reg_Bank/registers[21][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5408 )
         );
  MUX \Reg_Bank/U5486  ( .IN0(\Reg_Bank/registers[22][14] ), .IN1(
        \Reg_Bank/registers[23][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5407 )
         );
  MUX \Reg_Bank/U5485  ( .IN0(\Reg_Bank/n5405 ), .IN1(\Reg_Bank/n5402 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5406 ) );
  MUX \Reg_Bank/U5484  ( .IN0(\Reg_Bank/n5404 ), .IN1(\Reg_Bank/n5403 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5405 ) );
  MUX \Reg_Bank/U5483  ( .IN0(\Reg_Bank/registers[24][14] ), .IN1(
        \Reg_Bank/registers[25][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5404 )
         );
  MUX \Reg_Bank/U5482  ( .IN0(\Reg_Bank/registers[26][14] ), .IN1(
        \Reg_Bank/registers[27][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5403 )
         );
  MUX \Reg_Bank/U5481  ( .IN0(\Reg_Bank/n5401 ), .IN1(\Reg_Bank/n5400 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5402 ) );
  MUX \Reg_Bank/U5480  ( .IN0(\Reg_Bank/registers[28][14] ), .IN1(
        \Reg_Bank/registers[29][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5401 )
         );
  MUX \Reg_Bank/U5479  ( .IN0(\Reg_Bank/registers[30][14] ), .IN1(
        \Reg_Bank/registers[31][14] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5400 )
         );
  MUX \Reg_Bank/U5478  ( .IN0(\Reg_Bank/n5399 ), .IN1(\Reg_Bank/n5384 ), .SEL(
        rt_index[4]), .F(reg_target[13]) );
  MUX \Reg_Bank/U5477  ( .IN0(\Reg_Bank/n5398 ), .IN1(\Reg_Bank/n5391 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5399 ) );
  MUX \Reg_Bank/U5476  ( .IN0(\Reg_Bank/n5397 ), .IN1(\Reg_Bank/n5394 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5398 ) );
  MUX \Reg_Bank/U5475  ( .IN0(\Reg_Bank/n5396 ), .IN1(\Reg_Bank/n5395 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5397 ) );
  MUX \Reg_Bank/U5473  ( .IN0(\Reg_Bank/registers[2][13] ), .IN1(
        \Reg_Bank/registers[3][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5395 )
         );
  MUX \Reg_Bank/U5472  ( .IN0(\Reg_Bank/n5393 ), .IN1(\Reg_Bank/n5392 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5394 ) );
  MUX \Reg_Bank/U5471  ( .IN0(\Reg_Bank/registers[4][13] ), .IN1(
        \Reg_Bank/registers[5][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5393 )
         );
  MUX \Reg_Bank/U5470  ( .IN0(\Reg_Bank/registers[6][13] ), .IN1(
        \Reg_Bank/registers[7][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5392 )
         );
  MUX \Reg_Bank/U5469  ( .IN0(\Reg_Bank/n5390 ), .IN1(\Reg_Bank/n5387 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5391 ) );
  MUX \Reg_Bank/U5468  ( .IN0(\Reg_Bank/n5389 ), .IN1(\Reg_Bank/n5388 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5390 ) );
  MUX \Reg_Bank/U5467  ( .IN0(\Reg_Bank/registers[8][13] ), .IN1(
        \Reg_Bank/registers[9][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5389 )
         );
  MUX \Reg_Bank/U5466  ( .IN0(\Reg_Bank/registers[10][13] ), .IN1(
        \Reg_Bank/registers[11][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5388 )
         );
  MUX \Reg_Bank/U5465  ( .IN0(\Reg_Bank/n5386 ), .IN1(\Reg_Bank/n5385 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5387 ) );
  MUX \Reg_Bank/U5464  ( .IN0(\Reg_Bank/registers[12][13] ), .IN1(
        \Reg_Bank/registers[13][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5386 )
         );
  MUX \Reg_Bank/U5463  ( .IN0(\Reg_Bank/registers[14][13] ), .IN1(
        \Reg_Bank/registers[15][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5385 )
         );
  MUX \Reg_Bank/U5462  ( .IN0(\Reg_Bank/n5383 ), .IN1(\Reg_Bank/n5376 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5384 ) );
  MUX \Reg_Bank/U5461  ( .IN0(\Reg_Bank/n5382 ), .IN1(\Reg_Bank/n5379 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5383 ) );
  MUX \Reg_Bank/U5460  ( .IN0(\Reg_Bank/n5381 ), .IN1(\Reg_Bank/n5380 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5382 ) );
  MUX \Reg_Bank/U5459  ( .IN0(\Reg_Bank/registers[16][13] ), .IN1(
        \Reg_Bank/registers[17][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5381 )
         );
  MUX \Reg_Bank/U5458  ( .IN0(\Reg_Bank/registers[18][13] ), .IN1(
        \Reg_Bank/registers[19][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5380 )
         );
  MUX \Reg_Bank/U5457  ( .IN0(\Reg_Bank/n5378 ), .IN1(\Reg_Bank/n5377 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5379 ) );
  MUX \Reg_Bank/U5456  ( .IN0(\Reg_Bank/registers[20][13] ), .IN1(
        \Reg_Bank/registers[21][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5378 )
         );
  MUX \Reg_Bank/U5455  ( .IN0(\Reg_Bank/registers[22][13] ), .IN1(
        \Reg_Bank/registers[23][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5377 )
         );
  MUX \Reg_Bank/U5454  ( .IN0(\Reg_Bank/n5375 ), .IN1(\Reg_Bank/n5372 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5376 ) );
  MUX \Reg_Bank/U5453  ( .IN0(\Reg_Bank/n5374 ), .IN1(\Reg_Bank/n5373 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5375 ) );
  MUX \Reg_Bank/U5452  ( .IN0(\Reg_Bank/registers[24][13] ), .IN1(
        \Reg_Bank/registers[25][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5374 )
         );
  MUX \Reg_Bank/U5451  ( .IN0(\Reg_Bank/registers[26][13] ), .IN1(
        \Reg_Bank/registers[27][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5373 )
         );
  MUX \Reg_Bank/U5450  ( .IN0(\Reg_Bank/n5371 ), .IN1(\Reg_Bank/n5370 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5372 ) );
  MUX \Reg_Bank/U5449  ( .IN0(\Reg_Bank/registers[28][13] ), .IN1(
        \Reg_Bank/registers[29][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5371 )
         );
  MUX \Reg_Bank/U5448  ( .IN0(\Reg_Bank/registers[30][13] ), .IN1(
        \Reg_Bank/registers[31][13] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5370 )
         );
  MUX \Reg_Bank/U5447  ( .IN0(\Reg_Bank/n5369 ), .IN1(\Reg_Bank/n5354 ), .SEL(
        rt_index[4]), .F(reg_target[12]) );
  MUX \Reg_Bank/U5446  ( .IN0(\Reg_Bank/n5368 ), .IN1(\Reg_Bank/n5361 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5369 ) );
  MUX \Reg_Bank/U5445  ( .IN0(\Reg_Bank/n5367 ), .IN1(\Reg_Bank/n5364 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5368 ) );
  MUX \Reg_Bank/U5444  ( .IN0(\Reg_Bank/n5366 ), .IN1(\Reg_Bank/n5365 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5367 ) );
  MUX \Reg_Bank/U5442  ( .IN0(\Reg_Bank/registers[2][12] ), .IN1(
        \Reg_Bank/registers[3][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5365 )
         );
  MUX \Reg_Bank/U5441  ( .IN0(\Reg_Bank/n5363 ), .IN1(\Reg_Bank/n5362 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5364 ) );
  MUX \Reg_Bank/U5440  ( .IN0(\Reg_Bank/registers[4][12] ), .IN1(
        \Reg_Bank/registers[5][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5363 )
         );
  MUX \Reg_Bank/U5439  ( .IN0(\Reg_Bank/registers[6][12] ), .IN1(
        \Reg_Bank/registers[7][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5362 )
         );
  MUX \Reg_Bank/U5438  ( .IN0(\Reg_Bank/n5360 ), .IN1(\Reg_Bank/n5357 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5361 ) );
  MUX \Reg_Bank/U5437  ( .IN0(\Reg_Bank/n5359 ), .IN1(\Reg_Bank/n5358 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5360 ) );
  MUX \Reg_Bank/U5436  ( .IN0(\Reg_Bank/registers[8][12] ), .IN1(
        \Reg_Bank/registers[9][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5359 )
         );
  MUX \Reg_Bank/U5435  ( .IN0(\Reg_Bank/registers[10][12] ), .IN1(
        \Reg_Bank/registers[11][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5358 )
         );
  MUX \Reg_Bank/U5434  ( .IN0(\Reg_Bank/n5356 ), .IN1(\Reg_Bank/n5355 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5357 ) );
  MUX \Reg_Bank/U5433  ( .IN0(\Reg_Bank/registers[12][12] ), .IN1(
        \Reg_Bank/registers[13][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5356 )
         );
  MUX \Reg_Bank/U5432  ( .IN0(\Reg_Bank/registers[14][12] ), .IN1(
        \Reg_Bank/registers[15][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5355 )
         );
  MUX \Reg_Bank/U5431  ( .IN0(\Reg_Bank/n5353 ), .IN1(\Reg_Bank/n5346 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5354 ) );
  MUX \Reg_Bank/U5430  ( .IN0(\Reg_Bank/n5352 ), .IN1(\Reg_Bank/n5349 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5353 ) );
  MUX \Reg_Bank/U5429  ( .IN0(\Reg_Bank/n5351 ), .IN1(\Reg_Bank/n5350 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5352 ) );
  MUX \Reg_Bank/U5428  ( .IN0(\Reg_Bank/registers[16][12] ), .IN1(
        \Reg_Bank/registers[17][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5351 )
         );
  MUX \Reg_Bank/U5427  ( .IN0(\Reg_Bank/registers[18][12] ), .IN1(
        \Reg_Bank/registers[19][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5350 )
         );
  MUX \Reg_Bank/U5426  ( .IN0(\Reg_Bank/n5348 ), .IN1(\Reg_Bank/n5347 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5349 ) );
  MUX \Reg_Bank/U5425  ( .IN0(\Reg_Bank/registers[20][12] ), .IN1(
        \Reg_Bank/registers[21][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5348 )
         );
  MUX \Reg_Bank/U5424  ( .IN0(\Reg_Bank/registers[22][12] ), .IN1(
        \Reg_Bank/registers[23][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5347 )
         );
  MUX \Reg_Bank/U5423  ( .IN0(\Reg_Bank/n5345 ), .IN1(\Reg_Bank/n5342 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5346 ) );
  MUX \Reg_Bank/U5422  ( .IN0(\Reg_Bank/n5344 ), .IN1(\Reg_Bank/n5343 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5345 ) );
  MUX \Reg_Bank/U5421  ( .IN0(\Reg_Bank/registers[24][12] ), .IN1(
        \Reg_Bank/registers[25][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5344 )
         );
  MUX \Reg_Bank/U5420  ( .IN0(\Reg_Bank/registers[26][12] ), .IN1(
        \Reg_Bank/registers[27][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5343 )
         );
  MUX \Reg_Bank/U5419  ( .IN0(\Reg_Bank/n5341 ), .IN1(\Reg_Bank/n5340 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5342 ) );
  MUX \Reg_Bank/U5418  ( .IN0(\Reg_Bank/registers[28][12] ), .IN1(
        \Reg_Bank/registers[29][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5341 )
         );
  MUX \Reg_Bank/U5417  ( .IN0(\Reg_Bank/registers[30][12] ), .IN1(
        \Reg_Bank/registers[31][12] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5340 )
         );
  MUX \Reg_Bank/U5416  ( .IN0(\Reg_Bank/n5339 ), .IN1(\Reg_Bank/n5324 ), .SEL(
        rt_index[4]), .F(reg_target[11]) );
  MUX \Reg_Bank/U5415  ( .IN0(\Reg_Bank/n5338 ), .IN1(\Reg_Bank/n5331 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5339 ) );
  MUX \Reg_Bank/U5414  ( .IN0(\Reg_Bank/n5337 ), .IN1(\Reg_Bank/n5334 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5338 ) );
  MUX \Reg_Bank/U5413  ( .IN0(\Reg_Bank/n5336 ), .IN1(\Reg_Bank/n5335 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5337 ) );
  MUX \Reg_Bank/U5411  ( .IN0(\Reg_Bank/registers[2][11] ), .IN1(
        \Reg_Bank/registers[3][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5335 )
         );
  MUX \Reg_Bank/U5410  ( .IN0(\Reg_Bank/n5333 ), .IN1(\Reg_Bank/n5332 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5334 ) );
  MUX \Reg_Bank/U5409  ( .IN0(\Reg_Bank/registers[4][11] ), .IN1(
        \Reg_Bank/registers[5][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5333 )
         );
  MUX \Reg_Bank/U5408  ( .IN0(\Reg_Bank/registers[6][11] ), .IN1(
        \Reg_Bank/registers[7][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5332 )
         );
  MUX \Reg_Bank/U5407  ( .IN0(\Reg_Bank/n5330 ), .IN1(\Reg_Bank/n5327 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5331 ) );
  MUX \Reg_Bank/U5406  ( .IN0(\Reg_Bank/n5329 ), .IN1(\Reg_Bank/n5328 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5330 ) );
  MUX \Reg_Bank/U5405  ( .IN0(\Reg_Bank/registers[8][11] ), .IN1(
        \Reg_Bank/registers[9][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5329 )
         );
  MUX \Reg_Bank/U5404  ( .IN0(\Reg_Bank/registers[10][11] ), .IN1(
        \Reg_Bank/registers[11][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5328 )
         );
  MUX \Reg_Bank/U5403  ( .IN0(\Reg_Bank/n5326 ), .IN1(\Reg_Bank/n5325 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5327 ) );
  MUX \Reg_Bank/U5402  ( .IN0(\Reg_Bank/registers[12][11] ), .IN1(
        \Reg_Bank/registers[13][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5326 )
         );
  MUX \Reg_Bank/U5401  ( .IN0(\Reg_Bank/registers[14][11] ), .IN1(
        \Reg_Bank/registers[15][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5325 )
         );
  MUX \Reg_Bank/U5400  ( .IN0(\Reg_Bank/n5323 ), .IN1(\Reg_Bank/n5316 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5324 ) );
  MUX \Reg_Bank/U5399  ( .IN0(\Reg_Bank/n5322 ), .IN1(\Reg_Bank/n5319 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5323 ) );
  MUX \Reg_Bank/U5398  ( .IN0(\Reg_Bank/n5321 ), .IN1(\Reg_Bank/n5320 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5322 ) );
  MUX \Reg_Bank/U5397  ( .IN0(\Reg_Bank/registers[16][11] ), .IN1(
        \Reg_Bank/registers[17][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5321 )
         );
  MUX \Reg_Bank/U5396  ( .IN0(\Reg_Bank/registers[18][11] ), .IN1(
        \Reg_Bank/registers[19][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5320 )
         );
  MUX \Reg_Bank/U5395  ( .IN0(\Reg_Bank/n5318 ), .IN1(\Reg_Bank/n5317 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5319 ) );
  MUX \Reg_Bank/U5394  ( .IN0(\Reg_Bank/registers[20][11] ), .IN1(
        \Reg_Bank/registers[21][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5318 )
         );
  MUX \Reg_Bank/U5393  ( .IN0(\Reg_Bank/registers[22][11] ), .IN1(
        \Reg_Bank/registers[23][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5317 )
         );
  MUX \Reg_Bank/U5392  ( .IN0(\Reg_Bank/n5315 ), .IN1(\Reg_Bank/n5312 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5316 ) );
  MUX \Reg_Bank/U5391  ( .IN0(\Reg_Bank/n5314 ), .IN1(\Reg_Bank/n5313 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5315 ) );
  MUX \Reg_Bank/U5390  ( .IN0(\Reg_Bank/registers[24][11] ), .IN1(
        \Reg_Bank/registers[25][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5314 )
         );
  MUX \Reg_Bank/U5389  ( .IN0(\Reg_Bank/registers[26][11] ), .IN1(
        \Reg_Bank/registers[27][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5313 )
         );
  MUX \Reg_Bank/U5388  ( .IN0(\Reg_Bank/n5311 ), .IN1(\Reg_Bank/n5310 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5312 ) );
  MUX \Reg_Bank/U5387  ( .IN0(\Reg_Bank/registers[28][11] ), .IN1(
        \Reg_Bank/registers[29][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5311 )
         );
  MUX \Reg_Bank/U5386  ( .IN0(\Reg_Bank/registers[30][11] ), .IN1(
        \Reg_Bank/registers[31][11] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5310 )
         );
  MUX \Reg_Bank/U5385  ( .IN0(\Reg_Bank/n5309 ), .IN1(\Reg_Bank/n5294 ), .SEL(
        rt_index[4]), .F(reg_target[10]) );
  MUX \Reg_Bank/U5384  ( .IN0(\Reg_Bank/n5308 ), .IN1(\Reg_Bank/n5301 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5309 ) );
  MUX \Reg_Bank/U5383  ( .IN0(\Reg_Bank/n5307 ), .IN1(\Reg_Bank/n5304 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5308 ) );
  MUX \Reg_Bank/U5382  ( .IN0(\Reg_Bank/n5306 ), .IN1(\Reg_Bank/n5305 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5307 ) );
  MUX \Reg_Bank/U5380  ( .IN0(\Reg_Bank/registers[2][10] ), .IN1(
        \Reg_Bank/registers[3][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5305 )
         );
  MUX \Reg_Bank/U5379  ( .IN0(\Reg_Bank/n5303 ), .IN1(\Reg_Bank/n5302 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5304 ) );
  MUX \Reg_Bank/U5378  ( .IN0(\Reg_Bank/registers[4][10] ), .IN1(
        \Reg_Bank/registers[5][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5303 )
         );
  MUX \Reg_Bank/U5377  ( .IN0(\Reg_Bank/registers[6][10] ), .IN1(
        \Reg_Bank/registers[7][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5302 )
         );
  MUX \Reg_Bank/U5376  ( .IN0(\Reg_Bank/n5300 ), .IN1(\Reg_Bank/n5297 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5301 ) );
  MUX \Reg_Bank/U5375  ( .IN0(\Reg_Bank/n5299 ), .IN1(\Reg_Bank/n5298 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5300 ) );
  MUX \Reg_Bank/U5374  ( .IN0(\Reg_Bank/registers[8][10] ), .IN1(
        \Reg_Bank/registers[9][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5299 )
         );
  MUX \Reg_Bank/U5373  ( .IN0(\Reg_Bank/registers[10][10] ), .IN1(
        \Reg_Bank/registers[11][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5298 )
         );
  MUX \Reg_Bank/U5372  ( .IN0(\Reg_Bank/n5296 ), .IN1(\Reg_Bank/n5295 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5297 ) );
  MUX \Reg_Bank/U5371  ( .IN0(\Reg_Bank/registers[12][10] ), .IN1(
        \Reg_Bank/registers[13][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5296 )
         );
  MUX \Reg_Bank/U5370  ( .IN0(\Reg_Bank/registers[14][10] ), .IN1(
        \Reg_Bank/registers[15][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5295 )
         );
  MUX \Reg_Bank/U5369  ( .IN0(\Reg_Bank/n5293 ), .IN1(\Reg_Bank/n5286 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5294 ) );
  MUX \Reg_Bank/U5368  ( .IN0(\Reg_Bank/n5292 ), .IN1(\Reg_Bank/n5289 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5293 ) );
  MUX \Reg_Bank/U5367  ( .IN0(\Reg_Bank/n5291 ), .IN1(\Reg_Bank/n5290 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5292 ) );
  MUX \Reg_Bank/U5366  ( .IN0(\Reg_Bank/registers[16][10] ), .IN1(
        \Reg_Bank/registers[17][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5291 )
         );
  MUX \Reg_Bank/U5365  ( .IN0(\Reg_Bank/registers[18][10] ), .IN1(
        \Reg_Bank/registers[19][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5290 )
         );
  MUX \Reg_Bank/U5364  ( .IN0(\Reg_Bank/n5288 ), .IN1(\Reg_Bank/n5287 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5289 ) );
  MUX \Reg_Bank/U5363  ( .IN0(\Reg_Bank/registers[20][10] ), .IN1(
        \Reg_Bank/registers[21][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5288 )
         );
  MUX \Reg_Bank/U5362  ( .IN0(\Reg_Bank/registers[22][10] ), .IN1(
        \Reg_Bank/registers[23][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5287 )
         );
  MUX \Reg_Bank/U5361  ( .IN0(\Reg_Bank/n5285 ), .IN1(\Reg_Bank/n5282 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5286 ) );
  MUX \Reg_Bank/U5360  ( .IN0(\Reg_Bank/n5284 ), .IN1(\Reg_Bank/n5283 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5285 ) );
  MUX \Reg_Bank/U5359  ( .IN0(\Reg_Bank/registers[24][10] ), .IN1(
        \Reg_Bank/registers[25][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5284 )
         );
  MUX \Reg_Bank/U5358  ( .IN0(\Reg_Bank/registers[26][10] ), .IN1(
        \Reg_Bank/registers[27][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5283 )
         );
  MUX \Reg_Bank/U5357  ( .IN0(\Reg_Bank/n5281 ), .IN1(\Reg_Bank/n5280 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5282 ) );
  MUX \Reg_Bank/U5356  ( .IN0(\Reg_Bank/registers[28][10] ), .IN1(
        \Reg_Bank/registers[29][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5281 )
         );
  MUX \Reg_Bank/U5355  ( .IN0(\Reg_Bank/registers[30][10] ), .IN1(
        \Reg_Bank/registers[31][10] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5280 )
         );
  MUX \Reg_Bank/U5354  ( .IN0(\Reg_Bank/n5279 ), .IN1(\Reg_Bank/n5264 ), .SEL(
        rt_index[4]), .F(reg_target[9]) );
  MUX \Reg_Bank/U5353  ( .IN0(\Reg_Bank/n5278 ), .IN1(\Reg_Bank/n5271 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5279 ) );
  MUX \Reg_Bank/U5352  ( .IN0(\Reg_Bank/n5277 ), .IN1(\Reg_Bank/n5274 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5278 ) );
  MUX \Reg_Bank/U5351  ( .IN0(\Reg_Bank/n5276 ), .IN1(\Reg_Bank/n5275 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5277 ) );
  MUX \Reg_Bank/U5349  ( .IN0(\Reg_Bank/registers[2][9] ), .IN1(
        \Reg_Bank/registers[3][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5275 )
         );
  MUX \Reg_Bank/U5348  ( .IN0(\Reg_Bank/n5273 ), .IN1(\Reg_Bank/n5272 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5274 ) );
  MUX \Reg_Bank/U5347  ( .IN0(\Reg_Bank/registers[4][9] ), .IN1(
        \Reg_Bank/registers[5][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5273 )
         );
  MUX \Reg_Bank/U5346  ( .IN0(\Reg_Bank/registers[6][9] ), .IN1(
        \Reg_Bank/registers[7][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5272 )
         );
  MUX \Reg_Bank/U5345  ( .IN0(\Reg_Bank/n5270 ), .IN1(\Reg_Bank/n5267 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5271 ) );
  MUX \Reg_Bank/U5344  ( .IN0(\Reg_Bank/n5269 ), .IN1(\Reg_Bank/n5268 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5270 ) );
  MUX \Reg_Bank/U5343  ( .IN0(\Reg_Bank/registers[8][9] ), .IN1(
        \Reg_Bank/registers[9][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5269 )
         );
  MUX \Reg_Bank/U5342  ( .IN0(\Reg_Bank/registers[10][9] ), .IN1(
        \Reg_Bank/registers[11][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5268 )
         );
  MUX \Reg_Bank/U5341  ( .IN0(\Reg_Bank/n5266 ), .IN1(\Reg_Bank/n5265 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5267 ) );
  MUX \Reg_Bank/U5340  ( .IN0(\Reg_Bank/registers[12][9] ), .IN1(
        \Reg_Bank/registers[13][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5266 )
         );
  MUX \Reg_Bank/U5339  ( .IN0(\Reg_Bank/registers[14][9] ), .IN1(
        \Reg_Bank/registers[15][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5265 )
         );
  MUX \Reg_Bank/U5338  ( .IN0(\Reg_Bank/n5263 ), .IN1(\Reg_Bank/n5256 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5264 ) );
  MUX \Reg_Bank/U5337  ( .IN0(\Reg_Bank/n5262 ), .IN1(\Reg_Bank/n5259 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5263 ) );
  MUX \Reg_Bank/U5336  ( .IN0(\Reg_Bank/n5261 ), .IN1(\Reg_Bank/n5260 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5262 ) );
  MUX \Reg_Bank/U5335  ( .IN0(\Reg_Bank/registers[16][9] ), .IN1(
        \Reg_Bank/registers[17][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5261 )
         );
  MUX \Reg_Bank/U5334  ( .IN0(\Reg_Bank/registers[18][9] ), .IN1(
        \Reg_Bank/registers[19][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5260 )
         );
  MUX \Reg_Bank/U5333  ( .IN0(\Reg_Bank/n5258 ), .IN1(\Reg_Bank/n5257 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5259 ) );
  MUX \Reg_Bank/U5332  ( .IN0(\Reg_Bank/registers[20][9] ), .IN1(
        \Reg_Bank/registers[21][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5258 )
         );
  MUX \Reg_Bank/U5331  ( .IN0(\Reg_Bank/registers[22][9] ), .IN1(
        \Reg_Bank/registers[23][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5257 )
         );
  MUX \Reg_Bank/U5330  ( .IN0(\Reg_Bank/n5255 ), .IN1(\Reg_Bank/n5252 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5256 ) );
  MUX \Reg_Bank/U5329  ( .IN0(\Reg_Bank/n5254 ), .IN1(\Reg_Bank/n5253 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5255 ) );
  MUX \Reg_Bank/U5328  ( .IN0(\Reg_Bank/registers[24][9] ), .IN1(
        \Reg_Bank/registers[25][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5254 )
         );
  MUX \Reg_Bank/U5327  ( .IN0(\Reg_Bank/registers[26][9] ), .IN1(
        \Reg_Bank/registers[27][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5253 )
         );
  MUX \Reg_Bank/U5326  ( .IN0(\Reg_Bank/n5251 ), .IN1(\Reg_Bank/n5250 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5252 ) );
  MUX \Reg_Bank/U5325  ( .IN0(\Reg_Bank/registers[28][9] ), .IN1(
        \Reg_Bank/registers[29][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5251 )
         );
  MUX \Reg_Bank/U5324  ( .IN0(\Reg_Bank/registers[30][9] ), .IN1(
        \Reg_Bank/registers[31][9] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5250 )
         );
  MUX \Reg_Bank/U5323  ( .IN0(\Reg_Bank/n5249 ), .IN1(\Reg_Bank/n5234 ), .SEL(
        rt_index[4]), .F(reg_target[8]) );
  MUX \Reg_Bank/U5322  ( .IN0(\Reg_Bank/n5248 ), .IN1(\Reg_Bank/n5241 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5249 ) );
  MUX \Reg_Bank/U5321  ( .IN0(\Reg_Bank/n5247 ), .IN1(\Reg_Bank/n5244 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5248 ) );
  MUX \Reg_Bank/U5320  ( .IN0(\Reg_Bank/n5246 ), .IN1(\Reg_Bank/n5245 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5247 ) );
  MUX \Reg_Bank/U5318  ( .IN0(\Reg_Bank/registers[2][8] ), .IN1(
        \Reg_Bank/registers[3][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5245 )
         );
  MUX \Reg_Bank/U5317  ( .IN0(\Reg_Bank/n5243 ), .IN1(\Reg_Bank/n5242 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5244 ) );
  MUX \Reg_Bank/U5316  ( .IN0(\Reg_Bank/registers[4][8] ), .IN1(
        \Reg_Bank/registers[5][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5243 )
         );
  MUX \Reg_Bank/U5315  ( .IN0(\Reg_Bank/registers[6][8] ), .IN1(
        \Reg_Bank/registers[7][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5242 )
         );
  MUX \Reg_Bank/U5314  ( .IN0(\Reg_Bank/n5240 ), .IN1(\Reg_Bank/n5237 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5241 ) );
  MUX \Reg_Bank/U5313  ( .IN0(\Reg_Bank/n5239 ), .IN1(\Reg_Bank/n5238 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5240 ) );
  MUX \Reg_Bank/U5312  ( .IN0(\Reg_Bank/registers[8][8] ), .IN1(
        \Reg_Bank/registers[9][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5239 )
         );
  MUX \Reg_Bank/U5311  ( .IN0(\Reg_Bank/registers[10][8] ), .IN1(
        \Reg_Bank/registers[11][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5238 )
         );
  MUX \Reg_Bank/U5310  ( .IN0(\Reg_Bank/n5236 ), .IN1(\Reg_Bank/n5235 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5237 ) );
  MUX \Reg_Bank/U5309  ( .IN0(\Reg_Bank/registers[12][8] ), .IN1(
        \Reg_Bank/registers[13][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5236 )
         );
  MUX \Reg_Bank/U5308  ( .IN0(\Reg_Bank/registers[14][8] ), .IN1(
        \Reg_Bank/registers[15][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5235 )
         );
  MUX \Reg_Bank/U5307  ( .IN0(\Reg_Bank/n5233 ), .IN1(\Reg_Bank/n5226 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5234 ) );
  MUX \Reg_Bank/U5306  ( .IN0(\Reg_Bank/n5232 ), .IN1(\Reg_Bank/n5229 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5233 ) );
  MUX \Reg_Bank/U5305  ( .IN0(\Reg_Bank/n5231 ), .IN1(\Reg_Bank/n5230 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5232 ) );
  MUX \Reg_Bank/U5304  ( .IN0(\Reg_Bank/registers[16][8] ), .IN1(
        \Reg_Bank/registers[17][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5231 )
         );
  MUX \Reg_Bank/U5303  ( .IN0(\Reg_Bank/registers[18][8] ), .IN1(
        \Reg_Bank/registers[19][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5230 )
         );
  MUX \Reg_Bank/U5302  ( .IN0(\Reg_Bank/n5228 ), .IN1(\Reg_Bank/n5227 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5229 ) );
  MUX \Reg_Bank/U5301  ( .IN0(\Reg_Bank/registers[20][8] ), .IN1(
        \Reg_Bank/registers[21][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5228 )
         );
  MUX \Reg_Bank/U5300  ( .IN0(\Reg_Bank/registers[22][8] ), .IN1(
        \Reg_Bank/registers[23][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5227 )
         );
  MUX \Reg_Bank/U5299  ( .IN0(\Reg_Bank/n5225 ), .IN1(\Reg_Bank/n5222 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5226 ) );
  MUX \Reg_Bank/U5298  ( .IN0(\Reg_Bank/n5224 ), .IN1(\Reg_Bank/n5223 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5225 ) );
  MUX \Reg_Bank/U5297  ( .IN0(\Reg_Bank/registers[24][8] ), .IN1(
        \Reg_Bank/registers[25][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5224 )
         );
  MUX \Reg_Bank/U5296  ( .IN0(\Reg_Bank/registers[26][8] ), .IN1(
        \Reg_Bank/registers[27][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5223 )
         );
  MUX \Reg_Bank/U5295  ( .IN0(\Reg_Bank/n5221 ), .IN1(\Reg_Bank/n5220 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5222 ) );
  MUX \Reg_Bank/U5294  ( .IN0(\Reg_Bank/registers[28][8] ), .IN1(
        \Reg_Bank/registers[29][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5221 )
         );
  MUX \Reg_Bank/U5293  ( .IN0(\Reg_Bank/registers[30][8] ), .IN1(
        \Reg_Bank/registers[31][8] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5220 )
         );
  MUX \Reg_Bank/U5292  ( .IN0(\Reg_Bank/n5219 ), .IN1(\Reg_Bank/n5204 ), .SEL(
        rt_index[4]), .F(reg_target[7]) );
  MUX \Reg_Bank/U5291  ( .IN0(\Reg_Bank/n5218 ), .IN1(\Reg_Bank/n5211 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5219 ) );
  MUX \Reg_Bank/U5290  ( .IN0(\Reg_Bank/n5217 ), .IN1(\Reg_Bank/n5214 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5218 ) );
  MUX \Reg_Bank/U5289  ( .IN0(\Reg_Bank/n5216 ), .IN1(\Reg_Bank/n5215 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5217 ) );
  MUX \Reg_Bank/U5287  ( .IN0(\Reg_Bank/registers[2][7] ), .IN1(
        \Reg_Bank/registers[3][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5215 )
         );
  MUX \Reg_Bank/U5286  ( .IN0(\Reg_Bank/n5213 ), .IN1(\Reg_Bank/n5212 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5214 ) );
  MUX \Reg_Bank/U5285  ( .IN0(\Reg_Bank/registers[4][7] ), .IN1(
        \Reg_Bank/registers[5][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5213 )
         );
  MUX \Reg_Bank/U5284  ( .IN0(\Reg_Bank/registers[6][7] ), .IN1(
        \Reg_Bank/registers[7][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5212 )
         );
  MUX \Reg_Bank/U5283  ( .IN0(\Reg_Bank/n5210 ), .IN1(\Reg_Bank/n5207 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5211 ) );
  MUX \Reg_Bank/U5282  ( .IN0(\Reg_Bank/n5209 ), .IN1(\Reg_Bank/n5208 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5210 ) );
  MUX \Reg_Bank/U5281  ( .IN0(\Reg_Bank/registers[8][7] ), .IN1(
        \Reg_Bank/registers[9][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5209 )
         );
  MUX \Reg_Bank/U5280  ( .IN0(\Reg_Bank/registers[10][7] ), .IN1(
        \Reg_Bank/registers[11][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5208 )
         );
  MUX \Reg_Bank/U5279  ( .IN0(\Reg_Bank/n5206 ), .IN1(\Reg_Bank/n5205 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5207 ) );
  MUX \Reg_Bank/U5278  ( .IN0(\Reg_Bank/registers[12][7] ), .IN1(
        \Reg_Bank/registers[13][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5206 )
         );
  MUX \Reg_Bank/U5277  ( .IN0(\Reg_Bank/registers[14][7] ), .IN1(
        \Reg_Bank/registers[15][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5205 )
         );
  MUX \Reg_Bank/U5276  ( .IN0(\Reg_Bank/n5203 ), .IN1(\Reg_Bank/n5196 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5204 ) );
  MUX \Reg_Bank/U5275  ( .IN0(\Reg_Bank/n5202 ), .IN1(\Reg_Bank/n5199 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5203 ) );
  MUX \Reg_Bank/U5274  ( .IN0(\Reg_Bank/n5201 ), .IN1(\Reg_Bank/n5200 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5202 ) );
  MUX \Reg_Bank/U5273  ( .IN0(\Reg_Bank/registers[16][7] ), .IN1(
        \Reg_Bank/registers[17][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5201 )
         );
  MUX \Reg_Bank/U5272  ( .IN0(\Reg_Bank/registers[18][7] ), .IN1(
        \Reg_Bank/registers[19][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5200 )
         );
  MUX \Reg_Bank/U5271  ( .IN0(\Reg_Bank/n5198 ), .IN1(\Reg_Bank/n5197 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5199 ) );
  MUX \Reg_Bank/U5270  ( .IN0(\Reg_Bank/registers[20][7] ), .IN1(
        \Reg_Bank/registers[21][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5198 )
         );
  MUX \Reg_Bank/U5269  ( .IN0(\Reg_Bank/registers[22][7] ), .IN1(
        \Reg_Bank/registers[23][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5197 )
         );
  MUX \Reg_Bank/U5268  ( .IN0(\Reg_Bank/n5195 ), .IN1(\Reg_Bank/n5192 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5196 ) );
  MUX \Reg_Bank/U5267  ( .IN0(\Reg_Bank/n5194 ), .IN1(\Reg_Bank/n5193 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5195 ) );
  MUX \Reg_Bank/U5266  ( .IN0(\Reg_Bank/registers[24][7] ), .IN1(
        \Reg_Bank/registers[25][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5194 )
         );
  MUX \Reg_Bank/U5265  ( .IN0(\Reg_Bank/registers[26][7] ), .IN1(
        \Reg_Bank/registers[27][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5193 )
         );
  MUX \Reg_Bank/U5264  ( .IN0(\Reg_Bank/n5191 ), .IN1(\Reg_Bank/n5190 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5192 ) );
  MUX \Reg_Bank/U5263  ( .IN0(\Reg_Bank/registers[28][7] ), .IN1(
        \Reg_Bank/registers[29][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5191 )
         );
  MUX \Reg_Bank/U5262  ( .IN0(\Reg_Bank/registers[30][7] ), .IN1(
        \Reg_Bank/registers[31][7] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5190 )
         );
  MUX \Reg_Bank/U5261  ( .IN0(\Reg_Bank/n5189 ), .IN1(\Reg_Bank/n5174 ), .SEL(
        rt_index[4]), .F(reg_target[6]) );
  MUX \Reg_Bank/U5260  ( .IN0(\Reg_Bank/n5188 ), .IN1(\Reg_Bank/n5181 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5189 ) );
  MUX \Reg_Bank/U5259  ( .IN0(\Reg_Bank/n5187 ), .IN1(\Reg_Bank/n5184 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5188 ) );
  MUX \Reg_Bank/U5258  ( .IN0(\Reg_Bank/n5186 ), .IN1(\Reg_Bank/n5185 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5187 ) );
  MUX \Reg_Bank/U5256  ( .IN0(\Reg_Bank/registers[2][6] ), .IN1(
        \Reg_Bank/registers[3][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5185 )
         );
  MUX \Reg_Bank/U5255  ( .IN0(\Reg_Bank/n5183 ), .IN1(\Reg_Bank/n5182 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5184 ) );
  MUX \Reg_Bank/U5254  ( .IN0(\Reg_Bank/registers[4][6] ), .IN1(
        \Reg_Bank/registers[5][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5183 )
         );
  MUX \Reg_Bank/U5253  ( .IN0(\Reg_Bank/registers[6][6] ), .IN1(
        \Reg_Bank/registers[7][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5182 )
         );
  MUX \Reg_Bank/U5252  ( .IN0(\Reg_Bank/n5180 ), .IN1(\Reg_Bank/n5177 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5181 ) );
  MUX \Reg_Bank/U5251  ( .IN0(\Reg_Bank/n5179 ), .IN1(\Reg_Bank/n5178 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5180 ) );
  MUX \Reg_Bank/U5250  ( .IN0(\Reg_Bank/registers[8][6] ), .IN1(
        \Reg_Bank/registers[9][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5179 )
         );
  MUX \Reg_Bank/U5249  ( .IN0(\Reg_Bank/registers[10][6] ), .IN1(
        \Reg_Bank/registers[11][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5178 )
         );
  MUX \Reg_Bank/U5248  ( .IN0(\Reg_Bank/n5176 ), .IN1(\Reg_Bank/n5175 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5177 ) );
  MUX \Reg_Bank/U5247  ( .IN0(\Reg_Bank/registers[12][6] ), .IN1(
        \Reg_Bank/registers[13][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5176 )
         );
  MUX \Reg_Bank/U5246  ( .IN0(\Reg_Bank/registers[14][6] ), .IN1(
        \Reg_Bank/registers[15][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5175 )
         );
  MUX \Reg_Bank/U5245  ( .IN0(\Reg_Bank/n5173 ), .IN1(\Reg_Bank/n5166 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5174 ) );
  MUX \Reg_Bank/U5244  ( .IN0(\Reg_Bank/n5172 ), .IN1(\Reg_Bank/n5169 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5173 ) );
  MUX \Reg_Bank/U5243  ( .IN0(\Reg_Bank/n5171 ), .IN1(\Reg_Bank/n5170 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5172 ) );
  MUX \Reg_Bank/U5242  ( .IN0(\Reg_Bank/registers[16][6] ), .IN1(
        \Reg_Bank/registers[17][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5171 )
         );
  MUX \Reg_Bank/U5241  ( .IN0(\Reg_Bank/registers[18][6] ), .IN1(
        \Reg_Bank/registers[19][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5170 )
         );
  MUX \Reg_Bank/U5240  ( .IN0(\Reg_Bank/n5168 ), .IN1(\Reg_Bank/n5167 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5169 ) );
  MUX \Reg_Bank/U5239  ( .IN0(\Reg_Bank/registers[20][6] ), .IN1(
        \Reg_Bank/registers[21][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5168 )
         );
  MUX \Reg_Bank/U5238  ( .IN0(\Reg_Bank/registers[22][6] ), .IN1(
        \Reg_Bank/registers[23][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5167 )
         );
  MUX \Reg_Bank/U5237  ( .IN0(\Reg_Bank/n5165 ), .IN1(\Reg_Bank/n5162 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5166 ) );
  MUX \Reg_Bank/U5236  ( .IN0(\Reg_Bank/n5164 ), .IN1(\Reg_Bank/n5163 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5165 ) );
  MUX \Reg_Bank/U5235  ( .IN0(\Reg_Bank/registers[24][6] ), .IN1(
        \Reg_Bank/registers[25][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5164 )
         );
  MUX \Reg_Bank/U5234  ( .IN0(\Reg_Bank/registers[26][6] ), .IN1(
        \Reg_Bank/registers[27][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5163 )
         );
  MUX \Reg_Bank/U5233  ( .IN0(\Reg_Bank/n5161 ), .IN1(\Reg_Bank/n5160 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5162 ) );
  MUX \Reg_Bank/U5232  ( .IN0(\Reg_Bank/registers[28][6] ), .IN1(
        \Reg_Bank/registers[29][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5161 )
         );
  MUX \Reg_Bank/U5231  ( .IN0(\Reg_Bank/registers[30][6] ), .IN1(
        \Reg_Bank/registers[31][6] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5160 )
         );
  MUX \Reg_Bank/U5230  ( .IN0(\Reg_Bank/n5159 ), .IN1(\Reg_Bank/n5144 ), .SEL(
        rt_index[4]), .F(reg_target[5]) );
  MUX \Reg_Bank/U5229  ( .IN0(\Reg_Bank/n5158 ), .IN1(\Reg_Bank/n5151 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5159 ) );
  MUX \Reg_Bank/U5228  ( .IN0(\Reg_Bank/n5157 ), .IN1(\Reg_Bank/n5154 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5158 ) );
  MUX \Reg_Bank/U5227  ( .IN0(\Reg_Bank/n5156 ), .IN1(\Reg_Bank/n5155 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5157 ) );
  MUX \Reg_Bank/U5225  ( .IN0(\Reg_Bank/registers[2][5] ), .IN1(
        \Reg_Bank/registers[3][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5155 )
         );
  MUX \Reg_Bank/U5224  ( .IN0(\Reg_Bank/n5153 ), .IN1(\Reg_Bank/n5152 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5154 ) );
  MUX \Reg_Bank/U5223  ( .IN0(\Reg_Bank/registers[4][5] ), .IN1(
        \Reg_Bank/registers[5][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5153 )
         );
  MUX \Reg_Bank/U5222  ( .IN0(\Reg_Bank/registers[6][5] ), .IN1(
        \Reg_Bank/registers[7][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5152 )
         );
  MUX \Reg_Bank/U5221  ( .IN0(\Reg_Bank/n5150 ), .IN1(\Reg_Bank/n5147 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5151 ) );
  MUX \Reg_Bank/U5220  ( .IN0(\Reg_Bank/n5149 ), .IN1(\Reg_Bank/n5148 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5150 ) );
  MUX \Reg_Bank/U5219  ( .IN0(\Reg_Bank/registers[8][5] ), .IN1(
        \Reg_Bank/registers[9][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5149 )
         );
  MUX \Reg_Bank/U5218  ( .IN0(\Reg_Bank/registers[10][5] ), .IN1(
        \Reg_Bank/registers[11][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5148 )
         );
  MUX \Reg_Bank/U5217  ( .IN0(\Reg_Bank/n5146 ), .IN1(\Reg_Bank/n5145 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5147 ) );
  MUX \Reg_Bank/U5216  ( .IN0(\Reg_Bank/registers[12][5] ), .IN1(
        \Reg_Bank/registers[13][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5146 )
         );
  MUX \Reg_Bank/U5215  ( .IN0(\Reg_Bank/registers[14][5] ), .IN1(
        \Reg_Bank/registers[15][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5145 )
         );
  MUX \Reg_Bank/U5214  ( .IN0(\Reg_Bank/n5143 ), .IN1(\Reg_Bank/n5136 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5144 ) );
  MUX \Reg_Bank/U5213  ( .IN0(\Reg_Bank/n5142 ), .IN1(\Reg_Bank/n5139 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5143 ) );
  MUX \Reg_Bank/U5212  ( .IN0(\Reg_Bank/n5141 ), .IN1(\Reg_Bank/n5140 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5142 ) );
  MUX \Reg_Bank/U5211  ( .IN0(\Reg_Bank/registers[16][5] ), .IN1(
        \Reg_Bank/registers[17][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5141 )
         );
  MUX \Reg_Bank/U5210  ( .IN0(\Reg_Bank/registers[18][5] ), .IN1(
        \Reg_Bank/registers[19][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5140 )
         );
  MUX \Reg_Bank/U5209  ( .IN0(\Reg_Bank/n5138 ), .IN1(\Reg_Bank/n5137 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5139 ) );
  MUX \Reg_Bank/U5208  ( .IN0(\Reg_Bank/registers[20][5] ), .IN1(
        \Reg_Bank/registers[21][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5138 )
         );
  MUX \Reg_Bank/U5207  ( .IN0(\Reg_Bank/registers[22][5] ), .IN1(
        \Reg_Bank/registers[23][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5137 )
         );
  MUX \Reg_Bank/U5206  ( .IN0(\Reg_Bank/n5135 ), .IN1(\Reg_Bank/n5132 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5136 ) );
  MUX \Reg_Bank/U5205  ( .IN0(\Reg_Bank/n5134 ), .IN1(\Reg_Bank/n5133 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5135 ) );
  MUX \Reg_Bank/U5204  ( .IN0(\Reg_Bank/registers[24][5] ), .IN1(
        \Reg_Bank/registers[25][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5134 )
         );
  MUX \Reg_Bank/U5203  ( .IN0(\Reg_Bank/registers[26][5] ), .IN1(
        \Reg_Bank/registers[27][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5133 )
         );
  MUX \Reg_Bank/U5202  ( .IN0(\Reg_Bank/n5131 ), .IN1(\Reg_Bank/n5130 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5132 ) );
  MUX \Reg_Bank/U5201  ( .IN0(\Reg_Bank/registers[28][5] ), .IN1(
        \Reg_Bank/registers[29][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5131 )
         );
  MUX \Reg_Bank/U5200  ( .IN0(\Reg_Bank/registers[30][5] ), .IN1(
        \Reg_Bank/registers[31][5] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5130 )
         );
  MUX \Reg_Bank/U5199  ( .IN0(\Reg_Bank/n5129 ), .IN1(\Reg_Bank/n5114 ), .SEL(
        rt_index[4]), .F(reg_target[4]) );
  MUX \Reg_Bank/U5198  ( .IN0(\Reg_Bank/n5128 ), .IN1(\Reg_Bank/n5121 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5129 ) );
  MUX \Reg_Bank/U5197  ( .IN0(\Reg_Bank/n5127 ), .IN1(\Reg_Bank/n5124 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5128 ) );
  MUX \Reg_Bank/U5196  ( .IN0(\Reg_Bank/n5126 ), .IN1(\Reg_Bank/n5125 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5127 ) );
  MUX \Reg_Bank/U5194  ( .IN0(\Reg_Bank/registers[2][4] ), .IN1(
        \Reg_Bank/registers[3][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5125 )
         );
  MUX \Reg_Bank/U5193  ( .IN0(\Reg_Bank/n5123 ), .IN1(\Reg_Bank/n5122 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5124 ) );
  MUX \Reg_Bank/U5192  ( .IN0(\Reg_Bank/registers[4][4] ), .IN1(
        \Reg_Bank/registers[5][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5123 )
         );
  MUX \Reg_Bank/U5191  ( .IN0(\Reg_Bank/registers[6][4] ), .IN1(
        \Reg_Bank/registers[7][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5122 )
         );
  MUX \Reg_Bank/U5190  ( .IN0(\Reg_Bank/n5120 ), .IN1(\Reg_Bank/n5117 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5121 ) );
  MUX \Reg_Bank/U5189  ( .IN0(\Reg_Bank/n5119 ), .IN1(\Reg_Bank/n5118 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5120 ) );
  MUX \Reg_Bank/U5188  ( .IN0(\Reg_Bank/registers[8][4] ), .IN1(
        \Reg_Bank/registers[9][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5119 )
         );
  MUX \Reg_Bank/U5187  ( .IN0(\Reg_Bank/registers[10][4] ), .IN1(
        \Reg_Bank/registers[11][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5118 )
         );
  MUX \Reg_Bank/U5186  ( .IN0(\Reg_Bank/n5116 ), .IN1(\Reg_Bank/n5115 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5117 ) );
  MUX \Reg_Bank/U5185  ( .IN0(\Reg_Bank/registers[12][4] ), .IN1(
        \Reg_Bank/registers[13][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5116 )
         );
  MUX \Reg_Bank/U5184  ( .IN0(\Reg_Bank/registers[14][4] ), .IN1(
        \Reg_Bank/registers[15][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5115 )
         );
  MUX \Reg_Bank/U5183  ( .IN0(\Reg_Bank/n5113 ), .IN1(\Reg_Bank/n5106 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5114 ) );
  MUX \Reg_Bank/U5182  ( .IN0(\Reg_Bank/n5112 ), .IN1(\Reg_Bank/n5109 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5113 ) );
  MUX \Reg_Bank/U5181  ( .IN0(\Reg_Bank/n5111 ), .IN1(\Reg_Bank/n5110 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5112 ) );
  MUX \Reg_Bank/U5180  ( .IN0(\Reg_Bank/registers[16][4] ), .IN1(
        \Reg_Bank/registers[17][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5111 )
         );
  MUX \Reg_Bank/U5179  ( .IN0(\Reg_Bank/registers[18][4] ), .IN1(
        \Reg_Bank/registers[19][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5110 )
         );
  MUX \Reg_Bank/U5178  ( .IN0(\Reg_Bank/n5108 ), .IN1(\Reg_Bank/n5107 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5109 ) );
  MUX \Reg_Bank/U5177  ( .IN0(\Reg_Bank/registers[20][4] ), .IN1(
        \Reg_Bank/registers[21][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5108 )
         );
  MUX \Reg_Bank/U5176  ( .IN0(\Reg_Bank/registers[22][4] ), .IN1(
        \Reg_Bank/registers[23][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5107 )
         );
  MUX \Reg_Bank/U5175  ( .IN0(\Reg_Bank/n5105 ), .IN1(\Reg_Bank/n5102 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5106 ) );
  MUX \Reg_Bank/U5174  ( .IN0(\Reg_Bank/n5104 ), .IN1(\Reg_Bank/n5103 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5105 ) );
  MUX \Reg_Bank/U5173  ( .IN0(\Reg_Bank/registers[24][4] ), .IN1(
        \Reg_Bank/registers[25][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5104 )
         );
  MUX \Reg_Bank/U5172  ( .IN0(\Reg_Bank/registers[26][4] ), .IN1(
        \Reg_Bank/registers[27][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5103 )
         );
  MUX \Reg_Bank/U5171  ( .IN0(\Reg_Bank/n5101 ), .IN1(\Reg_Bank/n5100 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5102 ) );
  MUX \Reg_Bank/U5170  ( .IN0(\Reg_Bank/registers[28][4] ), .IN1(
        \Reg_Bank/registers[29][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5101 )
         );
  MUX \Reg_Bank/U5169  ( .IN0(\Reg_Bank/registers[30][4] ), .IN1(
        \Reg_Bank/registers[31][4] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5100 )
         );
  MUX \Reg_Bank/U5168  ( .IN0(\Reg_Bank/n5099 ), .IN1(\Reg_Bank/n5084 ), .SEL(
        rt_index[4]), .F(reg_target[3]) );
  MUX \Reg_Bank/U5167  ( .IN0(\Reg_Bank/n5098 ), .IN1(\Reg_Bank/n5091 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5099 ) );
  MUX \Reg_Bank/U5166  ( .IN0(\Reg_Bank/n5097 ), .IN1(\Reg_Bank/n5094 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5098 ) );
  MUX \Reg_Bank/U5165  ( .IN0(\Reg_Bank/n5096 ), .IN1(\Reg_Bank/n5095 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5097 ) );
  MUX \Reg_Bank/U5163  ( .IN0(\Reg_Bank/registers[2][3] ), .IN1(
        \Reg_Bank/registers[3][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5095 )
         );
  MUX \Reg_Bank/U5162  ( .IN0(\Reg_Bank/n5093 ), .IN1(\Reg_Bank/n5092 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5094 ) );
  MUX \Reg_Bank/U5161  ( .IN0(\Reg_Bank/registers[4][3] ), .IN1(
        \Reg_Bank/registers[5][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5093 )
         );
  MUX \Reg_Bank/U5160  ( .IN0(\Reg_Bank/registers[6][3] ), .IN1(
        \Reg_Bank/registers[7][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5092 )
         );
  MUX \Reg_Bank/U5159  ( .IN0(\Reg_Bank/n5090 ), .IN1(\Reg_Bank/n5087 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5091 ) );
  MUX \Reg_Bank/U5158  ( .IN0(\Reg_Bank/n5089 ), .IN1(\Reg_Bank/n5088 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5090 ) );
  MUX \Reg_Bank/U5157  ( .IN0(\Reg_Bank/registers[8][3] ), .IN1(
        \Reg_Bank/registers[9][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5089 )
         );
  MUX \Reg_Bank/U5156  ( .IN0(\Reg_Bank/registers[10][3] ), .IN1(
        \Reg_Bank/registers[11][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5088 )
         );
  MUX \Reg_Bank/U5155  ( .IN0(\Reg_Bank/n5086 ), .IN1(\Reg_Bank/n5085 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5087 ) );
  MUX \Reg_Bank/U5154  ( .IN0(\Reg_Bank/registers[12][3] ), .IN1(
        \Reg_Bank/registers[13][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5086 )
         );
  MUX \Reg_Bank/U5153  ( .IN0(\Reg_Bank/registers[14][3] ), .IN1(
        \Reg_Bank/registers[15][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5085 )
         );
  MUX \Reg_Bank/U5152  ( .IN0(\Reg_Bank/n5083 ), .IN1(\Reg_Bank/n5076 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5084 ) );
  MUX \Reg_Bank/U5151  ( .IN0(\Reg_Bank/n5082 ), .IN1(\Reg_Bank/n5079 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5083 ) );
  MUX \Reg_Bank/U5150  ( .IN0(\Reg_Bank/n5081 ), .IN1(\Reg_Bank/n5080 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5082 ) );
  MUX \Reg_Bank/U5149  ( .IN0(\Reg_Bank/registers[16][3] ), .IN1(
        \Reg_Bank/registers[17][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5081 )
         );
  MUX \Reg_Bank/U5148  ( .IN0(\Reg_Bank/registers[18][3] ), .IN1(
        \Reg_Bank/registers[19][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5080 )
         );
  MUX \Reg_Bank/U5147  ( .IN0(\Reg_Bank/n5078 ), .IN1(\Reg_Bank/n5077 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5079 ) );
  MUX \Reg_Bank/U5146  ( .IN0(\Reg_Bank/registers[20][3] ), .IN1(
        \Reg_Bank/registers[21][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5078 )
         );
  MUX \Reg_Bank/U5145  ( .IN0(\Reg_Bank/registers[22][3] ), .IN1(
        \Reg_Bank/registers[23][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5077 )
         );
  MUX \Reg_Bank/U5144  ( .IN0(\Reg_Bank/n5075 ), .IN1(\Reg_Bank/n5072 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5076 ) );
  MUX \Reg_Bank/U5143  ( .IN0(\Reg_Bank/n5074 ), .IN1(\Reg_Bank/n5073 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5075 ) );
  MUX \Reg_Bank/U5142  ( .IN0(\Reg_Bank/registers[24][3] ), .IN1(
        \Reg_Bank/registers[25][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5074 )
         );
  MUX \Reg_Bank/U5141  ( .IN0(\Reg_Bank/registers[26][3] ), .IN1(
        \Reg_Bank/registers[27][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5073 )
         );
  MUX \Reg_Bank/U5140  ( .IN0(\Reg_Bank/n5071 ), .IN1(\Reg_Bank/n5070 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5072 ) );
  MUX \Reg_Bank/U5139  ( .IN0(\Reg_Bank/registers[28][3] ), .IN1(
        \Reg_Bank/registers[29][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5071 )
         );
  MUX \Reg_Bank/U5138  ( .IN0(\Reg_Bank/registers[30][3] ), .IN1(
        \Reg_Bank/registers[31][3] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5070 )
         );
  MUX \Reg_Bank/U5137  ( .IN0(\Reg_Bank/n5069 ), .IN1(\Reg_Bank/n5054 ), .SEL(
        rt_index[4]), .F(reg_target[2]) );
  MUX \Reg_Bank/U5136  ( .IN0(\Reg_Bank/n5068 ), .IN1(\Reg_Bank/n5061 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5069 ) );
  MUX \Reg_Bank/U5135  ( .IN0(\Reg_Bank/n5067 ), .IN1(\Reg_Bank/n5064 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5068 ) );
  MUX \Reg_Bank/U5134  ( .IN0(\Reg_Bank/n5066 ), .IN1(\Reg_Bank/n5065 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5067 ) );
  MUX \Reg_Bank/U5132  ( .IN0(\Reg_Bank/registers[2][2] ), .IN1(
        \Reg_Bank/registers[3][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5065 )
         );
  MUX \Reg_Bank/U5131  ( .IN0(\Reg_Bank/n5063 ), .IN1(\Reg_Bank/n5062 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5064 ) );
  MUX \Reg_Bank/U5130  ( .IN0(\Reg_Bank/registers[4][2] ), .IN1(
        \Reg_Bank/registers[5][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5063 )
         );
  MUX \Reg_Bank/U5129  ( .IN0(\Reg_Bank/registers[6][2] ), .IN1(
        \Reg_Bank/registers[7][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5062 )
         );
  MUX \Reg_Bank/U5128  ( .IN0(\Reg_Bank/n5060 ), .IN1(\Reg_Bank/n5057 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5061 ) );
  MUX \Reg_Bank/U5127  ( .IN0(\Reg_Bank/n5059 ), .IN1(\Reg_Bank/n5058 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5060 ) );
  MUX \Reg_Bank/U5126  ( .IN0(\Reg_Bank/registers[8][2] ), .IN1(
        \Reg_Bank/registers[9][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5059 )
         );
  MUX \Reg_Bank/U5125  ( .IN0(\Reg_Bank/registers[10][2] ), .IN1(
        \Reg_Bank/registers[11][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5058 )
         );
  MUX \Reg_Bank/U5124  ( .IN0(\Reg_Bank/n5056 ), .IN1(\Reg_Bank/n5055 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5057 ) );
  MUX \Reg_Bank/U5123  ( .IN0(\Reg_Bank/registers[12][2] ), .IN1(
        \Reg_Bank/registers[13][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5056 )
         );
  MUX \Reg_Bank/U5122  ( .IN0(\Reg_Bank/registers[14][2] ), .IN1(
        \Reg_Bank/registers[15][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5055 )
         );
  MUX \Reg_Bank/U5121  ( .IN0(\Reg_Bank/n5053 ), .IN1(\Reg_Bank/n5046 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5054 ) );
  MUX \Reg_Bank/U5120  ( .IN0(\Reg_Bank/n5052 ), .IN1(\Reg_Bank/n5049 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5053 ) );
  MUX \Reg_Bank/U5119  ( .IN0(\Reg_Bank/n5051 ), .IN1(\Reg_Bank/n5050 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5052 ) );
  MUX \Reg_Bank/U5118  ( .IN0(\Reg_Bank/registers[16][2] ), .IN1(
        \Reg_Bank/registers[17][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5051 )
         );
  MUX \Reg_Bank/U5117  ( .IN0(\Reg_Bank/registers[18][2] ), .IN1(
        \Reg_Bank/registers[19][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5050 )
         );
  MUX \Reg_Bank/U5116  ( .IN0(\Reg_Bank/n5048 ), .IN1(\Reg_Bank/n5047 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5049 ) );
  MUX \Reg_Bank/U5115  ( .IN0(\Reg_Bank/registers[20][2] ), .IN1(
        \Reg_Bank/registers[21][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5048 )
         );
  MUX \Reg_Bank/U5114  ( .IN0(\Reg_Bank/registers[22][2] ), .IN1(
        \Reg_Bank/registers[23][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5047 )
         );
  MUX \Reg_Bank/U5113  ( .IN0(\Reg_Bank/n5045 ), .IN1(\Reg_Bank/n5042 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5046 ) );
  MUX \Reg_Bank/U5112  ( .IN0(\Reg_Bank/n5044 ), .IN1(\Reg_Bank/n5043 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5045 ) );
  MUX \Reg_Bank/U5111  ( .IN0(\Reg_Bank/registers[24][2] ), .IN1(
        \Reg_Bank/registers[25][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5044 )
         );
  MUX \Reg_Bank/U5110  ( .IN0(\Reg_Bank/registers[26][2] ), .IN1(
        \Reg_Bank/registers[27][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5043 )
         );
  MUX \Reg_Bank/U5109  ( .IN0(\Reg_Bank/n5041 ), .IN1(\Reg_Bank/n5040 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5042 ) );
  MUX \Reg_Bank/U5108  ( .IN0(\Reg_Bank/registers[28][2] ), .IN1(
        \Reg_Bank/registers[29][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5041 )
         );
  MUX \Reg_Bank/U5107  ( .IN0(\Reg_Bank/registers[30][2] ), .IN1(
        \Reg_Bank/registers[31][2] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5040 )
         );
  MUX \Reg_Bank/U5106  ( .IN0(\Reg_Bank/n5039 ), .IN1(\Reg_Bank/n5024 ), .SEL(
        rt_index[4]), .F(reg_target[1]) );
  MUX \Reg_Bank/U5105  ( .IN0(\Reg_Bank/n5038 ), .IN1(\Reg_Bank/n5031 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5039 ) );
  MUX \Reg_Bank/U5104  ( .IN0(\Reg_Bank/n5037 ), .IN1(\Reg_Bank/n5034 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5038 ) );
  MUX \Reg_Bank/U5103  ( .IN0(\Reg_Bank/n5036 ), .IN1(\Reg_Bank/n5035 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5037 ) );
  MUX \Reg_Bank/U5101  ( .IN0(\Reg_Bank/registers[2][1] ), .IN1(
        \Reg_Bank/registers[3][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5035 )
         );
  MUX \Reg_Bank/U5100  ( .IN0(\Reg_Bank/n5033 ), .IN1(\Reg_Bank/n5032 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5034 ) );
  MUX \Reg_Bank/U5099  ( .IN0(\Reg_Bank/registers[4][1] ), .IN1(
        \Reg_Bank/registers[5][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5033 )
         );
  MUX \Reg_Bank/U5098  ( .IN0(\Reg_Bank/registers[6][1] ), .IN1(
        \Reg_Bank/registers[7][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5032 )
         );
  MUX \Reg_Bank/U5097  ( .IN0(\Reg_Bank/n5030 ), .IN1(\Reg_Bank/n5027 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5031 ) );
  MUX \Reg_Bank/U5096  ( .IN0(\Reg_Bank/n5029 ), .IN1(\Reg_Bank/n5028 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5030 ) );
  MUX \Reg_Bank/U5095  ( .IN0(\Reg_Bank/registers[8][1] ), .IN1(
        \Reg_Bank/registers[9][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5029 )
         );
  MUX \Reg_Bank/U5094  ( .IN0(\Reg_Bank/registers[10][1] ), .IN1(
        \Reg_Bank/registers[11][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5028 )
         );
  MUX \Reg_Bank/U5093  ( .IN0(\Reg_Bank/n5026 ), .IN1(\Reg_Bank/n5025 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5027 ) );
  MUX \Reg_Bank/U5092  ( .IN0(\Reg_Bank/registers[12][1] ), .IN1(
        \Reg_Bank/registers[13][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5026 )
         );
  MUX \Reg_Bank/U5091  ( .IN0(\Reg_Bank/registers[14][1] ), .IN1(
        \Reg_Bank/registers[15][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5025 )
         );
  MUX \Reg_Bank/U5090  ( .IN0(\Reg_Bank/n5023 ), .IN1(\Reg_Bank/n5016 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5024 ) );
  MUX \Reg_Bank/U5089  ( .IN0(\Reg_Bank/n5022 ), .IN1(\Reg_Bank/n5019 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5023 ) );
  MUX \Reg_Bank/U5088  ( .IN0(\Reg_Bank/n5021 ), .IN1(\Reg_Bank/n5020 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5022 ) );
  MUX \Reg_Bank/U5087  ( .IN0(\Reg_Bank/registers[16][1] ), .IN1(
        \Reg_Bank/registers[17][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5021 )
         );
  MUX \Reg_Bank/U5086  ( .IN0(\Reg_Bank/registers[18][1] ), .IN1(
        \Reg_Bank/registers[19][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5020 )
         );
  MUX \Reg_Bank/U5085  ( .IN0(\Reg_Bank/n5018 ), .IN1(\Reg_Bank/n5017 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5019 ) );
  MUX \Reg_Bank/U5084  ( .IN0(\Reg_Bank/registers[20][1] ), .IN1(
        \Reg_Bank/registers[21][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5018 )
         );
  MUX \Reg_Bank/U5083  ( .IN0(\Reg_Bank/registers[22][1] ), .IN1(
        \Reg_Bank/registers[23][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5017 )
         );
  MUX \Reg_Bank/U5082  ( .IN0(\Reg_Bank/n5015 ), .IN1(\Reg_Bank/n5012 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5016 ) );
  MUX \Reg_Bank/U5081  ( .IN0(\Reg_Bank/n5014 ), .IN1(\Reg_Bank/n5013 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5015 ) );
  MUX \Reg_Bank/U5080  ( .IN0(\Reg_Bank/registers[24][1] ), .IN1(
        \Reg_Bank/registers[25][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5014 )
         );
  MUX \Reg_Bank/U5079  ( .IN0(\Reg_Bank/registers[26][1] ), .IN1(
        \Reg_Bank/registers[27][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5013 )
         );
  MUX \Reg_Bank/U5078  ( .IN0(\Reg_Bank/n5011 ), .IN1(\Reg_Bank/n5010 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5012 ) );
  MUX \Reg_Bank/U5077  ( .IN0(\Reg_Bank/registers[28][1] ), .IN1(
        \Reg_Bank/registers[29][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5011 )
         );
  MUX \Reg_Bank/U5076  ( .IN0(\Reg_Bank/registers[30][1] ), .IN1(
        \Reg_Bank/registers[31][1] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5010 )
         );
  MUX \Reg_Bank/U5075  ( .IN0(\Reg_Bank/n5009 ), .IN1(\Reg_Bank/n4994 ), .SEL(
        rt_index[4]), .F(reg_target[0]) );
  MUX \Reg_Bank/U5074  ( .IN0(\Reg_Bank/n5008 ), .IN1(\Reg_Bank/n5001 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n5009 ) );
  MUX \Reg_Bank/U5073  ( .IN0(\Reg_Bank/n5007 ), .IN1(\Reg_Bank/n5004 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5008 ) );
  MUX \Reg_Bank/U5072  ( .IN0(\Reg_Bank/n5006 ), .IN1(\Reg_Bank/n5005 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5007 ) );
  MUX \Reg_Bank/U5070  ( .IN0(\Reg_Bank/registers[2][0] ), .IN1(
        \Reg_Bank/registers[3][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5005 )
         );
  MUX \Reg_Bank/U5069  ( .IN0(\Reg_Bank/n5003 ), .IN1(\Reg_Bank/n5002 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5004 ) );
  MUX \Reg_Bank/U5068  ( .IN0(\Reg_Bank/registers[4][0] ), .IN1(
        \Reg_Bank/registers[5][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5003 )
         );
  MUX \Reg_Bank/U5067  ( .IN0(\Reg_Bank/registers[6][0] ), .IN1(
        \Reg_Bank/registers[7][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n5002 )
         );
  MUX \Reg_Bank/U5066  ( .IN0(\Reg_Bank/n5000 ), .IN1(\Reg_Bank/n4997 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n5001 ) );
  MUX \Reg_Bank/U5065  ( .IN0(\Reg_Bank/n4999 ), .IN1(\Reg_Bank/n4998 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n5000 ) );
  MUX \Reg_Bank/U5064  ( .IN0(\Reg_Bank/registers[8][0] ), .IN1(
        \Reg_Bank/registers[9][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4999 )
         );
  MUX \Reg_Bank/U5063  ( .IN0(\Reg_Bank/registers[10][0] ), .IN1(
        \Reg_Bank/registers[11][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4998 )
         );
  MUX \Reg_Bank/U5062  ( .IN0(\Reg_Bank/n4996 ), .IN1(\Reg_Bank/n4995 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n4997 ) );
  MUX \Reg_Bank/U5061  ( .IN0(\Reg_Bank/registers[12][0] ), .IN1(
        \Reg_Bank/registers[13][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4996 )
         );
  MUX \Reg_Bank/U5060  ( .IN0(\Reg_Bank/registers[14][0] ), .IN1(
        \Reg_Bank/registers[15][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4995 )
         );
  MUX \Reg_Bank/U5059  ( .IN0(\Reg_Bank/n4993 ), .IN1(\Reg_Bank/n4986 ), .SEL(
        rt_index[3]), .F(\Reg_Bank/n4994 ) );
  MUX \Reg_Bank/U5058  ( .IN0(\Reg_Bank/n4992 ), .IN1(\Reg_Bank/n4989 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n4993 ) );
  MUX \Reg_Bank/U5057  ( .IN0(\Reg_Bank/n4991 ), .IN1(\Reg_Bank/n4990 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n4992 ) );
  MUX \Reg_Bank/U5056  ( .IN0(\Reg_Bank/registers[16][0] ), .IN1(
        \Reg_Bank/registers[17][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4991 )
         );
  MUX \Reg_Bank/U5055  ( .IN0(\Reg_Bank/registers[18][0] ), .IN1(
        \Reg_Bank/registers[19][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4990 )
         );
  MUX \Reg_Bank/U5054  ( .IN0(\Reg_Bank/n4988 ), .IN1(\Reg_Bank/n4987 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n4989 ) );
  MUX \Reg_Bank/U5053  ( .IN0(\Reg_Bank/registers[20][0] ), .IN1(
        \Reg_Bank/registers[21][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4988 )
         );
  MUX \Reg_Bank/U5052  ( .IN0(\Reg_Bank/registers[22][0] ), .IN1(
        \Reg_Bank/registers[23][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4987 )
         );
  MUX \Reg_Bank/U5051  ( .IN0(\Reg_Bank/n4985 ), .IN1(\Reg_Bank/n4982 ), .SEL(
        rt_index[2]), .F(\Reg_Bank/n4986 ) );
  MUX \Reg_Bank/U5050  ( .IN0(\Reg_Bank/n4984 ), .IN1(\Reg_Bank/n4983 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n4985 ) );
  MUX \Reg_Bank/U5049  ( .IN0(\Reg_Bank/registers[24][0] ), .IN1(
        \Reg_Bank/registers[25][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4984 )
         );
  MUX \Reg_Bank/U5048  ( .IN0(\Reg_Bank/registers[26][0] ), .IN1(
        \Reg_Bank/registers[27][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4983 )
         );
  MUX \Reg_Bank/U5047  ( .IN0(\Reg_Bank/n4981 ), .IN1(\Reg_Bank/n4980 ), .SEL(
        rt_index[1]), .F(\Reg_Bank/n4982 ) );
  MUX \Reg_Bank/U5046  ( .IN0(\Reg_Bank/registers[28][0] ), .IN1(
        \Reg_Bank/registers[29][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4981 )
         );
  MUX \Reg_Bank/U5045  ( .IN0(\Reg_Bank/registers[30][0] ), .IN1(
        \Reg_Bank/registers[31][0] ), .SEL(rt_index[0]), .F(\Reg_Bank/n4980 )
         );
  MUX \Reg_Bank/U5044  ( .IN0(\Reg_Bank/n4979 ), .IN1(\Reg_Bank/n4964 ), .SEL(
        rs_index[4]), .F(reg_source[31]) );
  MUX \Reg_Bank/U5043  ( .IN0(\Reg_Bank/n4978 ), .IN1(\Reg_Bank/n4971 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4979 ) );
  MUX \Reg_Bank/U5042  ( .IN0(\Reg_Bank/n4977 ), .IN1(\Reg_Bank/n4974 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4978 ) );
  MUX \Reg_Bank/U5041  ( .IN0(\Reg_Bank/n4976 ), .IN1(\Reg_Bank/n4975 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4977 ) );
  MUX \Reg_Bank/U5039  ( .IN0(\Reg_Bank/registers[2][31] ), .IN1(
        \Reg_Bank/registers[3][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4975 )
         );
  MUX \Reg_Bank/U5038  ( .IN0(\Reg_Bank/n4973 ), .IN1(\Reg_Bank/n4972 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4974 ) );
  MUX \Reg_Bank/U5037  ( .IN0(\Reg_Bank/registers[4][31] ), .IN1(
        \Reg_Bank/registers[5][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4973 )
         );
  MUX \Reg_Bank/U5036  ( .IN0(\Reg_Bank/registers[6][31] ), .IN1(
        \Reg_Bank/registers[7][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4972 )
         );
  MUX \Reg_Bank/U5035  ( .IN0(\Reg_Bank/n4970 ), .IN1(\Reg_Bank/n4967 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4971 ) );
  MUX \Reg_Bank/U5034  ( .IN0(\Reg_Bank/n4969 ), .IN1(\Reg_Bank/n4968 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4970 ) );
  MUX \Reg_Bank/U5033  ( .IN0(\Reg_Bank/registers[8][31] ), .IN1(
        \Reg_Bank/registers[9][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4969 )
         );
  MUX \Reg_Bank/U5032  ( .IN0(\Reg_Bank/registers[10][31] ), .IN1(
        \Reg_Bank/registers[11][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4968 )
         );
  MUX \Reg_Bank/U5031  ( .IN0(\Reg_Bank/n4966 ), .IN1(\Reg_Bank/n4965 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4967 ) );
  MUX \Reg_Bank/U5030  ( .IN0(\Reg_Bank/registers[12][31] ), .IN1(
        \Reg_Bank/registers[13][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4966 )
         );
  MUX \Reg_Bank/U5029  ( .IN0(\Reg_Bank/registers[14][31] ), .IN1(
        \Reg_Bank/registers[15][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4965 )
         );
  MUX \Reg_Bank/U5028  ( .IN0(\Reg_Bank/n4963 ), .IN1(\Reg_Bank/n4956 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4964 ) );
  MUX \Reg_Bank/U5027  ( .IN0(\Reg_Bank/n4962 ), .IN1(\Reg_Bank/n4959 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4963 ) );
  MUX \Reg_Bank/U5026  ( .IN0(\Reg_Bank/n4961 ), .IN1(\Reg_Bank/n4960 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4962 ) );
  MUX \Reg_Bank/U5025  ( .IN0(\Reg_Bank/registers[16][31] ), .IN1(
        \Reg_Bank/registers[17][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4961 )
         );
  MUX \Reg_Bank/U5024  ( .IN0(\Reg_Bank/registers[18][31] ), .IN1(
        \Reg_Bank/registers[19][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4960 )
         );
  MUX \Reg_Bank/U5023  ( .IN0(\Reg_Bank/n4958 ), .IN1(\Reg_Bank/n4957 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4959 ) );
  MUX \Reg_Bank/U5022  ( .IN0(\Reg_Bank/registers[20][31] ), .IN1(
        \Reg_Bank/registers[21][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4958 )
         );
  MUX \Reg_Bank/U5021  ( .IN0(\Reg_Bank/registers[22][31] ), .IN1(
        \Reg_Bank/registers[23][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4957 )
         );
  MUX \Reg_Bank/U5020  ( .IN0(\Reg_Bank/n4955 ), .IN1(\Reg_Bank/n4952 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4956 ) );
  MUX \Reg_Bank/U5019  ( .IN0(\Reg_Bank/n4954 ), .IN1(\Reg_Bank/n4953 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4955 ) );
  MUX \Reg_Bank/U5018  ( .IN0(\Reg_Bank/registers[24][31] ), .IN1(
        \Reg_Bank/registers[25][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4954 )
         );
  MUX \Reg_Bank/U5017  ( .IN0(\Reg_Bank/registers[26][31] ), .IN1(
        \Reg_Bank/registers[27][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4953 )
         );
  MUX \Reg_Bank/U5016  ( .IN0(\Reg_Bank/n4951 ), .IN1(\Reg_Bank/n4950 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4952 ) );
  MUX \Reg_Bank/U5015  ( .IN0(\Reg_Bank/registers[28][31] ), .IN1(
        \Reg_Bank/registers[29][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4951 )
         );
  MUX \Reg_Bank/U5014  ( .IN0(\Reg_Bank/registers[30][31] ), .IN1(
        \Reg_Bank/registers[31][31] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4950 )
         );
  MUX \Reg_Bank/U5013  ( .IN0(\Reg_Bank/n4949 ), .IN1(\Reg_Bank/n4934 ), .SEL(
        rs_index[4]), .F(reg_source[30]) );
  MUX \Reg_Bank/U5012  ( .IN0(\Reg_Bank/n4948 ), .IN1(\Reg_Bank/n4941 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4949 ) );
  MUX \Reg_Bank/U5011  ( .IN0(\Reg_Bank/n4947 ), .IN1(\Reg_Bank/n4944 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4948 ) );
  MUX \Reg_Bank/U5010  ( .IN0(\Reg_Bank/n4946 ), .IN1(\Reg_Bank/n4945 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4947 ) );
  MUX \Reg_Bank/U5008  ( .IN0(\Reg_Bank/registers[2][30] ), .IN1(
        \Reg_Bank/registers[3][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4945 )
         );
  MUX \Reg_Bank/U5007  ( .IN0(\Reg_Bank/n4943 ), .IN1(\Reg_Bank/n4942 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4944 ) );
  MUX \Reg_Bank/U5006  ( .IN0(\Reg_Bank/registers[4][30] ), .IN1(
        \Reg_Bank/registers[5][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4943 )
         );
  MUX \Reg_Bank/U5005  ( .IN0(\Reg_Bank/registers[6][30] ), .IN1(
        \Reg_Bank/registers[7][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4942 )
         );
  MUX \Reg_Bank/U5004  ( .IN0(\Reg_Bank/n4940 ), .IN1(\Reg_Bank/n4937 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4941 ) );
  MUX \Reg_Bank/U5003  ( .IN0(\Reg_Bank/n4939 ), .IN1(\Reg_Bank/n4938 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4940 ) );
  MUX \Reg_Bank/U5002  ( .IN0(\Reg_Bank/registers[8][30] ), .IN1(
        \Reg_Bank/registers[9][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4939 )
         );
  MUX \Reg_Bank/U5001  ( .IN0(\Reg_Bank/registers[10][30] ), .IN1(
        \Reg_Bank/registers[11][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4938 )
         );
  MUX \Reg_Bank/U5000  ( .IN0(\Reg_Bank/n4936 ), .IN1(\Reg_Bank/n4935 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4937 ) );
  MUX \Reg_Bank/U4999  ( .IN0(\Reg_Bank/registers[12][30] ), .IN1(
        \Reg_Bank/registers[13][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4936 )
         );
  MUX \Reg_Bank/U4998  ( .IN0(\Reg_Bank/registers[14][30] ), .IN1(
        \Reg_Bank/registers[15][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4935 )
         );
  MUX \Reg_Bank/U4997  ( .IN0(\Reg_Bank/n4933 ), .IN1(\Reg_Bank/n4926 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4934 ) );
  MUX \Reg_Bank/U4996  ( .IN0(\Reg_Bank/n4932 ), .IN1(\Reg_Bank/n4929 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4933 ) );
  MUX \Reg_Bank/U4995  ( .IN0(\Reg_Bank/n4931 ), .IN1(\Reg_Bank/n4930 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4932 ) );
  MUX \Reg_Bank/U4994  ( .IN0(\Reg_Bank/registers[16][30] ), .IN1(
        \Reg_Bank/registers[17][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4931 )
         );
  MUX \Reg_Bank/U4993  ( .IN0(\Reg_Bank/registers[18][30] ), .IN1(
        \Reg_Bank/registers[19][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4930 )
         );
  MUX \Reg_Bank/U4992  ( .IN0(\Reg_Bank/n4928 ), .IN1(\Reg_Bank/n4927 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4929 ) );
  MUX \Reg_Bank/U4991  ( .IN0(\Reg_Bank/registers[20][30] ), .IN1(
        \Reg_Bank/registers[21][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4928 )
         );
  MUX \Reg_Bank/U4990  ( .IN0(\Reg_Bank/registers[22][30] ), .IN1(
        \Reg_Bank/registers[23][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4927 )
         );
  MUX \Reg_Bank/U4989  ( .IN0(\Reg_Bank/n4925 ), .IN1(\Reg_Bank/n4922 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4926 ) );
  MUX \Reg_Bank/U4988  ( .IN0(\Reg_Bank/n4924 ), .IN1(\Reg_Bank/n4923 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4925 ) );
  MUX \Reg_Bank/U4987  ( .IN0(\Reg_Bank/registers[24][30] ), .IN1(
        \Reg_Bank/registers[25][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4924 )
         );
  MUX \Reg_Bank/U4986  ( .IN0(\Reg_Bank/registers[26][30] ), .IN1(
        \Reg_Bank/registers[27][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4923 )
         );
  MUX \Reg_Bank/U4985  ( .IN0(\Reg_Bank/n4921 ), .IN1(\Reg_Bank/n4920 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4922 ) );
  MUX \Reg_Bank/U4984  ( .IN0(\Reg_Bank/registers[28][30] ), .IN1(
        \Reg_Bank/registers[29][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4921 )
         );
  MUX \Reg_Bank/U4983  ( .IN0(\Reg_Bank/registers[30][30] ), .IN1(
        \Reg_Bank/registers[31][30] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4920 )
         );
  MUX \Reg_Bank/U4982  ( .IN0(\Reg_Bank/n4919 ), .IN1(\Reg_Bank/n4904 ), .SEL(
        rs_index[4]), .F(reg_source[29]) );
  MUX \Reg_Bank/U4981  ( .IN0(\Reg_Bank/n4918 ), .IN1(\Reg_Bank/n4911 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4919 ) );
  MUX \Reg_Bank/U4980  ( .IN0(\Reg_Bank/n4917 ), .IN1(\Reg_Bank/n4914 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4918 ) );
  MUX \Reg_Bank/U4979  ( .IN0(\Reg_Bank/n4916 ), .IN1(\Reg_Bank/n4915 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4917 ) );
  MUX \Reg_Bank/U4977  ( .IN0(\Reg_Bank/registers[2][29] ), .IN1(
        \Reg_Bank/registers[3][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4915 )
         );
  MUX \Reg_Bank/U4976  ( .IN0(\Reg_Bank/n4913 ), .IN1(\Reg_Bank/n4912 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4914 ) );
  MUX \Reg_Bank/U4975  ( .IN0(\Reg_Bank/registers[4][29] ), .IN1(
        \Reg_Bank/registers[5][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4913 )
         );
  MUX \Reg_Bank/U4974  ( .IN0(\Reg_Bank/registers[6][29] ), .IN1(
        \Reg_Bank/registers[7][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4912 )
         );
  MUX \Reg_Bank/U4973  ( .IN0(\Reg_Bank/n4910 ), .IN1(\Reg_Bank/n4907 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4911 ) );
  MUX \Reg_Bank/U4972  ( .IN0(\Reg_Bank/n4909 ), .IN1(\Reg_Bank/n4908 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4910 ) );
  MUX \Reg_Bank/U4971  ( .IN0(\Reg_Bank/registers[8][29] ), .IN1(
        \Reg_Bank/registers[9][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4909 )
         );
  MUX \Reg_Bank/U4970  ( .IN0(\Reg_Bank/registers[10][29] ), .IN1(
        \Reg_Bank/registers[11][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4908 )
         );
  MUX \Reg_Bank/U4969  ( .IN0(\Reg_Bank/n4906 ), .IN1(\Reg_Bank/n4905 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4907 ) );
  MUX \Reg_Bank/U4968  ( .IN0(\Reg_Bank/registers[12][29] ), .IN1(
        \Reg_Bank/registers[13][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4906 )
         );
  MUX \Reg_Bank/U4967  ( .IN0(\Reg_Bank/registers[14][29] ), .IN1(
        \Reg_Bank/registers[15][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4905 )
         );
  MUX \Reg_Bank/U4966  ( .IN0(\Reg_Bank/n4903 ), .IN1(\Reg_Bank/n4896 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4904 ) );
  MUX \Reg_Bank/U4965  ( .IN0(\Reg_Bank/n4902 ), .IN1(\Reg_Bank/n4899 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4903 ) );
  MUX \Reg_Bank/U4964  ( .IN0(\Reg_Bank/n4901 ), .IN1(\Reg_Bank/n4900 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4902 ) );
  MUX \Reg_Bank/U4963  ( .IN0(\Reg_Bank/registers[16][29] ), .IN1(
        \Reg_Bank/registers[17][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4901 )
         );
  MUX \Reg_Bank/U4962  ( .IN0(\Reg_Bank/registers[18][29] ), .IN1(
        \Reg_Bank/registers[19][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4900 )
         );
  MUX \Reg_Bank/U4961  ( .IN0(\Reg_Bank/n4898 ), .IN1(\Reg_Bank/n4897 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4899 ) );
  MUX \Reg_Bank/U4960  ( .IN0(\Reg_Bank/registers[20][29] ), .IN1(
        \Reg_Bank/registers[21][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4898 )
         );
  MUX \Reg_Bank/U4959  ( .IN0(\Reg_Bank/registers[22][29] ), .IN1(
        \Reg_Bank/registers[23][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4897 )
         );
  MUX \Reg_Bank/U4958  ( .IN0(\Reg_Bank/n4895 ), .IN1(\Reg_Bank/n4892 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4896 ) );
  MUX \Reg_Bank/U4957  ( .IN0(\Reg_Bank/n4894 ), .IN1(\Reg_Bank/n4893 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4895 ) );
  MUX \Reg_Bank/U4956  ( .IN0(\Reg_Bank/registers[24][29] ), .IN1(
        \Reg_Bank/registers[25][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4894 )
         );
  MUX \Reg_Bank/U4955  ( .IN0(\Reg_Bank/registers[26][29] ), .IN1(
        \Reg_Bank/registers[27][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4893 )
         );
  MUX \Reg_Bank/U4954  ( .IN0(\Reg_Bank/n4891 ), .IN1(\Reg_Bank/n4890 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4892 ) );
  MUX \Reg_Bank/U4953  ( .IN0(\Reg_Bank/registers[28][29] ), .IN1(
        \Reg_Bank/registers[29][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4891 )
         );
  MUX \Reg_Bank/U4952  ( .IN0(\Reg_Bank/registers[30][29] ), .IN1(
        \Reg_Bank/registers[31][29] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4890 )
         );
  MUX \Reg_Bank/U4951  ( .IN0(\Reg_Bank/n4889 ), .IN1(\Reg_Bank/n4874 ), .SEL(
        rs_index[4]), .F(reg_source[28]) );
  MUX \Reg_Bank/U4950  ( .IN0(\Reg_Bank/n4888 ), .IN1(\Reg_Bank/n4881 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4889 ) );
  MUX \Reg_Bank/U4949  ( .IN0(\Reg_Bank/n4887 ), .IN1(\Reg_Bank/n4884 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4888 ) );
  MUX \Reg_Bank/U4948  ( .IN0(\Reg_Bank/n4886 ), .IN1(\Reg_Bank/n4885 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4887 ) );
  MUX \Reg_Bank/U4946  ( .IN0(\Reg_Bank/registers[2][28] ), .IN1(
        \Reg_Bank/registers[3][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4885 )
         );
  MUX \Reg_Bank/U4945  ( .IN0(\Reg_Bank/n4883 ), .IN1(\Reg_Bank/n4882 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4884 ) );
  MUX \Reg_Bank/U4944  ( .IN0(\Reg_Bank/registers[4][28] ), .IN1(
        \Reg_Bank/registers[5][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4883 )
         );
  MUX \Reg_Bank/U4943  ( .IN0(\Reg_Bank/registers[6][28] ), .IN1(
        \Reg_Bank/registers[7][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4882 )
         );
  MUX \Reg_Bank/U4942  ( .IN0(\Reg_Bank/n4880 ), .IN1(\Reg_Bank/n4877 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4881 ) );
  MUX \Reg_Bank/U4941  ( .IN0(\Reg_Bank/n4879 ), .IN1(\Reg_Bank/n4878 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4880 ) );
  MUX \Reg_Bank/U4940  ( .IN0(\Reg_Bank/registers[8][28] ), .IN1(
        \Reg_Bank/registers[9][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4879 )
         );
  MUX \Reg_Bank/U4939  ( .IN0(\Reg_Bank/registers[10][28] ), .IN1(
        \Reg_Bank/registers[11][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4878 )
         );
  MUX \Reg_Bank/U4938  ( .IN0(\Reg_Bank/n4876 ), .IN1(\Reg_Bank/n4875 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4877 ) );
  MUX \Reg_Bank/U4937  ( .IN0(\Reg_Bank/registers[12][28] ), .IN1(
        \Reg_Bank/registers[13][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4876 )
         );
  MUX \Reg_Bank/U4936  ( .IN0(\Reg_Bank/registers[14][28] ), .IN1(
        \Reg_Bank/registers[15][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4875 )
         );
  MUX \Reg_Bank/U4935  ( .IN0(\Reg_Bank/n4873 ), .IN1(\Reg_Bank/n4866 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4874 ) );
  MUX \Reg_Bank/U4934  ( .IN0(\Reg_Bank/n4872 ), .IN1(\Reg_Bank/n4869 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4873 ) );
  MUX \Reg_Bank/U4933  ( .IN0(\Reg_Bank/n4871 ), .IN1(\Reg_Bank/n4870 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4872 ) );
  MUX \Reg_Bank/U4932  ( .IN0(\Reg_Bank/registers[16][28] ), .IN1(
        \Reg_Bank/registers[17][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4871 )
         );
  MUX \Reg_Bank/U4931  ( .IN0(\Reg_Bank/registers[18][28] ), .IN1(
        \Reg_Bank/registers[19][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4870 )
         );
  MUX \Reg_Bank/U4930  ( .IN0(\Reg_Bank/n4868 ), .IN1(\Reg_Bank/n4867 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4869 ) );
  MUX \Reg_Bank/U4929  ( .IN0(\Reg_Bank/registers[20][28] ), .IN1(
        \Reg_Bank/registers[21][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4868 )
         );
  MUX \Reg_Bank/U4928  ( .IN0(\Reg_Bank/registers[22][28] ), .IN1(
        \Reg_Bank/registers[23][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4867 )
         );
  MUX \Reg_Bank/U4927  ( .IN0(\Reg_Bank/n4865 ), .IN1(\Reg_Bank/n4862 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4866 ) );
  MUX \Reg_Bank/U4926  ( .IN0(\Reg_Bank/n4864 ), .IN1(\Reg_Bank/n4863 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4865 ) );
  MUX \Reg_Bank/U4925  ( .IN0(\Reg_Bank/registers[24][28] ), .IN1(
        \Reg_Bank/registers[25][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4864 )
         );
  MUX \Reg_Bank/U4924  ( .IN0(\Reg_Bank/registers[26][28] ), .IN1(
        \Reg_Bank/registers[27][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4863 )
         );
  MUX \Reg_Bank/U4923  ( .IN0(\Reg_Bank/n4861 ), .IN1(\Reg_Bank/n4860 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4862 ) );
  MUX \Reg_Bank/U4922  ( .IN0(\Reg_Bank/registers[28][28] ), .IN1(
        \Reg_Bank/registers[29][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4861 )
         );
  MUX \Reg_Bank/U4921  ( .IN0(\Reg_Bank/registers[30][28] ), .IN1(
        \Reg_Bank/registers[31][28] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4860 )
         );
  MUX \Reg_Bank/U4920  ( .IN0(\Reg_Bank/n4859 ), .IN1(\Reg_Bank/n4844 ), .SEL(
        rs_index[4]), .F(reg_source[27]) );
  MUX \Reg_Bank/U4919  ( .IN0(\Reg_Bank/n4858 ), .IN1(\Reg_Bank/n4851 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4859 ) );
  MUX \Reg_Bank/U4918  ( .IN0(\Reg_Bank/n4857 ), .IN1(\Reg_Bank/n4854 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4858 ) );
  MUX \Reg_Bank/U4917  ( .IN0(\Reg_Bank/n4856 ), .IN1(\Reg_Bank/n4855 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4857 ) );
  MUX \Reg_Bank/U4915  ( .IN0(\Reg_Bank/registers[2][27] ), .IN1(
        \Reg_Bank/registers[3][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4855 )
         );
  MUX \Reg_Bank/U4914  ( .IN0(\Reg_Bank/n4853 ), .IN1(\Reg_Bank/n4852 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4854 ) );
  MUX \Reg_Bank/U4913  ( .IN0(\Reg_Bank/registers[4][27] ), .IN1(
        \Reg_Bank/registers[5][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4853 )
         );
  MUX \Reg_Bank/U4912  ( .IN0(\Reg_Bank/registers[6][27] ), .IN1(
        \Reg_Bank/registers[7][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4852 )
         );
  MUX \Reg_Bank/U4911  ( .IN0(\Reg_Bank/n4850 ), .IN1(\Reg_Bank/n4847 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4851 ) );
  MUX \Reg_Bank/U4910  ( .IN0(\Reg_Bank/n4849 ), .IN1(\Reg_Bank/n4848 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4850 ) );
  MUX \Reg_Bank/U4909  ( .IN0(\Reg_Bank/registers[8][27] ), .IN1(
        \Reg_Bank/registers[9][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4849 )
         );
  MUX \Reg_Bank/U4908  ( .IN0(\Reg_Bank/registers[10][27] ), .IN1(
        \Reg_Bank/registers[11][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4848 )
         );
  MUX \Reg_Bank/U4907  ( .IN0(\Reg_Bank/n4846 ), .IN1(\Reg_Bank/n4845 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4847 ) );
  MUX \Reg_Bank/U4906  ( .IN0(\Reg_Bank/registers[12][27] ), .IN1(
        \Reg_Bank/registers[13][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4846 )
         );
  MUX \Reg_Bank/U4905  ( .IN0(\Reg_Bank/registers[14][27] ), .IN1(
        \Reg_Bank/registers[15][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4845 )
         );
  MUX \Reg_Bank/U4904  ( .IN0(\Reg_Bank/n4843 ), .IN1(\Reg_Bank/n4836 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4844 ) );
  MUX \Reg_Bank/U4903  ( .IN0(\Reg_Bank/n4842 ), .IN1(\Reg_Bank/n4839 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4843 ) );
  MUX \Reg_Bank/U4902  ( .IN0(\Reg_Bank/n4841 ), .IN1(\Reg_Bank/n4840 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4842 ) );
  MUX \Reg_Bank/U4901  ( .IN0(\Reg_Bank/registers[16][27] ), .IN1(
        \Reg_Bank/registers[17][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4841 )
         );
  MUX \Reg_Bank/U4900  ( .IN0(\Reg_Bank/registers[18][27] ), .IN1(
        \Reg_Bank/registers[19][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4840 )
         );
  MUX \Reg_Bank/U4899  ( .IN0(\Reg_Bank/n4838 ), .IN1(\Reg_Bank/n4837 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4839 ) );
  MUX \Reg_Bank/U4898  ( .IN0(\Reg_Bank/registers[20][27] ), .IN1(
        \Reg_Bank/registers[21][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4838 )
         );
  MUX \Reg_Bank/U4897  ( .IN0(\Reg_Bank/registers[22][27] ), .IN1(
        \Reg_Bank/registers[23][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4837 )
         );
  MUX \Reg_Bank/U4896  ( .IN0(\Reg_Bank/n4835 ), .IN1(\Reg_Bank/n4832 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4836 ) );
  MUX \Reg_Bank/U4895  ( .IN0(\Reg_Bank/n4834 ), .IN1(\Reg_Bank/n4833 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4835 ) );
  MUX \Reg_Bank/U4894  ( .IN0(\Reg_Bank/registers[24][27] ), .IN1(
        \Reg_Bank/registers[25][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4834 )
         );
  MUX \Reg_Bank/U4893  ( .IN0(\Reg_Bank/registers[26][27] ), .IN1(
        \Reg_Bank/registers[27][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4833 )
         );
  MUX \Reg_Bank/U4892  ( .IN0(\Reg_Bank/n4831 ), .IN1(\Reg_Bank/n4830 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4832 ) );
  MUX \Reg_Bank/U4891  ( .IN0(\Reg_Bank/registers[28][27] ), .IN1(
        \Reg_Bank/registers[29][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4831 )
         );
  MUX \Reg_Bank/U4890  ( .IN0(\Reg_Bank/registers[30][27] ), .IN1(
        \Reg_Bank/registers[31][27] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4830 )
         );
  MUX \Reg_Bank/U4889  ( .IN0(\Reg_Bank/n4829 ), .IN1(\Reg_Bank/n4814 ), .SEL(
        rs_index[4]), .F(reg_source[26]) );
  MUX \Reg_Bank/U4888  ( .IN0(\Reg_Bank/n4828 ), .IN1(\Reg_Bank/n4821 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4829 ) );
  MUX \Reg_Bank/U4887  ( .IN0(\Reg_Bank/n4827 ), .IN1(\Reg_Bank/n4824 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4828 ) );
  MUX \Reg_Bank/U4886  ( .IN0(\Reg_Bank/n4826 ), .IN1(\Reg_Bank/n4825 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4827 ) );
  MUX \Reg_Bank/U4884  ( .IN0(\Reg_Bank/registers[2][26] ), .IN1(
        \Reg_Bank/registers[3][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4825 )
         );
  MUX \Reg_Bank/U4883  ( .IN0(\Reg_Bank/n4823 ), .IN1(\Reg_Bank/n4822 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4824 ) );
  MUX \Reg_Bank/U4882  ( .IN0(\Reg_Bank/registers[4][26] ), .IN1(
        \Reg_Bank/registers[5][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4823 )
         );
  MUX \Reg_Bank/U4881  ( .IN0(\Reg_Bank/registers[6][26] ), .IN1(
        \Reg_Bank/registers[7][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4822 )
         );
  MUX \Reg_Bank/U4880  ( .IN0(\Reg_Bank/n4820 ), .IN1(\Reg_Bank/n4817 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4821 ) );
  MUX \Reg_Bank/U4879  ( .IN0(\Reg_Bank/n4819 ), .IN1(\Reg_Bank/n4818 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4820 ) );
  MUX \Reg_Bank/U4878  ( .IN0(\Reg_Bank/registers[8][26] ), .IN1(
        \Reg_Bank/registers[9][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4819 )
         );
  MUX \Reg_Bank/U4877  ( .IN0(\Reg_Bank/registers[10][26] ), .IN1(
        \Reg_Bank/registers[11][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4818 )
         );
  MUX \Reg_Bank/U4876  ( .IN0(\Reg_Bank/n4816 ), .IN1(\Reg_Bank/n4815 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4817 ) );
  MUX \Reg_Bank/U4875  ( .IN0(\Reg_Bank/registers[12][26] ), .IN1(
        \Reg_Bank/registers[13][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4816 )
         );
  MUX \Reg_Bank/U4874  ( .IN0(\Reg_Bank/registers[14][26] ), .IN1(
        \Reg_Bank/registers[15][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4815 )
         );
  MUX \Reg_Bank/U4873  ( .IN0(\Reg_Bank/n4813 ), .IN1(\Reg_Bank/n4806 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4814 ) );
  MUX \Reg_Bank/U4872  ( .IN0(\Reg_Bank/n4812 ), .IN1(\Reg_Bank/n4809 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4813 ) );
  MUX \Reg_Bank/U4871  ( .IN0(\Reg_Bank/n4811 ), .IN1(\Reg_Bank/n4810 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4812 ) );
  MUX \Reg_Bank/U4870  ( .IN0(\Reg_Bank/registers[16][26] ), .IN1(
        \Reg_Bank/registers[17][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4811 )
         );
  MUX \Reg_Bank/U4869  ( .IN0(\Reg_Bank/registers[18][26] ), .IN1(
        \Reg_Bank/registers[19][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4810 )
         );
  MUX \Reg_Bank/U4868  ( .IN0(\Reg_Bank/n4808 ), .IN1(\Reg_Bank/n4807 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4809 ) );
  MUX \Reg_Bank/U4867  ( .IN0(\Reg_Bank/registers[20][26] ), .IN1(
        \Reg_Bank/registers[21][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4808 )
         );
  MUX \Reg_Bank/U4866  ( .IN0(\Reg_Bank/registers[22][26] ), .IN1(
        \Reg_Bank/registers[23][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4807 )
         );
  MUX \Reg_Bank/U4865  ( .IN0(\Reg_Bank/n4805 ), .IN1(\Reg_Bank/n4802 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4806 ) );
  MUX \Reg_Bank/U4864  ( .IN0(\Reg_Bank/n4804 ), .IN1(\Reg_Bank/n4803 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4805 ) );
  MUX \Reg_Bank/U4863  ( .IN0(\Reg_Bank/registers[24][26] ), .IN1(
        \Reg_Bank/registers[25][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4804 )
         );
  MUX \Reg_Bank/U4862  ( .IN0(\Reg_Bank/registers[26][26] ), .IN1(
        \Reg_Bank/registers[27][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4803 )
         );
  MUX \Reg_Bank/U4861  ( .IN0(\Reg_Bank/n4801 ), .IN1(\Reg_Bank/n4800 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4802 ) );
  MUX \Reg_Bank/U4860  ( .IN0(\Reg_Bank/registers[28][26] ), .IN1(
        \Reg_Bank/registers[29][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4801 )
         );
  MUX \Reg_Bank/U4859  ( .IN0(\Reg_Bank/registers[30][26] ), .IN1(
        \Reg_Bank/registers[31][26] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4800 )
         );
  MUX \Reg_Bank/U4858  ( .IN0(\Reg_Bank/n4799 ), .IN1(\Reg_Bank/n4784 ), .SEL(
        rs_index[4]), .F(reg_source[25]) );
  MUX \Reg_Bank/U4857  ( .IN0(\Reg_Bank/n4798 ), .IN1(\Reg_Bank/n4791 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4799 ) );
  MUX \Reg_Bank/U4856  ( .IN0(\Reg_Bank/n4797 ), .IN1(\Reg_Bank/n4794 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4798 ) );
  MUX \Reg_Bank/U4855  ( .IN0(\Reg_Bank/n4796 ), .IN1(\Reg_Bank/n4795 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4797 ) );
  MUX \Reg_Bank/U4853  ( .IN0(\Reg_Bank/registers[2][25] ), .IN1(
        \Reg_Bank/registers[3][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4795 )
         );
  MUX \Reg_Bank/U4852  ( .IN0(\Reg_Bank/n4793 ), .IN1(\Reg_Bank/n4792 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4794 ) );
  MUX \Reg_Bank/U4851  ( .IN0(\Reg_Bank/registers[4][25] ), .IN1(
        \Reg_Bank/registers[5][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4793 )
         );
  MUX \Reg_Bank/U4850  ( .IN0(\Reg_Bank/registers[6][25] ), .IN1(
        \Reg_Bank/registers[7][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4792 )
         );
  MUX \Reg_Bank/U4849  ( .IN0(\Reg_Bank/n4790 ), .IN1(\Reg_Bank/n4787 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4791 ) );
  MUX \Reg_Bank/U4848  ( .IN0(\Reg_Bank/n4789 ), .IN1(\Reg_Bank/n4788 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4790 ) );
  MUX \Reg_Bank/U4847  ( .IN0(\Reg_Bank/registers[8][25] ), .IN1(
        \Reg_Bank/registers[9][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4789 )
         );
  MUX \Reg_Bank/U4846  ( .IN0(\Reg_Bank/registers[10][25] ), .IN1(
        \Reg_Bank/registers[11][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4788 )
         );
  MUX \Reg_Bank/U4845  ( .IN0(\Reg_Bank/n4786 ), .IN1(\Reg_Bank/n4785 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4787 ) );
  MUX \Reg_Bank/U4844  ( .IN0(\Reg_Bank/registers[12][25] ), .IN1(
        \Reg_Bank/registers[13][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4786 )
         );
  MUX \Reg_Bank/U4843  ( .IN0(\Reg_Bank/registers[14][25] ), .IN1(
        \Reg_Bank/registers[15][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4785 )
         );
  MUX \Reg_Bank/U4842  ( .IN0(\Reg_Bank/n4783 ), .IN1(\Reg_Bank/n4776 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4784 ) );
  MUX \Reg_Bank/U4841  ( .IN0(\Reg_Bank/n4782 ), .IN1(\Reg_Bank/n4779 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4783 ) );
  MUX \Reg_Bank/U4840  ( .IN0(\Reg_Bank/n4781 ), .IN1(\Reg_Bank/n4780 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4782 ) );
  MUX \Reg_Bank/U4839  ( .IN0(\Reg_Bank/registers[16][25] ), .IN1(
        \Reg_Bank/registers[17][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4781 )
         );
  MUX \Reg_Bank/U4838  ( .IN0(\Reg_Bank/registers[18][25] ), .IN1(
        \Reg_Bank/registers[19][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4780 )
         );
  MUX \Reg_Bank/U4837  ( .IN0(\Reg_Bank/n4778 ), .IN1(\Reg_Bank/n4777 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4779 ) );
  MUX \Reg_Bank/U4836  ( .IN0(\Reg_Bank/registers[20][25] ), .IN1(
        \Reg_Bank/registers[21][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4778 )
         );
  MUX \Reg_Bank/U4835  ( .IN0(\Reg_Bank/registers[22][25] ), .IN1(
        \Reg_Bank/registers[23][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4777 )
         );
  MUX \Reg_Bank/U4834  ( .IN0(\Reg_Bank/n4775 ), .IN1(\Reg_Bank/n4772 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4776 ) );
  MUX \Reg_Bank/U4833  ( .IN0(\Reg_Bank/n4774 ), .IN1(\Reg_Bank/n4773 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4775 ) );
  MUX \Reg_Bank/U4832  ( .IN0(\Reg_Bank/registers[24][25] ), .IN1(
        \Reg_Bank/registers[25][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4774 )
         );
  MUX \Reg_Bank/U4831  ( .IN0(\Reg_Bank/registers[26][25] ), .IN1(
        \Reg_Bank/registers[27][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4773 )
         );
  MUX \Reg_Bank/U4830  ( .IN0(\Reg_Bank/n4771 ), .IN1(\Reg_Bank/n4770 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4772 ) );
  MUX \Reg_Bank/U4829  ( .IN0(\Reg_Bank/registers[28][25] ), .IN1(
        \Reg_Bank/registers[29][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4771 )
         );
  MUX \Reg_Bank/U4828  ( .IN0(\Reg_Bank/registers[30][25] ), .IN1(
        \Reg_Bank/registers[31][25] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4770 )
         );
  MUX \Reg_Bank/U4827  ( .IN0(\Reg_Bank/n4769 ), .IN1(\Reg_Bank/n4754 ), .SEL(
        rs_index[4]), .F(reg_source[24]) );
  MUX \Reg_Bank/U4826  ( .IN0(\Reg_Bank/n4768 ), .IN1(\Reg_Bank/n4761 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4769 ) );
  MUX \Reg_Bank/U4825  ( .IN0(\Reg_Bank/n4767 ), .IN1(\Reg_Bank/n4764 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4768 ) );
  MUX \Reg_Bank/U4824  ( .IN0(\Reg_Bank/n4766 ), .IN1(\Reg_Bank/n4765 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4767 ) );
  MUX \Reg_Bank/U4822  ( .IN0(\Reg_Bank/registers[2][24] ), .IN1(
        \Reg_Bank/registers[3][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4765 )
         );
  MUX \Reg_Bank/U4821  ( .IN0(\Reg_Bank/n4763 ), .IN1(\Reg_Bank/n4762 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4764 ) );
  MUX \Reg_Bank/U4820  ( .IN0(\Reg_Bank/registers[4][24] ), .IN1(
        \Reg_Bank/registers[5][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4763 )
         );
  MUX \Reg_Bank/U4819  ( .IN0(\Reg_Bank/registers[6][24] ), .IN1(
        \Reg_Bank/registers[7][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4762 )
         );
  MUX \Reg_Bank/U4818  ( .IN0(\Reg_Bank/n4760 ), .IN1(\Reg_Bank/n4757 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4761 ) );
  MUX \Reg_Bank/U4817  ( .IN0(\Reg_Bank/n4759 ), .IN1(\Reg_Bank/n4758 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4760 ) );
  MUX \Reg_Bank/U4816  ( .IN0(\Reg_Bank/registers[8][24] ), .IN1(
        \Reg_Bank/registers[9][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4759 )
         );
  MUX \Reg_Bank/U4815  ( .IN0(\Reg_Bank/registers[10][24] ), .IN1(
        \Reg_Bank/registers[11][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4758 )
         );
  MUX \Reg_Bank/U4814  ( .IN0(\Reg_Bank/n4756 ), .IN1(\Reg_Bank/n4755 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4757 ) );
  MUX \Reg_Bank/U4813  ( .IN0(\Reg_Bank/registers[12][24] ), .IN1(
        \Reg_Bank/registers[13][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4756 )
         );
  MUX \Reg_Bank/U4812  ( .IN0(\Reg_Bank/registers[14][24] ), .IN1(
        \Reg_Bank/registers[15][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4755 )
         );
  MUX \Reg_Bank/U4811  ( .IN0(\Reg_Bank/n4753 ), .IN1(\Reg_Bank/n4746 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4754 ) );
  MUX \Reg_Bank/U4810  ( .IN0(\Reg_Bank/n4752 ), .IN1(\Reg_Bank/n4749 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4753 ) );
  MUX \Reg_Bank/U4809  ( .IN0(\Reg_Bank/n4751 ), .IN1(\Reg_Bank/n4750 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4752 ) );
  MUX \Reg_Bank/U4808  ( .IN0(\Reg_Bank/registers[16][24] ), .IN1(
        \Reg_Bank/registers[17][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4751 )
         );
  MUX \Reg_Bank/U4807  ( .IN0(\Reg_Bank/registers[18][24] ), .IN1(
        \Reg_Bank/registers[19][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4750 )
         );
  MUX \Reg_Bank/U4806  ( .IN0(\Reg_Bank/n4748 ), .IN1(\Reg_Bank/n4747 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4749 ) );
  MUX \Reg_Bank/U4805  ( .IN0(\Reg_Bank/registers[20][24] ), .IN1(
        \Reg_Bank/registers[21][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4748 )
         );
  MUX \Reg_Bank/U4804  ( .IN0(\Reg_Bank/registers[22][24] ), .IN1(
        \Reg_Bank/registers[23][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4747 )
         );
  MUX \Reg_Bank/U4803  ( .IN0(\Reg_Bank/n4745 ), .IN1(\Reg_Bank/n4742 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4746 ) );
  MUX \Reg_Bank/U4802  ( .IN0(\Reg_Bank/n4744 ), .IN1(\Reg_Bank/n4743 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4745 ) );
  MUX \Reg_Bank/U4801  ( .IN0(\Reg_Bank/registers[24][24] ), .IN1(
        \Reg_Bank/registers[25][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4744 )
         );
  MUX \Reg_Bank/U4800  ( .IN0(\Reg_Bank/registers[26][24] ), .IN1(
        \Reg_Bank/registers[27][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4743 )
         );
  MUX \Reg_Bank/U4799  ( .IN0(\Reg_Bank/n4741 ), .IN1(\Reg_Bank/n4740 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4742 ) );
  MUX \Reg_Bank/U4798  ( .IN0(\Reg_Bank/registers[28][24] ), .IN1(
        \Reg_Bank/registers[29][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4741 )
         );
  MUX \Reg_Bank/U4797  ( .IN0(\Reg_Bank/registers[30][24] ), .IN1(
        \Reg_Bank/registers[31][24] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4740 )
         );
  MUX \Reg_Bank/U4796  ( .IN0(\Reg_Bank/n4739 ), .IN1(\Reg_Bank/n4724 ), .SEL(
        rs_index[4]), .F(reg_source[23]) );
  MUX \Reg_Bank/U4795  ( .IN0(\Reg_Bank/n4738 ), .IN1(\Reg_Bank/n4731 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4739 ) );
  MUX \Reg_Bank/U4794  ( .IN0(\Reg_Bank/n4737 ), .IN1(\Reg_Bank/n4734 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4738 ) );
  MUX \Reg_Bank/U4793  ( .IN0(\Reg_Bank/n4736 ), .IN1(\Reg_Bank/n4735 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4737 ) );
  MUX \Reg_Bank/U4791  ( .IN0(\Reg_Bank/registers[2][23] ), .IN1(
        \Reg_Bank/registers[3][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4735 )
         );
  MUX \Reg_Bank/U4790  ( .IN0(\Reg_Bank/n4733 ), .IN1(\Reg_Bank/n4732 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4734 ) );
  MUX \Reg_Bank/U4789  ( .IN0(\Reg_Bank/registers[4][23] ), .IN1(
        \Reg_Bank/registers[5][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4733 )
         );
  MUX \Reg_Bank/U4788  ( .IN0(\Reg_Bank/registers[6][23] ), .IN1(
        \Reg_Bank/registers[7][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4732 )
         );
  MUX \Reg_Bank/U4787  ( .IN0(\Reg_Bank/n4730 ), .IN1(\Reg_Bank/n4727 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4731 ) );
  MUX \Reg_Bank/U4786  ( .IN0(\Reg_Bank/n4729 ), .IN1(\Reg_Bank/n4728 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4730 ) );
  MUX \Reg_Bank/U4785  ( .IN0(\Reg_Bank/registers[8][23] ), .IN1(
        \Reg_Bank/registers[9][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4729 )
         );
  MUX \Reg_Bank/U4784  ( .IN0(\Reg_Bank/registers[10][23] ), .IN1(
        \Reg_Bank/registers[11][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4728 )
         );
  MUX \Reg_Bank/U4783  ( .IN0(\Reg_Bank/n4726 ), .IN1(\Reg_Bank/n4725 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4727 ) );
  MUX \Reg_Bank/U4782  ( .IN0(\Reg_Bank/registers[12][23] ), .IN1(
        \Reg_Bank/registers[13][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4726 )
         );
  MUX \Reg_Bank/U4781  ( .IN0(\Reg_Bank/registers[14][23] ), .IN1(
        \Reg_Bank/registers[15][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4725 )
         );
  MUX \Reg_Bank/U4780  ( .IN0(\Reg_Bank/n4723 ), .IN1(\Reg_Bank/n4716 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4724 ) );
  MUX \Reg_Bank/U4779  ( .IN0(\Reg_Bank/n4722 ), .IN1(\Reg_Bank/n4719 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4723 ) );
  MUX \Reg_Bank/U4778  ( .IN0(\Reg_Bank/n4721 ), .IN1(\Reg_Bank/n4720 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4722 ) );
  MUX \Reg_Bank/U4777  ( .IN0(\Reg_Bank/registers[16][23] ), .IN1(
        \Reg_Bank/registers[17][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4721 )
         );
  MUX \Reg_Bank/U4776  ( .IN0(\Reg_Bank/registers[18][23] ), .IN1(
        \Reg_Bank/registers[19][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4720 )
         );
  MUX \Reg_Bank/U4775  ( .IN0(\Reg_Bank/n4718 ), .IN1(\Reg_Bank/n4717 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4719 ) );
  MUX \Reg_Bank/U4774  ( .IN0(\Reg_Bank/registers[20][23] ), .IN1(
        \Reg_Bank/registers[21][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4718 )
         );
  MUX \Reg_Bank/U4773  ( .IN0(\Reg_Bank/registers[22][23] ), .IN1(
        \Reg_Bank/registers[23][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4717 )
         );
  MUX \Reg_Bank/U4772  ( .IN0(\Reg_Bank/n4715 ), .IN1(\Reg_Bank/n4712 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4716 ) );
  MUX \Reg_Bank/U4771  ( .IN0(\Reg_Bank/n4714 ), .IN1(\Reg_Bank/n4713 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4715 ) );
  MUX \Reg_Bank/U4770  ( .IN0(\Reg_Bank/registers[24][23] ), .IN1(
        \Reg_Bank/registers[25][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4714 )
         );
  MUX \Reg_Bank/U4769  ( .IN0(\Reg_Bank/registers[26][23] ), .IN1(
        \Reg_Bank/registers[27][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4713 )
         );
  MUX \Reg_Bank/U4768  ( .IN0(\Reg_Bank/n4711 ), .IN1(\Reg_Bank/n4710 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4712 ) );
  MUX \Reg_Bank/U4767  ( .IN0(\Reg_Bank/registers[28][23] ), .IN1(
        \Reg_Bank/registers[29][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4711 )
         );
  MUX \Reg_Bank/U4766  ( .IN0(\Reg_Bank/registers[30][23] ), .IN1(
        \Reg_Bank/registers[31][23] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4710 )
         );
  MUX \Reg_Bank/U4765  ( .IN0(\Reg_Bank/n4709 ), .IN1(\Reg_Bank/n4694 ), .SEL(
        rs_index[4]), .F(reg_source[22]) );
  MUX \Reg_Bank/U4764  ( .IN0(\Reg_Bank/n4708 ), .IN1(\Reg_Bank/n4701 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4709 ) );
  MUX \Reg_Bank/U4763  ( .IN0(\Reg_Bank/n4707 ), .IN1(\Reg_Bank/n4704 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4708 ) );
  MUX \Reg_Bank/U4762  ( .IN0(\Reg_Bank/n4706 ), .IN1(\Reg_Bank/n4705 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4707 ) );
  MUX \Reg_Bank/U4760  ( .IN0(\Reg_Bank/registers[2][22] ), .IN1(
        \Reg_Bank/registers[3][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4705 )
         );
  MUX \Reg_Bank/U4759  ( .IN0(\Reg_Bank/n4703 ), .IN1(\Reg_Bank/n4702 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4704 ) );
  MUX \Reg_Bank/U4758  ( .IN0(\Reg_Bank/registers[4][22] ), .IN1(
        \Reg_Bank/registers[5][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4703 )
         );
  MUX \Reg_Bank/U4757  ( .IN0(\Reg_Bank/registers[6][22] ), .IN1(
        \Reg_Bank/registers[7][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4702 )
         );
  MUX \Reg_Bank/U4756  ( .IN0(\Reg_Bank/n4700 ), .IN1(\Reg_Bank/n4697 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4701 ) );
  MUX \Reg_Bank/U4755  ( .IN0(\Reg_Bank/n4699 ), .IN1(\Reg_Bank/n4698 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4700 ) );
  MUX \Reg_Bank/U4754  ( .IN0(\Reg_Bank/registers[8][22] ), .IN1(
        \Reg_Bank/registers[9][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4699 )
         );
  MUX \Reg_Bank/U4753  ( .IN0(\Reg_Bank/registers[10][22] ), .IN1(
        \Reg_Bank/registers[11][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4698 )
         );
  MUX \Reg_Bank/U4752  ( .IN0(\Reg_Bank/n4696 ), .IN1(\Reg_Bank/n4695 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4697 ) );
  MUX \Reg_Bank/U4751  ( .IN0(\Reg_Bank/registers[12][22] ), .IN1(
        \Reg_Bank/registers[13][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4696 )
         );
  MUX \Reg_Bank/U4750  ( .IN0(\Reg_Bank/registers[14][22] ), .IN1(
        \Reg_Bank/registers[15][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4695 )
         );
  MUX \Reg_Bank/U4749  ( .IN0(\Reg_Bank/n4693 ), .IN1(\Reg_Bank/n4686 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4694 ) );
  MUX \Reg_Bank/U4748  ( .IN0(\Reg_Bank/n4692 ), .IN1(\Reg_Bank/n4689 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4693 ) );
  MUX \Reg_Bank/U4747  ( .IN0(\Reg_Bank/n4691 ), .IN1(\Reg_Bank/n4690 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4692 ) );
  MUX \Reg_Bank/U4746  ( .IN0(\Reg_Bank/registers[16][22] ), .IN1(
        \Reg_Bank/registers[17][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4691 )
         );
  MUX \Reg_Bank/U4745  ( .IN0(\Reg_Bank/registers[18][22] ), .IN1(
        \Reg_Bank/registers[19][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4690 )
         );
  MUX \Reg_Bank/U4744  ( .IN0(\Reg_Bank/n4688 ), .IN1(\Reg_Bank/n4687 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4689 ) );
  MUX \Reg_Bank/U4743  ( .IN0(\Reg_Bank/registers[20][22] ), .IN1(
        \Reg_Bank/registers[21][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4688 )
         );
  MUX \Reg_Bank/U4742  ( .IN0(\Reg_Bank/registers[22][22] ), .IN1(
        \Reg_Bank/registers[23][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4687 )
         );
  MUX \Reg_Bank/U4741  ( .IN0(\Reg_Bank/n4685 ), .IN1(\Reg_Bank/n4682 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4686 ) );
  MUX \Reg_Bank/U4740  ( .IN0(\Reg_Bank/n4684 ), .IN1(\Reg_Bank/n4683 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4685 ) );
  MUX \Reg_Bank/U4739  ( .IN0(\Reg_Bank/registers[24][22] ), .IN1(
        \Reg_Bank/registers[25][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4684 )
         );
  MUX \Reg_Bank/U4738  ( .IN0(\Reg_Bank/registers[26][22] ), .IN1(
        \Reg_Bank/registers[27][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4683 )
         );
  MUX \Reg_Bank/U4737  ( .IN0(\Reg_Bank/n4681 ), .IN1(\Reg_Bank/n4680 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4682 ) );
  MUX \Reg_Bank/U4736  ( .IN0(\Reg_Bank/registers[28][22] ), .IN1(
        \Reg_Bank/registers[29][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4681 )
         );
  MUX \Reg_Bank/U4735  ( .IN0(\Reg_Bank/registers[30][22] ), .IN1(
        \Reg_Bank/registers[31][22] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4680 )
         );
  MUX \Reg_Bank/U4734  ( .IN0(\Reg_Bank/n4679 ), .IN1(\Reg_Bank/n4664 ), .SEL(
        rs_index[4]), .F(reg_source[21]) );
  MUX \Reg_Bank/U4733  ( .IN0(\Reg_Bank/n4678 ), .IN1(\Reg_Bank/n4671 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4679 ) );
  MUX \Reg_Bank/U4732  ( .IN0(\Reg_Bank/n4677 ), .IN1(\Reg_Bank/n4674 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4678 ) );
  MUX \Reg_Bank/U4731  ( .IN0(\Reg_Bank/n4676 ), .IN1(\Reg_Bank/n4675 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4677 ) );
  MUX \Reg_Bank/U4729  ( .IN0(\Reg_Bank/registers[2][21] ), .IN1(
        \Reg_Bank/registers[3][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4675 )
         );
  MUX \Reg_Bank/U4728  ( .IN0(\Reg_Bank/n4673 ), .IN1(\Reg_Bank/n4672 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4674 ) );
  MUX \Reg_Bank/U4727  ( .IN0(\Reg_Bank/registers[4][21] ), .IN1(
        \Reg_Bank/registers[5][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4673 )
         );
  MUX \Reg_Bank/U4726  ( .IN0(\Reg_Bank/registers[6][21] ), .IN1(
        \Reg_Bank/registers[7][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4672 )
         );
  MUX \Reg_Bank/U4725  ( .IN0(\Reg_Bank/n4670 ), .IN1(\Reg_Bank/n4667 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4671 ) );
  MUX \Reg_Bank/U4724  ( .IN0(\Reg_Bank/n4669 ), .IN1(\Reg_Bank/n4668 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4670 ) );
  MUX \Reg_Bank/U4723  ( .IN0(\Reg_Bank/registers[8][21] ), .IN1(
        \Reg_Bank/registers[9][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4669 )
         );
  MUX \Reg_Bank/U4722  ( .IN0(\Reg_Bank/registers[10][21] ), .IN1(
        \Reg_Bank/registers[11][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4668 )
         );
  MUX \Reg_Bank/U4721  ( .IN0(\Reg_Bank/n4666 ), .IN1(\Reg_Bank/n4665 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4667 ) );
  MUX \Reg_Bank/U4720  ( .IN0(\Reg_Bank/registers[12][21] ), .IN1(
        \Reg_Bank/registers[13][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4666 )
         );
  MUX \Reg_Bank/U4719  ( .IN0(\Reg_Bank/registers[14][21] ), .IN1(
        \Reg_Bank/registers[15][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4665 )
         );
  MUX \Reg_Bank/U4718  ( .IN0(\Reg_Bank/n4663 ), .IN1(\Reg_Bank/n4656 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4664 ) );
  MUX \Reg_Bank/U4717  ( .IN0(\Reg_Bank/n4662 ), .IN1(\Reg_Bank/n4659 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4663 ) );
  MUX \Reg_Bank/U4716  ( .IN0(\Reg_Bank/n4661 ), .IN1(\Reg_Bank/n4660 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4662 ) );
  MUX \Reg_Bank/U4715  ( .IN0(\Reg_Bank/registers[16][21] ), .IN1(
        \Reg_Bank/registers[17][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4661 )
         );
  MUX \Reg_Bank/U4714  ( .IN0(\Reg_Bank/registers[18][21] ), .IN1(
        \Reg_Bank/registers[19][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4660 )
         );
  MUX \Reg_Bank/U4713  ( .IN0(\Reg_Bank/n4658 ), .IN1(\Reg_Bank/n4657 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4659 ) );
  MUX \Reg_Bank/U4712  ( .IN0(\Reg_Bank/registers[20][21] ), .IN1(
        \Reg_Bank/registers[21][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4658 )
         );
  MUX \Reg_Bank/U4711  ( .IN0(\Reg_Bank/registers[22][21] ), .IN1(
        \Reg_Bank/registers[23][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4657 )
         );
  MUX \Reg_Bank/U4710  ( .IN0(\Reg_Bank/n4655 ), .IN1(\Reg_Bank/n4652 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4656 ) );
  MUX \Reg_Bank/U4709  ( .IN0(\Reg_Bank/n4654 ), .IN1(\Reg_Bank/n4653 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4655 ) );
  MUX \Reg_Bank/U4708  ( .IN0(\Reg_Bank/registers[24][21] ), .IN1(
        \Reg_Bank/registers[25][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4654 )
         );
  MUX \Reg_Bank/U4707  ( .IN0(\Reg_Bank/registers[26][21] ), .IN1(
        \Reg_Bank/registers[27][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4653 )
         );
  MUX \Reg_Bank/U4706  ( .IN0(\Reg_Bank/n4651 ), .IN1(\Reg_Bank/n4650 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4652 ) );
  MUX \Reg_Bank/U4705  ( .IN0(\Reg_Bank/registers[28][21] ), .IN1(
        \Reg_Bank/registers[29][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4651 )
         );
  MUX \Reg_Bank/U4704  ( .IN0(\Reg_Bank/registers[30][21] ), .IN1(
        \Reg_Bank/registers[31][21] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4650 )
         );
  MUX \Reg_Bank/U4703  ( .IN0(\Reg_Bank/n4649 ), .IN1(\Reg_Bank/n4634 ), .SEL(
        rs_index[4]), .F(reg_source[20]) );
  MUX \Reg_Bank/U4702  ( .IN0(\Reg_Bank/n4648 ), .IN1(\Reg_Bank/n4641 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4649 ) );
  MUX \Reg_Bank/U4701  ( .IN0(\Reg_Bank/n4647 ), .IN1(\Reg_Bank/n4644 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4648 ) );
  MUX \Reg_Bank/U4700  ( .IN0(\Reg_Bank/n4646 ), .IN1(\Reg_Bank/n4645 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4647 ) );
  MUX \Reg_Bank/U4698  ( .IN0(\Reg_Bank/registers[2][20] ), .IN1(
        \Reg_Bank/registers[3][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4645 )
         );
  MUX \Reg_Bank/U4697  ( .IN0(\Reg_Bank/n4643 ), .IN1(\Reg_Bank/n4642 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4644 ) );
  MUX \Reg_Bank/U4696  ( .IN0(\Reg_Bank/registers[4][20] ), .IN1(
        \Reg_Bank/registers[5][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4643 )
         );
  MUX \Reg_Bank/U4695  ( .IN0(\Reg_Bank/registers[6][20] ), .IN1(
        \Reg_Bank/registers[7][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4642 )
         );
  MUX \Reg_Bank/U4694  ( .IN0(\Reg_Bank/n4640 ), .IN1(\Reg_Bank/n4637 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4641 ) );
  MUX \Reg_Bank/U4693  ( .IN0(\Reg_Bank/n4639 ), .IN1(\Reg_Bank/n4638 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4640 ) );
  MUX \Reg_Bank/U4692  ( .IN0(\Reg_Bank/registers[8][20] ), .IN1(
        \Reg_Bank/registers[9][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4639 )
         );
  MUX \Reg_Bank/U4691  ( .IN0(\Reg_Bank/registers[10][20] ), .IN1(
        \Reg_Bank/registers[11][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4638 )
         );
  MUX \Reg_Bank/U4690  ( .IN0(\Reg_Bank/n4636 ), .IN1(\Reg_Bank/n4635 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4637 ) );
  MUX \Reg_Bank/U4689  ( .IN0(\Reg_Bank/registers[12][20] ), .IN1(
        \Reg_Bank/registers[13][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4636 )
         );
  MUX \Reg_Bank/U4688  ( .IN0(\Reg_Bank/registers[14][20] ), .IN1(
        \Reg_Bank/registers[15][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4635 )
         );
  MUX \Reg_Bank/U4687  ( .IN0(\Reg_Bank/n4633 ), .IN1(\Reg_Bank/n4626 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4634 ) );
  MUX \Reg_Bank/U4686  ( .IN0(\Reg_Bank/n4632 ), .IN1(\Reg_Bank/n4629 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4633 ) );
  MUX \Reg_Bank/U4685  ( .IN0(\Reg_Bank/n4631 ), .IN1(\Reg_Bank/n4630 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4632 ) );
  MUX \Reg_Bank/U4684  ( .IN0(\Reg_Bank/registers[16][20] ), .IN1(
        \Reg_Bank/registers[17][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4631 )
         );
  MUX \Reg_Bank/U4683  ( .IN0(\Reg_Bank/registers[18][20] ), .IN1(
        \Reg_Bank/registers[19][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4630 )
         );
  MUX \Reg_Bank/U4682  ( .IN0(\Reg_Bank/n4628 ), .IN1(\Reg_Bank/n4627 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4629 ) );
  MUX \Reg_Bank/U4681  ( .IN0(\Reg_Bank/registers[20][20] ), .IN1(
        \Reg_Bank/registers[21][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4628 )
         );
  MUX \Reg_Bank/U4680  ( .IN0(\Reg_Bank/registers[22][20] ), .IN1(
        \Reg_Bank/registers[23][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4627 )
         );
  MUX \Reg_Bank/U4679  ( .IN0(\Reg_Bank/n4625 ), .IN1(\Reg_Bank/n4622 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4626 ) );
  MUX \Reg_Bank/U4678  ( .IN0(\Reg_Bank/n4624 ), .IN1(\Reg_Bank/n4623 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4625 ) );
  MUX \Reg_Bank/U4677  ( .IN0(\Reg_Bank/registers[24][20] ), .IN1(
        \Reg_Bank/registers[25][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4624 )
         );
  MUX \Reg_Bank/U4676  ( .IN0(\Reg_Bank/registers[26][20] ), .IN1(
        \Reg_Bank/registers[27][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4623 )
         );
  MUX \Reg_Bank/U4675  ( .IN0(\Reg_Bank/n4621 ), .IN1(\Reg_Bank/n4620 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4622 ) );
  MUX \Reg_Bank/U4674  ( .IN0(\Reg_Bank/registers[28][20] ), .IN1(
        \Reg_Bank/registers[29][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4621 )
         );
  MUX \Reg_Bank/U4673  ( .IN0(\Reg_Bank/registers[30][20] ), .IN1(
        \Reg_Bank/registers[31][20] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4620 )
         );
  MUX \Reg_Bank/U4672  ( .IN0(\Reg_Bank/n4619 ), .IN1(\Reg_Bank/n4604 ), .SEL(
        rs_index[4]), .F(reg_source[19]) );
  MUX \Reg_Bank/U4671  ( .IN0(\Reg_Bank/n4618 ), .IN1(\Reg_Bank/n4611 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4619 ) );
  MUX \Reg_Bank/U4670  ( .IN0(\Reg_Bank/n4617 ), .IN1(\Reg_Bank/n4614 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4618 ) );
  MUX \Reg_Bank/U4669  ( .IN0(\Reg_Bank/n4616 ), .IN1(\Reg_Bank/n4615 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4617 ) );
  MUX \Reg_Bank/U4667  ( .IN0(\Reg_Bank/registers[2][19] ), .IN1(
        \Reg_Bank/registers[3][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4615 )
         );
  MUX \Reg_Bank/U4666  ( .IN0(\Reg_Bank/n4613 ), .IN1(\Reg_Bank/n4612 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4614 ) );
  MUX \Reg_Bank/U4665  ( .IN0(\Reg_Bank/registers[4][19] ), .IN1(
        \Reg_Bank/registers[5][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4613 )
         );
  MUX \Reg_Bank/U4664  ( .IN0(\Reg_Bank/registers[6][19] ), .IN1(
        \Reg_Bank/registers[7][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4612 )
         );
  MUX \Reg_Bank/U4663  ( .IN0(\Reg_Bank/n4610 ), .IN1(\Reg_Bank/n4607 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4611 ) );
  MUX \Reg_Bank/U4662  ( .IN0(\Reg_Bank/n4609 ), .IN1(\Reg_Bank/n4608 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4610 ) );
  MUX \Reg_Bank/U4661  ( .IN0(\Reg_Bank/registers[8][19] ), .IN1(
        \Reg_Bank/registers[9][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4609 )
         );
  MUX \Reg_Bank/U4660  ( .IN0(\Reg_Bank/registers[10][19] ), .IN1(
        \Reg_Bank/registers[11][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4608 )
         );
  MUX \Reg_Bank/U4659  ( .IN0(\Reg_Bank/n4606 ), .IN1(\Reg_Bank/n4605 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4607 ) );
  MUX \Reg_Bank/U4658  ( .IN0(\Reg_Bank/registers[12][19] ), .IN1(
        \Reg_Bank/registers[13][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4606 )
         );
  MUX \Reg_Bank/U4657  ( .IN0(\Reg_Bank/registers[14][19] ), .IN1(
        \Reg_Bank/registers[15][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4605 )
         );
  MUX \Reg_Bank/U4656  ( .IN0(\Reg_Bank/n4603 ), .IN1(\Reg_Bank/n4596 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4604 ) );
  MUX \Reg_Bank/U4655  ( .IN0(\Reg_Bank/n4602 ), .IN1(\Reg_Bank/n4599 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4603 ) );
  MUX \Reg_Bank/U4654  ( .IN0(\Reg_Bank/n4601 ), .IN1(\Reg_Bank/n4600 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4602 ) );
  MUX \Reg_Bank/U4653  ( .IN0(\Reg_Bank/registers[16][19] ), .IN1(
        \Reg_Bank/registers[17][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4601 )
         );
  MUX \Reg_Bank/U4652  ( .IN0(\Reg_Bank/registers[18][19] ), .IN1(
        \Reg_Bank/registers[19][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4600 )
         );
  MUX \Reg_Bank/U4651  ( .IN0(\Reg_Bank/n4598 ), .IN1(\Reg_Bank/n4597 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4599 ) );
  MUX \Reg_Bank/U4650  ( .IN0(\Reg_Bank/registers[20][19] ), .IN1(
        \Reg_Bank/registers[21][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4598 )
         );
  MUX \Reg_Bank/U4649  ( .IN0(\Reg_Bank/registers[22][19] ), .IN1(
        \Reg_Bank/registers[23][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4597 )
         );
  MUX \Reg_Bank/U4648  ( .IN0(\Reg_Bank/n4595 ), .IN1(\Reg_Bank/n4592 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4596 ) );
  MUX \Reg_Bank/U4647  ( .IN0(\Reg_Bank/n4594 ), .IN1(\Reg_Bank/n4593 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4595 ) );
  MUX \Reg_Bank/U4646  ( .IN0(\Reg_Bank/registers[24][19] ), .IN1(
        \Reg_Bank/registers[25][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4594 )
         );
  MUX \Reg_Bank/U4645  ( .IN0(\Reg_Bank/registers[26][19] ), .IN1(
        \Reg_Bank/registers[27][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4593 )
         );
  MUX \Reg_Bank/U4644  ( .IN0(\Reg_Bank/n4591 ), .IN1(\Reg_Bank/n4590 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4592 ) );
  MUX \Reg_Bank/U4643  ( .IN0(\Reg_Bank/registers[28][19] ), .IN1(
        \Reg_Bank/registers[29][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4591 )
         );
  MUX \Reg_Bank/U4642  ( .IN0(\Reg_Bank/registers[30][19] ), .IN1(
        \Reg_Bank/registers[31][19] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4590 )
         );
  MUX \Reg_Bank/U4641  ( .IN0(\Reg_Bank/n4589 ), .IN1(\Reg_Bank/n4574 ), .SEL(
        rs_index[4]), .F(reg_source[18]) );
  MUX \Reg_Bank/U4640  ( .IN0(\Reg_Bank/n4588 ), .IN1(\Reg_Bank/n4581 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4589 ) );
  MUX \Reg_Bank/U4639  ( .IN0(\Reg_Bank/n4587 ), .IN1(\Reg_Bank/n4584 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4588 ) );
  MUX \Reg_Bank/U4638  ( .IN0(\Reg_Bank/n4586 ), .IN1(\Reg_Bank/n4585 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4587 ) );
  MUX \Reg_Bank/U4636  ( .IN0(\Reg_Bank/registers[2][18] ), .IN1(
        \Reg_Bank/registers[3][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4585 )
         );
  MUX \Reg_Bank/U4635  ( .IN0(\Reg_Bank/n4583 ), .IN1(\Reg_Bank/n4582 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4584 ) );
  MUX \Reg_Bank/U4634  ( .IN0(\Reg_Bank/registers[4][18] ), .IN1(
        \Reg_Bank/registers[5][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4583 )
         );
  MUX \Reg_Bank/U4633  ( .IN0(\Reg_Bank/registers[6][18] ), .IN1(
        \Reg_Bank/registers[7][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4582 )
         );
  MUX \Reg_Bank/U4632  ( .IN0(\Reg_Bank/n4580 ), .IN1(\Reg_Bank/n4577 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4581 ) );
  MUX \Reg_Bank/U4631  ( .IN0(\Reg_Bank/n4579 ), .IN1(\Reg_Bank/n4578 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4580 ) );
  MUX \Reg_Bank/U4630  ( .IN0(\Reg_Bank/registers[8][18] ), .IN1(
        \Reg_Bank/registers[9][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4579 )
         );
  MUX \Reg_Bank/U4629  ( .IN0(\Reg_Bank/registers[10][18] ), .IN1(
        \Reg_Bank/registers[11][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4578 )
         );
  MUX \Reg_Bank/U4628  ( .IN0(\Reg_Bank/n4576 ), .IN1(\Reg_Bank/n4575 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4577 ) );
  MUX \Reg_Bank/U4627  ( .IN0(\Reg_Bank/registers[12][18] ), .IN1(
        \Reg_Bank/registers[13][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4576 )
         );
  MUX \Reg_Bank/U4626  ( .IN0(\Reg_Bank/registers[14][18] ), .IN1(
        \Reg_Bank/registers[15][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4575 )
         );
  MUX \Reg_Bank/U4625  ( .IN0(\Reg_Bank/n4573 ), .IN1(\Reg_Bank/n4566 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4574 ) );
  MUX \Reg_Bank/U4624  ( .IN0(\Reg_Bank/n4572 ), .IN1(\Reg_Bank/n4569 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4573 ) );
  MUX \Reg_Bank/U4623  ( .IN0(\Reg_Bank/n4571 ), .IN1(\Reg_Bank/n4570 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4572 ) );
  MUX \Reg_Bank/U4622  ( .IN0(\Reg_Bank/registers[16][18] ), .IN1(
        \Reg_Bank/registers[17][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4571 )
         );
  MUX \Reg_Bank/U4621  ( .IN0(\Reg_Bank/registers[18][18] ), .IN1(
        \Reg_Bank/registers[19][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4570 )
         );
  MUX \Reg_Bank/U4620  ( .IN0(\Reg_Bank/n4568 ), .IN1(\Reg_Bank/n4567 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4569 ) );
  MUX \Reg_Bank/U4619  ( .IN0(\Reg_Bank/registers[20][18] ), .IN1(
        \Reg_Bank/registers[21][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4568 )
         );
  MUX \Reg_Bank/U4618  ( .IN0(\Reg_Bank/registers[22][18] ), .IN1(
        \Reg_Bank/registers[23][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4567 )
         );
  MUX \Reg_Bank/U4617  ( .IN0(\Reg_Bank/n4565 ), .IN1(\Reg_Bank/n4562 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4566 ) );
  MUX \Reg_Bank/U4616  ( .IN0(\Reg_Bank/n4564 ), .IN1(\Reg_Bank/n4563 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4565 ) );
  MUX \Reg_Bank/U4615  ( .IN0(\Reg_Bank/registers[24][18] ), .IN1(
        \Reg_Bank/registers[25][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4564 )
         );
  MUX \Reg_Bank/U4614  ( .IN0(\Reg_Bank/registers[26][18] ), .IN1(
        \Reg_Bank/registers[27][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4563 )
         );
  MUX \Reg_Bank/U4613  ( .IN0(\Reg_Bank/n4561 ), .IN1(\Reg_Bank/n4560 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4562 ) );
  MUX \Reg_Bank/U4612  ( .IN0(\Reg_Bank/registers[28][18] ), .IN1(
        \Reg_Bank/registers[29][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4561 )
         );
  MUX \Reg_Bank/U4611  ( .IN0(\Reg_Bank/registers[30][18] ), .IN1(
        \Reg_Bank/registers[31][18] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4560 )
         );
  MUX \Reg_Bank/U4610  ( .IN0(\Reg_Bank/n4559 ), .IN1(\Reg_Bank/n4544 ), .SEL(
        rs_index[4]), .F(reg_source[17]) );
  MUX \Reg_Bank/U4609  ( .IN0(\Reg_Bank/n4558 ), .IN1(\Reg_Bank/n4551 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4559 ) );
  MUX \Reg_Bank/U4608  ( .IN0(\Reg_Bank/n4557 ), .IN1(\Reg_Bank/n4554 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4558 ) );
  MUX \Reg_Bank/U4607  ( .IN0(\Reg_Bank/n4556 ), .IN1(\Reg_Bank/n4555 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4557 ) );
  MUX \Reg_Bank/U4605  ( .IN0(\Reg_Bank/registers[2][17] ), .IN1(
        \Reg_Bank/registers[3][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4555 )
         );
  MUX \Reg_Bank/U4604  ( .IN0(\Reg_Bank/n4553 ), .IN1(\Reg_Bank/n4552 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4554 ) );
  MUX \Reg_Bank/U4603  ( .IN0(\Reg_Bank/registers[4][17] ), .IN1(
        \Reg_Bank/registers[5][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4553 )
         );
  MUX \Reg_Bank/U4602  ( .IN0(\Reg_Bank/registers[6][17] ), .IN1(
        \Reg_Bank/registers[7][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4552 )
         );
  MUX \Reg_Bank/U4601  ( .IN0(\Reg_Bank/n4550 ), .IN1(\Reg_Bank/n4547 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4551 ) );
  MUX \Reg_Bank/U4600  ( .IN0(\Reg_Bank/n4549 ), .IN1(\Reg_Bank/n4548 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4550 ) );
  MUX \Reg_Bank/U4599  ( .IN0(\Reg_Bank/registers[8][17] ), .IN1(
        \Reg_Bank/registers[9][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4549 )
         );
  MUX \Reg_Bank/U4598  ( .IN0(\Reg_Bank/registers[10][17] ), .IN1(
        \Reg_Bank/registers[11][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4548 )
         );
  MUX \Reg_Bank/U4597  ( .IN0(\Reg_Bank/n4546 ), .IN1(\Reg_Bank/n4545 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4547 ) );
  MUX \Reg_Bank/U4596  ( .IN0(\Reg_Bank/registers[12][17] ), .IN1(
        \Reg_Bank/registers[13][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4546 )
         );
  MUX \Reg_Bank/U4595  ( .IN0(\Reg_Bank/registers[14][17] ), .IN1(
        \Reg_Bank/registers[15][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4545 )
         );
  MUX \Reg_Bank/U4594  ( .IN0(\Reg_Bank/n4543 ), .IN1(\Reg_Bank/n4536 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4544 ) );
  MUX \Reg_Bank/U4593  ( .IN0(\Reg_Bank/n4542 ), .IN1(\Reg_Bank/n4539 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4543 ) );
  MUX \Reg_Bank/U4592  ( .IN0(\Reg_Bank/n4541 ), .IN1(\Reg_Bank/n4540 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4542 ) );
  MUX \Reg_Bank/U4591  ( .IN0(\Reg_Bank/registers[16][17] ), .IN1(
        \Reg_Bank/registers[17][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4541 )
         );
  MUX \Reg_Bank/U4590  ( .IN0(\Reg_Bank/registers[18][17] ), .IN1(
        \Reg_Bank/registers[19][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4540 )
         );
  MUX \Reg_Bank/U4589  ( .IN0(\Reg_Bank/n4538 ), .IN1(\Reg_Bank/n4537 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4539 ) );
  MUX \Reg_Bank/U4588  ( .IN0(\Reg_Bank/registers[20][17] ), .IN1(
        \Reg_Bank/registers[21][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4538 )
         );
  MUX \Reg_Bank/U4587  ( .IN0(\Reg_Bank/registers[22][17] ), .IN1(
        \Reg_Bank/registers[23][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4537 )
         );
  MUX \Reg_Bank/U4586  ( .IN0(\Reg_Bank/n4535 ), .IN1(\Reg_Bank/n4532 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4536 ) );
  MUX \Reg_Bank/U4585  ( .IN0(\Reg_Bank/n4534 ), .IN1(\Reg_Bank/n4533 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4535 ) );
  MUX \Reg_Bank/U4584  ( .IN0(\Reg_Bank/registers[24][17] ), .IN1(
        \Reg_Bank/registers[25][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4534 )
         );
  MUX \Reg_Bank/U4583  ( .IN0(\Reg_Bank/registers[26][17] ), .IN1(
        \Reg_Bank/registers[27][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4533 )
         );
  MUX \Reg_Bank/U4582  ( .IN0(\Reg_Bank/n4531 ), .IN1(\Reg_Bank/n4530 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4532 ) );
  MUX \Reg_Bank/U4581  ( .IN0(\Reg_Bank/registers[28][17] ), .IN1(
        \Reg_Bank/registers[29][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4531 )
         );
  MUX \Reg_Bank/U4580  ( .IN0(\Reg_Bank/registers[30][17] ), .IN1(
        \Reg_Bank/registers[31][17] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4530 )
         );
  MUX \Reg_Bank/U4579  ( .IN0(\Reg_Bank/n4529 ), .IN1(\Reg_Bank/n4514 ), .SEL(
        rs_index[4]), .F(reg_source[16]) );
  MUX \Reg_Bank/U4578  ( .IN0(\Reg_Bank/n4528 ), .IN1(\Reg_Bank/n4521 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4529 ) );
  MUX \Reg_Bank/U4577  ( .IN0(\Reg_Bank/n4527 ), .IN1(\Reg_Bank/n4524 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4528 ) );
  MUX \Reg_Bank/U4576  ( .IN0(\Reg_Bank/n4526 ), .IN1(\Reg_Bank/n4525 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4527 ) );
  MUX \Reg_Bank/U4574  ( .IN0(\Reg_Bank/registers[2][16] ), .IN1(
        \Reg_Bank/registers[3][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4525 )
         );
  MUX \Reg_Bank/U4573  ( .IN0(\Reg_Bank/n4523 ), .IN1(\Reg_Bank/n4522 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4524 ) );
  MUX \Reg_Bank/U4572  ( .IN0(\Reg_Bank/registers[4][16] ), .IN1(
        \Reg_Bank/registers[5][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4523 )
         );
  MUX \Reg_Bank/U4571  ( .IN0(\Reg_Bank/registers[6][16] ), .IN1(
        \Reg_Bank/registers[7][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4522 )
         );
  MUX \Reg_Bank/U4570  ( .IN0(\Reg_Bank/n4520 ), .IN1(\Reg_Bank/n4517 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4521 ) );
  MUX \Reg_Bank/U4569  ( .IN0(\Reg_Bank/n4519 ), .IN1(\Reg_Bank/n4518 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4520 ) );
  MUX \Reg_Bank/U4568  ( .IN0(\Reg_Bank/registers[8][16] ), .IN1(
        \Reg_Bank/registers[9][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4519 )
         );
  MUX \Reg_Bank/U4567  ( .IN0(\Reg_Bank/registers[10][16] ), .IN1(
        \Reg_Bank/registers[11][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4518 )
         );
  MUX \Reg_Bank/U4566  ( .IN0(\Reg_Bank/n4516 ), .IN1(\Reg_Bank/n4515 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4517 ) );
  MUX \Reg_Bank/U4565  ( .IN0(\Reg_Bank/registers[12][16] ), .IN1(
        \Reg_Bank/registers[13][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4516 )
         );
  MUX \Reg_Bank/U4564  ( .IN0(\Reg_Bank/registers[14][16] ), .IN1(
        \Reg_Bank/registers[15][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4515 )
         );
  MUX \Reg_Bank/U4563  ( .IN0(\Reg_Bank/n4513 ), .IN1(\Reg_Bank/n4506 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4514 ) );
  MUX \Reg_Bank/U4562  ( .IN0(\Reg_Bank/n4512 ), .IN1(\Reg_Bank/n4509 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4513 ) );
  MUX \Reg_Bank/U4561  ( .IN0(\Reg_Bank/n4511 ), .IN1(\Reg_Bank/n4510 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4512 ) );
  MUX \Reg_Bank/U4560  ( .IN0(\Reg_Bank/registers[16][16] ), .IN1(
        \Reg_Bank/registers[17][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4511 )
         );
  MUX \Reg_Bank/U4559  ( .IN0(\Reg_Bank/registers[18][16] ), .IN1(
        \Reg_Bank/registers[19][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4510 )
         );
  MUX \Reg_Bank/U4558  ( .IN0(\Reg_Bank/n4508 ), .IN1(\Reg_Bank/n4507 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4509 ) );
  MUX \Reg_Bank/U4557  ( .IN0(\Reg_Bank/registers[20][16] ), .IN1(
        \Reg_Bank/registers[21][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4508 )
         );
  MUX \Reg_Bank/U4556  ( .IN0(\Reg_Bank/registers[22][16] ), .IN1(
        \Reg_Bank/registers[23][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4507 )
         );
  MUX \Reg_Bank/U4555  ( .IN0(\Reg_Bank/n4505 ), .IN1(\Reg_Bank/n4502 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4506 ) );
  MUX \Reg_Bank/U4554  ( .IN0(\Reg_Bank/n4504 ), .IN1(\Reg_Bank/n4503 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4505 ) );
  MUX \Reg_Bank/U4553  ( .IN0(\Reg_Bank/registers[24][16] ), .IN1(
        \Reg_Bank/registers[25][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4504 )
         );
  MUX \Reg_Bank/U4552  ( .IN0(\Reg_Bank/registers[26][16] ), .IN1(
        \Reg_Bank/registers[27][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4503 )
         );
  MUX \Reg_Bank/U4551  ( .IN0(\Reg_Bank/n4501 ), .IN1(\Reg_Bank/n4500 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4502 ) );
  MUX \Reg_Bank/U4550  ( .IN0(\Reg_Bank/registers[28][16] ), .IN1(
        \Reg_Bank/registers[29][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4501 )
         );
  MUX \Reg_Bank/U4549  ( .IN0(\Reg_Bank/registers[30][16] ), .IN1(
        \Reg_Bank/registers[31][16] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4500 )
         );
  MUX \Reg_Bank/U4548  ( .IN0(\Reg_Bank/n4499 ), .IN1(\Reg_Bank/n4484 ), .SEL(
        rs_index[4]), .F(reg_source[15]) );
  MUX \Reg_Bank/U4547  ( .IN0(\Reg_Bank/n4498 ), .IN1(\Reg_Bank/n4491 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4499 ) );
  MUX \Reg_Bank/U4546  ( .IN0(\Reg_Bank/n4497 ), .IN1(\Reg_Bank/n4494 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4498 ) );
  MUX \Reg_Bank/U4545  ( .IN0(\Reg_Bank/n4496 ), .IN1(\Reg_Bank/n4495 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4497 ) );
  MUX \Reg_Bank/U4543  ( .IN0(\Reg_Bank/registers[2][15] ), .IN1(
        \Reg_Bank/registers[3][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4495 )
         );
  MUX \Reg_Bank/U4542  ( .IN0(\Reg_Bank/n4493 ), .IN1(\Reg_Bank/n4492 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4494 ) );
  MUX \Reg_Bank/U4541  ( .IN0(\Reg_Bank/registers[4][15] ), .IN1(
        \Reg_Bank/registers[5][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4493 )
         );
  MUX \Reg_Bank/U4540  ( .IN0(\Reg_Bank/registers[6][15] ), .IN1(
        \Reg_Bank/registers[7][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4492 )
         );
  MUX \Reg_Bank/U4539  ( .IN0(\Reg_Bank/n4490 ), .IN1(\Reg_Bank/n4487 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4491 ) );
  MUX \Reg_Bank/U4538  ( .IN0(\Reg_Bank/n4489 ), .IN1(\Reg_Bank/n4488 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4490 ) );
  MUX \Reg_Bank/U4537  ( .IN0(\Reg_Bank/registers[8][15] ), .IN1(
        \Reg_Bank/registers[9][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4489 )
         );
  MUX \Reg_Bank/U4536  ( .IN0(\Reg_Bank/registers[10][15] ), .IN1(
        \Reg_Bank/registers[11][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4488 )
         );
  MUX \Reg_Bank/U4535  ( .IN0(\Reg_Bank/n4486 ), .IN1(\Reg_Bank/n4485 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4487 ) );
  MUX \Reg_Bank/U4534  ( .IN0(\Reg_Bank/registers[12][15] ), .IN1(
        \Reg_Bank/registers[13][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4486 )
         );
  MUX \Reg_Bank/U4533  ( .IN0(\Reg_Bank/registers[14][15] ), .IN1(
        \Reg_Bank/registers[15][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4485 )
         );
  MUX \Reg_Bank/U4532  ( .IN0(\Reg_Bank/n4483 ), .IN1(\Reg_Bank/n4476 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4484 ) );
  MUX \Reg_Bank/U4531  ( .IN0(\Reg_Bank/n4482 ), .IN1(\Reg_Bank/n4479 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4483 ) );
  MUX \Reg_Bank/U4530  ( .IN0(\Reg_Bank/n4481 ), .IN1(\Reg_Bank/n4480 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4482 ) );
  MUX \Reg_Bank/U4529  ( .IN0(\Reg_Bank/registers[16][15] ), .IN1(
        \Reg_Bank/registers[17][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4481 )
         );
  MUX \Reg_Bank/U4528  ( .IN0(\Reg_Bank/registers[18][15] ), .IN1(
        \Reg_Bank/registers[19][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4480 )
         );
  MUX \Reg_Bank/U4527  ( .IN0(\Reg_Bank/n4478 ), .IN1(\Reg_Bank/n4477 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4479 ) );
  MUX \Reg_Bank/U4526  ( .IN0(\Reg_Bank/registers[20][15] ), .IN1(
        \Reg_Bank/registers[21][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4478 )
         );
  MUX \Reg_Bank/U4525  ( .IN0(\Reg_Bank/registers[22][15] ), .IN1(
        \Reg_Bank/registers[23][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4477 )
         );
  MUX \Reg_Bank/U4524  ( .IN0(\Reg_Bank/n4475 ), .IN1(\Reg_Bank/n4472 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4476 ) );
  MUX \Reg_Bank/U4523  ( .IN0(\Reg_Bank/n4474 ), .IN1(\Reg_Bank/n4473 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4475 ) );
  MUX \Reg_Bank/U4522  ( .IN0(\Reg_Bank/registers[24][15] ), .IN1(
        \Reg_Bank/registers[25][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4474 )
         );
  MUX \Reg_Bank/U4521  ( .IN0(\Reg_Bank/registers[26][15] ), .IN1(
        \Reg_Bank/registers[27][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4473 )
         );
  MUX \Reg_Bank/U4520  ( .IN0(\Reg_Bank/n4471 ), .IN1(\Reg_Bank/n4470 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4472 ) );
  MUX \Reg_Bank/U4519  ( .IN0(\Reg_Bank/registers[28][15] ), .IN1(
        \Reg_Bank/registers[29][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4471 )
         );
  MUX \Reg_Bank/U4518  ( .IN0(\Reg_Bank/registers[30][15] ), .IN1(
        \Reg_Bank/registers[31][15] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4470 )
         );
  MUX \Reg_Bank/U4517  ( .IN0(\Reg_Bank/n4469 ), .IN1(\Reg_Bank/n4454 ), .SEL(
        rs_index[4]), .F(reg_source[14]) );
  MUX \Reg_Bank/U4516  ( .IN0(\Reg_Bank/n4468 ), .IN1(\Reg_Bank/n4461 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4469 ) );
  MUX \Reg_Bank/U4515  ( .IN0(\Reg_Bank/n4467 ), .IN1(\Reg_Bank/n4464 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4468 ) );
  MUX \Reg_Bank/U4514  ( .IN0(\Reg_Bank/n4466 ), .IN1(\Reg_Bank/n4465 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4467 ) );
  MUX \Reg_Bank/U4512  ( .IN0(\Reg_Bank/registers[2][14] ), .IN1(
        \Reg_Bank/registers[3][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4465 )
         );
  MUX \Reg_Bank/U4511  ( .IN0(\Reg_Bank/n4463 ), .IN1(\Reg_Bank/n4462 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4464 ) );
  MUX \Reg_Bank/U4510  ( .IN0(\Reg_Bank/registers[4][14] ), .IN1(
        \Reg_Bank/registers[5][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4463 )
         );
  MUX \Reg_Bank/U4509  ( .IN0(\Reg_Bank/registers[6][14] ), .IN1(
        \Reg_Bank/registers[7][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4462 )
         );
  MUX \Reg_Bank/U4508  ( .IN0(\Reg_Bank/n4460 ), .IN1(\Reg_Bank/n4457 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4461 ) );
  MUX \Reg_Bank/U4507  ( .IN0(\Reg_Bank/n4459 ), .IN1(\Reg_Bank/n4458 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4460 ) );
  MUX \Reg_Bank/U4506  ( .IN0(\Reg_Bank/registers[8][14] ), .IN1(
        \Reg_Bank/registers[9][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4459 )
         );
  MUX \Reg_Bank/U4505  ( .IN0(\Reg_Bank/registers[10][14] ), .IN1(
        \Reg_Bank/registers[11][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4458 )
         );
  MUX \Reg_Bank/U4504  ( .IN0(\Reg_Bank/n4456 ), .IN1(\Reg_Bank/n4455 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4457 ) );
  MUX \Reg_Bank/U4503  ( .IN0(\Reg_Bank/registers[12][14] ), .IN1(
        \Reg_Bank/registers[13][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4456 )
         );
  MUX \Reg_Bank/U4502  ( .IN0(\Reg_Bank/registers[14][14] ), .IN1(
        \Reg_Bank/registers[15][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4455 )
         );
  MUX \Reg_Bank/U4501  ( .IN0(\Reg_Bank/n4453 ), .IN1(\Reg_Bank/n4446 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4454 ) );
  MUX \Reg_Bank/U4500  ( .IN0(\Reg_Bank/n4452 ), .IN1(\Reg_Bank/n4449 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4453 ) );
  MUX \Reg_Bank/U4499  ( .IN0(\Reg_Bank/n4451 ), .IN1(\Reg_Bank/n4450 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4452 ) );
  MUX \Reg_Bank/U4498  ( .IN0(\Reg_Bank/registers[16][14] ), .IN1(
        \Reg_Bank/registers[17][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4451 )
         );
  MUX \Reg_Bank/U4497  ( .IN0(\Reg_Bank/registers[18][14] ), .IN1(
        \Reg_Bank/registers[19][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4450 )
         );
  MUX \Reg_Bank/U4496  ( .IN0(\Reg_Bank/n4448 ), .IN1(\Reg_Bank/n4447 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4449 ) );
  MUX \Reg_Bank/U4495  ( .IN0(\Reg_Bank/registers[20][14] ), .IN1(
        \Reg_Bank/registers[21][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4448 )
         );
  MUX \Reg_Bank/U4494  ( .IN0(\Reg_Bank/registers[22][14] ), .IN1(
        \Reg_Bank/registers[23][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4447 )
         );
  MUX \Reg_Bank/U4493  ( .IN0(\Reg_Bank/n4445 ), .IN1(\Reg_Bank/n4442 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4446 ) );
  MUX \Reg_Bank/U4492  ( .IN0(\Reg_Bank/n4444 ), .IN1(\Reg_Bank/n4443 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4445 ) );
  MUX \Reg_Bank/U4491  ( .IN0(\Reg_Bank/registers[24][14] ), .IN1(
        \Reg_Bank/registers[25][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4444 )
         );
  MUX \Reg_Bank/U4490  ( .IN0(\Reg_Bank/registers[26][14] ), .IN1(
        \Reg_Bank/registers[27][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4443 )
         );
  MUX \Reg_Bank/U4489  ( .IN0(\Reg_Bank/n4441 ), .IN1(\Reg_Bank/n4440 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4442 ) );
  MUX \Reg_Bank/U4488  ( .IN0(\Reg_Bank/registers[28][14] ), .IN1(
        \Reg_Bank/registers[29][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4441 )
         );
  MUX \Reg_Bank/U4487  ( .IN0(\Reg_Bank/registers[30][14] ), .IN1(
        \Reg_Bank/registers[31][14] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4440 )
         );
  MUX \Reg_Bank/U4486  ( .IN0(\Reg_Bank/n4439 ), .IN1(\Reg_Bank/n4424 ), .SEL(
        rs_index[4]), .F(reg_source[13]) );
  MUX \Reg_Bank/U4485  ( .IN0(\Reg_Bank/n4438 ), .IN1(\Reg_Bank/n4431 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4439 ) );
  MUX \Reg_Bank/U4484  ( .IN0(\Reg_Bank/n4437 ), .IN1(\Reg_Bank/n4434 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4438 ) );
  MUX \Reg_Bank/U4483  ( .IN0(\Reg_Bank/n4436 ), .IN1(\Reg_Bank/n4435 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4437 ) );
  MUX \Reg_Bank/U4481  ( .IN0(\Reg_Bank/registers[2][13] ), .IN1(
        \Reg_Bank/registers[3][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4435 )
         );
  MUX \Reg_Bank/U4480  ( .IN0(\Reg_Bank/n4433 ), .IN1(\Reg_Bank/n4432 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4434 ) );
  MUX \Reg_Bank/U4479  ( .IN0(\Reg_Bank/registers[4][13] ), .IN1(
        \Reg_Bank/registers[5][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4433 )
         );
  MUX \Reg_Bank/U4478  ( .IN0(\Reg_Bank/registers[6][13] ), .IN1(
        \Reg_Bank/registers[7][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4432 )
         );
  MUX \Reg_Bank/U4477  ( .IN0(\Reg_Bank/n4430 ), .IN1(\Reg_Bank/n4427 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4431 ) );
  MUX \Reg_Bank/U4476  ( .IN0(\Reg_Bank/n4429 ), .IN1(\Reg_Bank/n4428 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4430 ) );
  MUX \Reg_Bank/U4475  ( .IN0(\Reg_Bank/registers[8][13] ), .IN1(
        \Reg_Bank/registers[9][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4429 )
         );
  MUX \Reg_Bank/U4474  ( .IN0(\Reg_Bank/registers[10][13] ), .IN1(
        \Reg_Bank/registers[11][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4428 )
         );
  MUX \Reg_Bank/U4473  ( .IN0(\Reg_Bank/n4426 ), .IN1(\Reg_Bank/n4425 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4427 ) );
  MUX \Reg_Bank/U4472  ( .IN0(\Reg_Bank/registers[12][13] ), .IN1(
        \Reg_Bank/registers[13][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4426 )
         );
  MUX \Reg_Bank/U4471  ( .IN0(\Reg_Bank/registers[14][13] ), .IN1(
        \Reg_Bank/registers[15][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4425 )
         );
  MUX \Reg_Bank/U4470  ( .IN0(\Reg_Bank/n4423 ), .IN1(\Reg_Bank/n4416 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4424 ) );
  MUX \Reg_Bank/U4469  ( .IN0(\Reg_Bank/n4422 ), .IN1(\Reg_Bank/n4419 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4423 ) );
  MUX \Reg_Bank/U4468  ( .IN0(\Reg_Bank/n4421 ), .IN1(\Reg_Bank/n4420 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4422 ) );
  MUX \Reg_Bank/U4467  ( .IN0(\Reg_Bank/registers[16][13] ), .IN1(
        \Reg_Bank/registers[17][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4421 )
         );
  MUX \Reg_Bank/U4466  ( .IN0(\Reg_Bank/registers[18][13] ), .IN1(
        \Reg_Bank/registers[19][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4420 )
         );
  MUX \Reg_Bank/U4465  ( .IN0(\Reg_Bank/n4418 ), .IN1(\Reg_Bank/n4417 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4419 ) );
  MUX \Reg_Bank/U4464  ( .IN0(\Reg_Bank/registers[20][13] ), .IN1(
        \Reg_Bank/registers[21][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4418 )
         );
  MUX \Reg_Bank/U4463  ( .IN0(\Reg_Bank/registers[22][13] ), .IN1(
        \Reg_Bank/registers[23][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4417 )
         );
  MUX \Reg_Bank/U4462  ( .IN0(\Reg_Bank/n4415 ), .IN1(\Reg_Bank/n4412 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4416 ) );
  MUX \Reg_Bank/U4461  ( .IN0(\Reg_Bank/n4414 ), .IN1(\Reg_Bank/n4413 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4415 ) );
  MUX \Reg_Bank/U4460  ( .IN0(\Reg_Bank/registers[24][13] ), .IN1(
        \Reg_Bank/registers[25][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4414 )
         );
  MUX \Reg_Bank/U4459  ( .IN0(\Reg_Bank/registers[26][13] ), .IN1(
        \Reg_Bank/registers[27][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4413 )
         );
  MUX \Reg_Bank/U4458  ( .IN0(\Reg_Bank/n4411 ), .IN1(\Reg_Bank/n4410 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4412 ) );
  MUX \Reg_Bank/U4457  ( .IN0(\Reg_Bank/registers[28][13] ), .IN1(
        \Reg_Bank/registers[29][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4411 )
         );
  MUX \Reg_Bank/U4456  ( .IN0(\Reg_Bank/registers[30][13] ), .IN1(
        \Reg_Bank/registers[31][13] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4410 )
         );
  MUX \Reg_Bank/U4455  ( .IN0(\Reg_Bank/n4409 ), .IN1(\Reg_Bank/n4394 ), .SEL(
        rs_index[4]), .F(reg_source[12]) );
  MUX \Reg_Bank/U4454  ( .IN0(\Reg_Bank/n4408 ), .IN1(\Reg_Bank/n4401 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4409 ) );
  MUX \Reg_Bank/U4453  ( .IN0(\Reg_Bank/n4407 ), .IN1(\Reg_Bank/n4404 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4408 ) );
  MUX \Reg_Bank/U4452  ( .IN0(\Reg_Bank/n4406 ), .IN1(\Reg_Bank/n4405 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4407 ) );
  MUX \Reg_Bank/U4450  ( .IN0(\Reg_Bank/registers[2][12] ), .IN1(
        \Reg_Bank/registers[3][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4405 )
         );
  MUX \Reg_Bank/U4449  ( .IN0(\Reg_Bank/n4403 ), .IN1(\Reg_Bank/n4402 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4404 ) );
  MUX \Reg_Bank/U4448  ( .IN0(\Reg_Bank/registers[4][12] ), .IN1(
        \Reg_Bank/registers[5][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4403 )
         );
  MUX \Reg_Bank/U4447  ( .IN0(\Reg_Bank/registers[6][12] ), .IN1(
        \Reg_Bank/registers[7][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4402 )
         );
  MUX \Reg_Bank/U4446  ( .IN0(\Reg_Bank/n4400 ), .IN1(\Reg_Bank/n4397 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4401 ) );
  MUX \Reg_Bank/U4445  ( .IN0(\Reg_Bank/n4399 ), .IN1(\Reg_Bank/n4398 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4400 ) );
  MUX \Reg_Bank/U4444  ( .IN0(\Reg_Bank/registers[8][12] ), .IN1(
        \Reg_Bank/registers[9][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4399 )
         );
  MUX \Reg_Bank/U4443  ( .IN0(\Reg_Bank/registers[10][12] ), .IN1(
        \Reg_Bank/registers[11][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4398 )
         );
  MUX \Reg_Bank/U4442  ( .IN0(\Reg_Bank/n4396 ), .IN1(\Reg_Bank/n4395 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4397 ) );
  MUX \Reg_Bank/U4441  ( .IN0(\Reg_Bank/registers[12][12] ), .IN1(
        \Reg_Bank/registers[13][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4396 )
         );
  MUX \Reg_Bank/U4440  ( .IN0(\Reg_Bank/registers[14][12] ), .IN1(
        \Reg_Bank/registers[15][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4395 )
         );
  MUX \Reg_Bank/U4439  ( .IN0(\Reg_Bank/n4393 ), .IN1(\Reg_Bank/n4386 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4394 ) );
  MUX \Reg_Bank/U4438  ( .IN0(\Reg_Bank/n4392 ), .IN1(\Reg_Bank/n4389 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4393 ) );
  MUX \Reg_Bank/U4437  ( .IN0(\Reg_Bank/n4391 ), .IN1(\Reg_Bank/n4390 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4392 ) );
  MUX \Reg_Bank/U4436  ( .IN0(\Reg_Bank/registers[16][12] ), .IN1(
        \Reg_Bank/registers[17][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4391 )
         );
  MUX \Reg_Bank/U4435  ( .IN0(\Reg_Bank/registers[18][12] ), .IN1(
        \Reg_Bank/registers[19][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4390 )
         );
  MUX \Reg_Bank/U4434  ( .IN0(\Reg_Bank/n4388 ), .IN1(\Reg_Bank/n4387 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4389 ) );
  MUX \Reg_Bank/U4433  ( .IN0(\Reg_Bank/registers[20][12] ), .IN1(
        \Reg_Bank/registers[21][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4388 )
         );
  MUX \Reg_Bank/U4432  ( .IN0(\Reg_Bank/registers[22][12] ), .IN1(
        \Reg_Bank/registers[23][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4387 )
         );
  MUX \Reg_Bank/U4431  ( .IN0(\Reg_Bank/n4385 ), .IN1(\Reg_Bank/n4382 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4386 ) );
  MUX \Reg_Bank/U4430  ( .IN0(\Reg_Bank/n4384 ), .IN1(\Reg_Bank/n4383 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4385 ) );
  MUX \Reg_Bank/U4429  ( .IN0(\Reg_Bank/registers[24][12] ), .IN1(
        \Reg_Bank/registers[25][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4384 )
         );
  MUX \Reg_Bank/U4428  ( .IN0(\Reg_Bank/registers[26][12] ), .IN1(
        \Reg_Bank/registers[27][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4383 )
         );
  MUX \Reg_Bank/U4427  ( .IN0(\Reg_Bank/n4381 ), .IN1(\Reg_Bank/n4380 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4382 ) );
  MUX \Reg_Bank/U4426  ( .IN0(\Reg_Bank/registers[28][12] ), .IN1(
        \Reg_Bank/registers[29][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4381 )
         );
  MUX \Reg_Bank/U4425  ( .IN0(\Reg_Bank/registers[30][12] ), .IN1(
        \Reg_Bank/registers[31][12] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4380 )
         );
  MUX \Reg_Bank/U4424  ( .IN0(\Reg_Bank/n4379 ), .IN1(\Reg_Bank/n4364 ), .SEL(
        rs_index[4]), .F(reg_source[11]) );
  MUX \Reg_Bank/U4423  ( .IN0(\Reg_Bank/n4378 ), .IN1(\Reg_Bank/n4371 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4379 ) );
  MUX \Reg_Bank/U4422  ( .IN0(\Reg_Bank/n4377 ), .IN1(\Reg_Bank/n4374 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4378 ) );
  MUX \Reg_Bank/U4421  ( .IN0(\Reg_Bank/n4376 ), .IN1(\Reg_Bank/n4375 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4377 ) );
  MUX \Reg_Bank/U4419  ( .IN0(\Reg_Bank/registers[2][11] ), .IN1(
        \Reg_Bank/registers[3][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4375 )
         );
  MUX \Reg_Bank/U4418  ( .IN0(\Reg_Bank/n4373 ), .IN1(\Reg_Bank/n4372 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4374 ) );
  MUX \Reg_Bank/U4417  ( .IN0(\Reg_Bank/registers[4][11] ), .IN1(
        \Reg_Bank/registers[5][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4373 )
         );
  MUX \Reg_Bank/U4416  ( .IN0(\Reg_Bank/registers[6][11] ), .IN1(
        \Reg_Bank/registers[7][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4372 )
         );
  MUX \Reg_Bank/U4415  ( .IN0(\Reg_Bank/n4370 ), .IN1(\Reg_Bank/n4367 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4371 ) );
  MUX \Reg_Bank/U4414  ( .IN0(\Reg_Bank/n4369 ), .IN1(\Reg_Bank/n4368 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4370 ) );
  MUX \Reg_Bank/U4413  ( .IN0(\Reg_Bank/registers[8][11] ), .IN1(
        \Reg_Bank/registers[9][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4369 )
         );
  MUX \Reg_Bank/U4412  ( .IN0(\Reg_Bank/registers[10][11] ), .IN1(
        \Reg_Bank/registers[11][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4368 )
         );
  MUX \Reg_Bank/U4411  ( .IN0(\Reg_Bank/n4366 ), .IN1(\Reg_Bank/n4365 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4367 ) );
  MUX \Reg_Bank/U4410  ( .IN0(\Reg_Bank/registers[12][11] ), .IN1(
        \Reg_Bank/registers[13][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4366 )
         );
  MUX \Reg_Bank/U4409  ( .IN0(\Reg_Bank/registers[14][11] ), .IN1(
        \Reg_Bank/registers[15][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4365 )
         );
  MUX \Reg_Bank/U4408  ( .IN0(\Reg_Bank/n4363 ), .IN1(\Reg_Bank/n4356 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4364 ) );
  MUX \Reg_Bank/U4407  ( .IN0(\Reg_Bank/n4362 ), .IN1(\Reg_Bank/n4359 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4363 ) );
  MUX \Reg_Bank/U4406  ( .IN0(\Reg_Bank/n4361 ), .IN1(\Reg_Bank/n4360 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4362 ) );
  MUX \Reg_Bank/U4405  ( .IN0(\Reg_Bank/registers[16][11] ), .IN1(
        \Reg_Bank/registers[17][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4361 )
         );
  MUX \Reg_Bank/U4404  ( .IN0(\Reg_Bank/registers[18][11] ), .IN1(
        \Reg_Bank/registers[19][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4360 )
         );
  MUX \Reg_Bank/U4403  ( .IN0(\Reg_Bank/n4358 ), .IN1(\Reg_Bank/n4357 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4359 ) );
  MUX \Reg_Bank/U4402  ( .IN0(\Reg_Bank/registers[20][11] ), .IN1(
        \Reg_Bank/registers[21][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4358 )
         );
  MUX \Reg_Bank/U4401  ( .IN0(\Reg_Bank/registers[22][11] ), .IN1(
        \Reg_Bank/registers[23][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4357 )
         );
  MUX \Reg_Bank/U4400  ( .IN0(\Reg_Bank/n4355 ), .IN1(\Reg_Bank/n4352 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4356 ) );
  MUX \Reg_Bank/U4399  ( .IN0(\Reg_Bank/n4354 ), .IN1(\Reg_Bank/n4353 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4355 ) );
  MUX \Reg_Bank/U4398  ( .IN0(\Reg_Bank/registers[24][11] ), .IN1(
        \Reg_Bank/registers[25][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4354 )
         );
  MUX \Reg_Bank/U4397  ( .IN0(\Reg_Bank/registers[26][11] ), .IN1(
        \Reg_Bank/registers[27][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4353 )
         );
  MUX \Reg_Bank/U4396  ( .IN0(\Reg_Bank/n4351 ), .IN1(\Reg_Bank/n4350 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4352 ) );
  MUX \Reg_Bank/U4395  ( .IN0(\Reg_Bank/registers[28][11] ), .IN1(
        \Reg_Bank/registers[29][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4351 )
         );
  MUX \Reg_Bank/U4394  ( .IN0(\Reg_Bank/registers[30][11] ), .IN1(
        \Reg_Bank/registers[31][11] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4350 )
         );
  MUX \Reg_Bank/U4393  ( .IN0(\Reg_Bank/n4349 ), .IN1(\Reg_Bank/n4334 ), .SEL(
        rs_index[4]), .F(reg_source[10]) );
  MUX \Reg_Bank/U4392  ( .IN0(\Reg_Bank/n4348 ), .IN1(\Reg_Bank/n4341 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4349 ) );
  MUX \Reg_Bank/U4391  ( .IN0(\Reg_Bank/n4347 ), .IN1(\Reg_Bank/n4344 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4348 ) );
  MUX \Reg_Bank/U4390  ( .IN0(\Reg_Bank/n4346 ), .IN1(\Reg_Bank/n4345 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4347 ) );
  MUX \Reg_Bank/U4388  ( .IN0(\Reg_Bank/registers[2][10] ), .IN1(
        \Reg_Bank/registers[3][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4345 )
         );
  MUX \Reg_Bank/U4387  ( .IN0(\Reg_Bank/n4343 ), .IN1(\Reg_Bank/n4342 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4344 ) );
  MUX \Reg_Bank/U4386  ( .IN0(\Reg_Bank/registers[4][10] ), .IN1(
        \Reg_Bank/registers[5][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4343 )
         );
  MUX \Reg_Bank/U4385  ( .IN0(\Reg_Bank/registers[6][10] ), .IN1(
        \Reg_Bank/registers[7][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4342 )
         );
  MUX \Reg_Bank/U4384  ( .IN0(\Reg_Bank/n4340 ), .IN1(\Reg_Bank/n4337 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4341 ) );
  MUX \Reg_Bank/U4383  ( .IN0(\Reg_Bank/n4339 ), .IN1(\Reg_Bank/n4338 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4340 ) );
  MUX \Reg_Bank/U4382  ( .IN0(\Reg_Bank/registers[8][10] ), .IN1(
        \Reg_Bank/registers[9][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4339 )
         );
  MUX \Reg_Bank/U4381  ( .IN0(\Reg_Bank/registers[10][10] ), .IN1(
        \Reg_Bank/registers[11][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4338 )
         );
  MUX \Reg_Bank/U4380  ( .IN0(\Reg_Bank/n4336 ), .IN1(\Reg_Bank/n4335 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4337 ) );
  MUX \Reg_Bank/U4379  ( .IN0(\Reg_Bank/registers[12][10] ), .IN1(
        \Reg_Bank/registers[13][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4336 )
         );
  MUX \Reg_Bank/U4378  ( .IN0(\Reg_Bank/registers[14][10] ), .IN1(
        \Reg_Bank/registers[15][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4335 )
         );
  MUX \Reg_Bank/U4377  ( .IN0(\Reg_Bank/n4333 ), .IN1(\Reg_Bank/n4326 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4334 ) );
  MUX \Reg_Bank/U4376  ( .IN0(\Reg_Bank/n4332 ), .IN1(\Reg_Bank/n4329 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4333 ) );
  MUX \Reg_Bank/U4375  ( .IN0(\Reg_Bank/n4331 ), .IN1(\Reg_Bank/n4330 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4332 ) );
  MUX \Reg_Bank/U4374  ( .IN0(\Reg_Bank/registers[16][10] ), .IN1(
        \Reg_Bank/registers[17][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4331 )
         );
  MUX \Reg_Bank/U4373  ( .IN0(\Reg_Bank/registers[18][10] ), .IN1(
        \Reg_Bank/registers[19][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4330 )
         );
  MUX \Reg_Bank/U4372  ( .IN0(\Reg_Bank/n4328 ), .IN1(\Reg_Bank/n4327 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4329 ) );
  MUX \Reg_Bank/U4371  ( .IN0(\Reg_Bank/registers[20][10] ), .IN1(
        \Reg_Bank/registers[21][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4328 )
         );
  MUX \Reg_Bank/U4370  ( .IN0(\Reg_Bank/registers[22][10] ), .IN1(
        \Reg_Bank/registers[23][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4327 )
         );
  MUX \Reg_Bank/U4369  ( .IN0(\Reg_Bank/n4325 ), .IN1(\Reg_Bank/n4322 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4326 ) );
  MUX \Reg_Bank/U4368  ( .IN0(\Reg_Bank/n4324 ), .IN1(\Reg_Bank/n4323 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4325 ) );
  MUX \Reg_Bank/U4367  ( .IN0(\Reg_Bank/registers[24][10] ), .IN1(
        \Reg_Bank/registers[25][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4324 )
         );
  MUX \Reg_Bank/U4366  ( .IN0(\Reg_Bank/registers[26][10] ), .IN1(
        \Reg_Bank/registers[27][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4323 )
         );
  MUX \Reg_Bank/U4365  ( .IN0(\Reg_Bank/n4321 ), .IN1(\Reg_Bank/n4320 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4322 ) );
  MUX \Reg_Bank/U4364  ( .IN0(\Reg_Bank/registers[28][10] ), .IN1(
        \Reg_Bank/registers[29][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4321 )
         );
  MUX \Reg_Bank/U4363  ( .IN0(\Reg_Bank/registers[30][10] ), .IN1(
        \Reg_Bank/registers[31][10] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4320 )
         );
  MUX \Reg_Bank/U4362  ( .IN0(\Reg_Bank/n4319 ), .IN1(\Reg_Bank/n4304 ), .SEL(
        rs_index[4]), .F(reg_source[9]) );
  MUX \Reg_Bank/U4361  ( .IN0(\Reg_Bank/n4318 ), .IN1(\Reg_Bank/n4311 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4319 ) );
  MUX \Reg_Bank/U4360  ( .IN0(\Reg_Bank/n4317 ), .IN1(\Reg_Bank/n4314 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4318 ) );
  MUX \Reg_Bank/U4359  ( .IN0(\Reg_Bank/n4316 ), .IN1(\Reg_Bank/n4315 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4317 ) );
  MUX \Reg_Bank/U4357  ( .IN0(\Reg_Bank/registers[2][9] ), .IN1(
        \Reg_Bank/registers[3][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4315 )
         );
  MUX \Reg_Bank/U4356  ( .IN0(\Reg_Bank/n4313 ), .IN1(\Reg_Bank/n4312 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4314 ) );
  MUX \Reg_Bank/U4355  ( .IN0(\Reg_Bank/registers[4][9] ), .IN1(
        \Reg_Bank/registers[5][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4313 )
         );
  MUX \Reg_Bank/U4354  ( .IN0(\Reg_Bank/registers[6][9] ), .IN1(
        \Reg_Bank/registers[7][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4312 )
         );
  MUX \Reg_Bank/U4353  ( .IN0(\Reg_Bank/n4310 ), .IN1(\Reg_Bank/n4307 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4311 ) );
  MUX \Reg_Bank/U4352  ( .IN0(\Reg_Bank/n4309 ), .IN1(\Reg_Bank/n4308 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4310 ) );
  MUX \Reg_Bank/U4351  ( .IN0(\Reg_Bank/registers[8][9] ), .IN1(
        \Reg_Bank/registers[9][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4309 )
         );
  MUX \Reg_Bank/U4350  ( .IN0(\Reg_Bank/registers[10][9] ), .IN1(
        \Reg_Bank/registers[11][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4308 )
         );
  MUX \Reg_Bank/U4349  ( .IN0(\Reg_Bank/n4306 ), .IN1(\Reg_Bank/n4305 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4307 ) );
  MUX \Reg_Bank/U4348  ( .IN0(\Reg_Bank/registers[12][9] ), .IN1(
        \Reg_Bank/registers[13][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4306 )
         );
  MUX \Reg_Bank/U4347  ( .IN0(\Reg_Bank/registers[14][9] ), .IN1(
        \Reg_Bank/registers[15][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4305 )
         );
  MUX \Reg_Bank/U4346  ( .IN0(\Reg_Bank/n4303 ), .IN1(\Reg_Bank/n4296 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4304 ) );
  MUX \Reg_Bank/U4345  ( .IN0(\Reg_Bank/n4302 ), .IN1(\Reg_Bank/n4299 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4303 ) );
  MUX \Reg_Bank/U4344  ( .IN0(\Reg_Bank/n4301 ), .IN1(\Reg_Bank/n4300 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4302 ) );
  MUX \Reg_Bank/U4343  ( .IN0(\Reg_Bank/registers[16][9] ), .IN1(
        \Reg_Bank/registers[17][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4301 )
         );
  MUX \Reg_Bank/U4342  ( .IN0(\Reg_Bank/registers[18][9] ), .IN1(
        \Reg_Bank/registers[19][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4300 )
         );
  MUX \Reg_Bank/U4341  ( .IN0(\Reg_Bank/n4298 ), .IN1(\Reg_Bank/n4297 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4299 ) );
  MUX \Reg_Bank/U4340  ( .IN0(\Reg_Bank/registers[20][9] ), .IN1(
        \Reg_Bank/registers[21][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4298 )
         );
  MUX \Reg_Bank/U4339  ( .IN0(\Reg_Bank/registers[22][9] ), .IN1(
        \Reg_Bank/registers[23][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4297 )
         );
  MUX \Reg_Bank/U4338  ( .IN0(\Reg_Bank/n4295 ), .IN1(\Reg_Bank/n4292 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4296 ) );
  MUX \Reg_Bank/U4337  ( .IN0(\Reg_Bank/n4294 ), .IN1(\Reg_Bank/n4293 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4295 ) );
  MUX \Reg_Bank/U4336  ( .IN0(\Reg_Bank/registers[24][9] ), .IN1(
        \Reg_Bank/registers[25][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4294 )
         );
  MUX \Reg_Bank/U4335  ( .IN0(\Reg_Bank/registers[26][9] ), .IN1(
        \Reg_Bank/registers[27][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4293 )
         );
  MUX \Reg_Bank/U4334  ( .IN0(\Reg_Bank/n4291 ), .IN1(\Reg_Bank/n4290 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4292 ) );
  MUX \Reg_Bank/U4333  ( .IN0(\Reg_Bank/registers[28][9] ), .IN1(
        \Reg_Bank/registers[29][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4291 )
         );
  MUX \Reg_Bank/U4332  ( .IN0(\Reg_Bank/registers[30][9] ), .IN1(
        \Reg_Bank/registers[31][9] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4290 )
         );
  MUX \Reg_Bank/U4331  ( .IN0(\Reg_Bank/n4289 ), .IN1(\Reg_Bank/n4274 ), .SEL(
        rs_index[4]), .F(reg_source[8]) );
  MUX \Reg_Bank/U4330  ( .IN0(\Reg_Bank/n4288 ), .IN1(\Reg_Bank/n4281 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4289 ) );
  MUX \Reg_Bank/U4329  ( .IN0(\Reg_Bank/n4287 ), .IN1(\Reg_Bank/n4284 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4288 ) );
  MUX \Reg_Bank/U4328  ( .IN0(\Reg_Bank/n4286 ), .IN1(\Reg_Bank/n4285 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4287 ) );
  MUX \Reg_Bank/U4326  ( .IN0(\Reg_Bank/registers[2][8] ), .IN1(
        \Reg_Bank/registers[3][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4285 )
         );
  MUX \Reg_Bank/U4325  ( .IN0(\Reg_Bank/n4283 ), .IN1(\Reg_Bank/n4282 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4284 ) );
  MUX \Reg_Bank/U4324  ( .IN0(\Reg_Bank/registers[4][8] ), .IN1(
        \Reg_Bank/registers[5][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4283 )
         );
  MUX \Reg_Bank/U4323  ( .IN0(\Reg_Bank/registers[6][8] ), .IN1(
        \Reg_Bank/registers[7][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4282 )
         );
  MUX \Reg_Bank/U4322  ( .IN0(\Reg_Bank/n4280 ), .IN1(\Reg_Bank/n4277 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4281 ) );
  MUX \Reg_Bank/U4321  ( .IN0(\Reg_Bank/n4279 ), .IN1(\Reg_Bank/n4278 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4280 ) );
  MUX \Reg_Bank/U4320  ( .IN0(\Reg_Bank/registers[8][8] ), .IN1(
        \Reg_Bank/registers[9][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4279 )
         );
  MUX \Reg_Bank/U4319  ( .IN0(\Reg_Bank/registers[10][8] ), .IN1(
        \Reg_Bank/registers[11][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4278 )
         );
  MUX \Reg_Bank/U4318  ( .IN0(\Reg_Bank/n4276 ), .IN1(\Reg_Bank/n4275 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4277 ) );
  MUX \Reg_Bank/U4317  ( .IN0(\Reg_Bank/registers[12][8] ), .IN1(
        \Reg_Bank/registers[13][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4276 )
         );
  MUX \Reg_Bank/U4316  ( .IN0(\Reg_Bank/registers[14][8] ), .IN1(
        \Reg_Bank/registers[15][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4275 )
         );
  MUX \Reg_Bank/U4315  ( .IN0(\Reg_Bank/n4273 ), .IN1(\Reg_Bank/n4266 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4274 ) );
  MUX \Reg_Bank/U4314  ( .IN0(\Reg_Bank/n4272 ), .IN1(\Reg_Bank/n4269 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4273 ) );
  MUX \Reg_Bank/U4313  ( .IN0(\Reg_Bank/n4271 ), .IN1(\Reg_Bank/n4270 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4272 ) );
  MUX \Reg_Bank/U4312  ( .IN0(\Reg_Bank/registers[16][8] ), .IN1(
        \Reg_Bank/registers[17][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4271 )
         );
  MUX \Reg_Bank/U4311  ( .IN0(\Reg_Bank/registers[18][8] ), .IN1(
        \Reg_Bank/registers[19][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4270 )
         );
  MUX \Reg_Bank/U4310  ( .IN0(\Reg_Bank/n4268 ), .IN1(\Reg_Bank/n4267 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4269 ) );
  MUX \Reg_Bank/U4309  ( .IN0(\Reg_Bank/registers[20][8] ), .IN1(
        \Reg_Bank/registers[21][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4268 )
         );
  MUX \Reg_Bank/U4308  ( .IN0(\Reg_Bank/registers[22][8] ), .IN1(
        \Reg_Bank/registers[23][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4267 )
         );
  MUX \Reg_Bank/U4307  ( .IN0(\Reg_Bank/n4265 ), .IN1(\Reg_Bank/n4262 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4266 ) );
  MUX \Reg_Bank/U4306  ( .IN0(\Reg_Bank/n4264 ), .IN1(\Reg_Bank/n4263 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4265 ) );
  MUX \Reg_Bank/U4305  ( .IN0(\Reg_Bank/registers[24][8] ), .IN1(
        \Reg_Bank/registers[25][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4264 )
         );
  MUX \Reg_Bank/U4304  ( .IN0(\Reg_Bank/registers[26][8] ), .IN1(
        \Reg_Bank/registers[27][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4263 )
         );
  MUX \Reg_Bank/U4303  ( .IN0(\Reg_Bank/n4261 ), .IN1(\Reg_Bank/n4260 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4262 ) );
  MUX \Reg_Bank/U4302  ( .IN0(\Reg_Bank/registers[28][8] ), .IN1(
        \Reg_Bank/registers[29][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4261 )
         );
  MUX \Reg_Bank/U4301  ( .IN0(\Reg_Bank/registers[30][8] ), .IN1(
        \Reg_Bank/registers[31][8] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4260 )
         );
  MUX \Reg_Bank/U4300  ( .IN0(\Reg_Bank/n4259 ), .IN1(\Reg_Bank/n4244 ), .SEL(
        rs_index[4]), .F(reg_source[7]) );
  MUX \Reg_Bank/U4299  ( .IN0(\Reg_Bank/n4258 ), .IN1(\Reg_Bank/n4251 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4259 ) );
  MUX \Reg_Bank/U4298  ( .IN0(\Reg_Bank/n4257 ), .IN1(\Reg_Bank/n4254 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4258 ) );
  MUX \Reg_Bank/U4297  ( .IN0(\Reg_Bank/n4256 ), .IN1(\Reg_Bank/n4255 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4257 ) );
  MUX \Reg_Bank/U4295  ( .IN0(\Reg_Bank/registers[2][7] ), .IN1(
        \Reg_Bank/registers[3][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4255 )
         );
  MUX \Reg_Bank/U4294  ( .IN0(\Reg_Bank/n4253 ), .IN1(\Reg_Bank/n4252 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4254 ) );
  MUX \Reg_Bank/U4293  ( .IN0(\Reg_Bank/registers[4][7] ), .IN1(
        \Reg_Bank/registers[5][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4253 )
         );
  MUX \Reg_Bank/U4292  ( .IN0(\Reg_Bank/registers[6][7] ), .IN1(
        \Reg_Bank/registers[7][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4252 )
         );
  MUX \Reg_Bank/U4291  ( .IN0(\Reg_Bank/n4250 ), .IN1(\Reg_Bank/n4247 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4251 ) );
  MUX \Reg_Bank/U4290  ( .IN0(\Reg_Bank/n4249 ), .IN1(\Reg_Bank/n4248 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4250 ) );
  MUX \Reg_Bank/U4289  ( .IN0(\Reg_Bank/registers[8][7] ), .IN1(
        \Reg_Bank/registers[9][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4249 )
         );
  MUX \Reg_Bank/U4288  ( .IN0(\Reg_Bank/registers[10][7] ), .IN1(
        \Reg_Bank/registers[11][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4248 )
         );
  MUX \Reg_Bank/U4287  ( .IN0(\Reg_Bank/n4246 ), .IN1(\Reg_Bank/n4245 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4247 ) );
  MUX \Reg_Bank/U4286  ( .IN0(\Reg_Bank/registers[12][7] ), .IN1(
        \Reg_Bank/registers[13][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4246 )
         );
  MUX \Reg_Bank/U4285  ( .IN0(\Reg_Bank/registers[14][7] ), .IN1(
        \Reg_Bank/registers[15][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4245 )
         );
  MUX \Reg_Bank/U4284  ( .IN0(\Reg_Bank/n4243 ), .IN1(\Reg_Bank/n4236 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4244 ) );
  MUX \Reg_Bank/U4283  ( .IN0(\Reg_Bank/n4242 ), .IN1(\Reg_Bank/n4239 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4243 ) );
  MUX \Reg_Bank/U4282  ( .IN0(\Reg_Bank/n4241 ), .IN1(\Reg_Bank/n4240 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4242 ) );
  MUX \Reg_Bank/U4281  ( .IN0(\Reg_Bank/registers[16][7] ), .IN1(
        \Reg_Bank/registers[17][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4241 )
         );
  MUX \Reg_Bank/U4280  ( .IN0(\Reg_Bank/registers[18][7] ), .IN1(
        \Reg_Bank/registers[19][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4240 )
         );
  MUX \Reg_Bank/U4279  ( .IN0(\Reg_Bank/n4238 ), .IN1(\Reg_Bank/n4237 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4239 ) );
  MUX \Reg_Bank/U4278  ( .IN0(\Reg_Bank/registers[20][7] ), .IN1(
        \Reg_Bank/registers[21][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4238 )
         );
  MUX \Reg_Bank/U4277  ( .IN0(\Reg_Bank/registers[22][7] ), .IN1(
        \Reg_Bank/registers[23][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4237 )
         );
  MUX \Reg_Bank/U4276  ( .IN0(\Reg_Bank/n4235 ), .IN1(\Reg_Bank/n4232 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4236 ) );
  MUX \Reg_Bank/U4275  ( .IN0(\Reg_Bank/n4234 ), .IN1(\Reg_Bank/n4233 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4235 ) );
  MUX \Reg_Bank/U4274  ( .IN0(\Reg_Bank/registers[24][7] ), .IN1(
        \Reg_Bank/registers[25][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4234 )
         );
  MUX \Reg_Bank/U4273  ( .IN0(\Reg_Bank/registers[26][7] ), .IN1(
        \Reg_Bank/registers[27][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4233 )
         );
  MUX \Reg_Bank/U4272  ( .IN0(\Reg_Bank/n4231 ), .IN1(\Reg_Bank/n4230 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4232 ) );
  MUX \Reg_Bank/U4271  ( .IN0(\Reg_Bank/registers[28][7] ), .IN1(
        \Reg_Bank/registers[29][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4231 )
         );
  MUX \Reg_Bank/U4270  ( .IN0(\Reg_Bank/registers[30][7] ), .IN1(
        \Reg_Bank/registers[31][7] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4230 )
         );
  MUX \Reg_Bank/U4269  ( .IN0(\Reg_Bank/n4229 ), .IN1(\Reg_Bank/n4214 ), .SEL(
        rs_index[4]), .F(reg_source[6]) );
  MUX \Reg_Bank/U4268  ( .IN0(\Reg_Bank/n4228 ), .IN1(\Reg_Bank/n4221 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4229 ) );
  MUX \Reg_Bank/U4267  ( .IN0(\Reg_Bank/n4227 ), .IN1(\Reg_Bank/n4224 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4228 ) );
  MUX \Reg_Bank/U4266  ( .IN0(\Reg_Bank/n4226 ), .IN1(\Reg_Bank/n4225 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4227 ) );
  MUX \Reg_Bank/U4264  ( .IN0(\Reg_Bank/registers[2][6] ), .IN1(
        \Reg_Bank/registers[3][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4225 )
         );
  MUX \Reg_Bank/U4263  ( .IN0(\Reg_Bank/n4223 ), .IN1(\Reg_Bank/n4222 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4224 ) );
  MUX \Reg_Bank/U4262  ( .IN0(\Reg_Bank/registers[4][6] ), .IN1(
        \Reg_Bank/registers[5][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4223 )
         );
  MUX \Reg_Bank/U4261  ( .IN0(\Reg_Bank/registers[6][6] ), .IN1(
        \Reg_Bank/registers[7][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4222 )
         );
  MUX \Reg_Bank/U4260  ( .IN0(\Reg_Bank/n4220 ), .IN1(\Reg_Bank/n4217 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4221 ) );
  MUX \Reg_Bank/U4259  ( .IN0(\Reg_Bank/n4219 ), .IN1(\Reg_Bank/n4218 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4220 ) );
  MUX \Reg_Bank/U4258  ( .IN0(\Reg_Bank/registers[8][6] ), .IN1(
        \Reg_Bank/registers[9][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4219 )
         );
  MUX \Reg_Bank/U4257  ( .IN0(\Reg_Bank/registers[10][6] ), .IN1(
        \Reg_Bank/registers[11][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4218 )
         );
  MUX \Reg_Bank/U4256  ( .IN0(\Reg_Bank/n4216 ), .IN1(\Reg_Bank/n4215 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4217 ) );
  MUX \Reg_Bank/U4255  ( .IN0(\Reg_Bank/registers[12][6] ), .IN1(
        \Reg_Bank/registers[13][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4216 )
         );
  MUX \Reg_Bank/U4254  ( .IN0(\Reg_Bank/registers[14][6] ), .IN1(
        \Reg_Bank/registers[15][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4215 )
         );
  MUX \Reg_Bank/U4253  ( .IN0(\Reg_Bank/n4213 ), .IN1(\Reg_Bank/n4206 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4214 ) );
  MUX \Reg_Bank/U4252  ( .IN0(\Reg_Bank/n4212 ), .IN1(\Reg_Bank/n4209 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4213 ) );
  MUX \Reg_Bank/U4251  ( .IN0(\Reg_Bank/n4211 ), .IN1(\Reg_Bank/n4210 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4212 ) );
  MUX \Reg_Bank/U4250  ( .IN0(\Reg_Bank/registers[16][6] ), .IN1(
        \Reg_Bank/registers[17][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4211 )
         );
  MUX \Reg_Bank/U4249  ( .IN0(\Reg_Bank/registers[18][6] ), .IN1(
        \Reg_Bank/registers[19][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4210 )
         );
  MUX \Reg_Bank/U4248  ( .IN0(\Reg_Bank/n4208 ), .IN1(\Reg_Bank/n4207 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4209 ) );
  MUX \Reg_Bank/U4247  ( .IN0(\Reg_Bank/registers[20][6] ), .IN1(
        \Reg_Bank/registers[21][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4208 )
         );
  MUX \Reg_Bank/U4246  ( .IN0(\Reg_Bank/registers[22][6] ), .IN1(
        \Reg_Bank/registers[23][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4207 )
         );
  MUX \Reg_Bank/U4245  ( .IN0(\Reg_Bank/n4205 ), .IN1(\Reg_Bank/n4202 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4206 ) );
  MUX \Reg_Bank/U4244  ( .IN0(\Reg_Bank/n4204 ), .IN1(\Reg_Bank/n4203 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4205 ) );
  MUX \Reg_Bank/U4243  ( .IN0(\Reg_Bank/registers[24][6] ), .IN1(
        \Reg_Bank/registers[25][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4204 )
         );
  MUX \Reg_Bank/U4242  ( .IN0(\Reg_Bank/registers[26][6] ), .IN1(
        \Reg_Bank/registers[27][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4203 )
         );
  MUX \Reg_Bank/U4241  ( .IN0(\Reg_Bank/n4201 ), .IN1(\Reg_Bank/n4200 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4202 ) );
  MUX \Reg_Bank/U4240  ( .IN0(\Reg_Bank/registers[28][6] ), .IN1(
        \Reg_Bank/registers[29][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4201 )
         );
  MUX \Reg_Bank/U4239  ( .IN0(\Reg_Bank/registers[30][6] ), .IN1(
        \Reg_Bank/registers[31][6] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4200 )
         );
  MUX \Reg_Bank/U4238  ( .IN0(\Reg_Bank/n4199 ), .IN1(\Reg_Bank/n4184 ), .SEL(
        rs_index[4]), .F(reg_source[5]) );
  MUX \Reg_Bank/U4237  ( .IN0(\Reg_Bank/n4198 ), .IN1(\Reg_Bank/n4191 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4199 ) );
  MUX \Reg_Bank/U4236  ( .IN0(\Reg_Bank/n4197 ), .IN1(\Reg_Bank/n4194 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4198 ) );
  MUX \Reg_Bank/U4235  ( .IN0(\Reg_Bank/n4196 ), .IN1(\Reg_Bank/n4195 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4197 ) );
  MUX \Reg_Bank/U4233  ( .IN0(\Reg_Bank/registers[2][5] ), .IN1(
        \Reg_Bank/registers[3][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4195 )
         );
  MUX \Reg_Bank/U4232  ( .IN0(\Reg_Bank/n4193 ), .IN1(\Reg_Bank/n4192 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4194 ) );
  MUX \Reg_Bank/U4231  ( .IN0(\Reg_Bank/registers[4][5] ), .IN1(
        \Reg_Bank/registers[5][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4193 )
         );
  MUX \Reg_Bank/U4230  ( .IN0(\Reg_Bank/registers[6][5] ), .IN1(
        \Reg_Bank/registers[7][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4192 )
         );
  MUX \Reg_Bank/U4229  ( .IN0(\Reg_Bank/n4190 ), .IN1(\Reg_Bank/n4187 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4191 ) );
  MUX \Reg_Bank/U4228  ( .IN0(\Reg_Bank/n4189 ), .IN1(\Reg_Bank/n4188 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4190 ) );
  MUX \Reg_Bank/U4227  ( .IN0(\Reg_Bank/registers[8][5] ), .IN1(
        \Reg_Bank/registers[9][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4189 )
         );
  MUX \Reg_Bank/U4226  ( .IN0(\Reg_Bank/registers[10][5] ), .IN1(
        \Reg_Bank/registers[11][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4188 )
         );
  MUX \Reg_Bank/U4225  ( .IN0(\Reg_Bank/n4186 ), .IN1(\Reg_Bank/n4185 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4187 ) );
  MUX \Reg_Bank/U4224  ( .IN0(\Reg_Bank/registers[12][5] ), .IN1(
        \Reg_Bank/registers[13][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4186 )
         );
  MUX \Reg_Bank/U4223  ( .IN0(\Reg_Bank/registers[14][5] ), .IN1(
        \Reg_Bank/registers[15][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4185 )
         );
  MUX \Reg_Bank/U4222  ( .IN0(\Reg_Bank/n4183 ), .IN1(\Reg_Bank/n4176 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4184 ) );
  MUX \Reg_Bank/U4221  ( .IN0(\Reg_Bank/n4182 ), .IN1(\Reg_Bank/n4179 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4183 ) );
  MUX \Reg_Bank/U4220  ( .IN0(\Reg_Bank/n4181 ), .IN1(\Reg_Bank/n4180 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4182 ) );
  MUX \Reg_Bank/U4219  ( .IN0(\Reg_Bank/registers[16][5] ), .IN1(
        \Reg_Bank/registers[17][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4181 )
         );
  MUX \Reg_Bank/U4218  ( .IN0(\Reg_Bank/registers[18][5] ), .IN1(
        \Reg_Bank/registers[19][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4180 )
         );
  MUX \Reg_Bank/U4217  ( .IN0(\Reg_Bank/n4178 ), .IN1(\Reg_Bank/n4177 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4179 ) );
  MUX \Reg_Bank/U4216  ( .IN0(\Reg_Bank/registers[20][5] ), .IN1(
        \Reg_Bank/registers[21][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4178 )
         );
  MUX \Reg_Bank/U4215  ( .IN0(\Reg_Bank/registers[22][5] ), .IN1(
        \Reg_Bank/registers[23][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4177 )
         );
  MUX \Reg_Bank/U4214  ( .IN0(\Reg_Bank/n4175 ), .IN1(\Reg_Bank/n4172 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4176 ) );
  MUX \Reg_Bank/U4213  ( .IN0(\Reg_Bank/n4174 ), .IN1(\Reg_Bank/n4173 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4175 ) );
  MUX \Reg_Bank/U4212  ( .IN0(\Reg_Bank/registers[24][5] ), .IN1(
        \Reg_Bank/registers[25][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4174 )
         );
  MUX \Reg_Bank/U4211  ( .IN0(\Reg_Bank/registers[26][5] ), .IN1(
        \Reg_Bank/registers[27][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4173 )
         );
  MUX \Reg_Bank/U4210  ( .IN0(\Reg_Bank/n4171 ), .IN1(\Reg_Bank/n4170 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4172 ) );
  MUX \Reg_Bank/U4209  ( .IN0(\Reg_Bank/registers[28][5] ), .IN1(
        \Reg_Bank/registers[29][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4171 )
         );
  MUX \Reg_Bank/U4208  ( .IN0(\Reg_Bank/registers[30][5] ), .IN1(
        \Reg_Bank/registers[31][5] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4170 )
         );
  MUX \Reg_Bank/U4207  ( .IN0(\Reg_Bank/n4169 ), .IN1(\Reg_Bank/n4154 ), .SEL(
        rs_index[4]), .F(reg_source[4]) );
  MUX \Reg_Bank/U4206  ( .IN0(\Reg_Bank/n4168 ), .IN1(\Reg_Bank/n4161 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4169 ) );
  MUX \Reg_Bank/U4205  ( .IN0(\Reg_Bank/n4167 ), .IN1(\Reg_Bank/n4164 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4168 ) );
  MUX \Reg_Bank/U4204  ( .IN0(\Reg_Bank/n4166 ), .IN1(\Reg_Bank/n4165 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4167 ) );
  MUX \Reg_Bank/U4202  ( .IN0(\Reg_Bank/registers[2][4] ), .IN1(
        \Reg_Bank/registers[3][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4165 )
         );
  MUX \Reg_Bank/U4201  ( .IN0(\Reg_Bank/n4163 ), .IN1(\Reg_Bank/n4162 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4164 ) );
  MUX \Reg_Bank/U4200  ( .IN0(\Reg_Bank/registers[4][4] ), .IN1(
        \Reg_Bank/registers[5][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4163 )
         );
  MUX \Reg_Bank/U4199  ( .IN0(\Reg_Bank/registers[6][4] ), .IN1(
        \Reg_Bank/registers[7][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4162 )
         );
  MUX \Reg_Bank/U4198  ( .IN0(\Reg_Bank/n4160 ), .IN1(\Reg_Bank/n4157 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4161 ) );
  MUX \Reg_Bank/U4197  ( .IN0(\Reg_Bank/n4159 ), .IN1(\Reg_Bank/n4158 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4160 ) );
  MUX \Reg_Bank/U4196  ( .IN0(\Reg_Bank/registers[8][4] ), .IN1(
        \Reg_Bank/registers[9][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4159 )
         );
  MUX \Reg_Bank/U4195  ( .IN0(\Reg_Bank/registers[10][4] ), .IN1(
        \Reg_Bank/registers[11][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4158 )
         );
  MUX \Reg_Bank/U4194  ( .IN0(\Reg_Bank/n4156 ), .IN1(\Reg_Bank/n4155 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4157 ) );
  MUX \Reg_Bank/U4193  ( .IN0(\Reg_Bank/registers[12][4] ), .IN1(
        \Reg_Bank/registers[13][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4156 )
         );
  MUX \Reg_Bank/U4192  ( .IN0(\Reg_Bank/registers[14][4] ), .IN1(
        \Reg_Bank/registers[15][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4155 )
         );
  MUX \Reg_Bank/U4191  ( .IN0(\Reg_Bank/n4153 ), .IN1(\Reg_Bank/n4146 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4154 ) );
  MUX \Reg_Bank/U4190  ( .IN0(\Reg_Bank/n4152 ), .IN1(\Reg_Bank/n4149 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4153 ) );
  MUX \Reg_Bank/U4189  ( .IN0(\Reg_Bank/n4151 ), .IN1(\Reg_Bank/n4150 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4152 ) );
  MUX \Reg_Bank/U4188  ( .IN0(\Reg_Bank/registers[16][4] ), .IN1(
        \Reg_Bank/registers[17][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4151 )
         );
  MUX \Reg_Bank/U4187  ( .IN0(\Reg_Bank/registers[18][4] ), .IN1(
        \Reg_Bank/registers[19][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4150 )
         );
  MUX \Reg_Bank/U4186  ( .IN0(\Reg_Bank/n4148 ), .IN1(\Reg_Bank/n4147 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4149 ) );
  MUX \Reg_Bank/U4185  ( .IN0(\Reg_Bank/registers[20][4] ), .IN1(
        \Reg_Bank/registers[21][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4148 )
         );
  MUX \Reg_Bank/U4184  ( .IN0(\Reg_Bank/registers[22][4] ), .IN1(
        \Reg_Bank/registers[23][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4147 )
         );
  MUX \Reg_Bank/U4183  ( .IN0(\Reg_Bank/n4145 ), .IN1(\Reg_Bank/n4142 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4146 ) );
  MUX \Reg_Bank/U4182  ( .IN0(\Reg_Bank/n4144 ), .IN1(\Reg_Bank/n4143 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4145 ) );
  MUX \Reg_Bank/U4181  ( .IN0(\Reg_Bank/registers[24][4] ), .IN1(
        \Reg_Bank/registers[25][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4144 )
         );
  MUX \Reg_Bank/U4180  ( .IN0(\Reg_Bank/registers[26][4] ), .IN1(
        \Reg_Bank/registers[27][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4143 )
         );
  MUX \Reg_Bank/U4179  ( .IN0(\Reg_Bank/n4141 ), .IN1(\Reg_Bank/n4140 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4142 ) );
  MUX \Reg_Bank/U4178  ( .IN0(\Reg_Bank/registers[28][4] ), .IN1(
        \Reg_Bank/registers[29][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4141 )
         );
  MUX \Reg_Bank/U4177  ( .IN0(\Reg_Bank/registers[30][4] ), .IN1(
        \Reg_Bank/registers[31][4] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4140 )
         );
  MUX \Reg_Bank/U4176  ( .IN0(\Reg_Bank/n4139 ), .IN1(\Reg_Bank/n4124 ), .SEL(
        rs_index[4]), .F(reg_source[3]) );
  MUX \Reg_Bank/U4175  ( .IN0(\Reg_Bank/n4138 ), .IN1(\Reg_Bank/n4131 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4139 ) );
  MUX \Reg_Bank/U4174  ( .IN0(\Reg_Bank/n4137 ), .IN1(\Reg_Bank/n4134 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4138 ) );
  MUX \Reg_Bank/U4173  ( .IN0(\Reg_Bank/n4136 ), .IN1(\Reg_Bank/n4135 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4137 ) );
  MUX \Reg_Bank/U4171  ( .IN0(\Reg_Bank/registers[2][3] ), .IN1(
        \Reg_Bank/registers[3][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4135 )
         );
  MUX \Reg_Bank/U4170  ( .IN0(\Reg_Bank/n4133 ), .IN1(\Reg_Bank/n4132 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4134 ) );
  MUX \Reg_Bank/U4169  ( .IN0(\Reg_Bank/registers[4][3] ), .IN1(
        \Reg_Bank/registers[5][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4133 )
         );
  MUX \Reg_Bank/U4168  ( .IN0(\Reg_Bank/registers[6][3] ), .IN1(
        \Reg_Bank/registers[7][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4132 )
         );
  MUX \Reg_Bank/U4167  ( .IN0(\Reg_Bank/n4130 ), .IN1(\Reg_Bank/n4127 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4131 ) );
  MUX \Reg_Bank/U4166  ( .IN0(\Reg_Bank/n4129 ), .IN1(\Reg_Bank/n4128 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4130 ) );
  MUX \Reg_Bank/U4165  ( .IN0(\Reg_Bank/registers[8][3] ), .IN1(
        \Reg_Bank/registers[9][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4129 )
         );
  MUX \Reg_Bank/U4164  ( .IN0(\Reg_Bank/registers[10][3] ), .IN1(
        \Reg_Bank/registers[11][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4128 )
         );
  MUX \Reg_Bank/U4163  ( .IN0(\Reg_Bank/n4126 ), .IN1(\Reg_Bank/n4125 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4127 ) );
  MUX \Reg_Bank/U4162  ( .IN0(\Reg_Bank/registers[12][3] ), .IN1(
        \Reg_Bank/registers[13][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4126 )
         );
  MUX \Reg_Bank/U4161  ( .IN0(\Reg_Bank/registers[14][3] ), .IN1(
        \Reg_Bank/registers[15][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4125 )
         );
  MUX \Reg_Bank/U4160  ( .IN0(\Reg_Bank/n4123 ), .IN1(\Reg_Bank/n4116 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4124 ) );
  MUX \Reg_Bank/U4159  ( .IN0(\Reg_Bank/n4122 ), .IN1(\Reg_Bank/n4119 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4123 ) );
  MUX \Reg_Bank/U4158  ( .IN0(\Reg_Bank/n4121 ), .IN1(\Reg_Bank/n4120 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4122 ) );
  MUX \Reg_Bank/U4157  ( .IN0(\Reg_Bank/registers[16][3] ), .IN1(
        \Reg_Bank/registers[17][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4121 )
         );
  MUX \Reg_Bank/U4156  ( .IN0(\Reg_Bank/registers[18][3] ), .IN1(
        \Reg_Bank/registers[19][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4120 )
         );
  MUX \Reg_Bank/U4155  ( .IN0(\Reg_Bank/n4118 ), .IN1(\Reg_Bank/n4117 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4119 ) );
  MUX \Reg_Bank/U4154  ( .IN0(\Reg_Bank/registers[20][3] ), .IN1(
        \Reg_Bank/registers[21][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4118 )
         );
  MUX \Reg_Bank/U4153  ( .IN0(\Reg_Bank/registers[22][3] ), .IN1(
        \Reg_Bank/registers[23][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4117 )
         );
  MUX \Reg_Bank/U4152  ( .IN0(\Reg_Bank/n4115 ), .IN1(\Reg_Bank/n4112 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4116 ) );
  MUX \Reg_Bank/U4151  ( .IN0(\Reg_Bank/n4114 ), .IN1(\Reg_Bank/n4113 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4115 ) );
  MUX \Reg_Bank/U4150  ( .IN0(\Reg_Bank/registers[24][3] ), .IN1(
        \Reg_Bank/registers[25][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4114 )
         );
  MUX \Reg_Bank/U4149  ( .IN0(\Reg_Bank/registers[26][3] ), .IN1(
        \Reg_Bank/registers[27][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4113 )
         );
  MUX \Reg_Bank/U4148  ( .IN0(\Reg_Bank/n4111 ), .IN1(\Reg_Bank/n4110 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4112 ) );
  MUX \Reg_Bank/U4147  ( .IN0(\Reg_Bank/registers[28][3] ), .IN1(
        \Reg_Bank/registers[29][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4111 )
         );
  MUX \Reg_Bank/U4146  ( .IN0(\Reg_Bank/registers[30][3] ), .IN1(
        \Reg_Bank/registers[31][3] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4110 )
         );
  MUX \Reg_Bank/U4145  ( .IN0(\Reg_Bank/n4109 ), .IN1(\Reg_Bank/n4094 ), .SEL(
        rs_index[4]), .F(reg_source[2]) );
  MUX \Reg_Bank/U4144  ( .IN0(\Reg_Bank/n4108 ), .IN1(\Reg_Bank/n4101 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4109 ) );
  MUX \Reg_Bank/U4143  ( .IN0(\Reg_Bank/n4107 ), .IN1(\Reg_Bank/n4104 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4108 ) );
  MUX \Reg_Bank/U4142  ( .IN0(\Reg_Bank/n4106 ), .IN1(\Reg_Bank/n4105 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4107 ) );
  MUX \Reg_Bank/U4140  ( .IN0(\Reg_Bank/registers[2][2] ), .IN1(
        \Reg_Bank/registers[3][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4105 )
         );
  MUX \Reg_Bank/U4139  ( .IN0(\Reg_Bank/n4103 ), .IN1(\Reg_Bank/n4102 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4104 ) );
  MUX \Reg_Bank/U4138  ( .IN0(\Reg_Bank/registers[4][2] ), .IN1(
        \Reg_Bank/registers[5][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4103 )
         );
  MUX \Reg_Bank/U4137  ( .IN0(\Reg_Bank/registers[6][2] ), .IN1(
        \Reg_Bank/registers[7][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4102 )
         );
  MUX \Reg_Bank/U4136  ( .IN0(\Reg_Bank/n4100 ), .IN1(\Reg_Bank/n4097 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4101 ) );
  MUX \Reg_Bank/U4135  ( .IN0(\Reg_Bank/n4099 ), .IN1(\Reg_Bank/n4098 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4100 ) );
  MUX \Reg_Bank/U4134  ( .IN0(\Reg_Bank/registers[8][2] ), .IN1(
        \Reg_Bank/registers[9][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4099 )
         );
  MUX \Reg_Bank/U4133  ( .IN0(\Reg_Bank/registers[10][2] ), .IN1(
        \Reg_Bank/registers[11][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4098 )
         );
  MUX \Reg_Bank/U4132  ( .IN0(\Reg_Bank/n4096 ), .IN1(\Reg_Bank/n4095 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4097 ) );
  MUX \Reg_Bank/U4131  ( .IN0(\Reg_Bank/registers[12][2] ), .IN1(
        \Reg_Bank/registers[13][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4096 )
         );
  MUX \Reg_Bank/U4130  ( .IN0(\Reg_Bank/registers[14][2] ), .IN1(
        \Reg_Bank/registers[15][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4095 )
         );
  MUX \Reg_Bank/U4129  ( .IN0(\Reg_Bank/n4093 ), .IN1(\Reg_Bank/n4086 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4094 ) );
  MUX \Reg_Bank/U4128  ( .IN0(\Reg_Bank/n4092 ), .IN1(\Reg_Bank/n4089 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4093 ) );
  MUX \Reg_Bank/U4127  ( .IN0(\Reg_Bank/n4091 ), .IN1(\Reg_Bank/n4090 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4092 ) );
  MUX \Reg_Bank/U4126  ( .IN0(\Reg_Bank/registers[16][2] ), .IN1(
        \Reg_Bank/registers[17][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4091 )
         );
  MUX \Reg_Bank/U4125  ( .IN0(\Reg_Bank/registers[18][2] ), .IN1(
        \Reg_Bank/registers[19][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4090 )
         );
  MUX \Reg_Bank/U4124  ( .IN0(\Reg_Bank/n4088 ), .IN1(\Reg_Bank/n4087 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4089 ) );
  MUX \Reg_Bank/U4123  ( .IN0(\Reg_Bank/registers[20][2] ), .IN1(
        \Reg_Bank/registers[21][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4088 )
         );
  MUX \Reg_Bank/U4122  ( .IN0(\Reg_Bank/registers[22][2] ), .IN1(
        \Reg_Bank/registers[23][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4087 )
         );
  MUX \Reg_Bank/U4121  ( .IN0(\Reg_Bank/n4085 ), .IN1(\Reg_Bank/n4082 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4086 ) );
  MUX \Reg_Bank/U4120  ( .IN0(\Reg_Bank/n4084 ), .IN1(\Reg_Bank/n4083 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4085 ) );
  MUX \Reg_Bank/U4119  ( .IN0(\Reg_Bank/registers[24][2] ), .IN1(
        \Reg_Bank/registers[25][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4084 )
         );
  MUX \Reg_Bank/U4118  ( .IN0(\Reg_Bank/registers[26][2] ), .IN1(
        \Reg_Bank/registers[27][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4083 )
         );
  MUX \Reg_Bank/U4117  ( .IN0(\Reg_Bank/n4081 ), .IN1(\Reg_Bank/n4080 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4082 ) );
  MUX \Reg_Bank/U4116  ( .IN0(\Reg_Bank/registers[28][2] ), .IN1(
        \Reg_Bank/registers[29][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4081 )
         );
  MUX \Reg_Bank/U4115  ( .IN0(\Reg_Bank/registers[30][2] ), .IN1(
        \Reg_Bank/registers[31][2] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4080 )
         );
  MUX \Reg_Bank/U4114  ( .IN0(\Reg_Bank/n4079 ), .IN1(\Reg_Bank/n4064 ), .SEL(
        rs_index[4]), .F(reg_source[1]) );
  MUX \Reg_Bank/U4113  ( .IN0(\Reg_Bank/n4078 ), .IN1(\Reg_Bank/n4071 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4079 ) );
  MUX \Reg_Bank/U4112  ( .IN0(\Reg_Bank/n4077 ), .IN1(\Reg_Bank/n4074 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4078 ) );
  MUX \Reg_Bank/U4111  ( .IN0(\Reg_Bank/n4076 ), .IN1(\Reg_Bank/n4075 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4077 ) );
  MUX \Reg_Bank/U4109  ( .IN0(\Reg_Bank/registers[2][1] ), .IN1(
        \Reg_Bank/registers[3][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4075 )
         );
  MUX \Reg_Bank/U4108  ( .IN0(\Reg_Bank/n4073 ), .IN1(\Reg_Bank/n4072 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4074 ) );
  MUX \Reg_Bank/U4107  ( .IN0(\Reg_Bank/registers[4][1] ), .IN1(
        \Reg_Bank/registers[5][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4073 )
         );
  MUX \Reg_Bank/U4106  ( .IN0(\Reg_Bank/registers[6][1] ), .IN1(
        \Reg_Bank/registers[7][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4072 )
         );
  MUX \Reg_Bank/U4105  ( .IN0(\Reg_Bank/n4070 ), .IN1(\Reg_Bank/n4067 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4071 ) );
  MUX \Reg_Bank/U4104  ( .IN0(\Reg_Bank/n4069 ), .IN1(\Reg_Bank/n4068 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4070 ) );
  MUX \Reg_Bank/U4103  ( .IN0(\Reg_Bank/registers[8][1] ), .IN1(
        \Reg_Bank/registers[9][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4069 )
         );
  MUX \Reg_Bank/U4102  ( .IN0(\Reg_Bank/registers[10][1] ), .IN1(
        \Reg_Bank/registers[11][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4068 )
         );
  MUX \Reg_Bank/U4101  ( .IN0(\Reg_Bank/n4066 ), .IN1(\Reg_Bank/n4065 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4067 ) );
  MUX \Reg_Bank/U4100  ( .IN0(\Reg_Bank/registers[12][1] ), .IN1(
        \Reg_Bank/registers[13][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4066 )
         );
  MUX \Reg_Bank/U4099  ( .IN0(\Reg_Bank/registers[14][1] ), .IN1(
        \Reg_Bank/registers[15][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4065 )
         );
  MUX \Reg_Bank/U4098  ( .IN0(\Reg_Bank/n4063 ), .IN1(\Reg_Bank/n4056 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4064 ) );
  MUX \Reg_Bank/U4097  ( .IN0(\Reg_Bank/n4062 ), .IN1(\Reg_Bank/n4059 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4063 ) );
  MUX \Reg_Bank/U4096  ( .IN0(\Reg_Bank/n4061 ), .IN1(\Reg_Bank/n4060 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4062 ) );
  MUX \Reg_Bank/U4095  ( .IN0(\Reg_Bank/registers[16][1] ), .IN1(
        \Reg_Bank/registers[17][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4061 )
         );
  MUX \Reg_Bank/U4094  ( .IN0(\Reg_Bank/registers[18][1] ), .IN1(
        \Reg_Bank/registers[19][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4060 )
         );
  MUX \Reg_Bank/U4093  ( .IN0(\Reg_Bank/n4058 ), .IN1(\Reg_Bank/n4057 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4059 ) );
  MUX \Reg_Bank/U4092  ( .IN0(\Reg_Bank/registers[20][1] ), .IN1(
        \Reg_Bank/registers[21][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4058 )
         );
  MUX \Reg_Bank/U4091  ( .IN0(\Reg_Bank/registers[22][1] ), .IN1(
        \Reg_Bank/registers[23][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4057 )
         );
  MUX \Reg_Bank/U4090  ( .IN0(\Reg_Bank/n4055 ), .IN1(\Reg_Bank/n4052 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4056 ) );
  MUX \Reg_Bank/U4089  ( .IN0(\Reg_Bank/n4054 ), .IN1(\Reg_Bank/n4053 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4055 ) );
  MUX \Reg_Bank/U4088  ( .IN0(\Reg_Bank/registers[24][1] ), .IN1(
        \Reg_Bank/registers[25][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4054 )
         );
  MUX \Reg_Bank/U4087  ( .IN0(\Reg_Bank/registers[26][1] ), .IN1(
        \Reg_Bank/registers[27][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4053 )
         );
  MUX \Reg_Bank/U4086  ( .IN0(\Reg_Bank/n4051 ), .IN1(\Reg_Bank/n4050 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4052 ) );
  MUX \Reg_Bank/U4085  ( .IN0(\Reg_Bank/registers[28][1] ), .IN1(
        \Reg_Bank/registers[29][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4051 )
         );
  MUX \Reg_Bank/U4084  ( .IN0(\Reg_Bank/registers[30][1] ), .IN1(
        \Reg_Bank/registers[31][1] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4050 )
         );
  MUX \Reg_Bank/U4083  ( .IN0(\Reg_Bank/n4049 ), .IN1(\Reg_Bank/n4034 ), .SEL(
        rs_index[4]), .F(reg_source[0]) );
  MUX \Reg_Bank/U4082  ( .IN0(\Reg_Bank/n4048 ), .IN1(\Reg_Bank/n4041 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4049 ) );
  MUX \Reg_Bank/U4081  ( .IN0(\Reg_Bank/n4047 ), .IN1(\Reg_Bank/n4044 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4048 ) );
  MUX \Reg_Bank/U4080  ( .IN0(\Reg_Bank/n4046 ), .IN1(\Reg_Bank/n4045 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4047 ) );
  MUX \Reg_Bank/U4078  ( .IN0(\Reg_Bank/registers[2][0] ), .IN1(
        \Reg_Bank/registers[3][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4045 )
         );
  MUX \Reg_Bank/U4077  ( .IN0(\Reg_Bank/n4043 ), .IN1(\Reg_Bank/n4042 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4044 ) );
  MUX \Reg_Bank/U4076  ( .IN0(\Reg_Bank/registers[4][0] ), .IN1(
        \Reg_Bank/registers[5][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4043 )
         );
  MUX \Reg_Bank/U4075  ( .IN0(\Reg_Bank/registers[6][0] ), .IN1(
        \Reg_Bank/registers[7][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4042 )
         );
  MUX \Reg_Bank/U4074  ( .IN0(\Reg_Bank/n4040 ), .IN1(\Reg_Bank/n4037 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4041 ) );
  MUX \Reg_Bank/U4073  ( .IN0(\Reg_Bank/n4039 ), .IN1(\Reg_Bank/n4038 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4040 ) );
  MUX \Reg_Bank/U4072  ( .IN0(\Reg_Bank/registers[8][0] ), .IN1(
        \Reg_Bank/registers[9][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4039 )
         );
  MUX \Reg_Bank/U4071  ( .IN0(\Reg_Bank/registers[10][0] ), .IN1(
        \Reg_Bank/registers[11][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4038 )
         );
  MUX \Reg_Bank/U4070  ( .IN0(\Reg_Bank/n4036 ), .IN1(\Reg_Bank/n4035 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4037 ) );
  MUX \Reg_Bank/U4069  ( .IN0(\Reg_Bank/registers[12][0] ), .IN1(
        \Reg_Bank/registers[13][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4036 )
         );
  MUX \Reg_Bank/U4068  ( .IN0(\Reg_Bank/registers[14][0] ), .IN1(
        \Reg_Bank/registers[15][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4035 )
         );
  MUX \Reg_Bank/U4067  ( .IN0(\Reg_Bank/n4033 ), .IN1(\Reg_Bank/n4026 ), .SEL(
        rs_index[3]), .F(\Reg_Bank/n4034 ) );
  MUX \Reg_Bank/U4066  ( .IN0(\Reg_Bank/n4032 ), .IN1(\Reg_Bank/n4029 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4033 ) );
  MUX \Reg_Bank/U4065  ( .IN0(\Reg_Bank/n4031 ), .IN1(\Reg_Bank/n4030 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4032 ) );
  MUX \Reg_Bank/U4064  ( .IN0(\Reg_Bank/registers[16][0] ), .IN1(
        \Reg_Bank/registers[17][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4031 )
         );
  MUX \Reg_Bank/U4063  ( .IN0(\Reg_Bank/registers[18][0] ), .IN1(
        \Reg_Bank/registers[19][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4030 )
         );
  MUX \Reg_Bank/U4062  ( .IN0(\Reg_Bank/n4028 ), .IN1(\Reg_Bank/n4027 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4029 ) );
  MUX \Reg_Bank/U4061  ( .IN0(\Reg_Bank/registers[20][0] ), .IN1(
        \Reg_Bank/registers[21][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4028 )
         );
  MUX \Reg_Bank/U4060  ( .IN0(\Reg_Bank/registers[22][0] ), .IN1(
        \Reg_Bank/registers[23][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4027 )
         );
  MUX \Reg_Bank/U4059  ( .IN0(\Reg_Bank/n4025 ), .IN1(\Reg_Bank/n4022 ), .SEL(
        rs_index[2]), .F(\Reg_Bank/n4026 ) );
  MUX \Reg_Bank/U4058  ( .IN0(\Reg_Bank/n4024 ), .IN1(\Reg_Bank/n4023 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4025 ) );
  MUX \Reg_Bank/U4057  ( .IN0(\Reg_Bank/registers[24][0] ), .IN1(
        \Reg_Bank/registers[25][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4024 )
         );
  MUX \Reg_Bank/U4056  ( .IN0(\Reg_Bank/registers[26][0] ), .IN1(
        \Reg_Bank/registers[27][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4023 )
         );
  MUX \Reg_Bank/U4055  ( .IN0(\Reg_Bank/n4021 ), .IN1(\Reg_Bank/n4020 ), .SEL(
        rs_index[1]), .F(\Reg_Bank/n4022 ) );
  MUX \Reg_Bank/U4054  ( .IN0(\Reg_Bank/registers[28][0] ), .IN1(
        \Reg_Bank/registers[29][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4021 )
         );
  MUX \Reg_Bank/U4053  ( .IN0(\Reg_Bank/registers[30][0] ), .IN1(
        \Reg_Bank/registers[31][0] ), .SEL(rs_index[0]), .F(\Reg_Bank/n4020 )
         );
  DFF \Reg_Bank/registers_reg[1][0]  ( .D(\Reg_Bank/n3028 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][0] ) );
  DFF \Reg_Bank/registers_reg[1][1]  ( .D(\Reg_Bank/n3029 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][1] ) );
  DFF \Reg_Bank/registers_reg[1][2]  ( .D(\Reg_Bank/n3030 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][2] ) );
  DFF \Reg_Bank/registers_reg[1][3]  ( .D(\Reg_Bank/n3031 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][3] ) );
  DFF \Reg_Bank/registers_reg[1][4]  ( .D(\Reg_Bank/n3032 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][4] ) );
  DFF \Reg_Bank/registers_reg[1][5]  ( .D(\Reg_Bank/n3033 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][5] ) );
  DFF \Reg_Bank/registers_reg[1][6]  ( .D(\Reg_Bank/n3034 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][6] ) );
  DFF \Reg_Bank/registers_reg[1][7]  ( .D(\Reg_Bank/n3035 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][7] ) );
  DFF \Reg_Bank/registers_reg[1][8]  ( .D(\Reg_Bank/n3036 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][8] ) );
  DFF \Reg_Bank/registers_reg[1][9]  ( .D(\Reg_Bank/n3037 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][9] ) );
  DFF \Reg_Bank/registers_reg[1][10]  ( .D(\Reg_Bank/n3038 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][10] ) );
  DFF \Reg_Bank/registers_reg[1][11]  ( .D(\Reg_Bank/n3039 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][11] ) );
  DFF \Reg_Bank/registers_reg[1][12]  ( .D(\Reg_Bank/n3040 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][12] ) );
  DFF \Reg_Bank/registers_reg[1][13]  ( .D(\Reg_Bank/n3041 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][13] ) );
  DFF \Reg_Bank/registers_reg[1][14]  ( .D(\Reg_Bank/n3042 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][14] ) );
  DFF \Reg_Bank/registers_reg[1][15]  ( .D(\Reg_Bank/n3043 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][15] ) );
  DFF \Reg_Bank/registers_reg[1][16]  ( .D(\Reg_Bank/n3044 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][16] ) );
  DFF \Reg_Bank/registers_reg[1][17]  ( .D(\Reg_Bank/n3045 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][17] ) );
  DFF \Reg_Bank/registers_reg[1][18]  ( .D(\Reg_Bank/n3046 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][18] ) );
  DFF \Reg_Bank/registers_reg[1][19]  ( .D(\Reg_Bank/n3047 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][19] ) );
  DFF \Reg_Bank/registers_reg[1][20]  ( .D(\Reg_Bank/n3048 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][20] ) );
  DFF \Reg_Bank/registers_reg[1][21]  ( .D(\Reg_Bank/n3049 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][21] ) );
  DFF \Reg_Bank/registers_reg[1][22]  ( .D(\Reg_Bank/n3050 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][22] ) );
  DFF \Reg_Bank/registers_reg[1][23]  ( .D(\Reg_Bank/n3051 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][23] ) );
  DFF \Reg_Bank/registers_reg[1][24]  ( .D(\Reg_Bank/n3052 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][24] ) );
  DFF \Reg_Bank/registers_reg[1][25]  ( .D(\Reg_Bank/n3053 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][25] ) );
  DFF \Reg_Bank/registers_reg[1][26]  ( .D(\Reg_Bank/n3054 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][26] ) );
  DFF \Reg_Bank/registers_reg[1][27]  ( .D(\Reg_Bank/n3055 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][27] ) );
  DFF \Reg_Bank/registers_reg[1][28]  ( .D(\Reg_Bank/n3056 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][28] ) );
  DFF \Reg_Bank/registers_reg[1][29]  ( .D(\Reg_Bank/n3057 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][29] ) );
  DFF \Reg_Bank/registers_reg[1][30]  ( .D(\Reg_Bank/n3058 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][30] ) );
  DFF \Reg_Bank/registers_reg[1][31]  ( .D(\Reg_Bank/n3059 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[1][31] ) );
  DFF \Reg_Bank/registers_reg[2][0]  ( .D(\Reg_Bank/n3060 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][0] ) );
  DFF \Reg_Bank/registers_reg[2][1]  ( .D(\Reg_Bank/n3061 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][1] ) );
  DFF \Reg_Bank/registers_reg[2][2]  ( .D(\Reg_Bank/n3062 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][2] ) );
  DFF \Reg_Bank/registers_reg[2][3]  ( .D(\Reg_Bank/n3063 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][3] ) );
  DFF \Reg_Bank/registers_reg[2][4]  ( .D(\Reg_Bank/n3064 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][4] ) );
  DFF \Reg_Bank/registers_reg[2][5]  ( .D(\Reg_Bank/n3065 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][5] ) );
  DFF \Reg_Bank/registers_reg[2][6]  ( .D(\Reg_Bank/n3066 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][6] ) );
  DFF \Reg_Bank/registers_reg[2][7]  ( .D(\Reg_Bank/n3067 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][7] ) );
  DFF \Reg_Bank/registers_reg[2][8]  ( .D(\Reg_Bank/n3068 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][8] ) );
  DFF \Reg_Bank/registers_reg[2][9]  ( .D(\Reg_Bank/n3069 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][9] ) );
  DFF \Reg_Bank/registers_reg[2][10]  ( .D(\Reg_Bank/n3070 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][10] ) );
  DFF \Reg_Bank/registers_reg[2][11]  ( .D(\Reg_Bank/n3071 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][11] ) );
  DFF \Reg_Bank/registers_reg[2][12]  ( .D(\Reg_Bank/n3072 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][12] ) );
  DFF \Reg_Bank/registers_reg[2][13]  ( .D(\Reg_Bank/n3073 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][13] ) );
  DFF \Reg_Bank/registers_reg[2][14]  ( .D(\Reg_Bank/n3074 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][14] ) );
  DFF \Reg_Bank/registers_reg[2][15]  ( .D(\Reg_Bank/n3075 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][15] ) );
  DFF \Reg_Bank/registers_reg[2][16]  ( .D(\Reg_Bank/n3076 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][16] ) );
  DFF \Reg_Bank/registers_reg[2][17]  ( .D(\Reg_Bank/n3077 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][17] ) );
  DFF \Reg_Bank/registers_reg[2][18]  ( .D(\Reg_Bank/n3078 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][18] ) );
  DFF \Reg_Bank/registers_reg[2][19]  ( .D(\Reg_Bank/n3079 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][19] ) );
  DFF \Reg_Bank/registers_reg[2][20]  ( .D(\Reg_Bank/n3080 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][20] ) );
  DFF \Reg_Bank/registers_reg[2][21]  ( .D(\Reg_Bank/n3081 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][21] ) );
  DFF \Reg_Bank/registers_reg[2][22]  ( .D(\Reg_Bank/n3082 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][22] ) );
  DFF \Reg_Bank/registers_reg[2][23]  ( .D(\Reg_Bank/n3083 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][23] ) );
  DFF \Reg_Bank/registers_reg[2][24]  ( .D(\Reg_Bank/n3084 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][24] ) );
  DFF \Reg_Bank/registers_reg[2][25]  ( .D(\Reg_Bank/n3085 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][25] ) );
  DFF \Reg_Bank/registers_reg[2][26]  ( .D(\Reg_Bank/n3086 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][26] ) );
  DFF \Reg_Bank/registers_reg[2][27]  ( .D(\Reg_Bank/n3087 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][27] ) );
  DFF \Reg_Bank/registers_reg[2][28]  ( .D(\Reg_Bank/n3088 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][28] ) );
  DFF \Reg_Bank/registers_reg[2][29]  ( .D(\Reg_Bank/n3089 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][29] ) );
  DFF \Reg_Bank/registers_reg[2][30]  ( .D(\Reg_Bank/n3090 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][30] ) );
  DFF \Reg_Bank/registers_reg[2][31]  ( .D(\Reg_Bank/n3091 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[2][31] ) );
  DFF \Reg_Bank/registers_reg[3][0]  ( .D(\Reg_Bank/n3092 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][0] ) );
  DFF \Reg_Bank/registers_reg[3][1]  ( .D(\Reg_Bank/n3093 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][1] ) );
  DFF \Reg_Bank/registers_reg[3][2]  ( .D(\Reg_Bank/n3094 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][2] ) );
  DFF \Reg_Bank/registers_reg[3][3]  ( .D(\Reg_Bank/n3095 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][3] ) );
  DFF \Reg_Bank/registers_reg[3][4]  ( .D(\Reg_Bank/n3096 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][4] ) );
  DFF \Reg_Bank/registers_reg[3][5]  ( .D(\Reg_Bank/n3097 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][5] ) );
  DFF \Reg_Bank/registers_reg[3][6]  ( .D(\Reg_Bank/n3098 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][6] ) );
  DFF \Reg_Bank/registers_reg[3][7]  ( .D(\Reg_Bank/n3099 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][7] ) );
  DFF \Reg_Bank/registers_reg[3][8]  ( .D(\Reg_Bank/n3100 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][8] ) );
  DFF \Reg_Bank/registers_reg[3][9]  ( .D(\Reg_Bank/n3101 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][9] ) );
  DFF \Reg_Bank/registers_reg[3][10]  ( .D(\Reg_Bank/n3102 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][10] ) );
  DFF \Reg_Bank/registers_reg[3][11]  ( .D(\Reg_Bank/n3103 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][11] ) );
  DFF \Reg_Bank/registers_reg[3][12]  ( .D(\Reg_Bank/n3104 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][12] ) );
  DFF \Reg_Bank/registers_reg[3][13]  ( .D(\Reg_Bank/n3105 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][13] ) );
  DFF \Reg_Bank/registers_reg[3][14]  ( .D(\Reg_Bank/n3106 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][14] ) );
  DFF \Reg_Bank/registers_reg[3][15]  ( .D(\Reg_Bank/n3107 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][15] ) );
  DFF \Reg_Bank/registers_reg[3][16]  ( .D(\Reg_Bank/n3108 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][16] ) );
  DFF \Reg_Bank/registers_reg[3][17]  ( .D(\Reg_Bank/n3109 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][17] ) );
  DFF \Reg_Bank/registers_reg[3][18]  ( .D(\Reg_Bank/n3110 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][18] ) );
  DFF \Reg_Bank/registers_reg[3][19]  ( .D(\Reg_Bank/n3111 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][19] ) );
  DFF \Reg_Bank/registers_reg[3][20]  ( .D(\Reg_Bank/n3112 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][20] ) );
  DFF \Reg_Bank/registers_reg[3][21]  ( .D(\Reg_Bank/n3113 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][21] ) );
  DFF \Reg_Bank/registers_reg[3][22]  ( .D(\Reg_Bank/n3114 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][22] ) );
  DFF \Reg_Bank/registers_reg[3][23]  ( .D(\Reg_Bank/n3115 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][23] ) );
  DFF \Reg_Bank/registers_reg[3][24]  ( .D(\Reg_Bank/n3116 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][24] ) );
  DFF \Reg_Bank/registers_reg[3][25]  ( .D(\Reg_Bank/n3117 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][25] ) );
  DFF \Reg_Bank/registers_reg[3][26]  ( .D(\Reg_Bank/n3118 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][26] ) );
  DFF \Reg_Bank/registers_reg[3][27]  ( .D(\Reg_Bank/n3119 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][27] ) );
  DFF \Reg_Bank/registers_reg[3][28]  ( .D(\Reg_Bank/n3120 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][28] ) );
  DFF \Reg_Bank/registers_reg[3][29]  ( .D(\Reg_Bank/n3121 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][29] ) );
  DFF \Reg_Bank/registers_reg[3][30]  ( .D(\Reg_Bank/n3122 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][30] ) );
  DFF \Reg_Bank/registers_reg[3][31]  ( .D(\Reg_Bank/n3123 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[3][31] ) );
  DFF \Reg_Bank/registers_reg[4][0]  ( .D(\Reg_Bank/n3124 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][0] ) );
  DFF \Reg_Bank/registers_reg[4][1]  ( .D(\Reg_Bank/n3125 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][1] ) );
  DFF \Reg_Bank/registers_reg[4][2]  ( .D(\Reg_Bank/n3126 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][2] ) );
  DFF \Reg_Bank/registers_reg[4][3]  ( .D(\Reg_Bank/n3127 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][3] ) );
  DFF \Reg_Bank/registers_reg[4][4]  ( .D(\Reg_Bank/n3128 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][4] ) );
  DFF \Reg_Bank/registers_reg[4][5]  ( .D(\Reg_Bank/n3129 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][5] ) );
  DFF \Reg_Bank/registers_reg[4][6]  ( .D(\Reg_Bank/n3130 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][6] ) );
  DFF \Reg_Bank/registers_reg[4][7]  ( .D(\Reg_Bank/n3131 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][7] ) );
  DFF \Reg_Bank/registers_reg[4][8]  ( .D(\Reg_Bank/n3132 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][8] ) );
  DFF \Reg_Bank/registers_reg[4][9]  ( .D(\Reg_Bank/n3133 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][9] ) );
  DFF \Reg_Bank/registers_reg[4][10]  ( .D(\Reg_Bank/n3134 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][10] ) );
  DFF \Reg_Bank/registers_reg[4][11]  ( .D(\Reg_Bank/n3135 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][11] ) );
  DFF \Reg_Bank/registers_reg[4][12]  ( .D(\Reg_Bank/n3136 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][12] ) );
  DFF \Reg_Bank/registers_reg[4][13]  ( .D(\Reg_Bank/n3137 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][13] ) );
  DFF \Reg_Bank/registers_reg[4][14]  ( .D(\Reg_Bank/n3138 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][14] ) );
  DFF \Reg_Bank/registers_reg[4][15]  ( .D(\Reg_Bank/n3139 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][15] ) );
  DFF \Reg_Bank/registers_reg[4][16]  ( .D(\Reg_Bank/n3140 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][16] ) );
  DFF \Reg_Bank/registers_reg[4][17]  ( .D(\Reg_Bank/n3141 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][17] ) );
  DFF \Reg_Bank/registers_reg[4][18]  ( .D(\Reg_Bank/n3142 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][18] ) );
  DFF \Reg_Bank/registers_reg[4][19]  ( .D(\Reg_Bank/n3143 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][19] ) );
  DFF \Reg_Bank/registers_reg[4][20]  ( .D(\Reg_Bank/n3144 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][20] ) );
  DFF \Reg_Bank/registers_reg[4][21]  ( .D(\Reg_Bank/n3145 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][21] ) );
  DFF \Reg_Bank/registers_reg[4][22]  ( .D(\Reg_Bank/n3146 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][22] ) );
  DFF \Reg_Bank/registers_reg[4][23]  ( .D(\Reg_Bank/n3147 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][23] ) );
  DFF \Reg_Bank/registers_reg[4][24]  ( .D(\Reg_Bank/n3148 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][24] ) );
  DFF \Reg_Bank/registers_reg[4][25]  ( .D(\Reg_Bank/n3149 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][25] ) );
  DFF \Reg_Bank/registers_reg[4][26]  ( .D(\Reg_Bank/n3150 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][26] ) );
  DFF \Reg_Bank/registers_reg[4][27]  ( .D(\Reg_Bank/n3151 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][27] ) );
  DFF \Reg_Bank/registers_reg[4][28]  ( .D(\Reg_Bank/n3152 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][28] ) );
  DFF \Reg_Bank/registers_reg[4][29]  ( .D(\Reg_Bank/n3153 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][29] ) );
  DFF \Reg_Bank/registers_reg[4][30]  ( .D(\Reg_Bank/n3154 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][30] ) );
  DFF \Reg_Bank/registers_reg[4][31]  ( .D(\Reg_Bank/n3155 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[4][31] ) );
  DFF \Reg_Bank/registers_reg[5][0]  ( .D(\Reg_Bank/n3156 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][0] ) );
  DFF \Reg_Bank/registers_reg[5][1]  ( .D(\Reg_Bank/n3157 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][1] ) );
  DFF \Reg_Bank/registers_reg[5][2]  ( .D(\Reg_Bank/n3158 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][2] ) );
  DFF \Reg_Bank/registers_reg[5][3]  ( .D(\Reg_Bank/n3159 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][3] ) );
  DFF \Reg_Bank/registers_reg[5][4]  ( .D(\Reg_Bank/n3160 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][4] ) );
  DFF \Reg_Bank/registers_reg[5][5]  ( .D(\Reg_Bank/n3161 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][5] ) );
  DFF \Reg_Bank/registers_reg[5][6]  ( .D(\Reg_Bank/n3162 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][6] ) );
  DFF \Reg_Bank/registers_reg[5][7]  ( .D(\Reg_Bank/n3163 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][7] ) );
  DFF \Reg_Bank/registers_reg[5][8]  ( .D(\Reg_Bank/n3164 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][8] ) );
  DFF \Reg_Bank/registers_reg[5][9]  ( .D(\Reg_Bank/n3165 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][9] ) );
  DFF \Reg_Bank/registers_reg[5][10]  ( .D(\Reg_Bank/n3166 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][10] ) );
  DFF \Reg_Bank/registers_reg[5][11]  ( .D(\Reg_Bank/n3167 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][11] ) );
  DFF \Reg_Bank/registers_reg[5][12]  ( .D(\Reg_Bank/n3168 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][12] ) );
  DFF \Reg_Bank/registers_reg[5][13]  ( .D(\Reg_Bank/n3169 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][13] ) );
  DFF \Reg_Bank/registers_reg[5][14]  ( .D(\Reg_Bank/n3170 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][14] ) );
  DFF \Reg_Bank/registers_reg[5][15]  ( .D(\Reg_Bank/n3171 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][15] ) );
  DFF \Reg_Bank/registers_reg[5][16]  ( .D(\Reg_Bank/n3172 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][16] ) );
  DFF \Reg_Bank/registers_reg[5][17]  ( .D(\Reg_Bank/n3173 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][17] ) );
  DFF \Reg_Bank/registers_reg[5][18]  ( .D(\Reg_Bank/n3174 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][18] ) );
  DFF \Reg_Bank/registers_reg[5][19]  ( .D(\Reg_Bank/n3175 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][19] ) );
  DFF \Reg_Bank/registers_reg[5][20]  ( .D(\Reg_Bank/n3176 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][20] ) );
  DFF \Reg_Bank/registers_reg[5][21]  ( .D(\Reg_Bank/n3177 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][21] ) );
  DFF \Reg_Bank/registers_reg[5][22]  ( .D(\Reg_Bank/n3178 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][22] ) );
  DFF \Reg_Bank/registers_reg[5][23]  ( .D(\Reg_Bank/n3179 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][23] ) );
  DFF \Reg_Bank/registers_reg[5][24]  ( .D(\Reg_Bank/n3180 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][24] ) );
  DFF \Reg_Bank/registers_reg[5][25]  ( .D(\Reg_Bank/n3181 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][25] ) );
  DFF \Reg_Bank/registers_reg[5][26]  ( .D(\Reg_Bank/n3182 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][26] ) );
  DFF \Reg_Bank/registers_reg[5][27]  ( .D(\Reg_Bank/n3183 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][27] ) );
  DFF \Reg_Bank/registers_reg[5][28]  ( .D(\Reg_Bank/n3184 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][28] ) );
  DFF \Reg_Bank/registers_reg[5][29]  ( .D(\Reg_Bank/n3185 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][29] ) );
  DFF \Reg_Bank/registers_reg[5][30]  ( .D(\Reg_Bank/n3186 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][30] ) );
  DFF \Reg_Bank/registers_reg[5][31]  ( .D(\Reg_Bank/n3187 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[5][31] ) );
  DFF \Reg_Bank/registers_reg[6][0]  ( .D(\Reg_Bank/n3188 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][0] ) );
  DFF \Reg_Bank/registers_reg[6][1]  ( .D(\Reg_Bank/n3189 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][1] ) );
  DFF \Reg_Bank/registers_reg[6][2]  ( .D(\Reg_Bank/n3190 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][2] ) );
  DFF \Reg_Bank/registers_reg[6][3]  ( .D(\Reg_Bank/n3191 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][3] ) );
  DFF \Reg_Bank/registers_reg[6][4]  ( .D(\Reg_Bank/n3192 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][4] ) );
  DFF \Reg_Bank/registers_reg[6][5]  ( .D(\Reg_Bank/n3193 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][5] ) );
  DFF \Reg_Bank/registers_reg[6][6]  ( .D(\Reg_Bank/n3194 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][6] ) );
  DFF \Reg_Bank/registers_reg[6][7]  ( .D(\Reg_Bank/n3195 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][7] ) );
  DFF \Reg_Bank/registers_reg[6][8]  ( .D(\Reg_Bank/n3196 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][8] ) );
  DFF \Reg_Bank/registers_reg[6][9]  ( .D(\Reg_Bank/n3197 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][9] ) );
  DFF \Reg_Bank/registers_reg[6][10]  ( .D(\Reg_Bank/n3198 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][10] ) );
  DFF \Reg_Bank/registers_reg[6][11]  ( .D(\Reg_Bank/n3199 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][11] ) );
  DFF \Reg_Bank/registers_reg[6][12]  ( .D(\Reg_Bank/n3200 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][12] ) );
  DFF \Reg_Bank/registers_reg[6][13]  ( .D(\Reg_Bank/n3201 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][13] ) );
  DFF \Reg_Bank/registers_reg[6][14]  ( .D(\Reg_Bank/n3202 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][14] ) );
  DFF \Reg_Bank/registers_reg[6][15]  ( .D(\Reg_Bank/n3203 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][15] ) );
  DFF \Reg_Bank/registers_reg[6][16]  ( .D(\Reg_Bank/n3204 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][16] ) );
  DFF \Reg_Bank/registers_reg[6][17]  ( .D(\Reg_Bank/n3205 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][17] ) );
  DFF \Reg_Bank/registers_reg[6][18]  ( .D(\Reg_Bank/n3206 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][18] ) );
  DFF \Reg_Bank/registers_reg[6][19]  ( .D(\Reg_Bank/n3207 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][19] ) );
  DFF \Reg_Bank/registers_reg[6][20]  ( .D(\Reg_Bank/n3208 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][20] ) );
  DFF \Reg_Bank/registers_reg[6][21]  ( .D(\Reg_Bank/n3209 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][21] ) );
  DFF \Reg_Bank/registers_reg[6][22]  ( .D(\Reg_Bank/n3210 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][22] ) );
  DFF \Reg_Bank/registers_reg[6][23]  ( .D(\Reg_Bank/n3211 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][23] ) );
  DFF \Reg_Bank/registers_reg[6][24]  ( .D(\Reg_Bank/n3212 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][24] ) );
  DFF \Reg_Bank/registers_reg[6][25]  ( .D(\Reg_Bank/n3213 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][25] ) );
  DFF \Reg_Bank/registers_reg[6][26]  ( .D(\Reg_Bank/n3214 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][26] ) );
  DFF \Reg_Bank/registers_reg[6][27]  ( .D(\Reg_Bank/n3215 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][27] ) );
  DFF \Reg_Bank/registers_reg[6][28]  ( .D(\Reg_Bank/n3216 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][28] ) );
  DFF \Reg_Bank/registers_reg[6][29]  ( .D(\Reg_Bank/n3217 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][29] ) );
  DFF \Reg_Bank/registers_reg[6][30]  ( .D(\Reg_Bank/n3218 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][30] ) );
  DFF \Reg_Bank/registers_reg[6][31]  ( .D(\Reg_Bank/n3219 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[6][31] ) );
  DFF \Reg_Bank/registers_reg[7][0]  ( .D(\Reg_Bank/n3220 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][0] ) );
  DFF \Reg_Bank/registers_reg[7][1]  ( .D(\Reg_Bank/n3221 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][1] ) );
  DFF \Reg_Bank/registers_reg[7][2]  ( .D(\Reg_Bank/n3222 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][2] ) );
  DFF \Reg_Bank/registers_reg[7][3]  ( .D(\Reg_Bank/n3223 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][3] ) );
  DFF \Reg_Bank/registers_reg[7][4]  ( .D(\Reg_Bank/n3224 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][4] ) );
  DFF \Reg_Bank/registers_reg[7][5]  ( .D(\Reg_Bank/n3225 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][5] ) );
  DFF \Reg_Bank/registers_reg[7][6]  ( .D(\Reg_Bank/n3226 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][6] ) );
  DFF \Reg_Bank/registers_reg[7][7]  ( .D(\Reg_Bank/n3227 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][7] ) );
  DFF \Reg_Bank/registers_reg[7][8]  ( .D(\Reg_Bank/n3228 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][8] ) );
  DFF \Reg_Bank/registers_reg[7][9]  ( .D(\Reg_Bank/n3229 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][9] ) );
  DFF \Reg_Bank/registers_reg[7][10]  ( .D(\Reg_Bank/n3230 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][10] ) );
  DFF \Reg_Bank/registers_reg[7][11]  ( .D(\Reg_Bank/n3231 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][11] ) );
  DFF \Reg_Bank/registers_reg[7][12]  ( .D(\Reg_Bank/n3232 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][12] ) );
  DFF \Reg_Bank/registers_reg[7][13]  ( .D(\Reg_Bank/n3233 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][13] ) );
  DFF \Reg_Bank/registers_reg[7][14]  ( .D(\Reg_Bank/n3234 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][14] ) );
  DFF \Reg_Bank/registers_reg[7][15]  ( .D(\Reg_Bank/n3235 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][15] ) );
  DFF \Reg_Bank/registers_reg[7][16]  ( .D(\Reg_Bank/n3236 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][16] ) );
  DFF \Reg_Bank/registers_reg[7][17]  ( .D(\Reg_Bank/n3237 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][17] ) );
  DFF \Reg_Bank/registers_reg[7][18]  ( .D(\Reg_Bank/n3238 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][18] ) );
  DFF \Reg_Bank/registers_reg[7][19]  ( .D(\Reg_Bank/n3239 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][19] ) );
  DFF \Reg_Bank/registers_reg[7][20]  ( .D(\Reg_Bank/n3240 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][20] ) );
  DFF \Reg_Bank/registers_reg[7][21]  ( .D(\Reg_Bank/n3241 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][21] ) );
  DFF \Reg_Bank/registers_reg[7][22]  ( .D(\Reg_Bank/n3242 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][22] ) );
  DFF \Reg_Bank/registers_reg[7][23]  ( .D(\Reg_Bank/n3243 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][23] ) );
  DFF \Reg_Bank/registers_reg[7][24]  ( .D(\Reg_Bank/n3244 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][24] ) );
  DFF \Reg_Bank/registers_reg[7][25]  ( .D(\Reg_Bank/n3245 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][25] ) );
  DFF \Reg_Bank/registers_reg[7][26]  ( .D(\Reg_Bank/n3246 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][26] ) );
  DFF \Reg_Bank/registers_reg[7][27]  ( .D(\Reg_Bank/n3247 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][27] ) );
  DFF \Reg_Bank/registers_reg[7][28]  ( .D(\Reg_Bank/n3248 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][28] ) );
  DFF \Reg_Bank/registers_reg[7][29]  ( .D(\Reg_Bank/n3249 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][29] ) );
  DFF \Reg_Bank/registers_reg[7][30]  ( .D(\Reg_Bank/n3250 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][30] ) );
  DFF \Reg_Bank/registers_reg[7][31]  ( .D(\Reg_Bank/n3251 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[7][31] ) );
  DFF \Reg_Bank/registers_reg[8][0]  ( .D(\Reg_Bank/n3252 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][0] ) );
  DFF \Reg_Bank/registers_reg[8][1]  ( .D(\Reg_Bank/n3253 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][1] ) );
  DFF \Reg_Bank/registers_reg[8][2]  ( .D(\Reg_Bank/n3254 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][2] ) );
  DFF \Reg_Bank/registers_reg[8][3]  ( .D(\Reg_Bank/n3255 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][3] ) );
  DFF \Reg_Bank/registers_reg[8][4]  ( .D(\Reg_Bank/n3256 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][4] ) );
  DFF \Reg_Bank/registers_reg[8][5]  ( .D(\Reg_Bank/n3257 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][5] ) );
  DFF \Reg_Bank/registers_reg[8][6]  ( .D(\Reg_Bank/n3258 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][6] ) );
  DFF \Reg_Bank/registers_reg[8][7]  ( .D(\Reg_Bank/n3259 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][7] ) );
  DFF \Reg_Bank/registers_reg[8][8]  ( .D(\Reg_Bank/n3260 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][8] ) );
  DFF \Reg_Bank/registers_reg[8][9]  ( .D(\Reg_Bank/n3261 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][9] ) );
  DFF \Reg_Bank/registers_reg[8][10]  ( .D(\Reg_Bank/n3262 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][10] ) );
  DFF \Reg_Bank/registers_reg[8][11]  ( .D(\Reg_Bank/n3263 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][11] ) );
  DFF \Reg_Bank/registers_reg[8][12]  ( .D(\Reg_Bank/n3264 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][12] ) );
  DFF \Reg_Bank/registers_reg[8][13]  ( .D(\Reg_Bank/n3265 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][13] ) );
  DFF \Reg_Bank/registers_reg[8][14]  ( .D(\Reg_Bank/n3266 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][14] ) );
  DFF \Reg_Bank/registers_reg[8][15]  ( .D(\Reg_Bank/n3267 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][15] ) );
  DFF \Reg_Bank/registers_reg[8][16]  ( .D(\Reg_Bank/n3268 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][16] ) );
  DFF \Reg_Bank/registers_reg[8][17]  ( .D(\Reg_Bank/n3269 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][17] ) );
  DFF \Reg_Bank/registers_reg[8][18]  ( .D(\Reg_Bank/n3270 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][18] ) );
  DFF \Reg_Bank/registers_reg[8][19]  ( .D(\Reg_Bank/n3271 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][19] ) );
  DFF \Reg_Bank/registers_reg[8][20]  ( .D(\Reg_Bank/n3272 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][20] ) );
  DFF \Reg_Bank/registers_reg[8][21]  ( .D(\Reg_Bank/n3273 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][21] ) );
  DFF \Reg_Bank/registers_reg[8][22]  ( .D(\Reg_Bank/n3274 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][22] ) );
  DFF \Reg_Bank/registers_reg[8][23]  ( .D(\Reg_Bank/n3275 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][23] ) );
  DFF \Reg_Bank/registers_reg[8][24]  ( .D(\Reg_Bank/n3276 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][24] ) );
  DFF \Reg_Bank/registers_reg[8][25]  ( .D(\Reg_Bank/n3277 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][25] ) );
  DFF \Reg_Bank/registers_reg[8][26]  ( .D(\Reg_Bank/n3278 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][26] ) );
  DFF \Reg_Bank/registers_reg[8][27]  ( .D(\Reg_Bank/n3279 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][27] ) );
  DFF \Reg_Bank/registers_reg[8][28]  ( .D(\Reg_Bank/n3280 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][28] ) );
  DFF \Reg_Bank/registers_reg[8][29]  ( .D(\Reg_Bank/n3281 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][29] ) );
  DFF \Reg_Bank/registers_reg[8][30]  ( .D(\Reg_Bank/n3282 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][30] ) );
  DFF \Reg_Bank/registers_reg[8][31]  ( .D(\Reg_Bank/n3283 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[8][31] ) );
  DFF \Reg_Bank/registers_reg[9][0]  ( .D(\Reg_Bank/n3284 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][0] ) );
  DFF \Reg_Bank/registers_reg[9][1]  ( .D(\Reg_Bank/n3285 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][1] ) );
  DFF \Reg_Bank/registers_reg[9][2]  ( .D(\Reg_Bank/n3286 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][2] ) );
  DFF \Reg_Bank/registers_reg[9][3]  ( .D(\Reg_Bank/n3287 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][3] ) );
  DFF \Reg_Bank/registers_reg[9][4]  ( .D(\Reg_Bank/n3288 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][4] ) );
  DFF \Reg_Bank/registers_reg[9][5]  ( .D(\Reg_Bank/n3289 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][5] ) );
  DFF \Reg_Bank/registers_reg[9][6]  ( .D(\Reg_Bank/n3290 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][6] ) );
  DFF \Reg_Bank/registers_reg[9][7]  ( .D(\Reg_Bank/n3291 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][7] ) );
  DFF \Reg_Bank/registers_reg[9][8]  ( .D(\Reg_Bank/n3292 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][8] ) );
  DFF \Reg_Bank/registers_reg[9][9]  ( .D(\Reg_Bank/n3293 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][9] ) );
  DFF \Reg_Bank/registers_reg[9][10]  ( .D(\Reg_Bank/n3294 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][10] ) );
  DFF \Reg_Bank/registers_reg[9][11]  ( .D(\Reg_Bank/n3295 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][11] ) );
  DFF \Reg_Bank/registers_reg[9][12]  ( .D(\Reg_Bank/n3296 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][12] ) );
  DFF \Reg_Bank/registers_reg[9][13]  ( .D(\Reg_Bank/n3297 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][13] ) );
  DFF \Reg_Bank/registers_reg[9][14]  ( .D(\Reg_Bank/n3298 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][14] ) );
  DFF \Reg_Bank/registers_reg[9][15]  ( .D(\Reg_Bank/n3299 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][15] ) );
  DFF \Reg_Bank/registers_reg[9][16]  ( .D(\Reg_Bank/n3300 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][16] ) );
  DFF \Reg_Bank/registers_reg[9][17]  ( .D(\Reg_Bank/n3301 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][17] ) );
  DFF \Reg_Bank/registers_reg[9][18]  ( .D(\Reg_Bank/n3302 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][18] ) );
  DFF \Reg_Bank/registers_reg[9][19]  ( .D(\Reg_Bank/n3303 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][19] ) );
  DFF \Reg_Bank/registers_reg[9][20]  ( .D(\Reg_Bank/n3304 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][20] ) );
  DFF \Reg_Bank/registers_reg[9][21]  ( .D(\Reg_Bank/n3305 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][21] ) );
  DFF \Reg_Bank/registers_reg[9][22]  ( .D(\Reg_Bank/n3306 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][22] ) );
  DFF \Reg_Bank/registers_reg[9][23]  ( .D(\Reg_Bank/n3307 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][23] ) );
  DFF \Reg_Bank/registers_reg[9][24]  ( .D(\Reg_Bank/n3308 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][24] ) );
  DFF \Reg_Bank/registers_reg[9][25]  ( .D(\Reg_Bank/n3309 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][25] ) );
  DFF \Reg_Bank/registers_reg[9][26]  ( .D(\Reg_Bank/n3310 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][26] ) );
  DFF \Reg_Bank/registers_reg[9][27]  ( .D(\Reg_Bank/n3311 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][27] ) );
  DFF \Reg_Bank/registers_reg[9][28]  ( .D(\Reg_Bank/n3312 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][28] ) );
  DFF \Reg_Bank/registers_reg[9][29]  ( .D(\Reg_Bank/n3313 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][29] ) );
  DFF \Reg_Bank/registers_reg[9][30]  ( .D(\Reg_Bank/n3314 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][30] ) );
  DFF \Reg_Bank/registers_reg[9][31]  ( .D(\Reg_Bank/n3315 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[9][31] ) );
  DFF \Reg_Bank/registers_reg[10][0]  ( .D(\Reg_Bank/n3316 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][0] ) );
  DFF \Reg_Bank/registers_reg[10][1]  ( .D(\Reg_Bank/n3317 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][1] ) );
  DFF \Reg_Bank/registers_reg[10][2]  ( .D(\Reg_Bank/n3318 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][2] ) );
  DFF \Reg_Bank/registers_reg[10][3]  ( .D(\Reg_Bank/n3319 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][3] ) );
  DFF \Reg_Bank/registers_reg[10][4]  ( .D(\Reg_Bank/n3320 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][4] ) );
  DFF \Reg_Bank/registers_reg[10][5]  ( .D(\Reg_Bank/n3321 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][5] ) );
  DFF \Reg_Bank/registers_reg[10][6]  ( .D(\Reg_Bank/n3322 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][6] ) );
  DFF \Reg_Bank/registers_reg[10][7]  ( .D(\Reg_Bank/n3323 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][7] ) );
  DFF \Reg_Bank/registers_reg[10][8]  ( .D(\Reg_Bank/n3324 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][8] ) );
  DFF \Reg_Bank/registers_reg[10][9]  ( .D(\Reg_Bank/n3325 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[10][9] ) );
  DFF \Reg_Bank/registers_reg[10][10]  ( .D(\Reg_Bank/n3326 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][10] ) );
  DFF \Reg_Bank/registers_reg[10][11]  ( .D(\Reg_Bank/n3327 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][11] ) );
  DFF \Reg_Bank/registers_reg[10][12]  ( .D(\Reg_Bank/n3328 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][12] ) );
  DFF \Reg_Bank/registers_reg[10][13]  ( .D(\Reg_Bank/n3329 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][13] ) );
  DFF \Reg_Bank/registers_reg[10][14]  ( .D(\Reg_Bank/n3330 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][14] ) );
  DFF \Reg_Bank/registers_reg[10][15]  ( .D(\Reg_Bank/n3331 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][15] ) );
  DFF \Reg_Bank/registers_reg[10][16]  ( .D(\Reg_Bank/n3332 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][16] ) );
  DFF \Reg_Bank/registers_reg[10][17]  ( .D(\Reg_Bank/n3333 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][17] ) );
  DFF \Reg_Bank/registers_reg[10][18]  ( .D(\Reg_Bank/n3334 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][18] ) );
  DFF \Reg_Bank/registers_reg[10][19]  ( .D(\Reg_Bank/n3335 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][19] ) );
  DFF \Reg_Bank/registers_reg[10][20]  ( .D(\Reg_Bank/n3336 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][20] ) );
  DFF \Reg_Bank/registers_reg[10][21]  ( .D(\Reg_Bank/n3337 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][21] ) );
  DFF \Reg_Bank/registers_reg[10][22]  ( .D(\Reg_Bank/n3338 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][22] ) );
  DFF \Reg_Bank/registers_reg[10][23]  ( .D(\Reg_Bank/n3339 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][23] ) );
  DFF \Reg_Bank/registers_reg[10][24]  ( .D(\Reg_Bank/n3340 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][24] ) );
  DFF \Reg_Bank/registers_reg[10][25]  ( .D(\Reg_Bank/n3341 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][25] ) );
  DFF \Reg_Bank/registers_reg[10][26]  ( .D(\Reg_Bank/n3342 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][26] ) );
  DFF \Reg_Bank/registers_reg[10][27]  ( .D(\Reg_Bank/n3343 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][27] ) );
  DFF \Reg_Bank/registers_reg[10][28]  ( .D(\Reg_Bank/n3344 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][28] ) );
  DFF \Reg_Bank/registers_reg[10][29]  ( .D(\Reg_Bank/n3345 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][29] ) );
  DFF \Reg_Bank/registers_reg[10][30]  ( .D(\Reg_Bank/n3346 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][30] ) );
  DFF \Reg_Bank/registers_reg[10][31]  ( .D(\Reg_Bank/n3347 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[10][31] ) );
  DFF \Reg_Bank/registers_reg[11][0]  ( .D(\Reg_Bank/n3348 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][0] ) );
  DFF \Reg_Bank/registers_reg[11][1]  ( .D(\Reg_Bank/n3349 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][1] ) );
  DFF \Reg_Bank/registers_reg[11][2]  ( .D(\Reg_Bank/n3350 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][2] ) );
  DFF \Reg_Bank/registers_reg[11][3]  ( .D(\Reg_Bank/n3351 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][3] ) );
  DFF \Reg_Bank/registers_reg[11][4]  ( .D(\Reg_Bank/n3352 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][4] ) );
  DFF \Reg_Bank/registers_reg[11][5]  ( .D(\Reg_Bank/n3353 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][5] ) );
  DFF \Reg_Bank/registers_reg[11][6]  ( .D(\Reg_Bank/n3354 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][6] ) );
  DFF \Reg_Bank/registers_reg[11][7]  ( .D(\Reg_Bank/n3355 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][7] ) );
  DFF \Reg_Bank/registers_reg[11][8]  ( .D(\Reg_Bank/n3356 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][8] ) );
  DFF \Reg_Bank/registers_reg[11][9]  ( .D(\Reg_Bank/n3357 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[11][9] ) );
  DFF \Reg_Bank/registers_reg[11][10]  ( .D(\Reg_Bank/n3358 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][10] ) );
  DFF \Reg_Bank/registers_reg[11][11]  ( .D(\Reg_Bank/n3359 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][11] ) );
  DFF \Reg_Bank/registers_reg[11][12]  ( .D(\Reg_Bank/n3360 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][12] ) );
  DFF \Reg_Bank/registers_reg[11][13]  ( .D(\Reg_Bank/n3361 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][13] ) );
  DFF \Reg_Bank/registers_reg[11][14]  ( .D(\Reg_Bank/n3362 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][14] ) );
  DFF \Reg_Bank/registers_reg[11][15]  ( .D(\Reg_Bank/n3363 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][15] ) );
  DFF \Reg_Bank/registers_reg[11][16]  ( .D(\Reg_Bank/n3364 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][16] ) );
  DFF \Reg_Bank/registers_reg[11][17]  ( .D(\Reg_Bank/n3365 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][17] ) );
  DFF \Reg_Bank/registers_reg[11][18]  ( .D(\Reg_Bank/n3366 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][18] ) );
  DFF \Reg_Bank/registers_reg[11][19]  ( .D(\Reg_Bank/n3367 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][19] ) );
  DFF \Reg_Bank/registers_reg[11][20]  ( .D(\Reg_Bank/n3368 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][20] ) );
  DFF \Reg_Bank/registers_reg[11][21]  ( .D(\Reg_Bank/n3369 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][21] ) );
  DFF \Reg_Bank/registers_reg[11][22]  ( .D(\Reg_Bank/n3370 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][22] ) );
  DFF \Reg_Bank/registers_reg[11][23]  ( .D(\Reg_Bank/n3371 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][23] ) );
  DFF \Reg_Bank/registers_reg[11][24]  ( .D(\Reg_Bank/n3372 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][24] ) );
  DFF \Reg_Bank/registers_reg[11][25]  ( .D(\Reg_Bank/n3373 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][25] ) );
  DFF \Reg_Bank/registers_reg[11][26]  ( .D(\Reg_Bank/n3374 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][26] ) );
  DFF \Reg_Bank/registers_reg[11][27]  ( .D(\Reg_Bank/n3375 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][27] ) );
  DFF \Reg_Bank/registers_reg[11][28]  ( .D(\Reg_Bank/n3376 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][28] ) );
  DFF \Reg_Bank/registers_reg[11][29]  ( .D(\Reg_Bank/n3377 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][29] ) );
  DFF \Reg_Bank/registers_reg[11][30]  ( .D(\Reg_Bank/n3378 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][30] ) );
  DFF \Reg_Bank/registers_reg[11][31]  ( .D(\Reg_Bank/n3379 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[11][31] ) );
  DFF \Reg_Bank/registers_reg[12][0]  ( .D(\Reg_Bank/n3380 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][0] ) );
  DFF \Reg_Bank/registers_reg[12][1]  ( .D(\Reg_Bank/n3381 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][1] ) );
  DFF \Reg_Bank/registers_reg[12][2]  ( .D(\Reg_Bank/n3382 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][2] ) );
  DFF \Reg_Bank/registers_reg[12][3]  ( .D(\Reg_Bank/n3383 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][3] ) );
  DFF \Reg_Bank/registers_reg[12][4]  ( .D(\Reg_Bank/n3384 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][4] ) );
  DFF \Reg_Bank/registers_reg[12][5]  ( .D(\Reg_Bank/n3385 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][5] ) );
  DFF \Reg_Bank/registers_reg[12][6]  ( .D(\Reg_Bank/n3386 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][6] ) );
  DFF \Reg_Bank/registers_reg[12][7]  ( .D(\Reg_Bank/n3387 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][7] ) );
  DFF \Reg_Bank/registers_reg[12][8]  ( .D(\Reg_Bank/n3388 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][8] ) );
  DFF \Reg_Bank/registers_reg[12][9]  ( .D(\Reg_Bank/n3389 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[12][9] ) );
  DFF \Reg_Bank/registers_reg[12][10]  ( .D(\Reg_Bank/n3390 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][10] ) );
  DFF \Reg_Bank/registers_reg[12][11]  ( .D(\Reg_Bank/n3391 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][11] ) );
  DFF \Reg_Bank/registers_reg[12][12]  ( .D(\Reg_Bank/n3392 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][12] ) );
  DFF \Reg_Bank/registers_reg[12][13]  ( .D(\Reg_Bank/n3393 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][13] ) );
  DFF \Reg_Bank/registers_reg[12][14]  ( .D(\Reg_Bank/n3394 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][14] ) );
  DFF \Reg_Bank/registers_reg[12][15]  ( .D(\Reg_Bank/n3395 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][15] ) );
  DFF \Reg_Bank/registers_reg[12][16]  ( .D(\Reg_Bank/n3396 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][16] ) );
  DFF \Reg_Bank/registers_reg[12][17]  ( .D(\Reg_Bank/n3397 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][17] ) );
  DFF \Reg_Bank/registers_reg[12][18]  ( .D(\Reg_Bank/n3398 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][18] ) );
  DFF \Reg_Bank/registers_reg[12][19]  ( .D(\Reg_Bank/n3399 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][19] ) );
  DFF \Reg_Bank/registers_reg[12][20]  ( .D(\Reg_Bank/n3400 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][20] ) );
  DFF \Reg_Bank/registers_reg[12][21]  ( .D(\Reg_Bank/n3401 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][21] ) );
  DFF \Reg_Bank/registers_reg[12][22]  ( .D(\Reg_Bank/n3402 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][22] ) );
  DFF \Reg_Bank/registers_reg[12][23]  ( .D(\Reg_Bank/n3403 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][23] ) );
  DFF \Reg_Bank/registers_reg[12][24]  ( .D(\Reg_Bank/n3404 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][24] ) );
  DFF \Reg_Bank/registers_reg[12][25]  ( .D(\Reg_Bank/n3405 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][25] ) );
  DFF \Reg_Bank/registers_reg[12][26]  ( .D(\Reg_Bank/n3406 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][26] ) );
  DFF \Reg_Bank/registers_reg[12][27]  ( .D(\Reg_Bank/n3407 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][27] ) );
  DFF \Reg_Bank/registers_reg[12][28]  ( .D(\Reg_Bank/n3408 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][28] ) );
  DFF \Reg_Bank/registers_reg[12][29]  ( .D(\Reg_Bank/n3409 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][29] ) );
  DFF \Reg_Bank/registers_reg[12][30]  ( .D(\Reg_Bank/n3410 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][30] ) );
  DFF \Reg_Bank/registers_reg[12][31]  ( .D(\Reg_Bank/n3411 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[12][31] ) );
  DFF \Reg_Bank/registers_reg[13][0]  ( .D(\Reg_Bank/n3412 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][0] ) );
  DFF \Reg_Bank/registers_reg[13][1]  ( .D(\Reg_Bank/n3413 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][1] ) );
  DFF \Reg_Bank/registers_reg[13][2]  ( .D(\Reg_Bank/n3414 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][2] ) );
  DFF \Reg_Bank/registers_reg[13][3]  ( .D(\Reg_Bank/n3415 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][3] ) );
  DFF \Reg_Bank/registers_reg[13][4]  ( .D(\Reg_Bank/n3416 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][4] ) );
  DFF \Reg_Bank/registers_reg[13][5]  ( .D(\Reg_Bank/n3417 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][5] ) );
  DFF \Reg_Bank/registers_reg[13][6]  ( .D(\Reg_Bank/n3418 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][6] ) );
  DFF \Reg_Bank/registers_reg[13][7]  ( .D(\Reg_Bank/n3419 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][7] ) );
  DFF \Reg_Bank/registers_reg[13][8]  ( .D(\Reg_Bank/n3420 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][8] ) );
  DFF \Reg_Bank/registers_reg[13][9]  ( .D(\Reg_Bank/n3421 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[13][9] ) );
  DFF \Reg_Bank/registers_reg[13][10]  ( .D(\Reg_Bank/n3422 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][10] ) );
  DFF \Reg_Bank/registers_reg[13][11]  ( .D(\Reg_Bank/n3423 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][11] ) );
  DFF \Reg_Bank/registers_reg[13][12]  ( .D(\Reg_Bank/n3424 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][12] ) );
  DFF \Reg_Bank/registers_reg[13][13]  ( .D(\Reg_Bank/n3425 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][13] ) );
  DFF \Reg_Bank/registers_reg[13][14]  ( .D(\Reg_Bank/n3426 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][14] ) );
  DFF \Reg_Bank/registers_reg[13][15]  ( .D(\Reg_Bank/n3427 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][15] ) );
  DFF \Reg_Bank/registers_reg[13][16]  ( .D(\Reg_Bank/n3428 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][16] ) );
  DFF \Reg_Bank/registers_reg[13][17]  ( .D(\Reg_Bank/n3429 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][17] ) );
  DFF \Reg_Bank/registers_reg[13][18]  ( .D(\Reg_Bank/n3430 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][18] ) );
  DFF \Reg_Bank/registers_reg[13][19]  ( .D(\Reg_Bank/n3431 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][19] ) );
  DFF \Reg_Bank/registers_reg[13][20]  ( .D(\Reg_Bank/n3432 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][20] ) );
  DFF \Reg_Bank/registers_reg[13][21]  ( .D(\Reg_Bank/n3433 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][21] ) );
  DFF \Reg_Bank/registers_reg[13][22]  ( .D(\Reg_Bank/n3434 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][22] ) );
  DFF \Reg_Bank/registers_reg[13][23]  ( .D(\Reg_Bank/n3435 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][23] ) );
  DFF \Reg_Bank/registers_reg[13][24]  ( .D(\Reg_Bank/n3436 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][24] ) );
  DFF \Reg_Bank/registers_reg[13][25]  ( .D(\Reg_Bank/n3437 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][25] ) );
  DFF \Reg_Bank/registers_reg[13][26]  ( .D(\Reg_Bank/n3438 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][26] ) );
  DFF \Reg_Bank/registers_reg[13][27]  ( .D(\Reg_Bank/n3439 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][27] ) );
  DFF \Reg_Bank/registers_reg[13][28]  ( .D(\Reg_Bank/n3440 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][28] ) );
  DFF \Reg_Bank/registers_reg[13][29]  ( .D(\Reg_Bank/n3441 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][29] ) );
  DFF \Reg_Bank/registers_reg[13][30]  ( .D(\Reg_Bank/n3442 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][30] ) );
  DFF \Reg_Bank/registers_reg[13][31]  ( .D(\Reg_Bank/n3443 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[13][31] ) );
  DFF \Reg_Bank/registers_reg[14][0]  ( .D(\Reg_Bank/n3444 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][0] ) );
  DFF \Reg_Bank/registers_reg[14][1]  ( .D(\Reg_Bank/n3445 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][1] ) );
  DFF \Reg_Bank/registers_reg[14][2]  ( .D(\Reg_Bank/n3446 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][2] ) );
  DFF \Reg_Bank/registers_reg[14][3]  ( .D(\Reg_Bank/n3447 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][3] ) );
  DFF \Reg_Bank/registers_reg[14][4]  ( .D(\Reg_Bank/n3448 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][4] ) );
  DFF \Reg_Bank/registers_reg[14][5]  ( .D(\Reg_Bank/n3449 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][5] ) );
  DFF \Reg_Bank/registers_reg[14][6]  ( .D(\Reg_Bank/n3450 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][6] ) );
  DFF \Reg_Bank/registers_reg[14][7]  ( .D(\Reg_Bank/n3451 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][7] ) );
  DFF \Reg_Bank/registers_reg[14][8]  ( .D(\Reg_Bank/n3452 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][8] ) );
  DFF \Reg_Bank/registers_reg[14][9]  ( .D(\Reg_Bank/n3453 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[14][9] ) );
  DFF \Reg_Bank/registers_reg[14][10]  ( .D(\Reg_Bank/n3454 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][10] ) );
  DFF \Reg_Bank/registers_reg[14][11]  ( .D(\Reg_Bank/n3455 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][11] ) );
  DFF \Reg_Bank/registers_reg[14][12]  ( .D(\Reg_Bank/n3456 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][12] ) );
  DFF \Reg_Bank/registers_reg[14][13]  ( .D(\Reg_Bank/n3457 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][13] ) );
  DFF \Reg_Bank/registers_reg[14][14]  ( .D(\Reg_Bank/n3458 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][14] ) );
  DFF \Reg_Bank/registers_reg[14][15]  ( .D(\Reg_Bank/n3459 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][15] ) );
  DFF \Reg_Bank/registers_reg[14][16]  ( .D(\Reg_Bank/n3460 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][16] ) );
  DFF \Reg_Bank/registers_reg[14][17]  ( .D(\Reg_Bank/n3461 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][17] ) );
  DFF \Reg_Bank/registers_reg[14][18]  ( .D(\Reg_Bank/n3462 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][18] ) );
  DFF \Reg_Bank/registers_reg[14][19]  ( .D(\Reg_Bank/n3463 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][19] ) );
  DFF \Reg_Bank/registers_reg[14][20]  ( .D(\Reg_Bank/n3464 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][20] ) );
  DFF \Reg_Bank/registers_reg[14][21]  ( .D(\Reg_Bank/n3465 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][21] ) );
  DFF \Reg_Bank/registers_reg[14][22]  ( .D(\Reg_Bank/n3466 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][22] ) );
  DFF \Reg_Bank/registers_reg[14][23]  ( .D(\Reg_Bank/n3467 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][23] ) );
  DFF \Reg_Bank/registers_reg[14][24]  ( .D(\Reg_Bank/n3468 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][24] ) );
  DFF \Reg_Bank/registers_reg[14][25]  ( .D(\Reg_Bank/n3469 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][25] ) );
  DFF \Reg_Bank/registers_reg[14][26]  ( .D(\Reg_Bank/n3470 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][26] ) );
  DFF \Reg_Bank/registers_reg[14][27]  ( .D(\Reg_Bank/n3471 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][27] ) );
  DFF \Reg_Bank/registers_reg[14][28]  ( .D(\Reg_Bank/n3472 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][28] ) );
  DFF \Reg_Bank/registers_reg[14][29]  ( .D(\Reg_Bank/n3473 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][29] ) );
  DFF \Reg_Bank/registers_reg[14][30]  ( .D(\Reg_Bank/n3474 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][30] ) );
  DFF \Reg_Bank/registers_reg[14][31]  ( .D(\Reg_Bank/n3475 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[14][31] ) );
  DFF \Reg_Bank/registers_reg[15][0]  ( .D(\Reg_Bank/n3476 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][0] ) );
  DFF \Reg_Bank/registers_reg[15][1]  ( .D(\Reg_Bank/n3477 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][1] ) );
  DFF \Reg_Bank/registers_reg[15][2]  ( .D(\Reg_Bank/n3478 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][2] ) );
  DFF \Reg_Bank/registers_reg[15][3]  ( .D(\Reg_Bank/n3479 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][3] ) );
  DFF \Reg_Bank/registers_reg[15][4]  ( .D(\Reg_Bank/n3480 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][4] ) );
  DFF \Reg_Bank/registers_reg[15][5]  ( .D(\Reg_Bank/n3481 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][5] ) );
  DFF \Reg_Bank/registers_reg[15][6]  ( .D(\Reg_Bank/n3482 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][6] ) );
  DFF \Reg_Bank/registers_reg[15][7]  ( .D(\Reg_Bank/n3483 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][7] ) );
  DFF \Reg_Bank/registers_reg[15][8]  ( .D(\Reg_Bank/n3484 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][8] ) );
  DFF \Reg_Bank/registers_reg[15][9]  ( .D(\Reg_Bank/n3485 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[15][9] ) );
  DFF \Reg_Bank/registers_reg[15][10]  ( .D(\Reg_Bank/n3486 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][10] ) );
  DFF \Reg_Bank/registers_reg[15][11]  ( .D(\Reg_Bank/n3487 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][11] ) );
  DFF \Reg_Bank/registers_reg[15][12]  ( .D(\Reg_Bank/n3488 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][12] ) );
  DFF \Reg_Bank/registers_reg[15][13]  ( .D(\Reg_Bank/n3489 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][13] ) );
  DFF \Reg_Bank/registers_reg[15][14]  ( .D(\Reg_Bank/n3490 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][14] ) );
  DFF \Reg_Bank/registers_reg[15][15]  ( .D(\Reg_Bank/n3491 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][15] ) );
  DFF \Reg_Bank/registers_reg[15][16]  ( .D(\Reg_Bank/n3492 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][16] ) );
  DFF \Reg_Bank/registers_reg[15][17]  ( .D(\Reg_Bank/n3493 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][17] ) );
  DFF \Reg_Bank/registers_reg[15][18]  ( .D(\Reg_Bank/n3494 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][18] ) );
  DFF \Reg_Bank/registers_reg[15][19]  ( .D(\Reg_Bank/n3495 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][19] ) );
  DFF \Reg_Bank/registers_reg[15][20]  ( .D(\Reg_Bank/n3496 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][20] ) );
  DFF \Reg_Bank/registers_reg[15][21]  ( .D(\Reg_Bank/n3497 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][21] ) );
  DFF \Reg_Bank/registers_reg[15][22]  ( .D(\Reg_Bank/n3498 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][22] ) );
  DFF \Reg_Bank/registers_reg[15][23]  ( .D(\Reg_Bank/n3499 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][23] ) );
  DFF \Reg_Bank/registers_reg[15][24]  ( .D(\Reg_Bank/n3500 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][24] ) );
  DFF \Reg_Bank/registers_reg[15][25]  ( .D(\Reg_Bank/n3501 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][25] ) );
  DFF \Reg_Bank/registers_reg[15][26]  ( .D(\Reg_Bank/n3502 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][26] ) );
  DFF \Reg_Bank/registers_reg[15][27]  ( .D(\Reg_Bank/n3503 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][27] ) );
  DFF \Reg_Bank/registers_reg[15][28]  ( .D(\Reg_Bank/n3504 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][28] ) );
  DFF \Reg_Bank/registers_reg[15][29]  ( .D(\Reg_Bank/n3505 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][29] ) );
  DFF \Reg_Bank/registers_reg[15][30]  ( .D(\Reg_Bank/n3506 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][30] ) );
  DFF \Reg_Bank/registers_reg[15][31]  ( .D(\Reg_Bank/n3507 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[15][31] ) );
  DFF \Reg_Bank/registers_reg[16][0]  ( .D(\Reg_Bank/n3508 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][0] ) );
  DFF \Reg_Bank/registers_reg[16][1]  ( .D(\Reg_Bank/n3509 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][1] ) );
  DFF \Reg_Bank/registers_reg[16][2]  ( .D(\Reg_Bank/n3510 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][2] ) );
  DFF \Reg_Bank/registers_reg[16][3]  ( .D(\Reg_Bank/n3511 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][3] ) );
  DFF \Reg_Bank/registers_reg[16][4]  ( .D(\Reg_Bank/n3512 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][4] ) );
  DFF \Reg_Bank/registers_reg[16][5]  ( .D(\Reg_Bank/n3513 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][5] ) );
  DFF \Reg_Bank/registers_reg[16][6]  ( .D(\Reg_Bank/n3514 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][6] ) );
  DFF \Reg_Bank/registers_reg[16][7]  ( .D(\Reg_Bank/n3515 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][7] ) );
  DFF \Reg_Bank/registers_reg[16][8]  ( .D(\Reg_Bank/n3516 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][8] ) );
  DFF \Reg_Bank/registers_reg[16][9]  ( .D(\Reg_Bank/n3517 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[16][9] ) );
  DFF \Reg_Bank/registers_reg[16][10]  ( .D(\Reg_Bank/n3518 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][10] ) );
  DFF \Reg_Bank/registers_reg[16][11]  ( .D(\Reg_Bank/n3519 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][11] ) );
  DFF \Reg_Bank/registers_reg[16][12]  ( .D(\Reg_Bank/n3520 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][12] ) );
  DFF \Reg_Bank/registers_reg[16][13]  ( .D(\Reg_Bank/n3521 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][13] ) );
  DFF \Reg_Bank/registers_reg[16][14]  ( .D(\Reg_Bank/n3522 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][14] ) );
  DFF \Reg_Bank/registers_reg[16][15]  ( .D(\Reg_Bank/n3523 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][15] ) );
  DFF \Reg_Bank/registers_reg[16][16]  ( .D(\Reg_Bank/n3524 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][16] ) );
  DFF \Reg_Bank/registers_reg[16][17]  ( .D(\Reg_Bank/n3525 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][17] ) );
  DFF \Reg_Bank/registers_reg[16][18]  ( .D(\Reg_Bank/n3526 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][18] ) );
  DFF \Reg_Bank/registers_reg[16][19]  ( .D(\Reg_Bank/n3527 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][19] ) );
  DFF \Reg_Bank/registers_reg[16][20]  ( .D(\Reg_Bank/n3528 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][20] ) );
  DFF \Reg_Bank/registers_reg[16][21]  ( .D(\Reg_Bank/n3529 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][21] ) );
  DFF \Reg_Bank/registers_reg[16][22]  ( .D(\Reg_Bank/n3530 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][22] ) );
  DFF \Reg_Bank/registers_reg[16][23]  ( .D(\Reg_Bank/n3531 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][23] ) );
  DFF \Reg_Bank/registers_reg[16][24]  ( .D(\Reg_Bank/n3532 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][24] ) );
  DFF \Reg_Bank/registers_reg[16][25]  ( .D(\Reg_Bank/n3533 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][25] ) );
  DFF \Reg_Bank/registers_reg[16][26]  ( .D(\Reg_Bank/n3534 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][26] ) );
  DFF \Reg_Bank/registers_reg[16][27]  ( .D(\Reg_Bank/n3535 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][27] ) );
  DFF \Reg_Bank/registers_reg[16][28]  ( .D(\Reg_Bank/n3536 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][28] ) );
  DFF \Reg_Bank/registers_reg[16][29]  ( .D(\Reg_Bank/n3537 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][29] ) );
  DFF \Reg_Bank/registers_reg[16][30]  ( .D(\Reg_Bank/n3538 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][30] ) );
  DFF \Reg_Bank/registers_reg[16][31]  ( .D(\Reg_Bank/n3539 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[16][31] ) );
  DFF \Reg_Bank/registers_reg[17][0]  ( .D(\Reg_Bank/n3540 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][0] ) );
  DFF \Reg_Bank/registers_reg[17][1]  ( .D(\Reg_Bank/n3541 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][1] ) );
  DFF \Reg_Bank/registers_reg[17][2]  ( .D(\Reg_Bank/n3542 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][2] ) );
  DFF \Reg_Bank/registers_reg[17][3]  ( .D(\Reg_Bank/n3543 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][3] ) );
  DFF \Reg_Bank/registers_reg[17][4]  ( .D(\Reg_Bank/n3544 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][4] ) );
  DFF \Reg_Bank/registers_reg[17][5]  ( .D(\Reg_Bank/n3545 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][5] ) );
  DFF \Reg_Bank/registers_reg[17][6]  ( .D(\Reg_Bank/n3546 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][6] ) );
  DFF \Reg_Bank/registers_reg[17][7]  ( .D(\Reg_Bank/n3547 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][7] ) );
  DFF \Reg_Bank/registers_reg[17][8]  ( .D(\Reg_Bank/n3548 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][8] ) );
  DFF \Reg_Bank/registers_reg[17][9]  ( .D(\Reg_Bank/n3549 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[17][9] ) );
  DFF \Reg_Bank/registers_reg[17][10]  ( .D(\Reg_Bank/n3550 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][10] ) );
  DFF \Reg_Bank/registers_reg[17][11]  ( .D(\Reg_Bank/n3551 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][11] ) );
  DFF \Reg_Bank/registers_reg[17][12]  ( .D(\Reg_Bank/n3552 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][12] ) );
  DFF \Reg_Bank/registers_reg[17][13]  ( .D(\Reg_Bank/n3553 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][13] ) );
  DFF \Reg_Bank/registers_reg[17][14]  ( .D(\Reg_Bank/n3554 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][14] ) );
  DFF \Reg_Bank/registers_reg[17][15]  ( .D(\Reg_Bank/n3555 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][15] ) );
  DFF \Reg_Bank/registers_reg[17][16]  ( .D(\Reg_Bank/n3556 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][16] ) );
  DFF \Reg_Bank/registers_reg[17][17]  ( .D(\Reg_Bank/n3557 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][17] ) );
  DFF \Reg_Bank/registers_reg[17][18]  ( .D(\Reg_Bank/n3558 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][18] ) );
  DFF \Reg_Bank/registers_reg[17][19]  ( .D(\Reg_Bank/n3559 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][19] ) );
  DFF \Reg_Bank/registers_reg[17][20]  ( .D(\Reg_Bank/n3560 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][20] ) );
  DFF \Reg_Bank/registers_reg[17][21]  ( .D(\Reg_Bank/n3561 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][21] ) );
  DFF \Reg_Bank/registers_reg[17][22]  ( .D(\Reg_Bank/n3562 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][22] ) );
  DFF \Reg_Bank/registers_reg[17][23]  ( .D(\Reg_Bank/n3563 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][23] ) );
  DFF \Reg_Bank/registers_reg[17][24]  ( .D(\Reg_Bank/n3564 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][24] ) );
  DFF \Reg_Bank/registers_reg[17][25]  ( .D(\Reg_Bank/n3565 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][25] ) );
  DFF \Reg_Bank/registers_reg[17][26]  ( .D(\Reg_Bank/n3566 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][26] ) );
  DFF \Reg_Bank/registers_reg[17][27]  ( .D(\Reg_Bank/n3567 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][27] ) );
  DFF \Reg_Bank/registers_reg[17][28]  ( .D(\Reg_Bank/n3568 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][28] ) );
  DFF \Reg_Bank/registers_reg[17][29]  ( .D(\Reg_Bank/n3569 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][29] ) );
  DFF \Reg_Bank/registers_reg[17][30]  ( .D(\Reg_Bank/n3570 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][30] ) );
  DFF \Reg_Bank/registers_reg[17][31]  ( .D(\Reg_Bank/n3571 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[17][31] ) );
  DFF \Reg_Bank/registers_reg[18][0]  ( .D(\Reg_Bank/n3572 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][0] ) );
  DFF \Reg_Bank/registers_reg[18][1]  ( .D(\Reg_Bank/n3573 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][1] ) );
  DFF \Reg_Bank/registers_reg[18][2]  ( .D(\Reg_Bank/n3574 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][2] ) );
  DFF \Reg_Bank/registers_reg[18][3]  ( .D(\Reg_Bank/n3575 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][3] ) );
  DFF \Reg_Bank/registers_reg[18][4]  ( .D(\Reg_Bank/n3576 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][4] ) );
  DFF \Reg_Bank/registers_reg[18][5]  ( .D(\Reg_Bank/n3577 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][5] ) );
  DFF \Reg_Bank/registers_reg[18][6]  ( .D(\Reg_Bank/n3578 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][6] ) );
  DFF \Reg_Bank/registers_reg[18][7]  ( .D(\Reg_Bank/n3579 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][7] ) );
  DFF \Reg_Bank/registers_reg[18][8]  ( .D(\Reg_Bank/n3580 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][8] ) );
  DFF \Reg_Bank/registers_reg[18][9]  ( .D(\Reg_Bank/n3581 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[18][9] ) );
  DFF \Reg_Bank/registers_reg[18][10]  ( .D(\Reg_Bank/n3582 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][10] ) );
  DFF \Reg_Bank/registers_reg[18][11]  ( .D(\Reg_Bank/n3583 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][11] ) );
  DFF \Reg_Bank/registers_reg[18][12]  ( .D(\Reg_Bank/n3584 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][12] ) );
  DFF \Reg_Bank/registers_reg[18][13]  ( .D(\Reg_Bank/n3585 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][13] ) );
  DFF \Reg_Bank/registers_reg[18][14]  ( .D(\Reg_Bank/n3586 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][14] ) );
  DFF \Reg_Bank/registers_reg[18][15]  ( .D(\Reg_Bank/n3587 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][15] ) );
  DFF \Reg_Bank/registers_reg[18][16]  ( .D(\Reg_Bank/n3588 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][16] ) );
  DFF \Reg_Bank/registers_reg[18][17]  ( .D(\Reg_Bank/n3589 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][17] ) );
  DFF \Reg_Bank/registers_reg[18][18]  ( .D(\Reg_Bank/n3590 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][18] ) );
  DFF \Reg_Bank/registers_reg[18][19]  ( .D(\Reg_Bank/n3591 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][19] ) );
  DFF \Reg_Bank/registers_reg[18][20]  ( .D(\Reg_Bank/n3592 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][20] ) );
  DFF \Reg_Bank/registers_reg[18][21]  ( .D(\Reg_Bank/n3593 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][21] ) );
  DFF \Reg_Bank/registers_reg[18][22]  ( .D(\Reg_Bank/n3594 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][22] ) );
  DFF \Reg_Bank/registers_reg[18][23]  ( .D(\Reg_Bank/n3595 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][23] ) );
  DFF \Reg_Bank/registers_reg[18][24]  ( .D(\Reg_Bank/n3596 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][24] ) );
  DFF \Reg_Bank/registers_reg[18][25]  ( .D(\Reg_Bank/n3597 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][25] ) );
  DFF \Reg_Bank/registers_reg[18][26]  ( .D(\Reg_Bank/n3598 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][26] ) );
  DFF \Reg_Bank/registers_reg[18][27]  ( .D(\Reg_Bank/n3599 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][27] ) );
  DFF \Reg_Bank/registers_reg[18][28]  ( .D(\Reg_Bank/n3600 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][28] ) );
  DFF \Reg_Bank/registers_reg[18][29]  ( .D(\Reg_Bank/n3601 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][29] ) );
  DFF \Reg_Bank/registers_reg[18][30]  ( .D(\Reg_Bank/n3602 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][30] ) );
  DFF \Reg_Bank/registers_reg[18][31]  ( .D(\Reg_Bank/n3603 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[18][31] ) );
  DFF \Reg_Bank/registers_reg[19][0]  ( .D(\Reg_Bank/n3604 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][0] ) );
  DFF \Reg_Bank/registers_reg[19][1]  ( .D(\Reg_Bank/n3605 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][1] ) );
  DFF \Reg_Bank/registers_reg[19][2]  ( .D(\Reg_Bank/n3606 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][2] ) );
  DFF \Reg_Bank/registers_reg[19][3]  ( .D(\Reg_Bank/n3607 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][3] ) );
  DFF \Reg_Bank/registers_reg[19][4]  ( .D(\Reg_Bank/n3608 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][4] ) );
  DFF \Reg_Bank/registers_reg[19][5]  ( .D(\Reg_Bank/n3609 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][5] ) );
  DFF \Reg_Bank/registers_reg[19][6]  ( .D(\Reg_Bank/n3610 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][6] ) );
  DFF \Reg_Bank/registers_reg[19][7]  ( .D(\Reg_Bank/n3611 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][7] ) );
  DFF \Reg_Bank/registers_reg[19][8]  ( .D(\Reg_Bank/n3612 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][8] ) );
  DFF \Reg_Bank/registers_reg[19][9]  ( .D(\Reg_Bank/n3613 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[19][9] ) );
  DFF \Reg_Bank/registers_reg[19][10]  ( .D(\Reg_Bank/n3614 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][10] ) );
  DFF \Reg_Bank/registers_reg[19][11]  ( .D(\Reg_Bank/n3615 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][11] ) );
  DFF \Reg_Bank/registers_reg[19][12]  ( .D(\Reg_Bank/n3616 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][12] ) );
  DFF \Reg_Bank/registers_reg[19][13]  ( .D(\Reg_Bank/n3617 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][13] ) );
  DFF \Reg_Bank/registers_reg[19][14]  ( .D(\Reg_Bank/n3618 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][14] ) );
  DFF \Reg_Bank/registers_reg[19][15]  ( .D(\Reg_Bank/n3619 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][15] ) );
  DFF \Reg_Bank/registers_reg[19][16]  ( .D(\Reg_Bank/n3620 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][16] ) );
  DFF \Reg_Bank/registers_reg[19][17]  ( .D(\Reg_Bank/n3621 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][17] ) );
  DFF \Reg_Bank/registers_reg[19][18]  ( .D(\Reg_Bank/n3622 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][18] ) );
  DFF \Reg_Bank/registers_reg[19][19]  ( .D(\Reg_Bank/n3623 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][19] ) );
  DFF \Reg_Bank/registers_reg[19][20]  ( .D(\Reg_Bank/n3624 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][20] ) );
  DFF \Reg_Bank/registers_reg[19][21]  ( .D(\Reg_Bank/n3625 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][21] ) );
  DFF \Reg_Bank/registers_reg[19][22]  ( .D(\Reg_Bank/n3626 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][22] ) );
  DFF \Reg_Bank/registers_reg[19][23]  ( .D(\Reg_Bank/n3627 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][23] ) );
  DFF \Reg_Bank/registers_reg[19][24]  ( .D(\Reg_Bank/n3628 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][24] ) );
  DFF \Reg_Bank/registers_reg[19][25]  ( .D(\Reg_Bank/n3629 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][25] ) );
  DFF \Reg_Bank/registers_reg[19][26]  ( .D(\Reg_Bank/n3630 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][26] ) );
  DFF \Reg_Bank/registers_reg[19][27]  ( .D(\Reg_Bank/n3631 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][27] ) );
  DFF \Reg_Bank/registers_reg[19][28]  ( .D(\Reg_Bank/n3632 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][28] ) );
  DFF \Reg_Bank/registers_reg[19][29]  ( .D(\Reg_Bank/n3633 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][29] ) );
  DFF \Reg_Bank/registers_reg[19][30]  ( .D(\Reg_Bank/n3634 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][30] ) );
  DFF \Reg_Bank/registers_reg[19][31]  ( .D(\Reg_Bank/n3635 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[19][31] ) );
  DFF \Reg_Bank/registers_reg[20][0]  ( .D(\Reg_Bank/n3636 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][0] ) );
  DFF \Reg_Bank/registers_reg[20][1]  ( .D(\Reg_Bank/n3637 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][1] ) );
  DFF \Reg_Bank/registers_reg[20][2]  ( .D(\Reg_Bank/n3638 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][2] ) );
  DFF \Reg_Bank/registers_reg[20][3]  ( .D(\Reg_Bank/n3639 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][3] ) );
  DFF \Reg_Bank/registers_reg[20][4]  ( .D(\Reg_Bank/n3640 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][4] ) );
  DFF \Reg_Bank/registers_reg[20][5]  ( .D(\Reg_Bank/n3641 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][5] ) );
  DFF \Reg_Bank/registers_reg[20][6]  ( .D(\Reg_Bank/n3642 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][6] ) );
  DFF \Reg_Bank/registers_reg[20][7]  ( .D(\Reg_Bank/n3643 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][7] ) );
  DFF \Reg_Bank/registers_reg[20][8]  ( .D(\Reg_Bank/n3644 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][8] ) );
  DFF \Reg_Bank/registers_reg[20][9]  ( .D(\Reg_Bank/n3645 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[20][9] ) );
  DFF \Reg_Bank/registers_reg[20][10]  ( .D(\Reg_Bank/n3646 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][10] ) );
  DFF \Reg_Bank/registers_reg[20][11]  ( .D(\Reg_Bank/n3647 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][11] ) );
  DFF \Reg_Bank/registers_reg[20][12]  ( .D(\Reg_Bank/n3648 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][12] ) );
  DFF \Reg_Bank/registers_reg[20][13]  ( .D(\Reg_Bank/n3649 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][13] ) );
  DFF \Reg_Bank/registers_reg[20][14]  ( .D(\Reg_Bank/n3650 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][14] ) );
  DFF \Reg_Bank/registers_reg[20][15]  ( .D(\Reg_Bank/n3651 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][15] ) );
  DFF \Reg_Bank/registers_reg[20][16]  ( .D(\Reg_Bank/n3652 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][16] ) );
  DFF \Reg_Bank/registers_reg[20][17]  ( .D(\Reg_Bank/n3653 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][17] ) );
  DFF \Reg_Bank/registers_reg[20][18]  ( .D(\Reg_Bank/n3654 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][18] ) );
  DFF \Reg_Bank/registers_reg[20][19]  ( .D(\Reg_Bank/n3655 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][19] ) );
  DFF \Reg_Bank/registers_reg[20][20]  ( .D(\Reg_Bank/n3656 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][20] ) );
  DFF \Reg_Bank/registers_reg[20][21]  ( .D(\Reg_Bank/n3657 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][21] ) );
  DFF \Reg_Bank/registers_reg[20][22]  ( .D(\Reg_Bank/n3658 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][22] ) );
  DFF \Reg_Bank/registers_reg[20][23]  ( .D(\Reg_Bank/n3659 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][23] ) );
  DFF \Reg_Bank/registers_reg[20][24]  ( .D(\Reg_Bank/n3660 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][24] ) );
  DFF \Reg_Bank/registers_reg[20][25]  ( .D(\Reg_Bank/n3661 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][25] ) );
  DFF \Reg_Bank/registers_reg[20][26]  ( .D(\Reg_Bank/n3662 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][26] ) );
  DFF \Reg_Bank/registers_reg[20][27]  ( .D(\Reg_Bank/n3663 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][27] ) );
  DFF \Reg_Bank/registers_reg[20][28]  ( .D(\Reg_Bank/n3664 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][28] ) );
  DFF \Reg_Bank/registers_reg[20][29]  ( .D(\Reg_Bank/n3665 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][29] ) );
  DFF \Reg_Bank/registers_reg[20][30]  ( .D(\Reg_Bank/n3666 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][30] ) );
  DFF \Reg_Bank/registers_reg[20][31]  ( .D(\Reg_Bank/n3667 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[20][31] ) );
  DFF \Reg_Bank/registers_reg[21][0]  ( .D(\Reg_Bank/n3668 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][0] ) );
  DFF \Reg_Bank/registers_reg[21][1]  ( .D(\Reg_Bank/n3669 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][1] ) );
  DFF \Reg_Bank/registers_reg[21][2]  ( .D(\Reg_Bank/n3670 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][2] ) );
  DFF \Reg_Bank/registers_reg[21][3]  ( .D(\Reg_Bank/n3671 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][3] ) );
  DFF \Reg_Bank/registers_reg[21][4]  ( .D(\Reg_Bank/n3672 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][4] ) );
  DFF \Reg_Bank/registers_reg[21][5]  ( .D(\Reg_Bank/n3673 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][5] ) );
  DFF \Reg_Bank/registers_reg[21][6]  ( .D(\Reg_Bank/n3674 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][6] ) );
  DFF \Reg_Bank/registers_reg[21][7]  ( .D(\Reg_Bank/n3675 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][7] ) );
  DFF \Reg_Bank/registers_reg[21][8]  ( .D(\Reg_Bank/n3676 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][8] ) );
  DFF \Reg_Bank/registers_reg[21][9]  ( .D(\Reg_Bank/n3677 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[21][9] ) );
  DFF \Reg_Bank/registers_reg[21][10]  ( .D(\Reg_Bank/n3678 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][10] ) );
  DFF \Reg_Bank/registers_reg[21][11]  ( .D(\Reg_Bank/n3679 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][11] ) );
  DFF \Reg_Bank/registers_reg[21][12]  ( .D(\Reg_Bank/n3680 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][12] ) );
  DFF \Reg_Bank/registers_reg[21][13]  ( .D(\Reg_Bank/n3681 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][13] ) );
  DFF \Reg_Bank/registers_reg[21][14]  ( .D(\Reg_Bank/n3682 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][14] ) );
  DFF \Reg_Bank/registers_reg[21][15]  ( .D(\Reg_Bank/n3683 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][15] ) );
  DFF \Reg_Bank/registers_reg[21][16]  ( .D(\Reg_Bank/n3684 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][16] ) );
  DFF \Reg_Bank/registers_reg[21][17]  ( .D(\Reg_Bank/n3685 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][17] ) );
  DFF \Reg_Bank/registers_reg[21][18]  ( .D(\Reg_Bank/n3686 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][18] ) );
  DFF \Reg_Bank/registers_reg[21][19]  ( .D(\Reg_Bank/n3687 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][19] ) );
  DFF \Reg_Bank/registers_reg[21][20]  ( .D(\Reg_Bank/n3688 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][20] ) );
  DFF \Reg_Bank/registers_reg[21][21]  ( .D(\Reg_Bank/n3689 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][21] ) );
  DFF \Reg_Bank/registers_reg[21][22]  ( .D(\Reg_Bank/n3690 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][22] ) );
  DFF \Reg_Bank/registers_reg[21][23]  ( .D(\Reg_Bank/n3691 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][23] ) );
  DFF \Reg_Bank/registers_reg[21][24]  ( .D(\Reg_Bank/n3692 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][24] ) );
  DFF \Reg_Bank/registers_reg[21][25]  ( .D(\Reg_Bank/n3693 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][25] ) );
  DFF \Reg_Bank/registers_reg[21][26]  ( .D(\Reg_Bank/n3694 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][26] ) );
  DFF \Reg_Bank/registers_reg[21][27]  ( .D(\Reg_Bank/n3695 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][27] ) );
  DFF \Reg_Bank/registers_reg[21][28]  ( .D(\Reg_Bank/n3696 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][28] ) );
  DFF \Reg_Bank/registers_reg[21][29]  ( .D(\Reg_Bank/n3697 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][29] ) );
  DFF \Reg_Bank/registers_reg[21][30]  ( .D(\Reg_Bank/n3698 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][30] ) );
  DFF \Reg_Bank/registers_reg[21][31]  ( .D(\Reg_Bank/n3699 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[21][31] ) );
  DFF \Reg_Bank/registers_reg[22][0]  ( .D(\Reg_Bank/n3700 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][0] ) );
  DFF \Reg_Bank/registers_reg[22][1]  ( .D(\Reg_Bank/n3701 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][1] ) );
  DFF \Reg_Bank/registers_reg[22][2]  ( .D(\Reg_Bank/n3702 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][2] ) );
  DFF \Reg_Bank/registers_reg[22][3]  ( .D(\Reg_Bank/n3703 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][3] ) );
  DFF \Reg_Bank/registers_reg[22][4]  ( .D(\Reg_Bank/n3704 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][4] ) );
  DFF \Reg_Bank/registers_reg[22][5]  ( .D(\Reg_Bank/n3705 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][5] ) );
  DFF \Reg_Bank/registers_reg[22][6]  ( .D(\Reg_Bank/n3706 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][6] ) );
  DFF \Reg_Bank/registers_reg[22][7]  ( .D(\Reg_Bank/n3707 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][7] ) );
  DFF \Reg_Bank/registers_reg[22][8]  ( .D(\Reg_Bank/n3708 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][8] ) );
  DFF \Reg_Bank/registers_reg[22][9]  ( .D(\Reg_Bank/n3709 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[22][9] ) );
  DFF \Reg_Bank/registers_reg[22][10]  ( .D(\Reg_Bank/n3710 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][10] ) );
  DFF \Reg_Bank/registers_reg[22][11]  ( .D(\Reg_Bank/n3711 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][11] ) );
  DFF \Reg_Bank/registers_reg[22][12]  ( .D(\Reg_Bank/n3712 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][12] ) );
  DFF \Reg_Bank/registers_reg[22][13]  ( .D(\Reg_Bank/n3713 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][13] ) );
  DFF \Reg_Bank/registers_reg[22][14]  ( .D(\Reg_Bank/n3714 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][14] ) );
  DFF \Reg_Bank/registers_reg[22][15]  ( .D(\Reg_Bank/n3715 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][15] ) );
  DFF \Reg_Bank/registers_reg[22][16]  ( .D(\Reg_Bank/n3716 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][16] ) );
  DFF \Reg_Bank/registers_reg[22][17]  ( .D(\Reg_Bank/n3717 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][17] ) );
  DFF \Reg_Bank/registers_reg[22][18]  ( .D(\Reg_Bank/n3718 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][18] ) );
  DFF \Reg_Bank/registers_reg[22][19]  ( .D(\Reg_Bank/n3719 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][19] ) );
  DFF \Reg_Bank/registers_reg[22][20]  ( .D(\Reg_Bank/n3720 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][20] ) );
  DFF \Reg_Bank/registers_reg[22][21]  ( .D(\Reg_Bank/n3721 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][21] ) );
  DFF \Reg_Bank/registers_reg[22][22]  ( .D(\Reg_Bank/n3722 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][22] ) );
  DFF \Reg_Bank/registers_reg[22][23]  ( .D(\Reg_Bank/n3723 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][23] ) );
  DFF \Reg_Bank/registers_reg[22][24]  ( .D(\Reg_Bank/n3724 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][24] ) );
  DFF \Reg_Bank/registers_reg[22][25]  ( .D(\Reg_Bank/n3725 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][25] ) );
  DFF \Reg_Bank/registers_reg[22][26]  ( .D(\Reg_Bank/n3726 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][26] ) );
  DFF \Reg_Bank/registers_reg[22][27]  ( .D(\Reg_Bank/n3727 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][27] ) );
  DFF \Reg_Bank/registers_reg[22][28]  ( .D(\Reg_Bank/n3728 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][28] ) );
  DFF \Reg_Bank/registers_reg[22][29]  ( .D(\Reg_Bank/n3729 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][29] ) );
  DFF \Reg_Bank/registers_reg[22][30]  ( .D(\Reg_Bank/n3730 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][30] ) );
  DFF \Reg_Bank/registers_reg[22][31]  ( .D(\Reg_Bank/n3731 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[22][31] ) );
  DFF \Reg_Bank/registers_reg[23][0]  ( .D(\Reg_Bank/n3732 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][0] ) );
  DFF \Reg_Bank/registers_reg[23][1]  ( .D(\Reg_Bank/n3733 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][1] ) );
  DFF \Reg_Bank/registers_reg[23][2]  ( .D(\Reg_Bank/n3734 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][2] ) );
  DFF \Reg_Bank/registers_reg[23][3]  ( .D(\Reg_Bank/n3735 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][3] ) );
  DFF \Reg_Bank/registers_reg[23][4]  ( .D(\Reg_Bank/n3736 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][4] ) );
  DFF \Reg_Bank/registers_reg[23][5]  ( .D(\Reg_Bank/n3737 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][5] ) );
  DFF \Reg_Bank/registers_reg[23][6]  ( .D(\Reg_Bank/n3738 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][6] ) );
  DFF \Reg_Bank/registers_reg[23][7]  ( .D(\Reg_Bank/n3739 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][7] ) );
  DFF \Reg_Bank/registers_reg[23][8]  ( .D(\Reg_Bank/n3740 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][8] ) );
  DFF \Reg_Bank/registers_reg[23][9]  ( .D(\Reg_Bank/n3741 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[23][9] ) );
  DFF \Reg_Bank/registers_reg[23][10]  ( .D(\Reg_Bank/n3742 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][10] ) );
  DFF \Reg_Bank/registers_reg[23][11]  ( .D(\Reg_Bank/n3743 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][11] ) );
  DFF \Reg_Bank/registers_reg[23][12]  ( .D(\Reg_Bank/n3744 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][12] ) );
  DFF \Reg_Bank/registers_reg[23][13]  ( .D(\Reg_Bank/n3745 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][13] ) );
  DFF \Reg_Bank/registers_reg[23][14]  ( .D(\Reg_Bank/n3746 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][14] ) );
  DFF \Reg_Bank/registers_reg[23][15]  ( .D(\Reg_Bank/n3747 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][15] ) );
  DFF \Reg_Bank/registers_reg[23][16]  ( .D(\Reg_Bank/n3748 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][16] ) );
  DFF \Reg_Bank/registers_reg[23][17]  ( .D(\Reg_Bank/n3749 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][17] ) );
  DFF \Reg_Bank/registers_reg[23][18]  ( .D(\Reg_Bank/n3750 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][18] ) );
  DFF \Reg_Bank/registers_reg[23][19]  ( .D(\Reg_Bank/n3751 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][19] ) );
  DFF \Reg_Bank/registers_reg[23][20]  ( .D(\Reg_Bank/n3752 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][20] ) );
  DFF \Reg_Bank/registers_reg[23][21]  ( .D(\Reg_Bank/n3753 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][21] ) );
  DFF \Reg_Bank/registers_reg[23][22]  ( .D(\Reg_Bank/n3754 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][22] ) );
  DFF \Reg_Bank/registers_reg[23][23]  ( .D(\Reg_Bank/n3755 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][23] ) );
  DFF \Reg_Bank/registers_reg[23][24]  ( .D(\Reg_Bank/n3756 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][24] ) );
  DFF \Reg_Bank/registers_reg[23][25]  ( .D(\Reg_Bank/n3757 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][25] ) );
  DFF \Reg_Bank/registers_reg[23][26]  ( .D(\Reg_Bank/n3758 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][26] ) );
  DFF \Reg_Bank/registers_reg[23][27]  ( .D(\Reg_Bank/n3759 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][27] ) );
  DFF \Reg_Bank/registers_reg[23][28]  ( .D(\Reg_Bank/n3760 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][28] ) );
  DFF \Reg_Bank/registers_reg[23][29]  ( .D(\Reg_Bank/n3761 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][29] ) );
  DFF \Reg_Bank/registers_reg[23][30]  ( .D(\Reg_Bank/n3762 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][30] ) );
  DFF \Reg_Bank/registers_reg[23][31]  ( .D(\Reg_Bank/n3763 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[23][31] ) );
  DFF \Reg_Bank/registers_reg[24][0]  ( .D(\Reg_Bank/n3764 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][0] ) );
  DFF \Reg_Bank/registers_reg[24][1]  ( .D(\Reg_Bank/n3765 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][1] ) );
  DFF \Reg_Bank/registers_reg[24][2]  ( .D(\Reg_Bank/n3766 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][2] ) );
  DFF \Reg_Bank/registers_reg[24][3]  ( .D(\Reg_Bank/n3767 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][3] ) );
  DFF \Reg_Bank/registers_reg[24][4]  ( .D(\Reg_Bank/n3768 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][4] ) );
  DFF \Reg_Bank/registers_reg[24][5]  ( .D(\Reg_Bank/n3769 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][5] ) );
  DFF \Reg_Bank/registers_reg[24][6]  ( .D(\Reg_Bank/n3770 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][6] ) );
  DFF \Reg_Bank/registers_reg[24][7]  ( .D(\Reg_Bank/n3771 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][7] ) );
  DFF \Reg_Bank/registers_reg[24][8]  ( .D(\Reg_Bank/n3772 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][8] ) );
  DFF \Reg_Bank/registers_reg[24][9]  ( .D(\Reg_Bank/n3773 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[24][9] ) );
  DFF \Reg_Bank/registers_reg[24][10]  ( .D(\Reg_Bank/n3774 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][10] ) );
  DFF \Reg_Bank/registers_reg[24][11]  ( .D(\Reg_Bank/n3775 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][11] ) );
  DFF \Reg_Bank/registers_reg[24][12]  ( .D(\Reg_Bank/n3776 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][12] ) );
  DFF \Reg_Bank/registers_reg[24][13]  ( .D(\Reg_Bank/n3777 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][13] ) );
  DFF \Reg_Bank/registers_reg[24][14]  ( .D(\Reg_Bank/n3778 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][14] ) );
  DFF \Reg_Bank/registers_reg[24][15]  ( .D(\Reg_Bank/n3779 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][15] ) );
  DFF \Reg_Bank/registers_reg[24][16]  ( .D(\Reg_Bank/n3780 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][16] ) );
  DFF \Reg_Bank/registers_reg[24][17]  ( .D(\Reg_Bank/n3781 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][17] ) );
  DFF \Reg_Bank/registers_reg[24][18]  ( .D(\Reg_Bank/n3782 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][18] ) );
  DFF \Reg_Bank/registers_reg[24][19]  ( .D(\Reg_Bank/n3783 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][19] ) );
  DFF \Reg_Bank/registers_reg[24][20]  ( .D(\Reg_Bank/n3784 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][20] ) );
  DFF \Reg_Bank/registers_reg[24][21]  ( .D(\Reg_Bank/n3785 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][21] ) );
  DFF \Reg_Bank/registers_reg[24][22]  ( .D(\Reg_Bank/n3786 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][22] ) );
  DFF \Reg_Bank/registers_reg[24][23]  ( .D(\Reg_Bank/n3787 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][23] ) );
  DFF \Reg_Bank/registers_reg[24][24]  ( .D(\Reg_Bank/n3788 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][24] ) );
  DFF \Reg_Bank/registers_reg[24][25]  ( .D(\Reg_Bank/n3789 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][25] ) );
  DFF \Reg_Bank/registers_reg[24][26]  ( .D(\Reg_Bank/n3790 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][26] ) );
  DFF \Reg_Bank/registers_reg[24][27]  ( .D(\Reg_Bank/n3791 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][27] ) );
  DFF \Reg_Bank/registers_reg[24][28]  ( .D(\Reg_Bank/n3792 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][28] ) );
  DFF \Reg_Bank/registers_reg[24][29]  ( .D(\Reg_Bank/n3793 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][29] ) );
  DFF \Reg_Bank/registers_reg[24][30]  ( .D(\Reg_Bank/n3794 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][30] ) );
  DFF \Reg_Bank/registers_reg[24][31]  ( .D(\Reg_Bank/n3795 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[24][31] ) );
  DFF \Reg_Bank/registers_reg[25][0]  ( .D(\Reg_Bank/n3796 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][0] ) );
  DFF \Reg_Bank/registers_reg[25][1]  ( .D(\Reg_Bank/n3797 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][1] ) );
  DFF \Reg_Bank/registers_reg[25][2]  ( .D(\Reg_Bank/n3798 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][2] ) );
  DFF \Reg_Bank/registers_reg[25][3]  ( .D(\Reg_Bank/n3799 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][3] ) );
  DFF \Reg_Bank/registers_reg[25][4]  ( .D(\Reg_Bank/n3800 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][4] ) );
  DFF \Reg_Bank/registers_reg[25][5]  ( .D(\Reg_Bank/n3801 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][5] ) );
  DFF \Reg_Bank/registers_reg[25][6]  ( .D(\Reg_Bank/n3802 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][6] ) );
  DFF \Reg_Bank/registers_reg[25][7]  ( .D(\Reg_Bank/n3803 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][7] ) );
  DFF \Reg_Bank/registers_reg[25][8]  ( .D(\Reg_Bank/n3804 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][8] ) );
  DFF \Reg_Bank/registers_reg[25][9]  ( .D(\Reg_Bank/n3805 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[25][9] ) );
  DFF \Reg_Bank/registers_reg[25][10]  ( .D(\Reg_Bank/n3806 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][10] ) );
  DFF \Reg_Bank/registers_reg[25][11]  ( .D(\Reg_Bank/n3807 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][11] ) );
  DFF \Reg_Bank/registers_reg[25][12]  ( .D(\Reg_Bank/n3808 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][12] ) );
  DFF \Reg_Bank/registers_reg[25][13]  ( .D(\Reg_Bank/n3809 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][13] ) );
  DFF \Reg_Bank/registers_reg[25][14]  ( .D(\Reg_Bank/n3810 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][14] ) );
  DFF \Reg_Bank/registers_reg[25][15]  ( .D(\Reg_Bank/n3811 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][15] ) );
  DFF \Reg_Bank/registers_reg[25][16]  ( .D(\Reg_Bank/n3812 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][16] ) );
  DFF \Reg_Bank/registers_reg[25][17]  ( .D(\Reg_Bank/n3813 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][17] ) );
  DFF \Reg_Bank/registers_reg[25][18]  ( .D(\Reg_Bank/n3814 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][18] ) );
  DFF \Reg_Bank/registers_reg[25][19]  ( .D(\Reg_Bank/n3815 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][19] ) );
  DFF \Reg_Bank/registers_reg[25][20]  ( .D(\Reg_Bank/n3816 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][20] ) );
  DFF \Reg_Bank/registers_reg[25][21]  ( .D(\Reg_Bank/n3817 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][21] ) );
  DFF \Reg_Bank/registers_reg[25][22]  ( .D(\Reg_Bank/n3818 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][22] ) );
  DFF \Reg_Bank/registers_reg[25][23]  ( .D(\Reg_Bank/n3819 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][23] ) );
  DFF \Reg_Bank/registers_reg[25][24]  ( .D(\Reg_Bank/n3820 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][24] ) );
  DFF \Reg_Bank/registers_reg[25][25]  ( .D(\Reg_Bank/n3821 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][25] ) );
  DFF \Reg_Bank/registers_reg[25][26]  ( .D(\Reg_Bank/n3822 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][26] ) );
  DFF \Reg_Bank/registers_reg[25][27]  ( .D(\Reg_Bank/n3823 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][27] ) );
  DFF \Reg_Bank/registers_reg[25][28]  ( .D(\Reg_Bank/n3824 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][28] ) );
  DFF \Reg_Bank/registers_reg[25][29]  ( .D(\Reg_Bank/n3825 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][29] ) );
  DFF \Reg_Bank/registers_reg[25][30]  ( .D(\Reg_Bank/n3826 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][30] ) );
  DFF \Reg_Bank/registers_reg[25][31]  ( .D(\Reg_Bank/n3827 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[25][31] ) );
  DFF \Reg_Bank/registers_reg[26][0]  ( .D(\Reg_Bank/n3828 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][0] ) );
  DFF \Reg_Bank/registers_reg[26][1]  ( .D(\Reg_Bank/n3829 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][1] ) );
  DFF \Reg_Bank/registers_reg[26][2]  ( .D(\Reg_Bank/n3830 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][2] ) );
  DFF \Reg_Bank/registers_reg[26][3]  ( .D(\Reg_Bank/n3831 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][3] ) );
  DFF \Reg_Bank/registers_reg[26][4]  ( .D(\Reg_Bank/n3832 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][4] ) );
  DFF \Reg_Bank/registers_reg[26][5]  ( .D(\Reg_Bank/n3833 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][5] ) );
  DFF \Reg_Bank/registers_reg[26][6]  ( .D(\Reg_Bank/n3834 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][6] ) );
  DFF \Reg_Bank/registers_reg[26][7]  ( .D(\Reg_Bank/n3835 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][7] ) );
  DFF \Reg_Bank/registers_reg[26][8]  ( .D(\Reg_Bank/n3836 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][8] ) );
  DFF \Reg_Bank/registers_reg[26][9]  ( .D(\Reg_Bank/n3837 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[26][9] ) );
  DFF \Reg_Bank/registers_reg[26][10]  ( .D(\Reg_Bank/n3838 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][10] ) );
  DFF \Reg_Bank/registers_reg[26][11]  ( .D(\Reg_Bank/n3839 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][11] ) );
  DFF \Reg_Bank/registers_reg[26][12]  ( .D(\Reg_Bank/n3840 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][12] ) );
  DFF \Reg_Bank/registers_reg[26][13]  ( .D(\Reg_Bank/n3841 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][13] ) );
  DFF \Reg_Bank/registers_reg[26][14]  ( .D(\Reg_Bank/n3842 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][14] ) );
  DFF \Reg_Bank/registers_reg[26][15]  ( .D(\Reg_Bank/n3843 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][15] ) );
  DFF \Reg_Bank/registers_reg[26][16]  ( .D(\Reg_Bank/n3844 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][16] ) );
  DFF \Reg_Bank/registers_reg[26][17]  ( .D(\Reg_Bank/n3845 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][17] ) );
  DFF \Reg_Bank/registers_reg[26][18]  ( .D(\Reg_Bank/n3846 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][18] ) );
  DFF \Reg_Bank/registers_reg[26][19]  ( .D(\Reg_Bank/n3847 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][19] ) );
  DFF \Reg_Bank/registers_reg[26][20]  ( .D(\Reg_Bank/n3848 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][20] ) );
  DFF \Reg_Bank/registers_reg[26][21]  ( .D(\Reg_Bank/n3849 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][21] ) );
  DFF \Reg_Bank/registers_reg[26][22]  ( .D(\Reg_Bank/n3850 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][22] ) );
  DFF \Reg_Bank/registers_reg[26][23]  ( .D(\Reg_Bank/n3851 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][23] ) );
  DFF \Reg_Bank/registers_reg[26][24]  ( .D(\Reg_Bank/n3852 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][24] ) );
  DFF \Reg_Bank/registers_reg[26][25]  ( .D(\Reg_Bank/n3853 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][25] ) );
  DFF \Reg_Bank/registers_reg[26][26]  ( .D(\Reg_Bank/n3854 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][26] ) );
  DFF \Reg_Bank/registers_reg[26][27]  ( .D(\Reg_Bank/n3855 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][27] ) );
  DFF \Reg_Bank/registers_reg[26][28]  ( .D(\Reg_Bank/n3856 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][28] ) );
  DFF \Reg_Bank/registers_reg[26][29]  ( .D(\Reg_Bank/n3857 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][29] ) );
  DFF \Reg_Bank/registers_reg[26][30]  ( .D(\Reg_Bank/n3858 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][30] ) );
  DFF \Reg_Bank/registers_reg[26][31]  ( .D(\Reg_Bank/n3859 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[26][31] ) );
  DFF \Reg_Bank/registers_reg[27][0]  ( .D(\Reg_Bank/n3860 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][0] ) );
  DFF \Reg_Bank/registers_reg[27][1]  ( .D(\Reg_Bank/n3861 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][1] ) );
  DFF \Reg_Bank/registers_reg[27][2]  ( .D(\Reg_Bank/n3862 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][2] ) );
  DFF \Reg_Bank/registers_reg[27][3]  ( .D(\Reg_Bank/n3863 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][3] ) );
  DFF \Reg_Bank/registers_reg[27][4]  ( .D(\Reg_Bank/n3864 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][4] ) );
  DFF \Reg_Bank/registers_reg[27][5]  ( .D(\Reg_Bank/n3865 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][5] ) );
  DFF \Reg_Bank/registers_reg[27][6]  ( .D(\Reg_Bank/n3866 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][6] ) );
  DFF \Reg_Bank/registers_reg[27][7]  ( .D(\Reg_Bank/n3867 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][7] ) );
  DFF \Reg_Bank/registers_reg[27][8]  ( .D(\Reg_Bank/n3868 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][8] ) );
  DFF \Reg_Bank/registers_reg[27][9]  ( .D(\Reg_Bank/n3869 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[27][9] ) );
  DFF \Reg_Bank/registers_reg[27][10]  ( .D(\Reg_Bank/n3870 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][10] ) );
  DFF \Reg_Bank/registers_reg[27][11]  ( .D(\Reg_Bank/n3871 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][11] ) );
  DFF \Reg_Bank/registers_reg[27][12]  ( .D(\Reg_Bank/n3872 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][12] ) );
  DFF \Reg_Bank/registers_reg[27][13]  ( .D(\Reg_Bank/n3873 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][13] ) );
  DFF \Reg_Bank/registers_reg[27][14]  ( .D(\Reg_Bank/n3874 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][14] ) );
  DFF \Reg_Bank/registers_reg[27][15]  ( .D(\Reg_Bank/n3875 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][15] ) );
  DFF \Reg_Bank/registers_reg[27][16]  ( .D(\Reg_Bank/n3876 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][16] ) );
  DFF \Reg_Bank/registers_reg[27][17]  ( .D(\Reg_Bank/n3877 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][17] ) );
  DFF \Reg_Bank/registers_reg[27][18]  ( .D(\Reg_Bank/n3878 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][18] ) );
  DFF \Reg_Bank/registers_reg[27][19]  ( .D(\Reg_Bank/n3879 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][19] ) );
  DFF \Reg_Bank/registers_reg[27][20]  ( .D(\Reg_Bank/n3880 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][20] ) );
  DFF \Reg_Bank/registers_reg[27][21]  ( .D(\Reg_Bank/n3881 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][21] ) );
  DFF \Reg_Bank/registers_reg[27][22]  ( .D(\Reg_Bank/n3882 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][22] ) );
  DFF \Reg_Bank/registers_reg[27][23]  ( .D(\Reg_Bank/n3883 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][23] ) );
  DFF \Reg_Bank/registers_reg[27][24]  ( .D(\Reg_Bank/n3884 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][24] ) );
  DFF \Reg_Bank/registers_reg[27][25]  ( .D(\Reg_Bank/n3885 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][25] ) );
  DFF \Reg_Bank/registers_reg[27][26]  ( .D(\Reg_Bank/n3886 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][26] ) );
  DFF \Reg_Bank/registers_reg[27][27]  ( .D(\Reg_Bank/n3887 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][27] ) );
  DFF \Reg_Bank/registers_reg[27][28]  ( .D(\Reg_Bank/n3888 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][28] ) );
  DFF \Reg_Bank/registers_reg[27][29]  ( .D(\Reg_Bank/n3889 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][29] ) );
  DFF \Reg_Bank/registers_reg[27][30]  ( .D(\Reg_Bank/n3890 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][30] ) );
  DFF \Reg_Bank/registers_reg[27][31]  ( .D(\Reg_Bank/n3891 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[27][31] ) );
  DFF \Reg_Bank/registers_reg[28][0]  ( .D(\Reg_Bank/n3892 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][0] ) );
  DFF \Reg_Bank/registers_reg[28][1]  ( .D(\Reg_Bank/n3893 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][1] ) );
  DFF \Reg_Bank/registers_reg[28][2]  ( .D(\Reg_Bank/n3894 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][2] ) );
  DFF \Reg_Bank/registers_reg[28][3]  ( .D(\Reg_Bank/n3895 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][3] ) );
  DFF \Reg_Bank/registers_reg[28][4]  ( .D(\Reg_Bank/n3896 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][4] ) );
  DFF \Reg_Bank/registers_reg[28][5]  ( .D(\Reg_Bank/n3897 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][5] ) );
  DFF \Reg_Bank/registers_reg[28][6]  ( .D(\Reg_Bank/n3898 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][6] ) );
  DFF \Reg_Bank/registers_reg[28][7]  ( .D(\Reg_Bank/n3899 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][7] ) );
  DFF \Reg_Bank/registers_reg[28][8]  ( .D(\Reg_Bank/n3900 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][8] ) );
  DFF \Reg_Bank/registers_reg[28][9]  ( .D(\Reg_Bank/n3901 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[28][9] ) );
  DFF \Reg_Bank/registers_reg[28][10]  ( .D(\Reg_Bank/n3902 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][10] ) );
  DFF \Reg_Bank/registers_reg[28][11]  ( .D(\Reg_Bank/n3903 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][11] ) );
  DFF \Reg_Bank/registers_reg[28][12]  ( .D(\Reg_Bank/n3904 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][12] ) );
  DFF \Reg_Bank/registers_reg[28][13]  ( .D(\Reg_Bank/n3905 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][13] ) );
  DFF \Reg_Bank/registers_reg[28][14]  ( .D(\Reg_Bank/n3906 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][14] ) );
  DFF \Reg_Bank/registers_reg[28][15]  ( .D(\Reg_Bank/n3907 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][15] ) );
  DFF \Reg_Bank/registers_reg[28][16]  ( .D(\Reg_Bank/n3908 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][16] ) );
  DFF \Reg_Bank/registers_reg[28][17]  ( .D(\Reg_Bank/n3909 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][17] ) );
  DFF \Reg_Bank/registers_reg[28][18]  ( .D(\Reg_Bank/n3910 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][18] ) );
  DFF \Reg_Bank/registers_reg[28][19]  ( .D(\Reg_Bank/n3911 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][19] ) );
  DFF \Reg_Bank/registers_reg[28][20]  ( .D(\Reg_Bank/n3912 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][20] ) );
  DFF \Reg_Bank/registers_reg[28][21]  ( .D(\Reg_Bank/n3913 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][21] ) );
  DFF \Reg_Bank/registers_reg[28][22]  ( .D(\Reg_Bank/n3914 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][22] ) );
  DFF \Reg_Bank/registers_reg[28][23]  ( .D(\Reg_Bank/n3915 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][23] ) );
  DFF \Reg_Bank/registers_reg[28][24]  ( .D(\Reg_Bank/n3916 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][24] ) );
  DFF \Reg_Bank/registers_reg[28][25]  ( .D(\Reg_Bank/n3917 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][25] ) );
  DFF \Reg_Bank/registers_reg[28][26]  ( .D(\Reg_Bank/n3918 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][26] ) );
  DFF \Reg_Bank/registers_reg[28][27]  ( .D(\Reg_Bank/n3919 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][27] ) );
  DFF \Reg_Bank/registers_reg[28][28]  ( .D(\Reg_Bank/n3920 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][28] ) );
  DFF \Reg_Bank/registers_reg[28][29]  ( .D(\Reg_Bank/n3921 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][29] ) );
  DFF \Reg_Bank/registers_reg[28][30]  ( .D(\Reg_Bank/n3922 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][30] ) );
  DFF \Reg_Bank/registers_reg[28][31]  ( .D(\Reg_Bank/n3923 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[28][31] ) );
  DFF \Reg_Bank/registers_reg[29][0]  ( .D(\Reg_Bank/n3924 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][0] ) );
  DFF \Reg_Bank/registers_reg[29][1]  ( .D(\Reg_Bank/n3925 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][1] ) );
  DFF \Reg_Bank/registers_reg[29][2]  ( .D(\Reg_Bank/n3926 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][2] ) );
  DFF \Reg_Bank/registers_reg[29][3]  ( .D(\Reg_Bank/n3927 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][3] ) );
  DFF \Reg_Bank/registers_reg[29][4]  ( .D(\Reg_Bank/n3928 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][4] ) );
  DFF \Reg_Bank/registers_reg[29][5]  ( .D(\Reg_Bank/n3929 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][5] ) );
  DFF \Reg_Bank/registers_reg[29][6]  ( .D(\Reg_Bank/n3930 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][6] ) );
  DFF \Reg_Bank/registers_reg[29][7]  ( .D(\Reg_Bank/n3931 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][7] ) );
  DFF \Reg_Bank/registers_reg[29][8]  ( .D(\Reg_Bank/n3932 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][8] ) );
  DFF \Reg_Bank/registers_reg[29][9]  ( .D(\Reg_Bank/n3933 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[29][9] ) );
  DFF \Reg_Bank/registers_reg[29][10]  ( .D(\Reg_Bank/n3934 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][10] ) );
  DFF \Reg_Bank/registers_reg[29][11]  ( .D(\Reg_Bank/n3935 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][11] ) );
  DFF \Reg_Bank/registers_reg[29][12]  ( .D(\Reg_Bank/n3936 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][12] ) );
  DFF \Reg_Bank/registers_reg[29][13]  ( .D(\Reg_Bank/n3937 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][13] ) );
  DFF \Reg_Bank/registers_reg[29][14]  ( .D(\Reg_Bank/n3938 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][14] ) );
  DFF \Reg_Bank/registers_reg[29][15]  ( .D(\Reg_Bank/n3939 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][15] ) );
  DFF \Reg_Bank/registers_reg[29][16]  ( .D(\Reg_Bank/n3940 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][16] ) );
  DFF \Reg_Bank/registers_reg[29][17]  ( .D(\Reg_Bank/n3941 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][17] ) );
  DFF \Reg_Bank/registers_reg[29][18]  ( .D(\Reg_Bank/n3942 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][18] ) );
  DFF \Reg_Bank/registers_reg[29][19]  ( .D(\Reg_Bank/n3943 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][19] ) );
  DFF \Reg_Bank/registers_reg[29][20]  ( .D(\Reg_Bank/n3944 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][20] ) );
  DFF \Reg_Bank/registers_reg[29][21]  ( .D(\Reg_Bank/n3945 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][21] ) );
  DFF \Reg_Bank/registers_reg[29][22]  ( .D(\Reg_Bank/n3946 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][22] ) );
  DFF \Reg_Bank/registers_reg[29][23]  ( .D(\Reg_Bank/n3947 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][23] ) );
  DFF \Reg_Bank/registers_reg[29][24]  ( .D(\Reg_Bank/n3948 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][24] ) );
  DFF \Reg_Bank/registers_reg[29][25]  ( .D(\Reg_Bank/n3949 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][25] ) );
  DFF \Reg_Bank/registers_reg[29][26]  ( .D(\Reg_Bank/n3950 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][26] ) );
  DFF \Reg_Bank/registers_reg[29][27]  ( .D(\Reg_Bank/n3951 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][27] ) );
  DFF \Reg_Bank/registers_reg[29][28]  ( .D(\Reg_Bank/n3952 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][28] ) );
  DFF \Reg_Bank/registers_reg[29][29]  ( .D(\Reg_Bank/n3953 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][29] ) );
  DFF \Reg_Bank/registers_reg[29][30]  ( .D(\Reg_Bank/n3954 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][30] ) );
  DFF \Reg_Bank/registers_reg[29][31]  ( .D(\Reg_Bank/n3955 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[29][31] ) );
  DFF \Reg_Bank/registers_reg[30][0]  ( .D(\Reg_Bank/n3956 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][0] ) );
  DFF \Reg_Bank/registers_reg[30][1]  ( .D(\Reg_Bank/n3957 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][1] ) );
  DFF \Reg_Bank/registers_reg[30][2]  ( .D(\Reg_Bank/n3958 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][2] ) );
  DFF \Reg_Bank/registers_reg[30][3]  ( .D(\Reg_Bank/n3959 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][3] ) );
  DFF \Reg_Bank/registers_reg[30][4]  ( .D(\Reg_Bank/n3960 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][4] ) );
  DFF \Reg_Bank/registers_reg[30][5]  ( .D(\Reg_Bank/n3961 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][5] ) );
  DFF \Reg_Bank/registers_reg[30][6]  ( .D(\Reg_Bank/n3962 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][6] ) );
  DFF \Reg_Bank/registers_reg[30][7]  ( .D(\Reg_Bank/n3963 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][7] ) );
  DFF \Reg_Bank/registers_reg[30][8]  ( .D(\Reg_Bank/n3964 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][8] ) );
  DFF \Reg_Bank/registers_reg[30][9]  ( .D(\Reg_Bank/n3965 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[30][9] ) );
  DFF \Reg_Bank/registers_reg[30][10]  ( .D(\Reg_Bank/n3966 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][10] ) );
  DFF \Reg_Bank/registers_reg[30][11]  ( .D(\Reg_Bank/n3967 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][11] ) );
  DFF \Reg_Bank/registers_reg[30][12]  ( .D(\Reg_Bank/n3968 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][12] ) );
  DFF \Reg_Bank/registers_reg[30][13]  ( .D(\Reg_Bank/n3969 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][13] ) );
  DFF \Reg_Bank/registers_reg[30][14]  ( .D(\Reg_Bank/n3970 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][14] ) );
  DFF \Reg_Bank/registers_reg[30][15]  ( .D(\Reg_Bank/n3971 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][15] ) );
  DFF \Reg_Bank/registers_reg[30][16]  ( .D(\Reg_Bank/n3972 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][16] ) );
  DFF \Reg_Bank/registers_reg[30][17]  ( .D(\Reg_Bank/n3973 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][17] ) );
  DFF \Reg_Bank/registers_reg[30][18]  ( .D(\Reg_Bank/n3974 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][18] ) );
  DFF \Reg_Bank/registers_reg[30][19]  ( .D(\Reg_Bank/n3975 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][19] ) );
  DFF \Reg_Bank/registers_reg[30][20]  ( .D(\Reg_Bank/n3976 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][20] ) );
  DFF \Reg_Bank/registers_reg[30][21]  ( .D(\Reg_Bank/n3977 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][21] ) );
  DFF \Reg_Bank/registers_reg[30][22]  ( .D(\Reg_Bank/n3978 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][22] ) );
  DFF \Reg_Bank/registers_reg[30][23]  ( .D(\Reg_Bank/n3979 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][23] ) );
  DFF \Reg_Bank/registers_reg[30][24]  ( .D(\Reg_Bank/n3980 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][24] ) );
  DFF \Reg_Bank/registers_reg[30][25]  ( .D(\Reg_Bank/n3981 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][25] ) );
  DFF \Reg_Bank/registers_reg[30][26]  ( .D(\Reg_Bank/n3982 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][26] ) );
  DFF \Reg_Bank/registers_reg[30][27]  ( .D(\Reg_Bank/n3983 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][27] ) );
  DFF \Reg_Bank/registers_reg[30][28]  ( .D(\Reg_Bank/n3984 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][28] ) );
  DFF \Reg_Bank/registers_reg[30][29]  ( .D(\Reg_Bank/n3985 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][29] ) );
  DFF \Reg_Bank/registers_reg[30][30]  ( .D(\Reg_Bank/n3986 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][30] ) );
  DFF \Reg_Bank/registers_reg[30][31]  ( .D(\Reg_Bank/n3987 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[30][31] ) );
  DFF \Reg_Bank/registers_reg[31][0]  ( .D(\Reg_Bank/n3988 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][0] ) );
  DFF \Reg_Bank/registers_reg[31][1]  ( .D(\Reg_Bank/n3989 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][1] ) );
  DFF \Reg_Bank/registers_reg[31][2]  ( .D(\Reg_Bank/n3990 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][2] ) );
  DFF \Reg_Bank/registers_reg[31][3]  ( .D(\Reg_Bank/n3991 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][3] ) );
  DFF \Reg_Bank/registers_reg[31][4]  ( .D(\Reg_Bank/n3992 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][4] ) );
  DFF \Reg_Bank/registers_reg[31][5]  ( .D(\Reg_Bank/n3993 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][5] ) );
  DFF \Reg_Bank/registers_reg[31][6]  ( .D(\Reg_Bank/n3994 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][6] ) );
  DFF \Reg_Bank/registers_reg[31][7]  ( .D(\Reg_Bank/n3995 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][7] ) );
  DFF \Reg_Bank/registers_reg[31][8]  ( .D(\Reg_Bank/n3996 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][8] ) );
  DFF \Reg_Bank/registers_reg[31][9]  ( .D(\Reg_Bank/n3997 ), .CLK(clk), .RST(
        rst), .I(1'b0), .Q(\Reg_Bank/registers[31][9] ) );
  DFF \Reg_Bank/registers_reg[31][10]  ( .D(\Reg_Bank/n3998 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][10] ) );
  DFF \Reg_Bank/registers_reg[31][11]  ( .D(\Reg_Bank/n3999 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][11] ) );
  DFF \Reg_Bank/registers_reg[31][12]  ( .D(\Reg_Bank/n4000 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][12] ) );
  DFF \Reg_Bank/registers_reg[31][13]  ( .D(\Reg_Bank/n4001 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][13] ) );
  DFF \Reg_Bank/registers_reg[31][14]  ( .D(\Reg_Bank/n4002 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][14] ) );
  DFF \Reg_Bank/registers_reg[31][15]  ( .D(\Reg_Bank/n4003 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][15] ) );
  DFF \Reg_Bank/registers_reg[31][16]  ( .D(\Reg_Bank/n4004 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][16] ) );
  DFF \Reg_Bank/registers_reg[31][17]  ( .D(\Reg_Bank/n4005 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][17] ) );
  DFF \Reg_Bank/registers_reg[31][18]  ( .D(\Reg_Bank/n4006 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][18] ) );
  DFF \Reg_Bank/registers_reg[31][19]  ( .D(\Reg_Bank/n4007 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][19] ) );
  DFF \Reg_Bank/registers_reg[31][20]  ( .D(\Reg_Bank/n4008 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][20] ) );
  DFF \Reg_Bank/registers_reg[31][21]  ( .D(\Reg_Bank/n4009 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][21] ) );
  DFF \Reg_Bank/registers_reg[31][22]  ( .D(\Reg_Bank/n4010 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][22] ) );
  DFF \Reg_Bank/registers_reg[31][23]  ( .D(\Reg_Bank/n4011 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][23] ) );
  DFF \Reg_Bank/registers_reg[31][24]  ( .D(\Reg_Bank/n4012 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][24] ) );
  DFF \Reg_Bank/registers_reg[31][25]  ( .D(\Reg_Bank/n4013 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][25] ) );
  DFF \Reg_Bank/registers_reg[31][26]  ( .D(\Reg_Bank/n4014 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][26] ) );
  DFF \Reg_Bank/registers_reg[31][27]  ( .D(\Reg_Bank/n4015 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][27] ) );
  DFF \Reg_Bank/registers_reg[31][28]  ( .D(\Reg_Bank/n4016 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][28] ) );
  DFF \Reg_Bank/registers_reg[31][29]  ( .D(\Reg_Bank/n4017 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][29] ) );
  DFF \Reg_Bank/registers_reg[31][30]  ( .D(\Reg_Bank/n4018 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][30] ) );
  DFF \Reg_Bank/registers_reg[31][31]  ( .D(\Reg_Bank/n4019 ), .CLK(clk), 
        .RST(rst), .I(1'b0), .Q(\Reg_Bank/registers[31][31] ) );
  MUX \Shifter/sll_27/M1_0_1  ( .IN0(b_bus[1]), .IN1(b_bus[0]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][1] ) );
  MUX \Shifter/sll_27/M1_0_2  ( .IN0(b_bus[2]), .IN1(b_bus[1]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][2] ) );
  MUX \Shifter/sll_27/M1_0_3  ( .IN0(b_bus[3]), .IN1(b_bus[2]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][3] ) );
  MUX \Shifter/sll_27/M1_0_4  ( .IN0(b_bus[4]), .IN1(b_bus[3]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][4] ) );
  MUX \Shifter/sll_27/M1_0_5  ( .IN0(b_bus[5]), .IN1(b_bus[4]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][5] ) );
  MUX \Shifter/sll_27/M1_0_6  ( .IN0(b_bus[6]), .IN1(b_bus[5]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][6] ) );
  MUX \Shifter/sll_27/M1_0_7  ( .IN0(b_bus[7]), .IN1(b_bus[6]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][7] ) );
  MUX \Shifter/sll_27/M1_0_8  ( .IN0(b_bus[8]), .IN1(b_bus[7]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][8] ) );
  MUX \Shifter/sll_27/M1_0_9  ( .IN0(b_bus[9]), .IN1(b_bus[8]), .SEL(a_bus[0]), 
        .F(\Shifter/sll_27/ML_int[1][9] ) );
  MUX \Shifter/sll_27/M1_0_10  ( .IN0(b_bus[10]), .IN1(b_bus[9]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][10] ) );
  MUX \Shifter/sll_27/M1_0_11  ( .IN0(b_bus[11]), .IN1(b_bus[10]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][11] ) );
  MUX \Shifter/sll_27/M1_0_12  ( .IN0(b_bus[12]), .IN1(b_bus[11]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][12] ) );
  MUX \Shifter/sll_27/M1_0_13  ( .IN0(b_bus[13]), .IN1(b_bus[12]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][13] ) );
  MUX \Shifter/sll_27/M1_0_14  ( .IN0(b_bus[14]), .IN1(b_bus[13]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][14] ) );
  MUX \Shifter/sll_27/M1_0_15  ( .IN0(b_bus[15]), .IN1(b_bus[14]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][15] ) );
  MUX \Shifter/sll_27/M1_0_16  ( .IN0(b_bus[16]), .IN1(b_bus[15]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][16] ) );
  MUX \Shifter/sll_27/M1_0_17  ( .IN0(b_bus[17]), .IN1(b_bus[16]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][17] ) );
  MUX \Shifter/sll_27/M1_0_18  ( .IN0(b_bus[18]), .IN1(b_bus[17]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][18] ) );
  MUX \Shifter/sll_27/M1_0_19  ( .IN0(b_bus[19]), .IN1(b_bus[18]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][19] ) );
  MUX \Shifter/sll_27/M1_0_20  ( .IN0(b_bus[20]), .IN1(b_bus[19]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][20] ) );
  MUX \Shifter/sll_27/M1_0_21  ( .IN0(b_bus[21]), .IN1(b_bus[20]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][21] ) );
  MUX \Shifter/sll_27/M1_0_22  ( .IN0(b_bus[22]), .IN1(b_bus[21]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][22] ) );
  MUX \Shifter/sll_27/M1_0_23  ( .IN0(b_bus[23]), .IN1(b_bus[22]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][23] ) );
  MUX \Shifter/sll_27/M1_0_24  ( .IN0(b_bus[24]), .IN1(b_bus[23]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][24] ) );
  MUX \Shifter/sll_27/M1_0_25  ( .IN0(b_bus[25]), .IN1(b_bus[24]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][25] ) );
  MUX \Shifter/sll_27/M1_0_26  ( .IN0(b_bus[26]), .IN1(b_bus[25]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][26] ) );
  MUX \Shifter/sll_27/M1_0_27  ( .IN0(b_bus[27]), .IN1(b_bus[26]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][27] ) );
  MUX \Shifter/sll_27/M1_0_28  ( .IN0(b_bus[28]), .IN1(b_bus[27]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][28] ) );
  MUX \Shifter/sll_27/M1_0_29  ( .IN0(b_bus[29]), .IN1(b_bus[28]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][29] ) );
  MUX \Shifter/sll_27/M1_0_30  ( .IN0(b_bus[30]), .IN1(b_bus[29]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][30] ) );
  MUX \Shifter/sll_27/M1_0_31  ( .IN0(\Shifter/N75 ), .IN1(b_bus[30]), .SEL(
        a_bus[0]), .F(\Shifter/sll_27/ML_int[1][31] ) );
  MUX \Shifter/sll_27/M1_1_2  ( .IN0(\Shifter/sll_27/ML_int[1][2] ), .IN1(
        \Shifter/sll_27/ML_int[1][0] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][2] ) );
  MUX \Shifter/sll_27/M1_1_3  ( .IN0(\Shifter/sll_27/ML_int[1][3] ), .IN1(
        \Shifter/sll_27/ML_int[1][1] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][3] ) );
  MUX \Shifter/sll_27/M1_1_4  ( .IN0(\Shifter/sll_27/ML_int[1][4] ), .IN1(
        \Shifter/sll_27/ML_int[1][2] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][4] ) );
  MUX \Shifter/sll_27/M1_1_5  ( .IN0(\Shifter/sll_27/ML_int[1][5] ), .IN1(
        \Shifter/sll_27/ML_int[1][3] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][5] ) );
  MUX \Shifter/sll_27/M1_1_6  ( .IN0(\Shifter/sll_27/ML_int[1][6] ), .IN1(
        \Shifter/sll_27/ML_int[1][4] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][6] ) );
  MUX \Shifter/sll_27/M1_1_7  ( .IN0(\Shifter/sll_27/ML_int[1][7] ), .IN1(
        \Shifter/sll_27/ML_int[1][5] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][7] ) );
  MUX \Shifter/sll_27/M1_1_8  ( .IN0(\Shifter/sll_27/ML_int[1][8] ), .IN1(
        \Shifter/sll_27/ML_int[1][6] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][8] ) );
  MUX \Shifter/sll_27/M1_1_9  ( .IN0(\Shifter/sll_27/ML_int[1][9] ), .IN1(
        \Shifter/sll_27/ML_int[1][7] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][9] ) );
  MUX \Shifter/sll_27/M1_1_10  ( .IN0(\Shifter/sll_27/ML_int[1][10] ), .IN1(
        \Shifter/sll_27/ML_int[1][8] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][10] ) );
  MUX \Shifter/sll_27/M1_1_11  ( .IN0(\Shifter/sll_27/ML_int[1][11] ), .IN1(
        \Shifter/sll_27/ML_int[1][9] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][11] ) );
  MUX \Shifter/sll_27/M1_1_12  ( .IN0(\Shifter/sll_27/ML_int[1][12] ), .IN1(
        \Shifter/sll_27/ML_int[1][10] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][12] ) );
  MUX \Shifter/sll_27/M1_1_13  ( .IN0(\Shifter/sll_27/ML_int[1][13] ), .IN1(
        \Shifter/sll_27/ML_int[1][11] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][13] ) );
  MUX \Shifter/sll_27/M1_1_14  ( .IN0(\Shifter/sll_27/ML_int[1][14] ), .IN1(
        \Shifter/sll_27/ML_int[1][12] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][14] ) );
  MUX \Shifter/sll_27/M1_1_15  ( .IN0(\Shifter/sll_27/ML_int[1][15] ), .IN1(
        \Shifter/sll_27/ML_int[1][13] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][15] ) );
  MUX \Shifter/sll_27/M1_1_16  ( .IN0(\Shifter/sll_27/ML_int[1][16] ), .IN1(
        \Shifter/sll_27/ML_int[1][14] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][16] ) );
  MUX \Shifter/sll_27/M1_1_17  ( .IN0(\Shifter/sll_27/ML_int[1][17] ), .IN1(
        \Shifter/sll_27/ML_int[1][15] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][17] ) );
  MUX \Shifter/sll_27/M1_1_18  ( .IN0(\Shifter/sll_27/ML_int[1][18] ), .IN1(
        \Shifter/sll_27/ML_int[1][16] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][18] ) );
  MUX \Shifter/sll_27/M1_1_19  ( .IN0(\Shifter/sll_27/ML_int[1][19] ), .IN1(
        \Shifter/sll_27/ML_int[1][17] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][19] ) );
  MUX \Shifter/sll_27/M1_1_20  ( .IN0(\Shifter/sll_27/ML_int[1][20] ), .IN1(
        \Shifter/sll_27/ML_int[1][18] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][20] ) );
  MUX \Shifter/sll_27/M1_1_21  ( .IN0(\Shifter/sll_27/ML_int[1][21] ), .IN1(
        \Shifter/sll_27/ML_int[1][19] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][21] ) );
  MUX \Shifter/sll_27/M1_1_22  ( .IN0(\Shifter/sll_27/ML_int[1][22] ), .IN1(
        \Shifter/sll_27/ML_int[1][20] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][22] ) );
  MUX \Shifter/sll_27/M1_1_23  ( .IN0(\Shifter/sll_27/ML_int[1][23] ), .IN1(
        \Shifter/sll_27/ML_int[1][21] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][23] ) );
  MUX \Shifter/sll_27/M1_1_24  ( .IN0(\Shifter/sll_27/ML_int[1][24] ), .IN1(
        \Shifter/sll_27/ML_int[1][22] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][24] ) );
  MUX \Shifter/sll_27/M1_1_25  ( .IN0(\Shifter/sll_27/ML_int[1][25] ), .IN1(
        \Shifter/sll_27/ML_int[1][23] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][25] ) );
  MUX \Shifter/sll_27/M1_1_26  ( .IN0(\Shifter/sll_27/ML_int[1][26] ), .IN1(
        \Shifter/sll_27/ML_int[1][24] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][26] ) );
  MUX \Shifter/sll_27/M1_1_27  ( .IN0(\Shifter/sll_27/ML_int[1][27] ), .IN1(
        \Shifter/sll_27/ML_int[1][25] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][27] ) );
  MUX \Shifter/sll_27/M1_1_28  ( .IN0(\Shifter/sll_27/ML_int[1][28] ), .IN1(
        \Shifter/sll_27/ML_int[1][26] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][28] ) );
  MUX \Shifter/sll_27/M1_1_29  ( .IN0(\Shifter/sll_27/ML_int[1][29] ), .IN1(
        \Shifter/sll_27/ML_int[1][27] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][29] ) );
  MUX \Shifter/sll_27/M1_1_30  ( .IN0(\Shifter/sll_27/ML_int[1][30] ), .IN1(
        \Shifter/sll_27/ML_int[1][28] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][30] ) );
  MUX \Shifter/sll_27/M1_1_31  ( .IN0(\Shifter/sll_27/ML_int[1][31] ), .IN1(
        \Shifter/sll_27/ML_int[1][29] ), .SEL(a_bus[1]), .F(
        \Shifter/sll_27/ML_int[2][31] ) );
  MUX \Shifter/sll_27/M1_2_4  ( .IN0(\Shifter/sll_27/ML_int[2][4] ), .IN1(
        \Shifter/sll_27/ML_int[2][0] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][4] ) );
  MUX \Shifter/sll_27/M1_2_5  ( .IN0(\Shifter/sll_27/ML_int[2][5] ), .IN1(
        \Shifter/sll_27/ML_int[2][1] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][5] ) );
  MUX \Shifter/sll_27/M1_2_6  ( .IN0(\Shifter/sll_27/ML_int[2][6] ), .IN1(
        \Shifter/sll_27/ML_int[2][2] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][6] ) );
  MUX \Shifter/sll_27/M1_2_7  ( .IN0(\Shifter/sll_27/ML_int[2][7] ), .IN1(
        \Shifter/sll_27/ML_int[2][3] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][7] ) );
  MUX \Shifter/sll_27/M1_2_8  ( .IN0(\Shifter/sll_27/ML_int[2][8] ), .IN1(
        \Shifter/sll_27/ML_int[2][4] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][8] ) );
  MUX \Shifter/sll_27/M1_2_9  ( .IN0(\Shifter/sll_27/ML_int[2][9] ), .IN1(
        \Shifter/sll_27/ML_int[2][5] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][9] ) );
  MUX \Shifter/sll_27/M1_2_10  ( .IN0(\Shifter/sll_27/ML_int[2][10] ), .IN1(
        \Shifter/sll_27/ML_int[2][6] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][10] ) );
  MUX \Shifter/sll_27/M1_2_11  ( .IN0(\Shifter/sll_27/ML_int[2][11] ), .IN1(
        \Shifter/sll_27/ML_int[2][7] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][11] ) );
  MUX \Shifter/sll_27/M1_2_12  ( .IN0(\Shifter/sll_27/ML_int[2][12] ), .IN1(
        \Shifter/sll_27/ML_int[2][8] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][12] ) );
  MUX \Shifter/sll_27/M1_2_13  ( .IN0(\Shifter/sll_27/ML_int[2][13] ), .IN1(
        \Shifter/sll_27/ML_int[2][9] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][13] ) );
  MUX \Shifter/sll_27/M1_2_14  ( .IN0(\Shifter/sll_27/ML_int[2][14] ), .IN1(
        \Shifter/sll_27/ML_int[2][10] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][14] ) );
  MUX \Shifter/sll_27/M1_2_15  ( .IN0(\Shifter/sll_27/ML_int[2][15] ), .IN1(
        \Shifter/sll_27/ML_int[2][11] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][15] ) );
  MUX \Shifter/sll_27/M1_2_16  ( .IN0(\Shifter/sll_27/ML_int[2][16] ), .IN1(
        \Shifter/sll_27/ML_int[2][12] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][16] ) );
  MUX \Shifter/sll_27/M1_2_17  ( .IN0(\Shifter/sll_27/ML_int[2][17] ), .IN1(
        \Shifter/sll_27/ML_int[2][13] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][17] ) );
  MUX \Shifter/sll_27/M1_2_18  ( .IN0(\Shifter/sll_27/ML_int[2][18] ), .IN1(
        \Shifter/sll_27/ML_int[2][14] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][18] ) );
  MUX \Shifter/sll_27/M1_2_19  ( .IN0(\Shifter/sll_27/ML_int[2][19] ), .IN1(
        \Shifter/sll_27/ML_int[2][15] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][19] ) );
  MUX \Shifter/sll_27/M1_2_20  ( .IN0(\Shifter/sll_27/ML_int[2][20] ), .IN1(
        \Shifter/sll_27/ML_int[2][16] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][20] ) );
  MUX \Shifter/sll_27/M1_2_21  ( .IN0(\Shifter/sll_27/ML_int[2][21] ), .IN1(
        \Shifter/sll_27/ML_int[2][17] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][21] ) );
  MUX \Shifter/sll_27/M1_2_22  ( .IN0(\Shifter/sll_27/ML_int[2][22] ), .IN1(
        \Shifter/sll_27/ML_int[2][18] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][22] ) );
  MUX \Shifter/sll_27/M1_2_23  ( .IN0(\Shifter/sll_27/ML_int[2][23] ), .IN1(
        \Shifter/sll_27/ML_int[2][19] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][23] ) );
  MUX \Shifter/sll_27/M1_2_24  ( .IN0(\Shifter/sll_27/ML_int[2][24] ), .IN1(
        \Shifter/sll_27/ML_int[2][20] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][24] ) );
  MUX \Shifter/sll_27/M1_2_25  ( .IN0(\Shifter/sll_27/ML_int[2][25] ), .IN1(
        \Shifter/sll_27/ML_int[2][21] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][25] ) );
  MUX \Shifter/sll_27/M1_2_26  ( .IN0(\Shifter/sll_27/ML_int[2][26] ), .IN1(
        \Shifter/sll_27/ML_int[2][22] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][26] ) );
  MUX \Shifter/sll_27/M1_2_27  ( .IN0(\Shifter/sll_27/ML_int[2][27] ), .IN1(
        \Shifter/sll_27/ML_int[2][23] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][27] ) );
  MUX \Shifter/sll_27/M1_2_28  ( .IN0(\Shifter/sll_27/ML_int[2][28] ), .IN1(
        \Shifter/sll_27/ML_int[2][24] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][28] ) );
  MUX \Shifter/sll_27/M1_2_29  ( .IN0(\Shifter/sll_27/ML_int[2][29] ), .IN1(
        \Shifter/sll_27/ML_int[2][25] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][29] ) );
  MUX \Shifter/sll_27/M1_2_30  ( .IN0(\Shifter/sll_27/ML_int[2][30] ), .IN1(
        \Shifter/sll_27/ML_int[2][26] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][30] ) );
  MUX \Shifter/sll_27/M1_2_31  ( .IN0(\Shifter/sll_27/ML_int[2][31] ), .IN1(
        \Shifter/sll_27/ML_int[2][27] ), .SEL(a_bus[2]), .F(
        \Shifter/sll_27/ML_int[3][31] ) );
  MUX \Shifter/sll_27/M1_3_8  ( .IN0(\Shifter/sll_27/ML_int[3][8] ), .IN1(
        \Shifter/sll_27/ML_int[3][0] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][8] ) );
  MUX \Shifter/sll_27/M1_3_9  ( .IN0(\Shifter/sll_27/ML_int[3][9] ), .IN1(
        \Shifter/sll_27/ML_int[3][1] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][9] ) );
  MUX \Shifter/sll_27/M1_3_10  ( .IN0(\Shifter/sll_27/ML_int[3][10] ), .IN1(
        \Shifter/sll_27/ML_int[3][2] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][10] ) );
  MUX \Shifter/sll_27/M1_3_11  ( .IN0(\Shifter/sll_27/ML_int[3][11] ), .IN1(
        \Shifter/sll_27/ML_int[3][3] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][11] ) );
  MUX \Shifter/sll_27/M1_3_12  ( .IN0(\Shifter/sll_27/ML_int[3][12] ), .IN1(
        \Shifter/sll_27/ML_int[3][4] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][12] ) );
  MUX \Shifter/sll_27/M1_3_13  ( .IN0(\Shifter/sll_27/ML_int[3][13] ), .IN1(
        \Shifter/sll_27/ML_int[3][5] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][13] ) );
  MUX \Shifter/sll_27/M1_3_14  ( .IN0(\Shifter/sll_27/ML_int[3][14] ), .IN1(
        \Shifter/sll_27/ML_int[3][6] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][14] ) );
  MUX \Shifter/sll_27/M1_3_15  ( .IN0(\Shifter/sll_27/ML_int[3][15] ), .IN1(
        \Shifter/sll_27/ML_int[3][7] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][15] ) );
  MUX \Shifter/sll_27/M1_3_16  ( .IN0(\Shifter/sll_27/ML_int[3][16] ), .IN1(
        \Shifter/sll_27/ML_int[3][8] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][16] ) );
  MUX \Shifter/sll_27/M1_3_17  ( .IN0(\Shifter/sll_27/ML_int[3][17] ), .IN1(
        \Shifter/sll_27/ML_int[3][9] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][17] ) );
  MUX \Shifter/sll_27/M1_3_18  ( .IN0(\Shifter/sll_27/ML_int[3][18] ), .IN1(
        \Shifter/sll_27/ML_int[3][10] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][18] ) );
  MUX \Shifter/sll_27/M1_3_19  ( .IN0(\Shifter/sll_27/ML_int[3][19] ), .IN1(
        \Shifter/sll_27/ML_int[3][11] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][19] ) );
  MUX \Shifter/sll_27/M1_3_20  ( .IN0(\Shifter/sll_27/ML_int[3][20] ), .IN1(
        \Shifter/sll_27/ML_int[3][12] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][20] ) );
  MUX \Shifter/sll_27/M1_3_21  ( .IN0(\Shifter/sll_27/ML_int[3][21] ), .IN1(
        \Shifter/sll_27/ML_int[3][13] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][21] ) );
  MUX \Shifter/sll_27/M1_3_22  ( .IN0(\Shifter/sll_27/ML_int[3][22] ), .IN1(
        \Shifter/sll_27/ML_int[3][14] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][22] ) );
  MUX \Shifter/sll_27/M1_3_23  ( .IN0(\Shifter/sll_27/ML_int[3][23] ), .IN1(
        \Shifter/sll_27/ML_int[3][15] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][23] ) );
  MUX \Shifter/sll_27/M1_3_24  ( .IN0(\Shifter/sll_27/ML_int[3][24] ), .IN1(
        \Shifter/sll_27/ML_int[3][16] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][24] ) );
  MUX \Shifter/sll_27/M1_3_25  ( .IN0(\Shifter/sll_27/ML_int[3][25] ), .IN1(
        \Shifter/sll_27/ML_int[3][17] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][25] ) );
  MUX \Shifter/sll_27/M1_3_26  ( .IN0(\Shifter/sll_27/ML_int[3][26] ), .IN1(
        \Shifter/sll_27/ML_int[3][18] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][26] ) );
  MUX \Shifter/sll_27/M1_3_27  ( .IN0(\Shifter/sll_27/ML_int[3][27] ), .IN1(
        \Shifter/sll_27/ML_int[3][19] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][27] ) );
  MUX \Shifter/sll_27/M1_3_28  ( .IN0(\Shifter/sll_27/ML_int[3][28] ), .IN1(
        \Shifter/sll_27/ML_int[3][20] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][28] ) );
  MUX \Shifter/sll_27/M1_3_29  ( .IN0(\Shifter/sll_27/ML_int[3][29] ), .IN1(
        \Shifter/sll_27/ML_int[3][21] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][29] ) );
  MUX \Shifter/sll_27/M1_3_30  ( .IN0(\Shifter/sll_27/ML_int[3][30] ), .IN1(
        \Shifter/sll_27/ML_int[3][22] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][30] ) );
  MUX \Shifter/sll_27/M1_3_31  ( .IN0(\Shifter/sll_27/ML_int[3][31] ), .IN1(
        \Shifter/sll_27/ML_int[3][23] ), .SEL(a_bus[3]), .F(
        \Shifter/sll_27/ML_int[4][31] ) );
  MUX \Shifter/sll_27/M1_4_16  ( .IN0(\Shifter/sll_27/ML_int[4][16] ), .IN1(
        \Shifter/sll_27/ML_int[4][0] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][16] ) );
  MUX \Shifter/sll_27/M1_4_17  ( .IN0(\Shifter/sll_27/ML_int[4][17] ), .IN1(
        \Shifter/sll_27/ML_int[4][1] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][17] ) );
  MUX \Shifter/sll_27/M1_4_18  ( .IN0(\Shifter/sll_27/ML_int[4][18] ), .IN1(
        \Shifter/sll_27/ML_int[4][2] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][18] ) );
  MUX \Shifter/sll_27/M1_4_19  ( .IN0(\Shifter/sll_27/ML_int[4][19] ), .IN1(
        \Shifter/sll_27/ML_int[4][3] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][19] ) );
  MUX \Shifter/sll_27/M1_4_20  ( .IN0(\Shifter/sll_27/ML_int[4][20] ), .IN1(
        \Shifter/sll_27/ML_int[4][4] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][20] ) );
  MUX \Shifter/sll_27/M1_4_21  ( .IN0(\Shifter/sll_27/ML_int[4][21] ), .IN1(
        \Shifter/sll_27/ML_int[4][5] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][21] ) );
  MUX \Shifter/sll_27/M1_4_22  ( .IN0(\Shifter/sll_27/ML_int[4][22] ), .IN1(
        \Shifter/sll_27/ML_int[4][6] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][22] ) );
  MUX \Shifter/sll_27/M1_4_23  ( .IN0(\Shifter/sll_27/ML_int[4][23] ), .IN1(
        \Shifter/sll_27/ML_int[4][7] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][23] ) );
  MUX \Shifter/sll_27/M1_4_24  ( .IN0(\Shifter/sll_27/ML_int[4][24] ), .IN1(
        \Shifter/sll_27/ML_int[4][8] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][24] ) );
  MUX \Shifter/sll_27/M1_4_25  ( .IN0(\Shifter/sll_27/ML_int[4][25] ), .IN1(
        \Shifter/sll_27/ML_int[4][9] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][25] ) );
  MUX \Shifter/sll_27/M1_4_26  ( .IN0(\Shifter/sll_27/ML_int[4][26] ), .IN1(
        \Shifter/sll_27/ML_int[4][10] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][26] ) );
  MUX \Shifter/sll_27/M1_4_27  ( .IN0(\Shifter/sll_27/ML_int[4][27] ), .IN1(
        \Shifter/sll_27/ML_int[4][11] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][27] ) );
  MUX \Shifter/sll_27/M1_4_28  ( .IN0(\Shifter/sll_27/ML_int[4][28] ), .IN1(
        \Shifter/sll_27/ML_int[4][12] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][28] ) );
  MUX \Shifter/sll_27/M1_4_29  ( .IN0(\Shifter/sll_27/ML_int[4][29] ), .IN1(
        \Shifter/sll_27/ML_int[4][13] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][29] ) );
  MUX \Shifter/sll_27/M1_4_30  ( .IN0(\Shifter/sll_27/ML_int[4][30] ), .IN1(
        \Shifter/sll_27/ML_int[4][14] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][30] ) );
  MUX \Shifter/sll_27/M1_4_31  ( .IN0(\Shifter/sll_27/ML_int[4][31] ), .IN1(
        \Shifter/sll_27/ML_int[4][15] ), .SEL(a_bus[4]), .F(
        \Shifter/sll_27/ML_int[5][31] ) );
  HADDER \PC_Next/add_32/U1_1_1  ( .IN0(pc_current[3]), .IN1(pc_current[2]), 
        .COUT(\PC_Next/add_32/carry[2] ), .SUM(pc_plus4[3]) );
  HADDER \PC_Next/add_32/U1_1_2  ( .IN0(pc_current[4]), .IN1(
        \PC_Next/add_32/carry[2] ), .COUT(\PC_Next/add_32/carry[3] ), .SUM(
        pc_plus4[4]) );
  HADDER \PC_Next/add_32/U1_1_3  ( .IN0(pc_current[5]), .IN1(
        \PC_Next/add_32/carry[3] ), .COUT(\PC_Next/add_32/carry[4] ), .SUM(
        pc_plus4[5]) );
  HADDER \PC_Next/add_32/U1_1_4  ( .IN0(pc_current[6]), .IN1(
        \PC_Next/add_32/carry[4] ), .COUT(\PC_Next/add_32/carry[5] ), .SUM(
        pc_plus4[6]) );
  HADDER \PC_Next/add_32/U1_1_5  ( .IN0(pc_current[7]), .IN1(
        \PC_Next/add_32/carry[5] ), .COUT(\PC_Next/add_32/carry[6] ), .SUM(
        pc_plus4[7]) );
  HADDER \PC_Next/add_32/U1_1_6  ( .IN0(pc_current[8]), .IN1(
        \PC_Next/add_32/carry[6] ), .COUT(\PC_Next/add_32/carry[7] ), .SUM(
        pc_plus4[8]) );
  HADDER \PC_Next/add_32/U1_1_7  ( .IN0(pc_current[9]), .IN1(
        \PC_Next/add_32/carry[7] ), .COUT(\PC_Next/add_32/carry[8] ), .SUM(
        pc_plus4[9]) );
  HADDER \PC_Next/add_32/U1_1_8  ( .IN0(pc_current[10]), .IN1(
        \PC_Next/add_32/carry[8] ), .COUT(\PC_Next/add_32/carry[9] ), .SUM(
        pc_plus4[10]) );
  HADDER \PC_Next/add_32/U1_1_9  ( .IN0(pc_current[11]), .IN1(
        \PC_Next/add_32/carry[9] ), .COUT(\PC_Next/add_32/carry[10] ), .SUM(
        pc_plus4[11]) );
  HADDER \PC_Next/add_32/U1_1_10  ( .IN0(pc_current[12]), .IN1(
        \PC_Next/add_32/carry[10] ), .COUT(\PC_Next/add_32/carry[11] ), .SUM(
        pc_plus4[12]) );
  HADDER \PC_Next/add_32/U1_1_11  ( .IN0(pc_current[13]), .IN1(
        \PC_Next/add_32/carry[11] ), .COUT(\PC_Next/add_32/carry[12] ), .SUM(
        pc_plus4[13]) );
  HADDER \PC_Next/add_32/U1_1_12  ( .IN0(pc_current[14]), .IN1(
        \PC_Next/add_32/carry[12] ), .COUT(\PC_Next/add_32/carry[13] ), .SUM(
        pc_plus4[14]) );
  HADDER \PC_Next/add_32/U1_1_13  ( .IN0(pc_current[15]), .IN1(
        \PC_Next/add_32/carry[13] ), .COUT(\PC_Next/add_32/carry[14] ), .SUM(
        pc_plus4[15]) );
  HADDER \PC_Next/add_32/U1_1_14  ( .IN0(pc_current[16]), .IN1(
        \PC_Next/add_32/carry[14] ), .COUT(\PC_Next/add_32/carry[15] ), .SUM(
        pc_plus4[16]) );
  HADDER \PC_Next/add_32/U1_1_15  ( .IN0(pc_current[17]), .IN1(
        \PC_Next/add_32/carry[15] ), .COUT(\PC_Next/add_32/carry[16] ), .SUM(
        pc_plus4[17]) );
  HADDER \PC_Next/add_32/U1_1_16  ( .IN0(pc_current[18]), .IN1(
        \PC_Next/add_32/carry[16] ), .COUT(\PC_Next/add_32/carry[17] ), .SUM(
        pc_plus4[18]) );
  HADDER \PC_Next/add_32/U1_1_17  ( .IN0(pc_current[19]), .IN1(
        \PC_Next/add_32/carry[17] ), .COUT(\PC_Next/add_32/carry[18] ), .SUM(
        pc_plus4[19]) );
  HADDER \PC_Next/add_32/U1_1_18  ( .IN0(pc_current[20]), .IN1(
        \PC_Next/add_32/carry[18] ), .COUT(\PC_Next/add_32/carry[19] ), .SUM(
        pc_plus4[20]) );
  HADDER \PC_Next/add_32/U1_1_19  ( .IN0(pc_current[21]), .IN1(
        \PC_Next/add_32/carry[19] ), .COUT(\PC_Next/add_32/carry[20] ), .SUM(
        pc_plus4[21]) );
  HADDER \PC_Next/add_32/U1_1_20  ( .IN0(pc_current[22]), .IN1(
        \PC_Next/add_32/carry[20] ), .COUT(\PC_Next/add_32/carry[21] ), .SUM(
        pc_plus4[22]) );
  HADDER \PC_Next/add_32/U1_1_21  ( .IN0(pc_current[23]), .IN1(
        \PC_Next/add_32/carry[21] ), .COUT(\PC_Next/add_32/carry[22] ), .SUM(
        pc_plus4[23]) );
  HADDER \PC_Next/add_32/U1_1_22  ( .IN0(pc_current[24]), .IN1(
        \PC_Next/add_32/carry[22] ), .COUT(\PC_Next/add_32/carry[23] ), .SUM(
        pc_plus4[24]) );
  HADDER \PC_Next/add_32/U1_1_23  ( .IN0(pc_current[25]), .IN1(
        \PC_Next/add_32/carry[23] ), .COUT(\PC_Next/add_32/carry[24] ), .SUM(
        pc_plus4[25]) );
  HADDER \PC_Next/add_32/U1_1_24  ( .IN0(pc_current[26]), .IN1(
        \PC_Next/add_32/carry[24] ), .COUT(\PC_Next/add_32/carry[25] ), .SUM(
        pc_plus4[26]) );
  HADDER \PC_Next/add_32/U1_1_25  ( .IN0(pc_current[27]), .IN1(
        \PC_Next/add_32/carry[25] ), .COUT(\PC_Next/add_32/carry[26] ), .SUM(
        pc_plus4[27]) );
  HADDER \PC_Next/add_32/U1_1_26  ( .IN0(pc_current[28]), .IN1(
        \PC_Next/add_32/carry[26] ), .COUT(\PC_Next/add_32/carry[27] ), .SUM(
        pc_plus4[28]) );
  HADDER \PC_Next/add_32/U1_1_27  ( .IN0(pc_current[29]), .IN1(
        \PC_Next/add_32/carry[27] ), .COUT(\PC_Next/add_32/carry[28] ), .SUM(
        pc_plus4[29]) );
  HADDER \PC_Next/add_32/U1_1_28  ( .IN0(pc_current[30]), .IN1(
        \PC_Next/add_32/carry[28] ), .COUT(\PC_Next/add_32/carry[29] ), .SUM(
        pc_plus4[30]) );
  FADDER \PC_Next/add_48/U1_1  ( .CIN(pc_current[3]), .IN0(imm[1]), .IN1(
        \PC_Next/add_48/carry[1] ), .COUT(\PC_Next/add_48/carry[2] ), .SUM(
        \PC_Next/pc_jump[3] ) );
  FADDER \PC_Next/add_48/U1_2  ( .CIN(pc_current[4]), .IN0(imm[2]), .IN1(
        \PC_Next/add_48/carry[2] ), .COUT(\PC_Next/add_48/carry[3] ), .SUM(
        \PC_Next/pc_jump[4] ) );
  FADDER \PC_Next/add_48/U1_3  ( .CIN(pc_current[5]), .IN0(imm[3]), .IN1(
        \PC_Next/add_48/carry[3] ), .COUT(\PC_Next/add_48/carry[4] ), .SUM(
        \PC_Next/pc_jump[5] ) );
  FADDER \PC_Next/add_48/U1_4  ( .CIN(pc_current[6]), .IN0(imm[4]), .IN1(
        \PC_Next/add_48/carry[4] ), .COUT(\PC_Next/add_48/carry[5] ), .SUM(
        \PC_Next/pc_jump[6] ) );
  FADDER \PC_Next/add_48/U1_5  ( .CIN(pc_current[7]), .IN0(imm[5]), .IN1(
        \PC_Next/add_48/carry[5] ), .COUT(\PC_Next/add_48/carry[6] ), .SUM(
        \PC_Next/pc_jump[7] ) );
  FADDER \PC_Next/add_48/U1_6  ( .CIN(pc_current[8]), .IN0(imm[6]), .IN1(
        \PC_Next/add_48/carry[6] ), .COUT(\PC_Next/add_48/carry[7] ), .SUM(
        \PC_Next/pc_jump[8] ) );
  FADDER \PC_Next/add_48/U1_7  ( .CIN(pc_current[9]), .IN0(imm[7]), .IN1(
        \PC_Next/add_48/carry[7] ), .COUT(\PC_Next/add_48/carry[8] ), .SUM(
        \PC_Next/pc_jump[9] ) );
  FADDER \PC_Next/add_48/U1_8  ( .CIN(pc_current[10]), .IN0(imm[8]), .IN1(
        \PC_Next/add_48/carry[8] ), .COUT(\PC_Next/add_48/carry[9] ), .SUM(
        \PC_Next/pc_jump[10] ) );
  FADDER \PC_Next/add_48/U1_9  ( .CIN(pc_current[11]), .IN0(imm[9]), .IN1(
        \PC_Next/add_48/carry[9] ), .COUT(\PC_Next/add_48/carry[10] ), .SUM(
        \PC_Next/pc_jump[11] ) );
  FADDER \PC_Next/add_48/U1_10  ( .CIN(pc_current[12]), .IN0(imm[10]), .IN1(
        \PC_Next/add_48/carry[10] ), .COUT(\PC_Next/add_48/carry[11] ), .SUM(
        \PC_Next/pc_jump[12] ) );
  FADDER \PC_Next/add_48/U1_11  ( .CIN(pc_current[13]), .IN0(imm[11]), .IN1(
        \PC_Next/add_48/carry[11] ), .COUT(\PC_Next/add_48/carry[12] ), .SUM(
        \PC_Next/pc_jump[13] ) );
  FADDER \PC_Next/add_48/U1_12  ( .CIN(pc_current[14]), .IN0(imm[12]), .IN1(
        \PC_Next/add_48/carry[12] ), .COUT(\PC_Next/add_48/carry[13] ), .SUM(
        \PC_Next/pc_jump[14] ) );
  FADDER \PC_Next/add_48/U1_13  ( .CIN(pc_current[15]), .IN0(imm[13]), .IN1(
        \PC_Next/add_48/carry[13] ), .COUT(\PC_Next/add_48/carry[14] ), .SUM(
        \PC_Next/pc_jump[15] ) );
  FADDER \PC_Next/add_48/U1_14  ( .CIN(pc_current[16]), .IN0(imm[14]), .IN1(
        \PC_Next/add_48/carry[14] ), .COUT(\PC_Next/add_48/carry[15] ), .SUM(
        \PC_Next/pc_jump[16] ) );
  FADDER \PC_Next/add_48/U1_15  ( .CIN(pc_current[17]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[15] ), .COUT(\PC_Next/add_48/carry[16] ), .SUM(
        \PC_Next/pc_jump[17] ) );
  FADDER \PC_Next/add_48/U1_16  ( .CIN(pc_current[18]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[16] ), .COUT(\PC_Next/add_48/carry[17] ), .SUM(
        \PC_Next/pc_jump[18] ) );
  FADDER \PC_Next/add_48/U1_17  ( .CIN(pc_current[19]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[17] ), .COUT(\PC_Next/add_48/carry[18] ), .SUM(
        \PC_Next/pc_jump[19] ) );
  FADDER \PC_Next/add_48/U1_18  ( .CIN(pc_current[20]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[18] ), .COUT(\PC_Next/add_48/carry[19] ), .SUM(
        \PC_Next/pc_jump[20] ) );
  FADDER \PC_Next/add_48/U1_19  ( .CIN(pc_current[21]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[19] ), .COUT(\PC_Next/add_48/carry[20] ), .SUM(
        \PC_Next/pc_jump[21] ) );
  FADDER \PC_Next/add_48/U1_20  ( .CIN(pc_current[22]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[20] ), .COUT(\PC_Next/add_48/carry[21] ), .SUM(
        \PC_Next/pc_jump[22] ) );
  FADDER \PC_Next/add_48/U1_21  ( .CIN(pc_current[23]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[21] ), .COUT(\PC_Next/add_48/carry[22] ), .SUM(
        \PC_Next/pc_jump[23] ) );
  FADDER \PC_Next/add_48/U1_22  ( .CIN(pc_current[24]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[22] ), .COUT(\PC_Next/add_48/carry[23] ), .SUM(
        \PC_Next/pc_jump[24] ) );
  FADDER \PC_Next/add_48/U1_23  ( .CIN(pc_current[25]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[23] ), .COUT(\PC_Next/add_48/carry[24] ), .SUM(
        \PC_Next/pc_jump[25] ) );
  FADDER \PC_Next/add_48/U1_24  ( .CIN(pc_current[26]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[24] ), .COUT(\PC_Next/add_48/carry[25] ), .SUM(
        \PC_Next/pc_jump[26] ) );
  FADDER \PC_Next/add_48/U1_25  ( .CIN(pc_current[27]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[25] ), .COUT(\PC_Next/add_48/carry[26] ), .SUM(
        \PC_Next/pc_jump[27] ) );
  FADDER \PC_Next/add_48/U1_26  ( .CIN(pc_current[28]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[26] ), .COUT(\PC_Next/add_48/carry[27] ), .SUM(
        \PC_Next/pc_jump[28] ) );
  FADDER \PC_Next/add_48/U1_27  ( .CIN(pc_current[29]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[27] ), .COUT(\PC_Next/add_48/carry[28] ), .SUM(
        \PC_Next/pc_jump[29] ) );
  FADDER \PC_Next/add_48/U1_28  ( .CIN(pc_current[30]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[28] ), .COUT(\PC_Next/add_48/carry[29] ), .SUM(
        \PC_Next/pc_jump[30] ) );
  FADDER \PC_Next/add_48/U1_29  ( .CIN(pc_current[31]), .IN0(imm[15]), .IN1(
        \PC_Next/add_48/carry[29] ), .SUM(\PC_Next/pc_jump[31] ) );
  AND U34 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][31] ), .Z(
        \Reg_Bank/n5936 ) );
  AND U35 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][31] ), .Z(
        \Reg_Bank/n4976 ) );
  AND U36 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][30] ), .Z(
        \Reg_Bank/n5906 ) );
  AND U37 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][30] ), .Z(
        \Reg_Bank/n4946 ) );
  AND U38 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][29] ), .Z(
        \Reg_Bank/n5876 ) );
  AND U39 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][29] ), .Z(
        \Reg_Bank/n4916 ) );
  AND U40 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][28] ), .Z(
        \Reg_Bank/n5846 ) );
  AND U41 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][28] ), .Z(
        \Reg_Bank/n4886 ) );
  AND U42 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][27] ), .Z(
        \Reg_Bank/n5816 ) );
  AND U43 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][27] ), .Z(
        \Reg_Bank/n4856 ) );
  AND U44 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][26] ), .Z(
        \Reg_Bank/n5786 ) );
  AND U45 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][26] ), .Z(
        \Reg_Bank/n4826 ) );
  AND U46 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][25] ), .Z(
        \Reg_Bank/n5756 ) );
  AND U47 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][25] ), .Z(
        \Reg_Bank/n4796 ) );
  AND U48 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][24] ), .Z(
        \Reg_Bank/n5726 ) );
  AND U49 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][24] ), .Z(
        \Reg_Bank/n4766 ) );
  AND U50 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][23] ), .Z(
        \Reg_Bank/n5696 ) );
  AND U51 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][23] ), .Z(
        \Reg_Bank/n4736 ) );
  AND U52 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][22] ), .Z(
        \Reg_Bank/n5666 ) );
  AND U53 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][22] ), .Z(
        \Reg_Bank/n4706 ) );
  AND U54 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][21] ), .Z(
        \Reg_Bank/n5636 ) );
  AND U55 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][21] ), .Z(
        \Reg_Bank/n4676 ) );
  AND U56 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][20] ), .Z(
        \Reg_Bank/n5606 ) );
  AND U57 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][20] ), .Z(
        \Reg_Bank/n4646 ) );
  AND U58 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][19] ), .Z(
        \Reg_Bank/n5576 ) );
  AND U59 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][19] ), .Z(
        \Reg_Bank/n4616 ) );
  AND U60 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][18] ), .Z(
        \Reg_Bank/n5546 ) );
  AND U61 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][18] ), .Z(
        \Reg_Bank/n4586 ) );
  AND U62 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][17] ), .Z(
        \Reg_Bank/n5516 ) );
  AND U63 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][17] ), .Z(
        \Reg_Bank/n4556 ) );
  AND U64 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][16] ), .Z(
        \Reg_Bank/n5486 ) );
  AND U65 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][16] ), .Z(
        \Reg_Bank/n4526 ) );
  AND U66 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][15] ), .Z(
        \Reg_Bank/n5456 ) );
  AND U67 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][15] ), .Z(
        \Reg_Bank/n4496 ) );
  AND U68 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][14] ), .Z(
        \Reg_Bank/n5426 ) );
  AND U69 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][14] ), .Z(
        \Reg_Bank/n4466 ) );
  AND U70 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][13] ), .Z(
        \Reg_Bank/n5396 ) );
  AND U71 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][13] ), .Z(
        \Reg_Bank/n4436 ) );
  AND U72 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][12] ), .Z(
        \Reg_Bank/n5366 ) );
  AND U73 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][12] ), .Z(
        \Reg_Bank/n4406 ) );
  AND U74 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][11] ), .Z(
        \Reg_Bank/n5336 ) );
  AND U75 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][11] ), .Z(
        \Reg_Bank/n4376 ) );
  AND U76 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][10] ), .Z(
        \Reg_Bank/n5306 ) );
  AND U77 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][10] ), .Z(
        \Reg_Bank/n4346 ) );
  AND U78 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][9] ), .Z(
        \Reg_Bank/n5276 ) );
  AND U79 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][9] ), .Z(
        \Reg_Bank/n4316 ) );
  AND U80 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][8] ), .Z(
        \Reg_Bank/n5246 ) );
  AND U81 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][8] ), .Z(
        \Reg_Bank/n4286 ) );
  AND U82 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][7] ), .Z(
        \Reg_Bank/n5216 ) );
  AND U83 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][7] ), .Z(
        \Reg_Bank/n4256 ) );
  AND U84 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][6] ), .Z(
        \Reg_Bank/n5186 ) );
  AND U85 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][6] ), .Z(
        \Reg_Bank/n4226 ) );
  AND U86 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][5] ), .Z(
        \Reg_Bank/n5156 ) );
  AND U87 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][5] ), .Z(
        \Reg_Bank/n4196 ) );
  AND U88 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][4] ), .Z(
        \Reg_Bank/n5126 ) );
  AND U89 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][4] ), .Z(
        \Reg_Bank/n4166 ) );
  AND U90 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][3] ), .Z(
        \Reg_Bank/n5096 ) );
  AND U91 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][3] ), .Z(
        \Reg_Bank/n4136 ) );
  AND U92 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][2] ), .Z(
        \Reg_Bank/n5066 ) );
  AND U93 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][2] ), .Z(
        \Reg_Bank/n4106 ) );
  AND U94 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][1] ), .Z(
        \Reg_Bank/n5036 ) );
  AND U95 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][1] ), .Z(
        \Reg_Bank/n4076 ) );
  AND U96 ( .A(rt_index[0]), .B(\Reg_Bank/registers[1][0] ), .Z(
        \Reg_Bank/n5006 ) );
  AND U97 ( .A(rs_index[0]), .B(\Reg_Bank/registers[1][0] ), .Z(
        \Reg_Bank/n4046 ) );
  AND U98 ( .A(pc_current[2]), .B(imm[0]), .Z(\PC_Next/add_48/carry[1] ) );
  XOR U99 ( .A(imm[0]), .B(pc_current[2]), .Z(\PC_Next/pc_jump[2] ) );
  NAND U100 ( .A(n1), .B(n2), .Z(rt_index[4]) );
  NAND U101 ( .A(n3), .B(opcode[20]), .Z(n2) );
  AND U102 ( .A(n4), .B(n5), .Z(n1) );
  NANDN U103 ( .B(n6), .A(n7), .Z(n5) );
  NAND U104 ( .A(n8), .B(n9), .Z(n7) );
  NANDN U105 ( .B(n10), .A(n11), .Z(n9) );
  NAND U106 ( .A(n12), .B(n13), .Z(n11) );
  NANDN U107 ( .B(n14), .A(opcode[20]), .Z(n13) );
  NANDN U108 ( .B(n15), .A(opcode[20]), .Z(n12) );
  AND U109 ( .A(n16), .B(n17), .Z(n8) );
  NANDN U110 ( .B(n18), .A(n19), .Z(n17) );
  NAND U111 ( .A(n20), .B(n21), .Z(n19) );
  NANDN U112 ( .B(n22), .A(opcode[20]), .Z(n21) );
  NANDN U113 ( .B(n23), .A(opcode[20]), .Z(n20) );
  NAND U114 ( .A(n24), .B(opcode[20]), .Z(n16) );
  NAND U115 ( .A(n25), .B(n26), .Z(n4) );
  NAND U116 ( .A(n27), .B(n28), .Z(n25) );
  NAND U117 ( .A(n29), .B(opcode[20]), .Z(n28) );
  NAND U118 ( .A(n30), .B(opcode[20]), .Z(n27) );
  NAND U119 ( .A(n31), .B(n32), .Z(rt_index[3]) );
  NANDN U120 ( .B(n23), .A(n3), .Z(n32) );
  AND U121 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U122 ( .B(n6), .A(n35), .Z(n34) );
  NAND U123 ( .A(n36), .B(n37), .Z(n35) );
  NANDN U124 ( .B(n10), .A(n38), .Z(n37) );
  NAND U125 ( .A(n39), .B(n40), .Z(n38) );
  NANDN U126 ( .B(n23), .A(imm[1]), .Z(n40) );
  NANDN U127 ( .B(n15), .A(opcode[19]), .Z(n39) );
  AND U128 ( .A(n41), .B(n42), .Z(n36) );
  NANDN U129 ( .B(n23), .A(n43), .Z(n42) );
  NANDN U130 ( .B(n23), .A(n24), .Z(n41) );
  NAND U131 ( .A(n44), .B(n26), .Z(n33) );
  NAND U132 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U133 ( .B(n23), .A(n29), .Z(n46) );
  NANDN U134 ( .B(n23), .A(n30), .Z(n45) );
  NAND U135 ( .A(n47), .B(n48), .Z(rt_index[2]) );
  NANDN U136 ( .B(n49), .A(n3), .Z(n48) );
  AND U137 ( .A(n50), .B(n51), .Z(n47) );
  NANDN U138 ( .B(n6), .A(n52), .Z(n51) );
  NAND U139 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U140 ( .B(n10), .A(n55), .Z(n54) );
  NAND U141 ( .A(n56), .B(n57), .Z(n55) );
  NANDN U142 ( .B(n14), .A(opcode[18]), .Z(n57) );
  NANDN U143 ( .B(n15), .A(opcode[18]), .Z(n56) );
  AND U144 ( .A(n58), .B(n59), .Z(n53) );
  NANDN U145 ( .B(n18), .A(opcode[18]), .Z(n59) );
  NANDN U146 ( .B(n49), .A(n24), .Z(n58) );
  NAND U147 ( .A(n60), .B(n26), .Z(n50) );
  NAND U148 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U149 ( .B(n49), .A(n29), .Z(n62) );
  NANDN U150 ( .B(n49), .A(n30), .Z(n61) );
  NAND U151 ( .A(n63), .B(n64), .Z(rt_index[1]) );
  NANDN U152 ( .B(n65), .A(n3), .Z(n64) );
  AND U153 ( .A(n66), .B(n67), .Z(n63) );
  NANDN U154 ( .B(n6), .A(n68), .Z(n67) );
  NAND U155 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U156 ( .B(n10), .A(n71), .Z(n70) );
  NAND U157 ( .A(n72), .B(n73), .Z(n71) );
  NANDN U158 ( .B(n14), .A(opcode[17]), .Z(n73) );
  NANDN U159 ( .B(n15), .A(opcode[17]), .Z(n72) );
  AND U160 ( .A(n74), .B(n75), .Z(n69) );
  NANDN U161 ( .B(n18), .A(opcode[17]), .Z(n75) );
  NANDN U162 ( .B(n65), .A(n24), .Z(n74) );
  NAND U163 ( .A(n76), .B(n26), .Z(n66) );
  NAND U164 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U165 ( .B(n65), .A(n29), .Z(n78) );
  NANDN U166 ( .B(n65), .A(n30), .Z(n77) );
  NAND U167 ( .A(n79), .B(n80), .Z(rt_index[0]) );
  NANDN U168 ( .B(n81), .A(n3), .Z(n80) );
  AND U169 ( .A(n82), .B(n83), .Z(n79) );
  NANDN U170 ( .B(n6), .A(n84), .Z(n83) );
  NAND U171 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U172 ( .B(n10), .A(n87), .Z(n86) );
  NAND U173 ( .A(n88), .B(n89), .Z(n87) );
  NANDN U174 ( .B(n14), .A(opcode[16]), .Z(n89) );
  NANDN U175 ( .B(n15), .A(opcode[16]), .Z(n88) );
  AND U176 ( .A(n90), .B(n91), .Z(n85) );
  NANDN U177 ( .B(n18), .A(n92), .Z(n91) );
  NAND U178 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U179 ( .B(n22), .A(opcode[16]), .Z(n94) );
  NANDN U180 ( .B(n23), .A(opcode[16]), .Z(n93) );
  NANDN U181 ( .B(n81), .A(n24), .Z(n90) );
  NAND U182 ( .A(n95), .B(n96), .Z(n24) );
  NAND U183 ( .A(n97), .B(n26), .Z(n82) );
  NAND U184 ( .A(n98), .B(n99), .Z(n97) );
  NANDN U185 ( .B(n81), .A(n29), .Z(n99) );
  NANDN U186 ( .B(n81), .A(n30), .Z(n98) );
  NAND U187 ( .A(n100), .B(n101), .Z(rs_index[4]) );
  ANDN U188 ( .A(n102), .B(opcode[25]), .Z(n100) );
  NAND U189 ( .A(n103), .B(n104), .Z(n102) );
  MUX U190 ( .IN0(imm[15]), .IN1(opcode[20]), .SEL(opcode[23]), .F(n104) );
  NAND U191 ( .A(n105), .B(n106), .Z(rs_index[3]) );
  NAND U192 ( .A(n103), .B(n107), .Z(n106) );
  MUX U193 ( .IN0(imm[14]), .IN1(opcode[19]), .SEL(opcode[23]), .F(n107) );
  ANDN U194 ( .A(n101), .B(opcode[24]), .Z(n105) );
  NAND U195 ( .A(n108), .B(n109), .Z(rs_index[2]) );
  NANDN U196 ( .B(n6), .A(n110), .Z(n109) );
  NANDN U197 ( .B(opcode[23]), .A(n111), .Z(n110) );
  NAND U198 ( .A(n112), .B(n113), .Z(n111) );
  ANDN U199 ( .A(n114), .B(n10), .Z(n112) );
  AND U200 ( .A(n115), .B(n116), .Z(n108) );
  NAND U201 ( .A(n117), .B(n26), .Z(n116) );
  NAND U202 ( .A(n118), .B(n119), .Z(n117) );
  NANDN U203 ( .B(n10), .A(n120), .Z(n119) );
  NAND U204 ( .A(n121), .B(n122), .Z(n120) );
  NAND U205 ( .A(n123), .B(n124), .Z(n122) );
  MUX U206 ( .IN0(imm[13]), .IN1(opcode[18]), .SEL(opcode[23]), .F(n123) );
  NANDN U207 ( .B(n125), .A(n29), .Z(n121) );
  NANDN U208 ( .B(n126), .A(n127), .Z(n29) );
  NANDN U209 ( .B(n125), .A(n30), .Z(n118) );
  NAND U210 ( .A(n128), .B(n129), .Z(n30) );
  ANDN U211 ( .A(n18), .B(n130), .Z(n129) );
  NANDN U212 ( .B(n125), .A(n3), .Z(n115) );
  NAND U213 ( .A(n131), .B(n132), .Z(n3) );
  ANDN U214 ( .A(n133), .B(n134), .Z(n131) );
  NAND U215 ( .A(n135), .B(n136), .Z(rs_index[1]) );
  NAND U216 ( .A(n103), .B(n137), .Z(n136) );
  MUX U217 ( .IN0(imm[12]), .IN1(opcode[17]), .SEL(opcode[23]), .F(n137) );
  ANDN U218 ( .A(n101), .B(opcode[22]), .Z(n135) );
  NAND U219 ( .A(n138), .B(n139), .Z(rs_index[0]) );
  NAND U220 ( .A(n103), .B(n140), .Z(n139) );
  MUX U221 ( .IN0(imm[11]), .IN1(opcode[16]), .SEL(opcode[23]), .F(n140) );
  ANDN U222 ( .A(n101), .B(opcode[21]), .Z(n138) );
  NAND U223 ( .A(n141), .B(n142), .Z(n101) );
  ANDN U224 ( .A(n143), .B(n6), .Z(n142) );
  AND U225 ( .A(n114), .B(n113), .Z(n141) );
  MUX U226 ( .IN0(\Reg_Bank/registers[31][31] ), .IN1(n144), .SEL(n145), .F(
        \Reg_Bank/n4019 ) );
  MUX U227 ( .IN0(\Reg_Bank/registers[31][30] ), .IN1(n146), .SEL(n145), .F(
        \Reg_Bank/n4018 ) );
  MUX U228 ( .IN0(\Reg_Bank/registers[31][29] ), .IN1(n147), .SEL(n145), .F(
        \Reg_Bank/n4017 ) );
  MUX U229 ( .IN0(\Reg_Bank/registers[31][28] ), .IN1(n148), .SEL(n145), .F(
        \Reg_Bank/n4016 ) );
  MUX U230 ( .IN0(\Reg_Bank/registers[31][27] ), .IN1(n149), .SEL(n145), .F(
        \Reg_Bank/n4015 ) );
  MUX U231 ( .IN0(\Reg_Bank/registers[31][26] ), .IN1(n150), .SEL(n145), .F(
        \Reg_Bank/n4014 ) );
  MUX U232 ( .IN0(\Reg_Bank/registers[31][25] ), .IN1(n151), .SEL(n145), .F(
        \Reg_Bank/n4013 ) );
  MUX U233 ( .IN0(\Reg_Bank/registers[31][24] ), .IN1(n152), .SEL(n145), .F(
        \Reg_Bank/n4012 ) );
  MUX U234 ( .IN0(\Reg_Bank/registers[31][23] ), .IN1(n153), .SEL(n145), .F(
        \Reg_Bank/n4011 ) );
  MUX U235 ( .IN0(\Reg_Bank/registers[31][22] ), .IN1(n154), .SEL(n145), .F(
        \Reg_Bank/n4010 ) );
  MUX U236 ( .IN0(\Reg_Bank/registers[31][21] ), .IN1(n155), .SEL(n145), .F(
        \Reg_Bank/n4009 ) );
  MUX U237 ( .IN0(\Reg_Bank/registers[31][20] ), .IN1(n156), .SEL(n145), .F(
        \Reg_Bank/n4008 ) );
  MUX U238 ( .IN0(\Reg_Bank/registers[31][19] ), .IN1(n157), .SEL(n145), .F(
        \Reg_Bank/n4007 ) );
  MUX U239 ( .IN0(\Reg_Bank/registers[31][18] ), .IN1(n158), .SEL(n145), .F(
        \Reg_Bank/n4006 ) );
  MUX U240 ( .IN0(\Reg_Bank/registers[31][17] ), .IN1(n159), .SEL(n145), .F(
        \Reg_Bank/n4005 ) );
  MUX U241 ( .IN0(\Reg_Bank/registers[31][16] ), .IN1(n160), .SEL(n145), .F(
        \Reg_Bank/n4004 ) );
  MUX U242 ( .IN0(\Reg_Bank/registers[31][15] ), .IN1(n161), .SEL(n145), .F(
        \Reg_Bank/n4003 ) );
  MUX U243 ( .IN0(\Reg_Bank/registers[31][14] ), .IN1(n162), .SEL(n145), .F(
        \Reg_Bank/n4002 ) );
  MUX U244 ( .IN0(\Reg_Bank/registers[31][13] ), .IN1(n163), .SEL(n145), .F(
        \Reg_Bank/n4001 ) );
  MUX U245 ( .IN0(\Reg_Bank/registers[31][12] ), .IN1(n164), .SEL(n145), .F(
        \Reg_Bank/n4000 ) );
  MUX U246 ( .IN0(\Reg_Bank/registers[31][11] ), .IN1(n165), .SEL(n145), .F(
        \Reg_Bank/n3999 ) );
  MUX U247 ( .IN0(\Reg_Bank/registers[31][10] ), .IN1(n166), .SEL(n145), .F(
        \Reg_Bank/n3998 ) );
  MUX U248 ( .IN0(\Reg_Bank/registers[31][9] ), .IN1(n167), .SEL(n145), .F(
        \Reg_Bank/n3997 ) );
  MUX U249 ( .IN0(\Reg_Bank/registers[31][8] ), .IN1(n168), .SEL(n145), .F(
        \Reg_Bank/n3996 ) );
  MUX U250 ( .IN0(\Reg_Bank/registers[31][7] ), .IN1(n169), .SEL(n145), .F(
        \Reg_Bank/n3995 ) );
  MUX U251 ( .IN0(\Reg_Bank/registers[31][6] ), .IN1(n170), .SEL(n145), .F(
        \Reg_Bank/n3994 ) );
  MUX U252 ( .IN0(\Reg_Bank/registers[31][5] ), .IN1(n171), .SEL(n145), .F(
        \Reg_Bank/n3993 ) );
  MUX U253 ( .IN0(\Reg_Bank/registers[31][4] ), .IN1(n172), .SEL(n145), .F(
        \Reg_Bank/n3992 ) );
  MUX U254 ( .IN0(\Reg_Bank/registers[31][3] ), .IN1(n173), .SEL(n145), .F(
        \Reg_Bank/n3991 ) );
  MUX U255 ( .IN0(\Reg_Bank/registers[31][2] ), .IN1(n174), .SEL(n145), .F(
        \Reg_Bank/n3990 ) );
  IV U256 ( .A(n175), .Z(n145) );
  MUX U257 ( .IN0(n176), .IN1(\Reg_Bank/registers[31][1] ), .SEL(n175), .F(
        \Reg_Bank/n3989 ) );
  MUX U258 ( .IN0(n177), .IN1(\Reg_Bank/registers[31][0] ), .SEL(n175), .F(
        \Reg_Bank/n3988 ) );
  NANDN U259 ( .B(n178), .A(n179), .Z(n175) );
  MUX U260 ( .IN0(\Reg_Bank/registers[30][31] ), .IN1(n144), .SEL(n180), .F(
        \Reg_Bank/n3987 ) );
  MUX U261 ( .IN0(\Reg_Bank/registers[30][30] ), .IN1(n146), .SEL(n180), .F(
        \Reg_Bank/n3986 ) );
  MUX U262 ( .IN0(\Reg_Bank/registers[30][29] ), .IN1(n147), .SEL(n180), .F(
        \Reg_Bank/n3985 ) );
  MUX U263 ( .IN0(\Reg_Bank/registers[30][28] ), .IN1(n148), .SEL(n180), .F(
        \Reg_Bank/n3984 ) );
  MUX U264 ( .IN0(\Reg_Bank/registers[30][27] ), .IN1(n149), .SEL(n180), .F(
        \Reg_Bank/n3983 ) );
  MUX U265 ( .IN0(\Reg_Bank/registers[30][26] ), .IN1(n150), .SEL(n180), .F(
        \Reg_Bank/n3982 ) );
  MUX U266 ( .IN0(\Reg_Bank/registers[30][25] ), .IN1(n151), .SEL(n180), .F(
        \Reg_Bank/n3981 ) );
  MUX U267 ( .IN0(\Reg_Bank/registers[30][24] ), .IN1(n152), .SEL(n180), .F(
        \Reg_Bank/n3980 ) );
  MUX U268 ( .IN0(\Reg_Bank/registers[30][23] ), .IN1(n153), .SEL(n180), .F(
        \Reg_Bank/n3979 ) );
  MUX U269 ( .IN0(\Reg_Bank/registers[30][22] ), .IN1(n154), .SEL(n180), .F(
        \Reg_Bank/n3978 ) );
  MUX U270 ( .IN0(\Reg_Bank/registers[30][21] ), .IN1(n155), .SEL(n180), .F(
        \Reg_Bank/n3977 ) );
  MUX U271 ( .IN0(\Reg_Bank/registers[30][20] ), .IN1(n156), .SEL(n180), .F(
        \Reg_Bank/n3976 ) );
  MUX U272 ( .IN0(\Reg_Bank/registers[30][19] ), .IN1(n157), .SEL(n180), .F(
        \Reg_Bank/n3975 ) );
  MUX U273 ( .IN0(\Reg_Bank/registers[30][18] ), .IN1(n158), .SEL(n180), .F(
        \Reg_Bank/n3974 ) );
  MUX U274 ( .IN0(\Reg_Bank/registers[30][17] ), .IN1(n159), .SEL(n180), .F(
        \Reg_Bank/n3973 ) );
  MUX U275 ( .IN0(\Reg_Bank/registers[30][16] ), .IN1(n160), .SEL(n180), .F(
        \Reg_Bank/n3972 ) );
  MUX U276 ( .IN0(\Reg_Bank/registers[30][15] ), .IN1(n161), .SEL(n180), .F(
        \Reg_Bank/n3971 ) );
  MUX U277 ( .IN0(\Reg_Bank/registers[30][14] ), .IN1(n162), .SEL(n180), .F(
        \Reg_Bank/n3970 ) );
  MUX U278 ( .IN0(\Reg_Bank/registers[30][13] ), .IN1(n163), .SEL(n180), .F(
        \Reg_Bank/n3969 ) );
  MUX U279 ( .IN0(\Reg_Bank/registers[30][12] ), .IN1(n164), .SEL(n180), .F(
        \Reg_Bank/n3968 ) );
  MUX U280 ( .IN0(\Reg_Bank/registers[30][11] ), .IN1(n165), .SEL(n180), .F(
        \Reg_Bank/n3967 ) );
  MUX U281 ( .IN0(\Reg_Bank/registers[30][10] ), .IN1(n166), .SEL(n180), .F(
        \Reg_Bank/n3966 ) );
  MUX U282 ( .IN0(\Reg_Bank/registers[30][9] ), .IN1(n167), .SEL(n180), .F(
        \Reg_Bank/n3965 ) );
  MUX U283 ( .IN0(\Reg_Bank/registers[30][8] ), .IN1(n168), .SEL(n180), .F(
        \Reg_Bank/n3964 ) );
  MUX U284 ( .IN0(\Reg_Bank/registers[30][7] ), .IN1(n169), .SEL(n180), .F(
        \Reg_Bank/n3963 ) );
  MUX U285 ( .IN0(\Reg_Bank/registers[30][6] ), .IN1(n170), .SEL(n180), .F(
        \Reg_Bank/n3962 ) );
  MUX U286 ( .IN0(\Reg_Bank/registers[30][5] ), .IN1(n171), .SEL(n180), .F(
        \Reg_Bank/n3961 ) );
  MUX U287 ( .IN0(\Reg_Bank/registers[30][4] ), .IN1(n172), .SEL(n180), .F(
        \Reg_Bank/n3960 ) );
  MUX U288 ( .IN0(\Reg_Bank/registers[30][3] ), .IN1(n173), .SEL(n180), .F(
        \Reg_Bank/n3959 ) );
  MUX U289 ( .IN0(\Reg_Bank/registers[30][2] ), .IN1(n174), .SEL(n180), .F(
        \Reg_Bank/n3958 ) );
  IV U290 ( .A(n181), .Z(n180) );
  MUX U291 ( .IN0(n176), .IN1(\Reg_Bank/registers[30][1] ), .SEL(n181), .F(
        \Reg_Bank/n3957 ) );
  MUX U292 ( .IN0(n177), .IN1(\Reg_Bank/registers[30][0] ), .SEL(n181), .F(
        \Reg_Bank/n3956 ) );
  NAND U293 ( .A(n179), .B(n182), .Z(n181) );
  MUX U294 ( .IN0(\Reg_Bank/registers[29][31] ), .IN1(n144), .SEL(n183), .F(
        \Reg_Bank/n3955 ) );
  MUX U295 ( .IN0(\Reg_Bank/registers[29][30] ), .IN1(n146), .SEL(n183), .F(
        \Reg_Bank/n3954 ) );
  MUX U296 ( .IN0(\Reg_Bank/registers[29][29] ), .IN1(n147), .SEL(n183), .F(
        \Reg_Bank/n3953 ) );
  MUX U297 ( .IN0(\Reg_Bank/registers[29][28] ), .IN1(n148), .SEL(n183), .F(
        \Reg_Bank/n3952 ) );
  MUX U298 ( .IN0(\Reg_Bank/registers[29][27] ), .IN1(n149), .SEL(n183), .F(
        \Reg_Bank/n3951 ) );
  MUX U299 ( .IN0(\Reg_Bank/registers[29][26] ), .IN1(n150), .SEL(n183), .F(
        \Reg_Bank/n3950 ) );
  MUX U300 ( .IN0(\Reg_Bank/registers[29][25] ), .IN1(n151), .SEL(n183), .F(
        \Reg_Bank/n3949 ) );
  MUX U301 ( .IN0(\Reg_Bank/registers[29][24] ), .IN1(n152), .SEL(n183), .F(
        \Reg_Bank/n3948 ) );
  MUX U302 ( .IN0(\Reg_Bank/registers[29][23] ), .IN1(n153), .SEL(n183), .F(
        \Reg_Bank/n3947 ) );
  MUX U303 ( .IN0(\Reg_Bank/registers[29][22] ), .IN1(n154), .SEL(n183), .F(
        \Reg_Bank/n3946 ) );
  MUX U304 ( .IN0(\Reg_Bank/registers[29][21] ), .IN1(n155), .SEL(n183), .F(
        \Reg_Bank/n3945 ) );
  MUX U305 ( .IN0(\Reg_Bank/registers[29][20] ), .IN1(n156), .SEL(n183), .F(
        \Reg_Bank/n3944 ) );
  MUX U306 ( .IN0(\Reg_Bank/registers[29][19] ), .IN1(n157), .SEL(n183), .F(
        \Reg_Bank/n3943 ) );
  MUX U307 ( .IN0(\Reg_Bank/registers[29][18] ), .IN1(n158), .SEL(n183), .F(
        \Reg_Bank/n3942 ) );
  MUX U308 ( .IN0(\Reg_Bank/registers[29][17] ), .IN1(n159), .SEL(n183), .F(
        \Reg_Bank/n3941 ) );
  MUX U309 ( .IN0(\Reg_Bank/registers[29][16] ), .IN1(n160), .SEL(n183), .F(
        \Reg_Bank/n3940 ) );
  MUX U310 ( .IN0(\Reg_Bank/registers[29][15] ), .IN1(n161), .SEL(n183), .F(
        \Reg_Bank/n3939 ) );
  MUX U311 ( .IN0(\Reg_Bank/registers[29][14] ), .IN1(n162), .SEL(n183), .F(
        \Reg_Bank/n3938 ) );
  MUX U312 ( .IN0(\Reg_Bank/registers[29][13] ), .IN1(n163), .SEL(n183), .F(
        \Reg_Bank/n3937 ) );
  MUX U313 ( .IN0(\Reg_Bank/registers[29][12] ), .IN1(n164), .SEL(n183), .F(
        \Reg_Bank/n3936 ) );
  MUX U314 ( .IN0(\Reg_Bank/registers[29][11] ), .IN1(n165), .SEL(n183), .F(
        \Reg_Bank/n3935 ) );
  MUX U315 ( .IN0(\Reg_Bank/registers[29][10] ), .IN1(n166), .SEL(n183), .F(
        \Reg_Bank/n3934 ) );
  MUX U316 ( .IN0(\Reg_Bank/registers[29][9] ), .IN1(n167), .SEL(n183), .F(
        \Reg_Bank/n3933 ) );
  MUX U317 ( .IN0(\Reg_Bank/registers[29][8] ), .IN1(n168), .SEL(n183), .F(
        \Reg_Bank/n3932 ) );
  MUX U318 ( .IN0(\Reg_Bank/registers[29][7] ), .IN1(n169), .SEL(n183), .F(
        \Reg_Bank/n3931 ) );
  MUX U319 ( .IN0(\Reg_Bank/registers[29][6] ), .IN1(n170), .SEL(n183), .F(
        \Reg_Bank/n3930 ) );
  MUX U320 ( .IN0(\Reg_Bank/registers[29][5] ), .IN1(n171), .SEL(n183), .F(
        \Reg_Bank/n3929 ) );
  MUX U321 ( .IN0(\Reg_Bank/registers[29][4] ), .IN1(n172), .SEL(n183), .F(
        \Reg_Bank/n3928 ) );
  MUX U322 ( .IN0(\Reg_Bank/registers[29][3] ), .IN1(n173), .SEL(n183), .F(
        \Reg_Bank/n3927 ) );
  MUX U323 ( .IN0(\Reg_Bank/registers[29][2] ), .IN1(n174), .SEL(n183), .F(
        \Reg_Bank/n3926 ) );
  IV U324 ( .A(n184), .Z(n183) );
  MUX U325 ( .IN0(n176), .IN1(\Reg_Bank/registers[29][1] ), .SEL(n184), .F(
        \Reg_Bank/n3925 ) );
  MUX U326 ( .IN0(n177), .IN1(\Reg_Bank/registers[29][0] ), .SEL(n184), .F(
        \Reg_Bank/n3924 ) );
  NAND U327 ( .A(n179), .B(n185), .Z(n184) );
  MUX U328 ( .IN0(\Reg_Bank/registers[28][31] ), .IN1(n144), .SEL(n186), .F(
        \Reg_Bank/n3923 ) );
  MUX U329 ( .IN0(\Reg_Bank/registers[28][30] ), .IN1(n146), .SEL(n186), .F(
        \Reg_Bank/n3922 ) );
  MUX U330 ( .IN0(\Reg_Bank/registers[28][29] ), .IN1(n147), .SEL(n186), .F(
        \Reg_Bank/n3921 ) );
  MUX U331 ( .IN0(\Reg_Bank/registers[28][28] ), .IN1(n148), .SEL(n186), .F(
        \Reg_Bank/n3920 ) );
  MUX U332 ( .IN0(\Reg_Bank/registers[28][27] ), .IN1(n149), .SEL(n186), .F(
        \Reg_Bank/n3919 ) );
  MUX U333 ( .IN0(\Reg_Bank/registers[28][26] ), .IN1(n150), .SEL(n186), .F(
        \Reg_Bank/n3918 ) );
  MUX U334 ( .IN0(\Reg_Bank/registers[28][25] ), .IN1(n151), .SEL(n186), .F(
        \Reg_Bank/n3917 ) );
  MUX U335 ( .IN0(\Reg_Bank/registers[28][24] ), .IN1(n152), .SEL(n186), .F(
        \Reg_Bank/n3916 ) );
  MUX U336 ( .IN0(\Reg_Bank/registers[28][23] ), .IN1(n153), .SEL(n186), .F(
        \Reg_Bank/n3915 ) );
  MUX U337 ( .IN0(\Reg_Bank/registers[28][22] ), .IN1(n154), .SEL(n186), .F(
        \Reg_Bank/n3914 ) );
  MUX U338 ( .IN0(\Reg_Bank/registers[28][21] ), .IN1(n155), .SEL(n186), .F(
        \Reg_Bank/n3913 ) );
  MUX U339 ( .IN0(\Reg_Bank/registers[28][20] ), .IN1(n156), .SEL(n186), .F(
        \Reg_Bank/n3912 ) );
  MUX U340 ( .IN0(\Reg_Bank/registers[28][19] ), .IN1(n157), .SEL(n186), .F(
        \Reg_Bank/n3911 ) );
  MUX U341 ( .IN0(\Reg_Bank/registers[28][18] ), .IN1(n158), .SEL(n186), .F(
        \Reg_Bank/n3910 ) );
  MUX U342 ( .IN0(\Reg_Bank/registers[28][17] ), .IN1(n159), .SEL(n186), .F(
        \Reg_Bank/n3909 ) );
  MUX U343 ( .IN0(\Reg_Bank/registers[28][16] ), .IN1(n160), .SEL(n186), .F(
        \Reg_Bank/n3908 ) );
  MUX U344 ( .IN0(\Reg_Bank/registers[28][15] ), .IN1(n161), .SEL(n186), .F(
        \Reg_Bank/n3907 ) );
  MUX U345 ( .IN0(\Reg_Bank/registers[28][14] ), .IN1(n162), .SEL(n186), .F(
        \Reg_Bank/n3906 ) );
  MUX U346 ( .IN0(\Reg_Bank/registers[28][13] ), .IN1(n163), .SEL(n186), .F(
        \Reg_Bank/n3905 ) );
  MUX U347 ( .IN0(\Reg_Bank/registers[28][12] ), .IN1(n164), .SEL(n186), .F(
        \Reg_Bank/n3904 ) );
  MUX U348 ( .IN0(\Reg_Bank/registers[28][11] ), .IN1(n165), .SEL(n186), .F(
        \Reg_Bank/n3903 ) );
  MUX U349 ( .IN0(\Reg_Bank/registers[28][10] ), .IN1(n166), .SEL(n186), .F(
        \Reg_Bank/n3902 ) );
  MUX U350 ( .IN0(\Reg_Bank/registers[28][9] ), .IN1(n167), .SEL(n186), .F(
        \Reg_Bank/n3901 ) );
  MUX U351 ( .IN0(\Reg_Bank/registers[28][8] ), .IN1(n168), .SEL(n186), .F(
        \Reg_Bank/n3900 ) );
  MUX U352 ( .IN0(\Reg_Bank/registers[28][7] ), .IN1(n169), .SEL(n186), .F(
        \Reg_Bank/n3899 ) );
  MUX U353 ( .IN0(\Reg_Bank/registers[28][6] ), .IN1(n170), .SEL(n186), .F(
        \Reg_Bank/n3898 ) );
  MUX U354 ( .IN0(\Reg_Bank/registers[28][5] ), .IN1(n171), .SEL(n186), .F(
        \Reg_Bank/n3897 ) );
  MUX U355 ( .IN0(\Reg_Bank/registers[28][4] ), .IN1(n172), .SEL(n186), .F(
        \Reg_Bank/n3896 ) );
  MUX U356 ( .IN0(\Reg_Bank/registers[28][3] ), .IN1(n173), .SEL(n186), .F(
        \Reg_Bank/n3895 ) );
  MUX U357 ( .IN0(\Reg_Bank/registers[28][2] ), .IN1(n174), .SEL(n186), .F(
        \Reg_Bank/n3894 ) );
  IV U358 ( .A(n187), .Z(n186) );
  MUX U359 ( .IN0(n176), .IN1(\Reg_Bank/registers[28][1] ), .SEL(n187), .F(
        \Reg_Bank/n3893 ) );
  MUX U360 ( .IN0(n177), .IN1(\Reg_Bank/registers[28][0] ), .SEL(n187), .F(
        \Reg_Bank/n3892 ) );
  NAND U361 ( .A(n179), .B(n188), .Z(n187) );
  MUX U362 ( .IN0(\Reg_Bank/registers[27][31] ), .IN1(n144), .SEL(n189), .F(
        \Reg_Bank/n3891 ) );
  MUX U363 ( .IN0(\Reg_Bank/registers[27][30] ), .IN1(n146), .SEL(n189), .F(
        \Reg_Bank/n3890 ) );
  MUX U364 ( .IN0(\Reg_Bank/registers[27][29] ), .IN1(n147), .SEL(n189), .F(
        \Reg_Bank/n3889 ) );
  MUX U365 ( .IN0(\Reg_Bank/registers[27][28] ), .IN1(n148), .SEL(n189), .F(
        \Reg_Bank/n3888 ) );
  MUX U366 ( .IN0(\Reg_Bank/registers[27][27] ), .IN1(n149), .SEL(n189), .F(
        \Reg_Bank/n3887 ) );
  MUX U367 ( .IN0(\Reg_Bank/registers[27][26] ), .IN1(n150), .SEL(n189), .F(
        \Reg_Bank/n3886 ) );
  MUX U368 ( .IN0(\Reg_Bank/registers[27][25] ), .IN1(n151), .SEL(n189), .F(
        \Reg_Bank/n3885 ) );
  MUX U369 ( .IN0(\Reg_Bank/registers[27][24] ), .IN1(n152), .SEL(n189), .F(
        \Reg_Bank/n3884 ) );
  MUX U370 ( .IN0(\Reg_Bank/registers[27][23] ), .IN1(n153), .SEL(n189), .F(
        \Reg_Bank/n3883 ) );
  MUX U371 ( .IN0(\Reg_Bank/registers[27][22] ), .IN1(n154), .SEL(n189), .F(
        \Reg_Bank/n3882 ) );
  MUX U372 ( .IN0(\Reg_Bank/registers[27][21] ), .IN1(n155), .SEL(n189), .F(
        \Reg_Bank/n3881 ) );
  MUX U373 ( .IN0(\Reg_Bank/registers[27][20] ), .IN1(n156), .SEL(n189), .F(
        \Reg_Bank/n3880 ) );
  MUX U374 ( .IN0(\Reg_Bank/registers[27][19] ), .IN1(n157), .SEL(n189), .F(
        \Reg_Bank/n3879 ) );
  MUX U375 ( .IN0(\Reg_Bank/registers[27][18] ), .IN1(n158), .SEL(n189), .F(
        \Reg_Bank/n3878 ) );
  MUX U376 ( .IN0(\Reg_Bank/registers[27][17] ), .IN1(n159), .SEL(n189), .F(
        \Reg_Bank/n3877 ) );
  MUX U377 ( .IN0(\Reg_Bank/registers[27][16] ), .IN1(n160), .SEL(n189), .F(
        \Reg_Bank/n3876 ) );
  MUX U378 ( .IN0(\Reg_Bank/registers[27][15] ), .IN1(n161), .SEL(n189), .F(
        \Reg_Bank/n3875 ) );
  MUX U379 ( .IN0(\Reg_Bank/registers[27][14] ), .IN1(n162), .SEL(n189), .F(
        \Reg_Bank/n3874 ) );
  MUX U380 ( .IN0(\Reg_Bank/registers[27][13] ), .IN1(n163), .SEL(n189), .F(
        \Reg_Bank/n3873 ) );
  MUX U381 ( .IN0(\Reg_Bank/registers[27][12] ), .IN1(n164), .SEL(n189), .F(
        \Reg_Bank/n3872 ) );
  MUX U382 ( .IN0(\Reg_Bank/registers[27][11] ), .IN1(n165), .SEL(n189), .F(
        \Reg_Bank/n3871 ) );
  MUX U383 ( .IN0(\Reg_Bank/registers[27][10] ), .IN1(n166), .SEL(n189), .F(
        \Reg_Bank/n3870 ) );
  MUX U384 ( .IN0(\Reg_Bank/registers[27][9] ), .IN1(n167), .SEL(n189), .F(
        \Reg_Bank/n3869 ) );
  MUX U385 ( .IN0(\Reg_Bank/registers[27][8] ), .IN1(n168), .SEL(n189), .F(
        \Reg_Bank/n3868 ) );
  MUX U386 ( .IN0(\Reg_Bank/registers[27][7] ), .IN1(n169), .SEL(n189), .F(
        \Reg_Bank/n3867 ) );
  MUX U387 ( .IN0(\Reg_Bank/registers[27][6] ), .IN1(n170), .SEL(n189), .F(
        \Reg_Bank/n3866 ) );
  MUX U388 ( .IN0(\Reg_Bank/registers[27][5] ), .IN1(n171), .SEL(n189), .F(
        \Reg_Bank/n3865 ) );
  MUX U389 ( .IN0(\Reg_Bank/registers[27][4] ), .IN1(n172), .SEL(n189), .F(
        \Reg_Bank/n3864 ) );
  MUX U390 ( .IN0(\Reg_Bank/registers[27][3] ), .IN1(n173), .SEL(n189), .F(
        \Reg_Bank/n3863 ) );
  MUX U391 ( .IN0(\Reg_Bank/registers[27][2] ), .IN1(n174), .SEL(n189), .F(
        \Reg_Bank/n3862 ) );
  MUX U392 ( .IN0(\Reg_Bank/registers[27][1] ), .IN1(n176), .SEL(n189), .F(
        \Reg_Bank/n3861 ) );
  MUX U393 ( .IN0(\Reg_Bank/registers[27][0] ), .IN1(n177), .SEL(n189), .F(
        \Reg_Bank/n3860 ) );
  ANDN U394 ( .A(n179), .B(n190), .Z(n189) );
  MUX U395 ( .IN0(\Reg_Bank/registers[26][31] ), .IN1(n144), .SEL(n191), .F(
        \Reg_Bank/n3859 ) );
  MUX U396 ( .IN0(\Reg_Bank/registers[26][30] ), .IN1(n146), .SEL(n191), .F(
        \Reg_Bank/n3858 ) );
  MUX U397 ( .IN0(\Reg_Bank/registers[26][29] ), .IN1(n147), .SEL(n191), .F(
        \Reg_Bank/n3857 ) );
  MUX U398 ( .IN0(\Reg_Bank/registers[26][28] ), .IN1(n148), .SEL(n191), .F(
        \Reg_Bank/n3856 ) );
  MUX U399 ( .IN0(\Reg_Bank/registers[26][27] ), .IN1(n149), .SEL(n191), .F(
        \Reg_Bank/n3855 ) );
  MUX U400 ( .IN0(\Reg_Bank/registers[26][26] ), .IN1(n150), .SEL(n191), .F(
        \Reg_Bank/n3854 ) );
  MUX U401 ( .IN0(\Reg_Bank/registers[26][25] ), .IN1(n151), .SEL(n191), .F(
        \Reg_Bank/n3853 ) );
  MUX U402 ( .IN0(\Reg_Bank/registers[26][24] ), .IN1(n152), .SEL(n191), .F(
        \Reg_Bank/n3852 ) );
  MUX U403 ( .IN0(\Reg_Bank/registers[26][23] ), .IN1(n153), .SEL(n191), .F(
        \Reg_Bank/n3851 ) );
  MUX U404 ( .IN0(\Reg_Bank/registers[26][22] ), .IN1(n154), .SEL(n191), .F(
        \Reg_Bank/n3850 ) );
  MUX U405 ( .IN0(\Reg_Bank/registers[26][21] ), .IN1(n155), .SEL(n191), .F(
        \Reg_Bank/n3849 ) );
  MUX U406 ( .IN0(\Reg_Bank/registers[26][20] ), .IN1(n156), .SEL(n191), .F(
        \Reg_Bank/n3848 ) );
  MUX U407 ( .IN0(\Reg_Bank/registers[26][19] ), .IN1(n157), .SEL(n191), .F(
        \Reg_Bank/n3847 ) );
  MUX U408 ( .IN0(\Reg_Bank/registers[26][18] ), .IN1(n158), .SEL(n191), .F(
        \Reg_Bank/n3846 ) );
  MUX U409 ( .IN0(\Reg_Bank/registers[26][17] ), .IN1(n159), .SEL(n191), .F(
        \Reg_Bank/n3845 ) );
  MUX U410 ( .IN0(\Reg_Bank/registers[26][16] ), .IN1(n160), .SEL(n191), .F(
        \Reg_Bank/n3844 ) );
  MUX U411 ( .IN0(\Reg_Bank/registers[26][15] ), .IN1(n161), .SEL(n191), .F(
        \Reg_Bank/n3843 ) );
  MUX U412 ( .IN0(\Reg_Bank/registers[26][14] ), .IN1(n162), .SEL(n191), .F(
        \Reg_Bank/n3842 ) );
  MUX U413 ( .IN0(\Reg_Bank/registers[26][13] ), .IN1(n163), .SEL(n191), .F(
        \Reg_Bank/n3841 ) );
  MUX U414 ( .IN0(\Reg_Bank/registers[26][12] ), .IN1(n164), .SEL(n191), .F(
        \Reg_Bank/n3840 ) );
  MUX U415 ( .IN0(\Reg_Bank/registers[26][11] ), .IN1(n165), .SEL(n191), .F(
        \Reg_Bank/n3839 ) );
  MUX U416 ( .IN0(\Reg_Bank/registers[26][10] ), .IN1(n166), .SEL(n191), .F(
        \Reg_Bank/n3838 ) );
  MUX U417 ( .IN0(\Reg_Bank/registers[26][9] ), .IN1(n167), .SEL(n191), .F(
        \Reg_Bank/n3837 ) );
  MUX U418 ( .IN0(\Reg_Bank/registers[26][8] ), .IN1(n168), .SEL(n191), .F(
        \Reg_Bank/n3836 ) );
  MUX U419 ( .IN0(\Reg_Bank/registers[26][7] ), .IN1(n169), .SEL(n191), .F(
        \Reg_Bank/n3835 ) );
  MUX U420 ( .IN0(\Reg_Bank/registers[26][6] ), .IN1(n170), .SEL(n191), .F(
        \Reg_Bank/n3834 ) );
  MUX U421 ( .IN0(\Reg_Bank/registers[26][5] ), .IN1(n171), .SEL(n191), .F(
        \Reg_Bank/n3833 ) );
  MUX U422 ( .IN0(\Reg_Bank/registers[26][4] ), .IN1(n172), .SEL(n191), .F(
        \Reg_Bank/n3832 ) );
  MUX U423 ( .IN0(\Reg_Bank/registers[26][3] ), .IN1(n173), .SEL(n191), .F(
        \Reg_Bank/n3831 ) );
  MUX U424 ( .IN0(\Reg_Bank/registers[26][2] ), .IN1(n174), .SEL(n191), .F(
        \Reg_Bank/n3830 ) );
  MUX U425 ( .IN0(\Reg_Bank/registers[26][1] ), .IN1(n176), .SEL(n191), .F(
        \Reg_Bank/n3829 ) );
  MUX U426 ( .IN0(\Reg_Bank/registers[26][0] ), .IN1(n177), .SEL(n191), .F(
        \Reg_Bank/n3828 ) );
  ANDN U427 ( .A(n179), .B(n192), .Z(n191) );
  MUX U428 ( .IN0(\Reg_Bank/registers[25][31] ), .IN1(n144), .SEL(n193), .F(
        \Reg_Bank/n3827 ) );
  MUX U429 ( .IN0(\Reg_Bank/registers[25][30] ), .IN1(n146), .SEL(n193), .F(
        \Reg_Bank/n3826 ) );
  MUX U430 ( .IN0(\Reg_Bank/registers[25][29] ), .IN1(n147), .SEL(n193), .F(
        \Reg_Bank/n3825 ) );
  MUX U431 ( .IN0(\Reg_Bank/registers[25][28] ), .IN1(n148), .SEL(n193), .F(
        \Reg_Bank/n3824 ) );
  MUX U432 ( .IN0(\Reg_Bank/registers[25][27] ), .IN1(n149), .SEL(n193), .F(
        \Reg_Bank/n3823 ) );
  MUX U433 ( .IN0(\Reg_Bank/registers[25][26] ), .IN1(n150), .SEL(n193), .F(
        \Reg_Bank/n3822 ) );
  MUX U434 ( .IN0(\Reg_Bank/registers[25][25] ), .IN1(n151), .SEL(n193), .F(
        \Reg_Bank/n3821 ) );
  MUX U435 ( .IN0(\Reg_Bank/registers[25][24] ), .IN1(n152), .SEL(n193), .F(
        \Reg_Bank/n3820 ) );
  MUX U436 ( .IN0(\Reg_Bank/registers[25][23] ), .IN1(n153), .SEL(n193), .F(
        \Reg_Bank/n3819 ) );
  MUX U437 ( .IN0(\Reg_Bank/registers[25][22] ), .IN1(n154), .SEL(n193), .F(
        \Reg_Bank/n3818 ) );
  MUX U438 ( .IN0(\Reg_Bank/registers[25][21] ), .IN1(n155), .SEL(n193), .F(
        \Reg_Bank/n3817 ) );
  MUX U439 ( .IN0(\Reg_Bank/registers[25][20] ), .IN1(n156), .SEL(n193), .F(
        \Reg_Bank/n3816 ) );
  MUX U440 ( .IN0(\Reg_Bank/registers[25][19] ), .IN1(n157), .SEL(n193), .F(
        \Reg_Bank/n3815 ) );
  MUX U441 ( .IN0(\Reg_Bank/registers[25][18] ), .IN1(n158), .SEL(n193), .F(
        \Reg_Bank/n3814 ) );
  MUX U442 ( .IN0(\Reg_Bank/registers[25][17] ), .IN1(n159), .SEL(n193), .F(
        \Reg_Bank/n3813 ) );
  MUX U443 ( .IN0(\Reg_Bank/registers[25][16] ), .IN1(n160), .SEL(n193), .F(
        \Reg_Bank/n3812 ) );
  MUX U444 ( .IN0(\Reg_Bank/registers[25][15] ), .IN1(n161), .SEL(n193), .F(
        \Reg_Bank/n3811 ) );
  MUX U445 ( .IN0(\Reg_Bank/registers[25][14] ), .IN1(n162), .SEL(n193), .F(
        \Reg_Bank/n3810 ) );
  MUX U446 ( .IN0(\Reg_Bank/registers[25][13] ), .IN1(n163), .SEL(n193), .F(
        \Reg_Bank/n3809 ) );
  MUX U447 ( .IN0(\Reg_Bank/registers[25][12] ), .IN1(n164), .SEL(n193), .F(
        \Reg_Bank/n3808 ) );
  MUX U448 ( .IN0(\Reg_Bank/registers[25][11] ), .IN1(n165), .SEL(n193), .F(
        \Reg_Bank/n3807 ) );
  MUX U449 ( .IN0(\Reg_Bank/registers[25][10] ), .IN1(n166), .SEL(n193), .F(
        \Reg_Bank/n3806 ) );
  MUX U450 ( .IN0(\Reg_Bank/registers[25][9] ), .IN1(n167), .SEL(n193), .F(
        \Reg_Bank/n3805 ) );
  MUX U451 ( .IN0(\Reg_Bank/registers[25][8] ), .IN1(n168), .SEL(n193), .F(
        \Reg_Bank/n3804 ) );
  MUX U452 ( .IN0(\Reg_Bank/registers[25][7] ), .IN1(n169), .SEL(n193), .F(
        \Reg_Bank/n3803 ) );
  MUX U453 ( .IN0(\Reg_Bank/registers[25][6] ), .IN1(n170), .SEL(n193), .F(
        \Reg_Bank/n3802 ) );
  MUX U454 ( .IN0(\Reg_Bank/registers[25][5] ), .IN1(n171), .SEL(n193), .F(
        \Reg_Bank/n3801 ) );
  MUX U455 ( .IN0(\Reg_Bank/registers[25][4] ), .IN1(n172), .SEL(n193), .F(
        \Reg_Bank/n3800 ) );
  MUX U456 ( .IN0(\Reg_Bank/registers[25][3] ), .IN1(n173), .SEL(n193), .F(
        \Reg_Bank/n3799 ) );
  MUX U457 ( .IN0(\Reg_Bank/registers[25][2] ), .IN1(n174), .SEL(n193), .F(
        \Reg_Bank/n3798 ) );
  MUX U458 ( .IN0(\Reg_Bank/registers[25][1] ), .IN1(n176), .SEL(n193), .F(
        \Reg_Bank/n3797 ) );
  MUX U459 ( .IN0(\Reg_Bank/registers[25][0] ), .IN1(n177), .SEL(n193), .F(
        \Reg_Bank/n3796 ) );
  ANDN U460 ( .A(n179), .B(n194), .Z(n193) );
  MUX U461 ( .IN0(\Reg_Bank/registers[24][31] ), .IN1(n144), .SEL(n195), .F(
        \Reg_Bank/n3795 ) );
  MUX U462 ( .IN0(\Reg_Bank/registers[24][30] ), .IN1(n146), .SEL(n195), .F(
        \Reg_Bank/n3794 ) );
  MUX U463 ( .IN0(\Reg_Bank/registers[24][29] ), .IN1(n147), .SEL(n195), .F(
        \Reg_Bank/n3793 ) );
  MUX U464 ( .IN0(\Reg_Bank/registers[24][28] ), .IN1(n148), .SEL(n195), .F(
        \Reg_Bank/n3792 ) );
  MUX U465 ( .IN0(\Reg_Bank/registers[24][27] ), .IN1(n149), .SEL(n195), .F(
        \Reg_Bank/n3791 ) );
  MUX U466 ( .IN0(\Reg_Bank/registers[24][26] ), .IN1(n150), .SEL(n195), .F(
        \Reg_Bank/n3790 ) );
  MUX U467 ( .IN0(\Reg_Bank/registers[24][25] ), .IN1(n151), .SEL(n195), .F(
        \Reg_Bank/n3789 ) );
  MUX U468 ( .IN0(\Reg_Bank/registers[24][24] ), .IN1(n152), .SEL(n195), .F(
        \Reg_Bank/n3788 ) );
  MUX U469 ( .IN0(\Reg_Bank/registers[24][23] ), .IN1(n153), .SEL(n195), .F(
        \Reg_Bank/n3787 ) );
  MUX U470 ( .IN0(\Reg_Bank/registers[24][22] ), .IN1(n154), .SEL(n195), .F(
        \Reg_Bank/n3786 ) );
  MUX U471 ( .IN0(\Reg_Bank/registers[24][21] ), .IN1(n155), .SEL(n195), .F(
        \Reg_Bank/n3785 ) );
  MUX U472 ( .IN0(\Reg_Bank/registers[24][20] ), .IN1(n156), .SEL(n195), .F(
        \Reg_Bank/n3784 ) );
  MUX U473 ( .IN0(\Reg_Bank/registers[24][19] ), .IN1(n157), .SEL(n195), .F(
        \Reg_Bank/n3783 ) );
  MUX U474 ( .IN0(\Reg_Bank/registers[24][18] ), .IN1(n158), .SEL(n195), .F(
        \Reg_Bank/n3782 ) );
  MUX U475 ( .IN0(\Reg_Bank/registers[24][17] ), .IN1(n159), .SEL(n195), .F(
        \Reg_Bank/n3781 ) );
  MUX U476 ( .IN0(\Reg_Bank/registers[24][16] ), .IN1(n160), .SEL(n195), .F(
        \Reg_Bank/n3780 ) );
  MUX U477 ( .IN0(\Reg_Bank/registers[24][15] ), .IN1(n161), .SEL(n195), .F(
        \Reg_Bank/n3779 ) );
  MUX U478 ( .IN0(\Reg_Bank/registers[24][14] ), .IN1(n162), .SEL(n195), .F(
        \Reg_Bank/n3778 ) );
  MUX U479 ( .IN0(\Reg_Bank/registers[24][13] ), .IN1(n163), .SEL(n195), .F(
        \Reg_Bank/n3777 ) );
  MUX U480 ( .IN0(\Reg_Bank/registers[24][12] ), .IN1(n164), .SEL(n195), .F(
        \Reg_Bank/n3776 ) );
  MUX U481 ( .IN0(\Reg_Bank/registers[24][11] ), .IN1(n165), .SEL(n195), .F(
        \Reg_Bank/n3775 ) );
  MUX U482 ( .IN0(\Reg_Bank/registers[24][10] ), .IN1(n166), .SEL(n195), .F(
        \Reg_Bank/n3774 ) );
  MUX U483 ( .IN0(\Reg_Bank/registers[24][9] ), .IN1(n167), .SEL(n195), .F(
        \Reg_Bank/n3773 ) );
  MUX U484 ( .IN0(\Reg_Bank/registers[24][8] ), .IN1(n168), .SEL(n195), .F(
        \Reg_Bank/n3772 ) );
  MUX U485 ( .IN0(\Reg_Bank/registers[24][7] ), .IN1(n169), .SEL(n195), .F(
        \Reg_Bank/n3771 ) );
  MUX U486 ( .IN0(\Reg_Bank/registers[24][6] ), .IN1(n170), .SEL(n195), .F(
        \Reg_Bank/n3770 ) );
  MUX U487 ( .IN0(\Reg_Bank/registers[24][5] ), .IN1(n171), .SEL(n195), .F(
        \Reg_Bank/n3769 ) );
  MUX U488 ( .IN0(\Reg_Bank/registers[24][4] ), .IN1(n172), .SEL(n195), .F(
        \Reg_Bank/n3768 ) );
  MUX U489 ( .IN0(\Reg_Bank/registers[24][3] ), .IN1(n173), .SEL(n195), .F(
        \Reg_Bank/n3767 ) );
  MUX U490 ( .IN0(\Reg_Bank/registers[24][2] ), .IN1(n174), .SEL(n195), .F(
        \Reg_Bank/n3766 ) );
  MUX U491 ( .IN0(\Reg_Bank/registers[24][1] ), .IN1(n176), .SEL(n195), .F(
        \Reg_Bank/n3765 ) );
  MUX U492 ( .IN0(\Reg_Bank/registers[24][0] ), .IN1(n177), .SEL(n195), .F(
        \Reg_Bank/n3764 ) );
  ANDN U493 ( .A(n179), .B(n196), .Z(n195) );
  ANDN U494 ( .A(n197), .B(n198), .Z(n179) );
  MUX U495 ( .IN0(\Reg_Bank/registers[23][31] ), .IN1(n144), .SEL(n199), .F(
        \Reg_Bank/n3763 ) );
  MUX U496 ( .IN0(\Reg_Bank/registers[23][30] ), .IN1(n146), .SEL(n199), .F(
        \Reg_Bank/n3762 ) );
  MUX U497 ( .IN0(\Reg_Bank/registers[23][29] ), .IN1(n147), .SEL(n199), .F(
        \Reg_Bank/n3761 ) );
  MUX U498 ( .IN0(\Reg_Bank/registers[23][28] ), .IN1(n148), .SEL(n199), .F(
        \Reg_Bank/n3760 ) );
  MUX U499 ( .IN0(\Reg_Bank/registers[23][27] ), .IN1(n149), .SEL(n199), .F(
        \Reg_Bank/n3759 ) );
  MUX U500 ( .IN0(\Reg_Bank/registers[23][26] ), .IN1(n150), .SEL(n199), .F(
        \Reg_Bank/n3758 ) );
  MUX U501 ( .IN0(\Reg_Bank/registers[23][25] ), .IN1(n151), .SEL(n199), .F(
        \Reg_Bank/n3757 ) );
  MUX U502 ( .IN0(\Reg_Bank/registers[23][24] ), .IN1(n152), .SEL(n199), .F(
        \Reg_Bank/n3756 ) );
  MUX U503 ( .IN0(\Reg_Bank/registers[23][23] ), .IN1(n153), .SEL(n199), .F(
        \Reg_Bank/n3755 ) );
  MUX U504 ( .IN0(\Reg_Bank/registers[23][22] ), .IN1(n154), .SEL(n199), .F(
        \Reg_Bank/n3754 ) );
  MUX U505 ( .IN0(\Reg_Bank/registers[23][21] ), .IN1(n155), .SEL(n199), .F(
        \Reg_Bank/n3753 ) );
  MUX U506 ( .IN0(\Reg_Bank/registers[23][20] ), .IN1(n156), .SEL(n199), .F(
        \Reg_Bank/n3752 ) );
  MUX U507 ( .IN0(\Reg_Bank/registers[23][19] ), .IN1(n157), .SEL(n199), .F(
        \Reg_Bank/n3751 ) );
  MUX U508 ( .IN0(\Reg_Bank/registers[23][18] ), .IN1(n158), .SEL(n199), .F(
        \Reg_Bank/n3750 ) );
  MUX U509 ( .IN0(\Reg_Bank/registers[23][17] ), .IN1(n159), .SEL(n199), .F(
        \Reg_Bank/n3749 ) );
  MUX U510 ( .IN0(\Reg_Bank/registers[23][16] ), .IN1(n160), .SEL(n199), .F(
        \Reg_Bank/n3748 ) );
  MUX U511 ( .IN0(\Reg_Bank/registers[23][15] ), .IN1(n161), .SEL(n199), .F(
        \Reg_Bank/n3747 ) );
  MUX U512 ( .IN0(\Reg_Bank/registers[23][14] ), .IN1(n162), .SEL(n199), .F(
        \Reg_Bank/n3746 ) );
  MUX U513 ( .IN0(\Reg_Bank/registers[23][13] ), .IN1(n163), .SEL(n199), .F(
        \Reg_Bank/n3745 ) );
  MUX U514 ( .IN0(\Reg_Bank/registers[23][12] ), .IN1(n164), .SEL(n199), .F(
        \Reg_Bank/n3744 ) );
  MUX U515 ( .IN0(\Reg_Bank/registers[23][11] ), .IN1(n165), .SEL(n199), .F(
        \Reg_Bank/n3743 ) );
  MUX U516 ( .IN0(\Reg_Bank/registers[23][10] ), .IN1(n166), .SEL(n199), .F(
        \Reg_Bank/n3742 ) );
  MUX U517 ( .IN0(\Reg_Bank/registers[23][9] ), .IN1(n167), .SEL(n199), .F(
        \Reg_Bank/n3741 ) );
  MUX U518 ( .IN0(\Reg_Bank/registers[23][8] ), .IN1(n168), .SEL(n199), .F(
        \Reg_Bank/n3740 ) );
  MUX U519 ( .IN0(\Reg_Bank/registers[23][7] ), .IN1(n169), .SEL(n199), .F(
        \Reg_Bank/n3739 ) );
  MUX U520 ( .IN0(\Reg_Bank/registers[23][6] ), .IN1(n170), .SEL(n199), .F(
        \Reg_Bank/n3738 ) );
  MUX U521 ( .IN0(\Reg_Bank/registers[23][5] ), .IN1(n171), .SEL(n199), .F(
        \Reg_Bank/n3737 ) );
  MUX U522 ( .IN0(\Reg_Bank/registers[23][4] ), .IN1(n172), .SEL(n199), .F(
        \Reg_Bank/n3736 ) );
  MUX U523 ( .IN0(\Reg_Bank/registers[23][3] ), .IN1(n173), .SEL(n199), .F(
        \Reg_Bank/n3735 ) );
  MUX U524 ( .IN0(\Reg_Bank/registers[23][2] ), .IN1(n174), .SEL(n199), .F(
        \Reg_Bank/n3734 ) );
  MUX U525 ( .IN0(\Reg_Bank/registers[23][1] ), .IN1(n176), .SEL(n199), .F(
        \Reg_Bank/n3733 ) );
  MUX U526 ( .IN0(\Reg_Bank/registers[23][0] ), .IN1(n177), .SEL(n199), .F(
        \Reg_Bank/n3732 ) );
  ANDN U527 ( .A(n200), .B(n178), .Z(n199) );
  MUX U528 ( .IN0(\Reg_Bank/registers[22][31] ), .IN1(n144), .SEL(n201), .F(
        \Reg_Bank/n3731 ) );
  MUX U529 ( .IN0(\Reg_Bank/registers[22][30] ), .IN1(n146), .SEL(n201), .F(
        \Reg_Bank/n3730 ) );
  MUX U530 ( .IN0(\Reg_Bank/registers[22][29] ), .IN1(n147), .SEL(n201), .F(
        \Reg_Bank/n3729 ) );
  MUX U531 ( .IN0(\Reg_Bank/registers[22][28] ), .IN1(n148), .SEL(n201), .F(
        \Reg_Bank/n3728 ) );
  MUX U532 ( .IN0(\Reg_Bank/registers[22][27] ), .IN1(n149), .SEL(n201), .F(
        \Reg_Bank/n3727 ) );
  MUX U533 ( .IN0(\Reg_Bank/registers[22][26] ), .IN1(n150), .SEL(n201), .F(
        \Reg_Bank/n3726 ) );
  MUX U534 ( .IN0(\Reg_Bank/registers[22][25] ), .IN1(n151), .SEL(n201), .F(
        \Reg_Bank/n3725 ) );
  MUX U535 ( .IN0(\Reg_Bank/registers[22][24] ), .IN1(n152), .SEL(n201), .F(
        \Reg_Bank/n3724 ) );
  MUX U536 ( .IN0(\Reg_Bank/registers[22][23] ), .IN1(n153), .SEL(n201), .F(
        \Reg_Bank/n3723 ) );
  MUX U537 ( .IN0(\Reg_Bank/registers[22][22] ), .IN1(n154), .SEL(n201), .F(
        \Reg_Bank/n3722 ) );
  MUX U538 ( .IN0(\Reg_Bank/registers[22][21] ), .IN1(n155), .SEL(n201), .F(
        \Reg_Bank/n3721 ) );
  MUX U539 ( .IN0(\Reg_Bank/registers[22][20] ), .IN1(n156), .SEL(n201), .F(
        \Reg_Bank/n3720 ) );
  MUX U540 ( .IN0(\Reg_Bank/registers[22][19] ), .IN1(n157), .SEL(n201), .F(
        \Reg_Bank/n3719 ) );
  MUX U541 ( .IN0(\Reg_Bank/registers[22][18] ), .IN1(n158), .SEL(n201), .F(
        \Reg_Bank/n3718 ) );
  MUX U542 ( .IN0(\Reg_Bank/registers[22][17] ), .IN1(n159), .SEL(n201), .F(
        \Reg_Bank/n3717 ) );
  MUX U543 ( .IN0(\Reg_Bank/registers[22][16] ), .IN1(n160), .SEL(n201), .F(
        \Reg_Bank/n3716 ) );
  MUX U544 ( .IN0(\Reg_Bank/registers[22][15] ), .IN1(n161), .SEL(n201), .F(
        \Reg_Bank/n3715 ) );
  MUX U545 ( .IN0(\Reg_Bank/registers[22][14] ), .IN1(n162), .SEL(n201), .F(
        \Reg_Bank/n3714 ) );
  MUX U546 ( .IN0(\Reg_Bank/registers[22][13] ), .IN1(n163), .SEL(n201), .F(
        \Reg_Bank/n3713 ) );
  MUX U547 ( .IN0(\Reg_Bank/registers[22][12] ), .IN1(n164), .SEL(n201), .F(
        \Reg_Bank/n3712 ) );
  MUX U548 ( .IN0(\Reg_Bank/registers[22][11] ), .IN1(n165), .SEL(n201), .F(
        \Reg_Bank/n3711 ) );
  MUX U549 ( .IN0(\Reg_Bank/registers[22][10] ), .IN1(n166), .SEL(n201), .F(
        \Reg_Bank/n3710 ) );
  MUX U550 ( .IN0(\Reg_Bank/registers[22][9] ), .IN1(n167), .SEL(n201), .F(
        \Reg_Bank/n3709 ) );
  MUX U551 ( .IN0(\Reg_Bank/registers[22][8] ), .IN1(n168), .SEL(n201), .F(
        \Reg_Bank/n3708 ) );
  MUX U552 ( .IN0(\Reg_Bank/registers[22][7] ), .IN1(n169), .SEL(n201), .F(
        \Reg_Bank/n3707 ) );
  MUX U553 ( .IN0(\Reg_Bank/registers[22][6] ), .IN1(n170), .SEL(n201), .F(
        \Reg_Bank/n3706 ) );
  MUX U554 ( .IN0(\Reg_Bank/registers[22][5] ), .IN1(n171), .SEL(n201), .F(
        \Reg_Bank/n3705 ) );
  MUX U555 ( .IN0(\Reg_Bank/registers[22][4] ), .IN1(n172), .SEL(n201), .F(
        \Reg_Bank/n3704 ) );
  MUX U556 ( .IN0(\Reg_Bank/registers[22][3] ), .IN1(n173), .SEL(n201), .F(
        \Reg_Bank/n3703 ) );
  MUX U557 ( .IN0(\Reg_Bank/registers[22][2] ), .IN1(n174), .SEL(n201), .F(
        \Reg_Bank/n3702 ) );
  MUX U558 ( .IN0(\Reg_Bank/registers[22][1] ), .IN1(n176), .SEL(n201), .F(
        \Reg_Bank/n3701 ) );
  MUX U559 ( .IN0(\Reg_Bank/registers[22][0] ), .IN1(n177), .SEL(n201), .F(
        \Reg_Bank/n3700 ) );
  AND U560 ( .A(n182), .B(n200), .Z(n201) );
  MUX U561 ( .IN0(\Reg_Bank/registers[21][31] ), .IN1(n144), .SEL(n202), .F(
        \Reg_Bank/n3699 ) );
  MUX U562 ( .IN0(\Reg_Bank/registers[21][30] ), .IN1(n146), .SEL(n202), .F(
        \Reg_Bank/n3698 ) );
  MUX U563 ( .IN0(\Reg_Bank/registers[21][29] ), .IN1(n147), .SEL(n202), .F(
        \Reg_Bank/n3697 ) );
  MUX U564 ( .IN0(\Reg_Bank/registers[21][28] ), .IN1(n148), .SEL(n202), .F(
        \Reg_Bank/n3696 ) );
  MUX U565 ( .IN0(\Reg_Bank/registers[21][27] ), .IN1(n149), .SEL(n202), .F(
        \Reg_Bank/n3695 ) );
  MUX U566 ( .IN0(\Reg_Bank/registers[21][26] ), .IN1(n150), .SEL(n202), .F(
        \Reg_Bank/n3694 ) );
  MUX U567 ( .IN0(\Reg_Bank/registers[21][25] ), .IN1(n151), .SEL(n202), .F(
        \Reg_Bank/n3693 ) );
  MUX U568 ( .IN0(\Reg_Bank/registers[21][24] ), .IN1(n152), .SEL(n202), .F(
        \Reg_Bank/n3692 ) );
  MUX U569 ( .IN0(\Reg_Bank/registers[21][23] ), .IN1(n153), .SEL(n202), .F(
        \Reg_Bank/n3691 ) );
  MUX U570 ( .IN0(\Reg_Bank/registers[21][22] ), .IN1(n154), .SEL(n202), .F(
        \Reg_Bank/n3690 ) );
  MUX U571 ( .IN0(\Reg_Bank/registers[21][21] ), .IN1(n155), .SEL(n202), .F(
        \Reg_Bank/n3689 ) );
  MUX U572 ( .IN0(\Reg_Bank/registers[21][20] ), .IN1(n156), .SEL(n202), .F(
        \Reg_Bank/n3688 ) );
  MUX U573 ( .IN0(\Reg_Bank/registers[21][19] ), .IN1(n157), .SEL(n202), .F(
        \Reg_Bank/n3687 ) );
  MUX U574 ( .IN0(\Reg_Bank/registers[21][18] ), .IN1(n158), .SEL(n202), .F(
        \Reg_Bank/n3686 ) );
  MUX U575 ( .IN0(\Reg_Bank/registers[21][17] ), .IN1(n159), .SEL(n202), .F(
        \Reg_Bank/n3685 ) );
  MUX U576 ( .IN0(\Reg_Bank/registers[21][16] ), .IN1(n160), .SEL(n202), .F(
        \Reg_Bank/n3684 ) );
  MUX U577 ( .IN0(\Reg_Bank/registers[21][15] ), .IN1(n161), .SEL(n202), .F(
        \Reg_Bank/n3683 ) );
  MUX U578 ( .IN0(\Reg_Bank/registers[21][14] ), .IN1(n162), .SEL(n202), .F(
        \Reg_Bank/n3682 ) );
  MUX U579 ( .IN0(\Reg_Bank/registers[21][13] ), .IN1(n163), .SEL(n202), .F(
        \Reg_Bank/n3681 ) );
  MUX U580 ( .IN0(\Reg_Bank/registers[21][12] ), .IN1(n164), .SEL(n202), .F(
        \Reg_Bank/n3680 ) );
  MUX U581 ( .IN0(\Reg_Bank/registers[21][11] ), .IN1(n165), .SEL(n202), .F(
        \Reg_Bank/n3679 ) );
  MUX U582 ( .IN0(\Reg_Bank/registers[21][10] ), .IN1(n166), .SEL(n202), .F(
        \Reg_Bank/n3678 ) );
  MUX U583 ( .IN0(\Reg_Bank/registers[21][9] ), .IN1(n167), .SEL(n202), .F(
        \Reg_Bank/n3677 ) );
  MUX U584 ( .IN0(\Reg_Bank/registers[21][8] ), .IN1(n168), .SEL(n202), .F(
        \Reg_Bank/n3676 ) );
  MUX U585 ( .IN0(\Reg_Bank/registers[21][7] ), .IN1(n169), .SEL(n202), .F(
        \Reg_Bank/n3675 ) );
  MUX U586 ( .IN0(\Reg_Bank/registers[21][6] ), .IN1(n170), .SEL(n202), .F(
        \Reg_Bank/n3674 ) );
  MUX U587 ( .IN0(\Reg_Bank/registers[21][5] ), .IN1(n171), .SEL(n202), .F(
        \Reg_Bank/n3673 ) );
  MUX U588 ( .IN0(\Reg_Bank/registers[21][4] ), .IN1(n172), .SEL(n202), .F(
        \Reg_Bank/n3672 ) );
  MUX U589 ( .IN0(\Reg_Bank/registers[21][3] ), .IN1(n173), .SEL(n202), .F(
        \Reg_Bank/n3671 ) );
  MUX U590 ( .IN0(\Reg_Bank/registers[21][2] ), .IN1(n174), .SEL(n202), .F(
        \Reg_Bank/n3670 ) );
  MUX U591 ( .IN0(\Reg_Bank/registers[21][1] ), .IN1(n176), .SEL(n202), .F(
        \Reg_Bank/n3669 ) );
  MUX U592 ( .IN0(\Reg_Bank/registers[21][0] ), .IN1(n177), .SEL(n202), .F(
        \Reg_Bank/n3668 ) );
  AND U593 ( .A(n185), .B(n200), .Z(n202) );
  MUX U594 ( .IN0(\Reg_Bank/registers[20][31] ), .IN1(n144), .SEL(n203), .F(
        \Reg_Bank/n3667 ) );
  MUX U595 ( .IN0(\Reg_Bank/registers[20][30] ), .IN1(n146), .SEL(n203), .F(
        \Reg_Bank/n3666 ) );
  MUX U596 ( .IN0(\Reg_Bank/registers[20][29] ), .IN1(n147), .SEL(n203), .F(
        \Reg_Bank/n3665 ) );
  MUX U597 ( .IN0(\Reg_Bank/registers[20][28] ), .IN1(n148), .SEL(n203), .F(
        \Reg_Bank/n3664 ) );
  MUX U598 ( .IN0(\Reg_Bank/registers[20][27] ), .IN1(n149), .SEL(n203), .F(
        \Reg_Bank/n3663 ) );
  MUX U599 ( .IN0(\Reg_Bank/registers[20][26] ), .IN1(n150), .SEL(n203), .F(
        \Reg_Bank/n3662 ) );
  MUX U600 ( .IN0(\Reg_Bank/registers[20][25] ), .IN1(n151), .SEL(n203), .F(
        \Reg_Bank/n3661 ) );
  MUX U601 ( .IN0(\Reg_Bank/registers[20][24] ), .IN1(n152), .SEL(n203), .F(
        \Reg_Bank/n3660 ) );
  MUX U602 ( .IN0(\Reg_Bank/registers[20][23] ), .IN1(n153), .SEL(n203), .F(
        \Reg_Bank/n3659 ) );
  MUX U603 ( .IN0(\Reg_Bank/registers[20][22] ), .IN1(n154), .SEL(n203), .F(
        \Reg_Bank/n3658 ) );
  MUX U604 ( .IN0(\Reg_Bank/registers[20][21] ), .IN1(n155), .SEL(n203), .F(
        \Reg_Bank/n3657 ) );
  MUX U605 ( .IN0(\Reg_Bank/registers[20][20] ), .IN1(n156), .SEL(n203), .F(
        \Reg_Bank/n3656 ) );
  MUX U606 ( .IN0(\Reg_Bank/registers[20][19] ), .IN1(n157), .SEL(n203), .F(
        \Reg_Bank/n3655 ) );
  MUX U607 ( .IN0(\Reg_Bank/registers[20][18] ), .IN1(n158), .SEL(n203), .F(
        \Reg_Bank/n3654 ) );
  MUX U608 ( .IN0(\Reg_Bank/registers[20][17] ), .IN1(n159), .SEL(n203), .F(
        \Reg_Bank/n3653 ) );
  MUX U609 ( .IN0(\Reg_Bank/registers[20][16] ), .IN1(n160), .SEL(n203), .F(
        \Reg_Bank/n3652 ) );
  MUX U610 ( .IN0(\Reg_Bank/registers[20][15] ), .IN1(n161), .SEL(n203), .F(
        \Reg_Bank/n3651 ) );
  MUX U611 ( .IN0(\Reg_Bank/registers[20][14] ), .IN1(n162), .SEL(n203), .F(
        \Reg_Bank/n3650 ) );
  MUX U612 ( .IN0(\Reg_Bank/registers[20][13] ), .IN1(n163), .SEL(n203), .F(
        \Reg_Bank/n3649 ) );
  MUX U613 ( .IN0(\Reg_Bank/registers[20][12] ), .IN1(n164), .SEL(n203), .F(
        \Reg_Bank/n3648 ) );
  MUX U614 ( .IN0(\Reg_Bank/registers[20][11] ), .IN1(n165), .SEL(n203), .F(
        \Reg_Bank/n3647 ) );
  MUX U615 ( .IN0(\Reg_Bank/registers[20][10] ), .IN1(n166), .SEL(n203), .F(
        \Reg_Bank/n3646 ) );
  MUX U616 ( .IN0(\Reg_Bank/registers[20][9] ), .IN1(n167), .SEL(n203), .F(
        \Reg_Bank/n3645 ) );
  MUX U617 ( .IN0(\Reg_Bank/registers[20][8] ), .IN1(n168), .SEL(n203), .F(
        \Reg_Bank/n3644 ) );
  MUX U618 ( .IN0(\Reg_Bank/registers[20][7] ), .IN1(n169), .SEL(n203), .F(
        \Reg_Bank/n3643 ) );
  MUX U619 ( .IN0(\Reg_Bank/registers[20][6] ), .IN1(n170), .SEL(n203), .F(
        \Reg_Bank/n3642 ) );
  MUX U620 ( .IN0(\Reg_Bank/registers[20][5] ), .IN1(n171), .SEL(n203), .F(
        \Reg_Bank/n3641 ) );
  MUX U621 ( .IN0(\Reg_Bank/registers[20][4] ), .IN1(n172), .SEL(n203), .F(
        \Reg_Bank/n3640 ) );
  MUX U622 ( .IN0(\Reg_Bank/registers[20][3] ), .IN1(n173), .SEL(n203), .F(
        \Reg_Bank/n3639 ) );
  MUX U623 ( .IN0(\Reg_Bank/registers[20][2] ), .IN1(n174), .SEL(n203), .F(
        \Reg_Bank/n3638 ) );
  MUX U624 ( .IN0(\Reg_Bank/registers[20][1] ), .IN1(n176), .SEL(n203), .F(
        \Reg_Bank/n3637 ) );
  MUX U625 ( .IN0(\Reg_Bank/registers[20][0] ), .IN1(n177), .SEL(n203), .F(
        \Reg_Bank/n3636 ) );
  AND U626 ( .A(n188), .B(n200), .Z(n203) );
  MUX U627 ( .IN0(\Reg_Bank/registers[19][31] ), .IN1(n144), .SEL(n204), .F(
        \Reg_Bank/n3635 ) );
  MUX U628 ( .IN0(\Reg_Bank/registers[19][30] ), .IN1(n146), .SEL(n204), .F(
        \Reg_Bank/n3634 ) );
  MUX U629 ( .IN0(\Reg_Bank/registers[19][29] ), .IN1(n147), .SEL(n204), .F(
        \Reg_Bank/n3633 ) );
  MUX U630 ( .IN0(\Reg_Bank/registers[19][28] ), .IN1(n148), .SEL(n204), .F(
        \Reg_Bank/n3632 ) );
  MUX U631 ( .IN0(\Reg_Bank/registers[19][27] ), .IN1(n149), .SEL(n204), .F(
        \Reg_Bank/n3631 ) );
  MUX U632 ( .IN0(\Reg_Bank/registers[19][26] ), .IN1(n150), .SEL(n204), .F(
        \Reg_Bank/n3630 ) );
  MUX U633 ( .IN0(\Reg_Bank/registers[19][25] ), .IN1(n151), .SEL(n204), .F(
        \Reg_Bank/n3629 ) );
  MUX U634 ( .IN0(\Reg_Bank/registers[19][24] ), .IN1(n152), .SEL(n204), .F(
        \Reg_Bank/n3628 ) );
  MUX U635 ( .IN0(\Reg_Bank/registers[19][23] ), .IN1(n153), .SEL(n204), .F(
        \Reg_Bank/n3627 ) );
  MUX U636 ( .IN0(\Reg_Bank/registers[19][22] ), .IN1(n154), .SEL(n204), .F(
        \Reg_Bank/n3626 ) );
  MUX U637 ( .IN0(\Reg_Bank/registers[19][21] ), .IN1(n155), .SEL(n204), .F(
        \Reg_Bank/n3625 ) );
  MUX U638 ( .IN0(\Reg_Bank/registers[19][20] ), .IN1(n156), .SEL(n204), .F(
        \Reg_Bank/n3624 ) );
  MUX U639 ( .IN0(\Reg_Bank/registers[19][19] ), .IN1(n157), .SEL(n204), .F(
        \Reg_Bank/n3623 ) );
  MUX U640 ( .IN0(\Reg_Bank/registers[19][18] ), .IN1(n158), .SEL(n204), .F(
        \Reg_Bank/n3622 ) );
  MUX U641 ( .IN0(\Reg_Bank/registers[19][17] ), .IN1(n159), .SEL(n204), .F(
        \Reg_Bank/n3621 ) );
  MUX U642 ( .IN0(\Reg_Bank/registers[19][16] ), .IN1(n160), .SEL(n204), .F(
        \Reg_Bank/n3620 ) );
  MUX U643 ( .IN0(\Reg_Bank/registers[19][15] ), .IN1(n161), .SEL(n204), .F(
        \Reg_Bank/n3619 ) );
  MUX U644 ( .IN0(\Reg_Bank/registers[19][14] ), .IN1(n162), .SEL(n204), .F(
        \Reg_Bank/n3618 ) );
  MUX U645 ( .IN0(\Reg_Bank/registers[19][13] ), .IN1(n163), .SEL(n204), .F(
        \Reg_Bank/n3617 ) );
  MUX U646 ( .IN0(\Reg_Bank/registers[19][12] ), .IN1(n164), .SEL(n204), .F(
        \Reg_Bank/n3616 ) );
  MUX U647 ( .IN0(\Reg_Bank/registers[19][11] ), .IN1(n165), .SEL(n204), .F(
        \Reg_Bank/n3615 ) );
  MUX U648 ( .IN0(\Reg_Bank/registers[19][10] ), .IN1(n166), .SEL(n204), .F(
        \Reg_Bank/n3614 ) );
  MUX U649 ( .IN0(\Reg_Bank/registers[19][9] ), .IN1(n167), .SEL(n204), .F(
        \Reg_Bank/n3613 ) );
  MUX U650 ( .IN0(\Reg_Bank/registers[19][8] ), .IN1(n168), .SEL(n204), .F(
        \Reg_Bank/n3612 ) );
  MUX U651 ( .IN0(\Reg_Bank/registers[19][7] ), .IN1(n169), .SEL(n204), .F(
        \Reg_Bank/n3611 ) );
  MUX U652 ( .IN0(\Reg_Bank/registers[19][6] ), .IN1(n170), .SEL(n204), .F(
        \Reg_Bank/n3610 ) );
  MUX U653 ( .IN0(\Reg_Bank/registers[19][5] ), .IN1(n171), .SEL(n204), .F(
        \Reg_Bank/n3609 ) );
  MUX U654 ( .IN0(\Reg_Bank/registers[19][4] ), .IN1(n172), .SEL(n204), .F(
        \Reg_Bank/n3608 ) );
  MUX U655 ( .IN0(\Reg_Bank/registers[19][3] ), .IN1(n173), .SEL(n204), .F(
        \Reg_Bank/n3607 ) );
  MUX U656 ( .IN0(\Reg_Bank/registers[19][2] ), .IN1(n174), .SEL(n204), .F(
        \Reg_Bank/n3606 ) );
  MUX U657 ( .IN0(\Reg_Bank/registers[19][1] ), .IN1(n176), .SEL(n204), .F(
        \Reg_Bank/n3605 ) );
  MUX U658 ( .IN0(\Reg_Bank/registers[19][0] ), .IN1(n177), .SEL(n204), .F(
        \Reg_Bank/n3604 ) );
  ANDN U659 ( .A(n200), .B(n190), .Z(n204) );
  MUX U660 ( .IN0(\Reg_Bank/registers[18][31] ), .IN1(n144), .SEL(n205), .F(
        \Reg_Bank/n3603 ) );
  MUX U661 ( .IN0(\Reg_Bank/registers[18][30] ), .IN1(n146), .SEL(n205), .F(
        \Reg_Bank/n3602 ) );
  MUX U662 ( .IN0(\Reg_Bank/registers[18][29] ), .IN1(n147), .SEL(n205), .F(
        \Reg_Bank/n3601 ) );
  MUX U663 ( .IN0(\Reg_Bank/registers[18][28] ), .IN1(n148), .SEL(n205), .F(
        \Reg_Bank/n3600 ) );
  MUX U664 ( .IN0(\Reg_Bank/registers[18][27] ), .IN1(n149), .SEL(n205), .F(
        \Reg_Bank/n3599 ) );
  MUX U665 ( .IN0(\Reg_Bank/registers[18][26] ), .IN1(n150), .SEL(n205), .F(
        \Reg_Bank/n3598 ) );
  MUX U666 ( .IN0(\Reg_Bank/registers[18][25] ), .IN1(n151), .SEL(n205), .F(
        \Reg_Bank/n3597 ) );
  MUX U667 ( .IN0(\Reg_Bank/registers[18][24] ), .IN1(n152), .SEL(n205), .F(
        \Reg_Bank/n3596 ) );
  MUX U668 ( .IN0(\Reg_Bank/registers[18][23] ), .IN1(n153), .SEL(n205), .F(
        \Reg_Bank/n3595 ) );
  MUX U669 ( .IN0(\Reg_Bank/registers[18][22] ), .IN1(n154), .SEL(n205), .F(
        \Reg_Bank/n3594 ) );
  MUX U670 ( .IN0(\Reg_Bank/registers[18][21] ), .IN1(n155), .SEL(n205), .F(
        \Reg_Bank/n3593 ) );
  MUX U671 ( .IN0(\Reg_Bank/registers[18][20] ), .IN1(n156), .SEL(n205), .F(
        \Reg_Bank/n3592 ) );
  MUX U672 ( .IN0(\Reg_Bank/registers[18][19] ), .IN1(n157), .SEL(n205), .F(
        \Reg_Bank/n3591 ) );
  MUX U673 ( .IN0(\Reg_Bank/registers[18][18] ), .IN1(n158), .SEL(n205), .F(
        \Reg_Bank/n3590 ) );
  MUX U674 ( .IN0(\Reg_Bank/registers[18][17] ), .IN1(n159), .SEL(n205), .F(
        \Reg_Bank/n3589 ) );
  MUX U675 ( .IN0(\Reg_Bank/registers[18][16] ), .IN1(n160), .SEL(n205), .F(
        \Reg_Bank/n3588 ) );
  MUX U676 ( .IN0(\Reg_Bank/registers[18][15] ), .IN1(n161), .SEL(n205), .F(
        \Reg_Bank/n3587 ) );
  MUX U677 ( .IN0(\Reg_Bank/registers[18][14] ), .IN1(n162), .SEL(n205), .F(
        \Reg_Bank/n3586 ) );
  MUX U678 ( .IN0(\Reg_Bank/registers[18][13] ), .IN1(n163), .SEL(n205), .F(
        \Reg_Bank/n3585 ) );
  MUX U679 ( .IN0(\Reg_Bank/registers[18][12] ), .IN1(n164), .SEL(n205), .F(
        \Reg_Bank/n3584 ) );
  MUX U680 ( .IN0(\Reg_Bank/registers[18][11] ), .IN1(n165), .SEL(n205), .F(
        \Reg_Bank/n3583 ) );
  MUX U681 ( .IN0(\Reg_Bank/registers[18][10] ), .IN1(n166), .SEL(n205), .F(
        \Reg_Bank/n3582 ) );
  MUX U682 ( .IN0(\Reg_Bank/registers[18][9] ), .IN1(n167), .SEL(n205), .F(
        \Reg_Bank/n3581 ) );
  MUX U683 ( .IN0(\Reg_Bank/registers[18][8] ), .IN1(n168), .SEL(n205), .F(
        \Reg_Bank/n3580 ) );
  MUX U684 ( .IN0(\Reg_Bank/registers[18][7] ), .IN1(n169), .SEL(n205), .F(
        \Reg_Bank/n3579 ) );
  MUX U685 ( .IN0(\Reg_Bank/registers[18][6] ), .IN1(n170), .SEL(n205), .F(
        \Reg_Bank/n3578 ) );
  MUX U686 ( .IN0(\Reg_Bank/registers[18][5] ), .IN1(n171), .SEL(n205), .F(
        \Reg_Bank/n3577 ) );
  MUX U687 ( .IN0(\Reg_Bank/registers[18][4] ), .IN1(n172), .SEL(n205), .F(
        \Reg_Bank/n3576 ) );
  MUX U688 ( .IN0(\Reg_Bank/registers[18][3] ), .IN1(n173), .SEL(n205), .F(
        \Reg_Bank/n3575 ) );
  MUX U689 ( .IN0(\Reg_Bank/registers[18][2] ), .IN1(n174), .SEL(n205), .F(
        \Reg_Bank/n3574 ) );
  MUX U690 ( .IN0(\Reg_Bank/registers[18][1] ), .IN1(n176), .SEL(n205), .F(
        \Reg_Bank/n3573 ) );
  MUX U691 ( .IN0(\Reg_Bank/registers[18][0] ), .IN1(n177), .SEL(n205), .F(
        \Reg_Bank/n3572 ) );
  ANDN U692 ( .A(n200), .B(n192), .Z(n205) );
  MUX U693 ( .IN0(\Reg_Bank/registers[17][31] ), .IN1(n144), .SEL(n206), .F(
        \Reg_Bank/n3571 ) );
  MUX U694 ( .IN0(\Reg_Bank/registers[17][30] ), .IN1(n146), .SEL(n206), .F(
        \Reg_Bank/n3570 ) );
  MUX U695 ( .IN0(\Reg_Bank/registers[17][29] ), .IN1(n147), .SEL(n206), .F(
        \Reg_Bank/n3569 ) );
  MUX U696 ( .IN0(\Reg_Bank/registers[17][28] ), .IN1(n148), .SEL(n206), .F(
        \Reg_Bank/n3568 ) );
  MUX U697 ( .IN0(\Reg_Bank/registers[17][27] ), .IN1(n149), .SEL(n206), .F(
        \Reg_Bank/n3567 ) );
  MUX U698 ( .IN0(\Reg_Bank/registers[17][26] ), .IN1(n150), .SEL(n206), .F(
        \Reg_Bank/n3566 ) );
  MUX U699 ( .IN0(\Reg_Bank/registers[17][25] ), .IN1(n151), .SEL(n206), .F(
        \Reg_Bank/n3565 ) );
  MUX U700 ( .IN0(\Reg_Bank/registers[17][24] ), .IN1(n152), .SEL(n206), .F(
        \Reg_Bank/n3564 ) );
  MUX U701 ( .IN0(\Reg_Bank/registers[17][23] ), .IN1(n153), .SEL(n206), .F(
        \Reg_Bank/n3563 ) );
  MUX U702 ( .IN0(\Reg_Bank/registers[17][22] ), .IN1(n154), .SEL(n206), .F(
        \Reg_Bank/n3562 ) );
  MUX U703 ( .IN0(\Reg_Bank/registers[17][21] ), .IN1(n155), .SEL(n206), .F(
        \Reg_Bank/n3561 ) );
  MUX U704 ( .IN0(\Reg_Bank/registers[17][20] ), .IN1(n156), .SEL(n206), .F(
        \Reg_Bank/n3560 ) );
  MUX U705 ( .IN0(\Reg_Bank/registers[17][19] ), .IN1(n157), .SEL(n206), .F(
        \Reg_Bank/n3559 ) );
  MUX U706 ( .IN0(\Reg_Bank/registers[17][18] ), .IN1(n158), .SEL(n206), .F(
        \Reg_Bank/n3558 ) );
  MUX U707 ( .IN0(\Reg_Bank/registers[17][17] ), .IN1(n159), .SEL(n206), .F(
        \Reg_Bank/n3557 ) );
  MUX U708 ( .IN0(\Reg_Bank/registers[17][16] ), .IN1(n160), .SEL(n206), .F(
        \Reg_Bank/n3556 ) );
  MUX U709 ( .IN0(\Reg_Bank/registers[17][15] ), .IN1(n161), .SEL(n206), .F(
        \Reg_Bank/n3555 ) );
  MUX U710 ( .IN0(\Reg_Bank/registers[17][14] ), .IN1(n162), .SEL(n206), .F(
        \Reg_Bank/n3554 ) );
  MUX U711 ( .IN0(\Reg_Bank/registers[17][13] ), .IN1(n163), .SEL(n206), .F(
        \Reg_Bank/n3553 ) );
  MUX U712 ( .IN0(\Reg_Bank/registers[17][12] ), .IN1(n164), .SEL(n206), .F(
        \Reg_Bank/n3552 ) );
  MUX U713 ( .IN0(\Reg_Bank/registers[17][11] ), .IN1(n165), .SEL(n206), .F(
        \Reg_Bank/n3551 ) );
  MUX U714 ( .IN0(\Reg_Bank/registers[17][10] ), .IN1(n166), .SEL(n206), .F(
        \Reg_Bank/n3550 ) );
  MUX U715 ( .IN0(\Reg_Bank/registers[17][9] ), .IN1(n167), .SEL(n206), .F(
        \Reg_Bank/n3549 ) );
  MUX U716 ( .IN0(\Reg_Bank/registers[17][8] ), .IN1(n168), .SEL(n206), .F(
        \Reg_Bank/n3548 ) );
  MUX U717 ( .IN0(\Reg_Bank/registers[17][7] ), .IN1(n169), .SEL(n206), .F(
        \Reg_Bank/n3547 ) );
  MUX U718 ( .IN0(\Reg_Bank/registers[17][6] ), .IN1(n170), .SEL(n206), .F(
        \Reg_Bank/n3546 ) );
  MUX U719 ( .IN0(\Reg_Bank/registers[17][5] ), .IN1(n171), .SEL(n206), .F(
        \Reg_Bank/n3545 ) );
  MUX U720 ( .IN0(\Reg_Bank/registers[17][4] ), .IN1(n172), .SEL(n206), .F(
        \Reg_Bank/n3544 ) );
  MUX U721 ( .IN0(\Reg_Bank/registers[17][3] ), .IN1(n173), .SEL(n206), .F(
        \Reg_Bank/n3543 ) );
  MUX U722 ( .IN0(\Reg_Bank/registers[17][2] ), .IN1(n174), .SEL(n206), .F(
        \Reg_Bank/n3542 ) );
  MUX U723 ( .IN0(\Reg_Bank/registers[17][1] ), .IN1(n176), .SEL(n206), .F(
        \Reg_Bank/n3541 ) );
  MUX U724 ( .IN0(\Reg_Bank/registers[17][0] ), .IN1(n177), .SEL(n206), .F(
        \Reg_Bank/n3540 ) );
  ANDN U725 ( .A(n200), .B(n194), .Z(n206) );
  MUX U726 ( .IN0(\Reg_Bank/registers[16][31] ), .IN1(n144), .SEL(n207), .F(
        \Reg_Bank/n3539 ) );
  MUX U727 ( .IN0(\Reg_Bank/registers[16][30] ), .IN1(n146), .SEL(n207), .F(
        \Reg_Bank/n3538 ) );
  MUX U728 ( .IN0(\Reg_Bank/registers[16][29] ), .IN1(n147), .SEL(n207), .F(
        \Reg_Bank/n3537 ) );
  MUX U729 ( .IN0(\Reg_Bank/registers[16][28] ), .IN1(n148), .SEL(n207), .F(
        \Reg_Bank/n3536 ) );
  MUX U730 ( .IN0(\Reg_Bank/registers[16][27] ), .IN1(n149), .SEL(n207), .F(
        \Reg_Bank/n3535 ) );
  MUX U731 ( .IN0(\Reg_Bank/registers[16][26] ), .IN1(n150), .SEL(n207), .F(
        \Reg_Bank/n3534 ) );
  MUX U732 ( .IN0(\Reg_Bank/registers[16][25] ), .IN1(n151), .SEL(n207), .F(
        \Reg_Bank/n3533 ) );
  MUX U733 ( .IN0(\Reg_Bank/registers[16][24] ), .IN1(n152), .SEL(n207), .F(
        \Reg_Bank/n3532 ) );
  MUX U734 ( .IN0(\Reg_Bank/registers[16][23] ), .IN1(n153), .SEL(n207), .F(
        \Reg_Bank/n3531 ) );
  MUX U735 ( .IN0(\Reg_Bank/registers[16][22] ), .IN1(n154), .SEL(n207), .F(
        \Reg_Bank/n3530 ) );
  MUX U736 ( .IN0(\Reg_Bank/registers[16][21] ), .IN1(n155), .SEL(n207), .F(
        \Reg_Bank/n3529 ) );
  MUX U737 ( .IN0(\Reg_Bank/registers[16][20] ), .IN1(n156), .SEL(n207), .F(
        \Reg_Bank/n3528 ) );
  MUX U738 ( .IN0(\Reg_Bank/registers[16][19] ), .IN1(n157), .SEL(n207), .F(
        \Reg_Bank/n3527 ) );
  MUX U739 ( .IN0(\Reg_Bank/registers[16][18] ), .IN1(n158), .SEL(n207), .F(
        \Reg_Bank/n3526 ) );
  MUX U740 ( .IN0(\Reg_Bank/registers[16][17] ), .IN1(n159), .SEL(n207), .F(
        \Reg_Bank/n3525 ) );
  MUX U741 ( .IN0(\Reg_Bank/registers[16][16] ), .IN1(n160), .SEL(n207), .F(
        \Reg_Bank/n3524 ) );
  MUX U742 ( .IN0(\Reg_Bank/registers[16][15] ), .IN1(n161), .SEL(n207), .F(
        \Reg_Bank/n3523 ) );
  MUX U743 ( .IN0(\Reg_Bank/registers[16][14] ), .IN1(n162), .SEL(n207), .F(
        \Reg_Bank/n3522 ) );
  MUX U744 ( .IN0(\Reg_Bank/registers[16][13] ), .IN1(n163), .SEL(n207), .F(
        \Reg_Bank/n3521 ) );
  MUX U745 ( .IN0(\Reg_Bank/registers[16][12] ), .IN1(n164), .SEL(n207), .F(
        \Reg_Bank/n3520 ) );
  MUX U746 ( .IN0(\Reg_Bank/registers[16][11] ), .IN1(n165), .SEL(n207), .F(
        \Reg_Bank/n3519 ) );
  MUX U747 ( .IN0(\Reg_Bank/registers[16][10] ), .IN1(n166), .SEL(n207), .F(
        \Reg_Bank/n3518 ) );
  MUX U748 ( .IN0(\Reg_Bank/registers[16][9] ), .IN1(n167), .SEL(n207), .F(
        \Reg_Bank/n3517 ) );
  MUX U749 ( .IN0(\Reg_Bank/registers[16][8] ), .IN1(n168), .SEL(n207), .F(
        \Reg_Bank/n3516 ) );
  MUX U750 ( .IN0(\Reg_Bank/registers[16][7] ), .IN1(n169), .SEL(n207), .F(
        \Reg_Bank/n3515 ) );
  MUX U751 ( .IN0(\Reg_Bank/registers[16][6] ), .IN1(n170), .SEL(n207), .F(
        \Reg_Bank/n3514 ) );
  MUX U752 ( .IN0(\Reg_Bank/registers[16][5] ), .IN1(n171), .SEL(n207), .F(
        \Reg_Bank/n3513 ) );
  MUX U753 ( .IN0(\Reg_Bank/registers[16][4] ), .IN1(n172), .SEL(n207), .F(
        \Reg_Bank/n3512 ) );
  MUX U754 ( .IN0(\Reg_Bank/registers[16][3] ), .IN1(n173), .SEL(n207), .F(
        \Reg_Bank/n3511 ) );
  MUX U755 ( .IN0(\Reg_Bank/registers[16][2] ), .IN1(n174), .SEL(n207), .F(
        \Reg_Bank/n3510 ) );
  MUX U756 ( .IN0(\Reg_Bank/registers[16][1] ), .IN1(n176), .SEL(n207), .F(
        \Reg_Bank/n3509 ) );
  MUX U757 ( .IN0(\Reg_Bank/registers[16][0] ), .IN1(n177), .SEL(n207), .F(
        \Reg_Bank/n3508 ) );
  ANDN U758 ( .A(n200), .B(n196), .Z(n207) );
  IV U759 ( .A(n208), .Z(n196) );
  ANDN U760 ( .A(n197), .B(n209), .Z(n200) );
  IV U761 ( .A(n198), .Z(n209) );
  MUX U762 ( .IN0(\Reg_Bank/registers[15][31] ), .IN1(n144), .SEL(n210), .F(
        \Reg_Bank/n3507 ) );
  MUX U763 ( .IN0(\Reg_Bank/registers[15][30] ), .IN1(n146), .SEL(n210), .F(
        \Reg_Bank/n3506 ) );
  MUX U764 ( .IN0(\Reg_Bank/registers[15][29] ), .IN1(n147), .SEL(n210), .F(
        \Reg_Bank/n3505 ) );
  MUX U765 ( .IN0(\Reg_Bank/registers[15][28] ), .IN1(n148), .SEL(n210), .F(
        \Reg_Bank/n3504 ) );
  MUX U766 ( .IN0(\Reg_Bank/registers[15][27] ), .IN1(n149), .SEL(n210), .F(
        \Reg_Bank/n3503 ) );
  MUX U767 ( .IN0(\Reg_Bank/registers[15][26] ), .IN1(n150), .SEL(n210), .F(
        \Reg_Bank/n3502 ) );
  MUX U768 ( .IN0(\Reg_Bank/registers[15][25] ), .IN1(n151), .SEL(n210), .F(
        \Reg_Bank/n3501 ) );
  MUX U769 ( .IN0(\Reg_Bank/registers[15][24] ), .IN1(n152), .SEL(n210), .F(
        \Reg_Bank/n3500 ) );
  MUX U770 ( .IN0(\Reg_Bank/registers[15][23] ), .IN1(n153), .SEL(n210), .F(
        \Reg_Bank/n3499 ) );
  MUX U771 ( .IN0(\Reg_Bank/registers[15][22] ), .IN1(n154), .SEL(n210), .F(
        \Reg_Bank/n3498 ) );
  MUX U772 ( .IN0(\Reg_Bank/registers[15][21] ), .IN1(n155), .SEL(n210), .F(
        \Reg_Bank/n3497 ) );
  MUX U773 ( .IN0(\Reg_Bank/registers[15][20] ), .IN1(n156), .SEL(n210), .F(
        \Reg_Bank/n3496 ) );
  MUX U774 ( .IN0(\Reg_Bank/registers[15][19] ), .IN1(n157), .SEL(n210), .F(
        \Reg_Bank/n3495 ) );
  MUX U775 ( .IN0(\Reg_Bank/registers[15][18] ), .IN1(n158), .SEL(n210), .F(
        \Reg_Bank/n3494 ) );
  MUX U776 ( .IN0(\Reg_Bank/registers[15][17] ), .IN1(n159), .SEL(n210), .F(
        \Reg_Bank/n3493 ) );
  MUX U777 ( .IN0(\Reg_Bank/registers[15][16] ), .IN1(n160), .SEL(n210), .F(
        \Reg_Bank/n3492 ) );
  MUX U778 ( .IN0(\Reg_Bank/registers[15][15] ), .IN1(n161), .SEL(n210), .F(
        \Reg_Bank/n3491 ) );
  MUX U779 ( .IN0(\Reg_Bank/registers[15][14] ), .IN1(n162), .SEL(n210), .F(
        \Reg_Bank/n3490 ) );
  MUX U780 ( .IN0(\Reg_Bank/registers[15][13] ), .IN1(n163), .SEL(n210), .F(
        \Reg_Bank/n3489 ) );
  MUX U781 ( .IN0(\Reg_Bank/registers[15][12] ), .IN1(n164), .SEL(n210), .F(
        \Reg_Bank/n3488 ) );
  MUX U782 ( .IN0(\Reg_Bank/registers[15][11] ), .IN1(n165), .SEL(n210), .F(
        \Reg_Bank/n3487 ) );
  MUX U783 ( .IN0(\Reg_Bank/registers[15][10] ), .IN1(n166), .SEL(n210), .F(
        \Reg_Bank/n3486 ) );
  MUX U784 ( .IN0(\Reg_Bank/registers[15][9] ), .IN1(n167), .SEL(n210), .F(
        \Reg_Bank/n3485 ) );
  MUX U785 ( .IN0(\Reg_Bank/registers[15][8] ), .IN1(n168), .SEL(n210), .F(
        \Reg_Bank/n3484 ) );
  MUX U786 ( .IN0(\Reg_Bank/registers[15][7] ), .IN1(n169), .SEL(n210), .F(
        \Reg_Bank/n3483 ) );
  MUX U787 ( .IN0(\Reg_Bank/registers[15][6] ), .IN1(n170), .SEL(n210), .F(
        \Reg_Bank/n3482 ) );
  MUX U788 ( .IN0(\Reg_Bank/registers[15][5] ), .IN1(n171), .SEL(n210), .F(
        \Reg_Bank/n3481 ) );
  MUX U789 ( .IN0(\Reg_Bank/registers[15][4] ), .IN1(n172), .SEL(n210), .F(
        \Reg_Bank/n3480 ) );
  MUX U790 ( .IN0(\Reg_Bank/registers[15][3] ), .IN1(n173), .SEL(n210), .F(
        \Reg_Bank/n3479 ) );
  MUX U791 ( .IN0(\Reg_Bank/registers[15][2] ), .IN1(n174), .SEL(n210), .F(
        \Reg_Bank/n3478 ) );
  IV U792 ( .A(n211), .Z(n210) );
  MUX U793 ( .IN0(n176), .IN1(\Reg_Bank/registers[15][1] ), .SEL(n211), .F(
        \Reg_Bank/n3477 ) );
  MUX U794 ( .IN0(n177), .IN1(\Reg_Bank/registers[15][0] ), .SEL(n211), .F(
        \Reg_Bank/n3476 ) );
  OR U795 ( .A(n178), .B(n212), .Z(n211) );
  MUX U796 ( .IN0(\Reg_Bank/registers[14][31] ), .IN1(n144), .SEL(n213), .F(
        \Reg_Bank/n3475 ) );
  MUX U797 ( .IN0(\Reg_Bank/registers[14][30] ), .IN1(n146), .SEL(n213), .F(
        \Reg_Bank/n3474 ) );
  MUX U798 ( .IN0(\Reg_Bank/registers[14][29] ), .IN1(n147), .SEL(n213), .F(
        \Reg_Bank/n3473 ) );
  MUX U799 ( .IN0(\Reg_Bank/registers[14][28] ), .IN1(n148), .SEL(n213), .F(
        \Reg_Bank/n3472 ) );
  MUX U800 ( .IN0(\Reg_Bank/registers[14][27] ), .IN1(n149), .SEL(n213), .F(
        \Reg_Bank/n3471 ) );
  MUX U801 ( .IN0(\Reg_Bank/registers[14][26] ), .IN1(n150), .SEL(n213), .F(
        \Reg_Bank/n3470 ) );
  MUX U802 ( .IN0(\Reg_Bank/registers[14][25] ), .IN1(n151), .SEL(n213), .F(
        \Reg_Bank/n3469 ) );
  MUX U803 ( .IN0(\Reg_Bank/registers[14][24] ), .IN1(n152), .SEL(n213), .F(
        \Reg_Bank/n3468 ) );
  MUX U804 ( .IN0(\Reg_Bank/registers[14][23] ), .IN1(n153), .SEL(n213), .F(
        \Reg_Bank/n3467 ) );
  MUX U805 ( .IN0(\Reg_Bank/registers[14][22] ), .IN1(n154), .SEL(n213), .F(
        \Reg_Bank/n3466 ) );
  MUX U806 ( .IN0(\Reg_Bank/registers[14][21] ), .IN1(n155), .SEL(n213), .F(
        \Reg_Bank/n3465 ) );
  MUX U807 ( .IN0(\Reg_Bank/registers[14][20] ), .IN1(n156), .SEL(n213), .F(
        \Reg_Bank/n3464 ) );
  MUX U808 ( .IN0(\Reg_Bank/registers[14][19] ), .IN1(n157), .SEL(n213), .F(
        \Reg_Bank/n3463 ) );
  MUX U809 ( .IN0(\Reg_Bank/registers[14][18] ), .IN1(n158), .SEL(n213), .F(
        \Reg_Bank/n3462 ) );
  MUX U810 ( .IN0(\Reg_Bank/registers[14][17] ), .IN1(n159), .SEL(n213), .F(
        \Reg_Bank/n3461 ) );
  MUX U811 ( .IN0(\Reg_Bank/registers[14][16] ), .IN1(n160), .SEL(n213), .F(
        \Reg_Bank/n3460 ) );
  MUX U812 ( .IN0(\Reg_Bank/registers[14][15] ), .IN1(n161), .SEL(n213), .F(
        \Reg_Bank/n3459 ) );
  MUX U813 ( .IN0(\Reg_Bank/registers[14][14] ), .IN1(n162), .SEL(n213), .F(
        \Reg_Bank/n3458 ) );
  MUX U814 ( .IN0(\Reg_Bank/registers[14][13] ), .IN1(n163), .SEL(n213), .F(
        \Reg_Bank/n3457 ) );
  MUX U815 ( .IN0(\Reg_Bank/registers[14][12] ), .IN1(n164), .SEL(n213), .F(
        \Reg_Bank/n3456 ) );
  MUX U816 ( .IN0(\Reg_Bank/registers[14][11] ), .IN1(n165), .SEL(n213), .F(
        \Reg_Bank/n3455 ) );
  MUX U817 ( .IN0(\Reg_Bank/registers[14][10] ), .IN1(n166), .SEL(n213), .F(
        \Reg_Bank/n3454 ) );
  MUX U818 ( .IN0(\Reg_Bank/registers[14][9] ), .IN1(n167), .SEL(n213), .F(
        \Reg_Bank/n3453 ) );
  MUX U819 ( .IN0(\Reg_Bank/registers[14][8] ), .IN1(n168), .SEL(n213), .F(
        \Reg_Bank/n3452 ) );
  MUX U820 ( .IN0(\Reg_Bank/registers[14][7] ), .IN1(n169), .SEL(n213), .F(
        \Reg_Bank/n3451 ) );
  MUX U821 ( .IN0(\Reg_Bank/registers[14][6] ), .IN1(n170), .SEL(n213), .F(
        \Reg_Bank/n3450 ) );
  MUX U822 ( .IN0(\Reg_Bank/registers[14][5] ), .IN1(n171), .SEL(n213), .F(
        \Reg_Bank/n3449 ) );
  MUX U823 ( .IN0(\Reg_Bank/registers[14][4] ), .IN1(n172), .SEL(n213), .F(
        \Reg_Bank/n3448 ) );
  MUX U824 ( .IN0(\Reg_Bank/registers[14][3] ), .IN1(n173), .SEL(n213), .F(
        \Reg_Bank/n3447 ) );
  MUX U825 ( .IN0(\Reg_Bank/registers[14][2] ), .IN1(n174), .SEL(n213), .F(
        \Reg_Bank/n3446 ) );
  MUX U826 ( .IN0(\Reg_Bank/registers[14][1] ), .IN1(n176), .SEL(n213), .F(
        \Reg_Bank/n3445 ) );
  MUX U827 ( .IN0(\Reg_Bank/registers[14][0] ), .IN1(n177), .SEL(n213), .F(
        \Reg_Bank/n3444 ) );
  ANDN U828 ( .A(n182), .B(n212), .Z(n213) );
  MUX U829 ( .IN0(\Reg_Bank/registers[13][31] ), .IN1(n144), .SEL(n214), .F(
        \Reg_Bank/n3443 ) );
  MUX U830 ( .IN0(\Reg_Bank/registers[13][30] ), .IN1(n146), .SEL(n214), .F(
        \Reg_Bank/n3442 ) );
  MUX U831 ( .IN0(\Reg_Bank/registers[13][29] ), .IN1(n147), .SEL(n214), .F(
        \Reg_Bank/n3441 ) );
  MUX U832 ( .IN0(\Reg_Bank/registers[13][28] ), .IN1(n148), .SEL(n214), .F(
        \Reg_Bank/n3440 ) );
  MUX U833 ( .IN0(\Reg_Bank/registers[13][27] ), .IN1(n149), .SEL(n214), .F(
        \Reg_Bank/n3439 ) );
  MUX U834 ( .IN0(\Reg_Bank/registers[13][26] ), .IN1(n150), .SEL(n214), .F(
        \Reg_Bank/n3438 ) );
  MUX U835 ( .IN0(\Reg_Bank/registers[13][25] ), .IN1(n151), .SEL(n214), .F(
        \Reg_Bank/n3437 ) );
  MUX U836 ( .IN0(\Reg_Bank/registers[13][24] ), .IN1(n152), .SEL(n214), .F(
        \Reg_Bank/n3436 ) );
  MUX U837 ( .IN0(\Reg_Bank/registers[13][23] ), .IN1(n153), .SEL(n214), .F(
        \Reg_Bank/n3435 ) );
  MUX U838 ( .IN0(\Reg_Bank/registers[13][22] ), .IN1(n154), .SEL(n214), .F(
        \Reg_Bank/n3434 ) );
  MUX U839 ( .IN0(\Reg_Bank/registers[13][21] ), .IN1(n155), .SEL(n214), .F(
        \Reg_Bank/n3433 ) );
  MUX U840 ( .IN0(\Reg_Bank/registers[13][20] ), .IN1(n156), .SEL(n214), .F(
        \Reg_Bank/n3432 ) );
  MUX U841 ( .IN0(\Reg_Bank/registers[13][19] ), .IN1(n157), .SEL(n214), .F(
        \Reg_Bank/n3431 ) );
  MUX U842 ( .IN0(\Reg_Bank/registers[13][18] ), .IN1(n158), .SEL(n214), .F(
        \Reg_Bank/n3430 ) );
  MUX U843 ( .IN0(\Reg_Bank/registers[13][17] ), .IN1(n159), .SEL(n214), .F(
        \Reg_Bank/n3429 ) );
  MUX U844 ( .IN0(\Reg_Bank/registers[13][16] ), .IN1(n160), .SEL(n214), .F(
        \Reg_Bank/n3428 ) );
  MUX U845 ( .IN0(\Reg_Bank/registers[13][15] ), .IN1(n161), .SEL(n214), .F(
        \Reg_Bank/n3427 ) );
  MUX U846 ( .IN0(\Reg_Bank/registers[13][14] ), .IN1(n162), .SEL(n214), .F(
        \Reg_Bank/n3426 ) );
  MUX U847 ( .IN0(\Reg_Bank/registers[13][13] ), .IN1(n163), .SEL(n214), .F(
        \Reg_Bank/n3425 ) );
  MUX U848 ( .IN0(\Reg_Bank/registers[13][12] ), .IN1(n164), .SEL(n214), .F(
        \Reg_Bank/n3424 ) );
  MUX U849 ( .IN0(\Reg_Bank/registers[13][11] ), .IN1(n165), .SEL(n214), .F(
        \Reg_Bank/n3423 ) );
  MUX U850 ( .IN0(\Reg_Bank/registers[13][10] ), .IN1(n166), .SEL(n214), .F(
        \Reg_Bank/n3422 ) );
  MUX U851 ( .IN0(\Reg_Bank/registers[13][9] ), .IN1(n167), .SEL(n214), .F(
        \Reg_Bank/n3421 ) );
  MUX U852 ( .IN0(\Reg_Bank/registers[13][8] ), .IN1(n168), .SEL(n214), .F(
        \Reg_Bank/n3420 ) );
  MUX U853 ( .IN0(\Reg_Bank/registers[13][7] ), .IN1(n169), .SEL(n214), .F(
        \Reg_Bank/n3419 ) );
  MUX U854 ( .IN0(\Reg_Bank/registers[13][6] ), .IN1(n170), .SEL(n214), .F(
        \Reg_Bank/n3418 ) );
  MUX U855 ( .IN0(\Reg_Bank/registers[13][5] ), .IN1(n171), .SEL(n214), .F(
        \Reg_Bank/n3417 ) );
  MUX U856 ( .IN0(\Reg_Bank/registers[13][4] ), .IN1(n172), .SEL(n214), .F(
        \Reg_Bank/n3416 ) );
  MUX U857 ( .IN0(\Reg_Bank/registers[13][3] ), .IN1(n173), .SEL(n214), .F(
        \Reg_Bank/n3415 ) );
  MUX U858 ( .IN0(\Reg_Bank/registers[13][2] ), .IN1(n174), .SEL(n214), .F(
        \Reg_Bank/n3414 ) );
  MUX U859 ( .IN0(\Reg_Bank/registers[13][1] ), .IN1(n176), .SEL(n214), .F(
        \Reg_Bank/n3413 ) );
  MUX U860 ( .IN0(\Reg_Bank/registers[13][0] ), .IN1(n177), .SEL(n214), .F(
        \Reg_Bank/n3412 ) );
  ANDN U861 ( .A(n185), .B(n212), .Z(n214) );
  MUX U862 ( .IN0(\Reg_Bank/registers[12][31] ), .IN1(n144), .SEL(n215), .F(
        \Reg_Bank/n3411 ) );
  MUX U863 ( .IN0(\Reg_Bank/registers[12][30] ), .IN1(n146), .SEL(n215), .F(
        \Reg_Bank/n3410 ) );
  MUX U864 ( .IN0(\Reg_Bank/registers[12][29] ), .IN1(n147), .SEL(n215), .F(
        \Reg_Bank/n3409 ) );
  MUX U865 ( .IN0(\Reg_Bank/registers[12][28] ), .IN1(n148), .SEL(n215), .F(
        \Reg_Bank/n3408 ) );
  MUX U866 ( .IN0(\Reg_Bank/registers[12][27] ), .IN1(n149), .SEL(n215), .F(
        \Reg_Bank/n3407 ) );
  MUX U867 ( .IN0(\Reg_Bank/registers[12][26] ), .IN1(n150), .SEL(n215), .F(
        \Reg_Bank/n3406 ) );
  MUX U868 ( .IN0(\Reg_Bank/registers[12][25] ), .IN1(n151), .SEL(n215), .F(
        \Reg_Bank/n3405 ) );
  MUX U869 ( .IN0(\Reg_Bank/registers[12][24] ), .IN1(n152), .SEL(n215), .F(
        \Reg_Bank/n3404 ) );
  MUX U870 ( .IN0(\Reg_Bank/registers[12][23] ), .IN1(n153), .SEL(n215), .F(
        \Reg_Bank/n3403 ) );
  MUX U871 ( .IN0(\Reg_Bank/registers[12][22] ), .IN1(n154), .SEL(n215), .F(
        \Reg_Bank/n3402 ) );
  MUX U872 ( .IN0(\Reg_Bank/registers[12][21] ), .IN1(n155), .SEL(n215), .F(
        \Reg_Bank/n3401 ) );
  MUX U873 ( .IN0(\Reg_Bank/registers[12][20] ), .IN1(n156), .SEL(n215), .F(
        \Reg_Bank/n3400 ) );
  MUX U874 ( .IN0(\Reg_Bank/registers[12][19] ), .IN1(n157), .SEL(n215), .F(
        \Reg_Bank/n3399 ) );
  MUX U875 ( .IN0(\Reg_Bank/registers[12][18] ), .IN1(n158), .SEL(n215), .F(
        \Reg_Bank/n3398 ) );
  MUX U876 ( .IN0(\Reg_Bank/registers[12][17] ), .IN1(n159), .SEL(n215), .F(
        \Reg_Bank/n3397 ) );
  MUX U877 ( .IN0(\Reg_Bank/registers[12][16] ), .IN1(n160), .SEL(n215), .F(
        \Reg_Bank/n3396 ) );
  MUX U878 ( .IN0(\Reg_Bank/registers[12][15] ), .IN1(n161), .SEL(n215), .F(
        \Reg_Bank/n3395 ) );
  MUX U879 ( .IN0(\Reg_Bank/registers[12][14] ), .IN1(n162), .SEL(n215), .F(
        \Reg_Bank/n3394 ) );
  MUX U880 ( .IN0(\Reg_Bank/registers[12][13] ), .IN1(n163), .SEL(n215), .F(
        \Reg_Bank/n3393 ) );
  MUX U881 ( .IN0(\Reg_Bank/registers[12][12] ), .IN1(n164), .SEL(n215), .F(
        \Reg_Bank/n3392 ) );
  MUX U882 ( .IN0(\Reg_Bank/registers[12][11] ), .IN1(n165), .SEL(n215), .F(
        \Reg_Bank/n3391 ) );
  MUX U883 ( .IN0(\Reg_Bank/registers[12][10] ), .IN1(n166), .SEL(n215), .F(
        \Reg_Bank/n3390 ) );
  MUX U884 ( .IN0(\Reg_Bank/registers[12][9] ), .IN1(n167), .SEL(n215), .F(
        \Reg_Bank/n3389 ) );
  MUX U885 ( .IN0(\Reg_Bank/registers[12][8] ), .IN1(n168), .SEL(n215), .F(
        \Reg_Bank/n3388 ) );
  MUX U886 ( .IN0(\Reg_Bank/registers[12][7] ), .IN1(n169), .SEL(n215), .F(
        \Reg_Bank/n3387 ) );
  MUX U887 ( .IN0(\Reg_Bank/registers[12][6] ), .IN1(n170), .SEL(n215), .F(
        \Reg_Bank/n3386 ) );
  MUX U888 ( .IN0(\Reg_Bank/registers[12][5] ), .IN1(n171), .SEL(n215), .F(
        \Reg_Bank/n3385 ) );
  MUX U889 ( .IN0(\Reg_Bank/registers[12][4] ), .IN1(n172), .SEL(n215), .F(
        \Reg_Bank/n3384 ) );
  MUX U890 ( .IN0(\Reg_Bank/registers[12][3] ), .IN1(n173), .SEL(n215), .F(
        \Reg_Bank/n3383 ) );
  MUX U891 ( .IN0(\Reg_Bank/registers[12][2] ), .IN1(n174), .SEL(n215), .F(
        \Reg_Bank/n3382 ) );
  MUX U892 ( .IN0(\Reg_Bank/registers[12][1] ), .IN1(n176), .SEL(n215), .F(
        \Reg_Bank/n3381 ) );
  MUX U893 ( .IN0(\Reg_Bank/registers[12][0] ), .IN1(n177), .SEL(n215), .F(
        \Reg_Bank/n3380 ) );
  ANDN U894 ( .A(n188), .B(n212), .Z(n215) );
  MUX U895 ( .IN0(\Reg_Bank/registers[11][31] ), .IN1(n144), .SEL(n216), .F(
        \Reg_Bank/n3379 ) );
  MUX U896 ( .IN0(\Reg_Bank/registers[11][30] ), .IN1(n146), .SEL(n216), .F(
        \Reg_Bank/n3378 ) );
  MUX U897 ( .IN0(\Reg_Bank/registers[11][29] ), .IN1(n147), .SEL(n216), .F(
        \Reg_Bank/n3377 ) );
  MUX U898 ( .IN0(\Reg_Bank/registers[11][28] ), .IN1(n148), .SEL(n216), .F(
        \Reg_Bank/n3376 ) );
  MUX U899 ( .IN0(\Reg_Bank/registers[11][27] ), .IN1(n149), .SEL(n216), .F(
        \Reg_Bank/n3375 ) );
  MUX U900 ( .IN0(\Reg_Bank/registers[11][26] ), .IN1(n150), .SEL(n216), .F(
        \Reg_Bank/n3374 ) );
  MUX U901 ( .IN0(\Reg_Bank/registers[11][25] ), .IN1(n151), .SEL(n216), .F(
        \Reg_Bank/n3373 ) );
  MUX U902 ( .IN0(\Reg_Bank/registers[11][24] ), .IN1(n152), .SEL(n216), .F(
        \Reg_Bank/n3372 ) );
  MUX U903 ( .IN0(\Reg_Bank/registers[11][23] ), .IN1(n153), .SEL(n216), .F(
        \Reg_Bank/n3371 ) );
  MUX U904 ( .IN0(\Reg_Bank/registers[11][22] ), .IN1(n154), .SEL(n216), .F(
        \Reg_Bank/n3370 ) );
  MUX U905 ( .IN0(\Reg_Bank/registers[11][21] ), .IN1(n155), .SEL(n216), .F(
        \Reg_Bank/n3369 ) );
  MUX U906 ( .IN0(\Reg_Bank/registers[11][20] ), .IN1(n156), .SEL(n216), .F(
        \Reg_Bank/n3368 ) );
  MUX U907 ( .IN0(\Reg_Bank/registers[11][19] ), .IN1(n157), .SEL(n216), .F(
        \Reg_Bank/n3367 ) );
  MUX U908 ( .IN0(\Reg_Bank/registers[11][18] ), .IN1(n158), .SEL(n216), .F(
        \Reg_Bank/n3366 ) );
  MUX U909 ( .IN0(\Reg_Bank/registers[11][17] ), .IN1(n159), .SEL(n216), .F(
        \Reg_Bank/n3365 ) );
  MUX U910 ( .IN0(\Reg_Bank/registers[11][16] ), .IN1(n160), .SEL(n216), .F(
        \Reg_Bank/n3364 ) );
  MUX U911 ( .IN0(\Reg_Bank/registers[11][15] ), .IN1(n161), .SEL(n216), .F(
        \Reg_Bank/n3363 ) );
  MUX U912 ( .IN0(\Reg_Bank/registers[11][14] ), .IN1(n162), .SEL(n216), .F(
        \Reg_Bank/n3362 ) );
  MUX U913 ( .IN0(\Reg_Bank/registers[11][13] ), .IN1(n163), .SEL(n216), .F(
        \Reg_Bank/n3361 ) );
  MUX U914 ( .IN0(\Reg_Bank/registers[11][12] ), .IN1(n164), .SEL(n216), .F(
        \Reg_Bank/n3360 ) );
  MUX U915 ( .IN0(\Reg_Bank/registers[11][11] ), .IN1(n165), .SEL(n216), .F(
        \Reg_Bank/n3359 ) );
  MUX U916 ( .IN0(\Reg_Bank/registers[11][10] ), .IN1(n166), .SEL(n216), .F(
        \Reg_Bank/n3358 ) );
  MUX U917 ( .IN0(\Reg_Bank/registers[11][9] ), .IN1(n167), .SEL(n216), .F(
        \Reg_Bank/n3357 ) );
  MUX U918 ( .IN0(\Reg_Bank/registers[11][8] ), .IN1(n168), .SEL(n216), .F(
        \Reg_Bank/n3356 ) );
  MUX U919 ( .IN0(\Reg_Bank/registers[11][7] ), .IN1(n169), .SEL(n216), .F(
        \Reg_Bank/n3355 ) );
  MUX U920 ( .IN0(\Reg_Bank/registers[11][6] ), .IN1(n170), .SEL(n216), .F(
        \Reg_Bank/n3354 ) );
  MUX U921 ( .IN0(\Reg_Bank/registers[11][5] ), .IN1(n171), .SEL(n216), .F(
        \Reg_Bank/n3353 ) );
  MUX U922 ( .IN0(\Reg_Bank/registers[11][4] ), .IN1(n172), .SEL(n216), .F(
        \Reg_Bank/n3352 ) );
  MUX U923 ( .IN0(\Reg_Bank/registers[11][3] ), .IN1(n173), .SEL(n216), .F(
        \Reg_Bank/n3351 ) );
  MUX U924 ( .IN0(\Reg_Bank/registers[11][2] ), .IN1(n174), .SEL(n216), .F(
        \Reg_Bank/n3350 ) );
  MUX U925 ( .IN0(\Reg_Bank/registers[11][1] ), .IN1(n176), .SEL(n216), .F(
        \Reg_Bank/n3349 ) );
  MUX U926 ( .IN0(\Reg_Bank/registers[11][0] ), .IN1(n177), .SEL(n216), .F(
        \Reg_Bank/n3348 ) );
  ANDN U927 ( .A(n217), .B(n212), .Z(n216) );
  MUX U928 ( .IN0(\Reg_Bank/registers[10][31] ), .IN1(n144), .SEL(n218), .F(
        \Reg_Bank/n3347 ) );
  MUX U929 ( .IN0(\Reg_Bank/registers[10][30] ), .IN1(n146), .SEL(n218), .F(
        \Reg_Bank/n3346 ) );
  MUX U930 ( .IN0(\Reg_Bank/registers[10][29] ), .IN1(n147), .SEL(n218), .F(
        \Reg_Bank/n3345 ) );
  MUX U931 ( .IN0(\Reg_Bank/registers[10][28] ), .IN1(n148), .SEL(n218), .F(
        \Reg_Bank/n3344 ) );
  MUX U932 ( .IN0(\Reg_Bank/registers[10][27] ), .IN1(n149), .SEL(n218), .F(
        \Reg_Bank/n3343 ) );
  MUX U933 ( .IN0(\Reg_Bank/registers[10][26] ), .IN1(n150), .SEL(n218), .F(
        \Reg_Bank/n3342 ) );
  MUX U934 ( .IN0(\Reg_Bank/registers[10][25] ), .IN1(n151), .SEL(n218), .F(
        \Reg_Bank/n3341 ) );
  MUX U935 ( .IN0(\Reg_Bank/registers[10][24] ), .IN1(n152), .SEL(n218), .F(
        \Reg_Bank/n3340 ) );
  MUX U936 ( .IN0(\Reg_Bank/registers[10][23] ), .IN1(n153), .SEL(n218), .F(
        \Reg_Bank/n3339 ) );
  MUX U937 ( .IN0(\Reg_Bank/registers[10][22] ), .IN1(n154), .SEL(n218), .F(
        \Reg_Bank/n3338 ) );
  MUX U938 ( .IN0(\Reg_Bank/registers[10][21] ), .IN1(n155), .SEL(n218), .F(
        \Reg_Bank/n3337 ) );
  MUX U939 ( .IN0(\Reg_Bank/registers[10][20] ), .IN1(n156), .SEL(n218), .F(
        \Reg_Bank/n3336 ) );
  MUX U940 ( .IN0(\Reg_Bank/registers[10][19] ), .IN1(n157), .SEL(n218), .F(
        \Reg_Bank/n3335 ) );
  MUX U941 ( .IN0(\Reg_Bank/registers[10][18] ), .IN1(n158), .SEL(n218), .F(
        \Reg_Bank/n3334 ) );
  MUX U942 ( .IN0(\Reg_Bank/registers[10][17] ), .IN1(n159), .SEL(n218), .F(
        \Reg_Bank/n3333 ) );
  MUX U943 ( .IN0(\Reg_Bank/registers[10][16] ), .IN1(n160), .SEL(n218), .F(
        \Reg_Bank/n3332 ) );
  MUX U944 ( .IN0(\Reg_Bank/registers[10][15] ), .IN1(n161), .SEL(n218), .F(
        \Reg_Bank/n3331 ) );
  MUX U945 ( .IN0(\Reg_Bank/registers[10][14] ), .IN1(n162), .SEL(n218), .F(
        \Reg_Bank/n3330 ) );
  MUX U946 ( .IN0(\Reg_Bank/registers[10][13] ), .IN1(n163), .SEL(n218), .F(
        \Reg_Bank/n3329 ) );
  MUX U947 ( .IN0(\Reg_Bank/registers[10][12] ), .IN1(n164), .SEL(n218), .F(
        \Reg_Bank/n3328 ) );
  MUX U948 ( .IN0(\Reg_Bank/registers[10][11] ), .IN1(n165), .SEL(n218), .F(
        \Reg_Bank/n3327 ) );
  MUX U949 ( .IN0(\Reg_Bank/registers[10][10] ), .IN1(n166), .SEL(n218), .F(
        \Reg_Bank/n3326 ) );
  MUX U950 ( .IN0(\Reg_Bank/registers[10][9] ), .IN1(n167), .SEL(n218), .F(
        \Reg_Bank/n3325 ) );
  MUX U951 ( .IN0(\Reg_Bank/registers[10][8] ), .IN1(n168), .SEL(n218), .F(
        \Reg_Bank/n3324 ) );
  MUX U952 ( .IN0(\Reg_Bank/registers[10][7] ), .IN1(n169), .SEL(n218), .F(
        \Reg_Bank/n3323 ) );
  MUX U953 ( .IN0(\Reg_Bank/registers[10][6] ), .IN1(n170), .SEL(n218), .F(
        \Reg_Bank/n3322 ) );
  MUX U954 ( .IN0(\Reg_Bank/registers[10][5] ), .IN1(n171), .SEL(n218), .F(
        \Reg_Bank/n3321 ) );
  MUX U955 ( .IN0(\Reg_Bank/registers[10][4] ), .IN1(n172), .SEL(n218), .F(
        \Reg_Bank/n3320 ) );
  MUX U956 ( .IN0(\Reg_Bank/registers[10][3] ), .IN1(n173), .SEL(n218), .F(
        \Reg_Bank/n3319 ) );
  MUX U957 ( .IN0(\Reg_Bank/registers[10][2] ), .IN1(n174), .SEL(n218), .F(
        \Reg_Bank/n3318 ) );
  MUX U958 ( .IN0(\Reg_Bank/registers[10][1] ), .IN1(n176), .SEL(n218), .F(
        \Reg_Bank/n3317 ) );
  MUX U959 ( .IN0(\Reg_Bank/registers[10][0] ), .IN1(n177), .SEL(n218), .F(
        \Reg_Bank/n3316 ) );
  ANDN U960 ( .A(n219), .B(n212), .Z(n218) );
  MUX U961 ( .IN0(\Reg_Bank/registers[9][31] ), .IN1(n144), .SEL(n220), .F(
        \Reg_Bank/n3315 ) );
  MUX U962 ( .IN0(\Reg_Bank/registers[9][30] ), .IN1(n146), .SEL(n220), .F(
        \Reg_Bank/n3314 ) );
  MUX U963 ( .IN0(\Reg_Bank/registers[9][29] ), .IN1(n147), .SEL(n220), .F(
        \Reg_Bank/n3313 ) );
  MUX U964 ( .IN0(\Reg_Bank/registers[9][28] ), .IN1(n148), .SEL(n220), .F(
        \Reg_Bank/n3312 ) );
  MUX U965 ( .IN0(\Reg_Bank/registers[9][27] ), .IN1(n149), .SEL(n220), .F(
        \Reg_Bank/n3311 ) );
  MUX U966 ( .IN0(\Reg_Bank/registers[9][26] ), .IN1(n150), .SEL(n220), .F(
        \Reg_Bank/n3310 ) );
  MUX U967 ( .IN0(\Reg_Bank/registers[9][25] ), .IN1(n151), .SEL(n220), .F(
        \Reg_Bank/n3309 ) );
  MUX U968 ( .IN0(\Reg_Bank/registers[9][24] ), .IN1(n152), .SEL(n220), .F(
        \Reg_Bank/n3308 ) );
  MUX U969 ( .IN0(\Reg_Bank/registers[9][23] ), .IN1(n153), .SEL(n220), .F(
        \Reg_Bank/n3307 ) );
  MUX U970 ( .IN0(\Reg_Bank/registers[9][22] ), .IN1(n154), .SEL(n220), .F(
        \Reg_Bank/n3306 ) );
  MUX U971 ( .IN0(\Reg_Bank/registers[9][21] ), .IN1(n155), .SEL(n220), .F(
        \Reg_Bank/n3305 ) );
  MUX U972 ( .IN0(\Reg_Bank/registers[9][20] ), .IN1(n156), .SEL(n220), .F(
        \Reg_Bank/n3304 ) );
  MUX U973 ( .IN0(\Reg_Bank/registers[9][19] ), .IN1(n157), .SEL(n220), .F(
        \Reg_Bank/n3303 ) );
  MUX U974 ( .IN0(\Reg_Bank/registers[9][18] ), .IN1(n158), .SEL(n220), .F(
        \Reg_Bank/n3302 ) );
  MUX U975 ( .IN0(\Reg_Bank/registers[9][17] ), .IN1(n159), .SEL(n220), .F(
        \Reg_Bank/n3301 ) );
  MUX U976 ( .IN0(\Reg_Bank/registers[9][16] ), .IN1(n160), .SEL(n220), .F(
        \Reg_Bank/n3300 ) );
  MUX U977 ( .IN0(\Reg_Bank/registers[9][15] ), .IN1(n161), .SEL(n220), .F(
        \Reg_Bank/n3299 ) );
  MUX U978 ( .IN0(\Reg_Bank/registers[9][14] ), .IN1(n162), .SEL(n220), .F(
        \Reg_Bank/n3298 ) );
  MUX U979 ( .IN0(\Reg_Bank/registers[9][13] ), .IN1(n163), .SEL(n220), .F(
        \Reg_Bank/n3297 ) );
  MUX U980 ( .IN0(\Reg_Bank/registers[9][12] ), .IN1(n164), .SEL(n220), .F(
        \Reg_Bank/n3296 ) );
  MUX U981 ( .IN0(\Reg_Bank/registers[9][11] ), .IN1(n165), .SEL(n220), .F(
        \Reg_Bank/n3295 ) );
  MUX U982 ( .IN0(\Reg_Bank/registers[9][10] ), .IN1(n166), .SEL(n220), .F(
        \Reg_Bank/n3294 ) );
  MUX U983 ( .IN0(\Reg_Bank/registers[9][9] ), .IN1(n167), .SEL(n220), .F(
        \Reg_Bank/n3293 ) );
  MUX U984 ( .IN0(\Reg_Bank/registers[9][8] ), .IN1(n168), .SEL(n220), .F(
        \Reg_Bank/n3292 ) );
  MUX U985 ( .IN0(\Reg_Bank/registers[9][7] ), .IN1(n169), .SEL(n220), .F(
        \Reg_Bank/n3291 ) );
  MUX U986 ( .IN0(\Reg_Bank/registers[9][6] ), .IN1(n170), .SEL(n220), .F(
        \Reg_Bank/n3290 ) );
  MUX U987 ( .IN0(\Reg_Bank/registers[9][5] ), .IN1(n171), .SEL(n220), .F(
        \Reg_Bank/n3289 ) );
  MUX U988 ( .IN0(\Reg_Bank/registers[9][4] ), .IN1(n172), .SEL(n220), .F(
        \Reg_Bank/n3288 ) );
  MUX U989 ( .IN0(\Reg_Bank/registers[9][3] ), .IN1(n173), .SEL(n220), .F(
        \Reg_Bank/n3287 ) );
  MUX U990 ( .IN0(\Reg_Bank/registers[9][2] ), .IN1(n174), .SEL(n220), .F(
        \Reg_Bank/n3286 ) );
  MUX U991 ( .IN0(\Reg_Bank/registers[9][1] ), .IN1(n176), .SEL(n220), .F(
        \Reg_Bank/n3285 ) );
  MUX U992 ( .IN0(\Reg_Bank/registers[9][0] ), .IN1(n177), .SEL(n220), .F(
        \Reg_Bank/n3284 ) );
  ANDN U993 ( .A(n221), .B(n212), .Z(n220) );
  MUX U994 ( .IN0(\Reg_Bank/registers[8][31] ), .IN1(n144), .SEL(n222), .F(
        \Reg_Bank/n3283 ) );
  MUX U995 ( .IN0(\Reg_Bank/registers[8][30] ), .IN1(n146), .SEL(n222), .F(
        \Reg_Bank/n3282 ) );
  MUX U996 ( .IN0(\Reg_Bank/registers[8][29] ), .IN1(n147), .SEL(n222), .F(
        \Reg_Bank/n3281 ) );
  MUX U997 ( .IN0(\Reg_Bank/registers[8][28] ), .IN1(n148), .SEL(n222), .F(
        \Reg_Bank/n3280 ) );
  MUX U998 ( .IN0(\Reg_Bank/registers[8][27] ), .IN1(n149), .SEL(n222), .F(
        \Reg_Bank/n3279 ) );
  MUX U999 ( .IN0(\Reg_Bank/registers[8][26] ), .IN1(n150), .SEL(n222), .F(
        \Reg_Bank/n3278 ) );
  MUX U1000 ( .IN0(\Reg_Bank/registers[8][25] ), .IN1(n151), .SEL(n222), .F(
        \Reg_Bank/n3277 ) );
  MUX U1001 ( .IN0(\Reg_Bank/registers[8][24] ), .IN1(n152), .SEL(n222), .F(
        \Reg_Bank/n3276 ) );
  MUX U1002 ( .IN0(\Reg_Bank/registers[8][23] ), .IN1(n153), .SEL(n222), .F(
        \Reg_Bank/n3275 ) );
  MUX U1003 ( .IN0(\Reg_Bank/registers[8][22] ), .IN1(n154), .SEL(n222), .F(
        \Reg_Bank/n3274 ) );
  MUX U1004 ( .IN0(\Reg_Bank/registers[8][21] ), .IN1(n155), .SEL(n222), .F(
        \Reg_Bank/n3273 ) );
  MUX U1005 ( .IN0(\Reg_Bank/registers[8][20] ), .IN1(n156), .SEL(n222), .F(
        \Reg_Bank/n3272 ) );
  MUX U1006 ( .IN0(\Reg_Bank/registers[8][19] ), .IN1(n157), .SEL(n222), .F(
        \Reg_Bank/n3271 ) );
  MUX U1007 ( .IN0(\Reg_Bank/registers[8][18] ), .IN1(n158), .SEL(n222), .F(
        \Reg_Bank/n3270 ) );
  MUX U1008 ( .IN0(\Reg_Bank/registers[8][17] ), .IN1(n159), .SEL(n222), .F(
        \Reg_Bank/n3269 ) );
  MUX U1009 ( .IN0(\Reg_Bank/registers[8][16] ), .IN1(n160), .SEL(n222), .F(
        \Reg_Bank/n3268 ) );
  MUX U1010 ( .IN0(\Reg_Bank/registers[8][15] ), .IN1(n161), .SEL(n222), .F(
        \Reg_Bank/n3267 ) );
  MUX U1011 ( .IN0(\Reg_Bank/registers[8][14] ), .IN1(n162), .SEL(n222), .F(
        \Reg_Bank/n3266 ) );
  MUX U1012 ( .IN0(\Reg_Bank/registers[8][13] ), .IN1(n163), .SEL(n222), .F(
        \Reg_Bank/n3265 ) );
  MUX U1013 ( .IN0(\Reg_Bank/registers[8][12] ), .IN1(n164), .SEL(n222), .F(
        \Reg_Bank/n3264 ) );
  MUX U1014 ( .IN0(\Reg_Bank/registers[8][11] ), .IN1(n165), .SEL(n222), .F(
        \Reg_Bank/n3263 ) );
  MUX U1015 ( .IN0(\Reg_Bank/registers[8][10] ), .IN1(n166), .SEL(n222), .F(
        \Reg_Bank/n3262 ) );
  MUX U1016 ( .IN0(\Reg_Bank/registers[8][9] ), .IN1(n167), .SEL(n222), .F(
        \Reg_Bank/n3261 ) );
  MUX U1017 ( .IN0(\Reg_Bank/registers[8][8] ), .IN1(n168), .SEL(n222), .F(
        \Reg_Bank/n3260 ) );
  MUX U1018 ( .IN0(\Reg_Bank/registers[8][7] ), .IN1(n169), .SEL(n222), .F(
        \Reg_Bank/n3259 ) );
  MUX U1019 ( .IN0(\Reg_Bank/registers[8][6] ), .IN1(n170), .SEL(n222), .F(
        \Reg_Bank/n3258 ) );
  MUX U1020 ( .IN0(\Reg_Bank/registers[8][5] ), .IN1(n171), .SEL(n222), .F(
        \Reg_Bank/n3257 ) );
  MUX U1021 ( .IN0(\Reg_Bank/registers[8][4] ), .IN1(n172), .SEL(n222), .F(
        \Reg_Bank/n3256 ) );
  MUX U1022 ( .IN0(\Reg_Bank/registers[8][3] ), .IN1(n173), .SEL(n222), .F(
        \Reg_Bank/n3255 ) );
  MUX U1023 ( .IN0(\Reg_Bank/registers[8][2] ), .IN1(n174), .SEL(n222), .F(
        \Reg_Bank/n3254 ) );
  MUX U1024 ( .IN0(\Reg_Bank/registers[8][1] ), .IN1(n176), .SEL(n222), .F(
        \Reg_Bank/n3253 ) );
  MUX U1025 ( .IN0(\Reg_Bank/registers[8][0] ), .IN1(n177), .SEL(n222), .F(
        \Reg_Bank/n3252 ) );
  ANDN U1026 ( .A(n208), .B(n212), .Z(n222) );
  OR U1027 ( .A(n197), .B(n198), .Z(n212) );
  ANDN U1028 ( .A(n223), .B(n224), .Z(n208) );
  MUX U1029 ( .IN0(\Reg_Bank/registers[7][31] ), .IN1(n144), .SEL(n225), .F(
        \Reg_Bank/n3251 ) );
  MUX U1030 ( .IN0(\Reg_Bank/registers[7][30] ), .IN1(n146), .SEL(n225), .F(
        \Reg_Bank/n3250 ) );
  MUX U1031 ( .IN0(\Reg_Bank/registers[7][29] ), .IN1(n147), .SEL(n225), .F(
        \Reg_Bank/n3249 ) );
  MUX U1032 ( .IN0(\Reg_Bank/registers[7][28] ), .IN1(n148), .SEL(n225), .F(
        \Reg_Bank/n3248 ) );
  MUX U1033 ( .IN0(\Reg_Bank/registers[7][27] ), .IN1(n149), .SEL(n225), .F(
        \Reg_Bank/n3247 ) );
  MUX U1034 ( .IN0(\Reg_Bank/registers[7][26] ), .IN1(n150), .SEL(n225), .F(
        \Reg_Bank/n3246 ) );
  MUX U1035 ( .IN0(\Reg_Bank/registers[7][25] ), .IN1(n151), .SEL(n225), .F(
        \Reg_Bank/n3245 ) );
  MUX U1036 ( .IN0(\Reg_Bank/registers[7][24] ), .IN1(n152), .SEL(n225), .F(
        \Reg_Bank/n3244 ) );
  MUX U1037 ( .IN0(\Reg_Bank/registers[7][23] ), .IN1(n153), .SEL(n225), .F(
        \Reg_Bank/n3243 ) );
  MUX U1038 ( .IN0(\Reg_Bank/registers[7][22] ), .IN1(n154), .SEL(n225), .F(
        \Reg_Bank/n3242 ) );
  MUX U1039 ( .IN0(\Reg_Bank/registers[7][21] ), .IN1(n155), .SEL(n225), .F(
        \Reg_Bank/n3241 ) );
  MUX U1040 ( .IN0(\Reg_Bank/registers[7][20] ), .IN1(n156), .SEL(n225), .F(
        \Reg_Bank/n3240 ) );
  MUX U1041 ( .IN0(\Reg_Bank/registers[7][19] ), .IN1(n157), .SEL(n225), .F(
        \Reg_Bank/n3239 ) );
  MUX U1042 ( .IN0(\Reg_Bank/registers[7][18] ), .IN1(n158), .SEL(n225), .F(
        \Reg_Bank/n3238 ) );
  MUX U1043 ( .IN0(\Reg_Bank/registers[7][17] ), .IN1(n159), .SEL(n225), .F(
        \Reg_Bank/n3237 ) );
  MUX U1044 ( .IN0(\Reg_Bank/registers[7][16] ), .IN1(n160), .SEL(n225), .F(
        \Reg_Bank/n3236 ) );
  MUX U1045 ( .IN0(\Reg_Bank/registers[7][15] ), .IN1(n161), .SEL(n225), .F(
        \Reg_Bank/n3235 ) );
  MUX U1046 ( .IN0(\Reg_Bank/registers[7][14] ), .IN1(n162), .SEL(n225), .F(
        \Reg_Bank/n3234 ) );
  MUX U1047 ( .IN0(\Reg_Bank/registers[7][13] ), .IN1(n163), .SEL(n225), .F(
        \Reg_Bank/n3233 ) );
  MUX U1048 ( .IN0(\Reg_Bank/registers[7][12] ), .IN1(n164), .SEL(n225), .F(
        \Reg_Bank/n3232 ) );
  MUX U1049 ( .IN0(\Reg_Bank/registers[7][11] ), .IN1(n165), .SEL(n225), .F(
        \Reg_Bank/n3231 ) );
  MUX U1050 ( .IN0(\Reg_Bank/registers[7][10] ), .IN1(n166), .SEL(n225), .F(
        \Reg_Bank/n3230 ) );
  MUX U1051 ( .IN0(\Reg_Bank/registers[7][9] ), .IN1(n167), .SEL(n225), .F(
        \Reg_Bank/n3229 ) );
  MUX U1052 ( .IN0(\Reg_Bank/registers[7][8] ), .IN1(n168), .SEL(n225), .F(
        \Reg_Bank/n3228 ) );
  MUX U1053 ( .IN0(\Reg_Bank/registers[7][7] ), .IN1(n169), .SEL(n225), .F(
        \Reg_Bank/n3227 ) );
  MUX U1054 ( .IN0(\Reg_Bank/registers[7][6] ), .IN1(n170), .SEL(n225), .F(
        \Reg_Bank/n3226 ) );
  MUX U1055 ( .IN0(\Reg_Bank/registers[7][5] ), .IN1(n171), .SEL(n225), .F(
        \Reg_Bank/n3225 ) );
  MUX U1056 ( .IN0(\Reg_Bank/registers[7][4] ), .IN1(n172), .SEL(n225), .F(
        \Reg_Bank/n3224 ) );
  MUX U1057 ( .IN0(\Reg_Bank/registers[7][3] ), .IN1(n173), .SEL(n225), .F(
        \Reg_Bank/n3223 ) );
  MUX U1058 ( .IN0(\Reg_Bank/registers[7][2] ), .IN1(n174), .SEL(n225), .F(
        \Reg_Bank/n3222 ) );
  MUX U1059 ( .IN0(\Reg_Bank/registers[7][1] ), .IN1(n176), .SEL(n225), .F(
        \Reg_Bank/n3221 ) );
  MUX U1060 ( .IN0(\Reg_Bank/registers[7][0] ), .IN1(n177), .SEL(n225), .F(
        \Reg_Bank/n3220 ) );
  ANDN U1061 ( .A(n226), .B(n178), .Z(n225) );
  NAND U1062 ( .A(n224), .B(n227), .Z(n178) );
  MUX U1063 ( .IN0(\Reg_Bank/registers[6][31] ), .IN1(n144), .SEL(n228), .F(
        \Reg_Bank/n3219 ) );
  MUX U1064 ( .IN0(\Reg_Bank/registers[6][30] ), .IN1(n146), .SEL(n228), .F(
        \Reg_Bank/n3218 ) );
  MUX U1065 ( .IN0(\Reg_Bank/registers[6][29] ), .IN1(n147), .SEL(n228), .F(
        \Reg_Bank/n3217 ) );
  MUX U1066 ( .IN0(\Reg_Bank/registers[6][28] ), .IN1(n148), .SEL(n228), .F(
        \Reg_Bank/n3216 ) );
  MUX U1067 ( .IN0(\Reg_Bank/registers[6][27] ), .IN1(n149), .SEL(n228), .F(
        \Reg_Bank/n3215 ) );
  MUX U1068 ( .IN0(\Reg_Bank/registers[6][26] ), .IN1(n150), .SEL(n228), .F(
        \Reg_Bank/n3214 ) );
  MUX U1069 ( .IN0(\Reg_Bank/registers[6][25] ), .IN1(n151), .SEL(n228), .F(
        \Reg_Bank/n3213 ) );
  MUX U1070 ( .IN0(\Reg_Bank/registers[6][24] ), .IN1(n152), .SEL(n228), .F(
        \Reg_Bank/n3212 ) );
  MUX U1071 ( .IN0(\Reg_Bank/registers[6][23] ), .IN1(n153), .SEL(n228), .F(
        \Reg_Bank/n3211 ) );
  MUX U1072 ( .IN0(\Reg_Bank/registers[6][22] ), .IN1(n154), .SEL(n228), .F(
        \Reg_Bank/n3210 ) );
  MUX U1073 ( .IN0(\Reg_Bank/registers[6][21] ), .IN1(n155), .SEL(n228), .F(
        \Reg_Bank/n3209 ) );
  MUX U1074 ( .IN0(\Reg_Bank/registers[6][20] ), .IN1(n156), .SEL(n228), .F(
        \Reg_Bank/n3208 ) );
  MUX U1075 ( .IN0(\Reg_Bank/registers[6][19] ), .IN1(n157), .SEL(n228), .F(
        \Reg_Bank/n3207 ) );
  MUX U1076 ( .IN0(\Reg_Bank/registers[6][18] ), .IN1(n158), .SEL(n228), .F(
        \Reg_Bank/n3206 ) );
  MUX U1077 ( .IN0(\Reg_Bank/registers[6][17] ), .IN1(n159), .SEL(n228), .F(
        \Reg_Bank/n3205 ) );
  MUX U1078 ( .IN0(\Reg_Bank/registers[6][16] ), .IN1(n160), .SEL(n228), .F(
        \Reg_Bank/n3204 ) );
  MUX U1079 ( .IN0(\Reg_Bank/registers[6][15] ), .IN1(n161), .SEL(n228), .F(
        \Reg_Bank/n3203 ) );
  MUX U1080 ( .IN0(\Reg_Bank/registers[6][14] ), .IN1(n162), .SEL(n228), .F(
        \Reg_Bank/n3202 ) );
  MUX U1081 ( .IN0(\Reg_Bank/registers[6][13] ), .IN1(n163), .SEL(n228), .F(
        \Reg_Bank/n3201 ) );
  MUX U1082 ( .IN0(\Reg_Bank/registers[6][12] ), .IN1(n164), .SEL(n228), .F(
        \Reg_Bank/n3200 ) );
  MUX U1083 ( .IN0(\Reg_Bank/registers[6][11] ), .IN1(n165), .SEL(n228), .F(
        \Reg_Bank/n3199 ) );
  MUX U1084 ( .IN0(\Reg_Bank/registers[6][10] ), .IN1(n166), .SEL(n228), .F(
        \Reg_Bank/n3198 ) );
  MUX U1085 ( .IN0(\Reg_Bank/registers[6][9] ), .IN1(n167), .SEL(n228), .F(
        \Reg_Bank/n3197 ) );
  MUX U1086 ( .IN0(\Reg_Bank/registers[6][8] ), .IN1(n168), .SEL(n228), .F(
        \Reg_Bank/n3196 ) );
  MUX U1087 ( .IN0(\Reg_Bank/registers[6][7] ), .IN1(n169), .SEL(n228), .F(
        \Reg_Bank/n3195 ) );
  MUX U1088 ( .IN0(\Reg_Bank/registers[6][6] ), .IN1(n170), .SEL(n228), .F(
        \Reg_Bank/n3194 ) );
  MUX U1089 ( .IN0(\Reg_Bank/registers[6][5] ), .IN1(n171), .SEL(n228), .F(
        \Reg_Bank/n3193 ) );
  MUX U1090 ( .IN0(\Reg_Bank/registers[6][4] ), .IN1(n172), .SEL(n228), .F(
        \Reg_Bank/n3192 ) );
  MUX U1091 ( .IN0(\Reg_Bank/registers[6][3] ), .IN1(n173), .SEL(n228), .F(
        \Reg_Bank/n3191 ) );
  MUX U1092 ( .IN0(\Reg_Bank/registers[6][2] ), .IN1(n174), .SEL(n228), .F(
        \Reg_Bank/n3190 ) );
  MUX U1093 ( .IN0(\Reg_Bank/registers[6][1] ), .IN1(n176), .SEL(n228), .F(
        \Reg_Bank/n3189 ) );
  MUX U1094 ( .IN0(\Reg_Bank/registers[6][0] ), .IN1(n177), .SEL(n228), .F(
        \Reg_Bank/n3188 ) );
  AND U1095 ( .A(n182), .B(n226), .Z(n228) );
  AND U1096 ( .A(n224), .B(n229), .Z(n182) );
  MUX U1097 ( .IN0(\Reg_Bank/registers[5][31] ), .IN1(n144), .SEL(n230), .F(
        \Reg_Bank/n3187 ) );
  MUX U1098 ( .IN0(\Reg_Bank/registers[5][30] ), .IN1(n146), .SEL(n230), .F(
        \Reg_Bank/n3186 ) );
  MUX U1099 ( .IN0(\Reg_Bank/registers[5][29] ), .IN1(n147), .SEL(n230), .F(
        \Reg_Bank/n3185 ) );
  MUX U1100 ( .IN0(\Reg_Bank/registers[5][28] ), .IN1(n148), .SEL(n230), .F(
        \Reg_Bank/n3184 ) );
  MUX U1101 ( .IN0(\Reg_Bank/registers[5][27] ), .IN1(n149), .SEL(n230), .F(
        \Reg_Bank/n3183 ) );
  MUX U1102 ( .IN0(\Reg_Bank/registers[5][26] ), .IN1(n150), .SEL(n230), .F(
        \Reg_Bank/n3182 ) );
  MUX U1103 ( .IN0(\Reg_Bank/registers[5][25] ), .IN1(n151), .SEL(n230), .F(
        \Reg_Bank/n3181 ) );
  MUX U1104 ( .IN0(\Reg_Bank/registers[5][24] ), .IN1(n152), .SEL(n230), .F(
        \Reg_Bank/n3180 ) );
  MUX U1105 ( .IN0(\Reg_Bank/registers[5][23] ), .IN1(n153), .SEL(n230), .F(
        \Reg_Bank/n3179 ) );
  MUX U1106 ( .IN0(\Reg_Bank/registers[5][22] ), .IN1(n154), .SEL(n230), .F(
        \Reg_Bank/n3178 ) );
  MUX U1107 ( .IN0(\Reg_Bank/registers[5][21] ), .IN1(n155), .SEL(n230), .F(
        \Reg_Bank/n3177 ) );
  MUX U1108 ( .IN0(\Reg_Bank/registers[5][20] ), .IN1(n156), .SEL(n230), .F(
        \Reg_Bank/n3176 ) );
  MUX U1109 ( .IN0(\Reg_Bank/registers[5][19] ), .IN1(n157), .SEL(n230), .F(
        \Reg_Bank/n3175 ) );
  MUX U1110 ( .IN0(\Reg_Bank/registers[5][18] ), .IN1(n158), .SEL(n230), .F(
        \Reg_Bank/n3174 ) );
  MUX U1111 ( .IN0(\Reg_Bank/registers[5][17] ), .IN1(n159), .SEL(n230), .F(
        \Reg_Bank/n3173 ) );
  MUX U1112 ( .IN0(\Reg_Bank/registers[5][16] ), .IN1(n160), .SEL(n230), .F(
        \Reg_Bank/n3172 ) );
  MUX U1113 ( .IN0(\Reg_Bank/registers[5][15] ), .IN1(n161), .SEL(n230), .F(
        \Reg_Bank/n3171 ) );
  MUX U1114 ( .IN0(\Reg_Bank/registers[5][14] ), .IN1(n162), .SEL(n230), .F(
        \Reg_Bank/n3170 ) );
  MUX U1115 ( .IN0(\Reg_Bank/registers[5][13] ), .IN1(n163), .SEL(n230), .F(
        \Reg_Bank/n3169 ) );
  MUX U1116 ( .IN0(\Reg_Bank/registers[5][12] ), .IN1(n164), .SEL(n230), .F(
        \Reg_Bank/n3168 ) );
  MUX U1117 ( .IN0(\Reg_Bank/registers[5][11] ), .IN1(n165), .SEL(n230), .F(
        \Reg_Bank/n3167 ) );
  MUX U1118 ( .IN0(\Reg_Bank/registers[5][10] ), .IN1(n166), .SEL(n230), .F(
        \Reg_Bank/n3166 ) );
  MUX U1119 ( .IN0(\Reg_Bank/registers[5][9] ), .IN1(n167), .SEL(n230), .F(
        \Reg_Bank/n3165 ) );
  MUX U1120 ( .IN0(\Reg_Bank/registers[5][8] ), .IN1(n168), .SEL(n230), .F(
        \Reg_Bank/n3164 ) );
  MUX U1121 ( .IN0(\Reg_Bank/registers[5][7] ), .IN1(n169), .SEL(n230), .F(
        \Reg_Bank/n3163 ) );
  MUX U1122 ( .IN0(\Reg_Bank/registers[5][6] ), .IN1(n170), .SEL(n230), .F(
        \Reg_Bank/n3162 ) );
  MUX U1123 ( .IN0(\Reg_Bank/registers[5][5] ), .IN1(n171), .SEL(n230), .F(
        \Reg_Bank/n3161 ) );
  MUX U1124 ( .IN0(\Reg_Bank/registers[5][4] ), .IN1(n172), .SEL(n230), .F(
        \Reg_Bank/n3160 ) );
  MUX U1125 ( .IN0(\Reg_Bank/registers[5][3] ), .IN1(n173), .SEL(n230), .F(
        \Reg_Bank/n3159 ) );
  MUX U1126 ( .IN0(\Reg_Bank/registers[5][2] ), .IN1(n174), .SEL(n230), .F(
        \Reg_Bank/n3158 ) );
  MUX U1127 ( .IN0(\Reg_Bank/registers[5][1] ), .IN1(n176), .SEL(n230), .F(
        \Reg_Bank/n3157 ) );
  MUX U1128 ( .IN0(\Reg_Bank/registers[5][0] ), .IN1(n177), .SEL(n230), .F(
        \Reg_Bank/n3156 ) );
  AND U1129 ( .A(n185), .B(n226), .Z(n230) );
  AND U1130 ( .A(n224), .B(n231), .Z(n185) );
  MUX U1131 ( .IN0(\Reg_Bank/registers[4][31] ), .IN1(n144), .SEL(n232), .F(
        \Reg_Bank/n3155 ) );
  MUX U1132 ( .IN0(\Reg_Bank/registers[4][30] ), .IN1(n146), .SEL(n232), .F(
        \Reg_Bank/n3154 ) );
  MUX U1133 ( .IN0(\Reg_Bank/registers[4][29] ), .IN1(n147), .SEL(n232), .F(
        \Reg_Bank/n3153 ) );
  MUX U1134 ( .IN0(\Reg_Bank/registers[4][28] ), .IN1(n148), .SEL(n232), .F(
        \Reg_Bank/n3152 ) );
  MUX U1135 ( .IN0(\Reg_Bank/registers[4][27] ), .IN1(n149), .SEL(n232), .F(
        \Reg_Bank/n3151 ) );
  MUX U1136 ( .IN0(\Reg_Bank/registers[4][26] ), .IN1(n150), .SEL(n232), .F(
        \Reg_Bank/n3150 ) );
  MUX U1137 ( .IN0(\Reg_Bank/registers[4][25] ), .IN1(n151), .SEL(n232), .F(
        \Reg_Bank/n3149 ) );
  MUX U1138 ( .IN0(\Reg_Bank/registers[4][24] ), .IN1(n152), .SEL(n232), .F(
        \Reg_Bank/n3148 ) );
  MUX U1139 ( .IN0(\Reg_Bank/registers[4][23] ), .IN1(n153), .SEL(n232), .F(
        \Reg_Bank/n3147 ) );
  MUX U1140 ( .IN0(\Reg_Bank/registers[4][22] ), .IN1(n154), .SEL(n232), .F(
        \Reg_Bank/n3146 ) );
  MUX U1141 ( .IN0(\Reg_Bank/registers[4][21] ), .IN1(n155), .SEL(n232), .F(
        \Reg_Bank/n3145 ) );
  MUX U1142 ( .IN0(\Reg_Bank/registers[4][20] ), .IN1(n156), .SEL(n232), .F(
        \Reg_Bank/n3144 ) );
  MUX U1143 ( .IN0(\Reg_Bank/registers[4][19] ), .IN1(n157), .SEL(n232), .F(
        \Reg_Bank/n3143 ) );
  MUX U1144 ( .IN0(\Reg_Bank/registers[4][18] ), .IN1(n158), .SEL(n232), .F(
        \Reg_Bank/n3142 ) );
  MUX U1145 ( .IN0(\Reg_Bank/registers[4][17] ), .IN1(n159), .SEL(n232), .F(
        \Reg_Bank/n3141 ) );
  MUX U1146 ( .IN0(\Reg_Bank/registers[4][16] ), .IN1(n160), .SEL(n232), .F(
        \Reg_Bank/n3140 ) );
  MUX U1147 ( .IN0(\Reg_Bank/registers[4][15] ), .IN1(n161), .SEL(n232), .F(
        \Reg_Bank/n3139 ) );
  MUX U1148 ( .IN0(\Reg_Bank/registers[4][14] ), .IN1(n162), .SEL(n232), .F(
        \Reg_Bank/n3138 ) );
  MUX U1149 ( .IN0(\Reg_Bank/registers[4][13] ), .IN1(n163), .SEL(n232), .F(
        \Reg_Bank/n3137 ) );
  MUX U1150 ( .IN0(\Reg_Bank/registers[4][12] ), .IN1(n164), .SEL(n232), .F(
        \Reg_Bank/n3136 ) );
  MUX U1151 ( .IN0(\Reg_Bank/registers[4][11] ), .IN1(n165), .SEL(n232), .F(
        \Reg_Bank/n3135 ) );
  MUX U1152 ( .IN0(\Reg_Bank/registers[4][10] ), .IN1(n166), .SEL(n232), .F(
        \Reg_Bank/n3134 ) );
  MUX U1153 ( .IN0(\Reg_Bank/registers[4][9] ), .IN1(n167), .SEL(n232), .F(
        \Reg_Bank/n3133 ) );
  MUX U1154 ( .IN0(\Reg_Bank/registers[4][8] ), .IN1(n168), .SEL(n232), .F(
        \Reg_Bank/n3132 ) );
  MUX U1155 ( .IN0(\Reg_Bank/registers[4][7] ), .IN1(n169), .SEL(n232), .F(
        \Reg_Bank/n3131 ) );
  MUX U1156 ( .IN0(\Reg_Bank/registers[4][6] ), .IN1(n170), .SEL(n232), .F(
        \Reg_Bank/n3130 ) );
  MUX U1157 ( .IN0(\Reg_Bank/registers[4][5] ), .IN1(n171), .SEL(n232), .F(
        \Reg_Bank/n3129 ) );
  MUX U1158 ( .IN0(\Reg_Bank/registers[4][4] ), .IN1(n172), .SEL(n232), .F(
        \Reg_Bank/n3128 ) );
  MUX U1159 ( .IN0(\Reg_Bank/registers[4][3] ), .IN1(n173), .SEL(n232), .F(
        \Reg_Bank/n3127 ) );
  MUX U1160 ( .IN0(\Reg_Bank/registers[4][2] ), .IN1(n174), .SEL(n232), .F(
        \Reg_Bank/n3126 ) );
  MUX U1161 ( .IN0(\Reg_Bank/registers[4][1] ), .IN1(n176), .SEL(n232), .F(
        \Reg_Bank/n3125 ) );
  MUX U1162 ( .IN0(\Reg_Bank/registers[4][0] ), .IN1(n177), .SEL(n232), .F(
        \Reg_Bank/n3124 ) );
  AND U1163 ( .A(n188), .B(n226), .Z(n232) );
  AND U1164 ( .A(n224), .B(n223), .Z(n188) );
  ANDN U1165 ( .A(n233), .B(n234), .Z(n223) );
  MUX U1166 ( .IN0(\Reg_Bank/registers[3][31] ), .IN1(n144), .SEL(n235), .F(
        \Reg_Bank/n3123 ) );
  MUX U1167 ( .IN0(\Reg_Bank/registers[3][30] ), .IN1(n146), .SEL(n235), .F(
        \Reg_Bank/n3122 ) );
  MUX U1168 ( .IN0(\Reg_Bank/registers[3][29] ), .IN1(n147), .SEL(n235), .F(
        \Reg_Bank/n3121 ) );
  MUX U1169 ( .IN0(\Reg_Bank/registers[3][28] ), .IN1(n148), .SEL(n235), .F(
        \Reg_Bank/n3120 ) );
  MUX U1170 ( .IN0(\Reg_Bank/registers[3][27] ), .IN1(n149), .SEL(n235), .F(
        \Reg_Bank/n3119 ) );
  MUX U1171 ( .IN0(\Reg_Bank/registers[3][26] ), .IN1(n150), .SEL(n235), .F(
        \Reg_Bank/n3118 ) );
  MUX U1172 ( .IN0(\Reg_Bank/registers[3][25] ), .IN1(n151), .SEL(n235), .F(
        \Reg_Bank/n3117 ) );
  MUX U1173 ( .IN0(\Reg_Bank/registers[3][24] ), .IN1(n152), .SEL(n235), .F(
        \Reg_Bank/n3116 ) );
  MUX U1174 ( .IN0(\Reg_Bank/registers[3][23] ), .IN1(n153), .SEL(n235), .F(
        \Reg_Bank/n3115 ) );
  MUX U1175 ( .IN0(\Reg_Bank/registers[3][22] ), .IN1(n154), .SEL(n235), .F(
        \Reg_Bank/n3114 ) );
  MUX U1176 ( .IN0(\Reg_Bank/registers[3][21] ), .IN1(n155), .SEL(n235), .F(
        \Reg_Bank/n3113 ) );
  MUX U1177 ( .IN0(\Reg_Bank/registers[3][20] ), .IN1(n156), .SEL(n235), .F(
        \Reg_Bank/n3112 ) );
  MUX U1178 ( .IN0(\Reg_Bank/registers[3][19] ), .IN1(n157), .SEL(n235), .F(
        \Reg_Bank/n3111 ) );
  MUX U1179 ( .IN0(\Reg_Bank/registers[3][18] ), .IN1(n158), .SEL(n235), .F(
        \Reg_Bank/n3110 ) );
  MUX U1180 ( .IN0(\Reg_Bank/registers[3][17] ), .IN1(n159), .SEL(n235), .F(
        \Reg_Bank/n3109 ) );
  MUX U1181 ( .IN0(\Reg_Bank/registers[3][16] ), .IN1(n160), .SEL(n235), .F(
        \Reg_Bank/n3108 ) );
  MUX U1182 ( .IN0(\Reg_Bank/registers[3][15] ), .IN1(n161), .SEL(n235), .F(
        \Reg_Bank/n3107 ) );
  MUX U1183 ( .IN0(\Reg_Bank/registers[3][14] ), .IN1(n162), .SEL(n235), .F(
        \Reg_Bank/n3106 ) );
  MUX U1184 ( .IN0(\Reg_Bank/registers[3][13] ), .IN1(n163), .SEL(n235), .F(
        \Reg_Bank/n3105 ) );
  MUX U1185 ( .IN0(\Reg_Bank/registers[3][12] ), .IN1(n164), .SEL(n235), .F(
        \Reg_Bank/n3104 ) );
  MUX U1186 ( .IN0(\Reg_Bank/registers[3][11] ), .IN1(n165), .SEL(n235), .F(
        \Reg_Bank/n3103 ) );
  MUX U1187 ( .IN0(\Reg_Bank/registers[3][10] ), .IN1(n166), .SEL(n235), .F(
        \Reg_Bank/n3102 ) );
  MUX U1188 ( .IN0(\Reg_Bank/registers[3][9] ), .IN1(n167), .SEL(n235), .F(
        \Reg_Bank/n3101 ) );
  MUX U1189 ( .IN0(\Reg_Bank/registers[3][8] ), .IN1(n168), .SEL(n235), .F(
        \Reg_Bank/n3100 ) );
  MUX U1190 ( .IN0(\Reg_Bank/registers[3][7] ), .IN1(n169), .SEL(n235), .F(
        \Reg_Bank/n3099 ) );
  MUX U1191 ( .IN0(\Reg_Bank/registers[3][6] ), .IN1(n170), .SEL(n235), .F(
        \Reg_Bank/n3098 ) );
  MUX U1192 ( .IN0(\Reg_Bank/registers[3][5] ), .IN1(n171), .SEL(n235), .F(
        \Reg_Bank/n3097 ) );
  MUX U1193 ( .IN0(\Reg_Bank/registers[3][4] ), .IN1(n172), .SEL(n235), .F(
        \Reg_Bank/n3096 ) );
  MUX U1194 ( .IN0(\Reg_Bank/registers[3][3] ), .IN1(n173), .SEL(n235), .F(
        \Reg_Bank/n3095 ) );
  MUX U1195 ( .IN0(\Reg_Bank/registers[3][2] ), .IN1(n174), .SEL(n235), .F(
        \Reg_Bank/n3094 ) );
  MUX U1196 ( .IN0(\Reg_Bank/registers[3][1] ), .IN1(n176), .SEL(n235), .F(
        \Reg_Bank/n3093 ) );
  MUX U1197 ( .IN0(\Reg_Bank/registers[3][0] ), .IN1(n177), .SEL(n235), .F(
        \Reg_Bank/n3092 ) );
  ANDN U1198 ( .A(n226), .B(n190), .Z(n235) );
  IV U1199 ( .A(n217), .Z(n190) );
  ANDN U1200 ( .A(n227), .B(n224), .Z(n217) );
  AND U1201 ( .A(n234), .B(n236), .Z(n227) );
  MUX U1202 ( .IN0(\Reg_Bank/registers[2][31] ), .IN1(n144), .SEL(n237), .F(
        \Reg_Bank/n3091 ) );
  MUX U1203 ( .IN0(\Reg_Bank/registers[2][30] ), .IN1(n146), .SEL(n237), .F(
        \Reg_Bank/n3090 ) );
  MUX U1204 ( .IN0(\Reg_Bank/registers[2][29] ), .IN1(n147), .SEL(n237), .F(
        \Reg_Bank/n3089 ) );
  MUX U1205 ( .IN0(\Reg_Bank/registers[2][28] ), .IN1(n148), .SEL(n237), .F(
        \Reg_Bank/n3088 ) );
  MUX U1206 ( .IN0(\Reg_Bank/registers[2][27] ), .IN1(n149), .SEL(n237), .F(
        \Reg_Bank/n3087 ) );
  MUX U1207 ( .IN0(\Reg_Bank/registers[2][26] ), .IN1(n150), .SEL(n237), .F(
        \Reg_Bank/n3086 ) );
  MUX U1208 ( .IN0(\Reg_Bank/registers[2][25] ), .IN1(n151), .SEL(n237), .F(
        \Reg_Bank/n3085 ) );
  MUX U1209 ( .IN0(\Reg_Bank/registers[2][24] ), .IN1(n152), .SEL(n237), .F(
        \Reg_Bank/n3084 ) );
  MUX U1210 ( .IN0(\Reg_Bank/registers[2][23] ), .IN1(n153), .SEL(n237), .F(
        \Reg_Bank/n3083 ) );
  MUX U1211 ( .IN0(\Reg_Bank/registers[2][22] ), .IN1(n154), .SEL(n237), .F(
        \Reg_Bank/n3082 ) );
  MUX U1212 ( .IN0(\Reg_Bank/registers[2][21] ), .IN1(n155), .SEL(n237), .F(
        \Reg_Bank/n3081 ) );
  MUX U1213 ( .IN0(\Reg_Bank/registers[2][20] ), .IN1(n156), .SEL(n237), .F(
        \Reg_Bank/n3080 ) );
  MUX U1214 ( .IN0(\Reg_Bank/registers[2][19] ), .IN1(n157), .SEL(n237), .F(
        \Reg_Bank/n3079 ) );
  MUX U1215 ( .IN0(\Reg_Bank/registers[2][18] ), .IN1(n158), .SEL(n237), .F(
        \Reg_Bank/n3078 ) );
  MUX U1216 ( .IN0(\Reg_Bank/registers[2][17] ), .IN1(n159), .SEL(n237), .F(
        \Reg_Bank/n3077 ) );
  MUX U1217 ( .IN0(\Reg_Bank/registers[2][16] ), .IN1(n160), .SEL(n237), .F(
        \Reg_Bank/n3076 ) );
  MUX U1218 ( .IN0(\Reg_Bank/registers[2][15] ), .IN1(n161), .SEL(n237), .F(
        \Reg_Bank/n3075 ) );
  MUX U1219 ( .IN0(\Reg_Bank/registers[2][14] ), .IN1(n162), .SEL(n237), .F(
        \Reg_Bank/n3074 ) );
  MUX U1220 ( .IN0(\Reg_Bank/registers[2][13] ), .IN1(n163), .SEL(n237), .F(
        \Reg_Bank/n3073 ) );
  MUX U1221 ( .IN0(\Reg_Bank/registers[2][12] ), .IN1(n164), .SEL(n237), .F(
        \Reg_Bank/n3072 ) );
  MUX U1222 ( .IN0(\Reg_Bank/registers[2][11] ), .IN1(n165), .SEL(n237), .F(
        \Reg_Bank/n3071 ) );
  MUX U1223 ( .IN0(\Reg_Bank/registers[2][10] ), .IN1(n166), .SEL(n237), .F(
        \Reg_Bank/n3070 ) );
  MUX U1224 ( .IN0(\Reg_Bank/registers[2][9] ), .IN1(n167), .SEL(n237), .F(
        \Reg_Bank/n3069 ) );
  MUX U1225 ( .IN0(\Reg_Bank/registers[2][8] ), .IN1(n168), .SEL(n237), .F(
        \Reg_Bank/n3068 ) );
  MUX U1226 ( .IN0(\Reg_Bank/registers[2][7] ), .IN1(n169), .SEL(n237), .F(
        \Reg_Bank/n3067 ) );
  MUX U1227 ( .IN0(\Reg_Bank/registers[2][6] ), .IN1(n170), .SEL(n237), .F(
        \Reg_Bank/n3066 ) );
  MUX U1228 ( .IN0(\Reg_Bank/registers[2][5] ), .IN1(n171), .SEL(n237), .F(
        \Reg_Bank/n3065 ) );
  MUX U1229 ( .IN0(\Reg_Bank/registers[2][4] ), .IN1(n172), .SEL(n237), .F(
        \Reg_Bank/n3064 ) );
  MUX U1230 ( .IN0(\Reg_Bank/registers[2][3] ), .IN1(n173), .SEL(n237), .F(
        \Reg_Bank/n3063 ) );
  MUX U1231 ( .IN0(\Reg_Bank/registers[2][2] ), .IN1(n174), .SEL(n237), .F(
        \Reg_Bank/n3062 ) );
  MUX U1232 ( .IN0(\Reg_Bank/registers[2][1] ), .IN1(n176), .SEL(n237), .F(
        \Reg_Bank/n3061 ) );
  MUX U1233 ( .IN0(\Reg_Bank/registers[2][0] ), .IN1(n177), .SEL(n237), .F(
        \Reg_Bank/n3060 ) );
  ANDN U1234 ( .A(n226), .B(n192), .Z(n237) );
  IV U1235 ( .A(n219), .Z(n192) );
  ANDN U1236 ( .A(n229), .B(n224), .Z(n219) );
  ANDN U1237 ( .A(n234), .B(n236), .Z(n229) );
  MUX U1238 ( .IN0(\Reg_Bank/registers[1][31] ), .IN1(n144), .SEL(n238), .F(
        \Reg_Bank/n3059 ) );
  NAND U1239 ( .A(n239), .B(n240), .Z(n144) );
  AND U1240 ( .A(n241), .B(n242), .Z(n240) );
  NANDN U1241 ( .B(n243), .A(n244), .Z(n242) );
  AND U1242 ( .A(n245), .B(n246), .Z(n241) );
  NANDN U1243 ( .B(n247), .A(\Data_Mem/N714 ), .Z(n246) );
  OR U1244 ( .A(n248), .B(n249), .Z(n245) );
  AND U1245 ( .A(n250), .B(n251), .Z(n239) );
  NANDN U1246 ( .B(n252), .A(imm[15]), .Z(n251) );
  MUX U1247 ( .IN0(\Reg_Bank/registers[1][30] ), .IN1(n146), .SEL(n238), .F(
        \Reg_Bank/n3058 ) );
  NAND U1248 ( .A(n253), .B(n254), .Z(n146) );
  AND U1249 ( .A(n255), .B(n256), .Z(n254) );
  NANDN U1250 ( .B(n243), .A(pc_plus4[30]), .Z(n256) );
  AND U1251 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U1252 ( .B(n247), .A(\Data_Mem/N715 ), .Z(n258) );
  OR U1253 ( .A(n248), .B(n259), .Z(n257) );
  AND U1254 ( .A(n250), .B(n260), .Z(n253) );
  NANDN U1255 ( .B(n252), .A(imm[14]), .Z(n260) );
  MUX U1256 ( .IN0(\Reg_Bank/registers[1][29] ), .IN1(n147), .SEL(n238), .F(
        \Reg_Bank/n3057 ) );
  NAND U1257 ( .A(n261), .B(n262), .Z(n147) );
  AND U1258 ( .A(n263), .B(n264), .Z(n262) );
  NANDN U1259 ( .B(n243), .A(pc_plus4[29]), .Z(n264) );
  AND U1260 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U1261 ( .B(n247), .A(\Data_Mem/N716 ), .Z(n266) );
  OR U1262 ( .A(n248), .B(n267), .Z(n265) );
  AND U1263 ( .A(n250), .B(n268), .Z(n261) );
  NANDN U1264 ( .B(n252), .A(imm[13]), .Z(n268) );
  MUX U1265 ( .IN0(\Reg_Bank/registers[1][28] ), .IN1(n148), .SEL(n238), .F(
        \Reg_Bank/n3056 ) );
  NAND U1266 ( .A(n269), .B(n270), .Z(n148) );
  AND U1267 ( .A(n271), .B(n272), .Z(n270) );
  NANDN U1268 ( .B(n243), .A(pc_plus4[28]), .Z(n272) );
  AND U1269 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U1270 ( .B(n247), .A(\Data_Mem/N717 ), .Z(n274) );
  OR U1271 ( .A(n248), .B(n275), .Z(n273) );
  AND U1272 ( .A(n250), .B(n276), .Z(n269) );
  NANDN U1273 ( .B(n252), .A(imm[12]), .Z(n276) );
  MUX U1274 ( .IN0(\Reg_Bank/registers[1][27] ), .IN1(n149), .SEL(n238), .F(
        \Reg_Bank/n3055 ) );
  NAND U1275 ( .A(n277), .B(n278), .Z(n149) );
  AND U1276 ( .A(n279), .B(n280), .Z(n278) );
  NANDN U1277 ( .B(n243), .A(pc_plus4[27]), .Z(n280) );
  AND U1278 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U1279 ( .B(n247), .A(\Data_Mem/N718 ), .Z(n282) );
  OR U1280 ( .A(n248), .B(n283), .Z(n281) );
  AND U1281 ( .A(n250), .B(n284), .Z(n277) );
  NANDN U1282 ( .B(n252), .A(imm[11]), .Z(n284) );
  MUX U1283 ( .IN0(\Reg_Bank/registers[1][26] ), .IN1(n150), .SEL(n238), .F(
        \Reg_Bank/n3054 ) );
  NAND U1284 ( .A(n285), .B(n286), .Z(n150) );
  AND U1285 ( .A(n287), .B(n288), .Z(n286) );
  NANDN U1286 ( .B(n243), .A(pc_plus4[26]), .Z(n288) );
  AND U1287 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U1288 ( .B(n247), .A(\Data_Mem/N719 ), .Z(n290) );
  OR U1289 ( .A(n248), .B(n291), .Z(n289) );
  AND U1290 ( .A(n250), .B(n292), .Z(n285) );
  NANDN U1291 ( .B(n252), .A(imm[10]), .Z(n292) );
  MUX U1292 ( .IN0(\Reg_Bank/registers[1][25] ), .IN1(n151), .SEL(n238), .F(
        \Reg_Bank/n3053 ) );
  NAND U1293 ( .A(n293), .B(n294), .Z(n151) );
  AND U1294 ( .A(n295), .B(n296), .Z(n294) );
  NANDN U1295 ( .B(n243), .A(pc_plus4[25]), .Z(n296) );
  AND U1296 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U1297 ( .B(n247), .A(\Data_Mem/N720 ), .Z(n298) );
  OR U1298 ( .A(n248), .B(n299), .Z(n297) );
  AND U1299 ( .A(n250), .B(n300), .Z(n293) );
  NANDN U1300 ( .B(n252), .A(imm[9]), .Z(n300) );
  MUX U1301 ( .IN0(\Reg_Bank/registers[1][24] ), .IN1(n152), .SEL(n238), .F(
        \Reg_Bank/n3052 ) );
  NAND U1302 ( .A(n301), .B(n302), .Z(n152) );
  AND U1303 ( .A(n303), .B(n304), .Z(n302) );
  NANDN U1304 ( .B(n243), .A(pc_plus4[24]), .Z(n304) );
  AND U1305 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U1306 ( .B(n247), .A(\Data_Mem/N721 ), .Z(n306) );
  OR U1307 ( .A(n248), .B(n307), .Z(n305) );
  AND U1308 ( .A(n250), .B(n308), .Z(n301) );
  NANDN U1309 ( .B(n252), .A(imm[8]), .Z(n308) );
  MUX U1310 ( .IN0(\Reg_Bank/registers[1][23] ), .IN1(n153), .SEL(n238), .F(
        \Reg_Bank/n3051 ) );
  NAND U1311 ( .A(n309), .B(n310), .Z(n153) );
  AND U1312 ( .A(n311), .B(n312), .Z(n310) );
  NANDN U1313 ( .B(n243), .A(pc_plus4[23]), .Z(n312) );
  AND U1314 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U1315 ( .B(n247), .A(\Data_Mem/N722 ), .Z(n314) );
  OR U1316 ( .A(n248), .B(n315), .Z(n313) );
  AND U1317 ( .A(n250), .B(n316), .Z(n309) );
  NANDN U1318 ( .B(n252), .A(imm[7]), .Z(n316) );
  MUX U1319 ( .IN0(\Reg_Bank/registers[1][22] ), .IN1(n154), .SEL(n238), .F(
        \Reg_Bank/n3050 ) );
  NAND U1320 ( .A(n317), .B(n318), .Z(n154) );
  AND U1321 ( .A(n319), .B(n320), .Z(n318) );
  NANDN U1322 ( .B(n243), .A(pc_plus4[22]), .Z(n320) );
  AND U1323 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U1324 ( .B(n247), .A(\Data_Mem/N723 ), .Z(n322) );
  OR U1325 ( .A(n248), .B(n323), .Z(n321) );
  AND U1326 ( .A(n250), .B(n324), .Z(n317) );
  NANDN U1327 ( .B(n252), .A(imm[6]), .Z(n324) );
  MUX U1328 ( .IN0(\Reg_Bank/registers[1][21] ), .IN1(n155), .SEL(n238), .F(
        \Reg_Bank/n3049 ) );
  NAND U1329 ( .A(n325), .B(n326), .Z(n155) );
  AND U1330 ( .A(n327), .B(n328), .Z(n326) );
  NANDN U1331 ( .B(n243), .A(pc_plus4[21]), .Z(n328) );
  AND U1332 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U1333 ( .B(n247), .A(\Data_Mem/N724 ), .Z(n330) );
  OR U1334 ( .A(n248), .B(n331), .Z(n329) );
  AND U1335 ( .A(n250), .B(n332), .Z(n325) );
  NANDN U1336 ( .B(n252), .A(imm[5]), .Z(n332) );
  MUX U1337 ( .IN0(\Reg_Bank/registers[1][20] ), .IN1(n156), .SEL(n238), .F(
        \Reg_Bank/n3048 ) );
  NAND U1338 ( .A(n333), .B(n334), .Z(n156) );
  AND U1339 ( .A(n335), .B(n336), .Z(n334) );
  NANDN U1340 ( .B(n243), .A(pc_plus4[20]), .Z(n336) );
  AND U1341 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U1342 ( .B(n247), .A(\Data_Mem/N725 ), .Z(n338) );
  OR U1343 ( .A(n248), .B(n339), .Z(n337) );
  AND U1344 ( .A(n250), .B(n340), .Z(n333) );
  OR U1345 ( .A(n252), .B(n341), .Z(n340) );
  MUX U1346 ( .IN0(\Reg_Bank/registers[1][19] ), .IN1(n157), .SEL(n238), .F(
        \Reg_Bank/n3047 ) );
  NAND U1347 ( .A(n342), .B(n343), .Z(n157) );
  AND U1348 ( .A(n344), .B(n345), .Z(n343) );
  NANDN U1349 ( .B(n243), .A(pc_plus4[19]), .Z(n345) );
  AND U1350 ( .A(n346), .B(n347), .Z(n344) );
  NANDN U1351 ( .B(n247), .A(\Data_Mem/N726 ), .Z(n347) );
  OR U1352 ( .A(n248), .B(n348), .Z(n346) );
  AND U1353 ( .A(n250), .B(n349), .Z(n342) );
  OR U1354 ( .A(n252), .B(n350), .Z(n349) );
  MUX U1355 ( .IN0(\Reg_Bank/registers[1][18] ), .IN1(n158), .SEL(n238), .F(
        \Reg_Bank/n3046 ) );
  NAND U1356 ( .A(n351), .B(n352), .Z(n158) );
  AND U1357 ( .A(n353), .B(n354), .Z(n352) );
  NANDN U1358 ( .B(n243), .A(pc_plus4[18]), .Z(n354) );
  AND U1359 ( .A(n355), .B(n356), .Z(n353) );
  NANDN U1360 ( .B(n247), .A(\Data_Mem/N727 ), .Z(n356) );
  OR U1361 ( .A(n248), .B(n357), .Z(n355) );
  AND U1362 ( .A(n250), .B(n358), .Z(n351) );
  OR U1363 ( .A(n252), .B(n359), .Z(n358) );
  MUX U1364 ( .IN0(\Reg_Bank/registers[1][17] ), .IN1(n159), .SEL(n238), .F(
        \Reg_Bank/n3045 ) );
  NAND U1365 ( .A(n360), .B(n361), .Z(n159) );
  AND U1366 ( .A(n362), .B(n363), .Z(n361) );
  NANDN U1367 ( .B(n243), .A(pc_plus4[17]), .Z(n363) );
  AND U1368 ( .A(n364), .B(n365), .Z(n362) );
  NANDN U1369 ( .B(n247), .A(\Data_Mem/N728 ), .Z(n365) );
  OR U1370 ( .A(n248), .B(n366), .Z(n364) );
  AND U1371 ( .A(n250), .B(n367), .Z(n360) );
  OR U1372 ( .A(n252), .B(n14), .Z(n367) );
  MUX U1373 ( .IN0(\Reg_Bank/registers[1][16] ), .IN1(n160), .SEL(n238), .F(
        \Reg_Bank/n3044 ) );
  NAND U1374 ( .A(n368), .B(n369), .Z(n160) );
  AND U1375 ( .A(n370), .B(n371), .Z(n369) );
  NANDN U1376 ( .B(n243), .A(pc_plus4[16]), .Z(n371) );
  AND U1377 ( .A(n372), .B(n373), .Z(n370) );
  NANDN U1378 ( .B(n247), .A(\Data_Mem/N729 ), .Z(n373) );
  OR U1379 ( .A(n248), .B(n374), .Z(n372) );
  AND U1380 ( .A(n250), .B(n375), .Z(n368) );
  OR U1381 ( .A(n252), .B(n376), .Z(n375) );
  NAND U1382 ( .A(n377), .B(n378), .Z(n252) );
  AND U1383 ( .A(n379), .B(n380), .Z(n250) );
  IV U1384 ( .A(n381), .Z(n380) );
  NAND U1385 ( .A(n382), .B(n383), .Z(n379) );
  NANDN U1386 ( .B(n384), .A(n385), .Z(n382) );
  MUX U1387 ( .IN0(\Reg_Bank/registers[1][15] ), .IN1(n161), .SEL(n238), .F(
        \Reg_Bank/n3043 ) );
  NAND U1388 ( .A(n386), .B(n387), .Z(n161) );
  AND U1389 ( .A(n388), .B(n389), .Z(n387) );
  NANDN U1390 ( .B(n247), .A(\Data_Mem/N730 ), .Z(n389) );
  ANDN U1391 ( .A(n390), .B(n381), .Z(n388) );
  OR U1392 ( .A(n248), .B(n391), .Z(n390) );
  AND U1393 ( .A(n392), .B(n393), .Z(n386) );
  NANDN U1394 ( .B(n243), .A(pc_plus4[15]), .Z(n393) );
  AND U1395 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U1396 ( .B(n396), .A(n383), .Z(n395) );
  NANDN U1397 ( .B(n396), .A(n397), .Z(n394) );
  ANDN U1398 ( .A(n398), .B(n384), .Z(n396) );
  AND U1399 ( .A(\Data_Mem/N730 ), .B(n399), .Z(n384) );
  NANDN U1400 ( .B(n399), .A(\Data_Mem/N714 ), .Z(n398) );
  MUX U1401 ( .IN0(\Reg_Bank/registers[1][14] ), .IN1(n162), .SEL(n238), .F(
        \Reg_Bank/n3042 ) );
  NAND U1402 ( .A(n400), .B(n401), .Z(n162) );
  AND U1403 ( .A(n402), .B(n403), .Z(n401) );
  NANDN U1404 ( .B(n247), .A(\Data_Mem/N731 ), .Z(n403) );
  ANDN U1405 ( .A(n404), .B(n381), .Z(n402) );
  OR U1406 ( .A(n248), .B(n405), .Z(n404) );
  AND U1407 ( .A(n406), .B(n407), .Z(n400) );
  NANDN U1408 ( .B(n243), .A(pc_plus4[14]), .Z(n407) );
  AND U1409 ( .A(n408), .B(n409), .Z(n406) );
  NAND U1410 ( .A(n410), .B(n383), .Z(n409) );
  NAND U1411 ( .A(n410), .B(n397), .Z(n408) );
  MUX U1412 ( .IN0(\Data_Mem/N731 ), .IN1(\Data_Mem/N715 ), .SEL(n411), .F(
        n410) );
  MUX U1413 ( .IN0(\Reg_Bank/registers[1][13] ), .IN1(n163), .SEL(n238), .F(
        \Reg_Bank/n3041 ) );
  NAND U1414 ( .A(n412), .B(n413), .Z(n163) );
  AND U1415 ( .A(n414), .B(n415), .Z(n413) );
  NANDN U1416 ( .B(n247), .A(\Data_Mem/N732 ), .Z(n415) );
  ANDN U1417 ( .A(n416), .B(n381), .Z(n414) );
  OR U1418 ( .A(n248), .B(n417), .Z(n416) );
  AND U1419 ( .A(n418), .B(n419), .Z(n412) );
  NANDN U1420 ( .B(n243), .A(pc_plus4[13]), .Z(n419) );
  AND U1421 ( .A(n420), .B(n421), .Z(n418) );
  NAND U1422 ( .A(n422), .B(n383), .Z(n421) );
  NAND U1423 ( .A(n422), .B(n397), .Z(n420) );
  MUX U1424 ( .IN0(\Data_Mem/N732 ), .IN1(\Data_Mem/N716 ), .SEL(n411), .F(
        n422) );
  MUX U1425 ( .IN0(\Reg_Bank/registers[1][12] ), .IN1(n164), .SEL(n238), .F(
        \Reg_Bank/n3040 ) );
  NAND U1426 ( .A(n423), .B(n424), .Z(n164) );
  AND U1427 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U1428 ( .B(n247), .A(\Data_Mem/N733 ), .Z(n426) );
  ANDN U1429 ( .A(n427), .B(n381), .Z(n425) );
  OR U1430 ( .A(n248), .B(n428), .Z(n427) );
  AND U1431 ( .A(n429), .B(n430), .Z(n423) );
  NANDN U1432 ( .B(n243), .A(pc_plus4[12]), .Z(n430) );
  AND U1433 ( .A(n431), .B(n432), .Z(n429) );
  NAND U1434 ( .A(n433), .B(n383), .Z(n432) );
  NAND U1435 ( .A(n433), .B(n397), .Z(n431) );
  MUX U1436 ( .IN0(\Data_Mem/N733 ), .IN1(\Data_Mem/N717 ), .SEL(n411), .F(
        n433) );
  MUX U1437 ( .IN0(\Reg_Bank/registers[1][11] ), .IN1(n165), .SEL(n238), .F(
        \Reg_Bank/n3039 ) );
  NAND U1438 ( .A(n434), .B(n435), .Z(n165) );
  AND U1439 ( .A(n436), .B(n437), .Z(n435) );
  NANDN U1440 ( .B(n247), .A(\Data_Mem/N734 ), .Z(n437) );
  ANDN U1441 ( .A(n438), .B(n381), .Z(n436) );
  OR U1442 ( .A(n248), .B(n439), .Z(n438) );
  AND U1443 ( .A(n440), .B(n441), .Z(n434) );
  NANDN U1444 ( .B(n243), .A(pc_plus4[11]), .Z(n441) );
  AND U1445 ( .A(n442), .B(n443), .Z(n440) );
  NAND U1446 ( .A(n444), .B(n383), .Z(n443) );
  NAND U1447 ( .A(n444), .B(n397), .Z(n442) );
  MUX U1448 ( .IN0(\Data_Mem/N734 ), .IN1(\Data_Mem/N718 ), .SEL(n411), .F(
        n444) );
  MUX U1449 ( .IN0(\Reg_Bank/registers[1][10] ), .IN1(n166), .SEL(n238), .F(
        \Reg_Bank/n3038 ) );
  NAND U1450 ( .A(n445), .B(n446), .Z(n166) );
  AND U1451 ( .A(n447), .B(n448), .Z(n446) );
  NANDN U1452 ( .B(n247), .A(\Data_Mem/N735 ), .Z(n448) );
  ANDN U1453 ( .A(n449), .B(n381), .Z(n447) );
  OR U1454 ( .A(n248), .B(n450), .Z(n449) );
  AND U1455 ( .A(n451), .B(n452), .Z(n445) );
  NANDN U1456 ( .B(n243), .A(pc_plus4[10]), .Z(n452) );
  AND U1457 ( .A(n453), .B(n454), .Z(n451) );
  NAND U1458 ( .A(n455), .B(n383), .Z(n454) );
  NAND U1459 ( .A(n455), .B(n397), .Z(n453) );
  MUX U1460 ( .IN0(\Data_Mem/N735 ), .IN1(\Data_Mem/N719 ), .SEL(n411), .F(
        n455) );
  MUX U1461 ( .IN0(\Reg_Bank/registers[1][9] ), .IN1(n167), .SEL(n238), .F(
        \Reg_Bank/n3037 ) );
  NAND U1462 ( .A(n456), .B(n457), .Z(n167) );
  AND U1463 ( .A(n458), .B(n459), .Z(n457) );
  NANDN U1464 ( .B(n247), .A(\Data_Mem/N736 ), .Z(n459) );
  ANDN U1465 ( .A(n460), .B(n381), .Z(n458) );
  OR U1466 ( .A(n248), .B(n461), .Z(n460) );
  AND U1467 ( .A(n462), .B(n463), .Z(n456) );
  NANDN U1468 ( .B(n243), .A(pc_plus4[9]), .Z(n463) );
  AND U1469 ( .A(n464), .B(n465), .Z(n462) );
  NAND U1470 ( .A(n466), .B(n383), .Z(n465) );
  NAND U1471 ( .A(n466), .B(n397), .Z(n464) );
  MUX U1472 ( .IN0(\Data_Mem/N736 ), .IN1(\Data_Mem/N720 ), .SEL(n411), .F(
        n466) );
  MUX U1473 ( .IN0(\Reg_Bank/registers[1][8] ), .IN1(n168), .SEL(n238), .F(
        \Reg_Bank/n3036 ) );
  NAND U1474 ( .A(n467), .B(n468), .Z(n168) );
  AND U1475 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U1476 ( .B(n247), .A(\Data_Mem/N737 ), .Z(n470) );
  ANDN U1477 ( .A(n471), .B(n381), .Z(n469) );
  AND U1478 ( .A(n472), .B(\Data_Mem/N738 ), .Z(n381) );
  OR U1479 ( .A(n248), .B(n473), .Z(n471) );
  AND U1480 ( .A(n474), .B(n475), .Z(n467) );
  NANDN U1481 ( .B(n243), .A(pc_plus4[8]), .Z(n475) );
  AND U1482 ( .A(n476), .B(n477), .Z(n474) );
  NAND U1483 ( .A(n478), .B(n383), .Z(n477) );
  NAND U1484 ( .A(n478), .B(n397), .Z(n476) );
  MUX U1485 ( .IN0(\Data_Mem/N737 ), .IN1(\Data_Mem/N721 ), .SEL(n411), .F(
        n478) );
  MUX U1486 ( .IN0(\Reg_Bank/registers[1][7] ), .IN1(n169), .SEL(n238), .F(
        \Reg_Bank/n3035 ) );
  NAND U1487 ( .A(n479), .B(n480), .Z(n169) );
  AND U1488 ( .A(n481), .B(n482), .Z(n480) );
  AND U1489 ( .A(n483), .B(n484), .Z(n482) );
  OR U1490 ( .A(n248), .B(n485), .Z(n484) );
  NANDN U1491 ( .B(n247), .A(\Data_Mem/N738 ), .Z(n483) );
  AND U1492 ( .A(n486), .B(n487), .Z(n481) );
  NAND U1493 ( .A(n488), .B(n383), .Z(n487) );
  NANDN U1494 ( .B(n489), .A(n472), .Z(n486) );
  AND U1495 ( .A(n490), .B(n491), .Z(n479) );
  NANDN U1496 ( .B(n243), .A(pc_plus4[7]), .Z(n491) );
  AND U1497 ( .A(n492), .B(n493), .Z(n490) );
  OR U1498 ( .A(n494), .B(n489), .Z(n493) );
  AND U1499 ( .A(n495), .B(n496), .Z(n489) );
  AND U1500 ( .A(n497), .B(n498), .Z(n496) );
  NAND U1501 ( .A(\Data_Mem/N738 ), .B(n499), .Z(n498) );
  NAND U1502 ( .A(\Data_Mem/N730 ), .B(n500), .Z(n497) );
  AND U1503 ( .A(n501), .B(n502), .Z(n495) );
  NAND U1504 ( .A(\Data_Mem/N722 ), .B(n503), .Z(n502) );
  NAND U1505 ( .A(\Data_Mem/N714 ), .B(n504), .Z(n501) );
  NAND U1506 ( .A(n488), .B(n397), .Z(n492) );
  MUX U1507 ( .IN0(\Data_Mem/N738 ), .IN1(\Data_Mem/N722 ), .SEL(n411), .F(
        n488) );
  MUX U1508 ( .IN0(\Reg_Bank/registers[1][6] ), .IN1(n170), .SEL(n238), .F(
        \Reg_Bank/n3034 ) );
  NAND U1509 ( .A(n505), .B(n506), .Z(n170) );
  AND U1510 ( .A(n507), .B(n508), .Z(n506) );
  AND U1511 ( .A(n509), .B(n510), .Z(n508) );
  OR U1512 ( .A(n248), .B(n511), .Z(n510) );
  NANDN U1513 ( .B(n247), .A(\Data_Mem/N739 ), .Z(n509) );
  AND U1514 ( .A(n512), .B(n513), .Z(n507) );
  NAND U1515 ( .A(n514), .B(n383), .Z(n513) );
  NANDN U1516 ( .B(n515), .A(n472), .Z(n512) );
  AND U1517 ( .A(n516), .B(n517), .Z(n505) );
  NANDN U1518 ( .B(n243), .A(pc_plus4[6]), .Z(n517) );
  AND U1519 ( .A(n518), .B(n519), .Z(n516) );
  OR U1520 ( .A(n494), .B(n515), .Z(n519) );
  AND U1521 ( .A(n520), .B(n521), .Z(n515) );
  AND U1522 ( .A(n522), .B(n523), .Z(n521) );
  NAND U1523 ( .A(n499), .B(\Data_Mem/N739 ), .Z(n523) );
  NAND U1524 ( .A(\Data_Mem/N731 ), .B(n500), .Z(n522) );
  AND U1525 ( .A(n524), .B(n525), .Z(n520) );
  NAND U1526 ( .A(\Data_Mem/N723 ), .B(n503), .Z(n525) );
  NAND U1527 ( .A(\Data_Mem/N715 ), .B(n504), .Z(n524) );
  NAND U1528 ( .A(n514), .B(n397), .Z(n518) );
  MUX U1529 ( .IN0(\Data_Mem/N739 ), .IN1(\Data_Mem/N723 ), .SEL(n411), .F(
        n514) );
  MUX U1530 ( .IN0(\Reg_Bank/registers[1][5] ), .IN1(n171), .SEL(n238), .F(
        \Reg_Bank/n3033 ) );
  NAND U1531 ( .A(n526), .B(n527), .Z(n171) );
  AND U1532 ( .A(n528), .B(n529), .Z(n527) );
  AND U1533 ( .A(n530), .B(n531), .Z(n529) );
  OR U1534 ( .A(n248), .B(n532), .Z(n531) );
  NANDN U1535 ( .B(n247), .A(\Data_Mem/N740 ), .Z(n530) );
  AND U1536 ( .A(n533), .B(n534), .Z(n528) );
  NAND U1537 ( .A(n535), .B(n383), .Z(n534) );
  NANDN U1538 ( .B(n536), .A(n472), .Z(n533) );
  AND U1539 ( .A(n537), .B(n538), .Z(n526) );
  NANDN U1540 ( .B(n243), .A(pc_plus4[5]), .Z(n538) );
  AND U1541 ( .A(n539), .B(n540), .Z(n537) );
  OR U1542 ( .A(n494), .B(n536), .Z(n540) );
  AND U1543 ( .A(n541), .B(n542), .Z(n536) );
  AND U1544 ( .A(n543), .B(n544), .Z(n542) );
  NAND U1545 ( .A(n499), .B(\Data_Mem/N740 ), .Z(n544) );
  NAND U1546 ( .A(\Data_Mem/N732 ), .B(n500), .Z(n543) );
  AND U1547 ( .A(n545), .B(n546), .Z(n541) );
  NAND U1548 ( .A(\Data_Mem/N724 ), .B(n503), .Z(n546) );
  NAND U1549 ( .A(\Data_Mem/N716 ), .B(n504), .Z(n545) );
  NAND U1550 ( .A(n535), .B(n397), .Z(n539) );
  MUX U1551 ( .IN0(\Data_Mem/N740 ), .IN1(\Data_Mem/N724 ), .SEL(n411), .F(
        n535) );
  MUX U1552 ( .IN0(\Reg_Bank/registers[1][4] ), .IN1(n172), .SEL(n238), .F(
        \Reg_Bank/n3032 ) );
  NAND U1553 ( .A(n547), .B(n548), .Z(n172) );
  AND U1554 ( .A(n549), .B(n550), .Z(n548) );
  AND U1555 ( .A(n551), .B(n552), .Z(n550) );
  OR U1556 ( .A(n248), .B(n553), .Z(n552) );
  NANDN U1557 ( .B(n247), .A(\Data_Mem/N741 ), .Z(n551) );
  AND U1558 ( .A(n554), .B(n555), .Z(n549) );
  NAND U1559 ( .A(n556), .B(n383), .Z(n555) );
  NANDN U1560 ( .B(n557), .A(n472), .Z(n554) );
  AND U1561 ( .A(n558), .B(n559), .Z(n547) );
  NANDN U1562 ( .B(n243), .A(pc_plus4[4]), .Z(n559) );
  AND U1563 ( .A(n560), .B(n561), .Z(n558) );
  OR U1564 ( .A(n494), .B(n557), .Z(n561) );
  AND U1565 ( .A(n562), .B(n563), .Z(n557) );
  AND U1566 ( .A(n564), .B(n565), .Z(n563) );
  NAND U1567 ( .A(n499), .B(\Data_Mem/N741 ), .Z(n565) );
  NAND U1568 ( .A(\Data_Mem/N733 ), .B(n500), .Z(n564) );
  AND U1569 ( .A(n566), .B(n567), .Z(n562) );
  NAND U1570 ( .A(\Data_Mem/N725 ), .B(n503), .Z(n567) );
  NAND U1571 ( .A(\Data_Mem/N717 ), .B(n504), .Z(n566) );
  NAND U1572 ( .A(n556), .B(n397), .Z(n560) );
  MUX U1573 ( .IN0(\Data_Mem/N741 ), .IN1(\Data_Mem/N725 ), .SEL(n411), .F(
        n556) );
  MUX U1574 ( .IN0(\Reg_Bank/registers[1][3] ), .IN1(n173), .SEL(n238), .F(
        \Reg_Bank/n3031 ) );
  NAND U1575 ( .A(n568), .B(n569), .Z(n173) );
  AND U1576 ( .A(n570), .B(n571), .Z(n569) );
  AND U1577 ( .A(n572), .B(n573), .Z(n571) );
  OR U1578 ( .A(n248), .B(n574), .Z(n573) );
  NANDN U1579 ( .B(n247), .A(\Data_Mem/N742 ), .Z(n572) );
  AND U1580 ( .A(n575), .B(n576), .Z(n570) );
  NAND U1581 ( .A(n577), .B(n383), .Z(n576) );
  NANDN U1582 ( .B(n578), .A(n472), .Z(n575) );
  AND U1583 ( .A(n579), .B(n580), .Z(n568) );
  NANDN U1584 ( .B(n243), .A(pc_plus4[3]), .Z(n580) );
  AND U1585 ( .A(n581), .B(n582), .Z(n579) );
  OR U1586 ( .A(n494), .B(n578), .Z(n582) );
  AND U1587 ( .A(n583), .B(n584), .Z(n578) );
  AND U1588 ( .A(n585), .B(n586), .Z(n584) );
  NAND U1589 ( .A(n499), .B(\Data_Mem/N742 ), .Z(n586) );
  NAND U1590 ( .A(\Data_Mem/N734 ), .B(n500), .Z(n585) );
  AND U1591 ( .A(n587), .B(n588), .Z(n583) );
  NAND U1592 ( .A(\Data_Mem/N726 ), .B(n503), .Z(n588) );
  NAND U1593 ( .A(\Data_Mem/N718 ), .B(n504), .Z(n587) );
  NAND U1594 ( .A(n577), .B(n397), .Z(n581) );
  MUX U1595 ( .IN0(\Data_Mem/N742 ), .IN1(\Data_Mem/N726 ), .SEL(n411), .F(
        n577) );
  MUX U1596 ( .IN0(\Reg_Bank/registers[1][2] ), .IN1(n174), .SEL(n238), .F(
        \Reg_Bank/n3030 ) );
  NAND U1597 ( .A(n589), .B(n590), .Z(n174) );
  AND U1598 ( .A(n591), .B(n592), .Z(n590) );
  AND U1599 ( .A(n593), .B(n594), .Z(n592) );
  OR U1600 ( .A(n248), .B(n595), .Z(n594) );
  NANDN U1601 ( .B(n247), .A(\Data_Mem/N743 ), .Z(n593) );
  AND U1602 ( .A(n596), .B(n597), .Z(n591) );
  NAND U1603 ( .A(n598), .B(n383), .Z(n597) );
  NANDN U1604 ( .B(n599), .A(n472), .Z(n596) );
  AND U1605 ( .A(n600), .B(n601), .Z(n589) );
  NANDN U1606 ( .B(n243), .A(n602), .Z(n601) );
  NANDN U1607 ( .B(n377), .A(n378), .Z(n243) );
  AND U1608 ( .A(n603), .B(n604), .Z(n600) );
  OR U1609 ( .A(n494), .B(n599), .Z(n604) );
  AND U1610 ( .A(n605), .B(n606), .Z(n599) );
  AND U1611 ( .A(n607), .B(n608), .Z(n606) );
  NAND U1612 ( .A(n499), .B(\Data_Mem/N743 ), .Z(n608) );
  NAND U1613 ( .A(\Data_Mem/N735 ), .B(n500), .Z(n607) );
  AND U1614 ( .A(n609), .B(n610), .Z(n605) );
  NAND U1615 ( .A(\Data_Mem/N727 ), .B(n503), .Z(n610) );
  NAND U1616 ( .A(\Data_Mem/N719 ), .B(n504), .Z(n609) );
  NAND U1617 ( .A(n598), .B(n397), .Z(n603) );
  MUX U1618 ( .IN0(\Data_Mem/N743 ), .IN1(\Data_Mem/N727 ), .SEL(n411), .F(
        n598) );
  MUX U1619 ( .IN0(\Reg_Bank/registers[1][1] ), .IN1(n176), .SEL(n238), .F(
        \Reg_Bank/n3029 ) );
  NAND U1620 ( .A(n611), .B(n612), .Z(n176) );
  AND U1621 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U1622 ( .B(n615), .A(n472), .Z(n614) );
  AND U1623 ( .A(n616), .B(n617), .Z(n613) );
  NANDN U1624 ( .B(n247), .A(\Data_Mem/N744 ), .Z(n617) );
  NAND U1625 ( .A(n618), .B(n383), .Z(n616) );
  AND U1626 ( .A(n619), .B(n620), .Z(n611) );
  OR U1627 ( .A(n248), .B(n399), .Z(n620) );
  AND U1628 ( .A(n621), .B(n622), .Z(n619) );
  OR U1629 ( .A(n615), .B(n494), .Z(n622) );
  AND U1630 ( .A(n623), .B(n624), .Z(n615) );
  AND U1631 ( .A(n625), .B(n626), .Z(n624) );
  NAND U1632 ( .A(n499), .B(\Data_Mem/N744 ), .Z(n626) );
  NAND U1633 ( .A(\Data_Mem/N736 ), .B(n500), .Z(n625) );
  AND U1634 ( .A(n627), .B(n628), .Z(n623) );
  NAND U1635 ( .A(\Data_Mem/N728 ), .B(n503), .Z(n628) );
  NAND U1636 ( .A(\Data_Mem/N720 ), .B(n504), .Z(n627) );
  NAND U1637 ( .A(n618), .B(n397), .Z(n621) );
  MUX U1638 ( .IN0(\Data_Mem/N744 ), .IN1(\Data_Mem/N728 ), .SEL(n411), .F(
        n618) );
  MUX U1639 ( .IN0(\Reg_Bank/registers[1][0] ), .IN1(n177), .SEL(n238), .F(
        \Reg_Bank/n3028 ) );
  ANDN U1640 ( .A(n226), .B(n194), .Z(n238) );
  IV U1641 ( .A(n221), .Z(n194) );
  ANDN U1642 ( .A(n231), .B(n224), .Z(n221) );
  NAND U1643 ( .A(n629), .B(n630), .Z(n224) );
  AND U1644 ( .A(n631), .B(n632), .Z(n630) );
  OR U1645 ( .A(n633), .B(n49), .Z(n632) );
  NANDN U1646 ( .B(n6), .A(n634), .Z(n631) );
  NAND U1647 ( .A(n635), .B(n636), .Z(n634) );
  NANDN U1648 ( .B(n10), .A(n637), .Z(n636) );
  NAND U1649 ( .A(n638), .B(n639), .Z(n637) );
  AND U1650 ( .A(n640), .B(n641), .Z(n639) );
  NAND U1651 ( .A(n642), .B(n643), .Z(n641) );
  AND U1652 ( .A(imm[13]), .B(n644), .Z(n642) );
  AND U1653 ( .A(n645), .B(n646), .Z(n640) );
  NANDN U1654 ( .B(n647), .A(imm[13]), .Z(n646) );
  NANDN U1655 ( .B(n648), .A(imm[13]), .Z(n645) );
  AND U1656 ( .A(n649), .B(n650), .Z(n638) );
  NANDN U1657 ( .B(n651), .A(n652), .Z(n650) );
  AND U1658 ( .A(imm[13]), .B(n653), .Z(n652) );
  NAND U1659 ( .A(n654), .B(n113), .Z(n649) );
  NANDN U1660 ( .B(n114), .A(n655), .Z(n654) );
  NANDN U1661 ( .B(n656), .A(imm[13]), .Z(n655) );
  AND U1662 ( .A(n657), .B(n658), .Z(n629) );
  NAND U1663 ( .A(n103), .B(n659), .Z(n658) );
  MUX U1664 ( .IN0(opcode[18]), .IN1(imm[13]), .SEL(opcode[23]), .F(n659) );
  NANDN U1665 ( .B(n660), .A(n661), .Z(n657) );
  ANDN U1666 ( .A(n662), .B(n49), .Z(n661) );
  ANDN U1667 ( .A(n236), .B(n234), .Z(n231) );
  NAND U1668 ( .A(n663), .B(n664), .Z(n234) );
  AND U1669 ( .A(n665), .B(n666), .Z(n664) );
  OR U1670 ( .A(n633), .B(n65), .Z(n666) );
  NANDN U1671 ( .B(n6), .A(n667), .Z(n665) );
  NAND U1672 ( .A(n668), .B(n669), .Z(n667) );
  ANDN U1673 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U1674 ( .B(n10), .A(n672), .Z(n670) );
  NAND U1675 ( .A(n673), .B(n674), .Z(n672) );
  AND U1676 ( .A(n675), .B(n676), .Z(n674) );
  NAND U1677 ( .A(n677), .B(n643), .Z(n676) );
  AND U1678 ( .A(n644), .B(imm[12]), .Z(n677) );
  AND U1679 ( .A(n678), .B(n679), .Z(n675) );
  NANDN U1680 ( .B(n647), .A(imm[12]), .Z(n679) );
  NANDN U1681 ( .B(n648), .A(imm[12]), .Z(n678) );
  AND U1682 ( .A(n680), .B(n681), .Z(n673) );
  NANDN U1683 ( .B(n651), .A(n682), .Z(n681) );
  AND U1684 ( .A(n653), .B(imm[12]), .Z(n682) );
  NAND U1685 ( .A(n683), .B(n113), .Z(n680) );
  NANDN U1686 ( .B(n114), .A(n684), .Z(n683) );
  NANDN U1687 ( .B(n656), .A(imm[12]), .Z(n684) );
  AND U1688 ( .A(n685), .B(n686), .Z(n663) );
  NAND U1689 ( .A(n103), .B(n687), .Z(n686) );
  MUX U1690 ( .IN0(opcode[17]), .IN1(imm[12]), .SEL(opcode[23]), .F(n687) );
  NANDN U1691 ( .B(n660), .A(n688), .Z(n685) );
  ANDN U1692 ( .A(n662), .B(n65), .Z(n688) );
  IV U1693 ( .A(n233), .Z(n236) );
  AND U1694 ( .A(n689), .B(n690), .Z(n233) );
  AND U1695 ( .A(n691), .B(n692), .Z(n690) );
  OR U1696 ( .A(n633), .B(n81), .Z(n692) );
  NANDN U1697 ( .B(n6), .A(n693), .Z(n691) );
  NAND U1698 ( .A(n635), .B(n694), .Z(n693) );
  NANDN U1699 ( .B(n10), .A(n695), .Z(n694) );
  NAND U1700 ( .A(n696), .B(n697), .Z(n695) );
  AND U1701 ( .A(n698), .B(n699), .Z(n697) );
  NAND U1702 ( .A(n700), .B(n643), .Z(n699) );
  AND U1703 ( .A(n644), .B(imm[11]), .Z(n700) );
  AND U1704 ( .A(n701), .B(n702), .Z(n698) );
  NANDN U1705 ( .B(n647), .A(imm[11]), .Z(n702) );
  NANDN U1706 ( .B(n648), .A(imm[11]), .Z(n701) );
  AND U1707 ( .A(n703), .B(n704), .Z(n696) );
  NANDN U1708 ( .B(n651), .A(n705), .Z(n704) );
  AND U1709 ( .A(n653), .B(imm[11]), .Z(n705) );
  NANDN U1710 ( .B(n656), .A(n706), .Z(n703) );
  AND U1711 ( .A(n113), .B(imm[11]), .Z(n706) );
  AND U1712 ( .A(n707), .B(n708), .Z(n689) );
  NAND U1713 ( .A(n103), .B(n709), .Z(n708) );
  MUX U1714 ( .IN0(opcode[16]), .IN1(imm[11]), .SEL(opcode[23]), .F(n709) );
  NANDN U1715 ( .B(n660), .A(n710), .Z(n707) );
  ANDN U1716 ( .A(n662), .B(n81), .Z(n710) );
  ANDN U1717 ( .A(n198), .B(n197), .Z(n226) );
  NAND U1718 ( .A(n711), .B(n712), .Z(n197) );
  AND U1719 ( .A(n713), .B(n714), .Z(n712) );
  NANDN U1720 ( .B(n633), .A(opcode[20]), .Z(n714) );
  NANDN U1721 ( .B(n6), .A(n715), .Z(n713) );
  NAND U1722 ( .A(n635), .B(n716), .Z(n715) );
  NANDN U1723 ( .B(n10), .A(n717), .Z(n716) );
  NAND U1724 ( .A(n718), .B(n719), .Z(n717) );
  AND U1725 ( .A(n720), .B(n721), .Z(n719) );
  NAND U1726 ( .A(n722), .B(n643), .Z(n721) );
  AND U1727 ( .A(n644), .B(imm[15]), .Z(n722) );
  AND U1728 ( .A(n723), .B(n724), .Z(n720) );
  NANDN U1729 ( .B(n647), .A(imm[15]), .Z(n724) );
  NANDN U1730 ( .B(n648), .A(imm[15]), .Z(n723) );
  AND U1731 ( .A(n725), .B(n726), .Z(n718) );
  NANDN U1732 ( .B(n651), .A(n727), .Z(n726) );
  AND U1733 ( .A(n653), .B(imm[15]), .Z(n727) );
  NANDN U1734 ( .B(n656), .A(n728), .Z(n725) );
  AND U1735 ( .A(n113), .B(imm[15]), .Z(n728) );
  AND U1736 ( .A(n729), .B(n730), .Z(n711) );
  NAND U1737 ( .A(n103), .B(n731), .Z(n730) );
  MUX U1738 ( .IN0(opcode[20]), .IN1(imm[15]), .SEL(opcode[23]), .F(n731) );
  NANDN U1739 ( .B(n660), .A(n732), .Z(n729) );
  AND U1740 ( .A(n662), .B(opcode[20]), .Z(n732) );
  AND U1741 ( .A(n733), .B(n734), .Z(n198) );
  AND U1742 ( .A(n735), .B(n736), .Z(n734) );
  OR U1743 ( .A(n633), .B(n23), .Z(n736) );
  NANDN U1744 ( .B(n6), .A(n737), .Z(n735) );
  NAND U1745 ( .A(n635), .B(n738), .Z(n737) );
  NANDN U1746 ( .B(n10), .A(n739), .Z(n738) );
  NAND U1747 ( .A(n740), .B(n741), .Z(n739) );
  AND U1748 ( .A(n742), .B(n743), .Z(n741) );
  NAND U1749 ( .A(n744), .B(n643), .Z(n743) );
  ANDN U1750 ( .A(n350), .B(imm[5]), .Z(n643) );
  AND U1751 ( .A(n644), .B(imm[14]), .Z(n744) );
  NANDN U1752 ( .B(n745), .A(n746), .Z(n644) );
  OR U1753 ( .A(n747), .B(imm[0]), .Z(n746) );
  AND U1754 ( .A(n748), .B(n749), .Z(n742) );
  NANDN U1755 ( .B(n647), .A(imm[14]), .Z(n749) );
  NANDN U1756 ( .B(n648), .A(imm[14]), .Z(n748) );
  NAND U1757 ( .A(n750), .B(n751), .Z(n648) );
  OR U1758 ( .A(n752), .B(imm[1]), .Z(n750) );
  AND U1759 ( .A(n753), .B(n754), .Z(n740) );
  NANDN U1760 ( .B(n651), .A(n755), .Z(n754) );
  AND U1761 ( .A(n653), .B(imm[14]), .Z(n755) );
  OR U1762 ( .A(n756), .B(n745), .Z(n653) );
  NAND U1763 ( .A(n757), .B(n113), .Z(n753) );
  NANDN U1764 ( .B(n114), .A(n758), .Z(n757) );
  NANDN U1765 ( .B(n656), .A(imm[14]), .Z(n758) );
  AND U1766 ( .A(n759), .B(n760), .Z(n733) );
  NAND U1767 ( .A(n103), .B(n761), .Z(n760) );
  MUX U1768 ( .IN0(opcode[19]), .IN1(imm[14]), .SEL(opcode[23]), .F(n761) );
  NOR U1769 ( .A(n10), .B(n762), .Z(n103) );
  NAND U1770 ( .A(n26), .B(n124), .Z(n762) );
  ANDN U1771 ( .A(n127), .B(n126), .Z(n124) );
  NANDN U1772 ( .B(n660), .A(n763), .Z(n759) );
  ANDN U1773 ( .A(n662), .B(n23), .Z(n763) );
  NAND U1774 ( .A(n764), .B(n765), .Z(n177) );
  AND U1775 ( .A(n766), .B(n767), .Z(n765) );
  NANDN U1776 ( .B(n768), .A(n472), .Z(n767) );
  ANDN U1777 ( .A(n769), .B(n770), .Z(n472) );
  AND U1778 ( .A(n771), .B(n772), .Z(n766) );
  NANDN U1779 ( .B(n247), .A(\Data_Mem/N745 ), .Z(n772) );
  NANDN U1780 ( .B(n773), .A(n774), .Z(n247) );
  NAND U1781 ( .A(n775), .B(n383), .Z(n771) );
  ANDN U1782 ( .A(n769), .B(n776), .Z(n383) );
  AND U1783 ( .A(n777), .B(n778), .Z(n764) );
  NANDN U1784 ( .B(n248), .A(n779), .Z(n778) );
  NANDN U1785 ( .B(n378), .A(n377), .Z(n248) );
  NAND U1786 ( .A(n780), .B(n781), .Z(n377) );
  ANDN U1787 ( .A(n132), .B(n130), .Z(n781) );
  AND U1788 ( .A(n782), .B(n783), .Z(n780) );
  NANDN U1789 ( .B(n6), .A(n784), .Z(n783) );
  NAND U1790 ( .A(n785), .B(n786), .Z(n784) );
  AND U1791 ( .A(n787), .B(n788), .Z(n786) );
  NANDN U1792 ( .B(n18), .A(n789), .Z(n788) );
  NANDN U1793 ( .B(n790), .A(n22), .Z(n789) );
  NOR U1794 ( .A(n791), .B(n792), .Z(n787) );
  AND U1795 ( .A(n793), .B(n794), .Z(n785) );
  NANDN U1796 ( .B(n10), .A(n795), .Z(n794) );
  NAND U1797 ( .A(n796), .B(n15), .Z(n795) );
  NOR U1798 ( .A(imm[1]), .B(n797), .Z(n796) );
  NAND U1799 ( .A(n798), .B(n799), .Z(n378) );
  NANDN U1800 ( .B(n6), .A(n800), .Z(n799) );
  NAND U1801 ( .A(n635), .B(n801), .Z(n800) );
  NAND U1802 ( .A(n802), .B(n113), .Z(n801) );
  ANDN U1803 ( .A(n803), .B(n10), .Z(n802) );
  NANDN U1804 ( .B(n114), .A(n656), .Z(n803) );
  ANDN U1805 ( .A(n669), .B(n671), .Z(n635) );
  NANDN U1806 ( .B(n790), .A(n804), .Z(n669) );
  NOR U1807 ( .A(n18), .B(n805), .Z(n804) );
  NANDN U1808 ( .B(opcode[19]), .A(opcode[20]), .Z(n790) );
  OR U1809 ( .A(n633), .B(n806), .Z(n798) );
  AND U1810 ( .A(n807), .B(n808), .Z(n777) );
  OR U1811 ( .A(n768), .B(n494), .Z(n808) );
  NANDN U1812 ( .B(n809), .A(n810), .Z(n494) );
  ANDN U1813 ( .A(n774), .B(n769), .Z(n810) );
  AND U1814 ( .A(n811), .B(n812), .Z(n768) );
  AND U1815 ( .A(n813), .B(n814), .Z(n812) );
  NAND U1816 ( .A(n499), .B(\Data_Mem/N745 ), .Z(n814) );
  NAND U1817 ( .A(\Data_Mem/N737 ), .B(n500), .Z(n813) );
  AND U1818 ( .A(n815), .B(n816), .Z(n811) );
  NAND U1819 ( .A(\Data_Mem/N729 ), .B(n503), .Z(n816) );
  NAND U1820 ( .A(\Data_Mem/N721 ), .B(n504), .Z(n815) );
  NAND U1821 ( .A(n775), .B(n397), .Z(n807) );
  ANDN U1822 ( .A(n817), .B(n776), .Z(n397) );
  NANDN U1823 ( .B(n774), .A(n773), .Z(n776) );
  IV U1824 ( .A(n809), .Z(n773) );
  IV U1825 ( .A(n769), .Z(n817) );
  ANDN U1826 ( .A(n134), .B(n818), .Z(n769) );
  NAND U1827 ( .A(n819), .B(n385), .Z(n775) );
  NANDN U1828 ( .B(n399), .A(\Data_Mem/N729 ), .Z(n385) );
  NANDN U1829 ( .B(n411), .A(\Data_Mem/N745 ), .Z(n819) );
  NAND U1830 ( .A(n820), .B(n821), .Z(\PC_Next/pc_future[9] ) );
  AND U1831 ( .A(n822), .B(n823), .Z(n821) );
  NANDN U1832 ( .B(n824), .A(pc_plus4[9]), .Z(n823) );
  NANDN U1833 ( .B(n825), .A(imm[7]), .Z(n822) );
  AND U1834 ( .A(n826), .B(n827), .Z(n820) );
  NAND U1835 ( .A(n828), .B(n829), .Z(n827) );
  MUX U1836 ( .IN0(\PC_Next/pc_jump[9] ), .IN1(pc_plus4[9]), .SEL(n830), .F(
        n828) );
  NANDN U1837 ( .B(n461), .A(n831), .Z(n826) );
  IV U1838 ( .A(n832), .Z(n461) );
  NAND U1839 ( .A(n833), .B(n834), .Z(\PC_Next/pc_future[8] ) );
  AND U1840 ( .A(n835), .B(n836), .Z(n834) );
  NANDN U1841 ( .B(n824), .A(pc_plus4[8]), .Z(n836) );
  NANDN U1842 ( .B(n825), .A(imm[6]), .Z(n835) );
  AND U1843 ( .A(n837), .B(n838), .Z(n833) );
  NAND U1844 ( .A(n839), .B(n829), .Z(n838) );
  MUX U1845 ( .IN0(\PC_Next/pc_jump[8] ), .IN1(pc_plus4[8]), .SEL(n830), .F(
        n839) );
  NANDN U1846 ( .B(n473), .A(n831), .Z(n837) );
  NAND U1847 ( .A(n840), .B(n841), .Z(\PC_Next/pc_future[7] ) );
  AND U1848 ( .A(n842), .B(n843), .Z(n841) );
  NANDN U1849 ( .B(n824), .A(pc_plus4[7]), .Z(n843) );
  NANDN U1850 ( .B(n825), .A(imm[5]), .Z(n842) );
  AND U1851 ( .A(n844), .B(n845), .Z(n840) );
  NAND U1852 ( .A(n846), .B(n829), .Z(n845) );
  MUX U1853 ( .IN0(\PC_Next/pc_jump[7] ), .IN1(pc_plus4[7]), .SEL(n830), .F(
        n846) );
  NANDN U1854 ( .B(n485), .A(n831), .Z(n844) );
  NAND U1855 ( .A(n847), .B(n848), .Z(\PC_Next/pc_future[6] ) );
  AND U1856 ( .A(n849), .B(n850), .Z(n848) );
  NANDN U1857 ( .B(n824), .A(pc_plus4[6]), .Z(n850) );
  OR U1858 ( .A(n825), .B(n341), .Z(n849) );
  AND U1859 ( .A(n851), .B(n852), .Z(n847) );
  NAND U1860 ( .A(n853), .B(n829), .Z(n852) );
  MUX U1861 ( .IN0(\PC_Next/pc_jump[6] ), .IN1(pc_plus4[6]), .SEL(n830), .F(
        n853) );
  NANDN U1862 ( .B(n511), .A(n831), .Z(n851) );
  NAND U1863 ( .A(n854), .B(n855), .Z(\PC_Next/pc_future[5] ) );
  AND U1864 ( .A(n856), .B(n857), .Z(n855) );
  NANDN U1865 ( .B(n824), .A(pc_plus4[5]), .Z(n857) );
  OR U1866 ( .A(n825), .B(n350), .Z(n856) );
  AND U1867 ( .A(n858), .B(n859), .Z(n854) );
  NAND U1868 ( .A(n860), .B(n829), .Z(n859) );
  MUX U1869 ( .IN0(\PC_Next/pc_jump[5] ), .IN1(pc_plus4[5]), .SEL(n830), .F(
        n860) );
  NANDN U1870 ( .B(n532), .A(n831), .Z(n858) );
  NAND U1871 ( .A(n861), .B(n862), .Z(\PC_Next/pc_future[4] ) );
  AND U1872 ( .A(n863), .B(n864), .Z(n862) );
  NANDN U1873 ( .B(n824), .A(pc_plus4[4]), .Z(n864) );
  OR U1874 ( .A(n825), .B(n359), .Z(n863) );
  AND U1875 ( .A(n865), .B(n866), .Z(n861) );
  NAND U1876 ( .A(n867), .B(n829), .Z(n866) );
  MUX U1877 ( .IN0(\PC_Next/pc_jump[4] ), .IN1(pc_plus4[4]), .SEL(n830), .F(
        n867) );
  NANDN U1878 ( .B(n553), .A(n831), .Z(n865) );
  NAND U1879 ( .A(n868), .B(n869), .Z(\PC_Next/pc_future[3] ) );
  AND U1880 ( .A(n870), .B(n871), .Z(n869) );
  NANDN U1881 ( .B(n824), .A(pc_plus4[3]), .Z(n871) );
  OR U1882 ( .A(n825), .B(n14), .Z(n870) );
  AND U1883 ( .A(n872), .B(n873), .Z(n868) );
  NAND U1884 ( .A(n874), .B(n829), .Z(n873) );
  MUX U1885 ( .IN0(\PC_Next/pc_jump[3] ), .IN1(pc_plus4[3]), .SEL(n830), .F(
        n874) );
  NANDN U1886 ( .B(n574), .A(n831), .Z(n872) );
  NAND U1887 ( .A(n875), .B(n876), .Z(\PC_Next/pc_future[2] ) );
  AND U1888 ( .A(n877), .B(n878), .Z(n876) );
  OR U1889 ( .A(n824), .B(pc_current[2]), .Z(n878) );
  OR U1890 ( .A(n825), .B(n376), .Z(n877) );
  AND U1891 ( .A(n879), .B(n880), .Z(n875) );
  NAND U1892 ( .A(n881), .B(n829), .Z(n880) );
  MUX U1893 ( .IN0(\PC_Next/pc_jump[2] ), .IN1(n602), .SEL(n830), .F(n881) );
  IV U1894 ( .A(pc_current[2]), .Z(n602) );
  NANDN U1895 ( .B(n595), .A(n831), .Z(n879) );
  NAND U1896 ( .A(n882), .B(n883), .Z(\PC_Next/pc_future[27] ) );
  AND U1897 ( .A(n884), .B(n885), .Z(n883) );
  NANDN U1898 ( .B(n824), .A(pc_plus4[27]), .Z(n885) );
  OR U1899 ( .A(n825), .B(n886), .Z(n884) );
  AND U1900 ( .A(n887), .B(n888), .Z(n882) );
  NAND U1901 ( .A(n889), .B(n829), .Z(n888) );
  MUX U1902 ( .IN0(\PC_Next/pc_jump[27] ), .IN1(pc_plus4[27]), .SEL(n830), .F(
        n889) );
  NANDN U1903 ( .B(n283), .A(n831), .Z(n887) );
  NAND U1904 ( .A(n890), .B(n891), .Z(\PC_Next/pc_future[26] ) );
  AND U1905 ( .A(n892), .B(n893), .Z(n891) );
  NANDN U1906 ( .B(n824), .A(pc_plus4[26]), .Z(n893) );
  NANDN U1907 ( .B(n825), .A(opcode[24]), .Z(n892) );
  AND U1908 ( .A(n894), .B(n895), .Z(n890) );
  NAND U1909 ( .A(n896), .B(n829), .Z(n895) );
  MUX U1910 ( .IN0(\PC_Next/pc_jump[26] ), .IN1(pc_plus4[26]), .SEL(n830), .F(
        n896) );
  NANDN U1911 ( .B(n291), .A(n831), .Z(n894) );
  NAND U1912 ( .A(n897), .B(n898), .Z(\PC_Next/pc_future[25] ) );
  AND U1913 ( .A(n899), .B(n900), .Z(n898) );
  NANDN U1914 ( .B(n824), .A(pc_plus4[25]), .Z(n900) );
  OR U1915 ( .A(n825), .B(n125), .Z(n899) );
  IV U1916 ( .A(opcode[23]), .Z(n125) );
  AND U1917 ( .A(n901), .B(n902), .Z(n897) );
  NAND U1918 ( .A(n903), .B(n829), .Z(n902) );
  MUX U1919 ( .IN0(\PC_Next/pc_jump[25] ), .IN1(pc_plus4[25]), .SEL(n830), .F(
        n903) );
  NANDN U1920 ( .B(n299), .A(n831), .Z(n901) );
  NAND U1921 ( .A(n904), .B(n905), .Z(\PC_Next/pc_future[24] ) );
  AND U1922 ( .A(n906), .B(n907), .Z(n905) );
  NANDN U1923 ( .B(n824), .A(pc_plus4[24]), .Z(n907) );
  OR U1924 ( .A(n825), .B(n908), .Z(n906) );
  AND U1925 ( .A(n909), .B(n910), .Z(n904) );
  NAND U1926 ( .A(n911), .B(n829), .Z(n910) );
  MUX U1927 ( .IN0(\PC_Next/pc_jump[24] ), .IN1(pc_plus4[24]), .SEL(n830), .F(
        n911) );
  NANDN U1928 ( .B(n307), .A(n831), .Z(n909) );
  NAND U1929 ( .A(n912), .B(n913), .Z(\PC_Next/pc_future[23] ) );
  AND U1930 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U1931 ( .B(n824), .A(pc_plus4[23]), .Z(n915) );
  NANDN U1932 ( .B(n825), .A(opcode[21]), .Z(n914) );
  AND U1933 ( .A(n916), .B(n917), .Z(n912) );
  NAND U1934 ( .A(n918), .B(n829), .Z(n917) );
  MUX U1935 ( .IN0(\PC_Next/pc_jump[23] ), .IN1(pc_plus4[23]), .SEL(n830), .F(
        n918) );
  NANDN U1936 ( .B(n315), .A(n831), .Z(n916) );
  NAND U1937 ( .A(n919), .B(n920), .Z(\PC_Next/pc_future[22] ) );
  AND U1938 ( .A(n921), .B(n922), .Z(n920) );
  NANDN U1939 ( .B(n824), .A(pc_plus4[22]), .Z(n922) );
  NANDN U1940 ( .B(n825), .A(opcode[20]), .Z(n921) );
  AND U1941 ( .A(n923), .B(n924), .Z(n919) );
  NAND U1942 ( .A(n925), .B(n829), .Z(n924) );
  MUX U1943 ( .IN0(\PC_Next/pc_jump[22] ), .IN1(pc_plus4[22]), .SEL(n830), .F(
        n925) );
  NANDN U1944 ( .B(n323), .A(n831), .Z(n923) );
  NAND U1945 ( .A(n926), .B(n927), .Z(\PC_Next/pc_future[21] ) );
  AND U1946 ( .A(n928), .B(n929), .Z(n927) );
  NANDN U1947 ( .B(n824), .A(pc_plus4[21]), .Z(n929) );
  OR U1948 ( .A(n825), .B(n23), .Z(n928) );
  AND U1949 ( .A(n930), .B(n931), .Z(n926) );
  NAND U1950 ( .A(n932), .B(n829), .Z(n931) );
  MUX U1951 ( .IN0(\PC_Next/pc_jump[21] ), .IN1(pc_plus4[21]), .SEL(n830), .F(
        n932) );
  NANDN U1952 ( .B(n331), .A(n831), .Z(n930) );
  NAND U1953 ( .A(n933), .B(n934), .Z(\PC_Next/pc_future[20] ) );
  AND U1954 ( .A(n935), .B(n936), .Z(n934) );
  NANDN U1955 ( .B(n824), .A(pc_plus4[20]), .Z(n936) );
  OR U1956 ( .A(n825), .B(n49), .Z(n935) );
  AND U1957 ( .A(n937), .B(n938), .Z(n933) );
  NAND U1958 ( .A(n939), .B(n829), .Z(n938) );
  MUX U1959 ( .IN0(\PC_Next/pc_jump[20] ), .IN1(pc_plus4[20]), .SEL(n830), .F(
        n939) );
  NANDN U1960 ( .B(n339), .A(n831), .Z(n937) );
  NAND U1961 ( .A(n940), .B(n941), .Z(\PC_Next/pc_future[19] ) );
  AND U1962 ( .A(n942), .B(n943), .Z(n941) );
  NANDN U1963 ( .B(n824), .A(pc_plus4[19]), .Z(n943) );
  OR U1964 ( .A(n825), .B(n65), .Z(n942) );
  AND U1965 ( .A(n944), .B(n945), .Z(n940) );
  NAND U1966 ( .A(n946), .B(n829), .Z(n945) );
  MUX U1967 ( .IN0(\PC_Next/pc_jump[19] ), .IN1(pc_plus4[19]), .SEL(n830), .F(
        n946) );
  NANDN U1968 ( .B(n348), .A(n831), .Z(n944) );
  NAND U1969 ( .A(n947), .B(n948), .Z(\PC_Next/pc_future[18] ) );
  AND U1970 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U1971 ( .B(n824), .A(pc_plus4[18]), .Z(n950) );
  OR U1972 ( .A(n825), .B(n81), .Z(n949) );
  AND U1973 ( .A(n951), .B(n952), .Z(n947) );
  NAND U1974 ( .A(n953), .B(n829), .Z(n952) );
  MUX U1975 ( .IN0(\PC_Next/pc_jump[18] ), .IN1(pc_plus4[18]), .SEL(n830), .F(
        n953) );
  NANDN U1976 ( .B(n357), .A(n831), .Z(n951) );
  NAND U1977 ( .A(n954), .B(n955), .Z(\PC_Next/pc_future[17] ) );
  AND U1978 ( .A(n956), .B(n957), .Z(n955) );
  NANDN U1979 ( .B(n824), .A(pc_plus4[17]), .Z(n957) );
  NANDN U1980 ( .B(n825), .A(imm[15]), .Z(n956) );
  AND U1981 ( .A(n958), .B(n959), .Z(n954) );
  NAND U1982 ( .A(n960), .B(n829), .Z(n959) );
  MUX U1983 ( .IN0(\PC_Next/pc_jump[17] ), .IN1(pc_plus4[17]), .SEL(n830), .F(
        n960) );
  NANDN U1984 ( .B(n366), .A(n831), .Z(n958) );
  NAND U1985 ( .A(n961), .B(n962), .Z(\PC_Next/pc_future[16] ) );
  AND U1986 ( .A(n963), .B(n964), .Z(n962) );
  NANDN U1987 ( .B(n824), .A(pc_plus4[16]), .Z(n964) );
  NANDN U1988 ( .B(n825), .A(imm[14]), .Z(n963) );
  AND U1989 ( .A(n965), .B(n966), .Z(n961) );
  NAND U1990 ( .A(n967), .B(n829), .Z(n966) );
  MUX U1991 ( .IN0(\PC_Next/pc_jump[16] ), .IN1(pc_plus4[16]), .SEL(n830), .F(
        n967) );
  NANDN U1992 ( .B(n374), .A(n831), .Z(n965) );
  NAND U1993 ( .A(n968), .B(n969), .Z(\PC_Next/pc_future[15] ) );
  AND U1994 ( .A(n970), .B(n971), .Z(n969) );
  NANDN U1995 ( .B(n824), .A(pc_plus4[15]), .Z(n971) );
  NANDN U1996 ( .B(n825), .A(imm[13]), .Z(n970) );
  AND U1997 ( .A(n972), .B(n973), .Z(n968) );
  NAND U1998 ( .A(n974), .B(n829), .Z(n973) );
  MUX U1999 ( .IN0(\PC_Next/pc_jump[15] ), .IN1(pc_plus4[15]), .SEL(n830), .F(
        n974) );
  NANDN U2000 ( .B(n391), .A(n831), .Z(n972) );
  NAND U2001 ( .A(n975), .B(n976), .Z(\PC_Next/pc_future[14] ) );
  AND U2002 ( .A(n977), .B(n978), .Z(n976) );
  NANDN U2003 ( .B(n824), .A(pc_plus4[14]), .Z(n978) );
  NANDN U2004 ( .B(n825), .A(imm[12]), .Z(n977) );
  AND U2005 ( .A(n979), .B(n980), .Z(n975) );
  NAND U2006 ( .A(n981), .B(n829), .Z(n980) );
  MUX U2007 ( .IN0(\PC_Next/pc_jump[14] ), .IN1(pc_plus4[14]), .SEL(n830), .F(
        n981) );
  NANDN U2008 ( .B(n405), .A(n831), .Z(n979) );
  NAND U2009 ( .A(n982), .B(n983), .Z(\PC_Next/pc_future[13] ) );
  AND U2010 ( .A(n984), .B(n985), .Z(n983) );
  NANDN U2011 ( .B(n824), .A(pc_plus4[13]), .Z(n985) );
  NANDN U2012 ( .B(n825), .A(imm[11]), .Z(n984) );
  AND U2013 ( .A(n986), .B(n987), .Z(n982) );
  NAND U2014 ( .A(n988), .B(n829), .Z(n987) );
  MUX U2015 ( .IN0(\PC_Next/pc_jump[13] ), .IN1(pc_plus4[13]), .SEL(n830), .F(
        n988) );
  NANDN U2016 ( .B(n417), .A(n831), .Z(n986) );
  NAND U2017 ( .A(n989), .B(n990), .Z(\PC_Next/pc_future[12] ) );
  AND U2018 ( .A(n991), .B(n992), .Z(n990) );
  NANDN U2019 ( .B(n824), .A(pc_plus4[12]), .Z(n992) );
  NANDN U2020 ( .B(n825), .A(imm[10]), .Z(n991) );
  AND U2021 ( .A(n993), .B(n994), .Z(n989) );
  NAND U2022 ( .A(n995), .B(n829), .Z(n994) );
  MUX U2023 ( .IN0(\PC_Next/pc_jump[12] ), .IN1(pc_plus4[12]), .SEL(n830), .F(
        n995) );
  NANDN U2024 ( .B(n428), .A(n831), .Z(n993) );
  NAND U2025 ( .A(n996), .B(n997), .Z(\PC_Next/pc_future[11] ) );
  AND U2026 ( .A(n998), .B(n999), .Z(n997) );
  NANDN U2027 ( .B(n824), .A(pc_plus4[11]), .Z(n999) );
  NANDN U2028 ( .B(n825), .A(imm[9]), .Z(n998) );
  AND U2029 ( .A(n1000), .B(n1001), .Z(n996) );
  NAND U2030 ( .A(n1002), .B(n829), .Z(n1001) );
  MUX U2031 ( .IN0(\PC_Next/pc_jump[11] ), .IN1(pc_plus4[11]), .SEL(n830), .F(
        n1002) );
  NANDN U2032 ( .B(n439), .A(n831), .Z(n1000) );
  NAND U2033 ( .A(n1003), .B(n1004), .Z(\PC_Next/pc_future[10] ) );
  AND U2034 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U2035 ( .B(n824), .A(pc_plus4[10]), .Z(n1006) );
  NANDN U2036 ( .B(n825), .A(imm[8]), .Z(n1005) );
  AND U2037 ( .A(n1007), .B(n1008), .Z(n1003) );
  NAND U2038 ( .A(n1009), .B(n829), .Z(n1008) );
  MUX U2039 ( .IN0(\PC_Next/pc_jump[10] ), .IN1(pc_plus4[10]), .SEL(n830), .F(
        n1009) );
  NANDN U2040 ( .B(n450), .A(n831), .Z(n1007) );
  NAND U2041 ( .A(n1010), .B(n1011), .Z(\PC_Next/n311 ) );
  AND U2042 ( .A(n1012), .B(n1013), .Z(n1011) );
  NANDN U2043 ( .B(n825), .A(pc_current[28]), .Z(n1013) );
  NANDN U2044 ( .B(n824), .A(pc_plus4[28]), .Z(n1012) );
  AND U2045 ( .A(n1014), .B(n1015), .Z(n1010) );
  NAND U2046 ( .A(n1016), .B(n829), .Z(n1015) );
  MUX U2047 ( .IN0(\PC_Next/pc_jump[28] ), .IN1(pc_plus4[28]), .SEL(n830), .F(
        n1016) );
  IV U2048 ( .A(n1017), .Z(n830) );
  NANDN U2049 ( .B(n275), .A(n831), .Z(n1014) );
  NAND U2050 ( .A(n1018), .B(n1019), .Z(\PC_Next/n310 ) );
  AND U2051 ( .A(n1020), .B(n1021), .Z(n1019) );
  NANDN U2052 ( .B(n825), .A(pc_current[29]), .Z(n1021) );
  NANDN U2053 ( .B(n824), .A(pc_plus4[29]), .Z(n1020) );
  AND U2054 ( .A(n1022), .B(n1023), .Z(n1018) );
  NAND U2055 ( .A(n1024), .B(n829), .Z(n1023) );
  MUX U2056 ( .IN0(pc_plus4[29]), .IN1(\PC_Next/pc_jump[29] ), .SEL(n1017), 
        .F(n1024) );
  NANDN U2057 ( .B(n267), .A(n831), .Z(n1022) );
  NAND U2058 ( .A(n1025), .B(n1026), .Z(\PC_Next/n309 ) );
  AND U2059 ( .A(n1027), .B(n1028), .Z(n1026) );
  NANDN U2060 ( .B(n825), .A(pc_current[30]), .Z(n1028) );
  NANDN U2061 ( .B(n824), .A(pc_plus4[30]), .Z(n1027) );
  AND U2062 ( .A(n1029), .B(n1030), .Z(n1025) );
  NAND U2063 ( .A(n1031), .B(n829), .Z(n1030) );
  MUX U2064 ( .IN0(pc_plus4[30]), .IN1(\PC_Next/pc_jump[30] ), .SEL(n1017), 
        .F(n1031) );
  NANDN U2065 ( .B(n259), .A(n831), .Z(n1029) );
  NAND U2066 ( .A(n1032), .B(n1033), .Z(\PC_Next/n308 ) );
  AND U2067 ( .A(n1034), .B(n1035), .Z(n1033) );
  NANDN U2068 ( .B(n825), .A(pc_current[31]), .Z(n1035) );
  NANDN U2069 ( .B(n1036), .A(n1037), .Z(n825) );
  NANDN U2070 ( .B(n824), .A(n244), .Z(n1034) );
  NANDN U2071 ( .B(n1038), .A(n1037), .Z(n824) );
  AND U2072 ( .A(n1039), .B(n1040), .Z(n1032) );
  NAND U2073 ( .A(n1041), .B(n829), .Z(n1040) );
  ANDN U2074 ( .A(n1036), .B(n1037), .Z(n829) );
  IV U2075 ( .A(n1038), .Z(n1036) );
  MUX U2076 ( .IN0(n244), .IN1(\PC_Next/pc_jump[31] ), .SEL(n1017), .F(n1041)
         );
  NAND U2077 ( .A(n1042), .B(n1043), .Z(n1017) );
  AND U2078 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U2079 ( .A(n1046), .B(n249), .Z(n1045) );
  MUX U2080 ( .IN0(n1047), .IN1(n1048), .SEL(n1049), .F(n1044) );
  NAND U2081 ( .A(n1050), .B(n1051), .Z(n1048) );
  AND U2082 ( .A(n1052), .B(n1053), .Z(n1042) );
  MUX U2083 ( .IN0(n1054), .IN1(n1047), .SEL(n1050), .F(n1053) );
  OR U2084 ( .A(n1055), .B(n1056), .Z(n1047) );
  NANDN U2085 ( .B(n1057), .A(n1058), .Z(n1055) );
  OR U2086 ( .A(n1046), .B(n1059), .Z(n1054) );
  OR U2087 ( .A(n1058), .B(n1057), .Z(n1046) );
  MUX U2088 ( .IN0(n1060), .IN1(n1061), .SEL(n1050), .F(n1052) );
  AND U2089 ( .A(n1062), .B(n1063), .Z(n1050) );
  ANDN U2090 ( .A(n1064), .B(n791), .Z(n1063) );
  ANDN U2091 ( .A(n806), .B(n792), .Z(n1064) );
  IV U2092 ( .A(n130), .Z(n806) );
  AND U2093 ( .A(n1065), .B(n1066), .Z(n1062) );
  AND U2094 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U2095 ( .B(n18), .A(n1069), .Z(n1068) );
  NANDN U2096 ( .B(opcode[19]), .A(n22), .Z(n1069) );
  ANDN U2097 ( .A(n65), .B(opcode[18]), .Z(n22) );
  IV U2098 ( .A(opcode[17]), .Z(n65) );
  NANDN U2099 ( .B(n10), .A(n1070), .Z(n1067) );
  NANDN U2100 ( .B(imm[1]), .A(n15), .Z(n1070) );
  ANDN U2101 ( .A(n1071), .B(n350), .Z(n15) );
  ANDN U2102 ( .A(n341), .B(n1072), .Z(n1071) );
  IV U2103 ( .A(n651), .Z(n1072) );
  NANDN U2104 ( .B(n1073), .A(n1058), .Z(n1061) );
  NANDN U2105 ( .B(n1049), .A(n1051), .Z(n1060) );
  ANDN U2106 ( .A(n1057), .B(n1058), .Z(n1051) );
  NAND U2107 ( .A(n1074), .B(n1075), .Z(n1058) );
  ANDN U2108 ( .A(n1076), .B(n1077), .Z(n1075) );
  ANDN U2109 ( .A(n10), .B(n130), .Z(n1076) );
  AND U2110 ( .A(n1065), .B(n1078), .Z(n1074) );
  ANDN U2111 ( .A(n1079), .B(n671), .Z(n1078) );
  NANDN U2112 ( .B(n18), .A(n1080), .Z(n1079) );
  NAND U2113 ( .A(n1081), .B(n1082), .Z(n1080) );
  ANDN U2114 ( .A(n49), .B(opcode[19]), .Z(n1082) );
  ANDN U2115 ( .A(n81), .B(opcode[17]), .Z(n1081) );
  IV U2116 ( .A(opcode[16]), .Z(n81) );
  IV U2117 ( .A(n1073), .Z(n1057) );
  AND U2118 ( .A(n1083), .B(n1084), .Z(n1073) );
  NOR U2119 ( .A(n792), .B(n1085), .Z(n1084) );
  ANDN U2120 ( .A(n1065), .B(n1086), .Z(n1083) );
  AND U2121 ( .A(n782), .B(n1087), .Z(n1065) );
  ANDN U2122 ( .A(n132), .B(n134), .Z(n1087) );
  NAND U2123 ( .A(opcode[31]), .B(opcode[30]), .Z(n132) );
  ANDN U2124 ( .A(n133), .B(n26), .Z(n782) );
  IV U2125 ( .A(n1059), .Z(n1049) );
  NAND U2126 ( .A(n1088), .B(n1089), .Z(n1059) );
  AND U2127 ( .A(n1090), .B(n1091), .Z(n1089) );
  AND U2128 ( .A(n1092), .B(n1093), .Z(n1091) );
  AND U2129 ( .A(n1094), .B(n1095), .Z(n1093) );
  ANDN U2130 ( .A(n595), .B(N28), .Z(n1095) );
  ANDN U2131 ( .A(n553), .B(N26), .Z(n1094) );
  AND U2132 ( .A(n1096), .B(n1097), .Z(n1092) );
  ANDN U2133 ( .A(n511), .B(N24), .Z(n1097) );
  NOR U2134 ( .A(n411), .B(n779), .Z(n1096) );
  AND U2135 ( .A(n1098), .B(n1099), .Z(n1090) );
  AND U2136 ( .A(n1100), .B(n1101), .Z(n1099) );
  ANDN U2137 ( .A(n473), .B(n832), .Z(n1101) );
  NAND U2138 ( .A(n1102), .B(n1103), .Z(n832) );
  AND U2139 ( .A(n1104), .B(n1105), .Z(n1103) );
  AND U2140 ( .A(n1106), .B(n1107), .Z(n1105) );
  NAND U2141 ( .A(n1108), .B(n1109), .Z(n1107) );
  NAND U2142 ( .A(n1110), .B(n1111), .Z(n1108) );
  AND U2143 ( .A(n1112), .B(n1113), .Z(n1111) );
  AND U2144 ( .A(n1114), .B(n1115), .Z(n1112) );
  OR U2145 ( .A(n1116), .B(n1117), .Z(n1115) );
  NAND U2146 ( .A(n1118), .B(n1119), .Z(n1114) );
  NAND U2147 ( .A(n1120), .B(n1121), .Z(n1106) );
  NAND U2148 ( .A(n1110), .B(n1122), .Z(n1120) );
  AND U2149 ( .A(n1123), .B(n1113), .Z(n1122) );
  NAND U2150 ( .A(n1124), .B(n1125), .Z(n1113) );
  AND U2151 ( .A(n1126), .B(n1127), .Z(n1123) );
  OR U2152 ( .A(n1128), .B(n1117), .Z(n1127) );
  NAND U2153 ( .A(n1129), .B(n1119), .Z(n1126) );
  AND U2154 ( .A(n1130), .B(n1131), .Z(n1110) );
  NAND U2155 ( .A(n1132), .B(n1133), .Z(n1131) );
  NAND U2156 ( .A(n1134), .B(n1135), .Z(n1130) );
  AND U2157 ( .A(n1136), .B(n1137), .Z(n1104) );
  NAND U2158 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][9] ), .Z(n1137) );
  NAND U2159 ( .A(n1139), .B(n1140), .Z(n1136) );
  XNOR U2160 ( .A(n1141), .B(n1142), .Z(n1139) );
  AND U2161 ( .A(n1143), .B(n1144), .Z(n1102) );
  MUX U2162 ( .IN0(n1145), .IN1(n1146), .SEL(n1147), .F(n1144) );
  ANDN U2163 ( .A(n1142), .B(b_bus[9]), .Z(n1147) );
  AND U2164 ( .A(n1148), .B(n1149), .Z(n1143) );
  NAND U2165 ( .A(n1150), .B(n1151), .Z(n1149) );
  XNOR U2166 ( .A(n1142), .B(b_bus[9]), .Z(n1150) );
  IV U2167 ( .A(n1152), .Z(b_bus[9]) );
  NANDN U2168 ( .B(n1142), .A(n1153), .Z(n1148) );
  ANDN U2169 ( .A(n1154), .B(n1152), .Z(n1153) );
  AND U2170 ( .A(n1155), .B(n1156), .Z(n473) );
  AND U2171 ( .A(n1157), .B(n1158), .Z(n1156) );
  AND U2172 ( .A(n1159), .B(n1160), .Z(n1158) );
  NAND U2173 ( .A(n1161), .B(n1109), .Z(n1160) );
  NAND U2174 ( .A(n1162), .B(n1163), .Z(n1161) );
  AND U2175 ( .A(n1164), .B(n1165), .Z(n1163) );
  AND U2176 ( .A(n1166), .B(n1167), .Z(n1164) );
  OR U2177 ( .A(n1168), .B(n1117), .Z(n1167) );
  NAND U2178 ( .A(n1169), .B(n1118), .Z(n1166) );
  NAND U2179 ( .A(n1170), .B(n1121), .Z(n1159) );
  NAND U2180 ( .A(n1162), .B(n1171), .Z(n1170) );
  AND U2181 ( .A(n1172), .B(n1165), .Z(n1171) );
  NAND U2182 ( .A(n1124), .B(n1173), .Z(n1165) );
  AND U2183 ( .A(n1174), .B(n1175), .Z(n1172) );
  OR U2184 ( .A(n1176), .B(n1117), .Z(n1175) );
  NAND U2185 ( .A(n1169), .B(n1129), .Z(n1174) );
  AND U2186 ( .A(n1177), .B(n1178), .Z(n1162) );
  NAND U2187 ( .A(n1179), .B(n1132), .Z(n1178) );
  NAND U2188 ( .A(n1180), .B(n1134), .Z(n1177) );
  AND U2189 ( .A(n1181), .B(n1182), .Z(n1157) );
  NAND U2190 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][8] ), .Z(n1182) );
  NAND U2191 ( .A(n1183), .B(n1140), .Z(n1181) );
  XNOR U2192 ( .A(n1184), .B(n1185), .Z(n1183) );
  AND U2193 ( .A(n1186), .B(n1187), .Z(n1155) );
  MUX U2194 ( .IN0(n1145), .IN1(n1146), .SEL(n1188), .F(n1187) );
  ANDN U2195 ( .A(n1185), .B(b_bus[8]), .Z(n1188) );
  AND U2196 ( .A(n1189), .B(n1190), .Z(n1186) );
  NAND U2197 ( .A(n1191), .B(n1151), .Z(n1190) );
  XNOR U2198 ( .A(n1185), .B(b_bus[8]), .Z(n1191) );
  IV U2199 ( .A(n1192), .Z(b_bus[8]) );
  NANDN U2200 ( .B(n1185), .A(n1193), .Z(n1189) );
  ANDN U2201 ( .A(n1154), .B(n1192), .Z(n1193) );
  ANDN U2202 ( .A(n450), .B(n1194), .Z(n1100) );
  IV U2203 ( .A(n439), .Z(n1194) );
  AND U2204 ( .A(n1195), .B(n1196), .Z(n439) );
  AND U2205 ( .A(n1197), .B(n1198), .Z(n1196) );
  AND U2206 ( .A(n1199), .B(n1200), .Z(n1198) );
  NAND U2207 ( .A(n1201), .B(n1109), .Z(n1200) );
  NAND U2208 ( .A(n1202), .B(n1203), .Z(n1201) );
  AND U2209 ( .A(n1204), .B(n1205), .Z(n1203) );
  AND U2210 ( .A(n1206), .B(n1207), .Z(n1204) );
  NANDN U2211 ( .B(n1117), .A(n1208), .Z(n1207) );
  NAND U2212 ( .A(n1209), .B(n1118), .Z(n1206) );
  AND U2213 ( .A(n1210), .B(n1211), .Z(n1202) );
  NAND U2214 ( .A(n1212), .B(n1121), .Z(n1199) );
  NAND U2215 ( .A(n1213), .B(n1214), .Z(n1212) );
  AND U2216 ( .A(n1215), .B(n1211), .Z(n1214) );
  NAND U2217 ( .A(n1132), .B(n1216), .Z(n1211) );
  AND U2218 ( .A(n1210), .B(n1217), .Z(n1215) );
  NAND U2219 ( .A(n1209), .B(n1129), .Z(n1217) );
  NAND U2220 ( .A(n1218), .B(n1134), .Z(n1210) );
  AND U2221 ( .A(n1205), .B(n1219), .Z(n1213) );
  NANDN U2222 ( .B(n1220), .A(n1221), .Z(n1219) );
  ANDN U2223 ( .A(a_bus[4]), .B(a_bus[3]), .Z(n1221) );
  NAND U2224 ( .A(n1124), .B(n1222), .Z(n1205) );
  AND U2225 ( .A(n1223), .B(n1224), .Z(n1197) );
  NAND U2226 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][11] ), .Z(n1224) );
  NAND U2227 ( .A(n1225), .B(n1140), .Z(n1223) );
  XNOR U2228 ( .A(n1226), .B(n1227), .Z(n1225) );
  AND U2229 ( .A(n1228), .B(n1229), .Z(n1195) );
  MUX U2230 ( .IN0(n1145), .IN1(n1146), .SEL(n1230), .F(n1229) );
  ANDN U2231 ( .A(n1227), .B(b_bus[11]), .Z(n1230) );
  AND U2232 ( .A(n1231), .B(n1232), .Z(n1228) );
  NAND U2233 ( .A(n1233), .B(n1151), .Z(n1232) );
  XNOR U2234 ( .A(n1227), .B(b_bus[11]), .Z(n1233) );
  IV U2235 ( .A(n1234), .Z(b_bus[11]) );
  NANDN U2236 ( .B(n1227), .A(n1235), .Z(n1231) );
  ANDN U2237 ( .A(n1154), .B(n1234), .Z(n1235) );
  AND U2238 ( .A(n1236), .B(n1237), .Z(n450) );
  AND U2239 ( .A(n1238), .B(n1239), .Z(n1237) );
  AND U2240 ( .A(n1240), .B(n1241), .Z(n1239) );
  NAND U2241 ( .A(n1242), .B(n1109), .Z(n1241) );
  NAND U2242 ( .A(n1243), .B(n1244), .Z(n1242) );
  AND U2243 ( .A(n1245), .B(n1246), .Z(n1244) );
  AND U2244 ( .A(n1247), .B(n1248), .Z(n1245) );
  OR U2245 ( .A(n1249), .B(n1117), .Z(n1248) );
  NAND U2246 ( .A(n1250), .B(n1118), .Z(n1247) );
  NAND U2247 ( .A(n1251), .B(n1121), .Z(n1240) );
  NAND U2248 ( .A(n1243), .B(n1252), .Z(n1251) );
  AND U2249 ( .A(n1253), .B(n1246), .Z(n1252) );
  NAND U2250 ( .A(n1124), .B(n1254), .Z(n1246) );
  AND U2251 ( .A(n1255), .B(n1256), .Z(n1253) );
  OR U2252 ( .A(n1257), .B(n1117), .Z(n1256) );
  NAND U2253 ( .A(n1250), .B(n1129), .Z(n1255) );
  AND U2254 ( .A(n1258), .B(n1259), .Z(n1243) );
  NAND U2255 ( .A(n1132), .B(n1260), .Z(n1259) );
  NAND U2256 ( .A(n1261), .B(n1134), .Z(n1258) );
  AND U2257 ( .A(n1262), .B(n1263), .Z(n1238) );
  NAND U2258 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][10] ), .Z(n1263) );
  NAND U2259 ( .A(n1264), .B(n1140), .Z(n1262) );
  XNOR U2260 ( .A(n1265), .B(n1266), .Z(n1264) );
  AND U2261 ( .A(n1267), .B(n1268), .Z(n1236) );
  MUX U2262 ( .IN0(n1145), .IN1(n1146), .SEL(n1269), .F(n1268) );
  ANDN U2263 ( .A(n1266), .B(b_bus[10]), .Z(n1269) );
  AND U2264 ( .A(n1270), .B(n1271), .Z(n1267) );
  NAND U2265 ( .A(n1272), .B(n1151), .Z(n1271) );
  XNOR U2266 ( .A(n1266), .B(b_bus[10]), .Z(n1272) );
  IV U2267 ( .A(n1273), .Z(b_bus[10]) );
  NANDN U2268 ( .B(n1266), .A(n1274), .Z(n1270) );
  ANDN U2269 ( .A(n1154), .B(n1273), .Z(n1274) );
  AND U2270 ( .A(n1275), .B(n1276), .Z(n1098) );
  ANDN U2271 ( .A(n428), .B(n1277), .Z(n1276) );
  IV U2272 ( .A(n417), .Z(n1277) );
  AND U2273 ( .A(n1278), .B(n1279), .Z(n417) );
  AND U2274 ( .A(n1280), .B(n1281), .Z(n1279) );
  AND U2275 ( .A(n1282), .B(n1283), .Z(n1281) );
  NAND U2276 ( .A(n1284), .B(n1109), .Z(n1283) );
  NAND U2277 ( .A(n1285), .B(n1286), .Z(n1284) );
  AND U2278 ( .A(n1287), .B(n1288), .Z(n1286) );
  AND U2279 ( .A(n1289), .B(n1290), .Z(n1287) );
  OR U2280 ( .A(n1291), .B(n1117), .Z(n1290) );
  NAND U2281 ( .A(n1135), .B(n1118), .Z(n1289) );
  AND U2282 ( .A(n1292), .B(n1293), .Z(n1285) );
  NAND U2283 ( .A(n1294), .B(n1121), .Z(n1282) );
  NAND U2284 ( .A(n1295), .B(n1296), .Z(n1294) );
  AND U2285 ( .A(n1297), .B(n1293), .Z(n1296) );
  NAND U2286 ( .A(n1132), .B(n1125), .Z(n1293) );
  AND U2287 ( .A(n1292), .B(n1298), .Z(n1297) );
  NAND U2288 ( .A(n1135), .B(n1129), .Z(n1298) );
  NAND U2289 ( .A(n1133), .B(n1134), .Z(n1292) );
  AND U2290 ( .A(n1288), .B(n1299), .Z(n1295) );
  NAND U2291 ( .A(n1300), .B(n1301), .Z(n1299) );
  NAND U2292 ( .A(n1124), .B(n1302), .Z(n1288) );
  AND U2293 ( .A(n1303), .B(n1304), .Z(n1280) );
  NAND U2294 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][13] ), .Z(n1304) );
  NAND U2295 ( .A(n1305), .B(n1140), .Z(n1303) );
  XNOR U2296 ( .A(n1306), .B(n1307), .Z(n1305) );
  AND U2297 ( .A(n1308), .B(n1309), .Z(n1278) );
  MUX U2298 ( .IN0(n1145), .IN1(n1146), .SEL(n1310), .F(n1309) );
  ANDN U2299 ( .A(n1307), .B(b_bus[13]), .Z(n1310) );
  AND U2300 ( .A(n1311), .B(n1312), .Z(n1308) );
  NAND U2301 ( .A(n1313), .B(n1151), .Z(n1312) );
  XNOR U2302 ( .A(n1307), .B(b_bus[13]), .Z(n1313) );
  IV U2303 ( .A(n1314), .Z(b_bus[13]) );
  NANDN U2304 ( .B(n1307), .A(n1315), .Z(n1311) );
  ANDN U2305 ( .A(n1154), .B(n1314), .Z(n1315) );
  AND U2306 ( .A(n1316), .B(n1317), .Z(n428) );
  AND U2307 ( .A(n1318), .B(n1319), .Z(n1317) );
  AND U2308 ( .A(n1320), .B(n1321), .Z(n1319) );
  NAND U2309 ( .A(n1322), .B(n1109), .Z(n1321) );
  NAND U2310 ( .A(n1323), .B(n1324), .Z(n1322) );
  AND U2311 ( .A(n1325), .B(n1326), .Z(n1324) );
  AND U2312 ( .A(n1327), .B(n1328), .Z(n1325) );
  OR U2313 ( .A(n1329), .B(n1117), .Z(n1328) );
  NAND U2314 ( .A(n1180), .B(n1118), .Z(n1327) );
  AND U2315 ( .A(n1330), .B(n1331), .Z(n1323) );
  NAND U2316 ( .A(n1332), .B(n1121), .Z(n1320) );
  NAND U2317 ( .A(n1333), .B(n1334), .Z(n1332) );
  AND U2318 ( .A(n1335), .B(n1331), .Z(n1334) );
  NAND U2319 ( .A(n1173), .B(n1132), .Z(n1331) );
  AND U2320 ( .A(n1330), .B(n1336), .Z(n1335) );
  NAND U2321 ( .A(n1180), .B(n1129), .Z(n1336) );
  NAND U2322 ( .A(n1179), .B(n1134), .Z(n1330) );
  AND U2323 ( .A(n1326), .B(n1337), .Z(n1333) );
  NAND U2324 ( .A(n1338), .B(n1300), .Z(n1337) );
  NAND U2325 ( .A(n1124), .B(n1339), .Z(n1326) );
  AND U2326 ( .A(n1340), .B(n1341), .Z(n1318) );
  NAND U2327 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][12] ), .Z(n1341) );
  NAND U2328 ( .A(n1342), .B(n1140), .Z(n1340) );
  XNOR U2329 ( .A(n1343), .B(n1344), .Z(n1342) );
  AND U2330 ( .A(n1345), .B(n1346), .Z(n1316) );
  MUX U2331 ( .IN0(n1145), .IN1(n1146), .SEL(n1347), .F(n1346) );
  ANDN U2332 ( .A(n1344), .B(b_bus[12]), .Z(n1347) );
  AND U2333 ( .A(n1348), .B(n1349), .Z(n1345) );
  NAND U2334 ( .A(n1350), .B(n1151), .Z(n1349) );
  XNOR U2335 ( .A(n1344), .B(b_bus[12]), .Z(n1350) );
  IV U2336 ( .A(n1351), .Z(b_bus[12]) );
  NANDN U2337 ( .B(n1344), .A(n1352), .Z(n1348) );
  ANDN U2338 ( .A(n1154), .B(n1351), .Z(n1352) );
  ANDN U2339 ( .A(n405), .B(n1353), .Z(n1275) );
  IV U2340 ( .A(n391), .Z(n1353) );
  AND U2341 ( .A(n1354), .B(n1355), .Z(n391) );
  AND U2342 ( .A(n1356), .B(n1357), .Z(n1355) );
  AND U2343 ( .A(n1358), .B(n1359), .Z(n1357) );
  NAND U2344 ( .A(n1360), .B(n1109), .Z(n1359) );
  NAND U2345 ( .A(n1361), .B(n1362), .Z(n1360) );
  AND U2346 ( .A(n1363), .B(n1364), .Z(n1362) );
  AND U2347 ( .A(n1365), .B(n1366), .Z(n1363) );
  NAND U2348 ( .A(n1218), .B(n1118), .Z(n1366) );
  AND U2349 ( .A(n1367), .B(n1368), .Z(n1361) );
  NAND U2350 ( .A(n1124), .B(n1369), .Z(n1367) );
  NAND U2351 ( .A(n1370), .B(n1121), .Z(n1358) );
  NAND U2352 ( .A(n1371), .B(n1372), .Z(n1370) );
  AND U2353 ( .A(n1373), .B(n1368), .Z(n1372) );
  NAND U2354 ( .A(n1132), .B(n1222), .Z(n1368) );
  AND U2355 ( .A(n1364), .B(n1374), .Z(n1373) );
  NAND U2356 ( .A(n1218), .B(n1129), .Z(n1374) );
  NAND U2357 ( .A(n1216), .B(n1134), .Z(n1364) );
  AND U2358 ( .A(n1375), .B(n1376), .Z(n1371) );
  NANDN U2359 ( .B(n1377), .A(n1300), .Z(n1376) );
  NANDN U2360 ( .B(n1378), .A(n1124), .Z(n1375) );
  AND U2361 ( .A(n1379), .B(n1380), .Z(n1356) );
  NAND U2362 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][15] ), .Z(n1380) );
  NAND U2363 ( .A(n1381), .B(n1140), .Z(n1379) );
  XNOR U2364 ( .A(n1382), .B(n1383), .Z(n1381) );
  AND U2365 ( .A(n1384), .B(n1385), .Z(n1354) );
  MUX U2366 ( .IN0(n1145), .IN1(n1146), .SEL(n1386), .F(n1385) );
  ANDN U2367 ( .A(n1383), .B(b_bus[15]), .Z(n1386) );
  AND U2368 ( .A(n1387), .B(n1388), .Z(n1384) );
  NAND U2369 ( .A(n1389), .B(n1151), .Z(n1388) );
  XNOR U2370 ( .A(n1383), .B(b_bus[15]), .Z(n1389) );
  IV U2371 ( .A(n1390), .Z(b_bus[15]) );
  NANDN U2372 ( .B(n1383), .A(n1391), .Z(n1387) );
  ANDN U2373 ( .A(n1154), .B(n1390), .Z(n1391) );
  AND U2374 ( .A(n1392), .B(n1393), .Z(n405) );
  AND U2375 ( .A(n1394), .B(n1395), .Z(n1393) );
  AND U2376 ( .A(n1396), .B(n1397), .Z(n1395) );
  NAND U2377 ( .A(n1398), .B(n1109), .Z(n1397) );
  NAND U2378 ( .A(n1399), .B(n1400), .Z(n1398) );
  AND U2379 ( .A(n1401), .B(n1402), .Z(n1400) );
  AND U2380 ( .A(n1403), .B(n1404), .Z(n1401) );
  OR U2381 ( .A(n1405), .B(n1117), .Z(n1404) );
  NAND U2382 ( .A(n1261), .B(n1118), .Z(n1403) );
  AND U2383 ( .A(n1406), .B(n1407), .Z(n1399) );
  NAND U2384 ( .A(n1408), .B(n1121), .Z(n1396) );
  NAND U2385 ( .A(n1409), .B(n1410), .Z(n1408) );
  AND U2386 ( .A(n1411), .B(n1407), .Z(n1410) );
  NAND U2387 ( .A(n1132), .B(n1254), .Z(n1407) );
  AND U2388 ( .A(n1406), .B(n1412), .Z(n1411) );
  NAND U2389 ( .A(n1261), .B(n1129), .Z(n1412) );
  NAND U2390 ( .A(n1260), .B(n1134), .Z(n1406) );
  AND U2391 ( .A(n1402), .B(n1413), .Z(n1409) );
  NAND U2392 ( .A(n1300), .B(n1414), .Z(n1413) );
  AND U2393 ( .A(n1415), .B(a_bus[4]), .Z(n1300) );
  NAND U2394 ( .A(n1124), .B(n1416), .Z(n1402) );
  AND U2395 ( .A(n1417), .B(n1418), .Z(n1394) );
  NAND U2396 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][14] ), .Z(n1418) );
  NAND U2397 ( .A(n1419), .B(n1140), .Z(n1417) );
  XNOR U2398 ( .A(n1420), .B(n1421), .Z(n1419) );
  AND U2399 ( .A(n1422), .B(n1423), .Z(n1392) );
  MUX U2400 ( .IN0(n1145), .IN1(n1146), .SEL(n1424), .F(n1423) );
  ANDN U2401 ( .A(n1421), .B(b_bus[14]), .Z(n1424) );
  AND U2402 ( .A(n1425), .B(n1426), .Z(n1422) );
  NAND U2403 ( .A(n1427), .B(n1151), .Z(n1426) );
  XNOR U2404 ( .A(n1421), .B(b_bus[14]), .Z(n1427) );
  IV U2405 ( .A(n1428), .Z(b_bus[14]) );
  NANDN U2406 ( .B(n1421), .A(n1429), .Z(n1425) );
  ANDN U2407 ( .A(n1154), .B(n1428), .Z(n1429) );
  AND U2408 ( .A(n1430), .B(n1431), .Z(n1088) );
  AND U2409 ( .A(n1432), .B(n1433), .Z(n1431) );
  AND U2410 ( .A(n1434), .B(n1435), .Z(n1433) );
  ANDN U2411 ( .A(n374), .B(n1436), .Z(n1435) );
  IV U2412 ( .A(n366), .Z(n1436) );
  AND U2413 ( .A(n1437), .B(n1438), .Z(n366) );
  AND U2414 ( .A(n1439), .B(n1440), .Z(n1438) );
  AND U2415 ( .A(n1441), .B(n1442), .Z(n1440) );
  NAND U2416 ( .A(n1443), .B(n1109), .Z(n1442) );
  NAND U2417 ( .A(n1444), .B(n1365), .Z(n1443) );
  OR U2418 ( .A(n1445), .B(a_bus[4]), .Z(n1444) );
  NAND U2419 ( .A(n1446), .B(n1121), .Z(n1441) );
  NOR U2420 ( .A(a_bus[4]), .B(n1447), .Z(n1446) );
  AND U2421 ( .A(n1448), .B(n1449), .Z(n1439) );
  NANDN U2422 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][17] ), .Z(n1449) );
  NAND U2423 ( .A(n1451), .B(n1140), .Z(n1448) );
  XNOR U2424 ( .A(n1452), .B(n1453), .Z(n1451) );
  AND U2425 ( .A(n1454), .B(n1455), .Z(n1437) );
  MUX U2426 ( .IN0(n1145), .IN1(n1146), .SEL(n1456), .F(n1455) );
  ANDN U2427 ( .A(n1453), .B(b_bus[17]), .Z(n1456) );
  AND U2428 ( .A(n1457), .B(n1458), .Z(n1454) );
  NAND U2429 ( .A(n1459), .B(n1151), .Z(n1458) );
  XNOR U2430 ( .A(n1453), .B(b_bus[17]), .Z(n1459) );
  IV U2431 ( .A(n1460), .Z(b_bus[17]) );
  NANDN U2432 ( .B(n1453), .A(n1461), .Z(n1457) );
  ANDN U2433 ( .A(n1154), .B(n1460), .Z(n1461) );
  AND U2434 ( .A(n1462), .B(n1463), .Z(n374) );
  AND U2435 ( .A(n1464), .B(n1465), .Z(n1463) );
  AND U2436 ( .A(n1466), .B(n1467), .Z(n1465) );
  NAND U2437 ( .A(n1468), .B(n1109), .Z(n1467) );
  NAND U2438 ( .A(n1469), .B(n1365), .Z(n1468) );
  OR U2439 ( .A(n1470), .B(a_bus[4]), .Z(n1469) );
  NAND U2440 ( .A(n1471), .B(n1121), .Z(n1466) );
  NOR U2441 ( .A(a_bus[4]), .B(n1472), .Z(n1471) );
  AND U2442 ( .A(n1473), .B(n1474), .Z(n1464) );
  NANDN U2443 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][16] ), .Z(n1474) );
  NAND U2444 ( .A(n1475), .B(n1140), .Z(n1473) );
  XNOR U2445 ( .A(n1476), .B(n1477), .Z(n1475) );
  AND U2446 ( .A(n1478), .B(n1479), .Z(n1462) );
  MUX U2447 ( .IN0(n1145), .IN1(n1146), .SEL(n1480), .F(n1479) );
  ANDN U2448 ( .A(n1477), .B(b_bus[16]), .Z(n1480) );
  AND U2449 ( .A(n1481), .B(n1482), .Z(n1478) );
  NAND U2450 ( .A(n1483), .B(n1151), .Z(n1482) );
  XNOR U2451 ( .A(n1477), .B(b_bus[16]), .Z(n1483) );
  IV U2452 ( .A(n1484), .Z(b_bus[16]) );
  NANDN U2453 ( .B(n1477), .A(n1485), .Z(n1481) );
  ANDN U2454 ( .A(n1154), .B(n1484), .Z(n1485) );
  ANDN U2455 ( .A(n357), .B(n1486), .Z(n1434) );
  IV U2456 ( .A(n348), .Z(n1486) );
  AND U2457 ( .A(n1487), .B(n1488), .Z(n348) );
  AND U2458 ( .A(n1489), .B(n1490), .Z(n1488) );
  AND U2459 ( .A(n1491), .B(n1492), .Z(n1490) );
  NAND U2460 ( .A(n1493), .B(n1109), .Z(n1492) );
  NAND U2461 ( .A(n1494), .B(n1365), .Z(n1493) );
  OR U2462 ( .A(n1495), .B(a_bus[4]), .Z(n1494) );
  NAND U2463 ( .A(n1496), .B(n1121), .Z(n1491) );
  NOR U2464 ( .A(a_bus[4]), .B(n1497), .Z(n1496) );
  AND U2465 ( .A(n1498), .B(n1499), .Z(n1489) );
  NANDN U2466 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][19] ), .Z(n1499) );
  NAND U2467 ( .A(n1500), .B(n1140), .Z(n1498) );
  XNOR U2468 ( .A(n1501), .B(n1502), .Z(n1500) );
  AND U2469 ( .A(n1503), .B(n1504), .Z(n1487) );
  MUX U2470 ( .IN0(n1145), .IN1(n1146), .SEL(n1505), .F(n1504) );
  ANDN U2471 ( .A(n1502), .B(b_bus[19]), .Z(n1505) );
  AND U2472 ( .A(n1506), .B(n1507), .Z(n1503) );
  NAND U2473 ( .A(n1508), .B(n1151), .Z(n1507) );
  XNOR U2474 ( .A(n1502), .B(b_bus[19]), .Z(n1508) );
  IV U2475 ( .A(n1509), .Z(b_bus[19]) );
  NANDN U2476 ( .B(n1502), .A(n1510), .Z(n1506) );
  ANDN U2477 ( .A(n1154), .B(n1509), .Z(n1510) );
  AND U2478 ( .A(n1511), .B(n1512), .Z(n357) );
  AND U2479 ( .A(n1513), .B(n1514), .Z(n1512) );
  AND U2480 ( .A(n1515), .B(n1516), .Z(n1514) );
  NAND U2481 ( .A(n1517), .B(n1109), .Z(n1516) );
  NAND U2482 ( .A(n1518), .B(n1365), .Z(n1517) );
  OR U2483 ( .A(n1519), .B(a_bus[4]), .Z(n1518) );
  NAND U2484 ( .A(n1520), .B(n1121), .Z(n1515) );
  NOR U2485 ( .A(a_bus[4]), .B(n1521), .Z(n1520) );
  AND U2486 ( .A(n1522), .B(n1523), .Z(n1513) );
  NANDN U2487 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][18] ), .Z(n1523) );
  NAND U2488 ( .A(n1524), .B(n1140), .Z(n1522) );
  XNOR U2489 ( .A(n1525), .B(n1526), .Z(n1524) );
  AND U2490 ( .A(n1527), .B(n1528), .Z(n1511) );
  MUX U2491 ( .IN0(n1145), .IN1(n1146), .SEL(n1529), .F(n1528) );
  ANDN U2492 ( .A(n1526), .B(b_bus[18]), .Z(n1529) );
  AND U2493 ( .A(n1530), .B(n1531), .Z(n1527) );
  NAND U2494 ( .A(n1532), .B(n1151), .Z(n1531) );
  XNOR U2495 ( .A(n1526), .B(b_bus[18]), .Z(n1532) );
  IV U2496 ( .A(n1533), .Z(b_bus[18]) );
  NANDN U2497 ( .B(n1526), .A(n1534), .Z(n1530) );
  ANDN U2498 ( .A(n1154), .B(n1533), .Z(n1534) );
  AND U2499 ( .A(n1535), .B(n1536), .Z(n1432) );
  ANDN U2500 ( .A(n339), .B(n1537), .Z(n1536) );
  IV U2501 ( .A(n331), .Z(n1537) );
  AND U2502 ( .A(n1538), .B(n1539), .Z(n331) );
  AND U2503 ( .A(n1540), .B(n1541), .Z(n1539) );
  AND U2504 ( .A(n1542), .B(n1543), .Z(n1541) );
  NAND U2505 ( .A(n1544), .B(n1109), .Z(n1543) );
  NAND U2506 ( .A(n1545), .B(n1365), .Z(n1544) );
  OR U2507 ( .A(n1546), .B(a_bus[4]), .Z(n1545) );
  NAND U2508 ( .A(n1547), .B(n1121), .Z(n1542) );
  NOR U2509 ( .A(a_bus[4]), .B(n1548), .Z(n1547) );
  AND U2510 ( .A(n1549), .B(n1550), .Z(n1540) );
  NANDN U2511 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][21] ), .Z(n1550) );
  NAND U2512 ( .A(n1551), .B(n1140), .Z(n1549) );
  XNOR U2513 ( .A(n1552), .B(n1553), .Z(n1551) );
  AND U2514 ( .A(n1554), .B(n1555), .Z(n1538) );
  MUX U2515 ( .IN0(n1145), .IN1(n1146), .SEL(n1556), .F(n1555) );
  ANDN U2516 ( .A(n1553), .B(b_bus[21]), .Z(n1556) );
  AND U2517 ( .A(n1557), .B(n1558), .Z(n1554) );
  NAND U2518 ( .A(n1559), .B(n1151), .Z(n1558) );
  XNOR U2519 ( .A(n1553), .B(b_bus[21]), .Z(n1559) );
  IV U2520 ( .A(n1560), .Z(b_bus[21]) );
  NANDN U2521 ( .B(n1553), .A(n1561), .Z(n1557) );
  ANDN U2522 ( .A(n1154), .B(n1560), .Z(n1561) );
  AND U2523 ( .A(n1562), .B(n1563), .Z(n339) );
  AND U2524 ( .A(n1564), .B(n1565), .Z(n1563) );
  AND U2525 ( .A(n1566), .B(n1567), .Z(n1565) );
  NAND U2526 ( .A(n1568), .B(n1109), .Z(n1567) );
  NAND U2527 ( .A(n1569), .B(n1365), .Z(n1568) );
  OR U2528 ( .A(n1570), .B(a_bus[4]), .Z(n1569) );
  NAND U2529 ( .A(n1571), .B(n1121), .Z(n1566) );
  NOR U2530 ( .A(a_bus[4]), .B(n1572), .Z(n1571) );
  AND U2531 ( .A(n1573), .B(n1574), .Z(n1564) );
  NANDN U2532 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][20] ), .Z(n1574) );
  NAND U2533 ( .A(n1575), .B(n1140), .Z(n1573) );
  XNOR U2534 ( .A(n1576), .B(n1577), .Z(n1575) );
  AND U2535 ( .A(n1578), .B(n1579), .Z(n1562) );
  MUX U2536 ( .IN0(n1145), .IN1(n1146), .SEL(n1580), .F(n1579) );
  ANDN U2537 ( .A(n1577), .B(b_bus[20]), .Z(n1580) );
  AND U2538 ( .A(n1581), .B(n1582), .Z(n1578) );
  NAND U2539 ( .A(n1583), .B(n1151), .Z(n1582) );
  XNOR U2540 ( .A(n1577), .B(b_bus[20]), .Z(n1583) );
  IV U2541 ( .A(n1584), .Z(b_bus[20]) );
  NANDN U2542 ( .B(n1577), .A(n1585), .Z(n1581) );
  ANDN U2543 ( .A(n1154), .B(n1584), .Z(n1585) );
  ANDN U2544 ( .A(n323), .B(n1586), .Z(n1535) );
  IV U2545 ( .A(n315), .Z(n1586) );
  AND U2546 ( .A(n1587), .B(n1588), .Z(n315) );
  AND U2547 ( .A(n1589), .B(n1590), .Z(n1588) );
  AND U2548 ( .A(n1591), .B(n1592), .Z(n1590) );
  NAND U2549 ( .A(n1593), .B(n1109), .Z(n1592) );
  NAND U2550 ( .A(n1594), .B(n1365), .Z(n1593) );
  OR U2551 ( .A(n1595), .B(a_bus[4]), .Z(n1594) );
  NAND U2552 ( .A(n1596), .B(n1121), .Z(n1591) );
  NOR U2553 ( .A(a_bus[4]), .B(n1597), .Z(n1596) );
  AND U2554 ( .A(n1598), .B(n1599), .Z(n1589) );
  NANDN U2555 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][23] ), .Z(n1599) );
  NAND U2556 ( .A(n1600), .B(n1140), .Z(n1598) );
  XNOR U2557 ( .A(n1601), .B(n1602), .Z(n1600) );
  AND U2558 ( .A(n1603), .B(n1604), .Z(n1587) );
  MUX U2559 ( .IN0(n1145), .IN1(n1146), .SEL(n1605), .F(n1604) );
  ANDN U2560 ( .A(n1602), .B(b_bus[23]), .Z(n1605) );
  AND U2561 ( .A(n1606), .B(n1607), .Z(n1603) );
  NAND U2562 ( .A(n1608), .B(n1151), .Z(n1607) );
  XNOR U2563 ( .A(n1602), .B(b_bus[23]), .Z(n1608) );
  IV U2564 ( .A(n1609), .Z(b_bus[23]) );
  NANDN U2565 ( .B(n1602), .A(n1610), .Z(n1606) );
  ANDN U2566 ( .A(n1154), .B(n1609), .Z(n1610) );
  AND U2567 ( .A(n1611), .B(n1612), .Z(n323) );
  AND U2568 ( .A(n1613), .B(n1614), .Z(n1612) );
  AND U2569 ( .A(n1615), .B(n1616), .Z(n1614) );
  NAND U2570 ( .A(n1617), .B(n1109), .Z(n1616) );
  NAND U2571 ( .A(n1618), .B(n1365), .Z(n1617) );
  OR U2572 ( .A(n1619), .B(a_bus[4]), .Z(n1618) );
  NAND U2573 ( .A(n1620), .B(n1121), .Z(n1615) );
  NOR U2574 ( .A(a_bus[4]), .B(n1621), .Z(n1620) );
  AND U2575 ( .A(n1622), .B(n1623), .Z(n1613) );
  NANDN U2576 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][22] ), .Z(n1623) );
  NAND U2577 ( .A(n1624), .B(n1140), .Z(n1622) );
  XNOR U2578 ( .A(n1625), .B(n1626), .Z(n1624) );
  AND U2579 ( .A(n1627), .B(n1628), .Z(n1611) );
  MUX U2580 ( .IN0(n1145), .IN1(n1146), .SEL(n1629), .F(n1628) );
  ANDN U2581 ( .A(n1626), .B(b_bus[22]), .Z(n1629) );
  AND U2582 ( .A(n1630), .B(n1631), .Z(n1627) );
  NAND U2583 ( .A(n1632), .B(n1151), .Z(n1631) );
  XNOR U2584 ( .A(n1626), .B(b_bus[22]), .Z(n1632) );
  IV U2585 ( .A(n1633), .Z(b_bus[22]) );
  NANDN U2586 ( .B(n1626), .A(n1634), .Z(n1630) );
  ANDN U2587 ( .A(n1154), .B(n1633), .Z(n1634) );
  AND U2588 ( .A(n1635), .B(n1636), .Z(n1430) );
  AND U2589 ( .A(n1637), .B(n1638), .Z(n1636) );
  ANDN U2590 ( .A(n307), .B(n1639), .Z(n1638) );
  IV U2591 ( .A(n299), .Z(n1639) );
  AND U2592 ( .A(n1640), .B(n1641), .Z(n299) );
  AND U2593 ( .A(n1642), .B(n1643), .Z(n1641) );
  AND U2594 ( .A(n1644), .B(n1645), .Z(n1643) );
  NAND U2595 ( .A(n1646), .B(n1109), .Z(n1645) );
  NAND U2596 ( .A(n1647), .B(n1365), .Z(n1646) );
  OR U2597 ( .A(n1116), .B(a_bus[4]), .Z(n1647) );
  AND U2598 ( .A(n1648), .B(n1649), .Z(n1116) );
  NAND U2599 ( .A(n1302), .B(n1650), .Z(n1649) );
  ANDN U2600 ( .A(n1651), .B(n1652), .Z(n1648) );
  NAND U2601 ( .A(n1653), .B(n1654), .Z(n1651) );
  NAND U2602 ( .A(n1655), .B(n1121), .Z(n1644) );
  NOR U2603 ( .A(a_bus[4]), .B(n1128), .Z(n1655) );
  AND U2604 ( .A(n1656), .B(n1657), .Z(n1128) );
  NAND U2605 ( .A(n1415), .B(n1302), .Z(n1657) );
  NAND U2606 ( .A(n1301), .B(n1653), .Z(n1656) );
  AND U2607 ( .A(n1658), .B(n1659), .Z(n1642) );
  NANDN U2608 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][25] ), .Z(n1659) );
  NAND U2609 ( .A(n1660), .B(n1140), .Z(n1658) );
  XNOR U2610 ( .A(n1661), .B(n1662), .Z(n1660) );
  AND U2611 ( .A(n1663), .B(n1664), .Z(n1640) );
  MUX U2612 ( .IN0(n1145), .IN1(n1146), .SEL(n1665), .F(n1664) );
  ANDN U2613 ( .A(n1662), .B(b_bus[25]), .Z(n1665) );
  AND U2614 ( .A(n1666), .B(n1667), .Z(n1663) );
  NAND U2615 ( .A(n1668), .B(n1151), .Z(n1667) );
  XNOR U2616 ( .A(n1662), .B(b_bus[25]), .Z(n1668) );
  IV U2617 ( .A(n1669), .Z(b_bus[25]) );
  NANDN U2618 ( .B(n1662), .A(n1670), .Z(n1666) );
  ANDN U2619 ( .A(n1154), .B(n1669), .Z(n1670) );
  AND U2620 ( .A(n1671), .B(n1672), .Z(n307) );
  AND U2621 ( .A(n1673), .B(n1674), .Z(n1672) );
  AND U2622 ( .A(n1675), .B(n1676), .Z(n1674) );
  NAND U2623 ( .A(n1677), .B(n1109), .Z(n1676) );
  NAND U2624 ( .A(n1678), .B(n1365), .Z(n1677) );
  OR U2625 ( .A(n1168), .B(a_bus[4]), .Z(n1678) );
  AND U2626 ( .A(n1679), .B(n1680), .Z(n1168) );
  NAND U2627 ( .A(n1339), .B(n1650), .Z(n1680) );
  ANDN U2628 ( .A(n1681), .B(n1652), .Z(n1679) );
  NAND U2629 ( .A(n1682), .B(n1121), .Z(n1675) );
  NOR U2630 ( .A(a_bus[4]), .B(n1176), .Z(n1682) );
  AND U2631 ( .A(n1681), .B(n1683), .Z(n1176) );
  NAND U2632 ( .A(n1415), .B(n1339), .Z(n1683) );
  NAND U2633 ( .A(n1338), .B(n1653), .Z(n1681) );
  AND U2634 ( .A(n1684), .B(n1685), .Z(n1673) );
  NANDN U2635 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][24] ), .Z(n1685) );
  NAND U2636 ( .A(n1686), .B(n1140), .Z(n1684) );
  XNOR U2637 ( .A(n1687), .B(n1688), .Z(n1686) );
  AND U2638 ( .A(n1689), .B(n1690), .Z(n1671) );
  MUX U2639 ( .IN0(n1145), .IN1(n1146), .SEL(n1691), .F(n1690) );
  ANDN U2640 ( .A(n1688), .B(b_bus[24]), .Z(n1691) );
  AND U2641 ( .A(n1692), .B(n1693), .Z(n1689) );
  NAND U2642 ( .A(n1694), .B(n1151), .Z(n1693) );
  XNOR U2643 ( .A(n1688), .B(b_bus[24]), .Z(n1694) );
  IV U2644 ( .A(n1695), .Z(b_bus[24]) );
  NANDN U2645 ( .B(n1688), .A(n1696), .Z(n1692) );
  ANDN U2646 ( .A(n1154), .B(n1695), .Z(n1696) );
  ANDN U2647 ( .A(n291), .B(n1697), .Z(n1637) );
  IV U2648 ( .A(n283), .Z(n1697) );
  AND U2649 ( .A(n1698), .B(n1699), .Z(n283) );
  AND U2650 ( .A(n1700), .B(n1701), .Z(n1699) );
  AND U2651 ( .A(n1702), .B(n1703), .Z(n1701) );
  NAND U2652 ( .A(n1704), .B(n1109), .Z(n1703) );
  NAND U2653 ( .A(n1705), .B(n1365), .Z(n1704) );
  NANDN U2654 ( .B(a_bus[4]), .A(n1208), .Z(n1705) );
  NAND U2655 ( .A(n1706), .B(n1707), .Z(n1208) );
  NAND U2656 ( .A(n1369), .B(n1650), .Z(n1706) );
  NAND U2657 ( .A(n1708), .B(n1709), .Z(n1702) );
  ANDN U2658 ( .A(n1117), .B(a_bus[3]), .Z(n1709) );
  ANDN U2659 ( .A(n1121), .B(n1220), .Z(n1708) );
  AND U2660 ( .A(n1710), .B(n1711), .Z(n1700) );
  NANDN U2661 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][27] ), .Z(n1711) );
  NAND U2662 ( .A(n1712), .B(n1140), .Z(n1710) );
  XNOR U2663 ( .A(n1713), .B(n1714), .Z(n1712) );
  AND U2664 ( .A(n1715), .B(n1716), .Z(n1698) );
  MUX U2665 ( .IN0(n1145), .IN1(n1146), .SEL(n1717), .F(n1716) );
  ANDN U2666 ( .A(n1714), .B(b_bus[27]), .Z(n1717) );
  AND U2667 ( .A(n1718), .B(n1719), .Z(n1715) );
  NAND U2668 ( .A(n1720), .B(n1151), .Z(n1719) );
  XNOR U2669 ( .A(n1714), .B(b_bus[27]), .Z(n1720) );
  IV U2670 ( .A(n1721), .Z(b_bus[27]) );
  NANDN U2671 ( .B(n1714), .A(n1722), .Z(n1718) );
  ANDN U2672 ( .A(n1154), .B(n1721), .Z(n1722) );
  AND U2673 ( .A(n1723), .B(n1724), .Z(n291) );
  AND U2674 ( .A(n1725), .B(n1726), .Z(n1724) );
  AND U2675 ( .A(n1727), .B(n1728), .Z(n1726) );
  NAND U2676 ( .A(n1729), .B(n1109), .Z(n1728) );
  NAND U2677 ( .A(n1730), .B(n1365), .Z(n1729) );
  OR U2678 ( .A(n1249), .B(a_bus[4]), .Z(n1730) );
  AND U2679 ( .A(n1731), .B(n1732), .Z(n1249) );
  NAND U2680 ( .A(n1416), .B(n1650), .Z(n1732) );
  ANDN U2681 ( .A(n1733), .B(n1652), .Z(n1731) );
  NAND U2682 ( .A(n1734), .B(n1653), .Z(n1733) );
  NAND U2683 ( .A(n1735), .B(n1121), .Z(n1727) );
  NOR U2684 ( .A(a_bus[4]), .B(n1257), .Z(n1735) );
  AND U2685 ( .A(n1736), .B(n1737), .Z(n1257) );
  NAND U2686 ( .A(n1415), .B(n1416), .Z(n1737) );
  NAND U2687 ( .A(n1414), .B(n1653), .Z(n1736) );
  AND U2688 ( .A(n1738), .B(n1739), .Z(n1725) );
  NANDN U2689 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][26] ), .Z(n1739) );
  NAND U2690 ( .A(n1740), .B(n1140), .Z(n1738) );
  XNOR U2691 ( .A(n1741), .B(n1742), .Z(n1740) );
  AND U2692 ( .A(n1743), .B(n1744), .Z(n1723) );
  MUX U2693 ( .IN0(n1145), .IN1(n1146), .SEL(n1745), .F(n1744) );
  ANDN U2694 ( .A(n1742), .B(b_bus[26]), .Z(n1745) );
  AND U2695 ( .A(n1746), .B(n1747), .Z(n1743) );
  NAND U2696 ( .A(n1748), .B(n1151), .Z(n1747) );
  XNOR U2697 ( .A(n1742), .B(b_bus[26]), .Z(n1748) );
  IV U2698 ( .A(n1749), .Z(b_bus[26]) );
  NANDN U2699 ( .B(n1742), .A(n1750), .Z(n1746) );
  ANDN U2700 ( .A(n1154), .B(n1749), .Z(n1750) );
  AND U2701 ( .A(n1751), .B(n1752), .Z(n1635) );
  ANDN U2702 ( .A(n275), .B(n1753), .Z(n1752) );
  IV U2703 ( .A(n267), .Z(n1753) );
  AND U2704 ( .A(n1754), .B(n1755), .Z(n267) );
  AND U2705 ( .A(n1756), .B(n1757), .Z(n1755) );
  AND U2706 ( .A(n1758), .B(n1759), .Z(n1757) );
  NAND U2707 ( .A(n1760), .B(n1109), .Z(n1759) );
  NAND U2708 ( .A(n1761), .B(n1365), .Z(n1760) );
  OR U2709 ( .A(n1291), .B(a_bus[4]), .Z(n1761) );
  AND U2710 ( .A(n1762), .B(n1707), .Z(n1291) );
  NAND U2711 ( .A(n1654), .B(n1650), .Z(n1762) );
  NAND U2712 ( .A(n1763), .B(n1121), .Z(n1758) );
  AND U2713 ( .A(n1301), .B(n1129), .Z(n1763) );
  AND U2714 ( .A(n1764), .B(n1765), .Z(n1756) );
  NANDN U2715 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][29] ), .Z(n1765) );
  NAND U2716 ( .A(n1766), .B(n1140), .Z(n1764) );
  XNOR U2717 ( .A(n1767), .B(n1768), .Z(n1766) );
  AND U2718 ( .A(n1769), .B(n1770), .Z(n1754) );
  MUX U2719 ( .IN0(n1145), .IN1(n1146), .SEL(n1771), .F(n1770) );
  ANDN U2720 ( .A(n1768), .B(b_bus[29]), .Z(n1771) );
  AND U2721 ( .A(n1772), .B(n1773), .Z(n1769) );
  NAND U2722 ( .A(n1774), .B(n1151), .Z(n1773) );
  XNOR U2723 ( .A(n1768), .B(b_bus[29]), .Z(n1774) );
  IV U2724 ( .A(n1775), .Z(b_bus[29]) );
  NANDN U2725 ( .B(n1768), .A(n1776), .Z(n1772) );
  ANDN U2726 ( .A(n1154), .B(n1775), .Z(n1776) );
  AND U2727 ( .A(n1777), .B(n1778), .Z(n275) );
  AND U2728 ( .A(n1779), .B(n1780), .Z(n1778) );
  AND U2729 ( .A(n1781), .B(n1782), .Z(n1780) );
  NAND U2730 ( .A(n1783), .B(n1109), .Z(n1782) );
  NAND U2731 ( .A(n1784), .B(n1365), .Z(n1783) );
  OR U2732 ( .A(n1329), .B(a_bus[4]), .Z(n1784) );
  AND U2733 ( .A(n1707), .B(n1785), .Z(n1329) );
  NAND U2734 ( .A(n1338), .B(n1650), .Z(n1785) );
  NAND U2735 ( .A(n1786), .B(n1121), .Z(n1781) );
  AND U2736 ( .A(n1338), .B(n1129), .Z(n1786) );
  AND U2737 ( .A(n1787), .B(n1788), .Z(n1779) );
  NANDN U2738 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][28] ), .Z(n1788) );
  NAND U2739 ( .A(n1789), .B(n1140), .Z(n1787) );
  XNOR U2740 ( .A(n1790), .B(n1791), .Z(n1789) );
  AND U2741 ( .A(n1792), .B(n1793), .Z(n1777) );
  MUX U2742 ( .IN0(n1145), .IN1(n1146), .SEL(n1794), .F(n1793) );
  ANDN U2743 ( .A(n1791), .B(b_bus[28]), .Z(n1794) );
  AND U2744 ( .A(n1795), .B(n1796), .Z(n1792) );
  NAND U2745 ( .A(n1797), .B(n1151), .Z(n1796) );
  XNOR U2746 ( .A(n1791), .B(b_bus[28]), .Z(n1797) );
  IV U2747 ( .A(n1798), .Z(b_bus[28]) );
  NANDN U2748 ( .B(n1791), .A(n1799), .Z(n1795) );
  ANDN U2749 ( .A(n1154), .B(n1798), .Z(n1799) );
  ANDN U2750 ( .A(n259), .B(n1056), .Z(n1751) );
  IV U2751 ( .A(n249), .Z(n1056) );
  AND U2752 ( .A(n1800), .B(n1801), .Z(n259) );
  AND U2753 ( .A(n1802), .B(n1803), .Z(n1801) );
  AND U2754 ( .A(n1804), .B(n1805), .Z(n1803) );
  NAND U2755 ( .A(n1806), .B(n1109), .Z(n1805) );
  NAND U2756 ( .A(n1807), .B(n1365), .Z(n1806) );
  NAND U2757 ( .A(a_bus[4]), .B(\Shifter/N75 ), .Z(n1365) );
  OR U2758 ( .A(n1405), .B(a_bus[4]), .Z(n1807) );
  AND U2759 ( .A(n1808), .B(n1707), .Z(n1405) );
  ANDN U2760 ( .A(n1809), .B(n1652), .Z(n1707) );
  NANDN U2761 ( .B(n1810), .A(a_bus[2]), .Z(n1809) );
  NAND U2762 ( .A(n1734), .B(n1650), .Z(n1808) );
  NAND U2763 ( .A(n1811), .B(n1121), .Z(n1804) );
  AND U2764 ( .A(n1414), .B(n1129), .Z(n1811) );
  AND U2765 ( .A(n1812), .B(n1813), .Z(n1802) );
  NANDN U2766 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][30] ), .Z(n1813) );
  NAND U2767 ( .A(n1814), .B(n1140), .Z(n1812) );
  XNOR U2768 ( .A(n1815), .B(n1816), .Z(n1814) );
  AND U2769 ( .A(n1817), .B(n1818), .Z(n1800) );
  MUX U2770 ( .IN0(n1145), .IN1(n1146), .SEL(n1819), .F(n1818) );
  ANDN U2771 ( .A(n1816), .B(b_bus[30]), .Z(n1819) );
  AND U2772 ( .A(n1820), .B(n1821), .Z(n1817) );
  NAND U2773 ( .A(n1822), .B(n1151), .Z(n1821) );
  XNOR U2774 ( .A(n1816), .B(b_bus[30]), .Z(n1822) );
  NANDN U2775 ( .B(n1816), .A(n1823), .Z(n1820) );
  ANDN U2776 ( .A(n1154), .B(n1824), .Z(n1823) );
  XOR U2777 ( .A(pc_current[31]), .B(\PC_Next/add_32/carry[29] ), .Z(n244) );
  NANDN U2778 ( .B(n249), .A(n831), .Z(n1039) );
  ANDN U2779 ( .A(n1038), .B(n1037), .Z(n831) );
  NANDN U2780 ( .B(n6), .A(n1825), .Z(n1037) );
  NAND U2781 ( .A(n1826), .B(n1827), .Z(n1825) );
  AND U2782 ( .A(n1828), .B(n1829), .Z(n1826) );
  AND U2783 ( .A(n1830), .B(n1831), .Z(n1038) );
  NANDN U2784 ( .B(n1832), .A(n1829), .Z(n1830) );
  NAND U2785 ( .A(n143), .B(n1833), .Z(n1829) );
  AND U2786 ( .A(n1834), .B(n1835), .Z(n249) );
  AND U2787 ( .A(n1836), .B(n1837), .Z(n1835) );
  AND U2788 ( .A(n1838), .B(n1839), .Z(n1837) );
  NANDN U2789 ( .B(n1810), .A(n1109), .Z(n1839) );
  NANDN U2790 ( .B(n1377), .A(n1840), .Z(n1838) );
  AND U2791 ( .A(n1129), .B(n1121), .Z(n1840) );
  AND U2792 ( .A(n1841), .B(n1842), .Z(n1836) );
  NANDN U2793 ( .B(n1450), .A(\Shifter/sll_27/ML_int[5][31] ), .Z(n1842) );
  NAND U2794 ( .A(n1140), .B(n1843), .Z(n1841) );
  AND U2795 ( .A(n1844), .B(n1845), .Z(n1834) );
  MUX U2796 ( .IN0(n1145), .IN1(n1146), .SEL(n1846), .F(n1845) );
  ANDN U2797 ( .A(n1810), .B(n1847), .Z(n1846) );
  AND U2798 ( .A(n1848), .B(n1849), .Z(n1844) );
  NAND U2799 ( .A(n1850), .B(n1151), .Z(n1849) );
  XNOR U2800 ( .A(n1851), .B(\Shifter/N75 ), .Z(n1850) );
  NANDN U2801 ( .B(n1851), .A(n1852), .Z(n1848) );
  ANDN U2802 ( .A(n1154), .B(n1810), .Z(n1852) );
  IV U2803 ( .A(n553), .Z(N27) );
  IV U2804 ( .A(n485), .Z(N24) );
  MUX U2805 ( .IN0(n1853), .IN1(o[31]), .SEL(n1854), .F(\Data_Mem/n7760 ) );
  MUX U2806 ( .IN0(n1855), .IN1(o[30]), .SEL(n1854), .F(\Data_Mem/n7759 ) );
  MUX U2807 ( .IN0(n1856), .IN1(o[29]), .SEL(n1854), .F(\Data_Mem/n7758 ) );
  MUX U2808 ( .IN0(n1857), .IN1(o[28]), .SEL(n1854), .F(\Data_Mem/n7757 ) );
  MUX U2809 ( .IN0(n1858), .IN1(o[27]), .SEL(n1854), .F(\Data_Mem/n7756 ) );
  MUX U2810 ( .IN0(n1859), .IN1(o[26]), .SEL(n1854), .F(\Data_Mem/n7755 ) );
  MUX U2811 ( .IN0(n1860), .IN1(o[25]), .SEL(n1854), .F(\Data_Mem/n7754 ) );
  MUX U2812 ( .IN0(n1861), .IN1(o[24]), .SEL(n1854), .F(\Data_Mem/n7753 ) );
  ANDN U2813 ( .A(n1862), .B(n1863), .Z(n1854) );
  ANDN U2814 ( .A(n1864), .B(n1865), .Z(n1862) );
  OR U2815 ( .A(n1866), .B(n1867), .Z(n1864) );
  MUX U2816 ( .IN0(n1868), .IN1(o[23]), .SEL(n1869), .F(\Data_Mem/n7752 ) );
  MUX U2817 ( .IN0(n1870), .IN1(o[22]), .SEL(n1869), .F(\Data_Mem/n7751 ) );
  MUX U2818 ( .IN0(n1871), .IN1(o[21]), .SEL(n1869), .F(\Data_Mem/n7750 ) );
  MUX U2819 ( .IN0(n1872), .IN1(o[20]), .SEL(n1869), .F(\Data_Mem/n7749 ) );
  MUX U2820 ( .IN0(n1873), .IN1(o[19]), .SEL(n1869), .F(\Data_Mem/n7748 ) );
  IV U2821 ( .A(n1874), .Z(n1869) );
  MUX U2822 ( .IN0(o[18]), .IN1(n1875), .SEL(n1874), .F(\Data_Mem/n7747 ) );
  MUX U2823 ( .IN0(o[17]), .IN1(n1876), .SEL(n1874), .F(\Data_Mem/n7746 ) );
  MUX U2824 ( .IN0(o[16]), .IN1(n1877), .SEL(n1874), .F(\Data_Mem/n7745 ) );
  NAND U2825 ( .A(n1878), .B(n1879), .Z(n1874) );
  OR U2826 ( .A(n1866), .B(n1880), .Z(n1879) );
  NOR U2827 ( .A(n1863), .B(n1865), .Z(n1878) );
  ANDN U2828 ( .A(n1881), .B(n1882), .Z(n1865) );
  NOR U2829 ( .A(n399), .B(n1866), .Z(n1881) );
  MUX U2830 ( .IN0(n1883), .IN1(o[15]), .SEL(n1884), .F(\Data_Mem/n7744 ) );
  MUX U2831 ( .IN0(n1885), .IN1(o[14]), .SEL(n1884), .F(\Data_Mem/n7743 ) );
  MUX U2832 ( .IN0(n1886), .IN1(o[13]), .SEL(n1884), .F(\Data_Mem/n7742 ) );
  MUX U2833 ( .IN0(n1887), .IN1(o[12]), .SEL(n1884), .F(\Data_Mem/n7741 ) );
  MUX U2834 ( .IN0(n1888), .IN1(o[11]), .SEL(n1884), .F(\Data_Mem/n7740 ) );
  IV U2835 ( .A(n1889), .Z(n1884) );
  MUX U2836 ( .IN0(o[10]), .IN1(n1890), .SEL(n1889), .F(\Data_Mem/n7739 ) );
  MUX U2837 ( .IN0(o[9]), .IN1(n1891), .SEL(n1889), .F(\Data_Mem/n7738 ) );
  MUX U2838 ( .IN0(o[8]), .IN1(n1892), .SEL(n1889), .F(\Data_Mem/n7737 ) );
  NAND U2839 ( .A(n1893), .B(n1894), .Z(n1889) );
  OR U2840 ( .A(n1895), .B(n1866), .Z(n1894) );
  MUX U2841 ( .IN0(reg_target[7]), .IN1(o[7]), .SEL(n1896), .F(
        \Data_Mem/n7736 ) );
  MUX U2842 ( .IN0(reg_target[6]), .IN1(o[6]), .SEL(n1896), .F(
        \Data_Mem/n7735 ) );
  MUX U2843 ( .IN0(reg_target[5]), .IN1(o[5]), .SEL(n1896), .F(
        \Data_Mem/n7734 ) );
  MUX U2844 ( .IN0(reg_target[4]), .IN1(o[4]), .SEL(n1896), .F(
        \Data_Mem/n7733 ) );
  MUX U2845 ( .IN0(reg_target[3]), .IN1(o[3]), .SEL(n1896), .F(
        \Data_Mem/n7732 ) );
  IV U2846 ( .A(n1897), .Z(n1896) );
  MUX U2847 ( .IN0(o[2]), .IN1(reg_target[2]), .SEL(n1897), .F(
        \Data_Mem/n7731 ) );
  MUX U2848 ( .IN0(o[1]), .IN1(reg_target[1]), .SEL(n1897), .F(
        \Data_Mem/n7730 ) );
  MUX U2849 ( .IN0(o[0]), .IN1(reg_target[0]), .SEL(n1897), .F(
        \Data_Mem/n7729 ) );
  NAND U2850 ( .A(n1893), .B(n1898), .Z(n1897) );
  NANDN U2851 ( .B(n1866), .A(n1899), .Z(n1898) );
  NOR U2852 ( .A(n1863), .B(n1900), .Z(n1893) );
  ANDN U2853 ( .A(n1901), .B(n1882), .Z(n1900) );
  NOR U2854 ( .A(n411), .B(n1866), .Z(n1901) );
  ANDN U2855 ( .A(n1902), .B(n1866), .Z(n1863) );
  NAND U2856 ( .A(n1903), .B(n1904), .Z(n1866) );
  MUX U2857 ( .IN0(n1853), .IN1(o[63]), .SEL(n1905), .F(\Data_Mem/n7728 ) );
  MUX U2858 ( .IN0(n1855), .IN1(o[62]), .SEL(n1905), .F(\Data_Mem/n7727 ) );
  MUX U2859 ( .IN0(n1856), .IN1(o[61]), .SEL(n1905), .F(\Data_Mem/n7726 ) );
  MUX U2860 ( .IN0(n1857), .IN1(o[60]), .SEL(n1905), .F(\Data_Mem/n7725 ) );
  MUX U2861 ( .IN0(n1858), .IN1(o[59]), .SEL(n1905), .F(\Data_Mem/n7724 ) );
  MUX U2862 ( .IN0(n1859), .IN1(o[58]), .SEL(n1905), .F(\Data_Mem/n7723 ) );
  MUX U2863 ( .IN0(n1860), .IN1(o[57]), .SEL(n1905), .F(\Data_Mem/n7722 ) );
  MUX U2864 ( .IN0(n1861), .IN1(o[56]), .SEL(n1905), .F(\Data_Mem/n7721 ) );
  ANDN U2865 ( .A(n1906), .B(n1907), .Z(n1905) );
  AND U2866 ( .A(n1908), .B(n1909), .Z(n1906) );
  OR U2867 ( .A(n1867), .B(n1910), .Z(n1909) );
  MUX U2868 ( .IN0(n1868), .IN1(o[55]), .SEL(n1911), .F(\Data_Mem/n7720 ) );
  MUX U2869 ( .IN0(n1870), .IN1(o[54]), .SEL(n1911), .F(\Data_Mem/n7719 ) );
  MUX U2870 ( .IN0(n1871), .IN1(o[53]), .SEL(n1911), .F(\Data_Mem/n7718 ) );
  MUX U2871 ( .IN0(n1872), .IN1(o[52]), .SEL(n1911), .F(\Data_Mem/n7717 ) );
  MUX U2872 ( .IN0(n1873), .IN1(o[51]), .SEL(n1911), .F(\Data_Mem/n7716 ) );
  IV U2873 ( .A(n1912), .Z(n1911) );
  MUX U2874 ( .IN0(o[50]), .IN1(n1875), .SEL(n1912), .F(\Data_Mem/n7715 ) );
  MUX U2875 ( .IN0(o[49]), .IN1(n1876), .SEL(n1912), .F(\Data_Mem/n7714 ) );
  MUX U2876 ( .IN0(o[48]), .IN1(n1877), .SEL(n1912), .F(\Data_Mem/n7713 ) );
  NAND U2877 ( .A(n1913), .B(n1914), .Z(n1912) );
  OR U2878 ( .A(n1880), .B(n1910), .Z(n1914) );
  ANDN U2879 ( .A(n1908), .B(n1907), .Z(n1913) );
  NANDN U2880 ( .B(n1910), .A(n1915), .Z(n1908) );
  MUX U2881 ( .IN0(n1883), .IN1(o[47]), .SEL(n1916), .F(\Data_Mem/n7712 ) );
  MUX U2882 ( .IN0(n1885), .IN1(o[46]), .SEL(n1916), .F(\Data_Mem/n7711 ) );
  MUX U2883 ( .IN0(n1886), .IN1(o[45]), .SEL(n1916), .F(\Data_Mem/n7710 ) );
  MUX U2884 ( .IN0(n1887), .IN1(o[44]), .SEL(n1916), .F(\Data_Mem/n7709 ) );
  MUX U2885 ( .IN0(n1888), .IN1(o[43]), .SEL(n1916), .F(\Data_Mem/n7708 ) );
  IV U2886 ( .A(n1917), .Z(n1916) );
  MUX U2887 ( .IN0(o[42]), .IN1(n1890), .SEL(n1917), .F(\Data_Mem/n7707 ) );
  MUX U2888 ( .IN0(o[41]), .IN1(n1891), .SEL(n1917), .F(\Data_Mem/n7706 ) );
  MUX U2889 ( .IN0(o[40]), .IN1(n1892), .SEL(n1917), .F(\Data_Mem/n7705 ) );
  NAND U2890 ( .A(n1918), .B(n1919), .Z(n1917) );
  OR U2891 ( .A(n1895), .B(n1910), .Z(n1919) );
  MUX U2892 ( .IN0(reg_target[7]), .IN1(o[39]), .SEL(n1920), .F(
        \Data_Mem/n7704 ) );
  MUX U2893 ( .IN0(reg_target[6]), .IN1(o[38]), .SEL(n1920), .F(
        \Data_Mem/n7703 ) );
  MUX U2894 ( .IN0(reg_target[5]), .IN1(o[37]), .SEL(n1920), .F(
        \Data_Mem/n7702 ) );
  MUX U2895 ( .IN0(reg_target[4]), .IN1(o[36]), .SEL(n1920), .F(
        \Data_Mem/n7701 ) );
  MUX U2896 ( .IN0(reg_target[3]), .IN1(o[35]), .SEL(n1920), .F(
        \Data_Mem/n7700 ) );
  IV U2897 ( .A(n1921), .Z(n1920) );
  MUX U2898 ( .IN0(o[34]), .IN1(reg_target[2]), .SEL(n1921), .F(
        \Data_Mem/n7699 ) );
  MUX U2899 ( .IN0(o[33]), .IN1(reg_target[1]), .SEL(n1921), .F(
        \Data_Mem/n7698 ) );
  MUX U2900 ( .IN0(o[32]), .IN1(reg_target[0]), .SEL(n1921), .F(
        \Data_Mem/n7697 ) );
  NAND U2901 ( .A(n1918), .B(n1922), .Z(n1921) );
  NANDN U2902 ( .B(n1910), .A(n1899), .Z(n1922) );
  ANDN U2903 ( .A(n1923), .B(n1907), .Z(n1918) );
  ANDN U2904 ( .A(n1902), .B(n1910), .Z(n1907) );
  NANDN U2905 ( .B(n1910), .A(n1924), .Z(n1923) );
  NAND U2906 ( .A(n1904), .B(n1925), .Z(n1910) );
  MUX U2907 ( .IN0(n1853), .IN1(o[95]), .SEL(n1926), .F(\Data_Mem/n7696 ) );
  MUX U2908 ( .IN0(n1855), .IN1(o[94]), .SEL(n1926), .F(\Data_Mem/n7695 ) );
  MUX U2909 ( .IN0(n1856), .IN1(o[93]), .SEL(n1926), .F(\Data_Mem/n7694 ) );
  MUX U2910 ( .IN0(n1857), .IN1(o[92]), .SEL(n1926), .F(\Data_Mem/n7693 ) );
  MUX U2911 ( .IN0(n1858), .IN1(o[91]), .SEL(n1926), .F(\Data_Mem/n7692 ) );
  MUX U2912 ( .IN0(n1859), .IN1(o[90]), .SEL(n1926), .F(\Data_Mem/n7691 ) );
  MUX U2913 ( .IN0(n1860), .IN1(o[89]), .SEL(n1926), .F(\Data_Mem/n7690 ) );
  MUX U2914 ( .IN0(n1861), .IN1(o[88]), .SEL(n1926), .F(\Data_Mem/n7689 ) );
  ANDN U2915 ( .A(n1927), .B(n1928), .Z(n1926) );
  AND U2916 ( .A(n1929), .B(n1930), .Z(n1927) );
  OR U2917 ( .A(n1867), .B(n1931), .Z(n1930) );
  MUX U2918 ( .IN0(n1868), .IN1(o[87]), .SEL(n1932), .F(\Data_Mem/n7688 ) );
  MUX U2919 ( .IN0(n1870), .IN1(o[86]), .SEL(n1932), .F(\Data_Mem/n7687 ) );
  MUX U2920 ( .IN0(n1871), .IN1(o[85]), .SEL(n1932), .F(\Data_Mem/n7686 ) );
  MUX U2921 ( .IN0(n1872), .IN1(o[84]), .SEL(n1932), .F(\Data_Mem/n7685 ) );
  MUX U2922 ( .IN0(n1873), .IN1(o[83]), .SEL(n1932), .F(\Data_Mem/n7684 ) );
  IV U2923 ( .A(n1933), .Z(n1932) );
  MUX U2924 ( .IN0(o[82]), .IN1(n1875), .SEL(n1933), .F(\Data_Mem/n7683 ) );
  MUX U2925 ( .IN0(o[81]), .IN1(n1876), .SEL(n1933), .F(\Data_Mem/n7682 ) );
  MUX U2926 ( .IN0(o[80]), .IN1(n1877), .SEL(n1933), .F(\Data_Mem/n7681 ) );
  NAND U2927 ( .A(n1934), .B(n1935), .Z(n1933) );
  OR U2928 ( .A(n1880), .B(n1931), .Z(n1935) );
  ANDN U2929 ( .A(n1929), .B(n1928), .Z(n1934) );
  NANDN U2930 ( .B(n1931), .A(n1915), .Z(n1929) );
  MUX U2931 ( .IN0(n1883), .IN1(o[79]), .SEL(n1936), .F(\Data_Mem/n7680 ) );
  MUX U2932 ( .IN0(n1885), .IN1(o[78]), .SEL(n1936), .F(\Data_Mem/n7679 ) );
  MUX U2933 ( .IN0(n1886), .IN1(o[77]), .SEL(n1936), .F(\Data_Mem/n7678 ) );
  MUX U2934 ( .IN0(n1887), .IN1(o[76]), .SEL(n1936), .F(\Data_Mem/n7677 ) );
  MUX U2935 ( .IN0(n1888), .IN1(o[75]), .SEL(n1936), .F(\Data_Mem/n7676 ) );
  IV U2936 ( .A(n1937), .Z(n1936) );
  MUX U2937 ( .IN0(o[74]), .IN1(n1890), .SEL(n1937), .F(\Data_Mem/n7675 ) );
  MUX U2938 ( .IN0(o[73]), .IN1(n1891), .SEL(n1937), .F(\Data_Mem/n7674 ) );
  MUX U2939 ( .IN0(o[72]), .IN1(n1892), .SEL(n1937), .F(\Data_Mem/n7673 ) );
  NAND U2940 ( .A(n1938), .B(n1939), .Z(n1937) );
  OR U2941 ( .A(n1895), .B(n1931), .Z(n1939) );
  MUX U2942 ( .IN0(reg_target[7]), .IN1(o[71]), .SEL(n1940), .F(
        \Data_Mem/n7672 ) );
  MUX U2943 ( .IN0(reg_target[6]), .IN1(o[70]), .SEL(n1940), .F(
        \Data_Mem/n7671 ) );
  MUX U2944 ( .IN0(reg_target[5]), .IN1(o[69]), .SEL(n1940), .F(
        \Data_Mem/n7670 ) );
  MUX U2945 ( .IN0(reg_target[4]), .IN1(o[68]), .SEL(n1940), .F(
        \Data_Mem/n7669 ) );
  MUX U2946 ( .IN0(reg_target[3]), .IN1(o[67]), .SEL(n1940), .F(
        \Data_Mem/n7668 ) );
  IV U2947 ( .A(n1941), .Z(n1940) );
  MUX U2948 ( .IN0(o[66]), .IN1(reg_target[2]), .SEL(n1941), .F(
        \Data_Mem/n7667 ) );
  MUX U2949 ( .IN0(o[65]), .IN1(reg_target[1]), .SEL(n1941), .F(
        \Data_Mem/n7666 ) );
  MUX U2950 ( .IN0(o[64]), .IN1(reg_target[0]), .SEL(n1941), .F(
        \Data_Mem/n7665 ) );
  NAND U2951 ( .A(n1938), .B(n1942), .Z(n1941) );
  NANDN U2952 ( .B(n1931), .A(n1899), .Z(n1942) );
  ANDN U2953 ( .A(n1943), .B(n1928), .Z(n1938) );
  ANDN U2954 ( .A(n1902), .B(n1931), .Z(n1928) );
  NANDN U2955 ( .B(n1931), .A(n1924), .Z(n1943) );
  NAND U2956 ( .A(n1904), .B(n1944), .Z(n1931) );
  MUX U2957 ( .IN0(n1853), .IN1(o[127]), .SEL(n1945), .F(\Data_Mem/n7664 ) );
  MUX U2958 ( .IN0(n1855), .IN1(o[126]), .SEL(n1945), .F(\Data_Mem/n7663 ) );
  MUX U2959 ( .IN0(n1856), .IN1(o[125]), .SEL(n1945), .F(\Data_Mem/n7662 ) );
  MUX U2960 ( .IN0(n1857), .IN1(o[124]), .SEL(n1945), .F(\Data_Mem/n7661 ) );
  MUX U2961 ( .IN0(n1858), .IN1(o[123]), .SEL(n1945), .F(\Data_Mem/n7660 ) );
  MUX U2962 ( .IN0(n1859), .IN1(o[122]), .SEL(n1945), .F(\Data_Mem/n7659 ) );
  MUX U2963 ( .IN0(n1860), .IN1(o[121]), .SEL(n1945), .F(\Data_Mem/n7658 ) );
  MUX U2964 ( .IN0(n1861), .IN1(o[120]), .SEL(n1945), .F(\Data_Mem/n7657 ) );
  ANDN U2965 ( .A(n1946), .B(n1947), .Z(n1945) );
  AND U2966 ( .A(n1948), .B(n1949), .Z(n1946) );
  OR U2967 ( .A(n1867), .B(n1950), .Z(n1949) );
  MUX U2968 ( .IN0(n1868), .IN1(o[119]), .SEL(n1951), .F(\Data_Mem/n7656 ) );
  MUX U2969 ( .IN0(n1870), .IN1(o[118]), .SEL(n1951), .F(\Data_Mem/n7655 ) );
  MUX U2970 ( .IN0(n1871), .IN1(o[117]), .SEL(n1951), .F(\Data_Mem/n7654 ) );
  MUX U2971 ( .IN0(n1872), .IN1(o[116]), .SEL(n1951), .F(\Data_Mem/n7653 ) );
  MUX U2972 ( .IN0(n1873), .IN1(o[115]), .SEL(n1951), .F(\Data_Mem/n7652 ) );
  IV U2973 ( .A(n1952), .Z(n1951) );
  MUX U2974 ( .IN0(o[114]), .IN1(n1875), .SEL(n1952), .F(\Data_Mem/n7651 ) );
  MUX U2975 ( .IN0(o[113]), .IN1(n1876), .SEL(n1952), .F(\Data_Mem/n7650 ) );
  MUX U2976 ( .IN0(o[112]), .IN1(n1877), .SEL(n1952), .F(\Data_Mem/n7649 ) );
  NAND U2977 ( .A(n1953), .B(n1954), .Z(n1952) );
  OR U2978 ( .A(n1880), .B(n1950), .Z(n1954) );
  ANDN U2979 ( .A(n1948), .B(n1947), .Z(n1953) );
  NANDN U2980 ( .B(n1950), .A(n1915), .Z(n1948) );
  MUX U2981 ( .IN0(n1883), .IN1(o[111]), .SEL(n1955), .F(\Data_Mem/n7648 ) );
  MUX U2982 ( .IN0(n1885), .IN1(o[110]), .SEL(n1955), .F(\Data_Mem/n7647 ) );
  MUX U2983 ( .IN0(n1886), .IN1(o[109]), .SEL(n1955), .F(\Data_Mem/n7646 ) );
  MUX U2984 ( .IN0(n1887), .IN1(o[108]), .SEL(n1955), .F(\Data_Mem/n7645 ) );
  MUX U2985 ( .IN0(n1888), .IN1(o[107]), .SEL(n1955), .F(\Data_Mem/n7644 ) );
  IV U2986 ( .A(n1956), .Z(n1955) );
  MUX U2987 ( .IN0(o[106]), .IN1(n1890), .SEL(n1956), .F(\Data_Mem/n7643 ) );
  MUX U2988 ( .IN0(o[105]), .IN1(n1891), .SEL(n1956), .F(\Data_Mem/n7642 ) );
  MUX U2989 ( .IN0(o[104]), .IN1(n1892), .SEL(n1956), .F(\Data_Mem/n7641 ) );
  NAND U2990 ( .A(n1957), .B(n1958), .Z(n1956) );
  OR U2991 ( .A(n1895), .B(n1950), .Z(n1958) );
  MUX U2992 ( .IN0(reg_target[7]), .IN1(o[103]), .SEL(n1959), .F(
        \Data_Mem/n7640 ) );
  MUX U2993 ( .IN0(reg_target[6]), .IN1(o[102]), .SEL(n1959), .F(
        \Data_Mem/n7639 ) );
  MUX U2994 ( .IN0(reg_target[5]), .IN1(o[101]), .SEL(n1959), .F(
        \Data_Mem/n7638 ) );
  MUX U2995 ( .IN0(reg_target[4]), .IN1(o[100]), .SEL(n1959), .F(
        \Data_Mem/n7637 ) );
  MUX U2996 ( .IN0(reg_target[3]), .IN1(o[99]), .SEL(n1959), .F(
        \Data_Mem/n7636 ) );
  IV U2997 ( .A(n1960), .Z(n1959) );
  MUX U2998 ( .IN0(o[98]), .IN1(reg_target[2]), .SEL(n1960), .F(
        \Data_Mem/n7635 ) );
  MUX U2999 ( .IN0(o[97]), .IN1(reg_target[1]), .SEL(n1960), .F(
        \Data_Mem/n7634 ) );
  MUX U3000 ( .IN0(o[96]), .IN1(reg_target[0]), .SEL(n1960), .F(
        \Data_Mem/n7633 ) );
  NAND U3001 ( .A(n1957), .B(n1961), .Z(n1960) );
  NANDN U3002 ( .B(n1950), .A(n1899), .Z(n1961) );
  ANDN U3003 ( .A(n1962), .B(n1947), .Z(n1957) );
  ANDN U3004 ( .A(n1902), .B(n1950), .Z(n1947) );
  NANDN U3005 ( .B(n1950), .A(n1924), .Z(n1962) );
  NAND U3006 ( .A(n1904), .B(n1963), .Z(n1950) );
  MUX U3007 ( .IN0(n1853), .IN1(o[159]), .SEL(n1964), .F(\Data_Mem/n7632 ) );
  MUX U3008 ( .IN0(n1855), .IN1(o[158]), .SEL(n1964), .F(\Data_Mem/n7631 ) );
  MUX U3009 ( .IN0(n1856), .IN1(o[157]), .SEL(n1964), .F(\Data_Mem/n7630 ) );
  MUX U3010 ( .IN0(n1857), .IN1(o[156]), .SEL(n1964), .F(\Data_Mem/n7629 ) );
  MUX U3011 ( .IN0(n1858), .IN1(o[155]), .SEL(n1964), .F(\Data_Mem/n7628 ) );
  MUX U3012 ( .IN0(n1859), .IN1(o[154]), .SEL(n1964), .F(\Data_Mem/n7627 ) );
  MUX U3013 ( .IN0(n1860), .IN1(o[153]), .SEL(n1964), .F(\Data_Mem/n7626 ) );
  MUX U3014 ( .IN0(n1861), .IN1(o[152]), .SEL(n1964), .F(\Data_Mem/n7625 ) );
  ANDN U3015 ( .A(n1965), .B(n1966), .Z(n1964) );
  AND U3016 ( .A(n1967), .B(n1968), .Z(n1965) );
  OR U3017 ( .A(n1867), .B(n1969), .Z(n1968) );
  MUX U3018 ( .IN0(n1868), .IN1(o[151]), .SEL(n1970), .F(\Data_Mem/n7624 ) );
  MUX U3019 ( .IN0(n1870), .IN1(o[150]), .SEL(n1970), .F(\Data_Mem/n7623 ) );
  MUX U3020 ( .IN0(n1871), .IN1(o[149]), .SEL(n1970), .F(\Data_Mem/n7622 ) );
  MUX U3021 ( .IN0(n1872), .IN1(o[148]), .SEL(n1970), .F(\Data_Mem/n7621 ) );
  MUX U3022 ( .IN0(n1873), .IN1(o[147]), .SEL(n1970), .F(\Data_Mem/n7620 ) );
  IV U3023 ( .A(n1971), .Z(n1970) );
  MUX U3024 ( .IN0(o[146]), .IN1(n1875), .SEL(n1971), .F(\Data_Mem/n7619 ) );
  MUX U3025 ( .IN0(o[145]), .IN1(n1876), .SEL(n1971), .F(\Data_Mem/n7618 ) );
  MUX U3026 ( .IN0(o[144]), .IN1(n1877), .SEL(n1971), .F(\Data_Mem/n7617 ) );
  NAND U3027 ( .A(n1972), .B(n1973), .Z(n1971) );
  OR U3028 ( .A(n1880), .B(n1969), .Z(n1973) );
  ANDN U3029 ( .A(n1967), .B(n1966), .Z(n1972) );
  NANDN U3030 ( .B(n1969), .A(n1915), .Z(n1967) );
  MUX U3031 ( .IN0(n1883), .IN1(o[143]), .SEL(n1974), .F(\Data_Mem/n7616 ) );
  MUX U3032 ( .IN0(n1885), .IN1(o[142]), .SEL(n1974), .F(\Data_Mem/n7615 ) );
  MUX U3033 ( .IN0(n1886), .IN1(o[141]), .SEL(n1974), .F(\Data_Mem/n7614 ) );
  MUX U3034 ( .IN0(n1887), .IN1(o[140]), .SEL(n1974), .F(\Data_Mem/n7613 ) );
  MUX U3035 ( .IN0(n1888), .IN1(o[139]), .SEL(n1974), .F(\Data_Mem/n7612 ) );
  IV U3036 ( .A(n1975), .Z(n1974) );
  MUX U3037 ( .IN0(o[138]), .IN1(n1890), .SEL(n1975), .F(\Data_Mem/n7611 ) );
  MUX U3038 ( .IN0(o[137]), .IN1(n1891), .SEL(n1975), .F(\Data_Mem/n7610 ) );
  MUX U3039 ( .IN0(o[136]), .IN1(n1892), .SEL(n1975), .F(\Data_Mem/n7609 ) );
  NAND U3040 ( .A(n1976), .B(n1977), .Z(n1975) );
  OR U3041 ( .A(n1895), .B(n1969), .Z(n1977) );
  MUX U3042 ( .IN0(reg_target[7]), .IN1(o[135]), .SEL(n1978), .F(
        \Data_Mem/n7608 ) );
  MUX U3043 ( .IN0(reg_target[6]), .IN1(o[134]), .SEL(n1978), .F(
        \Data_Mem/n7607 ) );
  MUX U3044 ( .IN0(reg_target[5]), .IN1(o[133]), .SEL(n1978), .F(
        \Data_Mem/n7606 ) );
  MUX U3045 ( .IN0(reg_target[4]), .IN1(o[132]), .SEL(n1978), .F(
        \Data_Mem/n7605 ) );
  MUX U3046 ( .IN0(reg_target[3]), .IN1(o[131]), .SEL(n1978), .F(
        \Data_Mem/n7604 ) );
  IV U3047 ( .A(n1979), .Z(n1978) );
  MUX U3048 ( .IN0(o[130]), .IN1(reg_target[2]), .SEL(n1979), .F(
        \Data_Mem/n7603 ) );
  MUX U3049 ( .IN0(o[129]), .IN1(reg_target[1]), .SEL(n1979), .F(
        \Data_Mem/n7602 ) );
  MUX U3050 ( .IN0(o[128]), .IN1(reg_target[0]), .SEL(n1979), .F(
        \Data_Mem/n7601 ) );
  NAND U3051 ( .A(n1976), .B(n1980), .Z(n1979) );
  NANDN U3052 ( .B(n1969), .A(n1899), .Z(n1980) );
  ANDN U3053 ( .A(n1981), .B(n1966), .Z(n1976) );
  ANDN U3054 ( .A(n1902), .B(n1969), .Z(n1966) );
  NANDN U3055 ( .B(n1969), .A(n1924), .Z(n1981) );
  NAND U3056 ( .A(n1904), .B(n1982), .Z(n1969) );
  MUX U3057 ( .IN0(n1853), .IN1(o[191]), .SEL(n1983), .F(\Data_Mem/n7600 ) );
  MUX U3058 ( .IN0(n1855), .IN1(o[190]), .SEL(n1983), .F(\Data_Mem/n7599 ) );
  MUX U3059 ( .IN0(n1856), .IN1(o[189]), .SEL(n1983), .F(\Data_Mem/n7598 ) );
  MUX U3060 ( .IN0(n1857), .IN1(o[188]), .SEL(n1983), .F(\Data_Mem/n7597 ) );
  MUX U3061 ( .IN0(n1858), .IN1(o[187]), .SEL(n1983), .F(\Data_Mem/n7596 ) );
  MUX U3062 ( .IN0(n1859), .IN1(o[186]), .SEL(n1983), .F(\Data_Mem/n7595 ) );
  MUX U3063 ( .IN0(n1860), .IN1(o[185]), .SEL(n1983), .F(\Data_Mem/n7594 ) );
  MUX U3064 ( .IN0(n1861), .IN1(o[184]), .SEL(n1983), .F(\Data_Mem/n7593 ) );
  ANDN U3065 ( .A(n1984), .B(n1985), .Z(n1983) );
  AND U3066 ( .A(n1986), .B(n1987), .Z(n1984) );
  OR U3067 ( .A(n1867), .B(n1988), .Z(n1987) );
  MUX U3068 ( .IN0(n1868), .IN1(o[183]), .SEL(n1989), .F(\Data_Mem/n7592 ) );
  MUX U3069 ( .IN0(n1870), .IN1(o[182]), .SEL(n1989), .F(\Data_Mem/n7591 ) );
  MUX U3070 ( .IN0(n1871), .IN1(o[181]), .SEL(n1989), .F(\Data_Mem/n7590 ) );
  MUX U3071 ( .IN0(n1872), .IN1(o[180]), .SEL(n1989), .F(\Data_Mem/n7589 ) );
  MUX U3072 ( .IN0(n1873), .IN1(o[179]), .SEL(n1989), .F(\Data_Mem/n7588 ) );
  IV U3073 ( .A(n1990), .Z(n1989) );
  MUX U3074 ( .IN0(o[178]), .IN1(n1875), .SEL(n1990), .F(\Data_Mem/n7587 ) );
  MUX U3075 ( .IN0(o[177]), .IN1(n1876), .SEL(n1990), .F(\Data_Mem/n7586 ) );
  MUX U3076 ( .IN0(o[176]), .IN1(n1877), .SEL(n1990), .F(\Data_Mem/n7585 ) );
  NAND U3077 ( .A(n1991), .B(n1992), .Z(n1990) );
  OR U3078 ( .A(n1880), .B(n1988), .Z(n1992) );
  ANDN U3079 ( .A(n1986), .B(n1985), .Z(n1991) );
  NANDN U3080 ( .B(n1988), .A(n1915), .Z(n1986) );
  MUX U3081 ( .IN0(n1883), .IN1(o[175]), .SEL(n1993), .F(\Data_Mem/n7584 ) );
  MUX U3082 ( .IN0(n1885), .IN1(o[174]), .SEL(n1993), .F(\Data_Mem/n7583 ) );
  MUX U3083 ( .IN0(n1886), .IN1(o[173]), .SEL(n1993), .F(\Data_Mem/n7582 ) );
  MUX U3084 ( .IN0(n1887), .IN1(o[172]), .SEL(n1993), .F(\Data_Mem/n7581 ) );
  MUX U3085 ( .IN0(n1888), .IN1(o[171]), .SEL(n1993), .F(\Data_Mem/n7580 ) );
  IV U3086 ( .A(n1994), .Z(n1993) );
  MUX U3087 ( .IN0(o[170]), .IN1(n1890), .SEL(n1994), .F(\Data_Mem/n7579 ) );
  MUX U3088 ( .IN0(o[169]), .IN1(n1891), .SEL(n1994), .F(\Data_Mem/n7578 ) );
  MUX U3089 ( .IN0(o[168]), .IN1(n1892), .SEL(n1994), .F(\Data_Mem/n7577 ) );
  NAND U3090 ( .A(n1995), .B(n1996), .Z(n1994) );
  OR U3091 ( .A(n1895), .B(n1988), .Z(n1996) );
  MUX U3092 ( .IN0(reg_target[7]), .IN1(o[167]), .SEL(n1997), .F(
        \Data_Mem/n7576 ) );
  MUX U3093 ( .IN0(reg_target[6]), .IN1(o[166]), .SEL(n1997), .F(
        \Data_Mem/n7575 ) );
  MUX U3094 ( .IN0(reg_target[5]), .IN1(o[165]), .SEL(n1997), .F(
        \Data_Mem/n7574 ) );
  MUX U3095 ( .IN0(reg_target[4]), .IN1(o[164]), .SEL(n1997), .F(
        \Data_Mem/n7573 ) );
  MUX U3096 ( .IN0(reg_target[3]), .IN1(o[163]), .SEL(n1997), .F(
        \Data_Mem/n7572 ) );
  IV U3097 ( .A(n1998), .Z(n1997) );
  MUX U3098 ( .IN0(o[162]), .IN1(reg_target[2]), .SEL(n1998), .F(
        \Data_Mem/n7571 ) );
  MUX U3099 ( .IN0(o[161]), .IN1(reg_target[1]), .SEL(n1998), .F(
        \Data_Mem/n7570 ) );
  MUX U3100 ( .IN0(o[160]), .IN1(reg_target[0]), .SEL(n1998), .F(
        \Data_Mem/n7569 ) );
  NAND U3101 ( .A(n1995), .B(n1999), .Z(n1998) );
  NANDN U3102 ( .B(n1988), .A(n1899), .Z(n1999) );
  ANDN U3103 ( .A(n2000), .B(n1985), .Z(n1995) );
  ANDN U3104 ( .A(n1902), .B(n1988), .Z(n1985) );
  NANDN U3105 ( .B(n1988), .A(n1924), .Z(n2000) );
  NAND U3106 ( .A(n1904), .B(n2001), .Z(n1988) );
  MUX U3107 ( .IN0(n1853), .IN1(o[223]), .SEL(n2002), .F(\Data_Mem/n7568 ) );
  MUX U3108 ( .IN0(n1855), .IN1(o[222]), .SEL(n2002), .F(\Data_Mem/n7567 ) );
  MUX U3109 ( .IN0(n1856), .IN1(o[221]), .SEL(n2002), .F(\Data_Mem/n7566 ) );
  MUX U3110 ( .IN0(n1857), .IN1(o[220]), .SEL(n2002), .F(\Data_Mem/n7565 ) );
  MUX U3111 ( .IN0(n1858), .IN1(o[219]), .SEL(n2002), .F(\Data_Mem/n7564 ) );
  MUX U3112 ( .IN0(n1859), .IN1(o[218]), .SEL(n2002), .F(\Data_Mem/n7563 ) );
  MUX U3113 ( .IN0(n1860), .IN1(o[217]), .SEL(n2002), .F(\Data_Mem/n7562 ) );
  MUX U3114 ( .IN0(n1861), .IN1(o[216]), .SEL(n2002), .F(\Data_Mem/n7561 ) );
  ANDN U3115 ( .A(n2003), .B(n2004), .Z(n2002) );
  AND U3116 ( .A(n2005), .B(n2006), .Z(n2003) );
  OR U3117 ( .A(n1867), .B(n2007), .Z(n2006) );
  MUX U3118 ( .IN0(n1868), .IN1(o[215]), .SEL(n2008), .F(\Data_Mem/n7560 ) );
  MUX U3119 ( .IN0(n1870), .IN1(o[214]), .SEL(n2008), .F(\Data_Mem/n7559 ) );
  MUX U3120 ( .IN0(n1871), .IN1(o[213]), .SEL(n2008), .F(\Data_Mem/n7558 ) );
  MUX U3121 ( .IN0(n1872), .IN1(o[212]), .SEL(n2008), .F(\Data_Mem/n7557 ) );
  MUX U3122 ( .IN0(n1873), .IN1(o[211]), .SEL(n2008), .F(\Data_Mem/n7556 ) );
  IV U3123 ( .A(n2009), .Z(n2008) );
  MUX U3124 ( .IN0(o[210]), .IN1(n1875), .SEL(n2009), .F(\Data_Mem/n7555 ) );
  MUX U3125 ( .IN0(o[209]), .IN1(n1876), .SEL(n2009), .F(\Data_Mem/n7554 ) );
  MUX U3126 ( .IN0(o[208]), .IN1(n1877), .SEL(n2009), .F(\Data_Mem/n7553 ) );
  NAND U3127 ( .A(n2010), .B(n2011), .Z(n2009) );
  OR U3128 ( .A(n1880), .B(n2007), .Z(n2011) );
  ANDN U3129 ( .A(n2005), .B(n2004), .Z(n2010) );
  NANDN U3130 ( .B(n2007), .A(n1915), .Z(n2005) );
  MUX U3131 ( .IN0(n1883), .IN1(o[207]), .SEL(n2012), .F(\Data_Mem/n7552 ) );
  MUX U3132 ( .IN0(n1885), .IN1(o[206]), .SEL(n2012), .F(\Data_Mem/n7551 ) );
  MUX U3133 ( .IN0(n1886), .IN1(o[205]), .SEL(n2012), .F(\Data_Mem/n7550 ) );
  MUX U3134 ( .IN0(n1887), .IN1(o[204]), .SEL(n2012), .F(\Data_Mem/n7549 ) );
  MUX U3135 ( .IN0(n1888), .IN1(o[203]), .SEL(n2012), .F(\Data_Mem/n7548 ) );
  IV U3136 ( .A(n2013), .Z(n2012) );
  MUX U3137 ( .IN0(o[202]), .IN1(n1890), .SEL(n2013), .F(\Data_Mem/n7547 ) );
  MUX U3138 ( .IN0(o[201]), .IN1(n1891), .SEL(n2013), .F(\Data_Mem/n7546 ) );
  MUX U3139 ( .IN0(o[200]), .IN1(n1892), .SEL(n2013), .F(\Data_Mem/n7545 ) );
  NAND U3140 ( .A(n2014), .B(n2015), .Z(n2013) );
  OR U3141 ( .A(n1895), .B(n2007), .Z(n2015) );
  MUX U3142 ( .IN0(reg_target[7]), .IN1(o[199]), .SEL(n2016), .F(
        \Data_Mem/n7544 ) );
  MUX U3143 ( .IN0(reg_target[6]), .IN1(o[198]), .SEL(n2016), .F(
        \Data_Mem/n7543 ) );
  MUX U3144 ( .IN0(reg_target[5]), .IN1(o[197]), .SEL(n2016), .F(
        \Data_Mem/n7542 ) );
  MUX U3145 ( .IN0(reg_target[4]), .IN1(o[196]), .SEL(n2016), .F(
        \Data_Mem/n7541 ) );
  MUX U3146 ( .IN0(reg_target[3]), .IN1(o[195]), .SEL(n2016), .F(
        \Data_Mem/n7540 ) );
  IV U3147 ( .A(n2017), .Z(n2016) );
  MUX U3148 ( .IN0(o[194]), .IN1(reg_target[2]), .SEL(n2017), .F(
        \Data_Mem/n7539 ) );
  MUX U3149 ( .IN0(o[193]), .IN1(reg_target[1]), .SEL(n2017), .F(
        \Data_Mem/n7538 ) );
  MUX U3150 ( .IN0(o[192]), .IN1(reg_target[0]), .SEL(n2017), .F(
        \Data_Mem/n7537 ) );
  NAND U3151 ( .A(n2014), .B(n2018), .Z(n2017) );
  NANDN U3152 ( .B(n2007), .A(n1899), .Z(n2018) );
  ANDN U3153 ( .A(n2019), .B(n2004), .Z(n2014) );
  ANDN U3154 ( .A(n1902), .B(n2007), .Z(n2004) );
  NANDN U3155 ( .B(n2007), .A(n1924), .Z(n2019) );
  NAND U3156 ( .A(n1904), .B(n2020), .Z(n2007) );
  MUX U3157 ( .IN0(n1853), .IN1(o[255]), .SEL(n2021), .F(\Data_Mem/n7536 ) );
  MUX U3158 ( .IN0(n1855), .IN1(o[254]), .SEL(n2021), .F(\Data_Mem/n7535 ) );
  MUX U3159 ( .IN0(n1856), .IN1(o[253]), .SEL(n2021), .F(\Data_Mem/n7534 ) );
  MUX U3160 ( .IN0(n1857), .IN1(o[252]), .SEL(n2021), .F(\Data_Mem/n7533 ) );
  MUX U3161 ( .IN0(n1858), .IN1(o[251]), .SEL(n2021), .F(\Data_Mem/n7532 ) );
  MUX U3162 ( .IN0(n1859), .IN1(o[250]), .SEL(n2021), .F(\Data_Mem/n7531 ) );
  MUX U3163 ( .IN0(n1860), .IN1(o[249]), .SEL(n2021), .F(\Data_Mem/n7530 ) );
  MUX U3164 ( .IN0(n1861), .IN1(o[248]), .SEL(n2021), .F(\Data_Mem/n7529 ) );
  ANDN U3165 ( .A(n2022), .B(n2023), .Z(n2021) );
  AND U3166 ( .A(n2024), .B(n2025), .Z(n2022) );
  OR U3167 ( .A(n1867), .B(n2026), .Z(n2025) );
  MUX U3168 ( .IN0(n1868), .IN1(o[247]), .SEL(n2027), .F(\Data_Mem/n7528 ) );
  MUX U3169 ( .IN0(n1870), .IN1(o[246]), .SEL(n2027), .F(\Data_Mem/n7527 ) );
  MUX U3170 ( .IN0(n1871), .IN1(o[245]), .SEL(n2027), .F(\Data_Mem/n7526 ) );
  MUX U3171 ( .IN0(n1872), .IN1(o[244]), .SEL(n2027), .F(\Data_Mem/n7525 ) );
  MUX U3172 ( .IN0(n1873), .IN1(o[243]), .SEL(n2027), .F(\Data_Mem/n7524 ) );
  IV U3173 ( .A(n2028), .Z(n2027) );
  MUX U3174 ( .IN0(o[242]), .IN1(n1875), .SEL(n2028), .F(\Data_Mem/n7523 ) );
  MUX U3175 ( .IN0(o[241]), .IN1(n1876), .SEL(n2028), .F(\Data_Mem/n7522 ) );
  MUX U3176 ( .IN0(o[240]), .IN1(n1877), .SEL(n2028), .F(\Data_Mem/n7521 ) );
  NAND U3177 ( .A(n2029), .B(n2030), .Z(n2028) );
  OR U3178 ( .A(n1880), .B(n2026), .Z(n2030) );
  ANDN U3179 ( .A(n2024), .B(n2023), .Z(n2029) );
  NANDN U3180 ( .B(n2026), .A(n1915), .Z(n2024) );
  MUX U3181 ( .IN0(n1883), .IN1(o[239]), .SEL(n2031), .F(\Data_Mem/n7520 ) );
  MUX U3182 ( .IN0(n1885), .IN1(o[238]), .SEL(n2031), .F(\Data_Mem/n7519 ) );
  MUX U3183 ( .IN0(n1886), .IN1(o[237]), .SEL(n2031), .F(\Data_Mem/n7518 ) );
  MUX U3184 ( .IN0(n1887), .IN1(o[236]), .SEL(n2031), .F(\Data_Mem/n7517 ) );
  MUX U3185 ( .IN0(n1888), .IN1(o[235]), .SEL(n2031), .F(\Data_Mem/n7516 ) );
  IV U3186 ( .A(n2032), .Z(n2031) );
  MUX U3187 ( .IN0(o[234]), .IN1(n1890), .SEL(n2032), .F(\Data_Mem/n7515 ) );
  MUX U3188 ( .IN0(o[233]), .IN1(n1891), .SEL(n2032), .F(\Data_Mem/n7514 ) );
  MUX U3189 ( .IN0(o[232]), .IN1(n1892), .SEL(n2032), .F(\Data_Mem/n7513 ) );
  NAND U3190 ( .A(n2033), .B(n2034), .Z(n2032) );
  OR U3191 ( .A(n1895), .B(n2026), .Z(n2034) );
  MUX U3192 ( .IN0(reg_target[7]), .IN1(o[231]), .SEL(n2035), .F(
        \Data_Mem/n7512 ) );
  MUX U3193 ( .IN0(reg_target[6]), .IN1(o[230]), .SEL(n2035), .F(
        \Data_Mem/n7511 ) );
  MUX U3194 ( .IN0(reg_target[5]), .IN1(o[229]), .SEL(n2035), .F(
        \Data_Mem/n7510 ) );
  MUX U3195 ( .IN0(reg_target[4]), .IN1(o[228]), .SEL(n2035), .F(
        \Data_Mem/n7509 ) );
  MUX U3196 ( .IN0(reg_target[3]), .IN1(o[227]), .SEL(n2035), .F(
        \Data_Mem/n7508 ) );
  IV U3197 ( .A(n2036), .Z(n2035) );
  MUX U3198 ( .IN0(o[226]), .IN1(reg_target[2]), .SEL(n2036), .F(
        \Data_Mem/n7507 ) );
  MUX U3199 ( .IN0(o[225]), .IN1(reg_target[1]), .SEL(n2036), .F(
        \Data_Mem/n7506 ) );
  MUX U3200 ( .IN0(o[224]), .IN1(reg_target[0]), .SEL(n2036), .F(
        \Data_Mem/n7505 ) );
  NAND U3201 ( .A(n2033), .B(n2037), .Z(n2036) );
  NANDN U3202 ( .B(n2026), .A(n1899), .Z(n2037) );
  ANDN U3203 ( .A(n2038), .B(n2023), .Z(n2033) );
  ANDN U3204 ( .A(n1902), .B(n2026), .Z(n2023) );
  NANDN U3205 ( .B(n2026), .A(n1924), .Z(n2038) );
  NAND U3206 ( .A(n1904), .B(n2039), .Z(n2026) );
  AND U3207 ( .A(n2040), .B(n485), .Z(n1904) );
  MUX U3208 ( .IN0(n1853), .IN1(o[287]), .SEL(n2041), .F(\Data_Mem/n7504 ) );
  MUX U3209 ( .IN0(n1855), .IN1(o[286]), .SEL(n2041), .F(\Data_Mem/n7503 ) );
  MUX U3210 ( .IN0(n1856), .IN1(o[285]), .SEL(n2041), .F(\Data_Mem/n7502 ) );
  MUX U3211 ( .IN0(n1857), .IN1(o[284]), .SEL(n2041), .F(\Data_Mem/n7501 ) );
  MUX U3212 ( .IN0(n1858), .IN1(o[283]), .SEL(n2041), .F(\Data_Mem/n7500 ) );
  MUX U3213 ( .IN0(n1859), .IN1(o[282]), .SEL(n2041), .F(\Data_Mem/n7499 ) );
  MUX U3214 ( .IN0(n1860), .IN1(o[281]), .SEL(n2041), .F(\Data_Mem/n7498 ) );
  MUX U3215 ( .IN0(n1861), .IN1(o[280]), .SEL(n2041), .F(\Data_Mem/n7497 ) );
  ANDN U3216 ( .A(n2042), .B(n2043), .Z(n2041) );
  AND U3217 ( .A(n2044), .B(n2045), .Z(n2042) );
  OR U3218 ( .A(n1867), .B(n2046), .Z(n2045) );
  MUX U3219 ( .IN0(n1868), .IN1(o[279]), .SEL(n2047), .F(\Data_Mem/n7496 ) );
  MUX U3220 ( .IN0(n1870), .IN1(o[278]), .SEL(n2047), .F(\Data_Mem/n7495 ) );
  MUX U3221 ( .IN0(n1871), .IN1(o[277]), .SEL(n2047), .F(\Data_Mem/n7494 ) );
  MUX U3222 ( .IN0(n1872), .IN1(o[276]), .SEL(n2047), .F(\Data_Mem/n7493 ) );
  MUX U3223 ( .IN0(n1873), .IN1(o[275]), .SEL(n2047), .F(\Data_Mem/n7492 ) );
  IV U3224 ( .A(n2048), .Z(n2047) );
  MUX U3225 ( .IN0(o[274]), .IN1(n1875), .SEL(n2048), .F(\Data_Mem/n7491 ) );
  MUX U3226 ( .IN0(o[273]), .IN1(n1876), .SEL(n2048), .F(\Data_Mem/n7490 ) );
  MUX U3227 ( .IN0(o[272]), .IN1(n1877), .SEL(n2048), .F(\Data_Mem/n7489 ) );
  NAND U3228 ( .A(n2049), .B(n2050), .Z(n2048) );
  OR U3229 ( .A(n1880), .B(n2046), .Z(n2050) );
  ANDN U3230 ( .A(n2044), .B(n2043), .Z(n2049) );
  NANDN U3231 ( .B(n2046), .A(n1915), .Z(n2044) );
  MUX U3232 ( .IN0(n1883), .IN1(o[271]), .SEL(n2051), .F(\Data_Mem/n7488 ) );
  MUX U3233 ( .IN0(n1885), .IN1(o[270]), .SEL(n2051), .F(\Data_Mem/n7487 ) );
  MUX U3234 ( .IN0(n1886), .IN1(o[269]), .SEL(n2051), .F(\Data_Mem/n7486 ) );
  MUX U3235 ( .IN0(n1887), .IN1(o[268]), .SEL(n2051), .F(\Data_Mem/n7485 ) );
  MUX U3236 ( .IN0(n1888), .IN1(o[267]), .SEL(n2051), .F(\Data_Mem/n7484 ) );
  IV U3237 ( .A(n2052), .Z(n2051) );
  MUX U3238 ( .IN0(o[266]), .IN1(n1890), .SEL(n2052), .F(\Data_Mem/n7483 ) );
  MUX U3239 ( .IN0(o[265]), .IN1(n1891), .SEL(n2052), .F(\Data_Mem/n7482 ) );
  MUX U3240 ( .IN0(o[264]), .IN1(n1892), .SEL(n2052), .F(\Data_Mem/n7481 ) );
  NAND U3241 ( .A(n2053), .B(n2054), .Z(n2052) );
  OR U3242 ( .A(n1895), .B(n2046), .Z(n2054) );
  MUX U3243 ( .IN0(reg_target[7]), .IN1(o[263]), .SEL(n2055), .F(
        \Data_Mem/n7480 ) );
  MUX U3244 ( .IN0(reg_target[6]), .IN1(o[262]), .SEL(n2055), .F(
        \Data_Mem/n7479 ) );
  MUX U3245 ( .IN0(reg_target[5]), .IN1(o[261]), .SEL(n2055), .F(
        \Data_Mem/n7478 ) );
  MUX U3246 ( .IN0(reg_target[4]), .IN1(o[260]), .SEL(n2055), .F(
        \Data_Mem/n7477 ) );
  MUX U3247 ( .IN0(reg_target[3]), .IN1(o[259]), .SEL(n2055), .F(
        \Data_Mem/n7476 ) );
  IV U3248 ( .A(n2056), .Z(n2055) );
  MUX U3249 ( .IN0(o[258]), .IN1(reg_target[2]), .SEL(n2056), .F(
        \Data_Mem/n7475 ) );
  MUX U3250 ( .IN0(o[257]), .IN1(reg_target[1]), .SEL(n2056), .F(
        \Data_Mem/n7474 ) );
  MUX U3251 ( .IN0(o[256]), .IN1(reg_target[0]), .SEL(n2056), .F(
        \Data_Mem/n7473 ) );
  NAND U3252 ( .A(n2053), .B(n2057), .Z(n2056) );
  NANDN U3253 ( .B(n2046), .A(n1899), .Z(n2057) );
  ANDN U3254 ( .A(n2058), .B(n2043), .Z(n2053) );
  ANDN U3255 ( .A(n1902), .B(n2046), .Z(n2043) );
  NANDN U3256 ( .B(n2046), .A(n1924), .Z(n2058) );
  NAND U3257 ( .A(n1903), .B(n2059), .Z(n2046) );
  MUX U3258 ( .IN0(n1853), .IN1(o[319]), .SEL(n2060), .F(\Data_Mem/n7472 ) );
  MUX U3259 ( .IN0(n1855), .IN1(o[318]), .SEL(n2060), .F(\Data_Mem/n7471 ) );
  MUX U3260 ( .IN0(n1856), .IN1(o[317]), .SEL(n2060), .F(\Data_Mem/n7470 ) );
  MUX U3261 ( .IN0(n1857), .IN1(o[316]), .SEL(n2060), .F(\Data_Mem/n7469 ) );
  MUX U3262 ( .IN0(n1858), .IN1(o[315]), .SEL(n2060), .F(\Data_Mem/n7468 ) );
  MUX U3263 ( .IN0(n1859), .IN1(o[314]), .SEL(n2060), .F(\Data_Mem/n7467 ) );
  MUX U3264 ( .IN0(n1860), .IN1(o[313]), .SEL(n2060), .F(\Data_Mem/n7466 ) );
  MUX U3265 ( .IN0(n1861), .IN1(o[312]), .SEL(n2060), .F(\Data_Mem/n7465 ) );
  ANDN U3266 ( .A(n2061), .B(n2062), .Z(n2060) );
  AND U3267 ( .A(n2063), .B(n2064), .Z(n2061) );
  OR U3268 ( .A(n1867), .B(n2065), .Z(n2064) );
  MUX U3269 ( .IN0(n1868), .IN1(o[311]), .SEL(n2066), .F(\Data_Mem/n7464 ) );
  MUX U3270 ( .IN0(n1870), .IN1(o[310]), .SEL(n2066), .F(\Data_Mem/n7463 ) );
  MUX U3271 ( .IN0(n1871), .IN1(o[309]), .SEL(n2066), .F(\Data_Mem/n7462 ) );
  MUX U3272 ( .IN0(n1872), .IN1(o[308]), .SEL(n2066), .F(\Data_Mem/n7461 ) );
  MUX U3273 ( .IN0(n1873), .IN1(o[307]), .SEL(n2066), .F(\Data_Mem/n7460 ) );
  IV U3274 ( .A(n2067), .Z(n2066) );
  MUX U3275 ( .IN0(o[306]), .IN1(n1875), .SEL(n2067), .F(\Data_Mem/n7459 ) );
  MUX U3276 ( .IN0(o[305]), .IN1(n1876), .SEL(n2067), .F(\Data_Mem/n7458 ) );
  MUX U3277 ( .IN0(o[304]), .IN1(n1877), .SEL(n2067), .F(\Data_Mem/n7457 ) );
  NAND U3278 ( .A(n2068), .B(n2069), .Z(n2067) );
  OR U3279 ( .A(n1880), .B(n2065), .Z(n2069) );
  ANDN U3280 ( .A(n2063), .B(n2062), .Z(n2068) );
  NANDN U3281 ( .B(n2065), .A(n1915), .Z(n2063) );
  MUX U3282 ( .IN0(n1883), .IN1(o[303]), .SEL(n2070), .F(\Data_Mem/n7456 ) );
  MUX U3283 ( .IN0(n1885), .IN1(o[302]), .SEL(n2070), .F(\Data_Mem/n7455 ) );
  MUX U3284 ( .IN0(n1886), .IN1(o[301]), .SEL(n2070), .F(\Data_Mem/n7454 ) );
  MUX U3285 ( .IN0(n1887), .IN1(o[300]), .SEL(n2070), .F(\Data_Mem/n7453 ) );
  MUX U3286 ( .IN0(n1888), .IN1(o[299]), .SEL(n2070), .F(\Data_Mem/n7452 ) );
  IV U3287 ( .A(n2071), .Z(n2070) );
  MUX U3288 ( .IN0(o[298]), .IN1(n1890), .SEL(n2071), .F(\Data_Mem/n7451 ) );
  MUX U3289 ( .IN0(o[297]), .IN1(n1891), .SEL(n2071), .F(\Data_Mem/n7450 ) );
  MUX U3290 ( .IN0(o[296]), .IN1(n1892), .SEL(n2071), .F(\Data_Mem/n7449 ) );
  NAND U3291 ( .A(n2072), .B(n2073), .Z(n2071) );
  OR U3292 ( .A(n1895), .B(n2065), .Z(n2073) );
  MUX U3293 ( .IN0(reg_target[7]), .IN1(o[295]), .SEL(n2074), .F(
        \Data_Mem/n7448 ) );
  MUX U3294 ( .IN0(reg_target[6]), .IN1(o[294]), .SEL(n2074), .F(
        \Data_Mem/n7447 ) );
  MUX U3295 ( .IN0(reg_target[5]), .IN1(o[293]), .SEL(n2074), .F(
        \Data_Mem/n7446 ) );
  MUX U3296 ( .IN0(reg_target[4]), .IN1(o[292]), .SEL(n2074), .F(
        \Data_Mem/n7445 ) );
  MUX U3297 ( .IN0(reg_target[3]), .IN1(o[291]), .SEL(n2074), .F(
        \Data_Mem/n7444 ) );
  IV U3298 ( .A(n2075), .Z(n2074) );
  MUX U3299 ( .IN0(o[290]), .IN1(reg_target[2]), .SEL(n2075), .F(
        \Data_Mem/n7443 ) );
  MUX U3300 ( .IN0(o[289]), .IN1(reg_target[1]), .SEL(n2075), .F(
        \Data_Mem/n7442 ) );
  MUX U3301 ( .IN0(o[288]), .IN1(reg_target[0]), .SEL(n2075), .F(
        \Data_Mem/n7441 ) );
  NAND U3302 ( .A(n2072), .B(n2076), .Z(n2075) );
  NANDN U3303 ( .B(n2065), .A(n1899), .Z(n2076) );
  ANDN U3304 ( .A(n2077), .B(n2062), .Z(n2072) );
  ANDN U3305 ( .A(n1902), .B(n2065), .Z(n2062) );
  NANDN U3306 ( .B(n2065), .A(n1924), .Z(n2077) );
  NAND U3307 ( .A(n1925), .B(n2059), .Z(n2065) );
  MUX U3308 ( .IN0(n1853), .IN1(o[351]), .SEL(n2078), .F(\Data_Mem/n7440 ) );
  MUX U3309 ( .IN0(n1855), .IN1(o[350]), .SEL(n2078), .F(\Data_Mem/n7439 ) );
  MUX U3310 ( .IN0(n1856), .IN1(o[349]), .SEL(n2078), .F(\Data_Mem/n7438 ) );
  MUX U3311 ( .IN0(n1857), .IN1(o[348]), .SEL(n2078), .F(\Data_Mem/n7437 ) );
  MUX U3312 ( .IN0(n1858), .IN1(o[347]), .SEL(n2078), .F(\Data_Mem/n7436 ) );
  MUX U3313 ( .IN0(n1859), .IN1(o[346]), .SEL(n2078), .F(\Data_Mem/n7435 ) );
  MUX U3314 ( .IN0(n1860), .IN1(o[345]), .SEL(n2078), .F(\Data_Mem/n7434 ) );
  MUX U3315 ( .IN0(n1861), .IN1(o[344]), .SEL(n2078), .F(\Data_Mem/n7433 ) );
  ANDN U3316 ( .A(n2079), .B(n2080), .Z(n2078) );
  AND U3317 ( .A(n2081), .B(n2082), .Z(n2079) );
  OR U3318 ( .A(n1867), .B(n2083), .Z(n2082) );
  MUX U3319 ( .IN0(n1868), .IN1(o[343]), .SEL(n2084), .F(\Data_Mem/n7432 ) );
  MUX U3320 ( .IN0(n1870), .IN1(o[342]), .SEL(n2084), .F(\Data_Mem/n7431 ) );
  MUX U3321 ( .IN0(n1871), .IN1(o[341]), .SEL(n2084), .F(\Data_Mem/n7430 ) );
  MUX U3322 ( .IN0(n1872), .IN1(o[340]), .SEL(n2084), .F(\Data_Mem/n7429 ) );
  MUX U3323 ( .IN0(n1873), .IN1(o[339]), .SEL(n2084), .F(\Data_Mem/n7428 ) );
  IV U3324 ( .A(n2085), .Z(n2084) );
  MUX U3325 ( .IN0(o[338]), .IN1(n1875), .SEL(n2085), .F(\Data_Mem/n7427 ) );
  MUX U3326 ( .IN0(o[337]), .IN1(n1876), .SEL(n2085), .F(\Data_Mem/n7426 ) );
  MUX U3327 ( .IN0(o[336]), .IN1(n1877), .SEL(n2085), .F(\Data_Mem/n7425 ) );
  NAND U3328 ( .A(n2086), .B(n2087), .Z(n2085) );
  OR U3329 ( .A(n1880), .B(n2083), .Z(n2087) );
  ANDN U3330 ( .A(n2081), .B(n2080), .Z(n2086) );
  NANDN U3331 ( .B(n2083), .A(n1915), .Z(n2081) );
  MUX U3332 ( .IN0(n1883), .IN1(o[335]), .SEL(n2088), .F(\Data_Mem/n7424 ) );
  MUX U3333 ( .IN0(n1885), .IN1(o[334]), .SEL(n2088), .F(\Data_Mem/n7423 ) );
  MUX U3334 ( .IN0(n1886), .IN1(o[333]), .SEL(n2088), .F(\Data_Mem/n7422 ) );
  MUX U3335 ( .IN0(n1887), .IN1(o[332]), .SEL(n2088), .F(\Data_Mem/n7421 ) );
  MUX U3336 ( .IN0(n1888), .IN1(o[331]), .SEL(n2088), .F(\Data_Mem/n7420 ) );
  IV U3337 ( .A(n2089), .Z(n2088) );
  MUX U3338 ( .IN0(o[330]), .IN1(n1890), .SEL(n2089), .F(\Data_Mem/n7419 ) );
  MUX U3339 ( .IN0(o[329]), .IN1(n1891), .SEL(n2089), .F(\Data_Mem/n7418 ) );
  MUX U3340 ( .IN0(o[328]), .IN1(n1892), .SEL(n2089), .F(\Data_Mem/n7417 ) );
  NAND U3341 ( .A(n2090), .B(n2091), .Z(n2089) );
  OR U3342 ( .A(n1895), .B(n2083), .Z(n2091) );
  MUX U3343 ( .IN0(reg_target[7]), .IN1(o[327]), .SEL(n2092), .F(
        \Data_Mem/n7416 ) );
  MUX U3344 ( .IN0(reg_target[6]), .IN1(o[326]), .SEL(n2092), .F(
        \Data_Mem/n7415 ) );
  MUX U3345 ( .IN0(reg_target[5]), .IN1(o[325]), .SEL(n2092), .F(
        \Data_Mem/n7414 ) );
  MUX U3346 ( .IN0(reg_target[4]), .IN1(o[324]), .SEL(n2092), .F(
        \Data_Mem/n7413 ) );
  MUX U3347 ( .IN0(reg_target[3]), .IN1(o[323]), .SEL(n2092), .F(
        \Data_Mem/n7412 ) );
  IV U3348 ( .A(n2093), .Z(n2092) );
  MUX U3349 ( .IN0(o[322]), .IN1(reg_target[2]), .SEL(n2093), .F(
        \Data_Mem/n7411 ) );
  MUX U3350 ( .IN0(o[321]), .IN1(reg_target[1]), .SEL(n2093), .F(
        \Data_Mem/n7410 ) );
  MUX U3351 ( .IN0(o[320]), .IN1(reg_target[0]), .SEL(n2093), .F(
        \Data_Mem/n7409 ) );
  NAND U3352 ( .A(n2090), .B(n2094), .Z(n2093) );
  NANDN U3353 ( .B(n2083), .A(n1899), .Z(n2094) );
  ANDN U3354 ( .A(n2095), .B(n2080), .Z(n2090) );
  ANDN U3355 ( .A(n1902), .B(n2083), .Z(n2080) );
  NANDN U3356 ( .B(n2083), .A(n1924), .Z(n2095) );
  NAND U3357 ( .A(n1944), .B(n2059), .Z(n2083) );
  MUX U3358 ( .IN0(n1853), .IN1(o[383]), .SEL(n2096), .F(\Data_Mem/n7408 ) );
  MUX U3359 ( .IN0(n1855), .IN1(o[382]), .SEL(n2096), .F(\Data_Mem/n7407 ) );
  MUX U3360 ( .IN0(n1856), .IN1(o[381]), .SEL(n2096), .F(\Data_Mem/n7406 ) );
  MUX U3361 ( .IN0(n1857), .IN1(o[380]), .SEL(n2096), .F(\Data_Mem/n7405 ) );
  MUX U3362 ( .IN0(n1858), .IN1(o[379]), .SEL(n2096), .F(\Data_Mem/n7404 ) );
  MUX U3363 ( .IN0(n1859), .IN1(o[378]), .SEL(n2096), .F(\Data_Mem/n7403 ) );
  MUX U3364 ( .IN0(n1860), .IN1(o[377]), .SEL(n2096), .F(\Data_Mem/n7402 ) );
  MUX U3365 ( .IN0(n1861), .IN1(o[376]), .SEL(n2096), .F(\Data_Mem/n7401 ) );
  ANDN U3366 ( .A(n2097), .B(n2098), .Z(n2096) );
  AND U3367 ( .A(n2099), .B(n2100), .Z(n2097) );
  OR U3368 ( .A(n1867), .B(n2101), .Z(n2100) );
  MUX U3369 ( .IN0(n1868), .IN1(o[375]), .SEL(n2102), .F(\Data_Mem/n7400 ) );
  MUX U3370 ( .IN0(n1870), .IN1(o[374]), .SEL(n2102), .F(\Data_Mem/n7399 ) );
  MUX U3371 ( .IN0(n1871), .IN1(o[373]), .SEL(n2102), .F(\Data_Mem/n7398 ) );
  MUX U3372 ( .IN0(n1872), .IN1(o[372]), .SEL(n2102), .F(\Data_Mem/n7397 ) );
  MUX U3373 ( .IN0(n1873), .IN1(o[371]), .SEL(n2102), .F(\Data_Mem/n7396 ) );
  IV U3374 ( .A(n2103), .Z(n2102) );
  MUX U3375 ( .IN0(o[370]), .IN1(n1875), .SEL(n2103), .F(\Data_Mem/n7395 ) );
  MUX U3376 ( .IN0(o[369]), .IN1(n1876), .SEL(n2103), .F(\Data_Mem/n7394 ) );
  MUX U3377 ( .IN0(o[368]), .IN1(n1877), .SEL(n2103), .F(\Data_Mem/n7393 ) );
  NAND U3378 ( .A(n2104), .B(n2105), .Z(n2103) );
  OR U3379 ( .A(n1880), .B(n2101), .Z(n2105) );
  ANDN U3380 ( .A(n2099), .B(n2098), .Z(n2104) );
  NANDN U3381 ( .B(n2101), .A(n1915), .Z(n2099) );
  MUX U3382 ( .IN0(n1883), .IN1(o[367]), .SEL(n2106), .F(\Data_Mem/n7392 ) );
  MUX U3383 ( .IN0(n1885), .IN1(o[366]), .SEL(n2106), .F(\Data_Mem/n7391 ) );
  MUX U3384 ( .IN0(n1886), .IN1(o[365]), .SEL(n2106), .F(\Data_Mem/n7390 ) );
  MUX U3385 ( .IN0(n1887), .IN1(o[364]), .SEL(n2106), .F(\Data_Mem/n7389 ) );
  MUX U3386 ( .IN0(n1888), .IN1(o[363]), .SEL(n2106), .F(\Data_Mem/n7388 ) );
  IV U3387 ( .A(n2107), .Z(n2106) );
  MUX U3388 ( .IN0(o[362]), .IN1(n1890), .SEL(n2107), .F(\Data_Mem/n7387 ) );
  MUX U3389 ( .IN0(o[361]), .IN1(n1891), .SEL(n2107), .F(\Data_Mem/n7386 ) );
  MUX U3390 ( .IN0(o[360]), .IN1(n1892), .SEL(n2107), .F(\Data_Mem/n7385 ) );
  NAND U3391 ( .A(n2108), .B(n2109), .Z(n2107) );
  OR U3392 ( .A(n1895), .B(n2101), .Z(n2109) );
  MUX U3393 ( .IN0(reg_target[7]), .IN1(o[359]), .SEL(n2110), .F(
        \Data_Mem/n7384 ) );
  MUX U3394 ( .IN0(reg_target[6]), .IN1(o[358]), .SEL(n2110), .F(
        \Data_Mem/n7383 ) );
  MUX U3395 ( .IN0(reg_target[5]), .IN1(o[357]), .SEL(n2110), .F(
        \Data_Mem/n7382 ) );
  MUX U3396 ( .IN0(reg_target[4]), .IN1(o[356]), .SEL(n2110), .F(
        \Data_Mem/n7381 ) );
  MUX U3397 ( .IN0(reg_target[3]), .IN1(o[355]), .SEL(n2110), .F(
        \Data_Mem/n7380 ) );
  IV U3398 ( .A(n2111), .Z(n2110) );
  MUX U3399 ( .IN0(o[354]), .IN1(reg_target[2]), .SEL(n2111), .F(
        \Data_Mem/n7379 ) );
  MUX U3400 ( .IN0(o[353]), .IN1(reg_target[1]), .SEL(n2111), .F(
        \Data_Mem/n7378 ) );
  MUX U3401 ( .IN0(o[352]), .IN1(reg_target[0]), .SEL(n2111), .F(
        \Data_Mem/n7377 ) );
  NAND U3402 ( .A(n2108), .B(n2112), .Z(n2111) );
  NANDN U3403 ( .B(n2101), .A(n1899), .Z(n2112) );
  ANDN U3404 ( .A(n2113), .B(n2098), .Z(n2108) );
  ANDN U3405 ( .A(n1902), .B(n2101), .Z(n2098) );
  NANDN U3406 ( .B(n2101), .A(n1924), .Z(n2113) );
  NAND U3407 ( .A(n1963), .B(n2059), .Z(n2101) );
  MUX U3408 ( .IN0(n1853), .IN1(o[415]), .SEL(n2114), .F(\Data_Mem/n7376 ) );
  MUX U3409 ( .IN0(n1855), .IN1(o[414]), .SEL(n2114), .F(\Data_Mem/n7375 ) );
  MUX U3410 ( .IN0(n1856), .IN1(o[413]), .SEL(n2114), .F(\Data_Mem/n7374 ) );
  MUX U3411 ( .IN0(n1857), .IN1(o[412]), .SEL(n2114), .F(\Data_Mem/n7373 ) );
  MUX U3412 ( .IN0(n1858), .IN1(o[411]), .SEL(n2114), .F(\Data_Mem/n7372 ) );
  MUX U3413 ( .IN0(n1859), .IN1(o[410]), .SEL(n2114), .F(\Data_Mem/n7371 ) );
  MUX U3414 ( .IN0(n1860), .IN1(o[409]), .SEL(n2114), .F(\Data_Mem/n7370 ) );
  MUX U3415 ( .IN0(n1861), .IN1(o[408]), .SEL(n2114), .F(\Data_Mem/n7369 ) );
  ANDN U3416 ( .A(n2115), .B(n2116), .Z(n2114) );
  AND U3417 ( .A(n2117), .B(n2118), .Z(n2115) );
  OR U3418 ( .A(n1867), .B(n2119), .Z(n2118) );
  MUX U3419 ( .IN0(n1868), .IN1(o[407]), .SEL(n2120), .F(\Data_Mem/n7368 ) );
  MUX U3420 ( .IN0(n1870), .IN1(o[406]), .SEL(n2120), .F(\Data_Mem/n7367 ) );
  MUX U3421 ( .IN0(n1871), .IN1(o[405]), .SEL(n2120), .F(\Data_Mem/n7366 ) );
  MUX U3422 ( .IN0(n1872), .IN1(o[404]), .SEL(n2120), .F(\Data_Mem/n7365 ) );
  MUX U3423 ( .IN0(n1873), .IN1(o[403]), .SEL(n2120), .F(\Data_Mem/n7364 ) );
  IV U3424 ( .A(n2121), .Z(n2120) );
  MUX U3425 ( .IN0(o[402]), .IN1(n1875), .SEL(n2121), .F(\Data_Mem/n7363 ) );
  MUX U3426 ( .IN0(o[401]), .IN1(n1876), .SEL(n2121), .F(\Data_Mem/n7362 ) );
  MUX U3427 ( .IN0(o[400]), .IN1(n1877), .SEL(n2121), .F(\Data_Mem/n7361 ) );
  NAND U3428 ( .A(n2122), .B(n2123), .Z(n2121) );
  OR U3429 ( .A(n1880), .B(n2119), .Z(n2123) );
  ANDN U3430 ( .A(n2117), .B(n2116), .Z(n2122) );
  NANDN U3431 ( .B(n2119), .A(n1915), .Z(n2117) );
  MUX U3432 ( .IN0(n1883), .IN1(o[399]), .SEL(n2124), .F(\Data_Mem/n7360 ) );
  MUX U3433 ( .IN0(n1885), .IN1(o[398]), .SEL(n2124), .F(\Data_Mem/n7359 ) );
  MUX U3434 ( .IN0(n1886), .IN1(o[397]), .SEL(n2124), .F(\Data_Mem/n7358 ) );
  MUX U3435 ( .IN0(n1887), .IN1(o[396]), .SEL(n2124), .F(\Data_Mem/n7357 ) );
  MUX U3436 ( .IN0(n1888), .IN1(o[395]), .SEL(n2124), .F(\Data_Mem/n7356 ) );
  IV U3437 ( .A(n2125), .Z(n2124) );
  MUX U3438 ( .IN0(o[394]), .IN1(n1890), .SEL(n2125), .F(\Data_Mem/n7355 ) );
  MUX U3439 ( .IN0(o[393]), .IN1(n1891), .SEL(n2125), .F(\Data_Mem/n7354 ) );
  MUX U3440 ( .IN0(o[392]), .IN1(n1892), .SEL(n2125), .F(\Data_Mem/n7353 ) );
  NAND U3441 ( .A(n2126), .B(n2127), .Z(n2125) );
  OR U3442 ( .A(n1895), .B(n2119), .Z(n2127) );
  MUX U3443 ( .IN0(reg_target[7]), .IN1(o[391]), .SEL(n2128), .F(
        \Data_Mem/n7352 ) );
  MUX U3444 ( .IN0(reg_target[6]), .IN1(o[390]), .SEL(n2128), .F(
        \Data_Mem/n7351 ) );
  MUX U3445 ( .IN0(reg_target[5]), .IN1(o[389]), .SEL(n2128), .F(
        \Data_Mem/n7350 ) );
  MUX U3446 ( .IN0(reg_target[4]), .IN1(o[388]), .SEL(n2128), .F(
        \Data_Mem/n7349 ) );
  MUX U3447 ( .IN0(reg_target[3]), .IN1(o[387]), .SEL(n2128), .F(
        \Data_Mem/n7348 ) );
  IV U3448 ( .A(n2129), .Z(n2128) );
  MUX U3449 ( .IN0(o[386]), .IN1(reg_target[2]), .SEL(n2129), .F(
        \Data_Mem/n7347 ) );
  MUX U3450 ( .IN0(o[385]), .IN1(reg_target[1]), .SEL(n2129), .F(
        \Data_Mem/n7346 ) );
  MUX U3451 ( .IN0(o[384]), .IN1(reg_target[0]), .SEL(n2129), .F(
        \Data_Mem/n7345 ) );
  NAND U3452 ( .A(n2126), .B(n2130), .Z(n2129) );
  NANDN U3453 ( .B(n2119), .A(n1899), .Z(n2130) );
  ANDN U3454 ( .A(n2131), .B(n2116), .Z(n2126) );
  ANDN U3455 ( .A(n1902), .B(n2119), .Z(n2116) );
  NANDN U3456 ( .B(n2119), .A(n1924), .Z(n2131) );
  NAND U3457 ( .A(n1982), .B(n2059), .Z(n2119) );
  MUX U3458 ( .IN0(n1853), .IN1(o[447]), .SEL(n2132), .F(\Data_Mem/n7344 ) );
  MUX U3459 ( .IN0(n1855), .IN1(o[446]), .SEL(n2132), .F(\Data_Mem/n7343 ) );
  MUX U3460 ( .IN0(n1856), .IN1(o[445]), .SEL(n2132), .F(\Data_Mem/n7342 ) );
  MUX U3461 ( .IN0(n1857), .IN1(o[444]), .SEL(n2132), .F(\Data_Mem/n7341 ) );
  MUX U3462 ( .IN0(n1858), .IN1(o[443]), .SEL(n2132), .F(\Data_Mem/n7340 ) );
  MUX U3463 ( .IN0(n1859), .IN1(o[442]), .SEL(n2132), .F(\Data_Mem/n7339 ) );
  MUX U3464 ( .IN0(n1860), .IN1(o[441]), .SEL(n2132), .F(\Data_Mem/n7338 ) );
  MUX U3465 ( .IN0(n1861), .IN1(o[440]), .SEL(n2132), .F(\Data_Mem/n7337 ) );
  ANDN U3466 ( .A(n2133), .B(n2134), .Z(n2132) );
  AND U3467 ( .A(n2135), .B(n2136), .Z(n2133) );
  OR U3468 ( .A(n1867), .B(n2137), .Z(n2136) );
  MUX U3469 ( .IN0(n1868), .IN1(o[439]), .SEL(n2138), .F(\Data_Mem/n7336 ) );
  MUX U3470 ( .IN0(n1870), .IN1(o[438]), .SEL(n2138), .F(\Data_Mem/n7335 ) );
  MUX U3471 ( .IN0(n1871), .IN1(o[437]), .SEL(n2138), .F(\Data_Mem/n7334 ) );
  MUX U3472 ( .IN0(n1872), .IN1(o[436]), .SEL(n2138), .F(\Data_Mem/n7333 ) );
  MUX U3473 ( .IN0(n1873), .IN1(o[435]), .SEL(n2138), .F(\Data_Mem/n7332 ) );
  IV U3474 ( .A(n2139), .Z(n2138) );
  MUX U3475 ( .IN0(o[434]), .IN1(n1875), .SEL(n2139), .F(\Data_Mem/n7331 ) );
  MUX U3476 ( .IN0(o[433]), .IN1(n1876), .SEL(n2139), .F(\Data_Mem/n7330 ) );
  MUX U3477 ( .IN0(o[432]), .IN1(n1877), .SEL(n2139), .F(\Data_Mem/n7329 ) );
  NAND U3478 ( .A(n2140), .B(n2141), .Z(n2139) );
  OR U3479 ( .A(n1880), .B(n2137), .Z(n2141) );
  ANDN U3480 ( .A(n2135), .B(n2134), .Z(n2140) );
  NANDN U3481 ( .B(n2137), .A(n1915), .Z(n2135) );
  MUX U3482 ( .IN0(n1883), .IN1(o[431]), .SEL(n2142), .F(\Data_Mem/n7328 ) );
  MUX U3483 ( .IN0(n1885), .IN1(o[430]), .SEL(n2142), .F(\Data_Mem/n7327 ) );
  MUX U3484 ( .IN0(n1886), .IN1(o[429]), .SEL(n2142), .F(\Data_Mem/n7326 ) );
  MUX U3485 ( .IN0(n1887), .IN1(o[428]), .SEL(n2142), .F(\Data_Mem/n7325 ) );
  MUX U3486 ( .IN0(n1888), .IN1(o[427]), .SEL(n2142), .F(\Data_Mem/n7324 ) );
  IV U3487 ( .A(n2143), .Z(n2142) );
  MUX U3488 ( .IN0(o[426]), .IN1(n1890), .SEL(n2143), .F(\Data_Mem/n7323 ) );
  MUX U3489 ( .IN0(o[425]), .IN1(n1891), .SEL(n2143), .F(\Data_Mem/n7322 ) );
  MUX U3490 ( .IN0(o[424]), .IN1(n1892), .SEL(n2143), .F(\Data_Mem/n7321 ) );
  NAND U3491 ( .A(n2144), .B(n2145), .Z(n2143) );
  OR U3492 ( .A(n1895), .B(n2137), .Z(n2145) );
  MUX U3493 ( .IN0(reg_target[7]), .IN1(o[423]), .SEL(n2146), .F(
        \Data_Mem/n7320 ) );
  MUX U3494 ( .IN0(reg_target[6]), .IN1(o[422]), .SEL(n2146), .F(
        \Data_Mem/n7319 ) );
  MUX U3495 ( .IN0(reg_target[5]), .IN1(o[421]), .SEL(n2146), .F(
        \Data_Mem/n7318 ) );
  MUX U3496 ( .IN0(reg_target[4]), .IN1(o[420]), .SEL(n2146), .F(
        \Data_Mem/n7317 ) );
  MUX U3497 ( .IN0(reg_target[3]), .IN1(o[419]), .SEL(n2146), .F(
        \Data_Mem/n7316 ) );
  IV U3498 ( .A(n2147), .Z(n2146) );
  MUX U3499 ( .IN0(o[418]), .IN1(reg_target[2]), .SEL(n2147), .F(
        \Data_Mem/n7315 ) );
  MUX U3500 ( .IN0(o[417]), .IN1(reg_target[1]), .SEL(n2147), .F(
        \Data_Mem/n7314 ) );
  MUX U3501 ( .IN0(o[416]), .IN1(reg_target[0]), .SEL(n2147), .F(
        \Data_Mem/n7313 ) );
  NAND U3502 ( .A(n2144), .B(n2148), .Z(n2147) );
  NANDN U3503 ( .B(n2137), .A(n1899), .Z(n2148) );
  ANDN U3504 ( .A(n2149), .B(n2134), .Z(n2144) );
  ANDN U3505 ( .A(n1902), .B(n2137), .Z(n2134) );
  NANDN U3506 ( .B(n2137), .A(n1924), .Z(n2149) );
  NAND U3507 ( .A(n2001), .B(n2059), .Z(n2137) );
  MUX U3508 ( .IN0(n1853), .IN1(o[479]), .SEL(n2150), .F(\Data_Mem/n7312 ) );
  MUX U3509 ( .IN0(n1855), .IN1(o[478]), .SEL(n2150), .F(\Data_Mem/n7311 ) );
  MUX U3510 ( .IN0(n1856), .IN1(o[477]), .SEL(n2150), .F(\Data_Mem/n7310 ) );
  MUX U3511 ( .IN0(n1857), .IN1(o[476]), .SEL(n2150), .F(\Data_Mem/n7309 ) );
  MUX U3512 ( .IN0(n1858), .IN1(o[475]), .SEL(n2150), .F(\Data_Mem/n7308 ) );
  MUX U3513 ( .IN0(n1859), .IN1(o[474]), .SEL(n2150), .F(\Data_Mem/n7307 ) );
  MUX U3514 ( .IN0(n1860), .IN1(o[473]), .SEL(n2150), .F(\Data_Mem/n7306 ) );
  MUX U3515 ( .IN0(n1861), .IN1(o[472]), .SEL(n2150), .F(\Data_Mem/n7305 ) );
  ANDN U3516 ( .A(n2151), .B(n2152), .Z(n2150) );
  AND U3517 ( .A(n2153), .B(n2154), .Z(n2151) );
  OR U3518 ( .A(n1867), .B(n2155), .Z(n2154) );
  MUX U3519 ( .IN0(n1868), .IN1(o[471]), .SEL(n2156), .F(\Data_Mem/n7304 ) );
  MUX U3520 ( .IN0(n1870), .IN1(o[470]), .SEL(n2156), .F(\Data_Mem/n7303 ) );
  MUX U3521 ( .IN0(n1871), .IN1(o[469]), .SEL(n2156), .F(\Data_Mem/n7302 ) );
  MUX U3522 ( .IN0(n1872), .IN1(o[468]), .SEL(n2156), .F(\Data_Mem/n7301 ) );
  MUX U3523 ( .IN0(n1873), .IN1(o[467]), .SEL(n2156), .F(\Data_Mem/n7300 ) );
  IV U3524 ( .A(n2157), .Z(n2156) );
  MUX U3525 ( .IN0(o[466]), .IN1(n1875), .SEL(n2157), .F(\Data_Mem/n7299 ) );
  MUX U3526 ( .IN0(o[465]), .IN1(n1876), .SEL(n2157), .F(\Data_Mem/n7298 ) );
  MUX U3527 ( .IN0(o[464]), .IN1(n1877), .SEL(n2157), .F(\Data_Mem/n7297 ) );
  NAND U3528 ( .A(n2158), .B(n2159), .Z(n2157) );
  OR U3529 ( .A(n1880), .B(n2155), .Z(n2159) );
  ANDN U3530 ( .A(n2153), .B(n2152), .Z(n2158) );
  NANDN U3531 ( .B(n2155), .A(n1915), .Z(n2153) );
  MUX U3532 ( .IN0(n1883), .IN1(o[463]), .SEL(n2160), .F(\Data_Mem/n7296 ) );
  MUX U3533 ( .IN0(n1885), .IN1(o[462]), .SEL(n2160), .F(\Data_Mem/n7295 ) );
  MUX U3534 ( .IN0(n1886), .IN1(o[461]), .SEL(n2160), .F(\Data_Mem/n7294 ) );
  MUX U3535 ( .IN0(n1887), .IN1(o[460]), .SEL(n2160), .F(\Data_Mem/n7293 ) );
  MUX U3536 ( .IN0(n1888), .IN1(o[459]), .SEL(n2160), .F(\Data_Mem/n7292 ) );
  IV U3537 ( .A(n2161), .Z(n2160) );
  MUX U3538 ( .IN0(o[458]), .IN1(n1890), .SEL(n2161), .F(\Data_Mem/n7291 ) );
  MUX U3539 ( .IN0(o[457]), .IN1(n1891), .SEL(n2161), .F(\Data_Mem/n7290 ) );
  MUX U3540 ( .IN0(o[456]), .IN1(n1892), .SEL(n2161), .F(\Data_Mem/n7289 ) );
  NAND U3541 ( .A(n2162), .B(n2163), .Z(n2161) );
  OR U3542 ( .A(n1895), .B(n2155), .Z(n2163) );
  MUX U3543 ( .IN0(reg_target[7]), .IN1(o[455]), .SEL(n2164), .F(
        \Data_Mem/n7288 ) );
  MUX U3544 ( .IN0(reg_target[6]), .IN1(o[454]), .SEL(n2164), .F(
        \Data_Mem/n7287 ) );
  MUX U3545 ( .IN0(reg_target[5]), .IN1(o[453]), .SEL(n2164), .F(
        \Data_Mem/n7286 ) );
  MUX U3546 ( .IN0(reg_target[4]), .IN1(o[452]), .SEL(n2164), .F(
        \Data_Mem/n7285 ) );
  MUX U3547 ( .IN0(reg_target[3]), .IN1(o[451]), .SEL(n2164), .F(
        \Data_Mem/n7284 ) );
  IV U3548 ( .A(n2165), .Z(n2164) );
  MUX U3549 ( .IN0(o[450]), .IN1(reg_target[2]), .SEL(n2165), .F(
        \Data_Mem/n7283 ) );
  MUX U3550 ( .IN0(o[449]), .IN1(reg_target[1]), .SEL(n2165), .F(
        \Data_Mem/n7282 ) );
  MUX U3551 ( .IN0(o[448]), .IN1(reg_target[0]), .SEL(n2165), .F(
        \Data_Mem/n7281 ) );
  NAND U3552 ( .A(n2162), .B(n2166), .Z(n2165) );
  NANDN U3553 ( .B(n2155), .A(n1899), .Z(n2166) );
  ANDN U3554 ( .A(n2167), .B(n2152), .Z(n2162) );
  ANDN U3555 ( .A(n1902), .B(n2155), .Z(n2152) );
  NANDN U3556 ( .B(n2155), .A(n1924), .Z(n2167) );
  NAND U3557 ( .A(n2020), .B(n2059), .Z(n2155) );
  MUX U3558 ( .IN0(n1853), .IN1(o[511]), .SEL(n2168), .F(\Data_Mem/n7280 ) );
  MUX U3559 ( .IN0(n1855), .IN1(o[510]), .SEL(n2168), .F(\Data_Mem/n7279 ) );
  MUX U3560 ( .IN0(n1856), .IN1(o[509]), .SEL(n2168), .F(\Data_Mem/n7278 ) );
  MUX U3561 ( .IN0(n1857), .IN1(o[508]), .SEL(n2168), .F(\Data_Mem/n7277 ) );
  MUX U3562 ( .IN0(n1858), .IN1(o[507]), .SEL(n2168), .F(\Data_Mem/n7276 ) );
  MUX U3563 ( .IN0(n1859), .IN1(o[506]), .SEL(n2168), .F(\Data_Mem/n7275 ) );
  MUX U3564 ( .IN0(n1860), .IN1(o[505]), .SEL(n2168), .F(\Data_Mem/n7274 ) );
  MUX U3565 ( .IN0(n1861), .IN1(o[504]), .SEL(n2168), .F(\Data_Mem/n7273 ) );
  ANDN U3566 ( .A(n2169), .B(n2170), .Z(n2168) );
  AND U3567 ( .A(n2171), .B(n2172), .Z(n2169) );
  OR U3568 ( .A(n1867), .B(n2173), .Z(n2172) );
  MUX U3569 ( .IN0(n1868), .IN1(o[503]), .SEL(n2174), .F(\Data_Mem/n7272 ) );
  MUX U3570 ( .IN0(n1870), .IN1(o[502]), .SEL(n2174), .F(\Data_Mem/n7271 ) );
  MUX U3571 ( .IN0(n1871), .IN1(o[501]), .SEL(n2174), .F(\Data_Mem/n7270 ) );
  MUX U3572 ( .IN0(n1872), .IN1(o[500]), .SEL(n2174), .F(\Data_Mem/n7269 ) );
  MUX U3573 ( .IN0(n1873), .IN1(o[499]), .SEL(n2174), .F(\Data_Mem/n7268 ) );
  IV U3574 ( .A(n2175), .Z(n2174) );
  MUX U3575 ( .IN0(o[498]), .IN1(n1875), .SEL(n2175), .F(\Data_Mem/n7267 ) );
  MUX U3576 ( .IN0(o[497]), .IN1(n1876), .SEL(n2175), .F(\Data_Mem/n7266 ) );
  MUX U3577 ( .IN0(o[496]), .IN1(n1877), .SEL(n2175), .F(\Data_Mem/n7265 ) );
  NAND U3578 ( .A(n2176), .B(n2177), .Z(n2175) );
  OR U3579 ( .A(n1880), .B(n2173), .Z(n2177) );
  ANDN U3580 ( .A(n2171), .B(n2170), .Z(n2176) );
  NANDN U3581 ( .B(n2173), .A(n1915), .Z(n2171) );
  MUX U3582 ( .IN0(n1883), .IN1(o[495]), .SEL(n2178), .F(\Data_Mem/n7264 ) );
  MUX U3583 ( .IN0(n1885), .IN1(o[494]), .SEL(n2178), .F(\Data_Mem/n7263 ) );
  MUX U3584 ( .IN0(n1886), .IN1(o[493]), .SEL(n2178), .F(\Data_Mem/n7262 ) );
  MUX U3585 ( .IN0(n1887), .IN1(o[492]), .SEL(n2178), .F(\Data_Mem/n7261 ) );
  MUX U3586 ( .IN0(n1888), .IN1(o[491]), .SEL(n2178), .F(\Data_Mem/n7260 ) );
  IV U3587 ( .A(n2179), .Z(n2178) );
  MUX U3588 ( .IN0(o[490]), .IN1(n1890), .SEL(n2179), .F(\Data_Mem/n7259 ) );
  MUX U3589 ( .IN0(o[489]), .IN1(n1891), .SEL(n2179), .F(\Data_Mem/n7258 ) );
  MUX U3590 ( .IN0(o[488]), .IN1(n1892), .SEL(n2179), .F(\Data_Mem/n7257 ) );
  NAND U3591 ( .A(n2180), .B(n2181), .Z(n2179) );
  OR U3592 ( .A(n1895), .B(n2173), .Z(n2181) );
  MUX U3593 ( .IN0(reg_target[7]), .IN1(o[487]), .SEL(n2182), .F(
        \Data_Mem/n7256 ) );
  MUX U3594 ( .IN0(reg_target[6]), .IN1(o[486]), .SEL(n2182), .F(
        \Data_Mem/n7255 ) );
  MUX U3595 ( .IN0(reg_target[5]), .IN1(o[485]), .SEL(n2182), .F(
        \Data_Mem/n7254 ) );
  MUX U3596 ( .IN0(reg_target[4]), .IN1(o[484]), .SEL(n2182), .F(
        \Data_Mem/n7253 ) );
  MUX U3597 ( .IN0(reg_target[3]), .IN1(o[483]), .SEL(n2182), .F(
        \Data_Mem/n7252 ) );
  IV U3598 ( .A(n2183), .Z(n2182) );
  MUX U3599 ( .IN0(o[482]), .IN1(reg_target[2]), .SEL(n2183), .F(
        \Data_Mem/n7251 ) );
  MUX U3600 ( .IN0(o[481]), .IN1(reg_target[1]), .SEL(n2183), .F(
        \Data_Mem/n7250 ) );
  MUX U3601 ( .IN0(o[480]), .IN1(reg_target[0]), .SEL(n2183), .F(
        \Data_Mem/n7249 ) );
  NAND U3602 ( .A(n2180), .B(n2184), .Z(n2183) );
  NANDN U3603 ( .B(n2173), .A(n1899), .Z(n2184) );
  ANDN U3604 ( .A(n2185), .B(n2170), .Z(n2180) );
  ANDN U3605 ( .A(n1902), .B(n2173), .Z(n2170) );
  NANDN U3606 ( .B(n2173), .A(n1924), .Z(n2185) );
  NAND U3607 ( .A(n2059), .B(n2039), .Z(n2173) );
  AND U3608 ( .A(n2186), .B(n485), .Z(n2059) );
  MUX U3609 ( .IN0(n1853), .IN1(o[543]), .SEL(n2187), .F(\Data_Mem/n7248 ) );
  MUX U3610 ( .IN0(n1855), .IN1(o[542]), .SEL(n2187), .F(\Data_Mem/n7247 ) );
  MUX U3611 ( .IN0(n1856), .IN1(o[541]), .SEL(n2187), .F(\Data_Mem/n7246 ) );
  MUX U3612 ( .IN0(n1857), .IN1(o[540]), .SEL(n2187), .F(\Data_Mem/n7245 ) );
  MUX U3613 ( .IN0(n1858), .IN1(o[539]), .SEL(n2187), .F(\Data_Mem/n7244 ) );
  MUX U3614 ( .IN0(n1859), .IN1(o[538]), .SEL(n2187), .F(\Data_Mem/n7243 ) );
  MUX U3615 ( .IN0(n1860), .IN1(o[537]), .SEL(n2187), .F(\Data_Mem/n7242 ) );
  MUX U3616 ( .IN0(n1861), .IN1(o[536]), .SEL(n2187), .F(\Data_Mem/n7241 ) );
  ANDN U3617 ( .A(n2188), .B(n2189), .Z(n2187) );
  AND U3618 ( .A(n2190), .B(n2191), .Z(n2188) );
  OR U3619 ( .A(n1867), .B(n2192), .Z(n2191) );
  MUX U3620 ( .IN0(n1868), .IN1(o[535]), .SEL(n2193), .F(\Data_Mem/n7240 ) );
  MUX U3621 ( .IN0(n1870), .IN1(o[534]), .SEL(n2193), .F(\Data_Mem/n7239 ) );
  MUX U3622 ( .IN0(n1871), .IN1(o[533]), .SEL(n2193), .F(\Data_Mem/n7238 ) );
  MUX U3623 ( .IN0(n1872), .IN1(o[532]), .SEL(n2193), .F(\Data_Mem/n7237 ) );
  MUX U3624 ( .IN0(n1873), .IN1(o[531]), .SEL(n2193), .F(\Data_Mem/n7236 ) );
  IV U3625 ( .A(n2194), .Z(n2193) );
  MUX U3626 ( .IN0(o[530]), .IN1(n1875), .SEL(n2194), .F(\Data_Mem/n7235 ) );
  MUX U3627 ( .IN0(o[529]), .IN1(n1876), .SEL(n2194), .F(\Data_Mem/n7234 ) );
  MUX U3628 ( .IN0(o[528]), .IN1(n1877), .SEL(n2194), .F(\Data_Mem/n7233 ) );
  NAND U3629 ( .A(n2195), .B(n2196), .Z(n2194) );
  OR U3630 ( .A(n1880), .B(n2192), .Z(n2196) );
  ANDN U3631 ( .A(n2190), .B(n2189), .Z(n2195) );
  NANDN U3632 ( .B(n2192), .A(n1915), .Z(n2190) );
  MUX U3633 ( .IN0(n1883), .IN1(o[527]), .SEL(n2197), .F(\Data_Mem/n7232 ) );
  MUX U3634 ( .IN0(n1885), .IN1(o[526]), .SEL(n2197), .F(\Data_Mem/n7231 ) );
  MUX U3635 ( .IN0(n1886), .IN1(o[525]), .SEL(n2197), .F(\Data_Mem/n7230 ) );
  MUX U3636 ( .IN0(n1887), .IN1(o[524]), .SEL(n2197), .F(\Data_Mem/n7229 ) );
  MUX U3637 ( .IN0(n1888), .IN1(o[523]), .SEL(n2197), .F(\Data_Mem/n7228 ) );
  IV U3638 ( .A(n2198), .Z(n2197) );
  MUX U3639 ( .IN0(o[522]), .IN1(n1890), .SEL(n2198), .F(\Data_Mem/n7227 ) );
  MUX U3640 ( .IN0(o[521]), .IN1(n1891), .SEL(n2198), .F(\Data_Mem/n7226 ) );
  MUX U3641 ( .IN0(o[520]), .IN1(n1892), .SEL(n2198), .F(\Data_Mem/n7225 ) );
  NAND U3642 ( .A(n2199), .B(n2200), .Z(n2198) );
  OR U3643 ( .A(n1895), .B(n2192), .Z(n2200) );
  MUX U3644 ( .IN0(reg_target[7]), .IN1(o[519]), .SEL(n2201), .F(
        \Data_Mem/n7224 ) );
  MUX U3645 ( .IN0(reg_target[6]), .IN1(o[518]), .SEL(n2201), .F(
        \Data_Mem/n7223 ) );
  MUX U3646 ( .IN0(reg_target[5]), .IN1(o[517]), .SEL(n2201), .F(
        \Data_Mem/n7222 ) );
  MUX U3647 ( .IN0(reg_target[4]), .IN1(o[516]), .SEL(n2201), .F(
        \Data_Mem/n7221 ) );
  MUX U3648 ( .IN0(reg_target[3]), .IN1(o[515]), .SEL(n2201), .F(
        \Data_Mem/n7220 ) );
  IV U3649 ( .A(n2202), .Z(n2201) );
  MUX U3650 ( .IN0(o[514]), .IN1(reg_target[2]), .SEL(n2202), .F(
        \Data_Mem/n7219 ) );
  MUX U3651 ( .IN0(o[513]), .IN1(reg_target[1]), .SEL(n2202), .F(
        \Data_Mem/n7218 ) );
  MUX U3652 ( .IN0(o[512]), .IN1(reg_target[0]), .SEL(n2202), .F(
        \Data_Mem/n7217 ) );
  NAND U3653 ( .A(n2199), .B(n2203), .Z(n2202) );
  NANDN U3654 ( .B(n2192), .A(n1899), .Z(n2203) );
  ANDN U3655 ( .A(n2204), .B(n2189), .Z(n2199) );
  ANDN U3656 ( .A(n1902), .B(n2192), .Z(n2189) );
  NANDN U3657 ( .B(n2192), .A(n1924), .Z(n2204) );
  NAND U3658 ( .A(n1903), .B(n2205), .Z(n2192) );
  MUX U3659 ( .IN0(n1853), .IN1(o[575]), .SEL(n2206), .F(\Data_Mem/n7216 ) );
  MUX U3660 ( .IN0(n1855), .IN1(o[574]), .SEL(n2206), .F(\Data_Mem/n7215 ) );
  MUX U3661 ( .IN0(n1856), .IN1(o[573]), .SEL(n2206), .F(\Data_Mem/n7214 ) );
  MUX U3662 ( .IN0(n1857), .IN1(o[572]), .SEL(n2206), .F(\Data_Mem/n7213 ) );
  MUX U3663 ( .IN0(n1858), .IN1(o[571]), .SEL(n2206), .F(\Data_Mem/n7212 ) );
  MUX U3664 ( .IN0(n1859), .IN1(o[570]), .SEL(n2206), .F(\Data_Mem/n7211 ) );
  MUX U3665 ( .IN0(n1860), .IN1(o[569]), .SEL(n2206), .F(\Data_Mem/n7210 ) );
  MUX U3666 ( .IN0(n1861), .IN1(o[568]), .SEL(n2206), .F(\Data_Mem/n7209 ) );
  ANDN U3667 ( .A(n2207), .B(n2208), .Z(n2206) );
  AND U3668 ( .A(n2209), .B(n2210), .Z(n2207) );
  OR U3669 ( .A(n1867), .B(n2211), .Z(n2210) );
  MUX U3670 ( .IN0(n1868), .IN1(o[567]), .SEL(n2212), .F(\Data_Mem/n7208 ) );
  MUX U3671 ( .IN0(n1870), .IN1(o[566]), .SEL(n2212), .F(\Data_Mem/n7207 ) );
  MUX U3672 ( .IN0(n1871), .IN1(o[565]), .SEL(n2212), .F(\Data_Mem/n7206 ) );
  MUX U3673 ( .IN0(n1872), .IN1(o[564]), .SEL(n2212), .F(\Data_Mem/n7205 ) );
  MUX U3674 ( .IN0(n1873), .IN1(o[563]), .SEL(n2212), .F(\Data_Mem/n7204 ) );
  IV U3675 ( .A(n2213), .Z(n2212) );
  MUX U3676 ( .IN0(o[562]), .IN1(n1875), .SEL(n2213), .F(\Data_Mem/n7203 ) );
  MUX U3677 ( .IN0(o[561]), .IN1(n1876), .SEL(n2213), .F(\Data_Mem/n7202 ) );
  MUX U3678 ( .IN0(o[560]), .IN1(n1877), .SEL(n2213), .F(\Data_Mem/n7201 ) );
  NAND U3679 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U3680 ( .A(n1880), .B(n2211), .Z(n2215) );
  ANDN U3681 ( .A(n2209), .B(n2208), .Z(n2214) );
  NANDN U3682 ( .B(n2211), .A(n1915), .Z(n2209) );
  MUX U3683 ( .IN0(n1883), .IN1(o[559]), .SEL(n2216), .F(\Data_Mem/n7200 ) );
  MUX U3684 ( .IN0(n1885), .IN1(o[558]), .SEL(n2216), .F(\Data_Mem/n7199 ) );
  MUX U3685 ( .IN0(n1886), .IN1(o[557]), .SEL(n2216), .F(\Data_Mem/n7198 ) );
  MUX U3686 ( .IN0(n1887), .IN1(o[556]), .SEL(n2216), .F(\Data_Mem/n7197 ) );
  MUX U3687 ( .IN0(n1888), .IN1(o[555]), .SEL(n2216), .F(\Data_Mem/n7196 ) );
  IV U3688 ( .A(n2217), .Z(n2216) );
  MUX U3689 ( .IN0(o[554]), .IN1(n1890), .SEL(n2217), .F(\Data_Mem/n7195 ) );
  MUX U3690 ( .IN0(o[553]), .IN1(n1891), .SEL(n2217), .F(\Data_Mem/n7194 ) );
  MUX U3691 ( .IN0(o[552]), .IN1(n1892), .SEL(n2217), .F(\Data_Mem/n7193 ) );
  NAND U3692 ( .A(n2218), .B(n2219), .Z(n2217) );
  OR U3693 ( .A(n1895), .B(n2211), .Z(n2219) );
  MUX U3694 ( .IN0(reg_target[7]), .IN1(o[551]), .SEL(n2220), .F(
        \Data_Mem/n7192 ) );
  MUX U3695 ( .IN0(reg_target[6]), .IN1(o[550]), .SEL(n2220), .F(
        \Data_Mem/n7191 ) );
  MUX U3696 ( .IN0(reg_target[5]), .IN1(o[549]), .SEL(n2220), .F(
        \Data_Mem/n7190 ) );
  MUX U3697 ( .IN0(reg_target[4]), .IN1(o[548]), .SEL(n2220), .F(
        \Data_Mem/n7189 ) );
  MUX U3698 ( .IN0(reg_target[3]), .IN1(o[547]), .SEL(n2220), .F(
        \Data_Mem/n7188 ) );
  IV U3699 ( .A(n2221), .Z(n2220) );
  MUX U3700 ( .IN0(o[546]), .IN1(reg_target[2]), .SEL(n2221), .F(
        \Data_Mem/n7187 ) );
  MUX U3701 ( .IN0(o[545]), .IN1(reg_target[1]), .SEL(n2221), .F(
        \Data_Mem/n7186 ) );
  MUX U3702 ( .IN0(o[544]), .IN1(reg_target[0]), .SEL(n2221), .F(
        \Data_Mem/n7185 ) );
  NAND U3703 ( .A(n2218), .B(n2222), .Z(n2221) );
  NANDN U3704 ( .B(n2211), .A(n1899), .Z(n2222) );
  ANDN U3705 ( .A(n2223), .B(n2208), .Z(n2218) );
  ANDN U3706 ( .A(n1902), .B(n2211), .Z(n2208) );
  NANDN U3707 ( .B(n2211), .A(n1924), .Z(n2223) );
  NAND U3708 ( .A(n1925), .B(n2205), .Z(n2211) );
  MUX U3709 ( .IN0(n1853), .IN1(o[607]), .SEL(n2224), .F(\Data_Mem/n7184 ) );
  MUX U3710 ( .IN0(n1855), .IN1(o[606]), .SEL(n2224), .F(\Data_Mem/n7183 ) );
  MUX U3711 ( .IN0(n1856), .IN1(o[605]), .SEL(n2224), .F(\Data_Mem/n7182 ) );
  MUX U3712 ( .IN0(n1857), .IN1(o[604]), .SEL(n2224), .F(\Data_Mem/n7181 ) );
  MUX U3713 ( .IN0(n1858), .IN1(o[603]), .SEL(n2224), .F(\Data_Mem/n7180 ) );
  MUX U3714 ( .IN0(n1859), .IN1(o[602]), .SEL(n2224), .F(\Data_Mem/n7179 ) );
  MUX U3715 ( .IN0(n1860), .IN1(o[601]), .SEL(n2224), .F(\Data_Mem/n7178 ) );
  MUX U3716 ( .IN0(n1861), .IN1(o[600]), .SEL(n2224), .F(\Data_Mem/n7177 ) );
  ANDN U3717 ( .A(n2225), .B(n2226), .Z(n2224) );
  AND U3718 ( .A(n2227), .B(n2228), .Z(n2225) );
  OR U3719 ( .A(n1867), .B(n2229), .Z(n2228) );
  MUX U3720 ( .IN0(n1868), .IN1(o[599]), .SEL(n2230), .F(\Data_Mem/n7176 ) );
  MUX U3721 ( .IN0(n1870), .IN1(o[598]), .SEL(n2230), .F(\Data_Mem/n7175 ) );
  MUX U3722 ( .IN0(n1871), .IN1(o[597]), .SEL(n2230), .F(\Data_Mem/n7174 ) );
  MUX U3723 ( .IN0(n1872), .IN1(o[596]), .SEL(n2230), .F(\Data_Mem/n7173 ) );
  MUX U3724 ( .IN0(n1873), .IN1(o[595]), .SEL(n2230), .F(\Data_Mem/n7172 ) );
  IV U3725 ( .A(n2231), .Z(n2230) );
  MUX U3726 ( .IN0(o[594]), .IN1(n1875), .SEL(n2231), .F(\Data_Mem/n7171 ) );
  MUX U3727 ( .IN0(o[593]), .IN1(n1876), .SEL(n2231), .F(\Data_Mem/n7170 ) );
  MUX U3728 ( .IN0(o[592]), .IN1(n1877), .SEL(n2231), .F(\Data_Mem/n7169 ) );
  NAND U3729 ( .A(n2232), .B(n2233), .Z(n2231) );
  OR U3730 ( .A(n1880), .B(n2229), .Z(n2233) );
  ANDN U3731 ( .A(n2227), .B(n2226), .Z(n2232) );
  NANDN U3732 ( .B(n2229), .A(n1915), .Z(n2227) );
  MUX U3733 ( .IN0(n1883), .IN1(o[591]), .SEL(n2234), .F(\Data_Mem/n7168 ) );
  MUX U3734 ( .IN0(n1885), .IN1(o[590]), .SEL(n2234), .F(\Data_Mem/n7167 ) );
  MUX U3735 ( .IN0(n1886), .IN1(o[589]), .SEL(n2234), .F(\Data_Mem/n7166 ) );
  MUX U3736 ( .IN0(n1887), .IN1(o[588]), .SEL(n2234), .F(\Data_Mem/n7165 ) );
  MUX U3737 ( .IN0(n1888), .IN1(o[587]), .SEL(n2234), .F(\Data_Mem/n7164 ) );
  IV U3738 ( .A(n2235), .Z(n2234) );
  MUX U3739 ( .IN0(o[586]), .IN1(n1890), .SEL(n2235), .F(\Data_Mem/n7163 ) );
  MUX U3740 ( .IN0(o[585]), .IN1(n1891), .SEL(n2235), .F(\Data_Mem/n7162 ) );
  MUX U3741 ( .IN0(o[584]), .IN1(n1892), .SEL(n2235), .F(\Data_Mem/n7161 ) );
  NAND U3742 ( .A(n2236), .B(n2237), .Z(n2235) );
  OR U3743 ( .A(n1895), .B(n2229), .Z(n2237) );
  MUX U3744 ( .IN0(reg_target[7]), .IN1(o[583]), .SEL(n2238), .F(
        \Data_Mem/n7160 ) );
  MUX U3745 ( .IN0(reg_target[6]), .IN1(o[582]), .SEL(n2238), .F(
        \Data_Mem/n7159 ) );
  MUX U3746 ( .IN0(reg_target[5]), .IN1(o[581]), .SEL(n2238), .F(
        \Data_Mem/n7158 ) );
  MUX U3747 ( .IN0(reg_target[4]), .IN1(o[580]), .SEL(n2238), .F(
        \Data_Mem/n7157 ) );
  MUX U3748 ( .IN0(reg_target[3]), .IN1(o[579]), .SEL(n2238), .F(
        \Data_Mem/n7156 ) );
  IV U3749 ( .A(n2239), .Z(n2238) );
  MUX U3750 ( .IN0(o[578]), .IN1(reg_target[2]), .SEL(n2239), .F(
        \Data_Mem/n7155 ) );
  MUX U3751 ( .IN0(o[577]), .IN1(reg_target[1]), .SEL(n2239), .F(
        \Data_Mem/n7154 ) );
  MUX U3752 ( .IN0(o[576]), .IN1(reg_target[0]), .SEL(n2239), .F(
        \Data_Mem/n7153 ) );
  NAND U3753 ( .A(n2236), .B(n2240), .Z(n2239) );
  NANDN U3754 ( .B(n2229), .A(n1899), .Z(n2240) );
  ANDN U3755 ( .A(n2241), .B(n2226), .Z(n2236) );
  ANDN U3756 ( .A(n1902), .B(n2229), .Z(n2226) );
  NANDN U3757 ( .B(n2229), .A(n1924), .Z(n2241) );
  NAND U3758 ( .A(n1944), .B(n2205), .Z(n2229) );
  MUX U3759 ( .IN0(n1853), .IN1(o[639]), .SEL(n2242), .F(\Data_Mem/n7152 ) );
  MUX U3760 ( .IN0(n1855), .IN1(o[638]), .SEL(n2242), .F(\Data_Mem/n7151 ) );
  MUX U3761 ( .IN0(n1856), .IN1(o[637]), .SEL(n2242), .F(\Data_Mem/n7150 ) );
  MUX U3762 ( .IN0(n1857), .IN1(o[636]), .SEL(n2242), .F(\Data_Mem/n7149 ) );
  MUX U3763 ( .IN0(n1858), .IN1(o[635]), .SEL(n2242), .F(\Data_Mem/n7148 ) );
  MUX U3764 ( .IN0(n1859), .IN1(o[634]), .SEL(n2242), .F(\Data_Mem/n7147 ) );
  MUX U3765 ( .IN0(n1860), .IN1(o[633]), .SEL(n2242), .F(\Data_Mem/n7146 ) );
  MUX U3766 ( .IN0(n1861), .IN1(o[632]), .SEL(n2242), .F(\Data_Mem/n7145 ) );
  ANDN U3767 ( .A(n2243), .B(n2244), .Z(n2242) );
  AND U3768 ( .A(n2245), .B(n2246), .Z(n2243) );
  OR U3769 ( .A(n1867), .B(n2247), .Z(n2246) );
  MUX U3770 ( .IN0(n1868), .IN1(o[631]), .SEL(n2248), .F(\Data_Mem/n7144 ) );
  MUX U3771 ( .IN0(n1870), .IN1(o[630]), .SEL(n2248), .F(\Data_Mem/n7143 ) );
  MUX U3772 ( .IN0(n1871), .IN1(o[629]), .SEL(n2248), .F(\Data_Mem/n7142 ) );
  MUX U3773 ( .IN0(n1872), .IN1(o[628]), .SEL(n2248), .F(\Data_Mem/n7141 ) );
  MUX U3774 ( .IN0(n1873), .IN1(o[627]), .SEL(n2248), .F(\Data_Mem/n7140 ) );
  IV U3775 ( .A(n2249), .Z(n2248) );
  MUX U3776 ( .IN0(o[626]), .IN1(n1875), .SEL(n2249), .F(\Data_Mem/n7139 ) );
  MUX U3777 ( .IN0(o[625]), .IN1(n1876), .SEL(n2249), .F(\Data_Mem/n7138 ) );
  MUX U3778 ( .IN0(o[624]), .IN1(n1877), .SEL(n2249), .F(\Data_Mem/n7137 ) );
  NAND U3779 ( .A(n2250), .B(n2251), .Z(n2249) );
  OR U3780 ( .A(n1880), .B(n2247), .Z(n2251) );
  ANDN U3781 ( .A(n2245), .B(n2244), .Z(n2250) );
  NANDN U3782 ( .B(n2247), .A(n1915), .Z(n2245) );
  MUX U3783 ( .IN0(n1883), .IN1(o[623]), .SEL(n2252), .F(\Data_Mem/n7136 ) );
  MUX U3784 ( .IN0(n1885), .IN1(o[622]), .SEL(n2252), .F(\Data_Mem/n7135 ) );
  MUX U3785 ( .IN0(n1886), .IN1(o[621]), .SEL(n2252), .F(\Data_Mem/n7134 ) );
  MUX U3786 ( .IN0(n1887), .IN1(o[620]), .SEL(n2252), .F(\Data_Mem/n7133 ) );
  MUX U3787 ( .IN0(n1888), .IN1(o[619]), .SEL(n2252), .F(\Data_Mem/n7132 ) );
  IV U3788 ( .A(n2253), .Z(n2252) );
  MUX U3789 ( .IN0(o[618]), .IN1(n1890), .SEL(n2253), .F(\Data_Mem/n7131 ) );
  MUX U3790 ( .IN0(o[617]), .IN1(n1891), .SEL(n2253), .F(\Data_Mem/n7130 ) );
  MUX U3791 ( .IN0(o[616]), .IN1(n1892), .SEL(n2253), .F(\Data_Mem/n7129 ) );
  NAND U3792 ( .A(n2254), .B(n2255), .Z(n2253) );
  OR U3793 ( .A(n1895), .B(n2247), .Z(n2255) );
  MUX U3794 ( .IN0(reg_target[7]), .IN1(o[615]), .SEL(n2256), .F(
        \Data_Mem/n7128 ) );
  MUX U3795 ( .IN0(reg_target[6]), .IN1(o[614]), .SEL(n2256), .F(
        \Data_Mem/n7127 ) );
  MUX U3796 ( .IN0(reg_target[5]), .IN1(o[613]), .SEL(n2256), .F(
        \Data_Mem/n7126 ) );
  MUX U3797 ( .IN0(reg_target[4]), .IN1(o[612]), .SEL(n2256), .F(
        \Data_Mem/n7125 ) );
  MUX U3798 ( .IN0(reg_target[3]), .IN1(o[611]), .SEL(n2256), .F(
        \Data_Mem/n7124 ) );
  IV U3799 ( .A(n2257), .Z(n2256) );
  MUX U3800 ( .IN0(o[610]), .IN1(reg_target[2]), .SEL(n2257), .F(
        \Data_Mem/n7123 ) );
  MUX U3801 ( .IN0(o[609]), .IN1(reg_target[1]), .SEL(n2257), .F(
        \Data_Mem/n7122 ) );
  MUX U3802 ( .IN0(o[608]), .IN1(reg_target[0]), .SEL(n2257), .F(
        \Data_Mem/n7121 ) );
  NAND U3803 ( .A(n2254), .B(n2258), .Z(n2257) );
  NANDN U3804 ( .B(n2247), .A(n1899), .Z(n2258) );
  ANDN U3805 ( .A(n2259), .B(n2244), .Z(n2254) );
  ANDN U3806 ( .A(n1902), .B(n2247), .Z(n2244) );
  NANDN U3807 ( .B(n2247), .A(n1924), .Z(n2259) );
  NAND U3808 ( .A(n1963), .B(n2205), .Z(n2247) );
  MUX U3809 ( .IN0(n1853), .IN1(o[671]), .SEL(n2260), .F(\Data_Mem/n7120 ) );
  MUX U3810 ( .IN0(n1855), .IN1(o[670]), .SEL(n2260), .F(\Data_Mem/n7119 ) );
  MUX U3811 ( .IN0(n1856), .IN1(o[669]), .SEL(n2260), .F(\Data_Mem/n7118 ) );
  MUX U3812 ( .IN0(n1857), .IN1(o[668]), .SEL(n2260), .F(\Data_Mem/n7117 ) );
  MUX U3813 ( .IN0(n1858), .IN1(o[667]), .SEL(n2260), .F(\Data_Mem/n7116 ) );
  MUX U3814 ( .IN0(n1859), .IN1(o[666]), .SEL(n2260), .F(\Data_Mem/n7115 ) );
  MUX U3815 ( .IN0(n1860), .IN1(o[665]), .SEL(n2260), .F(\Data_Mem/n7114 ) );
  MUX U3816 ( .IN0(n1861), .IN1(o[664]), .SEL(n2260), .F(\Data_Mem/n7113 ) );
  ANDN U3817 ( .A(n2261), .B(n2262), .Z(n2260) );
  AND U3818 ( .A(n2263), .B(n2264), .Z(n2261) );
  OR U3819 ( .A(n1867), .B(n2265), .Z(n2264) );
  MUX U3820 ( .IN0(n1868), .IN1(o[663]), .SEL(n2266), .F(\Data_Mem/n7112 ) );
  MUX U3821 ( .IN0(n1870), .IN1(o[662]), .SEL(n2266), .F(\Data_Mem/n7111 ) );
  MUX U3822 ( .IN0(n1871), .IN1(o[661]), .SEL(n2266), .F(\Data_Mem/n7110 ) );
  MUX U3823 ( .IN0(n1872), .IN1(o[660]), .SEL(n2266), .F(\Data_Mem/n7109 ) );
  MUX U3824 ( .IN0(n1873), .IN1(o[659]), .SEL(n2266), .F(\Data_Mem/n7108 ) );
  IV U3825 ( .A(n2267), .Z(n2266) );
  MUX U3826 ( .IN0(o[658]), .IN1(n1875), .SEL(n2267), .F(\Data_Mem/n7107 ) );
  MUX U3827 ( .IN0(o[657]), .IN1(n1876), .SEL(n2267), .F(\Data_Mem/n7106 ) );
  MUX U3828 ( .IN0(o[656]), .IN1(n1877), .SEL(n2267), .F(\Data_Mem/n7105 ) );
  NAND U3829 ( .A(n2268), .B(n2269), .Z(n2267) );
  OR U3830 ( .A(n1880), .B(n2265), .Z(n2269) );
  ANDN U3831 ( .A(n2263), .B(n2262), .Z(n2268) );
  NANDN U3832 ( .B(n2265), .A(n1915), .Z(n2263) );
  MUX U3833 ( .IN0(n1883), .IN1(o[655]), .SEL(n2270), .F(\Data_Mem/n7104 ) );
  MUX U3834 ( .IN0(n1885), .IN1(o[654]), .SEL(n2270), .F(\Data_Mem/n7103 ) );
  MUX U3835 ( .IN0(n1886), .IN1(o[653]), .SEL(n2270), .F(\Data_Mem/n7102 ) );
  MUX U3836 ( .IN0(n1887), .IN1(o[652]), .SEL(n2270), .F(\Data_Mem/n7101 ) );
  MUX U3837 ( .IN0(n1888), .IN1(o[651]), .SEL(n2270), .F(\Data_Mem/n7100 ) );
  IV U3838 ( .A(n2271), .Z(n2270) );
  MUX U3839 ( .IN0(o[650]), .IN1(n1890), .SEL(n2271), .F(\Data_Mem/n7099 ) );
  MUX U3840 ( .IN0(o[649]), .IN1(n1891), .SEL(n2271), .F(\Data_Mem/n7098 ) );
  MUX U3841 ( .IN0(o[648]), .IN1(n1892), .SEL(n2271), .F(\Data_Mem/n7097 ) );
  NAND U3842 ( .A(n2272), .B(n2273), .Z(n2271) );
  OR U3843 ( .A(n1895), .B(n2265), .Z(n2273) );
  MUX U3844 ( .IN0(reg_target[7]), .IN1(o[647]), .SEL(n2274), .F(
        \Data_Mem/n7096 ) );
  MUX U3845 ( .IN0(reg_target[6]), .IN1(o[646]), .SEL(n2274), .F(
        \Data_Mem/n7095 ) );
  MUX U3846 ( .IN0(reg_target[5]), .IN1(o[645]), .SEL(n2274), .F(
        \Data_Mem/n7094 ) );
  MUX U3847 ( .IN0(reg_target[4]), .IN1(o[644]), .SEL(n2274), .F(
        \Data_Mem/n7093 ) );
  MUX U3848 ( .IN0(reg_target[3]), .IN1(o[643]), .SEL(n2274), .F(
        \Data_Mem/n7092 ) );
  IV U3849 ( .A(n2275), .Z(n2274) );
  MUX U3850 ( .IN0(o[642]), .IN1(reg_target[2]), .SEL(n2275), .F(
        \Data_Mem/n7091 ) );
  MUX U3851 ( .IN0(o[641]), .IN1(reg_target[1]), .SEL(n2275), .F(
        \Data_Mem/n7090 ) );
  MUX U3852 ( .IN0(o[640]), .IN1(reg_target[0]), .SEL(n2275), .F(
        \Data_Mem/n7089 ) );
  NAND U3853 ( .A(n2272), .B(n2276), .Z(n2275) );
  NANDN U3854 ( .B(n2265), .A(n1899), .Z(n2276) );
  ANDN U3855 ( .A(n2277), .B(n2262), .Z(n2272) );
  ANDN U3856 ( .A(n1902), .B(n2265), .Z(n2262) );
  NANDN U3857 ( .B(n2265), .A(n1924), .Z(n2277) );
  NAND U3858 ( .A(n1982), .B(n2205), .Z(n2265) );
  MUX U3859 ( .IN0(n1853), .IN1(o[703]), .SEL(n2278), .F(\Data_Mem/n7088 ) );
  MUX U3860 ( .IN0(n1855), .IN1(o[702]), .SEL(n2278), .F(\Data_Mem/n7087 ) );
  MUX U3861 ( .IN0(n1856), .IN1(o[701]), .SEL(n2278), .F(\Data_Mem/n7086 ) );
  MUX U3862 ( .IN0(n1857), .IN1(o[700]), .SEL(n2278), .F(\Data_Mem/n7085 ) );
  MUX U3863 ( .IN0(n1858), .IN1(o[699]), .SEL(n2278), .F(\Data_Mem/n7084 ) );
  MUX U3864 ( .IN0(n1859), .IN1(o[698]), .SEL(n2278), .F(\Data_Mem/n7083 ) );
  MUX U3865 ( .IN0(n1860), .IN1(o[697]), .SEL(n2278), .F(\Data_Mem/n7082 ) );
  MUX U3866 ( .IN0(n1861), .IN1(o[696]), .SEL(n2278), .F(\Data_Mem/n7081 ) );
  ANDN U3867 ( .A(n2279), .B(n2280), .Z(n2278) );
  AND U3868 ( .A(n2281), .B(n2282), .Z(n2279) );
  OR U3869 ( .A(n1867), .B(n2283), .Z(n2282) );
  MUX U3870 ( .IN0(n1868), .IN1(o[695]), .SEL(n2284), .F(\Data_Mem/n7080 ) );
  MUX U3871 ( .IN0(n1870), .IN1(o[694]), .SEL(n2284), .F(\Data_Mem/n7079 ) );
  MUX U3872 ( .IN0(n1871), .IN1(o[693]), .SEL(n2284), .F(\Data_Mem/n7078 ) );
  MUX U3873 ( .IN0(n1872), .IN1(o[692]), .SEL(n2284), .F(\Data_Mem/n7077 ) );
  MUX U3874 ( .IN0(n1873), .IN1(o[691]), .SEL(n2284), .F(\Data_Mem/n7076 ) );
  IV U3875 ( .A(n2285), .Z(n2284) );
  MUX U3876 ( .IN0(o[690]), .IN1(n1875), .SEL(n2285), .F(\Data_Mem/n7075 ) );
  MUX U3877 ( .IN0(o[689]), .IN1(n1876), .SEL(n2285), .F(\Data_Mem/n7074 ) );
  MUX U3878 ( .IN0(o[688]), .IN1(n1877), .SEL(n2285), .F(\Data_Mem/n7073 ) );
  NAND U3879 ( .A(n2286), .B(n2287), .Z(n2285) );
  OR U3880 ( .A(n1880), .B(n2283), .Z(n2287) );
  ANDN U3881 ( .A(n2281), .B(n2280), .Z(n2286) );
  NANDN U3882 ( .B(n2283), .A(n1915), .Z(n2281) );
  MUX U3883 ( .IN0(n1883), .IN1(o[687]), .SEL(n2288), .F(\Data_Mem/n7072 ) );
  MUX U3884 ( .IN0(n1885), .IN1(o[686]), .SEL(n2288), .F(\Data_Mem/n7071 ) );
  MUX U3885 ( .IN0(n1886), .IN1(o[685]), .SEL(n2288), .F(\Data_Mem/n7070 ) );
  MUX U3886 ( .IN0(n1887), .IN1(o[684]), .SEL(n2288), .F(\Data_Mem/n7069 ) );
  MUX U3887 ( .IN0(n1888), .IN1(o[683]), .SEL(n2288), .F(\Data_Mem/n7068 ) );
  IV U3888 ( .A(n2289), .Z(n2288) );
  MUX U3889 ( .IN0(o[682]), .IN1(n1890), .SEL(n2289), .F(\Data_Mem/n7067 ) );
  MUX U3890 ( .IN0(o[681]), .IN1(n1891), .SEL(n2289), .F(\Data_Mem/n7066 ) );
  MUX U3891 ( .IN0(o[680]), .IN1(n1892), .SEL(n2289), .F(\Data_Mem/n7065 ) );
  NAND U3892 ( .A(n2290), .B(n2291), .Z(n2289) );
  OR U3893 ( .A(n1895), .B(n2283), .Z(n2291) );
  MUX U3894 ( .IN0(reg_target[7]), .IN1(o[679]), .SEL(n2292), .F(
        \Data_Mem/n7064 ) );
  MUX U3895 ( .IN0(reg_target[6]), .IN1(o[678]), .SEL(n2292), .F(
        \Data_Mem/n7063 ) );
  MUX U3896 ( .IN0(reg_target[5]), .IN1(o[677]), .SEL(n2292), .F(
        \Data_Mem/n7062 ) );
  MUX U3897 ( .IN0(reg_target[4]), .IN1(o[676]), .SEL(n2292), .F(
        \Data_Mem/n7061 ) );
  MUX U3898 ( .IN0(reg_target[3]), .IN1(o[675]), .SEL(n2292), .F(
        \Data_Mem/n7060 ) );
  IV U3899 ( .A(n2293), .Z(n2292) );
  MUX U3900 ( .IN0(o[674]), .IN1(reg_target[2]), .SEL(n2293), .F(
        \Data_Mem/n7059 ) );
  MUX U3901 ( .IN0(o[673]), .IN1(reg_target[1]), .SEL(n2293), .F(
        \Data_Mem/n7058 ) );
  MUX U3902 ( .IN0(o[672]), .IN1(reg_target[0]), .SEL(n2293), .F(
        \Data_Mem/n7057 ) );
  NAND U3903 ( .A(n2290), .B(n2294), .Z(n2293) );
  NANDN U3904 ( .B(n2283), .A(n1899), .Z(n2294) );
  ANDN U3905 ( .A(n2295), .B(n2280), .Z(n2290) );
  ANDN U3906 ( .A(n1902), .B(n2283), .Z(n2280) );
  NANDN U3907 ( .B(n2283), .A(n1924), .Z(n2295) );
  NAND U3908 ( .A(n2001), .B(n2205), .Z(n2283) );
  MUX U3909 ( .IN0(n1853), .IN1(o[735]), .SEL(n2296), .F(\Data_Mem/n7056 ) );
  MUX U3910 ( .IN0(n1855), .IN1(o[734]), .SEL(n2296), .F(\Data_Mem/n7055 ) );
  MUX U3911 ( .IN0(n1856), .IN1(o[733]), .SEL(n2296), .F(\Data_Mem/n7054 ) );
  MUX U3912 ( .IN0(n1857), .IN1(o[732]), .SEL(n2296), .F(\Data_Mem/n7053 ) );
  MUX U3913 ( .IN0(n1858), .IN1(o[731]), .SEL(n2296), .F(\Data_Mem/n7052 ) );
  MUX U3914 ( .IN0(n1859), .IN1(o[730]), .SEL(n2296), .F(\Data_Mem/n7051 ) );
  MUX U3915 ( .IN0(n1860), .IN1(o[729]), .SEL(n2296), .F(\Data_Mem/n7050 ) );
  MUX U3916 ( .IN0(n1861), .IN1(o[728]), .SEL(n2296), .F(\Data_Mem/n7049 ) );
  ANDN U3917 ( .A(n2297), .B(n2298), .Z(n2296) );
  AND U3918 ( .A(n2299), .B(n2300), .Z(n2297) );
  OR U3919 ( .A(n1867), .B(n2301), .Z(n2300) );
  MUX U3920 ( .IN0(n1868), .IN1(o[727]), .SEL(n2302), .F(\Data_Mem/n7048 ) );
  MUX U3921 ( .IN0(n1870), .IN1(o[726]), .SEL(n2302), .F(\Data_Mem/n7047 ) );
  MUX U3922 ( .IN0(n1871), .IN1(o[725]), .SEL(n2302), .F(\Data_Mem/n7046 ) );
  MUX U3923 ( .IN0(n1872), .IN1(o[724]), .SEL(n2302), .F(\Data_Mem/n7045 ) );
  MUX U3924 ( .IN0(n1873), .IN1(o[723]), .SEL(n2302), .F(\Data_Mem/n7044 ) );
  IV U3925 ( .A(n2303), .Z(n2302) );
  MUX U3926 ( .IN0(o[722]), .IN1(n1875), .SEL(n2303), .F(\Data_Mem/n7043 ) );
  MUX U3927 ( .IN0(o[721]), .IN1(n1876), .SEL(n2303), .F(\Data_Mem/n7042 ) );
  MUX U3928 ( .IN0(o[720]), .IN1(n1877), .SEL(n2303), .F(\Data_Mem/n7041 ) );
  NAND U3929 ( .A(n2304), .B(n2305), .Z(n2303) );
  OR U3930 ( .A(n1880), .B(n2301), .Z(n2305) );
  ANDN U3931 ( .A(n2299), .B(n2298), .Z(n2304) );
  NANDN U3932 ( .B(n2301), .A(n1915), .Z(n2299) );
  MUX U3933 ( .IN0(n1883), .IN1(o[719]), .SEL(n2306), .F(\Data_Mem/n7040 ) );
  MUX U3934 ( .IN0(n1885), .IN1(o[718]), .SEL(n2306), .F(\Data_Mem/n7039 ) );
  MUX U3935 ( .IN0(n1886), .IN1(o[717]), .SEL(n2306), .F(\Data_Mem/n7038 ) );
  MUX U3936 ( .IN0(n1887), .IN1(o[716]), .SEL(n2306), .F(\Data_Mem/n7037 ) );
  MUX U3937 ( .IN0(n1888), .IN1(o[715]), .SEL(n2306), .F(\Data_Mem/n7036 ) );
  IV U3938 ( .A(n2307), .Z(n2306) );
  MUX U3939 ( .IN0(o[714]), .IN1(n1890), .SEL(n2307), .F(\Data_Mem/n7035 ) );
  MUX U3940 ( .IN0(o[713]), .IN1(n1891), .SEL(n2307), .F(\Data_Mem/n7034 ) );
  MUX U3941 ( .IN0(o[712]), .IN1(n1892), .SEL(n2307), .F(\Data_Mem/n7033 ) );
  NAND U3942 ( .A(n2308), .B(n2309), .Z(n2307) );
  OR U3943 ( .A(n1895), .B(n2301), .Z(n2309) );
  MUX U3944 ( .IN0(reg_target[7]), .IN1(o[711]), .SEL(n2310), .F(
        \Data_Mem/n7032 ) );
  MUX U3945 ( .IN0(reg_target[6]), .IN1(o[710]), .SEL(n2310), .F(
        \Data_Mem/n7031 ) );
  MUX U3946 ( .IN0(reg_target[5]), .IN1(o[709]), .SEL(n2310), .F(
        \Data_Mem/n7030 ) );
  MUX U3947 ( .IN0(reg_target[4]), .IN1(o[708]), .SEL(n2310), .F(
        \Data_Mem/n7029 ) );
  MUX U3948 ( .IN0(reg_target[3]), .IN1(o[707]), .SEL(n2310), .F(
        \Data_Mem/n7028 ) );
  IV U3949 ( .A(n2311), .Z(n2310) );
  MUX U3950 ( .IN0(o[706]), .IN1(reg_target[2]), .SEL(n2311), .F(
        \Data_Mem/n7027 ) );
  MUX U3951 ( .IN0(o[705]), .IN1(reg_target[1]), .SEL(n2311), .F(
        \Data_Mem/n7026 ) );
  MUX U3952 ( .IN0(o[704]), .IN1(reg_target[0]), .SEL(n2311), .F(
        \Data_Mem/n7025 ) );
  NAND U3953 ( .A(n2308), .B(n2312), .Z(n2311) );
  NANDN U3954 ( .B(n2301), .A(n1899), .Z(n2312) );
  ANDN U3955 ( .A(n2313), .B(n2298), .Z(n2308) );
  ANDN U3956 ( .A(n1902), .B(n2301), .Z(n2298) );
  NANDN U3957 ( .B(n2301), .A(n1924), .Z(n2313) );
  NAND U3958 ( .A(n2020), .B(n2205), .Z(n2301) );
  MUX U3959 ( .IN0(n1853), .IN1(o[767]), .SEL(n2314), .F(\Data_Mem/n7024 ) );
  MUX U3960 ( .IN0(n1855), .IN1(o[766]), .SEL(n2314), .F(\Data_Mem/n7023 ) );
  MUX U3961 ( .IN0(n1856), .IN1(o[765]), .SEL(n2314), .F(\Data_Mem/n7022 ) );
  MUX U3962 ( .IN0(n1857), .IN1(o[764]), .SEL(n2314), .F(\Data_Mem/n7021 ) );
  MUX U3963 ( .IN0(n1858), .IN1(o[763]), .SEL(n2314), .F(\Data_Mem/n7020 ) );
  MUX U3964 ( .IN0(n1859), .IN1(o[762]), .SEL(n2314), .F(\Data_Mem/n7019 ) );
  MUX U3965 ( .IN0(n1860), .IN1(o[761]), .SEL(n2314), .F(\Data_Mem/n7018 ) );
  MUX U3966 ( .IN0(n1861), .IN1(o[760]), .SEL(n2314), .F(\Data_Mem/n7017 ) );
  ANDN U3967 ( .A(n2315), .B(n2316), .Z(n2314) );
  AND U3968 ( .A(n2317), .B(n2318), .Z(n2315) );
  OR U3969 ( .A(n1867), .B(n2319), .Z(n2318) );
  MUX U3970 ( .IN0(n1868), .IN1(o[759]), .SEL(n2320), .F(\Data_Mem/n7016 ) );
  MUX U3971 ( .IN0(n1870), .IN1(o[758]), .SEL(n2320), .F(\Data_Mem/n7015 ) );
  MUX U3972 ( .IN0(n1871), .IN1(o[757]), .SEL(n2320), .F(\Data_Mem/n7014 ) );
  MUX U3973 ( .IN0(n1872), .IN1(o[756]), .SEL(n2320), .F(\Data_Mem/n7013 ) );
  MUX U3974 ( .IN0(n1873), .IN1(o[755]), .SEL(n2320), .F(\Data_Mem/n7012 ) );
  IV U3975 ( .A(n2321), .Z(n2320) );
  MUX U3976 ( .IN0(o[754]), .IN1(n1875), .SEL(n2321), .F(\Data_Mem/n7011 ) );
  MUX U3977 ( .IN0(o[753]), .IN1(n1876), .SEL(n2321), .F(\Data_Mem/n7010 ) );
  MUX U3978 ( .IN0(o[752]), .IN1(n1877), .SEL(n2321), .F(\Data_Mem/n7009 ) );
  NAND U3979 ( .A(n2322), .B(n2323), .Z(n2321) );
  OR U3980 ( .A(n1880), .B(n2319), .Z(n2323) );
  ANDN U3981 ( .A(n2317), .B(n2316), .Z(n2322) );
  NANDN U3982 ( .B(n2319), .A(n1915), .Z(n2317) );
  MUX U3983 ( .IN0(n1883), .IN1(o[751]), .SEL(n2324), .F(\Data_Mem/n7008 ) );
  MUX U3984 ( .IN0(n1885), .IN1(o[750]), .SEL(n2324), .F(\Data_Mem/n7007 ) );
  MUX U3985 ( .IN0(n1886), .IN1(o[749]), .SEL(n2324), .F(\Data_Mem/n7006 ) );
  MUX U3986 ( .IN0(n1887), .IN1(o[748]), .SEL(n2324), .F(\Data_Mem/n7005 ) );
  MUX U3987 ( .IN0(n1888), .IN1(o[747]), .SEL(n2324), .F(\Data_Mem/n7004 ) );
  IV U3988 ( .A(n2325), .Z(n2324) );
  MUX U3989 ( .IN0(o[746]), .IN1(n1890), .SEL(n2325), .F(\Data_Mem/n7003 ) );
  MUX U3990 ( .IN0(o[745]), .IN1(n1891), .SEL(n2325), .F(\Data_Mem/n7002 ) );
  MUX U3991 ( .IN0(o[744]), .IN1(n1892), .SEL(n2325), .F(\Data_Mem/n7001 ) );
  NAND U3992 ( .A(n2326), .B(n2327), .Z(n2325) );
  OR U3993 ( .A(n1895), .B(n2319), .Z(n2327) );
  MUX U3994 ( .IN0(reg_target[7]), .IN1(o[743]), .SEL(n2328), .F(
        \Data_Mem/n7000 ) );
  MUX U3995 ( .IN0(reg_target[6]), .IN1(o[742]), .SEL(n2328), .F(
        \Data_Mem/n6999 ) );
  MUX U3996 ( .IN0(reg_target[5]), .IN1(o[741]), .SEL(n2328), .F(
        \Data_Mem/n6998 ) );
  MUX U3997 ( .IN0(reg_target[4]), .IN1(o[740]), .SEL(n2328), .F(
        \Data_Mem/n6997 ) );
  MUX U3998 ( .IN0(reg_target[3]), .IN1(o[739]), .SEL(n2328), .F(
        \Data_Mem/n6996 ) );
  IV U3999 ( .A(n2329), .Z(n2328) );
  MUX U4000 ( .IN0(o[738]), .IN1(reg_target[2]), .SEL(n2329), .F(
        \Data_Mem/n6995 ) );
  MUX U4001 ( .IN0(o[737]), .IN1(reg_target[1]), .SEL(n2329), .F(
        \Data_Mem/n6994 ) );
  MUX U4002 ( .IN0(o[736]), .IN1(reg_target[0]), .SEL(n2329), .F(
        \Data_Mem/n6993 ) );
  NAND U4003 ( .A(n2326), .B(n2330), .Z(n2329) );
  NANDN U4004 ( .B(n2319), .A(n1899), .Z(n2330) );
  ANDN U4005 ( .A(n2331), .B(n2316), .Z(n2326) );
  ANDN U4006 ( .A(n1902), .B(n2319), .Z(n2316) );
  NANDN U4007 ( .B(n2319), .A(n1924), .Z(n2331) );
  NAND U4008 ( .A(n2205), .B(n2039), .Z(n2319) );
  AND U4009 ( .A(n2332), .B(n485), .Z(n2205) );
  MUX U4010 ( .IN0(n1853), .IN1(o[799]), .SEL(n2333), .F(\Data_Mem/n6992 ) );
  MUX U4011 ( .IN0(n1855), .IN1(o[798]), .SEL(n2333), .F(\Data_Mem/n6991 ) );
  MUX U4012 ( .IN0(n1856), .IN1(o[797]), .SEL(n2333), .F(\Data_Mem/n6990 ) );
  MUX U4013 ( .IN0(n1857), .IN1(o[796]), .SEL(n2333), .F(\Data_Mem/n6989 ) );
  MUX U4014 ( .IN0(n1858), .IN1(o[795]), .SEL(n2333), .F(\Data_Mem/n6988 ) );
  MUX U4015 ( .IN0(n1859), .IN1(o[794]), .SEL(n2333), .F(\Data_Mem/n6987 ) );
  MUX U4016 ( .IN0(n1860), .IN1(o[793]), .SEL(n2333), .F(\Data_Mem/n6986 ) );
  MUX U4017 ( .IN0(n1861), .IN1(o[792]), .SEL(n2333), .F(\Data_Mem/n6985 ) );
  ANDN U4018 ( .A(n2334), .B(n2335), .Z(n2333) );
  AND U4019 ( .A(n2336), .B(n2337), .Z(n2334) );
  OR U4020 ( .A(n1867), .B(n2338), .Z(n2337) );
  MUX U4021 ( .IN0(n1868), .IN1(o[791]), .SEL(n2339), .F(\Data_Mem/n6984 ) );
  MUX U4022 ( .IN0(n1870), .IN1(o[790]), .SEL(n2339), .F(\Data_Mem/n6983 ) );
  MUX U4023 ( .IN0(n1871), .IN1(o[789]), .SEL(n2339), .F(\Data_Mem/n6982 ) );
  MUX U4024 ( .IN0(n1872), .IN1(o[788]), .SEL(n2339), .F(\Data_Mem/n6981 ) );
  MUX U4025 ( .IN0(n1873), .IN1(o[787]), .SEL(n2339), .F(\Data_Mem/n6980 ) );
  IV U4026 ( .A(n2340), .Z(n2339) );
  MUX U4027 ( .IN0(o[786]), .IN1(n1875), .SEL(n2340), .F(\Data_Mem/n6979 ) );
  MUX U4028 ( .IN0(o[785]), .IN1(n1876), .SEL(n2340), .F(\Data_Mem/n6978 ) );
  MUX U4029 ( .IN0(o[784]), .IN1(n1877), .SEL(n2340), .F(\Data_Mem/n6977 ) );
  NAND U4030 ( .A(n2341), .B(n2342), .Z(n2340) );
  OR U4031 ( .A(n1880), .B(n2338), .Z(n2342) );
  ANDN U4032 ( .A(n2336), .B(n2335), .Z(n2341) );
  NANDN U4033 ( .B(n2338), .A(n1915), .Z(n2336) );
  MUX U4034 ( .IN0(n1883), .IN1(o[783]), .SEL(n2343), .F(\Data_Mem/n6976 ) );
  MUX U4035 ( .IN0(n1885), .IN1(o[782]), .SEL(n2343), .F(\Data_Mem/n6975 ) );
  MUX U4036 ( .IN0(n1886), .IN1(o[781]), .SEL(n2343), .F(\Data_Mem/n6974 ) );
  MUX U4037 ( .IN0(n1887), .IN1(o[780]), .SEL(n2343), .F(\Data_Mem/n6973 ) );
  MUX U4038 ( .IN0(n1888), .IN1(o[779]), .SEL(n2343), .F(\Data_Mem/n6972 ) );
  IV U4039 ( .A(n2344), .Z(n2343) );
  MUX U4040 ( .IN0(o[778]), .IN1(n1890), .SEL(n2344), .F(\Data_Mem/n6971 ) );
  MUX U4041 ( .IN0(o[777]), .IN1(n1891), .SEL(n2344), .F(\Data_Mem/n6970 ) );
  MUX U4042 ( .IN0(o[776]), .IN1(n1892), .SEL(n2344), .F(\Data_Mem/n6969 ) );
  NAND U4043 ( .A(n2345), .B(n2346), .Z(n2344) );
  OR U4044 ( .A(n1895), .B(n2338), .Z(n2346) );
  MUX U4045 ( .IN0(reg_target[7]), .IN1(o[775]), .SEL(n2347), .F(
        \Data_Mem/n6968 ) );
  MUX U4046 ( .IN0(reg_target[6]), .IN1(o[774]), .SEL(n2347), .F(
        \Data_Mem/n6967 ) );
  MUX U4047 ( .IN0(reg_target[5]), .IN1(o[773]), .SEL(n2347), .F(
        \Data_Mem/n6966 ) );
  MUX U4048 ( .IN0(reg_target[4]), .IN1(o[772]), .SEL(n2347), .F(
        \Data_Mem/n6965 ) );
  MUX U4049 ( .IN0(reg_target[3]), .IN1(o[771]), .SEL(n2347), .F(
        \Data_Mem/n6964 ) );
  IV U4050 ( .A(n2348), .Z(n2347) );
  MUX U4051 ( .IN0(o[770]), .IN1(reg_target[2]), .SEL(n2348), .F(
        \Data_Mem/n6963 ) );
  MUX U4052 ( .IN0(o[769]), .IN1(reg_target[1]), .SEL(n2348), .F(
        \Data_Mem/n6962 ) );
  MUX U4053 ( .IN0(o[768]), .IN1(reg_target[0]), .SEL(n2348), .F(
        \Data_Mem/n6961 ) );
  NAND U4054 ( .A(n2345), .B(n2349), .Z(n2348) );
  NANDN U4055 ( .B(n2338), .A(n1899), .Z(n2349) );
  ANDN U4056 ( .A(n2350), .B(n2335), .Z(n2345) );
  ANDN U4057 ( .A(n1902), .B(n2338), .Z(n2335) );
  NANDN U4058 ( .B(n2338), .A(n1924), .Z(n2350) );
  NAND U4059 ( .A(n1903), .B(n2351), .Z(n2338) );
  MUX U4060 ( .IN0(n1853), .IN1(o[831]), .SEL(n2352), .F(\Data_Mem/n6960 ) );
  MUX U4061 ( .IN0(n1855), .IN1(o[830]), .SEL(n2352), .F(\Data_Mem/n6959 ) );
  MUX U4062 ( .IN0(n1856), .IN1(o[829]), .SEL(n2352), .F(\Data_Mem/n6958 ) );
  MUX U4063 ( .IN0(n1857), .IN1(o[828]), .SEL(n2352), .F(\Data_Mem/n6957 ) );
  MUX U4064 ( .IN0(n1858), .IN1(o[827]), .SEL(n2352), .F(\Data_Mem/n6956 ) );
  MUX U4065 ( .IN0(n1859), .IN1(o[826]), .SEL(n2352), .F(\Data_Mem/n6955 ) );
  MUX U4066 ( .IN0(n1860), .IN1(o[825]), .SEL(n2352), .F(\Data_Mem/n6954 ) );
  MUX U4067 ( .IN0(n1861), .IN1(o[824]), .SEL(n2352), .F(\Data_Mem/n6953 ) );
  ANDN U4068 ( .A(n2353), .B(n2354), .Z(n2352) );
  AND U4069 ( .A(n2355), .B(n2356), .Z(n2353) );
  OR U4070 ( .A(n1867), .B(n2357), .Z(n2356) );
  MUX U4071 ( .IN0(n1868), .IN1(o[823]), .SEL(n2358), .F(\Data_Mem/n6952 ) );
  MUX U4072 ( .IN0(n1870), .IN1(o[822]), .SEL(n2358), .F(\Data_Mem/n6951 ) );
  MUX U4073 ( .IN0(n1871), .IN1(o[821]), .SEL(n2358), .F(\Data_Mem/n6950 ) );
  MUX U4074 ( .IN0(n1872), .IN1(o[820]), .SEL(n2358), .F(\Data_Mem/n6949 ) );
  MUX U4075 ( .IN0(n1873), .IN1(o[819]), .SEL(n2358), .F(\Data_Mem/n6948 ) );
  IV U4076 ( .A(n2359), .Z(n2358) );
  MUX U4077 ( .IN0(o[818]), .IN1(n1875), .SEL(n2359), .F(\Data_Mem/n6947 ) );
  MUX U4078 ( .IN0(o[817]), .IN1(n1876), .SEL(n2359), .F(\Data_Mem/n6946 ) );
  MUX U4079 ( .IN0(o[816]), .IN1(n1877), .SEL(n2359), .F(\Data_Mem/n6945 ) );
  NAND U4080 ( .A(n2360), .B(n2361), .Z(n2359) );
  OR U4081 ( .A(n1880), .B(n2357), .Z(n2361) );
  ANDN U4082 ( .A(n2355), .B(n2354), .Z(n2360) );
  NANDN U4083 ( .B(n2357), .A(n1915), .Z(n2355) );
  MUX U4084 ( .IN0(n1883), .IN1(o[815]), .SEL(n2362), .F(\Data_Mem/n6944 ) );
  MUX U4085 ( .IN0(n1885), .IN1(o[814]), .SEL(n2362), .F(\Data_Mem/n6943 ) );
  MUX U4086 ( .IN0(n1886), .IN1(o[813]), .SEL(n2362), .F(\Data_Mem/n6942 ) );
  MUX U4087 ( .IN0(n1887), .IN1(o[812]), .SEL(n2362), .F(\Data_Mem/n6941 ) );
  MUX U4088 ( .IN0(n1888), .IN1(o[811]), .SEL(n2362), .F(\Data_Mem/n6940 ) );
  IV U4089 ( .A(n2363), .Z(n2362) );
  MUX U4090 ( .IN0(o[810]), .IN1(n1890), .SEL(n2363), .F(\Data_Mem/n6939 ) );
  MUX U4091 ( .IN0(o[809]), .IN1(n1891), .SEL(n2363), .F(\Data_Mem/n6938 ) );
  MUX U4092 ( .IN0(o[808]), .IN1(n1892), .SEL(n2363), .F(\Data_Mem/n6937 ) );
  NAND U4093 ( .A(n2364), .B(n2365), .Z(n2363) );
  OR U4094 ( .A(n1895), .B(n2357), .Z(n2365) );
  MUX U4095 ( .IN0(reg_target[7]), .IN1(o[807]), .SEL(n2366), .F(
        \Data_Mem/n6936 ) );
  MUX U4096 ( .IN0(reg_target[6]), .IN1(o[806]), .SEL(n2366), .F(
        \Data_Mem/n6935 ) );
  MUX U4097 ( .IN0(reg_target[5]), .IN1(o[805]), .SEL(n2366), .F(
        \Data_Mem/n6934 ) );
  MUX U4098 ( .IN0(reg_target[4]), .IN1(o[804]), .SEL(n2366), .F(
        \Data_Mem/n6933 ) );
  MUX U4099 ( .IN0(reg_target[3]), .IN1(o[803]), .SEL(n2366), .F(
        \Data_Mem/n6932 ) );
  IV U4100 ( .A(n2367), .Z(n2366) );
  MUX U4101 ( .IN0(o[802]), .IN1(reg_target[2]), .SEL(n2367), .F(
        \Data_Mem/n6931 ) );
  MUX U4102 ( .IN0(o[801]), .IN1(reg_target[1]), .SEL(n2367), .F(
        \Data_Mem/n6930 ) );
  MUX U4103 ( .IN0(o[800]), .IN1(reg_target[0]), .SEL(n2367), .F(
        \Data_Mem/n6929 ) );
  NAND U4104 ( .A(n2364), .B(n2368), .Z(n2367) );
  NANDN U4105 ( .B(n2357), .A(n1899), .Z(n2368) );
  ANDN U4106 ( .A(n2369), .B(n2354), .Z(n2364) );
  ANDN U4107 ( .A(n1902), .B(n2357), .Z(n2354) );
  NANDN U4108 ( .B(n2357), .A(n1924), .Z(n2369) );
  NAND U4109 ( .A(n1925), .B(n2351), .Z(n2357) );
  MUX U4110 ( .IN0(n1853), .IN1(o[863]), .SEL(n2370), .F(\Data_Mem/n6928 ) );
  MUX U4111 ( .IN0(n1855), .IN1(o[862]), .SEL(n2370), .F(\Data_Mem/n6927 ) );
  MUX U4112 ( .IN0(n1856), .IN1(o[861]), .SEL(n2370), .F(\Data_Mem/n6926 ) );
  MUX U4113 ( .IN0(n1857), .IN1(o[860]), .SEL(n2370), .F(\Data_Mem/n6925 ) );
  MUX U4114 ( .IN0(n1858), .IN1(o[859]), .SEL(n2370), .F(\Data_Mem/n6924 ) );
  MUX U4115 ( .IN0(n1859), .IN1(o[858]), .SEL(n2370), .F(\Data_Mem/n6923 ) );
  MUX U4116 ( .IN0(n1860), .IN1(o[857]), .SEL(n2370), .F(\Data_Mem/n6922 ) );
  MUX U4117 ( .IN0(n1861), .IN1(o[856]), .SEL(n2370), .F(\Data_Mem/n6921 ) );
  ANDN U4118 ( .A(n2371), .B(n2372), .Z(n2370) );
  AND U4119 ( .A(n2373), .B(n2374), .Z(n2371) );
  OR U4120 ( .A(n1867), .B(n2375), .Z(n2374) );
  MUX U4121 ( .IN0(n1868), .IN1(o[855]), .SEL(n2376), .F(\Data_Mem/n6920 ) );
  MUX U4122 ( .IN0(n1870), .IN1(o[854]), .SEL(n2376), .F(\Data_Mem/n6919 ) );
  MUX U4123 ( .IN0(n1871), .IN1(o[853]), .SEL(n2376), .F(\Data_Mem/n6918 ) );
  MUX U4124 ( .IN0(n1872), .IN1(o[852]), .SEL(n2376), .F(\Data_Mem/n6917 ) );
  MUX U4125 ( .IN0(n1873), .IN1(o[851]), .SEL(n2376), .F(\Data_Mem/n6916 ) );
  IV U4126 ( .A(n2377), .Z(n2376) );
  MUX U4127 ( .IN0(o[850]), .IN1(n1875), .SEL(n2377), .F(\Data_Mem/n6915 ) );
  MUX U4128 ( .IN0(o[849]), .IN1(n1876), .SEL(n2377), .F(\Data_Mem/n6914 ) );
  MUX U4129 ( .IN0(o[848]), .IN1(n1877), .SEL(n2377), .F(\Data_Mem/n6913 ) );
  NAND U4130 ( .A(n2378), .B(n2379), .Z(n2377) );
  OR U4131 ( .A(n1880), .B(n2375), .Z(n2379) );
  ANDN U4132 ( .A(n2373), .B(n2372), .Z(n2378) );
  NANDN U4133 ( .B(n2375), .A(n1915), .Z(n2373) );
  MUX U4134 ( .IN0(n1883), .IN1(o[847]), .SEL(n2380), .F(\Data_Mem/n6912 ) );
  MUX U4135 ( .IN0(n1885), .IN1(o[846]), .SEL(n2380), .F(\Data_Mem/n6911 ) );
  MUX U4136 ( .IN0(n1886), .IN1(o[845]), .SEL(n2380), .F(\Data_Mem/n6910 ) );
  MUX U4137 ( .IN0(n1887), .IN1(o[844]), .SEL(n2380), .F(\Data_Mem/n6909 ) );
  MUX U4138 ( .IN0(n1888), .IN1(o[843]), .SEL(n2380), .F(\Data_Mem/n6908 ) );
  IV U4139 ( .A(n2381), .Z(n2380) );
  MUX U4140 ( .IN0(o[842]), .IN1(n1890), .SEL(n2381), .F(\Data_Mem/n6907 ) );
  MUX U4141 ( .IN0(o[841]), .IN1(n1891), .SEL(n2381), .F(\Data_Mem/n6906 ) );
  MUX U4142 ( .IN0(o[840]), .IN1(n1892), .SEL(n2381), .F(\Data_Mem/n6905 ) );
  NAND U4143 ( .A(n2382), .B(n2383), .Z(n2381) );
  OR U4144 ( .A(n1895), .B(n2375), .Z(n2383) );
  MUX U4145 ( .IN0(reg_target[7]), .IN1(o[839]), .SEL(n2384), .F(
        \Data_Mem/n6904 ) );
  MUX U4146 ( .IN0(reg_target[6]), .IN1(o[838]), .SEL(n2384), .F(
        \Data_Mem/n6903 ) );
  MUX U4147 ( .IN0(reg_target[5]), .IN1(o[837]), .SEL(n2384), .F(
        \Data_Mem/n6902 ) );
  MUX U4148 ( .IN0(reg_target[4]), .IN1(o[836]), .SEL(n2384), .F(
        \Data_Mem/n6901 ) );
  MUX U4149 ( .IN0(reg_target[3]), .IN1(o[835]), .SEL(n2384), .F(
        \Data_Mem/n6900 ) );
  IV U4150 ( .A(n2385), .Z(n2384) );
  MUX U4151 ( .IN0(o[834]), .IN1(reg_target[2]), .SEL(n2385), .F(
        \Data_Mem/n6899 ) );
  MUX U4152 ( .IN0(o[833]), .IN1(reg_target[1]), .SEL(n2385), .F(
        \Data_Mem/n6898 ) );
  MUX U4153 ( .IN0(o[832]), .IN1(reg_target[0]), .SEL(n2385), .F(
        \Data_Mem/n6897 ) );
  NAND U4154 ( .A(n2382), .B(n2386), .Z(n2385) );
  NANDN U4155 ( .B(n2375), .A(n1899), .Z(n2386) );
  ANDN U4156 ( .A(n2387), .B(n2372), .Z(n2382) );
  ANDN U4157 ( .A(n1902), .B(n2375), .Z(n2372) );
  NANDN U4158 ( .B(n2375), .A(n1924), .Z(n2387) );
  NAND U4159 ( .A(n1944), .B(n2351), .Z(n2375) );
  MUX U4160 ( .IN0(n1853), .IN1(o[895]), .SEL(n2388), .F(\Data_Mem/n6896 ) );
  MUX U4161 ( .IN0(n1855), .IN1(o[894]), .SEL(n2388), .F(\Data_Mem/n6895 ) );
  MUX U4162 ( .IN0(n1856), .IN1(o[893]), .SEL(n2388), .F(\Data_Mem/n6894 ) );
  MUX U4163 ( .IN0(n1857), .IN1(o[892]), .SEL(n2388), .F(\Data_Mem/n6893 ) );
  MUX U4164 ( .IN0(n1858), .IN1(o[891]), .SEL(n2388), .F(\Data_Mem/n6892 ) );
  MUX U4165 ( .IN0(n1859), .IN1(o[890]), .SEL(n2388), .F(\Data_Mem/n6891 ) );
  MUX U4166 ( .IN0(n1860), .IN1(o[889]), .SEL(n2388), .F(\Data_Mem/n6890 ) );
  MUX U4167 ( .IN0(n1861), .IN1(o[888]), .SEL(n2388), .F(\Data_Mem/n6889 ) );
  ANDN U4168 ( .A(n2389), .B(n2390), .Z(n2388) );
  AND U4169 ( .A(n2391), .B(n2392), .Z(n2389) );
  OR U4170 ( .A(n1867), .B(n2393), .Z(n2392) );
  MUX U4171 ( .IN0(n1868), .IN1(o[887]), .SEL(n2394), .F(\Data_Mem/n6888 ) );
  MUX U4172 ( .IN0(n1870), .IN1(o[886]), .SEL(n2394), .F(\Data_Mem/n6887 ) );
  MUX U4173 ( .IN0(n1871), .IN1(o[885]), .SEL(n2394), .F(\Data_Mem/n6886 ) );
  MUX U4174 ( .IN0(n1872), .IN1(o[884]), .SEL(n2394), .F(\Data_Mem/n6885 ) );
  MUX U4175 ( .IN0(n1873), .IN1(o[883]), .SEL(n2394), .F(\Data_Mem/n6884 ) );
  IV U4176 ( .A(n2395), .Z(n2394) );
  MUX U4177 ( .IN0(o[882]), .IN1(n1875), .SEL(n2395), .F(\Data_Mem/n6883 ) );
  MUX U4178 ( .IN0(o[881]), .IN1(n1876), .SEL(n2395), .F(\Data_Mem/n6882 ) );
  MUX U4179 ( .IN0(o[880]), .IN1(n1877), .SEL(n2395), .F(\Data_Mem/n6881 ) );
  NAND U4180 ( .A(n2396), .B(n2397), .Z(n2395) );
  OR U4181 ( .A(n1880), .B(n2393), .Z(n2397) );
  ANDN U4182 ( .A(n2391), .B(n2390), .Z(n2396) );
  NANDN U4183 ( .B(n2393), .A(n1915), .Z(n2391) );
  MUX U4184 ( .IN0(n1883), .IN1(o[879]), .SEL(n2398), .F(\Data_Mem/n6880 ) );
  MUX U4185 ( .IN0(n1885), .IN1(o[878]), .SEL(n2398), .F(\Data_Mem/n6879 ) );
  MUX U4186 ( .IN0(n1886), .IN1(o[877]), .SEL(n2398), .F(\Data_Mem/n6878 ) );
  MUX U4187 ( .IN0(n1887), .IN1(o[876]), .SEL(n2398), .F(\Data_Mem/n6877 ) );
  MUX U4188 ( .IN0(n1888), .IN1(o[875]), .SEL(n2398), .F(\Data_Mem/n6876 ) );
  IV U4189 ( .A(n2399), .Z(n2398) );
  MUX U4190 ( .IN0(o[874]), .IN1(n1890), .SEL(n2399), .F(\Data_Mem/n6875 ) );
  MUX U4191 ( .IN0(o[873]), .IN1(n1891), .SEL(n2399), .F(\Data_Mem/n6874 ) );
  MUX U4192 ( .IN0(o[872]), .IN1(n1892), .SEL(n2399), .F(\Data_Mem/n6873 ) );
  NAND U4193 ( .A(n2400), .B(n2401), .Z(n2399) );
  OR U4194 ( .A(n1895), .B(n2393), .Z(n2401) );
  MUX U4195 ( .IN0(reg_target[7]), .IN1(o[871]), .SEL(n2402), .F(
        \Data_Mem/n6872 ) );
  MUX U4196 ( .IN0(reg_target[6]), .IN1(o[870]), .SEL(n2402), .F(
        \Data_Mem/n6871 ) );
  MUX U4197 ( .IN0(reg_target[5]), .IN1(o[869]), .SEL(n2402), .F(
        \Data_Mem/n6870 ) );
  MUX U4198 ( .IN0(reg_target[4]), .IN1(o[868]), .SEL(n2402), .F(
        \Data_Mem/n6869 ) );
  MUX U4199 ( .IN0(reg_target[3]), .IN1(o[867]), .SEL(n2402), .F(
        \Data_Mem/n6868 ) );
  IV U4200 ( .A(n2403), .Z(n2402) );
  MUX U4201 ( .IN0(o[866]), .IN1(reg_target[2]), .SEL(n2403), .F(
        \Data_Mem/n6867 ) );
  MUX U4202 ( .IN0(o[865]), .IN1(reg_target[1]), .SEL(n2403), .F(
        \Data_Mem/n6866 ) );
  MUX U4203 ( .IN0(o[864]), .IN1(reg_target[0]), .SEL(n2403), .F(
        \Data_Mem/n6865 ) );
  NAND U4204 ( .A(n2400), .B(n2404), .Z(n2403) );
  NANDN U4205 ( .B(n2393), .A(n1899), .Z(n2404) );
  ANDN U4206 ( .A(n2405), .B(n2390), .Z(n2400) );
  ANDN U4207 ( .A(n1902), .B(n2393), .Z(n2390) );
  NANDN U4208 ( .B(n2393), .A(n1924), .Z(n2405) );
  NAND U4209 ( .A(n1963), .B(n2351), .Z(n2393) );
  MUX U4210 ( .IN0(n1853), .IN1(o[927]), .SEL(n2406), .F(\Data_Mem/n6864 ) );
  MUX U4211 ( .IN0(n1855), .IN1(o[926]), .SEL(n2406), .F(\Data_Mem/n6863 ) );
  MUX U4212 ( .IN0(n1856), .IN1(o[925]), .SEL(n2406), .F(\Data_Mem/n6862 ) );
  MUX U4213 ( .IN0(n1857), .IN1(o[924]), .SEL(n2406), .F(\Data_Mem/n6861 ) );
  MUX U4214 ( .IN0(n1858), .IN1(o[923]), .SEL(n2406), .F(\Data_Mem/n6860 ) );
  MUX U4215 ( .IN0(n1859), .IN1(o[922]), .SEL(n2406), .F(\Data_Mem/n6859 ) );
  MUX U4216 ( .IN0(n1860), .IN1(o[921]), .SEL(n2406), .F(\Data_Mem/n6858 ) );
  MUX U4217 ( .IN0(n1861), .IN1(o[920]), .SEL(n2406), .F(\Data_Mem/n6857 ) );
  ANDN U4218 ( .A(n2407), .B(n2408), .Z(n2406) );
  AND U4219 ( .A(n2409), .B(n2410), .Z(n2407) );
  OR U4220 ( .A(n1867), .B(n2411), .Z(n2410) );
  MUX U4221 ( .IN0(n1868), .IN1(o[919]), .SEL(n2412), .F(\Data_Mem/n6856 ) );
  MUX U4222 ( .IN0(n1870), .IN1(o[918]), .SEL(n2412), .F(\Data_Mem/n6855 ) );
  MUX U4223 ( .IN0(n1871), .IN1(o[917]), .SEL(n2412), .F(\Data_Mem/n6854 ) );
  MUX U4224 ( .IN0(n1872), .IN1(o[916]), .SEL(n2412), .F(\Data_Mem/n6853 ) );
  MUX U4225 ( .IN0(n1873), .IN1(o[915]), .SEL(n2412), .F(\Data_Mem/n6852 ) );
  IV U4226 ( .A(n2413), .Z(n2412) );
  MUX U4227 ( .IN0(o[914]), .IN1(n1875), .SEL(n2413), .F(\Data_Mem/n6851 ) );
  MUX U4228 ( .IN0(o[913]), .IN1(n1876), .SEL(n2413), .F(\Data_Mem/n6850 ) );
  MUX U4229 ( .IN0(o[912]), .IN1(n1877), .SEL(n2413), .F(\Data_Mem/n6849 ) );
  NAND U4230 ( .A(n2414), .B(n2415), .Z(n2413) );
  OR U4231 ( .A(n1880), .B(n2411), .Z(n2415) );
  ANDN U4232 ( .A(n2409), .B(n2408), .Z(n2414) );
  NANDN U4233 ( .B(n2411), .A(n1915), .Z(n2409) );
  MUX U4234 ( .IN0(n1883), .IN1(o[911]), .SEL(n2416), .F(\Data_Mem/n6848 ) );
  MUX U4235 ( .IN0(n1885), .IN1(o[910]), .SEL(n2416), .F(\Data_Mem/n6847 ) );
  MUX U4236 ( .IN0(n1886), .IN1(o[909]), .SEL(n2416), .F(\Data_Mem/n6846 ) );
  MUX U4237 ( .IN0(n1887), .IN1(o[908]), .SEL(n2416), .F(\Data_Mem/n6845 ) );
  MUX U4238 ( .IN0(n1888), .IN1(o[907]), .SEL(n2416), .F(\Data_Mem/n6844 ) );
  IV U4239 ( .A(n2417), .Z(n2416) );
  MUX U4240 ( .IN0(o[906]), .IN1(n1890), .SEL(n2417), .F(\Data_Mem/n6843 ) );
  MUX U4241 ( .IN0(o[905]), .IN1(n1891), .SEL(n2417), .F(\Data_Mem/n6842 ) );
  MUX U4242 ( .IN0(o[904]), .IN1(n1892), .SEL(n2417), .F(\Data_Mem/n6841 ) );
  NAND U4243 ( .A(n2418), .B(n2419), .Z(n2417) );
  OR U4244 ( .A(n1895), .B(n2411), .Z(n2419) );
  MUX U4245 ( .IN0(reg_target[7]), .IN1(o[903]), .SEL(n2420), .F(
        \Data_Mem/n6840 ) );
  MUX U4246 ( .IN0(reg_target[6]), .IN1(o[902]), .SEL(n2420), .F(
        \Data_Mem/n6839 ) );
  MUX U4247 ( .IN0(reg_target[5]), .IN1(o[901]), .SEL(n2420), .F(
        \Data_Mem/n6838 ) );
  MUX U4248 ( .IN0(reg_target[4]), .IN1(o[900]), .SEL(n2420), .F(
        \Data_Mem/n6837 ) );
  MUX U4249 ( .IN0(reg_target[3]), .IN1(o[899]), .SEL(n2420), .F(
        \Data_Mem/n6836 ) );
  IV U4250 ( .A(n2421), .Z(n2420) );
  MUX U4251 ( .IN0(o[898]), .IN1(reg_target[2]), .SEL(n2421), .F(
        \Data_Mem/n6835 ) );
  MUX U4252 ( .IN0(o[897]), .IN1(reg_target[1]), .SEL(n2421), .F(
        \Data_Mem/n6834 ) );
  MUX U4253 ( .IN0(o[896]), .IN1(reg_target[0]), .SEL(n2421), .F(
        \Data_Mem/n6833 ) );
  NAND U4254 ( .A(n2418), .B(n2422), .Z(n2421) );
  NANDN U4255 ( .B(n2411), .A(n1899), .Z(n2422) );
  ANDN U4256 ( .A(n2423), .B(n2408), .Z(n2418) );
  ANDN U4257 ( .A(n1902), .B(n2411), .Z(n2408) );
  NANDN U4258 ( .B(n2411), .A(n1924), .Z(n2423) );
  NAND U4259 ( .A(n1982), .B(n2351), .Z(n2411) );
  MUX U4260 ( .IN0(n1853), .IN1(o[959]), .SEL(n2424), .F(\Data_Mem/n6832 ) );
  MUX U4261 ( .IN0(n1855), .IN1(o[958]), .SEL(n2424), .F(\Data_Mem/n6831 ) );
  MUX U4262 ( .IN0(n1856), .IN1(o[957]), .SEL(n2424), .F(\Data_Mem/n6830 ) );
  MUX U4263 ( .IN0(n1857), .IN1(o[956]), .SEL(n2424), .F(\Data_Mem/n6829 ) );
  MUX U4264 ( .IN0(n1858), .IN1(o[955]), .SEL(n2424), .F(\Data_Mem/n6828 ) );
  MUX U4265 ( .IN0(n1859), .IN1(o[954]), .SEL(n2424), .F(\Data_Mem/n6827 ) );
  MUX U4266 ( .IN0(n1860), .IN1(o[953]), .SEL(n2424), .F(\Data_Mem/n6826 ) );
  MUX U4267 ( .IN0(n1861), .IN1(o[952]), .SEL(n2424), .F(\Data_Mem/n6825 ) );
  ANDN U4268 ( .A(n2425), .B(n2426), .Z(n2424) );
  AND U4269 ( .A(n2427), .B(n2428), .Z(n2425) );
  OR U4270 ( .A(n1867), .B(n2429), .Z(n2428) );
  MUX U4271 ( .IN0(n1868), .IN1(o[951]), .SEL(n2430), .F(\Data_Mem/n6824 ) );
  MUX U4272 ( .IN0(n1870), .IN1(o[950]), .SEL(n2430), .F(\Data_Mem/n6823 ) );
  MUX U4273 ( .IN0(n1871), .IN1(o[949]), .SEL(n2430), .F(\Data_Mem/n6822 ) );
  MUX U4274 ( .IN0(n1872), .IN1(o[948]), .SEL(n2430), .F(\Data_Mem/n6821 ) );
  MUX U4275 ( .IN0(n1873), .IN1(o[947]), .SEL(n2430), .F(\Data_Mem/n6820 ) );
  IV U4276 ( .A(n2431), .Z(n2430) );
  MUX U4277 ( .IN0(o[946]), .IN1(n1875), .SEL(n2431), .F(\Data_Mem/n6819 ) );
  MUX U4278 ( .IN0(o[945]), .IN1(n1876), .SEL(n2431), .F(\Data_Mem/n6818 ) );
  MUX U4279 ( .IN0(o[944]), .IN1(n1877), .SEL(n2431), .F(\Data_Mem/n6817 ) );
  NAND U4280 ( .A(n2432), .B(n2433), .Z(n2431) );
  OR U4281 ( .A(n1880), .B(n2429), .Z(n2433) );
  ANDN U4282 ( .A(n2427), .B(n2426), .Z(n2432) );
  NANDN U4283 ( .B(n2429), .A(n1915), .Z(n2427) );
  MUX U4284 ( .IN0(n1883), .IN1(o[943]), .SEL(n2434), .F(\Data_Mem/n6816 ) );
  MUX U4285 ( .IN0(n1885), .IN1(o[942]), .SEL(n2434), .F(\Data_Mem/n6815 ) );
  MUX U4286 ( .IN0(n1886), .IN1(o[941]), .SEL(n2434), .F(\Data_Mem/n6814 ) );
  MUX U4287 ( .IN0(n1887), .IN1(o[940]), .SEL(n2434), .F(\Data_Mem/n6813 ) );
  MUX U4288 ( .IN0(n1888), .IN1(o[939]), .SEL(n2434), .F(\Data_Mem/n6812 ) );
  IV U4289 ( .A(n2435), .Z(n2434) );
  MUX U4290 ( .IN0(o[938]), .IN1(n1890), .SEL(n2435), .F(\Data_Mem/n6811 ) );
  MUX U4291 ( .IN0(o[937]), .IN1(n1891), .SEL(n2435), .F(\Data_Mem/n6810 ) );
  MUX U4292 ( .IN0(o[936]), .IN1(n1892), .SEL(n2435), .F(\Data_Mem/n6809 ) );
  NAND U4293 ( .A(n2436), .B(n2437), .Z(n2435) );
  OR U4294 ( .A(n1895), .B(n2429), .Z(n2437) );
  MUX U4295 ( .IN0(reg_target[7]), .IN1(o[935]), .SEL(n2438), .F(
        \Data_Mem/n6808 ) );
  MUX U4296 ( .IN0(reg_target[6]), .IN1(o[934]), .SEL(n2438), .F(
        \Data_Mem/n6807 ) );
  MUX U4297 ( .IN0(reg_target[5]), .IN1(o[933]), .SEL(n2438), .F(
        \Data_Mem/n6806 ) );
  MUX U4298 ( .IN0(reg_target[4]), .IN1(o[932]), .SEL(n2438), .F(
        \Data_Mem/n6805 ) );
  MUX U4299 ( .IN0(reg_target[3]), .IN1(o[931]), .SEL(n2438), .F(
        \Data_Mem/n6804 ) );
  IV U4300 ( .A(n2439), .Z(n2438) );
  MUX U4301 ( .IN0(o[930]), .IN1(reg_target[2]), .SEL(n2439), .F(
        \Data_Mem/n6803 ) );
  MUX U4302 ( .IN0(o[929]), .IN1(reg_target[1]), .SEL(n2439), .F(
        \Data_Mem/n6802 ) );
  MUX U4303 ( .IN0(o[928]), .IN1(reg_target[0]), .SEL(n2439), .F(
        \Data_Mem/n6801 ) );
  NAND U4304 ( .A(n2436), .B(n2440), .Z(n2439) );
  NANDN U4305 ( .B(n2429), .A(n1899), .Z(n2440) );
  ANDN U4306 ( .A(n2441), .B(n2426), .Z(n2436) );
  ANDN U4307 ( .A(n1902), .B(n2429), .Z(n2426) );
  NANDN U4308 ( .B(n2429), .A(n1924), .Z(n2441) );
  NAND U4309 ( .A(n2001), .B(n2351), .Z(n2429) );
  MUX U4310 ( .IN0(n1853), .IN1(o[991]), .SEL(n2442), .F(\Data_Mem/n6800 ) );
  MUX U4311 ( .IN0(n1855), .IN1(o[990]), .SEL(n2442), .F(\Data_Mem/n6799 ) );
  MUX U4312 ( .IN0(n1856), .IN1(o[989]), .SEL(n2442), .F(\Data_Mem/n6798 ) );
  MUX U4313 ( .IN0(n1857), .IN1(o[988]), .SEL(n2442), .F(\Data_Mem/n6797 ) );
  MUX U4314 ( .IN0(n1858), .IN1(o[987]), .SEL(n2442), .F(\Data_Mem/n6796 ) );
  MUX U4315 ( .IN0(n1859), .IN1(o[986]), .SEL(n2442), .F(\Data_Mem/n6795 ) );
  MUX U4316 ( .IN0(n1860), .IN1(o[985]), .SEL(n2442), .F(\Data_Mem/n6794 ) );
  MUX U4317 ( .IN0(n1861), .IN1(o[984]), .SEL(n2442), .F(\Data_Mem/n6793 ) );
  ANDN U4318 ( .A(n2443), .B(n2444), .Z(n2442) );
  AND U4319 ( .A(n2445), .B(n2446), .Z(n2443) );
  OR U4320 ( .A(n1867), .B(n2447), .Z(n2446) );
  MUX U4321 ( .IN0(n1868), .IN1(o[983]), .SEL(n2448), .F(\Data_Mem/n6792 ) );
  MUX U4322 ( .IN0(n1870), .IN1(o[982]), .SEL(n2448), .F(\Data_Mem/n6791 ) );
  MUX U4323 ( .IN0(n1871), .IN1(o[981]), .SEL(n2448), .F(\Data_Mem/n6790 ) );
  MUX U4324 ( .IN0(n1872), .IN1(o[980]), .SEL(n2448), .F(\Data_Mem/n6789 ) );
  MUX U4325 ( .IN0(n1873), .IN1(o[979]), .SEL(n2448), .F(\Data_Mem/n6788 ) );
  IV U4326 ( .A(n2449), .Z(n2448) );
  MUX U4327 ( .IN0(o[978]), .IN1(n1875), .SEL(n2449), .F(\Data_Mem/n6787 ) );
  MUX U4328 ( .IN0(o[977]), .IN1(n1876), .SEL(n2449), .F(\Data_Mem/n6786 ) );
  MUX U4329 ( .IN0(o[976]), .IN1(n1877), .SEL(n2449), .F(\Data_Mem/n6785 ) );
  NAND U4330 ( .A(n2450), .B(n2451), .Z(n2449) );
  OR U4331 ( .A(n1880), .B(n2447), .Z(n2451) );
  ANDN U4332 ( .A(n2445), .B(n2444), .Z(n2450) );
  NANDN U4333 ( .B(n2447), .A(n1915), .Z(n2445) );
  MUX U4334 ( .IN0(n1883), .IN1(o[975]), .SEL(n2452), .F(\Data_Mem/n6784 ) );
  MUX U4335 ( .IN0(n1885), .IN1(o[974]), .SEL(n2452), .F(\Data_Mem/n6783 ) );
  MUX U4336 ( .IN0(n1886), .IN1(o[973]), .SEL(n2452), .F(\Data_Mem/n6782 ) );
  MUX U4337 ( .IN0(n1887), .IN1(o[972]), .SEL(n2452), .F(\Data_Mem/n6781 ) );
  MUX U4338 ( .IN0(n1888), .IN1(o[971]), .SEL(n2452), .F(\Data_Mem/n6780 ) );
  IV U4339 ( .A(n2453), .Z(n2452) );
  MUX U4340 ( .IN0(o[970]), .IN1(n1890), .SEL(n2453), .F(\Data_Mem/n6779 ) );
  MUX U4341 ( .IN0(o[969]), .IN1(n1891), .SEL(n2453), .F(\Data_Mem/n6778 ) );
  MUX U4342 ( .IN0(o[968]), .IN1(n1892), .SEL(n2453), .F(\Data_Mem/n6777 ) );
  NAND U4343 ( .A(n2454), .B(n2455), .Z(n2453) );
  OR U4344 ( .A(n1895), .B(n2447), .Z(n2455) );
  MUX U4345 ( .IN0(reg_target[7]), .IN1(o[967]), .SEL(n2456), .F(
        \Data_Mem/n6776 ) );
  MUX U4346 ( .IN0(reg_target[6]), .IN1(o[966]), .SEL(n2456), .F(
        \Data_Mem/n6775 ) );
  MUX U4347 ( .IN0(reg_target[5]), .IN1(o[965]), .SEL(n2456), .F(
        \Data_Mem/n6774 ) );
  MUX U4348 ( .IN0(reg_target[4]), .IN1(o[964]), .SEL(n2456), .F(
        \Data_Mem/n6773 ) );
  MUX U4349 ( .IN0(reg_target[3]), .IN1(o[963]), .SEL(n2456), .F(
        \Data_Mem/n6772 ) );
  IV U4350 ( .A(n2457), .Z(n2456) );
  MUX U4351 ( .IN0(o[962]), .IN1(reg_target[2]), .SEL(n2457), .F(
        \Data_Mem/n6771 ) );
  MUX U4352 ( .IN0(o[961]), .IN1(reg_target[1]), .SEL(n2457), .F(
        \Data_Mem/n6770 ) );
  MUX U4353 ( .IN0(o[960]), .IN1(reg_target[0]), .SEL(n2457), .F(
        \Data_Mem/n6769 ) );
  NAND U4354 ( .A(n2454), .B(n2458), .Z(n2457) );
  NANDN U4355 ( .B(n2447), .A(n1899), .Z(n2458) );
  ANDN U4356 ( .A(n2459), .B(n2444), .Z(n2454) );
  ANDN U4357 ( .A(n1902), .B(n2447), .Z(n2444) );
  NANDN U4358 ( .B(n2447), .A(n1924), .Z(n2459) );
  NAND U4359 ( .A(n2020), .B(n2351), .Z(n2447) );
  MUX U4360 ( .IN0(n1853), .IN1(o[1023]), .SEL(n2460), .F(\Data_Mem/n6768 ) );
  MUX U4361 ( .IN0(n1855), .IN1(o[1022]), .SEL(n2460), .F(\Data_Mem/n6767 ) );
  MUX U4362 ( .IN0(n1856), .IN1(o[1021]), .SEL(n2460), .F(\Data_Mem/n6766 ) );
  MUX U4363 ( .IN0(n1857), .IN1(o[1020]), .SEL(n2460), .F(\Data_Mem/n6765 ) );
  MUX U4364 ( .IN0(n1858), .IN1(o[1019]), .SEL(n2460), .F(\Data_Mem/n6764 ) );
  MUX U4365 ( .IN0(n1859), .IN1(o[1018]), .SEL(n2460), .F(\Data_Mem/n6763 ) );
  MUX U4366 ( .IN0(n1860), .IN1(o[1017]), .SEL(n2460), .F(\Data_Mem/n6762 ) );
  MUX U4367 ( .IN0(n1861), .IN1(o[1016]), .SEL(n2460), .F(\Data_Mem/n6761 ) );
  ANDN U4368 ( .A(n2461), .B(n2462), .Z(n2460) );
  AND U4369 ( .A(n2463), .B(n2464), .Z(n2461) );
  OR U4370 ( .A(n1867), .B(n2465), .Z(n2464) );
  MUX U4371 ( .IN0(n1868), .IN1(o[1015]), .SEL(n2466), .F(\Data_Mem/n6760 ) );
  MUX U4372 ( .IN0(n1870), .IN1(o[1014]), .SEL(n2466), .F(\Data_Mem/n6759 ) );
  MUX U4373 ( .IN0(n1871), .IN1(o[1013]), .SEL(n2466), .F(\Data_Mem/n6758 ) );
  MUX U4374 ( .IN0(n1872), .IN1(o[1012]), .SEL(n2466), .F(\Data_Mem/n6757 ) );
  MUX U4375 ( .IN0(n1873), .IN1(o[1011]), .SEL(n2466), .F(\Data_Mem/n6756 ) );
  IV U4376 ( .A(n2467), .Z(n2466) );
  MUX U4377 ( .IN0(o[1010]), .IN1(n1875), .SEL(n2467), .F(\Data_Mem/n6755 ) );
  MUX U4378 ( .IN0(o[1009]), .IN1(n1876), .SEL(n2467), .F(\Data_Mem/n6754 ) );
  MUX U4379 ( .IN0(o[1008]), .IN1(n1877), .SEL(n2467), .F(\Data_Mem/n6753 ) );
  NAND U4380 ( .A(n2468), .B(n2469), .Z(n2467) );
  OR U4381 ( .A(n1880), .B(n2465), .Z(n2469) );
  ANDN U4382 ( .A(n2463), .B(n2462), .Z(n2468) );
  NANDN U4383 ( .B(n2465), .A(n1915), .Z(n2463) );
  MUX U4384 ( .IN0(n1883), .IN1(o[1007]), .SEL(n2470), .F(\Data_Mem/n6752 ) );
  MUX U4385 ( .IN0(n1885), .IN1(o[1006]), .SEL(n2470), .F(\Data_Mem/n6751 ) );
  MUX U4386 ( .IN0(n1886), .IN1(o[1005]), .SEL(n2470), .F(\Data_Mem/n6750 ) );
  MUX U4387 ( .IN0(n1887), .IN1(o[1004]), .SEL(n2470), .F(\Data_Mem/n6749 ) );
  MUX U4388 ( .IN0(n1888), .IN1(o[1003]), .SEL(n2470), .F(\Data_Mem/n6748 ) );
  IV U4389 ( .A(n2471), .Z(n2470) );
  MUX U4390 ( .IN0(o[1002]), .IN1(n1890), .SEL(n2471), .F(\Data_Mem/n6747 ) );
  MUX U4391 ( .IN0(o[1001]), .IN1(n1891), .SEL(n2471), .F(\Data_Mem/n6746 ) );
  MUX U4392 ( .IN0(o[1000]), .IN1(n1892), .SEL(n2471), .F(\Data_Mem/n6745 ) );
  NAND U4393 ( .A(n2472), .B(n2473), .Z(n2471) );
  OR U4394 ( .A(n1895), .B(n2465), .Z(n2473) );
  MUX U4395 ( .IN0(reg_target[7]), .IN1(o[999]), .SEL(n2474), .F(
        \Data_Mem/n6744 ) );
  MUX U4396 ( .IN0(reg_target[6]), .IN1(o[998]), .SEL(n2474), .F(
        \Data_Mem/n6743 ) );
  MUX U4397 ( .IN0(reg_target[5]), .IN1(o[997]), .SEL(n2474), .F(
        \Data_Mem/n6742 ) );
  MUX U4398 ( .IN0(reg_target[4]), .IN1(o[996]), .SEL(n2474), .F(
        \Data_Mem/n6741 ) );
  MUX U4399 ( .IN0(reg_target[3]), .IN1(o[995]), .SEL(n2474), .F(
        \Data_Mem/n6740 ) );
  IV U4400 ( .A(n2475), .Z(n2474) );
  MUX U4401 ( .IN0(o[994]), .IN1(reg_target[2]), .SEL(n2475), .F(
        \Data_Mem/n6739 ) );
  MUX U4402 ( .IN0(o[993]), .IN1(reg_target[1]), .SEL(n2475), .F(
        \Data_Mem/n6738 ) );
  MUX U4403 ( .IN0(o[992]), .IN1(reg_target[0]), .SEL(n2475), .F(
        \Data_Mem/n6737 ) );
  NAND U4404 ( .A(n2472), .B(n2476), .Z(n2475) );
  NANDN U4405 ( .B(n2465), .A(n1899), .Z(n2476) );
  ANDN U4406 ( .A(n2477), .B(n2462), .Z(n2472) );
  ANDN U4407 ( .A(n1902), .B(n2465), .Z(n2462) );
  NANDN U4408 ( .B(n2465), .A(n1924), .Z(n2477) );
  NAND U4409 ( .A(n2351), .B(n2039), .Z(n2465) );
  AND U4410 ( .A(n2478), .B(n485), .Z(n2351) );
  MUX U4411 ( .IN0(n1853), .IN1(o[1055]), .SEL(n2479), .F(\Data_Mem/n6736 ) );
  MUX U4412 ( .IN0(n1855), .IN1(o[1054]), .SEL(n2479), .F(\Data_Mem/n6735 ) );
  MUX U4413 ( .IN0(n1856), .IN1(o[1053]), .SEL(n2479), .F(\Data_Mem/n6734 ) );
  MUX U4414 ( .IN0(n1857), .IN1(o[1052]), .SEL(n2479), .F(\Data_Mem/n6733 ) );
  MUX U4415 ( .IN0(n1858), .IN1(o[1051]), .SEL(n2479), .F(\Data_Mem/n6732 ) );
  MUX U4416 ( .IN0(n1859), .IN1(o[1050]), .SEL(n2479), .F(\Data_Mem/n6731 ) );
  MUX U4417 ( .IN0(n1860), .IN1(o[1049]), .SEL(n2479), .F(\Data_Mem/n6730 ) );
  MUX U4418 ( .IN0(n1861), .IN1(o[1048]), .SEL(n2479), .F(\Data_Mem/n6729 ) );
  ANDN U4419 ( .A(n2480), .B(n2481), .Z(n2479) );
  AND U4420 ( .A(n2482), .B(n2483), .Z(n2480) );
  OR U4421 ( .A(n1867), .B(n2484), .Z(n2483) );
  MUX U4422 ( .IN0(n1868), .IN1(o[1047]), .SEL(n2485), .F(\Data_Mem/n6728 ) );
  MUX U4423 ( .IN0(n1870), .IN1(o[1046]), .SEL(n2485), .F(\Data_Mem/n6727 ) );
  MUX U4424 ( .IN0(n1871), .IN1(o[1045]), .SEL(n2485), .F(\Data_Mem/n6726 ) );
  MUX U4425 ( .IN0(n1872), .IN1(o[1044]), .SEL(n2485), .F(\Data_Mem/n6725 ) );
  MUX U4426 ( .IN0(n1873), .IN1(o[1043]), .SEL(n2485), .F(\Data_Mem/n6724 ) );
  IV U4427 ( .A(n2486), .Z(n2485) );
  MUX U4428 ( .IN0(o[1042]), .IN1(n1875), .SEL(n2486), .F(\Data_Mem/n6723 ) );
  MUX U4429 ( .IN0(o[1041]), .IN1(n1876), .SEL(n2486), .F(\Data_Mem/n6722 ) );
  MUX U4430 ( .IN0(o[1040]), .IN1(n1877), .SEL(n2486), .F(\Data_Mem/n6721 ) );
  NAND U4431 ( .A(n2487), .B(n2488), .Z(n2486) );
  OR U4432 ( .A(n1880), .B(n2484), .Z(n2488) );
  ANDN U4433 ( .A(n2482), .B(n2481), .Z(n2487) );
  NANDN U4434 ( .B(n2484), .A(n1915), .Z(n2482) );
  MUX U4435 ( .IN0(n1883), .IN1(o[1039]), .SEL(n2489), .F(\Data_Mem/n6720 ) );
  MUX U4436 ( .IN0(n1885), .IN1(o[1038]), .SEL(n2489), .F(\Data_Mem/n6719 ) );
  MUX U4437 ( .IN0(n1886), .IN1(o[1037]), .SEL(n2489), .F(\Data_Mem/n6718 ) );
  MUX U4438 ( .IN0(n1887), .IN1(o[1036]), .SEL(n2489), .F(\Data_Mem/n6717 ) );
  MUX U4439 ( .IN0(n1888), .IN1(o[1035]), .SEL(n2489), .F(\Data_Mem/n6716 ) );
  IV U4440 ( .A(n2490), .Z(n2489) );
  MUX U4441 ( .IN0(o[1034]), .IN1(n1890), .SEL(n2490), .F(\Data_Mem/n6715 ) );
  MUX U4442 ( .IN0(o[1033]), .IN1(n1891), .SEL(n2490), .F(\Data_Mem/n6714 ) );
  MUX U4443 ( .IN0(o[1032]), .IN1(n1892), .SEL(n2490), .F(\Data_Mem/n6713 ) );
  NAND U4444 ( .A(n2491), .B(n2492), .Z(n2490) );
  OR U4445 ( .A(n1895), .B(n2484), .Z(n2492) );
  MUX U4446 ( .IN0(reg_target[7]), .IN1(o[1031]), .SEL(n2493), .F(
        \Data_Mem/n6712 ) );
  MUX U4447 ( .IN0(reg_target[6]), .IN1(o[1030]), .SEL(n2493), .F(
        \Data_Mem/n6711 ) );
  MUX U4448 ( .IN0(reg_target[5]), .IN1(o[1029]), .SEL(n2493), .F(
        \Data_Mem/n6710 ) );
  MUX U4449 ( .IN0(reg_target[4]), .IN1(o[1028]), .SEL(n2493), .F(
        \Data_Mem/n6709 ) );
  MUX U4450 ( .IN0(reg_target[3]), .IN1(o[1027]), .SEL(n2493), .F(
        \Data_Mem/n6708 ) );
  IV U4451 ( .A(n2494), .Z(n2493) );
  MUX U4452 ( .IN0(o[1026]), .IN1(reg_target[2]), .SEL(n2494), .F(
        \Data_Mem/n6707 ) );
  MUX U4453 ( .IN0(o[1025]), .IN1(reg_target[1]), .SEL(n2494), .F(
        \Data_Mem/n6706 ) );
  MUX U4454 ( .IN0(o[1024]), .IN1(reg_target[0]), .SEL(n2494), .F(
        \Data_Mem/n6705 ) );
  NAND U4455 ( .A(n2491), .B(n2495), .Z(n2494) );
  NANDN U4456 ( .B(n2484), .A(n1899), .Z(n2495) );
  ANDN U4457 ( .A(n2496), .B(n2481), .Z(n2491) );
  ANDN U4458 ( .A(n1902), .B(n2484), .Z(n2481) );
  NANDN U4459 ( .B(n2484), .A(n1924), .Z(n2496) );
  NAND U4460 ( .A(n1903), .B(n2497), .Z(n2484) );
  MUX U4461 ( .IN0(n1853), .IN1(o[1087]), .SEL(n2498), .F(\Data_Mem/n6704 ) );
  MUX U4462 ( .IN0(n1855), .IN1(o[1086]), .SEL(n2498), .F(\Data_Mem/n6703 ) );
  MUX U4463 ( .IN0(n1856), .IN1(o[1085]), .SEL(n2498), .F(\Data_Mem/n6702 ) );
  MUX U4464 ( .IN0(n1857), .IN1(o[1084]), .SEL(n2498), .F(\Data_Mem/n6701 ) );
  MUX U4465 ( .IN0(n1858), .IN1(o[1083]), .SEL(n2498), .F(\Data_Mem/n6700 ) );
  MUX U4466 ( .IN0(n1859), .IN1(o[1082]), .SEL(n2498), .F(\Data_Mem/n6699 ) );
  MUX U4467 ( .IN0(n1860), .IN1(o[1081]), .SEL(n2498), .F(\Data_Mem/n6698 ) );
  MUX U4468 ( .IN0(n1861), .IN1(o[1080]), .SEL(n2498), .F(\Data_Mem/n6697 ) );
  ANDN U4469 ( .A(n2499), .B(n2500), .Z(n2498) );
  AND U4470 ( .A(n2501), .B(n2502), .Z(n2499) );
  OR U4471 ( .A(n1867), .B(n2503), .Z(n2502) );
  MUX U4472 ( .IN0(n1868), .IN1(o[1079]), .SEL(n2504), .F(\Data_Mem/n6696 ) );
  MUX U4473 ( .IN0(n1870), .IN1(o[1078]), .SEL(n2504), .F(\Data_Mem/n6695 ) );
  MUX U4474 ( .IN0(n1871), .IN1(o[1077]), .SEL(n2504), .F(\Data_Mem/n6694 ) );
  MUX U4475 ( .IN0(n1872), .IN1(o[1076]), .SEL(n2504), .F(\Data_Mem/n6693 ) );
  MUX U4476 ( .IN0(n1873), .IN1(o[1075]), .SEL(n2504), .F(\Data_Mem/n6692 ) );
  IV U4477 ( .A(n2505), .Z(n2504) );
  MUX U4478 ( .IN0(o[1074]), .IN1(n1875), .SEL(n2505), .F(\Data_Mem/n6691 ) );
  MUX U4479 ( .IN0(o[1073]), .IN1(n1876), .SEL(n2505), .F(\Data_Mem/n6690 ) );
  MUX U4480 ( .IN0(o[1072]), .IN1(n1877), .SEL(n2505), .F(\Data_Mem/n6689 ) );
  NAND U4481 ( .A(n2506), .B(n2507), .Z(n2505) );
  OR U4482 ( .A(n1880), .B(n2503), .Z(n2507) );
  ANDN U4483 ( .A(n2501), .B(n2500), .Z(n2506) );
  NANDN U4484 ( .B(n2503), .A(n1915), .Z(n2501) );
  MUX U4485 ( .IN0(n1883), .IN1(o[1071]), .SEL(n2508), .F(\Data_Mem/n6688 ) );
  MUX U4486 ( .IN0(n1885), .IN1(o[1070]), .SEL(n2508), .F(\Data_Mem/n6687 ) );
  MUX U4487 ( .IN0(n1886), .IN1(o[1069]), .SEL(n2508), .F(\Data_Mem/n6686 ) );
  MUX U4488 ( .IN0(n1887), .IN1(o[1068]), .SEL(n2508), .F(\Data_Mem/n6685 ) );
  MUX U4489 ( .IN0(n1888), .IN1(o[1067]), .SEL(n2508), .F(\Data_Mem/n6684 ) );
  IV U4490 ( .A(n2509), .Z(n2508) );
  MUX U4491 ( .IN0(o[1066]), .IN1(n1890), .SEL(n2509), .F(\Data_Mem/n6683 ) );
  MUX U4492 ( .IN0(o[1065]), .IN1(n1891), .SEL(n2509), .F(\Data_Mem/n6682 ) );
  MUX U4493 ( .IN0(o[1064]), .IN1(n1892), .SEL(n2509), .F(\Data_Mem/n6681 ) );
  NAND U4494 ( .A(n2510), .B(n2511), .Z(n2509) );
  OR U4495 ( .A(n1895), .B(n2503), .Z(n2511) );
  MUX U4496 ( .IN0(reg_target[7]), .IN1(o[1063]), .SEL(n2512), .F(
        \Data_Mem/n6680 ) );
  MUX U4497 ( .IN0(reg_target[6]), .IN1(o[1062]), .SEL(n2512), .F(
        \Data_Mem/n6679 ) );
  MUX U4498 ( .IN0(reg_target[5]), .IN1(o[1061]), .SEL(n2512), .F(
        \Data_Mem/n6678 ) );
  MUX U4499 ( .IN0(reg_target[4]), .IN1(o[1060]), .SEL(n2512), .F(
        \Data_Mem/n6677 ) );
  MUX U4500 ( .IN0(reg_target[3]), .IN1(o[1059]), .SEL(n2512), .F(
        \Data_Mem/n6676 ) );
  IV U4501 ( .A(n2513), .Z(n2512) );
  MUX U4502 ( .IN0(o[1058]), .IN1(reg_target[2]), .SEL(n2513), .F(
        \Data_Mem/n6675 ) );
  MUX U4503 ( .IN0(o[1057]), .IN1(reg_target[1]), .SEL(n2513), .F(
        \Data_Mem/n6674 ) );
  MUX U4504 ( .IN0(o[1056]), .IN1(reg_target[0]), .SEL(n2513), .F(
        \Data_Mem/n6673 ) );
  NAND U4505 ( .A(n2510), .B(n2514), .Z(n2513) );
  NANDN U4506 ( .B(n2503), .A(n1899), .Z(n2514) );
  ANDN U4507 ( .A(n2515), .B(n2500), .Z(n2510) );
  ANDN U4508 ( .A(n1902), .B(n2503), .Z(n2500) );
  NANDN U4509 ( .B(n2503), .A(n1924), .Z(n2515) );
  NAND U4510 ( .A(n1925), .B(n2497), .Z(n2503) );
  MUX U4511 ( .IN0(n1853), .IN1(o[1119]), .SEL(n2516), .F(\Data_Mem/n6672 ) );
  MUX U4512 ( .IN0(n1855), .IN1(o[1118]), .SEL(n2516), .F(\Data_Mem/n6671 ) );
  MUX U4513 ( .IN0(n1856), .IN1(o[1117]), .SEL(n2516), .F(\Data_Mem/n6670 ) );
  MUX U4514 ( .IN0(n1857), .IN1(o[1116]), .SEL(n2516), .F(\Data_Mem/n6669 ) );
  MUX U4515 ( .IN0(n1858), .IN1(o[1115]), .SEL(n2516), .F(\Data_Mem/n6668 ) );
  MUX U4516 ( .IN0(n1859), .IN1(o[1114]), .SEL(n2516), .F(\Data_Mem/n6667 ) );
  MUX U4517 ( .IN0(n1860), .IN1(o[1113]), .SEL(n2516), .F(\Data_Mem/n6666 ) );
  MUX U4518 ( .IN0(n1861), .IN1(o[1112]), .SEL(n2516), .F(\Data_Mem/n6665 ) );
  ANDN U4519 ( .A(n2517), .B(n2518), .Z(n2516) );
  AND U4520 ( .A(n2519), .B(n2520), .Z(n2517) );
  OR U4521 ( .A(n1867), .B(n2521), .Z(n2520) );
  MUX U4522 ( .IN0(n1868), .IN1(o[1111]), .SEL(n2522), .F(\Data_Mem/n6664 ) );
  MUX U4523 ( .IN0(n1870), .IN1(o[1110]), .SEL(n2522), .F(\Data_Mem/n6663 ) );
  MUX U4524 ( .IN0(n1871), .IN1(o[1109]), .SEL(n2522), .F(\Data_Mem/n6662 ) );
  MUX U4525 ( .IN0(n1872), .IN1(o[1108]), .SEL(n2522), .F(\Data_Mem/n6661 ) );
  MUX U4526 ( .IN0(n1873), .IN1(o[1107]), .SEL(n2522), .F(\Data_Mem/n6660 ) );
  IV U4527 ( .A(n2523), .Z(n2522) );
  MUX U4528 ( .IN0(o[1106]), .IN1(n1875), .SEL(n2523), .F(\Data_Mem/n6659 ) );
  MUX U4529 ( .IN0(o[1105]), .IN1(n1876), .SEL(n2523), .F(\Data_Mem/n6658 ) );
  MUX U4530 ( .IN0(o[1104]), .IN1(n1877), .SEL(n2523), .F(\Data_Mem/n6657 ) );
  NAND U4531 ( .A(n2524), .B(n2525), .Z(n2523) );
  OR U4532 ( .A(n1880), .B(n2521), .Z(n2525) );
  ANDN U4533 ( .A(n2519), .B(n2518), .Z(n2524) );
  NANDN U4534 ( .B(n2521), .A(n1915), .Z(n2519) );
  MUX U4535 ( .IN0(n1883), .IN1(o[1103]), .SEL(n2526), .F(\Data_Mem/n6656 ) );
  MUX U4536 ( .IN0(n1885), .IN1(o[1102]), .SEL(n2526), .F(\Data_Mem/n6655 ) );
  MUX U4537 ( .IN0(n1886), .IN1(o[1101]), .SEL(n2526), .F(\Data_Mem/n6654 ) );
  MUX U4538 ( .IN0(n1887), .IN1(o[1100]), .SEL(n2526), .F(\Data_Mem/n6653 ) );
  MUX U4539 ( .IN0(n1888), .IN1(o[1099]), .SEL(n2526), .F(\Data_Mem/n6652 ) );
  IV U4540 ( .A(n2527), .Z(n2526) );
  MUX U4541 ( .IN0(o[1098]), .IN1(n1890), .SEL(n2527), .F(\Data_Mem/n6651 ) );
  MUX U4542 ( .IN0(o[1097]), .IN1(n1891), .SEL(n2527), .F(\Data_Mem/n6650 ) );
  MUX U4543 ( .IN0(o[1096]), .IN1(n1892), .SEL(n2527), .F(\Data_Mem/n6649 ) );
  NAND U4544 ( .A(n2528), .B(n2529), .Z(n2527) );
  OR U4545 ( .A(n1895), .B(n2521), .Z(n2529) );
  MUX U4546 ( .IN0(reg_target[7]), .IN1(o[1095]), .SEL(n2530), .F(
        \Data_Mem/n6648 ) );
  MUX U4547 ( .IN0(reg_target[6]), .IN1(o[1094]), .SEL(n2530), .F(
        \Data_Mem/n6647 ) );
  MUX U4548 ( .IN0(reg_target[5]), .IN1(o[1093]), .SEL(n2530), .F(
        \Data_Mem/n6646 ) );
  MUX U4549 ( .IN0(reg_target[4]), .IN1(o[1092]), .SEL(n2530), .F(
        \Data_Mem/n6645 ) );
  MUX U4550 ( .IN0(reg_target[3]), .IN1(o[1091]), .SEL(n2530), .F(
        \Data_Mem/n6644 ) );
  IV U4551 ( .A(n2531), .Z(n2530) );
  MUX U4552 ( .IN0(o[1090]), .IN1(reg_target[2]), .SEL(n2531), .F(
        \Data_Mem/n6643 ) );
  MUX U4553 ( .IN0(o[1089]), .IN1(reg_target[1]), .SEL(n2531), .F(
        \Data_Mem/n6642 ) );
  MUX U4554 ( .IN0(o[1088]), .IN1(reg_target[0]), .SEL(n2531), .F(
        \Data_Mem/n6641 ) );
  NAND U4555 ( .A(n2528), .B(n2532), .Z(n2531) );
  NANDN U4556 ( .B(n2521), .A(n1899), .Z(n2532) );
  ANDN U4557 ( .A(n2533), .B(n2518), .Z(n2528) );
  ANDN U4558 ( .A(n1902), .B(n2521), .Z(n2518) );
  NANDN U4559 ( .B(n2521), .A(n1924), .Z(n2533) );
  NAND U4560 ( .A(n1944), .B(n2497), .Z(n2521) );
  MUX U4561 ( .IN0(n1853), .IN1(o[1151]), .SEL(n2534), .F(\Data_Mem/n6640 ) );
  MUX U4562 ( .IN0(n1855), .IN1(o[1150]), .SEL(n2534), .F(\Data_Mem/n6639 ) );
  MUX U4563 ( .IN0(n1856), .IN1(o[1149]), .SEL(n2534), .F(\Data_Mem/n6638 ) );
  MUX U4564 ( .IN0(n1857), .IN1(o[1148]), .SEL(n2534), .F(\Data_Mem/n6637 ) );
  MUX U4565 ( .IN0(n1858), .IN1(o[1147]), .SEL(n2534), .F(\Data_Mem/n6636 ) );
  MUX U4566 ( .IN0(n1859), .IN1(o[1146]), .SEL(n2534), .F(\Data_Mem/n6635 ) );
  MUX U4567 ( .IN0(n1860), .IN1(o[1145]), .SEL(n2534), .F(\Data_Mem/n6634 ) );
  MUX U4568 ( .IN0(n1861), .IN1(o[1144]), .SEL(n2534), .F(\Data_Mem/n6633 ) );
  ANDN U4569 ( .A(n2535), .B(n2536), .Z(n2534) );
  AND U4570 ( .A(n2537), .B(n2538), .Z(n2535) );
  OR U4571 ( .A(n1867), .B(n2539), .Z(n2538) );
  MUX U4572 ( .IN0(n1868), .IN1(o[1143]), .SEL(n2540), .F(\Data_Mem/n6632 ) );
  MUX U4573 ( .IN0(n1870), .IN1(o[1142]), .SEL(n2540), .F(\Data_Mem/n6631 ) );
  MUX U4574 ( .IN0(n1871), .IN1(o[1141]), .SEL(n2540), .F(\Data_Mem/n6630 ) );
  MUX U4575 ( .IN0(n1872), .IN1(o[1140]), .SEL(n2540), .F(\Data_Mem/n6629 ) );
  MUX U4576 ( .IN0(n1873), .IN1(o[1139]), .SEL(n2540), .F(\Data_Mem/n6628 ) );
  IV U4577 ( .A(n2541), .Z(n2540) );
  MUX U4578 ( .IN0(o[1138]), .IN1(n1875), .SEL(n2541), .F(\Data_Mem/n6627 ) );
  MUX U4579 ( .IN0(o[1137]), .IN1(n1876), .SEL(n2541), .F(\Data_Mem/n6626 ) );
  MUX U4580 ( .IN0(o[1136]), .IN1(n1877), .SEL(n2541), .F(\Data_Mem/n6625 ) );
  NAND U4581 ( .A(n2542), .B(n2543), .Z(n2541) );
  OR U4582 ( .A(n1880), .B(n2539), .Z(n2543) );
  ANDN U4583 ( .A(n2537), .B(n2536), .Z(n2542) );
  NANDN U4584 ( .B(n2539), .A(n1915), .Z(n2537) );
  MUX U4585 ( .IN0(n1883), .IN1(o[1135]), .SEL(n2544), .F(\Data_Mem/n6624 ) );
  MUX U4586 ( .IN0(n1885), .IN1(o[1134]), .SEL(n2544), .F(\Data_Mem/n6623 ) );
  MUX U4587 ( .IN0(n1886), .IN1(o[1133]), .SEL(n2544), .F(\Data_Mem/n6622 ) );
  MUX U4588 ( .IN0(n1887), .IN1(o[1132]), .SEL(n2544), .F(\Data_Mem/n6621 ) );
  MUX U4589 ( .IN0(n1888), .IN1(o[1131]), .SEL(n2544), .F(\Data_Mem/n6620 ) );
  IV U4590 ( .A(n2545), .Z(n2544) );
  MUX U4591 ( .IN0(o[1130]), .IN1(n1890), .SEL(n2545), .F(\Data_Mem/n6619 ) );
  MUX U4592 ( .IN0(o[1129]), .IN1(n1891), .SEL(n2545), .F(\Data_Mem/n6618 ) );
  MUX U4593 ( .IN0(o[1128]), .IN1(n1892), .SEL(n2545), .F(\Data_Mem/n6617 ) );
  NAND U4594 ( .A(n2546), .B(n2547), .Z(n2545) );
  OR U4595 ( .A(n1895), .B(n2539), .Z(n2547) );
  MUX U4596 ( .IN0(reg_target[7]), .IN1(o[1127]), .SEL(n2548), .F(
        \Data_Mem/n6616 ) );
  MUX U4597 ( .IN0(reg_target[6]), .IN1(o[1126]), .SEL(n2548), .F(
        \Data_Mem/n6615 ) );
  MUX U4598 ( .IN0(reg_target[5]), .IN1(o[1125]), .SEL(n2548), .F(
        \Data_Mem/n6614 ) );
  MUX U4599 ( .IN0(reg_target[4]), .IN1(o[1124]), .SEL(n2548), .F(
        \Data_Mem/n6613 ) );
  MUX U4600 ( .IN0(reg_target[3]), .IN1(o[1123]), .SEL(n2548), .F(
        \Data_Mem/n6612 ) );
  IV U4601 ( .A(n2549), .Z(n2548) );
  MUX U4602 ( .IN0(o[1122]), .IN1(reg_target[2]), .SEL(n2549), .F(
        \Data_Mem/n6611 ) );
  MUX U4603 ( .IN0(o[1121]), .IN1(reg_target[1]), .SEL(n2549), .F(
        \Data_Mem/n6610 ) );
  MUX U4604 ( .IN0(o[1120]), .IN1(reg_target[0]), .SEL(n2549), .F(
        \Data_Mem/n6609 ) );
  NAND U4605 ( .A(n2546), .B(n2550), .Z(n2549) );
  NANDN U4606 ( .B(n2539), .A(n1899), .Z(n2550) );
  ANDN U4607 ( .A(n2551), .B(n2536), .Z(n2546) );
  ANDN U4608 ( .A(n1902), .B(n2539), .Z(n2536) );
  NANDN U4609 ( .B(n2539), .A(n1924), .Z(n2551) );
  NAND U4610 ( .A(n1963), .B(n2497), .Z(n2539) );
  MUX U4611 ( .IN0(n1853), .IN1(o[1183]), .SEL(n2552), .F(\Data_Mem/n6608 ) );
  MUX U4612 ( .IN0(n1855), .IN1(o[1182]), .SEL(n2552), .F(\Data_Mem/n6607 ) );
  MUX U4613 ( .IN0(n1856), .IN1(o[1181]), .SEL(n2552), .F(\Data_Mem/n6606 ) );
  MUX U4614 ( .IN0(n1857), .IN1(o[1180]), .SEL(n2552), .F(\Data_Mem/n6605 ) );
  MUX U4615 ( .IN0(n1858), .IN1(o[1179]), .SEL(n2552), .F(\Data_Mem/n6604 ) );
  MUX U4616 ( .IN0(n1859), .IN1(o[1178]), .SEL(n2552), .F(\Data_Mem/n6603 ) );
  MUX U4617 ( .IN0(n1860), .IN1(o[1177]), .SEL(n2552), .F(\Data_Mem/n6602 ) );
  MUX U4618 ( .IN0(n1861), .IN1(o[1176]), .SEL(n2552), .F(\Data_Mem/n6601 ) );
  ANDN U4619 ( .A(n2553), .B(n2554), .Z(n2552) );
  AND U4620 ( .A(n2555), .B(n2556), .Z(n2553) );
  OR U4621 ( .A(n1867), .B(n2557), .Z(n2556) );
  MUX U4622 ( .IN0(n1868), .IN1(o[1175]), .SEL(n2558), .F(\Data_Mem/n6600 ) );
  MUX U4623 ( .IN0(n1870), .IN1(o[1174]), .SEL(n2558), .F(\Data_Mem/n6599 ) );
  MUX U4624 ( .IN0(n1871), .IN1(o[1173]), .SEL(n2558), .F(\Data_Mem/n6598 ) );
  MUX U4625 ( .IN0(n1872), .IN1(o[1172]), .SEL(n2558), .F(\Data_Mem/n6597 ) );
  MUX U4626 ( .IN0(n1873), .IN1(o[1171]), .SEL(n2558), .F(\Data_Mem/n6596 ) );
  IV U4627 ( .A(n2559), .Z(n2558) );
  MUX U4628 ( .IN0(o[1170]), .IN1(n1875), .SEL(n2559), .F(\Data_Mem/n6595 ) );
  MUX U4629 ( .IN0(o[1169]), .IN1(n1876), .SEL(n2559), .F(\Data_Mem/n6594 ) );
  MUX U4630 ( .IN0(o[1168]), .IN1(n1877), .SEL(n2559), .F(\Data_Mem/n6593 ) );
  NAND U4631 ( .A(n2560), .B(n2561), .Z(n2559) );
  OR U4632 ( .A(n1880), .B(n2557), .Z(n2561) );
  ANDN U4633 ( .A(n2555), .B(n2554), .Z(n2560) );
  NANDN U4634 ( .B(n2557), .A(n1915), .Z(n2555) );
  MUX U4635 ( .IN0(n1883), .IN1(o[1167]), .SEL(n2562), .F(\Data_Mem/n6592 ) );
  MUX U4636 ( .IN0(n1885), .IN1(o[1166]), .SEL(n2562), .F(\Data_Mem/n6591 ) );
  MUX U4637 ( .IN0(n1886), .IN1(o[1165]), .SEL(n2562), .F(\Data_Mem/n6590 ) );
  MUX U4638 ( .IN0(n1887), .IN1(o[1164]), .SEL(n2562), .F(\Data_Mem/n6589 ) );
  MUX U4639 ( .IN0(n1888), .IN1(o[1163]), .SEL(n2562), .F(\Data_Mem/n6588 ) );
  IV U4640 ( .A(n2563), .Z(n2562) );
  MUX U4641 ( .IN0(o[1162]), .IN1(n1890), .SEL(n2563), .F(\Data_Mem/n6587 ) );
  MUX U4642 ( .IN0(o[1161]), .IN1(n1891), .SEL(n2563), .F(\Data_Mem/n6586 ) );
  MUX U4643 ( .IN0(o[1160]), .IN1(n1892), .SEL(n2563), .F(\Data_Mem/n6585 ) );
  NAND U4644 ( .A(n2564), .B(n2565), .Z(n2563) );
  OR U4645 ( .A(n1895), .B(n2557), .Z(n2565) );
  MUX U4646 ( .IN0(reg_target[7]), .IN1(o[1159]), .SEL(n2566), .F(
        \Data_Mem/n6584 ) );
  MUX U4647 ( .IN0(reg_target[6]), .IN1(o[1158]), .SEL(n2566), .F(
        \Data_Mem/n6583 ) );
  MUX U4648 ( .IN0(reg_target[5]), .IN1(o[1157]), .SEL(n2566), .F(
        \Data_Mem/n6582 ) );
  MUX U4649 ( .IN0(reg_target[4]), .IN1(o[1156]), .SEL(n2566), .F(
        \Data_Mem/n6581 ) );
  MUX U4650 ( .IN0(reg_target[3]), .IN1(o[1155]), .SEL(n2566), .F(
        \Data_Mem/n6580 ) );
  IV U4651 ( .A(n2567), .Z(n2566) );
  MUX U4652 ( .IN0(o[1154]), .IN1(reg_target[2]), .SEL(n2567), .F(
        \Data_Mem/n6579 ) );
  MUX U4653 ( .IN0(o[1153]), .IN1(reg_target[1]), .SEL(n2567), .F(
        \Data_Mem/n6578 ) );
  MUX U4654 ( .IN0(o[1152]), .IN1(reg_target[0]), .SEL(n2567), .F(
        \Data_Mem/n6577 ) );
  NAND U4655 ( .A(n2564), .B(n2568), .Z(n2567) );
  NANDN U4656 ( .B(n2557), .A(n1899), .Z(n2568) );
  ANDN U4657 ( .A(n2569), .B(n2554), .Z(n2564) );
  ANDN U4658 ( .A(n1902), .B(n2557), .Z(n2554) );
  NANDN U4659 ( .B(n2557), .A(n1924), .Z(n2569) );
  NAND U4660 ( .A(n1982), .B(n2497), .Z(n2557) );
  MUX U4661 ( .IN0(n1853), .IN1(o[1215]), .SEL(n2570), .F(\Data_Mem/n6576 ) );
  MUX U4662 ( .IN0(n1855), .IN1(o[1214]), .SEL(n2570), .F(\Data_Mem/n6575 ) );
  MUX U4663 ( .IN0(n1856), .IN1(o[1213]), .SEL(n2570), .F(\Data_Mem/n6574 ) );
  MUX U4664 ( .IN0(n1857), .IN1(o[1212]), .SEL(n2570), .F(\Data_Mem/n6573 ) );
  MUX U4665 ( .IN0(n1858), .IN1(o[1211]), .SEL(n2570), .F(\Data_Mem/n6572 ) );
  MUX U4666 ( .IN0(n1859), .IN1(o[1210]), .SEL(n2570), .F(\Data_Mem/n6571 ) );
  MUX U4667 ( .IN0(n1860), .IN1(o[1209]), .SEL(n2570), .F(\Data_Mem/n6570 ) );
  MUX U4668 ( .IN0(n1861), .IN1(o[1208]), .SEL(n2570), .F(\Data_Mem/n6569 ) );
  ANDN U4669 ( .A(n2571), .B(n2572), .Z(n2570) );
  AND U4670 ( .A(n2573), .B(n2574), .Z(n2571) );
  OR U4671 ( .A(n1867), .B(n2575), .Z(n2574) );
  MUX U4672 ( .IN0(n1868), .IN1(o[1207]), .SEL(n2576), .F(\Data_Mem/n6568 ) );
  MUX U4673 ( .IN0(n1870), .IN1(o[1206]), .SEL(n2576), .F(\Data_Mem/n6567 ) );
  MUX U4674 ( .IN0(n1871), .IN1(o[1205]), .SEL(n2576), .F(\Data_Mem/n6566 ) );
  MUX U4675 ( .IN0(n1872), .IN1(o[1204]), .SEL(n2576), .F(\Data_Mem/n6565 ) );
  MUX U4676 ( .IN0(n1873), .IN1(o[1203]), .SEL(n2576), .F(\Data_Mem/n6564 ) );
  IV U4677 ( .A(n2577), .Z(n2576) );
  MUX U4678 ( .IN0(o[1202]), .IN1(n1875), .SEL(n2577), .F(\Data_Mem/n6563 ) );
  MUX U4679 ( .IN0(o[1201]), .IN1(n1876), .SEL(n2577), .F(\Data_Mem/n6562 ) );
  MUX U4680 ( .IN0(o[1200]), .IN1(n1877), .SEL(n2577), .F(\Data_Mem/n6561 ) );
  NAND U4681 ( .A(n2578), .B(n2579), .Z(n2577) );
  OR U4682 ( .A(n1880), .B(n2575), .Z(n2579) );
  ANDN U4683 ( .A(n2573), .B(n2572), .Z(n2578) );
  NANDN U4684 ( .B(n2575), .A(n1915), .Z(n2573) );
  MUX U4685 ( .IN0(n1883), .IN1(o[1199]), .SEL(n2580), .F(\Data_Mem/n6560 ) );
  MUX U4686 ( .IN0(n1885), .IN1(o[1198]), .SEL(n2580), .F(\Data_Mem/n6559 ) );
  MUX U4687 ( .IN0(n1886), .IN1(o[1197]), .SEL(n2580), .F(\Data_Mem/n6558 ) );
  MUX U4688 ( .IN0(n1887), .IN1(o[1196]), .SEL(n2580), .F(\Data_Mem/n6557 ) );
  MUX U4689 ( .IN0(n1888), .IN1(o[1195]), .SEL(n2580), .F(\Data_Mem/n6556 ) );
  IV U4690 ( .A(n2581), .Z(n2580) );
  MUX U4691 ( .IN0(o[1194]), .IN1(n1890), .SEL(n2581), .F(\Data_Mem/n6555 ) );
  MUX U4692 ( .IN0(o[1193]), .IN1(n1891), .SEL(n2581), .F(\Data_Mem/n6554 ) );
  MUX U4693 ( .IN0(o[1192]), .IN1(n1892), .SEL(n2581), .F(\Data_Mem/n6553 ) );
  NAND U4694 ( .A(n2582), .B(n2583), .Z(n2581) );
  OR U4695 ( .A(n1895), .B(n2575), .Z(n2583) );
  MUX U4696 ( .IN0(reg_target[7]), .IN1(o[1191]), .SEL(n2584), .F(
        \Data_Mem/n6552 ) );
  MUX U4697 ( .IN0(reg_target[6]), .IN1(o[1190]), .SEL(n2584), .F(
        \Data_Mem/n6551 ) );
  MUX U4698 ( .IN0(reg_target[5]), .IN1(o[1189]), .SEL(n2584), .F(
        \Data_Mem/n6550 ) );
  MUX U4699 ( .IN0(reg_target[4]), .IN1(o[1188]), .SEL(n2584), .F(
        \Data_Mem/n6549 ) );
  MUX U4700 ( .IN0(reg_target[3]), .IN1(o[1187]), .SEL(n2584), .F(
        \Data_Mem/n6548 ) );
  IV U4701 ( .A(n2585), .Z(n2584) );
  MUX U4702 ( .IN0(o[1186]), .IN1(reg_target[2]), .SEL(n2585), .F(
        \Data_Mem/n6547 ) );
  MUX U4703 ( .IN0(o[1185]), .IN1(reg_target[1]), .SEL(n2585), .F(
        \Data_Mem/n6546 ) );
  MUX U4704 ( .IN0(o[1184]), .IN1(reg_target[0]), .SEL(n2585), .F(
        \Data_Mem/n6545 ) );
  NAND U4705 ( .A(n2582), .B(n2586), .Z(n2585) );
  NANDN U4706 ( .B(n2575), .A(n1899), .Z(n2586) );
  ANDN U4707 ( .A(n2587), .B(n2572), .Z(n2582) );
  ANDN U4708 ( .A(n1902), .B(n2575), .Z(n2572) );
  NANDN U4709 ( .B(n2575), .A(n1924), .Z(n2587) );
  NAND U4710 ( .A(n2001), .B(n2497), .Z(n2575) );
  MUX U4711 ( .IN0(n1853), .IN1(o[1247]), .SEL(n2588), .F(\Data_Mem/n6544 ) );
  MUX U4712 ( .IN0(n1855), .IN1(o[1246]), .SEL(n2588), .F(\Data_Mem/n6543 ) );
  MUX U4713 ( .IN0(n1856), .IN1(o[1245]), .SEL(n2588), .F(\Data_Mem/n6542 ) );
  MUX U4714 ( .IN0(n1857), .IN1(o[1244]), .SEL(n2588), .F(\Data_Mem/n6541 ) );
  MUX U4715 ( .IN0(n1858), .IN1(o[1243]), .SEL(n2588), .F(\Data_Mem/n6540 ) );
  MUX U4716 ( .IN0(n1859), .IN1(o[1242]), .SEL(n2588), .F(\Data_Mem/n6539 ) );
  MUX U4717 ( .IN0(n1860), .IN1(o[1241]), .SEL(n2588), .F(\Data_Mem/n6538 ) );
  MUX U4718 ( .IN0(n1861), .IN1(o[1240]), .SEL(n2588), .F(\Data_Mem/n6537 ) );
  ANDN U4719 ( .A(n2589), .B(n2590), .Z(n2588) );
  AND U4720 ( .A(n2591), .B(n2592), .Z(n2589) );
  OR U4721 ( .A(n1867), .B(n2593), .Z(n2592) );
  MUX U4722 ( .IN0(n1868), .IN1(o[1239]), .SEL(n2594), .F(\Data_Mem/n6536 ) );
  MUX U4723 ( .IN0(n1870), .IN1(o[1238]), .SEL(n2594), .F(\Data_Mem/n6535 ) );
  MUX U4724 ( .IN0(n1871), .IN1(o[1237]), .SEL(n2594), .F(\Data_Mem/n6534 ) );
  MUX U4725 ( .IN0(n1872), .IN1(o[1236]), .SEL(n2594), .F(\Data_Mem/n6533 ) );
  MUX U4726 ( .IN0(n1873), .IN1(o[1235]), .SEL(n2594), .F(\Data_Mem/n6532 ) );
  IV U4727 ( .A(n2595), .Z(n2594) );
  MUX U4728 ( .IN0(o[1234]), .IN1(n1875), .SEL(n2595), .F(\Data_Mem/n6531 ) );
  MUX U4729 ( .IN0(o[1233]), .IN1(n1876), .SEL(n2595), .F(\Data_Mem/n6530 ) );
  MUX U4730 ( .IN0(o[1232]), .IN1(n1877), .SEL(n2595), .F(\Data_Mem/n6529 ) );
  NAND U4731 ( .A(n2596), .B(n2597), .Z(n2595) );
  OR U4732 ( .A(n1880), .B(n2593), .Z(n2597) );
  ANDN U4733 ( .A(n2591), .B(n2590), .Z(n2596) );
  NANDN U4734 ( .B(n2593), .A(n1915), .Z(n2591) );
  MUX U4735 ( .IN0(n1883), .IN1(o[1231]), .SEL(n2598), .F(\Data_Mem/n6528 ) );
  MUX U4736 ( .IN0(n1885), .IN1(o[1230]), .SEL(n2598), .F(\Data_Mem/n6527 ) );
  MUX U4737 ( .IN0(n1886), .IN1(o[1229]), .SEL(n2598), .F(\Data_Mem/n6526 ) );
  MUX U4738 ( .IN0(n1887), .IN1(o[1228]), .SEL(n2598), .F(\Data_Mem/n6525 ) );
  MUX U4739 ( .IN0(n1888), .IN1(o[1227]), .SEL(n2598), .F(\Data_Mem/n6524 ) );
  IV U4740 ( .A(n2599), .Z(n2598) );
  MUX U4741 ( .IN0(o[1226]), .IN1(n1890), .SEL(n2599), .F(\Data_Mem/n6523 ) );
  MUX U4742 ( .IN0(o[1225]), .IN1(n1891), .SEL(n2599), .F(\Data_Mem/n6522 ) );
  MUX U4743 ( .IN0(o[1224]), .IN1(n1892), .SEL(n2599), .F(\Data_Mem/n6521 ) );
  NAND U4744 ( .A(n2600), .B(n2601), .Z(n2599) );
  OR U4745 ( .A(n1895), .B(n2593), .Z(n2601) );
  MUX U4746 ( .IN0(reg_target[7]), .IN1(o[1223]), .SEL(n2602), .F(
        \Data_Mem/n6520 ) );
  MUX U4747 ( .IN0(reg_target[6]), .IN1(o[1222]), .SEL(n2602), .F(
        \Data_Mem/n6519 ) );
  MUX U4748 ( .IN0(reg_target[5]), .IN1(o[1221]), .SEL(n2602), .F(
        \Data_Mem/n6518 ) );
  MUX U4749 ( .IN0(reg_target[4]), .IN1(o[1220]), .SEL(n2602), .F(
        \Data_Mem/n6517 ) );
  MUX U4750 ( .IN0(reg_target[3]), .IN1(o[1219]), .SEL(n2602), .F(
        \Data_Mem/n6516 ) );
  IV U4751 ( .A(n2603), .Z(n2602) );
  MUX U4752 ( .IN0(o[1218]), .IN1(reg_target[2]), .SEL(n2603), .F(
        \Data_Mem/n6515 ) );
  MUX U4753 ( .IN0(o[1217]), .IN1(reg_target[1]), .SEL(n2603), .F(
        \Data_Mem/n6514 ) );
  MUX U4754 ( .IN0(o[1216]), .IN1(reg_target[0]), .SEL(n2603), .F(
        \Data_Mem/n6513 ) );
  NAND U4755 ( .A(n2600), .B(n2604), .Z(n2603) );
  NANDN U4756 ( .B(n2593), .A(n1899), .Z(n2604) );
  ANDN U4757 ( .A(n2605), .B(n2590), .Z(n2600) );
  ANDN U4758 ( .A(n1902), .B(n2593), .Z(n2590) );
  NANDN U4759 ( .B(n2593), .A(n1924), .Z(n2605) );
  NAND U4760 ( .A(n2020), .B(n2497), .Z(n2593) );
  MUX U4761 ( .IN0(n1853), .IN1(o[1279]), .SEL(n2606), .F(\Data_Mem/n6512 ) );
  MUX U4762 ( .IN0(n1855), .IN1(o[1278]), .SEL(n2606), .F(\Data_Mem/n6511 ) );
  MUX U4763 ( .IN0(n1856), .IN1(o[1277]), .SEL(n2606), .F(\Data_Mem/n6510 ) );
  MUX U4764 ( .IN0(n1857), .IN1(o[1276]), .SEL(n2606), .F(\Data_Mem/n6509 ) );
  MUX U4765 ( .IN0(n1858), .IN1(o[1275]), .SEL(n2606), .F(\Data_Mem/n6508 ) );
  MUX U4766 ( .IN0(n1859), .IN1(o[1274]), .SEL(n2606), .F(\Data_Mem/n6507 ) );
  MUX U4767 ( .IN0(n1860), .IN1(o[1273]), .SEL(n2606), .F(\Data_Mem/n6506 ) );
  MUX U4768 ( .IN0(n1861), .IN1(o[1272]), .SEL(n2606), .F(\Data_Mem/n6505 ) );
  ANDN U4769 ( .A(n2607), .B(n2608), .Z(n2606) );
  AND U4770 ( .A(n2609), .B(n2610), .Z(n2607) );
  OR U4771 ( .A(n1867), .B(n2611), .Z(n2610) );
  MUX U4772 ( .IN0(n1868), .IN1(o[1271]), .SEL(n2612), .F(\Data_Mem/n6504 ) );
  MUX U4773 ( .IN0(n1870), .IN1(o[1270]), .SEL(n2612), .F(\Data_Mem/n6503 ) );
  MUX U4774 ( .IN0(n1871), .IN1(o[1269]), .SEL(n2612), .F(\Data_Mem/n6502 ) );
  MUX U4775 ( .IN0(n1872), .IN1(o[1268]), .SEL(n2612), .F(\Data_Mem/n6501 ) );
  MUX U4776 ( .IN0(n1873), .IN1(o[1267]), .SEL(n2612), .F(\Data_Mem/n6500 ) );
  IV U4777 ( .A(n2613), .Z(n2612) );
  MUX U4778 ( .IN0(o[1266]), .IN1(n1875), .SEL(n2613), .F(\Data_Mem/n6499 ) );
  MUX U4779 ( .IN0(o[1265]), .IN1(n1876), .SEL(n2613), .F(\Data_Mem/n6498 ) );
  MUX U4780 ( .IN0(o[1264]), .IN1(n1877), .SEL(n2613), .F(\Data_Mem/n6497 ) );
  NAND U4781 ( .A(n2614), .B(n2615), .Z(n2613) );
  OR U4782 ( .A(n1880), .B(n2611), .Z(n2615) );
  ANDN U4783 ( .A(n2609), .B(n2608), .Z(n2614) );
  NANDN U4784 ( .B(n2611), .A(n1915), .Z(n2609) );
  MUX U4785 ( .IN0(n1883), .IN1(o[1263]), .SEL(n2616), .F(\Data_Mem/n6496 ) );
  MUX U4786 ( .IN0(n1885), .IN1(o[1262]), .SEL(n2616), .F(\Data_Mem/n6495 ) );
  MUX U4787 ( .IN0(n1886), .IN1(o[1261]), .SEL(n2616), .F(\Data_Mem/n6494 ) );
  MUX U4788 ( .IN0(n1887), .IN1(o[1260]), .SEL(n2616), .F(\Data_Mem/n6493 ) );
  MUX U4789 ( .IN0(n1888), .IN1(o[1259]), .SEL(n2616), .F(\Data_Mem/n6492 ) );
  IV U4790 ( .A(n2617), .Z(n2616) );
  MUX U4791 ( .IN0(o[1258]), .IN1(n1890), .SEL(n2617), .F(\Data_Mem/n6491 ) );
  MUX U4792 ( .IN0(o[1257]), .IN1(n1891), .SEL(n2617), .F(\Data_Mem/n6490 ) );
  MUX U4793 ( .IN0(o[1256]), .IN1(n1892), .SEL(n2617), .F(\Data_Mem/n6489 ) );
  NAND U4794 ( .A(n2618), .B(n2619), .Z(n2617) );
  OR U4795 ( .A(n1895), .B(n2611), .Z(n2619) );
  MUX U4796 ( .IN0(reg_target[7]), .IN1(o[1255]), .SEL(n2620), .F(
        \Data_Mem/n6488 ) );
  MUX U4797 ( .IN0(reg_target[6]), .IN1(o[1254]), .SEL(n2620), .F(
        \Data_Mem/n6487 ) );
  MUX U4798 ( .IN0(reg_target[5]), .IN1(o[1253]), .SEL(n2620), .F(
        \Data_Mem/n6486 ) );
  MUX U4799 ( .IN0(reg_target[4]), .IN1(o[1252]), .SEL(n2620), .F(
        \Data_Mem/n6485 ) );
  MUX U4800 ( .IN0(reg_target[3]), .IN1(o[1251]), .SEL(n2620), .F(
        \Data_Mem/n6484 ) );
  IV U4801 ( .A(n2621), .Z(n2620) );
  MUX U4802 ( .IN0(o[1250]), .IN1(reg_target[2]), .SEL(n2621), .F(
        \Data_Mem/n6483 ) );
  MUX U4803 ( .IN0(o[1249]), .IN1(reg_target[1]), .SEL(n2621), .F(
        \Data_Mem/n6482 ) );
  MUX U4804 ( .IN0(o[1248]), .IN1(reg_target[0]), .SEL(n2621), .F(
        \Data_Mem/n6481 ) );
  NAND U4805 ( .A(n2618), .B(n2622), .Z(n2621) );
  NANDN U4806 ( .B(n2611), .A(n1899), .Z(n2622) );
  ANDN U4807 ( .A(n2623), .B(n2608), .Z(n2618) );
  ANDN U4808 ( .A(n1902), .B(n2611), .Z(n2608) );
  NANDN U4809 ( .B(n2611), .A(n1924), .Z(n2623) );
  NAND U4810 ( .A(n2497), .B(n2039), .Z(n2611) );
  ANDN U4811 ( .A(n2040), .B(n485), .Z(n2497) );
  AND U4812 ( .A(n532), .B(n511), .Z(n2040) );
  MUX U4813 ( .IN0(n1853), .IN1(o[1311]), .SEL(n2624), .F(\Data_Mem/n6480 ) );
  MUX U4814 ( .IN0(n1855), .IN1(o[1310]), .SEL(n2624), .F(\Data_Mem/n6479 ) );
  MUX U4815 ( .IN0(n1856), .IN1(o[1309]), .SEL(n2624), .F(\Data_Mem/n6478 ) );
  MUX U4816 ( .IN0(n1857), .IN1(o[1308]), .SEL(n2624), .F(\Data_Mem/n6477 ) );
  MUX U4817 ( .IN0(n1858), .IN1(o[1307]), .SEL(n2624), .F(\Data_Mem/n6476 ) );
  MUX U4818 ( .IN0(n1859), .IN1(o[1306]), .SEL(n2624), .F(\Data_Mem/n6475 ) );
  MUX U4819 ( .IN0(n1860), .IN1(o[1305]), .SEL(n2624), .F(\Data_Mem/n6474 ) );
  MUX U4820 ( .IN0(n1861), .IN1(o[1304]), .SEL(n2624), .F(\Data_Mem/n6473 ) );
  ANDN U4821 ( .A(n2625), .B(n2626), .Z(n2624) );
  AND U4822 ( .A(n2627), .B(n2628), .Z(n2625) );
  OR U4823 ( .A(n1867), .B(n2629), .Z(n2628) );
  MUX U4824 ( .IN0(n1868), .IN1(o[1303]), .SEL(n2630), .F(\Data_Mem/n6472 ) );
  MUX U4825 ( .IN0(n1870), .IN1(o[1302]), .SEL(n2630), .F(\Data_Mem/n6471 ) );
  MUX U4826 ( .IN0(n1871), .IN1(o[1301]), .SEL(n2630), .F(\Data_Mem/n6470 ) );
  MUX U4827 ( .IN0(n1872), .IN1(o[1300]), .SEL(n2630), .F(\Data_Mem/n6469 ) );
  MUX U4828 ( .IN0(n1873), .IN1(o[1299]), .SEL(n2630), .F(\Data_Mem/n6468 ) );
  IV U4829 ( .A(n2631), .Z(n2630) );
  MUX U4830 ( .IN0(o[1298]), .IN1(n1875), .SEL(n2631), .F(\Data_Mem/n6467 ) );
  MUX U4831 ( .IN0(o[1297]), .IN1(n1876), .SEL(n2631), .F(\Data_Mem/n6466 ) );
  MUX U4832 ( .IN0(o[1296]), .IN1(n1877), .SEL(n2631), .F(\Data_Mem/n6465 ) );
  NAND U4833 ( .A(n2632), .B(n2633), .Z(n2631) );
  OR U4834 ( .A(n1880), .B(n2629), .Z(n2633) );
  ANDN U4835 ( .A(n2627), .B(n2626), .Z(n2632) );
  NANDN U4836 ( .B(n2629), .A(n1915), .Z(n2627) );
  MUX U4837 ( .IN0(n1883), .IN1(o[1295]), .SEL(n2634), .F(\Data_Mem/n6464 ) );
  MUX U4838 ( .IN0(n1885), .IN1(o[1294]), .SEL(n2634), .F(\Data_Mem/n6463 ) );
  MUX U4839 ( .IN0(n1886), .IN1(o[1293]), .SEL(n2634), .F(\Data_Mem/n6462 ) );
  MUX U4840 ( .IN0(n1887), .IN1(o[1292]), .SEL(n2634), .F(\Data_Mem/n6461 ) );
  MUX U4841 ( .IN0(n1888), .IN1(o[1291]), .SEL(n2634), .F(\Data_Mem/n6460 ) );
  IV U4842 ( .A(n2635), .Z(n2634) );
  MUX U4843 ( .IN0(o[1290]), .IN1(n1890), .SEL(n2635), .F(\Data_Mem/n6459 ) );
  MUX U4844 ( .IN0(o[1289]), .IN1(n1891), .SEL(n2635), .F(\Data_Mem/n6458 ) );
  MUX U4845 ( .IN0(o[1288]), .IN1(n1892), .SEL(n2635), .F(\Data_Mem/n6457 ) );
  NAND U4846 ( .A(n2636), .B(n2637), .Z(n2635) );
  OR U4847 ( .A(n1895), .B(n2629), .Z(n2637) );
  MUX U4848 ( .IN0(reg_target[7]), .IN1(o[1287]), .SEL(n2638), .F(
        \Data_Mem/n6456 ) );
  MUX U4849 ( .IN0(reg_target[6]), .IN1(o[1286]), .SEL(n2638), .F(
        \Data_Mem/n6455 ) );
  MUX U4850 ( .IN0(reg_target[5]), .IN1(o[1285]), .SEL(n2638), .F(
        \Data_Mem/n6454 ) );
  MUX U4851 ( .IN0(reg_target[4]), .IN1(o[1284]), .SEL(n2638), .F(
        \Data_Mem/n6453 ) );
  MUX U4852 ( .IN0(reg_target[3]), .IN1(o[1283]), .SEL(n2638), .F(
        \Data_Mem/n6452 ) );
  IV U4853 ( .A(n2639), .Z(n2638) );
  MUX U4854 ( .IN0(o[1282]), .IN1(reg_target[2]), .SEL(n2639), .F(
        \Data_Mem/n6451 ) );
  MUX U4855 ( .IN0(o[1281]), .IN1(reg_target[1]), .SEL(n2639), .F(
        \Data_Mem/n6450 ) );
  MUX U4856 ( .IN0(o[1280]), .IN1(reg_target[0]), .SEL(n2639), .F(
        \Data_Mem/n6449 ) );
  NAND U4857 ( .A(n2636), .B(n2640), .Z(n2639) );
  NANDN U4858 ( .B(n2629), .A(n1899), .Z(n2640) );
  ANDN U4859 ( .A(n2641), .B(n2626), .Z(n2636) );
  ANDN U4860 ( .A(n1902), .B(n2629), .Z(n2626) );
  NANDN U4861 ( .B(n2629), .A(n1924), .Z(n2641) );
  NAND U4862 ( .A(n1903), .B(n2642), .Z(n2629) );
  MUX U4863 ( .IN0(n1853), .IN1(o[1343]), .SEL(n2643), .F(\Data_Mem/n6448 ) );
  MUX U4864 ( .IN0(n1855), .IN1(o[1342]), .SEL(n2643), .F(\Data_Mem/n6447 ) );
  MUX U4865 ( .IN0(n1856), .IN1(o[1341]), .SEL(n2643), .F(\Data_Mem/n6446 ) );
  MUX U4866 ( .IN0(n1857), .IN1(o[1340]), .SEL(n2643), .F(\Data_Mem/n6445 ) );
  MUX U4867 ( .IN0(n1858), .IN1(o[1339]), .SEL(n2643), .F(\Data_Mem/n6444 ) );
  MUX U4868 ( .IN0(n1859), .IN1(o[1338]), .SEL(n2643), .F(\Data_Mem/n6443 ) );
  MUX U4869 ( .IN0(n1860), .IN1(o[1337]), .SEL(n2643), .F(\Data_Mem/n6442 ) );
  MUX U4870 ( .IN0(n1861), .IN1(o[1336]), .SEL(n2643), .F(\Data_Mem/n6441 ) );
  ANDN U4871 ( .A(n2644), .B(n2645), .Z(n2643) );
  AND U4872 ( .A(n2646), .B(n2647), .Z(n2644) );
  OR U4873 ( .A(n1867), .B(n2648), .Z(n2647) );
  MUX U4874 ( .IN0(n1868), .IN1(o[1335]), .SEL(n2649), .F(\Data_Mem/n6440 ) );
  MUX U4875 ( .IN0(n1870), .IN1(o[1334]), .SEL(n2649), .F(\Data_Mem/n6439 ) );
  MUX U4876 ( .IN0(n1871), .IN1(o[1333]), .SEL(n2649), .F(\Data_Mem/n6438 ) );
  MUX U4877 ( .IN0(n1872), .IN1(o[1332]), .SEL(n2649), .F(\Data_Mem/n6437 ) );
  MUX U4878 ( .IN0(n1873), .IN1(o[1331]), .SEL(n2649), .F(\Data_Mem/n6436 ) );
  IV U4879 ( .A(n2650), .Z(n2649) );
  MUX U4880 ( .IN0(o[1330]), .IN1(n1875), .SEL(n2650), .F(\Data_Mem/n6435 ) );
  MUX U4881 ( .IN0(o[1329]), .IN1(n1876), .SEL(n2650), .F(\Data_Mem/n6434 ) );
  MUX U4882 ( .IN0(o[1328]), .IN1(n1877), .SEL(n2650), .F(\Data_Mem/n6433 ) );
  NAND U4883 ( .A(n2651), .B(n2652), .Z(n2650) );
  OR U4884 ( .A(n1880), .B(n2648), .Z(n2652) );
  ANDN U4885 ( .A(n2646), .B(n2645), .Z(n2651) );
  NANDN U4886 ( .B(n2648), .A(n1915), .Z(n2646) );
  MUX U4887 ( .IN0(n1883), .IN1(o[1327]), .SEL(n2653), .F(\Data_Mem/n6432 ) );
  MUX U4888 ( .IN0(n1885), .IN1(o[1326]), .SEL(n2653), .F(\Data_Mem/n6431 ) );
  MUX U4889 ( .IN0(n1886), .IN1(o[1325]), .SEL(n2653), .F(\Data_Mem/n6430 ) );
  MUX U4890 ( .IN0(n1887), .IN1(o[1324]), .SEL(n2653), .F(\Data_Mem/n6429 ) );
  MUX U4891 ( .IN0(n1888), .IN1(o[1323]), .SEL(n2653), .F(\Data_Mem/n6428 ) );
  IV U4892 ( .A(n2654), .Z(n2653) );
  MUX U4893 ( .IN0(o[1322]), .IN1(n1890), .SEL(n2654), .F(\Data_Mem/n6427 ) );
  MUX U4894 ( .IN0(o[1321]), .IN1(n1891), .SEL(n2654), .F(\Data_Mem/n6426 ) );
  MUX U4895 ( .IN0(o[1320]), .IN1(n1892), .SEL(n2654), .F(\Data_Mem/n6425 ) );
  NAND U4896 ( .A(n2655), .B(n2656), .Z(n2654) );
  OR U4897 ( .A(n1895), .B(n2648), .Z(n2656) );
  MUX U4898 ( .IN0(reg_target[7]), .IN1(o[1319]), .SEL(n2657), .F(
        \Data_Mem/n6424 ) );
  MUX U4899 ( .IN0(reg_target[6]), .IN1(o[1318]), .SEL(n2657), .F(
        \Data_Mem/n6423 ) );
  MUX U4900 ( .IN0(reg_target[5]), .IN1(o[1317]), .SEL(n2657), .F(
        \Data_Mem/n6422 ) );
  MUX U4901 ( .IN0(reg_target[4]), .IN1(o[1316]), .SEL(n2657), .F(
        \Data_Mem/n6421 ) );
  MUX U4902 ( .IN0(reg_target[3]), .IN1(o[1315]), .SEL(n2657), .F(
        \Data_Mem/n6420 ) );
  IV U4903 ( .A(n2658), .Z(n2657) );
  MUX U4904 ( .IN0(o[1314]), .IN1(reg_target[2]), .SEL(n2658), .F(
        \Data_Mem/n6419 ) );
  MUX U4905 ( .IN0(o[1313]), .IN1(reg_target[1]), .SEL(n2658), .F(
        \Data_Mem/n6418 ) );
  MUX U4906 ( .IN0(o[1312]), .IN1(reg_target[0]), .SEL(n2658), .F(
        \Data_Mem/n6417 ) );
  NAND U4907 ( .A(n2655), .B(n2659), .Z(n2658) );
  NANDN U4908 ( .B(n2648), .A(n1899), .Z(n2659) );
  ANDN U4909 ( .A(n2660), .B(n2645), .Z(n2655) );
  ANDN U4910 ( .A(n1902), .B(n2648), .Z(n2645) );
  NANDN U4911 ( .B(n2648), .A(n1924), .Z(n2660) );
  NAND U4912 ( .A(n1925), .B(n2642), .Z(n2648) );
  MUX U4913 ( .IN0(n1853), .IN1(o[1375]), .SEL(n2661), .F(\Data_Mem/n6416 ) );
  MUX U4914 ( .IN0(n1855), .IN1(o[1374]), .SEL(n2661), .F(\Data_Mem/n6415 ) );
  MUX U4915 ( .IN0(n1856), .IN1(o[1373]), .SEL(n2661), .F(\Data_Mem/n6414 ) );
  MUX U4916 ( .IN0(n1857), .IN1(o[1372]), .SEL(n2661), .F(\Data_Mem/n6413 ) );
  MUX U4917 ( .IN0(n1858), .IN1(o[1371]), .SEL(n2661), .F(\Data_Mem/n6412 ) );
  MUX U4918 ( .IN0(n1859), .IN1(o[1370]), .SEL(n2661), .F(\Data_Mem/n6411 ) );
  MUX U4919 ( .IN0(n1860), .IN1(o[1369]), .SEL(n2661), .F(\Data_Mem/n6410 ) );
  MUX U4920 ( .IN0(n1861), .IN1(o[1368]), .SEL(n2661), .F(\Data_Mem/n6409 ) );
  ANDN U4921 ( .A(n2662), .B(n2663), .Z(n2661) );
  AND U4922 ( .A(n2664), .B(n2665), .Z(n2662) );
  OR U4923 ( .A(n1867), .B(n2666), .Z(n2665) );
  MUX U4924 ( .IN0(n1868), .IN1(o[1367]), .SEL(n2667), .F(\Data_Mem/n6408 ) );
  MUX U4925 ( .IN0(n1870), .IN1(o[1366]), .SEL(n2667), .F(\Data_Mem/n6407 ) );
  MUX U4926 ( .IN0(n1871), .IN1(o[1365]), .SEL(n2667), .F(\Data_Mem/n6406 ) );
  MUX U4927 ( .IN0(n1872), .IN1(o[1364]), .SEL(n2667), .F(\Data_Mem/n6405 ) );
  MUX U4928 ( .IN0(n1873), .IN1(o[1363]), .SEL(n2667), .F(\Data_Mem/n6404 ) );
  IV U4929 ( .A(n2668), .Z(n2667) );
  MUX U4930 ( .IN0(o[1362]), .IN1(n1875), .SEL(n2668), .F(\Data_Mem/n6403 ) );
  MUX U4931 ( .IN0(o[1361]), .IN1(n1876), .SEL(n2668), .F(\Data_Mem/n6402 ) );
  MUX U4932 ( .IN0(o[1360]), .IN1(n1877), .SEL(n2668), .F(\Data_Mem/n6401 ) );
  NAND U4933 ( .A(n2669), .B(n2670), .Z(n2668) );
  OR U4934 ( .A(n1880), .B(n2666), .Z(n2670) );
  ANDN U4935 ( .A(n2664), .B(n2663), .Z(n2669) );
  NANDN U4936 ( .B(n2666), .A(n1915), .Z(n2664) );
  MUX U4937 ( .IN0(n1883), .IN1(o[1359]), .SEL(n2671), .F(\Data_Mem/n6400 ) );
  MUX U4938 ( .IN0(n1885), .IN1(o[1358]), .SEL(n2671), .F(\Data_Mem/n6399 ) );
  MUX U4939 ( .IN0(n1886), .IN1(o[1357]), .SEL(n2671), .F(\Data_Mem/n6398 ) );
  MUX U4940 ( .IN0(n1887), .IN1(o[1356]), .SEL(n2671), .F(\Data_Mem/n6397 ) );
  MUX U4941 ( .IN0(n1888), .IN1(o[1355]), .SEL(n2671), .F(\Data_Mem/n6396 ) );
  IV U4942 ( .A(n2672), .Z(n2671) );
  MUX U4943 ( .IN0(o[1354]), .IN1(n1890), .SEL(n2672), .F(\Data_Mem/n6395 ) );
  MUX U4944 ( .IN0(o[1353]), .IN1(n1891), .SEL(n2672), .F(\Data_Mem/n6394 ) );
  MUX U4945 ( .IN0(o[1352]), .IN1(n1892), .SEL(n2672), .F(\Data_Mem/n6393 ) );
  NAND U4946 ( .A(n2673), .B(n2674), .Z(n2672) );
  OR U4947 ( .A(n1895), .B(n2666), .Z(n2674) );
  MUX U4948 ( .IN0(reg_target[7]), .IN1(o[1351]), .SEL(n2675), .F(
        \Data_Mem/n6392 ) );
  MUX U4949 ( .IN0(reg_target[6]), .IN1(o[1350]), .SEL(n2675), .F(
        \Data_Mem/n6391 ) );
  MUX U4950 ( .IN0(reg_target[5]), .IN1(o[1349]), .SEL(n2675), .F(
        \Data_Mem/n6390 ) );
  MUX U4951 ( .IN0(reg_target[4]), .IN1(o[1348]), .SEL(n2675), .F(
        \Data_Mem/n6389 ) );
  MUX U4952 ( .IN0(reg_target[3]), .IN1(o[1347]), .SEL(n2675), .F(
        \Data_Mem/n6388 ) );
  IV U4953 ( .A(n2676), .Z(n2675) );
  MUX U4954 ( .IN0(o[1346]), .IN1(reg_target[2]), .SEL(n2676), .F(
        \Data_Mem/n6387 ) );
  MUX U4955 ( .IN0(o[1345]), .IN1(reg_target[1]), .SEL(n2676), .F(
        \Data_Mem/n6386 ) );
  MUX U4956 ( .IN0(o[1344]), .IN1(reg_target[0]), .SEL(n2676), .F(
        \Data_Mem/n6385 ) );
  NAND U4957 ( .A(n2673), .B(n2677), .Z(n2676) );
  NANDN U4958 ( .B(n2666), .A(n1899), .Z(n2677) );
  ANDN U4959 ( .A(n2678), .B(n2663), .Z(n2673) );
  ANDN U4960 ( .A(n1902), .B(n2666), .Z(n2663) );
  NANDN U4961 ( .B(n2666), .A(n1924), .Z(n2678) );
  NAND U4962 ( .A(n1944), .B(n2642), .Z(n2666) );
  MUX U4963 ( .IN0(n1853), .IN1(o[1407]), .SEL(n2679), .F(\Data_Mem/n6384 ) );
  MUX U4964 ( .IN0(n1855), .IN1(o[1406]), .SEL(n2679), .F(\Data_Mem/n6383 ) );
  MUX U4965 ( .IN0(n1856), .IN1(o[1405]), .SEL(n2679), .F(\Data_Mem/n6382 ) );
  MUX U4966 ( .IN0(n1857), .IN1(o[1404]), .SEL(n2679), .F(\Data_Mem/n6381 ) );
  MUX U4967 ( .IN0(n1858), .IN1(o[1403]), .SEL(n2679), .F(\Data_Mem/n6380 ) );
  MUX U4968 ( .IN0(n1859), .IN1(o[1402]), .SEL(n2679), .F(\Data_Mem/n6379 ) );
  MUX U4969 ( .IN0(n1860), .IN1(o[1401]), .SEL(n2679), .F(\Data_Mem/n6378 ) );
  MUX U4970 ( .IN0(n1861), .IN1(o[1400]), .SEL(n2679), .F(\Data_Mem/n6377 ) );
  ANDN U4971 ( .A(n2680), .B(n2681), .Z(n2679) );
  AND U4972 ( .A(n2682), .B(n2683), .Z(n2680) );
  OR U4973 ( .A(n1867), .B(n2684), .Z(n2683) );
  MUX U4974 ( .IN0(n1868), .IN1(o[1399]), .SEL(n2685), .F(\Data_Mem/n6376 ) );
  MUX U4975 ( .IN0(n1870), .IN1(o[1398]), .SEL(n2685), .F(\Data_Mem/n6375 ) );
  MUX U4976 ( .IN0(n1871), .IN1(o[1397]), .SEL(n2685), .F(\Data_Mem/n6374 ) );
  MUX U4977 ( .IN0(n1872), .IN1(o[1396]), .SEL(n2685), .F(\Data_Mem/n6373 ) );
  MUX U4978 ( .IN0(n1873), .IN1(o[1395]), .SEL(n2685), .F(\Data_Mem/n6372 ) );
  IV U4979 ( .A(n2686), .Z(n2685) );
  MUX U4980 ( .IN0(o[1394]), .IN1(n1875), .SEL(n2686), .F(\Data_Mem/n6371 ) );
  MUX U4981 ( .IN0(o[1393]), .IN1(n1876), .SEL(n2686), .F(\Data_Mem/n6370 ) );
  MUX U4982 ( .IN0(o[1392]), .IN1(n1877), .SEL(n2686), .F(\Data_Mem/n6369 ) );
  NAND U4983 ( .A(n2687), .B(n2688), .Z(n2686) );
  OR U4984 ( .A(n1880), .B(n2684), .Z(n2688) );
  ANDN U4985 ( .A(n2682), .B(n2681), .Z(n2687) );
  NANDN U4986 ( .B(n2684), .A(n1915), .Z(n2682) );
  MUX U4987 ( .IN0(n1883), .IN1(o[1391]), .SEL(n2689), .F(\Data_Mem/n6368 ) );
  MUX U4988 ( .IN0(n1885), .IN1(o[1390]), .SEL(n2689), .F(\Data_Mem/n6367 ) );
  MUX U4989 ( .IN0(n1886), .IN1(o[1389]), .SEL(n2689), .F(\Data_Mem/n6366 ) );
  MUX U4990 ( .IN0(n1887), .IN1(o[1388]), .SEL(n2689), .F(\Data_Mem/n6365 ) );
  MUX U4991 ( .IN0(n1888), .IN1(o[1387]), .SEL(n2689), .F(\Data_Mem/n6364 ) );
  IV U4992 ( .A(n2690), .Z(n2689) );
  MUX U4993 ( .IN0(o[1386]), .IN1(n1890), .SEL(n2690), .F(\Data_Mem/n6363 ) );
  MUX U4994 ( .IN0(o[1385]), .IN1(n1891), .SEL(n2690), .F(\Data_Mem/n6362 ) );
  MUX U4995 ( .IN0(o[1384]), .IN1(n1892), .SEL(n2690), .F(\Data_Mem/n6361 ) );
  NAND U4996 ( .A(n2691), .B(n2692), .Z(n2690) );
  OR U4997 ( .A(n1895), .B(n2684), .Z(n2692) );
  MUX U4998 ( .IN0(reg_target[7]), .IN1(o[1383]), .SEL(n2693), .F(
        \Data_Mem/n6360 ) );
  MUX U4999 ( .IN0(reg_target[6]), .IN1(o[1382]), .SEL(n2693), .F(
        \Data_Mem/n6359 ) );
  MUX U5000 ( .IN0(reg_target[5]), .IN1(o[1381]), .SEL(n2693), .F(
        \Data_Mem/n6358 ) );
  MUX U5001 ( .IN0(reg_target[4]), .IN1(o[1380]), .SEL(n2693), .F(
        \Data_Mem/n6357 ) );
  MUX U5002 ( .IN0(reg_target[3]), .IN1(o[1379]), .SEL(n2693), .F(
        \Data_Mem/n6356 ) );
  IV U5003 ( .A(n2694), .Z(n2693) );
  MUX U5004 ( .IN0(o[1378]), .IN1(reg_target[2]), .SEL(n2694), .F(
        \Data_Mem/n6355 ) );
  MUX U5005 ( .IN0(o[1377]), .IN1(reg_target[1]), .SEL(n2694), .F(
        \Data_Mem/n6354 ) );
  MUX U5006 ( .IN0(o[1376]), .IN1(reg_target[0]), .SEL(n2694), .F(
        \Data_Mem/n6353 ) );
  NAND U5007 ( .A(n2691), .B(n2695), .Z(n2694) );
  NANDN U5008 ( .B(n2684), .A(n1899), .Z(n2695) );
  ANDN U5009 ( .A(n2696), .B(n2681), .Z(n2691) );
  ANDN U5010 ( .A(n1902), .B(n2684), .Z(n2681) );
  NANDN U5011 ( .B(n2684), .A(n1924), .Z(n2696) );
  NAND U5012 ( .A(n1963), .B(n2642), .Z(n2684) );
  MUX U5013 ( .IN0(n1853), .IN1(o[1439]), .SEL(n2697), .F(\Data_Mem/n6352 ) );
  MUX U5014 ( .IN0(n1855), .IN1(o[1438]), .SEL(n2697), .F(\Data_Mem/n6351 ) );
  MUX U5015 ( .IN0(n1856), .IN1(o[1437]), .SEL(n2697), .F(\Data_Mem/n6350 ) );
  MUX U5016 ( .IN0(n1857), .IN1(o[1436]), .SEL(n2697), .F(\Data_Mem/n6349 ) );
  MUX U5017 ( .IN0(n1858), .IN1(o[1435]), .SEL(n2697), .F(\Data_Mem/n6348 ) );
  MUX U5018 ( .IN0(n1859), .IN1(o[1434]), .SEL(n2697), .F(\Data_Mem/n6347 ) );
  MUX U5019 ( .IN0(n1860), .IN1(o[1433]), .SEL(n2697), .F(\Data_Mem/n6346 ) );
  MUX U5020 ( .IN0(n1861), .IN1(o[1432]), .SEL(n2697), .F(\Data_Mem/n6345 ) );
  ANDN U5021 ( .A(n2698), .B(n2699), .Z(n2697) );
  AND U5022 ( .A(n2700), .B(n2701), .Z(n2698) );
  OR U5023 ( .A(n1867), .B(n2702), .Z(n2701) );
  MUX U5024 ( .IN0(n1868), .IN1(o[1431]), .SEL(n2703), .F(\Data_Mem/n6344 ) );
  MUX U5025 ( .IN0(n1870), .IN1(o[1430]), .SEL(n2703), .F(\Data_Mem/n6343 ) );
  MUX U5026 ( .IN0(n1871), .IN1(o[1429]), .SEL(n2703), .F(\Data_Mem/n6342 ) );
  MUX U5027 ( .IN0(n1872), .IN1(o[1428]), .SEL(n2703), .F(\Data_Mem/n6341 ) );
  MUX U5028 ( .IN0(n1873), .IN1(o[1427]), .SEL(n2703), .F(\Data_Mem/n6340 ) );
  IV U5029 ( .A(n2704), .Z(n2703) );
  MUX U5030 ( .IN0(o[1426]), .IN1(n1875), .SEL(n2704), .F(\Data_Mem/n6339 ) );
  MUX U5031 ( .IN0(o[1425]), .IN1(n1876), .SEL(n2704), .F(\Data_Mem/n6338 ) );
  MUX U5032 ( .IN0(o[1424]), .IN1(n1877), .SEL(n2704), .F(\Data_Mem/n6337 ) );
  NAND U5033 ( .A(n2705), .B(n2706), .Z(n2704) );
  OR U5034 ( .A(n1880), .B(n2702), .Z(n2706) );
  ANDN U5035 ( .A(n2700), .B(n2699), .Z(n2705) );
  NANDN U5036 ( .B(n2702), .A(n1915), .Z(n2700) );
  MUX U5037 ( .IN0(n1883), .IN1(o[1423]), .SEL(n2707), .F(\Data_Mem/n6336 ) );
  MUX U5038 ( .IN0(n1885), .IN1(o[1422]), .SEL(n2707), .F(\Data_Mem/n6335 ) );
  MUX U5039 ( .IN0(n1886), .IN1(o[1421]), .SEL(n2707), .F(\Data_Mem/n6334 ) );
  MUX U5040 ( .IN0(n1887), .IN1(o[1420]), .SEL(n2707), .F(\Data_Mem/n6333 ) );
  MUX U5041 ( .IN0(n1888), .IN1(o[1419]), .SEL(n2707), .F(\Data_Mem/n6332 ) );
  IV U5042 ( .A(n2708), .Z(n2707) );
  MUX U5043 ( .IN0(o[1418]), .IN1(n1890), .SEL(n2708), .F(\Data_Mem/n6331 ) );
  MUX U5044 ( .IN0(o[1417]), .IN1(n1891), .SEL(n2708), .F(\Data_Mem/n6330 ) );
  MUX U5045 ( .IN0(o[1416]), .IN1(n1892), .SEL(n2708), .F(\Data_Mem/n6329 ) );
  NAND U5046 ( .A(n2709), .B(n2710), .Z(n2708) );
  OR U5047 ( .A(n1895), .B(n2702), .Z(n2710) );
  MUX U5048 ( .IN0(reg_target[7]), .IN1(o[1415]), .SEL(n2711), .F(
        \Data_Mem/n6328 ) );
  MUX U5049 ( .IN0(reg_target[6]), .IN1(o[1414]), .SEL(n2711), .F(
        \Data_Mem/n6327 ) );
  MUX U5050 ( .IN0(reg_target[5]), .IN1(o[1413]), .SEL(n2711), .F(
        \Data_Mem/n6326 ) );
  MUX U5051 ( .IN0(reg_target[4]), .IN1(o[1412]), .SEL(n2711), .F(
        \Data_Mem/n6325 ) );
  MUX U5052 ( .IN0(reg_target[3]), .IN1(o[1411]), .SEL(n2711), .F(
        \Data_Mem/n6324 ) );
  IV U5053 ( .A(n2712), .Z(n2711) );
  MUX U5054 ( .IN0(o[1410]), .IN1(reg_target[2]), .SEL(n2712), .F(
        \Data_Mem/n6323 ) );
  MUX U5055 ( .IN0(o[1409]), .IN1(reg_target[1]), .SEL(n2712), .F(
        \Data_Mem/n6322 ) );
  MUX U5056 ( .IN0(o[1408]), .IN1(reg_target[0]), .SEL(n2712), .F(
        \Data_Mem/n6321 ) );
  NAND U5057 ( .A(n2709), .B(n2713), .Z(n2712) );
  NANDN U5058 ( .B(n2702), .A(n1899), .Z(n2713) );
  ANDN U5059 ( .A(n2714), .B(n2699), .Z(n2709) );
  ANDN U5060 ( .A(n1902), .B(n2702), .Z(n2699) );
  NANDN U5061 ( .B(n2702), .A(n1924), .Z(n2714) );
  NAND U5062 ( .A(n1982), .B(n2642), .Z(n2702) );
  MUX U5063 ( .IN0(n1853), .IN1(o[1471]), .SEL(n2715), .F(\Data_Mem/n6320 ) );
  MUX U5064 ( .IN0(n1855), .IN1(o[1470]), .SEL(n2715), .F(\Data_Mem/n6319 ) );
  MUX U5065 ( .IN0(n1856), .IN1(o[1469]), .SEL(n2715), .F(\Data_Mem/n6318 ) );
  MUX U5066 ( .IN0(n1857), .IN1(o[1468]), .SEL(n2715), .F(\Data_Mem/n6317 ) );
  MUX U5067 ( .IN0(n1858), .IN1(o[1467]), .SEL(n2715), .F(\Data_Mem/n6316 ) );
  MUX U5068 ( .IN0(n1859), .IN1(o[1466]), .SEL(n2715), .F(\Data_Mem/n6315 ) );
  MUX U5069 ( .IN0(n1860), .IN1(o[1465]), .SEL(n2715), .F(\Data_Mem/n6314 ) );
  MUX U5070 ( .IN0(n1861), .IN1(o[1464]), .SEL(n2715), .F(\Data_Mem/n6313 ) );
  ANDN U5071 ( .A(n2716), .B(n2717), .Z(n2715) );
  AND U5072 ( .A(n2718), .B(n2719), .Z(n2716) );
  OR U5073 ( .A(n1867), .B(n2720), .Z(n2719) );
  MUX U5074 ( .IN0(n1868), .IN1(o[1463]), .SEL(n2721), .F(\Data_Mem/n6312 ) );
  MUX U5075 ( .IN0(n1870), .IN1(o[1462]), .SEL(n2721), .F(\Data_Mem/n6311 ) );
  MUX U5076 ( .IN0(n1871), .IN1(o[1461]), .SEL(n2721), .F(\Data_Mem/n6310 ) );
  MUX U5077 ( .IN0(n1872), .IN1(o[1460]), .SEL(n2721), .F(\Data_Mem/n6309 ) );
  MUX U5078 ( .IN0(n1873), .IN1(o[1459]), .SEL(n2721), .F(\Data_Mem/n6308 ) );
  IV U5079 ( .A(n2722), .Z(n2721) );
  MUX U5080 ( .IN0(o[1458]), .IN1(n1875), .SEL(n2722), .F(\Data_Mem/n6307 ) );
  MUX U5081 ( .IN0(o[1457]), .IN1(n1876), .SEL(n2722), .F(\Data_Mem/n6306 ) );
  MUX U5082 ( .IN0(o[1456]), .IN1(n1877), .SEL(n2722), .F(\Data_Mem/n6305 ) );
  NAND U5083 ( .A(n2723), .B(n2724), .Z(n2722) );
  OR U5084 ( .A(n1880), .B(n2720), .Z(n2724) );
  ANDN U5085 ( .A(n2718), .B(n2717), .Z(n2723) );
  NANDN U5086 ( .B(n2720), .A(n1915), .Z(n2718) );
  MUX U5087 ( .IN0(n1883), .IN1(o[1455]), .SEL(n2725), .F(\Data_Mem/n6304 ) );
  MUX U5088 ( .IN0(n1885), .IN1(o[1454]), .SEL(n2725), .F(\Data_Mem/n6303 ) );
  MUX U5089 ( .IN0(n1886), .IN1(o[1453]), .SEL(n2725), .F(\Data_Mem/n6302 ) );
  MUX U5090 ( .IN0(n1887), .IN1(o[1452]), .SEL(n2725), .F(\Data_Mem/n6301 ) );
  MUX U5091 ( .IN0(n1888), .IN1(o[1451]), .SEL(n2725), .F(\Data_Mem/n6300 ) );
  IV U5092 ( .A(n2726), .Z(n2725) );
  MUX U5093 ( .IN0(o[1450]), .IN1(n1890), .SEL(n2726), .F(\Data_Mem/n6299 ) );
  MUX U5094 ( .IN0(o[1449]), .IN1(n1891), .SEL(n2726), .F(\Data_Mem/n6298 ) );
  MUX U5095 ( .IN0(o[1448]), .IN1(n1892), .SEL(n2726), .F(\Data_Mem/n6297 ) );
  NAND U5096 ( .A(n2727), .B(n2728), .Z(n2726) );
  OR U5097 ( .A(n1895), .B(n2720), .Z(n2728) );
  MUX U5098 ( .IN0(reg_target[7]), .IN1(o[1447]), .SEL(n2729), .F(
        \Data_Mem/n6296 ) );
  MUX U5099 ( .IN0(reg_target[6]), .IN1(o[1446]), .SEL(n2729), .F(
        \Data_Mem/n6295 ) );
  MUX U5100 ( .IN0(reg_target[5]), .IN1(o[1445]), .SEL(n2729), .F(
        \Data_Mem/n6294 ) );
  MUX U5101 ( .IN0(reg_target[4]), .IN1(o[1444]), .SEL(n2729), .F(
        \Data_Mem/n6293 ) );
  MUX U5102 ( .IN0(reg_target[3]), .IN1(o[1443]), .SEL(n2729), .F(
        \Data_Mem/n6292 ) );
  IV U5103 ( .A(n2730), .Z(n2729) );
  MUX U5104 ( .IN0(o[1442]), .IN1(reg_target[2]), .SEL(n2730), .F(
        \Data_Mem/n6291 ) );
  MUX U5105 ( .IN0(o[1441]), .IN1(reg_target[1]), .SEL(n2730), .F(
        \Data_Mem/n6290 ) );
  MUX U5106 ( .IN0(o[1440]), .IN1(reg_target[0]), .SEL(n2730), .F(
        \Data_Mem/n6289 ) );
  NAND U5107 ( .A(n2727), .B(n2731), .Z(n2730) );
  NANDN U5108 ( .B(n2720), .A(n1899), .Z(n2731) );
  ANDN U5109 ( .A(n2732), .B(n2717), .Z(n2727) );
  ANDN U5110 ( .A(n1902), .B(n2720), .Z(n2717) );
  NANDN U5111 ( .B(n2720), .A(n1924), .Z(n2732) );
  NAND U5112 ( .A(n2001), .B(n2642), .Z(n2720) );
  MUX U5113 ( .IN0(n1853), .IN1(o[1503]), .SEL(n2733), .F(\Data_Mem/n6288 ) );
  MUX U5114 ( .IN0(n1855), .IN1(o[1502]), .SEL(n2733), .F(\Data_Mem/n6287 ) );
  MUX U5115 ( .IN0(n1856), .IN1(o[1501]), .SEL(n2733), .F(\Data_Mem/n6286 ) );
  MUX U5116 ( .IN0(n1857), .IN1(o[1500]), .SEL(n2733), .F(\Data_Mem/n6285 ) );
  MUX U5117 ( .IN0(n1858), .IN1(o[1499]), .SEL(n2733), .F(\Data_Mem/n6284 ) );
  MUX U5118 ( .IN0(n1859), .IN1(o[1498]), .SEL(n2733), .F(\Data_Mem/n6283 ) );
  MUX U5119 ( .IN0(n1860), .IN1(o[1497]), .SEL(n2733), .F(\Data_Mem/n6282 ) );
  MUX U5120 ( .IN0(n1861), .IN1(o[1496]), .SEL(n2733), .F(\Data_Mem/n6281 ) );
  ANDN U5121 ( .A(n2734), .B(n2735), .Z(n2733) );
  AND U5122 ( .A(n2736), .B(n2737), .Z(n2734) );
  OR U5123 ( .A(n1867), .B(n2738), .Z(n2737) );
  MUX U5124 ( .IN0(n1868), .IN1(o[1495]), .SEL(n2739), .F(\Data_Mem/n6280 ) );
  MUX U5125 ( .IN0(n1870), .IN1(o[1494]), .SEL(n2739), .F(\Data_Mem/n6279 ) );
  MUX U5126 ( .IN0(n1871), .IN1(o[1493]), .SEL(n2739), .F(\Data_Mem/n6278 ) );
  MUX U5127 ( .IN0(n1872), .IN1(o[1492]), .SEL(n2739), .F(\Data_Mem/n6277 ) );
  MUX U5128 ( .IN0(n1873), .IN1(o[1491]), .SEL(n2739), .F(\Data_Mem/n6276 ) );
  IV U5129 ( .A(n2740), .Z(n2739) );
  MUX U5130 ( .IN0(o[1490]), .IN1(n1875), .SEL(n2740), .F(\Data_Mem/n6275 ) );
  MUX U5131 ( .IN0(o[1489]), .IN1(n1876), .SEL(n2740), .F(\Data_Mem/n6274 ) );
  MUX U5132 ( .IN0(o[1488]), .IN1(n1877), .SEL(n2740), .F(\Data_Mem/n6273 ) );
  NAND U5133 ( .A(n2741), .B(n2742), .Z(n2740) );
  OR U5134 ( .A(n1880), .B(n2738), .Z(n2742) );
  ANDN U5135 ( .A(n2736), .B(n2735), .Z(n2741) );
  NANDN U5136 ( .B(n2738), .A(n1915), .Z(n2736) );
  MUX U5137 ( .IN0(n1883), .IN1(o[1487]), .SEL(n2743), .F(\Data_Mem/n6272 ) );
  MUX U5138 ( .IN0(n1885), .IN1(o[1486]), .SEL(n2743), .F(\Data_Mem/n6271 ) );
  MUX U5139 ( .IN0(n1886), .IN1(o[1485]), .SEL(n2743), .F(\Data_Mem/n6270 ) );
  MUX U5140 ( .IN0(n1887), .IN1(o[1484]), .SEL(n2743), .F(\Data_Mem/n6269 ) );
  MUX U5141 ( .IN0(n1888), .IN1(o[1483]), .SEL(n2743), .F(\Data_Mem/n6268 ) );
  IV U5142 ( .A(n2744), .Z(n2743) );
  MUX U5143 ( .IN0(o[1482]), .IN1(n1890), .SEL(n2744), .F(\Data_Mem/n6267 ) );
  MUX U5144 ( .IN0(o[1481]), .IN1(n1891), .SEL(n2744), .F(\Data_Mem/n6266 ) );
  MUX U5145 ( .IN0(o[1480]), .IN1(n1892), .SEL(n2744), .F(\Data_Mem/n6265 ) );
  NAND U5146 ( .A(n2745), .B(n2746), .Z(n2744) );
  OR U5147 ( .A(n1895), .B(n2738), .Z(n2746) );
  MUX U5148 ( .IN0(reg_target[7]), .IN1(o[1479]), .SEL(n2747), .F(
        \Data_Mem/n6264 ) );
  MUX U5149 ( .IN0(reg_target[6]), .IN1(o[1478]), .SEL(n2747), .F(
        \Data_Mem/n6263 ) );
  MUX U5150 ( .IN0(reg_target[5]), .IN1(o[1477]), .SEL(n2747), .F(
        \Data_Mem/n6262 ) );
  MUX U5151 ( .IN0(reg_target[4]), .IN1(o[1476]), .SEL(n2747), .F(
        \Data_Mem/n6261 ) );
  MUX U5152 ( .IN0(reg_target[3]), .IN1(o[1475]), .SEL(n2747), .F(
        \Data_Mem/n6260 ) );
  IV U5153 ( .A(n2748), .Z(n2747) );
  MUX U5154 ( .IN0(o[1474]), .IN1(reg_target[2]), .SEL(n2748), .F(
        \Data_Mem/n6259 ) );
  MUX U5155 ( .IN0(o[1473]), .IN1(reg_target[1]), .SEL(n2748), .F(
        \Data_Mem/n6258 ) );
  MUX U5156 ( .IN0(o[1472]), .IN1(reg_target[0]), .SEL(n2748), .F(
        \Data_Mem/n6257 ) );
  NAND U5157 ( .A(n2745), .B(n2749), .Z(n2748) );
  NANDN U5158 ( .B(n2738), .A(n1899), .Z(n2749) );
  ANDN U5159 ( .A(n2750), .B(n2735), .Z(n2745) );
  ANDN U5160 ( .A(n1902), .B(n2738), .Z(n2735) );
  NANDN U5161 ( .B(n2738), .A(n1924), .Z(n2750) );
  NAND U5162 ( .A(n2020), .B(n2642), .Z(n2738) );
  MUX U5163 ( .IN0(n1853), .IN1(o[1535]), .SEL(n2751), .F(\Data_Mem/n6256 ) );
  MUX U5164 ( .IN0(n1855), .IN1(o[1534]), .SEL(n2751), .F(\Data_Mem/n6255 ) );
  MUX U5165 ( .IN0(n1856), .IN1(o[1533]), .SEL(n2751), .F(\Data_Mem/n6254 ) );
  MUX U5166 ( .IN0(n1857), .IN1(o[1532]), .SEL(n2751), .F(\Data_Mem/n6253 ) );
  MUX U5167 ( .IN0(n1858), .IN1(o[1531]), .SEL(n2751), .F(\Data_Mem/n6252 ) );
  MUX U5168 ( .IN0(n1859), .IN1(o[1530]), .SEL(n2751), .F(\Data_Mem/n6251 ) );
  MUX U5169 ( .IN0(n1860), .IN1(o[1529]), .SEL(n2751), .F(\Data_Mem/n6250 ) );
  MUX U5170 ( .IN0(n1861), .IN1(o[1528]), .SEL(n2751), .F(\Data_Mem/n6249 ) );
  ANDN U5171 ( .A(n2752), .B(n2753), .Z(n2751) );
  AND U5172 ( .A(n2754), .B(n2755), .Z(n2752) );
  OR U5173 ( .A(n1867), .B(n2756), .Z(n2755) );
  MUX U5174 ( .IN0(n1868), .IN1(o[1527]), .SEL(n2757), .F(\Data_Mem/n6248 ) );
  MUX U5175 ( .IN0(n1870), .IN1(o[1526]), .SEL(n2757), .F(\Data_Mem/n6247 ) );
  MUX U5176 ( .IN0(n1871), .IN1(o[1525]), .SEL(n2757), .F(\Data_Mem/n6246 ) );
  MUX U5177 ( .IN0(n1872), .IN1(o[1524]), .SEL(n2757), .F(\Data_Mem/n6245 ) );
  MUX U5178 ( .IN0(n1873), .IN1(o[1523]), .SEL(n2757), .F(\Data_Mem/n6244 ) );
  IV U5179 ( .A(n2758), .Z(n2757) );
  MUX U5180 ( .IN0(o[1522]), .IN1(n1875), .SEL(n2758), .F(\Data_Mem/n6243 ) );
  MUX U5181 ( .IN0(o[1521]), .IN1(n1876), .SEL(n2758), .F(\Data_Mem/n6242 ) );
  MUX U5182 ( .IN0(o[1520]), .IN1(n1877), .SEL(n2758), .F(\Data_Mem/n6241 ) );
  NAND U5183 ( .A(n2759), .B(n2760), .Z(n2758) );
  OR U5184 ( .A(n1880), .B(n2756), .Z(n2760) );
  ANDN U5185 ( .A(n2754), .B(n2753), .Z(n2759) );
  NANDN U5186 ( .B(n2756), .A(n1915), .Z(n2754) );
  MUX U5187 ( .IN0(n1883), .IN1(o[1519]), .SEL(n2761), .F(\Data_Mem/n6240 ) );
  MUX U5188 ( .IN0(n1885), .IN1(o[1518]), .SEL(n2761), .F(\Data_Mem/n6239 ) );
  MUX U5189 ( .IN0(n1886), .IN1(o[1517]), .SEL(n2761), .F(\Data_Mem/n6238 ) );
  MUX U5190 ( .IN0(n1887), .IN1(o[1516]), .SEL(n2761), .F(\Data_Mem/n6237 ) );
  MUX U5191 ( .IN0(n1888), .IN1(o[1515]), .SEL(n2761), .F(\Data_Mem/n6236 ) );
  IV U5192 ( .A(n2762), .Z(n2761) );
  MUX U5193 ( .IN0(o[1514]), .IN1(n1890), .SEL(n2762), .F(\Data_Mem/n6235 ) );
  MUX U5194 ( .IN0(o[1513]), .IN1(n1891), .SEL(n2762), .F(\Data_Mem/n6234 ) );
  MUX U5195 ( .IN0(o[1512]), .IN1(n1892), .SEL(n2762), .F(\Data_Mem/n6233 ) );
  NAND U5196 ( .A(n2763), .B(n2764), .Z(n2762) );
  OR U5197 ( .A(n1895), .B(n2756), .Z(n2764) );
  MUX U5198 ( .IN0(reg_target[7]), .IN1(o[1511]), .SEL(n2765), .F(
        \Data_Mem/n6232 ) );
  MUX U5199 ( .IN0(reg_target[6]), .IN1(o[1510]), .SEL(n2765), .F(
        \Data_Mem/n6231 ) );
  MUX U5200 ( .IN0(reg_target[5]), .IN1(o[1509]), .SEL(n2765), .F(
        \Data_Mem/n6230 ) );
  MUX U5201 ( .IN0(reg_target[4]), .IN1(o[1508]), .SEL(n2765), .F(
        \Data_Mem/n6229 ) );
  MUX U5202 ( .IN0(reg_target[3]), .IN1(o[1507]), .SEL(n2765), .F(
        \Data_Mem/n6228 ) );
  IV U5203 ( .A(n2766), .Z(n2765) );
  MUX U5204 ( .IN0(o[1506]), .IN1(reg_target[2]), .SEL(n2766), .F(
        \Data_Mem/n6227 ) );
  MUX U5205 ( .IN0(o[1505]), .IN1(reg_target[1]), .SEL(n2766), .F(
        \Data_Mem/n6226 ) );
  MUX U5206 ( .IN0(o[1504]), .IN1(reg_target[0]), .SEL(n2766), .F(
        \Data_Mem/n6225 ) );
  NAND U5207 ( .A(n2763), .B(n2767), .Z(n2766) );
  NANDN U5208 ( .B(n2756), .A(n1899), .Z(n2767) );
  ANDN U5209 ( .A(n2768), .B(n2753), .Z(n2763) );
  ANDN U5210 ( .A(n1902), .B(n2756), .Z(n2753) );
  NANDN U5211 ( .B(n2756), .A(n1924), .Z(n2768) );
  NAND U5212 ( .A(n2642), .B(n2039), .Z(n2756) );
  ANDN U5213 ( .A(n2186), .B(n485), .Z(n2642) );
  AND U5214 ( .A(n511), .B(N26), .Z(n2186) );
  MUX U5215 ( .IN0(n1853), .IN1(o[1567]), .SEL(n2769), .F(\Data_Mem/n6224 ) );
  MUX U5216 ( .IN0(n1855), .IN1(o[1566]), .SEL(n2769), .F(\Data_Mem/n6223 ) );
  MUX U5217 ( .IN0(n1856), .IN1(o[1565]), .SEL(n2769), .F(\Data_Mem/n6222 ) );
  MUX U5218 ( .IN0(n1857), .IN1(o[1564]), .SEL(n2769), .F(\Data_Mem/n6221 ) );
  MUX U5219 ( .IN0(n1858), .IN1(o[1563]), .SEL(n2769), .F(\Data_Mem/n6220 ) );
  MUX U5220 ( .IN0(n1859), .IN1(o[1562]), .SEL(n2769), .F(\Data_Mem/n6219 ) );
  MUX U5221 ( .IN0(n1860), .IN1(o[1561]), .SEL(n2769), .F(\Data_Mem/n6218 ) );
  MUX U5222 ( .IN0(n1861), .IN1(o[1560]), .SEL(n2769), .F(\Data_Mem/n6217 ) );
  ANDN U5223 ( .A(n2770), .B(n2771), .Z(n2769) );
  AND U5224 ( .A(n2772), .B(n2773), .Z(n2770) );
  OR U5225 ( .A(n1867), .B(n2774), .Z(n2773) );
  MUX U5226 ( .IN0(n1868), .IN1(o[1559]), .SEL(n2775), .F(\Data_Mem/n6216 ) );
  MUX U5227 ( .IN0(n1870), .IN1(o[1558]), .SEL(n2775), .F(\Data_Mem/n6215 ) );
  MUX U5228 ( .IN0(n1871), .IN1(o[1557]), .SEL(n2775), .F(\Data_Mem/n6214 ) );
  MUX U5229 ( .IN0(n1872), .IN1(o[1556]), .SEL(n2775), .F(\Data_Mem/n6213 ) );
  MUX U5230 ( .IN0(n1873), .IN1(o[1555]), .SEL(n2775), .F(\Data_Mem/n6212 ) );
  IV U5231 ( .A(n2776), .Z(n2775) );
  MUX U5232 ( .IN0(o[1554]), .IN1(n1875), .SEL(n2776), .F(\Data_Mem/n6211 ) );
  MUX U5233 ( .IN0(o[1553]), .IN1(n1876), .SEL(n2776), .F(\Data_Mem/n6210 ) );
  MUX U5234 ( .IN0(o[1552]), .IN1(n1877), .SEL(n2776), .F(\Data_Mem/n6209 ) );
  NAND U5235 ( .A(n2777), .B(n2778), .Z(n2776) );
  OR U5236 ( .A(n1880), .B(n2774), .Z(n2778) );
  ANDN U5237 ( .A(n2772), .B(n2771), .Z(n2777) );
  NANDN U5238 ( .B(n2774), .A(n1915), .Z(n2772) );
  MUX U5239 ( .IN0(n1883), .IN1(o[1551]), .SEL(n2779), .F(\Data_Mem/n6208 ) );
  MUX U5240 ( .IN0(n1885), .IN1(o[1550]), .SEL(n2779), .F(\Data_Mem/n6207 ) );
  MUX U5241 ( .IN0(n1886), .IN1(o[1549]), .SEL(n2779), .F(\Data_Mem/n6206 ) );
  MUX U5242 ( .IN0(n1887), .IN1(o[1548]), .SEL(n2779), .F(\Data_Mem/n6205 ) );
  MUX U5243 ( .IN0(n1888), .IN1(o[1547]), .SEL(n2779), .F(\Data_Mem/n6204 ) );
  IV U5244 ( .A(n2780), .Z(n2779) );
  MUX U5245 ( .IN0(o[1546]), .IN1(n1890), .SEL(n2780), .F(\Data_Mem/n6203 ) );
  MUX U5246 ( .IN0(o[1545]), .IN1(n1891), .SEL(n2780), .F(\Data_Mem/n6202 ) );
  MUX U5247 ( .IN0(o[1544]), .IN1(n1892), .SEL(n2780), .F(\Data_Mem/n6201 ) );
  NAND U5248 ( .A(n2781), .B(n2782), .Z(n2780) );
  OR U5249 ( .A(n1895), .B(n2774), .Z(n2782) );
  MUX U5250 ( .IN0(reg_target[7]), .IN1(o[1543]), .SEL(n2783), .F(
        \Data_Mem/n6200 ) );
  MUX U5251 ( .IN0(reg_target[6]), .IN1(o[1542]), .SEL(n2783), .F(
        \Data_Mem/n6199 ) );
  MUX U5252 ( .IN0(reg_target[5]), .IN1(o[1541]), .SEL(n2783), .F(
        \Data_Mem/n6198 ) );
  MUX U5253 ( .IN0(reg_target[4]), .IN1(o[1540]), .SEL(n2783), .F(
        \Data_Mem/n6197 ) );
  MUX U5254 ( .IN0(reg_target[3]), .IN1(o[1539]), .SEL(n2783), .F(
        \Data_Mem/n6196 ) );
  IV U5255 ( .A(n2784), .Z(n2783) );
  MUX U5256 ( .IN0(o[1538]), .IN1(reg_target[2]), .SEL(n2784), .F(
        \Data_Mem/n6195 ) );
  MUX U5257 ( .IN0(o[1537]), .IN1(reg_target[1]), .SEL(n2784), .F(
        \Data_Mem/n6194 ) );
  MUX U5258 ( .IN0(o[1536]), .IN1(reg_target[0]), .SEL(n2784), .F(
        \Data_Mem/n6193 ) );
  NAND U5259 ( .A(n2781), .B(n2785), .Z(n2784) );
  NANDN U5260 ( .B(n2774), .A(n1899), .Z(n2785) );
  ANDN U5261 ( .A(n2786), .B(n2771), .Z(n2781) );
  ANDN U5262 ( .A(n1902), .B(n2774), .Z(n2771) );
  NANDN U5263 ( .B(n2774), .A(n1924), .Z(n2786) );
  NAND U5264 ( .A(n1903), .B(n2787), .Z(n2774) );
  MUX U5265 ( .IN0(n1853), .IN1(o[1599]), .SEL(n2788), .F(\Data_Mem/n6192 ) );
  MUX U5266 ( .IN0(n1855), .IN1(o[1598]), .SEL(n2788), .F(\Data_Mem/n6191 ) );
  MUX U5267 ( .IN0(n1856), .IN1(o[1597]), .SEL(n2788), .F(\Data_Mem/n6190 ) );
  MUX U5268 ( .IN0(n1857), .IN1(o[1596]), .SEL(n2788), .F(\Data_Mem/n6189 ) );
  MUX U5269 ( .IN0(n1858), .IN1(o[1595]), .SEL(n2788), .F(\Data_Mem/n6188 ) );
  MUX U5270 ( .IN0(n1859), .IN1(o[1594]), .SEL(n2788), .F(\Data_Mem/n6187 ) );
  MUX U5271 ( .IN0(n1860), .IN1(o[1593]), .SEL(n2788), .F(\Data_Mem/n6186 ) );
  MUX U5272 ( .IN0(n1861), .IN1(o[1592]), .SEL(n2788), .F(\Data_Mem/n6185 ) );
  ANDN U5273 ( .A(n2789), .B(n2790), .Z(n2788) );
  AND U5274 ( .A(n2791), .B(n2792), .Z(n2789) );
  OR U5275 ( .A(n1867), .B(n2793), .Z(n2792) );
  MUX U5276 ( .IN0(n1868), .IN1(o[1591]), .SEL(n2794), .F(\Data_Mem/n6184 ) );
  MUX U5277 ( .IN0(n1870), .IN1(o[1590]), .SEL(n2794), .F(\Data_Mem/n6183 ) );
  MUX U5278 ( .IN0(n1871), .IN1(o[1589]), .SEL(n2794), .F(\Data_Mem/n6182 ) );
  MUX U5279 ( .IN0(n1872), .IN1(o[1588]), .SEL(n2794), .F(\Data_Mem/n6181 ) );
  MUX U5280 ( .IN0(n1873), .IN1(o[1587]), .SEL(n2794), .F(\Data_Mem/n6180 ) );
  IV U5281 ( .A(n2795), .Z(n2794) );
  MUX U5282 ( .IN0(o[1586]), .IN1(n1875), .SEL(n2795), .F(\Data_Mem/n6179 ) );
  MUX U5283 ( .IN0(o[1585]), .IN1(n1876), .SEL(n2795), .F(\Data_Mem/n6178 ) );
  MUX U5284 ( .IN0(o[1584]), .IN1(n1877), .SEL(n2795), .F(\Data_Mem/n6177 ) );
  NAND U5285 ( .A(n2796), .B(n2797), .Z(n2795) );
  OR U5286 ( .A(n1880), .B(n2793), .Z(n2797) );
  ANDN U5287 ( .A(n2791), .B(n2790), .Z(n2796) );
  NANDN U5288 ( .B(n2793), .A(n1915), .Z(n2791) );
  MUX U5289 ( .IN0(n1883), .IN1(o[1583]), .SEL(n2798), .F(\Data_Mem/n6176 ) );
  MUX U5290 ( .IN0(n1885), .IN1(o[1582]), .SEL(n2798), .F(\Data_Mem/n6175 ) );
  MUX U5291 ( .IN0(n1886), .IN1(o[1581]), .SEL(n2798), .F(\Data_Mem/n6174 ) );
  MUX U5292 ( .IN0(n1887), .IN1(o[1580]), .SEL(n2798), .F(\Data_Mem/n6173 ) );
  MUX U5293 ( .IN0(n1888), .IN1(o[1579]), .SEL(n2798), .F(\Data_Mem/n6172 ) );
  IV U5294 ( .A(n2799), .Z(n2798) );
  MUX U5295 ( .IN0(o[1578]), .IN1(n1890), .SEL(n2799), .F(\Data_Mem/n6171 ) );
  MUX U5296 ( .IN0(o[1577]), .IN1(n1891), .SEL(n2799), .F(\Data_Mem/n6170 ) );
  MUX U5297 ( .IN0(o[1576]), .IN1(n1892), .SEL(n2799), .F(\Data_Mem/n6169 ) );
  NAND U5298 ( .A(n2800), .B(n2801), .Z(n2799) );
  OR U5299 ( .A(n1895), .B(n2793), .Z(n2801) );
  MUX U5300 ( .IN0(reg_target[7]), .IN1(o[1575]), .SEL(n2802), .F(
        \Data_Mem/n6168 ) );
  MUX U5301 ( .IN0(reg_target[6]), .IN1(o[1574]), .SEL(n2802), .F(
        \Data_Mem/n6167 ) );
  MUX U5302 ( .IN0(reg_target[5]), .IN1(o[1573]), .SEL(n2802), .F(
        \Data_Mem/n6166 ) );
  MUX U5303 ( .IN0(reg_target[4]), .IN1(o[1572]), .SEL(n2802), .F(
        \Data_Mem/n6165 ) );
  MUX U5304 ( .IN0(reg_target[3]), .IN1(o[1571]), .SEL(n2802), .F(
        \Data_Mem/n6164 ) );
  IV U5305 ( .A(n2803), .Z(n2802) );
  MUX U5306 ( .IN0(o[1570]), .IN1(reg_target[2]), .SEL(n2803), .F(
        \Data_Mem/n6163 ) );
  MUX U5307 ( .IN0(o[1569]), .IN1(reg_target[1]), .SEL(n2803), .F(
        \Data_Mem/n6162 ) );
  MUX U5308 ( .IN0(o[1568]), .IN1(reg_target[0]), .SEL(n2803), .F(
        \Data_Mem/n6161 ) );
  NAND U5309 ( .A(n2800), .B(n2804), .Z(n2803) );
  NANDN U5310 ( .B(n2793), .A(n1899), .Z(n2804) );
  ANDN U5311 ( .A(n2805), .B(n2790), .Z(n2800) );
  ANDN U5312 ( .A(n1902), .B(n2793), .Z(n2790) );
  NANDN U5313 ( .B(n2793), .A(n1924), .Z(n2805) );
  NAND U5314 ( .A(n1925), .B(n2787), .Z(n2793) );
  MUX U5315 ( .IN0(n1853), .IN1(o[1631]), .SEL(n2806), .F(\Data_Mem/n6160 ) );
  MUX U5316 ( .IN0(n1855), .IN1(o[1630]), .SEL(n2806), .F(\Data_Mem/n6159 ) );
  MUX U5317 ( .IN0(n1856), .IN1(o[1629]), .SEL(n2806), .F(\Data_Mem/n6158 ) );
  MUX U5318 ( .IN0(n1857), .IN1(o[1628]), .SEL(n2806), .F(\Data_Mem/n6157 ) );
  MUX U5319 ( .IN0(n1858), .IN1(o[1627]), .SEL(n2806), .F(\Data_Mem/n6156 ) );
  MUX U5320 ( .IN0(n1859), .IN1(o[1626]), .SEL(n2806), .F(\Data_Mem/n6155 ) );
  MUX U5321 ( .IN0(n1860), .IN1(o[1625]), .SEL(n2806), .F(\Data_Mem/n6154 ) );
  MUX U5322 ( .IN0(n1861), .IN1(o[1624]), .SEL(n2806), .F(\Data_Mem/n6153 ) );
  ANDN U5323 ( .A(n2807), .B(n2808), .Z(n2806) );
  AND U5324 ( .A(n2809), .B(n2810), .Z(n2807) );
  OR U5325 ( .A(n1867), .B(n2811), .Z(n2810) );
  MUX U5326 ( .IN0(n1868), .IN1(o[1623]), .SEL(n2812), .F(\Data_Mem/n6152 ) );
  MUX U5327 ( .IN0(n1870), .IN1(o[1622]), .SEL(n2812), .F(\Data_Mem/n6151 ) );
  MUX U5328 ( .IN0(n1871), .IN1(o[1621]), .SEL(n2812), .F(\Data_Mem/n6150 ) );
  MUX U5329 ( .IN0(n1872), .IN1(o[1620]), .SEL(n2812), .F(\Data_Mem/n6149 ) );
  MUX U5330 ( .IN0(n1873), .IN1(o[1619]), .SEL(n2812), .F(\Data_Mem/n6148 ) );
  IV U5331 ( .A(n2813), .Z(n2812) );
  MUX U5332 ( .IN0(o[1618]), .IN1(n1875), .SEL(n2813), .F(\Data_Mem/n6147 ) );
  MUX U5333 ( .IN0(o[1617]), .IN1(n1876), .SEL(n2813), .F(\Data_Mem/n6146 ) );
  MUX U5334 ( .IN0(o[1616]), .IN1(n1877), .SEL(n2813), .F(\Data_Mem/n6145 ) );
  NAND U5335 ( .A(n2814), .B(n2815), .Z(n2813) );
  OR U5336 ( .A(n1880), .B(n2811), .Z(n2815) );
  ANDN U5337 ( .A(n2809), .B(n2808), .Z(n2814) );
  NANDN U5338 ( .B(n2811), .A(n1915), .Z(n2809) );
  MUX U5339 ( .IN0(n1883), .IN1(o[1615]), .SEL(n2816), .F(\Data_Mem/n6144 ) );
  MUX U5340 ( .IN0(n1885), .IN1(o[1614]), .SEL(n2816), .F(\Data_Mem/n6143 ) );
  MUX U5341 ( .IN0(n1886), .IN1(o[1613]), .SEL(n2816), .F(\Data_Mem/n6142 ) );
  MUX U5342 ( .IN0(n1887), .IN1(o[1612]), .SEL(n2816), .F(\Data_Mem/n6141 ) );
  MUX U5343 ( .IN0(n1888), .IN1(o[1611]), .SEL(n2816), .F(\Data_Mem/n6140 ) );
  IV U5344 ( .A(n2817), .Z(n2816) );
  MUX U5345 ( .IN0(o[1610]), .IN1(n1890), .SEL(n2817), .F(\Data_Mem/n6139 ) );
  MUX U5346 ( .IN0(o[1609]), .IN1(n1891), .SEL(n2817), .F(\Data_Mem/n6138 ) );
  MUX U5347 ( .IN0(o[1608]), .IN1(n1892), .SEL(n2817), .F(\Data_Mem/n6137 ) );
  NAND U5348 ( .A(n2818), .B(n2819), .Z(n2817) );
  OR U5349 ( .A(n1895), .B(n2811), .Z(n2819) );
  MUX U5350 ( .IN0(reg_target[7]), .IN1(o[1607]), .SEL(n2820), .F(
        \Data_Mem/n6136 ) );
  MUX U5351 ( .IN0(reg_target[6]), .IN1(o[1606]), .SEL(n2820), .F(
        \Data_Mem/n6135 ) );
  MUX U5352 ( .IN0(reg_target[5]), .IN1(o[1605]), .SEL(n2820), .F(
        \Data_Mem/n6134 ) );
  MUX U5353 ( .IN0(reg_target[4]), .IN1(o[1604]), .SEL(n2820), .F(
        \Data_Mem/n6133 ) );
  MUX U5354 ( .IN0(reg_target[3]), .IN1(o[1603]), .SEL(n2820), .F(
        \Data_Mem/n6132 ) );
  IV U5355 ( .A(n2821), .Z(n2820) );
  MUX U5356 ( .IN0(o[1602]), .IN1(reg_target[2]), .SEL(n2821), .F(
        \Data_Mem/n6131 ) );
  MUX U5357 ( .IN0(o[1601]), .IN1(reg_target[1]), .SEL(n2821), .F(
        \Data_Mem/n6130 ) );
  MUX U5358 ( .IN0(o[1600]), .IN1(reg_target[0]), .SEL(n2821), .F(
        \Data_Mem/n6129 ) );
  NAND U5359 ( .A(n2818), .B(n2822), .Z(n2821) );
  NANDN U5360 ( .B(n2811), .A(n1899), .Z(n2822) );
  ANDN U5361 ( .A(n2823), .B(n2808), .Z(n2818) );
  ANDN U5362 ( .A(n1902), .B(n2811), .Z(n2808) );
  NANDN U5363 ( .B(n2811), .A(n1924), .Z(n2823) );
  NAND U5364 ( .A(n1944), .B(n2787), .Z(n2811) );
  MUX U5365 ( .IN0(n1853), .IN1(o[1663]), .SEL(n2824), .F(\Data_Mem/n6128 ) );
  MUX U5366 ( .IN0(n1855), .IN1(o[1662]), .SEL(n2824), .F(\Data_Mem/n6127 ) );
  MUX U5367 ( .IN0(n1856), .IN1(o[1661]), .SEL(n2824), .F(\Data_Mem/n6126 ) );
  MUX U5368 ( .IN0(n1857), .IN1(o[1660]), .SEL(n2824), .F(\Data_Mem/n6125 ) );
  MUX U5369 ( .IN0(n1858), .IN1(o[1659]), .SEL(n2824), .F(\Data_Mem/n6124 ) );
  MUX U5370 ( .IN0(n1859), .IN1(o[1658]), .SEL(n2824), .F(\Data_Mem/n6123 ) );
  MUX U5371 ( .IN0(n1860), .IN1(o[1657]), .SEL(n2824), .F(\Data_Mem/n6122 ) );
  MUX U5372 ( .IN0(n1861), .IN1(o[1656]), .SEL(n2824), .F(\Data_Mem/n6121 ) );
  ANDN U5373 ( .A(n2825), .B(n2826), .Z(n2824) );
  AND U5374 ( .A(n2827), .B(n2828), .Z(n2825) );
  OR U5375 ( .A(n1867), .B(n2829), .Z(n2828) );
  MUX U5376 ( .IN0(n1868), .IN1(o[1655]), .SEL(n2830), .F(\Data_Mem/n6120 ) );
  MUX U5377 ( .IN0(n1870), .IN1(o[1654]), .SEL(n2830), .F(\Data_Mem/n6119 ) );
  MUX U5378 ( .IN0(n1871), .IN1(o[1653]), .SEL(n2830), .F(\Data_Mem/n6118 ) );
  MUX U5379 ( .IN0(n1872), .IN1(o[1652]), .SEL(n2830), .F(\Data_Mem/n6117 ) );
  MUX U5380 ( .IN0(n1873), .IN1(o[1651]), .SEL(n2830), .F(\Data_Mem/n6116 ) );
  IV U5381 ( .A(n2831), .Z(n2830) );
  MUX U5382 ( .IN0(o[1650]), .IN1(n1875), .SEL(n2831), .F(\Data_Mem/n6115 ) );
  MUX U5383 ( .IN0(o[1649]), .IN1(n1876), .SEL(n2831), .F(\Data_Mem/n6114 ) );
  MUX U5384 ( .IN0(o[1648]), .IN1(n1877), .SEL(n2831), .F(\Data_Mem/n6113 ) );
  NAND U5385 ( .A(n2832), .B(n2833), .Z(n2831) );
  OR U5386 ( .A(n1880), .B(n2829), .Z(n2833) );
  ANDN U5387 ( .A(n2827), .B(n2826), .Z(n2832) );
  NANDN U5388 ( .B(n2829), .A(n1915), .Z(n2827) );
  MUX U5389 ( .IN0(n1883), .IN1(o[1647]), .SEL(n2834), .F(\Data_Mem/n6112 ) );
  MUX U5390 ( .IN0(n1885), .IN1(o[1646]), .SEL(n2834), .F(\Data_Mem/n6111 ) );
  MUX U5391 ( .IN0(n1886), .IN1(o[1645]), .SEL(n2834), .F(\Data_Mem/n6110 ) );
  MUX U5392 ( .IN0(n1887), .IN1(o[1644]), .SEL(n2834), .F(\Data_Mem/n6109 ) );
  MUX U5393 ( .IN0(n1888), .IN1(o[1643]), .SEL(n2834), .F(\Data_Mem/n6108 ) );
  IV U5394 ( .A(n2835), .Z(n2834) );
  MUX U5395 ( .IN0(o[1642]), .IN1(n1890), .SEL(n2835), .F(\Data_Mem/n6107 ) );
  MUX U5396 ( .IN0(o[1641]), .IN1(n1891), .SEL(n2835), .F(\Data_Mem/n6106 ) );
  MUX U5397 ( .IN0(o[1640]), .IN1(n1892), .SEL(n2835), .F(\Data_Mem/n6105 ) );
  NAND U5398 ( .A(n2836), .B(n2837), .Z(n2835) );
  OR U5399 ( .A(n1895), .B(n2829), .Z(n2837) );
  MUX U5400 ( .IN0(reg_target[7]), .IN1(o[1639]), .SEL(n2838), .F(
        \Data_Mem/n6104 ) );
  MUX U5401 ( .IN0(reg_target[6]), .IN1(o[1638]), .SEL(n2838), .F(
        \Data_Mem/n6103 ) );
  MUX U5402 ( .IN0(reg_target[5]), .IN1(o[1637]), .SEL(n2838), .F(
        \Data_Mem/n6102 ) );
  MUX U5403 ( .IN0(reg_target[4]), .IN1(o[1636]), .SEL(n2838), .F(
        \Data_Mem/n6101 ) );
  MUX U5404 ( .IN0(reg_target[3]), .IN1(o[1635]), .SEL(n2838), .F(
        \Data_Mem/n6100 ) );
  IV U5405 ( .A(n2839), .Z(n2838) );
  MUX U5406 ( .IN0(o[1634]), .IN1(reg_target[2]), .SEL(n2839), .F(
        \Data_Mem/n6099 ) );
  MUX U5407 ( .IN0(o[1633]), .IN1(reg_target[1]), .SEL(n2839), .F(
        \Data_Mem/n6098 ) );
  MUX U5408 ( .IN0(o[1632]), .IN1(reg_target[0]), .SEL(n2839), .F(
        \Data_Mem/n6097 ) );
  NAND U5409 ( .A(n2836), .B(n2840), .Z(n2839) );
  NANDN U5410 ( .B(n2829), .A(n1899), .Z(n2840) );
  ANDN U5411 ( .A(n2841), .B(n2826), .Z(n2836) );
  ANDN U5412 ( .A(n1902), .B(n2829), .Z(n2826) );
  NANDN U5413 ( .B(n2829), .A(n1924), .Z(n2841) );
  NAND U5414 ( .A(n1963), .B(n2787), .Z(n2829) );
  MUX U5415 ( .IN0(n1853), .IN1(o[1695]), .SEL(n2842), .F(\Data_Mem/n6096 ) );
  MUX U5416 ( .IN0(n1855), .IN1(o[1694]), .SEL(n2842), .F(\Data_Mem/n6095 ) );
  MUX U5417 ( .IN0(n1856), .IN1(o[1693]), .SEL(n2842), .F(\Data_Mem/n6094 ) );
  MUX U5418 ( .IN0(n1857), .IN1(o[1692]), .SEL(n2842), .F(\Data_Mem/n6093 ) );
  MUX U5419 ( .IN0(n1858), .IN1(o[1691]), .SEL(n2842), .F(\Data_Mem/n6092 ) );
  MUX U5420 ( .IN0(n1859), .IN1(o[1690]), .SEL(n2842), .F(\Data_Mem/n6091 ) );
  MUX U5421 ( .IN0(n1860), .IN1(o[1689]), .SEL(n2842), .F(\Data_Mem/n6090 ) );
  MUX U5422 ( .IN0(n1861), .IN1(o[1688]), .SEL(n2842), .F(\Data_Mem/n6089 ) );
  ANDN U5423 ( .A(n2843), .B(n2844), .Z(n2842) );
  AND U5424 ( .A(n2845), .B(n2846), .Z(n2843) );
  OR U5425 ( .A(n1867), .B(n2847), .Z(n2846) );
  MUX U5426 ( .IN0(n1868), .IN1(o[1687]), .SEL(n2848), .F(\Data_Mem/n6088 ) );
  MUX U5427 ( .IN0(n1870), .IN1(o[1686]), .SEL(n2848), .F(\Data_Mem/n6087 ) );
  MUX U5428 ( .IN0(n1871), .IN1(o[1685]), .SEL(n2848), .F(\Data_Mem/n6086 ) );
  MUX U5429 ( .IN0(n1872), .IN1(o[1684]), .SEL(n2848), .F(\Data_Mem/n6085 ) );
  MUX U5430 ( .IN0(n1873), .IN1(o[1683]), .SEL(n2848), .F(\Data_Mem/n6084 ) );
  IV U5431 ( .A(n2849), .Z(n2848) );
  MUX U5432 ( .IN0(o[1682]), .IN1(n1875), .SEL(n2849), .F(\Data_Mem/n6083 ) );
  MUX U5433 ( .IN0(o[1681]), .IN1(n1876), .SEL(n2849), .F(\Data_Mem/n6082 ) );
  MUX U5434 ( .IN0(o[1680]), .IN1(n1877), .SEL(n2849), .F(\Data_Mem/n6081 ) );
  NAND U5435 ( .A(n2850), .B(n2851), .Z(n2849) );
  OR U5436 ( .A(n1880), .B(n2847), .Z(n2851) );
  ANDN U5437 ( .A(n2845), .B(n2844), .Z(n2850) );
  NANDN U5438 ( .B(n2847), .A(n1915), .Z(n2845) );
  MUX U5439 ( .IN0(n1883), .IN1(o[1679]), .SEL(n2852), .F(\Data_Mem/n6080 ) );
  MUX U5440 ( .IN0(n1885), .IN1(o[1678]), .SEL(n2852), .F(\Data_Mem/n6079 ) );
  MUX U5441 ( .IN0(n1886), .IN1(o[1677]), .SEL(n2852), .F(\Data_Mem/n6078 ) );
  MUX U5442 ( .IN0(n1887), .IN1(o[1676]), .SEL(n2852), .F(\Data_Mem/n6077 ) );
  MUX U5443 ( .IN0(n1888), .IN1(o[1675]), .SEL(n2852), .F(\Data_Mem/n6076 ) );
  IV U5444 ( .A(n2853), .Z(n2852) );
  MUX U5445 ( .IN0(o[1674]), .IN1(n1890), .SEL(n2853), .F(\Data_Mem/n6075 ) );
  MUX U5446 ( .IN0(o[1673]), .IN1(n1891), .SEL(n2853), .F(\Data_Mem/n6074 ) );
  MUX U5447 ( .IN0(o[1672]), .IN1(n1892), .SEL(n2853), .F(\Data_Mem/n6073 ) );
  NAND U5448 ( .A(n2854), .B(n2855), .Z(n2853) );
  OR U5449 ( .A(n1895), .B(n2847), .Z(n2855) );
  MUX U5450 ( .IN0(reg_target[7]), .IN1(o[1671]), .SEL(n2856), .F(
        \Data_Mem/n6072 ) );
  MUX U5451 ( .IN0(reg_target[6]), .IN1(o[1670]), .SEL(n2856), .F(
        \Data_Mem/n6071 ) );
  MUX U5452 ( .IN0(reg_target[5]), .IN1(o[1669]), .SEL(n2856), .F(
        \Data_Mem/n6070 ) );
  MUX U5453 ( .IN0(reg_target[4]), .IN1(o[1668]), .SEL(n2856), .F(
        \Data_Mem/n6069 ) );
  MUX U5454 ( .IN0(reg_target[3]), .IN1(o[1667]), .SEL(n2856), .F(
        \Data_Mem/n6068 ) );
  IV U5455 ( .A(n2857), .Z(n2856) );
  MUX U5456 ( .IN0(o[1666]), .IN1(reg_target[2]), .SEL(n2857), .F(
        \Data_Mem/n6067 ) );
  MUX U5457 ( .IN0(o[1665]), .IN1(reg_target[1]), .SEL(n2857), .F(
        \Data_Mem/n6066 ) );
  MUX U5458 ( .IN0(o[1664]), .IN1(reg_target[0]), .SEL(n2857), .F(
        \Data_Mem/n6065 ) );
  NAND U5459 ( .A(n2854), .B(n2858), .Z(n2857) );
  NANDN U5460 ( .B(n2847), .A(n1899), .Z(n2858) );
  ANDN U5461 ( .A(n2859), .B(n2844), .Z(n2854) );
  ANDN U5462 ( .A(n1902), .B(n2847), .Z(n2844) );
  NANDN U5463 ( .B(n2847), .A(n1924), .Z(n2859) );
  NAND U5464 ( .A(n1982), .B(n2787), .Z(n2847) );
  MUX U5465 ( .IN0(n1853), .IN1(o[1727]), .SEL(n2860), .F(\Data_Mem/n6064 ) );
  MUX U5466 ( .IN0(n1855), .IN1(o[1726]), .SEL(n2860), .F(\Data_Mem/n6063 ) );
  MUX U5467 ( .IN0(n1856), .IN1(o[1725]), .SEL(n2860), .F(\Data_Mem/n6062 ) );
  MUX U5468 ( .IN0(n1857), .IN1(o[1724]), .SEL(n2860), .F(\Data_Mem/n6061 ) );
  MUX U5469 ( .IN0(n1858), .IN1(o[1723]), .SEL(n2860), .F(\Data_Mem/n6060 ) );
  MUX U5470 ( .IN0(n1859), .IN1(o[1722]), .SEL(n2860), .F(\Data_Mem/n6059 ) );
  MUX U5471 ( .IN0(n1860), .IN1(o[1721]), .SEL(n2860), .F(\Data_Mem/n6058 ) );
  MUX U5472 ( .IN0(n1861), .IN1(o[1720]), .SEL(n2860), .F(\Data_Mem/n6057 ) );
  ANDN U5473 ( .A(n2861), .B(n2862), .Z(n2860) );
  AND U5474 ( .A(n2863), .B(n2864), .Z(n2861) );
  OR U5475 ( .A(n1867), .B(n2865), .Z(n2864) );
  MUX U5476 ( .IN0(n1868), .IN1(o[1719]), .SEL(n2866), .F(\Data_Mem/n6056 ) );
  MUX U5477 ( .IN0(n1870), .IN1(o[1718]), .SEL(n2866), .F(\Data_Mem/n6055 ) );
  MUX U5478 ( .IN0(n1871), .IN1(o[1717]), .SEL(n2866), .F(\Data_Mem/n6054 ) );
  MUX U5479 ( .IN0(n1872), .IN1(o[1716]), .SEL(n2866), .F(\Data_Mem/n6053 ) );
  MUX U5480 ( .IN0(n1873), .IN1(o[1715]), .SEL(n2866), .F(\Data_Mem/n6052 ) );
  IV U5481 ( .A(n2867), .Z(n2866) );
  MUX U5482 ( .IN0(o[1714]), .IN1(n1875), .SEL(n2867), .F(\Data_Mem/n6051 ) );
  MUX U5483 ( .IN0(o[1713]), .IN1(n1876), .SEL(n2867), .F(\Data_Mem/n6050 ) );
  MUX U5484 ( .IN0(o[1712]), .IN1(n1877), .SEL(n2867), .F(\Data_Mem/n6049 ) );
  NAND U5485 ( .A(n2868), .B(n2869), .Z(n2867) );
  OR U5486 ( .A(n1880), .B(n2865), .Z(n2869) );
  ANDN U5487 ( .A(n2863), .B(n2862), .Z(n2868) );
  NANDN U5488 ( .B(n2865), .A(n1915), .Z(n2863) );
  MUX U5489 ( .IN0(n1883), .IN1(o[1711]), .SEL(n2870), .F(\Data_Mem/n6048 ) );
  MUX U5490 ( .IN0(n1885), .IN1(o[1710]), .SEL(n2870), .F(\Data_Mem/n6047 ) );
  MUX U5491 ( .IN0(n1886), .IN1(o[1709]), .SEL(n2870), .F(\Data_Mem/n6046 ) );
  MUX U5492 ( .IN0(n1887), .IN1(o[1708]), .SEL(n2870), .F(\Data_Mem/n6045 ) );
  MUX U5493 ( .IN0(n1888), .IN1(o[1707]), .SEL(n2870), .F(\Data_Mem/n6044 ) );
  IV U5494 ( .A(n2871), .Z(n2870) );
  MUX U5495 ( .IN0(o[1706]), .IN1(n1890), .SEL(n2871), .F(\Data_Mem/n6043 ) );
  MUX U5496 ( .IN0(o[1705]), .IN1(n1891), .SEL(n2871), .F(\Data_Mem/n6042 ) );
  MUX U5497 ( .IN0(o[1704]), .IN1(n1892), .SEL(n2871), .F(\Data_Mem/n6041 ) );
  NAND U5498 ( .A(n2872), .B(n2873), .Z(n2871) );
  OR U5499 ( .A(n1895), .B(n2865), .Z(n2873) );
  MUX U5500 ( .IN0(reg_target[7]), .IN1(o[1703]), .SEL(n2874), .F(
        \Data_Mem/n6040 ) );
  MUX U5501 ( .IN0(reg_target[6]), .IN1(o[1702]), .SEL(n2874), .F(
        \Data_Mem/n6039 ) );
  MUX U5502 ( .IN0(reg_target[5]), .IN1(o[1701]), .SEL(n2874), .F(
        \Data_Mem/n6038 ) );
  MUX U5503 ( .IN0(reg_target[4]), .IN1(o[1700]), .SEL(n2874), .F(
        \Data_Mem/n6037 ) );
  MUX U5504 ( .IN0(reg_target[3]), .IN1(o[1699]), .SEL(n2874), .F(
        \Data_Mem/n6036 ) );
  IV U5505 ( .A(n2875), .Z(n2874) );
  MUX U5506 ( .IN0(o[1698]), .IN1(reg_target[2]), .SEL(n2875), .F(
        \Data_Mem/n6035 ) );
  MUX U5507 ( .IN0(o[1697]), .IN1(reg_target[1]), .SEL(n2875), .F(
        \Data_Mem/n6034 ) );
  MUX U5508 ( .IN0(o[1696]), .IN1(reg_target[0]), .SEL(n2875), .F(
        \Data_Mem/n6033 ) );
  NAND U5509 ( .A(n2872), .B(n2876), .Z(n2875) );
  NANDN U5510 ( .B(n2865), .A(n1899), .Z(n2876) );
  ANDN U5511 ( .A(n2877), .B(n2862), .Z(n2872) );
  ANDN U5512 ( .A(n1902), .B(n2865), .Z(n2862) );
  NANDN U5513 ( .B(n2865), .A(n1924), .Z(n2877) );
  NAND U5514 ( .A(n2001), .B(n2787), .Z(n2865) );
  MUX U5515 ( .IN0(n1853), .IN1(o[1759]), .SEL(n2878), .F(\Data_Mem/n6032 ) );
  MUX U5516 ( .IN0(n1855), .IN1(o[1758]), .SEL(n2878), .F(\Data_Mem/n6031 ) );
  MUX U5517 ( .IN0(n1856), .IN1(o[1757]), .SEL(n2878), .F(\Data_Mem/n6030 ) );
  MUX U5518 ( .IN0(n1857), .IN1(o[1756]), .SEL(n2878), .F(\Data_Mem/n6029 ) );
  MUX U5519 ( .IN0(n1858), .IN1(o[1755]), .SEL(n2878), .F(\Data_Mem/n6028 ) );
  MUX U5520 ( .IN0(n1859), .IN1(o[1754]), .SEL(n2878), .F(\Data_Mem/n6027 ) );
  MUX U5521 ( .IN0(n1860), .IN1(o[1753]), .SEL(n2878), .F(\Data_Mem/n6026 ) );
  MUX U5522 ( .IN0(n1861), .IN1(o[1752]), .SEL(n2878), .F(\Data_Mem/n6025 ) );
  ANDN U5523 ( .A(n2879), .B(n2880), .Z(n2878) );
  AND U5524 ( .A(n2881), .B(n2882), .Z(n2879) );
  OR U5525 ( .A(n1867), .B(n2883), .Z(n2882) );
  MUX U5526 ( .IN0(n1868), .IN1(o[1751]), .SEL(n2884), .F(\Data_Mem/n6024 ) );
  MUX U5527 ( .IN0(n1870), .IN1(o[1750]), .SEL(n2884), .F(\Data_Mem/n6023 ) );
  MUX U5528 ( .IN0(n1871), .IN1(o[1749]), .SEL(n2884), .F(\Data_Mem/n6022 ) );
  MUX U5529 ( .IN0(n1872), .IN1(o[1748]), .SEL(n2884), .F(\Data_Mem/n6021 ) );
  MUX U5530 ( .IN0(n1873), .IN1(o[1747]), .SEL(n2884), .F(\Data_Mem/n6020 ) );
  IV U5531 ( .A(n2885), .Z(n2884) );
  MUX U5532 ( .IN0(o[1746]), .IN1(n1875), .SEL(n2885), .F(\Data_Mem/n6019 ) );
  MUX U5533 ( .IN0(o[1745]), .IN1(n1876), .SEL(n2885), .F(\Data_Mem/n6018 ) );
  MUX U5534 ( .IN0(o[1744]), .IN1(n1877), .SEL(n2885), .F(\Data_Mem/n6017 ) );
  NAND U5535 ( .A(n2886), .B(n2887), .Z(n2885) );
  OR U5536 ( .A(n1880), .B(n2883), .Z(n2887) );
  ANDN U5537 ( .A(n2881), .B(n2880), .Z(n2886) );
  NANDN U5538 ( .B(n2883), .A(n1915), .Z(n2881) );
  MUX U5539 ( .IN0(n1883), .IN1(o[1743]), .SEL(n2888), .F(\Data_Mem/n6016 ) );
  MUX U5540 ( .IN0(n1885), .IN1(o[1742]), .SEL(n2888), .F(\Data_Mem/n6015 ) );
  MUX U5541 ( .IN0(n1886), .IN1(o[1741]), .SEL(n2888), .F(\Data_Mem/n6014 ) );
  MUX U5542 ( .IN0(n1887), .IN1(o[1740]), .SEL(n2888), .F(\Data_Mem/n6013 ) );
  MUX U5543 ( .IN0(n1888), .IN1(o[1739]), .SEL(n2888), .F(\Data_Mem/n6012 ) );
  IV U5544 ( .A(n2889), .Z(n2888) );
  MUX U5545 ( .IN0(o[1738]), .IN1(n1890), .SEL(n2889), .F(\Data_Mem/n6011 ) );
  MUX U5546 ( .IN0(o[1737]), .IN1(n1891), .SEL(n2889), .F(\Data_Mem/n6010 ) );
  MUX U5547 ( .IN0(o[1736]), .IN1(n1892), .SEL(n2889), .F(\Data_Mem/n6009 ) );
  NAND U5548 ( .A(n2890), .B(n2891), .Z(n2889) );
  OR U5549 ( .A(n1895), .B(n2883), .Z(n2891) );
  MUX U5550 ( .IN0(reg_target[7]), .IN1(o[1735]), .SEL(n2892), .F(
        \Data_Mem/n6008 ) );
  MUX U5551 ( .IN0(reg_target[6]), .IN1(o[1734]), .SEL(n2892), .F(
        \Data_Mem/n6007 ) );
  MUX U5552 ( .IN0(reg_target[5]), .IN1(o[1733]), .SEL(n2892), .F(
        \Data_Mem/n6006 ) );
  MUX U5553 ( .IN0(reg_target[4]), .IN1(o[1732]), .SEL(n2892), .F(
        \Data_Mem/n6005 ) );
  MUX U5554 ( .IN0(reg_target[3]), .IN1(o[1731]), .SEL(n2892), .F(
        \Data_Mem/n6004 ) );
  IV U5555 ( .A(n2893), .Z(n2892) );
  MUX U5556 ( .IN0(o[1730]), .IN1(reg_target[2]), .SEL(n2893), .F(
        \Data_Mem/n6003 ) );
  MUX U5557 ( .IN0(o[1729]), .IN1(reg_target[1]), .SEL(n2893), .F(
        \Data_Mem/n6002 ) );
  MUX U5558 ( .IN0(o[1728]), .IN1(reg_target[0]), .SEL(n2893), .F(
        \Data_Mem/n6001 ) );
  NAND U5559 ( .A(n2890), .B(n2894), .Z(n2893) );
  NANDN U5560 ( .B(n2883), .A(n1899), .Z(n2894) );
  ANDN U5561 ( .A(n2895), .B(n2880), .Z(n2890) );
  ANDN U5562 ( .A(n1902), .B(n2883), .Z(n2880) );
  NANDN U5563 ( .B(n2883), .A(n1924), .Z(n2895) );
  NAND U5564 ( .A(n2020), .B(n2787), .Z(n2883) );
  MUX U5565 ( .IN0(n1853), .IN1(o[1791]), .SEL(n2896), .F(\Data_Mem/n6000 ) );
  MUX U5566 ( .IN0(n1855), .IN1(o[1790]), .SEL(n2896), .F(\Data_Mem/n5999 ) );
  MUX U5567 ( .IN0(n1856), .IN1(o[1789]), .SEL(n2896), .F(\Data_Mem/n5998 ) );
  MUX U5568 ( .IN0(n1857), .IN1(o[1788]), .SEL(n2896), .F(\Data_Mem/n5997 ) );
  MUX U5569 ( .IN0(n1858), .IN1(o[1787]), .SEL(n2896), .F(\Data_Mem/n5996 ) );
  MUX U5570 ( .IN0(n1859), .IN1(o[1786]), .SEL(n2896), .F(\Data_Mem/n5995 ) );
  MUX U5571 ( .IN0(n1860), .IN1(o[1785]), .SEL(n2896), .F(\Data_Mem/n5994 ) );
  MUX U5572 ( .IN0(n1861), .IN1(o[1784]), .SEL(n2896), .F(\Data_Mem/n5993 ) );
  ANDN U5573 ( .A(n2897), .B(n2898), .Z(n2896) );
  AND U5574 ( .A(n2899), .B(n2900), .Z(n2897) );
  OR U5575 ( .A(n1867), .B(n2901), .Z(n2900) );
  MUX U5576 ( .IN0(n1868), .IN1(o[1783]), .SEL(n2902), .F(\Data_Mem/n5992 ) );
  MUX U5577 ( .IN0(n1870), .IN1(o[1782]), .SEL(n2902), .F(\Data_Mem/n5991 ) );
  MUX U5578 ( .IN0(n1871), .IN1(o[1781]), .SEL(n2902), .F(\Data_Mem/n5990 ) );
  MUX U5579 ( .IN0(n1872), .IN1(o[1780]), .SEL(n2902), .F(\Data_Mem/n5989 ) );
  MUX U5580 ( .IN0(n1873), .IN1(o[1779]), .SEL(n2902), .F(\Data_Mem/n5988 ) );
  IV U5581 ( .A(n2903), .Z(n2902) );
  MUX U5582 ( .IN0(o[1778]), .IN1(n1875), .SEL(n2903), .F(\Data_Mem/n5987 ) );
  MUX U5583 ( .IN0(o[1777]), .IN1(n1876), .SEL(n2903), .F(\Data_Mem/n5986 ) );
  MUX U5584 ( .IN0(o[1776]), .IN1(n1877), .SEL(n2903), .F(\Data_Mem/n5985 ) );
  NAND U5585 ( .A(n2904), .B(n2905), .Z(n2903) );
  OR U5586 ( .A(n1880), .B(n2901), .Z(n2905) );
  ANDN U5587 ( .A(n2899), .B(n2898), .Z(n2904) );
  NANDN U5588 ( .B(n2901), .A(n1915), .Z(n2899) );
  MUX U5589 ( .IN0(n1883), .IN1(o[1775]), .SEL(n2906), .F(\Data_Mem/n5984 ) );
  MUX U5590 ( .IN0(n1885), .IN1(o[1774]), .SEL(n2906), .F(\Data_Mem/n5983 ) );
  MUX U5591 ( .IN0(n1886), .IN1(o[1773]), .SEL(n2906), .F(\Data_Mem/n5982 ) );
  MUX U5592 ( .IN0(n1887), .IN1(o[1772]), .SEL(n2906), .F(\Data_Mem/n5981 ) );
  MUX U5593 ( .IN0(n1888), .IN1(o[1771]), .SEL(n2906), .F(\Data_Mem/n5980 ) );
  IV U5594 ( .A(n2907), .Z(n2906) );
  MUX U5595 ( .IN0(o[1770]), .IN1(n1890), .SEL(n2907), .F(\Data_Mem/n5979 ) );
  MUX U5596 ( .IN0(o[1769]), .IN1(n1891), .SEL(n2907), .F(\Data_Mem/n5978 ) );
  MUX U5597 ( .IN0(o[1768]), .IN1(n1892), .SEL(n2907), .F(\Data_Mem/n5977 ) );
  NAND U5598 ( .A(n2908), .B(n2909), .Z(n2907) );
  OR U5599 ( .A(n1895), .B(n2901), .Z(n2909) );
  MUX U5600 ( .IN0(reg_target[7]), .IN1(o[1767]), .SEL(n2910), .F(
        \Data_Mem/n5976 ) );
  MUX U5601 ( .IN0(reg_target[6]), .IN1(o[1766]), .SEL(n2910), .F(
        \Data_Mem/n5975 ) );
  MUX U5602 ( .IN0(reg_target[5]), .IN1(o[1765]), .SEL(n2910), .F(
        \Data_Mem/n5974 ) );
  MUX U5603 ( .IN0(reg_target[4]), .IN1(o[1764]), .SEL(n2910), .F(
        \Data_Mem/n5973 ) );
  MUX U5604 ( .IN0(reg_target[3]), .IN1(o[1763]), .SEL(n2910), .F(
        \Data_Mem/n5972 ) );
  IV U5605 ( .A(n2911), .Z(n2910) );
  MUX U5606 ( .IN0(o[1762]), .IN1(reg_target[2]), .SEL(n2911), .F(
        \Data_Mem/n5971 ) );
  MUX U5607 ( .IN0(o[1761]), .IN1(reg_target[1]), .SEL(n2911), .F(
        \Data_Mem/n5970 ) );
  MUX U5608 ( .IN0(o[1760]), .IN1(reg_target[0]), .SEL(n2911), .F(
        \Data_Mem/n5969 ) );
  NAND U5609 ( .A(n2908), .B(n2912), .Z(n2911) );
  NANDN U5610 ( .B(n2901), .A(n1899), .Z(n2912) );
  ANDN U5611 ( .A(n2913), .B(n2898), .Z(n2908) );
  ANDN U5612 ( .A(n1902), .B(n2901), .Z(n2898) );
  NANDN U5613 ( .B(n2901), .A(n1924), .Z(n2913) );
  NAND U5614 ( .A(n2787), .B(n2039), .Z(n2901) );
  ANDN U5615 ( .A(n2332), .B(n485), .Z(n2787) );
  AND U5616 ( .A(n532), .B(N25), .Z(n2332) );
  MUX U5617 ( .IN0(n1853), .IN1(o[1823]), .SEL(n2914), .F(\Data_Mem/n5968 ) );
  MUX U5618 ( .IN0(n1855), .IN1(o[1822]), .SEL(n2914), .F(\Data_Mem/n5967 ) );
  MUX U5619 ( .IN0(n1856), .IN1(o[1821]), .SEL(n2914), .F(\Data_Mem/n5966 ) );
  MUX U5620 ( .IN0(n1857), .IN1(o[1820]), .SEL(n2914), .F(\Data_Mem/n5965 ) );
  MUX U5621 ( .IN0(n1858), .IN1(o[1819]), .SEL(n2914), .F(\Data_Mem/n5964 ) );
  MUX U5622 ( .IN0(n1859), .IN1(o[1818]), .SEL(n2914), .F(\Data_Mem/n5963 ) );
  MUX U5623 ( .IN0(n1860), .IN1(o[1817]), .SEL(n2914), .F(\Data_Mem/n5962 ) );
  MUX U5624 ( .IN0(n1861), .IN1(o[1816]), .SEL(n2914), .F(\Data_Mem/n5961 ) );
  ANDN U5625 ( .A(n2915), .B(n2916), .Z(n2914) );
  AND U5626 ( .A(n2917), .B(n2918), .Z(n2915) );
  OR U5627 ( .A(n1867), .B(n2919), .Z(n2918) );
  MUX U5628 ( .IN0(n1868), .IN1(o[1815]), .SEL(n2920), .F(\Data_Mem/n5960 ) );
  MUX U5629 ( .IN0(n1870), .IN1(o[1814]), .SEL(n2920), .F(\Data_Mem/n5959 ) );
  MUX U5630 ( .IN0(n1871), .IN1(o[1813]), .SEL(n2920), .F(\Data_Mem/n5958 ) );
  MUX U5631 ( .IN0(n1872), .IN1(o[1812]), .SEL(n2920), .F(\Data_Mem/n5957 ) );
  MUX U5632 ( .IN0(n1873), .IN1(o[1811]), .SEL(n2920), .F(\Data_Mem/n5956 ) );
  IV U5633 ( .A(n2921), .Z(n2920) );
  MUX U5634 ( .IN0(o[1810]), .IN1(n1875), .SEL(n2921), .F(\Data_Mem/n5955 ) );
  MUX U5635 ( .IN0(o[1809]), .IN1(n1876), .SEL(n2921), .F(\Data_Mem/n5954 ) );
  MUX U5636 ( .IN0(o[1808]), .IN1(n1877), .SEL(n2921), .F(\Data_Mem/n5953 ) );
  NAND U5637 ( .A(n2922), .B(n2923), .Z(n2921) );
  OR U5638 ( .A(n1880), .B(n2919), .Z(n2923) );
  ANDN U5639 ( .A(n2917), .B(n2916), .Z(n2922) );
  NANDN U5640 ( .B(n2919), .A(n1915), .Z(n2917) );
  MUX U5641 ( .IN0(n1883), .IN1(o[1807]), .SEL(n2924), .F(\Data_Mem/n5952 ) );
  MUX U5642 ( .IN0(n1885), .IN1(o[1806]), .SEL(n2924), .F(\Data_Mem/n5951 ) );
  MUX U5643 ( .IN0(n1886), .IN1(o[1805]), .SEL(n2924), .F(\Data_Mem/n5950 ) );
  MUX U5644 ( .IN0(n1887), .IN1(o[1804]), .SEL(n2924), .F(\Data_Mem/n5949 ) );
  MUX U5645 ( .IN0(n1888), .IN1(o[1803]), .SEL(n2924), .F(\Data_Mem/n5948 ) );
  IV U5646 ( .A(n2925), .Z(n2924) );
  MUX U5647 ( .IN0(o[1802]), .IN1(n1890), .SEL(n2925), .F(\Data_Mem/n5947 ) );
  MUX U5648 ( .IN0(o[1801]), .IN1(n1891), .SEL(n2925), .F(\Data_Mem/n5946 ) );
  MUX U5649 ( .IN0(o[1800]), .IN1(n1892), .SEL(n2925), .F(\Data_Mem/n5945 ) );
  NAND U5650 ( .A(n2926), .B(n2927), .Z(n2925) );
  OR U5651 ( .A(n1895), .B(n2919), .Z(n2927) );
  MUX U5652 ( .IN0(reg_target[7]), .IN1(o[1799]), .SEL(n2928), .F(
        \Data_Mem/n5944 ) );
  MUX U5653 ( .IN0(reg_target[6]), .IN1(o[1798]), .SEL(n2928), .F(
        \Data_Mem/n5943 ) );
  MUX U5654 ( .IN0(reg_target[5]), .IN1(o[1797]), .SEL(n2928), .F(
        \Data_Mem/n5942 ) );
  MUX U5655 ( .IN0(reg_target[4]), .IN1(o[1796]), .SEL(n2928), .F(
        \Data_Mem/n5941 ) );
  MUX U5656 ( .IN0(reg_target[3]), .IN1(o[1795]), .SEL(n2928), .F(
        \Data_Mem/n5940 ) );
  IV U5657 ( .A(n2929), .Z(n2928) );
  MUX U5658 ( .IN0(o[1794]), .IN1(reg_target[2]), .SEL(n2929), .F(
        \Data_Mem/n5939 ) );
  MUX U5659 ( .IN0(o[1793]), .IN1(reg_target[1]), .SEL(n2929), .F(
        \Data_Mem/n5938 ) );
  MUX U5660 ( .IN0(o[1792]), .IN1(reg_target[0]), .SEL(n2929), .F(
        \Data_Mem/n5937 ) );
  NAND U5661 ( .A(n2926), .B(n2930), .Z(n2929) );
  NANDN U5662 ( .B(n2919), .A(n1899), .Z(n2930) );
  ANDN U5663 ( .A(n2931), .B(n2916), .Z(n2926) );
  ANDN U5664 ( .A(n1902), .B(n2919), .Z(n2916) );
  NANDN U5665 ( .B(n2919), .A(n1924), .Z(n2931) );
  NAND U5666 ( .A(n2932), .B(n1903), .Z(n2919) );
  AND U5667 ( .A(n2933), .B(n553), .Z(n1903) );
  MUX U5668 ( .IN0(n1853), .IN1(o[1855]), .SEL(n2934), .F(\Data_Mem/n5936 ) );
  MUX U5669 ( .IN0(n1855), .IN1(o[1854]), .SEL(n2934), .F(\Data_Mem/n5935 ) );
  MUX U5670 ( .IN0(n1856), .IN1(o[1853]), .SEL(n2934), .F(\Data_Mem/n5934 ) );
  MUX U5671 ( .IN0(n1857), .IN1(o[1852]), .SEL(n2934), .F(\Data_Mem/n5933 ) );
  MUX U5672 ( .IN0(n1858), .IN1(o[1851]), .SEL(n2934), .F(\Data_Mem/n5932 ) );
  MUX U5673 ( .IN0(n1859), .IN1(o[1850]), .SEL(n2934), .F(\Data_Mem/n5931 ) );
  MUX U5674 ( .IN0(n1860), .IN1(o[1849]), .SEL(n2934), .F(\Data_Mem/n5930 ) );
  MUX U5675 ( .IN0(n1861), .IN1(o[1848]), .SEL(n2934), .F(\Data_Mem/n5929 ) );
  ANDN U5676 ( .A(n2935), .B(n2936), .Z(n2934) );
  AND U5677 ( .A(n2937), .B(n2938), .Z(n2935) );
  OR U5678 ( .A(n1867), .B(n2939), .Z(n2938) );
  MUX U5679 ( .IN0(n1868), .IN1(o[1847]), .SEL(n2940), .F(\Data_Mem/n5928 ) );
  MUX U5680 ( .IN0(n1870), .IN1(o[1846]), .SEL(n2940), .F(\Data_Mem/n5927 ) );
  MUX U5681 ( .IN0(n1871), .IN1(o[1845]), .SEL(n2940), .F(\Data_Mem/n5926 ) );
  MUX U5682 ( .IN0(n1872), .IN1(o[1844]), .SEL(n2940), .F(\Data_Mem/n5925 ) );
  MUX U5683 ( .IN0(n1873), .IN1(o[1843]), .SEL(n2940), .F(\Data_Mem/n5924 ) );
  IV U5684 ( .A(n2941), .Z(n2940) );
  MUX U5685 ( .IN0(o[1842]), .IN1(n1875), .SEL(n2941), .F(\Data_Mem/n5923 ) );
  MUX U5686 ( .IN0(o[1841]), .IN1(n1876), .SEL(n2941), .F(\Data_Mem/n5922 ) );
  MUX U5687 ( .IN0(o[1840]), .IN1(n1877), .SEL(n2941), .F(\Data_Mem/n5921 ) );
  NAND U5688 ( .A(n2942), .B(n2943), .Z(n2941) );
  OR U5689 ( .A(n1880), .B(n2939), .Z(n2943) );
  ANDN U5690 ( .A(n2937), .B(n2936), .Z(n2942) );
  NANDN U5691 ( .B(n2939), .A(n1915), .Z(n2937) );
  MUX U5692 ( .IN0(n1883), .IN1(o[1839]), .SEL(n2944), .F(\Data_Mem/n5920 ) );
  MUX U5693 ( .IN0(n1885), .IN1(o[1838]), .SEL(n2944), .F(\Data_Mem/n5919 ) );
  MUX U5694 ( .IN0(n1886), .IN1(o[1837]), .SEL(n2944), .F(\Data_Mem/n5918 ) );
  MUX U5695 ( .IN0(n1887), .IN1(o[1836]), .SEL(n2944), .F(\Data_Mem/n5917 ) );
  MUX U5696 ( .IN0(n1888), .IN1(o[1835]), .SEL(n2944), .F(\Data_Mem/n5916 ) );
  IV U5697 ( .A(n2945), .Z(n2944) );
  MUX U5698 ( .IN0(o[1834]), .IN1(n1890), .SEL(n2945), .F(\Data_Mem/n5915 ) );
  MUX U5699 ( .IN0(o[1833]), .IN1(n1891), .SEL(n2945), .F(\Data_Mem/n5914 ) );
  MUX U5700 ( .IN0(o[1832]), .IN1(n1892), .SEL(n2945), .F(\Data_Mem/n5913 ) );
  NAND U5701 ( .A(n2946), .B(n2947), .Z(n2945) );
  OR U5702 ( .A(n1895), .B(n2939), .Z(n2947) );
  MUX U5703 ( .IN0(reg_target[7]), .IN1(o[1831]), .SEL(n2948), .F(
        \Data_Mem/n5912 ) );
  MUX U5704 ( .IN0(reg_target[6]), .IN1(o[1830]), .SEL(n2948), .F(
        \Data_Mem/n5911 ) );
  MUX U5705 ( .IN0(reg_target[5]), .IN1(o[1829]), .SEL(n2948), .F(
        \Data_Mem/n5910 ) );
  MUX U5706 ( .IN0(reg_target[4]), .IN1(o[1828]), .SEL(n2948), .F(
        \Data_Mem/n5909 ) );
  MUX U5707 ( .IN0(reg_target[3]), .IN1(o[1827]), .SEL(n2948), .F(
        \Data_Mem/n5908 ) );
  IV U5708 ( .A(n2949), .Z(n2948) );
  MUX U5709 ( .IN0(o[1826]), .IN1(reg_target[2]), .SEL(n2949), .F(
        \Data_Mem/n5907 ) );
  MUX U5710 ( .IN0(o[1825]), .IN1(reg_target[1]), .SEL(n2949), .F(
        \Data_Mem/n5906 ) );
  MUX U5711 ( .IN0(o[1824]), .IN1(reg_target[0]), .SEL(n2949), .F(
        \Data_Mem/n5905 ) );
  NAND U5712 ( .A(n2946), .B(n2950), .Z(n2949) );
  NANDN U5713 ( .B(n2939), .A(n1899), .Z(n2950) );
  ANDN U5714 ( .A(n2951), .B(n2936), .Z(n2946) );
  ANDN U5715 ( .A(n1902), .B(n2939), .Z(n2936) );
  NANDN U5716 ( .B(n2939), .A(n1924), .Z(n2951) );
  NAND U5717 ( .A(n1925), .B(n2932), .Z(n2939) );
  AND U5718 ( .A(n2952), .B(n553), .Z(n1925) );
  MUX U5719 ( .IN0(n1853), .IN1(o[1887]), .SEL(n2953), .F(\Data_Mem/n5904 ) );
  MUX U5720 ( .IN0(n1855), .IN1(o[1886]), .SEL(n2953), .F(\Data_Mem/n5903 ) );
  MUX U5721 ( .IN0(n1856), .IN1(o[1885]), .SEL(n2953), .F(\Data_Mem/n5902 ) );
  MUX U5722 ( .IN0(n1857), .IN1(o[1884]), .SEL(n2953), .F(\Data_Mem/n5901 ) );
  MUX U5723 ( .IN0(n1858), .IN1(o[1883]), .SEL(n2953), .F(\Data_Mem/n5900 ) );
  MUX U5724 ( .IN0(n1859), .IN1(o[1882]), .SEL(n2953), .F(\Data_Mem/n5899 ) );
  MUX U5725 ( .IN0(n1860), .IN1(o[1881]), .SEL(n2953), .F(\Data_Mem/n5898 ) );
  MUX U5726 ( .IN0(n1861), .IN1(o[1880]), .SEL(n2953), .F(\Data_Mem/n5897 ) );
  ANDN U5727 ( .A(n2954), .B(n2955), .Z(n2953) );
  AND U5728 ( .A(n2956), .B(n2957), .Z(n2954) );
  OR U5729 ( .A(n1867), .B(n2958), .Z(n2957) );
  MUX U5730 ( .IN0(n1868), .IN1(o[1879]), .SEL(n2959), .F(\Data_Mem/n5896 ) );
  MUX U5731 ( .IN0(n1870), .IN1(o[1878]), .SEL(n2959), .F(\Data_Mem/n5895 ) );
  MUX U5732 ( .IN0(n1871), .IN1(o[1877]), .SEL(n2959), .F(\Data_Mem/n5894 ) );
  MUX U5733 ( .IN0(n1872), .IN1(o[1876]), .SEL(n2959), .F(\Data_Mem/n5893 ) );
  MUX U5734 ( .IN0(n1873), .IN1(o[1875]), .SEL(n2959), .F(\Data_Mem/n5892 ) );
  IV U5735 ( .A(n2960), .Z(n2959) );
  MUX U5736 ( .IN0(o[1874]), .IN1(n1875), .SEL(n2960), .F(\Data_Mem/n5891 ) );
  MUX U5737 ( .IN0(o[1873]), .IN1(n1876), .SEL(n2960), .F(\Data_Mem/n5890 ) );
  MUX U5738 ( .IN0(o[1872]), .IN1(n1877), .SEL(n2960), .F(\Data_Mem/n5889 ) );
  NAND U5739 ( .A(n2961), .B(n2962), .Z(n2960) );
  OR U5740 ( .A(n1880), .B(n2958), .Z(n2962) );
  ANDN U5741 ( .A(n2956), .B(n2955), .Z(n2961) );
  NANDN U5742 ( .B(n2958), .A(n1915), .Z(n2956) );
  MUX U5743 ( .IN0(n1883), .IN1(o[1871]), .SEL(n2963), .F(\Data_Mem/n5888 ) );
  MUX U5744 ( .IN0(n1885), .IN1(o[1870]), .SEL(n2963), .F(\Data_Mem/n5887 ) );
  MUX U5745 ( .IN0(n1886), .IN1(o[1869]), .SEL(n2963), .F(\Data_Mem/n5886 ) );
  MUX U5746 ( .IN0(n1887), .IN1(o[1868]), .SEL(n2963), .F(\Data_Mem/n5885 ) );
  MUX U5747 ( .IN0(n1888), .IN1(o[1867]), .SEL(n2963), .F(\Data_Mem/n5884 ) );
  IV U5748 ( .A(n2964), .Z(n2963) );
  MUX U5749 ( .IN0(o[1866]), .IN1(n1890), .SEL(n2964), .F(\Data_Mem/n5883 ) );
  MUX U5750 ( .IN0(o[1865]), .IN1(n1891), .SEL(n2964), .F(\Data_Mem/n5882 ) );
  MUX U5751 ( .IN0(o[1864]), .IN1(n1892), .SEL(n2964), .F(\Data_Mem/n5881 ) );
  NAND U5752 ( .A(n2965), .B(n2966), .Z(n2964) );
  OR U5753 ( .A(n1895), .B(n2958), .Z(n2966) );
  MUX U5754 ( .IN0(reg_target[7]), .IN1(o[1863]), .SEL(n2967), .F(
        \Data_Mem/n5880 ) );
  MUX U5755 ( .IN0(reg_target[6]), .IN1(o[1862]), .SEL(n2967), .F(
        \Data_Mem/n5879 ) );
  MUX U5756 ( .IN0(reg_target[5]), .IN1(o[1861]), .SEL(n2967), .F(
        \Data_Mem/n5878 ) );
  MUX U5757 ( .IN0(reg_target[4]), .IN1(o[1860]), .SEL(n2967), .F(
        \Data_Mem/n5877 ) );
  MUX U5758 ( .IN0(reg_target[3]), .IN1(o[1859]), .SEL(n2967), .F(
        \Data_Mem/n5876 ) );
  IV U5759 ( .A(n2968), .Z(n2967) );
  MUX U5760 ( .IN0(o[1858]), .IN1(reg_target[2]), .SEL(n2968), .F(
        \Data_Mem/n5875 ) );
  MUX U5761 ( .IN0(o[1857]), .IN1(reg_target[1]), .SEL(n2968), .F(
        \Data_Mem/n5874 ) );
  MUX U5762 ( .IN0(o[1856]), .IN1(reg_target[0]), .SEL(n2968), .F(
        \Data_Mem/n5873 ) );
  NAND U5763 ( .A(n2965), .B(n2969), .Z(n2968) );
  NANDN U5764 ( .B(n2958), .A(n1899), .Z(n2969) );
  ANDN U5765 ( .A(n2970), .B(n2955), .Z(n2965) );
  ANDN U5766 ( .A(n1902), .B(n2958), .Z(n2955) );
  NANDN U5767 ( .B(n2958), .A(n1924), .Z(n2970) );
  NAND U5768 ( .A(n1944), .B(n2932), .Z(n2958) );
  AND U5769 ( .A(n2971), .B(n553), .Z(n1944) );
  MUX U5770 ( .IN0(n1853), .IN1(o[1919]), .SEL(n2972), .F(\Data_Mem/n5872 ) );
  MUX U5771 ( .IN0(n1855), .IN1(o[1918]), .SEL(n2972), .F(\Data_Mem/n5871 ) );
  MUX U5772 ( .IN0(n1856), .IN1(o[1917]), .SEL(n2972), .F(\Data_Mem/n5870 ) );
  MUX U5773 ( .IN0(n1857), .IN1(o[1916]), .SEL(n2972), .F(\Data_Mem/n5869 ) );
  MUX U5774 ( .IN0(n1858), .IN1(o[1915]), .SEL(n2972), .F(\Data_Mem/n5868 ) );
  MUX U5775 ( .IN0(n1859), .IN1(o[1914]), .SEL(n2972), .F(\Data_Mem/n5867 ) );
  MUX U5776 ( .IN0(n1860), .IN1(o[1913]), .SEL(n2972), .F(\Data_Mem/n5866 ) );
  MUX U5777 ( .IN0(n1861), .IN1(o[1912]), .SEL(n2972), .F(\Data_Mem/n5865 ) );
  ANDN U5778 ( .A(n2973), .B(n2974), .Z(n2972) );
  AND U5779 ( .A(n2975), .B(n2976), .Z(n2973) );
  OR U5780 ( .A(n1867), .B(n2977), .Z(n2976) );
  MUX U5781 ( .IN0(n1868), .IN1(o[1911]), .SEL(n2978), .F(\Data_Mem/n5864 ) );
  MUX U5782 ( .IN0(n1870), .IN1(o[1910]), .SEL(n2978), .F(\Data_Mem/n5863 ) );
  MUX U5783 ( .IN0(n1871), .IN1(o[1909]), .SEL(n2978), .F(\Data_Mem/n5862 ) );
  MUX U5784 ( .IN0(n1872), .IN1(o[1908]), .SEL(n2978), .F(\Data_Mem/n5861 ) );
  MUX U5785 ( .IN0(n1873), .IN1(o[1907]), .SEL(n2978), .F(\Data_Mem/n5860 ) );
  IV U5786 ( .A(n2979), .Z(n2978) );
  MUX U5787 ( .IN0(o[1906]), .IN1(n1875), .SEL(n2979), .F(\Data_Mem/n5859 ) );
  MUX U5788 ( .IN0(o[1905]), .IN1(n1876), .SEL(n2979), .F(\Data_Mem/n5858 ) );
  MUX U5789 ( .IN0(o[1904]), .IN1(n1877), .SEL(n2979), .F(\Data_Mem/n5857 ) );
  NAND U5790 ( .A(n2980), .B(n2981), .Z(n2979) );
  OR U5791 ( .A(n1880), .B(n2977), .Z(n2981) );
  ANDN U5792 ( .A(n2975), .B(n2974), .Z(n2980) );
  NANDN U5793 ( .B(n2977), .A(n1915), .Z(n2975) );
  MUX U5794 ( .IN0(n1883), .IN1(o[1903]), .SEL(n2982), .F(\Data_Mem/n5856 ) );
  MUX U5795 ( .IN0(n1885), .IN1(o[1902]), .SEL(n2982), .F(\Data_Mem/n5855 ) );
  MUX U5796 ( .IN0(n1886), .IN1(o[1901]), .SEL(n2982), .F(\Data_Mem/n5854 ) );
  MUX U5797 ( .IN0(n1887), .IN1(o[1900]), .SEL(n2982), .F(\Data_Mem/n5853 ) );
  MUX U5798 ( .IN0(n1888), .IN1(o[1899]), .SEL(n2982), .F(\Data_Mem/n5852 ) );
  IV U5799 ( .A(n2983), .Z(n2982) );
  MUX U5800 ( .IN0(o[1898]), .IN1(n1890), .SEL(n2983), .F(\Data_Mem/n5851 ) );
  MUX U5801 ( .IN0(o[1897]), .IN1(n1891), .SEL(n2983), .F(\Data_Mem/n5850 ) );
  MUX U5802 ( .IN0(o[1896]), .IN1(n1892), .SEL(n2983), .F(\Data_Mem/n5849 ) );
  NAND U5803 ( .A(n2984), .B(n2985), .Z(n2983) );
  OR U5804 ( .A(n1895), .B(n2977), .Z(n2985) );
  MUX U5805 ( .IN0(reg_target[7]), .IN1(o[1895]), .SEL(n2986), .F(
        \Data_Mem/n5848 ) );
  MUX U5806 ( .IN0(reg_target[6]), .IN1(o[1894]), .SEL(n2986), .F(
        \Data_Mem/n5847 ) );
  MUX U5807 ( .IN0(reg_target[5]), .IN1(o[1893]), .SEL(n2986), .F(
        \Data_Mem/n5846 ) );
  MUX U5808 ( .IN0(reg_target[4]), .IN1(o[1892]), .SEL(n2986), .F(
        \Data_Mem/n5845 ) );
  MUX U5809 ( .IN0(reg_target[3]), .IN1(o[1891]), .SEL(n2986), .F(
        \Data_Mem/n5844 ) );
  IV U5810 ( .A(n2987), .Z(n2986) );
  MUX U5811 ( .IN0(o[1890]), .IN1(reg_target[2]), .SEL(n2987), .F(
        \Data_Mem/n5843 ) );
  MUX U5812 ( .IN0(o[1889]), .IN1(reg_target[1]), .SEL(n2987), .F(
        \Data_Mem/n5842 ) );
  MUX U5813 ( .IN0(o[1888]), .IN1(reg_target[0]), .SEL(n2987), .F(
        \Data_Mem/n5841 ) );
  NAND U5814 ( .A(n2984), .B(n2988), .Z(n2987) );
  NANDN U5815 ( .B(n2977), .A(n1899), .Z(n2988) );
  ANDN U5816 ( .A(n2989), .B(n2974), .Z(n2984) );
  ANDN U5817 ( .A(n1902), .B(n2977), .Z(n2974) );
  NANDN U5818 ( .B(n2977), .A(n1924), .Z(n2989) );
  NAND U5819 ( .A(n1963), .B(n2932), .Z(n2977) );
  AND U5820 ( .A(n2990), .B(n553), .Z(n1963) );
  MUX U5821 ( .IN0(n1853), .IN1(o[1951]), .SEL(n2991), .F(\Data_Mem/n5840 ) );
  MUX U5822 ( .IN0(n1855), .IN1(o[1950]), .SEL(n2991), .F(\Data_Mem/n5839 ) );
  MUX U5823 ( .IN0(n1856), .IN1(o[1949]), .SEL(n2991), .F(\Data_Mem/n5838 ) );
  MUX U5824 ( .IN0(n1857), .IN1(o[1948]), .SEL(n2991), .F(\Data_Mem/n5837 ) );
  MUX U5825 ( .IN0(n1858), .IN1(o[1947]), .SEL(n2991), .F(\Data_Mem/n5836 ) );
  MUX U5826 ( .IN0(n1859), .IN1(o[1946]), .SEL(n2991), .F(\Data_Mem/n5835 ) );
  MUX U5827 ( .IN0(n1860), .IN1(o[1945]), .SEL(n2991), .F(\Data_Mem/n5834 ) );
  MUX U5828 ( .IN0(n1861), .IN1(o[1944]), .SEL(n2991), .F(\Data_Mem/n5833 ) );
  ANDN U5829 ( .A(n2992), .B(n2993), .Z(n2991) );
  AND U5830 ( .A(n2994), .B(n2995), .Z(n2992) );
  OR U5831 ( .A(n1867), .B(n2996), .Z(n2995) );
  MUX U5832 ( .IN0(n1868), .IN1(o[1943]), .SEL(n2997), .F(\Data_Mem/n5832 ) );
  MUX U5833 ( .IN0(n1870), .IN1(o[1942]), .SEL(n2997), .F(\Data_Mem/n5831 ) );
  MUX U5834 ( .IN0(n1871), .IN1(o[1941]), .SEL(n2997), .F(\Data_Mem/n5830 ) );
  MUX U5835 ( .IN0(n1872), .IN1(o[1940]), .SEL(n2997), .F(\Data_Mem/n5829 ) );
  MUX U5836 ( .IN0(n1873), .IN1(o[1939]), .SEL(n2997), .F(\Data_Mem/n5828 ) );
  IV U5837 ( .A(n2998), .Z(n2997) );
  MUX U5838 ( .IN0(o[1938]), .IN1(n1875), .SEL(n2998), .F(\Data_Mem/n5827 ) );
  MUX U5839 ( .IN0(o[1937]), .IN1(n1876), .SEL(n2998), .F(\Data_Mem/n5826 ) );
  MUX U5840 ( .IN0(o[1936]), .IN1(n1877), .SEL(n2998), .F(\Data_Mem/n5825 ) );
  NAND U5841 ( .A(n2999), .B(n3000), .Z(n2998) );
  OR U5842 ( .A(n1880), .B(n2996), .Z(n3000) );
  ANDN U5843 ( .A(n2994), .B(n2993), .Z(n2999) );
  NANDN U5844 ( .B(n2996), .A(n1915), .Z(n2994) );
  MUX U5845 ( .IN0(n1883), .IN1(o[1935]), .SEL(n3001), .F(\Data_Mem/n5824 ) );
  MUX U5846 ( .IN0(n1885), .IN1(o[1934]), .SEL(n3001), .F(\Data_Mem/n5823 ) );
  MUX U5847 ( .IN0(n1886), .IN1(o[1933]), .SEL(n3001), .F(\Data_Mem/n5822 ) );
  MUX U5848 ( .IN0(n1887), .IN1(o[1932]), .SEL(n3001), .F(\Data_Mem/n5821 ) );
  MUX U5849 ( .IN0(n1888), .IN1(o[1931]), .SEL(n3001), .F(\Data_Mem/n5820 ) );
  IV U5850 ( .A(n3002), .Z(n3001) );
  MUX U5851 ( .IN0(o[1930]), .IN1(n1890), .SEL(n3002), .F(\Data_Mem/n5819 ) );
  MUX U5852 ( .IN0(o[1929]), .IN1(n1891), .SEL(n3002), .F(\Data_Mem/n5818 ) );
  MUX U5853 ( .IN0(o[1928]), .IN1(n1892), .SEL(n3002), .F(\Data_Mem/n5817 ) );
  NAND U5854 ( .A(n3003), .B(n3004), .Z(n3002) );
  OR U5855 ( .A(n1895), .B(n2996), .Z(n3004) );
  MUX U5856 ( .IN0(reg_target[7]), .IN1(o[1927]), .SEL(n3005), .F(
        \Data_Mem/n5816 ) );
  MUX U5857 ( .IN0(reg_target[6]), .IN1(o[1926]), .SEL(n3005), .F(
        \Data_Mem/n5815 ) );
  MUX U5858 ( .IN0(reg_target[5]), .IN1(o[1925]), .SEL(n3005), .F(
        \Data_Mem/n5814 ) );
  MUX U5859 ( .IN0(reg_target[4]), .IN1(o[1924]), .SEL(n3005), .F(
        \Data_Mem/n5813 ) );
  MUX U5860 ( .IN0(reg_target[3]), .IN1(o[1923]), .SEL(n3005), .F(
        \Data_Mem/n5812 ) );
  IV U5861 ( .A(n3006), .Z(n3005) );
  MUX U5862 ( .IN0(o[1922]), .IN1(reg_target[2]), .SEL(n3006), .F(
        \Data_Mem/n5811 ) );
  MUX U5863 ( .IN0(o[1921]), .IN1(reg_target[1]), .SEL(n3006), .F(
        \Data_Mem/n5810 ) );
  MUX U5864 ( .IN0(o[1920]), .IN1(reg_target[0]), .SEL(n3006), .F(
        \Data_Mem/n5809 ) );
  NAND U5865 ( .A(n3003), .B(n3007), .Z(n3006) );
  NANDN U5866 ( .B(n2996), .A(n1899), .Z(n3007) );
  ANDN U5867 ( .A(n3008), .B(n2993), .Z(n3003) );
  ANDN U5868 ( .A(n1902), .B(n2996), .Z(n2993) );
  NANDN U5869 ( .B(n2996), .A(n1924), .Z(n3008) );
  NAND U5870 ( .A(n1982), .B(n2932), .Z(n2996) );
  ANDN U5871 ( .A(n2933), .B(n553), .Z(n1982) );
  AND U5872 ( .A(n595), .B(n574), .Z(n2933) );
  MUX U5873 ( .IN0(n1853), .IN1(o[1983]), .SEL(n3009), .F(\Data_Mem/n5808 ) );
  MUX U5874 ( .IN0(n1855), .IN1(o[1982]), .SEL(n3009), .F(\Data_Mem/n5807 ) );
  MUX U5875 ( .IN0(n1856), .IN1(o[1981]), .SEL(n3009), .F(\Data_Mem/n5806 ) );
  MUX U5876 ( .IN0(n1857), .IN1(o[1980]), .SEL(n3009), .F(\Data_Mem/n5805 ) );
  MUX U5877 ( .IN0(n1858), .IN1(o[1979]), .SEL(n3009), .F(\Data_Mem/n5804 ) );
  MUX U5878 ( .IN0(n1859), .IN1(o[1978]), .SEL(n3009), .F(\Data_Mem/n5803 ) );
  MUX U5879 ( .IN0(n1860), .IN1(o[1977]), .SEL(n3009), .F(\Data_Mem/n5802 ) );
  MUX U5880 ( .IN0(n1861), .IN1(o[1976]), .SEL(n3009), .F(\Data_Mem/n5801 ) );
  ANDN U5881 ( .A(n3010), .B(n3011), .Z(n3009) );
  AND U5882 ( .A(n3012), .B(n3013), .Z(n3010) );
  OR U5883 ( .A(n1867), .B(n3014), .Z(n3013) );
  MUX U5884 ( .IN0(n1868), .IN1(o[1975]), .SEL(n3015), .F(\Data_Mem/n5800 ) );
  MUX U5885 ( .IN0(n1870), .IN1(o[1974]), .SEL(n3015), .F(\Data_Mem/n5799 ) );
  MUX U5886 ( .IN0(n1871), .IN1(o[1973]), .SEL(n3015), .F(\Data_Mem/n5798 ) );
  MUX U5887 ( .IN0(n1872), .IN1(o[1972]), .SEL(n3015), .F(\Data_Mem/n5797 ) );
  MUX U5888 ( .IN0(n1873), .IN1(o[1971]), .SEL(n3015), .F(\Data_Mem/n5796 ) );
  IV U5889 ( .A(n3016), .Z(n3015) );
  MUX U5890 ( .IN0(o[1970]), .IN1(n1875), .SEL(n3016), .F(\Data_Mem/n5795 ) );
  MUX U5891 ( .IN0(o[1969]), .IN1(n1876), .SEL(n3016), .F(\Data_Mem/n5794 ) );
  MUX U5892 ( .IN0(o[1968]), .IN1(n1877), .SEL(n3016), .F(\Data_Mem/n5793 ) );
  NAND U5893 ( .A(n3017), .B(n3018), .Z(n3016) );
  OR U5894 ( .A(n1880), .B(n3014), .Z(n3018) );
  ANDN U5895 ( .A(n3012), .B(n3011), .Z(n3017) );
  NANDN U5896 ( .B(n3014), .A(n1915), .Z(n3012) );
  MUX U5897 ( .IN0(n1883), .IN1(o[1967]), .SEL(n3019), .F(\Data_Mem/n5792 ) );
  MUX U5898 ( .IN0(n1885), .IN1(o[1966]), .SEL(n3019), .F(\Data_Mem/n5791 ) );
  MUX U5899 ( .IN0(n1886), .IN1(o[1965]), .SEL(n3019), .F(\Data_Mem/n5790 ) );
  MUX U5900 ( .IN0(n1887), .IN1(o[1964]), .SEL(n3019), .F(\Data_Mem/n5789 ) );
  MUX U5901 ( .IN0(n1888), .IN1(o[1963]), .SEL(n3019), .F(\Data_Mem/n5788 ) );
  IV U5902 ( .A(n3020), .Z(n3019) );
  MUX U5903 ( .IN0(o[1962]), .IN1(n1890), .SEL(n3020), .F(\Data_Mem/n5787 ) );
  MUX U5904 ( .IN0(o[1961]), .IN1(n1891), .SEL(n3020), .F(\Data_Mem/n5786 ) );
  MUX U5905 ( .IN0(o[1960]), .IN1(n1892), .SEL(n3020), .F(\Data_Mem/n5785 ) );
  NAND U5906 ( .A(n3021), .B(n3022), .Z(n3020) );
  OR U5907 ( .A(n3014), .B(n1895), .Z(n3022) );
  MUX U5908 ( .IN0(reg_target[7]), .IN1(o[1959]), .SEL(n3023), .F(
        \Data_Mem/n5784 ) );
  MUX U5909 ( .IN0(reg_target[6]), .IN1(o[1958]), .SEL(n3023), .F(
        \Data_Mem/n5783 ) );
  MUX U5910 ( .IN0(reg_target[5]), .IN1(o[1957]), .SEL(n3023), .F(
        \Data_Mem/n5782 ) );
  MUX U5911 ( .IN0(reg_target[4]), .IN1(o[1956]), .SEL(n3023), .F(
        \Data_Mem/n5781 ) );
  MUX U5912 ( .IN0(reg_target[3]), .IN1(o[1955]), .SEL(n3023), .F(
        \Data_Mem/n5780 ) );
  IV U5913 ( .A(n3024), .Z(n3023) );
  MUX U5914 ( .IN0(o[1954]), .IN1(reg_target[2]), .SEL(n3024), .F(
        \Data_Mem/n5779 ) );
  MUX U5915 ( .IN0(o[1953]), .IN1(reg_target[1]), .SEL(n3024), .F(
        \Data_Mem/n5778 ) );
  MUX U5916 ( .IN0(o[1952]), .IN1(reg_target[0]), .SEL(n3024), .F(
        \Data_Mem/n5777 ) );
  NAND U5917 ( .A(n3021), .B(n3025), .Z(n3024) );
  NANDN U5918 ( .B(n3014), .A(n1899), .Z(n3025) );
  ANDN U5919 ( .A(n3026), .B(n3011), .Z(n3021) );
  ANDN U5920 ( .A(n1902), .B(n3014), .Z(n3011) );
  NANDN U5921 ( .B(n3014), .A(n1924), .Z(n3026) );
  NAND U5922 ( .A(n2001), .B(n2932), .Z(n3014) );
  ANDN U5923 ( .A(n2952), .B(n553), .Z(n2001) );
  AND U5924 ( .A(n574), .B(N29), .Z(n2952) );
  MUX U5925 ( .IN0(n1853), .IN1(o[2015]), .SEL(n3027), .F(\Data_Mem/n5776 ) );
  MUX U5926 ( .IN0(n1855), .IN1(o[2014]), .SEL(n3027), .F(\Data_Mem/n5775 ) );
  MUX U5927 ( .IN0(n1856), .IN1(o[2013]), .SEL(n3027), .F(\Data_Mem/n5774 ) );
  MUX U5928 ( .IN0(n1857), .IN1(o[2012]), .SEL(n3027), .F(\Data_Mem/n5773 ) );
  MUX U5929 ( .IN0(n1858), .IN1(o[2011]), .SEL(n3027), .F(\Data_Mem/n5772 ) );
  MUX U5930 ( .IN0(n1859), .IN1(o[2010]), .SEL(n3027), .F(\Data_Mem/n5771 ) );
  MUX U5931 ( .IN0(n1860), .IN1(o[2009]), .SEL(n3027), .F(\Data_Mem/n5770 ) );
  MUX U5932 ( .IN0(n1861), .IN1(o[2008]), .SEL(n3027), .F(\Data_Mem/n5769 ) );
  ANDN U5933 ( .A(n3028), .B(n3029), .Z(n3027) );
  ANDN U5934 ( .A(n3030), .B(n3031), .Z(n3028) );
  NANDN U5935 ( .B(n1867), .A(n3032), .Z(n3030) );
  NAND U5936 ( .A(n3033), .B(n504), .Z(n1867) );
  MUX U5937 ( .IN0(n1868), .IN1(o[2007]), .SEL(n3034), .F(\Data_Mem/n5768 ) );
  MUX U5938 ( .IN0(n1870), .IN1(o[2006]), .SEL(n3034), .F(\Data_Mem/n5767 ) );
  MUX U5939 ( .IN0(n1871), .IN1(o[2005]), .SEL(n3034), .F(\Data_Mem/n5766 ) );
  MUX U5940 ( .IN0(n1872), .IN1(o[2004]), .SEL(n3034), .F(\Data_Mem/n5765 ) );
  MUX U5941 ( .IN0(n1873), .IN1(o[2003]), .SEL(n3034), .F(\Data_Mem/n5764 ) );
  IV U5942 ( .A(n3035), .Z(n3034) );
  MUX U5943 ( .IN0(o[2002]), .IN1(n1875), .SEL(n3035), .F(\Data_Mem/n5763 ) );
  MUX U5944 ( .IN0(o[2001]), .IN1(n1876), .SEL(n3035), .F(\Data_Mem/n5762 ) );
  MUX U5945 ( .IN0(o[2000]), .IN1(n1877), .SEL(n3035), .F(\Data_Mem/n5761 ) );
  NAND U5946 ( .A(n3036), .B(n3037), .Z(n3035) );
  NANDN U5947 ( .B(n1880), .A(n3032), .Z(n3037) );
  NAND U5948 ( .A(n3033), .B(n503), .Z(n1880) );
  NOR U5949 ( .A(n3029), .B(n3031), .Z(n3036) );
  AND U5950 ( .A(n1915), .B(n3032), .Z(n3031) );
  MUX U5951 ( .IN0(n1883), .IN1(o[1999]), .SEL(n3038), .F(\Data_Mem/n5760 ) );
  MUX U5952 ( .IN0(n1885), .IN1(o[1998]), .SEL(n3038), .F(\Data_Mem/n5759 ) );
  MUX U5953 ( .IN0(n1886), .IN1(o[1997]), .SEL(n3038), .F(\Data_Mem/n5758 ) );
  MUX U5954 ( .IN0(n1887), .IN1(o[1996]), .SEL(n3038), .F(\Data_Mem/n5757 ) );
  MUX U5955 ( .IN0(n1888), .IN1(o[1995]), .SEL(n3038), .F(\Data_Mem/n5756 ) );
  IV U5956 ( .A(n3039), .Z(n3038) );
  MUX U5957 ( .IN0(o[1994]), .IN1(n1890), .SEL(n3039), .F(\Data_Mem/n5755 ) );
  MUX U5958 ( .IN0(o[1993]), .IN1(n1891), .SEL(n3039), .F(\Data_Mem/n5754 ) );
  MUX U5959 ( .IN0(o[1992]), .IN1(n1892), .SEL(n3039), .F(\Data_Mem/n5753 ) );
  NAND U5960 ( .A(n3040), .B(n3041), .Z(n3039) );
  NANDN U5961 ( .B(n1895), .A(n3032), .Z(n3041) );
  NAND U5962 ( .A(n3033), .B(n500), .Z(n1895) );
  MUX U5963 ( .IN0(reg_target[7]), .IN1(o[1991]), .SEL(n3042), .F(
        \Data_Mem/n5752 ) );
  MUX U5964 ( .IN0(reg_target[6]), .IN1(o[1990]), .SEL(n3042), .F(
        \Data_Mem/n5751 ) );
  MUX U5965 ( .IN0(reg_target[5]), .IN1(o[1989]), .SEL(n3042), .F(
        \Data_Mem/n5750 ) );
  MUX U5966 ( .IN0(reg_target[4]), .IN1(o[1988]), .SEL(n3042), .F(
        \Data_Mem/n5749 ) );
  MUX U5967 ( .IN0(reg_target[3]), .IN1(o[1987]), .SEL(n3042), .F(
        \Data_Mem/n5748 ) );
  IV U5968 ( .A(n3043), .Z(n3042) );
  MUX U5969 ( .IN0(o[1986]), .IN1(reg_target[2]), .SEL(n3043), .F(
        \Data_Mem/n5747 ) );
  MUX U5970 ( .IN0(o[1985]), .IN1(reg_target[1]), .SEL(n3043), .F(
        \Data_Mem/n5746 ) );
  MUX U5971 ( .IN0(o[1984]), .IN1(reg_target[0]), .SEL(n3043), .F(
        \Data_Mem/n5745 ) );
  NAND U5972 ( .A(n3040), .B(n3044), .Z(n3043) );
  NAND U5973 ( .A(n1899), .B(n3032), .Z(n3044) );
  NOR U5974 ( .A(n3029), .B(n3045), .Z(n3040) );
  AND U5975 ( .A(n1924), .B(n3032), .Z(n3045) );
  AND U5976 ( .A(n3032), .B(n1902), .Z(n3029) );
  AND U5977 ( .A(n2020), .B(n2932), .Z(n3032) );
  ANDN U5978 ( .A(n2971), .B(n553), .Z(n2020) );
  AND U5979 ( .A(n595), .B(N28), .Z(n2971) );
  MUX U5980 ( .IN0(n1853), .IN1(o[2047]), .SEL(n3046), .F(\Data_Mem/n5744 ) );
  NAND U5981 ( .A(n3047), .B(n3048), .Z(n1853) );
  NAND U5982 ( .A(n1902), .B(reg_target[31]), .Z(n3048) );
  AND U5983 ( .A(n3049), .B(n3050), .Z(n3047) );
  NANDN U5984 ( .B(n1882), .A(reg_target[15]), .Z(n3050) );
  MUX U5985 ( .IN0(n1855), .IN1(o[2046]), .SEL(n3046), .F(\Data_Mem/n5743 ) );
  NAND U5986 ( .A(n3051), .B(n3052), .Z(n1855) );
  NAND U5987 ( .A(n1902), .B(reg_target[30]), .Z(n3052) );
  AND U5988 ( .A(n3053), .B(n3054), .Z(n3051) );
  NANDN U5989 ( .B(n1882), .A(reg_target[14]), .Z(n3054) );
  MUX U5990 ( .IN0(n1856), .IN1(o[2045]), .SEL(n3046), .F(\Data_Mem/n5742 ) );
  NAND U5991 ( .A(n3055), .B(n3056), .Z(n1856) );
  NAND U5992 ( .A(n1902), .B(reg_target[29]), .Z(n3056) );
  AND U5993 ( .A(n3057), .B(n3058), .Z(n3055) );
  NANDN U5994 ( .B(n1882), .A(reg_target[13]), .Z(n3058) );
  MUX U5995 ( .IN0(n1857), .IN1(o[2044]), .SEL(n3046), .F(\Data_Mem/n5741 ) );
  NAND U5996 ( .A(n3059), .B(n3060), .Z(n1857) );
  NAND U5997 ( .A(n1902), .B(reg_target[28]), .Z(n3060) );
  AND U5998 ( .A(n3061), .B(n3062), .Z(n3059) );
  NANDN U5999 ( .B(n1882), .A(reg_target[12]), .Z(n3062) );
  MUX U6000 ( .IN0(n1858), .IN1(o[2043]), .SEL(n3046), .F(\Data_Mem/n5740 ) );
  NAND U6001 ( .A(n3063), .B(n3064), .Z(n1858) );
  NAND U6002 ( .A(n1902), .B(reg_target[27]), .Z(n3064) );
  AND U6003 ( .A(n3065), .B(n3066), .Z(n3063) );
  NANDN U6004 ( .B(n1882), .A(reg_target[11]), .Z(n3066) );
  MUX U6005 ( .IN0(n1859), .IN1(o[2042]), .SEL(n3046), .F(\Data_Mem/n5739 ) );
  NAND U6006 ( .A(n3067), .B(n3068), .Z(n1859) );
  NAND U6007 ( .A(n1902), .B(reg_target[26]), .Z(n3068) );
  AND U6008 ( .A(n3069), .B(n3070), .Z(n3067) );
  NANDN U6009 ( .B(n1882), .A(reg_target[10]), .Z(n3070) );
  MUX U6010 ( .IN0(n1860), .IN1(o[2041]), .SEL(n3046), .F(\Data_Mem/n5738 ) );
  NAND U6011 ( .A(n3071), .B(n3072), .Z(n1860) );
  NAND U6012 ( .A(n1902), .B(reg_target[25]), .Z(n3072) );
  AND U6013 ( .A(n3073), .B(n3074), .Z(n3071) );
  NANDN U6014 ( .B(n1882), .A(reg_target[9]), .Z(n3074) );
  MUX U6015 ( .IN0(n1861), .IN1(o[2040]), .SEL(n3046), .F(\Data_Mem/n5737 ) );
  ANDN U6016 ( .A(n3075), .B(n3076), .Z(n3046) );
  ANDN U6017 ( .A(n3077), .B(n3078), .Z(n3075) );
  NAND U6018 ( .A(n3079), .B(n504), .Z(n3077) );
  AND U6019 ( .A(n779), .B(n411), .Z(n504) );
  NAND U6020 ( .A(n3080), .B(n3081), .Z(n1861) );
  NAND U6021 ( .A(n1902), .B(reg_target[24]), .Z(n3081) );
  AND U6022 ( .A(n3082), .B(n3083), .Z(n3080) );
  NANDN U6023 ( .B(n1882), .A(reg_target[8]), .Z(n3083) );
  MUX U6024 ( .IN0(n1868), .IN1(o[2039]), .SEL(n3084), .F(\Data_Mem/n5736 ) );
  NAND U6025 ( .A(n3085), .B(n3086), .Z(n1868) );
  NAND U6026 ( .A(n3087), .B(reg_target[7]), .Z(n3086) );
  NAND U6027 ( .A(n1902), .B(reg_target[23]), .Z(n3085) );
  MUX U6028 ( .IN0(n1870), .IN1(o[2038]), .SEL(n3084), .F(\Data_Mem/n5735 ) );
  NAND U6029 ( .A(n3088), .B(n3089), .Z(n1870) );
  NAND U6030 ( .A(n3087), .B(reg_target[6]), .Z(n3089) );
  NAND U6031 ( .A(n1902), .B(reg_target[22]), .Z(n3088) );
  MUX U6032 ( .IN0(n1871), .IN1(o[2037]), .SEL(n3084), .F(\Data_Mem/n5734 ) );
  NAND U6033 ( .A(n3090), .B(n3091), .Z(n1871) );
  NAND U6034 ( .A(n3087), .B(reg_target[5]), .Z(n3091) );
  NAND U6035 ( .A(n1902), .B(reg_target[21]), .Z(n3090) );
  MUX U6036 ( .IN0(n1872), .IN1(o[2036]), .SEL(n3084), .F(\Data_Mem/n5733 ) );
  NAND U6037 ( .A(n3092), .B(n3093), .Z(n1872) );
  NAND U6038 ( .A(n3087), .B(reg_target[4]), .Z(n3093) );
  NAND U6039 ( .A(n1902), .B(reg_target[20]), .Z(n3092) );
  MUX U6040 ( .IN0(n1873), .IN1(o[2035]), .SEL(n3084), .F(\Data_Mem/n5732 ) );
  IV U6041 ( .A(n3094), .Z(n3084) );
  NAND U6042 ( .A(n3095), .B(n3096), .Z(n1873) );
  NAND U6043 ( .A(n3087), .B(reg_target[3]), .Z(n3096) );
  NAND U6044 ( .A(n1902), .B(reg_target[19]), .Z(n3095) );
  MUX U6045 ( .IN0(o[2034]), .IN1(n1875), .SEL(n3094), .F(\Data_Mem/n5731 ) );
  NAND U6046 ( .A(n3097), .B(n3098), .Z(n1875) );
  NAND U6047 ( .A(n3087), .B(reg_target[2]), .Z(n3098) );
  NAND U6048 ( .A(n1902), .B(reg_target[18]), .Z(n3097) );
  MUX U6049 ( .IN0(o[2033]), .IN1(n1876), .SEL(n3094), .F(\Data_Mem/n5730 ) );
  NAND U6050 ( .A(n3099), .B(n3100), .Z(n1876) );
  NAND U6051 ( .A(n3087), .B(reg_target[1]), .Z(n3100) );
  NAND U6052 ( .A(n1902), .B(reg_target[17]), .Z(n3099) );
  MUX U6053 ( .IN0(o[2032]), .IN1(n1877), .SEL(n3094), .F(\Data_Mem/n5729 ) );
  NAND U6054 ( .A(n3101), .B(n3102), .Z(n3094) );
  NAND U6055 ( .A(n3079), .B(n503), .Z(n3102) );
  ANDN U6056 ( .A(n411), .B(n779), .Z(n503) );
  NOR U6057 ( .A(n3076), .B(n3078), .Z(n3101) );
  ANDN U6058 ( .A(n1915), .B(n3103), .Z(n3078) );
  ANDN U6059 ( .A(n411), .B(n1882), .Z(n1915) );
  NAND U6060 ( .A(n3104), .B(n3105), .Z(n1877) );
  NAND U6061 ( .A(reg_target[0]), .B(n3087), .Z(n3105) );
  NANDN U6062 ( .B(n3033), .A(n1882), .Z(n3087) );
  NAND U6063 ( .A(n1902), .B(reg_target[16]), .Z(n3104) );
  MUX U6064 ( .IN0(n1883), .IN1(o[2031]), .SEL(n3106), .F(\Data_Mem/n5728 ) );
  NAND U6065 ( .A(n3049), .B(n3107), .Z(n1883) );
  NAND U6066 ( .A(n3108), .B(reg_target[15]), .Z(n3107) );
  NAND U6067 ( .A(n3033), .B(reg_target[7]), .Z(n3049) );
  MUX U6068 ( .IN0(n1885), .IN1(o[2030]), .SEL(n3106), .F(\Data_Mem/n5727 ) );
  NAND U6069 ( .A(n3053), .B(n3109), .Z(n1885) );
  NAND U6070 ( .A(n3108), .B(reg_target[14]), .Z(n3109) );
  NAND U6071 ( .A(n3033), .B(reg_target[6]), .Z(n3053) );
  MUX U6072 ( .IN0(n1886), .IN1(o[2029]), .SEL(n3106), .F(\Data_Mem/n5726 ) );
  NAND U6073 ( .A(n3057), .B(n3110), .Z(n1886) );
  NAND U6074 ( .A(n3108), .B(reg_target[13]), .Z(n3110) );
  NAND U6075 ( .A(n3033), .B(reg_target[5]), .Z(n3057) );
  MUX U6076 ( .IN0(n1887), .IN1(o[2028]), .SEL(n3106), .F(\Data_Mem/n5725 ) );
  NAND U6077 ( .A(n3061), .B(n3111), .Z(n1887) );
  NAND U6078 ( .A(n3108), .B(reg_target[12]), .Z(n3111) );
  NAND U6079 ( .A(n3033), .B(reg_target[4]), .Z(n3061) );
  MUX U6080 ( .IN0(n1888), .IN1(o[2027]), .SEL(n3106), .F(\Data_Mem/n5724 ) );
  IV U6081 ( .A(n3112), .Z(n3106) );
  NAND U6082 ( .A(n3065), .B(n3113), .Z(n1888) );
  NAND U6083 ( .A(n3108), .B(reg_target[11]), .Z(n3113) );
  NAND U6084 ( .A(n3033), .B(reg_target[3]), .Z(n3065) );
  MUX U6085 ( .IN0(o[2026]), .IN1(n1890), .SEL(n3112), .F(\Data_Mem/n5723 ) );
  NAND U6086 ( .A(n3069), .B(n3114), .Z(n1890) );
  NAND U6087 ( .A(n3108), .B(reg_target[10]), .Z(n3114) );
  NAND U6088 ( .A(n3033), .B(reg_target[2]), .Z(n3069) );
  MUX U6089 ( .IN0(o[2025]), .IN1(n1891), .SEL(n3112), .F(\Data_Mem/n5722 ) );
  NAND U6090 ( .A(n3073), .B(n3115), .Z(n1891) );
  NAND U6091 ( .A(n3108), .B(reg_target[9]), .Z(n3115) );
  NAND U6092 ( .A(n3033), .B(reg_target[1]), .Z(n3073) );
  MUX U6093 ( .IN0(o[2024]), .IN1(n1892), .SEL(n3112), .F(\Data_Mem/n5721 ) );
  NAND U6094 ( .A(n3116), .B(n3117), .Z(n3112) );
  NAND U6095 ( .A(n500), .B(n3079), .Z(n3117) );
  AND U6096 ( .A(n3033), .B(n3118), .Z(n3079) );
  ANDN U6097 ( .A(n779), .B(n411), .Z(n500) );
  IV U6098 ( .A(n399), .Z(n411) );
  NAND U6099 ( .A(n3082), .B(n3119), .Z(n1892) );
  NAND U6100 ( .A(reg_target[8]), .B(n3108), .Z(n3119) );
  NANDN U6101 ( .B(n1902), .A(n1882), .Z(n3108) );
  NAND U6102 ( .A(n3033), .B(reg_target[0]), .Z(n3082) );
  MUX U6103 ( .IN0(reg_target[7]), .IN1(o[2023]), .SEL(n3120), .F(
        \Data_Mem/n5720 ) );
  MUX U6104 ( .IN0(reg_target[6]), .IN1(o[2022]), .SEL(n3120), .F(
        \Data_Mem/n5719 ) );
  MUX U6105 ( .IN0(reg_target[5]), .IN1(o[2021]), .SEL(n3120), .F(
        \Data_Mem/n5718 ) );
  MUX U6106 ( .IN0(reg_target[4]), .IN1(o[2020]), .SEL(n3120), .F(
        \Data_Mem/n5717 ) );
  MUX U6107 ( .IN0(reg_target[3]), .IN1(o[2019]), .SEL(n3120), .F(
        \Data_Mem/n5716 ) );
  IV U6108 ( .A(n3121), .Z(n3120) );
  MUX U6109 ( .IN0(o[2018]), .IN1(reg_target[2]), .SEL(n3121), .F(
        \Data_Mem/n5715 ) );
  MUX U6110 ( .IN0(o[2017]), .IN1(reg_target[1]), .SEL(n3121), .F(
        \Data_Mem/n5714 ) );
  MUX U6111 ( .IN0(o[2016]), .IN1(reg_target[0]), .SEL(n3121), .F(
        \Data_Mem/n5713 ) );
  NAND U6112 ( .A(n3116), .B(n3122), .Z(n3121) );
  NANDN U6113 ( .B(n3103), .A(n1899), .Z(n3122) );
  AND U6114 ( .A(n499), .B(n3033), .Z(n1899) );
  ANDN U6115 ( .A(n3913), .B(n770), .Z(n3033) );
  NANDN U6116 ( .B(n809), .A(n774), .Z(n770) );
  ANDN U6117 ( .A(n399), .B(n779), .Z(n499) );
  NAND U6118 ( .A(n3123), .B(n3124), .Z(n779) );
  AND U6119 ( .A(n3125), .B(n3126), .Z(n3124) );
  AND U6120 ( .A(n3127), .B(n3128), .Z(n3126) );
  NAND U6121 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][0] ), .Z(n3128) );
  AND U6122 ( .A(\Shifter/sll_27/ML_int[3][0] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][0] ) );
  AND U6123 ( .A(\Shifter/sll_27/ML_int[2][0] ), .B(n3130), .Z(
        \Shifter/sll_27/ML_int[3][0] ) );
  AND U6124 ( .A(\Shifter/sll_27/ML_int[1][0] ), .B(n3131), .Z(
        \Shifter/sll_27/ML_int[2][0] ) );
  AND U6125 ( .A(b_bus[0]), .B(n3132), .Z(\Shifter/sll_27/ML_int[1][0] ) );
  AND U6126 ( .A(n3133), .B(n3134), .Z(n3127) );
  NAND U6127 ( .A(n3135), .B(n1109), .Z(n3134) );
  NAND U6128 ( .A(n3136), .B(n3137), .Z(n3135) );
  AND U6129 ( .A(n3138), .B(n3139), .Z(n3137) );
  AND U6130 ( .A(n3140), .B(n3141), .Z(n3138) );
  OR U6131 ( .A(n1470), .B(n1117), .Z(n3141) );
  AND U6132 ( .A(n3142), .B(n3143), .Z(n1470) );
  AND U6133 ( .A(n3144), .B(n3145), .Z(n3143) );
  NAND U6134 ( .A(n1179), .B(n1650), .Z(n3145) );
  AND U6135 ( .A(n3146), .B(n3147), .Z(n3136) );
  NAND U6136 ( .A(n3148), .B(n1118), .Z(n3147) );
  NAND U6137 ( .A(n3149), .B(n1121), .Z(n3133) );
  NAND U6138 ( .A(n3150), .B(n3151), .Z(n3149) );
  AND U6139 ( .A(n3152), .B(n3139), .Z(n3151) );
  NAND U6140 ( .A(n1132), .B(n1169), .Z(n3139) );
  AND U6141 ( .A(n3140), .B(n3153), .Z(n3152) );
  OR U6142 ( .A(n1472), .B(n1117), .Z(n3153) );
  AND U6143 ( .A(n3142), .B(n3154), .Z(n1472) );
  AND U6144 ( .A(n3144), .B(n3155), .Z(n3154) );
  NAND U6145 ( .A(n1415), .B(n1179), .Z(n3155) );
  NAND U6146 ( .A(n1173), .B(n1653), .Z(n3144) );
  AND U6147 ( .A(n3156), .B(n3157), .Z(n3142) );
  NAND U6148 ( .A(n1339), .B(n3158), .Z(n3157) );
  NAND U6149 ( .A(n1338), .B(n3159), .Z(n3156) );
  NANDN U6150 ( .B(n3160), .A(n1134), .Z(n3140) );
  AND U6151 ( .A(n3146), .B(n3161), .Z(n3150) );
  NAND U6152 ( .A(n3148), .B(n1129), .Z(n3161) );
  NAND U6153 ( .A(n3162), .B(n3163), .Z(n3148) );
  AND U6154 ( .A(n3164), .B(n3165), .Z(n3163) );
  OR U6155 ( .A(n3166), .B(n3167), .Z(n3165) );
  OR U6156 ( .A(n3168), .B(n3169), .Z(n3164) );
  AND U6157 ( .A(n3170), .B(n3171), .Z(n3162) );
  OR U6158 ( .A(n3172), .B(n3173), .Z(n3171) );
  OR U6159 ( .A(n3174), .B(n3175), .Z(n3170) );
  NAND U6160 ( .A(n1124), .B(n1180), .Z(n3146) );
  AND U6161 ( .A(n3176), .B(n3177), .Z(n3125) );
  NAND U6162 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U6163 ( .A(n3180), .B(n3181), .Z(n3178) );
  ANDN U6164 ( .A(n3182), .B(n3183), .Z(n3180) );
  XNOR U6165 ( .A(n3184), .B(n1851), .Z(n3182) );
  NAND U6166 ( .A(n3185), .B(n3186), .Z(n3176) );
  FADDER U6167 ( .CIN(n3187), .IN0(n1843), .IN1(n3188), .COUT(n3186) );
  NOR U6168 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U6169 ( .A(n3191), .B(n1847), .Z(n1843) );
  IV U6170 ( .A(n1851), .Z(n1847) );
  NANDN U6171 ( .B(n3192), .A(reg_source[31]), .Z(n1851) );
  IV U6172 ( .A(n3183), .Z(n3191) );
  XOR U6173 ( .A(n3193), .B(n3184), .Z(n3183) );
  IV U6174 ( .A(n3181), .Z(n3184) );
  XOR U6175 ( .A(n3194), .B(n3195), .Z(n3181) );
  AND U6176 ( .A(n1815), .B(n3196), .Z(n3195) );
  XNOR U6177 ( .A(n3197), .B(n1816), .Z(n3196) );
  NANDN U6178 ( .B(n3192), .A(reg_source[30]), .Z(n1816) );
  XNOR U6179 ( .A(n3198), .B(n3197), .Z(n1815) );
  IV U6180 ( .A(n3194), .Z(n3197) );
  XNOR U6181 ( .A(n3199), .B(n1824), .Z(n3198) );
  XOR U6182 ( .A(n3200), .B(n3201), .Z(n3194) );
  AND U6183 ( .A(n1767), .B(n3202), .Z(n3201) );
  XNOR U6184 ( .A(n3203), .B(n1768), .Z(n3202) );
  NANDN U6185 ( .B(n3192), .A(reg_source[29]), .Z(n1768) );
  XNOR U6186 ( .A(n3204), .B(n3203), .Z(n1767) );
  IV U6187 ( .A(n3200), .Z(n3203) );
  XNOR U6188 ( .A(n3199), .B(n1775), .Z(n3204) );
  XOR U6189 ( .A(n3205), .B(n3206), .Z(n3200) );
  AND U6190 ( .A(n1790), .B(n3207), .Z(n3206) );
  XNOR U6191 ( .A(n3208), .B(n1791), .Z(n3207) );
  NANDN U6192 ( .B(n3192), .A(reg_source[28]), .Z(n1791) );
  XNOR U6193 ( .A(n3209), .B(n3208), .Z(n1790) );
  IV U6194 ( .A(n3205), .Z(n3208) );
  XNOR U6195 ( .A(n3199), .B(n1798), .Z(n3209) );
  XOR U6196 ( .A(n3210), .B(n3211), .Z(n3205) );
  AND U6197 ( .A(n1713), .B(n3212), .Z(n3211) );
  XNOR U6198 ( .A(n3213), .B(n1714), .Z(n3212) );
  NANDN U6199 ( .B(n3192), .A(reg_source[27]), .Z(n1714) );
  XNOR U6200 ( .A(n3214), .B(n3213), .Z(n1713) );
  IV U6201 ( .A(n3210), .Z(n3213) );
  XNOR U6202 ( .A(n3199), .B(n1721), .Z(n3214) );
  XOR U6203 ( .A(n3215), .B(n3216), .Z(n3210) );
  AND U6204 ( .A(n1741), .B(n3217), .Z(n3216) );
  XNOR U6205 ( .A(n3218), .B(n1742), .Z(n3217) );
  NANDN U6206 ( .B(n3192), .A(reg_source[26]), .Z(n1742) );
  XNOR U6207 ( .A(n3219), .B(n3218), .Z(n1741) );
  IV U6208 ( .A(n3215), .Z(n3218) );
  XNOR U6209 ( .A(n3199), .B(n1749), .Z(n3219) );
  XOR U6210 ( .A(n3220), .B(n3221), .Z(n3215) );
  AND U6211 ( .A(n1661), .B(n3222), .Z(n3221) );
  XNOR U6212 ( .A(n3223), .B(n1662), .Z(n3222) );
  NANDN U6213 ( .B(n3192), .A(reg_source[25]), .Z(n1662) );
  XNOR U6214 ( .A(n3224), .B(n3223), .Z(n1661) );
  IV U6215 ( .A(n3220), .Z(n3223) );
  XNOR U6216 ( .A(n3199), .B(n1669), .Z(n3224) );
  XOR U6217 ( .A(n3225), .B(n3226), .Z(n3220) );
  AND U6218 ( .A(n1687), .B(n3227), .Z(n3226) );
  XNOR U6219 ( .A(n3228), .B(n1688), .Z(n3227) );
  NANDN U6220 ( .B(n3192), .A(reg_source[24]), .Z(n1688) );
  XNOR U6221 ( .A(n3229), .B(n3228), .Z(n1687) );
  IV U6222 ( .A(n3225), .Z(n3228) );
  XNOR U6223 ( .A(n3199), .B(n1695), .Z(n3229) );
  XOR U6224 ( .A(n3230), .B(n3231), .Z(n3225) );
  AND U6225 ( .A(n1601), .B(n3232), .Z(n3231) );
  XNOR U6226 ( .A(n3233), .B(n1602), .Z(n3232) );
  NANDN U6227 ( .B(n3192), .A(reg_source[23]), .Z(n1602) );
  XNOR U6228 ( .A(n3234), .B(n3233), .Z(n1601) );
  IV U6229 ( .A(n3230), .Z(n3233) );
  XNOR U6230 ( .A(n3199), .B(n1609), .Z(n3234) );
  XOR U6231 ( .A(n3235), .B(n3236), .Z(n3230) );
  AND U6232 ( .A(n1625), .B(n3237), .Z(n3236) );
  XNOR U6233 ( .A(n3238), .B(n1626), .Z(n3237) );
  NANDN U6234 ( .B(n3192), .A(reg_source[22]), .Z(n1626) );
  XNOR U6235 ( .A(n3239), .B(n3238), .Z(n1625) );
  IV U6236 ( .A(n3235), .Z(n3238) );
  XNOR U6237 ( .A(n3199), .B(n1633), .Z(n3239) );
  XOR U6238 ( .A(n3240), .B(n3241), .Z(n3235) );
  AND U6239 ( .A(n1552), .B(n3242), .Z(n3241) );
  XNOR U6240 ( .A(n3243), .B(n1553), .Z(n3242) );
  NANDN U6241 ( .B(n3192), .A(reg_source[21]), .Z(n1553) );
  XNOR U6242 ( .A(n3244), .B(n3243), .Z(n1552) );
  IV U6243 ( .A(n3240), .Z(n3243) );
  XNOR U6244 ( .A(n3199), .B(n1560), .Z(n3244) );
  XOR U6245 ( .A(n3245), .B(n3246), .Z(n3240) );
  AND U6246 ( .A(n1576), .B(n3247), .Z(n3246) );
  XNOR U6247 ( .A(n3248), .B(n1577), .Z(n3247) );
  NANDN U6248 ( .B(n3192), .A(reg_source[20]), .Z(n1577) );
  XNOR U6249 ( .A(n3249), .B(n3248), .Z(n1576) );
  IV U6250 ( .A(n3245), .Z(n3248) );
  XNOR U6251 ( .A(n3199), .B(n1584), .Z(n3249) );
  XOR U6252 ( .A(n3250), .B(n3251), .Z(n3245) );
  AND U6253 ( .A(n1501), .B(n3252), .Z(n3251) );
  XNOR U6254 ( .A(n3253), .B(n1502), .Z(n3252) );
  NANDN U6255 ( .B(n3192), .A(reg_source[19]), .Z(n1502) );
  XNOR U6256 ( .A(n3254), .B(n3253), .Z(n1501) );
  IV U6257 ( .A(n3250), .Z(n3253) );
  XNOR U6258 ( .A(n3199), .B(n1509), .Z(n3254) );
  XOR U6259 ( .A(n3255), .B(n3256), .Z(n3250) );
  AND U6260 ( .A(n1525), .B(n3257), .Z(n3256) );
  XNOR U6261 ( .A(n3258), .B(n1526), .Z(n3257) );
  NANDN U6262 ( .B(n3192), .A(reg_source[18]), .Z(n1526) );
  XNOR U6263 ( .A(n3259), .B(n3258), .Z(n1525) );
  IV U6264 ( .A(n3255), .Z(n3258) );
  XNOR U6265 ( .A(n3199), .B(n1533), .Z(n3259) );
  XOR U6266 ( .A(n3260), .B(n3261), .Z(n3255) );
  AND U6267 ( .A(n1452), .B(n3262), .Z(n3261) );
  XNOR U6268 ( .A(n3263), .B(n1453), .Z(n3262) );
  NANDN U6269 ( .B(n3192), .A(reg_source[17]), .Z(n1453) );
  XNOR U6270 ( .A(n3264), .B(n3263), .Z(n1452) );
  IV U6271 ( .A(n3260), .Z(n3263) );
  XNOR U6272 ( .A(n3199), .B(n1460), .Z(n3264) );
  XOR U6273 ( .A(n3265), .B(n3266), .Z(n3260) );
  AND U6274 ( .A(n1476), .B(n3267), .Z(n3266) );
  XNOR U6275 ( .A(n3268), .B(n1477), .Z(n3267) );
  NANDN U6276 ( .B(n3192), .A(reg_source[16]), .Z(n1477) );
  XNOR U6277 ( .A(n3269), .B(n3268), .Z(n1476) );
  IV U6278 ( .A(n3265), .Z(n3268) );
  XNOR U6279 ( .A(n3199), .B(n1484), .Z(n3269) );
  XOR U6280 ( .A(n3270), .B(n3271), .Z(n3265) );
  AND U6281 ( .A(n1382), .B(n3272), .Z(n3271) );
  XNOR U6282 ( .A(n3273), .B(n1383), .Z(n3272) );
  NANDN U6283 ( .B(n3192), .A(reg_source[15]), .Z(n1383) );
  XNOR U6284 ( .A(n3274), .B(n3273), .Z(n1382) );
  IV U6285 ( .A(n3270), .Z(n3273) );
  XNOR U6286 ( .A(n3199), .B(n1390), .Z(n3274) );
  XOR U6287 ( .A(n3275), .B(n3276), .Z(n3270) );
  AND U6288 ( .A(n1420), .B(n3277), .Z(n3276) );
  XNOR U6289 ( .A(n3278), .B(n1421), .Z(n3277) );
  NANDN U6290 ( .B(n3192), .A(reg_source[14]), .Z(n1421) );
  XNOR U6291 ( .A(n3279), .B(n3278), .Z(n1420) );
  IV U6292 ( .A(n3275), .Z(n3278) );
  XNOR U6293 ( .A(n3199), .B(n1428), .Z(n3279) );
  XOR U6294 ( .A(n3280), .B(n3281), .Z(n3275) );
  AND U6295 ( .A(n1306), .B(n3282), .Z(n3281) );
  XNOR U6296 ( .A(n3283), .B(n1307), .Z(n3282) );
  NANDN U6297 ( .B(n3192), .A(reg_source[13]), .Z(n1307) );
  XNOR U6298 ( .A(n3284), .B(n3283), .Z(n1306) );
  IV U6299 ( .A(n3280), .Z(n3283) );
  XNOR U6300 ( .A(n3199), .B(n1314), .Z(n3284) );
  XOR U6301 ( .A(n3285), .B(n3286), .Z(n3280) );
  AND U6302 ( .A(n1343), .B(n3287), .Z(n3286) );
  XNOR U6303 ( .A(n3288), .B(n1344), .Z(n3287) );
  NANDN U6304 ( .B(n3192), .A(reg_source[12]), .Z(n1344) );
  XNOR U6305 ( .A(n3289), .B(n3288), .Z(n1343) );
  IV U6306 ( .A(n3285), .Z(n3288) );
  XNOR U6307 ( .A(n3199), .B(n1351), .Z(n3289) );
  XOR U6308 ( .A(n3290), .B(n3291), .Z(n3285) );
  AND U6309 ( .A(n1226), .B(n3292), .Z(n3291) );
  XNOR U6310 ( .A(n3293), .B(n1227), .Z(n3292) );
  NANDN U6311 ( .B(n3192), .A(reg_source[11]), .Z(n1227) );
  XNOR U6312 ( .A(n3294), .B(n3293), .Z(n1226) );
  IV U6313 ( .A(n3290), .Z(n3293) );
  XNOR U6314 ( .A(n3199), .B(n1234), .Z(n3294) );
  XOR U6315 ( .A(n3295), .B(n3296), .Z(n3290) );
  AND U6316 ( .A(n1265), .B(n3297), .Z(n3296) );
  XNOR U6317 ( .A(n3298), .B(n1266), .Z(n3297) );
  NANDN U6318 ( .B(n3192), .A(reg_source[10]), .Z(n1266) );
  XNOR U6319 ( .A(n3299), .B(n3298), .Z(n1265) );
  IV U6320 ( .A(n3295), .Z(n3298) );
  XNOR U6321 ( .A(n3199), .B(n1273), .Z(n3299) );
  XOR U6322 ( .A(n3300), .B(n3301), .Z(n3295) );
  AND U6323 ( .A(n1141), .B(n3302), .Z(n3301) );
  XNOR U6324 ( .A(n3303), .B(n1142), .Z(n3302) );
  NANDN U6325 ( .B(n3192), .A(reg_source[9]), .Z(n1142) );
  XNOR U6326 ( .A(n3304), .B(n3303), .Z(n1141) );
  IV U6327 ( .A(n3300), .Z(n3303) );
  XNOR U6328 ( .A(n3199), .B(n1152), .Z(n3304) );
  XOR U6329 ( .A(n3305), .B(n3306), .Z(n3300) );
  AND U6330 ( .A(n1184), .B(n3307), .Z(n3306) );
  XNOR U6331 ( .A(n3308), .B(n1185), .Z(n3307) );
  NANDN U6332 ( .B(n3192), .A(reg_source[8]), .Z(n1185) );
  XNOR U6333 ( .A(n3309), .B(n3308), .Z(n1184) );
  IV U6334 ( .A(n3305), .Z(n3308) );
  XNOR U6335 ( .A(n3199), .B(n1192), .Z(n3309) );
  XOR U6336 ( .A(n3310), .B(n3311), .Z(n3305) );
  AND U6337 ( .A(n3312), .B(n3313), .Z(n3311) );
  XNOR U6338 ( .A(n3314), .B(n3315), .Z(n3313) );
  XNOR U6339 ( .A(n3199), .B(n1810), .Z(n3193) );
  ANDN U6340 ( .A(reg_source[31]), .B(n3192), .Z(n3187) );
  AND U6341 ( .A(n3316), .B(n3317), .Z(n3123) );
  AND U6342 ( .A(n3318), .B(n3319), .Z(n3317) );
  NAND U6343 ( .A(n3320), .B(n1140), .Z(n3319) );
  NAND U6344 ( .A(n3321), .B(n1154), .Z(n3318) );
  ANDN U6345 ( .A(b_bus[0]), .B(n3132), .Z(n3321) );
  AND U6346 ( .A(n3322), .B(n3323), .Z(n3316) );
  NAND U6347 ( .A(n3320), .B(n1151), .Z(n3323) );
  XNOR U6348 ( .A(n3132), .B(b_bus[0]), .Z(n3320) );
  IV U6349 ( .A(n3167), .Z(b_bus[0]) );
  MUX U6350 ( .IN0(n1145), .IN1(n1146), .SEL(n3324), .F(n3322) );
  ANDN U6351 ( .A(n3167), .B(a_bus[0]), .Z(n3324) );
  NOR U6352 ( .A(n3076), .B(n3325), .Z(n3116) );
  ANDN U6353 ( .A(n1924), .B(n3103), .Z(n3325) );
  ANDN U6354 ( .A(n399), .B(n1882), .Z(n1924) );
  OR U6355 ( .A(n774), .B(n3326), .Z(n1882) );
  NAND U6356 ( .A(n3327), .B(n3328), .Z(n774) );
  NAND U6357 ( .A(n3329), .B(n3330), .Z(n3328) );
  OR U6358 ( .A(n1086), .B(n671), .Z(n3329) );
  NANDN U6359 ( .B(n660), .A(n3331), .Z(n3327) );
  NAND U6360 ( .A(n3332), .B(n3333), .Z(n3331) );
  ANDN U6361 ( .A(n3334), .B(n671), .Z(n3333) );
  NOR U6362 ( .A(n791), .B(n1086), .Z(n3332) );
  NANDN U6363 ( .B(n143), .A(n3335), .Z(n1086) );
  AND U6364 ( .A(n3336), .B(n3337), .Z(n399) );
  AND U6365 ( .A(n3338), .B(n3339), .Z(n3337) );
  AND U6366 ( .A(n3340), .B(n3341), .Z(n3339) );
  NAND U6367 ( .A(n3342), .B(n1109), .Z(n3341) );
  NAND U6368 ( .A(n3343), .B(n3344), .Z(n3342) );
  AND U6369 ( .A(n3345), .B(n3346), .Z(n3344) );
  AND U6370 ( .A(n3347), .B(n3348), .Z(n3345) );
  OR U6371 ( .A(n1445), .B(n1117), .Z(n3348) );
  AND U6372 ( .A(n3349), .B(n3350), .Z(n1445) );
  AND U6373 ( .A(n3351), .B(n3352), .Z(n3350) );
  NAND U6374 ( .A(n1133), .B(n1650), .Z(n3352) );
  AND U6375 ( .A(n3353), .B(n3354), .Z(n3349) );
  NAND U6376 ( .A(n1654), .B(n3159), .Z(n3353) );
  AND U6377 ( .A(n3355), .B(n3356), .Z(n3343) );
  NAND U6378 ( .A(n3357), .B(n1118), .Z(n3356) );
  NAND U6379 ( .A(n3358), .B(n1121), .Z(n3340) );
  NAND U6380 ( .A(n3359), .B(n3360), .Z(n3358) );
  AND U6381 ( .A(n3361), .B(n3346), .Z(n3360) );
  NAND U6382 ( .A(n1119), .B(n1132), .Z(n3346) );
  AND U6383 ( .A(n3347), .B(n3362), .Z(n3361) );
  OR U6384 ( .A(n1447), .B(n1117), .Z(n3362) );
  AND U6385 ( .A(n3363), .B(n3364), .Z(n1447) );
  AND U6386 ( .A(n3351), .B(n3365), .Z(n3364) );
  NAND U6387 ( .A(n1415), .B(n1133), .Z(n3365) );
  NAND U6388 ( .A(n1125), .B(n1653), .Z(n3351) );
  AND U6389 ( .A(n3366), .B(n3354), .Z(n3363) );
  NAND U6390 ( .A(n1302), .B(n3158), .Z(n3354) );
  NAND U6391 ( .A(n1301), .B(n3159), .Z(n3366) );
  NANDN U6392 ( .B(n3367), .A(n1134), .Z(n3347) );
  AND U6393 ( .A(n3355), .B(n3368), .Z(n3359) );
  NAND U6394 ( .A(n3357), .B(n1129), .Z(n3368) );
  NAND U6395 ( .A(n3369), .B(n3370), .Z(n3357) );
  AND U6396 ( .A(n3371), .B(n3372), .Z(n3370) );
  OR U6397 ( .A(n3166), .B(n3169), .Z(n3372) );
  OR U6398 ( .A(n3168), .B(n3175), .Z(n3371) );
  AND U6399 ( .A(n3373), .B(n3374), .Z(n3369) );
  OR U6400 ( .A(n3172), .B(n3375), .Z(n3374) );
  OR U6401 ( .A(n3174), .B(n3173), .Z(n3373) );
  NAND U6402 ( .A(n1135), .B(n1124), .Z(n3355) );
  AND U6403 ( .A(n3376), .B(n3377), .Z(n3338) );
  NAND U6404 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][1] ), .Z(n3377) );
  AND U6405 ( .A(\Shifter/sll_27/ML_int[3][1] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][1] ) );
  AND U6406 ( .A(\Shifter/sll_27/ML_int[2][1] ), .B(n3130), .Z(
        \Shifter/sll_27/ML_int[3][1] ) );
  AND U6407 ( .A(\Shifter/sll_27/ML_int[1][1] ), .B(n3131), .Z(
        \Shifter/sll_27/ML_int[2][1] ) );
  NAND U6408 ( .A(n3378), .B(n1140), .Z(n3376) );
  XOR U6409 ( .A(n3379), .B(a_bus[1]), .Z(n3378) );
  AND U6410 ( .A(n3380), .B(n3381), .Z(n3336) );
  MUX U6411 ( .IN0(n1145), .IN1(n1146), .SEL(n3382), .F(n3381) );
  ANDN U6412 ( .A(n3169), .B(a_bus[1]), .Z(n3382) );
  AND U6413 ( .A(n3383), .B(n3384), .Z(n3380) );
  NAND U6414 ( .A(n3385), .B(n1151), .Z(n3384) );
  XNOR U6415 ( .A(n3131), .B(b_bus[1]), .Z(n3385) );
  NAND U6416 ( .A(n3386), .B(n1154), .Z(n3383) );
  ANDN U6417 ( .A(b_bus[1]), .B(n3131), .Z(n3386) );
  IV U6418 ( .A(n3169), .Z(b_bus[1]) );
  AND U6419 ( .A(n1902), .B(n3118), .Z(n3076) );
  IV U6420 ( .A(n3103), .Z(n3118) );
  NAND U6421 ( .A(n2039), .B(n2932), .Z(n3103) );
  ANDN U6422 ( .A(n2478), .B(n485), .Z(n2932) );
  AND U6423 ( .A(n3387), .B(n3388), .Z(n485) );
  AND U6424 ( .A(n3389), .B(n3390), .Z(n3388) );
  AND U6425 ( .A(n3391), .B(n3392), .Z(n3390) );
  NAND U6426 ( .A(n3393), .B(n1109), .Z(n3392) );
  NAND U6427 ( .A(n3394), .B(n3395), .Z(n3393) );
  AND U6428 ( .A(n3396), .B(n3397), .Z(n3395) );
  AND U6429 ( .A(n3398), .B(n3399), .Z(n3396) );
  OR U6430 ( .A(n1595), .B(n1117), .Z(n3399) );
  AND U6431 ( .A(n3400), .B(n3401), .Z(n1595) );
  NAND U6432 ( .A(n1222), .B(n1650), .Z(n3401) );
  ANDN U6433 ( .A(n3402), .B(n1652), .Z(n3400) );
  NAND U6434 ( .A(n1369), .B(n1653), .Z(n3402) );
  NANDN U6435 ( .B(n3403), .A(n1118), .Z(n3398) );
  NAND U6436 ( .A(n3404), .B(n1121), .Z(n3391) );
  NAND U6437 ( .A(n3394), .B(n3405), .Z(n3404) );
  AND U6438 ( .A(n3406), .B(n3397), .Z(n3405) );
  NAND U6439 ( .A(n1124), .B(n1216), .Z(n3397) );
  AND U6440 ( .A(n3407), .B(n3408), .Z(n3406) );
  OR U6441 ( .A(n1597), .B(n1117), .Z(n3408) );
  AND U6442 ( .A(n3409), .B(n3410), .Z(n1597) );
  NAND U6443 ( .A(n1415), .B(n1222), .Z(n3410) );
  AND U6444 ( .A(n3411), .B(n3412), .Z(n3409) );
  NANDN U6445 ( .B(n1378), .A(n1653), .Z(n3412) );
  NANDN U6446 ( .B(n1377), .A(n3158), .Z(n3411) );
  NANDN U6447 ( .B(n3403), .A(n1129), .Z(n3407) );
  AND U6448 ( .A(n3413), .B(n3414), .Z(n3394) );
  NAND U6449 ( .A(n1132), .B(n1218), .Z(n3414) );
  NAND U6450 ( .A(n1134), .B(n1209), .Z(n3413) );
  AND U6451 ( .A(n3415), .B(n3416), .Z(n3389) );
  NAND U6452 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][7] ), .Z(n3416) );
  AND U6453 ( .A(\Shifter/sll_27/ML_int[3][7] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][7] ) );
  NAND U6454 ( .A(n3417), .B(n1140), .Z(n3415) );
  XNOR U6455 ( .A(n3312), .B(n3315), .Z(n3417) );
  XNOR U6456 ( .A(n3418), .B(n3314), .Z(n3312) );
  IV U6457 ( .A(n3310), .Z(n3314) );
  XOR U6458 ( .A(n3419), .B(n3420), .Z(n3310) );
  AND U6459 ( .A(n3421), .B(n3422), .Z(n3420) );
  XNOR U6460 ( .A(n3423), .B(n3424), .Z(n3422) );
  XNOR U6461 ( .A(n3199), .B(n3425), .Z(n3418) );
  AND U6462 ( .A(n3426), .B(n3427), .Z(n3387) );
  MUX U6463 ( .IN0(n1145), .IN1(n1146), .SEL(n3428), .F(n3427) );
  ANDN U6464 ( .A(n3315), .B(b_bus[7]), .Z(n3428) );
  AND U6465 ( .A(n3429), .B(n3430), .Z(n3426) );
  NAND U6466 ( .A(n3431), .B(n1151), .Z(n3430) );
  XNOR U6467 ( .A(n3315), .B(b_bus[7]), .Z(n3431) );
  IV U6468 ( .A(n3425), .Z(b_bus[7]) );
  NANDN U6469 ( .B(n3315), .A(n3432), .Z(n3429) );
  ANDN U6470 ( .A(n1154), .B(n3425), .Z(n3432) );
  NANDN U6471 ( .B(n3192), .A(reg_source[7]), .Z(n3315) );
  AND U6472 ( .A(N25), .B(N26), .Z(n2478) );
  IV U6473 ( .A(n532), .Z(N26) );
  AND U6474 ( .A(n3433), .B(n3434), .Z(n532) );
  AND U6475 ( .A(n3435), .B(n3436), .Z(n3434) );
  AND U6476 ( .A(n3437), .B(n3438), .Z(n3436) );
  NAND U6477 ( .A(n3439), .B(n1109), .Z(n3438) );
  NAND U6478 ( .A(n3440), .B(n3441), .Z(n3439) );
  AND U6479 ( .A(n3442), .B(n3443), .Z(n3441) );
  AND U6480 ( .A(n3444), .B(n3445), .Z(n3442) );
  OR U6481 ( .A(n1546), .B(n1117), .Z(n3445) );
  AND U6482 ( .A(n3446), .B(n3447), .Z(n1546) );
  AND U6483 ( .A(n3448), .B(n3449), .Z(n3447) );
  NAND U6484 ( .A(n1125), .B(n1650), .Z(n3449) );
  AND U6485 ( .A(n3450), .B(n3451), .Z(n3446) );
  NAND U6486 ( .A(n3158), .B(n1654), .Z(n3450) );
  NAND U6487 ( .A(n3452), .B(n3453), .Z(n1654) );
  NANDN U6488 ( .B(n1810), .A(a_bus[1]), .Z(n3453) );
  AND U6489 ( .A(n3454), .B(n3455), .Z(n3452) );
  NANDN U6490 ( .B(n3367), .A(n1118), .Z(n3444) );
  NAND U6491 ( .A(n3456), .B(n1121), .Z(n3437) );
  NAND U6492 ( .A(n3440), .B(n3457), .Z(n3456) );
  AND U6493 ( .A(n3458), .B(n3443), .Z(n3457) );
  NAND U6494 ( .A(n1124), .B(n1133), .Z(n3443) );
  NAND U6495 ( .A(n3459), .B(n3460), .Z(n1133) );
  AND U6496 ( .A(n3461), .B(n3462), .Z(n3460) );
  OR U6497 ( .A(n3166), .B(n1460), .Z(n3462) );
  OR U6498 ( .A(n3168), .B(n1533), .Z(n3461) );
  AND U6499 ( .A(n3463), .B(n3464), .Z(n3459) );
  OR U6500 ( .A(n3172), .B(n1584), .Z(n3464) );
  OR U6501 ( .A(n3174), .B(n1509), .Z(n3463) );
  AND U6502 ( .A(n3465), .B(n3466), .Z(n3458) );
  OR U6503 ( .A(n1548), .B(n1117), .Z(n3466) );
  AND U6504 ( .A(n3467), .B(n3468), .Z(n1548) );
  NAND U6505 ( .A(n1415), .B(n1125), .Z(n3468) );
  NAND U6506 ( .A(n3469), .B(n3470), .Z(n1125) );
  AND U6507 ( .A(n3471), .B(n3472), .Z(n3470) );
  OR U6508 ( .A(n3166), .B(n1560), .Z(n3472) );
  OR U6509 ( .A(n3168), .B(n1633), .Z(n3471) );
  AND U6510 ( .A(n3473), .B(n3474), .Z(n3469) );
  OR U6511 ( .A(n3172), .B(n1695), .Z(n3474) );
  OR U6512 ( .A(n3174), .B(n1609), .Z(n3473) );
  AND U6513 ( .A(n3475), .B(n3451), .Z(n3467) );
  NAND U6514 ( .A(n1653), .B(n1302), .Z(n3451) );
  NAND U6515 ( .A(n3476), .B(n3477), .Z(n1302) );
  AND U6516 ( .A(n3478), .B(n3479), .Z(n3477) );
  OR U6517 ( .A(n3166), .B(n1669), .Z(n3479) );
  OR U6518 ( .A(n3168), .B(n1749), .Z(n3478) );
  AND U6519 ( .A(n3480), .B(n3481), .Z(n3476) );
  OR U6520 ( .A(n3172), .B(n1798), .Z(n3481) );
  OR U6521 ( .A(n3174), .B(n1721), .Z(n3480) );
  NAND U6522 ( .A(n1301), .B(n3158), .Z(n3475) );
  NAND U6523 ( .A(n3482), .B(n3455), .Z(n1301) );
  OR U6524 ( .A(n3166), .B(n1775), .Z(n3455) );
  AND U6525 ( .A(n3483), .B(n3454), .Z(n3482) );
  OR U6526 ( .A(n3168), .B(n1824), .Z(n3454) );
  OR U6527 ( .A(n3174), .B(n1810), .Z(n3483) );
  NANDN U6528 ( .B(n3367), .A(n1129), .Z(n3465) );
  AND U6529 ( .A(n3484), .B(n3485), .Z(n3367) );
  AND U6530 ( .A(n3486), .B(n3487), .Z(n3485) );
  OR U6531 ( .A(n3166), .B(n3488), .Z(n3487) );
  OR U6532 ( .A(n3168), .B(n3489), .Z(n3486) );
  AND U6533 ( .A(n3490), .B(n3491), .Z(n3484) );
  OR U6534 ( .A(n3172), .B(n1192), .Z(n3491) );
  OR U6535 ( .A(n3174), .B(n3425), .Z(n3490) );
  AND U6536 ( .A(n3492), .B(n3493), .Z(n3440) );
  NAND U6537 ( .A(n1132), .B(n1135), .Z(n3493) );
  NAND U6538 ( .A(n3494), .B(n3495), .Z(n1135) );
  AND U6539 ( .A(n3496), .B(n3497), .Z(n3495) );
  OR U6540 ( .A(n3166), .B(n1314), .Z(n3497) );
  OR U6541 ( .A(n3168), .B(n1428), .Z(n3496) );
  AND U6542 ( .A(n3498), .B(n3499), .Z(n3494) );
  OR U6543 ( .A(n3172), .B(n1484), .Z(n3499) );
  OR U6544 ( .A(n3174), .B(n1390), .Z(n3498) );
  NAND U6545 ( .A(n1134), .B(n1119), .Z(n3492) );
  NAND U6546 ( .A(n3500), .B(n3501), .Z(n1119) );
  AND U6547 ( .A(n3502), .B(n3503), .Z(n3501) );
  OR U6548 ( .A(n3166), .B(n1152), .Z(n3503) );
  OR U6549 ( .A(n3168), .B(n1273), .Z(n3502) );
  AND U6550 ( .A(n3504), .B(n3505), .Z(n3500) );
  OR U6551 ( .A(n3172), .B(n1351), .Z(n3505) );
  OR U6552 ( .A(n3174), .B(n1234), .Z(n3504) );
  AND U6553 ( .A(n3506), .B(n3507), .Z(n3435) );
  NAND U6554 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][5] ), .Z(n3507) );
  AND U6555 ( .A(\Shifter/sll_27/ML_int[3][5] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][5] ) );
  NAND U6556 ( .A(n3508), .B(n1140), .Z(n3506) );
  XNOR U6557 ( .A(n3509), .B(n3510), .Z(n3508) );
  AND U6558 ( .A(n3511), .B(n3512), .Z(n3433) );
  MUX U6559 ( .IN0(n1145), .IN1(n1146), .SEL(n3513), .F(n3512) );
  ANDN U6560 ( .A(n3510), .B(b_bus[5]), .Z(n3513) );
  AND U6561 ( .A(n3514), .B(n3515), .Z(n3511) );
  NAND U6562 ( .A(n3516), .B(n1151), .Z(n3515) );
  XNOR U6563 ( .A(n3510), .B(b_bus[5]), .Z(n3516) );
  IV U6564 ( .A(n3488), .Z(b_bus[5]) );
  NANDN U6565 ( .B(n3510), .A(n3517), .Z(n3514) );
  ANDN U6566 ( .A(n1154), .B(n3488), .Z(n3517) );
  IV U6567 ( .A(n511), .Z(N25) );
  AND U6568 ( .A(n3518), .B(n3519), .Z(n511) );
  AND U6569 ( .A(n3520), .B(n3521), .Z(n3519) );
  AND U6570 ( .A(n3522), .B(n3523), .Z(n3521) );
  NAND U6571 ( .A(n3524), .B(n1109), .Z(n3523) );
  NAND U6572 ( .A(n3525), .B(n3526), .Z(n3524) );
  AND U6573 ( .A(n3527), .B(n3528), .Z(n3526) );
  AND U6574 ( .A(n3529), .B(n3530), .Z(n3527) );
  OR U6575 ( .A(n1619), .B(n1117), .Z(n3530) );
  AND U6576 ( .A(n3531), .B(n3532), .Z(n1619) );
  AND U6577 ( .A(n3533), .B(n3534), .Z(n3532) );
  NAND U6578 ( .A(n1254), .B(n1650), .Z(n3534) );
  AND U6579 ( .A(n3448), .B(n3535), .Z(n3531) );
  NAND U6580 ( .A(n1734), .B(n3158), .Z(n3535) );
  NAND U6581 ( .A(n1118), .B(n3536), .Z(n3529) );
  NAND U6582 ( .A(n3537), .B(n1121), .Z(n3522) );
  NAND U6583 ( .A(n3525), .B(n3538), .Z(n3537) );
  AND U6584 ( .A(n3539), .B(n3528), .Z(n3538) );
  NAND U6585 ( .A(n1124), .B(n1260), .Z(n3528) );
  AND U6586 ( .A(n3540), .B(n3541), .Z(n3539) );
  OR U6587 ( .A(n1621), .B(n1117), .Z(n3541) );
  AND U6588 ( .A(n3542), .B(n3543), .Z(n1621) );
  NAND U6589 ( .A(n1415), .B(n1254), .Z(n3543) );
  AND U6590 ( .A(n3544), .B(n3533), .Z(n3542) );
  NAND U6591 ( .A(n1416), .B(n1653), .Z(n3533) );
  NAND U6592 ( .A(n1414), .B(n3158), .Z(n3544) );
  NAND U6593 ( .A(n1129), .B(n3536), .Z(n3540) );
  AND U6594 ( .A(n3545), .B(n3546), .Z(n3525) );
  NAND U6595 ( .A(n1132), .B(n1261), .Z(n3546) );
  NAND U6596 ( .A(n1134), .B(n1250), .Z(n3545) );
  AND U6597 ( .A(n3547), .B(n3548), .Z(n3520) );
  NAND U6598 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][6] ), .Z(n3548) );
  AND U6599 ( .A(\Shifter/sll_27/ML_int[3][6] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][6] ) );
  NAND U6600 ( .A(n3549), .B(n1140), .Z(n3547) );
  XNOR U6601 ( .A(n3421), .B(n3424), .Z(n3549) );
  XNOR U6602 ( .A(n3550), .B(n3423), .Z(n3421) );
  IV U6603 ( .A(n3419), .Z(n3423) );
  XOR U6604 ( .A(n3551), .B(n3552), .Z(n3419) );
  AND U6605 ( .A(n3509), .B(n3553), .Z(n3552) );
  XNOR U6606 ( .A(n3554), .B(n3510), .Z(n3553) );
  NANDN U6607 ( .B(n3192), .A(reg_source[5]), .Z(n3510) );
  XNOR U6608 ( .A(n3555), .B(n3554), .Z(n3509) );
  IV U6609 ( .A(n3551), .Z(n3554) );
  XNOR U6610 ( .A(n3199), .B(n3488), .Z(n3555) );
  XOR U6611 ( .A(n3556), .B(n3557), .Z(n3551) );
  AND U6612 ( .A(n3558), .B(n3559), .Z(n3557) );
  XNOR U6613 ( .A(n3560), .B(n1117), .Z(n3559) );
  XNOR U6614 ( .A(n3199), .B(n3489), .Z(n3550) );
  AND U6615 ( .A(n3561), .B(n3562), .Z(n3518) );
  MUX U6616 ( .IN0(n1145), .IN1(n1146), .SEL(n3563), .F(n3562) );
  ANDN U6617 ( .A(n3424), .B(b_bus[6]), .Z(n3563) );
  AND U6618 ( .A(n3564), .B(n3565), .Z(n3561) );
  NAND U6619 ( .A(n3566), .B(n1151), .Z(n3565) );
  XNOR U6620 ( .A(n3424), .B(b_bus[6]), .Z(n3566) );
  IV U6621 ( .A(n3489), .Z(b_bus[6]) );
  NANDN U6622 ( .B(n3424), .A(n3567), .Z(n3564) );
  ANDN U6623 ( .A(n1154), .B(n3489), .Z(n3567) );
  NANDN U6624 ( .B(n3192), .A(reg_source[6]), .Z(n3424) );
  ANDN U6625 ( .A(n2990), .B(n553), .Z(n2039) );
  AND U6626 ( .A(n3568), .B(n3569), .Z(n553) );
  AND U6627 ( .A(n3570), .B(n3571), .Z(n3569) );
  NAND U6628 ( .A(n3572), .B(n1140), .Z(n3571) );
  XOR U6629 ( .A(n3558), .B(a_bus[4]), .Z(n3572) );
  XNOR U6630 ( .A(n3573), .B(n3560), .Z(n3558) );
  IV U6631 ( .A(n3556), .Z(n3560) );
  XOR U6632 ( .A(n3574), .B(n3575), .Z(n3556) );
  AND U6633 ( .A(n3576), .B(n3577), .Z(n3575) );
  XNOR U6634 ( .A(n3578), .B(n3129), .Z(n3577) );
  XNOR U6635 ( .A(n3199), .B(n3375), .Z(n3573) );
  AND U6636 ( .A(n3579), .B(n3580), .Z(n3570) );
  NAND U6637 ( .A(n3581), .B(n1109), .Z(n3580) );
  NAND U6638 ( .A(n3582), .B(n3583), .Z(n3581) );
  AND U6639 ( .A(n3584), .B(n3585), .Z(n3583) );
  AND U6640 ( .A(n3586), .B(n3587), .Z(n3584) );
  OR U6641 ( .A(n1570), .B(n1117), .Z(n3587) );
  AND U6642 ( .A(n3588), .B(n3589), .Z(n1570) );
  AND U6643 ( .A(n3448), .B(n3590), .Z(n3589) );
  NAND U6644 ( .A(n1173), .B(n1650), .Z(n3590) );
  NANDN U6645 ( .B(n3160), .A(n1118), .Z(n3586) );
  NAND U6646 ( .A(n3591), .B(n1121), .Z(n3579) );
  NAND U6647 ( .A(n3582), .B(n3592), .Z(n3591) );
  AND U6648 ( .A(n3593), .B(n3585), .Z(n3592) );
  NAND U6649 ( .A(n1124), .B(n1179), .Z(n3585) );
  NAND U6650 ( .A(n3594), .B(n3595), .Z(n1179) );
  AND U6651 ( .A(n3596), .B(n3597), .Z(n3595) );
  OR U6652 ( .A(n3166), .B(n1484), .Z(n3597) );
  OR U6653 ( .A(n3168), .B(n1460), .Z(n3596) );
  AND U6654 ( .A(n3598), .B(n3599), .Z(n3594) );
  OR U6655 ( .A(n3172), .B(n1509), .Z(n3599) );
  OR U6656 ( .A(n3174), .B(n1533), .Z(n3598) );
  AND U6657 ( .A(n3600), .B(n3601), .Z(n3593) );
  OR U6658 ( .A(n1572), .B(n1117), .Z(n3601) );
  AND U6659 ( .A(n3588), .B(n3602), .Z(n1572) );
  NAND U6660 ( .A(n1415), .B(n1173), .Z(n3602) );
  NAND U6661 ( .A(n3603), .B(n3604), .Z(n1173) );
  AND U6662 ( .A(n3605), .B(n3606), .Z(n3604) );
  OR U6663 ( .A(n3166), .B(n1584), .Z(n3606) );
  OR U6664 ( .A(n3168), .B(n1560), .Z(n3605) );
  AND U6665 ( .A(n3607), .B(n3608), .Z(n3603) );
  OR U6666 ( .A(n3172), .B(n1609), .Z(n3608) );
  OR U6667 ( .A(n3174), .B(n1633), .Z(n3607) );
  AND U6668 ( .A(n3609), .B(n3610), .Z(n3588) );
  NAND U6669 ( .A(n1339), .B(n1653), .Z(n3610) );
  NAND U6670 ( .A(n3611), .B(n3612), .Z(n1339) );
  AND U6671 ( .A(n3613), .B(n3614), .Z(n3612) );
  OR U6672 ( .A(n3166), .B(n1695), .Z(n3614) );
  OR U6673 ( .A(n3168), .B(n1669), .Z(n3613) );
  AND U6674 ( .A(n3615), .B(n3616), .Z(n3611) );
  OR U6675 ( .A(n3172), .B(n1721), .Z(n3616) );
  OR U6676 ( .A(n3174), .B(n1749), .Z(n3615) );
  NAND U6677 ( .A(n3158), .B(n1338), .Z(n3609) );
  NAND U6678 ( .A(n3617), .B(n3618), .Z(n1338) );
  AND U6679 ( .A(n3619), .B(n3620), .Z(n3618) );
  OR U6680 ( .A(n3166), .B(n1798), .Z(n3620) );
  OR U6681 ( .A(n3168), .B(n1775), .Z(n3619) );
  AND U6682 ( .A(n3621), .B(n3622), .Z(n3617) );
  OR U6683 ( .A(n3172), .B(n1810), .Z(n3622) );
  OR U6684 ( .A(n3174), .B(n1824), .Z(n3621) );
  NANDN U6685 ( .B(n3160), .A(n1129), .Z(n3600) );
  AND U6686 ( .A(n3623), .B(n3624), .Z(n3160) );
  AND U6687 ( .A(n3625), .B(n3626), .Z(n3624) );
  OR U6688 ( .A(n3166), .B(n3375), .Z(n3626) );
  OR U6689 ( .A(n3168), .B(n3488), .Z(n3625) );
  AND U6690 ( .A(n3627), .B(n3628), .Z(n3623) );
  OR U6691 ( .A(n3172), .B(n3425), .Z(n3628) );
  OR U6692 ( .A(n3174), .B(n3489), .Z(n3627) );
  AND U6693 ( .A(n3629), .B(n3630), .Z(n3582) );
  NAND U6694 ( .A(n1132), .B(n1180), .Z(n3630) );
  NAND U6695 ( .A(n3631), .B(n3632), .Z(n1180) );
  AND U6696 ( .A(n3633), .B(n3634), .Z(n3632) );
  OR U6697 ( .A(n3166), .B(n1351), .Z(n3634) );
  OR U6698 ( .A(n3168), .B(n1314), .Z(n3633) );
  AND U6699 ( .A(n3635), .B(n3636), .Z(n3631) );
  OR U6700 ( .A(n3172), .B(n1390), .Z(n3636) );
  OR U6701 ( .A(n3174), .B(n1428), .Z(n3635) );
  NAND U6702 ( .A(n1134), .B(n1169), .Z(n3629) );
  NAND U6703 ( .A(n3637), .B(n3638), .Z(n1169) );
  AND U6704 ( .A(n3639), .B(n3640), .Z(n3638) );
  OR U6705 ( .A(n3166), .B(n1192), .Z(n3640) );
  OR U6706 ( .A(n3168), .B(n1152), .Z(n3639) );
  AND U6707 ( .A(n3641), .B(n3642), .Z(n3637) );
  OR U6708 ( .A(n3172), .B(n1234), .Z(n3642) );
  OR U6709 ( .A(n3174), .B(n1273), .Z(n3641) );
  AND U6710 ( .A(n3643), .B(n3644), .Z(n3568) );
  AND U6711 ( .A(n3645), .B(n3646), .Z(n3644) );
  NAND U6712 ( .A(n3647), .B(n1151), .Z(n3646) );
  XNOR U6713 ( .A(n1117), .B(b_bus[4]), .Z(n3647) );
  IV U6714 ( .A(n3375), .Z(b_bus[4]) );
  MUX U6715 ( .IN0(n1145), .IN1(n1146), .SEL(n3648), .F(n3645) );
  ANDN U6716 ( .A(n3375), .B(a_bus[4]), .Z(n3648) );
  MUX U6717 ( .IN0(n3649), .IN1(n3650), .SEL(n1117), .F(n3643) );
  NANDN U6718 ( .B(n1450), .A(\Shifter/sll_27/ML_int[4][4] ), .Z(n3650) );
  AND U6719 ( .A(\Shifter/sll_27/ML_int[3][4] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][4] ) );
  NANDN U6720 ( .B(n3375), .A(n1154), .Z(n3649) );
  AND U6721 ( .A(N28), .B(N29), .Z(n2990) );
  IV U6722 ( .A(n595), .Z(N29) );
  AND U6723 ( .A(n3651), .B(n3652), .Z(n595) );
  AND U6724 ( .A(n3653), .B(n3654), .Z(n3652) );
  AND U6725 ( .A(n3655), .B(n3656), .Z(n3654) );
  NAND U6726 ( .A(n3657), .B(n1109), .Z(n3656) );
  NAND U6727 ( .A(n3658), .B(n3659), .Z(n3657) );
  AND U6728 ( .A(n3660), .B(n3661), .Z(n3659) );
  AND U6729 ( .A(n3662), .B(n3663), .Z(n3660) );
  OR U6730 ( .A(n1519), .B(n1117), .Z(n3663) );
  AND U6731 ( .A(n3664), .B(n3665), .Z(n1519) );
  AND U6732 ( .A(n3666), .B(n3667), .Z(n3665) );
  NAND U6733 ( .A(n1260), .B(n1650), .Z(n3667) );
  AND U6734 ( .A(n3668), .B(n3669), .Z(n3664) );
  NAND U6735 ( .A(n3159), .B(n1734), .Z(n3668) );
  MUX U6736 ( .IN0(b_bus[30]), .IN1(\Shifter/N75 ), .SEL(n3166), .F(n1734) );
  IV U6737 ( .A(n1824), .Z(b_bus[30]) );
  AND U6738 ( .A(n3670), .B(n3671), .Z(n3658) );
  NAND U6739 ( .A(n3672), .B(n1118), .Z(n3671) );
  NAND U6740 ( .A(n3673), .B(n1121), .Z(n3655) );
  NAND U6741 ( .A(n3674), .B(n3675), .Z(n3673) );
  AND U6742 ( .A(n3676), .B(n3661), .Z(n3675) );
  NAND U6743 ( .A(n1250), .B(n1132), .Z(n3661) );
  NAND U6744 ( .A(n3677), .B(n3678), .Z(n1250) );
  AND U6745 ( .A(n3679), .B(n3680), .Z(n3678) );
  OR U6746 ( .A(n3166), .B(n1273), .Z(n3680) );
  OR U6747 ( .A(n3168), .B(n1234), .Z(n3679) );
  AND U6748 ( .A(n3681), .B(n3682), .Z(n3677) );
  OR U6749 ( .A(n3172), .B(n1314), .Z(n3682) );
  OR U6750 ( .A(n3174), .B(n1351), .Z(n3681) );
  AND U6751 ( .A(n3662), .B(n3683), .Z(n3676) );
  OR U6752 ( .A(n1521), .B(n1117), .Z(n3683) );
  AND U6753 ( .A(n3684), .B(n3685), .Z(n1521) );
  AND U6754 ( .A(n3666), .B(n3686), .Z(n3685) );
  NAND U6755 ( .A(n1415), .B(n1260), .Z(n3686) );
  NAND U6756 ( .A(n3687), .B(n3688), .Z(n1260) );
  AND U6757 ( .A(n3689), .B(n3690), .Z(n3688) );
  OR U6758 ( .A(n3166), .B(n1533), .Z(n3690) );
  OR U6759 ( .A(n3168), .B(n1509), .Z(n3689) );
  AND U6760 ( .A(n3691), .B(n3692), .Z(n3687) );
  OR U6761 ( .A(n3172), .B(n1560), .Z(n3692) );
  OR U6762 ( .A(n3174), .B(n1584), .Z(n3691) );
  NAND U6763 ( .A(n1254), .B(n1653), .Z(n3666) );
  NAND U6764 ( .A(n3693), .B(n3694), .Z(n1254) );
  AND U6765 ( .A(n3695), .B(n3696), .Z(n3694) );
  OR U6766 ( .A(n3166), .B(n1633), .Z(n3696) );
  OR U6767 ( .A(n3168), .B(n1609), .Z(n3695) );
  AND U6768 ( .A(n3697), .B(n3698), .Z(n3693) );
  OR U6769 ( .A(n3172), .B(n1669), .Z(n3698) );
  OR U6770 ( .A(n3174), .B(n1695), .Z(n3697) );
  AND U6771 ( .A(n3699), .B(n3669), .Z(n3684) );
  NAND U6772 ( .A(n3158), .B(n1416), .Z(n3669) );
  NAND U6773 ( .A(n3700), .B(n3701), .Z(n1416) );
  AND U6774 ( .A(n3702), .B(n3703), .Z(n3701) );
  OR U6775 ( .A(n3166), .B(n1749), .Z(n3703) );
  OR U6776 ( .A(n3168), .B(n1721), .Z(n3702) );
  AND U6777 ( .A(n3704), .B(n3705), .Z(n3700) );
  OR U6778 ( .A(n3172), .B(n1775), .Z(n3705) );
  OR U6779 ( .A(n3174), .B(n1798), .Z(n3704) );
  NAND U6780 ( .A(n1414), .B(n3159), .Z(n3699) );
  AND U6781 ( .A(a_bus[3]), .B(a_bus[2]), .Z(n3159) );
  NAND U6782 ( .A(n3706), .B(n3707), .Z(n1414) );
  OR U6783 ( .A(n3168), .B(n1810), .Z(n3707) );
  OR U6784 ( .A(n3166), .B(n1824), .Z(n3706) );
  NAND U6785 ( .A(n3536), .B(n1134), .Z(n3662) );
  NAND U6786 ( .A(n3708), .B(n3709), .Z(n3536) );
  AND U6787 ( .A(n3710), .B(n3711), .Z(n3709) );
  OR U6788 ( .A(n3166), .B(n3489), .Z(n3711) );
  OR U6789 ( .A(n3168), .B(n3425), .Z(n3710) );
  AND U6790 ( .A(n3712), .B(n3713), .Z(n3708) );
  OR U6791 ( .A(n3172), .B(n1152), .Z(n3713) );
  OR U6792 ( .A(n3174), .B(n1192), .Z(n3712) );
  AND U6793 ( .A(n3670), .B(n3714), .Z(n3674) );
  NAND U6794 ( .A(n3672), .B(n1129), .Z(n3714) );
  NAND U6795 ( .A(n3715), .B(n3716), .Z(n3672) );
  AND U6796 ( .A(n3717), .B(n3718), .Z(n3716) );
  OR U6797 ( .A(n3166), .B(n3175), .Z(n3718) );
  OR U6798 ( .A(n3168), .B(n3173), .Z(n3717) );
  AND U6799 ( .A(n3719), .B(n3720), .Z(n3715) );
  OR U6800 ( .A(n3172), .B(n3488), .Z(n3720) );
  OR U6801 ( .A(n3174), .B(n3375), .Z(n3719) );
  NAND U6802 ( .A(n1261), .B(n1124), .Z(n3670) );
  NAND U6803 ( .A(n3721), .B(n3722), .Z(n1261) );
  AND U6804 ( .A(n3723), .B(n3724), .Z(n3722) );
  OR U6805 ( .A(n3166), .B(n1428), .Z(n3724) );
  OR U6806 ( .A(n3168), .B(n1390), .Z(n3723) );
  AND U6807 ( .A(n3725), .B(n3726), .Z(n3721) );
  OR U6808 ( .A(n3172), .B(n1460), .Z(n3726) );
  OR U6809 ( .A(n3174), .B(n1484), .Z(n3725) );
  AND U6810 ( .A(n3727), .B(n3728), .Z(n3653) );
  NAND U6811 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][2] ), .Z(n3728) );
  AND U6812 ( .A(\Shifter/sll_27/ML_int[3][2] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][2] ) );
  AND U6813 ( .A(\Shifter/sll_27/ML_int[2][2] ), .B(n3130), .Z(
        \Shifter/sll_27/ML_int[3][2] ) );
  NAND U6814 ( .A(n3729), .B(n1140), .Z(n3727) );
  XOR U6815 ( .A(n3730), .B(a_bus[2]), .Z(n3729) );
  AND U6816 ( .A(n3731), .B(n3732), .Z(n3651) );
  MUX U6817 ( .IN0(n1145), .IN1(n1146), .SEL(n3733), .F(n3732) );
  ANDN U6818 ( .A(n3175), .B(a_bus[2]), .Z(n3733) );
  AND U6819 ( .A(n3734), .B(n3735), .Z(n3731) );
  NAND U6820 ( .A(n3736), .B(n1151), .Z(n3735) );
  XNOR U6821 ( .A(n3130), .B(b_bus[2]), .Z(n3736) );
  NAND U6822 ( .A(n3737), .B(n1154), .Z(n3734) );
  ANDN U6823 ( .A(b_bus[2]), .B(n3130), .Z(n3737) );
  IV U6824 ( .A(n3175), .Z(b_bus[2]) );
  IV U6825 ( .A(n574), .Z(N28) );
  AND U6826 ( .A(n3738), .B(n3739), .Z(n574) );
  AND U6827 ( .A(n3740), .B(n3741), .Z(n3739) );
  AND U6828 ( .A(n3742), .B(n3743), .Z(n3741) );
  NAND U6829 ( .A(n3744), .B(n1109), .Z(n3743) );
  ANDN U6830 ( .A(n3745), .B(n3746), .Z(n1109) );
  NAND U6831 ( .A(n3747), .B(n3748), .Z(n3744) );
  AND U6832 ( .A(n3749), .B(n3750), .Z(n3748) );
  AND U6833 ( .A(n3751), .B(n3752), .Z(n3749) );
  OR U6834 ( .A(n1495), .B(n1117), .Z(n3752) );
  AND U6835 ( .A(n3753), .B(n3754), .Z(n1495) );
  AND U6836 ( .A(n3448), .B(n3755), .Z(n3754) );
  NAND U6837 ( .A(n1216), .B(n1650), .Z(n3755) );
  NAND U6838 ( .A(a_bus[2]), .B(n1652), .Z(n3448) );
  AND U6839 ( .A(\Shifter/N75 ), .B(a_bus[3]), .Z(n1652) );
  IV U6840 ( .A(n1810), .Z(\Shifter/N75 ) );
  AND U6841 ( .A(n3756), .B(n3757), .Z(n3753) );
  NAND U6842 ( .A(n3158), .B(n1369), .Z(n3756) );
  NAND U6843 ( .A(n3758), .B(n3759), .Z(n1369) );
  AND U6844 ( .A(n3130), .B(a_bus[3]), .Z(n3158) );
  AND U6845 ( .A(n3760), .B(n3761), .Z(n3747) );
  NAND U6846 ( .A(n3762), .B(n1118), .Z(n3761) );
  AND U6847 ( .A(n1650), .B(n1117), .Z(n1118) );
  ANDN U6848 ( .A(n3130), .B(a_bus[3]), .Z(n1650) );
  NAND U6849 ( .A(n3763), .B(n1121), .Z(n3742) );
  NOR U6850 ( .A(n3745), .B(n3746), .Z(n1121) );
  NAND U6851 ( .A(n3764), .B(n3765), .Z(n3763) );
  AND U6852 ( .A(n3766), .B(n3750), .Z(n3765) );
  NAND U6853 ( .A(n1132), .B(n1209), .Z(n3750) );
  NAND U6854 ( .A(n3767), .B(n3768), .Z(n1209) );
  AND U6855 ( .A(n3769), .B(n3770), .Z(n3768) );
  OR U6856 ( .A(n3166), .B(n1234), .Z(n3770) );
  AND U6857 ( .A(n3771), .B(n3772), .Z(n1234) );
  NAND U6858 ( .A(n3773), .B(imm[11]), .Z(n3772) );
  NAND U6859 ( .A(n3774), .B(reg_target[11]), .Z(n3771) );
  OR U6860 ( .A(n3168), .B(n1351), .Z(n3769) );
  AND U6861 ( .A(n3775), .B(n3776), .Z(n1351) );
  NAND U6862 ( .A(n3773), .B(imm[12]), .Z(n3776) );
  NAND U6863 ( .A(n3774), .B(reg_target[12]), .Z(n3775) );
  AND U6864 ( .A(n3777), .B(n3778), .Z(n3767) );
  OR U6865 ( .A(n3172), .B(n1428), .Z(n3778) );
  AND U6866 ( .A(n3779), .B(n3780), .Z(n1428) );
  NAND U6867 ( .A(n3773), .B(imm[14]), .Z(n3780) );
  NAND U6868 ( .A(n3774), .B(reg_target[14]), .Z(n3779) );
  OR U6869 ( .A(n3174), .B(n1314), .Z(n3777) );
  AND U6870 ( .A(n3781), .B(n3782), .Z(n1314) );
  NAND U6871 ( .A(n3773), .B(imm[13]), .Z(n3782) );
  NAND U6872 ( .A(n3774), .B(reg_target[13]), .Z(n3781) );
  ANDN U6873 ( .A(n3783), .B(a_bus[2]), .Z(n1132) );
  AND U6874 ( .A(n3751), .B(n3784), .Z(n3766) );
  OR U6875 ( .A(n1497), .B(n1117), .Z(n3784) );
  AND U6876 ( .A(n3785), .B(n3786), .Z(n1497) );
  NANDN U6877 ( .B(n3129), .A(n3787), .Z(n3786) );
  IV U6878 ( .A(n1220), .Z(n3787) );
  MUX U6879 ( .IN0(n1377), .IN1(n1378), .SEL(n3130), .F(n1220) );
  AND U6880 ( .A(n3758), .B(n3759), .Z(n1378) );
  AND U6881 ( .A(n3788), .B(n3789), .Z(n3759) );
  OR U6882 ( .A(n3166), .B(n1721), .Z(n3789) );
  ANDN U6883 ( .A(n3790), .B(n3189), .Z(n1721) );
  NAND U6884 ( .A(n3774), .B(reg_target[27]), .Z(n3790) );
  OR U6885 ( .A(n3168), .B(n1798), .Z(n3788) );
  ANDN U6886 ( .A(n3791), .B(n3189), .Z(n1798) );
  NAND U6887 ( .A(n3774), .B(reg_target[28]), .Z(n3791) );
  AND U6888 ( .A(n3792), .B(n3793), .Z(n3758) );
  OR U6889 ( .A(n3172), .B(n1824), .Z(n3793) );
  ANDN U6890 ( .A(n3794), .B(n3189), .Z(n1824) );
  NAND U6891 ( .A(n3774), .B(reg_target[30]), .Z(n3794) );
  OR U6892 ( .A(n3174), .B(n1775), .Z(n3792) );
  ANDN U6893 ( .A(n3795), .B(n3189), .Z(n1775) );
  NAND U6894 ( .A(n3774), .B(reg_target[29]), .Z(n3795) );
  OR U6895 ( .A(n3166), .B(n1810), .Z(n1377) );
  ANDN U6896 ( .A(n3796), .B(n3190), .Z(n1810) );
  AND U6897 ( .A(n3774), .B(reg_target[31]), .Z(n3190) );
  AND U6898 ( .A(n3757), .B(n3797), .Z(n3785) );
  NAND U6899 ( .A(n1415), .B(n1216), .Z(n3797) );
  NAND U6900 ( .A(n3798), .B(n3799), .Z(n1216) );
  AND U6901 ( .A(n3800), .B(n3801), .Z(n3799) );
  OR U6902 ( .A(n3166), .B(n1509), .Z(n3801) );
  ANDN U6903 ( .A(n3802), .B(n3189), .Z(n1509) );
  NAND U6904 ( .A(n3774), .B(reg_target[19]), .Z(n3802) );
  OR U6905 ( .A(n3168), .B(n1584), .Z(n3800) );
  ANDN U6906 ( .A(n3803), .B(n3189), .Z(n1584) );
  NAND U6907 ( .A(n3774), .B(reg_target[20]), .Z(n3803) );
  AND U6908 ( .A(n3804), .B(n3805), .Z(n3798) );
  OR U6909 ( .A(n3172), .B(n1633), .Z(n3805) );
  ANDN U6910 ( .A(n3806), .B(n3189), .Z(n1633) );
  NAND U6911 ( .A(n3774), .B(reg_target[22]), .Z(n3806) );
  OR U6912 ( .A(n3174), .B(n1560), .Z(n3804) );
  ANDN U6913 ( .A(n3807), .B(n3189), .Z(n1560) );
  NAND U6914 ( .A(n3774), .B(reg_target[21]), .Z(n3807) );
  NAND U6915 ( .A(n1222), .B(n1653), .Z(n3757) );
  NAND U6916 ( .A(n3808), .B(n3809), .Z(n1222) );
  AND U6917 ( .A(n3810), .B(n3811), .Z(n3809) );
  OR U6918 ( .A(n3166), .B(n1609), .Z(n3811) );
  ANDN U6919 ( .A(n3812), .B(n3189), .Z(n1609) );
  NAND U6920 ( .A(n3774), .B(reg_target[23]), .Z(n3812) );
  OR U6921 ( .A(n3168), .B(n1695), .Z(n3810) );
  ANDN U6922 ( .A(n3813), .B(n3189), .Z(n1695) );
  NAND U6923 ( .A(n3774), .B(reg_target[24]), .Z(n3813) );
  AND U6924 ( .A(n3814), .B(n3815), .Z(n3808) );
  OR U6925 ( .A(n3172), .B(n1749), .Z(n3815) );
  ANDN U6926 ( .A(n3816), .B(n3189), .Z(n1749) );
  NAND U6927 ( .A(n3774), .B(reg_target[26]), .Z(n3816) );
  OR U6928 ( .A(n3174), .B(n1669), .Z(n3814) );
  ANDN U6929 ( .A(n3817), .B(n3189), .Z(n1669) );
  NAND U6930 ( .A(n3774), .B(reg_target[25]), .Z(n3817) );
  NANDN U6931 ( .B(n3403), .A(n1134), .Z(n3751) );
  AND U6932 ( .A(n1653), .B(n1117), .Z(n1134) );
  ANDN U6933 ( .A(a_bus[2]), .B(a_bus[3]), .Z(n1653) );
  AND U6934 ( .A(n3818), .B(n3819), .Z(n3403) );
  AND U6935 ( .A(n3820), .B(n3821), .Z(n3819) );
  OR U6936 ( .A(n3166), .B(n3425), .Z(n3821) );
  AND U6937 ( .A(n3822), .B(n3823), .Z(n3425) );
  NAND U6938 ( .A(n3773), .B(imm[7]), .Z(n3823) );
  NAND U6939 ( .A(n3774), .B(reg_target[7]), .Z(n3822) );
  OR U6940 ( .A(n3168), .B(n1192), .Z(n3820) );
  AND U6941 ( .A(n3824), .B(n3825), .Z(n1192) );
  NAND U6942 ( .A(n3773), .B(imm[8]), .Z(n3825) );
  NAND U6943 ( .A(n3774), .B(reg_target[8]), .Z(n3824) );
  AND U6944 ( .A(n3826), .B(n3827), .Z(n3818) );
  OR U6945 ( .A(n3172), .B(n1273), .Z(n3827) );
  AND U6946 ( .A(n3828), .B(n3829), .Z(n1273) );
  NAND U6947 ( .A(n3773), .B(imm[10]), .Z(n3829) );
  NAND U6948 ( .A(n3774), .B(reg_target[10]), .Z(n3828) );
  OR U6949 ( .A(n3174), .B(n1152), .Z(n3826) );
  AND U6950 ( .A(n3830), .B(n3831), .Z(n1152) );
  NAND U6951 ( .A(n3773), .B(imm[9]), .Z(n3831) );
  NAND U6952 ( .A(n3774), .B(reg_target[9]), .Z(n3830) );
  AND U6953 ( .A(n3760), .B(n3832), .Z(n3764) );
  NAND U6954 ( .A(n3762), .B(n1129), .Z(n3832) );
  AND U6955 ( .A(n1415), .B(n1117), .Z(n1129) );
  ANDN U6956 ( .A(n3129), .B(a_bus[2]), .Z(n1415) );
  NAND U6957 ( .A(n3833), .B(n3834), .Z(n3762) );
  AND U6958 ( .A(n3835), .B(n3836), .Z(n3834) );
  OR U6959 ( .A(n3166), .B(n3173), .Z(n3836) );
  OR U6960 ( .A(n3168), .B(n3375), .Z(n3835) );
  AND U6961 ( .A(n3837), .B(n3838), .Z(n3375) );
  NANDN U6962 ( .B(n341), .A(n3773), .Z(n3838) );
  NAND U6963 ( .A(n3774), .B(reg_target[4]), .Z(n3837) );
  AND U6964 ( .A(n3839), .B(n3840), .Z(n3833) );
  OR U6965 ( .A(n3172), .B(n3489), .Z(n3840) );
  AND U6966 ( .A(n3841), .B(n3842), .Z(n3489) );
  NAND U6967 ( .A(n3773), .B(imm[6]), .Z(n3842) );
  NAND U6968 ( .A(n3774), .B(reg_target[6]), .Z(n3841) );
  OR U6969 ( .A(n3174), .B(n3488), .Z(n3839) );
  AND U6970 ( .A(n3843), .B(n3844), .Z(n3488) );
  NAND U6971 ( .A(n3773), .B(imm[5]), .Z(n3844) );
  NAND U6972 ( .A(n3774), .B(reg_target[5]), .Z(n3843) );
  NAND U6973 ( .A(n1124), .B(n1218), .Z(n3760) );
  NAND U6974 ( .A(n3845), .B(n3846), .Z(n1218) );
  AND U6975 ( .A(n3847), .B(n3848), .Z(n3846) );
  OR U6976 ( .A(n3166), .B(n1390), .Z(n3848) );
  AND U6977 ( .A(n3849), .B(n3850), .Z(n1390) );
  NAND U6978 ( .A(n3773), .B(imm[15]), .Z(n3850) );
  NAND U6979 ( .A(n3774), .B(reg_target[15]), .Z(n3849) );
  NANDN U6980 ( .B(a_bus[1]), .A(n3132), .Z(n3166) );
  OR U6981 ( .A(n3168), .B(n1484), .Z(n3847) );
  ANDN U6982 ( .A(n3851), .B(n3189), .Z(n1484) );
  NAND U6983 ( .A(n3774), .B(reg_target[16]), .Z(n3851) );
  NANDN U6984 ( .B(a_bus[1]), .A(a_bus[0]), .Z(n3168) );
  AND U6985 ( .A(n3852), .B(n3853), .Z(n3845) );
  OR U6986 ( .A(n3172), .B(n1533), .Z(n3853) );
  ANDN U6987 ( .A(n3854), .B(n3189), .Z(n1533) );
  IV U6988 ( .A(n3796), .Z(n3189) );
  NANDN U6989 ( .B(n3855), .A(imm[15]), .Z(n3796) );
  NAND U6990 ( .A(n3774), .B(reg_target[18]), .Z(n3854) );
  NANDN U6991 ( .B(n3131), .A(a_bus[0]), .Z(n3172) );
  OR U6992 ( .A(n3174), .B(n1460), .Z(n3852) );
  AND U6993 ( .A(n3856), .B(n3857), .Z(n1460) );
  NANDN U6994 ( .B(n3858), .A(imm[15]), .Z(n3857) );
  NAND U6995 ( .A(n3774), .B(reg_target[17]), .Z(n3856) );
  NANDN U6996 ( .B(a_bus[0]), .A(a_bus[1]), .Z(n3174) );
  AND U6997 ( .A(n3783), .B(a_bus[2]), .Z(n1124) );
  AND U6998 ( .A(n1117), .B(a_bus[3]), .Z(n3783) );
  IV U6999 ( .A(a_bus[4]), .Z(n1117) );
  AND U7000 ( .A(n3859), .B(n3860), .Z(n3740) );
  NAND U7001 ( .A(n1138), .B(\Shifter/sll_27/ML_int[4][3] ), .Z(n3860) );
  AND U7002 ( .A(\Shifter/sll_27/ML_int[3][3] ), .B(n3129), .Z(
        \Shifter/sll_27/ML_int[4][3] ) );
  AND U7003 ( .A(\Shifter/sll_27/ML_int[2][3] ), .B(n3130), .Z(
        \Shifter/sll_27/ML_int[3][3] ) );
  NOR U7004 ( .A(a_bus[4]), .B(n1450), .Z(n1138) );
  NAND U7005 ( .A(n3746), .B(n3745), .Z(n1450) );
  AND U7006 ( .A(n3861), .B(n3862), .Z(n3745) );
  ANDN U7007 ( .A(n3863), .B(n6), .Z(n3861) );
  NANDN U7008 ( .B(n752), .A(n3864), .Z(n3863) );
  NANDN U7009 ( .B(n14), .A(imm[0]), .Z(n3864) );
  AND U7010 ( .A(n14), .B(n376), .Z(n752) );
  NANDN U7011 ( .B(n3865), .A(n3862), .Z(n3746) );
  MUX U7012 ( .IN0(reg_source[4]), .IN1(imm[10]), .SEL(n3192), .F(a_bus[4]) );
  NAND U7013 ( .A(n3866), .B(n1140), .Z(n3859) );
  NANDN U7014 ( .B(n3867), .A(n3868), .Z(n1140) );
  OR U7015 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U7016 ( .A(n3576), .B(a_bus[3]), .Z(n3866) );
  XNOR U7017 ( .A(n3871), .B(n3578), .Z(n3576) );
  IV U7018 ( .A(n3574), .Z(n3578) );
  XOR U7019 ( .A(n3872), .B(n3873), .Z(n3574) );
  AND U7020 ( .A(n3730), .B(n3874), .Z(n3873) );
  XNOR U7021 ( .A(n3875), .B(n3130), .Z(n3874) );
  IV U7022 ( .A(a_bus[2]), .Z(n3130) );
  MUX U7023 ( .IN0(reg_source[2]), .IN1(imm[8]), .SEL(n3192), .F(a_bus[2]) );
  XNOR U7024 ( .A(n3876), .B(n3875), .Z(n3730) );
  IV U7025 ( .A(n3872), .Z(n3875) );
  XNOR U7026 ( .A(n3199), .B(n3175), .Z(n3876) );
  AND U7027 ( .A(n3877), .B(n3878), .Z(n3175) );
  NANDN U7028 ( .B(n359), .A(n3773), .Z(n3878) );
  NAND U7029 ( .A(n3774), .B(reg_target[2]), .Z(n3877) );
  XOR U7030 ( .A(n3879), .B(n3880), .Z(n3872) );
  AND U7031 ( .A(n3379), .B(n3881), .Z(n3880) );
  XNOR U7032 ( .A(n3882), .B(n3131), .Z(n3881) );
  IV U7033 ( .A(a_bus[1]), .Z(n3131) );
  MUX U7034 ( .IN0(reg_source[1]), .IN1(imm[7]), .SEL(n3192), .F(a_bus[1]) );
  XNOR U7035 ( .A(n3883), .B(n3882), .Z(n3379) );
  IV U7036 ( .A(n3879), .Z(n3882) );
  XNOR U7037 ( .A(n3199), .B(n3169), .Z(n3883) );
  AND U7038 ( .A(n3884), .B(n3885), .Z(n3169) );
  NANDN U7039 ( .B(n14), .A(n3773), .Z(n3885) );
  NAND U7040 ( .A(n3774), .B(reg_target[1]), .Z(n3884) );
  XOR U7041 ( .A(n3199), .B(n3886), .Z(n3879) );
  ANDN U7042 ( .A(n3887), .B(n3167), .Z(n3886) );
  AND U7043 ( .A(n3888), .B(n3889), .Z(n3167) );
  NANDN U7044 ( .B(n376), .A(n3773), .Z(n3889) );
  NAND U7045 ( .A(reg_target[0]), .B(n3774), .Z(n3888) );
  XOR U7046 ( .A(n3132), .B(n3199), .Z(n3887) );
  IV U7047 ( .A(a_bus[0]), .Z(n3132) );
  MUX U7048 ( .IN0(reg_source[0]), .IN1(imm[6]), .SEL(n3192), .F(a_bus[0]) );
  XNOR U7049 ( .A(n3199), .B(n3173), .Z(n3871) );
  ANDN U7050 ( .A(n3890), .B(n3179), .Z(n3199) );
  ANDN U7051 ( .A(n3891), .B(n3892), .Z(n3179) );
  NOR U7052 ( .A(n3185), .B(n3867), .Z(n3890) );
  ANDN U7053 ( .A(n3891), .B(n3893), .Z(n3867) );
  ANDN U7054 ( .A(n3894), .B(n3895), .Z(n3185) );
  ANDN U7055 ( .A(n3896), .B(n3891), .Z(n3894) );
  AND U7056 ( .A(n3897), .B(n3898), .Z(n3738) );
  MUX U7057 ( .IN0(n1145), .IN1(n1146), .SEL(n3899), .F(n3898) );
  ANDN U7058 ( .A(n3173), .B(a_bus[3]), .Z(n3899) );
  NAND U7059 ( .A(n3900), .B(n3901), .Z(n1146) );
  ANDN U7060 ( .A(n3902), .B(n376), .Z(n3901) );
  ANDN U7061 ( .A(n143), .B(n359), .Z(n3902) );
  NOR U7062 ( .A(n3865), .B(n647), .Z(n3900) );
  NANDN U7063 ( .B(n14), .A(n1831), .Z(n3865) );
  NANDN U7064 ( .B(n3869), .A(n3870), .Z(n1145) );
  NANDN U7065 ( .B(n3903), .A(n3896), .Z(n3869) );
  AND U7066 ( .A(n3904), .B(n3905), .Z(n3897) );
  NAND U7067 ( .A(n3906), .B(n1151), .Z(n3905) );
  ANDN U7068 ( .A(n3870), .B(n3892), .Z(n1151) );
  NANDN U7069 ( .B(n3896), .A(n3895), .Z(n3892) );
  IV U7070 ( .A(n3903), .Z(n3895) );
  XNOR U7071 ( .A(n3129), .B(b_bus[3]), .Z(n3906) );
  NAND U7072 ( .A(n3907), .B(n1154), .Z(n3904) );
  ANDN U7073 ( .A(n3870), .B(n3893), .Z(n1154) );
  NANDN U7074 ( .B(n3896), .A(n3903), .Z(n3893) );
  AND U7075 ( .A(n3908), .B(n3909), .Z(n3903) );
  AND U7076 ( .A(n3910), .B(n3911), .Z(n3909) );
  ANDN U7077 ( .A(n3912), .B(n3913), .Z(n3911) );
  AND U7078 ( .A(n3914), .B(n3915), .Z(n3908) );
  NANDN U7079 ( .B(n6), .A(n3916), .Z(n3915) );
  NAND U7080 ( .A(n3917), .B(n1827), .Z(n3916) );
  AND U7081 ( .A(n1828), .B(n3918), .Z(n3917) );
  NANDN U7082 ( .B(n10), .A(n3919), .Z(n3918) );
  NAND U7083 ( .A(n3920), .B(n3921), .Z(n3919) );
  ANDN U7084 ( .A(n3922), .B(n1833), .Z(n3920) );
  NANDN U7085 ( .B(n647), .A(n3923), .Z(n3922) );
  NANDN U7086 ( .B(n3924), .A(n3925), .Z(n3923) );
  NANDN U7087 ( .B(imm[1]), .A(n359), .Z(n3925) );
  MUX U7088 ( .IN0(n14), .IN1(n3926), .SEL(n376), .F(n3924) );
  ANDN U7089 ( .A(imm[1]), .B(n359), .Z(n3926) );
  NANDN U7090 ( .B(n633), .A(n3927), .Z(n3914) );
  NAND U7091 ( .A(n3928), .B(n3929), .Z(n3927) );
  ANDN U7092 ( .A(n10), .B(n43), .Z(n3929) );
  ANDN U7093 ( .A(n3930), .B(n3931), .Z(n3928) );
  AND U7094 ( .A(n3932), .B(n3933), .Z(n3896) );
  NANDN U7095 ( .B(n633), .A(n3934), .Z(n3933) );
  OR U7096 ( .A(n1085), .B(n791), .Z(n3934) );
  NANDN U7097 ( .B(n6), .A(n3935), .Z(n3932) );
  NAND U7098 ( .A(n3936), .B(n96), .Z(n3935) );
  NANDN U7099 ( .B(n10), .A(n3937), .Z(n3936) );
  NAND U7100 ( .A(n3938), .B(n3921), .Z(n3937) );
  NANDN U7101 ( .B(n651), .A(n756), .Z(n3921) );
  ANDN U7102 ( .A(n3939), .B(n376), .Z(n756) );
  ANDN U7103 ( .A(n359), .B(n14), .Z(n3939) );
  NANDN U7104 ( .B(n647), .A(n3940), .Z(n3938) );
  NANDN U7105 ( .B(n3941), .A(n3942), .Z(n3940) );
  IV U7106 ( .A(n3891), .Z(n3870) );
  AND U7107 ( .A(n3943), .B(n3944), .Z(n3891) );
  NANDN U7108 ( .B(n6), .A(n3945), .Z(n3944) );
  NAND U7109 ( .A(n3946), .B(n1827), .Z(n3945) );
  AND U7110 ( .A(n3947), .B(n3948), .Z(n1827) );
  ANDN U7111 ( .A(n3334), .B(n130), .Z(n3947) );
  ANDN U7112 ( .A(n3949), .B(n3950), .Z(n130) );
  ANDN U7113 ( .A(opcode[26]), .B(n3951), .Z(n3949) );
  AND U7114 ( .A(n1828), .B(n3952), .Z(n3946) );
  NANDN U7115 ( .B(n10), .A(n3953), .Z(n3952) );
  NANDN U7116 ( .B(n1833), .A(n3954), .Z(n3953) );
  AND U7117 ( .A(n3955), .B(n3956), .Z(n3954) );
  NANDN U7118 ( .B(n647), .A(n3957), .Z(n3956) );
  NANDN U7119 ( .B(n114), .A(n3942), .Z(n3957) );
  NAND U7120 ( .A(n376), .B(imm[2]), .Z(n3942) );
  NAND U7121 ( .A(n3958), .B(imm[5]), .Z(n647) );
  ANDN U7122 ( .A(n350), .B(imm[4]), .Z(n3958) );
  NANDN U7123 ( .B(n651), .A(n745), .Z(n3955) );
  ANDN U7124 ( .A(n3959), .B(n14), .Z(n745) );
  ANDN U7125 ( .A(n376), .B(imm[2]), .Z(n3959) );
  NAND U7126 ( .A(n3960), .B(imm[5]), .Z(n651) );
  ANDN U7127 ( .A(n341), .B(n350), .Z(n3960) );
  AND U7128 ( .A(n3961), .B(n113), .Z(n1833) );
  AND U7129 ( .A(n3962), .B(imm[3]), .Z(n113) );
  NANDN U7130 ( .B(n797), .A(n3963), .Z(n3961) );
  ANDN U7131 ( .A(n656), .B(n114), .Z(n3963) );
  AND U7132 ( .A(n14), .B(imm[2]), .Z(n114) );
  OR U7133 ( .A(n747), .B(n376), .Z(n656) );
  IV U7134 ( .A(imm[0]), .Z(n376) );
  NOR U7135 ( .A(imm[0]), .B(n747), .Z(n797) );
  NANDN U7136 ( .B(imm[2]), .A(n14), .Z(n747) );
  IV U7137 ( .A(imm[1]), .Z(n14) );
  NANDN U7138 ( .B(n805), .A(n3964), .Z(n1828) );
  ANDN U7139 ( .A(n23), .B(n18), .Z(n3964) );
  IV U7140 ( .A(opcode[19]), .Z(n23) );
  NANDN U7141 ( .B(opcode[17]), .A(n49), .Z(n805) );
  IV U7142 ( .A(opcode[18]), .Z(n49) );
  AND U7143 ( .A(n3910), .B(n3965), .Z(n3943) );
  NANDN U7144 ( .B(n633), .A(n3966), .Z(n3965) );
  NANDN U7145 ( .B(n3931), .A(n793), .Z(n3966) );
  AND U7146 ( .A(n3334), .B(n3335), .Z(n793) );
  IV U7147 ( .A(n1077), .Z(n3335) );
  NAND U7148 ( .A(n3967), .B(n3968), .Z(n3910) );
  ANDN U7149 ( .A(n127), .B(n10), .Z(n3968) );
  ANDN U7150 ( .A(n908), .B(opcode[21]), .Z(n127) );
  IV U7151 ( .A(opcode[22]), .Z(n908) );
  ANDN U7152 ( .A(n26), .B(n126), .Z(n3967) );
  NANDN U7153 ( .B(opcode[24]), .A(n886), .Z(n126) );
  IV U7154 ( .A(opcode[25]), .Z(n886) );
  AND U7155 ( .A(n3969), .B(opcode[30]), .Z(n26) );
  ANDN U7156 ( .A(n3970), .B(opcode[29]), .Z(n3969) );
  ANDN U7157 ( .A(b_bus[3]), .B(n3129), .Z(n3907) );
  IV U7158 ( .A(a_bus[3]), .Z(n3129) );
  MUX U7159 ( .IN0(reg_source[3]), .IN1(imm[9]), .SEL(n3192), .F(a_bus[3]) );
  AND U7160 ( .A(n3971), .B(n3862), .Z(n3192) );
  AND U7161 ( .A(n751), .B(n143), .Z(n3862) );
  ANDN U7162 ( .A(n3962), .B(imm[3]), .Z(n751) );
  ANDN U7163 ( .A(n341), .B(imm[5]), .Z(n3962) );
  IV U7164 ( .A(imm[4]), .Z(n341) );
  ANDN U7165 ( .A(n3972), .B(n6), .Z(n3971) );
  IV U7166 ( .A(n1831), .Z(n6) );
  AND U7167 ( .A(n3973), .B(n133), .Z(n1831) );
  NANDN U7168 ( .B(n3941), .A(n3974), .Z(n3972) );
  NANDN U7169 ( .B(imm[0]), .A(n359), .Z(n3974) );
  AND U7170 ( .A(n359), .B(imm[1]), .Z(n3941) );
  IV U7171 ( .A(imm[2]), .Z(n359) );
  IV U7172 ( .A(n3173), .Z(b_bus[3]) );
  AND U7173 ( .A(n3975), .B(n3976), .Z(n3173) );
  NANDN U7174 ( .B(n350), .A(n3773), .Z(n3976) );
  NAND U7175 ( .A(n3977), .B(n3855), .Z(n3773) );
  NANDN U7176 ( .B(n3858), .A(n3978), .Z(n3855) );
  OR U7177 ( .A(n3978), .B(n3979), .Z(n3977) );
  IV U7178 ( .A(imm[3]), .Z(n350) );
  NAND U7179 ( .A(n3774), .B(reg_target[3]), .Z(n3975) );
  AND U7180 ( .A(n3978), .B(n3858), .Z(n3774) );
  IV U7181 ( .A(n3979), .Z(n3858) );
  NAND U7182 ( .A(n3980), .B(n3912), .Z(n3979) );
  NANDN U7183 ( .B(n660), .A(n662), .Z(n3912) );
  NANDN U7184 ( .B(n3981), .A(n128), .Z(n662) );
  NOR U7185 ( .A(n1832), .B(n3982), .Z(n128) );
  NANDN U7186 ( .B(n791), .A(n96), .Z(n3982) );
  ANDN U7187 ( .A(n3983), .B(n3913), .Z(n3980) );
  AND U7188 ( .A(n3984), .B(n3330), .Z(n3913) );
  NANDN U7189 ( .B(n633), .A(n3985), .Z(n3983) );
  OR U7190 ( .A(n3981), .B(n1077), .Z(n3985) );
  NANDN U7191 ( .B(n633), .A(n3986), .Z(n3978) );
  OR U7192 ( .A(n1085), .B(n3931), .Z(n3986) );
  IV U7193 ( .A(n3948), .Z(n3931) );
  ANDN U7194 ( .A(n3987), .B(n792), .Z(n3948) );
  IV U7195 ( .A(n791), .Z(n3987) );
  ANDN U7196 ( .A(n3988), .B(n3950), .Z(n791) );
  ANDN U7197 ( .A(n3989), .B(n3951), .Z(n3988) );
  NANDN U7198 ( .B(n671), .A(n3334), .Z(n1085) );
  NANDN U7199 ( .B(n133), .A(n3973), .Z(n633) );
  ANDN U7200 ( .A(n3970), .B(opcode[30]), .Z(n3973) );
  IV U7201 ( .A(opcode[31]), .Z(n3970) );
  AND U7202 ( .A(n809), .B(n3913), .Z(n1902) );
  NAND U7203 ( .A(n3984), .B(n3330), .Z(n3326) );
  OR U7204 ( .A(n3981), .B(n1832), .Z(n3984) );
  IV U7205 ( .A(n95), .Z(n1832) );
  ANDN U7206 ( .A(n3930), .B(n1077), .Z(n95) );
  ANDN U7207 ( .A(n3989), .B(n3990), .Z(n1077) );
  IV U7208 ( .A(n671), .Z(n3930) );
  NOR U7209 ( .A(n3989), .B(n3990), .Z(n671) );
  NANDN U7210 ( .B(n3951), .A(n3950), .Z(n3990) );
  IV U7211 ( .A(opcode[28]), .Z(n3950) );
  AND U7212 ( .A(n3991), .B(n3992), .Z(n809) );
  NANDN U7213 ( .B(n660), .A(n3993), .Z(n3992) );
  NANDN U7214 ( .B(n3981), .A(n96), .Z(n3993) );
  ANDN U7215 ( .A(n3334), .B(n792), .Z(n96) );
  NOR U7216 ( .A(n3989), .B(n3994), .Z(n792) );
  NANDN U7217 ( .B(n3994), .A(n3989), .Z(n3334) );
  NANDN U7218 ( .B(opcode[27]), .A(opcode[28]), .Z(n3994) );
  NANDN U7219 ( .B(n143), .A(n18), .Z(n3981) );
  IV U7220 ( .A(n134), .Z(n660) );
  AND U7221 ( .A(n3995), .B(n133), .Z(n134) );
  NANDN U7222 ( .B(n818), .A(n3330), .Z(n3991) );
  ANDN U7223 ( .A(n3995), .B(n133), .Z(n3330) );
  IV U7224 ( .A(opcode[29]), .Z(n133) );
  ANDN U7225 ( .A(opcode[31]), .B(opcode[30]), .Z(n3995) );
  AND U7226 ( .A(n18), .B(n10), .Z(n818) );
  IV U7227 ( .A(n143), .Z(n10) );
  ANDN U7228 ( .A(n3996), .B(opcode[26]), .Z(n143) );
  IV U7229 ( .A(n43), .Z(n18) );
  ANDN U7230 ( .A(n3996), .B(n3989), .Z(n43) );
  IV U7231 ( .A(opcode[26]), .Z(n3989) );
  ANDN U7232 ( .A(n3951), .B(opcode[28]), .Z(n3996) );
  IV U7233 ( .A(opcode[27]), .Z(n3951) );
endmodule

