module sum ( clk, rst, a, b, c );
input  [8191:0] a;
input  [8191:0] b;
output [8191:0] c;
input clk, rst;

wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
	n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, 
	n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
	n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
	n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, 
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
	n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
	n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
	n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
	n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
	n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
	n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
	n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
	n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
	n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
	n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
	n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
	n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
	n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
	n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
	n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
	n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
	n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
	n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
	n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
	n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
	n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
	n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, 
	n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
	n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
	n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
	n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
	n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
	n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, 
	n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
	n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
	n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
	n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
	n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
	n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
	n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
	n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
	n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, 
	n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
	n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
	n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, 
	n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
	n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
	n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
	n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
	n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, 
	n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, 
	n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
	n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
	n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
	n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
	n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, 
	n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, 
	n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
	n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
	n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
	n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
	n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
	n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, 
	n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
	n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
	n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
	n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
	n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
	n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, 
	n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
	n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
	n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
	n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
	n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
	n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
	n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
	n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
	n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, 
	n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
	n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
	n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, 
	n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, 
	n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
	n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
	n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
	n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, 
	n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, 
	n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
	n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
	n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
	n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
	n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, 
	n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, 
	n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
	n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
	n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
	n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
	n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
	n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
	n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
	n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
	n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
	n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
	n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
	n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
	n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
	n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
	n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
	n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
	n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
	n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
	n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
	n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
	n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
	n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
	n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
	n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
	n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
	n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
	n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
	n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
	n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
	n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
	n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
	n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
	n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
	n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
	n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
	n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
	n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
	n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
	n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
	n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
	n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
	n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
	n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
	n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
	n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
	n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
	n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
	n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
	n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
	n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
	n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
	n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
	n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
	n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
	n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
	n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
	n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
	n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
	n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
	n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
	n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
	n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
	n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
	n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
	n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
	n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
	n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
	n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
	n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
	n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
	n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
	n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
	n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
	n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
	n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
	n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
	n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
	n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
	n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
	n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
	n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
	n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, 
	n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, 
	n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
	n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
	n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
	n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
	n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
	n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
	n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
	n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
	n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
	n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
	n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
	n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
	n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
	n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
	n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
	n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
	n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
	n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
	n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
	n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
	n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
	n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
	n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
	n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
	n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
	n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
	n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
	n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
	n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
	n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
	n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
	n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
	n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
	n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
	n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
	n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
	n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
	n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
	n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, 
	n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, 
	n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
	n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
	n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, 
	n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, 
	n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, 
	n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, 
	n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, 
	n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, 
	n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, 
	n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, 
	n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, 
	n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, 
	n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, 
	n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, 
	n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, 
	n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, 
	n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
	n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
	n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
	n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, 
	n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
	n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
	n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
	n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, 
	n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, 
	n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
	n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
	n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, 
	n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, 
	n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, 
	n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
	n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, 
	n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, 
	n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, 
	n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
	n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, 
	n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, 
	n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, 
	n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, 
	n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, 
	n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, 
	n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
	n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, 
	n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, 
	n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, 
	n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, 
	n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, 
	n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, 
	n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
	n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
	n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, 
	n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, 
	n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
	n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, 
	n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, 
	n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, 
	n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, 
	n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, 
	n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, 
	n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, 
	n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, 
	n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, 
	n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, 
	n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, 
	n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
	n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
	n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, 
	n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, 
	n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, 
	n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, 
	n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, 
	n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, 
	n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, 
	n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
	n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
	n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
	n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, 
	n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, 
	n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, 
	n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, 
	n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, 
	n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, 
	n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, 
	n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, 
	n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, 
	n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, 
	n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, 
	n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
	n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, 
	n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, 
	n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, 
	n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, 
	n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, 
	n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, 
	n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, 
	n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, 
	n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, 
	n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, 
	n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, 
	n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, 
	n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, 
	n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
	n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, 
	n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, 
	n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, 
	n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, 
	n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, 
	n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, 
	n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, 
	n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, 
	n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, 
	n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, 
	n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, 
	n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, 
	n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, 
	n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, 
	n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, 
	n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, 
	n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, 
	n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, 
	n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, 
	n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, 
	n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, 
	n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, 
	n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, 
	n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, 
	n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, 
	n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
	n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, 
	n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, 
	n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, 
	n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, 
	n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, 
	n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
	n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, 
	n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, 
	n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, 
	n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, 
	n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, 
	n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, 
	n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, 
	n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, 
	n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, 
	n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, 
	n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, 
	n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, 
	n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, 
	n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, 
	n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, 
	n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, 
	n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
	n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, 
	n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, 
	n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, 
	n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, 
	n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, 
	n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, 
	n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, 
	n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, 
	n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, 
	n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, 
	n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, 
	n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
	n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
	n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, 
	n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, 
	n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, 
	n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, 
	n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, 
	n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, 
	n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, 
	n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, 
	n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, 
	n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
	n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, 
	n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, 
	n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, 
	n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, 
	n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, 
	n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, 
	n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, 
	n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, 
	n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, 
	n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, 
	n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, 
	n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, 
	n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, 
	n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, 
	n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, 
	n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, 
	n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, 
	n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, 
	n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, 
	n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, 
	n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, 
	n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, 
	n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, 
	n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, 
	n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, 
	n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, 
	n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, 
	n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, 
	n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, 
	n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, 
	n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, 
	n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, 
	n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, 
	n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, 
	n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, 
	n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, 
	n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, 
	n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, 
	n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, 
	n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, 
	n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, 
	n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, 
	n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, 
	n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, 
	n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, 
	n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, 
	n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, 
	n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, 
	n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, 
	n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, 
	n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, 
	n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, 
	n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, 
	n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, 
	n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, 
	n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, 
	n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, 
	n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, 
	n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, 
	n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, 
	n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, 
	n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, 
	n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, 
	n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, 
	n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, 
	n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, 
	n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, 
	n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, 
	n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, 
	n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, 
	n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, 
	n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, 
	n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, 
	n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, 
	n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, 
	n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, 
	n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, 
	n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, 
	n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, 
	n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, 
	n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, 
	n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
	n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, 
	n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, 
	n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, 
	n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, 
	n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, 
	n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, 
	n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, 
	n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, 
	n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, 
	n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, 
	n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, 
	n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, 
	n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, 
	n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, 
	n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, 
	n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
	n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, 
	n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, 
	n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, 
	n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, 
	n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, 
	n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, 
	n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, 
	n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, 
	n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, 
	n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, 
	n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, 
	n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, 
	n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, 
	n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, 
	n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, 
	n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, 
	n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, 
	n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, 
	n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, 
	n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
	n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, 
	n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, 
	n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, 
	n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, 
	n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, 
	n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, 
	n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, 
	n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
	n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, 
	n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
	n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, 
	n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
	n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, 
	n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
	n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
	n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
	n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
	n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
	n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
	n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
	n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
	n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
	n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
	n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
	n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
	n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
	n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
	n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
	n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, 
	n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, 
	n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, 
	n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
	n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, 
	n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
	n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
	n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
	n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
	n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
	n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
	n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
	n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, 
	n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, 
	n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
	n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, 
	n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
	n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, 
	n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, 
	n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, 
	n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, 
	n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, 
	n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, 
	n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, 
	n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, 
	n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, 
	n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, 
	n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
	n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, 
	n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, 
	n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, 
	n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, 
	n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, 
	n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, 
	n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, 
	n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
	n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, 
	n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, 
	n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, 
	n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
	n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, 
	n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, 
	n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, 
	n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, 
	n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, 
	n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, 
	n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, 
	n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, 
	n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
	n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
	n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
	n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
	n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
	n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
	n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, 
	n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, 
	n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, 
	n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, 
	n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, 
	n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, 
	n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, 
	n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, 
	n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, 
	n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
	n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, 
	n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
	n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, 
	n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
	n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, 
	n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, 
	n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, 
	n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
	n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, 
	n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, 
	n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, 
	n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, 
	n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, 
	n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, 
	n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, 
	n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, 
	n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, 
	n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, 
	n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, 
	n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, 
	n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, 
	n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, 
	n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, 
	n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, 
	n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
	n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, 
	n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, 
	n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, 
	n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, 
	n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, 
	n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, 
	n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, 
	n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, 
	n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, 
	n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, 
	n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, 
	n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, 
	n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, 
	n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, 
	n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, 
	n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, 
	n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, 
	n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, 
	n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, 
	n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, 
	n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, 
	n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, 
	n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, 
	n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, 
	n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, 
	n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, 
	n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, 
	n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, 
	n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, 
	n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, 
	n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, 
	n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, 
	n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, 
	n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, 
	n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, 
	n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, 
	n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, 
	n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, 
	n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, 
	n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, 
	n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, 
	n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, 
	n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, 
	n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, 
	n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, 
	n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, 
	n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, 
	n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, 
	n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, 
	n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, 
	n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, 
	n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, 
	n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, 
	n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, 
	n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, 
	n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, 
	n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, 
	n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, 
	n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, 
	n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, 
	n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, 
	n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, 
	n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, 
	n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, 
	n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, 
	n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
	n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
	n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, 
	n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
	n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, 
	n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
	n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, 
	n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, 
	n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, 
	n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
	n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, 
	n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, 
	n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, 
	n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, 
	n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, 
	n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, 
	n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, 
	n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, 
	n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, 
	n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, 
	n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, 
	n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, 
	n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, 
	n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, 
	n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, 
	n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, 
	n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, 
	n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, 
	n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, 
	n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, 
	n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, 
	n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, 
	n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, 
	n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, 
	n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, 
	n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, 
	n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, 
	n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, 
	n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, 
	n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, 
	n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, 
	n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, 
	n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, 
	n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, 
	n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, 
	n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, 
	n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, 
	n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, 
	n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, 
	n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, 
	n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, 
	n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, 
	n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, 
	n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, 
	n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, 
	n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, 
	n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, 
	n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, 
	n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, 
	n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, 
	n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, 
	n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, 
	n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, 
	n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, 
	n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, 
	n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, 
	n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, 
	n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, 
	n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, 
	n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, 
	n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, 
	n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, 
	n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, 
	n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, 
	n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, 
	n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, 
	n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, 
	n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, 
	n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, 
	n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, 
	n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, 
	n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, 
	n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, 
	n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, 
	n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, 
	n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, 
	n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, 
	n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, 
	n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, 
	n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, 
	n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, 
	n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, 
	n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, 
	n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, 
	n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, 
	n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, 
	n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, 
	n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, 
	n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, 
	n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, 
	n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, 
	n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, 
	n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, 
	n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, 
	n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, 
	n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, 
	n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, 
	n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, 
	n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, 
	n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, 
	n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, 
	n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, 
	n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, 
	n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, 
	n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, 
	n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, 
	n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, 
	n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, 
	n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, 
	n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, 
	n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, 
	n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, 
	n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, 
	n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, 
	n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, 
	n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, 
	n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, 
	n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, 
	n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, 
	n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, 
	n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, 
	n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, 
	n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, 
	n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, 
	n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, 
	n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, 
	n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, 
	n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, 
	n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, 
	n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, 
	n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, 
	n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, 
	n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, 
	n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, 
	n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, 
	n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, 
	n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, 
	n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, 
	n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, 
	n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, 
	n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, 
	n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, 
	n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, 
	n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, 
	n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, 
	n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, 
	n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, 
	n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, 
	n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, 
	n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, 
	n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, 
	n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, 
	n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, 
	n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, 
	n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, 
	n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, 
	n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, 
	n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, 
	n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, 
	n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, 
	n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, 
	n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, 
	n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, 
	n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, 
	n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, 
	n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, 
	n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, 
	n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, 
	n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, 
	n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, 
	n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, 
	n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, 
	n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, 
	n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, 
	n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, 
	n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, 
	n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, 
	n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, 
	n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, 
	n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, 
	n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, 
	n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, 
	n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, 
	n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, 
	n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, 
	n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, 
	n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, 
	n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, 
	n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, 
	n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, 
	n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, 
	n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, 
	n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, 
	n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, 
	n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, 
	n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, 
	n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, 
	n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, 
	n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, 
	n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, 
	n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, 
	n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, 
	n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, 
	n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, 
	n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, 
	n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, 
	n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, 
	n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, 
	n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, 
	n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, 
	n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, 
	n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, 
	n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, 
	n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, 
	n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, 
	n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, 
	n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, 
	n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, 
	n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, 
	n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, 
	n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, 
	n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, 
	n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, 
	n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, 
	n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, 
	n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, 
	n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, 
	n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, 
	n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, 
	n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, 
	n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, 
	n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, 
	n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, 
	n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, 
	n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, 
	n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, 
	n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, 
	n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, 
	n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, 
	n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, 
	n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, 
	n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, 
	n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, 
	n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, 
	n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, 
	n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, 
	n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, 
	n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, 
	n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, 
	n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, 
	n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, 
	n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, 
	n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, 
	n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, 
	n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, 
	n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, 
	n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, 
	n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, 
	n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, 
	n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, 
	n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, 
	n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, 
	n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, 
	n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, 
	n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, 
	n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, 
	n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, 
	n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, 
	n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, 
	n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, 
	n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, 
	n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, 
	n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, 
	n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, 
	n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, 
	n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, 
	n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, 
	n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, 
	n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, 
	n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, 
	n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, 
	n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, 
	n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, 
	n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, 
	n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, 
	n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, 
	n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, 
	n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, 
	n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, 
	n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, 
	n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, 
	n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, 
	n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, 
	n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, 
	n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, 
	n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, 
	n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, 
	n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, 
	n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, 
	n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, 
	n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, 
	n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, 
	n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, 
	n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
	n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, 
	n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, 
	n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, 
	n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, 
	n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, 
	n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, 
	n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, 
	n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, 
	n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
	n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, 
	n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, 
	n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, 
	n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
	n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, 
	n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, 
	n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, 
	n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, 
	n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, 
	n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, 
	n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, 
	n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, 
	n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, 
	n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, 
	n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
	n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, 
	n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, 
	n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
	n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, 
	n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, 
	n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, 
	n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, 
	n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, 
	n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, 
	n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
	n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, 
	n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
	n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, 
	n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, 
	n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, 
	n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, 
	n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, 
	n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, 
	n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, 
	n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, 
	n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, 
	n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, 
	n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, 
	n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, 
	n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, 
	n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, 
	n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, 
	n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, 
	n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, 
	n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, 
	n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, 
	n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, 
	n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
	n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, 
	n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, 
	n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, 
	n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, 
	n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, 
	n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, 
	n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, 
	n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, 
	n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, 
	n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, 
	n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, 
	n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, 
	n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, 
	n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, 
	n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, 
	n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, 
	n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, 
	n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, 
	n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, 
	n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, 
	n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, 
	n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, 
	n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, 
	n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, 
	n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, 
	n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, 
	n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, 
	n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, 
	n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, 
	n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, 
	n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, 
	n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, 
	n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
	n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, 
	n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, 
	n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, 
	n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
	n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, 
	n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, 
	n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, 
	n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, 
	n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, 
	n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, 
	n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, 
	n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, 
	n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, 
	n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, 
	n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, 
	n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, 
	n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, 
	n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, 
	n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, 
	n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, 
	n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, 
	n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, 
	n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, 
	n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, 
	n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, 
	n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, 
	n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, 
	n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, 
	n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, 
	n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, 
	n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, 
	n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, 
	n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, 
	n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, 
	n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, 
	n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, 
	n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, 
	n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, 
	n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, 
	n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, 
	n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, 
	n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, 
	n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, 
	n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, 
	n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, 
	n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, 
	n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, 
	n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, 
	n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, 
	n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, 
	n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, 
	n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, 
	n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, 
	n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, 
	n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, 
	n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, 
	n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, 
	n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
	n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, 
	n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, 
	n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, 
	n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, 
	n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
	n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, 
	n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, 
	n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, 
	n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, 
	n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, 
	n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, 
	n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, 
	n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, 
	n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, 
	n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, 
	n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, 
	n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, 
	n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
	n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, 
	n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, 
	n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, 
	n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, 
	n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, 
	n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, 
	n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, 
	n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, 
	n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, 
	n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, 
	n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, 
	n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, 
	n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, 
	n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, 
	n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, 
	n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, 
	n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, 
	n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, 
	n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, 
	n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, 
	n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, 
	n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, 
	n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, 
	n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, 
	n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, 
	n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, 
	n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, 
	n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, 
	n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, 
	n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, 
	n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, 
	n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
	n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, 
	n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, 
	n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, 
	n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, 
	n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, 
	n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, 
	n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, 
	n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, 
	n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, 
	n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, 
	n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, 
	n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, 
	n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, 
	n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, 
	n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, 
	n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, 
	n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, 
	n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, 
	n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, 
	n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, 
	n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, 
	n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, 
	n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, 
	n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, 
	n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, 
	n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, 
	n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, 
	n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, 
	n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, 
	n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, 
	n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, 
	n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, 
	n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, 
	n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, 
	n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, 
	n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, 
	n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, 
	n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, 
	n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, 
	n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, 
	n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
	n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, 
	n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, 
	n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, 
	n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, 
	n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, 
	n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, 
	n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, 
	n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, 
	n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, 
	n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, 
	n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, 
	n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, 
	n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, 
	n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, 
	n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, 
	n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, 
	n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, 
	n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, 
	n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, 
	n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, 
	n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, 
	n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, 
	n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, 
	n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, 
	n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, 
	n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, 
	n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, 
	n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, 
	n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, 
	n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, 
	n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, 
	n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, 
	n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, 
	n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, 
	n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, 
	n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, 
	n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, 
	n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, 
	n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, 
	n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, 
	n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, 
	n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, 
	n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, 
	n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, 
	n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, 
	n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, 
	n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, 
	n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, 
	n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, 
	n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, 
	n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, 
	n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, 
	n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, 
	n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, 
	n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, 
	n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, 
	n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, 
	n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, 
	n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, 
	n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, 
	n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, 
	n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, 
	n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, 
	n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, 
	n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, 
	n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, 
	n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, 
	n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, 
	n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, 
	n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, 
	n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, 
	n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, 
	n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, 
	n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, 
	n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, 
	n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, 
	n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, 
	n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, 
	n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, 
	n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, 
	n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, 
	n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, 
	n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, 
	n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, 
	n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, 
	n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, 
	n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, 
	n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, 
	n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, 
	n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, 
	n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, 
	n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, 
	n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, 
	n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, 
	n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, 
	n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, 
	n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, 
	n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, 
	n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, 
	n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, 
	n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, 
	n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, 
	n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, 
	n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, 
	n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, 
	n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, 
	n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, 
	n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, 
	n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, 
	n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, 
	n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, 
	n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, 
	n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, 
	n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, 
	n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, 
	n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, 
	n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, 
	n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, 
	n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, 
	n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, 
	n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, 
	n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, 
	n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, 
	n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, 
	n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, 
	n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, 
	n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, 
	n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, 
	n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, 
	n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, 
	n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, 
	n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, 
	n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, 
	n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, 
	n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, 
	n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, 
	n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, 
	n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, 
	n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, 
	n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, 
	n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, 
	n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, 
	n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, 
	n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, 
	n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, 
	n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, 
	n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, 
	n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, 
	n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, 
	n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, 
	n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
	n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, 
	n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, 
	n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, 
	n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, 
	n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, 
	n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, 
	n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, 
	n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, 
	n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, 
	n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, 
	n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, 
	n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, 
	n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, 
	n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, 
	n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, 
	n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, 
	n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, 
	n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, 
	n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, 
	n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, 
	n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, 
	n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, 
	n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
	n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, 
	n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, 
	n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, 
	n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, 
	n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, 
	n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, 
	n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, 
	n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, 
	n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, 
	n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, 
	n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, 
	n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, 
	n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, 
	n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, 
	n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, 
	n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, 
	n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, 
	n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, 
	n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, 
	n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, 
	n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, 
	n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, 
	n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, 
	n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, 
	n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, 
	n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, 
	n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, 
	n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, 
	n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, 
	n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, 
	n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, 
	n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, 
	n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, 
	n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, 
	n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, 
	n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, 
	n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, 
	n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, 
	n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, 
	n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, 
	n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, 
	n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, 
	n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, 
	n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, 
	n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, 
	n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, 
	n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, 
	n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, 
	n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, 
	n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, 
	n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, 
	n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, 
	n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, 
	n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, 
	n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, 
	n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
	n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, 
	n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, 
	n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, 
	n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, 
	n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, 
	n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, 
	n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, 
	n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, 
	n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, 
	n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, 
	n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, 
	n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, 
	n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, 
	n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, 
	n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, 
	n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, 
	n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, 
	n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, 
	n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, 
	n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, 
	n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, 
	n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, 
	n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, 
	n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, 
	n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, 
	n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, 
	n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, 
	n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, 
	n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, 
	n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, 
	n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, 
	n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, 
	n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, 
	n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, 
	n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, 
	n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, 
	n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, 
	n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, 
	n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, 
	n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, 
	n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, 
	n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, 
	n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, 
	n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, 
	n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, 
	n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, 
	n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, 
	n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, 
	n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, 
	n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, 
	n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, 
	n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, 
	n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, 
	n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, 
	n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, 
	n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, 
	n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, 
	n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
	n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, 
	n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, 
	n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, 
	n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, 
	n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, 
	n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, 
	n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, 
	n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, 
	n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, 
	n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, 
	n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, 
	n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, 
	n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, 
	n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, 
	n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, 
	n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, 
	n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, 
	n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, 
	n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, 
	n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, 
	n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, 
	n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, 
	n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, 
	n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, 
	n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, 
	n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, 
	n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, 
	n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, 
	n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, 
	n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, 
	n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, 
	n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, 
	n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, 
	n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, 
	n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, 
	n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, 
	n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, 
	n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, 
	n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, 
	n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, 
	n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, 
	n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, 
	n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, 
	n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, 
	n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, 
	n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, 
	n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, 
	n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, 
	n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, 
	n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, 
	n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, 
	n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, 
	n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, 
	n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, 
	n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, 
	n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, 
	n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
	n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, 
	n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, 
	n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, 
	n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, 
	n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, 
	n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, 
	n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, 
	n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, 
	n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, 
	n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, 
	n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, 
	n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, 
	n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, 
	n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, 
	n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, 
	n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, 
	n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, 
	n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, 
	n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, 
	n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, 
	n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, 
	n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, 
	n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, 
	n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, 
	n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, 
	n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, 
	n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, 
	n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, 
	n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, 
	n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, 
	n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, 
	n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, 
	n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, 
	n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, 
	n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, 
	n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, 
	n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, 
	n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, 
	n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, 
	n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, 
	n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, 
	n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, 
	n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, 
	n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, 
	n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, 
	n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, 
	n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, 
	n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, 
	n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, 
	n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, 
	n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, 
	n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, 
	n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, 
	n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, 
	n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, 
	n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, 
	n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, 
	n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, 
	n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, 
	n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, 
	n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, 
	n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, 
	n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, 
	n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, 
	n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, 
	n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, 
	n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, 
	n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, 
	n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, 
	n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, 
	n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, 
	n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, 
	n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, 
	n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, 
	n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, 
	n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, 
	n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, 
	n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, 
	n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, 
	n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, 
	n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, 
	n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, 
	n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, 
	n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, 
	n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, 
	n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, 
	n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, 
	n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, 
	n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, 
	n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, 
	n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, 
	n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, 
	n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, 
	n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, 
	n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, 
	n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, 
	n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, 
	n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, 
	n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, 
	n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, 
	n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, 
	n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, 
	n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, 
	n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, 
	n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, 
	n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, 
	n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, 
	n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, 
	n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, 
	n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, 
	n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, 
	n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, 
	n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, 
	n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, 
	n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, 
	n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, 
	n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, 
	n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, 
	n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, 
	n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, 
	n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, 
	n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, 
	n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, 
	n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, 
	n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, 
	n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, 
	n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, 
	n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, 
	n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, 
	n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, 
	n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, 
	n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, 
	n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, 
	n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, 
	n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, 
	n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, 
	n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, 
	n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, 
	n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, 
	n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, 
	n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, 
	n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, 
	n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, 
	n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, 
	n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, 
	n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, 
	n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, 
	n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, 
	n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, 
	n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, 
	n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, 
	n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, 
	n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, 
	n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, 
	n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, 
	n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, 
	n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, 
	n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, 
	n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, 
	n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, 
	n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, 
	n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, 
	n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, 
	n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, 
	n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, 
	n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, 
	n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, 
	n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, 
	n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, 
	n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, 
	n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, 
	n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, 
	n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, 
	n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, 
	n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, 
	n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, 
	n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, 
	n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, 
	n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, 
	n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, 
	n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, 
	n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, 
	n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, 
	n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, 
	n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, 
	n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, 
	n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, 
	n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, 
	n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, 
	n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, 
	n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, 
	n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, 
	n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, 
	n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, 
	n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, 
	n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, 
	n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, 
	n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, 
	n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, 
	n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, 
	n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, 
	n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, 
	n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, 
	n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, 
	n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, 
	n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, 
	n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, 
	n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, 
	n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, 
	n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, 
	n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, 
	n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, 
	n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, 
	n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, 
	n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, 
	n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, 
	n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, 
	n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, 
	n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, 
	n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, 
	n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, 
	n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, 
	n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, 
	n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, 
	n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, 
	n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, 
	n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, 
	n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, 
	n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, 
	n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, 
	n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, 
	n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, 
	n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, 
	n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, 
	n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, 
	n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, 
	n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, 
	n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, 
	n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, 
	n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, 
	n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, 
	n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, 
	n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, 
	n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, 
	n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, 
	n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, 
	n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, 
	n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, 
	n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, 
	n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, 
	n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, 
	n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, 
	n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, 
	n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, 
	n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, 
	n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, 
	n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, 
	n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, 
	n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, 
	n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, 
	n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, 
	n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, 
	n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, 
	n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, 
	n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, 
	n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, 
	n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, 
	n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, 
	n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, 
	n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, 
	n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, 
	n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, 
	n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, 
	n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, 
	n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, 
	n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, 
	n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, 
	n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, 
	n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, 
	n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, 
	n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, 
	n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, 
	n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, 
	n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, 
	n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, 
	n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, 
	n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, 
	n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, 
	n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, 
	n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, 
	n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, 
	n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, 
	n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, 
	n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, 
	n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, 
	n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, 
	n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, 
	n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, 
	n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, 
	n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, 
	n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, 
	n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, 
	n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, 
	n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, 
	n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, 
	n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, 
	n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, 
	n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, 
	n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, 
	n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, 
	n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, 
	n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, 
	n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, 
	n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, 
	n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, 
	n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, 
	n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, 
	n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, 
	n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, 
	n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, 
	n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, 
	n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, 
	n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, 
	n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, 
	n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, 
	n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, 
	n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, 
	n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, 
	n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, 
	n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, 
	n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, 
	n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, 
	n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, 
	n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, 
	n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, 
	n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, 
	n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, 
	n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, 
	n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, 
	n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, 
	n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, 
	n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, 
	n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, 
	n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, 
	n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, 
	n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, 
	n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, 
	n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, 
	n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, 
	n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, 
	n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, 
	n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, 
	n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, 
	n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, 
	n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, 
	n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, 
	n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, 
	n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, 
	n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, 
	n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, 
	n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, 
	n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, 
	n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, 
	n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, 
	n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, 
	n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, 
	n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, 
	n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, 
	n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, 
	n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, 
	n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, 
	n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, 
	n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, 
	n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, 
	n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, 
	n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, 
	n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, 
	n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, 
	n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, 
	n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, 
	n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, 
	n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, 
	n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, 
	n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, 
	n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, 
	n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, 
	n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, 
	n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, 
	n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, 
	n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, 
	n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, 
	n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, 
	n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, 
	n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, 
	n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, 
	n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, 
	n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, 
	n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, 
	n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, 
	n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, 
	n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, 
	n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, 
	n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, 
	n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, 
	n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, 
	n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, 
	n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, 
	n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, 
	n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, 
	n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, 
	n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, 
	n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, 
	n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, 
	n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, 
	n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, 
	n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, 
	n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, 
	n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, 
	n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, 
	n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, 
	n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, 
	n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, 
	n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, 
	n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, 
	n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, 
	n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, 
	n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, 
	n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, 
	n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, 
	n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, 
	n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, 
	n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, 
	n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, 
	n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, 
	n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, 
	n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, 
	n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, 
	n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, 
	n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, 
	n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, 
	n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, 
	n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, 
	n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, 
	n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, 
	n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, 
	n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, 
	n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, 
	n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, 
	n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, 
	n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, 
	n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, 
	n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, 
	n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, 
	n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, 
	n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, 
	n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, 
	n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, 
	n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, 
	n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, 
	n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, 
	n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, 
	n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, 
	n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, 
	n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, 
	n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, 
	n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, 
	n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, 
	n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, 
	n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, 
	n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, 
	n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, 
	n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, 
	n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, 
	n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, 
	n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, 
	n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, 
	n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, 
	n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, 
	n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, 
	n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, 
	n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, 
	n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, 
	n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, 
	n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, 
	n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, 
	n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, 
	n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, 
	n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, 
	n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, 
	n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, 
	n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, 
	n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, 
	n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, 
	n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, 
	n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, 
	n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, 
	n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, 
	n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, 
	n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, 
	n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, 
	n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, 
	n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, 
	n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, 
	n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, 
	n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, 
	n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, 
	n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, 
	n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, 
	n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, 
	n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, 
	n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, 
	n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, 
	n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, 
	n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, 
	n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, 
	n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, 
	n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, 
	n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, 
	n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, 
	n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, 
	n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, 
	n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, 
	n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, 
	n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, 
	n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, 
	n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, 
	n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, 
	n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, 
	n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, 
	n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, 
	n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, 
	n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, 
	n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, 
	n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, 
	n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, 
	n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, 
	n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, 
	n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, 
	n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, 
	n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, 
	n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, 
	n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, 
	n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, 
	n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, 
	n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, 
	n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, 
	n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, 
	n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, 
	n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, 
	n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, 
	n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, 
	n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, 
	n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, 
	n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, 
	n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, 
	n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, 
	n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, 
	n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, 
	n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, 
	n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, 
	n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, 
	n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, 
	n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, 
	n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, 
	n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, 
	n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, 
	n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, 
	n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, 
	n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, 
	n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, 
	n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, 
	n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, 
	n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, 
	n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, 
	n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, 
	n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, 
	n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, 
	n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, 
	n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, 
	n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, 
	n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, 
	n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, 
	n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, 
	n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, 
	n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, 
	n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, 
	n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, 
	n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, 
	n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, 
	n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, 
	n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, 
	n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, 
	n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, 
	n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, 
	n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, 
	n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, 
	n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, 
	n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, 
	n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, 
	n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, 
	n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, 
	n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, 
	n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, 
	n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, 
	n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, 
	n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, 
	n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, 
	n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, 
	n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, 
	n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, 
	n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, 
	n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, 
	n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, 
	n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, 
	n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, 
	n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, 
	n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, 
	n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, 
	n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, 
	n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, 
	n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, 
	n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, 
	n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, 
	n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, 
	n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, 
	n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, 
	n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, 
	n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, 
	n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, 
	n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, 
	n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, 
	n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, 
	n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, 
	n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, 
	n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, 
	n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, 
	n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, 
	n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, 
	n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, 
	n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, 
	n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, 
	n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, 
	n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, 
	n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, 
	n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, 
	n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, 
	n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, 
	n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, 
	n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, 
	n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, 
	n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, 
	n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, 
	n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, 
	n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, 
	n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, 
	n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, 
	n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, 
	n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, 
	n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, 
	n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, 
	n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, 
	n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, 
	n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, 
	n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, 
	n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, 
	n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, 
	n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, 
	n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, 
	n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, 
	n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, 
	n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, 
	n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, 
	n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, 
	n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, 
	n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, 
	n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, 
	n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, 
	n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, 
	n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, 
	n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, 
	n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, 
	n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, 
	n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, 
	n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, 
	n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, 
	n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, 
	n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, 
	n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, 
	n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, 
	n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, 
	n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, 
	n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, 
	n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, 
	n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, 
	n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, 
	n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, 
	n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, 
	n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, 
	n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, 
	n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, 
	n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, 
	n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, 
	n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, 
	n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, 
	n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, 
	n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, 
	n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, 
	n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, 
	n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, 
	n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, 
	n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, 
	n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, 
	n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, 
	n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, 
	n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, 
	n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, 
	n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, 
	n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, 
	n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, 
	n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, 
	n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, 
	n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, 
	n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, 
	n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, 
	n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, 
	n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, 
	n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, 
	n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, 
	n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, 
	n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, 
	n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, 
	n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, 
	n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, 
	n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, 
	n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, 
	n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, 
	n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, 
	n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, 
	n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, 
	n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, 
	n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, 
	n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, 
	n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, 
	n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, 
	n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, 
	n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, 
	n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, 
	n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, 
	n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, 
	n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, 
	n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, 
	n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, 
	n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, 
	n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, 
	n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, 
	n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, 
	n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, 
	n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, 
	n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, 
	n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, 
	n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, 
	n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, 
	n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, 
	n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, 
	n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, 
	n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, 
	n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, 
	n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, 
	n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, 
	n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, 
	n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, 
	n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, 
	n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, 
	n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, 
	n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, 
	n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, 
	n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, 
	n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, 
	n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, 
	n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, 
	n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, 
	n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, 
	n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, 
	n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, 
	n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, 
	n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, 
	n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, 
	n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, 
	n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, 
	n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, 
	n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, 
	n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, 
	n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, 
	n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, 
	n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, 
	n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, 
	n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, 
	n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, 
	n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, 
	n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, 
	n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, 
	n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, 
	n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, 
	n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, 
	n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, 
	n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, 
	n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, 
	n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, 
	n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, 
	n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, 
	n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, 
	n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, 
	n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, 
	n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, 
	n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, 
	n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, 
	n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, 
	n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, 
	n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, 
	n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, 
	n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, 
	n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, 
	n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, 
	n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, 
	n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, 
	n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, 
	n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, 
	n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, 
	n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, 
	n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, 
	n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, 
	n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, 
	n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, 
	n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, 
	n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, 
	n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, 
	n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, 
	n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, 
	n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, 
	n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, 
	n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, 
	n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, 
	n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, 
	n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, 
	n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, 
	n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, 
	n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, 
	n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, 
	n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, 
	n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, 
	n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, 
	n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, 
	n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, 
	n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, 
	n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, 
	n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, 
	n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, 
	n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, 
	n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, 
	n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, 
	n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, 
	n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, 
	n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, 
	n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, 
	n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, 
	n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, 
	n24570, n24571, n24572, n24573, n24574, n24575;

wire c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, 
	c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, 
	c20, c21, c22, c23, c24, c25, c26, c27, c28, c29, 
	c30, c31, c32, c33, c34, c35, c36, c37, c38, c39, 
	c40, c41, c42, c43, c44, c45, c46, c47, c48, c49, 
	c50, c51, c52, c53, c54, c55, c56, c57, c58, c59, 
	c60, c61, c62, c63, c64, c65, c66, c67, c68, c69, 
	c70, c71, c72, c73, c74, c75, c76, c77, c78, c79, 
	c80, c81, c82, c83, c84, c85, c86, c87, c88, c89, 
	c90, c91, c92, c93, c94, c95, c96, c97, c98, c99, 
	c100, c101, c102, c103, c104, c105, c106, c107, c108, c109, 
	c110, c111, c112, c113, c114, c115, c116, c117, c118, c119, 
	c120, c121, c122, c123, c124, c125, c126, c127, c128, c129, 
	c130, c131, c132, c133, c134, c135, c136, c137, c138, c139, 
	c140, c141, c142, c143, c144, c145, c146, c147, c148, c149, 
	c150, c151, c152, c153, c154, c155, c156, c157, c158, c159, 
	c160, c161, c162, c163, c164, c165, c166, c167, c168, c169, 
	c170, c171, c172, c173, c174, c175, c176, c177, c178, c179, 
	c180, c181, c182, c183, c184, c185, c186, c187, c188, c189, 
	c190, c191, c192, c193, c194, c195, c196, c197, c198, c199, 
	c200, c201, c202, c203, c204, c205, c206, c207, c208, c209, 
	c210, c211, c212, c213, c214, c215, c216, c217, c218, c219, 
	c220, c221, c222, c223, c224, c225, c226, c227, c228, c229, 
	c230, c231, c232, c233, c234, c235, c236, c237, c238, c239, 
	c240, c241, c242, c243, c244, c245, c246, c247, c248, c249, 
	c250, c251, c252, c253, c254, c255, c256, c257, c258, c259, 
	c260, c261, c262, c263, c264, c265, c266, c267, c268, c269, 
	c270, c271, c272, c273, c274, c275, c276, c277, c278, c279, 
	c280, c281, c282, c283, c284, c285, c286, c287, c288, c289, 
	c290, c291, c292, c293, c294, c295, c296, c297, c298, c299, 
	c300, c301, c302, c303, c304, c305, c306, c307, c308, c309, 
	c310, c311, c312, c313, c314, c315, c316, c317, c318, c319, 
	c320, c321, c322, c323, c324, c325, c326, c327, c328, c329, 
	c330, c331, c332, c333, c334, c335, c336, c337, c338, c339, 
	c340, c341, c342, c343, c344, c345, c346, c347, c348, c349, 
	c350, c351, c352, c353, c354, c355, c356, c357, c358, c359, 
	c360, c361, c362, c363, c364, c365, c366, c367, c368, c369, 
	c370, c371, c372, c373, c374, c375, c376, c377, c378, c379, 
	c380, c381, c382, c383, c384, c385, c386, c387, c388, c389, 
	c390, c391, c392, c393, c394, c395, c396, c397, c398, c399, 
	c400, c401, c402, c403, c404, c405, c406, c407, c408, c409, 
	c410, c411, c412, c413, c414, c415, c416, c417, c418, c419, 
	c420, c421, c422, c423, c424, c425, c426, c427, c428, c429, 
	c430, c431, c432, c433, c434, c435, c436, c437, c438, c439, 
	c440, c441, c442, c443, c444, c445, c446, c447, c448, c449, 
	c450, c451, c452, c453, c454, c455, c456, c457, c458, c459, 
	c460, c461, c462, c463, c464, c465, c466, c467, c468, c469, 
	c470, c471, c472, c473, c474, c475, c476, c477, c478, c479, 
	c480, c481, c482, c483, c484, c485, c486, c487, c488, c489, 
	c490, c491, c492, c493, c494, c495, c496, c497, c498, c499, 
	c500, c501, c502, c503, c504, c505, c506, c507, c508, c509, 
	c510, c511, c512, c513, c514, c515, c516, c517, c518, c519, 
	c520, c521, c522, c523, c524, c525, c526, c527, c528, c529, 
	c530, c531, c532, c533, c534, c535, c536, c537, c538, c539, 
	c540, c541, c542, c543, c544, c545, c546, c547, c548, c549, 
	c550, c551, c552, c553, c554, c555, c556, c557, c558, c559, 
	c560, c561, c562, c563, c564, c565, c566, c567, c568, c569, 
	c570, c571, c572, c573, c574, c575, c576, c577, c578, c579, 
	c580, c581, c582, c583, c584, c585, c586, c587, c588, c589, 
	c590, c591, c592, c593, c594, c595, c596, c597, c598, c599, 
	c600, c601, c602, c603, c604, c605, c606, c607, c608, c609, 
	c610, c611, c612, c613, c614, c615, c616, c617, c618, c619, 
	c620, c621, c622, c623, c624, c625, c626, c627, c628, c629, 
	c630, c631, c632, c633, c634, c635, c636, c637, c638, c639, 
	c640, c641, c642, c643, c644, c645, c646, c647, c648, c649, 
	c650, c651, c652, c653, c654, c655, c656, c657, c658, c659, 
	c660, c661, c662, c663, c664, c665, c666, c667, c668, c669, 
	c670, c671, c672, c673, c674, c675, c676, c677, c678, c679, 
	c680, c681, c682, c683, c684, c685, c686, c687, c688, c689, 
	c690, c691, c692, c693, c694, c695, c696, c697, c698, c699, 
	c700, c701, c702, c703, c704, c705, c706, c707, c708, c709, 
	c710, c711, c712, c713, c714, c715, c716, c717, c718, c719, 
	c720, c721, c722, c723, c724, c725, c726, c727, c728, c729, 
	c730, c731, c732, c733, c734, c735, c736, c737, c738, c739, 
	c740, c741, c742, c743, c744, c745, c746, c747, c748, c749, 
	c750, c751, c752, c753, c754, c755, c756, c757, c758, c759, 
	c760, c761, c762, c763, c764, c765, c766, c767, c768, c769, 
	c770, c771, c772, c773, c774, c775, c776, c777, c778, c779, 
	c780, c781, c782, c783, c784, c785, c786, c787, c788, c789, 
	c790, c791, c792, c793, c794, c795, c796, c797, c798, c799, 
	c800, c801, c802, c803, c804, c805, c806, c807, c808, c809, 
	c810, c811, c812, c813, c814, c815, c816, c817, c818, c819, 
	c820, c821, c822, c823, c824, c825, c826, c827, c828, c829, 
	c830, c831, c832, c833, c834, c835, c836, c837, c838, c839, 
	c840, c841, c842, c843, c844, c845, c846, c847, c848, c849, 
	c850, c851, c852, c853, c854, c855, c856, c857, c858, c859, 
	c860, c861, c862, c863, c864, c865, c866, c867, c868, c869, 
	c870, c871, c872, c873, c874, c875, c876, c877, c878, c879, 
	c880, c881, c882, c883, c884, c885, c886, c887, c888, c889, 
	c890, c891, c892, c893, c894, c895, c896, c897, c898, c899, 
	c900, c901, c902, c903, c904, c905, c906, c907, c908, c909, 
	c910, c911, c912, c913, c914, c915, c916, c917, c918, c919, 
	c920, c921, c922, c923, c924, c925, c926, c927, c928, c929, 
	c930, c931, c932, c933, c934, c935, c936, c937, c938, c939, 
	c940, c941, c942, c943, c944, c945, c946, c947, c948, c949, 
	c950, c951, c952, c953, c954, c955, c956, c957, c958, c959, 
	c960, c961, c962, c963, c964, c965, c966, c967, c968, c969, 
	c970, c971, c972, c973, c974, c975, c976, c977, c978, c979, 
	c980, c981, c982, c983, c984, c985, c986, c987, c988, c989, 
	c990, c991, c992, c993, c994, c995, c996, c997, c998, c999, 
	c1000, c1001, c1002, c1003, c1004, c1005, c1006, c1007, c1008, c1009, 
	c1010, c1011, c1012, c1013, c1014, c1015, c1016, c1017, c1018, c1019, 
	c1020, c1021, c1022, c1023, c1024, c1025, c1026, c1027, c1028, c1029, 
	c1030, c1031, c1032, c1033, c1034, c1035, c1036, c1037, c1038, c1039, 
	c1040, c1041, c1042, c1043, c1044, c1045, c1046, c1047, c1048, c1049, 
	c1050, c1051, c1052, c1053, c1054, c1055, c1056, c1057, c1058, c1059, 
	c1060, c1061, c1062, c1063, c1064, c1065, c1066, c1067, c1068, c1069, 
	c1070, c1071, c1072, c1073, c1074, c1075, c1076, c1077, c1078, c1079, 
	c1080, c1081, c1082, c1083, c1084, c1085, c1086, c1087, c1088, c1089, 
	c1090, c1091, c1092, c1093, c1094, c1095, c1096, c1097, c1098, c1099, 
	c1100, c1101, c1102, c1103, c1104, c1105, c1106, c1107, c1108, c1109, 
	c1110, c1111, c1112, c1113, c1114, c1115, c1116, c1117, c1118, c1119, 
	c1120, c1121, c1122, c1123, c1124, c1125, c1126, c1127, c1128, c1129, 
	c1130, c1131, c1132, c1133, c1134, c1135, c1136, c1137, c1138, c1139, 
	c1140, c1141, c1142, c1143, c1144, c1145, c1146, c1147, c1148, c1149, 
	c1150, c1151, c1152, c1153, c1154, c1155, c1156, c1157, c1158, c1159, 
	c1160, c1161, c1162, c1163, c1164, c1165, c1166, c1167, c1168, c1169, 
	c1170, c1171, c1172, c1173, c1174, c1175, c1176, c1177, c1178, c1179, 
	c1180, c1181, c1182, c1183, c1184, c1185, c1186, c1187, c1188, c1189, 
	c1190, c1191, c1192, c1193, c1194, c1195, c1196, c1197, c1198, c1199, 
	c1200, c1201, c1202, c1203, c1204, c1205, c1206, c1207, c1208, c1209, 
	c1210, c1211, c1212, c1213, c1214, c1215, c1216, c1217, c1218, c1219, 
	c1220, c1221, c1222, c1223, c1224, c1225, c1226, c1227, c1228, c1229, 
	c1230, c1231, c1232, c1233, c1234, c1235, c1236, c1237, c1238, c1239, 
	c1240, c1241, c1242, c1243, c1244, c1245, c1246, c1247, c1248, c1249, 
	c1250, c1251, c1252, c1253, c1254, c1255, c1256, c1257, c1258, c1259, 
	c1260, c1261, c1262, c1263, c1264, c1265, c1266, c1267, c1268, c1269, 
	c1270, c1271, c1272, c1273, c1274, c1275, c1276, c1277, c1278, c1279, 
	c1280, c1281, c1282, c1283, c1284, c1285, c1286, c1287, c1288, c1289, 
	c1290, c1291, c1292, c1293, c1294, c1295, c1296, c1297, c1298, c1299, 
	c1300, c1301, c1302, c1303, c1304, c1305, c1306, c1307, c1308, c1309, 
	c1310, c1311, c1312, c1313, c1314, c1315, c1316, c1317, c1318, c1319, 
	c1320, c1321, c1322, c1323, c1324, c1325, c1326, c1327, c1328, c1329, 
	c1330, c1331, c1332, c1333, c1334, c1335, c1336, c1337, c1338, c1339, 
	c1340, c1341, c1342, c1343, c1344, c1345, c1346, c1347, c1348, c1349, 
	c1350, c1351, c1352, c1353, c1354, c1355, c1356, c1357, c1358, c1359, 
	c1360, c1361, c1362, c1363, c1364, c1365, c1366, c1367, c1368, c1369, 
	c1370, c1371, c1372, c1373, c1374, c1375, c1376, c1377, c1378, c1379, 
	c1380, c1381, c1382, c1383, c1384, c1385, c1386, c1387, c1388, c1389, 
	c1390, c1391, c1392, c1393, c1394, c1395, c1396, c1397, c1398, c1399, 
	c1400, c1401, c1402, c1403, c1404, c1405, c1406, c1407, c1408, c1409, 
	c1410, c1411, c1412, c1413, c1414, c1415, c1416, c1417, c1418, c1419, 
	c1420, c1421, c1422, c1423, c1424, c1425, c1426, c1427, c1428, c1429, 
	c1430, c1431, c1432, c1433, c1434, c1435, c1436, c1437, c1438, c1439, 
	c1440, c1441, c1442, c1443, c1444, c1445, c1446, c1447, c1448, c1449, 
	c1450, c1451, c1452, c1453, c1454, c1455, c1456, c1457, c1458, c1459, 
	c1460, c1461, c1462, c1463, c1464, c1465, c1466, c1467, c1468, c1469, 
	c1470, c1471, c1472, c1473, c1474, c1475, c1476, c1477, c1478, c1479, 
	c1480, c1481, c1482, c1483, c1484, c1485, c1486, c1487, c1488, c1489, 
	c1490, c1491, c1492, c1493, c1494, c1495, c1496, c1497, c1498, c1499, 
	c1500, c1501, c1502, c1503, c1504, c1505, c1506, c1507, c1508, c1509, 
	c1510, c1511, c1512, c1513, c1514, c1515, c1516, c1517, c1518, c1519, 
	c1520, c1521, c1522, c1523, c1524, c1525, c1526, c1527, c1528, c1529, 
	c1530, c1531, c1532, c1533, c1534, c1535, c1536, c1537, c1538, c1539, 
	c1540, c1541, c1542, c1543, c1544, c1545, c1546, c1547, c1548, c1549, 
	c1550, c1551, c1552, c1553, c1554, c1555, c1556, c1557, c1558, c1559, 
	c1560, c1561, c1562, c1563, c1564, c1565, c1566, c1567, c1568, c1569, 
	c1570, c1571, c1572, c1573, c1574, c1575, c1576, c1577, c1578, c1579, 
	c1580, c1581, c1582, c1583, c1584, c1585, c1586, c1587, c1588, c1589, 
	c1590, c1591, c1592, c1593, c1594, c1595, c1596, c1597, c1598, c1599, 
	c1600, c1601, c1602, c1603, c1604, c1605, c1606, c1607, c1608, c1609, 
	c1610, c1611, c1612, c1613, c1614, c1615, c1616, c1617, c1618, c1619, 
	c1620, c1621, c1622, c1623, c1624, c1625, c1626, c1627, c1628, c1629, 
	c1630, c1631, c1632, c1633, c1634, c1635, c1636, c1637, c1638, c1639, 
	c1640, c1641, c1642, c1643, c1644, c1645, c1646, c1647, c1648, c1649, 
	c1650, c1651, c1652, c1653, c1654, c1655, c1656, c1657, c1658, c1659, 
	c1660, c1661, c1662, c1663, c1664, c1665, c1666, c1667, c1668, c1669, 
	c1670, c1671, c1672, c1673, c1674, c1675, c1676, c1677, c1678, c1679, 
	c1680, c1681, c1682, c1683, c1684, c1685, c1686, c1687, c1688, c1689, 
	c1690, c1691, c1692, c1693, c1694, c1695, c1696, c1697, c1698, c1699, 
	c1700, c1701, c1702, c1703, c1704, c1705, c1706, c1707, c1708, c1709, 
	c1710, c1711, c1712, c1713, c1714, c1715, c1716, c1717, c1718, c1719, 
	c1720, c1721, c1722, c1723, c1724, c1725, c1726, c1727, c1728, c1729, 
	c1730, c1731, c1732, c1733, c1734, c1735, c1736, c1737, c1738, c1739, 
	c1740, c1741, c1742, c1743, c1744, c1745, c1746, c1747, c1748, c1749, 
	c1750, c1751, c1752, c1753, c1754, c1755, c1756, c1757, c1758, c1759, 
	c1760, c1761, c1762, c1763, c1764, c1765, c1766, c1767, c1768, c1769, 
	c1770, c1771, c1772, c1773, c1774, c1775, c1776, c1777, c1778, c1779, 
	c1780, c1781, c1782, c1783, c1784, c1785, c1786, c1787, c1788, c1789, 
	c1790, c1791, c1792, c1793, c1794, c1795, c1796, c1797, c1798, c1799, 
	c1800, c1801, c1802, c1803, c1804, c1805, c1806, c1807, c1808, c1809, 
	c1810, c1811, c1812, c1813, c1814, c1815, c1816, c1817, c1818, c1819, 
	c1820, c1821, c1822, c1823, c1824, c1825, c1826, c1827, c1828, c1829, 
	c1830, c1831, c1832, c1833, c1834, c1835, c1836, c1837, c1838, c1839, 
	c1840, c1841, c1842, c1843, c1844, c1845, c1846, c1847, c1848, c1849, 
	c1850, c1851, c1852, c1853, c1854, c1855, c1856, c1857, c1858, c1859, 
	c1860, c1861, c1862, c1863, c1864, c1865, c1866, c1867, c1868, c1869, 
	c1870, c1871, c1872, c1873, c1874, c1875, c1876, c1877, c1878, c1879, 
	c1880, c1881, c1882, c1883, c1884, c1885, c1886, c1887, c1888, c1889, 
	c1890, c1891, c1892, c1893, c1894, c1895, c1896, c1897, c1898, c1899, 
	c1900, c1901, c1902, c1903, c1904, c1905, c1906, c1907, c1908, c1909, 
	c1910, c1911, c1912, c1913, c1914, c1915, c1916, c1917, c1918, c1919, 
	c1920, c1921, c1922, c1923, c1924, c1925, c1926, c1927, c1928, c1929, 
	c1930, c1931, c1932, c1933, c1934, c1935, c1936, c1937, c1938, c1939, 
	c1940, c1941, c1942, c1943, c1944, c1945, c1946, c1947, c1948, c1949, 
	c1950, c1951, c1952, c1953, c1954, c1955, c1956, c1957, c1958, c1959, 
	c1960, c1961, c1962, c1963, c1964, c1965, c1966, c1967, c1968, c1969, 
	c1970, c1971, c1972, c1973, c1974, c1975, c1976, c1977, c1978, c1979, 
	c1980, c1981, c1982, c1983, c1984, c1985, c1986, c1987, c1988, c1989, 
	c1990, c1991, c1992, c1993, c1994, c1995, c1996, c1997, c1998, c1999, 
	c2000, c2001, c2002, c2003, c2004, c2005, c2006, c2007, c2008, c2009, 
	c2010, c2011, c2012, c2013, c2014, c2015, c2016, c2017, c2018, c2019, 
	c2020, c2021, c2022, c2023, c2024, c2025, c2026, c2027, c2028, c2029, 
	c2030, c2031, c2032, c2033, c2034, c2035, c2036, c2037, c2038, c2039, 
	c2040, c2041, c2042, c2043, c2044, c2045, c2046, c2047, c2048, c2049, 
	c2050, c2051, c2052, c2053, c2054, c2055, c2056, c2057, c2058, c2059, 
	c2060, c2061, c2062, c2063, c2064, c2065, c2066, c2067, c2068, c2069, 
	c2070, c2071, c2072, c2073, c2074, c2075, c2076, c2077, c2078, c2079, 
	c2080, c2081, c2082, c2083, c2084, c2085, c2086, c2087, c2088, c2089, 
	c2090, c2091, c2092, c2093, c2094, c2095, c2096, c2097, c2098, c2099, 
	c2100, c2101, c2102, c2103, c2104, c2105, c2106, c2107, c2108, c2109, 
	c2110, c2111, c2112, c2113, c2114, c2115, c2116, c2117, c2118, c2119, 
	c2120, c2121, c2122, c2123, c2124, c2125, c2126, c2127, c2128, c2129, 
	c2130, c2131, c2132, c2133, c2134, c2135, c2136, c2137, c2138, c2139, 
	c2140, c2141, c2142, c2143, c2144, c2145, c2146, c2147, c2148, c2149, 
	c2150, c2151, c2152, c2153, c2154, c2155, c2156, c2157, c2158, c2159, 
	c2160, c2161, c2162, c2163, c2164, c2165, c2166, c2167, c2168, c2169, 
	c2170, c2171, c2172, c2173, c2174, c2175, c2176, c2177, c2178, c2179, 
	c2180, c2181, c2182, c2183, c2184, c2185, c2186, c2187, c2188, c2189, 
	c2190, c2191, c2192, c2193, c2194, c2195, c2196, c2197, c2198, c2199, 
	c2200, c2201, c2202, c2203, c2204, c2205, c2206, c2207, c2208, c2209, 
	c2210, c2211, c2212, c2213, c2214, c2215, c2216, c2217, c2218, c2219, 
	c2220, c2221, c2222, c2223, c2224, c2225, c2226, c2227, c2228, c2229, 
	c2230, c2231, c2232, c2233, c2234, c2235, c2236, c2237, c2238, c2239, 
	c2240, c2241, c2242, c2243, c2244, c2245, c2246, c2247, c2248, c2249, 
	c2250, c2251, c2252, c2253, c2254, c2255, c2256, c2257, c2258, c2259, 
	c2260, c2261, c2262, c2263, c2264, c2265, c2266, c2267, c2268, c2269, 
	c2270, c2271, c2272, c2273, c2274, c2275, c2276, c2277, c2278, c2279, 
	c2280, c2281, c2282, c2283, c2284, c2285, c2286, c2287, c2288, c2289, 
	c2290, c2291, c2292, c2293, c2294, c2295, c2296, c2297, c2298, c2299, 
	c2300, c2301, c2302, c2303, c2304, c2305, c2306, c2307, c2308, c2309, 
	c2310, c2311, c2312, c2313, c2314, c2315, c2316, c2317, c2318, c2319, 
	c2320, c2321, c2322, c2323, c2324, c2325, c2326, c2327, c2328, c2329, 
	c2330, c2331, c2332, c2333, c2334, c2335, c2336, c2337, c2338, c2339, 
	c2340, c2341, c2342, c2343, c2344, c2345, c2346, c2347, c2348, c2349, 
	c2350, c2351, c2352, c2353, c2354, c2355, c2356, c2357, c2358, c2359, 
	c2360, c2361, c2362, c2363, c2364, c2365, c2366, c2367, c2368, c2369, 
	c2370, c2371, c2372, c2373, c2374, c2375, c2376, c2377, c2378, c2379, 
	c2380, c2381, c2382, c2383, c2384, c2385, c2386, c2387, c2388, c2389, 
	c2390, c2391, c2392, c2393, c2394, c2395, c2396, c2397, c2398, c2399, 
	c2400, c2401, c2402, c2403, c2404, c2405, c2406, c2407, c2408, c2409, 
	c2410, c2411, c2412, c2413, c2414, c2415, c2416, c2417, c2418, c2419, 
	c2420, c2421, c2422, c2423, c2424, c2425, c2426, c2427, c2428, c2429, 
	c2430, c2431, c2432, c2433, c2434, c2435, c2436, c2437, c2438, c2439, 
	c2440, c2441, c2442, c2443, c2444, c2445, c2446, c2447, c2448, c2449, 
	c2450, c2451, c2452, c2453, c2454, c2455, c2456, c2457, c2458, c2459, 
	c2460, c2461, c2462, c2463, c2464, c2465, c2466, c2467, c2468, c2469, 
	c2470, c2471, c2472, c2473, c2474, c2475, c2476, c2477, c2478, c2479, 
	c2480, c2481, c2482, c2483, c2484, c2485, c2486, c2487, c2488, c2489, 
	c2490, c2491, c2492, c2493, c2494, c2495, c2496, c2497, c2498, c2499, 
	c2500, c2501, c2502, c2503, c2504, c2505, c2506, c2507, c2508, c2509, 
	c2510, c2511, c2512, c2513, c2514, c2515, c2516, c2517, c2518, c2519, 
	c2520, c2521, c2522, c2523, c2524, c2525, c2526, c2527, c2528, c2529, 
	c2530, c2531, c2532, c2533, c2534, c2535, c2536, c2537, c2538, c2539, 
	c2540, c2541, c2542, c2543, c2544, c2545, c2546, c2547, c2548, c2549, 
	c2550, c2551, c2552, c2553, c2554, c2555, c2556, c2557, c2558, c2559, 
	c2560, c2561, c2562, c2563, c2564, c2565, c2566, c2567, c2568, c2569, 
	c2570, c2571, c2572, c2573, c2574, c2575, c2576, c2577, c2578, c2579, 
	c2580, c2581, c2582, c2583, c2584, c2585, c2586, c2587, c2588, c2589, 
	c2590, c2591, c2592, c2593, c2594, c2595, c2596, c2597, c2598, c2599, 
	c2600, c2601, c2602, c2603, c2604, c2605, c2606, c2607, c2608, c2609, 
	c2610, c2611, c2612, c2613, c2614, c2615, c2616, c2617, c2618, c2619, 
	c2620, c2621, c2622, c2623, c2624, c2625, c2626, c2627, c2628, c2629, 
	c2630, c2631, c2632, c2633, c2634, c2635, c2636, c2637, c2638, c2639, 
	c2640, c2641, c2642, c2643, c2644, c2645, c2646, c2647, c2648, c2649, 
	c2650, c2651, c2652, c2653, c2654, c2655, c2656, c2657, c2658, c2659, 
	c2660, c2661, c2662, c2663, c2664, c2665, c2666, c2667, c2668, c2669, 
	c2670, c2671, c2672, c2673, c2674, c2675, c2676, c2677, c2678, c2679, 
	c2680, c2681, c2682, c2683, c2684, c2685, c2686, c2687, c2688, c2689, 
	c2690, c2691, c2692, c2693, c2694, c2695, c2696, c2697, c2698, c2699, 
	c2700, c2701, c2702, c2703, c2704, c2705, c2706, c2707, c2708, c2709, 
	c2710, c2711, c2712, c2713, c2714, c2715, c2716, c2717, c2718, c2719, 
	c2720, c2721, c2722, c2723, c2724, c2725, c2726, c2727, c2728, c2729, 
	c2730, c2731, c2732, c2733, c2734, c2735, c2736, c2737, c2738, c2739, 
	c2740, c2741, c2742, c2743, c2744, c2745, c2746, c2747, c2748, c2749, 
	c2750, c2751, c2752, c2753, c2754, c2755, c2756, c2757, c2758, c2759, 
	c2760, c2761, c2762, c2763, c2764, c2765, c2766, c2767, c2768, c2769, 
	c2770, c2771, c2772, c2773, c2774, c2775, c2776, c2777, c2778, c2779, 
	c2780, c2781, c2782, c2783, c2784, c2785, c2786, c2787, c2788, c2789, 
	c2790, c2791, c2792, c2793, c2794, c2795, c2796, c2797, c2798, c2799, 
	c2800, c2801, c2802, c2803, c2804, c2805, c2806, c2807, c2808, c2809, 
	c2810, c2811, c2812, c2813, c2814, c2815, c2816, c2817, c2818, c2819, 
	c2820, c2821, c2822, c2823, c2824, c2825, c2826, c2827, c2828, c2829, 
	c2830, c2831, c2832, c2833, c2834, c2835, c2836, c2837, c2838, c2839, 
	c2840, c2841, c2842, c2843, c2844, c2845, c2846, c2847, c2848, c2849, 
	c2850, c2851, c2852, c2853, c2854, c2855, c2856, c2857, c2858, c2859, 
	c2860, c2861, c2862, c2863, c2864, c2865, c2866, c2867, c2868, c2869, 
	c2870, c2871, c2872, c2873, c2874, c2875, c2876, c2877, c2878, c2879, 
	c2880, c2881, c2882, c2883, c2884, c2885, c2886, c2887, c2888, c2889, 
	c2890, c2891, c2892, c2893, c2894, c2895, c2896, c2897, c2898, c2899, 
	c2900, c2901, c2902, c2903, c2904, c2905, c2906, c2907, c2908, c2909, 
	c2910, c2911, c2912, c2913, c2914, c2915, c2916, c2917, c2918, c2919, 
	c2920, c2921, c2922, c2923, c2924, c2925, c2926, c2927, c2928, c2929, 
	c2930, c2931, c2932, c2933, c2934, c2935, c2936, c2937, c2938, c2939, 
	c2940, c2941, c2942, c2943, c2944, c2945, c2946, c2947, c2948, c2949, 
	c2950, c2951, c2952, c2953, c2954, c2955, c2956, c2957, c2958, c2959, 
	c2960, c2961, c2962, c2963, c2964, c2965, c2966, c2967, c2968, c2969, 
	c2970, c2971, c2972, c2973, c2974, c2975, c2976, c2977, c2978, c2979, 
	c2980, c2981, c2982, c2983, c2984, c2985, c2986, c2987, c2988, c2989, 
	c2990, c2991, c2992, c2993, c2994, c2995, c2996, c2997, c2998, c2999, 
	c3000, c3001, c3002, c3003, c3004, c3005, c3006, c3007, c3008, c3009, 
	c3010, c3011, c3012, c3013, c3014, c3015, c3016, c3017, c3018, c3019, 
	c3020, c3021, c3022, c3023, c3024, c3025, c3026, c3027, c3028, c3029, 
	c3030, c3031, c3032, c3033, c3034, c3035, c3036, c3037, c3038, c3039, 
	c3040, c3041, c3042, c3043, c3044, c3045, c3046, c3047, c3048, c3049, 
	c3050, c3051, c3052, c3053, c3054, c3055, c3056, c3057, c3058, c3059, 
	c3060, c3061, c3062, c3063, c3064, c3065, c3066, c3067, c3068, c3069, 
	c3070, c3071, c3072, c3073, c3074, c3075, c3076, c3077, c3078, c3079, 
	c3080, c3081, c3082, c3083, c3084, c3085, c3086, c3087, c3088, c3089, 
	c3090, c3091, c3092, c3093, c3094, c3095, c3096, c3097, c3098, c3099, 
	c3100, c3101, c3102, c3103, c3104, c3105, c3106, c3107, c3108, c3109, 
	c3110, c3111, c3112, c3113, c3114, c3115, c3116, c3117, c3118, c3119, 
	c3120, c3121, c3122, c3123, c3124, c3125, c3126, c3127, c3128, c3129, 
	c3130, c3131, c3132, c3133, c3134, c3135, c3136, c3137, c3138, c3139, 
	c3140, c3141, c3142, c3143, c3144, c3145, c3146, c3147, c3148, c3149, 
	c3150, c3151, c3152, c3153, c3154, c3155, c3156, c3157, c3158, c3159, 
	c3160, c3161, c3162, c3163, c3164, c3165, c3166, c3167, c3168, c3169, 
	c3170, c3171, c3172, c3173, c3174, c3175, c3176, c3177, c3178, c3179, 
	c3180, c3181, c3182, c3183, c3184, c3185, c3186, c3187, c3188, c3189, 
	c3190, c3191, c3192, c3193, c3194, c3195, c3196, c3197, c3198, c3199, 
	c3200, c3201, c3202, c3203, c3204, c3205, c3206, c3207, c3208, c3209, 
	c3210, c3211, c3212, c3213, c3214, c3215, c3216, c3217, c3218, c3219, 
	c3220, c3221, c3222, c3223, c3224, c3225, c3226, c3227, c3228, c3229, 
	c3230, c3231, c3232, c3233, c3234, c3235, c3236, c3237, c3238, c3239, 
	c3240, c3241, c3242, c3243, c3244, c3245, c3246, c3247, c3248, c3249, 
	c3250, c3251, c3252, c3253, c3254, c3255, c3256, c3257, c3258, c3259, 
	c3260, c3261, c3262, c3263, c3264, c3265, c3266, c3267, c3268, c3269, 
	c3270, c3271, c3272, c3273, c3274, c3275, c3276, c3277, c3278, c3279, 
	c3280, c3281, c3282, c3283, c3284, c3285, c3286, c3287, c3288, c3289, 
	c3290, c3291, c3292, c3293, c3294, c3295, c3296, c3297, c3298, c3299, 
	c3300, c3301, c3302, c3303, c3304, c3305, c3306, c3307, c3308, c3309, 
	c3310, c3311, c3312, c3313, c3314, c3315, c3316, c3317, c3318, c3319, 
	c3320, c3321, c3322, c3323, c3324, c3325, c3326, c3327, c3328, c3329, 
	c3330, c3331, c3332, c3333, c3334, c3335, c3336, c3337, c3338, c3339, 
	c3340, c3341, c3342, c3343, c3344, c3345, c3346, c3347, c3348, c3349, 
	c3350, c3351, c3352, c3353, c3354, c3355, c3356, c3357, c3358, c3359, 
	c3360, c3361, c3362, c3363, c3364, c3365, c3366, c3367, c3368, c3369, 
	c3370, c3371, c3372, c3373, c3374, c3375, c3376, c3377, c3378, c3379, 
	c3380, c3381, c3382, c3383, c3384, c3385, c3386, c3387, c3388, c3389, 
	c3390, c3391, c3392, c3393, c3394, c3395, c3396, c3397, c3398, c3399, 
	c3400, c3401, c3402, c3403, c3404, c3405, c3406, c3407, c3408, c3409, 
	c3410, c3411, c3412, c3413, c3414, c3415, c3416, c3417, c3418, c3419, 
	c3420, c3421, c3422, c3423, c3424, c3425, c3426, c3427, c3428, c3429, 
	c3430, c3431, c3432, c3433, c3434, c3435, c3436, c3437, c3438, c3439, 
	c3440, c3441, c3442, c3443, c3444, c3445, c3446, c3447, c3448, c3449, 
	c3450, c3451, c3452, c3453, c3454, c3455, c3456, c3457, c3458, c3459, 
	c3460, c3461, c3462, c3463, c3464, c3465, c3466, c3467, c3468, c3469, 
	c3470, c3471, c3472, c3473, c3474, c3475, c3476, c3477, c3478, c3479, 
	c3480, c3481, c3482, c3483, c3484, c3485, c3486, c3487, c3488, c3489, 
	c3490, c3491, c3492, c3493, c3494, c3495, c3496, c3497, c3498, c3499, 
	c3500, c3501, c3502, c3503, c3504, c3505, c3506, c3507, c3508, c3509, 
	c3510, c3511, c3512, c3513, c3514, c3515, c3516, c3517, c3518, c3519, 
	c3520, c3521, c3522, c3523, c3524, c3525, c3526, c3527, c3528, c3529, 
	c3530, c3531, c3532, c3533, c3534, c3535, c3536, c3537, c3538, c3539, 
	c3540, c3541, c3542, c3543, c3544, c3545, c3546, c3547, c3548, c3549, 
	c3550, c3551, c3552, c3553, c3554, c3555, c3556, c3557, c3558, c3559, 
	c3560, c3561, c3562, c3563, c3564, c3565, c3566, c3567, c3568, c3569, 
	c3570, c3571, c3572, c3573, c3574, c3575, c3576, c3577, c3578, c3579, 
	c3580, c3581, c3582, c3583, c3584, c3585, c3586, c3587, c3588, c3589, 
	c3590, c3591, c3592, c3593, c3594, c3595, c3596, c3597, c3598, c3599, 
	c3600, c3601, c3602, c3603, c3604, c3605, c3606, c3607, c3608, c3609, 
	c3610, c3611, c3612, c3613, c3614, c3615, c3616, c3617, c3618, c3619, 
	c3620, c3621, c3622, c3623, c3624, c3625, c3626, c3627, c3628, c3629, 
	c3630, c3631, c3632, c3633, c3634, c3635, c3636, c3637, c3638, c3639, 
	c3640, c3641, c3642, c3643, c3644, c3645, c3646, c3647, c3648, c3649, 
	c3650, c3651, c3652, c3653, c3654, c3655, c3656, c3657, c3658, c3659, 
	c3660, c3661, c3662, c3663, c3664, c3665, c3666, c3667, c3668, c3669, 
	c3670, c3671, c3672, c3673, c3674, c3675, c3676, c3677, c3678, c3679, 
	c3680, c3681, c3682, c3683, c3684, c3685, c3686, c3687, c3688, c3689, 
	c3690, c3691, c3692, c3693, c3694, c3695, c3696, c3697, c3698, c3699, 
	c3700, c3701, c3702, c3703, c3704, c3705, c3706, c3707, c3708, c3709, 
	c3710, c3711, c3712, c3713, c3714, c3715, c3716, c3717, c3718, c3719, 
	c3720, c3721, c3722, c3723, c3724, c3725, c3726, c3727, c3728, c3729, 
	c3730, c3731, c3732, c3733, c3734, c3735, c3736, c3737, c3738, c3739, 
	c3740, c3741, c3742, c3743, c3744, c3745, c3746, c3747, c3748, c3749, 
	c3750, c3751, c3752, c3753, c3754, c3755, c3756, c3757, c3758, c3759, 
	c3760, c3761, c3762, c3763, c3764, c3765, c3766, c3767, c3768, c3769, 
	c3770, c3771, c3772, c3773, c3774, c3775, c3776, c3777, c3778, c3779, 
	c3780, c3781, c3782, c3783, c3784, c3785, c3786, c3787, c3788, c3789, 
	c3790, c3791, c3792, c3793, c3794, c3795, c3796, c3797, c3798, c3799, 
	c3800, c3801, c3802, c3803, c3804, c3805, c3806, c3807, c3808, c3809, 
	c3810, c3811, c3812, c3813, c3814, c3815, c3816, c3817, c3818, c3819, 
	c3820, c3821, c3822, c3823, c3824, c3825, c3826, c3827, c3828, c3829, 
	c3830, c3831, c3832, c3833, c3834, c3835, c3836, c3837, c3838, c3839, 
	c3840, c3841, c3842, c3843, c3844, c3845, c3846, c3847, c3848, c3849, 
	c3850, c3851, c3852, c3853, c3854, c3855, c3856, c3857, c3858, c3859, 
	c3860, c3861, c3862, c3863, c3864, c3865, c3866, c3867, c3868, c3869, 
	c3870, c3871, c3872, c3873, c3874, c3875, c3876, c3877, c3878, c3879, 
	c3880, c3881, c3882, c3883, c3884, c3885, c3886, c3887, c3888, c3889, 
	c3890, c3891, c3892, c3893, c3894, c3895, c3896, c3897, c3898, c3899, 
	c3900, c3901, c3902, c3903, c3904, c3905, c3906, c3907, c3908, c3909, 
	c3910, c3911, c3912, c3913, c3914, c3915, c3916, c3917, c3918, c3919, 
	c3920, c3921, c3922, c3923, c3924, c3925, c3926, c3927, c3928, c3929, 
	c3930, c3931, c3932, c3933, c3934, c3935, c3936, c3937, c3938, c3939, 
	c3940, c3941, c3942, c3943, c3944, c3945, c3946, c3947, c3948, c3949, 
	c3950, c3951, c3952, c3953, c3954, c3955, c3956, c3957, c3958, c3959, 
	c3960, c3961, c3962, c3963, c3964, c3965, c3966, c3967, c3968, c3969, 
	c3970, c3971, c3972, c3973, c3974, c3975, c3976, c3977, c3978, c3979, 
	c3980, c3981, c3982, c3983, c3984, c3985, c3986, c3987, c3988, c3989, 
	c3990, c3991, c3992, c3993, c3994, c3995, c3996, c3997, c3998, c3999, 
	c4000, c4001, c4002, c4003, c4004, c4005, c4006, c4007, c4008, c4009, 
	c4010, c4011, c4012, c4013, c4014, c4015, c4016, c4017, c4018, c4019, 
	c4020, c4021, c4022, c4023, c4024, c4025, c4026, c4027, c4028, c4029, 
	c4030, c4031, c4032, c4033, c4034, c4035, c4036, c4037, c4038, c4039, 
	c4040, c4041, c4042, c4043, c4044, c4045, c4046, c4047, c4048, c4049, 
	c4050, c4051, c4052, c4053, c4054, c4055, c4056, c4057, c4058, c4059, 
	c4060, c4061, c4062, c4063, c4064, c4065, c4066, c4067, c4068, c4069, 
	c4070, c4071, c4072, c4073, c4074, c4075, c4076, c4077, c4078, c4079, 
	c4080, c4081, c4082, c4083, c4084, c4085, c4086, c4087, c4088, c4089, 
	c4090, c4091, c4092, c4093, c4094, c4095, c4096, c4097, c4098, c4099, 
	c4100, c4101, c4102, c4103, c4104, c4105, c4106, c4107, c4108, c4109, 
	c4110, c4111, c4112, c4113, c4114, c4115, c4116, c4117, c4118, c4119, 
	c4120, c4121, c4122, c4123, c4124, c4125, c4126, c4127, c4128, c4129, 
	c4130, c4131, c4132, c4133, c4134, c4135, c4136, c4137, c4138, c4139, 
	c4140, c4141, c4142, c4143, c4144, c4145, c4146, c4147, c4148, c4149, 
	c4150, c4151, c4152, c4153, c4154, c4155, c4156, c4157, c4158, c4159, 
	c4160, c4161, c4162, c4163, c4164, c4165, c4166, c4167, c4168, c4169, 
	c4170, c4171, c4172, c4173, c4174, c4175, c4176, c4177, c4178, c4179, 
	c4180, c4181, c4182, c4183, c4184, c4185, c4186, c4187, c4188, c4189, 
	c4190, c4191, c4192, c4193, c4194, c4195, c4196, c4197, c4198, c4199, 
	c4200, c4201, c4202, c4203, c4204, c4205, c4206, c4207, c4208, c4209, 
	c4210, c4211, c4212, c4213, c4214, c4215, c4216, c4217, c4218, c4219, 
	c4220, c4221, c4222, c4223, c4224, c4225, c4226, c4227, c4228, c4229, 
	c4230, c4231, c4232, c4233, c4234, c4235, c4236, c4237, c4238, c4239, 
	c4240, c4241, c4242, c4243, c4244, c4245, c4246, c4247, c4248, c4249, 
	c4250, c4251, c4252, c4253, c4254, c4255, c4256, c4257, c4258, c4259, 
	c4260, c4261, c4262, c4263, c4264, c4265, c4266, c4267, c4268, c4269, 
	c4270, c4271, c4272, c4273, c4274, c4275, c4276, c4277, c4278, c4279, 
	c4280, c4281, c4282, c4283, c4284, c4285, c4286, c4287, c4288, c4289, 
	c4290, c4291, c4292, c4293, c4294, c4295, c4296, c4297, c4298, c4299, 
	c4300, c4301, c4302, c4303, c4304, c4305, c4306, c4307, c4308, c4309, 
	c4310, c4311, c4312, c4313, c4314, c4315, c4316, c4317, c4318, c4319, 
	c4320, c4321, c4322, c4323, c4324, c4325, c4326, c4327, c4328, c4329, 
	c4330, c4331, c4332, c4333, c4334, c4335, c4336, c4337, c4338, c4339, 
	c4340, c4341, c4342, c4343, c4344, c4345, c4346, c4347, c4348, c4349, 
	c4350, c4351, c4352, c4353, c4354, c4355, c4356, c4357, c4358, c4359, 
	c4360, c4361, c4362, c4363, c4364, c4365, c4366, c4367, c4368, c4369, 
	c4370, c4371, c4372, c4373, c4374, c4375, c4376, c4377, c4378, c4379, 
	c4380, c4381, c4382, c4383, c4384, c4385, c4386, c4387, c4388, c4389, 
	c4390, c4391, c4392, c4393, c4394, c4395, c4396, c4397, c4398, c4399, 
	c4400, c4401, c4402, c4403, c4404, c4405, c4406, c4407, c4408, c4409, 
	c4410, c4411, c4412, c4413, c4414, c4415, c4416, c4417, c4418, c4419, 
	c4420, c4421, c4422, c4423, c4424, c4425, c4426, c4427, c4428, c4429, 
	c4430, c4431, c4432, c4433, c4434, c4435, c4436, c4437, c4438, c4439, 
	c4440, c4441, c4442, c4443, c4444, c4445, c4446, c4447, c4448, c4449, 
	c4450, c4451, c4452, c4453, c4454, c4455, c4456, c4457, c4458, c4459, 
	c4460, c4461, c4462, c4463, c4464, c4465, c4466, c4467, c4468, c4469, 
	c4470, c4471, c4472, c4473, c4474, c4475, c4476, c4477, c4478, c4479, 
	c4480, c4481, c4482, c4483, c4484, c4485, c4486, c4487, c4488, c4489, 
	c4490, c4491, c4492, c4493, c4494, c4495, c4496, c4497, c4498, c4499, 
	c4500, c4501, c4502, c4503, c4504, c4505, c4506, c4507, c4508, c4509, 
	c4510, c4511, c4512, c4513, c4514, c4515, c4516, c4517, c4518, c4519, 
	c4520, c4521, c4522, c4523, c4524, c4525, c4526, c4527, c4528, c4529, 
	c4530, c4531, c4532, c4533, c4534, c4535, c4536, c4537, c4538, c4539, 
	c4540, c4541, c4542, c4543, c4544, c4545, c4546, c4547, c4548, c4549, 
	c4550, c4551, c4552, c4553, c4554, c4555, c4556, c4557, c4558, c4559, 
	c4560, c4561, c4562, c4563, c4564, c4565, c4566, c4567, c4568, c4569, 
	c4570, c4571, c4572, c4573, c4574, c4575, c4576, c4577, c4578, c4579, 
	c4580, c4581, c4582, c4583, c4584, c4585, c4586, c4587, c4588, c4589, 
	c4590, c4591, c4592, c4593, c4594, c4595, c4596, c4597, c4598, c4599, 
	c4600, c4601, c4602, c4603, c4604, c4605, c4606, c4607, c4608, c4609, 
	c4610, c4611, c4612, c4613, c4614, c4615, c4616, c4617, c4618, c4619, 
	c4620, c4621, c4622, c4623, c4624, c4625, c4626, c4627, c4628, c4629, 
	c4630, c4631, c4632, c4633, c4634, c4635, c4636, c4637, c4638, c4639, 
	c4640, c4641, c4642, c4643, c4644, c4645, c4646, c4647, c4648, c4649, 
	c4650, c4651, c4652, c4653, c4654, c4655, c4656, c4657, c4658, c4659, 
	c4660, c4661, c4662, c4663, c4664, c4665, c4666, c4667, c4668, c4669, 
	c4670, c4671, c4672, c4673, c4674, c4675, c4676, c4677, c4678, c4679, 
	c4680, c4681, c4682, c4683, c4684, c4685, c4686, c4687, c4688, c4689, 
	c4690, c4691, c4692, c4693, c4694, c4695, c4696, c4697, c4698, c4699, 
	c4700, c4701, c4702, c4703, c4704, c4705, c4706, c4707, c4708, c4709, 
	c4710, c4711, c4712, c4713, c4714, c4715, c4716, c4717, c4718, c4719, 
	c4720, c4721, c4722, c4723, c4724, c4725, c4726, c4727, c4728, c4729, 
	c4730, c4731, c4732, c4733, c4734, c4735, c4736, c4737, c4738, c4739, 
	c4740, c4741, c4742, c4743, c4744, c4745, c4746, c4747, c4748, c4749, 
	c4750, c4751, c4752, c4753, c4754, c4755, c4756, c4757, c4758, c4759, 
	c4760, c4761, c4762, c4763, c4764, c4765, c4766, c4767, c4768, c4769, 
	c4770, c4771, c4772, c4773, c4774, c4775, c4776, c4777, c4778, c4779, 
	c4780, c4781, c4782, c4783, c4784, c4785, c4786, c4787, c4788, c4789, 
	c4790, c4791, c4792, c4793, c4794, c4795, c4796, c4797, c4798, c4799, 
	c4800, c4801, c4802, c4803, c4804, c4805, c4806, c4807, c4808, c4809, 
	c4810, c4811, c4812, c4813, c4814, c4815, c4816, c4817, c4818, c4819, 
	c4820, c4821, c4822, c4823, c4824, c4825, c4826, c4827, c4828, c4829, 
	c4830, c4831, c4832, c4833, c4834, c4835, c4836, c4837, c4838, c4839, 
	c4840, c4841, c4842, c4843, c4844, c4845, c4846, c4847, c4848, c4849, 
	c4850, c4851, c4852, c4853, c4854, c4855, c4856, c4857, c4858, c4859, 
	c4860, c4861, c4862, c4863, c4864, c4865, c4866, c4867, c4868, c4869, 
	c4870, c4871, c4872, c4873, c4874, c4875, c4876, c4877, c4878, c4879, 
	c4880, c4881, c4882, c4883, c4884, c4885, c4886, c4887, c4888, c4889, 
	c4890, c4891, c4892, c4893, c4894, c4895, c4896, c4897, c4898, c4899, 
	c4900, c4901, c4902, c4903, c4904, c4905, c4906, c4907, c4908, c4909, 
	c4910, c4911, c4912, c4913, c4914, c4915, c4916, c4917, c4918, c4919, 
	c4920, c4921, c4922, c4923, c4924, c4925, c4926, c4927, c4928, c4929, 
	c4930, c4931, c4932, c4933, c4934, c4935, c4936, c4937, c4938, c4939, 
	c4940, c4941, c4942, c4943, c4944, c4945, c4946, c4947, c4948, c4949, 
	c4950, c4951, c4952, c4953, c4954, c4955, c4956, c4957, c4958, c4959, 
	c4960, c4961, c4962, c4963, c4964, c4965, c4966, c4967, c4968, c4969, 
	c4970, c4971, c4972, c4973, c4974, c4975, c4976, c4977, c4978, c4979, 
	c4980, c4981, c4982, c4983, c4984, c4985, c4986, c4987, c4988, c4989, 
	c4990, c4991, c4992, c4993, c4994, c4995, c4996, c4997, c4998, c4999, 
	c5000, c5001, c5002, c5003, c5004, c5005, c5006, c5007, c5008, c5009, 
	c5010, c5011, c5012, c5013, c5014, c5015, c5016, c5017, c5018, c5019, 
	c5020, c5021, c5022, c5023, c5024, c5025, c5026, c5027, c5028, c5029, 
	c5030, c5031, c5032, c5033, c5034, c5035, c5036, c5037, c5038, c5039, 
	c5040, c5041, c5042, c5043, c5044, c5045, c5046, c5047, c5048, c5049, 
	c5050, c5051, c5052, c5053, c5054, c5055, c5056, c5057, c5058, c5059, 
	c5060, c5061, c5062, c5063, c5064, c5065, c5066, c5067, c5068, c5069, 
	c5070, c5071, c5072, c5073, c5074, c5075, c5076, c5077, c5078, c5079, 
	c5080, c5081, c5082, c5083, c5084, c5085, c5086, c5087, c5088, c5089, 
	c5090, c5091, c5092, c5093, c5094, c5095, c5096, c5097, c5098, c5099, 
	c5100, c5101, c5102, c5103, c5104, c5105, c5106, c5107, c5108, c5109, 
	c5110, c5111, c5112, c5113, c5114, c5115, c5116, c5117, c5118, c5119, 
	c5120, c5121, c5122, c5123, c5124, c5125, c5126, c5127, c5128, c5129, 
	c5130, c5131, c5132, c5133, c5134, c5135, c5136, c5137, c5138, c5139, 
	c5140, c5141, c5142, c5143, c5144, c5145, c5146, c5147, c5148, c5149, 
	c5150, c5151, c5152, c5153, c5154, c5155, c5156, c5157, c5158, c5159, 
	c5160, c5161, c5162, c5163, c5164, c5165, c5166, c5167, c5168, c5169, 
	c5170, c5171, c5172, c5173, c5174, c5175, c5176, c5177, c5178, c5179, 
	c5180, c5181, c5182, c5183, c5184, c5185, c5186, c5187, c5188, c5189, 
	c5190, c5191, c5192, c5193, c5194, c5195, c5196, c5197, c5198, c5199, 
	c5200, c5201, c5202, c5203, c5204, c5205, c5206, c5207, c5208, c5209, 
	c5210, c5211, c5212, c5213, c5214, c5215, c5216, c5217, c5218, c5219, 
	c5220, c5221, c5222, c5223, c5224, c5225, c5226, c5227, c5228, c5229, 
	c5230, c5231, c5232, c5233, c5234, c5235, c5236, c5237, c5238, c5239, 
	c5240, c5241, c5242, c5243, c5244, c5245, c5246, c5247, c5248, c5249, 
	c5250, c5251, c5252, c5253, c5254, c5255, c5256, c5257, c5258, c5259, 
	c5260, c5261, c5262, c5263, c5264, c5265, c5266, c5267, c5268, c5269, 
	c5270, c5271, c5272, c5273, c5274, c5275, c5276, c5277, c5278, c5279, 
	c5280, c5281, c5282, c5283, c5284, c5285, c5286, c5287, c5288, c5289, 
	c5290, c5291, c5292, c5293, c5294, c5295, c5296, c5297, c5298, c5299, 
	c5300, c5301, c5302, c5303, c5304, c5305, c5306, c5307, c5308, c5309, 
	c5310, c5311, c5312, c5313, c5314, c5315, c5316, c5317, c5318, c5319, 
	c5320, c5321, c5322, c5323, c5324, c5325, c5326, c5327, c5328, c5329, 
	c5330, c5331, c5332, c5333, c5334, c5335, c5336, c5337, c5338, c5339, 
	c5340, c5341, c5342, c5343, c5344, c5345, c5346, c5347, c5348, c5349, 
	c5350, c5351, c5352, c5353, c5354, c5355, c5356, c5357, c5358, c5359, 
	c5360, c5361, c5362, c5363, c5364, c5365, c5366, c5367, c5368, c5369, 
	c5370, c5371, c5372, c5373, c5374, c5375, c5376, c5377, c5378, c5379, 
	c5380, c5381, c5382, c5383, c5384, c5385, c5386, c5387, c5388, c5389, 
	c5390, c5391, c5392, c5393, c5394, c5395, c5396, c5397, c5398, c5399, 
	c5400, c5401, c5402, c5403, c5404, c5405, c5406, c5407, c5408, c5409, 
	c5410, c5411, c5412, c5413, c5414, c5415, c5416, c5417, c5418, c5419, 
	c5420, c5421, c5422, c5423, c5424, c5425, c5426, c5427, c5428, c5429, 
	c5430, c5431, c5432, c5433, c5434, c5435, c5436, c5437, c5438, c5439, 
	c5440, c5441, c5442, c5443, c5444, c5445, c5446, c5447, c5448, c5449, 
	c5450, c5451, c5452, c5453, c5454, c5455, c5456, c5457, c5458, c5459, 
	c5460, c5461, c5462, c5463, c5464, c5465, c5466, c5467, c5468, c5469, 
	c5470, c5471, c5472, c5473, c5474, c5475, c5476, c5477, c5478, c5479, 
	c5480, c5481, c5482, c5483, c5484, c5485, c5486, c5487, c5488, c5489, 
	c5490, c5491, c5492, c5493, c5494, c5495, c5496, c5497, c5498, c5499, 
	c5500, c5501, c5502, c5503, c5504, c5505, c5506, c5507, c5508, c5509, 
	c5510, c5511, c5512, c5513, c5514, c5515, c5516, c5517, c5518, c5519, 
	c5520, c5521, c5522, c5523, c5524, c5525, c5526, c5527, c5528, c5529, 
	c5530, c5531, c5532, c5533, c5534, c5535, c5536, c5537, c5538, c5539, 
	c5540, c5541, c5542, c5543, c5544, c5545, c5546, c5547, c5548, c5549, 
	c5550, c5551, c5552, c5553, c5554, c5555, c5556, c5557, c5558, c5559, 
	c5560, c5561, c5562, c5563, c5564, c5565, c5566, c5567, c5568, c5569, 
	c5570, c5571, c5572, c5573, c5574, c5575, c5576, c5577, c5578, c5579, 
	c5580, c5581, c5582, c5583, c5584, c5585, c5586, c5587, c5588, c5589, 
	c5590, c5591, c5592, c5593, c5594, c5595, c5596, c5597, c5598, c5599, 
	c5600, c5601, c5602, c5603, c5604, c5605, c5606, c5607, c5608, c5609, 
	c5610, c5611, c5612, c5613, c5614, c5615, c5616, c5617, c5618, c5619, 
	c5620, c5621, c5622, c5623, c5624, c5625, c5626, c5627, c5628, c5629, 
	c5630, c5631, c5632, c5633, c5634, c5635, c5636, c5637, c5638, c5639, 
	c5640, c5641, c5642, c5643, c5644, c5645, c5646, c5647, c5648, c5649, 
	c5650, c5651, c5652, c5653, c5654, c5655, c5656, c5657, c5658, c5659, 
	c5660, c5661, c5662, c5663, c5664, c5665, c5666, c5667, c5668, c5669, 
	c5670, c5671, c5672, c5673, c5674, c5675, c5676, c5677, c5678, c5679, 
	c5680, c5681, c5682, c5683, c5684, c5685, c5686, c5687, c5688, c5689, 
	c5690, c5691, c5692, c5693, c5694, c5695, c5696, c5697, c5698, c5699, 
	c5700, c5701, c5702, c5703, c5704, c5705, c5706, c5707, c5708, c5709, 
	c5710, c5711, c5712, c5713, c5714, c5715, c5716, c5717, c5718, c5719, 
	c5720, c5721, c5722, c5723, c5724, c5725, c5726, c5727, c5728, c5729, 
	c5730, c5731, c5732, c5733, c5734, c5735, c5736, c5737, c5738, c5739, 
	c5740, c5741, c5742, c5743, c5744, c5745, c5746, c5747, c5748, c5749, 
	c5750, c5751, c5752, c5753, c5754, c5755, c5756, c5757, c5758, c5759, 
	c5760, c5761, c5762, c5763, c5764, c5765, c5766, c5767, c5768, c5769, 
	c5770, c5771, c5772, c5773, c5774, c5775, c5776, c5777, c5778, c5779, 
	c5780, c5781, c5782, c5783, c5784, c5785, c5786, c5787, c5788, c5789, 
	c5790, c5791, c5792, c5793, c5794, c5795, c5796, c5797, c5798, c5799, 
	c5800, c5801, c5802, c5803, c5804, c5805, c5806, c5807, c5808, c5809, 
	c5810, c5811, c5812, c5813, c5814, c5815, c5816, c5817, c5818, c5819, 
	c5820, c5821, c5822, c5823, c5824, c5825, c5826, c5827, c5828, c5829, 
	c5830, c5831, c5832, c5833, c5834, c5835, c5836, c5837, c5838, c5839, 
	c5840, c5841, c5842, c5843, c5844, c5845, c5846, c5847, c5848, c5849, 
	c5850, c5851, c5852, c5853, c5854, c5855, c5856, c5857, c5858, c5859, 
	c5860, c5861, c5862, c5863, c5864, c5865, c5866, c5867, c5868, c5869, 
	c5870, c5871, c5872, c5873, c5874, c5875, c5876, c5877, c5878, c5879, 
	c5880, c5881, c5882, c5883, c5884, c5885, c5886, c5887, c5888, c5889, 
	c5890, c5891, c5892, c5893, c5894, c5895, c5896, c5897, c5898, c5899, 
	c5900, c5901, c5902, c5903, c5904, c5905, c5906, c5907, c5908, c5909, 
	c5910, c5911, c5912, c5913, c5914, c5915, c5916, c5917, c5918, c5919, 
	c5920, c5921, c5922, c5923, c5924, c5925, c5926, c5927, c5928, c5929, 
	c5930, c5931, c5932, c5933, c5934, c5935, c5936, c5937, c5938, c5939, 
	c5940, c5941, c5942, c5943, c5944, c5945, c5946, c5947, c5948, c5949, 
	c5950, c5951, c5952, c5953, c5954, c5955, c5956, c5957, c5958, c5959, 
	c5960, c5961, c5962, c5963, c5964, c5965, c5966, c5967, c5968, c5969, 
	c5970, c5971, c5972, c5973, c5974, c5975, c5976, c5977, c5978, c5979, 
	c5980, c5981, c5982, c5983, c5984, c5985, c5986, c5987, c5988, c5989, 
	c5990, c5991, c5992, c5993, c5994, c5995, c5996, c5997, c5998, c5999, 
	c6000, c6001, c6002, c6003, c6004, c6005, c6006, c6007, c6008, c6009, 
	c6010, c6011, c6012, c6013, c6014, c6015, c6016, c6017, c6018, c6019, 
	c6020, c6021, c6022, c6023, c6024, c6025, c6026, c6027, c6028, c6029, 
	c6030, c6031, c6032, c6033, c6034, c6035, c6036, c6037, c6038, c6039, 
	c6040, c6041, c6042, c6043, c6044, c6045, c6046, c6047, c6048, c6049, 
	c6050, c6051, c6052, c6053, c6054, c6055, c6056, c6057, c6058, c6059, 
	c6060, c6061, c6062, c6063, c6064, c6065, c6066, c6067, c6068, c6069, 
	c6070, c6071, c6072, c6073, c6074, c6075, c6076, c6077, c6078, c6079, 
	c6080, c6081, c6082, c6083, c6084, c6085, c6086, c6087, c6088, c6089, 
	c6090, c6091, c6092, c6093, c6094, c6095, c6096, c6097, c6098, c6099, 
	c6100, c6101, c6102, c6103, c6104, c6105, c6106, c6107, c6108, c6109, 
	c6110, c6111, c6112, c6113, c6114, c6115, c6116, c6117, c6118, c6119, 
	c6120, c6121, c6122, c6123, c6124, c6125, c6126, c6127, c6128, c6129, 
	c6130, c6131, c6132, c6133, c6134, c6135, c6136, c6137, c6138, c6139, 
	c6140, c6141, c6142, c6143, c6144, c6145, c6146, c6147, c6148, c6149, 
	c6150, c6151, c6152, c6153, c6154, c6155, c6156, c6157, c6158, c6159, 
	c6160, c6161, c6162, c6163, c6164, c6165, c6166, c6167, c6168, c6169, 
	c6170, c6171, c6172, c6173, c6174, c6175, c6176, c6177, c6178, c6179, 
	c6180, c6181, c6182, c6183, c6184, c6185, c6186, c6187, c6188, c6189, 
	c6190, c6191, c6192, c6193, c6194, c6195, c6196, c6197, c6198, c6199, 
	c6200, c6201, c6202, c6203, c6204, c6205, c6206, c6207, c6208, c6209, 
	c6210, c6211, c6212, c6213, c6214, c6215, c6216, c6217, c6218, c6219, 
	c6220, c6221, c6222, c6223, c6224, c6225, c6226, c6227, c6228, c6229, 
	c6230, c6231, c6232, c6233, c6234, c6235, c6236, c6237, c6238, c6239, 
	c6240, c6241, c6242, c6243, c6244, c6245, c6246, c6247, c6248, c6249, 
	c6250, c6251, c6252, c6253, c6254, c6255, c6256, c6257, c6258, c6259, 
	c6260, c6261, c6262, c6263, c6264, c6265, c6266, c6267, c6268, c6269, 
	c6270, c6271, c6272, c6273, c6274, c6275, c6276, c6277, c6278, c6279, 
	c6280, c6281, c6282, c6283, c6284, c6285, c6286, c6287, c6288, c6289, 
	c6290, c6291, c6292, c6293, c6294, c6295, c6296, c6297, c6298, c6299, 
	c6300, c6301, c6302, c6303, c6304, c6305, c6306, c6307, c6308, c6309, 
	c6310, c6311, c6312, c6313, c6314, c6315, c6316, c6317, c6318, c6319, 
	c6320, c6321, c6322, c6323, c6324, c6325, c6326, c6327, c6328, c6329, 
	c6330, c6331, c6332, c6333, c6334, c6335, c6336, c6337, c6338, c6339, 
	c6340, c6341, c6342, c6343, c6344, c6345, c6346, c6347, c6348, c6349, 
	c6350, c6351, c6352, c6353, c6354, c6355, c6356, c6357, c6358, c6359, 
	c6360, c6361, c6362, c6363, c6364, c6365, c6366, c6367, c6368, c6369, 
	c6370, c6371, c6372, c6373, c6374, c6375, c6376, c6377, c6378, c6379, 
	c6380, c6381, c6382, c6383, c6384, c6385, c6386, c6387, c6388, c6389, 
	c6390, c6391, c6392, c6393, c6394, c6395, c6396, c6397, c6398, c6399, 
	c6400, c6401, c6402, c6403, c6404, c6405, c6406, c6407, c6408, c6409, 
	c6410, c6411, c6412, c6413, c6414, c6415, c6416, c6417, c6418, c6419, 
	c6420, c6421, c6422, c6423, c6424, c6425, c6426, c6427, c6428, c6429, 
	c6430, c6431, c6432, c6433, c6434, c6435, c6436, c6437, c6438, c6439, 
	c6440, c6441, c6442, c6443, c6444, c6445, c6446, c6447, c6448, c6449, 
	c6450, c6451, c6452, c6453, c6454, c6455, c6456, c6457, c6458, c6459, 
	c6460, c6461, c6462, c6463, c6464, c6465, c6466, c6467, c6468, c6469, 
	c6470, c6471, c6472, c6473, c6474, c6475, c6476, c6477, c6478, c6479, 
	c6480, c6481, c6482, c6483, c6484, c6485, c6486, c6487, c6488, c6489, 
	c6490, c6491, c6492, c6493, c6494, c6495, c6496, c6497, c6498, c6499, 
	c6500, c6501, c6502, c6503, c6504, c6505, c6506, c6507, c6508, c6509, 
	c6510, c6511, c6512, c6513, c6514, c6515, c6516, c6517, c6518, c6519, 
	c6520, c6521, c6522, c6523, c6524, c6525, c6526, c6527, c6528, c6529, 
	c6530, c6531, c6532, c6533, c6534, c6535, c6536, c6537, c6538, c6539, 
	c6540, c6541, c6542, c6543, c6544, c6545, c6546, c6547, c6548, c6549, 
	c6550, c6551, c6552, c6553, c6554, c6555, c6556, c6557, c6558, c6559, 
	c6560, c6561, c6562, c6563, c6564, c6565, c6566, c6567, c6568, c6569, 
	c6570, c6571, c6572, c6573, c6574, c6575, c6576, c6577, c6578, c6579, 
	c6580, c6581, c6582, c6583, c6584, c6585, c6586, c6587, c6588, c6589, 
	c6590, c6591, c6592, c6593, c6594, c6595, c6596, c6597, c6598, c6599, 
	c6600, c6601, c6602, c6603, c6604, c6605, c6606, c6607, c6608, c6609, 
	c6610, c6611, c6612, c6613, c6614, c6615, c6616, c6617, c6618, c6619, 
	c6620, c6621, c6622, c6623, c6624, c6625, c6626, c6627, c6628, c6629, 
	c6630, c6631, c6632, c6633, c6634, c6635, c6636, c6637, c6638, c6639, 
	c6640, c6641, c6642, c6643, c6644, c6645, c6646, c6647, c6648, c6649, 
	c6650, c6651, c6652, c6653, c6654, c6655, c6656, c6657, c6658, c6659, 
	c6660, c6661, c6662, c6663, c6664, c6665, c6666, c6667, c6668, c6669, 
	c6670, c6671, c6672, c6673, c6674, c6675, c6676, c6677, c6678, c6679, 
	c6680, c6681, c6682, c6683, c6684, c6685, c6686, c6687, c6688, c6689, 
	c6690, c6691, c6692, c6693, c6694, c6695, c6696, c6697, c6698, c6699, 
	c6700, c6701, c6702, c6703, c6704, c6705, c6706, c6707, c6708, c6709, 
	c6710, c6711, c6712, c6713, c6714, c6715, c6716, c6717, c6718, c6719, 
	c6720, c6721, c6722, c6723, c6724, c6725, c6726, c6727, c6728, c6729, 
	c6730, c6731, c6732, c6733, c6734, c6735, c6736, c6737, c6738, c6739, 
	c6740, c6741, c6742, c6743, c6744, c6745, c6746, c6747, c6748, c6749, 
	c6750, c6751, c6752, c6753, c6754, c6755, c6756, c6757, c6758, c6759, 
	c6760, c6761, c6762, c6763, c6764, c6765, c6766, c6767, c6768, c6769, 
	c6770, c6771, c6772, c6773, c6774, c6775, c6776, c6777, c6778, c6779, 
	c6780, c6781, c6782, c6783, c6784, c6785, c6786, c6787, c6788, c6789, 
	c6790, c6791, c6792, c6793, c6794, c6795, c6796, c6797, c6798, c6799, 
	c6800, c6801, c6802, c6803, c6804, c6805, c6806, c6807, c6808, c6809, 
	c6810, c6811, c6812, c6813, c6814, c6815, c6816, c6817, c6818, c6819, 
	c6820, c6821, c6822, c6823, c6824, c6825, c6826, c6827, c6828, c6829, 
	c6830, c6831, c6832, c6833, c6834, c6835, c6836, c6837, c6838, c6839, 
	c6840, c6841, c6842, c6843, c6844, c6845, c6846, c6847, c6848, c6849, 
	c6850, c6851, c6852, c6853, c6854, c6855, c6856, c6857, c6858, c6859, 
	c6860, c6861, c6862, c6863, c6864, c6865, c6866, c6867, c6868, c6869, 
	c6870, c6871, c6872, c6873, c6874, c6875, c6876, c6877, c6878, c6879, 
	c6880, c6881, c6882, c6883, c6884, c6885, c6886, c6887, c6888, c6889, 
	c6890, c6891, c6892, c6893, c6894, c6895, c6896, c6897, c6898, c6899, 
	c6900, c6901, c6902, c6903, c6904, c6905, c6906, c6907, c6908, c6909, 
	c6910, c6911, c6912, c6913, c6914, c6915, c6916, c6917, c6918, c6919, 
	c6920, c6921, c6922, c6923, c6924, c6925, c6926, c6927, c6928, c6929, 
	c6930, c6931, c6932, c6933, c6934, c6935, c6936, c6937, c6938, c6939, 
	c6940, c6941, c6942, c6943, c6944, c6945, c6946, c6947, c6948, c6949, 
	c6950, c6951, c6952, c6953, c6954, c6955, c6956, c6957, c6958, c6959, 
	c6960, c6961, c6962, c6963, c6964, c6965, c6966, c6967, c6968, c6969, 
	c6970, c6971, c6972, c6973, c6974, c6975, c6976, c6977, c6978, c6979, 
	c6980, c6981, c6982, c6983, c6984, c6985, c6986, c6987, c6988, c6989, 
	c6990, c6991, c6992, c6993, c6994, c6995, c6996, c6997, c6998, c6999, 
	c7000, c7001, c7002, c7003, c7004, c7005, c7006, c7007, c7008, c7009, 
	c7010, c7011, c7012, c7013, c7014, c7015, c7016, c7017, c7018, c7019, 
	c7020, c7021, c7022, c7023, c7024, c7025, c7026, c7027, c7028, c7029, 
	c7030, c7031, c7032, c7033, c7034, c7035, c7036, c7037, c7038, c7039, 
	c7040, c7041, c7042, c7043, c7044, c7045, c7046, c7047, c7048, c7049, 
	c7050, c7051, c7052, c7053, c7054, c7055, c7056, c7057, c7058, c7059, 
	c7060, c7061, c7062, c7063, c7064, c7065, c7066, c7067, c7068, c7069, 
	c7070, c7071, c7072, c7073, c7074, c7075, c7076, c7077, c7078, c7079, 
	c7080, c7081, c7082, c7083, c7084, c7085, c7086, c7087, c7088, c7089, 
	c7090, c7091, c7092, c7093, c7094, c7095, c7096, c7097, c7098, c7099, 
	c7100, c7101, c7102, c7103, c7104, c7105, c7106, c7107, c7108, c7109, 
	c7110, c7111, c7112, c7113, c7114, c7115, c7116, c7117, c7118, c7119, 
	c7120, c7121, c7122, c7123, c7124, c7125, c7126, c7127, c7128, c7129, 
	c7130, c7131, c7132, c7133, c7134, c7135, c7136, c7137, c7138, c7139, 
	c7140, c7141, c7142, c7143, c7144, c7145, c7146, c7147, c7148, c7149, 
	c7150, c7151, c7152, c7153, c7154, c7155, c7156, c7157, c7158, c7159, 
	c7160, c7161, c7162, c7163, c7164, c7165, c7166, c7167, c7168, c7169, 
	c7170, c7171, c7172, c7173, c7174, c7175, c7176, c7177, c7178, c7179, 
	c7180, c7181, c7182, c7183, c7184, c7185, c7186, c7187, c7188, c7189, 
	c7190, c7191, c7192, c7193, c7194, c7195, c7196, c7197, c7198, c7199, 
	c7200, c7201, c7202, c7203, c7204, c7205, c7206, c7207, c7208, c7209, 
	c7210, c7211, c7212, c7213, c7214, c7215, c7216, c7217, c7218, c7219, 
	c7220, c7221, c7222, c7223, c7224, c7225, c7226, c7227, c7228, c7229, 
	c7230, c7231, c7232, c7233, c7234, c7235, c7236, c7237, c7238, c7239, 
	c7240, c7241, c7242, c7243, c7244, c7245, c7246, c7247, c7248, c7249, 
	c7250, c7251, c7252, c7253, c7254, c7255, c7256, c7257, c7258, c7259, 
	c7260, c7261, c7262, c7263, c7264, c7265, c7266, c7267, c7268, c7269, 
	c7270, c7271, c7272, c7273, c7274, c7275, c7276, c7277, c7278, c7279, 
	c7280, c7281, c7282, c7283, c7284, c7285, c7286, c7287, c7288, c7289, 
	c7290, c7291, c7292, c7293, c7294, c7295, c7296, c7297, c7298, c7299, 
	c7300, c7301, c7302, c7303, c7304, c7305, c7306, c7307, c7308, c7309, 
	c7310, c7311, c7312, c7313, c7314, c7315, c7316, c7317, c7318, c7319, 
	c7320, c7321, c7322, c7323, c7324, c7325, c7326, c7327, c7328, c7329, 
	c7330, c7331, c7332, c7333, c7334, c7335, c7336, c7337, c7338, c7339, 
	c7340, c7341, c7342, c7343, c7344, c7345, c7346, c7347, c7348, c7349, 
	c7350, c7351, c7352, c7353, c7354, c7355, c7356, c7357, c7358, c7359, 
	c7360, c7361, c7362, c7363, c7364, c7365, c7366, c7367, c7368, c7369, 
	c7370, c7371, c7372, c7373, c7374, c7375, c7376, c7377, c7378, c7379, 
	c7380, c7381, c7382, c7383, c7384, c7385, c7386, c7387, c7388, c7389, 
	c7390, c7391, c7392, c7393, c7394, c7395, c7396, c7397, c7398, c7399, 
	c7400, c7401, c7402, c7403, c7404, c7405, c7406, c7407, c7408, c7409, 
	c7410, c7411, c7412, c7413, c7414, c7415, c7416, c7417, c7418, c7419, 
	c7420, c7421, c7422, c7423, c7424, c7425, c7426, c7427, c7428, c7429, 
	c7430, c7431, c7432, c7433, c7434, c7435, c7436, c7437, c7438, c7439, 
	c7440, c7441, c7442, c7443, c7444, c7445, c7446, c7447, c7448, c7449, 
	c7450, c7451, c7452, c7453, c7454, c7455, c7456, c7457, c7458, c7459, 
	c7460, c7461, c7462, c7463, c7464, c7465, c7466, c7467, c7468, c7469, 
	c7470, c7471, c7472, c7473, c7474, c7475, c7476, c7477, c7478, c7479, 
	c7480, c7481, c7482, c7483, c7484, c7485, c7486, c7487, c7488, c7489, 
	c7490, c7491, c7492, c7493, c7494, c7495, c7496, c7497, c7498, c7499, 
	c7500, c7501, c7502, c7503, c7504, c7505, c7506, c7507, c7508, c7509, 
	c7510, c7511, c7512, c7513, c7514, c7515, c7516, c7517, c7518, c7519, 
	c7520, c7521, c7522, c7523, c7524, c7525, c7526, c7527, c7528, c7529, 
	c7530, c7531, c7532, c7533, c7534, c7535, c7536, c7537, c7538, c7539, 
	c7540, c7541, c7542, c7543, c7544, c7545, c7546, c7547, c7548, c7549, 
	c7550, c7551, c7552, c7553, c7554, c7555, c7556, c7557, c7558, c7559, 
	c7560, c7561, c7562, c7563, c7564, c7565, c7566, c7567, c7568, c7569, 
	c7570, c7571, c7572, c7573, c7574, c7575, c7576, c7577, c7578, c7579, 
	c7580, c7581, c7582, c7583, c7584, c7585, c7586, c7587, c7588, c7589, 
	c7590, c7591, c7592, c7593, c7594, c7595, c7596, c7597, c7598, c7599, 
	c7600, c7601, c7602, c7603, c7604, c7605, c7606, c7607, c7608, c7609, 
	c7610, c7611, c7612, c7613, c7614, c7615, c7616, c7617, c7618, c7619, 
	c7620, c7621, c7622, c7623, c7624, c7625, c7626, c7627, c7628, c7629, 
	c7630, c7631, c7632, c7633, c7634, c7635, c7636, c7637, c7638, c7639, 
	c7640, c7641, c7642, c7643, c7644, c7645, c7646, c7647, c7648, c7649, 
	c7650, c7651, c7652, c7653, c7654, c7655, c7656, c7657, c7658, c7659, 
	c7660, c7661, c7662, c7663, c7664, c7665, c7666, c7667, c7668, c7669, 
	c7670, c7671, c7672, c7673, c7674, c7675, c7676, c7677, c7678, c7679, 
	c7680, c7681, c7682, c7683, c7684, c7685, c7686, c7687, c7688, c7689, 
	c7690, c7691, c7692, c7693, c7694, c7695, c7696, c7697, c7698, c7699, 
	c7700, c7701, c7702, c7703, c7704, c7705, c7706, c7707, c7708, c7709, 
	c7710, c7711, c7712, c7713, c7714, c7715, c7716, c7717, c7718, c7719, 
	c7720, c7721, c7722, c7723, c7724, c7725, c7726, c7727, c7728, c7729, 
	c7730, c7731, c7732, c7733, c7734, c7735, c7736, c7737, c7738, c7739, 
	c7740, c7741, c7742, c7743, c7744, c7745, c7746, c7747, c7748, c7749, 
	c7750, c7751, c7752, c7753, c7754, c7755, c7756, c7757, c7758, c7759, 
	c7760, c7761, c7762, c7763, c7764, c7765, c7766, c7767, c7768, c7769, 
	c7770, c7771, c7772, c7773, c7774, c7775, c7776, c7777, c7778, c7779, 
	c7780, c7781, c7782, c7783, c7784, c7785, c7786, c7787, c7788, c7789, 
	c7790, c7791, c7792, c7793, c7794, c7795, c7796, c7797, c7798, c7799, 
	c7800, c7801, c7802, c7803, c7804, c7805, c7806, c7807, c7808, c7809, 
	c7810, c7811, c7812, c7813, c7814, c7815, c7816, c7817, c7818, c7819, 
	c7820, c7821, c7822, c7823, c7824, c7825, c7826, c7827, c7828, c7829, 
	c7830, c7831, c7832, c7833, c7834, c7835, c7836, c7837, c7838, c7839, 
	c7840, c7841, c7842, c7843, c7844, c7845, c7846, c7847, c7848, c7849, 
	c7850, c7851, c7852, c7853, c7854, c7855, c7856, c7857, c7858, c7859, 
	c7860, c7861, c7862, c7863, c7864, c7865, c7866, c7867, c7868, c7869, 
	c7870, c7871, c7872, c7873, c7874, c7875, c7876, c7877, c7878, c7879, 
	c7880, c7881, c7882, c7883, c7884, c7885, c7886, c7887, c7888, c7889, 
	c7890, c7891, c7892, c7893, c7894, c7895, c7896, c7897, c7898, c7899, 
	c7900, c7901, c7902, c7903, c7904, c7905, c7906, c7907, c7908, c7909, 
	c7910, c7911, c7912, c7913, c7914, c7915, c7916, c7917, c7918, c7919, 
	c7920, c7921, c7922, c7923, c7924, c7925, c7926, c7927, c7928, c7929, 
	c7930, c7931, c7932, c7933, c7934, c7935, c7936, c7937, c7938, c7939, 
	c7940, c7941, c7942, c7943, c7944, c7945, c7946, c7947, c7948, c7949, 
	c7950, c7951, c7952, c7953, c7954, c7955, c7956, c7957, c7958, c7959, 
	c7960, c7961, c7962, c7963, c7964, c7965, c7966, c7967, c7968, c7969, 
	c7970, c7971, c7972, c7973, c7974, c7975, c7976, c7977, c7978, c7979, 
	c7980, c7981, c7982, c7983, c7984, c7985, c7986, c7987, c7988, c7989, 
	c7990, c7991, c7992, c7993, c7994, c7995, c7996, c7997, c7998, c7999, 
	c8000, c8001, c8002, c8003, c8004, c8005, c8006, c8007, c8008, c8009, 
	c8010, c8011, c8012, c8013, c8014, c8015, c8016, c8017, c8018, c8019, 
	c8020, c8021, c8022, c8023, c8024, c8025, c8026, c8027, c8028, c8029, 
	c8030, c8031, c8032, c8033, c8034, c8035, c8036, c8037, c8038, c8039, 
	c8040, c8041, c8042, c8043, c8044, c8045, c8046, c8047, c8048, c8049, 
	c8050, c8051, c8052, c8053, c8054, c8055, c8056, c8057, c8058, c8059, 
	c8060, c8061, c8062, c8063, c8064, c8065, c8066, c8067, c8068, c8069, 
	c8070, c8071, c8072, c8073, c8074, c8075, c8076, c8077, c8078, c8079, 
	c8080, c8081, c8082, c8083, c8084, c8085, c8086, c8087, c8088, c8089, 
	c8090, c8091, c8092, c8093, c8094, c8095, c8096, c8097, c8098, c8099, 
	c8100, c8101, c8102, c8103, c8104, c8105, c8106, c8107, c8108, c8109, 
	c8110, c8111, c8112, c8113, c8114, c8115, c8116, c8117, c8118, c8119, 
	c8120, c8121, c8122, c8123, c8124, c8125, c8126, c8127, c8128, c8129, 
	c8130, c8131, c8132, c8133, c8134, c8135, c8136, c8137, c8138, c8139, 
	c8140, c8141, c8142, c8143, c8144, c8145, c8146, c8147, c8148, c8149, 
	c8150, c8151, c8152, c8153, c8154, c8155, c8156, c8157, c8158, c8159, 
	c8160, c8161, c8162, c8163, c8164, c8165, c8166, c8167, c8168, c8169, 
	c8170, c8171, c8172, c8173, c8174, c8175, c8176, c8177, c8178, c8179, 
	c8180, c8181, c8182, c8183, c8184, c8185, c8186, c8187, c8188, c8189, 
	c8190, c8191;

DFF carry_on_reg ( .D(c8191), .CLK(clk), .RST(rst), .Q(c0) );

XOR U0 ( .A(c0), .B(n0), .Z(c1) );
ANDN U1 ( .B(n1), .A(n2), .Z(n0) );
XOR U2 ( .A(c0), .B(b[0]), .Z(n1) );
XNOR U3 ( .A(b[0]), .B(n2), .Z(c[0]) );
XNOR U4 ( .A(a[0]), .B(c0), .Z(n2) );
XOR U5 ( .A(c1), .B(n3), .Z(c2) );
ANDN U6 ( .B(n4), .A(n5), .Z(n3) );
XOR U7 ( .A(c1), .B(b[1]), .Z(n4) );
XNOR U8 ( .A(b[1]), .B(n5), .Z(c[1]) );
XNOR U9 ( .A(a[1]), .B(c1), .Z(n5) );
XOR U10 ( .A(c2), .B(n6), .Z(c3) );
ANDN U11 ( .B(n7), .A(n8), .Z(n6) );
XOR U12 ( .A(c2), .B(b[2]), .Z(n7) );
XNOR U13 ( .A(b[2]), .B(n8), .Z(c[2]) );
XNOR U14 ( .A(a[2]), .B(c2), .Z(n8) );
XOR U15 ( .A(c3), .B(n9), .Z(c4) );
ANDN U16 ( .B(n10), .A(n11), .Z(n9) );
XOR U17 ( .A(c3), .B(b[3]), .Z(n10) );
XNOR U18 ( .A(b[3]), .B(n11), .Z(c[3]) );
XNOR U19 ( .A(a[3]), .B(c3), .Z(n11) );
XOR U20 ( .A(c4), .B(n12), .Z(c5) );
ANDN U21 ( .B(n13), .A(n14), .Z(n12) );
XOR U22 ( .A(c4), .B(b[4]), .Z(n13) );
XNOR U23 ( .A(b[4]), .B(n14), .Z(c[4]) );
XNOR U24 ( .A(a[4]), .B(c4), .Z(n14) );
XOR U25 ( .A(c5), .B(n15), .Z(c6) );
ANDN U26 ( .B(n16), .A(n17), .Z(n15) );
XOR U27 ( .A(c5), .B(b[5]), .Z(n16) );
XNOR U28 ( .A(b[5]), .B(n17), .Z(c[5]) );
XNOR U29 ( .A(a[5]), .B(c5), .Z(n17) );
XOR U30 ( .A(c6), .B(n18), .Z(c7) );
ANDN U31 ( .B(n19), .A(n20), .Z(n18) );
XOR U32 ( .A(c6), .B(b[6]), .Z(n19) );
XNOR U33 ( .A(b[6]), .B(n20), .Z(c[6]) );
XNOR U34 ( .A(a[6]), .B(c6), .Z(n20) );
XOR U35 ( .A(c7), .B(n21), .Z(c8) );
ANDN U36 ( .B(n22), .A(n23), .Z(n21) );
XOR U37 ( .A(c7), .B(b[7]), .Z(n22) );
XNOR U38 ( .A(b[7]), .B(n23), .Z(c[7]) );
XNOR U39 ( .A(a[7]), .B(c7), .Z(n23) );
XOR U40 ( .A(c8), .B(n24), .Z(c9) );
ANDN U41 ( .B(n25), .A(n26), .Z(n24) );
XOR U42 ( .A(c8), .B(b[8]), .Z(n25) );
XNOR U43 ( .A(b[8]), .B(n26), .Z(c[8]) );
XNOR U44 ( .A(a[8]), .B(c8), .Z(n26) );
XOR U45 ( .A(c9), .B(n27), .Z(c10) );
ANDN U46 ( .B(n28), .A(n29), .Z(n27) );
XOR U47 ( .A(c9), .B(b[9]), .Z(n28) );
XNOR U48 ( .A(b[9]), .B(n29), .Z(c[9]) );
XNOR U49 ( .A(a[9]), .B(c9), .Z(n29) );
XOR U50 ( .A(c10), .B(n30), .Z(c11) );
ANDN U51 ( .B(n31), .A(n32), .Z(n30) );
XOR U52 ( .A(c10), .B(b[10]), .Z(n31) );
XNOR U53 ( .A(b[10]), .B(n32), .Z(c[10]) );
XNOR U54 ( .A(a[10]), .B(c10), .Z(n32) );
XOR U55 ( .A(c11), .B(n33), .Z(c12) );
ANDN U56 ( .B(n34), .A(n35), .Z(n33) );
XOR U57 ( .A(c11), .B(b[11]), .Z(n34) );
XNOR U58 ( .A(b[11]), .B(n35), .Z(c[11]) );
XNOR U59 ( .A(a[11]), .B(c11), .Z(n35) );
XOR U60 ( .A(c12), .B(n36), .Z(c13) );
ANDN U61 ( .B(n37), .A(n38), .Z(n36) );
XOR U62 ( .A(c12), .B(b[12]), .Z(n37) );
XNOR U63 ( .A(b[12]), .B(n38), .Z(c[12]) );
XNOR U64 ( .A(a[12]), .B(c12), .Z(n38) );
XOR U65 ( .A(c13), .B(n39), .Z(c14) );
ANDN U66 ( .B(n40), .A(n41), .Z(n39) );
XOR U67 ( .A(c13), .B(b[13]), .Z(n40) );
XNOR U68 ( .A(b[13]), .B(n41), .Z(c[13]) );
XNOR U69 ( .A(a[13]), .B(c13), .Z(n41) );
XOR U70 ( .A(c14), .B(n42), .Z(c15) );
ANDN U71 ( .B(n43), .A(n44), .Z(n42) );
XOR U72 ( .A(c14), .B(b[14]), .Z(n43) );
XNOR U73 ( .A(b[14]), .B(n44), .Z(c[14]) );
XNOR U74 ( .A(a[14]), .B(c14), .Z(n44) );
XOR U75 ( .A(c15), .B(n45), .Z(c16) );
ANDN U76 ( .B(n46), .A(n47), .Z(n45) );
XOR U77 ( .A(c15), .B(b[15]), .Z(n46) );
XNOR U78 ( .A(b[15]), .B(n47), .Z(c[15]) );
XNOR U79 ( .A(a[15]), .B(c15), .Z(n47) );
XOR U80 ( .A(c16), .B(n48), .Z(c17) );
ANDN U81 ( .B(n49), .A(n50), .Z(n48) );
XOR U82 ( .A(c16), .B(b[16]), .Z(n49) );
XNOR U83 ( .A(b[16]), .B(n50), .Z(c[16]) );
XNOR U84 ( .A(a[16]), .B(c16), .Z(n50) );
XOR U85 ( .A(c17), .B(n51), .Z(c18) );
ANDN U86 ( .B(n52), .A(n53), .Z(n51) );
XOR U87 ( .A(c17), .B(b[17]), .Z(n52) );
XNOR U88 ( .A(b[17]), .B(n53), .Z(c[17]) );
XNOR U89 ( .A(a[17]), .B(c17), .Z(n53) );
XOR U90 ( .A(c18), .B(n54), .Z(c19) );
ANDN U91 ( .B(n55), .A(n56), .Z(n54) );
XOR U92 ( .A(c18), .B(b[18]), .Z(n55) );
XNOR U93 ( .A(b[18]), .B(n56), .Z(c[18]) );
XNOR U94 ( .A(a[18]), .B(c18), .Z(n56) );
XOR U95 ( .A(c19), .B(n57), .Z(c20) );
ANDN U96 ( .B(n58), .A(n59), .Z(n57) );
XOR U97 ( .A(c19), .B(b[19]), .Z(n58) );
XNOR U98 ( .A(b[19]), .B(n59), .Z(c[19]) );
XNOR U99 ( .A(a[19]), .B(c19), .Z(n59) );
XOR U100 ( .A(c20), .B(n60), .Z(c21) );
ANDN U101 ( .B(n61), .A(n62), .Z(n60) );
XOR U102 ( .A(c20), .B(b[20]), .Z(n61) );
XNOR U103 ( .A(b[20]), .B(n62), .Z(c[20]) );
XNOR U104 ( .A(a[20]), .B(c20), .Z(n62) );
XOR U105 ( .A(c21), .B(n63), .Z(c22) );
ANDN U106 ( .B(n64), .A(n65), .Z(n63) );
XOR U107 ( .A(c21), .B(b[21]), .Z(n64) );
XNOR U108 ( .A(b[21]), .B(n65), .Z(c[21]) );
XNOR U109 ( .A(a[21]), .B(c21), .Z(n65) );
XOR U110 ( .A(c22), .B(n66), .Z(c23) );
ANDN U111 ( .B(n67), .A(n68), .Z(n66) );
XOR U112 ( .A(c22), .B(b[22]), .Z(n67) );
XNOR U113 ( .A(b[22]), .B(n68), .Z(c[22]) );
XNOR U114 ( .A(a[22]), .B(c22), .Z(n68) );
XOR U115 ( .A(c23), .B(n69), .Z(c24) );
ANDN U116 ( .B(n70), .A(n71), .Z(n69) );
XOR U117 ( .A(c23), .B(b[23]), .Z(n70) );
XNOR U118 ( .A(b[23]), .B(n71), .Z(c[23]) );
XNOR U119 ( .A(a[23]), .B(c23), .Z(n71) );
XOR U120 ( .A(c24), .B(n72), .Z(c25) );
ANDN U121 ( .B(n73), .A(n74), .Z(n72) );
XOR U122 ( .A(c24), .B(b[24]), .Z(n73) );
XNOR U123 ( .A(b[24]), .B(n74), .Z(c[24]) );
XNOR U124 ( .A(a[24]), .B(c24), .Z(n74) );
XOR U125 ( .A(c25), .B(n75), .Z(c26) );
ANDN U126 ( .B(n76), .A(n77), .Z(n75) );
XOR U127 ( .A(c25), .B(b[25]), .Z(n76) );
XNOR U128 ( .A(b[25]), .B(n77), .Z(c[25]) );
XNOR U129 ( .A(a[25]), .B(c25), .Z(n77) );
XOR U130 ( .A(c26), .B(n78), .Z(c27) );
ANDN U131 ( .B(n79), .A(n80), .Z(n78) );
XOR U132 ( .A(c26), .B(b[26]), .Z(n79) );
XNOR U133 ( .A(b[26]), .B(n80), .Z(c[26]) );
XNOR U134 ( .A(a[26]), .B(c26), .Z(n80) );
XOR U135 ( .A(c27), .B(n81), .Z(c28) );
ANDN U136 ( .B(n82), .A(n83), .Z(n81) );
XOR U137 ( .A(c27), .B(b[27]), .Z(n82) );
XNOR U138 ( .A(b[27]), .B(n83), .Z(c[27]) );
XNOR U139 ( .A(a[27]), .B(c27), .Z(n83) );
XOR U140 ( .A(c28), .B(n84), .Z(c29) );
ANDN U141 ( .B(n85), .A(n86), .Z(n84) );
XOR U142 ( .A(c28), .B(b[28]), .Z(n85) );
XNOR U143 ( .A(b[28]), .B(n86), .Z(c[28]) );
XNOR U144 ( .A(a[28]), .B(c28), .Z(n86) );
XOR U145 ( .A(c29), .B(n87), .Z(c30) );
ANDN U146 ( .B(n88), .A(n89), .Z(n87) );
XOR U147 ( .A(c29), .B(b[29]), .Z(n88) );
XNOR U148 ( .A(b[29]), .B(n89), .Z(c[29]) );
XNOR U149 ( .A(a[29]), .B(c29), .Z(n89) );
XOR U150 ( .A(c30), .B(n90), .Z(c31) );
ANDN U151 ( .B(n91), .A(n92), .Z(n90) );
XOR U152 ( .A(c30), .B(b[30]), .Z(n91) );
XNOR U153 ( .A(b[30]), .B(n92), .Z(c[30]) );
XNOR U154 ( .A(a[30]), .B(c30), .Z(n92) );
XOR U155 ( .A(c31), .B(n93), .Z(c32) );
ANDN U156 ( .B(n94), .A(n95), .Z(n93) );
XOR U157 ( .A(c31), .B(b[31]), .Z(n94) );
XNOR U158 ( .A(b[31]), .B(n95), .Z(c[31]) );
XNOR U159 ( .A(a[31]), .B(c31), .Z(n95) );
XOR U160 ( .A(c32), .B(n96), .Z(c33) );
ANDN U161 ( .B(n97), .A(n98), .Z(n96) );
XOR U162 ( .A(c32), .B(b[32]), .Z(n97) );
XNOR U163 ( .A(b[32]), .B(n98), .Z(c[32]) );
XNOR U164 ( .A(a[32]), .B(c32), .Z(n98) );
XOR U165 ( .A(c33), .B(n99), .Z(c34) );
ANDN U166 ( .B(n100), .A(n101), .Z(n99) );
XOR U167 ( .A(c33), .B(b[33]), .Z(n100) );
XNOR U168 ( .A(b[33]), .B(n101), .Z(c[33]) );
XNOR U169 ( .A(a[33]), .B(c33), .Z(n101) );
XOR U170 ( .A(c34), .B(n102), .Z(c35) );
ANDN U171 ( .B(n103), .A(n104), .Z(n102) );
XOR U172 ( .A(c34), .B(b[34]), .Z(n103) );
XNOR U173 ( .A(b[34]), .B(n104), .Z(c[34]) );
XNOR U174 ( .A(a[34]), .B(c34), .Z(n104) );
XOR U175 ( .A(c35), .B(n105), .Z(c36) );
ANDN U176 ( .B(n106), .A(n107), .Z(n105) );
XOR U177 ( .A(c35), .B(b[35]), .Z(n106) );
XNOR U178 ( .A(b[35]), .B(n107), .Z(c[35]) );
XNOR U179 ( .A(a[35]), .B(c35), .Z(n107) );
XOR U180 ( .A(c36), .B(n108), .Z(c37) );
ANDN U181 ( .B(n109), .A(n110), .Z(n108) );
XOR U182 ( .A(c36), .B(b[36]), .Z(n109) );
XNOR U183 ( .A(b[36]), .B(n110), .Z(c[36]) );
XNOR U184 ( .A(a[36]), .B(c36), .Z(n110) );
XOR U185 ( .A(c37), .B(n111), .Z(c38) );
ANDN U186 ( .B(n112), .A(n113), .Z(n111) );
XOR U187 ( .A(c37), .B(b[37]), .Z(n112) );
XNOR U188 ( .A(b[37]), .B(n113), .Z(c[37]) );
XNOR U189 ( .A(a[37]), .B(c37), .Z(n113) );
XOR U190 ( .A(c38), .B(n114), .Z(c39) );
ANDN U191 ( .B(n115), .A(n116), .Z(n114) );
XOR U192 ( .A(c38), .B(b[38]), .Z(n115) );
XNOR U193 ( .A(b[38]), .B(n116), .Z(c[38]) );
XNOR U194 ( .A(a[38]), .B(c38), .Z(n116) );
XOR U195 ( .A(c39), .B(n117), .Z(c40) );
ANDN U196 ( .B(n118), .A(n119), .Z(n117) );
XOR U197 ( .A(c39), .B(b[39]), .Z(n118) );
XNOR U198 ( .A(b[39]), .B(n119), .Z(c[39]) );
XNOR U199 ( .A(a[39]), .B(c39), .Z(n119) );
XOR U200 ( .A(c40), .B(n120), .Z(c41) );
ANDN U201 ( .B(n121), .A(n122), .Z(n120) );
XOR U202 ( .A(c40), .B(b[40]), .Z(n121) );
XNOR U203 ( .A(b[40]), .B(n122), .Z(c[40]) );
XNOR U204 ( .A(a[40]), .B(c40), .Z(n122) );
XOR U205 ( .A(c41), .B(n123), .Z(c42) );
ANDN U206 ( .B(n124), .A(n125), .Z(n123) );
XOR U207 ( .A(c41), .B(b[41]), .Z(n124) );
XNOR U208 ( .A(b[41]), .B(n125), .Z(c[41]) );
XNOR U209 ( .A(a[41]), .B(c41), .Z(n125) );
XOR U210 ( .A(c42), .B(n126), .Z(c43) );
ANDN U211 ( .B(n127), .A(n128), .Z(n126) );
XOR U212 ( .A(c42), .B(b[42]), .Z(n127) );
XNOR U213 ( .A(b[42]), .B(n128), .Z(c[42]) );
XNOR U214 ( .A(a[42]), .B(c42), .Z(n128) );
XOR U215 ( .A(c43), .B(n129), .Z(c44) );
ANDN U216 ( .B(n130), .A(n131), .Z(n129) );
XOR U217 ( .A(c43), .B(b[43]), .Z(n130) );
XNOR U218 ( .A(b[43]), .B(n131), .Z(c[43]) );
XNOR U219 ( .A(a[43]), .B(c43), .Z(n131) );
XOR U220 ( .A(c44), .B(n132), .Z(c45) );
ANDN U221 ( .B(n133), .A(n134), .Z(n132) );
XOR U222 ( .A(c44), .B(b[44]), .Z(n133) );
XNOR U223 ( .A(b[44]), .B(n134), .Z(c[44]) );
XNOR U224 ( .A(a[44]), .B(c44), .Z(n134) );
XOR U225 ( .A(c45), .B(n135), .Z(c46) );
ANDN U226 ( .B(n136), .A(n137), .Z(n135) );
XOR U227 ( .A(c45), .B(b[45]), .Z(n136) );
XNOR U228 ( .A(b[45]), .B(n137), .Z(c[45]) );
XNOR U229 ( .A(a[45]), .B(c45), .Z(n137) );
XOR U230 ( .A(c46), .B(n138), .Z(c47) );
ANDN U231 ( .B(n139), .A(n140), .Z(n138) );
XOR U232 ( .A(c46), .B(b[46]), .Z(n139) );
XNOR U233 ( .A(b[46]), .B(n140), .Z(c[46]) );
XNOR U234 ( .A(a[46]), .B(c46), .Z(n140) );
XOR U235 ( .A(c47), .B(n141), .Z(c48) );
ANDN U236 ( .B(n142), .A(n143), .Z(n141) );
XOR U237 ( .A(c47), .B(b[47]), .Z(n142) );
XNOR U238 ( .A(b[47]), .B(n143), .Z(c[47]) );
XNOR U239 ( .A(a[47]), .B(c47), .Z(n143) );
XOR U240 ( .A(c48), .B(n144), .Z(c49) );
ANDN U241 ( .B(n145), .A(n146), .Z(n144) );
XOR U242 ( .A(c48), .B(b[48]), .Z(n145) );
XNOR U243 ( .A(b[48]), .B(n146), .Z(c[48]) );
XNOR U244 ( .A(a[48]), .B(c48), .Z(n146) );
XOR U245 ( .A(c49), .B(n147), .Z(c50) );
ANDN U246 ( .B(n148), .A(n149), .Z(n147) );
XOR U247 ( .A(c49), .B(b[49]), .Z(n148) );
XNOR U248 ( .A(b[49]), .B(n149), .Z(c[49]) );
XNOR U249 ( .A(a[49]), .B(c49), .Z(n149) );
XOR U250 ( .A(c50), .B(n150), .Z(c51) );
ANDN U251 ( .B(n151), .A(n152), .Z(n150) );
XOR U252 ( .A(c50), .B(b[50]), .Z(n151) );
XNOR U253 ( .A(b[50]), .B(n152), .Z(c[50]) );
XNOR U254 ( .A(a[50]), .B(c50), .Z(n152) );
XOR U255 ( .A(c51), .B(n153), .Z(c52) );
ANDN U256 ( .B(n154), .A(n155), .Z(n153) );
XOR U257 ( .A(c51), .B(b[51]), .Z(n154) );
XNOR U258 ( .A(b[51]), .B(n155), .Z(c[51]) );
XNOR U259 ( .A(a[51]), .B(c51), .Z(n155) );
XOR U260 ( .A(c52), .B(n156), .Z(c53) );
ANDN U261 ( .B(n157), .A(n158), .Z(n156) );
XOR U262 ( .A(c52), .B(b[52]), .Z(n157) );
XNOR U263 ( .A(b[52]), .B(n158), .Z(c[52]) );
XNOR U264 ( .A(a[52]), .B(c52), .Z(n158) );
XOR U265 ( .A(c53), .B(n159), .Z(c54) );
ANDN U266 ( .B(n160), .A(n161), .Z(n159) );
XOR U267 ( .A(c53), .B(b[53]), .Z(n160) );
XNOR U268 ( .A(b[53]), .B(n161), .Z(c[53]) );
XNOR U269 ( .A(a[53]), .B(c53), .Z(n161) );
XOR U270 ( .A(c54), .B(n162), .Z(c55) );
ANDN U271 ( .B(n163), .A(n164), .Z(n162) );
XOR U272 ( .A(c54), .B(b[54]), .Z(n163) );
XNOR U273 ( .A(b[54]), .B(n164), .Z(c[54]) );
XNOR U274 ( .A(a[54]), .B(c54), .Z(n164) );
XOR U275 ( .A(c55), .B(n165), .Z(c56) );
ANDN U276 ( .B(n166), .A(n167), .Z(n165) );
XOR U277 ( .A(c55), .B(b[55]), .Z(n166) );
XNOR U278 ( .A(b[55]), .B(n167), .Z(c[55]) );
XNOR U279 ( .A(a[55]), .B(c55), .Z(n167) );
XOR U280 ( .A(c56), .B(n168), .Z(c57) );
ANDN U281 ( .B(n169), .A(n170), .Z(n168) );
XOR U282 ( .A(c56), .B(b[56]), .Z(n169) );
XNOR U283 ( .A(b[56]), .B(n170), .Z(c[56]) );
XNOR U284 ( .A(a[56]), .B(c56), .Z(n170) );
XOR U285 ( .A(c57), .B(n171), .Z(c58) );
ANDN U286 ( .B(n172), .A(n173), .Z(n171) );
XOR U287 ( .A(c57), .B(b[57]), .Z(n172) );
XNOR U288 ( .A(b[57]), .B(n173), .Z(c[57]) );
XNOR U289 ( .A(a[57]), .B(c57), .Z(n173) );
XOR U290 ( .A(c58), .B(n174), .Z(c59) );
ANDN U291 ( .B(n175), .A(n176), .Z(n174) );
XOR U292 ( .A(c58), .B(b[58]), .Z(n175) );
XNOR U293 ( .A(b[58]), .B(n176), .Z(c[58]) );
XNOR U294 ( .A(a[58]), .B(c58), .Z(n176) );
XOR U295 ( .A(c59), .B(n177), .Z(c60) );
ANDN U296 ( .B(n178), .A(n179), .Z(n177) );
XOR U297 ( .A(c59), .B(b[59]), .Z(n178) );
XNOR U298 ( .A(b[59]), .B(n179), .Z(c[59]) );
XNOR U299 ( .A(a[59]), .B(c59), .Z(n179) );
XOR U300 ( .A(c60), .B(n180), .Z(c61) );
ANDN U301 ( .B(n181), .A(n182), .Z(n180) );
XOR U302 ( .A(c60), .B(b[60]), .Z(n181) );
XNOR U303 ( .A(b[60]), .B(n182), .Z(c[60]) );
XNOR U304 ( .A(a[60]), .B(c60), .Z(n182) );
XOR U305 ( .A(c61), .B(n183), .Z(c62) );
ANDN U306 ( .B(n184), .A(n185), .Z(n183) );
XOR U307 ( .A(c61), .B(b[61]), .Z(n184) );
XNOR U308 ( .A(b[61]), .B(n185), .Z(c[61]) );
XNOR U309 ( .A(a[61]), .B(c61), .Z(n185) );
XOR U310 ( .A(c62), .B(n186), .Z(c63) );
ANDN U311 ( .B(n187), .A(n188), .Z(n186) );
XOR U312 ( .A(c62), .B(b[62]), .Z(n187) );
XNOR U313 ( .A(b[62]), .B(n188), .Z(c[62]) );
XNOR U314 ( .A(a[62]), .B(c62), .Z(n188) );
XOR U315 ( .A(c63), .B(n189), .Z(c64) );
ANDN U316 ( .B(n190), .A(n191), .Z(n189) );
XOR U317 ( .A(c63), .B(b[63]), .Z(n190) );
XNOR U318 ( .A(b[63]), .B(n191), .Z(c[63]) );
XNOR U319 ( .A(a[63]), .B(c63), .Z(n191) );
XOR U320 ( .A(c64), .B(n192), .Z(c65) );
ANDN U321 ( .B(n193), .A(n194), .Z(n192) );
XOR U322 ( .A(c64), .B(b[64]), .Z(n193) );
XNOR U323 ( .A(b[64]), .B(n194), .Z(c[64]) );
XNOR U324 ( .A(a[64]), .B(c64), .Z(n194) );
XOR U325 ( .A(c65), .B(n195), .Z(c66) );
ANDN U326 ( .B(n196), .A(n197), .Z(n195) );
XOR U327 ( .A(c65), .B(b[65]), .Z(n196) );
XNOR U328 ( .A(b[65]), .B(n197), .Z(c[65]) );
XNOR U329 ( .A(a[65]), .B(c65), .Z(n197) );
XOR U330 ( .A(c66), .B(n198), .Z(c67) );
ANDN U331 ( .B(n199), .A(n200), .Z(n198) );
XOR U332 ( .A(c66), .B(b[66]), .Z(n199) );
XNOR U333 ( .A(b[66]), .B(n200), .Z(c[66]) );
XNOR U334 ( .A(a[66]), .B(c66), .Z(n200) );
XOR U335 ( .A(c67), .B(n201), .Z(c68) );
ANDN U336 ( .B(n202), .A(n203), .Z(n201) );
XOR U337 ( .A(c67), .B(b[67]), .Z(n202) );
XNOR U338 ( .A(b[67]), .B(n203), .Z(c[67]) );
XNOR U339 ( .A(a[67]), .B(c67), .Z(n203) );
XOR U340 ( .A(c68), .B(n204), .Z(c69) );
ANDN U341 ( .B(n205), .A(n206), .Z(n204) );
XOR U342 ( .A(c68), .B(b[68]), .Z(n205) );
XNOR U343 ( .A(b[68]), .B(n206), .Z(c[68]) );
XNOR U344 ( .A(a[68]), .B(c68), .Z(n206) );
XOR U345 ( .A(c69), .B(n207), .Z(c70) );
ANDN U346 ( .B(n208), .A(n209), .Z(n207) );
XOR U347 ( .A(c69), .B(b[69]), .Z(n208) );
XNOR U348 ( .A(b[69]), .B(n209), .Z(c[69]) );
XNOR U349 ( .A(a[69]), .B(c69), .Z(n209) );
XOR U350 ( .A(c70), .B(n210), .Z(c71) );
ANDN U351 ( .B(n211), .A(n212), .Z(n210) );
XOR U352 ( .A(c70), .B(b[70]), .Z(n211) );
XNOR U353 ( .A(b[70]), .B(n212), .Z(c[70]) );
XNOR U354 ( .A(a[70]), .B(c70), .Z(n212) );
XOR U355 ( .A(c71), .B(n213), .Z(c72) );
ANDN U356 ( .B(n214), .A(n215), .Z(n213) );
XOR U357 ( .A(c71), .B(b[71]), .Z(n214) );
XNOR U358 ( .A(b[71]), .B(n215), .Z(c[71]) );
XNOR U359 ( .A(a[71]), .B(c71), .Z(n215) );
XOR U360 ( .A(c72), .B(n216), .Z(c73) );
ANDN U361 ( .B(n217), .A(n218), .Z(n216) );
XOR U362 ( .A(c72), .B(b[72]), .Z(n217) );
XNOR U363 ( .A(b[72]), .B(n218), .Z(c[72]) );
XNOR U364 ( .A(a[72]), .B(c72), .Z(n218) );
XOR U365 ( .A(c73), .B(n219), .Z(c74) );
ANDN U366 ( .B(n220), .A(n221), .Z(n219) );
XOR U367 ( .A(c73), .B(b[73]), .Z(n220) );
XNOR U368 ( .A(b[73]), .B(n221), .Z(c[73]) );
XNOR U369 ( .A(a[73]), .B(c73), .Z(n221) );
XOR U370 ( .A(c74), .B(n222), .Z(c75) );
ANDN U371 ( .B(n223), .A(n224), .Z(n222) );
XOR U372 ( .A(c74), .B(b[74]), .Z(n223) );
XNOR U373 ( .A(b[74]), .B(n224), .Z(c[74]) );
XNOR U374 ( .A(a[74]), .B(c74), .Z(n224) );
XOR U375 ( .A(c75), .B(n225), .Z(c76) );
ANDN U376 ( .B(n226), .A(n227), .Z(n225) );
XOR U377 ( .A(c75), .B(b[75]), .Z(n226) );
XNOR U378 ( .A(b[75]), .B(n227), .Z(c[75]) );
XNOR U379 ( .A(a[75]), .B(c75), .Z(n227) );
XOR U380 ( .A(c76), .B(n228), .Z(c77) );
ANDN U381 ( .B(n229), .A(n230), .Z(n228) );
XOR U382 ( .A(c76), .B(b[76]), .Z(n229) );
XNOR U383 ( .A(b[76]), .B(n230), .Z(c[76]) );
XNOR U384 ( .A(a[76]), .B(c76), .Z(n230) );
XOR U385 ( .A(c77), .B(n231), .Z(c78) );
ANDN U386 ( .B(n232), .A(n233), .Z(n231) );
XOR U387 ( .A(c77), .B(b[77]), .Z(n232) );
XNOR U388 ( .A(b[77]), .B(n233), .Z(c[77]) );
XNOR U389 ( .A(a[77]), .B(c77), .Z(n233) );
XOR U390 ( .A(c78), .B(n234), .Z(c79) );
ANDN U391 ( .B(n235), .A(n236), .Z(n234) );
XOR U392 ( .A(c78), .B(b[78]), .Z(n235) );
XNOR U393 ( .A(b[78]), .B(n236), .Z(c[78]) );
XNOR U394 ( .A(a[78]), .B(c78), .Z(n236) );
XOR U395 ( .A(c79), .B(n237), .Z(c80) );
ANDN U396 ( .B(n238), .A(n239), .Z(n237) );
XOR U397 ( .A(c79), .B(b[79]), .Z(n238) );
XNOR U398 ( .A(b[79]), .B(n239), .Z(c[79]) );
XNOR U399 ( .A(a[79]), .B(c79), .Z(n239) );
XOR U400 ( .A(c80), .B(n240), .Z(c81) );
ANDN U401 ( .B(n241), .A(n242), .Z(n240) );
XOR U402 ( .A(c80), .B(b[80]), .Z(n241) );
XNOR U403 ( .A(b[80]), .B(n242), .Z(c[80]) );
XNOR U404 ( .A(a[80]), .B(c80), .Z(n242) );
XOR U405 ( .A(c81), .B(n243), .Z(c82) );
ANDN U406 ( .B(n244), .A(n245), .Z(n243) );
XOR U407 ( .A(c81), .B(b[81]), .Z(n244) );
XNOR U408 ( .A(b[81]), .B(n245), .Z(c[81]) );
XNOR U409 ( .A(a[81]), .B(c81), .Z(n245) );
XOR U410 ( .A(c82), .B(n246), .Z(c83) );
ANDN U411 ( .B(n247), .A(n248), .Z(n246) );
XOR U412 ( .A(c82), .B(b[82]), .Z(n247) );
XNOR U413 ( .A(b[82]), .B(n248), .Z(c[82]) );
XNOR U414 ( .A(a[82]), .B(c82), .Z(n248) );
XOR U415 ( .A(c83), .B(n249), .Z(c84) );
ANDN U416 ( .B(n250), .A(n251), .Z(n249) );
XOR U417 ( .A(c83), .B(b[83]), .Z(n250) );
XNOR U418 ( .A(b[83]), .B(n251), .Z(c[83]) );
XNOR U419 ( .A(a[83]), .B(c83), .Z(n251) );
XOR U420 ( .A(c84), .B(n252), .Z(c85) );
ANDN U421 ( .B(n253), .A(n254), .Z(n252) );
XOR U422 ( .A(c84), .B(b[84]), .Z(n253) );
XNOR U423 ( .A(b[84]), .B(n254), .Z(c[84]) );
XNOR U424 ( .A(a[84]), .B(c84), .Z(n254) );
XOR U425 ( .A(c85), .B(n255), .Z(c86) );
ANDN U426 ( .B(n256), .A(n257), .Z(n255) );
XOR U427 ( .A(c85), .B(b[85]), .Z(n256) );
XNOR U428 ( .A(b[85]), .B(n257), .Z(c[85]) );
XNOR U429 ( .A(a[85]), .B(c85), .Z(n257) );
XOR U430 ( .A(c86), .B(n258), .Z(c87) );
ANDN U431 ( .B(n259), .A(n260), .Z(n258) );
XOR U432 ( .A(c86), .B(b[86]), .Z(n259) );
XNOR U433 ( .A(b[86]), .B(n260), .Z(c[86]) );
XNOR U434 ( .A(a[86]), .B(c86), .Z(n260) );
XOR U435 ( .A(c87), .B(n261), .Z(c88) );
ANDN U436 ( .B(n262), .A(n263), .Z(n261) );
XOR U437 ( .A(c87), .B(b[87]), .Z(n262) );
XNOR U438 ( .A(b[87]), .B(n263), .Z(c[87]) );
XNOR U439 ( .A(a[87]), .B(c87), .Z(n263) );
XOR U440 ( .A(c88), .B(n264), .Z(c89) );
ANDN U441 ( .B(n265), .A(n266), .Z(n264) );
XOR U442 ( .A(c88), .B(b[88]), .Z(n265) );
XNOR U443 ( .A(b[88]), .B(n266), .Z(c[88]) );
XNOR U444 ( .A(a[88]), .B(c88), .Z(n266) );
XOR U445 ( .A(c89), .B(n267), .Z(c90) );
ANDN U446 ( .B(n268), .A(n269), .Z(n267) );
XOR U447 ( .A(c89), .B(b[89]), .Z(n268) );
XNOR U448 ( .A(b[89]), .B(n269), .Z(c[89]) );
XNOR U449 ( .A(a[89]), .B(c89), .Z(n269) );
XOR U450 ( .A(c90), .B(n270), .Z(c91) );
ANDN U451 ( .B(n271), .A(n272), .Z(n270) );
XOR U452 ( .A(c90), .B(b[90]), .Z(n271) );
XNOR U453 ( .A(b[90]), .B(n272), .Z(c[90]) );
XNOR U454 ( .A(a[90]), .B(c90), .Z(n272) );
XOR U455 ( .A(c91), .B(n273), .Z(c92) );
ANDN U456 ( .B(n274), .A(n275), .Z(n273) );
XOR U457 ( .A(c91), .B(b[91]), .Z(n274) );
XNOR U458 ( .A(b[91]), .B(n275), .Z(c[91]) );
XNOR U459 ( .A(a[91]), .B(c91), .Z(n275) );
XOR U460 ( .A(c92), .B(n276), .Z(c93) );
ANDN U461 ( .B(n277), .A(n278), .Z(n276) );
XOR U462 ( .A(c92), .B(b[92]), .Z(n277) );
XNOR U463 ( .A(b[92]), .B(n278), .Z(c[92]) );
XNOR U464 ( .A(a[92]), .B(c92), .Z(n278) );
XOR U465 ( .A(c93), .B(n279), .Z(c94) );
ANDN U466 ( .B(n280), .A(n281), .Z(n279) );
XOR U467 ( .A(c93), .B(b[93]), .Z(n280) );
XNOR U468 ( .A(b[93]), .B(n281), .Z(c[93]) );
XNOR U469 ( .A(a[93]), .B(c93), .Z(n281) );
XOR U470 ( .A(c94), .B(n282), .Z(c95) );
ANDN U471 ( .B(n283), .A(n284), .Z(n282) );
XOR U472 ( .A(c94), .B(b[94]), .Z(n283) );
XNOR U473 ( .A(b[94]), .B(n284), .Z(c[94]) );
XNOR U474 ( .A(a[94]), .B(c94), .Z(n284) );
XOR U475 ( .A(c95), .B(n285), .Z(c96) );
ANDN U476 ( .B(n286), .A(n287), .Z(n285) );
XOR U477 ( .A(c95), .B(b[95]), .Z(n286) );
XNOR U478 ( .A(b[95]), .B(n287), .Z(c[95]) );
XNOR U479 ( .A(a[95]), .B(c95), .Z(n287) );
XOR U480 ( .A(c96), .B(n288), .Z(c97) );
ANDN U481 ( .B(n289), .A(n290), .Z(n288) );
XOR U482 ( .A(c96), .B(b[96]), .Z(n289) );
XNOR U483 ( .A(b[96]), .B(n290), .Z(c[96]) );
XNOR U484 ( .A(a[96]), .B(c96), .Z(n290) );
XOR U485 ( .A(c97), .B(n291), .Z(c98) );
ANDN U486 ( .B(n292), .A(n293), .Z(n291) );
XOR U487 ( .A(c97), .B(b[97]), .Z(n292) );
XNOR U488 ( .A(b[97]), .B(n293), .Z(c[97]) );
XNOR U489 ( .A(a[97]), .B(c97), .Z(n293) );
XOR U490 ( .A(c98), .B(n294), .Z(c99) );
ANDN U491 ( .B(n295), .A(n296), .Z(n294) );
XOR U492 ( .A(c98), .B(b[98]), .Z(n295) );
XNOR U493 ( .A(b[98]), .B(n296), .Z(c[98]) );
XNOR U494 ( .A(a[98]), .B(c98), .Z(n296) );
XOR U495 ( .A(c99), .B(n297), .Z(c100) );
ANDN U496 ( .B(n298), .A(n299), .Z(n297) );
XOR U497 ( .A(c99), .B(b[99]), .Z(n298) );
XNOR U498 ( .A(b[99]), .B(n299), .Z(c[99]) );
XNOR U499 ( .A(a[99]), .B(c99), .Z(n299) );
XOR U500 ( .A(c100), .B(n300), .Z(c101) );
ANDN U501 ( .B(n301), .A(n302), .Z(n300) );
XOR U502 ( .A(c100), .B(b[100]), .Z(n301) );
XNOR U503 ( .A(b[100]), .B(n302), .Z(c[100]) );
XNOR U504 ( .A(a[100]), .B(c100), .Z(n302) );
XOR U505 ( .A(c101), .B(n303), .Z(c102) );
ANDN U506 ( .B(n304), .A(n305), .Z(n303) );
XOR U507 ( .A(c101), .B(b[101]), .Z(n304) );
XNOR U508 ( .A(b[101]), .B(n305), .Z(c[101]) );
XNOR U509 ( .A(a[101]), .B(c101), .Z(n305) );
XOR U510 ( .A(c102), .B(n306), .Z(c103) );
ANDN U511 ( .B(n307), .A(n308), .Z(n306) );
XOR U512 ( .A(c102), .B(b[102]), .Z(n307) );
XNOR U513 ( .A(b[102]), .B(n308), .Z(c[102]) );
XNOR U514 ( .A(a[102]), .B(c102), .Z(n308) );
XOR U515 ( .A(c103), .B(n309), .Z(c104) );
ANDN U516 ( .B(n310), .A(n311), .Z(n309) );
XOR U517 ( .A(c103), .B(b[103]), .Z(n310) );
XNOR U518 ( .A(b[103]), .B(n311), .Z(c[103]) );
XNOR U519 ( .A(a[103]), .B(c103), .Z(n311) );
XOR U520 ( .A(c104), .B(n312), .Z(c105) );
ANDN U521 ( .B(n313), .A(n314), .Z(n312) );
XOR U522 ( .A(c104), .B(b[104]), .Z(n313) );
XNOR U523 ( .A(b[104]), .B(n314), .Z(c[104]) );
XNOR U524 ( .A(a[104]), .B(c104), .Z(n314) );
XOR U525 ( .A(c105), .B(n315), .Z(c106) );
ANDN U526 ( .B(n316), .A(n317), .Z(n315) );
XOR U527 ( .A(c105), .B(b[105]), .Z(n316) );
XNOR U528 ( .A(b[105]), .B(n317), .Z(c[105]) );
XNOR U529 ( .A(a[105]), .B(c105), .Z(n317) );
XOR U530 ( .A(c106), .B(n318), .Z(c107) );
ANDN U531 ( .B(n319), .A(n320), .Z(n318) );
XOR U532 ( .A(c106), .B(b[106]), .Z(n319) );
XNOR U533 ( .A(b[106]), .B(n320), .Z(c[106]) );
XNOR U534 ( .A(a[106]), .B(c106), .Z(n320) );
XOR U535 ( .A(c107), .B(n321), .Z(c108) );
ANDN U536 ( .B(n322), .A(n323), .Z(n321) );
XOR U537 ( .A(c107), .B(b[107]), .Z(n322) );
XNOR U538 ( .A(b[107]), .B(n323), .Z(c[107]) );
XNOR U539 ( .A(a[107]), .B(c107), .Z(n323) );
XOR U540 ( .A(c108), .B(n324), .Z(c109) );
ANDN U541 ( .B(n325), .A(n326), .Z(n324) );
XOR U542 ( .A(c108), .B(b[108]), .Z(n325) );
XNOR U543 ( .A(b[108]), .B(n326), .Z(c[108]) );
XNOR U544 ( .A(a[108]), .B(c108), .Z(n326) );
XOR U545 ( .A(c109), .B(n327), .Z(c110) );
ANDN U546 ( .B(n328), .A(n329), .Z(n327) );
XOR U547 ( .A(c109), .B(b[109]), .Z(n328) );
XNOR U548 ( .A(b[109]), .B(n329), .Z(c[109]) );
XNOR U549 ( .A(a[109]), .B(c109), .Z(n329) );
XOR U550 ( .A(c110), .B(n330), .Z(c111) );
ANDN U551 ( .B(n331), .A(n332), .Z(n330) );
XOR U552 ( .A(c110), .B(b[110]), .Z(n331) );
XNOR U553 ( .A(b[110]), .B(n332), .Z(c[110]) );
XNOR U554 ( .A(a[110]), .B(c110), .Z(n332) );
XOR U555 ( .A(c111), .B(n333), .Z(c112) );
ANDN U556 ( .B(n334), .A(n335), .Z(n333) );
XOR U557 ( .A(c111), .B(b[111]), .Z(n334) );
XNOR U558 ( .A(b[111]), .B(n335), .Z(c[111]) );
XNOR U559 ( .A(a[111]), .B(c111), .Z(n335) );
XOR U560 ( .A(c112), .B(n336), .Z(c113) );
ANDN U561 ( .B(n337), .A(n338), .Z(n336) );
XOR U562 ( .A(c112), .B(b[112]), .Z(n337) );
XNOR U563 ( .A(b[112]), .B(n338), .Z(c[112]) );
XNOR U564 ( .A(a[112]), .B(c112), .Z(n338) );
XOR U565 ( .A(c113), .B(n339), .Z(c114) );
ANDN U566 ( .B(n340), .A(n341), .Z(n339) );
XOR U567 ( .A(c113), .B(b[113]), .Z(n340) );
XNOR U568 ( .A(b[113]), .B(n341), .Z(c[113]) );
XNOR U569 ( .A(a[113]), .B(c113), .Z(n341) );
XOR U570 ( .A(c114), .B(n342), .Z(c115) );
ANDN U571 ( .B(n343), .A(n344), .Z(n342) );
XOR U572 ( .A(c114), .B(b[114]), .Z(n343) );
XNOR U573 ( .A(b[114]), .B(n344), .Z(c[114]) );
XNOR U574 ( .A(a[114]), .B(c114), .Z(n344) );
XOR U575 ( .A(c115), .B(n345), .Z(c116) );
ANDN U576 ( .B(n346), .A(n347), .Z(n345) );
XOR U577 ( .A(c115), .B(b[115]), .Z(n346) );
XNOR U578 ( .A(b[115]), .B(n347), .Z(c[115]) );
XNOR U579 ( .A(a[115]), .B(c115), .Z(n347) );
XOR U580 ( .A(c116), .B(n348), .Z(c117) );
ANDN U581 ( .B(n349), .A(n350), .Z(n348) );
XOR U582 ( .A(c116), .B(b[116]), .Z(n349) );
XNOR U583 ( .A(b[116]), .B(n350), .Z(c[116]) );
XNOR U584 ( .A(a[116]), .B(c116), .Z(n350) );
XOR U585 ( .A(c117), .B(n351), .Z(c118) );
ANDN U586 ( .B(n352), .A(n353), .Z(n351) );
XOR U587 ( .A(c117), .B(b[117]), .Z(n352) );
XNOR U588 ( .A(b[117]), .B(n353), .Z(c[117]) );
XNOR U589 ( .A(a[117]), .B(c117), .Z(n353) );
XOR U590 ( .A(c118), .B(n354), .Z(c119) );
ANDN U591 ( .B(n355), .A(n356), .Z(n354) );
XOR U592 ( .A(c118), .B(b[118]), .Z(n355) );
XNOR U593 ( .A(b[118]), .B(n356), .Z(c[118]) );
XNOR U594 ( .A(a[118]), .B(c118), .Z(n356) );
XOR U595 ( .A(c119), .B(n357), .Z(c120) );
ANDN U596 ( .B(n358), .A(n359), .Z(n357) );
XOR U597 ( .A(c119), .B(b[119]), .Z(n358) );
XNOR U598 ( .A(b[119]), .B(n359), .Z(c[119]) );
XNOR U599 ( .A(a[119]), .B(c119), .Z(n359) );
XOR U600 ( .A(c120), .B(n360), .Z(c121) );
ANDN U601 ( .B(n361), .A(n362), .Z(n360) );
XOR U602 ( .A(c120), .B(b[120]), .Z(n361) );
XNOR U603 ( .A(b[120]), .B(n362), .Z(c[120]) );
XNOR U604 ( .A(a[120]), .B(c120), .Z(n362) );
XOR U605 ( .A(c121), .B(n363), .Z(c122) );
ANDN U606 ( .B(n364), .A(n365), .Z(n363) );
XOR U607 ( .A(c121), .B(b[121]), .Z(n364) );
XNOR U608 ( .A(b[121]), .B(n365), .Z(c[121]) );
XNOR U609 ( .A(a[121]), .B(c121), .Z(n365) );
XOR U610 ( .A(c122), .B(n366), .Z(c123) );
ANDN U611 ( .B(n367), .A(n368), .Z(n366) );
XOR U612 ( .A(c122), .B(b[122]), .Z(n367) );
XNOR U613 ( .A(b[122]), .B(n368), .Z(c[122]) );
XNOR U614 ( .A(a[122]), .B(c122), .Z(n368) );
XOR U615 ( .A(c123), .B(n369), .Z(c124) );
ANDN U616 ( .B(n370), .A(n371), .Z(n369) );
XOR U617 ( .A(c123), .B(b[123]), .Z(n370) );
XNOR U618 ( .A(b[123]), .B(n371), .Z(c[123]) );
XNOR U619 ( .A(a[123]), .B(c123), .Z(n371) );
XOR U620 ( .A(c124), .B(n372), .Z(c125) );
ANDN U621 ( .B(n373), .A(n374), .Z(n372) );
XOR U622 ( .A(c124), .B(b[124]), .Z(n373) );
XNOR U623 ( .A(b[124]), .B(n374), .Z(c[124]) );
XNOR U624 ( .A(a[124]), .B(c124), .Z(n374) );
XOR U625 ( .A(c125), .B(n375), .Z(c126) );
ANDN U626 ( .B(n376), .A(n377), .Z(n375) );
XOR U627 ( .A(c125), .B(b[125]), .Z(n376) );
XNOR U628 ( .A(b[125]), .B(n377), .Z(c[125]) );
XNOR U629 ( .A(a[125]), .B(c125), .Z(n377) );
XOR U630 ( .A(c126), .B(n378), .Z(c127) );
ANDN U631 ( .B(n379), .A(n380), .Z(n378) );
XOR U632 ( .A(c126), .B(b[126]), .Z(n379) );
XNOR U633 ( .A(b[126]), .B(n380), .Z(c[126]) );
XNOR U634 ( .A(a[126]), .B(c126), .Z(n380) );
XOR U635 ( .A(c127), .B(n381), .Z(c128) );
ANDN U636 ( .B(n382), .A(n383), .Z(n381) );
XOR U637 ( .A(c127), .B(b[127]), .Z(n382) );
XNOR U638 ( .A(b[127]), .B(n383), .Z(c[127]) );
XNOR U639 ( .A(a[127]), .B(c127), .Z(n383) );
XOR U640 ( .A(c128), .B(n384), .Z(c129) );
ANDN U641 ( .B(n385), .A(n386), .Z(n384) );
XOR U642 ( .A(c128), .B(b[128]), .Z(n385) );
XNOR U643 ( .A(b[128]), .B(n386), .Z(c[128]) );
XNOR U644 ( .A(a[128]), .B(c128), .Z(n386) );
XOR U645 ( .A(c129), .B(n387), .Z(c130) );
ANDN U646 ( .B(n388), .A(n389), .Z(n387) );
XOR U647 ( .A(c129), .B(b[129]), .Z(n388) );
XNOR U648 ( .A(b[129]), .B(n389), .Z(c[129]) );
XNOR U649 ( .A(a[129]), .B(c129), .Z(n389) );
XOR U650 ( .A(c130), .B(n390), .Z(c131) );
ANDN U651 ( .B(n391), .A(n392), .Z(n390) );
XOR U652 ( .A(c130), .B(b[130]), .Z(n391) );
XNOR U653 ( .A(b[130]), .B(n392), .Z(c[130]) );
XNOR U654 ( .A(a[130]), .B(c130), .Z(n392) );
XOR U655 ( .A(c131), .B(n393), .Z(c132) );
ANDN U656 ( .B(n394), .A(n395), .Z(n393) );
XOR U657 ( .A(c131), .B(b[131]), .Z(n394) );
XNOR U658 ( .A(b[131]), .B(n395), .Z(c[131]) );
XNOR U659 ( .A(a[131]), .B(c131), .Z(n395) );
XOR U660 ( .A(c132), .B(n396), .Z(c133) );
ANDN U661 ( .B(n397), .A(n398), .Z(n396) );
XOR U662 ( .A(c132), .B(b[132]), .Z(n397) );
XNOR U663 ( .A(b[132]), .B(n398), .Z(c[132]) );
XNOR U664 ( .A(a[132]), .B(c132), .Z(n398) );
XOR U665 ( .A(c133), .B(n399), .Z(c134) );
ANDN U666 ( .B(n400), .A(n401), .Z(n399) );
XOR U667 ( .A(c133), .B(b[133]), .Z(n400) );
XNOR U668 ( .A(b[133]), .B(n401), .Z(c[133]) );
XNOR U669 ( .A(a[133]), .B(c133), .Z(n401) );
XOR U670 ( .A(c134), .B(n402), .Z(c135) );
ANDN U671 ( .B(n403), .A(n404), .Z(n402) );
XOR U672 ( .A(c134), .B(b[134]), .Z(n403) );
XNOR U673 ( .A(b[134]), .B(n404), .Z(c[134]) );
XNOR U674 ( .A(a[134]), .B(c134), .Z(n404) );
XOR U675 ( .A(c135), .B(n405), .Z(c136) );
ANDN U676 ( .B(n406), .A(n407), .Z(n405) );
XOR U677 ( .A(c135), .B(b[135]), .Z(n406) );
XNOR U678 ( .A(b[135]), .B(n407), .Z(c[135]) );
XNOR U679 ( .A(a[135]), .B(c135), .Z(n407) );
XOR U680 ( .A(c136), .B(n408), .Z(c137) );
ANDN U681 ( .B(n409), .A(n410), .Z(n408) );
XOR U682 ( .A(c136), .B(b[136]), .Z(n409) );
XNOR U683 ( .A(b[136]), .B(n410), .Z(c[136]) );
XNOR U684 ( .A(a[136]), .B(c136), .Z(n410) );
XOR U685 ( .A(c137), .B(n411), .Z(c138) );
ANDN U686 ( .B(n412), .A(n413), .Z(n411) );
XOR U687 ( .A(c137), .B(b[137]), .Z(n412) );
XNOR U688 ( .A(b[137]), .B(n413), .Z(c[137]) );
XNOR U689 ( .A(a[137]), .B(c137), .Z(n413) );
XOR U690 ( .A(c138), .B(n414), .Z(c139) );
ANDN U691 ( .B(n415), .A(n416), .Z(n414) );
XOR U692 ( .A(c138), .B(b[138]), .Z(n415) );
XNOR U693 ( .A(b[138]), .B(n416), .Z(c[138]) );
XNOR U694 ( .A(a[138]), .B(c138), .Z(n416) );
XOR U695 ( .A(c139), .B(n417), .Z(c140) );
ANDN U696 ( .B(n418), .A(n419), .Z(n417) );
XOR U697 ( .A(c139), .B(b[139]), .Z(n418) );
XNOR U698 ( .A(b[139]), .B(n419), .Z(c[139]) );
XNOR U699 ( .A(a[139]), .B(c139), .Z(n419) );
XOR U700 ( .A(c140), .B(n420), .Z(c141) );
ANDN U701 ( .B(n421), .A(n422), .Z(n420) );
XOR U702 ( .A(c140), .B(b[140]), .Z(n421) );
XNOR U703 ( .A(b[140]), .B(n422), .Z(c[140]) );
XNOR U704 ( .A(a[140]), .B(c140), .Z(n422) );
XOR U705 ( .A(c141), .B(n423), .Z(c142) );
ANDN U706 ( .B(n424), .A(n425), .Z(n423) );
XOR U707 ( .A(c141), .B(b[141]), .Z(n424) );
XNOR U708 ( .A(b[141]), .B(n425), .Z(c[141]) );
XNOR U709 ( .A(a[141]), .B(c141), .Z(n425) );
XOR U710 ( .A(c142), .B(n426), .Z(c143) );
ANDN U711 ( .B(n427), .A(n428), .Z(n426) );
XOR U712 ( .A(c142), .B(b[142]), .Z(n427) );
XNOR U713 ( .A(b[142]), .B(n428), .Z(c[142]) );
XNOR U714 ( .A(a[142]), .B(c142), .Z(n428) );
XOR U715 ( .A(c143), .B(n429), .Z(c144) );
ANDN U716 ( .B(n430), .A(n431), .Z(n429) );
XOR U717 ( .A(c143), .B(b[143]), .Z(n430) );
XNOR U718 ( .A(b[143]), .B(n431), .Z(c[143]) );
XNOR U719 ( .A(a[143]), .B(c143), .Z(n431) );
XOR U720 ( .A(c144), .B(n432), .Z(c145) );
ANDN U721 ( .B(n433), .A(n434), .Z(n432) );
XOR U722 ( .A(c144), .B(b[144]), .Z(n433) );
XNOR U723 ( .A(b[144]), .B(n434), .Z(c[144]) );
XNOR U724 ( .A(a[144]), .B(c144), .Z(n434) );
XOR U725 ( .A(c145), .B(n435), .Z(c146) );
ANDN U726 ( .B(n436), .A(n437), .Z(n435) );
XOR U727 ( .A(c145), .B(b[145]), .Z(n436) );
XNOR U728 ( .A(b[145]), .B(n437), .Z(c[145]) );
XNOR U729 ( .A(a[145]), .B(c145), .Z(n437) );
XOR U730 ( .A(c146), .B(n438), .Z(c147) );
ANDN U731 ( .B(n439), .A(n440), .Z(n438) );
XOR U732 ( .A(c146), .B(b[146]), .Z(n439) );
XNOR U733 ( .A(b[146]), .B(n440), .Z(c[146]) );
XNOR U734 ( .A(a[146]), .B(c146), .Z(n440) );
XOR U735 ( .A(c147), .B(n441), .Z(c148) );
ANDN U736 ( .B(n442), .A(n443), .Z(n441) );
XOR U737 ( .A(c147), .B(b[147]), .Z(n442) );
XNOR U738 ( .A(b[147]), .B(n443), .Z(c[147]) );
XNOR U739 ( .A(a[147]), .B(c147), .Z(n443) );
XOR U740 ( .A(c148), .B(n444), .Z(c149) );
ANDN U741 ( .B(n445), .A(n446), .Z(n444) );
XOR U742 ( .A(c148), .B(b[148]), .Z(n445) );
XNOR U743 ( .A(b[148]), .B(n446), .Z(c[148]) );
XNOR U744 ( .A(a[148]), .B(c148), .Z(n446) );
XOR U745 ( .A(c149), .B(n447), .Z(c150) );
ANDN U746 ( .B(n448), .A(n449), .Z(n447) );
XOR U747 ( .A(c149), .B(b[149]), .Z(n448) );
XNOR U748 ( .A(b[149]), .B(n449), .Z(c[149]) );
XNOR U749 ( .A(a[149]), .B(c149), .Z(n449) );
XOR U750 ( .A(c150), .B(n450), .Z(c151) );
ANDN U751 ( .B(n451), .A(n452), .Z(n450) );
XOR U752 ( .A(c150), .B(b[150]), .Z(n451) );
XNOR U753 ( .A(b[150]), .B(n452), .Z(c[150]) );
XNOR U754 ( .A(a[150]), .B(c150), .Z(n452) );
XOR U755 ( .A(c151), .B(n453), .Z(c152) );
ANDN U756 ( .B(n454), .A(n455), .Z(n453) );
XOR U757 ( .A(c151), .B(b[151]), .Z(n454) );
XNOR U758 ( .A(b[151]), .B(n455), .Z(c[151]) );
XNOR U759 ( .A(a[151]), .B(c151), .Z(n455) );
XOR U760 ( .A(c152), .B(n456), .Z(c153) );
ANDN U761 ( .B(n457), .A(n458), .Z(n456) );
XOR U762 ( .A(c152), .B(b[152]), .Z(n457) );
XNOR U763 ( .A(b[152]), .B(n458), .Z(c[152]) );
XNOR U764 ( .A(a[152]), .B(c152), .Z(n458) );
XOR U765 ( .A(c153), .B(n459), .Z(c154) );
ANDN U766 ( .B(n460), .A(n461), .Z(n459) );
XOR U767 ( .A(c153), .B(b[153]), .Z(n460) );
XNOR U768 ( .A(b[153]), .B(n461), .Z(c[153]) );
XNOR U769 ( .A(a[153]), .B(c153), .Z(n461) );
XOR U770 ( .A(c154), .B(n462), .Z(c155) );
ANDN U771 ( .B(n463), .A(n464), .Z(n462) );
XOR U772 ( .A(c154), .B(b[154]), .Z(n463) );
XNOR U773 ( .A(b[154]), .B(n464), .Z(c[154]) );
XNOR U774 ( .A(a[154]), .B(c154), .Z(n464) );
XOR U775 ( .A(c155), .B(n465), .Z(c156) );
ANDN U776 ( .B(n466), .A(n467), .Z(n465) );
XOR U777 ( .A(c155), .B(b[155]), .Z(n466) );
XNOR U778 ( .A(b[155]), .B(n467), .Z(c[155]) );
XNOR U779 ( .A(a[155]), .B(c155), .Z(n467) );
XOR U780 ( .A(c156), .B(n468), .Z(c157) );
ANDN U781 ( .B(n469), .A(n470), .Z(n468) );
XOR U782 ( .A(c156), .B(b[156]), .Z(n469) );
XNOR U783 ( .A(b[156]), .B(n470), .Z(c[156]) );
XNOR U784 ( .A(a[156]), .B(c156), .Z(n470) );
XOR U785 ( .A(c157), .B(n471), .Z(c158) );
ANDN U786 ( .B(n472), .A(n473), .Z(n471) );
XOR U787 ( .A(c157), .B(b[157]), .Z(n472) );
XNOR U788 ( .A(b[157]), .B(n473), .Z(c[157]) );
XNOR U789 ( .A(a[157]), .B(c157), .Z(n473) );
XOR U790 ( .A(c158), .B(n474), .Z(c159) );
ANDN U791 ( .B(n475), .A(n476), .Z(n474) );
XOR U792 ( .A(c158), .B(b[158]), .Z(n475) );
XNOR U793 ( .A(b[158]), .B(n476), .Z(c[158]) );
XNOR U794 ( .A(a[158]), .B(c158), .Z(n476) );
XOR U795 ( .A(c159), .B(n477), .Z(c160) );
ANDN U796 ( .B(n478), .A(n479), .Z(n477) );
XOR U797 ( .A(c159), .B(b[159]), .Z(n478) );
XNOR U798 ( .A(b[159]), .B(n479), .Z(c[159]) );
XNOR U799 ( .A(a[159]), .B(c159), .Z(n479) );
XOR U800 ( .A(c160), .B(n480), .Z(c161) );
ANDN U801 ( .B(n481), .A(n482), .Z(n480) );
XOR U802 ( .A(c160), .B(b[160]), .Z(n481) );
XNOR U803 ( .A(b[160]), .B(n482), .Z(c[160]) );
XNOR U804 ( .A(a[160]), .B(c160), .Z(n482) );
XOR U805 ( .A(c161), .B(n483), .Z(c162) );
ANDN U806 ( .B(n484), .A(n485), .Z(n483) );
XOR U807 ( .A(c161), .B(b[161]), .Z(n484) );
XNOR U808 ( .A(b[161]), .B(n485), .Z(c[161]) );
XNOR U809 ( .A(a[161]), .B(c161), .Z(n485) );
XOR U810 ( .A(c162), .B(n486), .Z(c163) );
ANDN U811 ( .B(n487), .A(n488), .Z(n486) );
XOR U812 ( .A(c162), .B(b[162]), .Z(n487) );
XNOR U813 ( .A(b[162]), .B(n488), .Z(c[162]) );
XNOR U814 ( .A(a[162]), .B(c162), .Z(n488) );
XOR U815 ( .A(c163), .B(n489), .Z(c164) );
ANDN U816 ( .B(n490), .A(n491), .Z(n489) );
XOR U817 ( .A(c163), .B(b[163]), .Z(n490) );
XNOR U818 ( .A(b[163]), .B(n491), .Z(c[163]) );
XNOR U819 ( .A(a[163]), .B(c163), .Z(n491) );
XOR U820 ( .A(c164), .B(n492), .Z(c165) );
ANDN U821 ( .B(n493), .A(n494), .Z(n492) );
XOR U822 ( .A(c164), .B(b[164]), .Z(n493) );
XNOR U823 ( .A(b[164]), .B(n494), .Z(c[164]) );
XNOR U824 ( .A(a[164]), .B(c164), .Z(n494) );
XOR U825 ( .A(c165), .B(n495), .Z(c166) );
ANDN U826 ( .B(n496), .A(n497), .Z(n495) );
XOR U827 ( .A(c165), .B(b[165]), .Z(n496) );
XNOR U828 ( .A(b[165]), .B(n497), .Z(c[165]) );
XNOR U829 ( .A(a[165]), .B(c165), .Z(n497) );
XOR U830 ( .A(c166), .B(n498), .Z(c167) );
ANDN U831 ( .B(n499), .A(n500), .Z(n498) );
XOR U832 ( .A(c166), .B(b[166]), .Z(n499) );
XNOR U833 ( .A(b[166]), .B(n500), .Z(c[166]) );
XNOR U834 ( .A(a[166]), .B(c166), .Z(n500) );
XOR U835 ( .A(c167), .B(n501), .Z(c168) );
ANDN U836 ( .B(n502), .A(n503), .Z(n501) );
XOR U837 ( .A(c167), .B(b[167]), .Z(n502) );
XNOR U838 ( .A(b[167]), .B(n503), .Z(c[167]) );
XNOR U839 ( .A(a[167]), .B(c167), .Z(n503) );
XOR U840 ( .A(c168), .B(n504), .Z(c169) );
ANDN U841 ( .B(n505), .A(n506), .Z(n504) );
XOR U842 ( .A(c168), .B(b[168]), .Z(n505) );
XNOR U843 ( .A(b[168]), .B(n506), .Z(c[168]) );
XNOR U844 ( .A(a[168]), .B(c168), .Z(n506) );
XOR U845 ( .A(c169), .B(n507), .Z(c170) );
ANDN U846 ( .B(n508), .A(n509), .Z(n507) );
XOR U847 ( .A(c169), .B(b[169]), .Z(n508) );
XNOR U848 ( .A(b[169]), .B(n509), .Z(c[169]) );
XNOR U849 ( .A(a[169]), .B(c169), .Z(n509) );
XOR U850 ( .A(c170), .B(n510), .Z(c171) );
ANDN U851 ( .B(n511), .A(n512), .Z(n510) );
XOR U852 ( .A(c170), .B(b[170]), .Z(n511) );
XNOR U853 ( .A(b[170]), .B(n512), .Z(c[170]) );
XNOR U854 ( .A(a[170]), .B(c170), .Z(n512) );
XOR U855 ( .A(c171), .B(n513), .Z(c172) );
ANDN U856 ( .B(n514), .A(n515), .Z(n513) );
XOR U857 ( .A(c171), .B(b[171]), .Z(n514) );
XNOR U858 ( .A(b[171]), .B(n515), .Z(c[171]) );
XNOR U859 ( .A(a[171]), .B(c171), .Z(n515) );
XOR U860 ( .A(c172), .B(n516), .Z(c173) );
ANDN U861 ( .B(n517), .A(n518), .Z(n516) );
XOR U862 ( .A(c172), .B(b[172]), .Z(n517) );
XNOR U863 ( .A(b[172]), .B(n518), .Z(c[172]) );
XNOR U864 ( .A(a[172]), .B(c172), .Z(n518) );
XOR U865 ( .A(c173), .B(n519), .Z(c174) );
ANDN U866 ( .B(n520), .A(n521), .Z(n519) );
XOR U867 ( .A(c173), .B(b[173]), .Z(n520) );
XNOR U868 ( .A(b[173]), .B(n521), .Z(c[173]) );
XNOR U869 ( .A(a[173]), .B(c173), .Z(n521) );
XOR U870 ( .A(c174), .B(n522), .Z(c175) );
ANDN U871 ( .B(n523), .A(n524), .Z(n522) );
XOR U872 ( .A(c174), .B(b[174]), .Z(n523) );
XNOR U873 ( .A(b[174]), .B(n524), .Z(c[174]) );
XNOR U874 ( .A(a[174]), .B(c174), .Z(n524) );
XOR U875 ( .A(c175), .B(n525), .Z(c176) );
ANDN U876 ( .B(n526), .A(n527), .Z(n525) );
XOR U877 ( .A(c175), .B(b[175]), .Z(n526) );
XNOR U878 ( .A(b[175]), .B(n527), .Z(c[175]) );
XNOR U879 ( .A(a[175]), .B(c175), .Z(n527) );
XOR U880 ( .A(c176), .B(n528), .Z(c177) );
ANDN U881 ( .B(n529), .A(n530), .Z(n528) );
XOR U882 ( .A(c176), .B(b[176]), .Z(n529) );
XNOR U883 ( .A(b[176]), .B(n530), .Z(c[176]) );
XNOR U884 ( .A(a[176]), .B(c176), .Z(n530) );
XOR U885 ( .A(c177), .B(n531), .Z(c178) );
ANDN U886 ( .B(n532), .A(n533), .Z(n531) );
XOR U887 ( .A(c177), .B(b[177]), .Z(n532) );
XNOR U888 ( .A(b[177]), .B(n533), .Z(c[177]) );
XNOR U889 ( .A(a[177]), .B(c177), .Z(n533) );
XOR U890 ( .A(c178), .B(n534), .Z(c179) );
ANDN U891 ( .B(n535), .A(n536), .Z(n534) );
XOR U892 ( .A(c178), .B(b[178]), .Z(n535) );
XNOR U893 ( .A(b[178]), .B(n536), .Z(c[178]) );
XNOR U894 ( .A(a[178]), .B(c178), .Z(n536) );
XOR U895 ( .A(c179), .B(n537), .Z(c180) );
ANDN U896 ( .B(n538), .A(n539), .Z(n537) );
XOR U897 ( .A(c179), .B(b[179]), .Z(n538) );
XNOR U898 ( .A(b[179]), .B(n539), .Z(c[179]) );
XNOR U899 ( .A(a[179]), .B(c179), .Z(n539) );
XOR U900 ( .A(c180), .B(n540), .Z(c181) );
ANDN U901 ( .B(n541), .A(n542), .Z(n540) );
XOR U902 ( .A(c180), .B(b[180]), .Z(n541) );
XNOR U903 ( .A(b[180]), .B(n542), .Z(c[180]) );
XNOR U904 ( .A(a[180]), .B(c180), .Z(n542) );
XOR U905 ( .A(c181), .B(n543), .Z(c182) );
ANDN U906 ( .B(n544), .A(n545), .Z(n543) );
XOR U907 ( .A(c181), .B(b[181]), .Z(n544) );
XNOR U908 ( .A(b[181]), .B(n545), .Z(c[181]) );
XNOR U909 ( .A(a[181]), .B(c181), .Z(n545) );
XOR U910 ( .A(c182), .B(n546), .Z(c183) );
ANDN U911 ( .B(n547), .A(n548), .Z(n546) );
XOR U912 ( .A(c182), .B(b[182]), .Z(n547) );
XNOR U913 ( .A(b[182]), .B(n548), .Z(c[182]) );
XNOR U914 ( .A(a[182]), .B(c182), .Z(n548) );
XOR U915 ( .A(c183), .B(n549), .Z(c184) );
ANDN U916 ( .B(n550), .A(n551), .Z(n549) );
XOR U917 ( .A(c183), .B(b[183]), .Z(n550) );
XNOR U918 ( .A(b[183]), .B(n551), .Z(c[183]) );
XNOR U919 ( .A(a[183]), .B(c183), .Z(n551) );
XOR U920 ( .A(c184), .B(n552), .Z(c185) );
ANDN U921 ( .B(n553), .A(n554), .Z(n552) );
XOR U922 ( .A(c184), .B(b[184]), .Z(n553) );
XNOR U923 ( .A(b[184]), .B(n554), .Z(c[184]) );
XNOR U924 ( .A(a[184]), .B(c184), .Z(n554) );
XOR U925 ( .A(c185), .B(n555), .Z(c186) );
ANDN U926 ( .B(n556), .A(n557), .Z(n555) );
XOR U927 ( .A(c185), .B(b[185]), .Z(n556) );
XNOR U928 ( .A(b[185]), .B(n557), .Z(c[185]) );
XNOR U929 ( .A(a[185]), .B(c185), .Z(n557) );
XOR U930 ( .A(c186), .B(n558), .Z(c187) );
ANDN U931 ( .B(n559), .A(n560), .Z(n558) );
XOR U932 ( .A(c186), .B(b[186]), .Z(n559) );
XNOR U933 ( .A(b[186]), .B(n560), .Z(c[186]) );
XNOR U934 ( .A(a[186]), .B(c186), .Z(n560) );
XOR U935 ( .A(c187), .B(n561), .Z(c188) );
ANDN U936 ( .B(n562), .A(n563), .Z(n561) );
XOR U937 ( .A(c187), .B(b[187]), .Z(n562) );
XNOR U938 ( .A(b[187]), .B(n563), .Z(c[187]) );
XNOR U939 ( .A(a[187]), .B(c187), .Z(n563) );
XOR U940 ( .A(c188), .B(n564), .Z(c189) );
ANDN U941 ( .B(n565), .A(n566), .Z(n564) );
XOR U942 ( .A(c188), .B(b[188]), .Z(n565) );
XNOR U943 ( .A(b[188]), .B(n566), .Z(c[188]) );
XNOR U944 ( .A(a[188]), .B(c188), .Z(n566) );
XOR U945 ( .A(c189), .B(n567), .Z(c190) );
ANDN U946 ( .B(n568), .A(n569), .Z(n567) );
XOR U947 ( .A(c189), .B(b[189]), .Z(n568) );
XNOR U948 ( .A(b[189]), .B(n569), .Z(c[189]) );
XNOR U949 ( .A(a[189]), .B(c189), .Z(n569) );
XOR U950 ( .A(c190), .B(n570), .Z(c191) );
ANDN U951 ( .B(n571), .A(n572), .Z(n570) );
XOR U952 ( .A(c190), .B(b[190]), .Z(n571) );
XNOR U953 ( .A(b[190]), .B(n572), .Z(c[190]) );
XNOR U954 ( .A(a[190]), .B(c190), .Z(n572) );
XOR U955 ( .A(c191), .B(n573), .Z(c192) );
ANDN U956 ( .B(n574), .A(n575), .Z(n573) );
XOR U957 ( .A(c191), .B(b[191]), .Z(n574) );
XNOR U958 ( .A(b[191]), .B(n575), .Z(c[191]) );
XNOR U959 ( .A(a[191]), .B(c191), .Z(n575) );
XOR U960 ( .A(c192), .B(n576), .Z(c193) );
ANDN U961 ( .B(n577), .A(n578), .Z(n576) );
XOR U962 ( .A(c192), .B(b[192]), .Z(n577) );
XNOR U963 ( .A(b[192]), .B(n578), .Z(c[192]) );
XNOR U964 ( .A(a[192]), .B(c192), .Z(n578) );
XOR U965 ( .A(c193), .B(n579), .Z(c194) );
ANDN U966 ( .B(n580), .A(n581), .Z(n579) );
XOR U967 ( .A(c193), .B(b[193]), .Z(n580) );
XNOR U968 ( .A(b[193]), .B(n581), .Z(c[193]) );
XNOR U969 ( .A(a[193]), .B(c193), .Z(n581) );
XOR U970 ( .A(c194), .B(n582), .Z(c195) );
ANDN U971 ( .B(n583), .A(n584), .Z(n582) );
XOR U972 ( .A(c194), .B(b[194]), .Z(n583) );
XNOR U973 ( .A(b[194]), .B(n584), .Z(c[194]) );
XNOR U974 ( .A(a[194]), .B(c194), .Z(n584) );
XOR U975 ( .A(c195), .B(n585), .Z(c196) );
ANDN U976 ( .B(n586), .A(n587), .Z(n585) );
XOR U977 ( .A(c195), .B(b[195]), .Z(n586) );
XNOR U978 ( .A(b[195]), .B(n587), .Z(c[195]) );
XNOR U979 ( .A(a[195]), .B(c195), .Z(n587) );
XOR U980 ( .A(c196), .B(n588), .Z(c197) );
ANDN U981 ( .B(n589), .A(n590), .Z(n588) );
XOR U982 ( .A(c196), .B(b[196]), .Z(n589) );
XNOR U983 ( .A(b[196]), .B(n590), .Z(c[196]) );
XNOR U984 ( .A(a[196]), .B(c196), .Z(n590) );
XOR U985 ( .A(c197), .B(n591), .Z(c198) );
ANDN U986 ( .B(n592), .A(n593), .Z(n591) );
XOR U987 ( .A(c197), .B(b[197]), .Z(n592) );
XNOR U988 ( .A(b[197]), .B(n593), .Z(c[197]) );
XNOR U989 ( .A(a[197]), .B(c197), .Z(n593) );
XOR U990 ( .A(c198), .B(n594), .Z(c199) );
ANDN U991 ( .B(n595), .A(n596), .Z(n594) );
XOR U992 ( .A(c198), .B(b[198]), .Z(n595) );
XNOR U993 ( .A(b[198]), .B(n596), .Z(c[198]) );
XNOR U994 ( .A(a[198]), .B(c198), .Z(n596) );
XOR U995 ( .A(c199), .B(n597), .Z(c200) );
ANDN U996 ( .B(n598), .A(n599), .Z(n597) );
XOR U997 ( .A(c199), .B(b[199]), .Z(n598) );
XNOR U998 ( .A(b[199]), .B(n599), .Z(c[199]) );
XNOR U999 ( .A(a[199]), .B(c199), .Z(n599) );
XOR U1000 ( .A(c200), .B(n600), .Z(c201) );
ANDN U1001 ( .B(n601), .A(n602), .Z(n600) );
XOR U1002 ( .A(c200), .B(b[200]), .Z(n601) );
XNOR U1003 ( .A(b[200]), .B(n602), .Z(c[200]) );
XNOR U1004 ( .A(a[200]), .B(c200), .Z(n602) );
XOR U1005 ( .A(c201), .B(n603), .Z(c202) );
ANDN U1006 ( .B(n604), .A(n605), .Z(n603) );
XOR U1007 ( .A(c201), .B(b[201]), .Z(n604) );
XNOR U1008 ( .A(b[201]), .B(n605), .Z(c[201]) );
XNOR U1009 ( .A(a[201]), .B(c201), .Z(n605) );
XOR U1010 ( .A(c202), .B(n606), .Z(c203) );
ANDN U1011 ( .B(n607), .A(n608), .Z(n606) );
XOR U1012 ( .A(c202), .B(b[202]), .Z(n607) );
XNOR U1013 ( .A(b[202]), .B(n608), .Z(c[202]) );
XNOR U1014 ( .A(a[202]), .B(c202), .Z(n608) );
XOR U1015 ( .A(c203), .B(n609), .Z(c204) );
ANDN U1016 ( .B(n610), .A(n611), .Z(n609) );
XOR U1017 ( .A(c203), .B(b[203]), .Z(n610) );
XNOR U1018 ( .A(b[203]), .B(n611), .Z(c[203]) );
XNOR U1019 ( .A(a[203]), .B(c203), .Z(n611) );
XOR U1020 ( .A(c204), .B(n612), .Z(c205) );
ANDN U1021 ( .B(n613), .A(n614), .Z(n612) );
XOR U1022 ( .A(c204), .B(b[204]), .Z(n613) );
XNOR U1023 ( .A(b[204]), .B(n614), .Z(c[204]) );
XNOR U1024 ( .A(a[204]), .B(c204), .Z(n614) );
XOR U1025 ( .A(c205), .B(n615), .Z(c206) );
ANDN U1026 ( .B(n616), .A(n617), .Z(n615) );
XOR U1027 ( .A(c205), .B(b[205]), .Z(n616) );
XNOR U1028 ( .A(b[205]), .B(n617), .Z(c[205]) );
XNOR U1029 ( .A(a[205]), .B(c205), .Z(n617) );
XOR U1030 ( .A(c206), .B(n618), .Z(c207) );
ANDN U1031 ( .B(n619), .A(n620), .Z(n618) );
XOR U1032 ( .A(c206), .B(b[206]), .Z(n619) );
XNOR U1033 ( .A(b[206]), .B(n620), .Z(c[206]) );
XNOR U1034 ( .A(a[206]), .B(c206), .Z(n620) );
XOR U1035 ( .A(c207), .B(n621), .Z(c208) );
ANDN U1036 ( .B(n622), .A(n623), .Z(n621) );
XOR U1037 ( .A(c207), .B(b[207]), .Z(n622) );
XNOR U1038 ( .A(b[207]), .B(n623), .Z(c[207]) );
XNOR U1039 ( .A(a[207]), .B(c207), .Z(n623) );
XOR U1040 ( .A(c208), .B(n624), .Z(c209) );
ANDN U1041 ( .B(n625), .A(n626), .Z(n624) );
XOR U1042 ( .A(c208), .B(b[208]), .Z(n625) );
XNOR U1043 ( .A(b[208]), .B(n626), .Z(c[208]) );
XNOR U1044 ( .A(a[208]), .B(c208), .Z(n626) );
XOR U1045 ( .A(c209), .B(n627), .Z(c210) );
ANDN U1046 ( .B(n628), .A(n629), .Z(n627) );
XOR U1047 ( .A(c209), .B(b[209]), .Z(n628) );
XNOR U1048 ( .A(b[209]), .B(n629), .Z(c[209]) );
XNOR U1049 ( .A(a[209]), .B(c209), .Z(n629) );
XOR U1050 ( .A(c210), .B(n630), .Z(c211) );
ANDN U1051 ( .B(n631), .A(n632), .Z(n630) );
XOR U1052 ( .A(c210), .B(b[210]), .Z(n631) );
XNOR U1053 ( .A(b[210]), .B(n632), .Z(c[210]) );
XNOR U1054 ( .A(a[210]), .B(c210), .Z(n632) );
XOR U1055 ( .A(c211), .B(n633), .Z(c212) );
ANDN U1056 ( .B(n634), .A(n635), .Z(n633) );
XOR U1057 ( .A(c211), .B(b[211]), .Z(n634) );
XNOR U1058 ( .A(b[211]), .B(n635), .Z(c[211]) );
XNOR U1059 ( .A(a[211]), .B(c211), .Z(n635) );
XOR U1060 ( .A(c212), .B(n636), .Z(c213) );
ANDN U1061 ( .B(n637), .A(n638), .Z(n636) );
XOR U1062 ( .A(c212), .B(b[212]), .Z(n637) );
XNOR U1063 ( .A(b[212]), .B(n638), .Z(c[212]) );
XNOR U1064 ( .A(a[212]), .B(c212), .Z(n638) );
XOR U1065 ( .A(c213), .B(n639), .Z(c214) );
ANDN U1066 ( .B(n640), .A(n641), .Z(n639) );
XOR U1067 ( .A(c213), .B(b[213]), .Z(n640) );
XNOR U1068 ( .A(b[213]), .B(n641), .Z(c[213]) );
XNOR U1069 ( .A(a[213]), .B(c213), .Z(n641) );
XOR U1070 ( .A(c214), .B(n642), .Z(c215) );
ANDN U1071 ( .B(n643), .A(n644), .Z(n642) );
XOR U1072 ( .A(c214), .B(b[214]), .Z(n643) );
XNOR U1073 ( .A(b[214]), .B(n644), .Z(c[214]) );
XNOR U1074 ( .A(a[214]), .B(c214), .Z(n644) );
XOR U1075 ( .A(c215), .B(n645), .Z(c216) );
ANDN U1076 ( .B(n646), .A(n647), .Z(n645) );
XOR U1077 ( .A(c215), .B(b[215]), .Z(n646) );
XNOR U1078 ( .A(b[215]), .B(n647), .Z(c[215]) );
XNOR U1079 ( .A(a[215]), .B(c215), .Z(n647) );
XOR U1080 ( .A(c216), .B(n648), .Z(c217) );
ANDN U1081 ( .B(n649), .A(n650), .Z(n648) );
XOR U1082 ( .A(c216), .B(b[216]), .Z(n649) );
XNOR U1083 ( .A(b[216]), .B(n650), .Z(c[216]) );
XNOR U1084 ( .A(a[216]), .B(c216), .Z(n650) );
XOR U1085 ( .A(c217), .B(n651), .Z(c218) );
ANDN U1086 ( .B(n652), .A(n653), .Z(n651) );
XOR U1087 ( .A(c217), .B(b[217]), .Z(n652) );
XNOR U1088 ( .A(b[217]), .B(n653), .Z(c[217]) );
XNOR U1089 ( .A(a[217]), .B(c217), .Z(n653) );
XOR U1090 ( .A(c218), .B(n654), .Z(c219) );
ANDN U1091 ( .B(n655), .A(n656), .Z(n654) );
XOR U1092 ( .A(c218), .B(b[218]), .Z(n655) );
XNOR U1093 ( .A(b[218]), .B(n656), .Z(c[218]) );
XNOR U1094 ( .A(a[218]), .B(c218), .Z(n656) );
XOR U1095 ( .A(c219), .B(n657), .Z(c220) );
ANDN U1096 ( .B(n658), .A(n659), .Z(n657) );
XOR U1097 ( .A(c219), .B(b[219]), .Z(n658) );
XNOR U1098 ( .A(b[219]), .B(n659), .Z(c[219]) );
XNOR U1099 ( .A(a[219]), .B(c219), .Z(n659) );
XOR U1100 ( .A(c220), .B(n660), .Z(c221) );
ANDN U1101 ( .B(n661), .A(n662), .Z(n660) );
XOR U1102 ( .A(c220), .B(b[220]), .Z(n661) );
XNOR U1103 ( .A(b[220]), .B(n662), .Z(c[220]) );
XNOR U1104 ( .A(a[220]), .B(c220), .Z(n662) );
XOR U1105 ( .A(c221), .B(n663), .Z(c222) );
ANDN U1106 ( .B(n664), .A(n665), .Z(n663) );
XOR U1107 ( .A(c221), .B(b[221]), .Z(n664) );
XNOR U1108 ( .A(b[221]), .B(n665), .Z(c[221]) );
XNOR U1109 ( .A(a[221]), .B(c221), .Z(n665) );
XOR U1110 ( .A(c222), .B(n666), .Z(c223) );
ANDN U1111 ( .B(n667), .A(n668), .Z(n666) );
XOR U1112 ( .A(c222), .B(b[222]), .Z(n667) );
XNOR U1113 ( .A(b[222]), .B(n668), .Z(c[222]) );
XNOR U1114 ( .A(a[222]), .B(c222), .Z(n668) );
XOR U1115 ( .A(c223), .B(n669), .Z(c224) );
ANDN U1116 ( .B(n670), .A(n671), .Z(n669) );
XOR U1117 ( .A(c223), .B(b[223]), .Z(n670) );
XNOR U1118 ( .A(b[223]), .B(n671), .Z(c[223]) );
XNOR U1119 ( .A(a[223]), .B(c223), .Z(n671) );
XOR U1120 ( .A(c224), .B(n672), .Z(c225) );
ANDN U1121 ( .B(n673), .A(n674), .Z(n672) );
XOR U1122 ( .A(c224), .B(b[224]), .Z(n673) );
XNOR U1123 ( .A(b[224]), .B(n674), .Z(c[224]) );
XNOR U1124 ( .A(a[224]), .B(c224), .Z(n674) );
XOR U1125 ( .A(c225), .B(n675), .Z(c226) );
ANDN U1126 ( .B(n676), .A(n677), .Z(n675) );
XOR U1127 ( .A(c225), .B(b[225]), .Z(n676) );
XNOR U1128 ( .A(b[225]), .B(n677), .Z(c[225]) );
XNOR U1129 ( .A(a[225]), .B(c225), .Z(n677) );
XOR U1130 ( .A(c226), .B(n678), .Z(c227) );
ANDN U1131 ( .B(n679), .A(n680), .Z(n678) );
XOR U1132 ( .A(c226), .B(b[226]), .Z(n679) );
XNOR U1133 ( .A(b[226]), .B(n680), .Z(c[226]) );
XNOR U1134 ( .A(a[226]), .B(c226), .Z(n680) );
XOR U1135 ( .A(c227), .B(n681), .Z(c228) );
ANDN U1136 ( .B(n682), .A(n683), .Z(n681) );
XOR U1137 ( .A(c227), .B(b[227]), .Z(n682) );
XNOR U1138 ( .A(b[227]), .B(n683), .Z(c[227]) );
XNOR U1139 ( .A(a[227]), .B(c227), .Z(n683) );
XOR U1140 ( .A(c228), .B(n684), .Z(c229) );
ANDN U1141 ( .B(n685), .A(n686), .Z(n684) );
XOR U1142 ( .A(c228), .B(b[228]), .Z(n685) );
XNOR U1143 ( .A(b[228]), .B(n686), .Z(c[228]) );
XNOR U1144 ( .A(a[228]), .B(c228), .Z(n686) );
XOR U1145 ( .A(c229), .B(n687), .Z(c230) );
ANDN U1146 ( .B(n688), .A(n689), .Z(n687) );
XOR U1147 ( .A(c229), .B(b[229]), .Z(n688) );
XNOR U1148 ( .A(b[229]), .B(n689), .Z(c[229]) );
XNOR U1149 ( .A(a[229]), .B(c229), .Z(n689) );
XOR U1150 ( .A(c230), .B(n690), .Z(c231) );
ANDN U1151 ( .B(n691), .A(n692), .Z(n690) );
XOR U1152 ( .A(c230), .B(b[230]), .Z(n691) );
XNOR U1153 ( .A(b[230]), .B(n692), .Z(c[230]) );
XNOR U1154 ( .A(a[230]), .B(c230), .Z(n692) );
XOR U1155 ( .A(c231), .B(n693), .Z(c232) );
ANDN U1156 ( .B(n694), .A(n695), .Z(n693) );
XOR U1157 ( .A(c231), .B(b[231]), .Z(n694) );
XNOR U1158 ( .A(b[231]), .B(n695), .Z(c[231]) );
XNOR U1159 ( .A(a[231]), .B(c231), .Z(n695) );
XOR U1160 ( .A(c232), .B(n696), .Z(c233) );
ANDN U1161 ( .B(n697), .A(n698), .Z(n696) );
XOR U1162 ( .A(c232), .B(b[232]), .Z(n697) );
XNOR U1163 ( .A(b[232]), .B(n698), .Z(c[232]) );
XNOR U1164 ( .A(a[232]), .B(c232), .Z(n698) );
XOR U1165 ( .A(c233), .B(n699), .Z(c234) );
ANDN U1166 ( .B(n700), .A(n701), .Z(n699) );
XOR U1167 ( .A(c233), .B(b[233]), .Z(n700) );
XNOR U1168 ( .A(b[233]), .B(n701), .Z(c[233]) );
XNOR U1169 ( .A(a[233]), .B(c233), .Z(n701) );
XOR U1170 ( .A(c234), .B(n702), .Z(c235) );
ANDN U1171 ( .B(n703), .A(n704), .Z(n702) );
XOR U1172 ( .A(c234), .B(b[234]), .Z(n703) );
XNOR U1173 ( .A(b[234]), .B(n704), .Z(c[234]) );
XNOR U1174 ( .A(a[234]), .B(c234), .Z(n704) );
XOR U1175 ( .A(c235), .B(n705), .Z(c236) );
ANDN U1176 ( .B(n706), .A(n707), .Z(n705) );
XOR U1177 ( .A(c235), .B(b[235]), .Z(n706) );
XNOR U1178 ( .A(b[235]), .B(n707), .Z(c[235]) );
XNOR U1179 ( .A(a[235]), .B(c235), .Z(n707) );
XOR U1180 ( .A(c236), .B(n708), .Z(c237) );
ANDN U1181 ( .B(n709), .A(n710), .Z(n708) );
XOR U1182 ( .A(c236), .B(b[236]), .Z(n709) );
XNOR U1183 ( .A(b[236]), .B(n710), .Z(c[236]) );
XNOR U1184 ( .A(a[236]), .B(c236), .Z(n710) );
XOR U1185 ( .A(c237), .B(n711), .Z(c238) );
ANDN U1186 ( .B(n712), .A(n713), .Z(n711) );
XOR U1187 ( .A(c237), .B(b[237]), .Z(n712) );
XNOR U1188 ( .A(b[237]), .B(n713), .Z(c[237]) );
XNOR U1189 ( .A(a[237]), .B(c237), .Z(n713) );
XOR U1190 ( .A(c238), .B(n714), .Z(c239) );
ANDN U1191 ( .B(n715), .A(n716), .Z(n714) );
XOR U1192 ( .A(c238), .B(b[238]), .Z(n715) );
XNOR U1193 ( .A(b[238]), .B(n716), .Z(c[238]) );
XNOR U1194 ( .A(a[238]), .B(c238), .Z(n716) );
XOR U1195 ( .A(c239), .B(n717), .Z(c240) );
ANDN U1196 ( .B(n718), .A(n719), .Z(n717) );
XOR U1197 ( .A(c239), .B(b[239]), .Z(n718) );
XNOR U1198 ( .A(b[239]), .B(n719), .Z(c[239]) );
XNOR U1199 ( .A(a[239]), .B(c239), .Z(n719) );
XOR U1200 ( .A(c240), .B(n720), .Z(c241) );
ANDN U1201 ( .B(n721), .A(n722), .Z(n720) );
XOR U1202 ( .A(c240), .B(b[240]), .Z(n721) );
XNOR U1203 ( .A(b[240]), .B(n722), .Z(c[240]) );
XNOR U1204 ( .A(a[240]), .B(c240), .Z(n722) );
XOR U1205 ( .A(c241), .B(n723), .Z(c242) );
ANDN U1206 ( .B(n724), .A(n725), .Z(n723) );
XOR U1207 ( .A(c241), .B(b[241]), .Z(n724) );
XNOR U1208 ( .A(b[241]), .B(n725), .Z(c[241]) );
XNOR U1209 ( .A(a[241]), .B(c241), .Z(n725) );
XOR U1210 ( .A(c242), .B(n726), .Z(c243) );
ANDN U1211 ( .B(n727), .A(n728), .Z(n726) );
XOR U1212 ( .A(c242), .B(b[242]), .Z(n727) );
XNOR U1213 ( .A(b[242]), .B(n728), .Z(c[242]) );
XNOR U1214 ( .A(a[242]), .B(c242), .Z(n728) );
XOR U1215 ( .A(c243), .B(n729), .Z(c244) );
ANDN U1216 ( .B(n730), .A(n731), .Z(n729) );
XOR U1217 ( .A(c243), .B(b[243]), .Z(n730) );
XNOR U1218 ( .A(b[243]), .B(n731), .Z(c[243]) );
XNOR U1219 ( .A(a[243]), .B(c243), .Z(n731) );
XOR U1220 ( .A(c244), .B(n732), .Z(c245) );
ANDN U1221 ( .B(n733), .A(n734), .Z(n732) );
XOR U1222 ( .A(c244), .B(b[244]), .Z(n733) );
XNOR U1223 ( .A(b[244]), .B(n734), .Z(c[244]) );
XNOR U1224 ( .A(a[244]), .B(c244), .Z(n734) );
XOR U1225 ( .A(c245), .B(n735), .Z(c246) );
ANDN U1226 ( .B(n736), .A(n737), .Z(n735) );
XOR U1227 ( .A(c245), .B(b[245]), .Z(n736) );
XNOR U1228 ( .A(b[245]), .B(n737), .Z(c[245]) );
XNOR U1229 ( .A(a[245]), .B(c245), .Z(n737) );
XOR U1230 ( .A(c246), .B(n738), .Z(c247) );
ANDN U1231 ( .B(n739), .A(n740), .Z(n738) );
XOR U1232 ( .A(c246), .B(b[246]), .Z(n739) );
XNOR U1233 ( .A(b[246]), .B(n740), .Z(c[246]) );
XNOR U1234 ( .A(a[246]), .B(c246), .Z(n740) );
XOR U1235 ( .A(c247), .B(n741), .Z(c248) );
ANDN U1236 ( .B(n742), .A(n743), .Z(n741) );
XOR U1237 ( .A(c247), .B(b[247]), .Z(n742) );
XNOR U1238 ( .A(b[247]), .B(n743), .Z(c[247]) );
XNOR U1239 ( .A(a[247]), .B(c247), .Z(n743) );
XOR U1240 ( .A(c248), .B(n744), .Z(c249) );
ANDN U1241 ( .B(n745), .A(n746), .Z(n744) );
XOR U1242 ( .A(c248), .B(b[248]), .Z(n745) );
XNOR U1243 ( .A(b[248]), .B(n746), .Z(c[248]) );
XNOR U1244 ( .A(a[248]), .B(c248), .Z(n746) );
XOR U1245 ( .A(c249), .B(n747), .Z(c250) );
ANDN U1246 ( .B(n748), .A(n749), .Z(n747) );
XOR U1247 ( .A(c249), .B(b[249]), .Z(n748) );
XNOR U1248 ( .A(b[249]), .B(n749), .Z(c[249]) );
XNOR U1249 ( .A(a[249]), .B(c249), .Z(n749) );
XOR U1250 ( .A(c250), .B(n750), .Z(c251) );
ANDN U1251 ( .B(n751), .A(n752), .Z(n750) );
XOR U1252 ( .A(c250), .B(b[250]), .Z(n751) );
XNOR U1253 ( .A(b[250]), .B(n752), .Z(c[250]) );
XNOR U1254 ( .A(a[250]), .B(c250), .Z(n752) );
XOR U1255 ( .A(c251), .B(n753), .Z(c252) );
ANDN U1256 ( .B(n754), .A(n755), .Z(n753) );
XOR U1257 ( .A(c251), .B(b[251]), .Z(n754) );
XNOR U1258 ( .A(b[251]), .B(n755), .Z(c[251]) );
XNOR U1259 ( .A(a[251]), .B(c251), .Z(n755) );
XOR U1260 ( .A(c252), .B(n756), .Z(c253) );
ANDN U1261 ( .B(n757), .A(n758), .Z(n756) );
XOR U1262 ( .A(c252), .B(b[252]), .Z(n757) );
XNOR U1263 ( .A(b[252]), .B(n758), .Z(c[252]) );
XNOR U1264 ( .A(a[252]), .B(c252), .Z(n758) );
XOR U1265 ( .A(c253), .B(n759), .Z(c254) );
ANDN U1266 ( .B(n760), .A(n761), .Z(n759) );
XOR U1267 ( .A(c253), .B(b[253]), .Z(n760) );
XNOR U1268 ( .A(b[253]), .B(n761), .Z(c[253]) );
XNOR U1269 ( .A(a[253]), .B(c253), .Z(n761) );
XOR U1270 ( .A(c254), .B(n762), .Z(c255) );
ANDN U1271 ( .B(n763), .A(n764), .Z(n762) );
XOR U1272 ( .A(c254), .B(b[254]), .Z(n763) );
XNOR U1273 ( .A(b[254]), .B(n764), .Z(c[254]) );
XNOR U1274 ( .A(a[254]), .B(c254), .Z(n764) );
XOR U1275 ( .A(c255), .B(n765), .Z(c256) );
ANDN U1276 ( .B(n766), .A(n767), .Z(n765) );
XOR U1277 ( .A(c255), .B(b[255]), .Z(n766) );
XNOR U1278 ( .A(b[255]), .B(n767), .Z(c[255]) );
XNOR U1279 ( .A(a[255]), .B(c255), .Z(n767) );
XOR U1280 ( .A(c256), .B(n768), .Z(c257) );
ANDN U1281 ( .B(n769), .A(n770), .Z(n768) );
XOR U1282 ( .A(c256), .B(b[256]), .Z(n769) );
XNOR U1283 ( .A(b[256]), .B(n770), .Z(c[256]) );
XNOR U1284 ( .A(a[256]), .B(c256), .Z(n770) );
XOR U1285 ( .A(c257), .B(n771), .Z(c258) );
ANDN U1286 ( .B(n772), .A(n773), .Z(n771) );
XOR U1287 ( .A(c257), .B(b[257]), .Z(n772) );
XNOR U1288 ( .A(b[257]), .B(n773), .Z(c[257]) );
XNOR U1289 ( .A(a[257]), .B(c257), .Z(n773) );
XOR U1290 ( .A(c258), .B(n774), .Z(c259) );
ANDN U1291 ( .B(n775), .A(n776), .Z(n774) );
XOR U1292 ( .A(c258), .B(b[258]), .Z(n775) );
XNOR U1293 ( .A(b[258]), .B(n776), .Z(c[258]) );
XNOR U1294 ( .A(a[258]), .B(c258), .Z(n776) );
XOR U1295 ( .A(c259), .B(n777), .Z(c260) );
ANDN U1296 ( .B(n778), .A(n779), .Z(n777) );
XOR U1297 ( .A(c259), .B(b[259]), .Z(n778) );
XNOR U1298 ( .A(b[259]), .B(n779), .Z(c[259]) );
XNOR U1299 ( .A(a[259]), .B(c259), .Z(n779) );
XOR U1300 ( .A(c260), .B(n780), .Z(c261) );
ANDN U1301 ( .B(n781), .A(n782), .Z(n780) );
XOR U1302 ( .A(c260), .B(b[260]), .Z(n781) );
XNOR U1303 ( .A(b[260]), .B(n782), .Z(c[260]) );
XNOR U1304 ( .A(a[260]), .B(c260), .Z(n782) );
XOR U1305 ( .A(c261), .B(n783), .Z(c262) );
ANDN U1306 ( .B(n784), .A(n785), .Z(n783) );
XOR U1307 ( .A(c261), .B(b[261]), .Z(n784) );
XNOR U1308 ( .A(b[261]), .B(n785), .Z(c[261]) );
XNOR U1309 ( .A(a[261]), .B(c261), .Z(n785) );
XOR U1310 ( .A(c262), .B(n786), .Z(c263) );
ANDN U1311 ( .B(n787), .A(n788), .Z(n786) );
XOR U1312 ( .A(c262), .B(b[262]), .Z(n787) );
XNOR U1313 ( .A(b[262]), .B(n788), .Z(c[262]) );
XNOR U1314 ( .A(a[262]), .B(c262), .Z(n788) );
XOR U1315 ( .A(c263), .B(n789), .Z(c264) );
ANDN U1316 ( .B(n790), .A(n791), .Z(n789) );
XOR U1317 ( .A(c263), .B(b[263]), .Z(n790) );
XNOR U1318 ( .A(b[263]), .B(n791), .Z(c[263]) );
XNOR U1319 ( .A(a[263]), .B(c263), .Z(n791) );
XOR U1320 ( .A(c264), .B(n792), .Z(c265) );
ANDN U1321 ( .B(n793), .A(n794), .Z(n792) );
XOR U1322 ( .A(c264), .B(b[264]), .Z(n793) );
XNOR U1323 ( .A(b[264]), .B(n794), .Z(c[264]) );
XNOR U1324 ( .A(a[264]), .B(c264), .Z(n794) );
XOR U1325 ( .A(c265), .B(n795), .Z(c266) );
ANDN U1326 ( .B(n796), .A(n797), .Z(n795) );
XOR U1327 ( .A(c265), .B(b[265]), .Z(n796) );
XNOR U1328 ( .A(b[265]), .B(n797), .Z(c[265]) );
XNOR U1329 ( .A(a[265]), .B(c265), .Z(n797) );
XOR U1330 ( .A(c266), .B(n798), .Z(c267) );
ANDN U1331 ( .B(n799), .A(n800), .Z(n798) );
XOR U1332 ( .A(c266), .B(b[266]), .Z(n799) );
XNOR U1333 ( .A(b[266]), .B(n800), .Z(c[266]) );
XNOR U1334 ( .A(a[266]), .B(c266), .Z(n800) );
XOR U1335 ( .A(c267), .B(n801), .Z(c268) );
ANDN U1336 ( .B(n802), .A(n803), .Z(n801) );
XOR U1337 ( .A(c267), .B(b[267]), .Z(n802) );
XNOR U1338 ( .A(b[267]), .B(n803), .Z(c[267]) );
XNOR U1339 ( .A(a[267]), .B(c267), .Z(n803) );
XOR U1340 ( .A(c268), .B(n804), .Z(c269) );
ANDN U1341 ( .B(n805), .A(n806), .Z(n804) );
XOR U1342 ( .A(c268), .B(b[268]), .Z(n805) );
XNOR U1343 ( .A(b[268]), .B(n806), .Z(c[268]) );
XNOR U1344 ( .A(a[268]), .B(c268), .Z(n806) );
XOR U1345 ( .A(c269), .B(n807), .Z(c270) );
ANDN U1346 ( .B(n808), .A(n809), .Z(n807) );
XOR U1347 ( .A(c269), .B(b[269]), .Z(n808) );
XNOR U1348 ( .A(b[269]), .B(n809), .Z(c[269]) );
XNOR U1349 ( .A(a[269]), .B(c269), .Z(n809) );
XOR U1350 ( .A(c270), .B(n810), .Z(c271) );
ANDN U1351 ( .B(n811), .A(n812), .Z(n810) );
XOR U1352 ( .A(c270), .B(b[270]), .Z(n811) );
XNOR U1353 ( .A(b[270]), .B(n812), .Z(c[270]) );
XNOR U1354 ( .A(a[270]), .B(c270), .Z(n812) );
XOR U1355 ( .A(c271), .B(n813), .Z(c272) );
ANDN U1356 ( .B(n814), .A(n815), .Z(n813) );
XOR U1357 ( .A(c271), .B(b[271]), .Z(n814) );
XNOR U1358 ( .A(b[271]), .B(n815), .Z(c[271]) );
XNOR U1359 ( .A(a[271]), .B(c271), .Z(n815) );
XOR U1360 ( .A(c272), .B(n816), .Z(c273) );
ANDN U1361 ( .B(n817), .A(n818), .Z(n816) );
XOR U1362 ( .A(c272), .B(b[272]), .Z(n817) );
XNOR U1363 ( .A(b[272]), .B(n818), .Z(c[272]) );
XNOR U1364 ( .A(a[272]), .B(c272), .Z(n818) );
XOR U1365 ( .A(c273), .B(n819), .Z(c274) );
ANDN U1366 ( .B(n820), .A(n821), .Z(n819) );
XOR U1367 ( .A(c273), .B(b[273]), .Z(n820) );
XNOR U1368 ( .A(b[273]), .B(n821), .Z(c[273]) );
XNOR U1369 ( .A(a[273]), .B(c273), .Z(n821) );
XOR U1370 ( .A(c274), .B(n822), .Z(c275) );
ANDN U1371 ( .B(n823), .A(n824), .Z(n822) );
XOR U1372 ( .A(c274), .B(b[274]), .Z(n823) );
XNOR U1373 ( .A(b[274]), .B(n824), .Z(c[274]) );
XNOR U1374 ( .A(a[274]), .B(c274), .Z(n824) );
XOR U1375 ( .A(c275), .B(n825), .Z(c276) );
ANDN U1376 ( .B(n826), .A(n827), .Z(n825) );
XOR U1377 ( .A(c275), .B(b[275]), .Z(n826) );
XNOR U1378 ( .A(b[275]), .B(n827), .Z(c[275]) );
XNOR U1379 ( .A(a[275]), .B(c275), .Z(n827) );
XOR U1380 ( .A(c276), .B(n828), .Z(c277) );
ANDN U1381 ( .B(n829), .A(n830), .Z(n828) );
XOR U1382 ( .A(c276), .B(b[276]), .Z(n829) );
XNOR U1383 ( .A(b[276]), .B(n830), .Z(c[276]) );
XNOR U1384 ( .A(a[276]), .B(c276), .Z(n830) );
XOR U1385 ( .A(c277), .B(n831), .Z(c278) );
ANDN U1386 ( .B(n832), .A(n833), .Z(n831) );
XOR U1387 ( .A(c277), .B(b[277]), .Z(n832) );
XNOR U1388 ( .A(b[277]), .B(n833), .Z(c[277]) );
XNOR U1389 ( .A(a[277]), .B(c277), .Z(n833) );
XOR U1390 ( .A(c278), .B(n834), .Z(c279) );
ANDN U1391 ( .B(n835), .A(n836), .Z(n834) );
XOR U1392 ( .A(c278), .B(b[278]), .Z(n835) );
XNOR U1393 ( .A(b[278]), .B(n836), .Z(c[278]) );
XNOR U1394 ( .A(a[278]), .B(c278), .Z(n836) );
XOR U1395 ( .A(c279), .B(n837), .Z(c280) );
ANDN U1396 ( .B(n838), .A(n839), .Z(n837) );
XOR U1397 ( .A(c279), .B(b[279]), .Z(n838) );
XNOR U1398 ( .A(b[279]), .B(n839), .Z(c[279]) );
XNOR U1399 ( .A(a[279]), .B(c279), .Z(n839) );
XOR U1400 ( .A(c280), .B(n840), .Z(c281) );
ANDN U1401 ( .B(n841), .A(n842), .Z(n840) );
XOR U1402 ( .A(c280), .B(b[280]), .Z(n841) );
XNOR U1403 ( .A(b[280]), .B(n842), .Z(c[280]) );
XNOR U1404 ( .A(a[280]), .B(c280), .Z(n842) );
XOR U1405 ( .A(c281), .B(n843), .Z(c282) );
ANDN U1406 ( .B(n844), .A(n845), .Z(n843) );
XOR U1407 ( .A(c281), .B(b[281]), .Z(n844) );
XNOR U1408 ( .A(b[281]), .B(n845), .Z(c[281]) );
XNOR U1409 ( .A(a[281]), .B(c281), .Z(n845) );
XOR U1410 ( .A(c282), .B(n846), .Z(c283) );
ANDN U1411 ( .B(n847), .A(n848), .Z(n846) );
XOR U1412 ( .A(c282), .B(b[282]), .Z(n847) );
XNOR U1413 ( .A(b[282]), .B(n848), .Z(c[282]) );
XNOR U1414 ( .A(a[282]), .B(c282), .Z(n848) );
XOR U1415 ( .A(c283), .B(n849), .Z(c284) );
ANDN U1416 ( .B(n850), .A(n851), .Z(n849) );
XOR U1417 ( .A(c283), .B(b[283]), .Z(n850) );
XNOR U1418 ( .A(b[283]), .B(n851), .Z(c[283]) );
XNOR U1419 ( .A(a[283]), .B(c283), .Z(n851) );
XOR U1420 ( .A(c284), .B(n852), .Z(c285) );
ANDN U1421 ( .B(n853), .A(n854), .Z(n852) );
XOR U1422 ( .A(c284), .B(b[284]), .Z(n853) );
XNOR U1423 ( .A(b[284]), .B(n854), .Z(c[284]) );
XNOR U1424 ( .A(a[284]), .B(c284), .Z(n854) );
XOR U1425 ( .A(c285), .B(n855), .Z(c286) );
ANDN U1426 ( .B(n856), .A(n857), .Z(n855) );
XOR U1427 ( .A(c285), .B(b[285]), .Z(n856) );
XNOR U1428 ( .A(b[285]), .B(n857), .Z(c[285]) );
XNOR U1429 ( .A(a[285]), .B(c285), .Z(n857) );
XOR U1430 ( .A(c286), .B(n858), .Z(c287) );
ANDN U1431 ( .B(n859), .A(n860), .Z(n858) );
XOR U1432 ( .A(c286), .B(b[286]), .Z(n859) );
XNOR U1433 ( .A(b[286]), .B(n860), .Z(c[286]) );
XNOR U1434 ( .A(a[286]), .B(c286), .Z(n860) );
XOR U1435 ( .A(c287), .B(n861), .Z(c288) );
ANDN U1436 ( .B(n862), .A(n863), .Z(n861) );
XOR U1437 ( .A(c287), .B(b[287]), .Z(n862) );
XNOR U1438 ( .A(b[287]), .B(n863), .Z(c[287]) );
XNOR U1439 ( .A(a[287]), .B(c287), .Z(n863) );
XOR U1440 ( .A(c288), .B(n864), .Z(c289) );
ANDN U1441 ( .B(n865), .A(n866), .Z(n864) );
XOR U1442 ( .A(c288), .B(b[288]), .Z(n865) );
XNOR U1443 ( .A(b[288]), .B(n866), .Z(c[288]) );
XNOR U1444 ( .A(a[288]), .B(c288), .Z(n866) );
XOR U1445 ( .A(c289), .B(n867), .Z(c290) );
ANDN U1446 ( .B(n868), .A(n869), .Z(n867) );
XOR U1447 ( .A(c289), .B(b[289]), .Z(n868) );
XNOR U1448 ( .A(b[289]), .B(n869), .Z(c[289]) );
XNOR U1449 ( .A(a[289]), .B(c289), .Z(n869) );
XOR U1450 ( .A(c290), .B(n870), .Z(c291) );
ANDN U1451 ( .B(n871), .A(n872), .Z(n870) );
XOR U1452 ( .A(c290), .B(b[290]), .Z(n871) );
XNOR U1453 ( .A(b[290]), .B(n872), .Z(c[290]) );
XNOR U1454 ( .A(a[290]), .B(c290), .Z(n872) );
XOR U1455 ( .A(c291), .B(n873), .Z(c292) );
ANDN U1456 ( .B(n874), .A(n875), .Z(n873) );
XOR U1457 ( .A(c291), .B(b[291]), .Z(n874) );
XNOR U1458 ( .A(b[291]), .B(n875), .Z(c[291]) );
XNOR U1459 ( .A(a[291]), .B(c291), .Z(n875) );
XOR U1460 ( .A(c292), .B(n876), .Z(c293) );
ANDN U1461 ( .B(n877), .A(n878), .Z(n876) );
XOR U1462 ( .A(c292), .B(b[292]), .Z(n877) );
XNOR U1463 ( .A(b[292]), .B(n878), .Z(c[292]) );
XNOR U1464 ( .A(a[292]), .B(c292), .Z(n878) );
XOR U1465 ( .A(c293), .B(n879), .Z(c294) );
ANDN U1466 ( .B(n880), .A(n881), .Z(n879) );
XOR U1467 ( .A(c293), .B(b[293]), .Z(n880) );
XNOR U1468 ( .A(b[293]), .B(n881), .Z(c[293]) );
XNOR U1469 ( .A(a[293]), .B(c293), .Z(n881) );
XOR U1470 ( .A(c294), .B(n882), .Z(c295) );
ANDN U1471 ( .B(n883), .A(n884), .Z(n882) );
XOR U1472 ( .A(c294), .B(b[294]), .Z(n883) );
XNOR U1473 ( .A(b[294]), .B(n884), .Z(c[294]) );
XNOR U1474 ( .A(a[294]), .B(c294), .Z(n884) );
XOR U1475 ( .A(c295), .B(n885), .Z(c296) );
ANDN U1476 ( .B(n886), .A(n887), .Z(n885) );
XOR U1477 ( .A(c295), .B(b[295]), .Z(n886) );
XNOR U1478 ( .A(b[295]), .B(n887), .Z(c[295]) );
XNOR U1479 ( .A(a[295]), .B(c295), .Z(n887) );
XOR U1480 ( .A(c296), .B(n888), .Z(c297) );
ANDN U1481 ( .B(n889), .A(n890), .Z(n888) );
XOR U1482 ( .A(c296), .B(b[296]), .Z(n889) );
XNOR U1483 ( .A(b[296]), .B(n890), .Z(c[296]) );
XNOR U1484 ( .A(a[296]), .B(c296), .Z(n890) );
XOR U1485 ( .A(c297), .B(n891), .Z(c298) );
ANDN U1486 ( .B(n892), .A(n893), .Z(n891) );
XOR U1487 ( .A(c297), .B(b[297]), .Z(n892) );
XNOR U1488 ( .A(b[297]), .B(n893), .Z(c[297]) );
XNOR U1489 ( .A(a[297]), .B(c297), .Z(n893) );
XOR U1490 ( .A(c298), .B(n894), .Z(c299) );
ANDN U1491 ( .B(n895), .A(n896), .Z(n894) );
XOR U1492 ( .A(c298), .B(b[298]), .Z(n895) );
XNOR U1493 ( .A(b[298]), .B(n896), .Z(c[298]) );
XNOR U1494 ( .A(a[298]), .B(c298), .Z(n896) );
XOR U1495 ( .A(c299), .B(n897), .Z(c300) );
ANDN U1496 ( .B(n898), .A(n899), .Z(n897) );
XOR U1497 ( .A(c299), .B(b[299]), .Z(n898) );
XNOR U1498 ( .A(b[299]), .B(n899), .Z(c[299]) );
XNOR U1499 ( .A(a[299]), .B(c299), .Z(n899) );
XOR U1500 ( .A(c300), .B(n900), .Z(c301) );
ANDN U1501 ( .B(n901), .A(n902), .Z(n900) );
XOR U1502 ( .A(c300), .B(b[300]), .Z(n901) );
XNOR U1503 ( .A(b[300]), .B(n902), .Z(c[300]) );
XNOR U1504 ( .A(a[300]), .B(c300), .Z(n902) );
XOR U1505 ( .A(c301), .B(n903), .Z(c302) );
ANDN U1506 ( .B(n904), .A(n905), .Z(n903) );
XOR U1507 ( .A(c301), .B(b[301]), .Z(n904) );
XNOR U1508 ( .A(b[301]), .B(n905), .Z(c[301]) );
XNOR U1509 ( .A(a[301]), .B(c301), .Z(n905) );
XOR U1510 ( .A(c302), .B(n906), .Z(c303) );
ANDN U1511 ( .B(n907), .A(n908), .Z(n906) );
XOR U1512 ( .A(c302), .B(b[302]), .Z(n907) );
XNOR U1513 ( .A(b[302]), .B(n908), .Z(c[302]) );
XNOR U1514 ( .A(a[302]), .B(c302), .Z(n908) );
XOR U1515 ( .A(c303), .B(n909), .Z(c304) );
ANDN U1516 ( .B(n910), .A(n911), .Z(n909) );
XOR U1517 ( .A(c303), .B(b[303]), .Z(n910) );
XNOR U1518 ( .A(b[303]), .B(n911), .Z(c[303]) );
XNOR U1519 ( .A(a[303]), .B(c303), .Z(n911) );
XOR U1520 ( .A(c304), .B(n912), .Z(c305) );
ANDN U1521 ( .B(n913), .A(n914), .Z(n912) );
XOR U1522 ( .A(c304), .B(b[304]), .Z(n913) );
XNOR U1523 ( .A(b[304]), .B(n914), .Z(c[304]) );
XNOR U1524 ( .A(a[304]), .B(c304), .Z(n914) );
XOR U1525 ( .A(c305), .B(n915), .Z(c306) );
ANDN U1526 ( .B(n916), .A(n917), .Z(n915) );
XOR U1527 ( .A(c305), .B(b[305]), .Z(n916) );
XNOR U1528 ( .A(b[305]), .B(n917), .Z(c[305]) );
XNOR U1529 ( .A(a[305]), .B(c305), .Z(n917) );
XOR U1530 ( .A(c306), .B(n918), .Z(c307) );
ANDN U1531 ( .B(n919), .A(n920), .Z(n918) );
XOR U1532 ( .A(c306), .B(b[306]), .Z(n919) );
XNOR U1533 ( .A(b[306]), .B(n920), .Z(c[306]) );
XNOR U1534 ( .A(a[306]), .B(c306), .Z(n920) );
XOR U1535 ( .A(c307), .B(n921), .Z(c308) );
ANDN U1536 ( .B(n922), .A(n923), .Z(n921) );
XOR U1537 ( .A(c307), .B(b[307]), .Z(n922) );
XNOR U1538 ( .A(b[307]), .B(n923), .Z(c[307]) );
XNOR U1539 ( .A(a[307]), .B(c307), .Z(n923) );
XOR U1540 ( .A(c308), .B(n924), .Z(c309) );
ANDN U1541 ( .B(n925), .A(n926), .Z(n924) );
XOR U1542 ( .A(c308), .B(b[308]), .Z(n925) );
XNOR U1543 ( .A(b[308]), .B(n926), .Z(c[308]) );
XNOR U1544 ( .A(a[308]), .B(c308), .Z(n926) );
XOR U1545 ( .A(c309), .B(n927), .Z(c310) );
ANDN U1546 ( .B(n928), .A(n929), .Z(n927) );
XOR U1547 ( .A(c309), .B(b[309]), .Z(n928) );
XNOR U1548 ( .A(b[309]), .B(n929), .Z(c[309]) );
XNOR U1549 ( .A(a[309]), .B(c309), .Z(n929) );
XOR U1550 ( .A(c310), .B(n930), .Z(c311) );
ANDN U1551 ( .B(n931), .A(n932), .Z(n930) );
XOR U1552 ( .A(c310), .B(b[310]), .Z(n931) );
XNOR U1553 ( .A(b[310]), .B(n932), .Z(c[310]) );
XNOR U1554 ( .A(a[310]), .B(c310), .Z(n932) );
XOR U1555 ( .A(c311), .B(n933), .Z(c312) );
ANDN U1556 ( .B(n934), .A(n935), .Z(n933) );
XOR U1557 ( .A(c311), .B(b[311]), .Z(n934) );
XNOR U1558 ( .A(b[311]), .B(n935), .Z(c[311]) );
XNOR U1559 ( .A(a[311]), .B(c311), .Z(n935) );
XOR U1560 ( .A(c312), .B(n936), .Z(c313) );
ANDN U1561 ( .B(n937), .A(n938), .Z(n936) );
XOR U1562 ( .A(c312), .B(b[312]), .Z(n937) );
XNOR U1563 ( .A(b[312]), .B(n938), .Z(c[312]) );
XNOR U1564 ( .A(a[312]), .B(c312), .Z(n938) );
XOR U1565 ( .A(c313), .B(n939), .Z(c314) );
ANDN U1566 ( .B(n940), .A(n941), .Z(n939) );
XOR U1567 ( .A(c313), .B(b[313]), .Z(n940) );
XNOR U1568 ( .A(b[313]), .B(n941), .Z(c[313]) );
XNOR U1569 ( .A(a[313]), .B(c313), .Z(n941) );
XOR U1570 ( .A(c314), .B(n942), .Z(c315) );
ANDN U1571 ( .B(n943), .A(n944), .Z(n942) );
XOR U1572 ( .A(c314), .B(b[314]), .Z(n943) );
XNOR U1573 ( .A(b[314]), .B(n944), .Z(c[314]) );
XNOR U1574 ( .A(a[314]), .B(c314), .Z(n944) );
XOR U1575 ( .A(c315), .B(n945), .Z(c316) );
ANDN U1576 ( .B(n946), .A(n947), .Z(n945) );
XOR U1577 ( .A(c315), .B(b[315]), .Z(n946) );
XNOR U1578 ( .A(b[315]), .B(n947), .Z(c[315]) );
XNOR U1579 ( .A(a[315]), .B(c315), .Z(n947) );
XOR U1580 ( .A(c316), .B(n948), .Z(c317) );
ANDN U1581 ( .B(n949), .A(n950), .Z(n948) );
XOR U1582 ( .A(c316), .B(b[316]), .Z(n949) );
XNOR U1583 ( .A(b[316]), .B(n950), .Z(c[316]) );
XNOR U1584 ( .A(a[316]), .B(c316), .Z(n950) );
XOR U1585 ( .A(c317), .B(n951), .Z(c318) );
ANDN U1586 ( .B(n952), .A(n953), .Z(n951) );
XOR U1587 ( .A(c317), .B(b[317]), .Z(n952) );
XNOR U1588 ( .A(b[317]), .B(n953), .Z(c[317]) );
XNOR U1589 ( .A(a[317]), .B(c317), .Z(n953) );
XOR U1590 ( .A(c318), .B(n954), .Z(c319) );
ANDN U1591 ( .B(n955), .A(n956), .Z(n954) );
XOR U1592 ( .A(c318), .B(b[318]), .Z(n955) );
XNOR U1593 ( .A(b[318]), .B(n956), .Z(c[318]) );
XNOR U1594 ( .A(a[318]), .B(c318), .Z(n956) );
XOR U1595 ( .A(c319), .B(n957), .Z(c320) );
ANDN U1596 ( .B(n958), .A(n959), .Z(n957) );
XOR U1597 ( .A(c319), .B(b[319]), .Z(n958) );
XNOR U1598 ( .A(b[319]), .B(n959), .Z(c[319]) );
XNOR U1599 ( .A(a[319]), .B(c319), .Z(n959) );
XOR U1600 ( .A(c320), .B(n960), .Z(c321) );
ANDN U1601 ( .B(n961), .A(n962), .Z(n960) );
XOR U1602 ( .A(c320), .B(b[320]), .Z(n961) );
XNOR U1603 ( .A(b[320]), .B(n962), .Z(c[320]) );
XNOR U1604 ( .A(a[320]), .B(c320), .Z(n962) );
XOR U1605 ( .A(c321), .B(n963), .Z(c322) );
ANDN U1606 ( .B(n964), .A(n965), .Z(n963) );
XOR U1607 ( .A(c321), .B(b[321]), .Z(n964) );
XNOR U1608 ( .A(b[321]), .B(n965), .Z(c[321]) );
XNOR U1609 ( .A(a[321]), .B(c321), .Z(n965) );
XOR U1610 ( .A(c322), .B(n966), .Z(c323) );
ANDN U1611 ( .B(n967), .A(n968), .Z(n966) );
XOR U1612 ( .A(c322), .B(b[322]), .Z(n967) );
XNOR U1613 ( .A(b[322]), .B(n968), .Z(c[322]) );
XNOR U1614 ( .A(a[322]), .B(c322), .Z(n968) );
XOR U1615 ( .A(c323), .B(n969), .Z(c324) );
ANDN U1616 ( .B(n970), .A(n971), .Z(n969) );
XOR U1617 ( .A(c323), .B(b[323]), .Z(n970) );
XNOR U1618 ( .A(b[323]), .B(n971), .Z(c[323]) );
XNOR U1619 ( .A(a[323]), .B(c323), .Z(n971) );
XOR U1620 ( .A(c324), .B(n972), .Z(c325) );
ANDN U1621 ( .B(n973), .A(n974), .Z(n972) );
XOR U1622 ( .A(c324), .B(b[324]), .Z(n973) );
XNOR U1623 ( .A(b[324]), .B(n974), .Z(c[324]) );
XNOR U1624 ( .A(a[324]), .B(c324), .Z(n974) );
XOR U1625 ( .A(c325), .B(n975), .Z(c326) );
ANDN U1626 ( .B(n976), .A(n977), .Z(n975) );
XOR U1627 ( .A(c325), .B(b[325]), .Z(n976) );
XNOR U1628 ( .A(b[325]), .B(n977), .Z(c[325]) );
XNOR U1629 ( .A(a[325]), .B(c325), .Z(n977) );
XOR U1630 ( .A(c326), .B(n978), .Z(c327) );
ANDN U1631 ( .B(n979), .A(n980), .Z(n978) );
XOR U1632 ( .A(c326), .B(b[326]), .Z(n979) );
XNOR U1633 ( .A(b[326]), .B(n980), .Z(c[326]) );
XNOR U1634 ( .A(a[326]), .B(c326), .Z(n980) );
XOR U1635 ( .A(c327), .B(n981), .Z(c328) );
ANDN U1636 ( .B(n982), .A(n983), .Z(n981) );
XOR U1637 ( .A(c327), .B(b[327]), .Z(n982) );
XNOR U1638 ( .A(b[327]), .B(n983), .Z(c[327]) );
XNOR U1639 ( .A(a[327]), .B(c327), .Z(n983) );
XOR U1640 ( .A(c328), .B(n984), .Z(c329) );
ANDN U1641 ( .B(n985), .A(n986), .Z(n984) );
XOR U1642 ( .A(c328), .B(b[328]), .Z(n985) );
XNOR U1643 ( .A(b[328]), .B(n986), .Z(c[328]) );
XNOR U1644 ( .A(a[328]), .B(c328), .Z(n986) );
XOR U1645 ( .A(c329), .B(n987), .Z(c330) );
ANDN U1646 ( .B(n988), .A(n989), .Z(n987) );
XOR U1647 ( .A(c329), .B(b[329]), .Z(n988) );
XNOR U1648 ( .A(b[329]), .B(n989), .Z(c[329]) );
XNOR U1649 ( .A(a[329]), .B(c329), .Z(n989) );
XOR U1650 ( .A(c330), .B(n990), .Z(c331) );
ANDN U1651 ( .B(n991), .A(n992), .Z(n990) );
XOR U1652 ( .A(c330), .B(b[330]), .Z(n991) );
XNOR U1653 ( .A(b[330]), .B(n992), .Z(c[330]) );
XNOR U1654 ( .A(a[330]), .B(c330), .Z(n992) );
XOR U1655 ( .A(c331), .B(n993), .Z(c332) );
ANDN U1656 ( .B(n994), .A(n995), .Z(n993) );
XOR U1657 ( .A(c331), .B(b[331]), .Z(n994) );
XNOR U1658 ( .A(b[331]), .B(n995), .Z(c[331]) );
XNOR U1659 ( .A(a[331]), .B(c331), .Z(n995) );
XOR U1660 ( .A(c332), .B(n996), .Z(c333) );
ANDN U1661 ( .B(n997), .A(n998), .Z(n996) );
XOR U1662 ( .A(c332), .B(b[332]), .Z(n997) );
XNOR U1663 ( .A(b[332]), .B(n998), .Z(c[332]) );
XNOR U1664 ( .A(a[332]), .B(c332), .Z(n998) );
XOR U1665 ( .A(c333), .B(n999), .Z(c334) );
ANDN U1666 ( .B(n1000), .A(n1001), .Z(n999) );
XOR U1667 ( .A(c333), .B(b[333]), .Z(n1000) );
XNOR U1668 ( .A(b[333]), .B(n1001), .Z(c[333]) );
XNOR U1669 ( .A(a[333]), .B(c333), .Z(n1001) );
XOR U1670 ( .A(c334), .B(n1002), .Z(c335) );
ANDN U1671 ( .B(n1003), .A(n1004), .Z(n1002) );
XOR U1672 ( .A(c334), .B(b[334]), .Z(n1003) );
XNOR U1673 ( .A(b[334]), .B(n1004), .Z(c[334]) );
XNOR U1674 ( .A(a[334]), .B(c334), .Z(n1004) );
XOR U1675 ( .A(c335), .B(n1005), .Z(c336) );
ANDN U1676 ( .B(n1006), .A(n1007), .Z(n1005) );
XOR U1677 ( .A(c335), .B(b[335]), .Z(n1006) );
XNOR U1678 ( .A(b[335]), .B(n1007), .Z(c[335]) );
XNOR U1679 ( .A(a[335]), .B(c335), .Z(n1007) );
XOR U1680 ( .A(c336), .B(n1008), .Z(c337) );
ANDN U1681 ( .B(n1009), .A(n1010), .Z(n1008) );
XOR U1682 ( .A(c336), .B(b[336]), .Z(n1009) );
XNOR U1683 ( .A(b[336]), .B(n1010), .Z(c[336]) );
XNOR U1684 ( .A(a[336]), .B(c336), .Z(n1010) );
XOR U1685 ( .A(c337), .B(n1011), .Z(c338) );
ANDN U1686 ( .B(n1012), .A(n1013), .Z(n1011) );
XOR U1687 ( .A(c337), .B(b[337]), .Z(n1012) );
XNOR U1688 ( .A(b[337]), .B(n1013), .Z(c[337]) );
XNOR U1689 ( .A(a[337]), .B(c337), .Z(n1013) );
XOR U1690 ( .A(c338), .B(n1014), .Z(c339) );
ANDN U1691 ( .B(n1015), .A(n1016), .Z(n1014) );
XOR U1692 ( .A(c338), .B(b[338]), .Z(n1015) );
XNOR U1693 ( .A(b[338]), .B(n1016), .Z(c[338]) );
XNOR U1694 ( .A(a[338]), .B(c338), .Z(n1016) );
XOR U1695 ( .A(c339), .B(n1017), .Z(c340) );
ANDN U1696 ( .B(n1018), .A(n1019), .Z(n1017) );
XOR U1697 ( .A(c339), .B(b[339]), .Z(n1018) );
XNOR U1698 ( .A(b[339]), .B(n1019), .Z(c[339]) );
XNOR U1699 ( .A(a[339]), .B(c339), .Z(n1019) );
XOR U1700 ( .A(c340), .B(n1020), .Z(c341) );
ANDN U1701 ( .B(n1021), .A(n1022), .Z(n1020) );
XOR U1702 ( .A(c340), .B(b[340]), .Z(n1021) );
XNOR U1703 ( .A(b[340]), .B(n1022), .Z(c[340]) );
XNOR U1704 ( .A(a[340]), .B(c340), .Z(n1022) );
XOR U1705 ( .A(c341), .B(n1023), .Z(c342) );
ANDN U1706 ( .B(n1024), .A(n1025), .Z(n1023) );
XOR U1707 ( .A(c341), .B(b[341]), .Z(n1024) );
XNOR U1708 ( .A(b[341]), .B(n1025), .Z(c[341]) );
XNOR U1709 ( .A(a[341]), .B(c341), .Z(n1025) );
XOR U1710 ( .A(c342), .B(n1026), .Z(c343) );
ANDN U1711 ( .B(n1027), .A(n1028), .Z(n1026) );
XOR U1712 ( .A(c342), .B(b[342]), .Z(n1027) );
XNOR U1713 ( .A(b[342]), .B(n1028), .Z(c[342]) );
XNOR U1714 ( .A(a[342]), .B(c342), .Z(n1028) );
XOR U1715 ( .A(c343), .B(n1029), .Z(c344) );
ANDN U1716 ( .B(n1030), .A(n1031), .Z(n1029) );
XOR U1717 ( .A(c343), .B(b[343]), .Z(n1030) );
XNOR U1718 ( .A(b[343]), .B(n1031), .Z(c[343]) );
XNOR U1719 ( .A(a[343]), .B(c343), .Z(n1031) );
XOR U1720 ( .A(c344), .B(n1032), .Z(c345) );
ANDN U1721 ( .B(n1033), .A(n1034), .Z(n1032) );
XOR U1722 ( .A(c344), .B(b[344]), .Z(n1033) );
XNOR U1723 ( .A(b[344]), .B(n1034), .Z(c[344]) );
XNOR U1724 ( .A(a[344]), .B(c344), .Z(n1034) );
XOR U1725 ( .A(c345), .B(n1035), .Z(c346) );
ANDN U1726 ( .B(n1036), .A(n1037), .Z(n1035) );
XOR U1727 ( .A(c345), .B(b[345]), .Z(n1036) );
XNOR U1728 ( .A(b[345]), .B(n1037), .Z(c[345]) );
XNOR U1729 ( .A(a[345]), .B(c345), .Z(n1037) );
XOR U1730 ( .A(c346), .B(n1038), .Z(c347) );
ANDN U1731 ( .B(n1039), .A(n1040), .Z(n1038) );
XOR U1732 ( .A(c346), .B(b[346]), .Z(n1039) );
XNOR U1733 ( .A(b[346]), .B(n1040), .Z(c[346]) );
XNOR U1734 ( .A(a[346]), .B(c346), .Z(n1040) );
XOR U1735 ( .A(c347), .B(n1041), .Z(c348) );
ANDN U1736 ( .B(n1042), .A(n1043), .Z(n1041) );
XOR U1737 ( .A(c347), .B(b[347]), .Z(n1042) );
XNOR U1738 ( .A(b[347]), .B(n1043), .Z(c[347]) );
XNOR U1739 ( .A(a[347]), .B(c347), .Z(n1043) );
XOR U1740 ( .A(c348), .B(n1044), .Z(c349) );
ANDN U1741 ( .B(n1045), .A(n1046), .Z(n1044) );
XOR U1742 ( .A(c348), .B(b[348]), .Z(n1045) );
XNOR U1743 ( .A(b[348]), .B(n1046), .Z(c[348]) );
XNOR U1744 ( .A(a[348]), .B(c348), .Z(n1046) );
XOR U1745 ( .A(c349), .B(n1047), .Z(c350) );
ANDN U1746 ( .B(n1048), .A(n1049), .Z(n1047) );
XOR U1747 ( .A(c349), .B(b[349]), .Z(n1048) );
XNOR U1748 ( .A(b[349]), .B(n1049), .Z(c[349]) );
XNOR U1749 ( .A(a[349]), .B(c349), .Z(n1049) );
XOR U1750 ( .A(c350), .B(n1050), .Z(c351) );
ANDN U1751 ( .B(n1051), .A(n1052), .Z(n1050) );
XOR U1752 ( .A(c350), .B(b[350]), .Z(n1051) );
XNOR U1753 ( .A(b[350]), .B(n1052), .Z(c[350]) );
XNOR U1754 ( .A(a[350]), .B(c350), .Z(n1052) );
XOR U1755 ( .A(c351), .B(n1053), .Z(c352) );
ANDN U1756 ( .B(n1054), .A(n1055), .Z(n1053) );
XOR U1757 ( .A(c351), .B(b[351]), .Z(n1054) );
XNOR U1758 ( .A(b[351]), .B(n1055), .Z(c[351]) );
XNOR U1759 ( .A(a[351]), .B(c351), .Z(n1055) );
XOR U1760 ( .A(c352), .B(n1056), .Z(c353) );
ANDN U1761 ( .B(n1057), .A(n1058), .Z(n1056) );
XOR U1762 ( .A(c352), .B(b[352]), .Z(n1057) );
XNOR U1763 ( .A(b[352]), .B(n1058), .Z(c[352]) );
XNOR U1764 ( .A(a[352]), .B(c352), .Z(n1058) );
XOR U1765 ( .A(c353), .B(n1059), .Z(c354) );
ANDN U1766 ( .B(n1060), .A(n1061), .Z(n1059) );
XOR U1767 ( .A(c353), .B(b[353]), .Z(n1060) );
XNOR U1768 ( .A(b[353]), .B(n1061), .Z(c[353]) );
XNOR U1769 ( .A(a[353]), .B(c353), .Z(n1061) );
XOR U1770 ( .A(c354), .B(n1062), .Z(c355) );
ANDN U1771 ( .B(n1063), .A(n1064), .Z(n1062) );
XOR U1772 ( .A(c354), .B(b[354]), .Z(n1063) );
XNOR U1773 ( .A(b[354]), .B(n1064), .Z(c[354]) );
XNOR U1774 ( .A(a[354]), .B(c354), .Z(n1064) );
XOR U1775 ( .A(c355), .B(n1065), .Z(c356) );
ANDN U1776 ( .B(n1066), .A(n1067), .Z(n1065) );
XOR U1777 ( .A(c355), .B(b[355]), .Z(n1066) );
XNOR U1778 ( .A(b[355]), .B(n1067), .Z(c[355]) );
XNOR U1779 ( .A(a[355]), .B(c355), .Z(n1067) );
XOR U1780 ( .A(c356), .B(n1068), .Z(c357) );
ANDN U1781 ( .B(n1069), .A(n1070), .Z(n1068) );
XOR U1782 ( .A(c356), .B(b[356]), .Z(n1069) );
XNOR U1783 ( .A(b[356]), .B(n1070), .Z(c[356]) );
XNOR U1784 ( .A(a[356]), .B(c356), .Z(n1070) );
XOR U1785 ( .A(c357), .B(n1071), .Z(c358) );
ANDN U1786 ( .B(n1072), .A(n1073), .Z(n1071) );
XOR U1787 ( .A(c357), .B(b[357]), .Z(n1072) );
XNOR U1788 ( .A(b[357]), .B(n1073), .Z(c[357]) );
XNOR U1789 ( .A(a[357]), .B(c357), .Z(n1073) );
XOR U1790 ( .A(c358), .B(n1074), .Z(c359) );
ANDN U1791 ( .B(n1075), .A(n1076), .Z(n1074) );
XOR U1792 ( .A(c358), .B(b[358]), .Z(n1075) );
XNOR U1793 ( .A(b[358]), .B(n1076), .Z(c[358]) );
XNOR U1794 ( .A(a[358]), .B(c358), .Z(n1076) );
XOR U1795 ( .A(c359), .B(n1077), .Z(c360) );
ANDN U1796 ( .B(n1078), .A(n1079), .Z(n1077) );
XOR U1797 ( .A(c359), .B(b[359]), .Z(n1078) );
XNOR U1798 ( .A(b[359]), .B(n1079), .Z(c[359]) );
XNOR U1799 ( .A(a[359]), .B(c359), .Z(n1079) );
XOR U1800 ( .A(c360), .B(n1080), .Z(c361) );
ANDN U1801 ( .B(n1081), .A(n1082), .Z(n1080) );
XOR U1802 ( .A(c360), .B(b[360]), .Z(n1081) );
XNOR U1803 ( .A(b[360]), .B(n1082), .Z(c[360]) );
XNOR U1804 ( .A(a[360]), .B(c360), .Z(n1082) );
XOR U1805 ( .A(c361), .B(n1083), .Z(c362) );
ANDN U1806 ( .B(n1084), .A(n1085), .Z(n1083) );
XOR U1807 ( .A(c361), .B(b[361]), .Z(n1084) );
XNOR U1808 ( .A(b[361]), .B(n1085), .Z(c[361]) );
XNOR U1809 ( .A(a[361]), .B(c361), .Z(n1085) );
XOR U1810 ( .A(c362), .B(n1086), .Z(c363) );
ANDN U1811 ( .B(n1087), .A(n1088), .Z(n1086) );
XOR U1812 ( .A(c362), .B(b[362]), .Z(n1087) );
XNOR U1813 ( .A(b[362]), .B(n1088), .Z(c[362]) );
XNOR U1814 ( .A(a[362]), .B(c362), .Z(n1088) );
XOR U1815 ( .A(c363), .B(n1089), .Z(c364) );
ANDN U1816 ( .B(n1090), .A(n1091), .Z(n1089) );
XOR U1817 ( .A(c363), .B(b[363]), .Z(n1090) );
XNOR U1818 ( .A(b[363]), .B(n1091), .Z(c[363]) );
XNOR U1819 ( .A(a[363]), .B(c363), .Z(n1091) );
XOR U1820 ( .A(c364), .B(n1092), .Z(c365) );
ANDN U1821 ( .B(n1093), .A(n1094), .Z(n1092) );
XOR U1822 ( .A(c364), .B(b[364]), .Z(n1093) );
XNOR U1823 ( .A(b[364]), .B(n1094), .Z(c[364]) );
XNOR U1824 ( .A(a[364]), .B(c364), .Z(n1094) );
XOR U1825 ( .A(c365), .B(n1095), .Z(c366) );
ANDN U1826 ( .B(n1096), .A(n1097), .Z(n1095) );
XOR U1827 ( .A(c365), .B(b[365]), .Z(n1096) );
XNOR U1828 ( .A(b[365]), .B(n1097), .Z(c[365]) );
XNOR U1829 ( .A(a[365]), .B(c365), .Z(n1097) );
XOR U1830 ( .A(c366), .B(n1098), .Z(c367) );
ANDN U1831 ( .B(n1099), .A(n1100), .Z(n1098) );
XOR U1832 ( .A(c366), .B(b[366]), .Z(n1099) );
XNOR U1833 ( .A(b[366]), .B(n1100), .Z(c[366]) );
XNOR U1834 ( .A(a[366]), .B(c366), .Z(n1100) );
XOR U1835 ( .A(c367), .B(n1101), .Z(c368) );
ANDN U1836 ( .B(n1102), .A(n1103), .Z(n1101) );
XOR U1837 ( .A(c367), .B(b[367]), .Z(n1102) );
XNOR U1838 ( .A(b[367]), .B(n1103), .Z(c[367]) );
XNOR U1839 ( .A(a[367]), .B(c367), .Z(n1103) );
XOR U1840 ( .A(c368), .B(n1104), .Z(c369) );
ANDN U1841 ( .B(n1105), .A(n1106), .Z(n1104) );
XOR U1842 ( .A(c368), .B(b[368]), .Z(n1105) );
XNOR U1843 ( .A(b[368]), .B(n1106), .Z(c[368]) );
XNOR U1844 ( .A(a[368]), .B(c368), .Z(n1106) );
XOR U1845 ( .A(c369), .B(n1107), .Z(c370) );
ANDN U1846 ( .B(n1108), .A(n1109), .Z(n1107) );
XOR U1847 ( .A(c369), .B(b[369]), .Z(n1108) );
XNOR U1848 ( .A(b[369]), .B(n1109), .Z(c[369]) );
XNOR U1849 ( .A(a[369]), .B(c369), .Z(n1109) );
XOR U1850 ( .A(c370), .B(n1110), .Z(c371) );
ANDN U1851 ( .B(n1111), .A(n1112), .Z(n1110) );
XOR U1852 ( .A(c370), .B(b[370]), .Z(n1111) );
XNOR U1853 ( .A(b[370]), .B(n1112), .Z(c[370]) );
XNOR U1854 ( .A(a[370]), .B(c370), .Z(n1112) );
XOR U1855 ( .A(c371), .B(n1113), .Z(c372) );
ANDN U1856 ( .B(n1114), .A(n1115), .Z(n1113) );
XOR U1857 ( .A(c371), .B(b[371]), .Z(n1114) );
XNOR U1858 ( .A(b[371]), .B(n1115), .Z(c[371]) );
XNOR U1859 ( .A(a[371]), .B(c371), .Z(n1115) );
XOR U1860 ( .A(c372), .B(n1116), .Z(c373) );
ANDN U1861 ( .B(n1117), .A(n1118), .Z(n1116) );
XOR U1862 ( .A(c372), .B(b[372]), .Z(n1117) );
XNOR U1863 ( .A(b[372]), .B(n1118), .Z(c[372]) );
XNOR U1864 ( .A(a[372]), .B(c372), .Z(n1118) );
XOR U1865 ( .A(c373), .B(n1119), .Z(c374) );
ANDN U1866 ( .B(n1120), .A(n1121), .Z(n1119) );
XOR U1867 ( .A(c373), .B(b[373]), .Z(n1120) );
XNOR U1868 ( .A(b[373]), .B(n1121), .Z(c[373]) );
XNOR U1869 ( .A(a[373]), .B(c373), .Z(n1121) );
XOR U1870 ( .A(c374), .B(n1122), .Z(c375) );
ANDN U1871 ( .B(n1123), .A(n1124), .Z(n1122) );
XOR U1872 ( .A(c374), .B(b[374]), .Z(n1123) );
XNOR U1873 ( .A(b[374]), .B(n1124), .Z(c[374]) );
XNOR U1874 ( .A(a[374]), .B(c374), .Z(n1124) );
XOR U1875 ( .A(c375), .B(n1125), .Z(c376) );
ANDN U1876 ( .B(n1126), .A(n1127), .Z(n1125) );
XOR U1877 ( .A(c375), .B(b[375]), .Z(n1126) );
XNOR U1878 ( .A(b[375]), .B(n1127), .Z(c[375]) );
XNOR U1879 ( .A(a[375]), .B(c375), .Z(n1127) );
XOR U1880 ( .A(c376), .B(n1128), .Z(c377) );
ANDN U1881 ( .B(n1129), .A(n1130), .Z(n1128) );
XOR U1882 ( .A(c376), .B(b[376]), .Z(n1129) );
XNOR U1883 ( .A(b[376]), .B(n1130), .Z(c[376]) );
XNOR U1884 ( .A(a[376]), .B(c376), .Z(n1130) );
XOR U1885 ( .A(c377), .B(n1131), .Z(c378) );
ANDN U1886 ( .B(n1132), .A(n1133), .Z(n1131) );
XOR U1887 ( .A(c377), .B(b[377]), .Z(n1132) );
XNOR U1888 ( .A(b[377]), .B(n1133), .Z(c[377]) );
XNOR U1889 ( .A(a[377]), .B(c377), .Z(n1133) );
XOR U1890 ( .A(c378), .B(n1134), .Z(c379) );
ANDN U1891 ( .B(n1135), .A(n1136), .Z(n1134) );
XOR U1892 ( .A(c378), .B(b[378]), .Z(n1135) );
XNOR U1893 ( .A(b[378]), .B(n1136), .Z(c[378]) );
XNOR U1894 ( .A(a[378]), .B(c378), .Z(n1136) );
XOR U1895 ( .A(c379), .B(n1137), .Z(c380) );
ANDN U1896 ( .B(n1138), .A(n1139), .Z(n1137) );
XOR U1897 ( .A(c379), .B(b[379]), .Z(n1138) );
XNOR U1898 ( .A(b[379]), .B(n1139), .Z(c[379]) );
XNOR U1899 ( .A(a[379]), .B(c379), .Z(n1139) );
XOR U1900 ( .A(c380), .B(n1140), .Z(c381) );
ANDN U1901 ( .B(n1141), .A(n1142), .Z(n1140) );
XOR U1902 ( .A(c380), .B(b[380]), .Z(n1141) );
XNOR U1903 ( .A(b[380]), .B(n1142), .Z(c[380]) );
XNOR U1904 ( .A(a[380]), .B(c380), .Z(n1142) );
XOR U1905 ( .A(c381), .B(n1143), .Z(c382) );
ANDN U1906 ( .B(n1144), .A(n1145), .Z(n1143) );
XOR U1907 ( .A(c381), .B(b[381]), .Z(n1144) );
XNOR U1908 ( .A(b[381]), .B(n1145), .Z(c[381]) );
XNOR U1909 ( .A(a[381]), .B(c381), .Z(n1145) );
XOR U1910 ( .A(c382), .B(n1146), .Z(c383) );
ANDN U1911 ( .B(n1147), .A(n1148), .Z(n1146) );
XOR U1912 ( .A(c382), .B(b[382]), .Z(n1147) );
XNOR U1913 ( .A(b[382]), .B(n1148), .Z(c[382]) );
XNOR U1914 ( .A(a[382]), .B(c382), .Z(n1148) );
XOR U1915 ( .A(c383), .B(n1149), .Z(c384) );
ANDN U1916 ( .B(n1150), .A(n1151), .Z(n1149) );
XOR U1917 ( .A(c383), .B(b[383]), .Z(n1150) );
XNOR U1918 ( .A(b[383]), .B(n1151), .Z(c[383]) );
XNOR U1919 ( .A(a[383]), .B(c383), .Z(n1151) );
XOR U1920 ( .A(c384), .B(n1152), .Z(c385) );
ANDN U1921 ( .B(n1153), .A(n1154), .Z(n1152) );
XOR U1922 ( .A(c384), .B(b[384]), .Z(n1153) );
XNOR U1923 ( .A(b[384]), .B(n1154), .Z(c[384]) );
XNOR U1924 ( .A(a[384]), .B(c384), .Z(n1154) );
XOR U1925 ( .A(c385), .B(n1155), .Z(c386) );
ANDN U1926 ( .B(n1156), .A(n1157), .Z(n1155) );
XOR U1927 ( .A(c385), .B(b[385]), .Z(n1156) );
XNOR U1928 ( .A(b[385]), .B(n1157), .Z(c[385]) );
XNOR U1929 ( .A(a[385]), .B(c385), .Z(n1157) );
XOR U1930 ( .A(c386), .B(n1158), .Z(c387) );
ANDN U1931 ( .B(n1159), .A(n1160), .Z(n1158) );
XOR U1932 ( .A(c386), .B(b[386]), .Z(n1159) );
XNOR U1933 ( .A(b[386]), .B(n1160), .Z(c[386]) );
XNOR U1934 ( .A(a[386]), .B(c386), .Z(n1160) );
XOR U1935 ( .A(c387), .B(n1161), .Z(c388) );
ANDN U1936 ( .B(n1162), .A(n1163), .Z(n1161) );
XOR U1937 ( .A(c387), .B(b[387]), .Z(n1162) );
XNOR U1938 ( .A(b[387]), .B(n1163), .Z(c[387]) );
XNOR U1939 ( .A(a[387]), .B(c387), .Z(n1163) );
XOR U1940 ( .A(c388), .B(n1164), .Z(c389) );
ANDN U1941 ( .B(n1165), .A(n1166), .Z(n1164) );
XOR U1942 ( .A(c388), .B(b[388]), .Z(n1165) );
XNOR U1943 ( .A(b[388]), .B(n1166), .Z(c[388]) );
XNOR U1944 ( .A(a[388]), .B(c388), .Z(n1166) );
XOR U1945 ( .A(c389), .B(n1167), .Z(c390) );
ANDN U1946 ( .B(n1168), .A(n1169), .Z(n1167) );
XOR U1947 ( .A(c389), .B(b[389]), .Z(n1168) );
XNOR U1948 ( .A(b[389]), .B(n1169), .Z(c[389]) );
XNOR U1949 ( .A(a[389]), .B(c389), .Z(n1169) );
XOR U1950 ( .A(c390), .B(n1170), .Z(c391) );
ANDN U1951 ( .B(n1171), .A(n1172), .Z(n1170) );
XOR U1952 ( .A(c390), .B(b[390]), .Z(n1171) );
XNOR U1953 ( .A(b[390]), .B(n1172), .Z(c[390]) );
XNOR U1954 ( .A(a[390]), .B(c390), .Z(n1172) );
XOR U1955 ( .A(c391), .B(n1173), .Z(c392) );
ANDN U1956 ( .B(n1174), .A(n1175), .Z(n1173) );
XOR U1957 ( .A(c391), .B(b[391]), .Z(n1174) );
XNOR U1958 ( .A(b[391]), .B(n1175), .Z(c[391]) );
XNOR U1959 ( .A(a[391]), .B(c391), .Z(n1175) );
XOR U1960 ( .A(c392), .B(n1176), .Z(c393) );
ANDN U1961 ( .B(n1177), .A(n1178), .Z(n1176) );
XOR U1962 ( .A(c392), .B(b[392]), .Z(n1177) );
XNOR U1963 ( .A(b[392]), .B(n1178), .Z(c[392]) );
XNOR U1964 ( .A(a[392]), .B(c392), .Z(n1178) );
XOR U1965 ( .A(c393), .B(n1179), .Z(c394) );
ANDN U1966 ( .B(n1180), .A(n1181), .Z(n1179) );
XOR U1967 ( .A(c393), .B(b[393]), .Z(n1180) );
XNOR U1968 ( .A(b[393]), .B(n1181), .Z(c[393]) );
XNOR U1969 ( .A(a[393]), .B(c393), .Z(n1181) );
XOR U1970 ( .A(c394), .B(n1182), .Z(c395) );
ANDN U1971 ( .B(n1183), .A(n1184), .Z(n1182) );
XOR U1972 ( .A(c394), .B(b[394]), .Z(n1183) );
XNOR U1973 ( .A(b[394]), .B(n1184), .Z(c[394]) );
XNOR U1974 ( .A(a[394]), .B(c394), .Z(n1184) );
XOR U1975 ( .A(c395), .B(n1185), .Z(c396) );
ANDN U1976 ( .B(n1186), .A(n1187), .Z(n1185) );
XOR U1977 ( .A(c395), .B(b[395]), .Z(n1186) );
XNOR U1978 ( .A(b[395]), .B(n1187), .Z(c[395]) );
XNOR U1979 ( .A(a[395]), .B(c395), .Z(n1187) );
XOR U1980 ( .A(c396), .B(n1188), .Z(c397) );
ANDN U1981 ( .B(n1189), .A(n1190), .Z(n1188) );
XOR U1982 ( .A(c396), .B(b[396]), .Z(n1189) );
XNOR U1983 ( .A(b[396]), .B(n1190), .Z(c[396]) );
XNOR U1984 ( .A(a[396]), .B(c396), .Z(n1190) );
XOR U1985 ( .A(c397), .B(n1191), .Z(c398) );
ANDN U1986 ( .B(n1192), .A(n1193), .Z(n1191) );
XOR U1987 ( .A(c397), .B(b[397]), .Z(n1192) );
XNOR U1988 ( .A(b[397]), .B(n1193), .Z(c[397]) );
XNOR U1989 ( .A(a[397]), .B(c397), .Z(n1193) );
XOR U1990 ( .A(c398), .B(n1194), .Z(c399) );
ANDN U1991 ( .B(n1195), .A(n1196), .Z(n1194) );
XOR U1992 ( .A(c398), .B(b[398]), .Z(n1195) );
XNOR U1993 ( .A(b[398]), .B(n1196), .Z(c[398]) );
XNOR U1994 ( .A(a[398]), .B(c398), .Z(n1196) );
XOR U1995 ( .A(c399), .B(n1197), .Z(c400) );
ANDN U1996 ( .B(n1198), .A(n1199), .Z(n1197) );
XOR U1997 ( .A(c399), .B(b[399]), .Z(n1198) );
XNOR U1998 ( .A(b[399]), .B(n1199), .Z(c[399]) );
XNOR U1999 ( .A(a[399]), .B(c399), .Z(n1199) );
XOR U2000 ( .A(c400), .B(n1200), .Z(c401) );
ANDN U2001 ( .B(n1201), .A(n1202), .Z(n1200) );
XOR U2002 ( .A(c400), .B(b[400]), .Z(n1201) );
XNOR U2003 ( .A(b[400]), .B(n1202), .Z(c[400]) );
XNOR U2004 ( .A(a[400]), .B(c400), .Z(n1202) );
XOR U2005 ( .A(c401), .B(n1203), .Z(c402) );
ANDN U2006 ( .B(n1204), .A(n1205), .Z(n1203) );
XOR U2007 ( .A(c401), .B(b[401]), .Z(n1204) );
XNOR U2008 ( .A(b[401]), .B(n1205), .Z(c[401]) );
XNOR U2009 ( .A(a[401]), .B(c401), .Z(n1205) );
XOR U2010 ( .A(c402), .B(n1206), .Z(c403) );
ANDN U2011 ( .B(n1207), .A(n1208), .Z(n1206) );
XOR U2012 ( .A(c402), .B(b[402]), .Z(n1207) );
XNOR U2013 ( .A(b[402]), .B(n1208), .Z(c[402]) );
XNOR U2014 ( .A(a[402]), .B(c402), .Z(n1208) );
XOR U2015 ( .A(c403), .B(n1209), .Z(c404) );
ANDN U2016 ( .B(n1210), .A(n1211), .Z(n1209) );
XOR U2017 ( .A(c403), .B(b[403]), .Z(n1210) );
XNOR U2018 ( .A(b[403]), .B(n1211), .Z(c[403]) );
XNOR U2019 ( .A(a[403]), .B(c403), .Z(n1211) );
XOR U2020 ( .A(c404), .B(n1212), .Z(c405) );
ANDN U2021 ( .B(n1213), .A(n1214), .Z(n1212) );
XOR U2022 ( .A(c404), .B(b[404]), .Z(n1213) );
XNOR U2023 ( .A(b[404]), .B(n1214), .Z(c[404]) );
XNOR U2024 ( .A(a[404]), .B(c404), .Z(n1214) );
XOR U2025 ( .A(c405), .B(n1215), .Z(c406) );
ANDN U2026 ( .B(n1216), .A(n1217), .Z(n1215) );
XOR U2027 ( .A(c405), .B(b[405]), .Z(n1216) );
XNOR U2028 ( .A(b[405]), .B(n1217), .Z(c[405]) );
XNOR U2029 ( .A(a[405]), .B(c405), .Z(n1217) );
XOR U2030 ( .A(c406), .B(n1218), .Z(c407) );
ANDN U2031 ( .B(n1219), .A(n1220), .Z(n1218) );
XOR U2032 ( .A(c406), .B(b[406]), .Z(n1219) );
XNOR U2033 ( .A(b[406]), .B(n1220), .Z(c[406]) );
XNOR U2034 ( .A(a[406]), .B(c406), .Z(n1220) );
XOR U2035 ( .A(c407), .B(n1221), .Z(c408) );
ANDN U2036 ( .B(n1222), .A(n1223), .Z(n1221) );
XOR U2037 ( .A(c407), .B(b[407]), .Z(n1222) );
XNOR U2038 ( .A(b[407]), .B(n1223), .Z(c[407]) );
XNOR U2039 ( .A(a[407]), .B(c407), .Z(n1223) );
XOR U2040 ( .A(c408), .B(n1224), .Z(c409) );
ANDN U2041 ( .B(n1225), .A(n1226), .Z(n1224) );
XOR U2042 ( .A(c408), .B(b[408]), .Z(n1225) );
XNOR U2043 ( .A(b[408]), .B(n1226), .Z(c[408]) );
XNOR U2044 ( .A(a[408]), .B(c408), .Z(n1226) );
XOR U2045 ( .A(c409), .B(n1227), .Z(c410) );
ANDN U2046 ( .B(n1228), .A(n1229), .Z(n1227) );
XOR U2047 ( .A(c409), .B(b[409]), .Z(n1228) );
XNOR U2048 ( .A(b[409]), .B(n1229), .Z(c[409]) );
XNOR U2049 ( .A(a[409]), .B(c409), .Z(n1229) );
XOR U2050 ( .A(c410), .B(n1230), .Z(c411) );
ANDN U2051 ( .B(n1231), .A(n1232), .Z(n1230) );
XOR U2052 ( .A(c410), .B(b[410]), .Z(n1231) );
XNOR U2053 ( .A(b[410]), .B(n1232), .Z(c[410]) );
XNOR U2054 ( .A(a[410]), .B(c410), .Z(n1232) );
XOR U2055 ( .A(c411), .B(n1233), .Z(c412) );
ANDN U2056 ( .B(n1234), .A(n1235), .Z(n1233) );
XOR U2057 ( .A(c411), .B(b[411]), .Z(n1234) );
XNOR U2058 ( .A(b[411]), .B(n1235), .Z(c[411]) );
XNOR U2059 ( .A(a[411]), .B(c411), .Z(n1235) );
XOR U2060 ( .A(c412), .B(n1236), .Z(c413) );
ANDN U2061 ( .B(n1237), .A(n1238), .Z(n1236) );
XOR U2062 ( .A(c412), .B(b[412]), .Z(n1237) );
XNOR U2063 ( .A(b[412]), .B(n1238), .Z(c[412]) );
XNOR U2064 ( .A(a[412]), .B(c412), .Z(n1238) );
XOR U2065 ( .A(c413), .B(n1239), .Z(c414) );
ANDN U2066 ( .B(n1240), .A(n1241), .Z(n1239) );
XOR U2067 ( .A(c413), .B(b[413]), .Z(n1240) );
XNOR U2068 ( .A(b[413]), .B(n1241), .Z(c[413]) );
XNOR U2069 ( .A(a[413]), .B(c413), .Z(n1241) );
XOR U2070 ( .A(c414), .B(n1242), .Z(c415) );
ANDN U2071 ( .B(n1243), .A(n1244), .Z(n1242) );
XOR U2072 ( .A(c414), .B(b[414]), .Z(n1243) );
XNOR U2073 ( .A(b[414]), .B(n1244), .Z(c[414]) );
XNOR U2074 ( .A(a[414]), .B(c414), .Z(n1244) );
XOR U2075 ( .A(c415), .B(n1245), .Z(c416) );
ANDN U2076 ( .B(n1246), .A(n1247), .Z(n1245) );
XOR U2077 ( .A(c415), .B(b[415]), .Z(n1246) );
XNOR U2078 ( .A(b[415]), .B(n1247), .Z(c[415]) );
XNOR U2079 ( .A(a[415]), .B(c415), .Z(n1247) );
XOR U2080 ( .A(c416), .B(n1248), .Z(c417) );
ANDN U2081 ( .B(n1249), .A(n1250), .Z(n1248) );
XOR U2082 ( .A(c416), .B(b[416]), .Z(n1249) );
XNOR U2083 ( .A(b[416]), .B(n1250), .Z(c[416]) );
XNOR U2084 ( .A(a[416]), .B(c416), .Z(n1250) );
XOR U2085 ( .A(c417), .B(n1251), .Z(c418) );
ANDN U2086 ( .B(n1252), .A(n1253), .Z(n1251) );
XOR U2087 ( .A(c417), .B(b[417]), .Z(n1252) );
XNOR U2088 ( .A(b[417]), .B(n1253), .Z(c[417]) );
XNOR U2089 ( .A(a[417]), .B(c417), .Z(n1253) );
XOR U2090 ( .A(c418), .B(n1254), .Z(c419) );
ANDN U2091 ( .B(n1255), .A(n1256), .Z(n1254) );
XOR U2092 ( .A(c418), .B(b[418]), .Z(n1255) );
XNOR U2093 ( .A(b[418]), .B(n1256), .Z(c[418]) );
XNOR U2094 ( .A(a[418]), .B(c418), .Z(n1256) );
XOR U2095 ( .A(c419), .B(n1257), .Z(c420) );
ANDN U2096 ( .B(n1258), .A(n1259), .Z(n1257) );
XOR U2097 ( .A(c419), .B(b[419]), .Z(n1258) );
XNOR U2098 ( .A(b[419]), .B(n1259), .Z(c[419]) );
XNOR U2099 ( .A(a[419]), .B(c419), .Z(n1259) );
XOR U2100 ( .A(c420), .B(n1260), .Z(c421) );
ANDN U2101 ( .B(n1261), .A(n1262), .Z(n1260) );
XOR U2102 ( .A(c420), .B(b[420]), .Z(n1261) );
XNOR U2103 ( .A(b[420]), .B(n1262), .Z(c[420]) );
XNOR U2104 ( .A(a[420]), .B(c420), .Z(n1262) );
XOR U2105 ( .A(c421), .B(n1263), .Z(c422) );
ANDN U2106 ( .B(n1264), .A(n1265), .Z(n1263) );
XOR U2107 ( .A(c421), .B(b[421]), .Z(n1264) );
XNOR U2108 ( .A(b[421]), .B(n1265), .Z(c[421]) );
XNOR U2109 ( .A(a[421]), .B(c421), .Z(n1265) );
XOR U2110 ( .A(c422), .B(n1266), .Z(c423) );
ANDN U2111 ( .B(n1267), .A(n1268), .Z(n1266) );
XOR U2112 ( .A(c422), .B(b[422]), .Z(n1267) );
XNOR U2113 ( .A(b[422]), .B(n1268), .Z(c[422]) );
XNOR U2114 ( .A(a[422]), .B(c422), .Z(n1268) );
XOR U2115 ( .A(c423), .B(n1269), .Z(c424) );
ANDN U2116 ( .B(n1270), .A(n1271), .Z(n1269) );
XOR U2117 ( .A(c423), .B(b[423]), .Z(n1270) );
XNOR U2118 ( .A(b[423]), .B(n1271), .Z(c[423]) );
XNOR U2119 ( .A(a[423]), .B(c423), .Z(n1271) );
XOR U2120 ( .A(c424), .B(n1272), .Z(c425) );
ANDN U2121 ( .B(n1273), .A(n1274), .Z(n1272) );
XOR U2122 ( .A(c424), .B(b[424]), .Z(n1273) );
XNOR U2123 ( .A(b[424]), .B(n1274), .Z(c[424]) );
XNOR U2124 ( .A(a[424]), .B(c424), .Z(n1274) );
XOR U2125 ( .A(c425), .B(n1275), .Z(c426) );
ANDN U2126 ( .B(n1276), .A(n1277), .Z(n1275) );
XOR U2127 ( .A(c425), .B(b[425]), .Z(n1276) );
XNOR U2128 ( .A(b[425]), .B(n1277), .Z(c[425]) );
XNOR U2129 ( .A(a[425]), .B(c425), .Z(n1277) );
XOR U2130 ( .A(c426), .B(n1278), .Z(c427) );
ANDN U2131 ( .B(n1279), .A(n1280), .Z(n1278) );
XOR U2132 ( .A(c426), .B(b[426]), .Z(n1279) );
XNOR U2133 ( .A(b[426]), .B(n1280), .Z(c[426]) );
XNOR U2134 ( .A(a[426]), .B(c426), .Z(n1280) );
XOR U2135 ( .A(c427), .B(n1281), .Z(c428) );
ANDN U2136 ( .B(n1282), .A(n1283), .Z(n1281) );
XOR U2137 ( .A(c427), .B(b[427]), .Z(n1282) );
XNOR U2138 ( .A(b[427]), .B(n1283), .Z(c[427]) );
XNOR U2139 ( .A(a[427]), .B(c427), .Z(n1283) );
XOR U2140 ( .A(c428), .B(n1284), .Z(c429) );
ANDN U2141 ( .B(n1285), .A(n1286), .Z(n1284) );
XOR U2142 ( .A(c428), .B(b[428]), .Z(n1285) );
XNOR U2143 ( .A(b[428]), .B(n1286), .Z(c[428]) );
XNOR U2144 ( .A(a[428]), .B(c428), .Z(n1286) );
XOR U2145 ( .A(c429), .B(n1287), .Z(c430) );
ANDN U2146 ( .B(n1288), .A(n1289), .Z(n1287) );
XOR U2147 ( .A(c429), .B(b[429]), .Z(n1288) );
XNOR U2148 ( .A(b[429]), .B(n1289), .Z(c[429]) );
XNOR U2149 ( .A(a[429]), .B(c429), .Z(n1289) );
XOR U2150 ( .A(c430), .B(n1290), .Z(c431) );
ANDN U2151 ( .B(n1291), .A(n1292), .Z(n1290) );
XOR U2152 ( .A(c430), .B(b[430]), .Z(n1291) );
XNOR U2153 ( .A(b[430]), .B(n1292), .Z(c[430]) );
XNOR U2154 ( .A(a[430]), .B(c430), .Z(n1292) );
XOR U2155 ( .A(c431), .B(n1293), .Z(c432) );
ANDN U2156 ( .B(n1294), .A(n1295), .Z(n1293) );
XOR U2157 ( .A(c431), .B(b[431]), .Z(n1294) );
XNOR U2158 ( .A(b[431]), .B(n1295), .Z(c[431]) );
XNOR U2159 ( .A(a[431]), .B(c431), .Z(n1295) );
XOR U2160 ( .A(c432), .B(n1296), .Z(c433) );
ANDN U2161 ( .B(n1297), .A(n1298), .Z(n1296) );
XOR U2162 ( .A(c432), .B(b[432]), .Z(n1297) );
XNOR U2163 ( .A(b[432]), .B(n1298), .Z(c[432]) );
XNOR U2164 ( .A(a[432]), .B(c432), .Z(n1298) );
XOR U2165 ( .A(c433), .B(n1299), .Z(c434) );
ANDN U2166 ( .B(n1300), .A(n1301), .Z(n1299) );
XOR U2167 ( .A(c433), .B(b[433]), .Z(n1300) );
XNOR U2168 ( .A(b[433]), .B(n1301), .Z(c[433]) );
XNOR U2169 ( .A(a[433]), .B(c433), .Z(n1301) );
XOR U2170 ( .A(c434), .B(n1302), .Z(c435) );
ANDN U2171 ( .B(n1303), .A(n1304), .Z(n1302) );
XOR U2172 ( .A(c434), .B(b[434]), .Z(n1303) );
XNOR U2173 ( .A(b[434]), .B(n1304), .Z(c[434]) );
XNOR U2174 ( .A(a[434]), .B(c434), .Z(n1304) );
XOR U2175 ( .A(c435), .B(n1305), .Z(c436) );
ANDN U2176 ( .B(n1306), .A(n1307), .Z(n1305) );
XOR U2177 ( .A(c435), .B(b[435]), .Z(n1306) );
XNOR U2178 ( .A(b[435]), .B(n1307), .Z(c[435]) );
XNOR U2179 ( .A(a[435]), .B(c435), .Z(n1307) );
XOR U2180 ( .A(c436), .B(n1308), .Z(c437) );
ANDN U2181 ( .B(n1309), .A(n1310), .Z(n1308) );
XOR U2182 ( .A(c436), .B(b[436]), .Z(n1309) );
XNOR U2183 ( .A(b[436]), .B(n1310), .Z(c[436]) );
XNOR U2184 ( .A(a[436]), .B(c436), .Z(n1310) );
XOR U2185 ( .A(c437), .B(n1311), .Z(c438) );
ANDN U2186 ( .B(n1312), .A(n1313), .Z(n1311) );
XOR U2187 ( .A(c437), .B(b[437]), .Z(n1312) );
XNOR U2188 ( .A(b[437]), .B(n1313), .Z(c[437]) );
XNOR U2189 ( .A(a[437]), .B(c437), .Z(n1313) );
XOR U2190 ( .A(c438), .B(n1314), .Z(c439) );
ANDN U2191 ( .B(n1315), .A(n1316), .Z(n1314) );
XOR U2192 ( .A(c438), .B(b[438]), .Z(n1315) );
XNOR U2193 ( .A(b[438]), .B(n1316), .Z(c[438]) );
XNOR U2194 ( .A(a[438]), .B(c438), .Z(n1316) );
XOR U2195 ( .A(c439), .B(n1317), .Z(c440) );
ANDN U2196 ( .B(n1318), .A(n1319), .Z(n1317) );
XOR U2197 ( .A(c439), .B(b[439]), .Z(n1318) );
XNOR U2198 ( .A(b[439]), .B(n1319), .Z(c[439]) );
XNOR U2199 ( .A(a[439]), .B(c439), .Z(n1319) );
XOR U2200 ( .A(c440), .B(n1320), .Z(c441) );
ANDN U2201 ( .B(n1321), .A(n1322), .Z(n1320) );
XOR U2202 ( .A(c440), .B(b[440]), .Z(n1321) );
XNOR U2203 ( .A(b[440]), .B(n1322), .Z(c[440]) );
XNOR U2204 ( .A(a[440]), .B(c440), .Z(n1322) );
XOR U2205 ( .A(c441), .B(n1323), .Z(c442) );
ANDN U2206 ( .B(n1324), .A(n1325), .Z(n1323) );
XOR U2207 ( .A(c441), .B(b[441]), .Z(n1324) );
XNOR U2208 ( .A(b[441]), .B(n1325), .Z(c[441]) );
XNOR U2209 ( .A(a[441]), .B(c441), .Z(n1325) );
XOR U2210 ( .A(c442), .B(n1326), .Z(c443) );
ANDN U2211 ( .B(n1327), .A(n1328), .Z(n1326) );
XOR U2212 ( .A(c442), .B(b[442]), .Z(n1327) );
XNOR U2213 ( .A(b[442]), .B(n1328), .Z(c[442]) );
XNOR U2214 ( .A(a[442]), .B(c442), .Z(n1328) );
XOR U2215 ( .A(c443), .B(n1329), .Z(c444) );
ANDN U2216 ( .B(n1330), .A(n1331), .Z(n1329) );
XOR U2217 ( .A(c443), .B(b[443]), .Z(n1330) );
XNOR U2218 ( .A(b[443]), .B(n1331), .Z(c[443]) );
XNOR U2219 ( .A(a[443]), .B(c443), .Z(n1331) );
XOR U2220 ( .A(c444), .B(n1332), .Z(c445) );
ANDN U2221 ( .B(n1333), .A(n1334), .Z(n1332) );
XOR U2222 ( .A(c444), .B(b[444]), .Z(n1333) );
XNOR U2223 ( .A(b[444]), .B(n1334), .Z(c[444]) );
XNOR U2224 ( .A(a[444]), .B(c444), .Z(n1334) );
XOR U2225 ( .A(c445), .B(n1335), .Z(c446) );
ANDN U2226 ( .B(n1336), .A(n1337), .Z(n1335) );
XOR U2227 ( .A(c445), .B(b[445]), .Z(n1336) );
XNOR U2228 ( .A(b[445]), .B(n1337), .Z(c[445]) );
XNOR U2229 ( .A(a[445]), .B(c445), .Z(n1337) );
XOR U2230 ( .A(c446), .B(n1338), .Z(c447) );
ANDN U2231 ( .B(n1339), .A(n1340), .Z(n1338) );
XOR U2232 ( .A(c446), .B(b[446]), .Z(n1339) );
XNOR U2233 ( .A(b[446]), .B(n1340), .Z(c[446]) );
XNOR U2234 ( .A(a[446]), .B(c446), .Z(n1340) );
XOR U2235 ( .A(c447), .B(n1341), .Z(c448) );
ANDN U2236 ( .B(n1342), .A(n1343), .Z(n1341) );
XOR U2237 ( .A(c447), .B(b[447]), .Z(n1342) );
XNOR U2238 ( .A(b[447]), .B(n1343), .Z(c[447]) );
XNOR U2239 ( .A(a[447]), .B(c447), .Z(n1343) );
XOR U2240 ( .A(c448), .B(n1344), .Z(c449) );
ANDN U2241 ( .B(n1345), .A(n1346), .Z(n1344) );
XOR U2242 ( .A(c448), .B(b[448]), .Z(n1345) );
XNOR U2243 ( .A(b[448]), .B(n1346), .Z(c[448]) );
XNOR U2244 ( .A(a[448]), .B(c448), .Z(n1346) );
XOR U2245 ( .A(c449), .B(n1347), .Z(c450) );
ANDN U2246 ( .B(n1348), .A(n1349), .Z(n1347) );
XOR U2247 ( .A(c449), .B(b[449]), .Z(n1348) );
XNOR U2248 ( .A(b[449]), .B(n1349), .Z(c[449]) );
XNOR U2249 ( .A(a[449]), .B(c449), .Z(n1349) );
XOR U2250 ( .A(c450), .B(n1350), .Z(c451) );
ANDN U2251 ( .B(n1351), .A(n1352), .Z(n1350) );
XOR U2252 ( .A(c450), .B(b[450]), .Z(n1351) );
XNOR U2253 ( .A(b[450]), .B(n1352), .Z(c[450]) );
XNOR U2254 ( .A(a[450]), .B(c450), .Z(n1352) );
XOR U2255 ( .A(c451), .B(n1353), .Z(c452) );
ANDN U2256 ( .B(n1354), .A(n1355), .Z(n1353) );
XOR U2257 ( .A(c451), .B(b[451]), .Z(n1354) );
XNOR U2258 ( .A(b[451]), .B(n1355), .Z(c[451]) );
XNOR U2259 ( .A(a[451]), .B(c451), .Z(n1355) );
XOR U2260 ( .A(c452), .B(n1356), .Z(c453) );
ANDN U2261 ( .B(n1357), .A(n1358), .Z(n1356) );
XOR U2262 ( .A(c452), .B(b[452]), .Z(n1357) );
XNOR U2263 ( .A(b[452]), .B(n1358), .Z(c[452]) );
XNOR U2264 ( .A(a[452]), .B(c452), .Z(n1358) );
XOR U2265 ( .A(c453), .B(n1359), .Z(c454) );
ANDN U2266 ( .B(n1360), .A(n1361), .Z(n1359) );
XOR U2267 ( .A(c453), .B(b[453]), .Z(n1360) );
XNOR U2268 ( .A(b[453]), .B(n1361), .Z(c[453]) );
XNOR U2269 ( .A(a[453]), .B(c453), .Z(n1361) );
XOR U2270 ( .A(c454), .B(n1362), .Z(c455) );
ANDN U2271 ( .B(n1363), .A(n1364), .Z(n1362) );
XOR U2272 ( .A(c454), .B(b[454]), .Z(n1363) );
XNOR U2273 ( .A(b[454]), .B(n1364), .Z(c[454]) );
XNOR U2274 ( .A(a[454]), .B(c454), .Z(n1364) );
XOR U2275 ( .A(c455), .B(n1365), .Z(c456) );
ANDN U2276 ( .B(n1366), .A(n1367), .Z(n1365) );
XOR U2277 ( .A(c455), .B(b[455]), .Z(n1366) );
XNOR U2278 ( .A(b[455]), .B(n1367), .Z(c[455]) );
XNOR U2279 ( .A(a[455]), .B(c455), .Z(n1367) );
XOR U2280 ( .A(c456), .B(n1368), .Z(c457) );
ANDN U2281 ( .B(n1369), .A(n1370), .Z(n1368) );
XOR U2282 ( .A(c456), .B(b[456]), .Z(n1369) );
XNOR U2283 ( .A(b[456]), .B(n1370), .Z(c[456]) );
XNOR U2284 ( .A(a[456]), .B(c456), .Z(n1370) );
XOR U2285 ( .A(c457), .B(n1371), .Z(c458) );
ANDN U2286 ( .B(n1372), .A(n1373), .Z(n1371) );
XOR U2287 ( .A(c457), .B(b[457]), .Z(n1372) );
XNOR U2288 ( .A(b[457]), .B(n1373), .Z(c[457]) );
XNOR U2289 ( .A(a[457]), .B(c457), .Z(n1373) );
XOR U2290 ( .A(c458), .B(n1374), .Z(c459) );
ANDN U2291 ( .B(n1375), .A(n1376), .Z(n1374) );
XOR U2292 ( .A(c458), .B(b[458]), .Z(n1375) );
XNOR U2293 ( .A(b[458]), .B(n1376), .Z(c[458]) );
XNOR U2294 ( .A(a[458]), .B(c458), .Z(n1376) );
XOR U2295 ( .A(c459), .B(n1377), .Z(c460) );
ANDN U2296 ( .B(n1378), .A(n1379), .Z(n1377) );
XOR U2297 ( .A(c459), .B(b[459]), .Z(n1378) );
XNOR U2298 ( .A(b[459]), .B(n1379), .Z(c[459]) );
XNOR U2299 ( .A(a[459]), .B(c459), .Z(n1379) );
XOR U2300 ( .A(c460), .B(n1380), .Z(c461) );
ANDN U2301 ( .B(n1381), .A(n1382), .Z(n1380) );
XOR U2302 ( .A(c460), .B(b[460]), .Z(n1381) );
XNOR U2303 ( .A(b[460]), .B(n1382), .Z(c[460]) );
XNOR U2304 ( .A(a[460]), .B(c460), .Z(n1382) );
XOR U2305 ( .A(c461), .B(n1383), .Z(c462) );
ANDN U2306 ( .B(n1384), .A(n1385), .Z(n1383) );
XOR U2307 ( .A(c461), .B(b[461]), .Z(n1384) );
XNOR U2308 ( .A(b[461]), .B(n1385), .Z(c[461]) );
XNOR U2309 ( .A(a[461]), .B(c461), .Z(n1385) );
XOR U2310 ( .A(c462), .B(n1386), .Z(c463) );
ANDN U2311 ( .B(n1387), .A(n1388), .Z(n1386) );
XOR U2312 ( .A(c462), .B(b[462]), .Z(n1387) );
XNOR U2313 ( .A(b[462]), .B(n1388), .Z(c[462]) );
XNOR U2314 ( .A(a[462]), .B(c462), .Z(n1388) );
XOR U2315 ( .A(c463), .B(n1389), .Z(c464) );
ANDN U2316 ( .B(n1390), .A(n1391), .Z(n1389) );
XOR U2317 ( .A(c463), .B(b[463]), .Z(n1390) );
XNOR U2318 ( .A(b[463]), .B(n1391), .Z(c[463]) );
XNOR U2319 ( .A(a[463]), .B(c463), .Z(n1391) );
XOR U2320 ( .A(c464), .B(n1392), .Z(c465) );
ANDN U2321 ( .B(n1393), .A(n1394), .Z(n1392) );
XOR U2322 ( .A(c464), .B(b[464]), .Z(n1393) );
XNOR U2323 ( .A(b[464]), .B(n1394), .Z(c[464]) );
XNOR U2324 ( .A(a[464]), .B(c464), .Z(n1394) );
XOR U2325 ( .A(c465), .B(n1395), .Z(c466) );
ANDN U2326 ( .B(n1396), .A(n1397), .Z(n1395) );
XOR U2327 ( .A(c465), .B(b[465]), .Z(n1396) );
XNOR U2328 ( .A(b[465]), .B(n1397), .Z(c[465]) );
XNOR U2329 ( .A(a[465]), .B(c465), .Z(n1397) );
XOR U2330 ( .A(c466), .B(n1398), .Z(c467) );
ANDN U2331 ( .B(n1399), .A(n1400), .Z(n1398) );
XOR U2332 ( .A(c466), .B(b[466]), .Z(n1399) );
XNOR U2333 ( .A(b[466]), .B(n1400), .Z(c[466]) );
XNOR U2334 ( .A(a[466]), .B(c466), .Z(n1400) );
XOR U2335 ( .A(c467), .B(n1401), .Z(c468) );
ANDN U2336 ( .B(n1402), .A(n1403), .Z(n1401) );
XOR U2337 ( .A(c467), .B(b[467]), .Z(n1402) );
XNOR U2338 ( .A(b[467]), .B(n1403), .Z(c[467]) );
XNOR U2339 ( .A(a[467]), .B(c467), .Z(n1403) );
XOR U2340 ( .A(c468), .B(n1404), .Z(c469) );
ANDN U2341 ( .B(n1405), .A(n1406), .Z(n1404) );
XOR U2342 ( .A(c468), .B(b[468]), .Z(n1405) );
XNOR U2343 ( .A(b[468]), .B(n1406), .Z(c[468]) );
XNOR U2344 ( .A(a[468]), .B(c468), .Z(n1406) );
XOR U2345 ( .A(c469), .B(n1407), .Z(c470) );
ANDN U2346 ( .B(n1408), .A(n1409), .Z(n1407) );
XOR U2347 ( .A(c469), .B(b[469]), .Z(n1408) );
XNOR U2348 ( .A(b[469]), .B(n1409), .Z(c[469]) );
XNOR U2349 ( .A(a[469]), .B(c469), .Z(n1409) );
XOR U2350 ( .A(c470), .B(n1410), .Z(c471) );
ANDN U2351 ( .B(n1411), .A(n1412), .Z(n1410) );
XOR U2352 ( .A(c470), .B(b[470]), .Z(n1411) );
XNOR U2353 ( .A(b[470]), .B(n1412), .Z(c[470]) );
XNOR U2354 ( .A(a[470]), .B(c470), .Z(n1412) );
XOR U2355 ( .A(c471), .B(n1413), .Z(c472) );
ANDN U2356 ( .B(n1414), .A(n1415), .Z(n1413) );
XOR U2357 ( .A(c471), .B(b[471]), .Z(n1414) );
XNOR U2358 ( .A(b[471]), .B(n1415), .Z(c[471]) );
XNOR U2359 ( .A(a[471]), .B(c471), .Z(n1415) );
XOR U2360 ( .A(c472), .B(n1416), .Z(c473) );
ANDN U2361 ( .B(n1417), .A(n1418), .Z(n1416) );
XOR U2362 ( .A(c472), .B(b[472]), .Z(n1417) );
XNOR U2363 ( .A(b[472]), .B(n1418), .Z(c[472]) );
XNOR U2364 ( .A(a[472]), .B(c472), .Z(n1418) );
XOR U2365 ( .A(c473), .B(n1419), .Z(c474) );
ANDN U2366 ( .B(n1420), .A(n1421), .Z(n1419) );
XOR U2367 ( .A(c473), .B(b[473]), .Z(n1420) );
XNOR U2368 ( .A(b[473]), .B(n1421), .Z(c[473]) );
XNOR U2369 ( .A(a[473]), .B(c473), .Z(n1421) );
XOR U2370 ( .A(c474), .B(n1422), .Z(c475) );
ANDN U2371 ( .B(n1423), .A(n1424), .Z(n1422) );
XOR U2372 ( .A(c474), .B(b[474]), .Z(n1423) );
XNOR U2373 ( .A(b[474]), .B(n1424), .Z(c[474]) );
XNOR U2374 ( .A(a[474]), .B(c474), .Z(n1424) );
XOR U2375 ( .A(c475), .B(n1425), .Z(c476) );
ANDN U2376 ( .B(n1426), .A(n1427), .Z(n1425) );
XOR U2377 ( .A(c475), .B(b[475]), .Z(n1426) );
XNOR U2378 ( .A(b[475]), .B(n1427), .Z(c[475]) );
XNOR U2379 ( .A(a[475]), .B(c475), .Z(n1427) );
XOR U2380 ( .A(c476), .B(n1428), .Z(c477) );
ANDN U2381 ( .B(n1429), .A(n1430), .Z(n1428) );
XOR U2382 ( .A(c476), .B(b[476]), .Z(n1429) );
XNOR U2383 ( .A(b[476]), .B(n1430), .Z(c[476]) );
XNOR U2384 ( .A(a[476]), .B(c476), .Z(n1430) );
XOR U2385 ( .A(c477), .B(n1431), .Z(c478) );
ANDN U2386 ( .B(n1432), .A(n1433), .Z(n1431) );
XOR U2387 ( .A(c477), .B(b[477]), .Z(n1432) );
XNOR U2388 ( .A(b[477]), .B(n1433), .Z(c[477]) );
XNOR U2389 ( .A(a[477]), .B(c477), .Z(n1433) );
XOR U2390 ( .A(c478), .B(n1434), .Z(c479) );
ANDN U2391 ( .B(n1435), .A(n1436), .Z(n1434) );
XOR U2392 ( .A(c478), .B(b[478]), .Z(n1435) );
XNOR U2393 ( .A(b[478]), .B(n1436), .Z(c[478]) );
XNOR U2394 ( .A(a[478]), .B(c478), .Z(n1436) );
XOR U2395 ( .A(c479), .B(n1437), .Z(c480) );
ANDN U2396 ( .B(n1438), .A(n1439), .Z(n1437) );
XOR U2397 ( .A(c479), .B(b[479]), .Z(n1438) );
XNOR U2398 ( .A(b[479]), .B(n1439), .Z(c[479]) );
XNOR U2399 ( .A(a[479]), .B(c479), .Z(n1439) );
XOR U2400 ( .A(c480), .B(n1440), .Z(c481) );
ANDN U2401 ( .B(n1441), .A(n1442), .Z(n1440) );
XOR U2402 ( .A(c480), .B(b[480]), .Z(n1441) );
XNOR U2403 ( .A(b[480]), .B(n1442), .Z(c[480]) );
XNOR U2404 ( .A(a[480]), .B(c480), .Z(n1442) );
XOR U2405 ( .A(c481), .B(n1443), .Z(c482) );
ANDN U2406 ( .B(n1444), .A(n1445), .Z(n1443) );
XOR U2407 ( .A(c481), .B(b[481]), .Z(n1444) );
XNOR U2408 ( .A(b[481]), .B(n1445), .Z(c[481]) );
XNOR U2409 ( .A(a[481]), .B(c481), .Z(n1445) );
XOR U2410 ( .A(c482), .B(n1446), .Z(c483) );
ANDN U2411 ( .B(n1447), .A(n1448), .Z(n1446) );
XOR U2412 ( .A(c482), .B(b[482]), .Z(n1447) );
XNOR U2413 ( .A(b[482]), .B(n1448), .Z(c[482]) );
XNOR U2414 ( .A(a[482]), .B(c482), .Z(n1448) );
XOR U2415 ( .A(c483), .B(n1449), .Z(c484) );
ANDN U2416 ( .B(n1450), .A(n1451), .Z(n1449) );
XOR U2417 ( .A(c483), .B(b[483]), .Z(n1450) );
XNOR U2418 ( .A(b[483]), .B(n1451), .Z(c[483]) );
XNOR U2419 ( .A(a[483]), .B(c483), .Z(n1451) );
XOR U2420 ( .A(c484), .B(n1452), .Z(c485) );
ANDN U2421 ( .B(n1453), .A(n1454), .Z(n1452) );
XOR U2422 ( .A(c484), .B(b[484]), .Z(n1453) );
XNOR U2423 ( .A(b[484]), .B(n1454), .Z(c[484]) );
XNOR U2424 ( .A(a[484]), .B(c484), .Z(n1454) );
XOR U2425 ( .A(c485), .B(n1455), .Z(c486) );
ANDN U2426 ( .B(n1456), .A(n1457), .Z(n1455) );
XOR U2427 ( .A(c485), .B(b[485]), .Z(n1456) );
XNOR U2428 ( .A(b[485]), .B(n1457), .Z(c[485]) );
XNOR U2429 ( .A(a[485]), .B(c485), .Z(n1457) );
XOR U2430 ( .A(c486), .B(n1458), .Z(c487) );
ANDN U2431 ( .B(n1459), .A(n1460), .Z(n1458) );
XOR U2432 ( .A(c486), .B(b[486]), .Z(n1459) );
XNOR U2433 ( .A(b[486]), .B(n1460), .Z(c[486]) );
XNOR U2434 ( .A(a[486]), .B(c486), .Z(n1460) );
XOR U2435 ( .A(c487), .B(n1461), .Z(c488) );
ANDN U2436 ( .B(n1462), .A(n1463), .Z(n1461) );
XOR U2437 ( .A(c487), .B(b[487]), .Z(n1462) );
XNOR U2438 ( .A(b[487]), .B(n1463), .Z(c[487]) );
XNOR U2439 ( .A(a[487]), .B(c487), .Z(n1463) );
XOR U2440 ( .A(c488), .B(n1464), .Z(c489) );
ANDN U2441 ( .B(n1465), .A(n1466), .Z(n1464) );
XOR U2442 ( .A(c488), .B(b[488]), .Z(n1465) );
XNOR U2443 ( .A(b[488]), .B(n1466), .Z(c[488]) );
XNOR U2444 ( .A(a[488]), .B(c488), .Z(n1466) );
XOR U2445 ( .A(c489), .B(n1467), .Z(c490) );
ANDN U2446 ( .B(n1468), .A(n1469), .Z(n1467) );
XOR U2447 ( .A(c489), .B(b[489]), .Z(n1468) );
XNOR U2448 ( .A(b[489]), .B(n1469), .Z(c[489]) );
XNOR U2449 ( .A(a[489]), .B(c489), .Z(n1469) );
XOR U2450 ( .A(c490), .B(n1470), .Z(c491) );
ANDN U2451 ( .B(n1471), .A(n1472), .Z(n1470) );
XOR U2452 ( .A(c490), .B(b[490]), .Z(n1471) );
XNOR U2453 ( .A(b[490]), .B(n1472), .Z(c[490]) );
XNOR U2454 ( .A(a[490]), .B(c490), .Z(n1472) );
XOR U2455 ( .A(c491), .B(n1473), .Z(c492) );
ANDN U2456 ( .B(n1474), .A(n1475), .Z(n1473) );
XOR U2457 ( .A(c491), .B(b[491]), .Z(n1474) );
XNOR U2458 ( .A(b[491]), .B(n1475), .Z(c[491]) );
XNOR U2459 ( .A(a[491]), .B(c491), .Z(n1475) );
XOR U2460 ( .A(c492), .B(n1476), .Z(c493) );
ANDN U2461 ( .B(n1477), .A(n1478), .Z(n1476) );
XOR U2462 ( .A(c492), .B(b[492]), .Z(n1477) );
XNOR U2463 ( .A(b[492]), .B(n1478), .Z(c[492]) );
XNOR U2464 ( .A(a[492]), .B(c492), .Z(n1478) );
XOR U2465 ( .A(c493), .B(n1479), .Z(c494) );
ANDN U2466 ( .B(n1480), .A(n1481), .Z(n1479) );
XOR U2467 ( .A(c493), .B(b[493]), .Z(n1480) );
XNOR U2468 ( .A(b[493]), .B(n1481), .Z(c[493]) );
XNOR U2469 ( .A(a[493]), .B(c493), .Z(n1481) );
XOR U2470 ( .A(c494), .B(n1482), .Z(c495) );
ANDN U2471 ( .B(n1483), .A(n1484), .Z(n1482) );
XOR U2472 ( .A(c494), .B(b[494]), .Z(n1483) );
XNOR U2473 ( .A(b[494]), .B(n1484), .Z(c[494]) );
XNOR U2474 ( .A(a[494]), .B(c494), .Z(n1484) );
XOR U2475 ( .A(c495), .B(n1485), .Z(c496) );
ANDN U2476 ( .B(n1486), .A(n1487), .Z(n1485) );
XOR U2477 ( .A(c495), .B(b[495]), .Z(n1486) );
XNOR U2478 ( .A(b[495]), .B(n1487), .Z(c[495]) );
XNOR U2479 ( .A(a[495]), .B(c495), .Z(n1487) );
XOR U2480 ( .A(c496), .B(n1488), .Z(c497) );
ANDN U2481 ( .B(n1489), .A(n1490), .Z(n1488) );
XOR U2482 ( .A(c496), .B(b[496]), .Z(n1489) );
XNOR U2483 ( .A(b[496]), .B(n1490), .Z(c[496]) );
XNOR U2484 ( .A(a[496]), .B(c496), .Z(n1490) );
XOR U2485 ( .A(c497), .B(n1491), .Z(c498) );
ANDN U2486 ( .B(n1492), .A(n1493), .Z(n1491) );
XOR U2487 ( .A(c497), .B(b[497]), .Z(n1492) );
XNOR U2488 ( .A(b[497]), .B(n1493), .Z(c[497]) );
XNOR U2489 ( .A(a[497]), .B(c497), .Z(n1493) );
XOR U2490 ( .A(c498), .B(n1494), .Z(c499) );
ANDN U2491 ( .B(n1495), .A(n1496), .Z(n1494) );
XOR U2492 ( .A(c498), .B(b[498]), .Z(n1495) );
XNOR U2493 ( .A(b[498]), .B(n1496), .Z(c[498]) );
XNOR U2494 ( .A(a[498]), .B(c498), .Z(n1496) );
XOR U2495 ( .A(c499), .B(n1497), .Z(c500) );
ANDN U2496 ( .B(n1498), .A(n1499), .Z(n1497) );
XOR U2497 ( .A(c499), .B(b[499]), .Z(n1498) );
XNOR U2498 ( .A(b[499]), .B(n1499), .Z(c[499]) );
XNOR U2499 ( .A(a[499]), .B(c499), .Z(n1499) );
XOR U2500 ( .A(c500), .B(n1500), .Z(c501) );
ANDN U2501 ( .B(n1501), .A(n1502), .Z(n1500) );
XOR U2502 ( .A(c500), .B(b[500]), .Z(n1501) );
XNOR U2503 ( .A(b[500]), .B(n1502), .Z(c[500]) );
XNOR U2504 ( .A(a[500]), .B(c500), .Z(n1502) );
XOR U2505 ( .A(c501), .B(n1503), .Z(c502) );
ANDN U2506 ( .B(n1504), .A(n1505), .Z(n1503) );
XOR U2507 ( .A(c501), .B(b[501]), .Z(n1504) );
XNOR U2508 ( .A(b[501]), .B(n1505), .Z(c[501]) );
XNOR U2509 ( .A(a[501]), .B(c501), .Z(n1505) );
XOR U2510 ( .A(c502), .B(n1506), .Z(c503) );
ANDN U2511 ( .B(n1507), .A(n1508), .Z(n1506) );
XOR U2512 ( .A(c502), .B(b[502]), .Z(n1507) );
XNOR U2513 ( .A(b[502]), .B(n1508), .Z(c[502]) );
XNOR U2514 ( .A(a[502]), .B(c502), .Z(n1508) );
XOR U2515 ( .A(c503), .B(n1509), .Z(c504) );
ANDN U2516 ( .B(n1510), .A(n1511), .Z(n1509) );
XOR U2517 ( .A(c503), .B(b[503]), .Z(n1510) );
XNOR U2518 ( .A(b[503]), .B(n1511), .Z(c[503]) );
XNOR U2519 ( .A(a[503]), .B(c503), .Z(n1511) );
XOR U2520 ( .A(c504), .B(n1512), .Z(c505) );
ANDN U2521 ( .B(n1513), .A(n1514), .Z(n1512) );
XOR U2522 ( .A(c504), .B(b[504]), .Z(n1513) );
XNOR U2523 ( .A(b[504]), .B(n1514), .Z(c[504]) );
XNOR U2524 ( .A(a[504]), .B(c504), .Z(n1514) );
XOR U2525 ( .A(c505), .B(n1515), .Z(c506) );
ANDN U2526 ( .B(n1516), .A(n1517), .Z(n1515) );
XOR U2527 ( .A(c505), .B(b[505]), .Z(n1516) );
XNOR U2528 ( .A(b[505]), .B(n1517), .Z(c[505]) );
XNOR U2529 ( .A(a[505]), .B(c505), .Z(n1517) );
XOR U2530 ( .A(c506), .B(n1518), .Z(c507) );
ANDN U2531 ( .B(n1519), .A(n1520), .Z(n1518) );
XOR U2532 ( .A(c506), .B(b[506]), .Z(n1519) );
XNOR U2533 ( .A(b[506]), .B(n1520), .Z(c[506]) );
XNOR U2534 ( .A(a[506]), .B(c506), .Z(n1520) );
XOR U2535 ( .A(c507), .B(n1521), .Z(c508) );
ANDN U2536 ( .B(n1522), .A(n1523), .Z(n1521) );
XOR U2537 ( .A(c507), .B(b[507]), .Z(n1522) );
XNOR U2538 ( .A(b[507]), .B(n1523), .Z(c[507]) );
XNOR U2539 ( .A(a[507]), .B(c507), .Z(n1523) );
XOR U2540 ( .A(c508), .B(n1524), .Z(c509) );
ANDN U2541 ( .B(n1525), .A(n1526), .Z(n1524) );
XOR U2542 ( .A(c508), .B(b[508]), .Z(n1525) );
XNOR U2543 ( .A(b[508]), .B(n1526), .Z(c[508]) );
XNOR U2544 ( .A(a[508]), .B(c508), .Z(n1526) );
XOR U2545 ( .A(c509), .B(n1527), .Z(c510) );
ANDN U2546 ( .B(n1528), .A(n1529), .Z(n1527) );
XOR U2547 ( .A(c509), .B(b[509]), .Z(n1528) );
XNOR U2548 ( .A(b[509]), .B(n1529), .Z(c[509]) );
XNOR U2549 ( .A(a[509]), .B(c509), .Z(n1529) );
XOR U2550 ( .A(c510), .B(n1530), .Z(c511) );
ANDN U2551 ( .B(n1531), .A(n1532), .Z(n1530) );
XOR U2552 ( .A(c510), .B(b[510]), .Z(n1531) );
XNOR U2553 ( .A(b[510]), .B(n1532), .Z(c[510]) );
XNOR U2554 ( .A(a[510]), .B(c510), .Z(n1532) );
XOR U2555 ( .A(c511), .B(n1533), .Z(c512) );
ANDN U2556 ( .B(n1534), .A(n1535), .Z(n1533) );
XOR U2557 ( .A(c511), .B(b[511]), .Z(n1534) );
XNOR U2558 ( .A(b[511]), .B(n1535), .Z(c[511]) );
XNOR U2559 ( .A(a[511]), .B(c511), .Z(n1535) );
XOR U2560 ( .A(c512), .B(n1536), .Z(c513) );
ANDN U2561 ( .B(n1537), .A(n1538), .Z(n1536) );
XOR U2562 ( .A(c512), .B(b[512]), .Z(n1537) );
XNOR U2563 ( .A(b[512]), .B(n1538), .Z(c[512]) );
XNOR U2564 ( .A(a[512]), .B(c512), .Z(n1538) );
XOR U2565 ( .A(c513), .B(n1539), .Z(c514) );
ANDN U2566 ( .B(n1540), .A(n1541), .Z(n1539) );
XOR U2567 ( .A(c513), .B(b[513]), .Z(n1540) );
XNOR U2568 ( .A(b[513]), .B(n1541), .Z(c[513]) );
XNOR U2569 ( .A(a[513]), .B(c513), .Z(n1541) );
XOR U2570 ( .A(c514), .B(n1542), .Z(c515) );
ANDN U2571 ( .B(n1543), .A(n1544), .Z(n1542) );
XOR U2572 ( .A(c514), .B(b[514]), .Z(n1543) );
XNOR U2573 ( .A(b[514]), .B(n1544), .Z(c[514]) );
XNOR U2574 ( .A(a[514]), .B(c514), .Z(n1544) );
XOR U2575 ( .A(c515), .B(n1545), .Z(c516) );
ANDN U2576 ( .B(n1546), .A(n1547), .Z(n1545) );
XOR U2577 ( .A(c515), .B(b[515]), .Z(n1546) );
XNOR U2578 ( .A(b[515]), .B(n1547), .Z(c[515]) );
XNOR U2579 ( .A(a[515]), .B(c515), .Z(n1547) );
XOR U2580 ( .A(c516), .B(n1548), .Z(c517) );
ANDN U2581 ( .B(n1549), .A(n1550), .Z(n1548) );
XOR U2582 ( .A(c516), .B(b[516]), .Z(n1549) );
XNOR U2583 ( .A(b[516]), .B(n1550), .Z(c[516]) );
XNOR U2584 ( .A(a[516]), .B(c516), .Z(n1550) );
XOR U2585 ( .A(c517), .B(n1551), .Z(c518) );
ANDN U2586 ( .B(n1552), .A(n1553), .Z(n1551) );
XOR U2587 ( .A(c517), .B(b[517]), .Z(n1552) );
XNOR U2588 ( .A(b[517]), .B(n1553), .Z(c[517]) );
XNOR U2589 ( .A(a[517]), .B(c517), .Z(n1553) );
XOR U2590 ( .A(c518), .B(n1554), .Z(c519) );
ANDN U2591 ( .B(n1555), .A(n1556), .Z(n1554) );
XOR U2592 ( .A(c518), .B(b[518]), .Z(n1555) );
XNOR U2593 ( .A(b[518]), .B(n1556), .Z(c[518]) );
XNOR U2594 ( .A(a[518]), .B(c518), .Z(n1556) );
XOR U2595 ( .A(c519), .B(n1557), .Z(c520) );
ANDN U2596 ( .B(n1558), .A(n1559), .Z(n1557) );
XOR U2597 ( .A(c519), .B(b[519]), .Z(n1558) );
XNOR U2598 ( .A(b[519]), .B(n1559), .Z(c[519]) );
XNOR U2599 ( .A(a[519]), .B(c519), .Z(n1559) );
XOR U2600 ( .A(c520), .B(n1560), .Z(c521) );
ANDN U2601 ( .B(n1561), .A(n1562), .Z(n1560) );
XOR U2602 ( .A(c520), .B(b[520]), .Z(n1561) );
XNOR U2603 ( .A(b[520]), .B(n1562), .Z(c[520]) );
XNOR U2604 ( .A(a[520]), .B(c520), .Z(n1562) );
XOR U2605 ( .A(c521), .B(n1563), .Z(c522) );
ANDN U2606 ( .B(n1564), .A(n1565), .Z(n1563) );
XOR U2607 ( .A(c521), .B(b[521]), .Z(n1564) );
XNOR U2608 ( .A(b[521]), .B(n1565), .Z(c[521]) );
XNOR U2609 ( .A(a[521]), .B(c521), .Z(n1565) );
XOR U2610 ( .A(c522), .B(n1566), .Z(c523) );
ANDN U2611 ( .B(n1567), .A(n1568), .Z(n1566) );
XOR U2612 ( .A(c522), .B(b[522]), .Z(n1567) );
XNOR U2613 ( .A(b[522]), .B(n1568), .Z(c[522]) );
XNOR U2614 ( .A(a[522]), .B(c522), .Z(n1568) );
XOR U2615 ( .A(c523), .B(n1569), .Z(c524) );
ANDN U2616 ( .B(n1570), .A(n1571), .Z(n1569) );
XOR U2617 ( .A(c523), .B(b[523]), .Z(n1570) );
XNOR U2618 ( .A(b[523]), .B(n1571), .Z(c[523]) );
XNOR U2619 ( .A(a[523]), .B(c523), .Z(n1571) );
XOR U2620 ( .A(c524), .B(n1572), .Z(c525) );
ANDN U2621 ( .B(n1573), .A(n1574), .Z(n1572) );
XOR U2622 ( .A(c524), .B(b[524]), .Z(n1573) );
XNOR U2623 ( .A(b[524]), .B(n1574), .Z(c[524]) );
XNOR U2624 ( .A(a[524]), .B(c524), .Z(n1574) );
XOR U2625 ( .A(c525), .B(n1575), .Z(c526) );
ANDN U2626 ( .B(n1576), .A(n1577), .Z(n1575) );
XOR U2627 ( .A(c525), .B(b[525]), .Z(n1576) );
XNOR U2628 ( .A(b[525]), .B(n1577), .Z(c[525]) );
XNOR U2629 ( .A(a[525]), .B(c525), .Z(n1577) );
XOR U2630 ( .A(c526), .B(n1578), .Z(c527) );
ANDN U2631 ( .B(n1579), .A(n1580), .Z(n1578) );
XOR U2632 ( .A(c526), .B(b[526]), .Z(n1579) );
XNOR U2633 ( .A(b[526]), .B(n1580), .Z(c[526]) );
XNOR U2634 ( .A(a[526]), .B(c526), .Z(n1580) );
XOR U2635 ( .A(c527), .B(n1581), .Z(c528) );
ANDN U2636 ( .B(n1582), .A(n1583), .Z(n1581) );
XOR U2637 ( .A(c527), .B(b[527]), .Z(n1582) );
XNOR U2638 ( .A(b[527]), .B(n1583), .Z(c[527]) );
XNOR U2639 ( .A(a[527]), .B(c527), .Z(n1583) );
XOR U2640 ( .A(c528), .B(n1584), .Z(c529) );
ANDN U2641 ( .B(n1585), .A(n1586), .Z(n1584) );
XOR U2642 ( .A(c528), .B(b[528]), .Z(n1585) );
XNOR U2643 ( .A(b[528]), .B(n1586), .Z(c[528]) );
XNOR U2644 ( .A(a[528]), .B(c528), .Z(n1586) );
XOR U2645 ( .A(c529), .B(n1587), .Z(c530) );
ANDN U2646 ( .B(n1588), .A(n1589), .Z(n1587) );
XOR U2647 ( .A(c529), .B(b[529]), .Z(n1588) );
XNOR U2648 ( .A(b[529]), .B(n1589), .Z(c[529]) );
XNOR U2649 ( .A(a[529]), .B(c529), .Z(n1589) );
XOR U2650 ( .A(c530), .B(n1590), .Z(c531) );
ANDN U2651 ( .B(n1591), .A(n1592), .Z(n1590) );
XOR U2652 ( .A(c530), .B(b[530]), .Z(n1591) );
XNOR U2653 ( .A(b[530]), .B(n1592), .Z(c[530]) );
XNOR U2654 ( .A(a[530]), .B(c530), .Z(n1592) );
XOR U2655 ( .A(c531), .B(n1593), .Z(c532) );
ANDN U2656 ( .B(n1594), .A(n1595), .Z(n1593) );
XOR U2657 ( .A(c531), .B(b[531]), .Z(n1594) );
XNOR U2658 ( .A(b[531]), .B(n1595), .Z(c[531]) );
XNOR U2659 ( .A(a[531]), .B(c531), .Z(n1595) );
XOR U2660 ( .A(c532), .B(n1596), .Z(c533) );
ANDN U2661 ( .B(n1597), .A(n1598), .Z(n1596) );
XOR U2662 ( .A(c532), .B(b[532]), .Z(n1597) );
XNOR U2663 ( .A(b[532]), .B(n1598), .Z(c[532]) );
XNOR U2664 ( .A(a[532]), .B(c532), .Z(n1598) );
XOR U2665 ( .A(c533), .B(n1599), .Z(c534) );
ANDN U2666 ( .B(n1600), .A(n1601), .Z(n1599) );
XOR U2667 ( .A(c533), .B(b[533]), .Z(n1600) );
XNOR U2668 ( .A(b[533]), .B(n1601), .Z(c[533]) );
XNOR U2669 ( .A(a[533]), .B(c533), .Z(n1601) );
XOR U2670 ( .A(c534), .B(n1602), .Z(c535) );
ANDN U2671 ( .B(n1603), .A(n1604), .Z(n1602) );
XOR U2672 ( .A(c534), .B(b[534]), .Z(n1603) );
XNOR U2673 ( .A(b[534]), .B(n1604), .Z(c[534]) );
XNOR U2674 ( .A(a[534]), .B(c534), .Z(n1604) );
XOR U2675 ( .A(c535), .B(n1605), .Z(c536) );
ANDN U2676 ( .B(n1606), .A(n1607), .Z(n1605) );
XOR U2677 ( .A(c535), .B(b[535]), .Z(n1606) );
XNOR U2678 ( .A(b[535]), .B(n1607), .Z(c[535]) );
XNOR U2679 ( .A(a[535]), .B(c535), .Z(n1607) );
XOR U2680 ( .A(c536), .B(n1608), .Z(c537) );
ANDN U2681 ( .B(n1609), .A(n1610), .Z(n1608) );
XOR U2682 ( .A(c536), .B(b[536]), .Z(n1609) );
XNOR U2683 ( .A(b[536]), .B(n1610), .Z(c[536]) );
XNOR U2684 ( .A(a[536]), .B(c536), .Z(n1610) );
XOR U2685 ( .A(c537), .B(n1611), .Z(c538) );
ANDN U2686 ( .B(n1612), .A(n1613), .Z(n1611) );
XOR U2687 ( .A(c537), .B(b[537]), .Z(n1612) );
XNOR U2688 ( .A(b[537]), .B(n1613), .Z(c[537]) );
XNOR U2689 ( .A(a[537]), .B(c537), .Z(n1613) );
XOR U2690 ( .A(c538), .B(n1614), .Z(c539) );
ANDN U2691 ( .B(n1615), .A(n1616), .Z(n1614) );
XOR U2692 ( .A(c538), .B(b[538]), .Z(n1615) );
XNOR U2693 ( .A(b[538]), .B(n1616), .Z(c[538]) );
XNOR U2694 ( .A(a[538]), .B(c538), .Z(n1616) );
XOR U2695 ( .A(c539), .B(n1617), .Z(c540) );
ANDN U2696 ( .B(n1618), .A(n1619), .Z(n1617) );
XOR U2697 ( .A(c539), .B(b[539]), .Z(n1618) );
XNOR U2698 ( .A(b[539]), .B(n1619), .Z(c[539]) );
XNOR U2699 ( .A(a[539]), .B(c539), .Z(n1619) );
XOR U2700 ( .A(c540), .B(n1620), .Z(c541) );
ANDN U2701 ( .B(n1621), .A(n1622), .Z(n1620) );
XOR U2702 ( .A(c540), .B(b[540]), .Z(n1621) );
XNOR U2703 ( .A(b[540]), .B(n1622), .Z(c[540]) );
XNOR U2704 ( .A(a[540]), .B(c540), .Z(n1622) );
XOR U2705 ( .A(c541), .B(n1623), .Z(c542) );
ANDN U2706 ( .B(n1624), .A(n1625), .Z(n1623) );
XOR U2707 ( .A(c541), .B(b[541]), .Z(n1624) );
XNOR U2708 ( .A(b[541]), .B(n1625), .Z(c[541]) );
XNOR U2709 ( .A(a[541]), .B(c541), .Z(n1625) );
XOR U2710 ( .A(c542), .B(n1626), .Z(c543) );
ANDN U2711 ( .B(n1627), .A(n1628), .Z(n1626) );
XOR U2712 ( .A(c542), .B(b[542]), .Z(n1627) );
XNOR U2713 ( .A(b[542]), .B(n1628), .Z(c[542]) );
XNOR U2714 ( .A(a[542]), .B(c542), .Z(n1628) );
XOR U2715 ( .A(c543), .B(n1629), .Z(c544) );
ANDN U2716 ( .B(n1630), .A(n1631), .Z(n1629) );
XOR U2717 ( .A(c543), .B(b[543]), .Z(n1630) );
XNOR U2718 ( .A(b[543]), .B(n1631), .Z(c[543]) );
XNOR U2719 ( .A(a[543]), .B(c543), .Z(n1631) );
XOR U2720 ( .A(c544), .B(n1632), .Z(c545) );
ANDN U2721 ( .B(n1633), .A(n1634), .Z(n1632) );
XOR U2722 ( .A(c544), .B(b[544]), .Z(n1633) );
XNOR U2723 ( .A(b[544]), .B(n1634), .Z(c[544]) );
XNOR U2724 ( .A(a[544]), .B(c544), .Z(n1634) );
XOR U2725 ( .A(c545), .B(n1635), .Z(c546) );
ANDN U2726 ( .B(n1636), .A(n1637), .Z(n1635) );
XOR U2727 ( .A(c545), .B(b[545]), .Z(n1636) );
XNOR U2728 ( .A(b[545]), .B(n1637), .Z(c[545]) );
XNOR U2729 ( .A(a[545]), .B(c545), .Z(n1637) );
XOR U2730 ( .A(c546), .B(n1638), .Z(c547) );
ANDN U2731 ( .B(n1639), .A(n1640), .Z(n1638) );
XOR U2732 ( .A(c546), .B(b[546]), .Z(n1639) );
XNOR U2733 ( .A(b[546]), .B(n1640), .Z(c[546]) );
XNOR U2734 ( .A(a[546]), .B(c546), .Z(n1640) );
XOR U2735 ( .A(c547), .B(n1641), .Z(c548) );
ANDN U2736 ( .B(n1642), .A(n1643), .Z(n1641) );
XOR U2737 ( .A(c547), .B(b[547]), .Z(n1642) );
XNOR U2738 ( .A(b[547]), .B(n1643), .Z(c[547]) );
XNOR U2739 ( .A(a[547]), .B(c547), .Z(n1643) );
XOR U2740 ( .A(c548), .B(n1644), .Z(c549) );
ANDN U2741 ( .B(n1645), .A(n1646), .Z(n1644) );
XOR U2742 ( .A(c548), .B(b[548]), .Z(n1645) );
XNOR U2743 ( .A(b[548]), .B(n1646), .Z(c[548]) );
XNOR U2744 ( .A(a[548]), .B(c548), .Z(n1646) );
XOR U2745 ( .A(c549), .B(n1647), .Z(c550) );
ANDN U2746 ( .B(n1648), .A(n1649), .Z(n1647) );
XOR U2747 ( .A(c549), .B(b[549]), .Z(n1648) );
XNOR U2748 ( .A(b[549]), .B(n1649), .Z(c[549]) );
XNOR U2749 ( .A(a[549]), .B(c549), .Z(n1649) );
XOR U2750 ( .A(c550), .B(n1650), .Z(c551) );
ANDN U2751 ( .B(n1651), .A(n1652), .Z(n1650) );
XOR U2752 ( .A(c550), .B(b[550]), .Z(n1651) );
XNOR U2753 ( .A(b[550]), .B(n1652), .Z(c[550]) );
XNOR U2754 ( .A(a[550]), .B(c550), .Z(n1652) );
XOR U2755 ( .A(c551), .B(n1653), .Z(c552) );
ANDN U2756 ( .B(n1654), .A(n1655), .Z(n1653) );
XOR U2757 ( .A(c551), .B(b[551]), .Z(n1654) );
XNOR U2758 ( .A(b[551]), .B(n1655), .Z(c[551]) );
XNOR U2759 ( .A(a[551]), .B(c551), .Z(n1655) );
XOR U2760 ( .A(c552), .B(n1656), .Z(c553) );
ANDN U2761 ( .B(n1657), .A(n1658), .Z(n1656) );
XOR U2762 ( .A(c552), .B(b[552]), .Z(n1657) );
XNOR U2763 ( .A(b[552]), .B(n1658), .Z(c[552]) );
XNOR U2764 ( .A(a[552]), .B(c552), .Z(n1658) );
XOR U2765 ( .A(c553), .B(n1659), .Z(c554) );
ANDN U2766 ( .B(n1660), .A(n1661), .Z(n1659) );
XOR U2767 ( .A(c553), .B(b[553]), .Z(n1660) );
XNOR U2768 ( .A(b[553]), .B(n1661), .Z(c[553]) );
XNOR U2769 ( .A(a[553]), .B(c553), .Z(n1661) );
XOR U2770 ( .A(c554), .B(n1662), .Z(c555) );
ANDN U2771 ( .B(n1663), .A(n1664), .Z(n1662) );
XOR U2772 ( .A(c554), .B(b[554]), .Z(n1663) );
XNOR U2773 ( .A(b[554]), .B(n1664), .Z(c[554]) );
XNOR U2774 ( .A(a[554]), .B(c554), .Z(n1664) );
XOR U2775 ( .A(c555), .B(n1665), .Z(c556) );
ANDN U2776 ( .B(n1666), .A(n1667), .Z(n1665) );
XOR U2777 ( .A(c555), .B(b[555]), .Z(n1666) );
XNOR U2778 ( .A(b[555]), .B(n1667), .Z(c[555]) );
XNOR U2779 ( .A(a[555]), .B(c555), .Z(n1667) );
XOR U2780 ( .A(c556), .B(n1668), .Z(c557) );
ANDN U2781 ( .B(n1669), .A(n1670), .Z(n1668) );
XOR U2782 ( .A(c556), .B(b[556]), .Z(n1669) );
XNOR U2783 ( .A(b[556]), .B(n1670), .Z(c[556]) );
XNOR U2784 ( .A(a[556]), .B(c556), .Z(n1670) );
XOR U2785 ( .A(c557), .B(n1671), .Z(c558) );
ANDN U2786 ( .B(n1672), .A(n1673), .Z(n1671) );
XOR U2787 ( .A(c557), .B(b[557]), .Z(n1672) );
XNOR U2788 ( .A(b[557]), .B(n1673), .Z(c[557]) );
XNOR U2789 ( .A(a[557]), .B(c557), .Z(n1673) );
XOR U2790 ( .A(c558), .B(n1674), .Z(c559) );
ANDN U2791 ( .B(n1675), .A(n1676), .Z(n1674) );
XOR U2792 ( .A(c558), .B(b[558]), .Z(n1675) );
XNOR U2793 ( .A(b[558]), .B(n1676), .Z(c[558]) );
XNOR U2794 ( .A(a[558]), .B(c558), .Z(n1676) );
XOR U2795 ( .A(c559), .B(n1677), .Z(c560) );
ANDN U2796 ( .B(n1678), .A(n1679), .Z(n1677) );
XOR U2797 ( .A(c559), .B(b[559]), .Z(n1678) );
XNOR U2798 ( .A(b[559]), .B(n1679), .Z(c[559]) );
XNOR U2799 ( .A(a[559]), .B(c559), .Z(n1679) );
XOR U2800 ( .A(c560), .B(n1680), .Z(c561) );
ANDN U2801 ( .B(n1681), .A(n1682), .Z(n1680) );
XOR U2802 ( .A(c560), .B(b[560]), .Z(n1681) );
XNOR U2803 ( .A(b[560]), .B(n1682), .Z(c[560]) );
XNOR U2804 ( .A(a[560]), .B(c560), .Z(n1682) );
XOR U2805 ( .A(c561), .B(n1683), .Z(c562) );
ANDN U2806 ( .B(n1684), .A(n1685), .Z(n1683) );
XOR U2807 ( .A(c561), .B(b[561]), .Z(n1684) );
XNOR U2808 ( .A(b[561]), .B(n1685), .Z(c[561]) );
XNOR U2809 ( .A(a[561]), .B(c561), .Z(n1685) );
XOR U2810 ( .A(c562), .B(n1686), .Z(c563) );
ANDN U2811 ( .B(n1687), .A(n1688), .Z(n1686) );
XOR U2812 ( .A(c562), .B(b[562]), .Z(n1687) );
XNOR U2813 ( .A(b[562]), .B(n1688), .Z(c[562]) );
XNOR U2814 ( .A(a[562]), .B(c562), .Z(n1688) );
XOR U2815 ( .A(c563), .B(n1689), .Z(c564) );
ANDN U2816 ( .B(n1690), .A(n1691), .Z(n1689) );
XOR U2817 ( .A(c563), .B(b[563]), .Z(n1690) );
XNOR U2818 ( .A(b[563]), .B(n1691), .Z(c[563]) );
XNOR U2819 ( .A(a[563]), .B(c563), .Z(n1691) );
XOR U2820 ( .A(c564), .B(n1692), .Z(c565) );
ANDN U2821 ( .B(n1693), .A(n1694), .Z(n1692) );
XOR U2822 ( .A(c564), .B(b[564]), .Z(n1693) );
XNOR U2823 ( .A(b[564]), .B(n1694), .Z(c[564]) );
XNOR U2824 ( .A(a[564]), .B(c564), .Z(n1694) );
XOR U2825 ( .A(c565), .B(n1695), .Z(c566) );
ANDN U2826 ( .B(n1696), .A(n1697), .Z(n1695) );
XOR U2827 ( .A(c565), .B(b[565]), .Z(n1696) );
XNOR U2828 ( .A(b[565]), .B(n1697), .Z(c[565]) );
XNOR U2829 ( .A(a[565]), .B(c565), .Z(n1697) );
XOR U2830 ( .A(c566), .B(n1698), .Z(c567) );
ANDN U2831 ( .B(n1699), .A(n1700), .Z(n1698) );
XOR U2832 ( .A(c566), .B(b[566]), .Z(n1699) );
XNOR U2833 ( .A(b[566]), .B(n1700), .Z(c[566]) );
XNOR U2834 ( .A(a[566]), .B(c566), .Z(n1700) );
XOR U2835 ( .A(c567), .B(n1701), .Z(c568) );
ANDN U2836 ( .B(n1702), .A(n1703), .Z(n1701) );
XOR U2837 ( .A(c567), .B(b[567]), .Z(n1702) );
XNOR U2838 ( .A(b[567]), .B(n1703), .Z(c[567]) );
XNOR U2839 ( .A(a[567]), .B(c567), .Z(n1703) );
XOR U2840 ( .A(c568), .B(n1704), .Z(c569) );
ANDN U2841 ( .B(n1705), .A(n1706), .Z(n1704) );
XOR U2842 ( .A(c568), .B(b[568]), .Z(n1705) );
XNOR U2843 ( .A(b[568]), .B(n1706), .Z(c[568]) );
XNOR U2844 ( .A(a[568]), .B(c568), .Z(n1706) );
XOR U2845 ( .A(c569), .B(n1707), .Z(c570) );
ANDN U2846 ( .B(n1708), .A(n1709), .Z(n1707) );
XOR U2847 ( .A(c569), .B(b[569]), .Z(n1708) );
XNOR U2848 ( .A(b[569]), .B(n1709), .Z(c[569]) );
XNOR U2849 ( .A(a[569]), .B(c569), .Z(n1709) );
XOR U2850 ( .A(c570), .B(n1710), .Z(c571) );
ANDN U2851 ( .B(n1711), .A(n1712), .Z(n1710) );
XOR U2852 ( .A(c570), .B(b[570]), .Z(n1711) );
XNOR U2853 ( .A(b[570]), .B(n1712), .Z(c[570]) );
XNOR U2854 ( .A(a[570]), .B(c570), .Z(n1712) );
XOR U2855 ( .A(c571), .B(n1713), .Z(c572) );
ANDN U2856 ( .B(n1714), .A(n1715), .Z(n1713) );
XOR U2857 ( .A(c571), .B(b[571]), .Z(n1714) );
XNOR U2858 ( .A(b[571]), .B(n1715), .Z(c[571]) );
XNOR U2859 ( .A(a[571]), .B(c571), .Z(n1715) );
XOR U2860 ( .A(c572), .B(n1716), .Z(c573) );
ANDN U2861 ( .B(n1717), .A(n1718), .Z(n1716) );
XOR U2862 ( .A(c572), .B(b[572]), .Z(n1717) );
XNOR U2863 ( .A(b[572]), .B(n1718), .Z(c[572]) );
XNOR U2864 ( .A(a[572]), .B(c572), .Z(n1718) );
XOR U2865 ( .A(c573), .B(n1719), .Z(c574) );
ANDN U2866 ( .B(n1720), .A(n1721), .Z(n1719) );
XOR U2867 ( .A(c573), .B(b[573]), .Z(n1720) );
XNOR U2868 ( .A(b[573]), .B(n1721), .Z(c[573]) );
XNOR U2869 ( .A(a[573]), .B(c573), .Z(n1721) );
XOR U2870 ( .A(c574), .B(n1722), .Z(c575) );
ANDN U2871 ( .B(n1723), .A(n1724), .Z(n1722) );
XOR U2872 ( .A(c574), .B(b[574]), .Z(n1723) );
XNOR U2873 ( .A(b[574]), .B(n1724), .Z(c[574]) );
XNOR U2874 ( .A(a[574]), .B(c574), .Z(n1724) );
XOR U2875 ( .A(c575), .B(n1725), .Z(c576) );
ANDN U2876 ( .B(n1726), .A(n1727), .Z(n1725) );
XOR U2877 ( .A(c575), .B(b[575]), .Z(n1726) );
XNOR U2878 ( .A(b[575]), .B(n1727), .Z(c[575]) );
XNOR U2879 ( .A(a[575]), .B(c575), .Z(n1727) );
XOR U2880 ( .A(c576), .B(n1728), .Z(c577) );
ANDN U2881 ( .B(n1729), .A(n1730), .Z(n1728) );
XOR U2882 ( .A(c576), .B(b[576]), .Z(n1729) );
XNOR U2883 ( .A(b[576]), .B(n1730), .Z(c[576]) );
XNOR U2884 ( .A(a[576]), .B(c576), .Z(n1730) );
XOR U2885 ( .A(c577), .B(n1731), .Z(c578) );
ANDN U2886 ( .B(n1732), .A(n1733), .Z(n1731) );
XOR U2887 ( .A(c577), .B(b[577]), .Z(n1732) );
XNOR U2888 ( .A(b[577]), .B(n1733), .Z(c[577]) );
XNOR U2889 ( .A(a[577]), .B(c577), .Z(n1733) );
XOR U2890 ( .A(c578), .B(n1734), .Z(c579) );
ANDN U2891 ( .B(n1735), .A(n1736), .Z(n1734) );
XOR U2892 ( .A(c578), .B(b[578]), .Z(n1735) );
XNOR U2893 ( .A(b[578]), .B(n1736), .Z(c[578]) );
XNOR U2894 ( .A(a[578]), .B(c578), .Z(n1736) );
XOR U2895 ( .A(c579), .B(n1737), .Z(c580) );
ANDN U2896 ( .B(n1738), .A(n1739), .Z(n1737) );
XOR U2897 ( .A(c579), .B(b[579]), .Z(n1738) );
XNOR U2898 ( .A(b[579]), .B(n1739), .Z(c[579]) );
XNOR U2899 ( .A(a[579]), .B(c579), .Z(n1739) );
XOR U2900 ( .A(c580), .B(n1740), .Z(c581) );
ANDN U2901 ( .B(n1741), .A(n1742), .Z(n1740) );
XOR U2902 ( .A(c580), .B(b[580]), .Z(n1741) );
XNOR U2903 ( .A(b[580]), .B(n1742), .Z(c[580]) );
XNOR U2904 ( .A(a[580]), .B(c580), .Z(n1742) );
XOR U2905 ( .A(c581), .B(n1743), .Z(c582) );
ANDN U2906 ( .B(n1744), .A(n1745), .Z(n1743) );
XOR U2907 ( .A(c581), .B(b[581]), .Z(n1744) );
XNOR U2908 ( .A(b[581]), .B(n1745), .Z(c[581]) );
XNOR U2909 ( .A(a[581]), .B(c581), .Z(n1745) );
XOR U2910 ( .A(c582), .B(n1746), .Z(c583) );
ANDN U2911 ( .B(n1747), .A(n1748), .Z(n1746) );
XOR U2912 ( .A(c582), .B(b[582]), .Z(n1747) );
XNOR U2913 ( .A(b[582]), .B(n1748), .Z(c[582]) );
XNOR U2914 ( .A(a[582]), .B(c582), .Z(n1748) );
XOR U2915 ( .A(c583), .B(n1749), .Z(c584) );
ANDN U2916 ( .B(n1750), .A(n1751), .Z(n1749) );
XOR U2917 ( .A(c583), .B(b[583]), .Z(n1750) );
XNOR U2918 ( .A(b[583]), .B(n1751), .Z(c[583]) );
XNOR U2919 ( .A(a[583]), .B(c583), .Z(n1751) );
XOR U2920 ( .A(c584), .B(n1752), .Z(c585) );
ANDN U2921 ( .B(n1753), .A(n1754), .Z(n1752) );
XOR U2922 ( .A(c584), .B(b[584]), .Z(n1753) );
XNOR U2923 ( .A(b[584]), .B(n1754), .Z(c[584]) );
XNOR U2924 ( .A(a[584]), .B(c584), .Z(n1754) );
XOR U2925 ( .A(c585), .B(n1755), .Z(c586) );
ANDN U2926 ( .B(n1756), .A(n1757), .Z(n1755) );
XOR U2927 ( .A(c585), .B(b[585]), .Z(n1756) );
XNOR U2928 ( .A(b[585]), .B(n1757), .Z(c[585]) );
XNOR U2929 ( .A(a[585]), .B(c585), .Z(n1757) );
XOR U2930 ( .A(c586), .B(n1758), .Z(c587) );
ANDN U2931 ( .B(n1759), .A(n1760), .Z(n1758) );
XOR U2932 ( .A(c586), .B(b[586]), .Z(n1759) );
XNOR U2933 ( .A(b[586]), .B(n1760), .Z(c[586]) );
XNOR U2934 ( .A(a[586]), .B(c586), .Z(n1760) );
XOR U2935 ( .A(c587), .B(n1761), .Z(c588) );
ANDN U2936 ( .B(n1762), .A(n1763), .Z(n1761) );
XOR U2937 ( .A(c587), .B(b[587]), .Z(n1762) );
XNOR U2938 ( .A(b[587]), .B(n1763), .Z(c[587]) );
XNOR U2939 ( .A(a[587]), .B(c587), .Z(n1763) );
XOR U2940 ( .A(c588), .B(n1764), .Z(c589) );
ANDN U2941 ( .B(n1765), .A(n1766), .Z(n1764) );
XOR U2942 ( .A(c588), .B(b[588]), .Z(n1765) );
XNOR U2943 ( .A(b[588]), .B(n1766), .Z(c[588]) );
XNOR U2944 ( .A(a[588]), .B(c588), .Z(n1766) );
XOR U2945 ( .A(c589), .B(n1767), .Z(c590) );
ANDN U2946 ( .B(n1768), .A(n1769), .Z(n1767) );
XOR U2947 ( .A(c589), .B(b[589]), .Z(n1768) );
XNOR U2948 ( .A(b[589]), .B(n1769), .Z(c[589]) );
XNOR U2949 ( .A(a[589]), .B(c589), .Z(n1769) );
XOR U2950 ( .A(c590), .B(n1770), .Z(c591) );
ANDN U2951 ( .B(n1771), .A(n1772), .Z(n1770) );
XOR U2952 ( .A(c590), .B(b[590]), .Z(n1771) );
XNOR U2953 ( .A(b[590]), .B(n1772), .Z(c[590]) );
XNOR U2954 ( .A(a[590]), .B(c590), .Z(n1772) );
XOR U2955 ( .A(c591), .B(n1773), .Z(c592) );
ANDN U2956 ( .B(n1774), .A(n1775), .Z(n1773) );
XOR U2957 ( .A(c591), .B(b[591]), .Z(n1774) );
XNOR U2958 ( .A(b[591]), .B(n1775), .Z(c[591]) );
XNOR U2959 ( .A(a[591]), .B(c591), .Z(n1775) );
XOR U2960 ( .A(c592), .B(n1776), .Z(c593) );
ANDN U2961 ( .B(n1777), .A(n1778), .Z(n1776) );
XOR U2962 ( .A(c592), .B(b[592]), .Z(n1777) );
XNOR U2963 ( .A(b[592]), .B(n1778), .Z(c[592]) );
XNOR U2964 ( .A(a[592]), .B(c592), .Z(n1778) );
XOR U2965 ( .A(c593), .B(n1779), .Z(c594) );
ANDN U2966 ( .B(n1780), .A(n1781), .Z(n1779) );
XOR U2967 ( .A(c593), .B(b[593]), .Z(n1780) );
XNOR U2968 ( .A(b[593]), .B(n1781), .Z(c[593]) );
XNOR U2969 ( .A(a[593]), .B(c593), .Z(n1781) );
XOR U2970 ( .A(c594), .B(n1782), .Z(c595) );
ANDN U2971 ( .B(n1783), .A(n1784), .Z(n1782) );
XOR U2972 ( .A(c594), .B(b[594]), .Z(n1783) );
XNOR U2973 ( .A(b[594]), .B(n1784), .Z(c[594]) );
XNOR U2974 ( .A(a[594]), .B(c594), .Z(n1784) );
XOR U2975 ( .A(c595), .B(n1785), .Z(c596) );
ANDN U2976 ( .B(n1786), .A(n1787), .Z(n1785) );
XOR U2977 ( .A(c595), .B(b[595]), .Z(n1786) );
XNOR U2978 ( .A(b[595]), .B(n1787), .Z(c[595]) );
XNOR U2979 ( .A(a[595]), .B(c595), .Z(n1787) );
XOR U2980 ( .A(c596), .B(n1788), .Z(c597) );
ANDN U2981 ( .B(n1789), .A(n1790), .Z(n1788) );
XOR U2982 ( .A(c596), .B(b[596]), .Z(n1789) );
XNOR U2983 ( .A(b[596]), .B(n1790), .Z(c[596]) );
XNOR U2984 ( .A(a[596]), .B(c596), .Z(n1790) );
XOR U2985 ( .A(c597), .B(n1791), .Z(c598) );
ANDN U2986 ( .B(n1792), .A(n1793), .Z(n1791) );
XOR U2987 ( .A(c597), .B(b[597]), .Z(n1792) );
XNOR U2988 ( .A(b[597]), .B(n1793), .Z(c[597]) );
XNOR U2989 ( .A(a[597]), .B(c597), .Z(n1793) );
XOR U2990 ( .A(c598), .B(n1794), .Z(c599) );
ANDN U2991 ( .B(n1795), .A(n1796), .Z(n1794) );
XOR U2992 ( .A(c598), .B(b[598]), .Z(n1795) );
XNOR U2993 ( .A(b[598]), .B(n1796), .Z(c[598]) );
XNOR U2994 ( .A(a[598]), .B(c598), .Z(n1796) );
XOR U2995 ( .A(c599), .B(n1797), .Z(c600) );
ANDN U2996 ( .B(n1798), .A(n1799), .Z(n1797) );
XOR U2997 ( .A(c599), .B(b[599]), .Z(n1798) );
XNOR U2998 ( .A(b[599]), .B(n1799), .Z(c[599]) );
XNOR U2999 ( .A(a[599]), .B(c599), .Z(n1799) );
XOR U3000 ( .A(c600), .B(n1800), .Z(c601) );
ANDN U3001 ( .B(n1801), .A(n1802), .Z(n1800) );
XOR U3002 ( .A(c600), .B(b[600]), .Z(n1801) );
XNOR U3003 ( .A(b[600]), .B(n1802), .Z(c[600]) );
XNOR U3004 ( .A(a[600]), .B(c600), .Z(n1802) );
XOR U3005 ( .A(c601), .B(n1803), .Z(c602) );
ANDN U3006 ( .B(n1804), .A(n1805), .Z(n1803) );
XOR U3007 ( .A(c601), .B(b[601]), .Z(n1804) );
XNOR U3008 ( .A(b[601]), .B(n1805), .Z(c[601]) );
XNOR U3009 ( .A(a[601]), .B(c601), .Z(n1805) );
XOR U3010 ( .A(c602), .B(n1806), .Z(c603) );
ANDN U3011 ( .B(n1807), .A(n1808), .Z(n1806) );
XOR U3012 ( .A(c602), .B(b[602]), .Z(n1807) );
XNOR U3013 ( .A(b[602]), .B(n1808), .Z(c[602]) );
XNOR U3014 ( .A(a[602]), .B(c602), .Z(n1808) );
XOR U3015 ( .A(c603), .B(n1809), .Z(c604) );
ANDN U3016 ( .B(n1810), .A(n1811), .Z(n1809) );
XOR U3017 ( .A(c603), .B(b[603]), .Z(n1810) );
XNOR U3018 ( .A(b[603]), .B(n1811), .Z(c[603]) );
XNOR U3019 ( .A(a[603]), .B(c603), .Z(n1811) );
XOR U3020 ( .A(c604), .B(n1812), .Z(c605) );
ANDN U3021 ( .B(n1813), .A(n1814), .Z(n1812) );
XOR U3022 ( .A(c604), .B(b[604]), .Z(n1813) );
XNOR U3023 ( .A(b[604]), .B(n1814), .Z(c[604]) );
XNOR U3024 ( .A(a[604]), .B(c604), .Z(n1814) );
XOR U3025 ( .A(c605), .B(n1815), .Z(c606) );
ANDN U3026 ( .B(n1816), .A(n1817), .Z(n1815) );
XOR U3027 ( .A(c605), .B(b[605]), .Z(n1816) );
XNOR U3028 ( .A(b[605]), .B(n1817), .Z(c[605]) );
XNOR U3029 ( .A(a[605]), .B(c605), .Z(n1817) );
XOR U3030 ( .A(c606), .B(n1818), .Z(c607) );
ANDN U3031 ( .B(n1819), .A(n1820), .Z(n1818) );
XOR U3032 ( .A(c606), .B(b[606]), .Z(n1819) );
XNOR U3033 ( .A(b[606]), .B(n1820), .Z(c[606]) );
XNOR U3034 ( .A(a[606]), .B(c606), .Z(n1820) );
XOR U3035 ( .A(c607), .B(n1821), .Z(c608) );
ANDN U3036 ( .B(n1822), .A(n1823), .Z(n1821) );
XOR U3037 ( .A(c607), .B(b[607]), .Z(n1822) );
XNOR U3038 ( .A(b[607]), .B(n1823), .Z(c[607]) );
XNOR U3039 ( .A(a[607]), .B(c607), .Z(n1823) );
XOR U3040 ( .A(c608), .B(n1824), .Z(c609) );
ANDN U3041 ( .B(n1825), .A(n1826), .Z(n1824) );
XOR U3042 ( .A(c608), .B(b[608]), .Z(n1825) );
XNOR U3043 ( .A(b[608]), .B(n1826), .Z(c[608]) );
XNOR U3044 ( .A(a[608]), .B(c608), .Z(n1826) );
XOR U3045 ( .A(c609), .B(n1827), .Z(c610) );
ANDN U3046 ( .B(n1828), .A(n1829), .Z(n1827) );
XOR U3047 ( .A(c609), .B(b[609]), .Z(n1828) );
XNOR U3048 ( .A(b[609]), .B(n1829), .Z(c[609]) );
XNOR U3049 ( .A(a[609]), .B(c609), .Z(n1829) );
XOR U3050 ( .A(c610), .B(n1830), .Z(c611) );
ANDN U3051 ( .B(n1831), .A(n1832), .Z(n1830) );
XOR U3052 ( .A(c610), .B(b[610]), .Z(n1831) );
XNOR U3053 ( .A(b[610]), .B(n1832), .Z(c[610]) );
XNOR U3054 ( .A(a[610]), .B(c610), .Z(n1832) );
XOR U3055 ( .A(c611), .B(n1833), .Z(c612) );
ANDN U3056 ( .B(n1834), .A(n1835), .Z(n1833) );
XOR U3057 ( .A(c611), .B(b[611]), .Z(n1834) );
XNOR U3058 ( .A(b[611]), .B(n1835), .Z(c[611]) );
XNOR U3059 ( .A(a[611]), .B(c611), .Z(n1835) );
XOR U3060 ( .A(c612), .B(n1836), .Z(c613) );
ANDN U3061 ( .B(n1837), .A(n1838), .Z(n1836) );
XOR U3062 ( .A(c612), .B(b[612]), .Z(n1837) );
XNOR U3063 ( .A(b[612]), .B(n1838), .Z(c[612]) );
XNOR U3064 ( .A(a[612]), .B(c612), .Z(n1838) );
XOR U3065 ( .A(c613), .B(n1839), .Z(c614) );
ANDN U3066 ( .B(n1840), .A(n1841), .Z(n1839) );
XOR U3067 ( .A(c613), .B(b[613]), .Z(n1840) );
XNOR U3068 ( .A(b[613]), .B(n1841), .Z(c[613]) );
XNOR U3069 ( .A(a[613]), .B(c613), .Z(n1841) );
XOR U3070 ( .A(c614), .B(n1842), .Z(c615) );
ANDN U3071 ( .B(n1843), .A(n1844), .Z(n1842) );
XOR U3072 ( .A(c614), .B(b[614]), .Z(n1843) );
XNOR U3073 ( .A(b[614]), .B(n1844), .Z(c[614]) );
XNOR U3074 ( .A(a[614]), .B(c614), .Z(n1844) );
XOR U3075 ( .A(c615), .B(n1845), .Z(c616) );
ANDN U3076 ( .B(n1846), .A(n1847), .Z(n1845) );
XOR U3077 ( .A(c615), .B(b[615]), .Z(n1846) );
XNOR U3078 ( .A(b[615]), .B(n1847), .Z(c[615]) );
XNOR U3079 ( .A(a[615]), .B(c615), .Z(n1847) );
XOR U3080 ( .A(c616), .B(n1848), .Z(c617) );
ANDN U3081 ( .B(n1849), .A(n1850), .Z(n1848) );
XOR U3082 ( .A(c616), .B(b[616]), .Z(n1849) );
XNOR U3083 ( .A(b[616]), .B(n1850), .Z(c[616]) );
XNOR U3084 ( .A(a[616]), .B(c616), .Z(n1850) );
XOR U3085 ( .A(c617), .B(n1851), .Z(c618) );
ANDN U3086 ( .B(n1852), .A(n1853), .Z(n1851) );
XOR U3087 ( .A(c617), .B(b[617]), .Z(n1852) );
XNOR U3088 ( .A(b[617]), .B(n1853), .Z(c[617]) );
XNOR U3089 ( .A(a[617]), .B(c617), .Z(n1853) );
XOR U3090 ( .A(c618), .B(n1854), .Z(c619) );
ANDN U3091 ( .B(n1855), .A(n1856), .Z(n1854) );
XOR U3092 ( .A(c618), .B(b[618]), .Z(n1855) );
XNOR U3093 ( .A(b[618]), .B(n1856), .Z(c[618]) );
XNOR U3094 ( .A(a[618]), .B(c618), .Z(n1856) );
XOR U3095 ( .A(c619), .B(n1857), .Z(c620) );
ANDN U3096 ( .B(n1858), .A(n1859), .Z(n1857) );
XOR U3097 ( .A(c619), .B(b[619]), .Z(n1858) );
XNOR U3098 ( .A(b[619]), .B(n1859), .Z(c[619]) );
XNOR U3099 ( .A(a[619]), .B(c619), .Z(n1859) );
XOR U3100 ( .A(c620), .B(n1860), .Z(c621) );
ANDN U3101 ( .B(n1861), .A(n1862), .Z(n1860) );
XOR U3102 ( .A(c620), .B(b[620]), .Z(n1861) );
XNOR U3103 ( .A(b[620]), .B(n1862), .Z(c[620]) );
XNOR U3104 ( .A(a[620]), .B(c620), .Z(n1862) );
XOR U3105 ( .A(c621), .B(n1863), .Z(c622) );
ANDN U3106 ( .B(n1864), .A(n1865), .Z(n1863) );
XOR U3107 ( .A(c621), .B(b[621]), .Z(n1864) );
XNOR U3108 ( .A(b[621]), .B(n1865), .Z(c[621]) );
XNOR U3109 ( .A(a[621]), .B(c621), .Z(n1865) );
XOR U3110 ( .A(c622), .B(n1866), .Z(c623) );
ANDN U3111 ( .B(n1867), .A(n1868), .Z(n1866) );
XOR U3112 ( .A(c622), .B(b[622]), .Z(n1867) );
XNOR U3113 ( .A(b[622]), .B(n1868), .Z(c[622]) );
XNOR U3114 ( .A(a[622]), .B(c622), .Z(n1868) );
XOR U3115 ( .A(c623), .B(n1869), .Z(c624) );
ANDN U3116 ( .B(n1870), .A(n1871), .Z(n1869) );
XOR U3117 ( .A(c623), .B(b[623]), .Z(n1870) );
XNOR U3118 ( .A(b[623]), .B(n1871), .Z(c[623]) );
XNOR U3119 ( .A(a[623]), .B(c623), .Z(n1871) );
XOR U3120 ( .A(c624), .B(n1872), .Z(c625) );
ANDN U3121 ( .B(n1873), .A(n1874), .Z(n1872) );
XOR U3122 ( .A(c624), .B(b[624]), .Z(n1873) );
XNOR U3123 ( .A(b[624]), .B(n1874), .Z(c[624]) );
XNOR U3124 ( .A(a[624]), .B(c624), .Z(n1874) );
XOR U3125 ( .A(c625), .B(n1875), .Z(c626) );
ANDN U3126 ( .B(n1876), .A(n1877), .Z(n1875) );
XOR U3127 ( .A(c625), .B(b[625]), .Z(n1876) );
XNOR U3128 ( .A(b[625]), .B(n1877), .Z(c[625]) );
XNOR U3129 ( .A(a[625]), .B(c625), .Z(n1877) );
XOR U3130 ( .A(c626), .B(n1878), .Z(c627) );
ANDN U3131 ( .B(n1879), .A(n1880), .Z(n1878) );
XOR U3132 ( .A(c626), .B(b[626]), .Z(n1879) );
XNOR U3133 ( .A(b[626]), .B(n1880), .Z(c[626]) );
XNOR U3134 ( .A(a[626]), .B(c626), .Z(n1880) );
XOR U3135 ( .A(c627), .B(n1881), .Z(c628) );
ANDN U3136 ( .B(n1882), .A(n1883), .Z(n1881) );
XOR U3137 ( .A(c627), .B(b[627]), .Z(n1882) );
XNOR U3138 ( .A(b[627]), .B(n1883), .Z(c[627]) );
XNOR U3139 ( .A(a[627]), .B(c627), .Z(n1883) );
XOR U3140 ( .A(c628), .B(n1884), .Z(c629) );
ANDN U3141 ( .B(n1885), .A(n1886), .Z(n1884) );
XOR U3142 ( .A(c628), .B(b[628]), .Z(n1885) );
XNOR U3143 ( .A(b[628]), .B(n1886), .Z(c[628]) );
XNOR U3144 ( .A(a[628]), .B(c628), .Z(n1886) );
XOR U3145 ( .A(c629), .B(n1887), .Z(c630) );
ANDN U3146 ( .B(n1888), .A(n1889), .Z(n1887) );
XOR U3147 ( .A(c629), .B(b[629]), .Z(n1888) );
XNOR U3148 ( .A(b[629]), .B(n1889), .Z(c[629]) );
XNOR U3149 ( .A(a[629]), .B(c629), .Z(n1889) );
XOR U3150 ( .A(c630), .B(n1890), .Z(c631) );
ANDN U3151 ( .B(n1891), .A(n1892), .Z(n1890) );
XOR U3152 ( .A(c630), .B(b[630]), .Z(n1891) );
XNOR U3153 ( .A(b[630]), .B(n1892), .Z(c[630]) );
XNOR U3154 ( .A(a[630]), .B(c630), .Z(n1892) );
XOR U3155 ( .A(c631), .B(n1893), .Z(c632) );
ANDN U3156 ( .B(n1894), .A(n1895), .Z(n1893) );
XOR U3157 ( .A(c631), .B(b[631]), .Z(n1894) );
XNOR U3158 ( .A(b[631]), .B(n1895), .Z(c[631]) );
XNOR U3159 ( .A(a[631]), .B(c631), .Z(n1895) );
XOR U3160 ( .A(c632), .B(n1896), .Z(c633) );
ANDN U3161 ( .B(n1897), .A(n1898), .Z(n1896) );
XOR U3162 ( .A(c632), .B(b[632]), .Z(n1897) );
XNOR U3163 ( .A(b[632]), .B(n1898), .Z(c[632]) );
XNOR U3164 ( .A(a[632]), .B(c632), .Z(n1898) );
XOR U3165 ( .A(c633), .B(n1899), .Z(c634) );
ANDN U3166 ( .B(n1900), .A(n1901), .Z(n1899) );
XOR U3167 ( .A(c633), .B(b[633]), .Z(n1900) );
XNOR U3168 ( .A(b[633]), .B(n1901), .Z(c[633]) );
XNOR U3169 ( .A(a[633]), .B(c633), .Z(n1901) );
XOR U3170 ( .A(c634), .B(n1902), .Z(c635) );
ANDN U3171 ( .B(n1903), .A(n1904), .Z(n1902) );
XOR U3172 ( .A(c634), .B(b[634]), .Z(n1903) );
XNOR U3173 ( .A(b[634]), .B(n1904), .Z(c[634]) );
XNOR U3174 ( .A(a[634]), .B(c634), .Z(n1904) );
XOR U3175 ( .A(c635), .B(n1905), .Z(c636) );
ANDN U3176 ( .B(n1906), .A(n1907), .Z(n1905) );
XOR U3177 ( .A(c635), .B(b[635]), .Z(n1906) );
XNOR U3178 ( .A(b[635]), .B(n1907), .Z(c[635]) );
XNOR U3179 ( .A(a[635]), .B(c635), .Z(n1907) );
XOR U3180 ( .A(c636), .B(n1908), .Z(c637) );
ANDN U3181 ( .B(n1909), .A(n1910), .Z(n1908) );
XOR U3182 ( .A(c636), .B(b[636]), .Z(n1909) );
XNOR U3183 ( .A(b[636]), .B(n1910), .Z(c[636]) );
XNOR U3184 ( .A(a[636]), .B(c636), .Z(n1910) );
XOR U3185 ( .A(c637), .B(n1911), .Z(c638) );
ANDN U3186 ( .B(n1912), .A(n1913), .Z(n1911) );
XOR U3187 ( .A(c637), .B(b[637]), .Z(n1912) );
XNOR U3188 ( .A(b[637]), .B(n1913), .Z(c[637]) );
XNOR U3189 ( .A(a[637]), .B(c637), .Z(n1913) );
XOR U3190 ( .A(c638), .B(n1914), .Z(c639) );
ANDN U3191 ( .B(n1915), .A(n1916), .Z(n1914) );
XOR U3192 ( .A(c638), .B(b[638]), .Z(n1915) );
XNOR U3193 ( .A(b[638]), .B(n1916), .Z(c[638]) );
XNOR U3194 ( .A(a[638]), .B(c638), .Z(n1916) );
XOR U3195 ( .A(c639), .B(n1917), .Z(c640) );
ANDN U3196 ( .B(n1918), .A(n1919), .Z(n1917) );
XOR U3197 ( .A(c639), .B(b[639]), .Z(n1918) );
XNOR U3198 ( .A(b[639]), .B(n1919), .Z(c[639]) );
XNOR U3199 ( .A(a[639]), .B(c639), .Z(n1919) );
XOR U3200 ( .A(c640), .B(n1920), .Z(c641) );
ANDN U3201 ( .B(n1921), .A(n1922), .Z(n1920) );
XOR U3202 ( .A(c640), .B(b[640]), .Z(n1921) );
XNOR U3203 ( .A(b[640]), .B(n1922), .Z(c[640]) );
XNOR U3204 ( .A(a[640]), .B(c640), .Z(n1922) );
XOR U3205 ( .A(c641), .B(n1923), .Z(c642) );
ANDN U3206 ( .B(n1924), .A(n1925), .Z(n1923) );
XOR U3207 ( .A(c641), .B(b[641]), .Z(n1924) );
XNOR U3208 ( .A(b[641]), .B(n1925), .Z(c[641]) );
XNOR U3209 ( .A(a[641]), .B(c641), .Z(n1925) );
XOR U3210 ( .A(c642), .B(n1926), .Z(c643) );
ANDN U3211 ( .B(n1927), .A(n1928), .Z(n1926) );
XOR U3212 ( .A(c642), .B(b[642]), .Z(n1927) );
XNOR U3213 ( .A(b[642]), .B(n1928), .Z(c[642]) );
XNOR U3214 ( .A(a[642]), .B(c642), .Z(n1928) );
XOR U3215 ( .A(c643), .B(n1929), .Z(c644) );
ANDN U3216 ( .B(n1930), .A(n1931), .Z(n1929) );
XOR U3217 ( .A(c643), .B(b[643]), .Z(n1930) );
XNOR U3218 ( .A(b[643]), .B(n1931), .Z(c[643]) );
XNOR U3219 ( .A(a[643]), .B(c643), .Z(n1931) );
XOR U3220 ( .A(c644), .B(n1932), .Z(c645) );
ANDN U3221 ( .B(n1933), .A(n1934), .Z(n1932) );
XOR U3222 ( .A(c644), .B(b[644]), .Z(n1933) );
XNOR U3223 ( .A(b[644]), .B(n1934), .Z(c[644]) );
XNOR U3224 ( .A(a[644]), .B(c644), .Z(n1934) );
XOR U3225 ( .A(c645), .B(n1935), .Z(c646) );
ANDN U3226 ( .B(n1936), .A(n1937), .Z(n1935) );
XOR U3227 ( .A(c645), .B(b[645]), .Z(n1936) );
XNOR U3228 ( .A(b[645]), .B(n1937), .Z(c[645]) );
XNOR U3229 ( .A(a[645]), .B(c645), .Z(n1937) );
XOR U3230 ( .A(c646), .B(n1938), .Z(c647) );
ANDN U3231 ( .B(n1939), .A(n1940), .Z(n1938) );
XOR U3232 ( .A(c646), .B(b[646]), .Z(n1939) );
XNOR U3233 ( .A(b[646]), .B(n1940), .Z(c[646]) );
XNOR U3234 ( .A(a[646]), .B(c646), .Z(n1940) );
XOR U3235 ( .A(c647), .B(n1941), .Z(c648) );
ANDN U3236 ( .B(n1942), .A(n1943), .Z(n1941) );
XOR U3237 ( .A(c647), .B(b[647]), .Z(n1942) );
XNOR U3238 ( .A(b[647]), .B(n1943), .Z(c[647]) );
XNOR U3239 ( .A(a[647]), .B(c647), .Z(n1943) );
XOR U3240 ( .A(c648), .B(n1944), .Z(c649) );
ANDN U3241 ( .B(n1945), .A(n1946), .Z(n1944) );
XOR U3242 ( .A(c648), .B(b[648]), .Z(n1945) );
XNOR U3243 ( .A(b[648]), .B(n1946), .Z(c[648]) );
XNOR U3244 ( .A(a[648]), .B(c648), .Z(n1946) );
XOR U3245 ( .A(c649), .B(n1947), .Z(c650) );
ANDN U3246 ( .B(n1948), .A(n1949), .Z(n1947) );
XOR U3247 ( .A(c649), .B(b[649]), .Z(n1948) );
XNOR U3248 ( .A(b[649]), .B(n1949), .Z(c[649]) );
XNOR U3249 ( .A(a[649]), .B(c649), .Z(n1949) );
XOR U3250 ( .A(c650), .B(n1950), .Z(c651) );
ANDN U3251 ( .B(n1951), .A(n1952), .Z(n1950) );
XOR U3252 ( .A(c650), .B(b[650]), .Z(n1951) );
XNOR U3253 ( .A(b[650]), .B(n1952), .Z(c[650]) );
XNOR U3254 ( .A(a[650]), .B(c650), .Z(n1952) );
XOR U3255 ( .A(c651), .B(n1953), .Z(c652) );
ANDN U3256 ( .B(n1954), .A(n1955), .Z(n1953) );
XOR U3257 ( .A(c651), .B(b[651]), .Z(n1954) );
XNOR U3258 ( .A(b[651]), .B(n1955), .Z(c[651]) );
XNOR U3259 ( .A(a[651]), .B(c651), .Z(n1955) );
XOR U3260 ( .A(c652), .B(n1956), .Z(c653) );
ANDN U3261 ( .B(n1957), .A(n1958), .Z(n1956) );
XOR U3262 ( .A(c652), .B(b[652]), .Z(n1957) );
XNOR U3263 ( .A(b[652]), .B(n1958), .Z(c[652]) );
XNOR U3264 ( .A(a[652]), .B(c652), .Z(n1958) );
XOR U3265 ( .A(c653), .B(n1959), .Z(c654) );
ANDN U3266 ( .B(n1960), .A(n1961), .Z(n1959) );
XOR U3267 ( .A(c653), .B(b[653]), .Z(n1960) );
XNOR U3268 ( .A(b[653]), .B(n1961), .Z(c[653]) );
XNOR U3269 ( .A(a[653]), .B(c653), .Z(n1961) );
XOR U3270 ( .A(c654), .B(n1962), .Z(c655) );
ANDN U3271 ( .B(n1963), .A(n1964), .Z(n1962) );
XOR U3272 ( .A(c654), .B(b[654]), .Z(n1963) );
XNOR U3273 ( .A(b[654]), .B(n1964), .Z(c[654]) );
XNOR U3274 ( .A(a[654]), .B(c654), .Z(n1964) );
XOR U3275 ( .A(c655), .B(n1965), .Z(c656) );
ANDN U3276 ( .B(n1966), .A(n1967), .Z(n1965) );
XOR U3277 ( .A(c655), .B(b[655]), .Z(n1966) );
XNOR U3278 ( .A(b[655]), .B(n1967), .Z(c[655]) );
XNOR U3279 ( .A(a[655]), .B(c655), .Z(n1967) );
XOR U3280 ( .A(c656), .B(n1968), .Z(c657) );
ANDN U3281 ( .B(n1969), .A(n1970), .Z(n1968) );
XOR U3282 ( .A(c656), .B(b[656]), .Z(n1969) );
XNOR U3283 ( .A(b[656]), .B(n1970), .Z(c[656]) );
XNOR U3284 ( .A(a[656]), .B(c656), .Z(n1970) );
XOR U3285 ( .A(c657), .B(n1971), .Z(c658) );
ANDN U3286 ( .B(n1972), .A(n1973), .Z(n1971) );
XOR U3287 ( .A(c657), .B(b[657]), .Z(n1972) );
XNOR U3288 ( .A(b[657]), .B(n1973), .Z(c[657]) );
XNOR U3289 ( .A(a[657]), .B(c657), .Z(n1973) );
XOR U3290 ( .A(c658), .B(n1974), .Z(c659) );
ANDN U3291 ( .B(n1975), .A(n1976), .Z(n1974) );
XOR U3292 ( .A(c658), .B(b[658]), .Z(n1975) );
XNOR U3293 ( .A(b[658]), .B(n1976), .Z(c[658]) );
XNOR U3294 ( .A(a[658]), .B(c658), .Z(n1976) );
XOR U3295 ( .A(c659), .B(n1977), .Z(c660) );
ANDN U3296 ( .B(n1978), .A(n1979), .Z(n1977) );
XOR U3297 ( .A(c659), .B(b[659]), .Z(n1978) );
XNOR U3298 ( .A(b[659]), .B(n1979), .Z(c[659]) );
XNOR U3299 ( .A(a[659]), .B(c659), .Z(n1979) );
XOR U3300 ( .A(c660), .B(n1980), .Z(c661) );
ANDN U3301 ( .B(n1981), .A(n1982), .Z(n1980) );
XOR U3302 ( .A(c660), .B(b[660]), .Z(n1981) );
XNOR U3303 ( .A(b[660]), .B(n1982), .Z(c[660]) );
XNOR U3304 ( .A(a[660]), .B(c660), .Z(n1982) );
XOR U3305 ( .A(c661), .B(n1983), .Z(c662) );
ANDN U3306 ( .B(n1984), .A(n1985), .Z(n1983) );
XOR U3307 ( .A(c661), .B(b[661]), .Z(n1984) );
XNOR U3308 ( .A(b[661]), .B(n1985), .Z(c[661]) );
XNOR U3309 ( .A(a[661]), .B(c661), .Z(n1985) );
XOR U3310 ( .A(c662), .B(n1986), .Z(c663) );
ANDN U3311 ( .B(n1987), .A(n1988), .Z(n1986) );
XOR U3312 ( .A(c662), .B(b[662]), .Z(n1987) );
XNOR U3313 ( .A(b[662]), .B(n1988), .Z(c[662]) );
XNOR U3314 ( .A(a[662]), .B(c662), .Z(n1988) );
XOR U3315 ( .A(c663), .B(n1989), .Z(c664) );
ANDN U3316 ( .B(n1990), .A(n1991), .Z(n1989) );
XOR U3317 ( .A(c663), .B(b[663]), .Z(n1990) );
XNOR U3318 ( .A(b[663]), .B(n1991), .Z(c[663]) );
XNOR U3319 ( .A(a[663]), .B(c663), .Z(n1991) );
XOR U3320 ( .A(c664), .B(n1992), .Z(c665) );
ANDN U3321 ( .B(n1993), .A(n1994), .Z(n1992) );
XOR U3322 ( .A(c664), .B(b[664]), .Z(n1993) );
XNOR U3323 ( .A(b[664]), .B(n1994), .Z(c[664]) );
XNOR U3324 ( .A(a[664]), .B(c664), .Z(n1994) );
XOR U3325 ( .A(c665), .B(n1995), .Z(c666) );
ANDN U3326 ( .B(n1996), .A(n1997), .Z(n1995) );
XOR U3327 ( .A(c665), .B(b[665]), .Z(n1996) );
XNOR U3328 ( .A(b[665]), .B(n1997), .Z(c[665]) );
XNOR U3329 ( .A(a[665]), .B(c665), .Z(n1997) );
XOR U3330 ( .A(c666), .B(n1998), .Z(c667) );
ANDN U3331 ( .B(n1999), .A(n2000), .Z(n1998) );
XOR U3332 ( .A(c666), .B(b[666]), .Z(n1999) );
XNOR U3333 ( .A(b[666]), .B(n2000), .Z(c[666]) );
XNOR U3334 ( .A(a[666]), .B(c666), .Z(n2000) );
XOR U3335 ( .A(c667), .B(n2001), .Z(c668) );
ANDN U3336 ( .B(n2002), .A(n2003), .Z(n2001) );
XOR U3337 ( .A(c667), .B(b[667]), .Z(n2002) );
XNOR U3338 ( .A(b[667]), .B(n2003), .Z(c[667]) );
XNOR U3339 ( .A(a[667]), .B(c667), .Z(n2003) );
XOR U3340 ( .A(c668), .B(n2004), .Z(c669) );
ANDN U3341 ( .B(n2005), .A(n2006), .Z(n2004) );
XOR U3342 ( .A(c668), .B(b[668]), .Z(n2005) );
XNOR U3343 ( .A(b[668]), .B(n2006), .Z(c[668]) );
XNOR U3344 ( .A(a[668]), .B(c668), .Z(n2006) );
XOR U3345 ( .A(c669), .B(n2007), .Z(c670) );
ANDN U3346 ( .B(n2008), .A(n2009), .Z(n2007) );
XOR U3347 ( .A(c669), .B(b[669]), .Z(n2008) );
XNOR U3348 ( .A(b[669]), .B(n2009), .Z(c[669]) );
XNOR U3349 ( .A(a[669]), .B(c669), .Z(n2009) );
XOR U3350 ( .A(c670), .B(n2010), .Z(c671) );
ANDN U3351 ( .B(n2011), .A(n2012), .Z(n2010) );
XOR U3352 ( .A(c670), .B(b[670]), .Z(n2011) );
XNOR U3353 ( .A(b[670]), .B(n2012), .Z(c[670]) );
XNOR U3354 ( .A(a[670]), .B(c670), .Z(n2012) );
XOR U3355 ( .A(c671), .B(n2013), .Z(c672) );
ANDN U3356 ( .B(n2014), .A(n2015), .Z(n2013) );
XOR U3357 ( .A(c671), .B(b[671]), .Z(n2014) );
XNOR U3358 ( .A(b[671]), .B(n2015), .Z(c[671]) );
XNOR U3359 ( .A(a[671]), .B(c671), .Z(n2015) );
XOR U3360 ( .A(c672), .B(n2016), .Z(c673) );
ANDN U3361 ( .B(n2017), .A(n2018), .Z(n2016) );
XOR U3362 ( .A(c672), .B(b[672]), .Z(n2017) );
XNOR U3363 ( .A(b[672]), .B(n2018), .Z(c[672]) );
XNOR U3364 ( .A(a[672]), .B(c672), .Z(n2018) );
XOR U3365 ( .A(c673), .B(n2019), .Z(c674) );
ANDN U3366 ( .B(n2020), .A(n2021), .Z(n2019) );
XOR U3367 ( .A(c673), .B(b[673]), .Z(n2020) );
XNOR U3368 ( .A(b[673]), .B(n2021), .Z(c[673]) );
XNOR U3369 ( .A(a[673]), .B(c673), .Z(n2021) );
XOR U3370 ( .A(c674), .B(n2022), .Z(c675) );
ANDN U3371 ( .B(n2023), .A(n2024), .Z(n2022) );
XOR U3372 ( .A(c674), .B(b[674]), .Z(n2023) );
XNOR U3373 ( .A(b[674]), .B(n2024), .Z(c[674]) );
XNOR U3374 ( .A(a[674]), .B(c674), .Z(n2024) );
XOR U3375 ( .A(c675), .B(n2025), .Z(c676) );
ANDN U3376 ( .B(n2026), .A(n2027), .Z(n2025) );
XOR U3377 ( .A(c675), .B(b[675]), .Z(n2026) );
XNOR U3378 ( .A(b[675]), .B(n2027), .Z(c[675]) );
XNOR U3379 ( .A(a[675]), .B(c675), .Z(n2027) );
XOR U3380 ( .A(c676), .B(n2028), .Z(c677) );
ANDN U3381 ( .B(n2029), .A(n2030), .Z(n2028) );
XOR U3382 ( .A(c676), .B(b[676]), .Z(n2029) );
XNOR U3383 ( .A(b[676]), .B(n2030), .Z(c[676]) );
XNOR U3384 ( .A(a[676]), .B(c676), .Z(n2030) );
XOR U3385 ( .A(c677), .B(n2031), .Z(c678) );
ANDN U3386 ( .B(n2032), .A(n2033), .Z(n2031) );
XOR U3387 ( .A(c677), .B(b[677]), .Z(n2032) );
XNOR U3388 ( .A(b[677]), .B(n2033), .Z(c[677]) );
XNOR U3389 ( .A(a[677]), .B(c677), .Z(n2033) );
XOR U3390 ( .A(c678), .B(n2034), .Z(c679) );
ANDN U3391 ( .B(n2035), .A(n2036), .Z(n2034) );
XOR U3392 ( .A(c678), .B(b[678]), .Z(n2035) );
XNOR U3393 ( .A(b[678]), .B(n2036), .Z(c[678]) );
XNOR U3394 ( .A(a[678]), .B(c678), .Z(n2036) );
XOR U3395 ( .A(c679), .B(n2037), .Z(c680) );
ANDN U3396 ( .B(n2038), .A(n2039), .Z(n2037) );
XOR U3397 ( .A(c679), .B(b[679]), .Z(n2038) );
XNOR U3398 ( .A(b[679]), .B(n2039), .Z(c[679]) );
XNOR U3399 ( .A(a[679]), .B(c679), .Z(n2039) );
XOR U3400 ( .A(c680), .B(n2040), .Z(c681) );
ANDN U3401 ( .B(n2041), .A(n2042), .Z(n2040) );
XOR U3402 ( .A(c680), .B(b[680]), .Z(n2041) );
XNOR U3403 ( .A(b[680]), .B(n2042), .Z(c[680]) );
XNOR U3404 ( .A(a[680]), .B(c680), .Z(n2042) );
XOR U3405 ( .A(c681), .B(n2043), .Z(c682) );
ANDN U3406 ( .B(n2044), .A(n2045), .Z(n2043) );
XOR U3407 ( .A(c681), .B(b[681]), .Z(n2044) );
XNOR U3408 ( .A(b[681]), .B(n2045), .Z(c[681]) );
XNOR U3409 ( .A(a[681]), .B(c681), .Z(n2045) );
XOR U3410 ( .A(c682), .B(n2046), .Z(c683) );
ANDN U3411 ( .B(n2047), .A(n2048), .Z(n2046) );
XOR U3412 ( .A(c682), .B(b[682]), .Z(n2047) );
XNOR U3413 ( .A(b[682]), .B(n2048), .Z(c[682]) );
XNOR U3414 ( .A(a[682]), .B(c682), .Z(n2048) );
XOR U3415 ( .A(c683), .B(n2049), .Z(c684) );
ANDN U3416 ( .B(n2050), .A(n2051), .Z(n2049) );
XOR U3417 ( .A(c683), .B(b[683]), .Z(n2050) );
XNOR U3418 ( .A(b[683]), .B(n2051), .Z(c[683]) );
XNOR U3419 ( .A(a[683]), .B(c683), .Z(n2051) );
XOR U3420 ( .A(c684), .B(n2052), .Z(c685) );
ANDN U3421 ( .B(n2053), .A(n2054), .Z(n2052) );
XOR U3422 ( .A(c684), .B(b[684]), .Z(n2053) );
XNOR U3423 ( .A(b[684]), .B(n2054), .Z(c[684]) );
XNOR U3424 ( .A(a[684]), .B(c684), .Z(n2054) );
XOR U3425 ( .A(c685), .B(n2055), .Z(c686) );
ANDN U3426 ( .B(n2056), .A(n2057), .Z(n2055) );
XOR U3427 ( .A(c685), .B(b[685]), .Z(n2056) );
XNOR U3428 ( .A(b[685]), .B(n2057), .Z(c[685]) );
XNOR U3429 ( .A(a[685]), .B(c685), .Z(n2057) );
XOR U3430 ( .A(c686), .B(n2058), .Z(c687) );
ANDN U3431 ( .B(n2059), .A(n2060), .Z(n2058) );
XOR U3432 ( .A(c686), .B(b[686]), .Z(n2059) );
XNOR U3433 ( .A(b[686]), .B(n2060), .Z(c[686]) );
XNOR U3434 ( .A(a[686]), .B(c686), .Z(n2060) );
XOR U3435 ( .A(c687), .B(n2061), .Z(c688) );
ANDN U3436 ( .B(n2062), .A(n2063), .Z(n2061) );
XOR U3437 ( .A(c687), .B(b[687]), .Z(n2062) );
XNOR U3438 ( .A(b[687]), .B(n2063), .Z(c[687]) );
XNOR U3439 ( .A(a[687]), .B(c687), .Z(n2063) );
XOR U3440 ( .A(c688), .B(n2064), .Z(c689) );
ANDN U3441 ( .B(n2065), .A(n2066), .Z(n2064) );
XOR U3442 ( .A(c688), .B(b[688]), .Z(n2065) );
XNOR U3443 ( .A(b[688]), .B(n2066), .Z(c[688]) );
XNOR U3444 ( .A(a[688]), .B(c688), .Z(n2066) );
XOR U3445 ( .A(c689), .B(n2067), .Z(c690) );
ANDN U3446 ( .B(n2068), .A(n2069), .Z(n2067) );
XOR U3447 ( .A(c689), .B(b[689]), .Z(n2068) );
XNOR U3448 ( .A(b[689]), .B(n2069), .Z(c[689]) );
XNOR U3449 ( .A(a[689]), .B(c689), .Z(n2069) );
XOR U3450 ( .A(c690), .B(n2070), .Z(c691) );
ANDN U3451 ( .B(n2071), .A(n2072), .Z(n2070) );
XOR U3452 ( .A(c690), .B(b[690]), .Z(n2071) );
XNOR U3453 ( .A(b[690]), .B(n2072), .Z(c[690]) );
XNOR U3454 ( .A(a[690]), .B(c690), .Z(n2072) );
XOR U3455 ( .A(c691), .B(n2073), .Z(c692) );
ANDN U3456 ( .B(n2074), .A(n2075), .Z(n2073) );
XOR U3457 ( .A(c691), .B(b[691]), .Z(n2074) );
XNOR U3458 ( .A(b[691]), .B(n2075), .Z(c[691]) );
XNOR U3459 ( .A(a[691]), .B(c691), .Z(n2075) );
XOR U3460 ( .A(c692), .B(n2076), .Z(c693) );
ANDN U3461 ( .B(n2077), .A(n2078), .Z(n2076) );
XOR U3462 ( .A(c692), .B(b[692]), .Z(n2077) );
XNOR U3463 ( .A(b[692]), .B(n2078), .Z(c[692]) );
XNOR U3464 ( .A(a[692]), .B(c692), .Z(n2078) );
XOR U3465 ( .A(c693), .B(n2079), .Z(c694) );
ANDN U3466 ( .B(n2080), .A(n2081), .Z(n2079) );
XOR U3467 ( .A(c693), .B(b[693]), .Z(n2080) );
XNOR U3468 ( .A(b[693]), .B(n2081), .Z(c[693]) );
XNOR U3469 ( .A(a[693]), .B(c693), .Z(n2081) );
XOR U3470 ( .A(c694), .B(n2082), .Z(c695) );
ANDN U3471 ( .B(n2083), .A(n2084), .Z(n2082) );
XOR U3472 ( .A(c694), .B(b[694]), .Z(n2083) );
XNOR U3473 ( .A(b[694]), .B(n2084), .Z(c[694]) );
XNOR U3474 ( .A(a[694]), .B(c694), .Z(n2084) );
XOR U3475 ( .A(c695), .B(n2085), .Z(c696) );
ANDN U3476 ( .B(n2086), .A(n2087), .Z(n2085) );
XOR U3477 ( .A(c695), .B(b[695]), .Z(n2086) );
XNOR U3478 ( .A(b[695]), .B(n2087), .Z(c[695]) );
XNOR U3479 ( .A(a[695]), .B(c695), .Z(n2087) );
XOR U3480 ( .A(c696), .B(n2088), .Z(c697) );
ANDN U3481 ( .B(n2089), .A(n2090), .Z(n2088) );
XOR U3482 ( .A(c696), .B(b[696]), .Z(n2089) );
XNOR U3483 ( .A(b[696]), .B(n2090), .Z(c[696]) );
XNOR U3484 ( .A(a[696]), .B(c696), .Z(n2090) );
XOR U3485 ( .A(c697), .B(n2091), .Z(c698) );
ANDN U3486 ( .B(n2092), .A(n2093), .Z(n2091) );
XOR U3487 ( .A(c697), .B(b[697]), .Z(n2092) );
XNOR U3488 ( .A(b[697]), .B(n2093), .Z(c[697]) );
XNOR U3489 ( .A(a[697]), .B(c697), .Z(n2093) );
XOR U3490 ( .A(c698), .B(n2094), .Z(c699) );
ANDN U3491 ( .B(n2095), .A(n2096), .Z(n2094) );
XOR U3492 ( .A(c698), .B(b[698]), .Z(n2095) );
XNOR U3493 ( .A(b[698]), .B(n2096), .Z(c[698]) );
XNOR U3494 ( .A(a[698]), .B(c698), .Z(n2096) );
XOR U3495 ( .A(c699), .B(n2097), .Z(c700) );
ANDN U3496 ( .B(n2098), .A(n2099), .Z(n2097) );
XOR U3497 ( .A(c699), .B(b[699]), .Z(n2098) );
XNOR U3498 ( .A(b[699]), .B(n2099), .Z(c[699]) );
XNOR U3499 ( .A(a[699]), .B(c699), .Z(n2099) );
XOR U3500 ( .A(c700), .B(n2100), .Z(c701) );
ANDN U3501 ( .B(n2101), .A(n2102), .Z(n2100) );
XOR U3502 ( .A(c700), .B(b[700]), .Z(n2101) );
XNOR U3503 ( .A(b[700]), .B(n2102), .Z(c[700]) );
XNOR U3504 ( .A(a[700]), .B(c700), .Z(n2102) );
XOR U3505 ( .A(c701), .B(n2103), .Z(c702) );
ANDN U3506 ( .B(n2104), .A(n2105), .Z(n2103) );
XOR U3507 ( .A(c701), .B(b[701]), .Z(n2104) );
XNOR U3508 ( .A(b[701]), .B(n2105), .Z(c[701]) );
XNOR U3509 ( .A(a[701]), .B(c701), .Z(n2105) );
XOR U3510 ( .A(c702), .B(n2106), .Z(c703) );
ANDN U3511 ( .B(n2107), .A(n2108), .Z(n2106) );
XOR U3512 ( .A(c702), .B(b[702]), .Z(n2107) );
XNOR U3513 ( .A(b[702]), .B(n2108), .Z(c[702]) );
XNOR U3514 ( .A(a[702]), .B(c702), .Z(n2108) );
XOR U3515 ( .A(c703), .B(n2109), .Z(c704) );
ANDN U3516 ( .B(n2110), .A(n2111), .Z(n2109) );
XOR U3517 ( .A(c703), .B(b[703]), .Z(n2110) );
XNOR U3518 ( .A(b[703]), .B(n2111), .Z(c[703]) );
XNOR U3519 ( .A(a[703]), .B(c703), .Z(n2111) );
XOR U3520 ( .A(c704), .B(n2112), .Z(c705) );
ANDN U3521 ( .B(n2113), .A(n2114), .Z(n2112) );
XOR U3522 ( .A(c704), .B(b[704]), .Z(n2113) );
XNOR U3523 ( .A(b[704]), .B(n2114), .Z(c[704]) );
XNOR U3524 ( .A(a[704]), .B(c704), .Z(n2114) );
XOR U3525 ( .A(c705), .B(n2115), .Z(c706) );
ANDN U3526 ( .B(n2116), .A(n2117), .Z(n2115) );
XOR U3527 ( .A(c705), .B(b[705]), .Z(n2116) );
XNOR U3528 ( .A(b[705]), .B(n2117), .Z(c[705]) );
XNOR U3529 ( .A(a[705]), .B(c705), .Z(n2117) );
XOR U3530 ( .A(c706), .B(n2118), .Z(c707) );
ANDN U3531 ( .B(n2119), .A(n2120), .Z(n2118) );
XOR U3532 ( .A(c706), .B(b[706]), .Z(n2119) );
XNOR U3533 ( .A(b[706]), .B(n2120), .Z(c[706]) );
XNOR U3534 ( .A(a[706]), .B(c706), .Z(n2120) );
XOR U3535 ( .A(c707), .B(n2121), .Z(c708) );
ANDN U3536 ( .B(n2122), .A(n2123), .Z(n2121) );
XOR U3537 ( .A(c707), .B(b[707]), .Z(n2122) );
XNOR U3538 ( .A(b[707]), .B(n2123), .Z(c[707]) );
XNOR U3539 ( .A(a[707]), .B(c707), .Z(n2123) );
XOR U3540 ( .A(c708), .B(n2124), .Z(c709) );
ANDN U3541 ( .B(n2125), .A(n2126), .Z(n2124) );
XOR U3542 ( .A(c708), .B(b[708]), .Z(n2125) );
XNOR U3543 ( .A(b[708]), .B(n2126), .Z(c[708]) );
XNOR U3544 ( .A(a[708]), .B(c708), .Z(n2126) );
XOR U3545 ( .A(c709), .B(n2127), .Z(c710) );
ANDN U3546 ( .B(n2128), .A(n2129), .Z(n2127) );
XOR U3547 ( .A(c709), .B(b[709]), .Z(n2128) );
XNOR U3548 ( .A(b[709]), .B(n2129), .Z(c[709]) );
XNOR U3549 ( .A(a[709]), .B(c709), .Z(n2129) );
XOR U3550 ( .A(c710), .B(n2130), .Z(c711) );
ANDN U3551 ( .B(n2131), .A(n2132), .Z(n2130) );
XOR U3552 ( .A(c710), .B(b[710]), .Z(n2131) );
XNOR U3553 ( .A(b[710]), .B(n2132), .Z(c[710]) );
XNOR U3554 ( .A(a[710]), .B(c710), .Z(n2132) );
XOR U3555 ( .A(c711), .B(n2133), .Z(c712) );
ANDN U3556 ( .B(n2134), .A(n2135), .Z(n2133) );
XOR U3557 ( .A(c711), .B(b[711]), .Z(n2134) );
XNOR U3558 ( .A(b[711]), .B(n2135), .Z(c[711]) );
XNOR U3559 ( .A(a[711]), .B(c711), .Z(n2135) );
XOR U3560 ( .A(c712), .B(n2136), .Z(c713) );
ANDN U3561 ( .B(n2137), .A(n2138), .Z(n2136) );
XOR U3562 ( .A(c712), .B(b[712]), .Z(n2137) );
XNOR U3563 ( .A(b[712]), .B(n2138), .Z(c[712]) );
XNOR U3564 ( .A(a[712]), .B(c712), .Z(n2138) );
XOR U3565 ( .A(c713), .B(n2139), .Z(c714) );
ANDN U3566 ( .B(n2140), .A(n2141), .Z(n2139) );
XOR U3567 ( .A(c713), .B(b[713]), .Z(n2140) );
XNOR U3568 ( .A(b[713]), .B(n2141), .Z(c[713]) );
XNOR U3569 ( .A(a[713]), .B(c713), .Z(n2141) );
XOR U3570 ( .A(c714), .B(n2142), .Z(c715) );
ANDN U3571 ( .B(n2143), .A(n2144), .Z(n2142) );
XOR U3572 ( .A(c714), .B(b[714]), .Z(n2143) );
XNOR U3573 ( .A(b[714]), .B(n2144), .Z(c[714]) );
XNOR U3574 ( .A(a[714]), .B(c714), .Z(n2144) );
XOR U3575 ( .A(c715), .B(n2145), .Z(c716) );
ANDN U3576 ( .B(n2146), .A(n2147), .Z(n2145) );
XOR U3577 ( .A(c715), .B(b[715]), .Z(n2146) );
XNOR U3578 ( .A(b[715]), .B(n2147), .Z(c[715]) );
XNOR U3579 ( .A(a[715]), .B(c715), .Z(n2147) );
XOR U3580 ( .A(c716), .B(n2148), .Z(c717) );
ANDN U3581 ( .B(n2149), .A(n2150), .Z(n2148) );
XOR U3582 ( .A(c716), .B(b[716]), .Z(n2149) );
XNOR U3583 ( .A(b[716]), .B(n2150), .Z(c[716]) );
XNOR U3584 ( .A(a[716]), .B(c716), .Z(n2150) );
XOR U3585 ( .A(c717), .B(n2151), .Z(c718) );
ANDN U3586 ( .B(n2152), .A(n2153), .Z(n2151) );
XOR U3587 ( .A(c717), .B(b[717]), .Z(n2152) );
XNOR U3588 ( .A(b[717]), .B(n2153), .Z(c[717]) );
XNOR U3589 ( .A(a[717]), .B(c717), .Z(n2153) );
XOR U3590 ( .A(c718), .B(n2154), .Z(c719) );
ANDN U3591 ( .B(n2155), .A(n2156), .Z(n2154) );
XOR U3592 ( .A(c718), .B(b[718]), .Z(n2155) );
XNOR U3593 ( .A(b[718]), .B(n2156), .Z(c[718]) );
XNOR U3594 ( .A(a[718]), .B(c718), .Z(n2156) );
XOR U3595 ( .A(c719), .B(n2157), .Z(c720) );
ANDN U3596 ( .B(n2158), .A(n2159), .Z(n2157) );
XOR U3597 ( .A(c719), .B(b[719]), .Z(n2158) );
XNOR U3598 ( .A(b[719]), .B(n2159), .Z(c[719]) );
XNOR U3599 ( .A(a[719]), .B(c719), .Z(n2159) );
XOR U3600 ( .A(c720), .B(n2160), .Z(c721) );
ANDN U3601 ( .B(n2161), .A(n2162), .Z(n2160) );
XOR U3602 ( .A(c720), .B(b[720]), .Z(n2161) );
XNOR U3603 ( .A(b[720]), .B(n2162), .Z(c[720]) );
XNOR U3604 ( .A(a[720]), .B(c720), .Z(n2162) );
XOR U3605 ( .A(c721), .B(n2163), .Z(c722) );
ANDN U3606 ( .B(n2164), .A(n2165), .Z(n2163) );
XOR U3607 ( .A(c721), .B(b[721]), .Z(n2164) );
XNOR U3608 ( .A(b[721]), .B(n2165), .Z(c[721]) );
XNOR U3609 ( .A(a[721]), .B(c721), .Z(n2165) );
XOR U3610 ( .A(c722), .B(n2166), .Z(c723) );
ANDN U3611 ( .B(n2167), .A(n2168), .Z(n2166) );
XOR U3612 ( .A(c722), .B(b[722]), .Z(n2167) );
XNOR U3613 ( .A(b[722]), .B(n2168), .Z(c[722]) );
XNOR U3614 ( .A(a[722]), .B(c722), .Z(n2168) );
XOR U3615 ( .A(c723), .B(n2169), .Z(c724) );
ANDN U3616 ( .B(n2170), .A(n2171), .Z(n2169) );
XOR U3617 ( .A(c723), .B(b[723]), .Z(n2170) );
XNOR U3618 ( .A(b[723]), .B(n2171), .Z(c[723]) );
XNOR U3619 ( .A(a[723]), .B(c723), .Z(n2171) );
XOR U3620 ( .A(c724), .B(n2172), .Z(c725) );
ANDN U3621 ( .B(n2173), .A(n2174), .Z(n2172) );
XOR U3622 ( .A(c724), .B(b[724]), .Z(n2173) );
XNOR U3623 ( .A(b[724]), .B(n2174), .Z(c[724]) );
XNOR U3624 ( .A(a[724]), .B(c724), .Z(n2174) );
XOR U3625 ( .A(c725), .B(n2175), .Z(c726) );
ANDN U3626 ( .B(n2176), .A(n2177), .Z(n2175) );
XOR U3627 ( .A(c725), .B(b[725]), .Z(n2176) );
XNOR U3628 ( .A(b[725]), .B(n2177), .Z(c[725]) );
XNOR U3629 ( .A(a[725]), .B(c725), .Z(n2177) );
XOR U3630 ( .A(c726), .B(n2178), .Z(c727) );
ANDN U3631 ( .B(n2179), .A(n2180), .Z(n2178) );
XOR U3632 ( .A(c726), .B(b[726]), .Z(n2179) );
XNOR U3633 ( .A(b[726]), .B(n2180), .Z(c[726]) );
XNOR U3634 ( .A(a[726]), .B(c726), .Z(n2180) );
XOR U3635 ( .A(c727), .B(n2181), .Z(c728) );
ANDN U3636 ( .B(n2182), .A(n2183), .Z(n2181) );
XOR U3637 ( .A(c727), .B(b[727]), .Z(n2182) );
XNOR U3638 ( .A(b[727]), .B(n2183), .Z(c[727]) );
XNOR U3639 ( .A(a[727]), .B(c727), .Z(n2183) );
XOR U3640 ( .A(c728), .B(n2184), .Z(c729) );
ANDN U3641 ( .B(n2185), .A(n2186), .Z(n2184) );
XOR U3642 ( .A(c728), .B(b[728]), .Z(n2185) );
XNOR U3643 ( .A(b[728]), .B(n2186), .Z(c[728]) );
XNOR U3644 ( .A(a[728]), .B(c728), .Z(n2186) );
XOR U3645 ( .A(c729), .B(n2187), .Z(c730) );
ANDN U3646 ( .B(n2188), .A(n2189), .Z(n2187) );
XOR U3647 ( .A(c729), .B(b[729]), .Z(n2188) );
XNOR U3648 ( .A(b[729]), .B(n2189), .Z(c[729]) );
XNOR U3649 ( .A(a[729]), .B(c729), .Z(n2189) );
XOR U3650 ( .A(c730), .B(n2190), .Z(c731) );
ANDN U3651 ( .B(n2191), .A(n2192), .Z(n2190) );
XOR U3652 ( .A(c730), .B(b[730]), .Z(n2191) );
XNOR U3653 ( .A(b[730]), .B(n2192), .Z(c[730]) );
XNOR U3654 ( .A(a[730]), .B(c730), .Z(n2192) );
XOR U3655 ( .A(c731), .B(n2193), .Z(c732) );
ANDN U3656 ( .B(n2194), .A(n2195), .Z(n2193) );
XOR U3657 ( .A(c731), .B(b[731]), .Z(n2194) );
XNOR U3658 ( .A(b[731]), .B(n2195), .Z(c[731]) );
XNOR U3659 ( .A(a[731]), .B(c731), .Z(n2195) );
XOR U3660 ( .A(c732), .B(n2196), .Z(c733) );
ANDN U3661 ( .B(n2197), .A(n2198), .Z(n2196) );
XOR U3662 ( .A(c732), .B(b[732]), .Z(n2197) );
XNOR U3663 ( .A(b[732]), .B(n2198), .Z(c[732]) );
XNOR U3664 ( .A(a[732]), .B(c732), .Z(n2198) );
XOR U3665 ( .A(c733), .B(n2199), .Z(c734) );
ANDN U3666 ( .B(n2200), .A(n2201), .Z(n2199) );
XOR U3667 ( .A(c733), .B(b[733]), .Z(n2200) );
XNOR U3668 ( .A(b[733]), .B(n2201), .Z(c[733]) );
XNOR U3669 ( .A(a[733]), .B(c733), .Z(n2201) );
XOR U3670 ( .A(c734), .B(n2202), .Z(c735) );
ANDN U3671 ( .B(n2203), .A(n2204), .Z(n2202) );
XOR U3672 ( .A(c734), .B(b[734]), .Z(n2203) );
XNOR U3673 ( .A(b[734]), .B(n2204), .Z(c[734]) );
XNOR U3674 ( .A(a[734]), .B(c734), .Z(n2204) );
XOR U3675 ( .A(c735), .B(n2205), .Z(c736) );
ANDN U3676 ( .B(n2206), .A(n2207), .Z(n2205) );
XOR U3677 ( .A(c735), .B(b[735]), .Z(n2206) );
XNOR U3678 ( .A(b[735]), .B(n2207), .Z(c[735]) );
XNOR U3679 ( .A(a[735]), .B(c735), .Z(n2207) );
XOR U3680 ( .A(c736), .B(n2208), .Z(c737) );
ANDN U3681 ( .B(n2209), .A(n2210), .Z(n2208) );
XOR U3682 ( .A(c736), .B(b[736]), .Z(n2209) );
XNOR U3683 ( .A(b[736]), .B(n2210), .Z(c[736]) );
XNOR U3684 ( .A(a[736]), .B(c736), .Z(n2210) );
XOR U3685 ( .A(c737), .B(n2211), .Z(c738) );
ANDN U3686 ( .B(n2212), .A(n2213), .Z(n2211) );
XOR U3687 ( .A(c737), .B(b[737]), .Z(n2212) );
XNOR U3688 ( .A(b[737]), .B(n2213), .Z(c[737]) );
XNOR U3689 ( .A(a[737]), .B(c737), .Z(n2213) );
XOR U3690 ( .A(c738), .B(n2214), .Z(c739) );
ANDN U3691 ( .B(n2215), .A(n2216), .Z(n2214) );
XOR U3692 ( .A(c738), .B(b[738]), .Z(n2215) );
XNOR U3693 ( .A(b[738]), .B(n2216), .Z(c[738]) );
XNOR U3694 ( .A(a[738]), .B(c738), .Z(n2216) );
XOR U3695 ( .A(c739), .B(n2217), .Z(c740) );
ANDN U3696 ( .B(n2218), .A(n2219), .Z(n2217) );
XOR U3697 ( .A(c739), .B(b[739]), .Z(n2218) );
XNOR U3698 ( .A(b[739]), .B(n2219), .Z(c[739]) );
XNOR U3699 ( .A(a[739]), .B(c739), .Z(n2219) );
XOR U3700 ( .A(c740), .B(n2220), .Z(c741) );
ANDN U3701 ( .B(n2221), .A(n2222), .Z(n2220) );
XOR U3702 ( .A(c740), .B(b[740]), .Z(n2221) );
XNOR U3703 ( .A(b[740]), .B(n2222), .Z(c[740]) );
XNOR U3704 ( .A(a[740]), .B(c740), .Z(n2222) );
XOR U3705 ( .A(c741), .B(n2223), .Z(c742) );
ANDN U3706 ( .B(n2224), .A(n2225), .Z(n2223) );
XOR U3707 ( .A(c741), .B(b[741]), .Z(n2224) );
XNOR U3708 ( .A(b[741]), .B(n2225), .Z(c[741]) );
XNOR U3709 ( .A(a[741]), .B(c741), .Z(n2225) );
XOR U3710 ( .A(c742), .B(n2226), .Z(c743) );
ANDN U3711 ( .B(n2227), .A(n2228), .Z(n2226) );
XOR U3712 ( .A(c742), .B(b[742]), .Z(n2227) );
XNOR U3713 ( .A(b[742]), .B(n2228), .Z(c[742]) );
XNOR U3714 ( .A(a[742]), .B(c742), .Z(n2228) );
XOR U3715 ( .A(c743), .B(n2229), .Z(c744) );
ANDN U3716 ( .B(n2230), .A(n2231), .Z(n2229) );
XOR U3717 ( .A(c743), .B(b[743]), .Z(n2230) );
XNOR U3718 ( .A(b[743]), .B(n2231), .Z(c[743]) );
XNOR U3719 ( .A(a[743]), .B(c743), .Z(n2231) );
XOR U3720 ( .A(c744), .B(n2232), .Z(c745) );
ANDN U3721 ( .B(n2233), .A(n2234), .Z(n2232) );
XOR U3722 ( .A(c744), .B(b[744]), .Z(n2233) );
XNOR U3723 ( .A(b[744]), .B(n2234), .Z(c[744]) );
XNOR U3724 ( .A(a[744]), .B(c744), .Z(n2234) );
XOR U3725 ( .A(c745), .B(n2235), .Z(c746) );
ANDN U3726 ( .B(n2236), .A(n2237), .Z(n2235) );
XOR U3727 ( .A(c745), .B(b[745]), .Z(n2236) );
XNOR U3728 ( .A(b[745]), .B(n2237), .Z(c[745]) );
XNOR U3729 ( .A(a[745]), .B(c745), .Z(n2237) );
XOR U3730 ( .A(c746), .B(n2238), .Z(c747) );
ANDN U3731 ( .B(n2239), .A(n2240), .Z(n2238) );
XOR U3732 ( .A(c746), .B(b[746]), .Z(n2239) );
XNOR U3733 ( .A(b[746]), .B(n2240), .Z(c[746]) );
XNOR U3734 ( .A(a[746]), .B(c746), .Z(n2240) );
XOR U3735 ( .A(c747), .B(n2241), .Z(c748) );
ANDN U3736 ( .B(n2242), .A(n2243), .Z(n2241) );
XOR U3737 ( .A(c747), .B(b[747]), .Z(n2242) );
XNOR U3738 ( .A(b[747]), .B(n2243), .Z(c[747]) );
XNOR U3739 ( .A(a[747]), .B(c747), .Z(n2243) );
XOR U3740 ( .A(c748), .B(n2244), .Z(c749) );
ANDN U3741 ( .B(n2245), .A(n2246), .Z(n2244) );
XOR U3742 ( .A(c748), .B(b[748]), .Z(n2245) );
XNOR U3743 ( .A(b[748]), .B(n2246), .Z(c[748]) );
XNOR U3744 ( .A(a[748]), .B(c748), .Z(n2246) );
XOR U3745 ( .A(c749), .B(n2247), .Z(c750) );
ANDN U3746 ( .B(n2248), .A(n2249), .Z(n2247) );
XOR U3747 ( .A(c749), .B(b[749]), .Z(n2248) );
XNOR U3748 ( .A(b[749]), .B(n2249), .Z(c[749]) );
XNOR U3749 ( .A(a[749]), .B(c749), .Z(n2249) );
XOR U3750 ( .A(c750), .B(n2250), .Z(c751) );
ANDN U3751 ( .B(n2251), .A(n2252), .Z(n2250) );
XOR U3752 ( .A(c750), .B(b[750]), .Z(n2251) );
XNOR U3753 ( .A(b[750]), .B(n2252), .Z(c[750]) );
XNOR U3754 ( .A(a[750]), .B(c750), .Z(n2252) );
XOR U3755 ( .A(c751), .B(n2253), .Z(c752) );
ANDN U3756 ( .B(n2254), .A(n2255), .Z(n2253) );
XOR U3757 ( .A(c751), .B(b[751]), .Z(n2254) );
XNOR U3758 ( .A(b[751]), .B(n2255), .Z(c[751]) );
XNOR U3759 ( .A(a[751]), .B(c751), .Z(n2255) );
XOR U3760 ( .A(c752), .B(n2256), .Z(c753) );
ANDN U3761 ( .B(n2257), .A(n2258), .Z(n2256) );
XOR U3762 ( .A(c752), .B(b[752]), .Z(n2257) );
XNOR U3763 ( .A(b[752]), .B(n2258), .Z(c[752]) );
XNOR U3764 ( .A(a[752]), .B(c752), .Z(n2258) );
XOR U3765 ( .A(c753), .B(n2259), .Z(c754) );
ANDN U3766 ( .B(n2260), .A(n2261), .Z(n2259) );
XOR U3767 ( .A(c753), .B(b[753]), .Z(n2260) );
XNOR U3768 ( .A(b[753]), .B(n2261), .Z(c[753]) );
XNOR U3769 ( .A(a[753]), .B(c753), .Z(n2261) );
XOR U3770 ( .A(c754), .B(n2262), .Z(c755) );
ANDN U3771 ( .B(n2263), .A(n2264), .Z(n2262) );
XOR U3772 ( .A(c754), .B(b[754]), .Z(n2263) );
XNOR U3773 ( .A(b[754]), .B(n2264), .Z(c[754]) );
XNOR U3774 ( .A(a[754]), .B(c754), .Z(n2264) );
XOR U3775 ( .A(c755), .B(n2265), .Z(c756) );
ANDN U3776 ( .B(n2266), .A(n2267), .Z(n2265) );
XOR U3777 ( .A(c755), .B(b[755]), .Z(n2266) );
XNOR U3778 ( .A(b[755]), .B(n2267), .Z(c[755]) );
XNOR U3779 ( .A(a[755]), .B(c755), .Z(n2267) );
XOR U3780 ( .A(c756), .B(n2268), .Z(c757) );
ANDN U3781 ( .B(n2269), .A(n2270), .Z(n2268) );
XOR U3782 ( .A(c756), .B(b[756]), .Z(n2269) );
XNOR U3783 ( .A(b[756]), .B(n2270), .Z(c[756]) );
XNOR U3784 ( .A(a[756]), .B(c756), .Z(n2270) );
XOR U3785 ( .A(c757), .B(n2271), .Z(c758) );
ANDN U3786 ( .B(n2272), .A(n2273), .Z(n2271) );
XOR U3787 ( .A(c757), .B(b[757]), .Z(n2272) );
XNOR U3788 ( .A(b[757]), .B(n2273), .Z(c[757]) );
XNOR U3789 ( .A(a[757]), .B(c757), .Z(n2273) );
XOR U3790 ( .A(c758), .B(n2274), .Z(c759) );
ANDN U3791 ( .B(n2275), .A(n2276), .Z(n2274) );
XOR U3792 ( .A(c758), .B(b[758]), .Z(n2275) );
XNOR U3793 ( .A(b[758]), .B(n2276), .Z(c[758]) );
XNOR U3794 ( .A(a[758]), .B(c758), .Z(n2276) );
XOR U3795 ( .A(c759), .B(n2277), .Z(c760) );
ANDN U3796 ( .B(n2278), .A(n2279), .Z(n2277) );
XOR U3797 ( .A(c759), .B(b[759]), .Z(n2278) );
XNOR U3798 ( .A(b[759]), .B(n2279), .Z(c[759]) );
XNOR U3799 ( .A(a[759]), .B(c759), .Z(n2279) );
XOR U3800 ( .A(c760), .B(n2280), .Z(c761) );
ANDN U3801 ( .B(n2281), .A(n2282), .Z(n2280) );
XOR U3802 ( .A(c760), .B(b[760]), .Z(n2281) );
XNOR U3803 ( .A(b[760]), .B(n2282), .Z(c[760]) );
XNOR U3804 ( .A(a[760]), .B(c760), .Z(n2282) );
XOR U3805 ( .A(c761), .B(n2283), .Z(c762) );
ANDN U3806 ( .B(n2284), .A(n2285), .Z(n2283) );
XOR U3807 ( .A(c761), .B(b[761]), .Z(n2284) );
XNOR U3808 ( .A(b[761]), .B(n2285), .Z(c[761]) );
XNOR U3809 ( .A(a[761]), .B(c761), .Z(n2285) );
XOR U3810 ( .A(c762), .B(n2286), .Z(c763) );
ANDN U3811 ( .B(n2287), .A(n2288), .Z(n2286) );
XOR U3812 ( .A(c762), .B(b[762]), .Z(n2287) );
XNOR U3813 ( .A(b[762]), .B(n2288), .Z(c[762]) );
XNOR U3814 ( .A(a[762]), .B(c762), .Z(n2288) );
XOR U3815 ( .A(c763), .B(n2289), .Z(c764) );
ANDN U3816 ( .B(n2290), .A(n2291), .Z(n2289) );
XOR U3817 ( .A(c763), .B(b[763]), .Z(n2290) );
XNOR U3818 ( .A(b[763]), .B(n2291), .Z(c[763]) );
XNOR U3819 ( .A(a[763]), .B(c763), .Z(n2291) );
XOR U3820 ( .A(c764), .B(n2292), .Z(c765) );
ANDN U3821 ( .B(n2293), .A(n2294), .Z(n2292) );
XOR U3822 ( .A(c764), .B(b[764]), .Z(n2293) );
XNOR U3823 ( .A(b[764]), .B(n2294), .Z(c[764]) );
XNOR U3824 ( .A(a[764]), .B(c764), .Z(n2294) );
XOR U3825 ( .A(c765), .B(n2295), .Z(c766) );
ANDN U3826 ( .B(n2296), .A(n2297), .Z(n2295) );
XOR U3827 ( .A(c765), .B(b[765]), .Z(n2296) );
XNOR U3828 ( .A(b[765]), .B(n2297), .Z(c[765]) );
XNOR U3829 ( .A(a[765]), .B(c765), .Z(n2297) );
XOR U3830 ( .A(c766), .B(n2298), .Z(c767) );
ANDN U3831 ( .B(n2299), .A(n2300), .Z(n2298) );
XOR U3832 ( .A(c766), .B(b[766]), .Z(n2299) );
XNOR U3833 ( .A(b[766]), .B(n2300), .Z(c[766]) );
XNOR U3834 ( .A(a[766]), .B(c766), .Z(n2300) );
XOR U3835 ( .A(c767), .B(n2301), .Z(c768) );
ANDN U3836 ( .B(n2302), .A(n2303), .Z(n2301) );
XOR U3837 ( .A(c767), .B(b[767]), .Z(n2302) );
XNOR U3838 ( .A(b[767]), .B(n2303), .Z(c[767]) );
XNOR U3839 ( .A(a[767]), .B(c767), .Z(n2303) );
XOR U3840 ( .A(c768), .B(n2304), .Z(c769) );
ANDN U3841 ( .B(n2305), .A(n2306), .Z(n2304) );
XOR U3842 ( .A(c768), .B(b[768]), .Z(n2305) );
XNOR U3843 ( .A(b[768]), .B(n2306), .Z(c[768]) );
XNOR U3844 ( .A(a[768]), .B(c768), .Z(n2306) );
XOR U3845 ( .A(c769), .B(n2307), .Z(c770) );
ANDN U3846 ( .B(n2308), .A(n2309), .Z(n2307) );
XOR U3847 ( .A(c769), .B(b[769]), .Z(n2308) );
XNOR U3848 ( .A(b[769]), .B(n2309), .Z(c[769]) );
XNOR U3849 ( .A(a[769]), .B(c769), .Z(n2309) );
XOR U3850 ( .A(c770), .B(n2310), .Z(c771) );
ANDN U3851 ( .B(n2311), .A(n2312), .Z(n2310) );
XOR U3852 ( .A(c770), .B(b[770]), .Z(n2311) );
XNOR U3853 ( .A(b[770]), .B(n2312), .Z(c[770]) );
XNOR U3854 ( .A(a[770]), .B(c770), .Z(n2312) );
XOR U3855 ( .A(c771), .B(n2313), .Z(c772) );
ANDN U3856 ( .B(n2314), .A(n2315), .Z(n2313) );
XOR U3857 ( .A(c771), .B(b[771]), .Z(n2314) );
XNOR U3858 ( .A(b[771]), .B(n2315), .Z(c[771]) );
XNOR U3859 ( .A(a[771]), .B(c771), .Z(n2315) );
XOR U3860 ( .A(c772), .B(n2316), .Z(c773) );
ANDN U3861 ( .B(n2317), .A(n2318), .Z(n2316) );
XOR U3862 ( .A(c772), .B(b[772]), .Z(n2317) );
XNOR U3863 ( .A(b[772]), .B(n2318), .Z(c[772]) );
XNOR U3864 ( .A(a[772]), .B(c772), .Z(n2318) );
XOR U3865 ( .A(c773), .B(n2319), .Z(c774) );
ANDN U3866 ( .B(n2320), .A(n2321), .Z(n2319) );
XOR U3867 ( .A(c773), .B(b[773]), .Z(n2320) );
XNOR U3868 ( .A(b[773]), .B(n2321), .Z(c[773]) );
XNOR U3869 ( .A(a[773]), .B(c773), .Z(n2321) );
XOR U3870 ( .A(c774), .B(n2322), .Z(c775) );
ANDN U3871 ( .B(n2323), .A(n2324), .Z(n2322) );
XOR U3872 ( .A(c774), .B(b[774]), .Z(n2323) );
XNOR U3873 ( .A(b[774]), .B(n2324), .Z(c[774]) );
XNOR U3874 ( .A(a[774]), .B(c774), .Z(n2324) );
XOR U3875 ( .A(c775), .B(n2325), .Z(c776) );
ANDN U3876 ( .B(n2326), .A(n2327), .Z(n2325) );
XOR U3877 ( .A(c775), .B(b[775]), .Z(n2326) );
XNOR U3878 ( .A(b[775]), .B(n2327), .Z(c[775]) );
XNOR U3879 ( .A(a[775]), .B(c775), .Z(n2327) );
XOR U3880 ( .A(c776), .B(n2328), .Z(c777) );
ANDN U3881 ( .B(n2329), .A(n2330), .Z(n2328) );
XOR U3882 ( .A(c776), .B(b[776]), .Z(n2329) );
XNOR U3883 ( .A(b[776]), .B(n2330), .Z(c[776]) );
XNOR U3884 ( .A(a[776]), .B(c776), .Z(n2330) );
XOR U3885 ( .A(c777), .B(n2331), .Z(c778) );
ANDN U3886 ( .B(n2332), .A(n2333), .Z(n2331) );
XOR U3887 ( .A(c777), .B(b[777]), .Z(n2332) );
XNOR U3888 ( .A(b[777]), .B(n2333), .Z(c[777]) );
XNOR U3889 ( .A(a[777]), .B(c777), .Z(n2333) );
XOR U3890 ( .A(c778), .B(n2334), .Z(c779) );
ANDN U3891 ( .B(n2335), .A(n2336), .Z(n2334) );
XOR U3892 ( .A(c778), .B(b[778]), .Z(n2335) );
XNOR U3893 ( .A(b[778]), .B(n2336), .Z(c[778]) );
XNOR U3894 ( .A(a[778]), .B(c778), .Z(n2336) );
XOR U3895 ( .A(c779), .B(n2337), .Z(c780) );
ANDN U3896 ( .B(n2338), .A(n2339), .Z(n2337) );
XOR U3897 ( .A(c779), .B(b[779]), .Z(n2338) );
XNOR U3898 ( .A(b[779]), .B(n2339), .Z(c[779]) );
XNOR U3899 ( .A(a[779]), .B(c779), .Z(n2339) );
XOR U3900 ( .A(c780), .B(n2340), .Z(c781) );
ANDN U3901 ( .B(n2341), .A(n2342), .Z(n2340) );
XOR U3902 ( .A(c780), .B(b[780]), .Z(n2341) );
XNOR U3903 ( .A(b[780]), .B(n2342), .Z(c[780]) );
XNOR U3904 ( .A(a[780]), .B(c780), .Z(n2342) );
XOR U3905 ( .A(c781), .B(n2343), .Z(c782) );
ANDN U3906 ( .B(n2344), .A(n2345), .Z(n2343) );
XOR U3907 ( .A(c781), .B(b[781]), .Z(n2344) );
XNOR U3908 ( .A(b[781]), .B(n2345), .Z(c[781]) );
XNOR U3909 ( .A(a[781]), .B(c781), .Z(n2345) );
XOR U3910 ( .A(c782), .B(n2346), .Z(c783) );
ANDN U3911 ( .B(n2347), .A(n2348), .Z(n2346) );
XOR U3912 ( .A(c782), .B(b[782]), .Z(n2347) );
XNOR U3913 ( .A(b[782]), .B(n2348), .Z(c[782]) );
XNOR U3914 ( .A(a[782]), .B(c782), .Z(n2348) );
XOR U3915 ( .A(c783), .B(n2349), .Z(c784) );
ANDN U3916 ( .B(n2350), .A(n2351), .Z(n2349) );
XOR U3917 ( .A(c783), .B(b[783]), .Z(n2350) );
XNOR U3918 ( .A(b[783]), .B(n2351), .Z(c[783]) );
XNOR U3919 ( .A(a[783]), .B(c783), .Z(n2351) );
XOR U3920 ( .A(c784), .B(n2352), .Z(c785) );
ANDN U3921 ( .B(n2353), .A(n2354), .Z(n2352) );
XOR U3922 ( .A(c784), .B(b[784]), .Z(n2353) );
XNOR U3923 ( .A(b[784]), .B(n2354), .Z(c[784]) );
XNOR U3924 ( .A(a[784]), .B(c784), .Z(n2354) );
XOR U3925 ( .A(c785), .B(n2355), .Z(c786) );
ANDN U3926 ( .B(n2356), .A(n2357), .Z(n2355) );
XOR U3927 ( .A(c785), .B(b[785]), .Z(n2356) );
XNOR U3928 ( .A(b[785]), .B(n2357), .Z(c[785]) );
XNOR U3929 ( .A(a[785]), .B(c785), .Z(n2357) );
XOR U3930 ( .A(c786), .B(n2358), .Z(c787) );
ANDN U3931 ( .B(n2359), .A(n2360), .Z(n2358) );
XOR U3932 ( .A(c786), .B(b[786]), .Z(n2359) );
XNOR U3933 ( .A(b[786]), .B(n2360), .Z(c[786]) );
XNOR U3934 ( .A(a[786]), .B(c786), .Z(n2360) );
XOR U3935 ( .A(c787), .B(n2361), .Z(c788) );
ANDN U3936 ( .B(n2362), .A(n2363), .Z(n2361) );
XOR U3937 ( .A(c787), .B(b[787]), .Z(n2362) );
XNOR U3938 ( .A(b[787]), .B(n2363), .Z(c[787]) );
XNOR U3939 ( .A(a[787]), .B(c787), .Z(n2363) );
XOR U3940 ( .A(c788), .B(n2364), .Z(c789) );
ANDN U3941 ( .B(n2365), .A(n2366), .Z(n2364) );
XOR U3942 ( .A(c788), .B(b[788]), .Z(n2365) );
XNOR U3943 ( .A(b[788]), .B(n2366), .Z(c[788]) );
XNOR U3944 ( .A(a[788]), .B(c788), .Z(n2366) );
XOR U3945 ( .A(c789), .B(n2367), .Z(c790) );
ANDN U3946 ( .B(n2368), .A(n2369), .Z(n2367) );
XOR U3947 ( .A(c789), .B(b[789]), .Z(n2368) );
XNOR U3948 ( .A(b[789]), .B(n2369), .Z(c[789]) );
XNOR U3949 ( .A(a[789]), .B(c789), .Z(n2369) );
XOR U3950 ( .A(c790), .B(n2370), .Z(c791) );
ANDN U3951 ( .B(n2371), .A(n2372), .Z(n2370) );
XOR U3952 ( .A(c790), .B(b[790]), .Z(n2371) );
XNOR U3953 ( .A(b[790]), .B(n2372), .Z(c[790]) );
XNOR U3954 ( .A(a[790]), .B(c790), .Z(n2372) );
XOR U3955 ( .A(c791), .B(n2373), .Z(c792) );
ANDN U3956 ( .B(n2374), .A(n2375), .Z(n2373) );
XOR U3957 ( .A(c791), .B(b[791]), .Z(n2374) );
XNOR U3958 ( .A(b[791]), .B(n2375), .Z(c[791]) );
XNOR U3959 ( .A(a[791]), .B(c791), .Z(n2375) );
XOR U3960 ( .A(c792), .B(n2376), .Z(c793) );
ANDN U3961 ( .B(n2377), .A(n2378), .Z(n2376) );
XOR U3962 ( .A(c792), .B(b[792]), .Z(n2377) );
XNOR U3963 ( .A(b[792]), .B(n2378), .Z(c[792]) );
XNOR U3964 ( .A(a[792]), .B(c792), .Z(n2378) );
XOR U3965 ( .A(c793), .B(n2379), .Z(c794) );
ANDN U3966 ( .B(n2380), .A(n2381), .Z(n2379) );
XOR U3967 ( .A(c793), .B(b[793]), .Z(n2380) );
XNOR U3968 ( .A(b[793]), .B(n2381), .Z(c[793]) );
XNOR U3969 ( .A(a[793]), .B(c793), .Z(n2381) );
XOR U3970 ( .A(c794), .B(n2382), .Z(c795) );
ANDN U3971 ( .B(n2383), .A(n2384), .Z(n2382) );
XOR U3972 ( .A(c794), .B(b[794]), .Z(n2383) );
XNOR U3973 ( .A(b[794]), .B(n2384), .Z(c[794]) );
XNOR U3974 ( .A(a[794]), .B(c794), .Z(n2384) );
XOR U3975 ( .A(c795), .B(n2385), .Z(c796) );
ANDN U3976 ( .B(n2386), .A(n2387), .Z(n2385) );
XOR U3977 ( .A(c795), .B(b[795]), .Z(n2386) );
XNOR U3978 ( .A(b[795]), .B(n2387), .Z(c[795]) );
XNOR U3979 ( .A(a[795]), .B(c795), .Z(n2387) );
XOR U3980 ( .A(c796), .B(n2388), .Z(c797) );
ANDN U3981 ( .B(n2389), .A(n2390), .Z(n2388) );
XOR U3982 ( .A(c796), .B(b[796]), .Z(n2389) );
XNOR U3983 ( .A(b[796]), .B(n2390), .Z(c[796]) );
XNOR U3984 ( .A(a[796]), .B(c796), .Z(n2390) );
XOR U3985 ( .A(c797), .B(n2391), .Z(c798) );
ANDN U3986 ( .B(n2392), .A(n2393), .Z(n2391) );
XOR U3987 ( .A(c797), .B(b[797]), .Z(n2392) );
XNOR U3988 ( .A(b[797]), .B(n2393), .Z(c[797]) );
XNOR U3989 ( .A(a[797]), .B(c797), .Z(n2393) );
XOR U3990 ( .A(c798), .B(n2394), .Z(c799) );
ANDN U3991 ( .B(n2395), .A(n2396), .Z(n2394) );
XOR U3992 ( .A(c798), .B(b[798]), .Z(n2395) );
XNOR U3993 ( .A(b[798]), .B(n2396), .Z(c[798]) );
XNOR U3994 ( .A(a[798]), .B(c798), .Z(n2396) );
XOR U3995 ( .A(c799), .B(n2397), .Z(c800) );
ANDN U3996 ( .B(n2398), .A(n2399), .Z(n2397) );
XOR U3997 ( .A(c799), .B(b[799]), .Z(n2398) );
XNOR U3998 ( .A(b[799]), .B(n2399), .Z(c[799]) );
XNOR U3999 ( .A(a[799]), .B(c799), .Z(n2399) );
XOR U4000 ( .A(c800), .B(n2400), .Z(c801) );
ANDN U4001 ( .B(n2401), .A(n2402), .Z(n2400) );
XOR U4002 ( .A(c800), .B(b[800]), .Z(n2401) );
XNOR U4003 ( .A(b[800]), .B(n2402), .Z(c[800]) );
XNOR U4004 ( .A(a[800]), .B(c800), .Z(n2402) );
XOR U4005 ( .A(c801), .B(n2403), .Z(c802) );
ANDN U4006 ( .B(n2404), .A(n2405), .Z(n2403) );
XOR U4007 ( .A(c801), .B(b[801]), .Z(n2404) );
XNOR U4008 ( .A(b[801]), .B(n2405), .Z(c[801]) );
XNOR U4009 ( .A(a[801]), .B(c801), .Z(n2405) );
XOR U4010 ( .A(c802), .B(n2406), .Z(c803) );
ANDN U4011 ( .B(n2407), .A(n2408), .Z(n2406) );
XOR U4012 ( .A(c802), .B(b[802]), .Z(n2407) );
XNOR U4013 ( .A(b[802]), .B(n2408), .Z(c[802]) );
XNOR U4014 ( .A(a[802]), .B(c802), .Z(n2408) );
XOR U4015 ( .A(c803), .B(n2409), .Z(c804) );
ANDN U4016 ( .B(n2410), .A(n2411), .Z(n2409) );
XOR U4017 ( .A(c803), .B(b[803]), .Z(n2410) );
XNOR U4018 ( .A(b[803]), .B(n2411), .Z(c[803]) );
XNOR U4019 ( .A(a[803]), .B(c803), .Z(n2411) );
XOR U4020 ( .A(c804), .B(n2412), .Z(c805) );
ANDN U4021 ( .B(n2413), .A(n2414), .Z(n2412) );
XOR U4022 ( .A(c804), .B(b[804]), .Z(n2413) );
XNOR U4023 ( .A(b[804]), .B(n2414), .Z(c[804]) );
XNOR U4024 ( .A(a[804]), .B(c804), .Z(n2414) );
XOR U4025 ( .A(c805), .B(n2415), .Z(c806) );
ANDN U4026 ( .B(n2416), .A(n2417), .Z(n2415) );
XOR U4027 ( .A(c805), .B(b[805]), .Z(n2416) );
XNOR U4028 ( .A(b[805]), .B(n2417), .Z(c[805]) );
XNOR U4029 ( .A(a[805]), .B(c805), .Z(n2417) );
XOR U4030 ( .A(c806), .B(n2418), .Z(c807) );
ANDN U4031 ( .B(n2419), .A(n2420), .Z(n2418) );
XOR U4032 ( .A(c806), .B(b[806]), .Z(n2419) );
XNOR U4033 ( .A(b[806]), .B(n2420), .Z(c[806]) );
XNOR U4034 ( .A(a[806]), .B(c806), .Z(n2420) );
XOR U4035 ( .A(c807), .B(n2421), .Z(c808) );
ANDN U4036 ( .B(n2422), .A(n2423), .Z(n2421) );
XOR U4037 ( .A(c807), .B(b[807]), .Z(n2422) );
XNOR U4038 ( .A(b[807]), .B(n2423), .Z(c[807]) );
XNOR U4039 ( .A(a[807]), .B(c807), .Z(n2423) );
XOR U4040 ( .A(c808), .B(n2424), .Z(c809) );
ANDN U4041 ( .B(n2425), .A(n2426), .Z(n2424) );
XOR U4042 ( .A(c808), .B(b[808]), .Z(n2425) );
XNOR U4043 ( .A(b[808]), .B(n2426), .Z(c[808]) );
XNOR U4044 ( .A(a[808]), .B(c808), .Z(n2426) );
XOR U4045 ( .A(c809), .B(n2427), .Z(c810) );
ANDN U4046 ( .B(n2428), .A(n2429), .Z(n2427) );
XOR U4047 ( .A(c809), .B(b[809]), .Z(n2428) );
XNOR U4048 ( .A(b[809]), .B(n2429), .Z(c[809]) );
XNOR U4049 ( .A(a[809]), .B(c809), .Z(n2429) );
XOR U4050 ( .A(c810), .B(n2430), .Z(c811) );
ANDN U4051 ( .B(n2431), .A(n2432), .Z(n2430) );
XOR U4052 ( .A(c810), .B(b[810]), .Z(n2431) );
XNOR U4053 ( .A(b[810]), .B(n2432), .Z(c[810]) );
XNOR U4054 ( .A(a[810]), .B(c810), .Z(n2432) );
XOR U4055 ( .A(c811), .B(n2433), .Z(c812) );
ANDN U4056 ( .B(n2434), .A(n2435), .Z(n2433) );
XOR U4057 ( .A(c811), .B(b[811]), .Z(n2434) );
XNOR U4058 ( .A(b[811]), .B(n2435), .Z(c[811]) );
XNOR U4059 ( .A(a[811]), .B(c811), .Z(n2435) );
XOR U4060 ( .A(c812), .B(n2436), .Z(c813) );
ANDN U4061 ( .B(n2437), .A(n2438), .Z(n2436) );
XOR U4062 ( .A(c812), .B(b[812]), .Z(n2437) );
XNOR U4063 ( .A(b[812]), .B(n2438), .Z(c[812]) );
XNOR U4064 ( .A(a[812]), .B(c812), .Z(n2438) );
XOR U4065 ( .A(c813), .B(n2439), .Z(c814) );
ANDN U4066 ( .B(n2440), .A(n2441), .Z(n2439) );
XOR U4067 ( .A(c813), .B(b[813]), .Z(n2440) );
XNOR U4068 ( .A(b[813]), .B(n2441), .Z(c[813]) );
XNOR U4069 ( .A(a[813]), .B(c813), .Z(n2441) );
XOR U4070 ( .A(c814), .B(n2442), .Z(c815) );
ANDN U4071 ( .B(n2443), .A(n2444), .Z(n2442) );
XOR U4072 ( .A(c814), .B(b[814]), .Z(n2443) );
XNOR U4073 ( .A(b[814]), .B(n2444), .Z(c[814]) );
XNOR U4074 ( .A(a[814]), .B(c814), .Z(n2444) );
XOR U4075 ( .A(c815), .B(n2445), .Z(c816) );
ANDN U4076 ( .B(n2446), .A(n2447), .Z(n2445) );
XOR U4077 ( .A(c815), .B(b[815]), .Z(n2446) );
XNOR U4078 ( .A(b[815]), .B(n2447), .Z(c[815]) );
XNOR U4079 ( .A(a[815]), .B(c815), .Z(n2447) );
XOR U4080 ( .A(c816), .B(n2448), .Z(c817) );
ANDN U4081 ( .B(n2449), .A(n2450), .Z(n2448) );
XOR U4082 ( .A(c816), .B(b[816]), .Z(n2449) );
XNOR U4083 ( .A(b[816]), .B(n2450), .Z(c[816]) );
XNOR U4084 ( .A(a[816]), .B(c816), .Z(n2450) );
XOR U4085 ( .A(c817), .B(n2451), .Z(c818) );
ANDN U4086 ( .B(n2452), .A(n2453), .Z(n2451) );
XOR U4087 ( .A(c817), .B(b[817]), .Z(n2452) );
XNOR U4088 ( .A(b[817]), .B(n2453), .Z(c[817]) );
XNOR U4089 ( .A(a[817]), .B(c817), .Z(n2453) );
XOR U4090 ( .A(c818), .B(n2454), .Z(c819) );
ANDN U4091 ( .B(n2455), .A(n2456), .Z(n2454) );
XOR U4092 ( .A(c818), .B(b[818]), .Z(n2455) );
XNOR U4093 ( .A(b[818]), .B(n2456), .Z(c[818]) );
XNOR U4094 ( .A(a[818]), .B(c818), .Z(n2456) );
XOR U4095 ( .A(c819), .B(n2457), .Z(c820) );
ANDN U4096 ( .B(n2458), .A(n2459), .Z(n2457) );
XOR U4097 ( .A(c819), .B(b[819]), .Z(n2458) );
XNOR U4098 ( .A(b[819]), .B(n2459), .Z(c[819]) );
XNOR U4099 ( .A(a[819]), .B(c819), .Z(n2459) );
XOR U4100 ( .A(c820), .B(n2460), .Z(c821) );
ANDN U4101 ( .B(n2461), .A(n2462), .Z(n2460) );
XOR U4102 ( .A(c820), .B(b[820]), .Z(n2461) );
XNOR U4103 ( .A(b[820]), .B(n2462), .Z(c[820]) );
XNOR U4104 ( .A(a[820]), .B(c820), .Z(n2462) );
XOR U4105 ( .A(c821), .B(n2463), .Z(c822) );
ANDN U4106 ( .B(n2464), .A(n2465), .Z(n2463) );
XOR U4107 ( .A(c821), .B(b[821]), .Z(n2464) );
XNOR U4108 ( .A(b[821]), .B(n2465), .Z(c[821]) );
XNOR U4109 ( .A(a[821]), .B(c821), .Z(n2465) );
XOR U4110 ( .A(c822), .B(n2466), .Z(c823) );
ANDN U4111 ( .B(n2467), .A(n2468), .Z(n2466) );
XOR U4112 ( .A(c822), .B(b[822]), .Z(n2467) );
XNOR U4113 ( .A(b[822]), .B(n2468), .Z(c[822]) );
XNOR U4114 ( .A(a[822]), .B(c822), .Z(n2468) );
XOR U4115 ( .A(c823), .B(n2469), .Z(c824) );
ANDN U4116 ( .B(n2470), .A(n2471), .Z(n2469) );
XOR U4117 ( .A(c823), .B(b[823]), .Z(n2470) );
XNOR U4118 ( .A(b[823]), .B(n2471), .Z(c[823]) );
XNOR U4119 ( .A(a[823]), .B(c823), .Z(n2471) );
XOR U4120 ( .A(c824), .B(n2472), .Z(c825) );
ANDN U4121 ( .B(n2473), .A(n2474), .Z(n2472) );
XOR U4122 ( .A(c824), .B(b[824]), .Z(n2473) );
XNOR U4123 ( .A(b[824]), .B(n2474), .Z(c[824]) );
XNOR U4124 ( .A(a[824]), .B(c824), .Z(n2474) );
XOR U4125 ( .A(c825), .B(n2475), .Z(c826) );
ANDN U4126 ( .B(n2476), .A(n2477), .Z(n2475) );
XOR U4127 ( .A(c825), .B(b[825]), .Z(n2476) );
XNOR U4128 ( .A(b[825]), .B(n2477), .Z(c[825]) );
XNOR U4129 ( .A(a[825]), .B(c825), .Z(n2477) );
XOR U4130 ( .A(c826), .B(n2478), .Z(c827) );
ANDN U4131 ( .B(n2479), .A(n2480), .Z(n2478) );
XOR U4132 ( .A(c826), .B(b[826]), .Z(n2479) );
XNOR U4133 ( .A(b[826]), .B(n2480), .Z(c[826]) );
XNOR U4134 ( .A(a[826]), .B(c826), .Z(n2480) );
XOR U4135 ( .A(c827), .B(n2481), .Z(c828) );
ANDN U4136 ( .B(n2482), .A(n2483), .Z(n2481) );
XOR U4137 ( .A(c827), .B(b[827]), .Z(n2482) );
XNOR U4138 ( .A(b[827]), .B(n2483), .Z(c[827]) );
XNOR U4139 ( .A(a[827]), .B(c827), .Z(n2483) );
XOR U4140 ( .A(c828), .B(n2484), .Z(c829) );
ANDN U4141 ( .B(n2485), .A(n2486), .Z(n2484) );
XOR U4142 ( .A(c828), .B(b[828]), .Z(n2485) );
XNOR U4143 ( .A(b[828]), .B(n2486), .Z(c[828]) );
XNOR U4144 ( .A(a[828]), .B(c828), .Z(n2486) );
XOR U4145 ( .A(c829), .B(n2487), .Z(c830) );
ANDN U4146 ( .B(n2488), .A(n2489), .Z(n2487) );
XOR U4147 ( .A(c829), .B(b[829]), .Z(n2488) );
XNOR U4148 ( .A(b[829]), .B(n2489), .Z(c[829]) );
XNOR U4149 ( .A(a[829]), .B(c829), .Z(n2489) );
XOR U4150 ( .A(c830), .B(n2490), .Z(c831) );
ANDN U4151 ( .B(n2491), .A(n2492), .Z(n2490) );
XOR U4152 ( .A(c830), .B(b[830]), .Z(n2491) );
XNOR U4153 ( .A(b[830]), .B(n2492), .Z(c[830]) );
XNOR U4154 ( .A(a[830]), .B(c830), .Z(n2492) );
XOR U4155 ( .A(c831), .B(n2493), .Z(c832) );
ANDN U4156 ( .B(n2494), .A(n2495), .Z(n2493) );
XOR U4157 ( .A(c831), .B(b[831]), .Z(n2494) );
XNOR U4158 ( .A(b[831]), .B(n2495), .Z(c[831]) );
XNOR U4159 ( .A(a[831]), .B(c831), .Z(n2495) );
XOR U4160 ( .A(c832), .B(n2496), .Z(c833) );
ANDN U4161 ( .B(n2497), .A(n2498), .Z(n2496) );
XOR U4162 ( .A(c832), .B(b[832]), .Z(n2497) );
XNOR U4163 ( .A(b[832]), .B(n2498), .Z(c[832]) );
XNOR U4164 ( .A(a[832]), .B(c832), .Z(n2498) );
XOR U4165 ( .A(c833), .B(n2499), .Z(c834) );
ANDN U4166 ( .B(n2500), .A(n2501), .Z(n2499) );
XOR U4167 ( .A(c833), .B(b[833]), .Z(n2500) );
XNOR U4168 ( .A(b[833]), .B(n2501), .Z(c[833]) );
XNOR U4169 ( .A(a[833]), .B(c833), .Z(n2501) );
XOR U4170 ( .A(c834), .B(n2502), .Z(c835) );
ANDN U4171 ( .B(n2503), .A(n2504), .Z(n2502) );
XOR U4172 ( .A(c834), .B(b[834]), .Z(n2503) );
XNOR U4173 ( .A(b[834]), .B(n2504), .Z(c[834]) );
XNOR U4174 ( .A(a[834]), .B(c834), .Z(n2504) );
XOR U4175 ( .A(c835), .B(n2505), .Z(c836) );
ANDN U4176 ( .B(n2506), .A(n2507), .Z(n2505) );
XOR U4177 ( .A(c835), .B(b[835]), .Z(n2506) );
XNOR U4178 ( .A(b[835]), .B(n2507), .Z(c[835]) );
XNOR U4179 ( .A(a[835]), .B(c835), .Z(n2507) );
XOR U4180 ( .A(c836), .B(n2508), .Z(c837) );
ANDN U4181 ( .B(n2509), .A(n2510), .Z(n2508) );
XOR U4182 ( .A(c836), .B(b[836]), .Z(n2509) );
XNOR U4183 ( .A(b[836]), .B(n2510), .Z(c[836]) );
XNOR U4184 ( .A(a[836]), .B(c836), .Z(n2510) );
XOR U4185 ( .A(c837), .B(n2511), .Z(c838) );
ANDN U4186 ( .B(n2512), .A(n2513), .Z(n2511) );
XOR U4187 ( .A(c837), .B(b[837]), .Z(n2512) );
XNOR U4188 ( .A(b[837]), .B(n2513), .Z(c[837]) );
XNOR U4189 ( .A(a[837]), .B(c837), .Z(n2513) );
XOR U4190 ( .A(c838), .B(n2514), .Z(c839) );
ANDN U4191 ( .B(n2515), .A(n2516), .Z(n2514) );
XOR U4192 ( .A(c838), .B(b[838]), .Z(n2515) );
XNOR U4193 ( .A(b[838]), .B(n2516), .Z(c[838]) );
XNOR U4194 ( .A(a[838]), .B(c838), .Z(n2516) );
XOR U4195 ( .A(c839), .B(n2517), .Z(c840) );
ANDN U4196 ( .B(n2518), .A(n2519), .Z(n2517) );
XOR U4197 ( .A(c839), .B(b[839]), .Z(n2518) );
XNOR U4198 ( .A(b[839]), .B(n2519), .Z(c[839]) );
XNOR U4199 ( .A(a[839]), .B(c839), .Z(n2519) );
XOR U4200 ( .A(c840), .B(n2520), .Z(c841) );
ANDN U4201 ( .B(n2521), .A(n2522), .Z(n2520) );
XOR U4202 ( .A(c840), .B(b[840]), .Z(n2521) );
XNOR U4203 ( .A(b[840]), .B(n2522), .Z(c[840]) );
XNOR U4204 ( .A(a[840]), .B(c840), .Z(n2522) );
XOR U4205 ( .A(c841), .B(n2523), .Z(c842) );
ANDN U4206 ( .B(n2524), .A(n2525), .Z(n2523) );
XOR U4207 ( .A(c841), .B(b[841]), .Z(n2524) );
XNOR U4208 ( .A(b[841]), .B(n2525), .Z(c[841]) );
XNOR U4209 ( .A(a[841]), .B(c841), .Z(n2525) );
XOR U4210 ( .A(c842), .B(n2526), .Z(c843) );
ANDN U4211 ( .B(n2527), .A(n2528), .Z(n2526) );
XOR U4212 ( .A(c842), .B(b[842]), .Z(n2527) );
XNOR U4213 ( .A(b[842]), .B(n2528), .Z(c[842]) );
XNOR U4214 ( .A(a[842]), .B(c842), .Z(n2528) );
XOR U4215 ( .A(c843), .B(n2529), .Z(c844) );
ANDN U4216 ( .B(n2530), .A(n2531), .Z(n2529) );
XOR U4217 ( .A(c843), .B(b[843]), .Z(n2530) );
XNOR U4218 ( .A(b[843]), .B(n2531), .Z(c[843]) );
XNOR U4219 ( .A(a[843]), .B(c843), .Z(n2531) );
XOR U4220 ( .A(c844), .B(n2532), .Z(c845) );
ANDN U4221 ( .B(n2533), .A(n2534), .Z(n2532) );
XOR U4222 ( .A(c844), .B(b[844]), .Z(n2533) );
XNOR U4223 ( .A(b[844]), .B(n2534), .Z(c[844]) );
XNOR U4224 ( .A(a[844]), .B(c844), .Z(n2534) );
XOR U4225 ( .A(c845), .B(n2535), .Z(c846) );
ANDN U4226 ( .B(n2536), .A(n2537), .Z(n2535) );
XOR U4227 ( .A(c845), .B(b[845]), .Z(n2536) );
XNOR U4228 ( .A(b[845]), .B(n2537), .Z(c[845]) );
XNOR U4229 ( .A(a[845]), .B(c845), .Z(n2537) );
XOR U4230 ( .A(c846), .B(n2538), .Z(c847) );
ANDN U4231 ( .B(n2539), .A(n2540), .Z(n2538) );
XOR U4232 ( .A(c846), .B(b[846]), .Z(n2539) );
XNOR U4233 ( .A(b[846]), .B(n2540), .Z(c[846]) );
XNOR U4234 ( .A(a[846]), .B(c846), .Z(n2540) );
XOR U4235 ( .A(c847), .B(n2541), .Z(c848) );
ANDN U4236 ( .B(n2542), .A(n2543), .Z(n2541) );
XOR U4237 ( .A(c847), .B(b[847]), .Z(n2542) );
XNOR U4238 ( .A(b[847]), .B(n2543), .Z(c[847]) );
XNOR U4239 ( .A(a[847]), .B(c847), .Z(n2543) );
XOR U4240 ( .A(c848), .B(n2544), .Z(c849) );
ANDN U4241 ( .B(n2545), .A(n2546), .Z(n2544) );
XOR U4242 ( .A(c848), .B(b[848]), .Z(n2545) );
XNOR U4243 ( .A(b[848]), .B(n2546), .Z(c[848]) );
XNOR U4244 ( .A(a[848]), .B(c848), .Z(n2546) );
XOR U4245 ( .A(c849), .B(n2547), .Z(c850) );
ANDN U4246 ( .B(n2548), .A(n2549), .Z(n2547) );
XOR U4247 ( .A(c849), .B(b[849]), .Z(n2548) );
XNOR U4248 ( .A(b[849]), .B(n2549), .Z(c[849]) );
XNOR U4249 ( .A(a[849]), .B(c849), .Z(n2549) );
XOR U4250 ( .A(c850), .B(n2550), .Z(c851) );
ANDN U4251 ( .B(n2551), .A(n2552), .Z(n2550) );
XOR U4252 ( .A(c850), .B(b[850]), .Z(n2551) );
XNOR U4253 ( .A(b[850]), .B(n2552), .Z(c[850]) );
XNOR U4254 ( .A(a[850]), .B(c850), .Z(n2552) );
XOR U4255 ( .A(c851), .B(n2553), .Z(c852) );
ANDN U4256 ( .B(n2554), .A(n2555), .Z(n2553) );
XOR U4257 ( .A(c851), .B(b[851]), .Z(n2554) );
XNOR U4258 ( .A(b[851]), .B(n2555), .Z(c[851]) );
XNOR U4259 ( .A(a[851]), .B(c851), .Z(n2555) );
XOR U4260 ( .A(c852), .B(n2556), .Z(c853) );
ANDN U4261 ( .B(n2557), .A(n2558), .Z(n2556) );
XOR U4262 ( .A(c852), .B(b[852]), .Z(n2557) );
XNOR U4263 ( .A(b[852]), .B(n2558), .Z(c[852]) );
XNOR U4264 ( .A(a[852]), .B(c852), .Z(n2558) );
XOR U4265 ( .A(c853), .B(n2559), .Z(c854) );
ANDN U4266 ( .B(n2560), .A(n2561), .Z(n2559) );
XOR U4267 ( .A(c853), .B(b[853]), .Z(n2560) );
XNOR U4268 ( .A(b[853]), .B(n2561), .Z(c[853]) );
XNOR U4269 ( .A(a[853]), .B(c853), .Z(n2561) );
XOR U4270 ( .A(c854), .B(n2562), .Z(c855) );
ANDN U4271 ( .B(n2563), .A(n2564), .Z(n2562) );
XOR U4272 ( .A(c854), .B(b[854]), .Z(n2563) );
XNOR U4273 ( .A(b[854]), .B(n2564), .Z(c[854]) );
XNOR U4274 ( .A(a[854]), .B(c854), .Z(n2564) );
XOR U4275 ( .A(c855), .B(n2565), .Z(c856) );
ANDN U4276 ( .B(n2566), .A(n2567), .Z(n2565) );
XOR U4277 ( .A(c855), .B(b[855]), .Z(n2566) );
XNOR U4278 ( .A(b[855]), .B(n2567), .Z(c[855]) );
XNOR U4279 ( .A(a[855]), .B(c855), .Z(n2567) );
XOR U4280 ( .A(c856), .B(n2568), .Z(c857) );
ANDN U4281 ( .B(n2569), .A(n2570), .Z(n2568) );
XOR U4282 ( .A(c856), .B(b[856]), .Z(n2569) );
XNOR U4283 ( .A(b[856]), .B(n2570), .Z(c[856]) );
XNOR U4284 ( .A(a[856]), .B(c856), .Z(n2570) );
XOR U4285 ( .A(c857), .B(n2571), .Z(c858) );
ANDN U4286 ( .B(n2572), .A(n2573), .Z(n2571) );
XOR U4287 ( .A(c857), .B(b[857]), .Z(n2572) );
XNOR U4288 ( .A(b[857]), .B(n2573), .Z(c[857]) );
XNOR U4289 ( .A(a[857]), .B(c857), .Z(n2573) );
XOR U4290 ( .A(c858), .B(n2574), .Z(c859) );
ANDN U4291 ( .B(n2575), .A(n2576), .Z(n2574) );
XOR U4292 ( .A(c858), .B(b[858]), .Z(n2575) );
XNOR U4293 ( .A(b[858]), .B(n2576), .Z(c[858]) );
XNOR U4294 ( .A(a[858]), .B(c858), .Z(n2576) );
XOR U4295 ( .A(c859), .B(n2577), .Z(c860) );
ANDN U4296 ( .B(n2578), .A(n2579), .Z(n2577) );
XOR U4297 ( .A(c859), .B(b[859]), .Z(n2578) );
XNOR U4298 ( .A(b[859]), .B(n2579), .Z(c[859]) );
XNOR U4299 ( .A(a[859]), .B(c859), .Z(n2579) );
XOR U4300 ( .A(c860), .B(n2580), .Z(c861) );
ANDN U4301 ( .B(n2581), .A(n2582), .Z(n2580) );
XOR U4302 ( .A(c860), .B(b[860]), .Z(n2581) );
XNOR U4303 ( .A(b[860]), .B(n2582), .Z(c[860]) );
XNOR U4304 ( .A(a[860]), .B(c860), .Z(n2582) );
XOR U4305 ( .A(c861), .B(n2583), .Z(c862) );
ANDN U4306 ( .B(n2584), .A(n2585), .Z(n2583) );
XOR U4307 ( .A(c861), .B(b[861]), .Z(n2584) );
XNOR U4308 ( .A(b[861]), .B(n2585), .Z(c[861]) );
XNOR U4309 ( .A(a[861]), .B(c861), .Z(n2585) );
XOR U4310 ( .A(c862), .B(n2586), .Z(c863) );
ANDN U4311 ( .B(n2587), .A(n2588), .Z(n2586) );
XOR U4312 ( .A(c862), .B(b[862]), .Z(n2587) );
XNOR U4313 ( .A(b[862]), .B(n2588), .Z(c[862]) );
XNOR U4314 ( .A(a[862]), .B(c862), .Z(n2588) );
XOR U4315 ( .A(c863), .B(n2589), .Z(c864) );
ANDN U4316 ( .B(n2590), .A(n2591), .Z(n2589) );
XOR U4317 ( .A(c863), .B(b[863]), .Z(n2590) );
XNOR U4318 ( .A(b[863]), .B(n2591), .Z(c[863]) );
XNOR U4319 ( .A(a[863]), .B(c863), .Z(n2591) );
XOR U4320 ( .A(c864), .B(n2592), .Z(c865) );
ANDN U4321 ( .B(n2593), .A(n2594), .Z(n2592) );
XOR U4322 ( .A(c864), .B(b[864]), .Z(n2593) );
XNOR U4323 ( .A(b[864]), .B(n2594), .Z(c[864]) );
XNOR U4324 ( .A(a[864]), .B(c864), .Z(n2594) );
XOR U4325 ( .A(c865), .B(n2595), .Z(c866) );
ANDN U4326 ( .B(n2596), .A(n2597), .Z(n2595) );
XOR U4327 ( .A(c865), .B(b[865]), .Z(n2596) );
XNOR U4328 ( .A(b[865]), .B(n2597), .Z(c[865]) );
XNOR U4329 ( .A(a[865]), .B(c865), .Z(n2597) );
XOR U4330 ( .A(c866), .B(n2598), .Z(c867) );
ANDN U4331 ( .B(n2599), .A(n2600), .Z(n2598) );
XOR U4332 ( .A(c866), .B(b[866]), .Z(n2599) );
XNOR U4333 ( .A(b[866]), .B(n2600), .Z(c[866]) );
XNOR U4334 ( .A(a[866]), .B(c866), .Z(n2600) );
XOR U4335 ( .A(c867), .B(n2601), .Z(c868) );
ANDN U4336 ( .B(n2602), .A(n2603), .Z(n2601) );
XOR U4337 ( .A(c867), .B(b[867]), .Z(n2602) );
XNOR U4338 ( .A(b[867]), .B(n2603), .Z(c[867]) );
XNOR U4339 ( .A(a[867]), .B(c867), .Z(n2603) );
XOR U4340 ( .A(c868), .B(n2604), .Z(c869) );
ANDN U4341 ( .B(n2605), .A(n2606), .Z(n2604) );
XOR U4342 ( .A(c868), .B(b[868]), .Z(n2605) );
XNOR U4343 ( .A(b[868]), .B(n2606), .Z(c[868]) );
XNOR U4344 ( .A(a[868]), .B(c868), .Z(n2606) );
XOR U4345 ( .A(c869), .B(n2607), .Z(c870) );
ANDN U4346 ( .B(n2608), .A(n2609), .Z(n2607) );
XOR U4347 ( .A(c869), .B(b[869]), .Z(n2608) );
XNOR U4348 ( .A(b[869]), .B(n2609), .Z(c[869]) );
XNOR U4349 ( .A(a[869]), .B(c869), .Z(n2609) );
XOR U4350 ( .A(c870), .B(n2610), .Z(c871) );
ANDN U4351 ( .B(n2611), .A(n2612), .Z(n2610) );
XOR U4352 ( .A(c870), .B(b[870]), .Z(n2611) );
XNOR U4353 ( .A(b[870]), .B(n2612), .Z(c[870]) );
XNOR U4354 ( .A(a[870]), .B(c870), .Z(n2612) );
XOR U4355 ( .A(c871), .B(n2613), .Z(c872) );
ANDN U4356 ( .B(n2614), .A(n2615), .Z(n2613) );
XOR U4357 ( .A(c871), .B(b[871]), .Z(n2614) );
XNOR U4358 ( .A(b[871]), .B(n2615), .Z(c[871]) );
XNOR U4359 ( .A(a[871]), .B(c871), .Z(n2615) );
XOR U4360 ( .A(c872), .B(n2616), .Z(c873) );
ANDN U4361 ( .B(n2617), .A(n2618), .Z(n2616) );
XOR U4362 ( .A(c872), .B(b[872]), .Z(n2617) );
XNOR U4363 ( .A(b[872]), .B(n2618), .Z(c[872]) );
XNOR U4364 ( .A(a[872]), .B(c872), .Z(n2618) );
XOR U4365 ( .A(c873), .B(n2619), .Z(c874) );
ANDN U4366 ( .B(n2620), .A(n2621), .Z(n2619) );
XOR U4367 ( .A(c873), .B(b[873]), .Z(n2620) );
XNOR U4368 ( .A(b[873]), .B(n2621), .Z(c[873]) );
XNOR U4369 ( .A(a[873]), .B(c873), .Z(n2621) );
XOR U4370 ( .A(c874), .B(n2622), .Z(c875) );
ANDN U4371 ( .B(n2623), .A(n2624), .Z(n2622) );
XOR U4372 ( .A(c874), .B(b[874]), .Z(n2623) );
XNOR U4373 ( .A(b[874]), .B(n2624), .Z(c[874]) );
XNOR U4374 ( .A(a[874]), .B(c874), .Z(n2624) );
XOR U4375 ( .A(c875), .B(n2625), .Z(c876) );
ANDN U4376 ( .B(n2626), .A(n2627), .Z(n2625) );
XOR U4377 ( .A(c875), .B(b[875]), .Z(n2626) );
XNOR U4378 ( .A(b[875]), .B(n2627), .Z(c[875]) );
XNOR U4379 ( .A(a[875]), .B(c875), .Z(n2627) );
XOR U4380 ( .A(c876), .B(n2628), .Z(c877) );
ANDN U4381 ( .B(n2629), .A(n2630), .Z(n2628) );
XOR U4382 ( .A(c876), .B(b[876]), .Z(n2629) );
XNOR U4383 ( .A(b[876]), .B(n2630), .Z(c[876]) );
XNOR U4384 ( .A(a[876]), .B(c876), .Z(n2630) );
XOR U4385 ( .A(c877), .B(n2631), .Z(c878) );
ANDN U4386 ( .B(n2632), .A(n2633), .Z(n2631) );
XOR U4387 ( .A(c877), .B(b[877]), .Z(n2632) );
XNOR U4388 ( .A(b[877]), .B(n2633), .Z(c[877]) );
XNOR U4389 ( .A(a[877]), .B(c877), .Z(n2633) );
XOR U4390 ( .A(c878), .B(n2634), .Z(c879) );
ANDN U4391 ( .B(n2635), .A(n2636), .Z(n2634) );
XOR U4392 ( .A(c878), .B(b[878]), .Z(n2635) );
XNOR U4393 ( .A(b[878]), .B(n2636), .Z(c[878]) );
XNOR U4394 ( .A(a[878]), .B(c878), .Z(n2636) );
XOR U4395 ( .A(c879), .B(n2637), .Z(c880) );
ANDN U4396 ( .B(n2638), .A(n2639), .Z(n2637) );
XOR U4397 ( .A(c879), .B(b[879]), .Z(n2638) );
XNOR U4398 ( .A(b[879]), .B(n2639), .Z(c[879]) );
XNOR U4399 ( .A(a[879]), .B(c879), .Z(n2639) );
XOR U4400 ( .A(c880), .B(n2640), .Z(c881) );
ANDN U4401 ( .B(n2641), .A(n2642), .Z(n2640) );
XOR U4402 ( .A(c880), .B(b[880]), .Z(n2641) );
XNOR U4403 ( .A(b[880]), .B(n2642), .Z(c[880]) );
XNOR U4404 ( .A(a[880]), .B(c880), .Z(n2642) );
XOR U4405 ( .A(c881), .B(n2643), .Z(c882) );
ANDN U4406 ( .B(n2644), .A(n2645), .Z(n2643) );
XOR U4407 ( .A(c881), .B(b[881]), .Z(n2644) );
XNOR U4408 ( .A(b[881]), .B(n2645), .Z(c[881]) );
XNOR U4409 ( .A(a[881]), .B(c881), .Z(n2645) );
XOR U4410 ( .A(c882), .B(n2646), .Z(c883) );
ANDN U4411 ( .B(n2647), .A(n2648), .Z(n2646) );
XOR U4412 ( .A(c882), .B(b[882]), .Z(n2647) );
XNOR U4413 ( .A(b[882]), .B(n2648), .Z(c[882]) );
XNOR U4414 ( .A(a[882]), .B(c882), .Z(n2648) );
XOR U4415 ( .A(c883), .B(n2649), .Z(c884) );
ANDN U4416 ( .B(n2650), .A(n2651), .Z(n2649) );
XOR U4417 ( .A(c883), .B(b[883]), .Z(n2650) );
XNOR U4418 ( .A(b[883]), .B(n2651), .Z(c[883]) );
XNOR U4419 ( .A(a[883]), .B(c883), .Z(n2651) );
XOR U4420 ( .A(c884), .B(n2652), .Z(c885) );
ANDN U4421 ( .B(n2653), .A(n2654), .Z(n2652) );
XOR U4422 ( .A(c884), .B(b[884]), .Z(n2653) );
XNOR U4423 ( .A(b[884]), .B(n2654), .Z(c[884]) );
XNOR U4424 ( .A(a[884]), .B(c884), .Z(n2654) );
XOR U4425 ( .A(c885), .B(n2655), .Z(c886) );
ANDN U4426 ( .B(n2656), .A(n2657), .Z(n2655) );
XOR U4427 ( .A(c885), .B(b[885]), .Z(n2656) );
XNOR U4428 ( .A(b[885]), .B(n2657), .Z(c[885]) );
XNOR U4429 ( .A(a[885]), .B(c885), .Z(n2657) );
XOR U4430 ( .A(c886), .B(n2658), .Z(c887) );
ANDN U4431 ( .B(n2659), .A(n2660), .Z(n2658) );
XOR U4432 ( .A(c886), .B(b[886]), .Z(n2659) );
XNOR U4433 ( .A(b[886]), .B(n2660), .Z(c[886]) );
XNOR U4434 ( .A(a[886]), .B(c886), .Z(n2660) );
XOR U4435 ( .A(c887), .B(n2661), .Z(c888) );
ANDN U4436 ( .B(n2662), .A(n2663), .Z(n2661) );
XOR U4437 ( .A(c887), .B(b[887]), .Z(n2662) );
XNOR U4438 ( .A(b[887]), .B(n2663), .Z(c[887]) );
XNOR U4439 ( .A(a[887]), .B(c887), .Z(n2663) );
XOR U4440 ( .A(c888), .B(n2664), .Z(c889) );
ANDN U4441 ( .B(n2665), .A(n2666), .Z(n2664) );
XOR U4442 ( .A(c888), .B(b[888]), .Z(n2665) );
XNOR U4443 ( .A(b[888]), .B(n2666), .Z(c[888]) );
XNOR U4444 ( .A(a[888]), .B(c888), .Z(n2666) );
XOR U4445 ( .A(c889), .B(n2667), .Z(c890) );
ANDN U4446 ( .B(n2668), .A(n2669), .Z(n2667) );
XOR U4447 ( .A(c889), .B(b[889]), .Z(n2668) );
XNOR U4448 ( .A(b[889]), .B(n2669), .Z(c[889]) );
XNOR U4449 ( .A(a[889]), .B(c889), .Z(n2669) );
XOR U4450 ( .A(c890), .B(n2670), .Z(c891) );
ANDN U4451 ( .B(n2671), .A(n2672), .Z(n2670) );
XOR U4452 ( .A(c890), .B(b[890]), .Z(n2671) );
XNOR U4453 ( .A(b[890]), .B(n2672), .Z(c[890]) );
XNOR U4454 ( .A(a[890]), .B(c890), .Z(n2672) );
XOR U4455 ( .A(c891), .B(n2673), .Z(c892) );
ANDN U4456 ( .B(n2674), .A(n2675), .Z(n2673) );
XOR U4457 ( .A(c891), .B(b[891]), .Z(n2674) );
XNOR U4458 ( .A(b[891]), .B(n2675), .Z(c[891]) );
XNOR U4459 ( .A(a[891]), .B(c891), .Z(n2675) );
XOR U4460 ( .A(c892), .B(n2676), .Z(c893) );
ANDN U4461 ( .B(n2677), .A(n2678), .Z(n2676) );
XOR U4462 ( .A(c892), .B(b[892]), .Z(n2677) );
XNOR U4463 ( .A(b[892]), .B(n2678), .Z(c[892]) );
XNOR U4464 ( .A(a[892]), .B(c892), .Z(n2678) );
XOR U4465 ( .A(c893), .B(n2679), .Z(c894) );
ANDN U4466 ( .B(n2680), .A(n2681), .Z(n2679) );
XOR U4467 ( .A(c893), .B(b[893]), .Z(n2680) );
XNOR U4468 ( .A(b[893]), .B(n2681), .Z(c[893]) );
XNOR U4469 ( .A(a[893]), .B(c893), .Z(n2681) );
XOR U4470 ( .A(c894), .B(n2682), .Z(c895) );
ANDN U4471 ( .B(n2683), .A(n2684), .Z(n2682) );
XOR U4472 ( .A(c894), .B(b[894]), .Z(n2683) );
XNOR U4473 ( .A(b[894]), .B(n2684), .Z(c[894]) );
XNOR U4474 ( .A(a[894]), .B(c894), .Z(n2684) );
XOR U4475 ( .A(c895), .B(n2685), .Z(c896) );
ANDN U4476 ( .B(n2686), .A(n2687), .Z(n2685) );
XOR U4477 ( .A(c895), .B(b[895]), .Z(n2686) );
XNOR U4478 ( .A(b[895]), .B(n2687), .Z(c[895]) );
XNOR U4479 ( .A(a[895]), .B(c895), .Z(n2687) );
XOR U4480 ( .A(c896), .B(n2688), .Z(c897) );
ANDN U4481 ( .B(n2689), .A(n2690), .Z(n2688) );
XOR U4482 ( .A(c896), .B(b[896]), .Z(n2689) );
XNOR U4483 ( .A(b[896]), .B(n2690), .Z(c[896]) );
XNOR U4484 ( .A(a[896]), .B(c896), .Z(n2690) );
XOR U4485 ( .A(c897), .B(n2691), .Z(c898) );
ANDN U4486 ( .B(n2692), .A(n2693), .Z(n2691) );
XOR U4487 ( .A(c897), .B(b[897]), .Z(n2692) );
XNOR U4488 ( .A(b[897]), .B(n2693), .Z(c[897]) );
XNOR U4489 ( .A(a[897]), .B(c897), .Z(n2693) );
XOR U4490 ( .A(c898), .B(n2694), .Z(c899) );
ANDN U4491 ( .B(n2695), .A(n2696), .Z(n2694) );
XOR U4492 ( .A(c898), .B(b[898]), .Z(n2695) );
XNOR U4493 ( .A(b[898]), .B(n2696), .Z(c[898]) );
XNOR U4494 ( .A(a[898]), .B(c898), .Z(n2696) );
XOR U4495 ( .A(c899), .B(n2697), .Z(c900) );
ANDN U4496 ( .B(n2698), .A(n2699), .Z(n2697) );
XOR U4497 ( .A(c899), .B(b[899]), .Z(n2698) );
XNOR U4498 ( .A(b[899]), .B(n2699), .Z(c[899]) );
XNOR U4499 ( .A(a[899]), .B(c899), .Z(n2699) );
XOR U4500 ( .A(c900), .B(n2700), .Z(c901) );
ANDN U4501 ( .B(n2701), .A(n2702), .Z(n2700) );
XOR U4502 ( .A(c900), .B(b[900]), .Z(n2701) );
XNOR U4503 ( .A(b[900]), .B(n2702), .Z(c[900]) );
XNOR U4504 ( .A(a[900]), .B(c900), .Z(n2702) );
XOR U4505 ( .A(c901), .B(n2703), .Z(c902) );
ANDN U4506 ( .B(n2704), .A(n2705), .Z(n2703) );
XOR U4507 ( .A(c901), .B(b[901]), .Z(n2704) );
XNOR U4508 ( .A(b[901]), .B(n2705), .Z(c[901]) );
XNOR U4509 ( .A(a[901]), .B(c901), .Z(n2705) );
XOR U4510 ( .A(c902), .B(n2706), .Z(c903) );
ANDN U4511 ( .B(n2707), .A(n2708), .Z(n2706) );
XOR U4512 ( .A(c902), .B(b[902]), .Z(n2707) );
XNOR U4513 ( .A(b[902]), .B(n2708), .Z(c[902]) );
XNOR U4514 ( .A(a[902]), .B(c902), .Z(n2708) );
XOR U4515 ( .A(c903), .B(n2709), .Z(c904) );
ANDN U4516 ( .B(n2710), .A(n2711), .Z(n2709) );
XOR U4517 ( .A(c903), .B(b[903]), .Z(n2710) );
XNOR U4518 ( .A(b[903]), .B(n2711), .Z(c[903]) );
XNOR U4519 ( .A(a[903]), .B(c903), .Z(n2711) );
XOR U4520 ( .A(c904), .B(n2712), .Z(c905) );
ANDN U4521 ( .B(n2713), .A(n2714), .Z(n2712) );
XOR U4522 ( .A(c904), .B(b[904]), .Z(n2713) );
XNOR U4523 ( .A(b[904]), .B(n2714), .Z(c[904]) );
XNOR U4524 ( .A(a[904]), .B(c904), .Z(n2714) );
XOR U4525 ( .A(c905), .B(n2715), .Z(c906) );
ANDN U4526 ( .B(n2716), .A(n2717), .Z(n2715) );
XOR U4527 ( .A(c905), .B(b[905]), .Z(n2716) );
XNOR U4528 ( .A(b[905]), .B(n2717), .Z(c[905]) );
XNOR U4529 ( .A(a[905]), .B(c905), .Z(n2717) );
XOR U4530 ( .A(c906), .B(n2718), .Z(c907) );
ANDN U4531 ( .B(n2719), .A(n2720), .Z(n2718) );
XOR U4532 ( .A(c906), .B(b[906]), .Z(n2719) );
XNOR U4533 ( .A(b[906]), .B(n2720), .Z(c[906]) );
XNOR U4534 ( .A(a[906]), .B(c906), .Z(n2720) );
XOR U4535 ( .A(c907), .B(n2721), .Z(c908) );
ANDN U4536 ( .B(n2722), .A(n2723), .Z(n2721) );
XOR U4537 ( .A(c907), .B(b[907]), .Z(n2722) );
XNOR U4538 ( .A(b[907]), .B(n2723), .Z(c[907]) );
XNOR U4539 ( .A(a[907]), .B(c907), .Z(n2723) );
XOR U4540 ( .A(c908), .B(n2724), .Z(c909) );
ANDN U4541 ( .B(n2725), .A(n2726), .Z(n2724) );
XOR U4542 ( .A(c908), .B(b[908]), .Z(n2725) );
XNOR U4543 ( .A(b[908]), .B(n2726), .Z(c[908]) );
XNOR U4544 ( .A(a[908]), .B(c908), .Z(n2726) );
XOR U4545 ( .A(c909), .B(n2727), .Z(c910) );
ANDN U4546 ( .B(n2728), .A(n2729), .Z(n2727) );
XOR U4547 ( .A(c909), .B(b[909]), .Z(n2728) );
XNOR U4548 ( .A(b[909]), .B(n2729), .Z(c[909]) );
XNOR U4549 ( .A(a[909]), .B(c909), .Z(n2729) );
XOR U4550 ( .A(c910), .B(n2730), .Z(c911) );
ANDN U4551 ( .B(n2731), .A(n2732), .Z(n2730) );
XOR U4552 ( .A(c910), .B(b[910]), .Z(n2731) );
XNOR U4553 ( .A(b[910]), .B(n2732), .Z(c[910]) );
XNOR U4554 ( .A(a[910]), .B(c910), .Z(n2732) );
XOR U4555 ( .A(c911), .B(n2733), .Z(c912) );
ANDN U4556 ( .B(n2734), .A(n2735), .Z(n2733) );
XOR U4557 ( .A(c911), .B(b[911]), .Z(n2734) );
XNOR U4558 ( .A(b[911]), .B(n2735), .Z(c[911]) );
XNOR U4559 ( .A(a[911]), .B(c911), .Z(n2735) );
XOR U4560 ( .A(c912), .B(n2736), .Z(c913) );
ANDN U4561 ( .B(n2737), .A(n2738), .Z(n2736) );
XOR U4562 ( .A(c912), .B(b[912]), .Z(n2737) );
XNOR U4563 ( .A(b[912]), .B(n2738), .Z(c[912]) );
XNOR U4564 ( .A(a[912]), .B(c912), .Z(n2738) );
XOR U4565 ( .A(c913), .B(n2739), .Z(c914) );
ANDN U4566 ( .B(n2740), .A(n2741), .Z(n2739) );
XOR U4567 ( .A(c913), .B(b[913]), .Z(n2740) );
XNOR U4568 ( .A(b[913]), .B(n2741), .Z(c[913]) );
XNOR U4569 ( .A(a[913]), .B(c913), .Z(n2741) );
XOR U4570 ( .A(c914), .B(n2742), .Z(c915) );
ANDN U4571 ( .B(n2743), .A(n2744), .Z(n2742) );
XOR U4572 ( .A(c914), .B(b[914]), .Z(n2743) );
XNOR U4573 ( .A(b[914]), .B(n2744), .Z(c[914]) );
XNOR U4574 ( .A(a[914]), .B(c914), .Z(n2744) );
XOR U4575 ( .A(c915), .B(n2745), .Z(c916) );
ANDN U4576 ( .B(n2746), .A(n2747), .Z(n2745) );
XOR U4577 ( .A(c915), .B(b[915]), .Z(n2746) );
XNOR U4578 ( .A(b[915]), .B(n2747), .Z(c[915]) );
XNOR U4579 ( .A(a[915]), .B(c915), .Z(n2747) );
XOR U4580 ( .A(c916), .B(n2748), .Z(c917) );
ANDN U4581 ( .B(n2749), .A(n2750), .Z(n2748) );
XOR U4582 ( .A(c916), .B(b[916]), .Z(n2749) );
XNOR U4583 ( .A(b[916]), .B(n2750), .Z(c[916]) );
XNOR U4584 ( .A(a[916]), .B(c916), .Z(n2750) );
XOR U4585 ( .A(c917), .B(n2751), .Z(c918) );
ANDN U4586 ( .B(n2752), .A(n2753), .Z(n2751) );
XOR U4587 ( .A(c917), .B(b[917]), .Z(n2752) );
XNOR U4588 ( .A(b[917]), .B(n2753), .Z(c[917]) );
XNOR U4589 ( .A(a[917]), .B(c917), .Z(n2753) );
XOR U4590 ( .A(c918), .B(n2754), .Z(c919) );
ANDN U4591 ( .B(n2755), .A(n2756), .Z(n2754) );
XOR U4592 ( .A(c918), .B(b[918]), .Z(n2755) );
XNOR U4593 ( .A(b[918]), .B(n2756), .Z(c[918]) );
XNOR U4594 ( .A(a[918]), .B(c918), .Z(n2756) );
XOR U4595 ( .A(c919), .B(n2757), .Z(c920) );
ANDN U4596 ( .B(n2758), .A(n2759), .Z(n2757) );
XOR U4597 ( .A(c919), .B(b[919]), .Z(n2758) );
XNOR U4598 ( .A(b[919]), .B(n2759), .Z(c[919]) );
XNOR U4599 ( .A(a[919]), .B(c919), .Z(n2759) );
XOR U4600 ( .A(c920), .B(n2760), .Z(c921) );
ANDN U4601 ( .B(n2761), .A(n2762), .Z(n2760) );
XOR U4602 ( .A(c920), .B(b[920]), .Z(n2761) );
XNOR U4603 ( .A(b[920]), .B(n2762), .Z(c[920]) );
XNOR U4604 ( .A(a[920]), .B(c920), .Z(n2762) );
XOR U4605 ( .A(c921), .B(n2763), .Z(c922) );
ANDN U4606 ( .B(n2764), .A(n2765), .Z(n2763) );
XOR U4607 ( .A(c921), .B(b[921]), .Z(n2764) );
XNOR U4608 ( .A(b[921]), .B(n2765), .Z(c[921]) );
XNOR U4609 ( .A(a[921]), .B(c921), .Z(n2765) );
XOR U4610 ( .A(c922), .B(n2766), .Z(c923) );
ANDN U4611 ( .B(n2767), .A(n2768), .Z(n2766) );
XOR U4612 ( .A(c922), .B(b[922]), .Z(n2767) );
XNOR U4613 ( .A(b[922]), .B(n2768), .Z(c[922]) );
XNOR U4614 ( .A(a[922]), .B(c922), .Z(n2768) );
XOR U4615 ( .A(c923), .B(n2769), .Z(c924) );
ANDN U4616 ( .B(n2770), .A(n2771), .Z(n2769) );
XOR U4617 ( .A(c923), .B(b[923]), .Z(n2770) );
XNOR U4618 ( .A(b[923]), .B(n2771), .Z(c[923]) );
XNOR U4619 ( .A(a[923]), .B(c923), .Z(n2771) );
XOR U4620 ( .A(c924), .B(n2772), .Z(c925) );
ANDN U4621 ( .B(n2773), .A(n2774), .Z(n2772) );
XOR U4622 ( .A(c924), .B(b[924]), .Z(n2773) );
XNOR U4623 ( .A(b[924]), .B(n2774), .Z(c[924]) );
XNOR U4624 ( .A(a[924]), .B(c924), .Z(n2774) );
XOR U4625 ( .A(c925), .B(n2775), .Z(c926) );
ANDN U4626 ( .B(n2776), .A(n2777), .Z(n2775) );
XOR U4627 ( .A(c925), .B(b[925]), .Z(n2776) );
XNOR U4628 ( .A(b[925]), .B(n2777), .Z(c[925]) );
XNOR U4629 ( .A(a[925]), .B(c925), .Z(n2777) );
XOR U4630 ( .A(c926), .B(n2778), .Z(c927) );
ANDN U4631 ( .B(n2779), .A(n2780), .Z(n2778) );
XOR U4632 ( .A(c926), .B(b[926]), .Z(n2779) );
XNOR U4633 ( .A(b[926]), .B(n2780), .Z(c[926]) );
XNOR U4634 ( .A(a[926]), .B(c926), .Z(n2780) );
XOR U4635 ( .A(c927), .B(n2781), .Z(c928) );
ANDN U4636 ( .B(n2782), .A(n2783), .Z(n2781) );
XOR U4637 ( .A(c927), .B(b[927]), .Z(n2782) );
XNOR U4638 ( .A(b[927]), .B(n2783), .Z(c[927]) );
XNOR U4639 ( .A(a[927]), .B(c927), .Z(n2783) );
XOR U4640 ( .A(c928), .B(n2784), .Z(c929) );
ANDN U4641 ( .B(n2785), .A(n2786), .Z(n2784) );
XOR U4642 ( .A(c928), .B(b[928]), .Z(n2785) );
XNOR U4643 ( .A(b[928]), .B(n2786), .Z(c[928]) );
XNOR U4644 ( .A(a[928]), .B(c928), .Z(n2786) );
XOR U4645 ( .A(c929), .B(n2787), .Z(c930) );
ANDN U4646 ( .B(n2788), .A(n2789), .Z(n2787) );
XOR U4647 ( .A(c929), .B(b[929]), .Z(n2788) );
XNOR U4648 ( .A(b[929]), .B(n2789), .Z(c[929]) );
XNOR U4649 ( .A(a[929]), .B(c929), .Z(n2789) );
XOR U4650 ( .A(c930), .B(n2790), .Z(c931) );
ANDN U4651 ( .B(n2791), .A(n2792), .Z(n2790) );
XOR U4652 ( .A(c930), .B(b[930]), .Z(n2791) );
XNOR U4653 ( .A(b[930]), .B(n2792), .Z(c[930]) );
XNOR U4654 ( .A(a[930]), .B(c930), .Z(n2792) );
XOR U4655 ( .A(c931), .B(n2793), .Z(c932) );
ANDN U4656 ( .B(n2794), .A(n2795), .Z(n2793) );
XOR U4657 ( .A(c931), .B(b[931]), .Z(n2794) );
XNOR U4658 ( .A(b[931]), .B(n2795), .Z(c[931]) );
XNOR U4659 ( .A(a[931]), .B(c931), .Z(n2795) );
XOR U4660 ( .A(c932), .B(n2796), .Z(c933) );
ANDN U4661 ( .B(n2797), .A(n2798), .Z(n2796) );
XOR U4662 ( .A(c932), .B(b[932]), .Z(n2797) );
XNOR U4663 ( .A(b[932]), .B(n2798), .Z(c[932]) );
XNOR U4664 ( .A(a[932]), .B(c932), .Z(n2798) );
XOR U4665 ( .A(c933), .B(n2799), .Z(c934) );
ANDN U4666 ( .B(n2800), .A(n2801), .Z(n2799) );
XOR U4667 ( .A(c933), .B(b[933]), .Z(n2800) );
XNOR U4668 ( .A(b[933]), .B(n2801), .Z(c[933]) );
XNOR U4669 ( .A(a[933]), .B(c933), .Z(n2801) );
XOR U4670 ( .A(c934), .B(n2802), .Z(c935) );
ANDN U4671 ( .B(n2803), .A(n2804), .Z(n2802) );
XOR U4672 ( .A(c934), .B(b[934]), .Z(n2803) );
XNOR U4673 ( .A(b[934]), .B(n2804), .Z(c[934]) );
XNOR U4674 ( .A(a[934]), .B(c934), .Z(n2804) );
XOR U4675 ( .A(c935), .B(n2805), .Z(c936) );
ANDN U4676 ( .B(n2806), .A(n2807), .Z(n2805) );
XOR U4677 ( .A(c935), .B(b[935]), .Z(n2806) );
XNOR U4678 ( .A(b[935]), .B(n2807), .Z(c[935]) );
XNOR U4679 ( .A(a[935]), .B(c935), .Z(n2807) );
XOR U4680 ( .A(c936), .B(n2808), .Z(c937) );
ANDN U4681 ( .B(n2809), .A(n2810), .Z(n2808) );
XOR U4682 ( .A(c936), .B(b[936]), .Z(n2809) );
XNOR U4683 ( .A(b[936]), .B(n2810), .Z(c[936]) );
XNOR U4684 ( .A(a[936]), .B(c936), .Z(n2810) );
XOR U4685 ( .A(c937), .B(n2811), .Z(c938) );
ANDN U4686 ( .B(n2812), .A(n2813), .Z(n2811) );
XOR U4687 ( .A(c937), .B(b[937]), .Z(n2812) );
XNOR U4688 ( .A(b[937]), .B(n2813), .Z(c[937]) );
XNOR U4689 ( .A(a[937]), .B(c937), .Z(n2813) );
XOR U4690 ( .A(c938), .B(n2814), .Z(c939) );
ANDN U4691 ( .B(n2815), .A(n2816), .Z(n2814) );
XOR U4692 ( .A(c938), .B(b[938]), .Z(n2815) );
XNOR U4693 ( .A(b[938]), .B(n2816), .Z(c[938]) );
XNOR U4694 ( .A(a[938]), .B(c938), .Z(n2816) );
XOR U4695 ( .A(c939), .B(n2817), .Z(c940) );
ANDN U4696 ( .B(n2818), .A(n2819), .Z(n2817) );
XOR U4697 ( .A(c939), .B(b[939]), .Z(n2818) );
XNOR U4698 ( .A(b[939]), .B(n2819), .Z(c[939]) );
XNOR U4699 ( .A(a[939]), .B(c939), .Z(n2819) );
XOR U4700 ( .A(c940), .B(n2820), .Z(c941) );
ANDN U4701 ( .B(n2821), .A(n2822), .Z(n2820) );
XOR U4702 ( .A(c940), .B(b[940]), .Z(n2821) );
XNOR U4703 ( .A(b[940]), .B(n2822), .Z(c[940]) );
XNOR U4704 ( .A(a[940]), .B(c940), .Z(n2822) );
XOR U4705 ( .A(c941), .B(n2823), .Z(c942) );
ANDN U4706 ( .B(n2824), .A(n2825), .Z(n2823) );
XOR U4707 ( .A(c941), .B(b[941]), .Z(n2824) );
XNOR U4708 ( .A(b[941]), .B(n2825), .Z(c[941]) );
XNOR U4709 ( .A(a[941]), .B(c941), .Z(n2825) );
XOR U4710 ( .A(c942), .B(n2826), .Z(c943) );
ANDN U4711 ( .B(n2827), .A(n2828), .Z(n2826) );
XOR U4712 ( .A(c942), .B(b[942]), .Z(n2827) );
XNOR U4713 ( .A(b[942]), .B(n2828), .Z(c[942]) );
XNOR U4714 ( .A(a[942]), .B(c942), .Z(n2828) );
XOR U4715 ( .A(c943), .B(n2829), .Z(c944) );
ANDN U4716 ( .B(n2830), .A(n2831), .Z(n2829) );
XOR U4717 ( .A(c943), .B(b[943]), .Z(n2830) );
XNOR U4718 ( .A(b[943]), .B(n2831), .Z(c[943]) );
XNOR U4719 ( .A(a[943]), .B(c943), .Z(n2831) );
XOR U4720 ( .A(c944), .B(n2832), .Z(c945) );
ANDN U4721 ( .B(n2833), .A(n2834), .Z(n2832) );
XOR U4722 ( .A(c944), .B(b[944]), .Z(n2833) );
XNOR U4723 ( .A(b[944]), .B(n2834), .Z(c[944]) );
XNOR U4724 ( .A(a[944]), .B(c944), .Z(n2834) );
XOR U4725 ( .A(c945), .B(n2835), .Z(c946) );
ANDN U4726 ( .B(n2836), .A(n2837), .Z(n2835) );
XOR U4727 ( .A(c945), .B(b[945]), .Z(n2836) );
XNOR U4728 ( .A(b[945]), .B(n2837), .Z(c[945]) );
XNOR U4729 ( .A(a[945]), .B(c945), .Z(n2837) );
XOR U4730 ( .A(c946), .B(n2838), .Z(c947) );
ANDN U4731 ( .B(n2839), .A(n2840), .Z(n2838) );
XOR U4732 ( .A(c946), .B(b[946]), .Z(n2839) );
XNOR U4733 ( .A(b[946]), .B(n2840), .Z(c[946]) );
XNOR U4734 ( .A(a[946]), .B(c946), .Z(n2840) );
XOR U4735 ( .A(c947), .B(n2841), .Z(c948) );
ANDN U4736 ( .B(n2842), .A(n2843), .Z(n2841) );
XOR U4737 ( .A(c947), .B(b[947]), .Z(n2842) );
XNOR U4738 ( .A(b[947]), .B(n2843), .Z(c[947]) );
XNOR U4739 ( .A(a[947]), .B(c947), .Z(n2843) );
XOR U4740 ( .A(c948), .B(n2844), .Z(c949) );
ANDN U4741 ( .B(n2845), .A(n2846), .Z(n2844) );
XOR U4742 ( .A(c948), .B(b[948]), .Z(n2845) );
XNOR U4743 ( .A(b[948]), .B(n2846), .Z(c[948]) );
XNOR U4744 ( .A(a[948]), .B(c948), .Z(n2846) );
XOR U4745 ( .A(c949), .B(n2847), .Z(c950) );
ANDN U4746 ( .B(n2848), .A(n2849), .Z(n2847) );
XOR U4747 ( .A(c949), .B(b[949]), .Z(n2848) );
XNOR U4748 ( .A(b[949]), .B(n2849), .Z(c[949]) );
XNOR U4749 ( .A(a[949]), .B(c949), .Z(n2849) );
XOR U4750 ( .A(c950), .B(n2850), .Z(c951) );
ANDN U4751 ( .B(n2851), .A(n2852), .Z(n2850) );
XOR U4752 ( .A(c950), .B(b[950]), .Z(n2851) );
XNOR U4753 ( .A(b[950]), .B(n2852), .Z(c[950]) );
XNOR U4754 ( .A(a[950]), .B(c950), .Z(n2852) );
XOR U4755 ( .A(c951), .B(n2853), .Z(c952) );
ANDN U4756 ( .B(n2854), .A(n2855), .Z(n2853) );
XOR U4757 ( .A(c951), .B(b[951]), .Z(n2854) );
XNOR U4758 ( .A(b[951]), .B(n2855), .Z(c[951]) );
XNOR U4759 ( .A(a[951]), .B(c951), .Z(n2855) );
XOR U4760 ( .A(c952), .B(n2856), .Z(c953) );
ANDN U4761 ( .B(n2857), .A(n2858), .Z(n2856) );
XOR U4762 ( .A(c952), .B(b[952]), .Z(n2857) );
XNOR U4763 ( .A(b[952]), .B(n2858), .Z(c[952]) );
XNOR U4764 ( .A(a[952]), .B(c952), .Z(n2858) );
XOR U4765 ( .A(c953), .B(n2859), .Z(c954) );
ANDN U4766 ( .B(n2860), .A(n2861), .Z(n2859) );
XOR U4767 ( .A(c953), .B(b[953]), .Z(n2860) );
XNOR U4768 ( .A(b[953]), .B(n2861), .Z(c[953]) );
XNOR U4769 ( .A(a[953]), .B(c953), .Z(n2861) );
XOR U4770 ( .A(c954), .B(n2862), .Z(c955) );
ANDN U4771 ( .B(n2863), .A(n2864), .Z(n2862) );
XOR U4772 ( .A(c954), .B(b[954]), .Z(n2863) );
XNOR U4773 ( .A(b[954]), .B(n2864), .Z(c[954]) );
XNOR U4774 ( .A(a[954]), .B(c954), .Z(n2864) );
XOR U4775 ( .A(c955), .B(n2865), .Z(c956) );
ANDN U4776 ( .B(n2866), .A(n2867), .Z(n2865) );
XOR U4777 ( .A(c955), .B(b[955]), .Z(n2866) );
XNOR U4778 ( .A(b[955]), .B(n2867), .Z(c[955]) );
XNOR U4779 ( .A(a[955]), .B(c955), .Z(n2867) );
XOR U4780 ( .A(c956), .B(n2868), .Z(c957) );
ANDN U4781 ( .B(n2869), .A(n2870), .Z(n2868) );
XOR U4782 ( .A(c956), .B(b[956]), .Z(n2869) );
XNOR U4783 ( .A(b[956]), .B(n2870), .Z(c[956]) );
XNOR U4784 ( .A(a[956]), .B(c956), .Z(n2870) );
XOR U4785 ( .A(c957), .B(n2871), .Z(c958) );
ANDN U4786 ( .B(n2872), .A(n2873), .Z(n2871) );
XOR U4787 ( .A(c957), .B(b[957]), .Z(n2872) );
XNOR U4788 ( .A(b[957]), .B(n2873), .Z(c[957]) );
XNOR U4789 ( .A(a[957]), .B(c957), .Z(n2873) );
XOR U4790 ( .A(c958), .B(n2874), .Z(c959) );
ANDN U4791 ( .B(n2875), .A(n2876), .Z(n2874) );
XOR U4792 ( .A(c958), .B(b[958]), .Z(n2875) );
XNOR U4793 ( .A(b[958]), .B(n2876), .Z(c[958]) );
XNOR U4794 ( .A(a[958]), .B(c958), .Z(n2876) );
XOR U4795 ( .A(c959), .B(n2877), .Z(c960) );
ANDN U4796 ( .B(n2878), .A(n2879), .Z(n2877) );
XOR U4797 ( .A(c959), .B(b[959]), .Z(n2878) );
XNOR U4798 ( .A(b[959]), .B(n2879), .Z(c[959]) );
XNOR U4799 ( .A(a[959]), .B(c959), .Z(n2879) );
XOR U4800 ( .A(c960), .B(n2880), .Z(c961) );
ANDN U4801 ( .B(n2881), .A(n2882), .Z(n2880) );
XOR U4802 ( .A(c960), .B(b[960]), .Z(n2881) );
XNOR U4803 ( .A(b[960]), .B(n2882), .Z(c[960]) );
XNOR U4804 ( .A(a[960]), .B(c960), .Z(n2882) );
XOR U4805 ( .A(c961), .B(n2883), .Z(c962) );
ANDN U4806 ( .B(n2884), .A(n2885), .Z(n2883) );
XOR U4807 ( .A(c961), .B(b[961]), .Z(n2884) );
XNOR U4808 ( .A(b[961]), .B(n2885), .Z(c[961]) );
XNOR U4809 ( .A(a[961]), .B(c961), .Z(n2885) );
XOR U4810 ( .A(c962), .B(n2886), .Z(c963) );
ANDN U4811 ( .B(n2887), .A(n2888), .Z(n2886) );
XOR U4812 ( .A(c962), .B(b[962]), .Z(n2887) );
XNOR U4813 ( .A(b[962]), .B(n2888), .Z(c[962]) );
XNOR U4814 ( .A(a[962]), .B(c962), .Z(n2888) );
XOR U4815 ( .A(c963), .B(n2889), .Z(c964) );
ANDN U4816 ( .B(n2890), .A(n2891), .Z(n2889) );
XOR U4817 ( .A(c963), .B(b[963]), .Z(n2890) );
XNOR U4818 ( .A(b[963]), .B(n2891), .Z(c[963]) );
XNOR U4819 ( .A(a[963]), .B(c963), .Z(n2891) );
XOR U4820 ( .A(c964), .B(n2892), .Z(c965) );
ANDN U4821 ( .B(n2893), .A(n2894), .Z(n2892) );
XOR U4822 ( .A(c964), .B(b[964]), .Z(n2893) );
XNOR U4823 ( .A(b[964]), .B(n2894), .Z(c[964]) );
XNOR U4824 ( .A(a[964]), .B(c964), .Z(n2894) );
XOR U4825 ( .A(c965), .B(n2895), .Z(c966) );
ANDN U4826 ( .B(n2896), .A(n2897), .Z(n2895) );
XOR U4827 ( .A(c965), .B(b[965]), .Z(n2896) );
XNOR U4828 ( .A(b[965]), .B(n2897), .Z(c[965]) );
XNOR U4829 ( .A(a[965]), .B(c965), .Z(n2897) );
XOR U4830 ( .A(c966), .B(n2898), .Z(c967) );
ANDN U4831 ( .B(n2899), .A(n2900), .Z(n2898) );
XOR U4832 ( .A(c966), .B(b[966]), .Z(n2899) );
XNOR U4833 ( .A(b[966]), .B(n2900), .Z(c[966]) );
XNOR U4834 ( .A(a[966]), .B(c966), .Z(n2900) );
XOR U4835 ( .A(c967), .B(n2901), .Z(c968) );
ANDN U4836 ( .B(n2902), .A(n2903), .Z(n2901) );
XOR U4837 ( .A(c967), .B(b[967]), .Z(n2902) );
XNOR U4838 ( .A(b[967]), .B(n2903), .Z(c[967]) );
XNOR U4839 ( .A(a[967]), .B(c967), .Z(n2903) );
XOR U4840 ( .A(c968), .B(n2904), .Z(c969) );
ANDN U4841 ( .B(n2905), .A(n2906), .Z(n2904) );
XOR U4842 ( .A(c968), .B(b[968]), .Z(n2905) );
XNOR U4843 ( .A(b[968]), .B(n2906), .Z(c[968]) );
XNOR U4844 ( .A(a[968]), .B(c968), .Z(n2906) );
XOR U4845 ( .A(c969), .B(n2907), .Z(c970) );
ANDN U4846 ( .B(n2908), .A(n2909), .Z(n2907) );
XOR U4847 ( .A(c969), .B(b[969]), .Z(n2908) );
XNOR U4848 ( .A(b[969]), .B(n2909), .Z(c[969]) );
XNOR U4849 ( .A(a[969]), .B(c969), .Z(n2909) );
XOR U4850 ( .A(c970), .B(n2910), .Z(c971) );
ANDN U4851 ( .B(n2911), .A(n2912), .Z(n2910) );
XOR U4852 ( .A(c970), .B(b[970]), .Z(n2911) );
XNOR U4853 ( .A(b[970]), .B(n2912), .Z(c[970]) );
XNOR U4854 ( .A(a[970]), .B(c970), .Z(n2912) );
XOR U4855 ( .A(c971), .B(n2913), .Z(c972) );
ANDN U4856 ( .B(n2914), .A(n2915), .Z(n2913) );
XOR U4857 ( .A(c971), .B(b[971]), .Z(n2914) );
XNOR U4858 ( .A(b[971]), .B(n2915), .Z(c[971]) );
XNOR U4859 ( .A(a[971]), .B(c971), .Z(n2915) );
XOR U4860 ( .A(c972), .B(n2916), .Z(c973) );
ANDN U4861 ( .B(n2917), .A(n2918), .Z(n2916) );
XOR U4862 ( .A(c972), .B(b[972]), .Z(n2917) );
XNOR U4863 ( .A(b[972]), .B(n2918), .Z(c[972]) );
XNOR U4864 ( .A(a[972]), .B(c972), .Z(n2918) );
XOR U4865 ( .A(c973), .B(n2919), .Z(c974) );
ANDN U4866 ( .B(n2920), .A(n2921), .Z(n2919) );
XOR U4867 ( .A(c973), .B(b[973]), .Z(n2920) );
XNOR U4868 ( .A(b[973]), .B(n2921), .Z(c[973]) );
XNOR U4869 ( .A(a[973]), .B(c973), .Z(n2921) );
XOR U4870 ( .A(c974), .B(n2922), .Z(c975) );
ANDN U4871 ( .B(n2923), .A(n2924), .Z(n2922) );
XOR U4872 ( .A(c974), .B(b[974]), .Z(n2923) );
XNOR U4873 ( .A(b[974]), .B(n2924), .Z(c[974]) );
XNOR U4874 ( .A(a[974]), .B(c974), .Z(n2924) );
XOR U4875 ( .A(c975), .B(n2925), .Z(c976) );
ANDN U4876 ( .B(n2926), .A(n2927), .Z(n2925) );
XOR U4877 ( .A(c975), .B(b[975]), .Z(n2926) );
XNOR U4878 ( .A(b[975]), .B(n2927), .Z(c[975]) );
XNOR U4879 ( .A(a[975]), .B(c975), .Z(n2927) );
XOR U4880 ( .A(c976), .B(n2928), .Z(c977) );
ANDN U4881 ( .B(n2929), .A(n2930), .Z(n2928) );
XOR U4882 ( .A(c976), .B(b[976]), .Z(n2929) );
XNOR U4883 ( .A(b[976]), .B(n2930), .Z(c[976]) );
XNOR U4884 ( .A(a[976]), .B(c976), .Z(n2930) );
XOR U4885 ( .A(c977), .B(n2931), .Z(c978) );
ANDN U4886 ( .B(n2932), .A(n2933), .Z(n2931) );
XOR U4887 ( .A(c977), .B(b[977]), .Z(n2932) );
XNOR U4888 ( .A(b[977]), .B(n2933), .Z(c[977]) );
XNOR U4889 ( .A(a[977]), .B(c977), .Z(n2933) );
XOR U4890 ( .A(c978), .B(n2934), .Z(c979) );
ANDN U4891 ( .B(n2935), .A(n2936), .Z(n2934) );
XOR U4892 ( .A(c978), .B(b[978]), .Z(n2935) );
XNOR U4893 ( .A(b[978]), .B(n2936), .Z(c[978]) );
XNOR U4894 ( .A(a[978]), .B(c978), .Z(n2936) );
XOR U4895 ( .A(c979), .B(n2937), .Z(c980) );
ANDN U4896 ( .B(n2938), .A(n2939), .Z(n2937) );
XOR U4897 ( .A(c979), .B(b[979]), .Z(n2938) );
XNOR U4898 ( .A(b[979]), .B(n2939), .Z(c[979]) );
XNOR U4899 ( .A(a[979]), .B(c979), .Z(n2939) );
XOR U4900 ( .A(c980), .B(n2940), .Z(c981) );
ANDN U4901 ( .B(n2941), .A(n2942), .Z(n2940) );
XOR U4902 ( .A(c980), .B(b[980]), .Z(n2941) );
XNOR U4903 ( .A(b[980]), .B(n2942), .Z(c[980]) );
XNOR U4904 ( .A(a[980]), .B(c980), .Z(n2942) );
XOR U4905 ( .A(c981), .B(n2943), .Z(c982) );
ANDN U4906 ( .B(n2944), .A(n2945), .Z(n2943) );
XOR U4907 ( .A(c981), .B(b[981]), .Z(n2944) );
XNOR U4908 ( .A(b[981]), .B(n2945), .Z(c[981]) );
XNOR U4909 ( .A(a[981]), .B(c981), .Z(n2945) );
XOR U4910 ( .A(c982), .B(n2946), .Z(c983) );
ANDN U4911 ( .B(n2947), .A(n2948), .Z(n2946) );
XOR U4912 ( .A(c982), .B(b[982]), .Z(n2947) );
XNOR U4913 ( .A(b[982]), .B(n2948), .Z(c[982]) );
XNOR U4914 ( .A(a[982]), .B(c982), .Z(n2948) );
XOR U4915 ( .A(c983), .B(n2949), .Z(c984) );
ANDN U4916 ( .B(n2950), .A(n2951), .Z(n2949) );
XOR U4917 ( .A(c983), .B(b[983]), .Z(n2950) );
XNOR U4918 ( .A(b[983]), .B(n2951), .Z(c[983]) );
XNOR U4919 ( .A(a[983]), .B(c983), .Z(n2951) );
XOR U4920 ( .A(c984), .B(n2952), .Z(c985) );
ANDN U4921 ( .B(n2953), .A(n2954), .Z(n2952) );
XOR U4922 ( .A(c984), .B(b[984]), .Z(n2953) );
XNOR U4923 ( .A(b[984]), .B(n2954), .Z(c[984]) );
XNOR U4924 ( .A(a[984]), .B(c984), .Z(n2954) );
XOR U4925 ( .A(c985), .B(n2955), .Z(c986) );
ANDN U4926 ( .B(n2956), .A(n2957), .Z(n2955) );
XOR U4927 ( .A(c985), .B(b[985]), .Z(n2956) );
XNOR U4928 ( .A(b[985]), .B(n2957), .Z(c[985]) );
XNOR U4929 ( .A(a[985]), .B(c985), .Z(n2957) );
XOR U4930 ( .A(c986), .B(n2958), .Z(c987) );
ANDN U4931 ( .B(n2959), .A(n2960), .Z(n2958) );
XOR U4932 ( .A(c986), .B(b[986]), .Z(n2959) );
XNOR U4933 ( .A(b[986]), .B(n2960), .Z(c[986]) );
XNOR U4934 ( .A(a[986]), .B(c986), .Z(n2960) );
XOR U4935 ( .A(c987), .B(n2961), .Z(c988) );
ANDN U4936 ( .B(n2962), .A(n2963), .Z(n2961) );
XOR U4937 ( .A(c987), .B(b[987]), .Z(n2962) );
XNOR U4938 ( .A(b[987]), .B(n2963), .Z(c[987]) );
XNOR U4939 ( .A(a[987]), .B(c987), .Z(n2963) );
XOR U4940 ( .A(c988), .B(n2964), .Z(c989) );
ANDN U4941 ( .B(n2965), .A(n2966), .Z(n2964) );
XOR U4942 ( .A(c988), .B(b[988]), .Z(n2965) );
XNOR U4943 ( .A(b[988]), .B(n2966), .Z(c[988]) );
XNOR U4944 ( .A(a[988]), .B(c988), .Z(n2966) );
XOR U4945 ( .A(c989), .B(n2967), .Z(c990) );
ANDN U4946 ( .B(n2968), .A(n2969), .Z(n2967) );
XOR U4947 ( .A(c989), .B(b[989]), .Z(n2968) );
XNOR U4948 ( .A(b[989]), .B(n2969), .Z(c[989]) );
XNOR U4949 ( .A(a[989]), .B(c989), .Z(n2969) );
XOR U4950 ( .A(c990), .B(n2970), .Z(c991) );
ANDN U4951 ( .B(n2971), .A(n2972), .Z(n2970) );
XOR U4952 ( .A(c990), .B(b[990]), .Z(n2971) );
XNOR U4953 ( .A(b[990]), .B(n2972), .Z(c[990]) );
XNOR U4954 ( .A(a[990]), .B(c990), .Z(n2972) );
XOR U4955 ( .A(c991), .B(n2973), .Z(c992) );
ANDN U4956 ( .B(n2974), .A(n2975), .Z(n2973) );
XOR U4957 ( .A(c991), .B(b[991]), .Z(n2974) );
XNOR U4958 ( .A(b[991]), .B(n2975), .Z(c[991]) );
XNOR U4959 ( .A(a[991]), .B(c991), .Z(n2975) );
XOR U4960 ( .A(c992), .B(n2976), .Z(c993) );
ANDN U4961 ( .B(n2977), .A(n2978), .Z(n2976) );
XOR U4962 ( .A(c992), .B(b[992]), .Z(n2977) );
XNOR U4963 ( .A(b[992]), .B(n2978), .Z(c[992]) );
XNOR U4964 ( .A(a[992]), .B(c992), .Z(n2978) );
XOR U4965 ( .A(c993), .B(n2979), .Z(c994) );
ANDN U4966 ( .B(n2980), .A(n2981), .Z(n2979) );
XOR U4967 ( .A(c993), .B(b[993]), .Z(n2980) );
XNOR U4968 ( .A(b[993]), .B(n2981), .Z(c[993]) );
XNOR U4969 ( .A(a[993]), .B(c993), .Z(n2981) );
XOR U4970 ( .A(c994), .B(n2982), .Z(c995) );
ANDN U4971 ( .B(n2983), .A(n2984), .Z(n2982) );
XOR U4972 ( .A(c994), .B(b[994]), .Z(n2983) );
XNOR U4973 ( .A(b[994]), .B(n2984), .Z(c[994]) );
XNOR U4974 ( .A(a[994]), .B(c994), .Z(n2984) );
XOR U4975 ( .A(c995), .B(n2985), .Z(c996) );
ANDN U4976 ( .B(n2986), .A(n2987), .Z(n2985) );
XOR U4977 ( .A(c995), .B(b[995]), .Z(n2986) );
XNOR U4978 ( .A(b[995]), .B(n2987), .Z(c[995]) );
XNOR U4979 ( .A(a[995]), .B(c995), .Z(n2987) );
XOR U4980 ( .A(c996), .B(n2988), .Z(c997) );
ANDN U4981 ( .B(n2989), .A(n2990), .Z(n2988) );
XOR U4982 ( .A(c996), .B(b[996]), .Z(n2989) );
XNOR U4983 ( .A(b[996]), .B(n2990), .Z(c[996]) );
XNOR U4984 ( .A(a[996]), .B(c996), .Z(n2990) );
XOR U4985 ( .A(c997), .B(n2991), .Z(c998) );
ANDN U4986 ( .B(n2992), .A(n2993), .Z(n2991) );
XOR U4987 ( .A(c997), .B(b[997]), .Z(n2992) );
XNOR U4988 ( .A(b[997]), .B(n2993), .Z(c[997]) );
XNOR U4989 ( .A(a[997]), .B(c997), .Z(n2993) );
XOR U4990 ( .A(c998), .B(n2994), .Z(c999) );
ANDN U4991 ( .B(n2995), .A(n2996), .Z(n2994) );
XOR U4992 ( .A(c998), .B(b[998]), .Z(n2995) );
XNOR U4993 ( .A(b[998]), .B(n2996), .Z(c[998]) );
XNOR U4994 ( .A(a[998]), .B(c998), .Z(n2996) );
XOR U4995 ( .A(c999), .B(n2997), .Z(c1000) );
ANDN U4996 ( .B(n2998), .A(n2999), .Z(n2997) );
XOR U4997 ( .A(c999), .B(b[999]), .Z(n2998) );
XNOR U4998 ( .A(b[999]), .B(n2999), .Z(c[999]) );
XNOR U4999 ( .A(a[999]), .B(c999), .Z(n2999) );
XOR U5000 ( .A(c1000), .B(n3000), .Z(c1001) );
ANDN U5001 ( .B(n3001), .A(n3002), .Z(n3000) );
XOR U5002 ( .A(c1000), .B(b[1000]), .Z(n3001) );
XNOR U5003 ( .A(b[1000]), .B(n3002), .Z(c[1000]) );
XNOR U5004 ( .A(a[1000]), .B(c1000), .Z(n3002) );
XOR U5005 ( .A(c1001), .B(n3003), .Z(c1002) );
ANDN U5006 ( .B(n3004), .A(n3005), .Z(n3003) );
XOR U5007 ( .A(c1001), .B(b[1001]), .Z(n3004) );
XNOR U5008 ( .A(b[1001]), .B(n3005), .Z(c[1001]) );
XNOR U5009 ( .A(a[1001]), .B(c1001), .Z(n3005) );
XOR U5010 ( .A(c1002), .B(n3006), .Z(c1003) );
ANDN U5011 ( .B(n3007), .A(n3008), .Z(n3006) );
XOR U5012 ( .A(c1002), .B(b[1002]), .Z(n3007) );
XNOR U5013 ( .A(b[1002]), .B(n3008), .Z(c[1002]) );
XNOR U5014 ( .A(a[1002]), .B(c1002), .Z(n3008) );
XOR U5015 ( .A(c1003), .B(n3009), .Z(c1004) );
ANDN U5016 ( .B(n3010), .A(n3011), .Z(n3009) );
XOR U5017 ( .A(c1003), .B(b[1003]), .Z(n3010) );
XNOR U5018 ( .A(b[1003]), .B(n3011), .Z(c[1003]) );
XNOR U5019 ( .A(a[1003]), .B(c1003), .Z(n3011) );
XOR U5020 ( .A(c1004), .B(n3012), .Z(c1005) );
ANDN U5021 ( .B(n3013), .A(n3014), .Z(n3012) );
XOR U5022 ( .A(c1004), .B(b[1004]), .Z(n3013) );
XNOR U5023 ( .A(b[1004]), .B(n3014), .Z(c[1004]) );
XNOR U5024 ( .A(a[1004]), .B(c1004), .Z(n3014) );
XOR U5025 ( .A(c1005), .B(n3015), .Z(c1006) );
ANDN U5026 ( .B(n3016), .A(n3017), .Z(n3015) );
XOR U5027 ( .A(c1005), .B(b[1005]), .Z(n3016) );
XNOR U5028 ( .A(b[1005]), .B(n3017), .Z(c[1005]) );
XNOR U5029 ( .A(a[1005]), .B(c1005), .Z(n3017) );
XOR U5030 ( .A(c1006), .B(n3018), .Z(c1007) );
ANDN U5031 ( .B(n3019), .A(n3020), .Z(n3018) );
XOR U5032 ( .A(c1006), .B(b[1006]), .Z(n3019) );
XNOR U5033 ( .A(b[1006]), .B(n3020), .Z(c[1006]) );
XNOR U5034 ( .A(a[1006]), .B(c1006), .Z(n3020) );
XOR U5035 ( .A(c1007), .B(n3021), .Z(c1008) );
ANDN U5036 ( .B(n3022), .A(n3023), .Z(n3021) );
XOR U5037 ( .A(c1007), .B(b[1007]), .Z(n3022) );
XNOR U5038 ( .A(b[1007]), .B(n3023), .Z(c[1007]) );
XNOR U5039 ( .A(a[1007]), .B(c1007), .Z(n3023) );
XOR U5040 ( .A(c1008), .B(n3024), .Z(c1009) );
ANDN U5041 ( .B(n3025), .A(n3026), .Z(n3024) );
XOR U5042 ( .A(c1008), .B(b[1008]), .Z(n3025) );
XNOR U5043 ( .A(b[1008]), .B(n3026), .Z(c[1008]) );
XNOR U5044 ( .A(a[1008]), .B(c1008), .Z(n3026) );
XOR U5045 ( .A(c1009), .B(n3027), .Z(c1010) );
ANDN U5046 ( .B(n3028), .A(n3029), .Z(n3027) );
XOR U5047 ( .A(c1009), .B(b[1009]), .Z(n3028) );
XNOR U5048 ( .A(b[1009]), .B(n3029), .Z(c[1009]) );
XNOR U5049 ( .A(a[1009]), .B(c1009), .Z(n3029) );
XOR U5050 ( .A(c1010), .B(n3030), .Z(c1011) );
ANDN U5051 ( .B(n3031), .A(n3032), .Z(n3030) );
XOR U5052 ( .A(c1010), .B(b[1010]), .Z(n3031) );
XNOR U5053 ( .A(b[1010]), .B(n3032), .Z(c[1010]) );
XNOR U5054 ( .A(a[1010]), .B(c1010), .Z(n3032) );
XOR U5055 ( .A(c1011), .B(n3033), .Z(c1012) );
ANDN U5056 ( .B(n3034), .A(n3035), .Z(n3033) );
XOR U5057 ( .A(c1011), .B(b[1011]), .Z(n3034) );
XNOR U5058 ( .A(b[1011]), .B(n3035), .Z(c[1011]) );
XNOR U5059 ( .A(a[1011]), .B(c1011), .Z(n3035) );
XOR U5060 ( .A(c1012), .B(n3036), .Z(c1013) );
ANDN U5061 ( .B(n3037), .A(n3038), .Z(n3036) );
XOR U5062 ( .A(c1012), .B(b[1012]), .Z(n3037) );
XNOR U5063 ( .A(b[1012]), .B(n3038), .Z(c[1012]) );
XNOR U5064 ( .A(a[1012]), .B(c1012), .Z(n3038) );
XOR U5065 ( .A(c1013), .B(n3039), .Z(c1014) );
ANDN U5066 ( .B(n3040), .A(n3041), .Z(n3039) );
XOR U5067 ( .A(c1013), .B(b[1013]), .Z(n3040) );
XNOR U5068 ( .A(b[1013]), .B(n3041), .Z(c[1013]) );
XNOR U5069 ( .A(a[1013]), .B(c1013), .Z(n3041) );
XOR U5070 ( .A(c1014), .B(n3042), .Z(c1015) );
ANDN U5071 ( .B(n3043), .A(n3044), .Z(n3042) );
XOR U5072 ( .A(c1014), .B(b[1014]), .Z(n3043) );
XNOR U5073 ( .A(b[1014]), .B(n3044), .Z(c[1014]) );
XNOR U5074 ( .A(a[1014]), .B(c1014), .Z(n3044) );
XOR U5075 ( .A(c1015), .B(n3045), .Z(c1016) );
ANDN U5076 ( .B(n3046), .A(n3047), .Z(n3045) );
XOR U5077 ( .A(c1015), .B(b[1015]), .Z(n3046) );
XNOR U5078 ( .A(b[1015]), .B(n3047), .Z(c[1015]) );
XNOR U5079 ( .A(a[1015]), .B(c1015), .Z(n3047) );
XOR U5080 ( .A(c1016), .B(n3048), .Z(c1017) );
ANDN U5081 ( .B(n3049), .A(n3050), .Z(n3048) );
XOR U5082 ( .A(c1016), .B(b[1016]), .Z(n3049) );
XNOR U5083 ( .A(b[1016]), .B(n3050), .Z(c[1016]) );
XNOR U5084 ( .A(a[1016]), .B(c1016), .Z(n3050) );
XOR U5085 ( .A(c1017), .B(n3051), .Z(c1018) );
ANDN U5086 ( .B(n3052), .A(n3053), .Z(n3051) );
XOR U5087 ( .A(c1017), .B(b[1017]), .Z(n3052) );
XNOR U5088 ( .A(b[1017]), .B(n3053), .Z(c[1017]) );
XNOR U5089 ( .A(a[1017]), .B(c1017), .Z(n3053) );
XOR U5090 ( .A(c1018), .B(n3054), .Z(c1019) );
ANDN U5091 ( .B(n3055), .A(n3056), .Z(n3054) );
XOR U5092 ( .A(c1018), .B(b[1018]), .Z(n3055) );
XNOR U5093 ( .A(b[1018]), .B(n3056), .Z(c[1018]) );
XNOR U5094 ( .A(a[1018]), .B(c1018), .Z(n3056) );
XOR U5095 ( .A(c1019), .B(n3057), .Z(c1020) );
ANDN U5096 ( .B(n3058), .A(n3059), .Z(n3057) );
XOR U5097 ( .A(c1019), .B(b[1019]), .Z(n3058) );
XNOR U5098 ( .A(b[1019]), .B(n3059), .Z(c[1019]) );
XNOR U5099 ( .A(a[1019]), .B(c1019), .Z(n3059) );
XOR U5100 ( .A(c1020), .B(n3060), .Z(c1021) );
ANDN U5101 ( .B(n3061), .A(n3062), .Z(n3060) );
XOR U5102 ( .A(c1020), .B(b[1020]), .Z(n3061) );
XNOR U5103 ( .A(b[1020]), .B(n3062), .Z(c[1020]) );
XNOR U5104 ( .A(a[1020]), .B(c1020), .Z(n3062) );
XOR U5105 ( .A(c1021), .B(n3063), .Z(c1022) );
ANDN U5106 ( .B(n3064), .A(n3065), .Z(n3063) );
XOR U5107 ( .A(c1021), .B(b[1021]), .Z(n3064) );
XNOR U5108 ( .A(b[1021]), .B(n3065), .Z(c[1021]) );
XNOR U5109 ( .A(a[1021]), .B(c1021), .Z(n3065) );
XOR U5110 ( .A(c1022), .B(n3066), .Z(c1023) );
ANDN U5111 ( .B(n3067), .A(n3068), .Z(n3066) );
XOR U5112 ( .A(c1022), .B(b[1022]), .Z(n3067) );
XNOR U5113 ( .A(b[1022]), .B(n3068), .Z(c[1022]) );
XNOR U5114 ( .A(a[1022]), .B(c1022), .Z(n3068) );
XOR U5115 ( .A(c1023), .B(n3069), .Z(c1024) );
ANDN U5116 ( .B(n3070), .A(n3071), .Z(n3069) );
XOR U5117 ( .A(c1023), .B(b[1023]), .Z(n3070) );
XNOR U5118 ( .A(b[1023]), .B(n3071), .Z(c[1023]) );
XNOR U5119 ( .A(a[1023]), .B(c1023), .Z(n3071) );
XOR U5120 ( .A(c1024), .B(n3072), .Z(c1025) );
ANDN U5121 ( .B(n3073), .A(n3074), .Z(n3072) );
XOR U5122 ( .A(c1024), .B(b[1024]), .Z(n3073) );
XNOR U5123 ( .A(b[1024]), .B(n3074), .Z(c[1024]) );
XNOR U5124 ( .A(a[1024]), .B(c1024), .Z(n3074) );
XOR U5125 ( .A(c1025), .B(n3075), .Z(c1026) );
ANDN U5126 ( .B(n3076), .A(n3077), .Z(n3075) );
XOR U5127 ( .A(c1025), .B(b[1025]), .Z(n3076) );
XNOR U5128 ( .A(b[1025]), .B(n3077), .Z(c[1025]) );
XNOR U5129 ( .A(a[1025]), .B(c1025), .Z(n3077) );
XOR U5130 ( .A(c1026), .B(n3078), .Z(c1027) );
ANDN U5131 ( .B(n3079), .A(n3080), .Z(n3078) );
XOR U5132 ( .A(c1026), .B(b[1026]), .Z(n3079) );
XNOR U5133 ( .A(b[1026]), .B(n3080), .Z(c[1026]) );
XNOR U5134 ( .A(a[1026]), .B(c1026), .Z(n3080) );
XOR U5135 ( .A(c1027), .B(n3081), .Z(c1028) );
ANDN U5136 ( .B(n3082), .A(n3083), .Z(n3081) );
XOR U5137 ( .A(c1027), .B(b[1027]), .Z(n3082) );
XNOR U5138 ( .A(b[1027]), .B(n3083), .Z(c[1027]) );
XNOR U5139 ( .A(a[1027]), .B(c1027), .Z(n3083) );
XOR U5140 ( .A(c1028), .B(n3084), .Z(c1029) );
ANDN U5141 ( .B(n3085), .A(n3086), .Z(n3084) );
XOR U5142 ( .A(c1028), .B(b[1028]), .Z(n3085) );
XNOR U5143 ( .A(b[1028]), .B(n3086), .Z(c[1028]) );
XNOR U5144 ( .A(a[1028]), .B(c1028), .Z(n3086) );
XOR U5145 ( .A(c1029), .B(n3087), .Z(c1030) );
ANDN U5146 ( .B(n3088), .A(n3089), .Z(n3087) );
XOR U5147 ( .A(c1029), .B(b[1029]), .Z(n3088) );
XNOR U5148 ( .A(b[1029]), .B(n3089), .Z(c[1029]) );
XNOR U5149 ( .A(a[1029]), .B(c1029), .Z(n3089) );
XOR U5150 ( .A(c1030), .B(n3090), .Z(c1031) );
ANDN U5151 ( .B(n3091), .A(n3092), .Z(n3090) );
XOR U5152 ( .A(c1030), .B(b[1030]), .Z(n3091) );
XNOR U5153 ( .A(b[1030]), .B(n3092), .Z(c[1030]) );
XNOR U5154 ( .A(a[1030]), .B(c1030), .Z(n3092) );
XOR U5155 ( .A(c1031), .B(n3093), .Z(c1032) );
ANDN U5156 ( .B(n3094), .A(n3095), .Z(n3093) );
XOR U5157 ( .A(c1031), .B(b[1031]), .Z(n3094) );
XNOR U5158 ( .A(b[1031]), .B(n3095), .Z(c[1031]) );
XNOR U5159 ( .A(a[1031]), .B(c1031), .Z(n3095) );
XOR U5160 ( .A(c1032), .B(n3096), .Z(c1033) );
ANDN U5161 ( .B(n3097), .A(n3098), .Z(n3096) );
XOR U5162 ( .A(c1032), .B(b[1032]), .Z(n3097) );
XNOR U5163 ( .A(b[1032]), .B(n3098), .Z(c[1032]) );
XNOR U5164 ( .A(a[1032]), .B(c1032), .Z(n3098) );
XOR U5165 ( .A(c1033), .B(n3099), .Z(c1034) );
ANDN U5166 ( .B(n3100), .A(n3101), .Z(n3099) );
XOR U5167 ( .A(c1033), .B(b[1033]), .Z(n3100) );
XNOR U5168 ( .A(b[1033]), .B(n3101), .Z(c[1033]) );
XNOR U5169 ( .A(a[1033]), .B(c1033), .Z(n3101) );
XOR U5170 ( .A(c1034), .B(n3102), .Z(c1035) );
ANDN U5171 ( .B(n3103), .A(n3104), .Z(n3102) );
XOR U5172 ( .A(c1034), .B(b[1034]), .Z(n3103) );
XNOR U5173 ( .A(b[1034]), .B(n3104), .Z(c[1034]) );
XNOR U5174 ( .A(a[1034]), .B(c1034), .Z(n3104) );
XOR U5175 ( .A(c1035), .B(n3105), .Z(c1036) );
ANDN U5176 ( .B(n3106), .A(n3107), .Z(n3105) );
XOR U5177 ( .A(c1035), .B(b[1035]), .Z(n3106) );
XNOR U5178 ( .A(b[1035]), .B(n3107), .Z(c[1035]) );
XNOR U5179 ( .A(a[1035]), .B(c1035), .Z(n3107) );
XOR U5180 ( .A(c1036), .B(n3108), .Z(c1037) );
ANDN U5181 ( .B(n3109), .A(n3110), .Z(n3108) );
XOR U5182 ( .A(c1036), .B(b[1036]), .Z(n3109) );
XNOR U5183 ( .A(b[1036]), .B(n3110), .Z(c[1036]) );
XNOR U5184 ( .A(a[1036]), .B(c1036), .Z(n3110) );
XOR U5185 ( .A(c1037), .B(n3111), .Z(c1038) );
ANDN U5186 ( .B(n3112), .A(n3113), .Z(n3111) );
XOR U5187 ( .A(c1037), .B(b[1037]), .Z(n3112) );
XNOR U5188 ( .A(b[1037]), .B(n3113), .Z(c[1037]) );
XNOR U5189 ( .A(a[1037]), .B(c1037), .Z(n3113) );
XOR U5190 ( .A(c1038), .B(n3114), .Z(c1039) );
ANDN U5191 ( .B(n3115), .A(n3116), .Z(n3114) );
XOR U5192 ( .A(c1038), .B(b[1038]), .Z(n3115) );
XNOR U5193 ( .A(b[1038]), .B(n3116), .Z(c[1038]) );
XNOR U5194 ( .A(a[1038]), .B(c1038), .Z(n3116) );
XOR U5195 ( .A(c1039), .B(n3117), .Z(c1040) );
ANDN U5196 ( .B(n3118), .A(n3119), .Z(n3117) );
XOR U5197 ( .A(c1039), .B(b[1039]), .Z(n3118) );
XNOR U5198 ( .A(b[1039]), .B(n3119), .Z(c[1039]) );
XNOR U5199 ( .A(a[1039]), .B(c1039), .Z(n3119) );
XOR U5200 ( .A(c1040), .B(n3120), .Z(c1041) );
ANDN U5201 ( .B(n3121), .A(n3122), .Z(n3120) );
XOR U5202 ( .A(c1040), .B(b[1040]), .Z(n3121) );
XNOR U5203 ( .A(b[1040]), .B(n3122), .Z(c[1040]) );
XNOR U5204 ( .A(a[1040]), .B(c1040), .Z(n3122) );
XOR U5205 ( .A(c1041), .B(n3123), .Z(c1042) );
ANDN U5206 ( .B(n3124), .A(n3125), .Z(n3123) );
XOR U5207 ( .A(c1041), .B(b[1041]), .Z(n3124) );
XNOR U5208 ( .A(b[1041]), .B(n3125), .Z(c[1041]) );
XNOR U5209 ( .A(a[1041]), .B(c1041), .Z(n3125) );
XOR U5210 ( .A(c1042), .B(n3126), .Z(c1043) );
ANDN U5211 ( .B(n3127), .A(n3128), .Z(n3126) );
XOR U5212 ( .A(c1042), .B(b[1042]), .Z(n3127) );
XNOR U5213 ( .A(b[1042]), .B(n3128), .Z(c[1042]) );
XNOR U5214 ( .A(a[1042]), .B(c1042), .Z(n3128) );
XOR U5215 ( .A(c1043), .B(n3129), .Z(c1044) );
ANDN U5216 ( .B(n3130), .A(n3131), .Z(n3129) );
XOR U5217 ( .A(c1043), .B(b[1043]), .Z(n3130) );
XNOR U5218 ( .A(b[1043]), .B(n3131), .Z(c[1043]) );
XNOR U5219 ( .A(a[1043]), .B(c1043), .Z(n3131) );
XOR U5220 ( .A(c1044), .B(n3132), .Z(c1045) );
ANDN U5221 ( .B(n3133), .A(n3134), .Z(n3132) );
XOR U5222 ( .A(c1044), .B(b[1044]), .Z(n3133) );
XNOR U5223 ( .A(b[1044]), .B(n3134), .Z(c[1044]) );
XNOR U5224 ( .A(a[1044]), .B(c1044), .Z(n3134) );
XOR U5225 ( .A(c1045), .B(n3135), .Z(c1046) );
ANDN U5226 ( .B(n3136), .A(n3137), .Z(n3135) );
XOR U5227 ( .A(c1045), .B(b[1045]), .Z(n3136) );
XNOR U5228 ( .A(b[1045]), .B(n3137), .Z(c[1045]) );
XNOR U5229 ( .A(a[1045]), .B(c1045), .Z(n3137) );
XOR U5230 ( .A(c1046), .B(n3138), .Z(c1047) );
ANDN U5231 ( .B(n3139), .A(n3140), .Z(n3138) );
XOR U5232 ( .A(c1046), .B(b[1046]), .Z(n3139) );
XNOR U5233 ( .A(b[1046]), .B(n3140), .Z(c[1046]) );
XNOR U5234 ( .A(a[1046]), .B(c1046), .Z(n3140) );
XOR U5235 ( .A(c1047), .B(n3141), .Z(c1048) );
ANDN U5236 ( .B(n3142), .A(n3143), .Z(n3141) );
XOR U5237 ( .A(c1047), .B(b[1047]), .Z(n3142) );
XNOR U5238 ( .A(b[1047]), .B(n3143), .Z(c[1047]) );
XNOR U5239 ( .A(a[1047]), .B(c1047), .Z(n3143) );
XOR U5240 ( .A(c1048), .B(n3144), .Z(c1049) );
ANDN U5241 ( .B(n3145), .A(n3146), .Z(n3144) );
XOR U5242 ( .A(c1048), .B(b[1048]), .Z(n3145) );
XNOR U5243 ( .A(b[1048]), .B(n3146), .Z(c[1048]) );
XNOR U5244 ( .A(a[1048]), .B(c1048), .Z(n3146) );
XOR U5245 ( .A(c1049), .B(n3147), .Z(c1050) );
ANDN U5246 ( .B(n3148), .A(n3149), .Z(n3147) );
XOR U5247 ( .A(c1049), .B(b[1049]), .Z(n3148) );
XNOR U5248 ( .A(b[1049]), .B(n3149), .Z(c[1049]) );
XNOR U5249 ( .A(a[1049]), .B(c1049), .Z(n3149) );
XOR U5250 ( .A(c1050), .B(n3150), .Z(c1051) );
ANDN U5251 ( .B(n3151), .A(n3152), .Z(n3150) );
XOR U5252 ( .A(c1050), .B(b[1050]), .Z(n3151) );
XNOR U5253 ( .A(b[1050]), .B(n3152), .Z(c[1050]) );
XNOR U5254 ( .A(a[1050]), .B(c1050), .Z(n3152) );
XOR U5255 ( .A(c1051), .B(n3153), .Z(c1052) );
ANDN U5256 ( .B(n3154), .A(n3155), .Z(n3153) );
XOR U5257 ( .A(c1051), .B(b[1051]), .Z(n3154) );
XNOR U5258 ( .A(b[1051]), .B(n3155), .Z(c[1051]) );
XNOR U5259 ( .A(a[1051]), .B(c1051), .Z(n3155) );
XOR U5260 ( .A(c1052), .B(n3156), .Z(c1053) );
ANDN U5261 ( .B(n3157), .A(n3158), .Z(n3156) );
XOR U5262 ( .A(c1052), .B(b[1052]), .Z(n3157) );
XNOR U5263 ( .A(b[1052]), .B(n3158), .Z(c[1052]) );
XNOR U5264 ( .A(a[1052]), .B(c1052), .Z(n3158) );
XOR U5265 ( .A(c1053), .B(n3159), .Z(c1054) );
ANDN U5266 ( .B(n3160), .A(n3161), .Z(n3159) );
XOR U5267 ( .A(c1053), .B(b[1053]), .Z(n3160) );
XNOR U5268 ( .A(b[1053]), .B(n3161), .Z(c[1053]) );
XNOR U5269 ( .A(a[1053]), .B(c1053), .Z(n3161) );
XOR U5270 ( .A(c1054), .B(n3162), .Z(c1055) );
ANDN U5271 ( .B(n3163), .A(n3164), .Z(n3162) );
XOR U5272 ( .A(c1054), .B(b[1054]), .Z(n3163) );
XNOR U5273 ( .A(b[1054]), .B(n3164), .Z(c[1054]) );
XNOR U5274 ( .A(a[1054]), .B(c1054), .Z(n3164) );
XOR U5275 ( .A(c1055), .B(n3165), .Z(c1056) );
ANDN U5276 ( .B(n3166), .A(n3167), .Z(n3165) );
XOR U5277 ( .A(c1055), .B(b[1055]), .Z(n3166) );
XNOR U5278 ( .A(b[1055]), .B(n3167), .Z(c[1055]) );
XNOR U5279 ( .A(a[1055]), .B(c1055), .Z(n3167) );
XOR U5280 ( .A(c1056), .B(n3168), .Z(c1057) );
ANDN U5281 ( .B(n3169), .A(n3170), .Z(n3168) );
XOR U5282 ( .A(c1056), .B(b[1056]), .Z(n3169) );
XNOR U5283 ( .A(b[1056]), .B(n3170), .Z(c[1056]) );
XNOR U5284 ( .A(a[1056]), .B(c1056), .Z(n3170) );
XOR U5285 ( .A(c1057), .B(n3171), .Z(c1058) );
ANDN U5286 ( .B(n3172), .A(n3173), .Z(n3171) );
XOR U5287 ( .A(c1057), .B(b[1057]), .Z(n3172) );
XNOR U5288 ( .A(b[1057]), .B(n3173), .Z(c[1057]) );
XNOR U5289 ( .A(a[1057]), .B(c1057), .Z(n3173) );
XOR U5290 ( .A(c1058), .B(n3174), .Z(c1059) );
ANDN U5291 ( .B(n3175), .A(n3176), .Z(n3174) );
XOR U5292 ( .A(c1058), .B(b[1058]), .Z(n3175) );
XNOR U5293 ( .A(b[1058]), .B(n3176), .Z(c[1058]) );
XNOR U5294 ( .A(a[1058]), .B(c1058), .Z(n3176) );
XOR U5295 ( .A(c1059), .B(n3177), .Z(c1060) );
ANDN U5296 ( .B(n3178), .A(n3179), .Z(n3177) );
XOR U5297 ( .A(c1059), .B(b[1059]), .Z(n3178) );
XNOR U5298 ( .A(b[1059]), .B(n3179), .Z(c[1059]) );
XNOR U5299 ( .A(a[1059]), .B(c1059), .Z(n3179) );
XOR U5300 ( .A(c1060), .B(n3180), .Z(c1061) );
ANDN U5301 ( .B(n3181), .A(n3182), .Z(n3180) );
XOR U5302 ( .A(c1060), .B(b[1060]), .Z(n3181) );
XNOR U5303 ( .A(b[1060]), .B(n3182), .Z(c[1060]) );
XNOR U5304 ( .A(a[1060]), .B(c1060), .Z(n3182) );
XOR U5305 ( .A(c1061), .B(n3183), .Z(c1062) );
ANDN U5306 ( .B(n3184), .A(n3185), .Z(n3183) );
XOR U5307 ( .A(c1061), .B(b[1061]), .Z(n3184) );
XNOR U5308 ( .A(b[1061]), .B(n3185), .Z(c[1061]) );
XNOR U5309 ( .A(a[1061]), .B(c1061), .Z(n3185) );
XOR U5310 ( .A(c1062), .B(n3186), .Z(c1063) );
ANDN U5311 ( .B(n3187), .A(n3188), .Z(n3186) );
XOR U5312 ( .A(c1062), .B(b[1062]), .Z(n3187) );
XNOR U5313 ( .A(b[1062]), .B(n3188), .Z(c[1062]) );
XNOR U5314 ( .A(a[1062]), .B(c1062), .Z(n3188) );
XOR U5315 ( .A(c1063), .B(n3189), .Z(c1064) );
ANDN U5316 ( .B(n3190), .A(n3191), .Z(n3189) );
XOR U5317 ( .A(c1063), .B(b[1063]), .Z(n3190) );
XNOR U5318 ( .A(b[1063]), .B(n3191), .Z(c[1063]) );
XNOR U5319 ( .A(a[1063]), .B(c1063), .Z(n3191) );
XOR U5320 ( .A(c1064), .B(n3192), .Z(c1065) );
ANDN U5321 ( .B(n3193), .A(n3194), .Z(n3192) );
XOR U5322 ( .A(c1064), .B(b[1064]), .Z(n3193) );
XNOR U5323 ( .A(b[1064]), .B(n3194), .Z(c[1064]) );
XNOR U5324 ( .A(a[1064]), .B(c1064), .Z(n3194) );
XOR U5325 ( .A(c1065), .B(n3195), .Z(c1066) );
ANDN U5326 ( .B(n3196), .A(n3197), .Z(n3195) );
XOR U5327 ( .A(c1065), .B(b[1065]), .Z(n3196) );
XNOR U5328 ( .A(b[1065]), .B(n3197), .Z(c[1065]) );
XNOR U5329 ( .A(a[1065]), .B(c1065), .Z(n3197) );
XOR U5330 ( .A(c1066), .B(n3198), .Z(c1067) );
ANDN U5331 ( .B(n3199), .A(n3200), .Z(n3198) );
XOR U5332 ( .A(c1066), .B(b[1066]), .Z(n3199) );
XNOR U5333 ( .A(b[1066]), .B(n3200), .Z(c[1066]) );
XNOR U5334 ( .A(a[1066]), .B(c1066), .Z(n3200) );
XOR U5335 ( .A(c1067), .B(n3201), .Z(c1068) );
ANDN U5336 ( .B(n3202), .A(n3203), .Z(n3201) );
XOR U5337 ( .A(c1067), .B(b[1067]), .Z(n3202) );
XNOR U5338 ( .A(b[1067]), .B(n3203), .Z(c[1067]) );
XNOR U5339 ( .A(a[1067]), .B(c1067), .Z(n3203) );
XOR U5340 ( .A(c1068), .B(n3204), .Z(c1069) );
ANDN U5341 ( .B(n3205), .A(n3206), .Z(n3204) );
XOR U5342 ( .A(c1068), .B(b[1068]), .Z(n3205) );
XNOR U5343 ( .A(b[1068]), .B(n3206), .Z(c[1068]) );
XNOR U5344 ( .A(a[1068]), .B(c1068), .Z(n3206) );
XOR U5345 ( .A(c1069), .B(n3207), .Z(c1070) );
ANDN U5346 ( .B(n3208), .A(n3209), .Z(n3207) );
XOR U5347 ( .A(c1069), .B(b[1069]), .Z(n3208) );
XNOR U5348 ( .A(b[1069]), .B(n3209), .Z(c[1069]) );
XNOR U5349 ( .A(a[1069]), .B(c1069), .Z(n3209) );
XOR U5350 ( .A(c1070), .B(n3210), .Z(c1071) );
ANDN U5351 ( .B(n3211), .A(n3212), .Z(n3210) );
XOR U5352 ( .A(c1070), .B(b[1070]), .Z(n3211) );
XNOR U5353 ( .A(b[1070]), .B(n3212), .Z(c[1070]) );
XNOR U5354 ( .A(a[1070]), .B(c1070), .Z(n3212) );
XOR U5355 ( .A(c1071), .B(n3213), .Z(c1072) );
ANDN U5356 ( .B(n3214), .A(n3215), .Z(n3213) );
XOR U5357 ( .A(c1071), .B(b[1071]), .Z(n3214) );
XNOR U5358 ( .A(b[1071]), .B(n3215), .Z(c[1071]) );
XNOR U5359 ( .A(a[1071]), .B(c1071), .Z(n3215) );
XOR U5360 ( .A(c1072), .B(n3216), .Z(c1073) );
ANDN U5361 ( .B(n3217), .A(n3218), .Z(n3216) );
XOR U5362 ( .A(c1072), .B(b[1072]), .Z(n3217) );
XNOR U5363 ( .A(b[1072]), .B(n3218), .Z(c[1072]) );
XNOR U5364 ( .A(a[1072]), .B(c1072), .Z(n3218) );
XOR U5365 ( .A(c1073), .B(n3219), .Z(c1074) );
ANDN U5366 ( .B(n3220), .A(n3221), .Z(n3219) );
XOR U5367 ( .A(c1073), .B(b[1073]), .Z(n3220) );
XNOR U5368 ( .A(b[1073]), .B(n3221), .Z(c[1073]) );
XNOR U5369 ( .A(a[1073]), .B(c1073), .Z(n3221) );
XOR U5370 ( .A(c1074), .B(n3222), .Z(c1075) );
ANDN U5371 ( .B(n3223), .A(n3224), .Z(n3222) );
XOR U5372 ( .A(c1074), .B(b[1074]), .Z(n3223) );
XNOR U5373 ( .A(b[1074]), .B(n3224), .Z(c[1074]) );
XNOR U5374 ( .A(a[1074]), .B(c1074), .Z(n3224) );
XOR U5375 ( .A(c1075), .B(n3225), .Z(c1076) );
ANDN U5376 ( .B(n3226), .A(n3227), .Z(n3225) );
XOR U5377 ( .A(c1075), .B(b[1075]), .Z(n3226) );
XNOR U5378 ( .A(b[1075]), .B(n3227), .Z(c[1075]) );
XNOR U5379 ( .A(a[1075]), .B(c1075), .Z(n3227) );
XOR U5380 ( .A(c1076), .B(n3228), .Z(c1077) );
ANDN U5381 ( .B(n3229), .A(n3230), .Z(n3228) );
XOR U5382 ( .A(c1076), .B(b[1076]), .Z(n3229) );
XNOR U5383 ( .A(b[1076]), .B(n3230), .Z(c[1076]) );
XNOR U5384 ( .A(a[1076]), .B(c1076), .Z(n3230) );
XOR U5385 ( .A(c1077), .B(n3231), .Z(c1078) );
ANDN U5386 ( .B(n3232), .A(n3233), .Z(n3231) );
XOR U5387 ( .A(c1077), .B(b[1077]), .Z(n3232) );
XNOR U5388 ( .A(b[1077]), .B(n3233), .Z(c[1077]) );
XNOR U5389 ( .A(a[1077]), .B(c1077), .Z(n3233) );
XOR U5390 ( .A(c1078), .B(n3234), .Z(c1079) );
ANDN U5391 ( .B(n3235), .A(n3236), .Z(n3234) );
XOR U5392 ( .A(c1078), .B(b[1078]), .Z(n3235) );
XNOR U5393 ( .A(b[1078]), .B(n3236), .Z(c[1078]) );
XNOR U5394 ( .A(a[1078]), .B(c1078), .Z(n3236) );
XOR U5395 ( .A(c1079), .B(n3237), .Z(c1080) );
ANDN U5396 ( .B(n3238), .A(n3239), .Z(n3237) );
XOR U5397 ( .A(c1079), .B(b[1079]), .Z(n3238) );
XNOR U5398 ( .A(b[1079]), .B(n3239), .Z(c[1079]) );
XNOR U5399 ( .A(a[1079]), .B(c1079), .Z(n3239) );
XOR U5400 ( .A(c1080), .B(n3240), .Z(c1081) );
ANDN U5401 ( .B(n3241), .A(n3242), .Z(n3240) );
XOR U5402 ( .A(c1080), .B(b[1080]), .Z(n3241) );
XNOR U5403 ( .A(b[1080]), .B(n3242), .Z(c[1080]) );
XNOR U5404 ( .A(a[1080]), .B(c1080), .Z(n3242) );
XOR U5405 ( .A(c1081), .B(n3243), .Z(c1082) );
ANDN U5406 ( .B(n3244), .A(n3245), .Z(n3243) );
XOR U5407 ( .A(c1081), .B(b[1081]), .Z(n3244) );
XNOR U5408 ( .A(b[1081]), .B(n3245), .Z(c[1081]) );
XNOR U5409 ( .A(a[1081]), .B(c1081), .Z(n3245) );
XOR U5410 ( .A(c1082), .B(n3246), .Z(c1083) );
ANDN U5411 ( .B(n3247), .A(n3248), .Z(n3246) );
XOR U5412 ( .A(c1082), .B(b[1082]), .Z(n3247) );
XNOR U5413 ( .A(b[1082]), .B(n3248), .Z(c[1082]) );
XNOR U5414 ( .A(a[1082]), .B(c1082), .Z(n3248) );
XOR U5415 ( .A(c1083), .B(n3249), .Z(c1084) );
ANDN U5416 ( .B(n3250), .A(n3251), .Z(n3249) );
XOR U5417 ( .A(c1083), .B(b[1083]), .Z(n3250) );
XNOR U5418 ( .A(b[1083]), .B(n3251), .Z(c[1083]) );
XNOR U5419 ( .A(a[1083]), .B(c1083), .Z(n3251) );
XOR U5420 ( .A(c1084), .B(n3252), .Z(c1085) );
ANDN U5421 ( .B(n3253), .A(n3254), .Z(n3252) );
XOR U5422 ( .A(c1084), .B(b[1084]), .Z(n3253) );
XNOR U5423 ( .A(b[1084]), .B(n3254), .Z(c[1084]) );
XNOR U5424 ( .A(a[1084]), .B(c1084), .Z(n3254) );
XOR U5425 ( .A(c1085), .B(n3255), .Z(c1086) );
ANDN U5426 ( .B(n3256), .A(n3257), .Z(n3255) );
XOR U5427 ( .A(c1085), .B(b[1085]), .Z(n3256) );
XNOR U5428 ( .A(b[1085]), .B(n3257), .Z(c[1085]) );
XNOR U5429 ( .A(a[1085]), .B(c1085), .Z(n3257) );
XOR U5430 ( .A(c1086), .B(n3258), .Z(c1087) );
ANDN U5431 ( .B(n3259), .A(n3260), .Z(n3258) );
XOR U5432 ( .A(c1086), .B(b[1086]), .Z(n3259) );
XNOR U5433 ( .A(b[1086]), .B(n3260), .Z(c[1086]) );
XNOR U5434 ( .A(a[1086]), .B(c1086), .Z(n3260) );
XOR U5435 ( .A(c1087), .B(n3261), .Z(c1088) );
ANDN U5436 ( .B(n3262), .A(n3263), .Z(n3261) );
XOR U5437 ( .A(c1087), .B(b[1087]), .Z(n3262) );
XNOR U5438 ( .A(b[1087]), .B(n3263), .Z(c[1087]) );
XNOR U5439 ( .A(a[1087]), .B(c1087), .Z(n3263) );
XOR U5440 ( .A(c1088), .B(n3264), .Z(c1089) );
ANDN U5441 ( .B(n3265), .A(n3266), .Z(n3264) );
XOR U5442 ( .A(c1088), .B(b[1088]), .Z(n3265) );
XNOR U5443 ( .A(b[1088]), .B(n3266), .Z(c[1088]) );
XNOR U5444 ( .A(a[1088]), .B(c1088), .Z(n3266) );
XOR U5445 ( .A(c1089), .B(n3267), .Z(c1090) );
ANDN U5446 ( .B(n3268), .A(n3269), .Z(n3267) );
XOR U5447 ( .A(c1089), .B(b[1089]), .Z(n3268) );
XNOR U5448 ( .A(b[1089]), .B(n3269), .Z(c[1089]) );
XNOR U5449 ( .A(a[1089]), .B(c1089), .Z(n3269) );
XOR U5450 ( .A(c1090), .B(n3270), .Z(c1091) );
ANDN U5451 ( .B(n3271), .A(n3272), .Z(n3270) );
XOR U5452 ( .A(c1090), .B(b[1090]), .Z(n3271) );
XNOR U5453 ( .A(b[1090]), .B(n3272), .Z(c[1090]) );
XNOR U5454 ( .A(a[1090]), .B(c1090), .Z(n3272) );
XOR U5455 ( .A(c1091), .B(n3273), .Z(c1092) );
ANDN U5456 ( .B(n3274), .A(n3275), .Z(n3273) );
XOR U5457 ( .A(c1091), .B(b[1091]), .Z(n3274) );
XNOR U5458 ( .A(b[1091]), .B(n3275), .Z(c[1091]) );
XNOR U5459 ( .A(a[1091]), .B(c1091), .Z(n3275) );
XOR U5460 ( .A(c1092), .B(n3276), .Z(c1093) );
ANDN U5461 ( .B(n3277), .A(n3278), .Z(n3276) );
XOR U5462 ( .A(c1092), .B(b[1092]), .Z(n3277) );
XNOR U5463 ( .A(b[1092]), .B(n3278), .Z(c[1092]) );
XNOR U5464 ( .A(a[1092]), .B(c1092), .Z(n3278) );
XOR U5465 ( .A(c1093), .B(n3279), .Z(c1094) );
ANDN U5466 ( .B(n3280), .A(n3281), .Z(n3279) );
XOR U5467 ( .A(c1093), .B(b[1093]), .Z(n3280) );
XNOR U5468 ( .A(b[1093]), .B(n3281), .Z(c[1093]) );
XNOR U5469 ( .A(a[1093]), .B(c1093), .Z(n3281) );
XOR U5470 ( .A(c1094), .B(n3282), .Z(c1095) );
ANDN U5471 ( .B(n3283), .A(n3284), .Z(n3282) );
XOR U5472 ( .A(c1094), .B(b[1094]), .Z(n3283) );
XNOR U5473 ( .A(b[1094]), .B(n3284), .Z(c[1094]) );
XNOR U5474 ( .A(a[1094]), .B(c1094), .Z(n3284) );
XOR U5475 ( .A(c1095), .B(n3285), .Z(c1096) );
ANDN U5476 ( .B(n3286), .A(n3287), .Z(n3285) );
XOR U5477 ( .A(c1095), .B(b[1095]), .Z(n3286) );
XNOR U5478 ( .A(b[1095]), .B(n3287), .Z(c[1095]) );
XNOR U5479 ( .A(a[1095]), .B(c1095), .Z(n3287) );
XOR U5480 ( .A(c1096), .B(n3288), .Z(c1097) );
ANDN U5481 ( .B(n3289), .A(n3290), .Z(n3288) );
XOR U5482 ( .A(c1096), .B(b[1096]), .Z(n3289) );
XNOR U5483 ( .A(b[1096]), .B(n3290), .Z(c[1096]) );
XNOR U5484 ( .A(a[1096]), .B(c1096), .Z(n3290) );
XOR U5485 ( .A(c1097), .B(n3291), .Z(c1098) );
ANDN U5486 ( .B(n3292), .A(n3293), .Z(n3291) );
XOR U5487 ( .A(c1097), .B(b[1097]), .Z(n3292) );
XNOR U5488 ( .A(b[1097]), .B(n3293), .Z(c[1097]) );
XNOR U5489 ( .A(a[1097]), .B(c1097), .Z(n3293) );
XOR U5490 ( .A(c1098), .B(n3294), .Z(c1099) );
ANDN U5491 ( .B(n3295), .A(n3296), .Z(n3294) );
XOR U5492 ( .A(c1098), .B(b[1098]), .Z(n3295) );
XNOR U5493 ( .A(b[1098]), .B(n3296), .Z(c[1098]) );
XNOR U5494 ( .A(a[1098]), .B(c1098), .Z(n3296) );
XOR U5495 ( .A(c1099), .B(n3297), .Z(c1100) );
ANDN U5496 ( .B(n3298), .A(n3299), .Z(n3297) );
XOR U5497 ( .A(c1099), .B(b[1099]), .Z(n3298) );
XNOR U5498 ( .A(b[1099]), .B(n3299), .Z(c[1099]) );
XNOR U5499 ( .A(a[1099]), .B(c1099), .Z(n3299) );
XOR U5500 ( .A(c1100), .B(n3300), .Z(c1101) );
ANDN U5501 ( .B(n3301), .A(n3302), .Z(n3300) );
XOR U5502 ( .A(c1100), .B(b[1100]), .Z(n3301) );
XNOR U5503 ( .A(b[1100]), .B(n3302), .Z(c[1100]) );
XNOR U5504 ( .A(a[1100]), .B(c1100), .Z(n3302) );
XOR U5505 ( .A(c1101), .B(n3303), .Z(c1102) );
ANDN U5506 ( .B(n3304), .A(n3305), .Z(n3303) );
XOR U5507 ( .A(c1101), .B(b[1101]), .Z(n3304) );
XNOR U5508 ( .A(b[1101]), .B(n3305), .Z(c[1101]) );
XNOR U5509 ( .A(a[1101]), .B(c1101), .Z(n3305) );
XOR U5510 ( .A(c1102), .B(n3306), .Z(c1103) );
ANDN U5511 ( .B(n3307), .A(n3308), .Z(n3306) );
XOR U5512 ( .A(c1102), .B(b[1102]), .Z(n3307) );
XNOR U5513 ( .A(b[1102]), .B(n3308), .Z(c[1102]) );
XNOR U5514 ( .A(a[1102]), .B(c1102), .Z(n3308) );
XOR U5515 ( .A(c1103), .B(n3309), .Z(c1104) );
ANDN U5516 ( .B(n3310), .A(n3311), .Z(n3309) );
XOR U5517 ( .A(c1103), .B(b[1103]), .Z(n3310) );
XNOR U5518 ( .A(b[1103]), .B(n3311), .Z(c[1103]) );
XNOR U5519 ( .A(a[1103]), .B(c1103), .Z(n3311) );
XOR U5520 ( .A(c1104), .B(n3312), .Z(c1105) );
ANDN U5521 ( .B(n3313), .A(n3314), .Z(n3312) );
XOR U5522 ( .A(c1104), .B(b[1104]), .Z(n3313) );
XNOR U5523 ( .A(b[1104]), .B(n3314), .Z(c[1104]) );
XNOR U5524 ( .A(a[1104]), .B(c1104), .Z(n3314) );
XOR U5525 ( .A(c1105), .B(n3315), .Z(c1106) );
ANDN U5526 ( .B(n3316), .A(n3317), .Z(n3315) );
XOR U5527 ( .A(c1105), .B(b[1105]), .Z(n3316) );
XNOR U5528 ( .A(b[1105]), .B(n3317), .Z(c[1105]) );
XNOR U5529 ( .A(a[1105]), .B(c1105), .Z(n3317) );
XOR U5530 ( .A(c1106), .B(n3318), .Z(c1107) );
ANDN U5531 ( .B(n3319), .A(n3320), .Z(n3318) );
XOR U5532 ( .A(c1106), .B(b[1106]), .Z(n3319) );
XNOR U5533 ( .A(b[1106]), .B(n3320), .Z(c[1106]) );
XNOR U5534 ( .A(a[1106]), .B(c1106), .Z(n3320) );
XOR U5535 ( .A(c1107), .B(n3321), .Z(c1108) );
ANDN U5536 ( .B(n3322), .A(n3323), .Z(n3321) );
XOR U5537 ( .A(c1107), .B(b[1107]), .Z(n3322) );
XNOR U5538 ( .A(b[1107]), .B(n3323), .Z(c[1107]) );
XNOR U5539 ( .A(a[1107]), .B(c1107), .Z(n3323) );
XOR U5540 ( .A(c1108), .B(n3324), .Z(c1109) );
ANDN U5541 ( .B(n3325), .A(n3326), .Z(n3324) );
XOR U5542 ( .A(c1108), .B(b[1108]), .Z(n3325) );
XNOR U5543 ( .A(b[1108]), .B(n3326), .Z(c[1108]) );
XNOR U5544 ( .A(a[1108]), .B(c1108), .Z(n3326) );
XOR U5545 ( .A(c1109), .B(n3327), .Z(c1110) );
ANDN U5546 ( .B(n3328), .A(n3329), .Z(n3327) );
XOR U5547 ( .A(c1109), .B(b[1109]), .Z(n3328) );
XNOR U5548 ( .A(b[1109]), .B(n3329), .Z(c[1109]) );
XNOR U5549 ( .A(a[1109]), .B(c1109), .Z(n3329) );
XOR U5550 ( .A(c1110), .B(n3330), .Z(c1111) );
ANDN U5551 ( .B(n3331), .A(n3332), .Z(n3330) );
XOR U5552 ( .A(c1110), .B(b[1110]), .Z(n3331) );
XNOR U5553 ( .A(b[1110]), .B(n3332), .Z(c[1110]) );
XNOR U5554 ( .A(a[1110]), .B(c1110), .Z(n3332) );
XOR U5555 ( .A(c1111), .B(n3333), .Z(c1112) );
ANDN U5556 ( .B(n3334), .A(n3335), .Z(n3333) );
XOR U5557 ( .A(c1111), .B(b[1111]), .Z(n3334) );
XNOR U5558 ( .A(b[1111]), .B(n3335), .Z(c[1111]) );
XNOR U5559 ( .A(a[1111]), .B(c1111), .Z(n3335) );
XOR U5560 ( .A(c1112), .B(n3336), .Z(c1113) );
ANDN U5561 ( .B(n3337), .A(n3338), .Z(n3336) );
XOR U5562 ( .A(c1112), .B(b[1112]), .Z(n3337) );
XNOR U5563 ( .A(b[1112]), .B(n3338), .Z(c[1112]) );
XNOR U5564 ( .A(a[1112]), .B(c1112), .Z(n3338) );
XOR U5565 ( .A(c1113), .B(n3339), .Z(c1114) );
ANDN U5566 ( .B(n3340), .A(n3341), .Z(n3339) );
XOR U5567 ( .A(c1113), .B(b[1113]), .Z(n3340) );
XNOR U5568 ( .A(b[1113]), .B(n3341), .Z(c[1113]) );
XNOR U5569 ( .A(a[1113]), .B(c1113), .Z(n3341) );
XOR U5570 ( .A(c1114), .B(n3342), .Z(c1115) );
ANDN U5571 ( .B(n3343), .A(n3344), .Z(n3342) );
XOR U5572 ( .A(c1114), .B(b[1114]), .Z(n3343) );
XNOR U5573 ( .A(b[1114]), .B(n3344), .Z(c[1114]) );
XNOR U5574 ( .A(a[1114]), .B(c1114), .Z(n3344) );
XOR U5575 ( .A(c1115), .B(n3345), .Z(c1116) );
ANDN U5576 ( .B(n3346), .A(n3347), .Z(n3345) );
XOR U5577 ( .A(c1115), .B(b[1115]), .Z(n3346) );
XNOR U5578 ( .A(b[1115]), .B(n3347), .Z(c[1115]) );
XNOR U5579 ( .A(a[1115]), .B(c1115), .Z(n3347) );
XOR U5580 ( .A(c1116), .B(n3348), .Z(c1117) );
ANDN U5581 ( .B(n3349), .A(n3350), .Z(n3348) );
XOR U5582 ( .A(c1116), .B(b[1116]), .Z(n3349) );
XNOR U5583 ( .A(b[1116]), .B(n3350), .Z(c[1116]) );
XNOR U5584 ( .A(a[1116]), .B(c1116), .Z(n3350) );
XOR U5585 ( .A(c1117), .B(n3351), .Z(c1118) );
ANDN U5586 ( .B(n3352), .A(n3353), .Z(n3351) );
XOR U5587 ( .A(c1117), .B(b[1117]), .Z(n3352) );
XNOR U5588 ( .A(b[1117]), .B(n3353), .Z(c[1117]) );
XNOR U5589 ( .A(a[1117]), .B(c1117), .Z(n3353) );
XOR U5590 ( .A(c1118), .B(n3354), .Z(c1119) );
ANDN U5591 ( .B(n3355), .A(n3356), .Z(n3354) );
XOR U5592 ( .A(c1118), .B(b[1118]), .Z(n3355) );
XNOR U5593 ( .A(b[1118]), .B(n3356), .Z(c[1118]) );
XNOR U5594 ( .A(a[1118]), .B(c1118), .Z(n3356) );
XOR U5595 ( .A(c1119), .B(n3357), .Z(c1120) );
ANDN U5596 ( .B(n3358), .A(n3359), .Z(n3357) );
XOR U5597 ( .A(c1119), .B(b[1119]), .Z(n3358) );
XNOR U5598 ( .A(b[1119]), .B(n3359), .Z(c[1119]) );
XNOR U5599 ( .A(a[1119]), .B(c1119), .Z(n3359) );
XOR U5600 ( .A(c1120), .B(n3360), .Z(c1121) );
ANDN U5601 ( .B(n3361), .A(n3362), .Z(n3360) );
XOR U5602 ( .A(c1120), .B(b[1120]), .Z(n3361) );
XNOR U5603 ( .A(b[1120]), .B(n3362), .Z(c[1120]) );
XNOR U5604 ( .A(a[1120]), .B(c1120), .Z(n3362) );
XOR U5605 ( .A(c1121), .B(n3363), .Z(c1122) );
ANDN U5606 ( .B(n3364), .A(n3365), .Z(n3363) );
XOR U5607 ( .A(c1121), .B(b[1121]), .Z(n3364) );
XNOR U5608 ( .A(b[1121]), .B(n3365), .Z(c[1121]) );
XNOR U5609 ( .A(a[1121]), .B(c1121), .Z(n3365) );
XOR U5610 ( .A(c1122), .B(n3366), .Z(c1123) );
ANDN U5611 ( .B(n3367), .A(n3368), .Z(n3366) );
XOR U5612 ( .A(c1122), .B(b[1122]), .Z(n3367) );
XNOR U5613 ( .A(b[1122]), .B(n3368), .Z(c[1122]) );
XNOR U5614 ( .A(a[1122]), .B(c1122), .Z(n3368) );
XOR U5615 ( .A(c1123), .B(n3369), .Z(c1124) );
ANDN U5616 ( .B(n3370), .A(n3371), .Z(n3369) );
XOR U5617 ( .A(c1123), .B(b[1123]), .Z(n3370) );
XNOR U5618 ( .A(b[1123]), .B(n3371), .Z(c[1123]) );
XNOR U5619 ( .A(a[1123]), .B(c1123), .Z(n3371) );
XOR U5620 ( .A(c1124), .B(n3372), .Z(c1125) );
ANDN U5621 ( .B(n3373), .A(n3374), .Z(n3372) );
XOR U5622 ( .A(c1124), .B(b[1124]), .Z(n3373) );
XNOR U5623 ( .A(b[1124]), .B(n3374), .Z(c[1124]) );
XNOR U5624 ( .A(a[1124]), .B(c1124), .Z(n3374) );
XOR U5625 ( .A(c1125), .B(n3375), .Z(c1126) );
ANDN U5626 ( .B(n3376), .A(n3377), .Z(n3375) );
XOR U5627 ( .A(c1125), .B(b[1125]), .Z(n3376) );
XNOR U5628 ( .A(b[1125]), .B(n3377), .Z(c[1125]) );
XNOR U5629 ( .A(a[1125]), .B(c1125), .Z(n3377) );
XOR U5630 ( .A(c1126), .B(n3378), .Z(c1127) );
ANDN U5631 ( .B(n3379), .A(n3380), .Z(n3378) );
XOR U5632 ( .A(c1126), .B(b[1126]), .Z(n3379) );
XNOR U5633 ( .A(b[1126]), .B(n3380), .Z(c[1126]) );
XNOR U5634 ( .A(a[1126]), .B(c1126), .Z(n3380) );
XOR U5635 ( .A(c1127), .B(n3381), .Z(c1128) );
ANDN U5636 ( .B(n3382), .A(n3383), .Z(n3381) );
XOR U5637 ( .A(c1127), .B(b[1127]), .Z(n3382) );
XNOR U5638 ( .A(b[1127]), .B(n3383), .Z(c[1127]) );
XNOR U5639 ( .A(a[1127]), .B(c1127), .Z(n3383) );
XOR U5640 ( .A(c1128), .B(n3384), .Z(c1129) );
ANDN U5641 ( .B(n3385), .A(n3386), .Z(n3384) );
XOR U5642 ( .A(c1128), .B(b[1128]), .Z(n3385) );
XNOR U5643 ( .A(b[1128]), .B(n3386), .Z(c[1128]) );
XNOR U5644 ( .A(a[1128]), .B(c1128), .Z(n3386) );
XOR U5645 ( .A(c1129), .B(n3387), .Z(c1130) );
ANDN U5646 ( .B(n3388), .A(n3389), .Z(n3387) );
XOR U5647 ( .A(c1129), .B(b[1129]), .Z(n3388) );
XNOR U5648 ( .A(b[1129]), .B(n3389), .Z(c[1129]) );
XNOR U5649 ( .A(a[1129]), .B(c1129), .Z(n3389) );
XOR U5650 ( .A(c1130), .B(n3390), .Z(c1131) );
ANDN U5651 ( .B(n3391), .A(n3392), .Z(n3390) );
XOR U5652 ( .A(c1130), .B(b[1130]), .Z(n3391) );
XNOR U5653 ( .A(b[1130]), .B(n3392), .Z(c[1130]) );
XNOR U5654 ( .A(a[1130]), .B(c1130), .Z(n3392) );
XOR U5655 ( .A(c1131), .B(n3393), .Z(c1132) );
ANDN U5656 ( .B(n3394), .A(n3395), .Z(n3393) );
XOR U5657 ( .A(c1131), .B(b[1131]), .Z(n3394) );
XNOR U5658 ( .A(b[1131]), .B(n3395), .Z(c[1131]) );
XNOR U5659 ( .A(a[1131]), .B(c1131), .Z(n3395) );
XOR U5660 ( .A(c1132), .B(n3396), .Z(c1133) );
ANDN U5661 ( .B(n3397), .A(n3398), .Z(n3396) );
XOR U5662 ( .A(c1132), .B(b[1132]), .Z(n3397) );
XNOR U5663 ( .A(b[1132]), .B(n3398), .Z(c[1132]) );
XNOR U5664 ( .A(a[1132]), .B(c1132), .Z(n3398) );
XOR U5665 ( .A(c1133), .B(n3399), .Z(c1134) );
ANDN U5666 ( .B(n3400), .A(n3401), .Z(n3399) );
XOR U5667 ( .A(c1133), .B(b[1133]), .Z(n3400) );
XNOR U5668 ( .A(b[1133]), .B(n3401), .Z(c[1133]) );
XNOR U5669 ( .A(a[1133]), .B(c1133), .Z(n3401) );
XOR U5670 ( .A(c1134), .B(n3402), .Z(c1135) );
ANDN U5671 ( .B(n3403), .A(n3404), .Z(n3402) );
XOR U5672 ( .A(c1134), .B(b[1134]), .Z(n3403) );
XNOR U5673 ( .A(b[1134]), .B(n3404), .Z(c[1134]) );
XNOR U5674 ( .A(a[1134]), .B(c1134), .Z(n3404) );
XOR U5675 ( .A(c1135), .B(n3405), .Z(c1136) );
ANDN U5676 ( .B(n3406), .A(n3407), .Z(n3405) );
XOR U5677 ( .A(c1135), .B(b[1135]), .Z(n3406) );
XNOR U5678 ( .A(b[1135]), .B(n3407), .Z(c[1135]) );
XNOR U5679 ( .A(a[1135]), .B(c1135), .Z(n3407) );
XOR U5680 ( .A(c1136), .B(n3408), .Z(c1137) );
ANDN U5681 ( .B(n3409), .A(n3410), .Z(n3408) );
XOR U5682 ( .A(c1136), .B(b[1136]), .Z(n3409) );
XNOR U5683 ( .A(b[1136]), .B(n3410), .Z(c[1136]) );
XNOR U5684 ( .A(a[1136]), .B(c1136), .Z(n3410) );
XOR U5685 ( .A(c1137), .B(n3411), .Z(c1138) );
ANDN U5686 ( .B(n3412), .A(n3413), .Z(n3411) );
XOR U5687 ( .A(c1137), .B(b[1137]), .Z(n3412) );
XNOR U5688 ( .A(b[1137]), .B(n3413), .Z(c[1137]) );
XNOR U5689 ( .A(a[1137]), .B(c1137), .Z(n3413) );
XOR U5690 ( .A(c1138), .B(n3414), .Z(c1139) );
ANDN U5691 ( .B(n3415), .A(n3416), .Z(n3414) );
XOR U5692 ( .A(c1138), .B(b[1138]), .Z(n3415) );
XNOR U5693 ( .A(b[1138]), .B(n3416), .Z(c[1138]) );
XNOR U5694 ( .A(a[1138]), .B(c1138), .Z(n3416) );
XOR U5695 ( .A(c1139), .B(n3417), .Z(c1140) );
ANDN U5696 ( .B(n3418), .A(n3419), .Z(n3417) );
XOR U5697 ( .A(c1139), .B(b[1139]), .Z(n3418) );
XNOR U5698 ( .A(b[1139]), .B(n3419), .Z(c[1139]) );
XNOR U5699 ( .A(a[1139]), .B(c1139), .Z(n3419) );
XOR U5700 ( .A(c1140), .B(n3420), .Z(c1141) );
ANDN U5701 ( .B(n3421), .A(n3422), .Z(n3420) );
XOR U5702 ( .A(c1140), .B(b[1140]), .Z(n3421) );
XNOR U5703 ( .A(b[1140]), .B(n3422), .Z(c[1140]) );
XNOR U5704 ( .A(a[1140]), .B(c1140), .Z(n3422) );
XOR U5705 ( .A(c1141), .B(n3423), .Z(c1142) );
ANDN U5706 ( .B(n3424), .A(n3425), .Z(n3423) );
XOR U5707 ( .A(c1141), .B(b[1141]), .Z(n3424) );
XNOR U5708 ( .A(b[1141]), .B(n3425), .Z(c[1141]) );
XNOR U5709 ( .A(a[1141]), .B(c1141), .Z(n3425) );
XOR U5710 ( .A(c1142), .B(n3426), .Z(c1143) );
ANDN U5711 ( .B(n3427), .A(n3428), .Z(n3426) );
XOR U5712 ( .A(c1142), .B(b[1142]), .Z(n3427) );
XNOR U5713 ( .A(b[1142]), .B(n3428), .Z(c[1142]) );
XNOR U5714 ( .A(a[1142]), .B(c1142), .Z(n3428) );
XOR U5715 ( .A(c1143), .B(n3429), .Z(c1144) );
ANDN U5716 ( .B(n3430), .A(n3431), .Z(n3429) );
XOR U5717 ( .A(c1143), .B(b[1143]), .Z(n3430) );
XNOR U5718 ( .A(b[1143]), .B(n3431), .Z(c[1143]) );
XNOR U5719 ( .A(a[1143]), .B(c1143), .Z(n3431) );
XOR U5720 ( .A(c1144), .B(n3432), .Z(c1145) );
ANDN U5721 ( .B(n3433), .A(n3434), .Z(n3432) );
XOR U5722 ( .A(c1144), .B(b[1144]), .Z(n3433) );
XNOR U5723 ( .A(b[1144]), .B(n3434), .Z(c[1144]) );
XNOR U5724 ( .A(a[1144]), .B(c1144), .Z(n3434) );
XOR U5725 ( .A(c1145), .B(n3435), .Z(c1146) );
ANDN U5726 ( .B(n3436), .A(n3437), .Z(n3435) );
XOR U5727 ( .A(c1145), .B(b[1145]), .Z(n3436) );
XNOR U5728 ( .A(b[1145]), .B(n3437), .Z(c[1145]) );
XNOR U5729 ( .A(a[1145]), .B(c1145), .Z(n3437) );
XOR U5730 ( .A(c1146), .B(n3438), .Z(c1147) );
ANDN U5731 ( .B(n3439), .A(n3440), .Z(n3438) );
XOR U5732 ( .A(c1146), .B(b[1146]), .Z(n3439) );
XNOR U5733 ( .A(b[1146]), .B(n3440), .Z(c[1146]) );
XNOR U5734 ( .A(a[1146]), .B(c1146), .Z(n3440) );
XOR U5735 ( .A(c1147), .B(n3441), .Z(c1148) );
ANDN U5736 ( .B(n3442), .A(n3443), .Z(n3441) );
XOR U5737 ( .A(c1147), .B(b[1147]), .Z(n3442) );
XNOR U5738 ( .A(b[1147]), .B(n3443), .Z(c[1147]) );
XNOR U5739 ( .A(a[1147]), .B(c1147), .Z(n3443) );
XOR U5740 ( .A(c1148), .B(n3444), .Z(c1149) );
ANDN U5741 ( .B(n3445), .A(n3446), .Z(n3444) );
XOR U5742 ( .A(c1148), .B(b[1148]), .Z(n3445) );
XNOR U5743 ( .A(b[1148]), .B(n3446), .Z(c[1148]) );
XNOR U5744 ( .A(a[1148]), .B(c1148), .Z(n3446) );
XOR U5745 ( .A(c1149), .B(n3447), .Z(c1150) );
ANDN U5746 ( .B(n3448), .A(n3449), .Z(n3447) );
XOR U5747 ( .A(c1149), .B(b[1149]), .Z(n3448) );
XNOR U5748 ( .A(b[1149]), .B(n3449), .Z(c[1149]) );
XNOR U5749 ( .A(a[1149]), .B(c1149), .Z(n3449) );
XOR U5750 ( .A(c1150), .B(n3450), .Z(c1151) );
ANDN U5751 ( .B(n3451), .A(n3452), .Z(n3450) );
XOR U5752 ( .A(c1150), .B(b[1150]), .Z(n3451) );
XNOR U5753 ( .A(b[1150]), .B(n3452), .Z(c[1150]) );
XNOR U5754 ( .A(a[1150]), .B(c1150), .Z(n3452) );
XOR U5755 ( .A(c1151), .B(n3453), .Z(c1152) );
ANDN U5756 ( .B(n3454), .A(n3455), .Z(n3453) );
XOR U5757 ( .A(c1151), .B(b[1151]), .Z(n3454) );
XNOR U5758 ( .A(b[1151]), .B(n3455), .Z(c[1151]) );
XNOR U5759 ( .A(a[1151]), .B(c1151), .Z(n3455) );
XOR U5760 ( .A(c1152), .B(n3456), .Z(c1153) );
ANDN U5761 ( .B(n3457), .A(n3458), .Z(n3456) );
XOR U5762 ( .A(c1152), .B(b[1152]), .Z(n3457) );
XNOR U5763 ( .A(b[1152]), .B(n3458), .Z(c[1152]) );
XNOR U5764 ( .A(a[1152]), .B(c1152), .Z(n3458) );
XOR U5765 ( .A(c1153), .B(n3459), .Z(c1154) );
ANDN U5766 ( .B(n3460), .A(n3461), .Z(n3459) );
XOR U5767 ( .A(c1153), .B(b[1153]), .Z(n3460) );
XNOR U5768 ( .A(b[1153]), .B(n3461), .Z(c[1153]) );
XNOR U5769 ( .A(a[1153]), .B(c1153), .Z(n3461) );
XOR U5770 ( .A(c1154), .B(n3462), .Z(c1155) );
ANDN U5771 ( .B(n3463), .A(n3464), .Z(n3462) );
XOR U5772 ( .A(c1154), .B(b[1154]), .Z(n3463) );
XNOR U5773 ( .A(b[1154]), .B(n3464), .Z(c[1154]) );
XNOR U5774 ( .A(a[1154]), .B(c1154), .Z(n3464) );
XOR U5775 ( .A(c1155), .B(n3465), .Z(c1156) );
ANDN U5776 ( .B(n3466), .A(n3467), .Z(n3465) );
XOR U5777 ( .A(c1155), .B(b[1155]), .Z(n3466) );
XNOR U5778 ( .A(b[1155]), .B(n3467), .Z(c[1155]) );
XNOR U5779 ( .A(a[1155]), .B(c1155), .Z(n3467) );
XOR U5780 ( .A(c1156), .B(n3468), .Z(c1157) );
ANDN U5781 ( .B(n3469), .A(n3470), .Z(n3468) );
XOR U5782 ( .A(c1156), .B(b[1156]), .Z(n3469) );
XNOR U5783 ( .A(b[1156]), .B(n3470), .Z(c[1156]) );
XNOR U5784 ( .A(a[1156]), .B(c1156), .Z(n3470) );
XOR U5785 ( .A(c1157), .B(n3471), .Z(c1158) );
ANDN U5786 ( .B(n3472), .A(n3473), .Z(n3471) );
XOR U5787 ( .A(c1157), .B(b[1157]), .Z(n3472) );
XNOR U5788 ( .A(b[1157]), .B(n3473), .Z(c[1157]) );
XNOR U5789 ( .A(a[1157]), .B(c1157), .Z(n3473) );
XOR U5790 ( .A(c1158), .B(n3474), .Z(c1159) );
ANDN U5791 ( .B(n3475), .A(n3476), .Z(n3474) );
XOR U5792 ( .A(c1158), .B(b[1158]), .Z(n3475) );
XNOR U5793 ( .A(b[1158]), .B(n3476), .Z(c[1158]) );
XNOR U5794 ( .A(a[1158]), .B(c1158), .Z(n3476) );
XOR U5795 ( .A(c1159), .B(n3477), .Z(c1160) );
ANDN U5796 ( .B(n3478), .A(n3479), .Z(n3477) );
XOR U5797 ( .A(c1159), .B(b[1159]), .Z(n3478) );
XNOR U5798 ( .A(b[1159]), .B(n3479), .Z(c[1159]) );
XNOR U5799 ( .A(a[1159]), .B(c1159), .Z(n3479) );
XOR U5800 ( .A(c1160), .B(n3480), .Z(c1161) );
ANDN U5801 ( .B(n3481), .A(n3482), .Z(n3480) );
XOR U5802 ( .A(c1160), .B(b[1160]), .Z(n3481) );
XNOR U5803 ( .A(b[1160]), .B(n3482), .Z(c[1160]) );
XNOR U5804 ( .A(a[1160]), .B(c1160), .Z(n3482) );
XOR U5805 ( .A(c1161), .B(n3483), .Z(c1162) );
ANDN U5806 ( .B(n3484), .A(n3485), .Z(n3483) );
XOR U5807 ( .A(c1161), .B(b[1161]), .Z(n3484) );
XNOR U5808 ( .A(b[1161]), .B(n3485), .Z(c[1161]) );
XNOR U5809 ( .A(a[1161]), .B(c1161), .Z(n3485) );
XOR U5810 ( .A(c1162), .B(n3486), .Z(c1163) );
ANDN U5811 ( .B(n3487), .A(n3488), .Z(n3486) );
XOR U5812 ( .A(c1162), .B(b[1162]), .Z(n3487) );
XNOR U5813 ( .A(b[1162]), .B(n3488), .Z(c[1162]) );
XNOR U5814 ( .A(a[1162]), .B(c1162), .Z(n3488) );
XOR U5815 ( .A(c1163), .B(n3489), .Z(c1164) );
ANDN U5816 ( .B(n3490), .A(n3491), .Z(n3489) );
XOR U5817 ( .A(c1163), .B(b[1163]), .Z(n3490) );
XNOR U5818 ( .A(b[1163]), .B(n3491), .Z(c[1163]) );
XNOR U5819 ( .A(a[1163]), .B(c1163), .Z(n3491) );
XOR U5820 ( .A(c1164), .B(n3492), .Z(c1165) );
ANDN U5821 ( .B(n3493), .A(n3494), .Z(n3492) );
XOR U5822 ( .A(c1164), .B(b[1164]), .Z(n3493) );
XNOR U5823 ( .A(b[1164]), .B(n3494), .Z(c[1164]) );
XNOR U5824 ( .A(a[1164]), .B(c1164), .Z(n3494) );
XOR U5825 ( .A(c1165), .B(n3495), .Z(c1166) );
ANDN U5826 ( .B(n3496), .A(n3497), .Z(n3495) );
XOR U5827 ( .A(c1165), .B(b[1165]), .Z(n3496) );
XNOR U5828 ( .A(b[1165]), .B(n3497), .Z(c[1165]) );
XNOR U5829 ( .A(a[1165]), .B(c1165), .Z(n3497) );
XOR U5830 ( .A(c1166), .B(n3498), .Z(c1167) );
ANDN U5831 ( .B(n3499), .A(n3500), .Z(n3498) );
XOR U5832 ( .A(c1166), .B(b[1166]), .Z(n3499) );
XNOR U5833 ( .A(b[1166]), .B(n3500), .Z(c[1166]) );
XNOR U5834 ( .A(a[1166]), .B(c1166), .Z(n3500) );
XOR U5835 ( .A(c1167), .B(n3501), .Z(c1168) );
ANDN U5836 ( .B(n3502), .A(n3503), .Z(n3501) );
XOR U5837 ( .A(c1167), .B(b[1167]), .Z(n3502) );
XNOR U5838 ( .A(b[1167]), .B(n3503), .Z(c[1167]) );
XNOR U5839 ( .A(a[1167]), .B(c1167), .Z(n3503) );
XOR U5840 ( .A(c1168), .B(n3504), .Z(c1169) );
ANDN U5841 ( .B(n3505), .A(n3506), .Z(n3504) );
XOR U5842 ( .A(c1168), .B(b[1168]), .Z(n3505) );
XNOR U5843 ( .A(b[1168]), .B(n3506), .Z(c[1168]) );
XNOR U5844 ( .A(a[1168]), .B(c1168), .Z(n3506) );
XOR U5845 ( .A(c1169), .B(n3507), .Z(c1170) );
ANDN U5846 ( .B(n3508), .A(n3509), .Z(n3507) );
XOR U5847 ( .A(c1169), .B(b[1169]), .Z(n3508) );
XNOR U5848 ( .A(b[1169]), .B(n3509), .Z(c[1169]) );
XNOR U5849 ( .A(a[1169]), .B(c1169), .Z(n3509) );
XOR U5850 ( .A(c1170), .B(n3510), .Z(c1171) );
ANDN U5851 ( .B(n3511), .A(n3512), .Z(n3510) );
XOR U5852 ( .A(c1170), .B(b[1170]), .Z(n3511) );
XNOR U5853 ( .A(b[1170]), .B(n3512), .Z(c[1170]) );
XNOR U5854 ( .A(a[1170]), .B(c1170), .Z(n3512) );
XOR U5855 ( .A(c1171), .B(n3513), .Z(c1172) );
ANDN U5856 ( .B(n3514), .A(n3515), .Z(n3513) );
XOR U5857 ( .A(c1171), .B(b[1171]), .Z(n3514) );
XNOR U5858 ( .A(b[1171]), .B(n3515), .Z(c[1171]) );
XNOR U5859 ( .A(a[1171]), .B(c1171), .Z(n3515) );
XOR U5860 ( .A(c1172), .B(n3516), .Z(c1173) );
ANDN U5861 ( .B(n3517), .A(n3518), .Z(n3516) );
XOR U5862 ( .A(c1172), .B(b[1172]), .Z(n3517) );
XNOR U5863 ( .A(b[1172]), .B(n3518), .Z(c[1172]) );
XNOR U5864 ( .A(a[1172]), .B(c1172), .Z(n3518) );
XOR U5865 ( .A(c1173), .B(n3519), .Z(c1174) );
ANDN U5866 ( .B(n3520), .A(n3521), .Z(n3519) );
XOR U5867 ( .A(c1173), .B(b[1173]), .Z(n3520) );
XNOR U5868 ( .A(b[1173]), .B(n3521), .Z(c[1173]) );
XNOR U5869 ( .A(a[1173]), .B(c1173), .Z(n3521) );
XOR U5870 ( .A(c1174), .B(n3522), .Z(c1175) );
ANDN U5871 ( .B(n3523), .A(n3524), .Z(n3522) );
XOR U5872 ( .A(c1174), .B(b[1174]), .Z(n3523) );
XNOR U5873 ( .A(b[1174]), .B(n3524), .Z(c[1174]) );
XNOR U5874 ( .A(a[1174]), .B(c1174), .Z(n3524) );
XOR U5875 ( .A(c1175), .B(n3525), .Z(c1176) );
ANDN U5876 ( .B(n3526), .A(n3527), .Z(n3525) );
XOR U5877 ( .A(c1175), .B(b[1175]), .Z(n3526) );
XNOR U5878 ( .A(b[1175]), .B(n3527), .Z(c[1175]) );
XNOR U5879 ( .A(a[1175]), .B(c1175), .Z(n3527) );
XOR U5880 ( .A(c1176), .B(n3528), .Z(c1177) );
ANDN U5881 ( .B(n3529), .A(n3530), .Z(n3528) );
XOR U5882 ( .A(c1176), .B(b[1176]), .Z(n3529) );
XNOR U5883 ( .A(b[1176]), .B(n3530), .Z(c[1176]) );
XNOR U5884 ( .A(a[1176]), .B(c1176), .Z(n3530) );
XOR U5885 ( .A(c1177), .B(n3531), .Z(c1178) );
ANDN U5886 ( .B(n3532), .A(n3533), .Z(n3531) );
XOR U5887 ( .A(c1177), .B(b[1177]), .Z(n3532) );
XNOR U5888 ( .A(b[1177]), .B(n3533), .Z(c[1177]) );
XNOR U5889 ( .A(a[1177]), .B(c1177), .Z(n3533) );
XOR U5890 ( .A(c1178), .B(n3534), .Z(c1179) );
ANDN U5891 ( .B(n3535), .A(n3536), .Z(n3534) );
XOR U5892 ( .A(c1178), .B(b[1178]), .Z(n3535) );
XNOR U5893 ( .A(b[1178]), .B(n3536), .Z(c[1178]) );
XNOR U5894 ( .A(a[1178]), .B(c1178), .Z(n3536) );
XOR U5895 ( .A(c1179), .B(n3537), .Z(c1180) );
ANDN U5896 ( .B(n3538), .A(n3539), .Z(n3537) );
XOR U5897 ( .A(c1179), .B(b[1179]), .Z(n3538) );
XNOR U5898 ( .A(b[1179]), .B(n3539), .Z(c[1179]) );
XNOR U5899 ( .A(a[1179]), .B(c1179), .Z(n3539) );
XOR U5900 ( .A(c1180), .B(n3540), .Z(c1181) );
ANDN U5901 ( .B(n3541), .A(n3542), .Z(n3540) );
XOR U5902 ( .A(c1180), .B(b[1180]), .Z(n3541) );
XNOR U5903 ( .A(b[1180]), .B(n3542), .Z(c[1180]) );
XNOR U5904 ( .A(a[1180]), .B(c1180), .Z(n3542) );
XOR U5905 ( .A(c1181), .B(n3543), .Z(c1182) );
ANDN U5906 ( .B(n3544), .A(n3545), .Z(n3543) );
XOR U5907 ( .A(c1181), .B(b[1181]), .Z(n3544) );
XNOR U5908 ( .A(b[1181]), .B(n3545), .Z(c[1181]) );
XNOR U5909 ( .A(a[1181]), .B(c1181), .Z(n3545) );
XOR U5910 ( .A(c1182), .B(n3546), .Z(c1183) );
ANDN U5911 ( .B(n3547), .A(n3548), .Z(n3546) );
XOR U5912 ( .A(c1182), .B(b[1182]), .Z(n3547) );
XNOR U5913 ( .A(b[1182]), .B(n3548), .Z(c[1182]) );
XNOR U5914 ( .A(a[1182]), .B(c1182), .Z(n3548) );
XOR U5915 ( .A(c1183), .B(n3549), .Z(c1184) );
ANDN U5916 ( .B(n3550), .A(n3551), .Z(n3549) );
XOR U5917 ( .A(c1183), .B(b[1183]), .Z(n3550) );
XNOR U5918 ( .A(b[1183]), .B(n3551), .Z(c[1183]) );
XNOR U5919 ( .A(a[1183]), .B(c1183), .Z(n3551) );
XOR U5920 ( .A(c1184), .B(n3552), .Z(c1185) );
ANDN U5921 ( .B(n3553), .A(n3554), .Z(n3552) );
XOR U5922 ( .A(c1184), .B(b[1184]), .Z(n3553) );
XNOR U5923 ( .A(b[1184]), .B(n3554), .Z(c[1184]) );
XNOR U5924 ( .A(a[1184]), .B(c1184), .Z(n3554) );
XOR U5925 ( .A(c1185), .B(n3555), .Z(c1186) );
ANDN U5926 ( .B(n3556), .A(n3557), .Z(n3555) );
XOR U5927 ( .A(c1185), .B(b[1185]), .Z(n3556) );
XNOR U5928 ( .A(b[1185]), .B(n3557), .Z(c[1185]) );
XNOR U5929 ( .A(a[1185]), .B(c1185), .Z(n3557) );
XOR U5930 ( .A(c1186), .B(n3558), .Z(c1187) );
ANDN U5931 ( .B(n3559), .A(n3560), .Z(n3558) );
XOR U5932 ( .A(c1186), .B(b[1186]), .Z(n3559) );
XNOR U5933 ( .A(b[1186]), .B(n3560), .Z(c[1186]) );
XNOR U5934 ( .A(a[1186]), .B(c1186), .Z(n3560) );
XOR U5935 ( .A(c1187), .B(n3561), .Z(c1188) );
ANDN U5936 ( .B(n3562), .A(n3563), .Z(n3561) );
XOR U5937 ( .A(c1187), .B(b[1187]), .Z(n3562) );
XNOR U5938 ( .A(b[1187]), .B(n3563), .Z(c[1187]) );
XNOR U5939 ( .A(a[1187]), .B(c1187), .Z(n3563) );
XOR U5940 ( .A(c1188), .B(n3564), .Z(c1189) );
ANDN U5941 ( .B(n3565), .A(n3566), .Z(n3564) );
XOR U5942 ( .A(c1188), .B(b[1188]), .Z(n3565) );
XNOR U5943 ( .A(b[1188]), .B(n3566), .Z(c[1188]) );
XNOR U5944 ( .A(a[1188]), .B(c1188), .Z(n3566) );
XOR U5945 ( .A(c1189), .B(n3567), .Z(c1190) );
ANDN U5946 ( .B(n3568), .A(n3569), .Z(n3567) );
XOR U5947 ( .A(c1189), .B(b[1189]), .Z(n3568) );
XNOR U5948 ( .A(b[1189]), .B(n3569), .Z(c[1189]) );
XNOR U5949 ( .A(a[1189]), .B(c1189), .Z(n3569) );
XOR U5950 ( .A(c1190), .B(n3570), .Z(c1191) );
ANDN U5951 ( .B(n3571), .A(n3572), .Z(n3570) );
XOR U5952 ( .A(c1190), .B(b[1190]), .Z(n3571) );
XNOR U5953 ( .A(b[1190]), .B(n3572), .Z(c[1190]) );
XNOR U5954 ( .A(a[1190]), .B(c1190), .Z(n3572) );
XOR U5955 ( .A(c1191), .B(n3573), .Z(c1192) );
ANDN U5956 ( .B(n3574), .A(n3575), .Z(n3573) );
XOR U5957 ( .A(c1191), .B(b[1191]), .Z(n3574) );
XNOR U5958 ( .A(b[1191]), .B(n3575), .Z(c[1191]) );
XNOR U5959 ( .A(a[1191]), .B(c1191), .Z(n3575) );
XOR U5960 ( .A(c1192), .B(n3576), .Z(c1193) );
ANDN U5961 ( .B(n3577), .A(n3578), .Z(n3576) );
XOR U5962 ( .A(c1192), .B(b[1192]), .Z(n3577) );
XNOR U5963 ( .A(b[1192]), .B(n3578), .Z(c[1192]) );
XNOR U5964 ( .A(a[1192]), .B(c1192), .Z(n3578) );
XOR U5965 ( .A(c1193), .B(n3579), .Z(c1194) );
ANDN U5966 ( .B(n3580), .A(n3581), .Z(n3579) );
XOR U5967 ( .A(c1193), .B(b[1193]), .Z(n3580) );
XNOR U5968 ( .A(b[1193]), .B(n3581), .Z(c[1193]) );
XNOR U5969 ( .A(a[1193]), .B(c1193), .Z(n3581) );
XOR U5970 ( .A(c1194), .B(n3582), .Z(c1195) );
ANDN U5971 ( .B(n3583), .A(n3584), .Z(n3582) );
XOR U5972 ( .A(c1194), .B(b[1194]), .Z(n3583) );
XNOR U5973 ( .A(b[1194]), .B(n3584), .Z(c[1194]) );
XNOR U5974 ( .A(a[1194]), .B(c1194), .Z(n3584) );
XOR U5975 ( .A(c1195), .B(n3585), .Z(c1196) );
ANDN U5976 ( .B(n3586), .A(n3587), .Z(n3585) );
XOR U5977 ( .A(c1195), .B(b[1195]), .Z(n3586) );
XNOR U5978 ( .A(b[1195]), .B(n3587), .Z(c[1195]) );
XNOR U5979 ( .A(a[1195]), .B(c1195), .Z(n3587) );
XOR U5980 ( .A(c1196), .B(n3588), .Z(c1197) );
ANDN U5981 ( .B(n3589), .A(n3590), .Z(n3588) );
XOR U5982 ( .A(c1196), .B(b[1196]), .Z(n3589) );
XNOR U5983 ( .A(b[1196]), .B(n3590), .Z(c[1196]) );
XNOR U5984 ( .A(a[1196]), .B(c1196), .Z(n3590) );
XOR U5985 ( .A(c1197), .B(n3591), .Z(c1198) );
ANDN U5986 ( .B(n3592), .A(n3593), .Z(n3591) );
XOR U5987 ( .A(c1197), .B(b[1197]), .Z(n3592) );
XNOR U5988 ( .A(b[1197]), .B(n3593), .Z(c[1197]) );
XNOR U5989 ( .A(a[1197]), .B(c1197), .Z(n3593) );
XOR U5990 ( .A(c1198), .B(n3594), .Z(c1199) );
ANDN U5991 ( .B(n3595), .A(n3596), .Z(n3594) );
XOR U5992 ( .A(c1198), .B(b[1198]), .Z(n3595) );
XNOR U5993 ( .A(b[1198]), .B(n3596), .Z(c[1198]) );
XNOR U5994 ( .A(a[1198]), .B(c1198), .Z(n3596) );
XOR U5995 ( .A(c1199), .B(n3597), .Z(c1200) );
ANDN U5996 ( .B(n3598), .A(n3599), .Z(n3597) );
XOR U5997 ( .A(c1199), .B(b[1199]), .Z(n3598) );
XNOR U5998 ( .A(b[1199]), .B(n3599), .Z(c[1199]) );
XNOR U5999 ( .A(a[1199]), .B(c1199), .Z(n3599) );
XOR U6000 ( .A(c1200), .B(n3600), .Z(c1201) );
ANDN U6001 ( .B(n3601), .A(n3602), .Z(n3600) );
XOR U6002 ( .A(c1200), .B(b[1200]), .Z(n3601) );
XNOR U6003 ( .A(b[1200]), .B(n3602), .Z(c[1200]) );
XNOR U6004 ( .A(a[1200]), .B(c1200), .Z(n3602) );
XOR U6005 ( .A(c1201), .B(n3603), .Z(c1202) );
ANDN U6006 ( .B(n3604), .A(n3605), .Z(n3603) );
XOR U6007 ( .A(c1201), .B(b[1201]), .Z(n3604) );
XNOR U6008 ( .A(b[1201]), .B(n3605), .Z(c[1201]) );
XNOR U6009 ( .A(a[1201]), .B(c1201), .Z(n3605) );
XOR U6010 ( .A(c1202), .B(n3606), .Z(c1203) );
ANDN U6011 ( .B(n3607), .A(n3608), .Z(n3606) );
XOR U6012 ( .A(c1202), .B(b[1202]), .Z(n3607) );
XNOR U6013 ( .A(b[1202]), .B(n3608), .Z(c[1202]) );
XNOR U6014 ( .A(a[1202]), .B(c1202), .Z(n3608) );
XOR U6015 ( .A(c1203), .B(n3609), .Z(c1204) );
ANDN U6016 ( .B(n3610), .A(n3611), .Z(n3609) );
XOR U6017 ( .A(c1203), .B(b[1203]), .Z(n3610) );
XNOR U6018 ( .A(b[1203]), .B(n3611), .Z(c[1203]) );
XNOR U6019 ( .A(a[1203]), .B(c1203), .Z(n3611) );
XOR U6020 ( .A(c1204), .B(n3612), .Z(c1205) );
ANDN U6021 ( .B(n3613), .A(n3614), .Z(n3612) );
XOR U6022 ( .A(c1204), .B(b[1204]), .Z(n3613) );
XNOR U6023 ( .A(b[1204]), .B(n3614), .Z(c[1204]) );
XNOR U6024 ( .A(a[1204]), .B(c1204), .Z(n3614) );
XOR U6025 ( .A(c1205), .B(n3615), .Z(c1206) );
ANDN U6026 ( .B(n3616), .A(n3617), .Z(n3615) );
XOR U6027 ( .A(c1205), .B(b[1205]), .Z(n3616) );
XNOR U6028 ( .A(b[1205]), .B(n3617), .Z(c[1205]) );
XNOR U6029 ( .A(a[1205]), .B(c1205), .Z(n3617) );
XOR U6030 ( .A(c1206), .B(n3618), .Z(c1207) );
ANDN U6031 ( .B(n3619), .A(n3620), .Z(n3618) );
XOR U6032 ( .A(c1206), .B(b[1206]), .Z(n3619) );
XNOR U6033 ( .A(b[1206]), .B(n3620), .Z(c[1206]) );
XNOR U6034 ( .A(a[1206]), .B(c1206), .Z(n3620) );
XOR U6035 ( .A(c1207), .B(n3621), .Z(c1208) );
ANDN U6036 ( .B(n3622), .A(n3623), .Z(n3621) );
XOR U6037 ( .A(c1207), .B(b[1207]), .Z(n3622) );
XNOR U6038 ( .A(b[1207]), .B(n3623), .Z(c[1207]) );
XNOR U6039 ( .A(a[1207]), .B(c1207), .Z(n3623) );
XOR U6040 ( .A(c1208), .B(n3624), .Z(c1209) );
ANDN U6041 ( .B(n3625), .A(n3626), .Z(n3624) );
XOR U6042 ( .A(c1208), .B(b[1208]), .Z(n3625) );
XNOR U6043 ( .A(b[1208]), .B(n3626), .Z(c[1208]) );
XNOR U6044 ( .A(a[1208]), .B(c1208), .Z(n3626) );
XOR U6045 ( .A(c1209), .B(n3627), .Z(c1210) );
ANDN U6046 ( .B(n3628), .A(n3629), .Z(n3627) );
XOR U6047 ( .A(c1209), .B(b[1209]), .Z(n3628) );
XNOR U6048 ( .A(b[1209]), .B(n3629), .Z(c[1209]) );
XNOR U6049 ( .A(a[1209]), .B(c1209), .Z(n3629) );
XOR U6050 ( .A(c1210), .B(n3630), .Z(c1211) );
ANDN U6051 ( .B(n3631), .A(n3632), .Z(n3630) );
XOR U6052 ( .A(c1210), .B(b[1210]), .Z(n3631) );
XNOR U6053 ( .A(b[1210]), .B(n3632), .Z(c[1210]) );
XNOR U6054 ( .A(a[1210]), .B(c1210), .Z(n3632) );
XOR U6055 ( .A(c1211), .B(n3633), .Z(c1212) );
ANDN U6056 ( .B(n3634), .A(n3635), .Z(n3633) );
XOR U6057 ( .A(c1211), .B(b[1211]), .Z(n3634) );
XNOR U6058 ( .A(b[1211]), .B(n3635), .Z(c[1211]) );
XNOR U6059 ( .A(a[1211]), .B(c1211), .Z(n3635) );
XOR U6060 ( .A(c1212), .B(n3636), .Z(c1213) );
ANDN U6061 ( .B(n3637), .A(n3638), .Z(n3636) );
XOR U6062 ( .A(c1212), .B(b[1212]), .Z(n3637) );
XNOR U6063 ( .A(b[1212]), .B(n3638), .Z(c[1212]) );
XNOR U6064 ( .A(a[1212]), .B(c1212), .Z(n3638) );
XOR U6065 ( .A(c1213), .B(n3639), .Z(c1214) );
ANDN U6066 ( .B(n3640), .A(n3641), .Z(n3639) );
XOR U6067 ( .A(c1213), .B(b[1213]), .Z(n3640) );
XNOR U6068 ( .A(b[1213]), .B(n3641), .Z(c[1213]) );
XNOR U6069 ( .A(a[1213]), .B(c1213), .Z(n3641) );
XOR U6070 ( .A(c1214), .B(n3642), .Z(c1215) );
ANDN U6071 ( .B(n3643), .A(n3644), .Z(n3642) );
XOR U6072 ( .A(c1214), .B(b[1214]), .Z(n3643) );
XNOR U6073 ( .A(b[1214]), .B(n3644), .Z(c[1214]) );
XNOR U6074 ( .A(a[1214]), .B(c1214), .Z(n3644) );
XOR U6075 ( .A(c1215), .B(n3645), .Z(c1216) );
ANDN U6076 ( .B(n3646), .A(n3647), .Z(n3645) );
XOR U6077 ( .A(c1215), .B(b[1215]), .Z(n3646) );
XNOR U6078 ( .A(b[1215]), .B(n3647), .Z(c[1215]) );
XNOR U6079 ( .A(a[1215]), .B(c1215), .Z(n3647) );
XOR U6080 ( .A(c1216), .B(n3648), .Z(c1217) );
ANDN U6081 ( .B(n3649), .A(n3650), .Z(n3648) );
XOR U6082 ( .A(c1216), .B(b[1216]), .Z(n3649) );
XNOR U6083 ( .A(b[1216]), .B(n3650), .Z(c[1216]) );
XNOR U6084 ( .A(a[1216]), .B(c1216), .Z(n3650) );
XOR U6085 ( .A(c1217), .B(n3651), .Z(c1218) );
ANDN U6086 ( .B(n3652), .A(n3653), .Z(n3651) );
XOR U6087 ( .A(c1217), .B(b[1217]), .Z(n3652) );
XNOR U6088 ( .A(b[1217]), .B(n3653), .Z(c[1217]) );
XNOR U6089 ( .A(a[1217]), .B(c1217), .Z(n3653) );
XOR U6090 ( .A(c1218), .B(n3654), .Z(c1219) );
ANDN U6091 ( .B(n3655), .A(n3656), .Z(n3654) );
XOR U6092 ( .A(c1218), .B(b[1218]), .Z(n3655) );
XNOR U6093 ( .A(b[1218]), .B(n3656), .Z(c[1218]) );
XNOR U6094 ( .A(a[1218]), .B(c1218), .Z(n3656) );
XOR U6095 ( .A(c1219), .B(n3657), .Z(c1220) );
ANDN U6096 ( .B(n3658), .A(n3659), .Z(n3657) );
XOR U6097 ( .A(c1219), .B(b[1219]), .Z(n3658) );
XNOR U6098 ( .A(b[1219]), .B(n3659), .Z(c[1219]) );
XNOR U6099 ( .A(a[1219]), .B(c1219), .Z(n3659) );
XOR U6100 ( .A(c1220), .B(n3660), .Z(c1221) );
ANDN U6101 ( .B(n3661), .A(n3662), .Z(n3660) );
XOR U6102 ( .A(c1220), .B(b[1220]), .Z(n3661) );
XNOR U6103 ( .A(b[1220]), .B(n3662), .Z(c[1220]) );
XNOR U6104 ( .A(a[1220]), .B(c1220), .Z(n3662) );
XOR U6105 ( .A(c1221), .B(n3663), .Z(c1222) );
ANDN U6106 ( .B(n3664), .A(n3665), .Z(n3663) );
XOR U6107 ( .A(c1221), .B(b[1221]), .Z(n3664) );
XNOR U6108 ( .A(b[1221]), .B(n3665), .Z(c[1221]) );
XNOR U6109 ( .A(a[1221]), .B(c1221), .Z(n3665) );
XOR U6110 ( .A(c1222), .B(n3666), .Z(c1223) );
ANDN U6111 ( .B(n3667), .A(n3668), .Z(n3666) );
XOR U6112 ( .A(c1222), .B(b[1222]), .Z(n3667) );
XNOR U6113 ( .A(b[1222]), .B(n3668), .Z(c[1222]) );
XNOR U6114 ( .A(a[1222]), .B(c1222), .Z(n3668) );
XOR U6115 ( .A(c1223), .B(n3669), .Z(c1224) );
ANDN U6116 ( .B(n3670), .A(n3671), .Z(n3669) );
XOR U6117 ( .A(c1223), .B(b[1223]), .Z(n3670) );
XNOR U6118 ( .A(b[1223]), .B(n3671), .Z(c[1223]) );
XNOR U6119 ( .A(a[1223]), .B(c1223), .Z(n3671) );
XOR U6120 ( .A(c1224), .B(n3672), .Z(c1225) );
ANDN U6121 ( .B(n3673), .A(n3674), .Z(n3672) );
XOR U6122 ( .A(c1224), .B(b[1224]), .Z(n3673) );
XNOR U6123 ( .A(b[1224]), .B(n3674), .Z(c[1224]) );
XNOR U6124 ( .A(a[1224]), .B(c1224), .Z(n3674) );
XOR U6125 ( .A(c1225), .B(n3675), .Z(c1226) );
ANDN U6126 ( .B(n3676), .A(n3677), .Z(n3675) );
XOR U6127 ( .A(c1225), .B(b[1225]), .Z(n3676) );
XNOR U6128 ( .A(b[1225]), .B(n3677), .Z(c[1225]) );
XNOR U6129 ( .A(a[1225]), .B(c1225), .Z(n3677) );
XOR U6130 ( .A(c1226), .B(n3678), .Z(c1227) );
ANDN U6131 ( .B(n3679), .A(n3680), .Z(n3678) );
XOR U6132 ( .A(c1226), .B(b[1226]), .Z(n3679) );
XNOR U6133 ( .A(b[1226]), .B(n3680), .Z(c[1226]) );
XNOR U6134 ( .A(a[1226]), .B(c1226), .Z(n3680) );
XOR U6135 ( .A(c1227), .B(n3681), .Z(c1228) );
ANDN U6136 ( .B(n3682), .A(n3683), .Z(n3681) );
XOR U6137 ( .A(c1227), .B(b[1227]), .Z(n3682) );
XNOR U6138 ( .A(b[1227]), .B(n3683), .Z(c[1227]) );
XNOR U6139 ( .A(a[1227]), .B(c1227), .Z(n3683) );
XOR U6140 ( .A(c1228), .B(n3684), .Z(c1229) );
ANDN U6141 ( .B(n3685), .A(n3686), .Z(n3684) );
XOR U6142 ( .A(c1228), .B(b[1228]), .Z(n3685) );
XNOR U6143 ( .A(b[1228]), .B(n3686), .Z(c[1228]) );
XNOR U6144 ( .A(a[1228]), .B(c1228), .Z(n3686) );
XOR U6145 ( .A(c1229), .B(n3687), .Z(c1230) );
ANDN U6146 ( .B(n3688), .A(n3689), .Z(n3687) );
XOR U6147 ( .A(c1229), .B(b[1229]), .Z(n3688) );
XNOR U6148 ( .A(b[1229]), .B(n3689), .Z(c[1229]) );
XNOR U6149 ( .A(a[1229]), .B(c1229), .Z(n3689) );
XOR U6150 ( .A(c1230), .B(n3690), .Z(c1231) );
ANDN U6151 ( .B(n3691), .A(n3692), .Z(n3690) );
XOR U6152 ( .A(c1230), .B(b[1230]), .Z(n3691) );
XNOR U6153 ( .A(b[1230]), .B(n3692), .Z(c[1230]) );
XNOR U6154 ( .A(a[1230]), .B(c1230), .Z(n3692) );
XOR U6155 ( .A(c1231), .B(n3693), .Z(c1232) );
ANDN U6156 ( .B(n3694), .A(n3695), .Z(n3693) );
XOR U6157 ( .A(c1231), .B(b[1231]), .Z(n3694) );
XNOR U6158 ( .A(b[1231]), .B(n3695), .Z(c[1231]) );
XNOR U6159 ( .A(a[1231]), .B(c1231), .Z(n3695) );
XOR U6160 ( .A(c1232), .B(n3696), .Z(c1233) );
ANDN U6161 ( .B(n3697), .A(n3698), .Z(n3696) );
XOR U6162 ( .A(c1232), .B(b[1232]), .Z(n3697) );
XNOR U6163 ( .A(b[1232]), .B(n3698), .Z(c[1232]) );
XNOR U6164 ( .A(a[1232]), .B(c1232), .Z(n3698) );
XOR U6165 ( .A(c1233), .B(n3699), .Z(c1234) );
ANDN U6166 ( .B(n3700), .A(n3701), .Z(n3699) );
XOR U6167 ( .A(c1233), .B(b[1233]), .Z(n3700) );
XNOR U6168 ( .A(b[1233]), .B(n3701), .Z(c[1233]) );
XNOR U6169 ( .A(a[1233]), .B(c1233), .Z(n3701) );
XOR U6170 ( .A(c1234), .B(n3702), .Z(c1235) );
ANDN U6171 ( .B(n3703), .A(n3704), .Z(n3702) );
XOR U6172 ( .A(c1234), .B(b[1234]), .Z(n3703) );
XNOR U6173 ( .A(b[1234]), .B(n3704), .Z(c[1234]) );
XNOR U6174 ( .A(a[1234]), .B(c1234), .Z(n3704) );
XOR U6175 ( .A(c1235), .B(n3705), .Z(c1236) );
ANDN U6176 ( .B(n3706), .A(n3707), .Z(n3705) );
XOR U6177 ( .A(c1235), .B(b[1235]), .Z(n3706) );
XNOR U6178 ( .A(b[1235]), .B(n3707), .Z(c[1235]) );
XNOR U6179 ( .A(a[1235]), .B(c1235), .Z(n3707) );
XOR U6180 ( .A(c1236), .B(n3708), .Z(c1237) );
ANDN U6181 ( .B(n3709), .A(n3710), .Z(n3708) );
XOR U6182 ( .A(c1236), .B(b[1236]), .Z(n3709) );
XNOR U6183 ( .A(b[1236]), .B(n3710), .Z(c[1236]) );
XNOR U6184 ( .A(a[1236]), .B(c1236), .Z(n3710) );
XOR U6185 ( .A(c1237), .B(n3711), .Z(c1238) );
ANDN U6186 ( .B(n3712), .A(n3713), .Z(n3711) );
XOR U6187 ( .A(c1237), .B(b[1237]), .Z(n3712) );
XNOR U6188 ( .A(b[1237]), .B(n3713), .Z(c[1237]) );
XNOR U6189 ( .A(a[1237]), .B(c1237), .Z(n3713) );
XOR U6190 ( .A(c1238), .B(n3714), .Z(c1239) );
ANDN U6191 ( .B(n3715), .A(n3716), .Z(n3714) );
XOR U6192 ( .A(c1238), .B(b[1238]), .Z(n3715) );
XNOR U6193 ( .A(b[1238]), .B(n3716), .Z(c[1238]) );
XNOR U6194 ( .A(a[1238]), .B(c1238), .Z(n3716) );
XOR U6195 ( .A(c1239), .B(n3717), .Z(c1240) );
ANDN U6196 ( .B(n3718), .A(n3719), .Z(n3717) );
XOR U6197 ( .A(c1239), .B(b[1239]), .Z(n3718) );
XNOR U6198 ( .A(b[1239]), .B(n3719), .Z(c[1239]) );
XNOR U6199 ( .A(a[1239]), .B(c1239), .Z(n3719) );
XOR U6200 ( .A(c1240), .B(n3720), .Z(c1241) );
ANDN U6201 ( .B(n3721), .A(n3722), .Z(n3720) );
XOR U6202 ( .A(c1240), .B(b[1240]), .Z(n3721) );
XNOR U6203 ( .A(b[1240]), .B(n3722), .Z(c[1240]) );
XNOR U6204 ( .A(a[1240]), .B(c1240), .Z(n3722) );
XOR U6205 ( .A(c1241), .B(n3723), .Z(c1242) );
ANDN U6206 ( .B(n3724), .A(n3725), .Z(n3723) );
XOR U6207 ( .A(c1241), .B(b[1241]), .Z(n3724) );
XNOR U6208 ( .A(b[1241]), .B(n3725), .Z(c[1241]) );
XNOR U6209 ( .A(a[1241]), .B(c1241), .Z(n3725) );
XOR U6210 ( .A(c1242), .B(n3726), .Z(c1243) );
ANDN U6211 ( .B(n3727), .A(n3728), .Z(n3726) );
XOR U6212 ( .A(c1242), .B(b[1242]), .Z(n3727) );
XNOR U6213 ( .A(b[1242]), .B(n3728), .Z(c[1242]) );
XNOR U6214 ( .A(a[1242]), .B(c1242), .Z(n3728) );
XOR U6215 ( .A(c1243), .B(n3729), .Z(c1244) );
ANDN U6216 ( .B(n3730), .A(n3731), .Z(n3729) );
XOR U6217 ( .A(c1243), .B(b[1243]), .Z(n3730) );
XNOR U6218 ( .A(b[1243]), .B(n3731), .Z(c[1243]) );
XNOR U6219 ( .A(a[1243]), .B(c1243), .Z(n3731) );
XOR U6220 ( .A(c1244), .B(n3732), .Z(c1245) );
ANDN U6221 ( .B(n3733), .A(n3734), .Z(n3732) );
XOR U6222 ( .A(c1244), .B(b[1244]), .Z(n3733) );
XNOR U6223 ( .A(b[1244]), .B(n3734), .Z(c[1244]) );
XNOR U6224 ( .A(a[1244]), .B(c1244), .Z(n3734) );
XOR U6225 ( .A(c1245), .B(n3735), .Z(c1246) );
ANDN U6226 ( .B(n3736), .A(n3737), .Z(n3735) );
XOR U6227 ( .A(c1245), .B(b[1245]), .Z(n3736) );
XNOR U6228 ( .A(b[1245]), .B(n3737), .Z(c[1245]) );
XNOR U6229 ( .A(a[1245]), .B(c1245), .Z(n3737) );
XOR U6230 ( .A(c1246), .B(n3738), .Z(c1247) );
ANDN U6231 ( .B(n3739), .A(n3740), .Z(n3738) );
XOR U6232 ( .A(c1246), .B(b[1246]), .Z(n3739) );
XNOR U6233 ( .A(b[1246]), .B(n3740), .Z(c[1246]) );
XNOR U6234 ( .A(a[1246]), .B(c1246), .Z(n3740) );
XOR U6235 ( .A(c1247), .B(n3741), .Z(c1248) );
ANDN U6236 ( .B(n3742), .A(n3743), .Z(n3741) );
XOR U6237 ( .A(c1247), .B(b[1247]), .Z(n3742) );
XNOR U6238 ( .A(b[1247]), .B(n3743), .Z(c[1247]) );
XNOR U6239 ( .A(a[1247]), .B(c1247), .Z(n3743) );
XOR U6240 ( .A(c1248), .B(n3744), .Z(c1249) );
ANDN U6241 ( .B(n3745), .A(n3746), .Z(n3744) );
XOR U6242 ( .A(c1248), .B(b[1248]), .Z(n3745) );
XNOR U6243 ( .A(b[1248]), .B(n3746), .Z(c[1248]) );
XNOR U6244 ( .A(a[1248]), .B(c1248), .Z(n3746) );
XOR U6245 ( .A(c1249), .B(n3747), .Z(c1250) );
ANDN U6246 ( .B(n3748), .A(n3749), .Z(n3747) );
XOR U6247 ( .A(c1249), .B(b[1249]), .Z(n3748) );
XNOR U6248 ( .A(b[1249]), .B(n3749), .Z(c[1249]) );
XNOR U6249 ( .A(a[1249]), .B(c1249), .Z(n3749) );
XOR U6250 ( .A(c1250), .B(n3750), .Z(c1251) );
ANDN U6251 ( .B(n3751), .A(n3752), .Z(n3750) );
XOR U6252 ( .A(c1250), .B(b[1250]), .Z(n3751) );
XNOR U6253 ( .A(b[1250]), .B(n3752), .Z(c[1250]) );
XNOR U6254 ( .A(a[1250]), .B(c1250), .Z(n3752) );
XOR U6255 ( .A(c1251), .B(n3753), .Z(c1252) );
ANDN U6256 ( .B(n3754), .A(n3755), .Z(n3753) );
XOR U6257 ( .A(c1251), .B(b[1251]), .Z(n3754) );
XNOR U6258 ( .A(b[1251]), .B(n3755), .Z(c[1251]) );
XNOR U6259 ( .A(a[1251]), .B(c1251), .Z(n3755) );
XOR U6260 ( .A(c1252), .B(n3756), .Z(c1253) );
ANDN U6261 ( .B(n3757), .A(n3758), .Z(n3756) );
XOR U6262 ( .A(c1252), .B(b[1252]), .Z(n3757) );
XNOR U6263 ( .A(b[1252]), .B(n3758), .Z(c[1252]) );
XNOR U6264 ( .A(a[1252]), .B(c1252), .Z(n3758) );
XOR U6265 ( .A(c1253), .B(n3759), .Z(c1254) );
ANDN U6266 ( .B(n3760), .A(n3761), .Z(n3759) );
XOR U6267 ( .A(c1253), .B(b[1253]), .Z(n3760) );
XNOR U6268 ( .A(b[1253]), .B(n3761), .Z(c[1253]) );
XNOR U6269 ( .A(a[1253]), .B(c1253), .Z(n3761) );
XOR U6270 ( .A(c1254), .B(n3762), .Z(c1255) );
ANDN U6271 ( .B(n3763), .A(n3764), .Z(n3762) );
XOR U6272 ( .A(c1254), .B(b[1254]), .Z(n3763) );
XNOR U6273 ( .A(b[1254]), .B(n3764), .Z(c[1254]) );
XNOR U6274 ( .A(a[1254]), .B(c1254), .Z(n3764) );
XOR U6275 ( .A(c1255), .B(n3765), .Z(c1256) );
ANDN U6276 ( .B(n3766), .A(n3767), .Z(n3765) );
XOR U6277 ( .A(c1255), .B(b[1255]), .Z(n3766) );
XNOR U6278 ( .A(b[1255]), .B(n3767), .Z(c[1255]) );
XNOR U6279 ( .A(a[1255]), .B(c1255), .Z(n3767) );
XOR U6280 ( .A(c1256), .B(n3768), .Z(c1257) );
ANDN U6281 ( .B(n3769), .A(n3770), .Z(n3768) );
XOR U6282 ( .A(c1256), .B(b[1256]), .Z(n3769) );
XNOR U6283 ( .A(b[1256]), .B(n3770), .Z(c[1256]) );
XNOR U6284 ( .A(a[1256]), .B(c1256), .Z(n3770) );
XOR U6285 ( .A(c1257), .B(n3771), .Z(c1258) );
ANDN U6286 ( .B(n3772), .A(n3773), .Z(n3771) );
XOR U6287 ( .A(c1257), .B(b[1257]), .Z(n3772) );
XNOR U6288 ( .A(b[1257]), .B(n3773), .Z(c[1257]) );
XNOR U6289 ( .A(a[1257]), .B(c1257), .Z(n3773) );
XOR U6290 ( .A(c1258), .B(n3774), .Z(c1259) );
ANDN U6291 ( .B(n3775), .A(n3776), .Z(n3774) );
XOR U6292 ( .A(c1258), .B(b[1258]), .Z(n3775) );
XNOR U6293 ( .A(b[1258]), .B(n3776), .Z(c[1258]) );
XNOR U6294 ( .A(a[1258]), .B(c1258), .Z(n3776) );
XOR U6295 ( .A(c1259), .B(n3777), .Z(c1260) );
ANDN U6296 ( .B(n3778), .A(n3779), .Z(n3777) );
XOR U6297 ( .A(c1259), .B(b[1259]), .Z(n3778) );
XNOR U6298 ( .A(b[1259]), .B(n3779), .Z(c[1259]) );
XNOR U6299 ( .A(a[1259]), .B(c1259), .Z(n3779) );
XOR U6300 ( .A(c1260), .B(n3780), .Z(c1261) );
ANDN U6301 ( .B(n3781), .A(n3782), .Z(n3780) );
XOR U6302 ( .A(c1260), .B(b[1260]), .Z(n3781) );
XNOR U6303 ( .A(b[1260]), .B(n3782), .Z(c[1260]) );
XNOR U6304 ( .A(a[1260]), .B(c1260), .Z(n3782) );
XOR U6305 ( .A(c1261), .B(n3783), .Z(c1262) );
ANDN U6306 ( .B(n3784), .A(n3785), .Z(n3783) );
XOR U6307 ( .A(c1261), .B(b[1261]), .Z(n3784) );
XNOR U6308 ( .A(b[1261]), .B(n3785), .Z(c[1261]) );
XNOR U6309 ( .A(a[1261]), .B(c1261), .Z(n3785) );
XOR U6310 ( .A(c1262), .B(n3786), .Z(c1263) );
ANDN U6311 ( .B(n3787), .A(n3788), .Z(n3786) );
XOR U6312 ( .A(c1262), .B(b[1262]), .Z(n3787) );
XNOR U6313 ( .A(b[1262]), .B(n3788), .Z(c[1262]) );
XNOR U6314 ( .A(a[1262]), .B(c1262), .Z(n3788) );
XOR U6315 ( .A(c1263), .B(n3789), .Z(c1264) );
ANDN U6316 ( .B(n3790), .A(n3791), .Z(n3789) );
XOR U6317 ( .A(c1263), .B(b[1263]), .Z(n3790) );
XNOR U6318 ( .A(b[1263]), .B(n3791), .Z(c[1263]) );
XNOR U6319 ( .A(a[1263]), .B(c1263), .Z(n3791) );
XOR U6320 ( .A(c1264), .B(n3792), .Z(c1265) );
ANDN U6321 ( .B(n3793), .A(n3794), .Z(n3792) );
XOR U6322 ( .A(c1264), .B(b[1264]), .Z(n3793) );
XNOR U6323 ( .A(b[1264]), .B(n3794), .Z(c[1264]) );
XNOR U6324 ( .A(a[1264]), .B(c1264), .Z(n3794) );
XOR U6325 ( .A(c1265), .B(n3795), .Z(c1266) );
ANDN U6326 ( .B(n3796), .A(n3797), .Z(n3795) );
XOR U6327 ( .A(c1265), .B(b[1265]), .Z(n3796) );
XNOR U6328 ( .A(b[1265]), .B(n3797), .Z(c[1265]) );
XNOR U6329 ( .A(a[1265]), .B(c1265), .Z(n3797) );
XOR U6330 ( .A(c1266), .B(n3798), .Z(c1267) );
ANDN U6331 ( .B(n3799), .A(n3800), .Z(n3798) );
XOR U6332 ( .A(c1266), .B(b[1266]), .Z(n3799) );
XNOR U6333 ( .A(b[1266]), .B(n3800), .Z(c[1266]) );
XNOR U6334 ( .A(a[1266]), .B(c1266), .Z(n3800) );
XOR U6335 ( .A(c1267), .B(n3801), .Z(c1268) );
ANDN U6336 ( .B(n3802), .A(n3803), .Z(n3801) );
XOR U6337 ( .A(c1267), .B(b[1267]), .Z(n3802) );
XNOR U6338 ( .A(b[1267]), .B(n3803), .Z(c[1267]) );
XNOR U6339 ( .A(a[1267]), .B(c1267), .Z(n3803) );
XOR U6340 ( .A(c1268), .B(n3804), .Z(c1269) );
ANDN U6341 ( .B(n3805), .A(n3806), .Z(n3804) );
XOR U6342 ( .A(c1268), .B(b[1268]), .Z(n3805) );
XNOR U6343 ( .A(b[1268]), .B(n3806), .Z(c[1268]) );
XNOR U6344 ( .A(a[1268]), .B(c1268), .Z(n3806) );
XOR U6345 ( .A(c1269), .B(n3807), .Z(c1270) );
ANDN U6346 ( .B(n3808), .A(n3809), .Z(n3807) );
XOR U6347 ( .A(c1269), .B(b[1269]), .Z(n3808) );
XNOR U6348 ( .A(b[1269]), .B(n3809), .Z(c[1269]) );
XNOR U6349 ( .A(a[1269]), .B(c1269), .Z(n3809) );
XOR U6350 ( .A(c1270), .B(n3810), .Z(c1271) );
ANDN U6351 ( .B(n3811), .A(n3812), .Z(n3810) );
XOR U6352 ( .A(c1270), .B(b[1270]), .Z(n3811) );
XNOR U6353 ( .A(b[1270]), .B(n3812), .Z(c[1270]) );
XNOR U6354 ( .A(a[1270]), .B(c1270), .Z(n3812) );
XOR U6355 ( .A(c1271), .B(n3813), .Z(c1272) );
ANDN U6356 ( .B(n3814), .A(n3815), .Z(n3813) );
XOR U6357 ( .A(c1271), .B(b[1271]), .Z(n3814) );
XNOR U6358 ( .A(b[1271]), .B(n3815), .Z(c[1271]) );
XNOR U6359 ( .A(a[1271]), .B(c1271), .Z(n3815) );
XOR U6360 ( .A(c1272), .B(n3816), .Z(c1273) );
ANDN U6361 ( .B(n3817), .A(n3818), .Z(n3816) );
XOR U6362 ( .A(c1272), .B(b[1272]), .Z(n3817) );
XNOR U6363 ( .A(b[1272]), .B(n3818), .Z(c[1272]) );
XNOR U6364 ( .A(a[1272]), .B(c1272), .Z(n3818) );
XOR U6365 ( .A(c1273), .B(n3819), .Z(c1274) );
ANDN U6366 ( .B(n3820), .A(n3821), .Z(n3819) );
XOR U6367 ( .A(c1273), .B(b[1273]), .Z(n3820) );
XNOR U6368 ( .A(b[1273]), .B(n3821), .Z(c[1273]) );
XNOR U6369 ( .A(a[1273]), .B(c1273), .Z(n3821) );
XOR U6370 ( .A(c1274), .B(n3822), .Z(c1275) );
ANDN U6371 ( .B(n3823), .A(n3824), .Z(n3822) );
XOR U6372 ( .A(c1274), .B(b[1274]), .Z(n3823) );
XNOR U6373 ( .A(b[1274]), .B(n3824), .Z(c[1274]) );
XNOR U6374 ( .A(a[1274]), .B(c1274), .Z(n3824) );
XOR U6375 ( .A(c1275), .B(n3825), .Z(c1276) );
ANDN U6376 ( .B(n3826), .A(n3827), .Z(n3825) );
XOR U6377 ( .A(c1275), .B(b[1275]), .Z(n3826) );
XNOR U6378 ( .A(b[1275]), .B(n3827), .Z(c[1275]) );
XNOR U6379 ( .A(a[1275]), .B(c1275), .Z(n3827) );
XOR U6380 ( .A(c1276), .B(n3828), .Z(c1277) );
ANDN U6381 ( .B(n3829), .A(n3830), .Z(n3828) );
XOR U6382 ( .A(c1276), .B(b[1276]), .Z(n3829) );
XNOR U6383 ( .A(b[1276]), .B(n3830), .Z(c[1276]) );
XNOR U6384 ( .A(a[1276]), .B(c1276), .Z(n3830) );
XOR U6385 ( .A(c1277), .B(n3831), .Z(c1278) );
ANDN U6386 ( .B(n3832), .A(n3833), .Z(n3831) );
XOR U6387 ( .A(c1277), .B(b[1277]), .Z(n3832) );
XNOR U6388 ( .A(b[1277]), .B(n3833), .Z(c[1277]) );
XNOR U6389 ( .A(a[1277]), .B(c1277), .Z(n3833) );
XOR U6390 ( .A(c1278), .B(n3834), .Z(c1279) );
ANDN U6391 ( .B(n3835), .A(n3836), .Z(n3834) );
XOR U6392 ( .A(c1278), .B(b[1278]), .Z(n3835) );
XNOR U6393 ( .A(b[1278]), .B(n3836), .Z(c[1278]) );
XNOR U6394 ( .A(a[1278]), .B(c1278), .Z(n3836) );
XOR U6395 ( .A(c1279), .B(n3837), .Z(c1280) );
ANDN U6396 ( .B(n3838), .A(n3839), .Z(n3837) );
XOR U6397 ( .A(c1279), .B(b[1279]), .Z(n3838) );
XNOR U6398 ( .A(b[1279]), .B(n3839), .Z(c[1279]) );
XNOR U6399 ( .A(a[1279]), .B(c1279), .Z(n3839) );
XOR U6400 ( .A(c1280), .B(n3840), .Z(c1281) );
ANDN U6401 ( .B(n3841), .A(n3842), .Z(n3840) );
XOR U6402 ( .A(c1280), .B(b[1280]), .Z(n3841) );
XNOR U6403 ( .A(b[1280]), .B(n3842), .Z(c[1280]) );
XNOR U6404 ( .A(a[1280]), .B(c1280), .Z(n3842) );
XOR U6405 ( .A(c1281), .B(n3843), .Z(c1282) );
ANDN U6406 ( .B(n3844), .A(n3845), .Z(n3843) );
XOR U6407 ( .A(c1281), .B(b[1281]), .Z(n3844) );
XNOR U6408 ( .A(b[1281]), .B(n3845), .Z(c[1281]) );
XNOR U6409 ( .A(a[1281]), .B(c1281), .Z(n3845) );
XOR U6410 ( .A(c1282), .B(n3846), .Z(c1283) );
ANDN U6411 ( .B(n3847), .A(n3848), .Z(n3846) );
XOR U6412 ( .A(c1282), .B(b[1282]), .Z(n3847) );
XNOR U6413 ( .A(b[1282]), .B(n3848), .Z(c[1282]) );
XNOR U6414 ( .A(a[1282]), .B(c1282), .Z(n3848) );
XOR U6415 ( .A(c1283), .B(n3849), .Z(c1284) );
ANDN U6416 ( .B(n3850), .A(n3851), .Z(n3849) );
XOR U6417 ( .A(c1283), .B(b[1283]), .Z(n3850) );
XNOR U6418 ( .A(b[1283]), .B(n3851), .Z(c[1283]) );
XNOR U6419 ( .A(a[1283]), .B(c1283), .Z(n3851) );
XOR U6420 ( .A(c1284), .B(n3852), .Z(c1285) );
ANDN U6421 ( .B(n3853), .A(n3854), .Z(n3852) );
XOR U6422 ( .A(c1284), .B(b[1284]), .Z(n3853) );
XNOR U6423 ( .A(b[1284]), .B(n3854), .Z(c[1284]) );
XNOR U6424 ( .A(a[1284]), .B(c1284), .Z(n3854) );
XOR U6425 ( .A(c1285), .B(n3855), .Z(c1286) );
ANDN U6426 ( .B(n3856), .A(n3857), .Z(n3855) );
XOR U6427 ( .A(c1285), .B(b[1285]), .Z(n3856) );
XNOR U6428 ( .A(b[1285]), .B(n3857), .Z(c[1285]) );
XNOR U6429 ( .A(a[1285]), .B(c1285), .Z(n3857) );
XOR U6430 ( .A(c1286), .B(n3858), .Z(c1287) );
ANDN U6431 ( .B(n3859), .A(n3860), .Z(n3858) );
XOR U6432 ( .A(c1286), .B(b[1286]), .Z(n3859) );
XNOR U6433 ( .A(b[1286]), .B(n3860), .Z(c[1286]) );
XNOR U6434 ( .A(a[1286]), .B(c1286), .Z(n3860) );
XOR U6435 ( .A(c1287), .B(n3861), .Z(c1288) );
ANDN U6436 ( .B(n3862), .A(n3863), .Z(n3861) );
XOR U6437 ( .A(c1287), .B(b[1287]), .Z(n3862) );
XNOR U6438 ( .A(b[1287]), .B(n3863), .Z(c[1287]) );
XNOR U6439 ( .A(a[1287]), .B(c1287), .Z(n3863) );
XOR U6440 ( .A(c1288), .B(n3864), .Z(c1289) );
ANDN U6441 ( .B(n3865), .A(n3866), .Z(n3864) );
XOR U6442 ( .A(c1288), .B(b[1288]), .Z(n3865) );
XNOR U6443 ( .A(b[1288]), .B(n3866), .Z(c[1288]) );
XNOR U6444 ( .A(a[1288]), .B(c1288), .Z(n3866) );
XOR U6445 ( .A(c1289), .B(n3867), .Z(c1290) );
ANDN U6446 ( .B(n3868), .A(n3869), .Z(n3867) );
XOR U6447 ( .A(c1289), .B(b[1289]), .Z(n3868) );
XNOR U6448 ( .A(b[1289]), .B(n3869), .Z(c[1289]) );
XNOR U6449 ( .A(a[1289]), .B(c1289), .Z(n3869) );
XOR U6450 ( .A(c1290), .B(n3870), .Z(c1291) );
ANDN U6451 ( .B(n3871), .A(n3872), .Z(n3870) );
XOR U6452 ( .A(c1290), .B(b[1290]), .Z(n3871) );
XNOR U6453 ( .A(b[1290]), .B(n3872), .Z(c[1290]) );
XNOR U6454 ( .A(a[1290]), .B(c1290), .Z(n3872) );
XOR U6455 ( .A(c1291), .B(n3873), .Z(c1292) );
ANDN U6456 ( .B(n3874), .A(n3875), .Z(n3873) );
XOR U6457 ( .A(c1291), .B(b[1291]), .Z(n3874) );
XNOR U6458 ( .A(b[1291]), .B(n3875), .Z(c[1291]) );
XNOR U6459 ( .A(a[1291]), .B(c1291), .Z(n3875) );
XOR U6460 ( .A(c1292), .B(n3876), .Z(c1293) );
ANDN U6461 ( .B(n3877), .A(n3878), .Z(n3876) );
XOR U6462 ( .A(c1292), .B(b[1292]), .Z(n3877) );
XNOR U6463 ( .A(b[1292]), .B(n3878), .Z(c[1292]) );
XNOR U6464 ( .A(a[1292]), .B(c1292), .Z(n3878) );
XOR U6465 ( .A(c1293), .B(n3879), .Z(c1294) );
ANDN U6466 ( .B(n3880), .A(n3881), .Z(n3879) );
XOR U6467 ( .A(c1293), .B(b[1293]), .Z(n3880) );
XNOR U6468 ( .A(b[1293]), .B(n3881), .Z(c[1293]) );
XNOR U6469 ( .A(a[1293]), .B(c1293), .Z(n3881) );
XOR U6470 ( .A(c1294), .B(n3882), .Z(c1295) );
ANDN U6471 ( .B(n3883), .A(n3884), .Z(n3882) );
XOR U6472 ( .A(c1294), .B(b[1294]), .Z(n3883) );
XNOR U6473 ( .A(b[1294]), .B(n3884), .Z(c[1294]) );
XNOR U6474 ( .A(a[1294]), .B(c1294), .Z(n3884) );
XOR U6475 ( .A(c1295), .B(n3885), .Z(c1296) );
ANDN U6476 ( .B(n3886), .A(n3887), .Z(n3885) );
XOR U6477 ( .A(c1295), .B(b[1295]), .Z(n3886) );
XNOR U6478 ( .A(b[1295]), .B(n3887), .Z(c[1295]) );
XNOR U6479 ( .A(a[1295]), .B(c1295), .Z(n3887) );
XOR U6480 ( .A(c1296), .B(n3888), .Z(c1297) );
ANDN U6481 ( .B(n3889), .A(n3890), .Z(n3888) );
XOR U6482 ( .A(c1296), .B(b[1296]), .Z(n3889) );
XNOR U6483 ( .A(b[1296]), .B(n3890), .Z(c[1296]) );
XNOR U6484 ( .A(a[1296]), .B(c1296), .Z(n3890) );
XOR U6485 ( .A(c1297), .B(n3891), .Z(c1298) );
ANDN U6486 ( .B(n3892), .A(n3893), .Z(n3891) );
XOR U6487 ( .A(c1297), .B(b[1297]), .Z(n3892) );
XNOR U6488 ( .A(b[1297]), .B(n3893), .Z(c[1297]) );
XNOR U6489 ( .A(a[1297]), .B(c1297), .Z(n3893) );
XOR U6490 ( .A(c1298), .B(n3894), .Z(c1299) );
ANDN U6491 ( .B(n3895), .A(n3896), .Z(n3894) );
XOR U6492 ( .A(c1298), .B(b[1298]), .Z(n3895) );
XNOR U6493 ( .A(b[1298]), .B(n3896), .Z(c[1298]) );
XNOR U6494 ( .A(a[1298]), .B(c1298), .Z(n3896) );
XOR U6495 ( .A(c1299), .B(n3897), .Z(c1300) );
ANDN U6496 ( .B(n3898), .A(n3899), .Z(n3897) );
XOR U6497 ( .A(c1299), .B(b[1299]), .Z(n3898) );
XNOR U6498 ( .A(b[1299]), .B(n3899), .Z(c[1299]) );
XNOR U6499 ( .A(a[1299]), .B(c1299), .Z(n3899) );
XOR U6500 ( .A(c1300), .B(n3900), .Z(c1301) );
ANDN U6501 ( .B(n3901), .A(n3902), .Z(n3900) );
XOR U6502 ( .A(c1300), .B(b[1300]), .Z(n3901) );
XNOR U6503 ( .A(b[1300]), .B(n3902), .Z(c[1300]) );
XNOR U6504 ( .A(a[1300]), .B(c1300), .Z(n3902) );
XOR U6505 ( .A(c1301), .B(n3903), .Z(c1302) );
ANDN U6506 ( .B(n3904), .A(n3905), .Z(n3903) );
XOR U6507 ( .A(c1301), .B(b[1301]), .Z(n3904) );
XNOR U6508 ( .A(b[1301]), .B(n3905), .Z(c[1301]) );
XNOR U6509 ( .A(a[1301]), .B(c1301), .Z(n3905) );
XOR U6510 ( .A(c1302), .B(n3906), .Z(c1303) );
ANDN U6511 ( .B(n3907), .A(n3908), .Z(n3906) );
XOR U6512 ( .A(c1302), .B(b[1302]), .Z(n3907) );
XNOR U6513 ( .A(b[1302]), .B(n3908), .Z(c[1302]) );
XNOR U6514 ( .A(a[1302]), .B(c1302), .Z(n3908) );
XOR U6515 ( .A(c1303), .B(n3909), .Z(c1304) );
ANDN U6516 ( .B(n3910), .A(n3911), .Z(n3909) );
XOR U6517 ( .A(c1303), .B(b[1303]), .Z(n3910) );
XNOR U6518 ( .A(b[1303]), .B(n3911), .Z(c[1303]) );
XNOR U6519 ( .A(a[1303]), .B(c1303), .Z(n3911) );
XOR U6520 ( .A(c1304), .B(n3912), .Z(c1305) );
ANDN U6521 ( .B(n3913), .A(n3914), .Z(n3912) );
XOR U6522 ( .A(c1304), .B(b[1304]), .Z(n3913) );
XNOR U6523 ( .A(b[1304]), .B(n3914), .Z(c[1304]) );
XNOR U6524 ( .A(a[1304]), .B(c1304), .Z(n3914) );
XOR U6525 ( .A(c1305), .B(n3915), .Z(c1306) );
ANDN U6526 ( .B(n3916), .A(n3917), .Z(n3915) );
XOR U6527 ( .A(c1305), .B(b[1305]), .Z(n3916) );
XNOR U6528 ( .A(b[1305]), .B(n3917), .Z(c[1305]) );
XNOR U6529 ( .A(a[1305]), .B(c1305), .Z(n3917) );
XOR U6530 ( .A(c1306), .B(n3918), .Z(c1307) );
ANDN U6531 ( .B(n3919), .A(n3920), .Z(n3918) );
XOR U6532 ( .A(c1306), .B(b[1306]), .Z(n3919) );
XNOR U6533 ( .A(b[1306]), .B(n3920), .Z(c[1306]) );
XNOR U6534 ( .A(a[1306]), .B(c1306), .Z(n3920) );
XOR U6535 ( .A(c1307), .B(n3921), .Z(c1308) );
ANDN U6536 ( .B(n3922), .A(n3923), .Z(n3921) );
XOR U6537 ( .A(c1307), .B(b[1307]), .Z(n3922) );
XNOR U6538 ( .A(b[1307]), .B(n3923), .Z(c[1307]) );
XNOR U6539 ( .A(a[1307]), .B(c1307), .Z(n3923) );
XOR U6540 ( .A(c1308), .B(n3924), .Z(c1309) );
ANDN U6541 ( .B(n3925), .A(n3926), .Z(n3924) );
XOR U6542 ( .A(c1308), .B(b[1308]), .Z(n3925) );
XNOR U6543 ( .A(b[1308]), .B(n3926), .Z(c[1308]) );
XNOR U6544 ( .A(a[1308]), .B(c1308), .Z(n3926) );
XOR U6545 ( .A(c1309), .B(n3927), .Z(c1310) );
ANDN U6546 ( .B(n3928), .A(n3929), .Z(n3927) );
XOR U6547 ( .A(c1309), .B(b[1309]), .Z(n3928) );
XNOR U6548 ( .A(b[1309]), .B(n3929), .Z(c[1309]) );
XNOR U6549 ( .A(a[1309]), .B(c1309), .Z(n3929) );
XOR U6550 ( .A(c1310), .B(n3930), .Z(c1311) );
ANDN U6551 ( .B(n3931), .A(n3932), .Z(n3930) );
XOR U6552 ( .A(c1310), .B(b[1310]), .Z(n3931) );
XNOR U6553 ( .A(b[1310]), .B(n3932), .Z(c[1310]) );
XNOR U6554 ( .A(a[1310]), .B(c1310), .Z(n3932) );
XOR U6555 ( .A(c1311), .B(n3933), .Z(c1312) );
ANDN U6556 ( .B(n3934), .A(n3935), .Z(n3933) );
XOR U6557 ( .A(c1311), .B(b[1311]), .Z(n3934) );
XNOR U6558 ( .A(b[1311]), .B(n3935), .Z(c[1311]) );
XNOR U6559 ( .A(a[1311]), .B(c1311), .Z(n3935) );
XOR U6560 ( .A(c1312), .B(n3936), .Z(c1313) );
ANDN U6561 ( .B(n3937), .A(n3938), .Z(n3936) );
XOR U6562 ( .A(c1312), .B(b[1312]), .Z(n3937) );
XNOR U6563 ( .A(b[1312]), .B(n3938), .Z(c[1312]) );
XNOR U6564 ( .A(a[1312]), .B(c1312), .Z(n3938) );
XOR U6565 ( .A(c1313), .B(n3939), .Z(c1314) );
ANDN U6566 ( .B(n3940), .A(n3941), .Z(n3939) );
XOR U6567 ( .A(c1313), .B(b[1313]), .Z(n3940) );
XNOR U6568 ( .A(b[1313]), .B(n3941), .Z(c[1313]) );
XNOR U6569 ( .A(a[1313]), .B(c1313), .Z(n3941) );
XOR U6570 ( .A(c1314), .B(n3942), .Z(c1315) );
ANDN U6571 ( .B(n3943), .A(n3944), .Z(n3942) );
XOR U6572 ( .A(c1314), .B(b[1314]), .Z(n3943) );
XNOR U6573 ( .A(b[1314]), .B(n3944), .Z(c[1314]) );
XNOR U6574 ( .A(a[1314]), .B(c1314), .Z(n3944) );
XOR U6575 ( .A(c1315), .B(n3945), .Z(c1316) );
ANDN U6576 ( .B(n3946), .A(n3947), .Z(n3945) );
XOR U6577 ( .A(c1315), .B(b[1315]), .Z(n3946) );
XNOR U6578 ( .A(b[1315]), .B(n3947), .Z(c[1315]) );
XNOR U6579 ( .A(a[1315]), .B(c1315), .Z(n3947) );
XOR U6580 ( .A(c1316), .B(n3948), .Z(c1317) );
ANDN U6581 ( .B(n3949), .A(n3950), .Z(n3948) );
XOR U6582 ( .A(c1316), .B(b[1316]), .Z(n3949) );
XNOR U6583 ( .A(b[1316]), .B(n3950), .Z(c[1316]) );
XNOR U6584 ( .A(a[1316]), .B(c1316), .Z(n3950) );
XOR U6585 ( .A(c1317), .B(n3951), .Z(c1318) );
ANDN U6586 ( .B(n3952), .A(n3953), .Z(n3951) );
XOR U6587 ( .A(c1317), .B(b[1317]), .Z(n3952) );
XNOR U6588 ( .A(b[1317]), .B(n3953), .Z(c[1317]) );
XNOR U6589 ( .A(a[1317]), .B(c1317), .Z(n3953) );
XOR U6590 ( .A(c1318), .B(n3954), .Z(c1319) );
ANDN U6591 ( .B(n3955), .A(n3956), .Z(n3954) );
XOR U6592 ( .A(c1318), .B(b[1318]), .Z(n3955) );
XNOR U6593 ( .A(b[1318]), .B(n3956), .Z(c[1318]) );
XNOR U6594 ( .A(a[1318]), .B(c1318), .Z(n3956) );
XOR U6595 ( .A(c1319), .B(n3957), .Z(c1320) );
ANDN U6596 ( .B(n3958), .A(n3959), .Z(n3957) );
XOR U6597 ( .A(c1319), .B(b[1319]), .Z(n3958) );
XNOR U6598 ( .A(b[1319]), .B(n3959), .Z(c[1319]) );
XNOR U6599 ( .A(a[1319]), .B(c1319), .Z(n3959) );
XOR U6600 ( .A(c1320), .B(n3960), .Z(c1321) );
ANDN U6601 ( .B(n3961), .A(n3962), .Z(n3960) );
XOR U6602 ( .A(c1320), .B(b[1320]), .Z(n3961) );
XNOR U6603 ( .A(b[1320]), .B(n3962), .Z(c[1320]) );
XNOR U6604 ( .A(a[1320]), .B(c1320), .Z(n3962) );
XOR U6605 ( .A(c1321), .B(n3963), .Z(c1322) );
ANDN U6606 ( .B(n3964), .A(n3965), .Z(n3963) );
XOR U6607 ( .A(c1321), .B(b[1321]), .Z(n3964) );
XNOR U6608 ( .A(b[1321]), .B(n3965), .Z(c[1321]) );
XNOR U6609 ( .A(a[1321]), .B(c1321), .Z(n3965) );
XOR U6610 ( .A(c1322), .B(n3966), .Z(c1323) );
ANDN U6611 ( .B(n3967), .A(n3968), .Z(n3966) );
XOR U6612 ( .A(c1322), .B(b[1322]), .Z(n3967) );
XNOR U6613 ( .A(b[1322]), .B(n3968), .Z(c[1322]) );
XNOR U6614 ( .A(a[1322]), .B(c1322), .Z(n3968) );
XOR U6615 ( .A(c1323), .B(n3969), .Z(c1324) );
ANDN U6616 ( .B(n3970), .A(n3971), .Z(n3969) );
XOR U6617 ( .A(c1323), .B(b[1323]), .Z(n3970) );
XNOR U6618 ( .A(b[1323]), .B(n3971), .Z(c[1323]) );
XNOR U6619 ( .A(a[1323]), .B(c1323), .Z(n3971) );
XOR U6620 ( .A(c1324), .B(n3972), .Z(c1325) );
ANDN U6621 ( .B(n3973), .A(n3974), .Z(n3972) );
XOR U6622 ( .A(c1324), .B(b[1324]), .Z(n3973) );
XNOR U6623 ( .A(b[1324]), .B(n3974), .Z(c[1324]) );
XNOR U6624 ( .A(a[1324]), .B(c1324), .Z(n3974) );
XOR U6625 ( .A(c1325), .B(n3975), .Z(c1326) );
ANDN U6626 ( .B(n3976), .A(n3977), .Z(n3975) );
XOR U6627 ( .A(c1325), .B(b[1325]), .Z(n3976) );
XNOR U6628 ( .A(b[1325]), .B(n3977), .Z(c[1325]) );
XNOR U6629 ( .A(a[1325]), .B(c1325), .Z(n3977) );
XOR U6630 ( .A(c1326), .B(n3978), .Z(c1327) );
ANDN U6631 ( .B(n3979), .A(n3980), .Z(n3978) );
XOR U6632 ( .A(c1326), .B(b[1326]), .Z(n3979) );
XNOR U6633 ( .A(b[1326]), .B(n3980), .Z(c[1326]) );
XNOR U6634 ( .A(a[1326]), .B(c1326), .Z(n3980) );
XOR U6635 ( .A(c1327), .B(n3981), .Z(c1328) );
ANDN U6636 ( .B(n3982), .A(n3983), .Z(n3981) );
XOR U6637 ( .A(c1327), .B(b[1327]), .Z(n3982) );
XNOR U6638 ( .A(b[1327]), .B(n3983), .Z(c[1327]) );
XNOR U6639 ( .A(a[1327]), .B(c1327), .Z(n3983) );
XOR U6640 ( .A(c1328), .B(n3984), .Z(c1329) );
ANDN U6641 ( .B(n3985), .A(n3986), .Z(n3984) );
XOR U6642 ( .A(c1328), .B(b[1328]), .Z(n3985) );
XNOR U6643 ( .A(b[1328]), .B(n3986), .Z(c[1328]) );
XNOR U6644 ( .A(a[1328]), .B(c1328), .Z(n3986) );
XOR U6645 ( .A(c1329), .B(n3987), .Z(c1330) );
ANDN U6646 ( .B(n3988), .A(n3989), .Z(n3987) );
XOR U6647 ( .A(c1329), .B(b[1329]), .Z(n3988) );
XNOR U6648 ( .A(b[1329]), .B(n3989), .Z(c[1329]) );
XNOR U6649 ( .A(a[1329]), .B(c1329), .Z(n3989) );
XOR U6650 ( .A(c1330), .B(n3990), .Z(c1331) );
ANDN U6651 ( .B(n3991), .A(n3992), .Z(n3990) );
XOR U6652 ( .A(c1330), .B(b[1330]), .Z(n3991) );
XNOR U6653 ( .A(b[1330]), .B(n3992), .Z(c[1330]) );
XNOR U6654 ( .A(a[1330]), .B(c1330), .Z(n3992) );
XOR U6655 ( .A(c1331), .B(n3993), .Z(c1332) );
ANDN U6656 ( .B(n3994), .A(n3995), .Z(n3993) );
XOR U6657 ( .A(c1331), .B(b[1331]), .Z(n3994) );
XNOR U6658 ( .A(b[1331]), .B(n3995), .Z(c[1331]) );
XNOR U6659 ( .A(a[1331]), .B(c1331), .Z(n3995) );
XOR U6660 ( .A(c1332), .B(n3996), .Z(c1333) );
ANDN U6661 ( .B(n3997), .A(n3998), .Z(n3996) );
XOR U6662 ( .A(c1332), .B(b[1332]), .Z(n3997) );
XNOR U6663 ( .A(b[1332]), .B(n3998), .Z(c[1332]) );
XNOR U6664 ( .A(a[1332]), .B(c1332), .Z(n3998) );
XOR U6665 ( .A(c1333), .B(n3999), .Z(c1334) );
ANDN U6666 ( .B(n4000), .A(n4001), .Z(n3999) );
XOR U6667 ( .A(c1333), .B(b[1333]), .Z(n4000) );
XNOR U6668 ( .A(b[1333]), .B(n4001), .Z(c[1333]) );
XNOR U6669 ( .A(a[1333]), .B(c1333), .Z(n4001) );
XOR U6670 ( .A(c1334), .B(n4002), .Z(c1335) );
ANDN U6671 ( .B(n4003), .A(n4004), .Z(n4002) );
XOR U6672 ( .A(c1334), .B(b[1334]), .Z(n4003) );
XNOR U6673 ( .A(b[1334]), .B(n4004), .Z(c[1334]) );
XNOR U6674 ( .A(a[1334]), .B(c1334), .Z(n4004) );
XOR U6675 ( .A(c1335), .B(n4005), .Z(c1336) );
ANDN U6676 ( .B(n4006), .A(n4007), .Z(n4005) );
XOR U6677 ( .A(c1335), .B(b[1335]), .Z(n4006) );
XNOR U6678 ( .A(b[1335]), .B(n4007), .Z(c[1335]) );
XNOR U6679 ( .A(a[1335]), .B(c1335), .Z(n4007) );
XOR U6680 ( .A(c1336), .B(n4008), .Z(c1337) );
ANDN U6681 ( .B(n4009), .A(n4010), .Z(n4008) );
XOR U6682 ( .A(c1336), .B(b[1336]), .Z(n4009) );
XNOR U6683 ( .A(b[1336]), .B(n4010), .Z(c[1336]) );
XNOR U6684 ( .A(a[1336]), .B(c1336), .Z(n4010) );
XOR U6685 ( .A(c1337), .B(n4011), .Z(c1338) );
ANDN U6686 ( .B(n4012), .A(n4013), .Z(n4011) );
XOR U6687 ( .A(c1337), .B(b[1337]), .Z(n4012) );
XNOR U6688 ( .A(b[1337]), .B(n4013), .Z(c[1337]) );
XNOR U6689 ( .A(a[1337]), .B(c1337), .Z(n4013) );
XOR U6690 ( .A(c1338), .B(n4014), .Z(c1339) );
ANDN U6691 ( .B(n4015), .A(n4016), .Z(n4014) );
XOR U6692 ( .A(c1338), .B(b[1338]), .Z(n4015) );
XNOR U6693 ( .A(b[1338]), .B(n4016), .Z(c[1338]) );
XNOR U6694 ( .A(a[1338]), .B(c1338), .Z(n4016) );
XOR U6695 ( .A(c1339), .B(n4017), .Z(c1340) );
ANDN U6696 ( .B(n4018), .A(n4019), .Z(n4017) );
XOR U6697 ( .A(c1339), .B(b[1339]), .Z(n4018) );
XNOR U6698 ( .A(b[1339]), .B(n4019), .Z(c[1339]) );
XNOR U6699 ( .A(a[1339]), .B(c1339), .Z(n4019) );
XOR U6700 ( .A(c1340), .B(n4020), .Z(c1341) );
ANDN U6701 ( .B(n4021), .A(n4022), .Z(n4020) );
XOR U6702 ( .A(c1340), .B(b[1340]), .Z(n4021) );
XNOR U6703 ( .A(b[1340]), .B(n4022), .Z(c[1340]) );
XNOR U6704 ( .A(a[1340]), .B(c1340), .Z(n4022) );
XOR U6705 ( .A(c1341), .B(n4023), .Z(c1342) );
ANDN U6706 ( .B(n4024), .A(n4025), .Z(n4023) );
XOR U6707 ( .A(c1341), .B(b[1341]), .Z(n4024) );
XNOR U6708 ( .A(b[1341]), .B(n4025), .Z(c[1341]) );
XNOR U6709 ( .A(a[1341]), .B(c1341), .Z(n4025) );
XOR U6710 ( .A(c1342), .B(n4026), .Z(c1343) );
ANDN U6711 ( .B(n4027), .A(n4028), .Z(n4026) );
XOR U6712 ( .A(c1342), .B(b[1342]), .Z(n4027) );
XNOR U6713 ( .A(b[1342]), .B(n4028), .Z(c[1342]) );
XNOR U6714 ( .A(a[1342]), .B(c1342), .Z(n4028) );
XOR U6715 ( .A(c1343), .B(n4029), .Z(c1344) );
ANDN U6716 ( .B(n4030), .A(n4031), .Z(n4029) );
XOR U6717 ( .A(c1343), .B(b[1343]), .Z(n4030) );
XNOR U6718 ( .A(b[1343]), .B(n4031), .Z(c[1343]) );
XNOR U6719 ( .A(a[1343]), .B(c1343), .Z(n4031) );
XOR U6720 ( .A(c1344), .B(n4032), .Z(c1345) );
ANDN U6721 ( .B(n4033), .A(n4034), .Z(n4032) );
XOR U6722 ( .A(c1344), .B(b[1344]), .Z(n4033) );
XNOR U6723 ( .A(b[1344]), .B(n4034), .Z(c[1344]) );
XNOR U6724 ( .A(a[1344]), .B(c1344), .Z(n4034) );
XOR U6725 ( .A(c1345), .B(n4035), .Z(c1346) );
ANDN U6726 ( .B(n4036), .A(n4037), .Z(n4035) );
XOR U6727 ( .A(c1345), .B(b[1345]), .Z(n4036) );
XNOR U6728 ( .A(b[1345]), .B(n4037), .Z(c[1345]) );
XNOR U6729 ( .A(a[1345]), .B(c1345), .Z(n4037) );
XOR U6730 ( .A(c1346), .B(n4038), .Z(c1347) );
ANDN U6731 ( .B(n4039), .A(n4040), .Z(n4038) );
XOR U6732 ( .A(c1346), .B(b[1346]), .Z(n4039) );
XNOR U6733 ( .A(b[1346]), .B(n4040), .Z(c[1346]) );
XNOR U6734 ( .A(a[1346]), .B(c1346), .Z(n4040) );
XOR U6735 ( .A(c1347), .B(n4041), .Z(c1348) );
ANDN U6736 ( .B(n4042), .A(n4043), .Z(n4041) );
XOR U6737 ( .A(c1347), .B(b[1347]), .Z(n4042) );
XNOR U6738 ( .A(b[1347]), .B(n4043), .Z(c[1347]) );
XNOR U6739 ( .A(a[1347]), .B(c1347), .Z(n4043) );
XOR U6740 ( .A(c1348), .B(n4044), .Z(c1349) );
ANDN U6741 ( .B(n4045), .A(n4046), .Z(n4044) );
XOR U6742 ( .A(c1348), .B(b[1348]), .Z(n4045) );
XNOR U6743 ( .A(b[1348]), .B(n4046), .Z(c[1348]) );
XNOR U6744 ( .A(a[1348]), .B(c1348), .Z(n4046) );
XOR U6745 ( .A(c1349), .B(n4047), .Z(c1350) );
ANDN U6746 ( .B(n4048), .A(n4049), .Z(n4047) );
XOR U6747 ( .A(c1349), .B(b[1349]), .Z(n4048) );
XNOR U6748 ( .A(b[1349]), .B(n4049), .Z(c[1349]) );
XNOR U6749 ( .A(a[1349]), .B(c1349), .Z(n4049) );
XOR U6750 ( .A(c1350), .B(n4050), .Z(c1351) );
ANDN U6751 ( .B(n4051), .A(n4052), .Z(n4050) );
XOR U6752 ( .A(c1350), .B(b[1350]), .Z(n4051) );
XNOR U6753 ( .A(b[1350]), .B(n4052), .Z(c[1350]) );
XNOR U6754 ( .A(a[1350]), .B(c1350), .Z(n4052) );
XOR U6755 ( .A(c1351), .B(n4053), .Z(c1352) );
ANDN U6756 ( .B(n4054), .A(n4055), .Z(n4053) );
XOR U6757 ( .A(c1351), .B(b[1351]), .Z(n4054) );
XNOR U6758 ( .A(b[1351]), .B(n4055), .Z(c[1351]) );
XNOR U6759 ( .A(a[1351]), .B(c1351), .Z(n4055) );
XOR U6760 ( .A(c1352), .B(n4056), .Z(c1353) );
ANDN U6761 ( .B(n4057), .A(n4058), .Z(n4056) );
XOR U6762 ( .A(c1352), .B(b[1352]), .Z(n4057) );
XNOR U6763 ( .A(b[1352]), .B(n4058), .Z(c[1352]) );
XNOR U6764 ( .A(a[1352]), .B(c1352), .Z(n4058) );
XOR U6765 ( .A(c1353), .B(n4059), .Z(c1354) );
ANDN U6766 ( .B(n4060), .A(n4061), .Z(n4059) );
XOR U6767 ( .A(c1353), .B(b[1353]), .Z(n4060) );
XNOR U6768 ( .A(b[1353]), .B(n4061), .Z(c[1353]) );
XNOR U6769 ( .A(a[1353]), .B(c1353), .Z(n4061) );
XOR U6770 ( .A(c1354), .B(n4062), .Z(c1355) );
ANDN U6771 ( .B(n4063), .A(n4064), .Z(n4062) );
XOR U6772 ( .A(c1354), .B(b[1354]), .Z(n4063) );
XNOR U6773 ( .A(b[1354]), .B(n4064), .Z(c[1354]) );
XNOR U6774 ( .A(a[1354]), .B(c1354), .Z(n4064) );
XOR U6775 ( .A(c1355), .B(n4065), .Z(c1356) );
ANDN U6776 ( .B(n4066), .A(n4067), .Z(n4065) );
XOR U6777 ( .A(c1355), .B(b[1355]), .Z(n4066) );
XNOR U6778 ( .A(b[1355]), .B(n4067), .Z(c[1355]) );
XNOR U6779 ( .A(a[1355]), .B(c1355), .Z(n4067) );
XOR U6780 ( .A(c1356), .B(n4068), .Z(c1357) );
ANDN U6781 ( .B(n4069), .A(n4070), .Z(n4068) );
XOR U6782 ( .A(c1356), .B(b[1356]), .Z(n4069) );
XNOR U6783 ( .A(b[1356]), .B(n4070), .Z(c[1356]) );
XNOR U6784 ( .A(a[1356]), .B(c1356), .Z(n4070) );
XOR U6785 ( .A(c1357), .B(n4071), .Z(c1358) );
ANDN U6786 ( .B(n4072), .A(n4073), .Z(n4071) );
XOR U6787 ( .A(c1357), .B(b[1357]), .Z(n4072) );
XNOR U6788 ( .A(b[1357]), .B(n4073), .Z(c[1357]) );
XNOR U6789 ( .A(a[1357]), .B(c1357), .Z(n4073) );
XOR U6790 ( .A(c1358), .B(n4074), .Z(c1359) );
ANDN U6791 ( .B(n4075), .A(n4076), .Z(n4074) );
XOR U6792 ( .A(c1358), .B(b[1358]), .Z(n4075) );
XNOR U6793 ( .A(b[1358]), .B(n4076), .Z(c[1358]) );
XNOR U6794 ( .A(a[1358]), .B(c1358), .Z(n4076) );
XOR U6795 ( .A(c1359), .B(n4077), .Z(c1360) );
ANDN U6796 ( .B(n4078), .A(n4079), .Z(n4077) );
XOR U6797 ( .A(c1359), .B(b[1359]), .Z(n4078) );
XNOR U6798 ( .A(b[1359]), .B(n4079), .Z(c[1359]) );
XNOR U6799 ( .A(a[1359]), .B(c1359), .Z(n4079) );
XOR U6800 ( .A(c1360), .B(n4080), .Z(c1361) );
ANDN U6801 ( .B(n4081), .A(n4082), .Z(n4080) );
XOR U6802 ( .A(c1360), .B(b[1360]), .Z(n4081) );
XNOR U6803 ( .A(b[1360]), .B(n4082), .Z(c[1360]) );
XNOR U6804 ( .A(a[1360]), .B(c1360), .Z(n4082) );
XOR U6805 ( .A(c1361), .B(n4083), .Z(c1362) );
ANDN U6806 ( .B(n4084), .A(n4085), .Z(n4083) );
XOR U6807 ( .A(c1361), .B(b[1361]), .Z(n4084) );
XNOR U6808 ( .A(b[1361]), .B(n4085), .Z(c[1361]) );
XNOR U6809 ( .A(a[1361]), .B(c1361), .Z(n4085) );
XOR U6810 ( .A(c1362), .B(n4086), .Z(c1363) );
ANDN U6811 ( .B(n4087), .A(n4088), .Z(n4086) );
XOR U6812 ( .A(c1362), .B(b[1362]), .Z(n4087) );
XNOR U6813 ( .A(b[1362]), .B(n4088), .Z(c[1362]) );
XNOR U6814 ( .A(a[1362]), .B(c1362), .Z(n4088) );
XOR U6815 ( .A(c1363), .B(n4089), .Z(c1364) );
ANDN U6816 ( .B(n4090), .A(n4091), .Z(n4089) );
XOR U6817 ( .A(c1363), .B(b[1363]), .Z(n4090) );
XNOR U6818 ( .A(b[1363]), .B(n4091), .Z(c[1363]) );
XNOR U6819 ( .A(a[1363]), .B(c1363), .Z(n4091) );
XOR U6820 ( .A(c1364), .B(n4092), .Z(c1365) );
ANDN U6821 ( .B(n4093), .A(n4094), .Z(n4092) );
XOR U6822 ( .A(c1364), .B(b[1364]), .Z(n4093) );
XNOR U6823 ( .A(b[1364]), .B(n4094), .Z(c[1364]) );
XNOR U6824 ( .A(a[1364]), .B(c1364), .Z(n4094) );
XOR U6825 ( .A(c1365), .B(n4095), .Z(c1366) );
ANDN U6826 ( .B(n4096), .A(n4097), .Z(n4095) );
XOR U6827 ( .A(c1365), .B(b[1365]), .Z(n4096) );
XNOR U6828 ( .A(b[1365]), .B(n4097), .Z(c[1365]) );
XNOR U6829 ( .A(a[1365]), .B(c1365), .Z(n4097) );
XOR U6830 ( .A(c1366), .B(n4098), .Z(c1367) );
ANDN U6831 ( .B(n4099), .A(n4100), .Z(n4098) );
XOR U6832 ( .A(c1366), .B(b[1366]), .Z(n4099) );
XNOR U6833 ( .A(b[1366]), .B(n4100), .Z(c[1366]) );
XNOR U6834 ( .A(a[1366]), .B(c1366), .Z(n4100) );
XOR U6835 ( .A(c1367), .B(n4101), .Z(c1368) );
ANDN U6836 ( .B(n4102), .A(n4103), .Z(n4101) );
XOR U6837 ( .A(c1367), .B(b[1367]), .Z(n4102) );
XNOR U6838 ( .A(b[1367]), .B(n4103), .Z(c[1367]) );
XNOR U6839 ( .A(a[1367]), .B(c1367), .Z(n4103) );
XOR U6840 ( .A(c1368), .B(n4104), .Z(c1369) );
ANDN U6841 ( .B(n4105), .A(n4106), .Z(n4104) );
XOR U6842 ( .A(c1368), .B(b[1368]), .Z(n4105) );
XNOR U6843 ( .A(b[1368]), .B(n4106), .Z(c[1368]) );
XNOR U6844 ( .A(a[1368]), .B(c1368), .Z(n4106) );
XOR U6845 ( .A(c1369), .B(n4107), .Z(c1370) );
ANDN U6846 ( .B(n4108), .A(n4109), .Z(n4107) );
XOR U6847 ( .A(c1369), .B(b[1369]), .Z(n4108) );
XNOR U6848 ( .A(b[1369]), .B(n4109), .Z(c[1369]) );
XNOR U6849 ( .A(a[1369]), .B(c1369), .Z(n4109) );
XOR U6850 ( .A(c1370), .B(n4110), .Z(c1371) );
ANDN U6851 ( .B(n4111), .A(n4112), .Z(n4110) );
XOR U6852 ( .A(c1370), .B(b[1370]), .Z(n4111) );
XNOR U6853 ( .A(b[1370]), .B(n4112), .Z(c[1370]) );
XNOR U6854 ( .A(a[1370]), .B(c1370), .Z(n4112) );
XOR U6855 ( .A(c1371), .B(n4113), .Z(c1372) );
ANDN U6856 ( .B(n4114), .A(n4115), .Z(n4113) );
XOR U6857 ( .A(c1371), .B(b[1371]), .Z(n4114) );
XNOR U6858 ( .A(b[1371]), .B(n4115), .Z(c[1371]) );
XNOR U6859 ( .A(a[1371]), .B(c1371), .Z(n4115) );
XOR U6860 ( .A(c1372), .B(n4116), .Z(c1373) );
ANDN U6861 ( .B(n4117), .A(n4118), .Z(n4116) );
XOR U6862 ( .A(c1372), .B(b[1372]), .Z(n4117) );
XNOR U6863 ( .A(b[1372]), .B(n4118), .Z(c[1372]) );
XNOR U6864 ( .A(a[1372]), .B(c1372), .Z(n4118) );
XOR U6865 ( .A(c1373), .B(n4119), .Z(c1374) );
ANDN U6866 ( .B(n4120), .A(n4121), .Z(n4119) );
XOR U6867 ( .A(c1373), .B(b[1373]), .Z(n4120) );
XNOR U6868 ( .A(b[1373]), .B(n4121), .Z(c[1373]) );
XNOR U6869 ( .A(a[1373]), .B(c1373), .Z(n4121) );
XOR U6870 ( .A(c1374), .B(n4122), .Z(c1375) );
ANDN U6871 ( .B(n4123), .A(n4124), .Z(n4122) );
XOR U6872 ( .A(c1374), .B(b[1374]), .Z(n4123) );
XNOR U6873 ( .A(b[1374]), .B(n4124), .Z(c[1374]) );
XNOR U6874 ( .A(a[1374]), .B(c1374), .Z(n4124) );
XOR U6875 ( .A(c1375), .B(n4125), .Z(c1376) );
ANDN U6876 ( .B(n4126), .A(n4127), .Z(n4125) );
XOR U6877 ( .A(c1375), .B(b[1375]), .Z(n4126) );
XNOR U6878 ( .A(b[1375]), .B(n4127), .Z(c[1375]) );
XNOR U6879 ( .A(a[1375]), .B(c1375), .Z(n4127) );
XOR U6880 ( .A(c1376), .B(n4128), .Z(c1377) );
ANDN U6881 ( .B(n4129), .A(n4130), .Z(n4128) );
XOR U6882 ( .A(c1376), .B(b[1376]), .Z(n4129) );
XNOR U6883 ( .A(b[1376]), .B(n4130), .Z(c[1376]) );
XNOR U6884 ( .A(a[1376]), .B(c1376), .Z(n4130) );
XOR U6885 ( .A(c1377), .B(n4131), .Z(c1378) );
ANDN U6886 ( .B(n4132), .A(n4133), .Z(n4131) );
XOR U6887 ( .A(c1377), .B(b[1377]), .Z(n4132) );
XNOR U6888 ( .A(b[1377]), .B(n4133), .Z(c[1377]) );
XNOR U6889 ( .A(a[1377]), .B(c1377), .Z(n4133) );
XOR U6890 ( .A(c1378), .B(n4134), .Z(c1379) );
ANDN U6891 ( .B(n4135), .A(n4136), .Z(n4134) );
XOR U6892 ( .A(c1378), .B(b[1378]), .Z(n4135) );
XNOR U6893 ( .A(b[1378]), .B(n4136), .Z(c[1378]) );
XNOR U6894 ( .A(a[1378]), .B(c1378), .Z(n4136) );
XOR U6895 ( .A(c1379), .B(n4137), .Z(c1380) );
ANDN U6896 ( .B(n4138), .A(n4139), .Z(n4137) );
XOR U6897 ( .A(c1379), .B(b[1379]), .Z(n4138) );
XNOR U6898 ( .A(b[1379]), .B(n4139), .Z(c[1379]) );
XNOR U6899 ( .A(a[1379]), .B(c1379), .Z(n4139) );
XOR U6900 ( .A(c1380), .B(n4140), .Z(c1381) );
ANDN U6901 ( .B(n4141), .A(n4142), .Z(n4140) );
XOR U6902 ( .A(c1380), .B(b[1380]), .Z(n4141) );
XNOR U6903 ( .A(b[1380]), .B(n4142), .Z(c[1380]) );
XNOR U6904 ( .A(a[1380]), .B(c1380), .Z(n4142) );
XOR U6905 ( .A(c1381), .B(n4143), .Z(c1382) );
ANDN U6906 ( .B(n4144), .A(n4145), .Z(n4143) );
XOR U6907 ( .A(c1381), .B(b[1381]), .Z(n4144) );
XNOR U6908 ( .A(b[1381]), .B(n4145), .Z(c[1381]) );
XNOR U6909 ( .A(a[1381]), .B(c1381), .Z(n4145) );
XOR U6910 ( .A(c1382), .B(n4146), .Z(c1383) );
ANDN U6911 ( .B(n4147), .A(n4148), .Z(n4146) );
XOR U6912 ( .A(c1382), .B(b[1382]), .Z(n4147) );
XNOR U6913 ( .A(b[1382]), .B(n4148), .Z(c[1382]) );
XNOR U6914 ( .A(a[1382]), .B(c1382), .Z(n4148) );
XOR U6915 ( .A(c1383), .B(n4149), .Z(c1384) );
ANDN U6916 ( .B(n4150), .A(n4151), .Z(n4149) );
XOR U6917 ( .A(c1383), .B(b[1383]), .Z(n4150) );
XNOR U6918 ( .A(b[1383]), .B(n4151), .Z(c[1383]) );
XNOR U6919 ( .A(a[1383]), .B(c1383), .Z(n4151) );
XOR U6920 ( .A(c1384), .B(n4152), .Z(c1385) );
ANDN U6921 ( .B(n4153), .A(n4154), .Z(n4152) );
XOR U6922 ( .A(c1384), .B(b[1384]), .Z(n4153) );
XNOR U6923 ( .A(b[1384]), .B(n4154), .Z(c[1384]) );
XNOR U6924 ( .A(a[1384]), .B(c1384), .Z(n4154) );
XOR U6925 ( .A(c1385), .B(n4155), .Z(c1386) );
ANDN U6926 ( .B(n4156), .A(n4157), .Z(n4155) );
XOR U6927 ( .A(c1385), .B(b[1385]), .Z(n4156) );
XNOR U6928 ( .A(b[1385]), .B(n4157), .Z(c[1385]) );
XNOR U6929 ( .A(a[1385]), .B(c1385), .Z(n4157) );
XOR U6930 ( .A(c1386), .B(n4158), .Z(c1387) );
ANDN U6931 ( .B(n4159), .A(n4160), .Z(n4158) );
XOR U6932 ( .A(c1386), .B(b[1386]), .Z(n4159) );
XNOR U6933 ( .A(b[1386]), .B(n4160), .Z(c[1386]) );
XNOR U6934 ( .A(a[1386]), .B(c1386), .Z(n4160) );
XOR U6935 ( .A(c1387), .B(n4161), .Z(c1388) );
ANDN U6936 ( .B(n4162), .A(n4163), .Z(n4161) );
XOR U6937 ( .A(c1387), .B(b[1387]), .Z(n4162) );
XNOR U6938 ( .A(b[1387]), .B(n4163), .Z(c[1387]) );
XNOR U6939 ( .A(a[1387]), .B(c1387), .Z(n4163) );
XOR U6940 ( .A(c1388), .B(n4164), .Z(c1389) );
ANDN U6941 ( .B(n4165), .A(n4166), .Z(n4164) );
XOR U6942 ( .A(c1388), .B(b[1388]), .Z(n4165) );
XNOR U6943 ( .A(b[1388]), .B(n4166), .Z(c[1388]) );
XNOR U6944 ( .A(a[1388]), .B(c1388), .Z(n4166) );
XOR U6945 ( .A(c1389), .B(n4167), .Z(c1390) );
ANDN U6946 ( .B(n4168), .A(n4169), .Z(n4167) );
XOR U6947 ( .A(c1389), .B(b[1389]), .Z(n4168) );
XNOR U6948 ( .A(b[1389]), .B(n4169), .Z(c[1389]) );
XNOR U6949 ( .A(a[1389]), .B(c1389), .Z(n4169) );
XOR U6950 ( .A(c1390), .B(n4170), .Z(c1391) );
ANDN U6951 ( .B(n4171), .A(n4172), .Z(n4170) );
XOR U6952 ( .A(c1390), .B(b[1390]), .Z(n4171) );
XNOR U6953 ( .A(b[1390]), .B(n4172), .Z(c[1390]) );
XNOR U6954 ( .A(a[1390]), .B(c1390), .Z(n4172) );
XOR U6955 ( .A(c1391), .B(n4173), .Z(c1392) );
ANDN U6956 ( .B(n4174), .A(n4175), .Z(n4173) );
XOR U6957 ( .A(c1391), .B(b[1391]), .Z(n4174) );
XNOR U6958 ( .A(b[1391]), .B(n4175), .Z(c[1391]) );
XNOR U6959 ( .A(a[1391]), .B(c1391), .Z(n4175) );
XOR U6960 ( .A(c1392), .B(n4176), .Z(c1393) );
ANDN U6961 ( .B(n4177), .A(n4178), .Z(n4176) );
XOR U6962 ( .A(c1392), .B(b[1392]), .Z(n4177) );
XNOR U6963 ( .A(b[1392]), .B(n4178), .Z(c[1392]) );
XNOR U6964 ( .A(a[1392]), .B(c1392), .Z(n4178) );
XOR U6965 ( .A(c1393), .B(n4179), .Z(c1394) );
ANDN U6966 ( .B(n4180), .A(n4181), .Z(n4179) );
XOR U6967 ( .A(c1393), .B(b[1393]), .Z(n4180) );
XNOR U6968 ( .A(b[1393]), .B(n4181), .Z(c[1393]) );
XNOR U6969 ( .A(a[1393]), .B(c1393), .Z(n4181) );
XOR U6970 ( .A(c1394), .B(n4182), .Z(c1395) );
ANDN U6971 ( .B(n4183), .A(n4184), .Z(n4182) );
XOR U6972 ( .A(c1394), .B(b[1394]), .Z(n4183) );
XNOR U6973 ( .A(b[1394]), .B(n4184), .Z(c[1394]) );
XNOR U6974 ( .A(a[1394]), .B(c1394), .Z(n4184) );
XOR U6975 ( .A(c1395), .B(n4185), .Z(c1396) );
ANDN U6976 ( .B(n4186), .A(n4187), .Z(n4185) );
XOR U6977 ( .A(c1395), .B(b[1395]), .Z(n4186) );
XNOR U6978 ( .A(b[1395]), .B(n4187), .Z(c[1395]) );
XNOR U6979 ( .A(a[1395]), .B(c1395), .Z(n4187) );
XOR U6980 ( .A(c1396), .B(n4188), .Z(c1397) );
ANDN U6981 ( .B(n4189), .A(n4190), .Z(n4188) );
XOR U6982 ( .A(c1396), .B(b[1396]), .Z(n4189) );
XNOR U6983 ( .A(b[1396]), .B(n4190), .Z(c[1396]) );
XNOR U6984 ( .A(a[1396]), .B(c1396), .Z(n4190) );
XOR U6985 ( .A(c1397), .B(n4191), .Z(c1398) );
ANDN U6986 ( .B(n4192), .A(n4193), .Z(n4191) );
XOR U6987 ( .A(c1397), .B(b[1397]), .Z(n4192) );
XNOR U6988 ( .A(b[1397]), .B(n4193), .Z(c[1397]) );
XNOR U6989 ( .A(a[1397]), .B(c1397), .Z(n4193) );
XOR U6990 ( .A(c1398), .B(n4194), .Z(c1399) );
ANDN U6991 ( .B(n4195), .A(n4196), .Z(n4194) );
XOR U6992 ( .A(c1398), .B(b[1398]), .Z(n4195) );
XNOR U6993 ( .A(b[1398]), .B(n4196), .Z(c[1398]) );
XNOR U6994 ( .A(a[1398]), .B(c1398), .Z(n4196) );
XOR U6995 ( .A(c1399), .B(n4197), .Z(c1400) );
ANDN U6996 ( .B(n4198), .A(n4199), .Z(n4197) );
XOR U6997 ( .A(c1399), .B(b[1399]), .Z(n4198) );
XNOR U6998 ( .A(b[1399]), .B(n4199), .Z(c[1399]) );
XNOR U6999 ( .A(a[1399]), .B(c1399), .Z(n4199) );
XOR U7000 ( .A(c1400), .B(n4200), .Z(c1401) );
ANDN U7001 ( .B(n4201), .A(n4202), .Z(n4200) );
XOR U7002 ( .A(c1400), .B(b[1400]), .Z(n4201) );
XNOR U7003 ( .A(b[1400]), .B(n4202), .Z(c[1400]) );
XNOR U7004 ( .A(a[1400]), .B(c1400), .Z(n4202) );
XOR U7005 ( .A(c1401), .B(n4203), .Z(c1402) );
ANDN U7006 ( .B(n4204), .A(n4205), .Z(n4203) );
XOR U7007 ( .A(c1401), .B(b[1401]), .Z(n4204) );
XNOR U7008 ( .A(b[1401]), .B(n4205), .Z(c[1401]) );
XNOR U7009 ( .A(a[1401]), .B(c1401), .Z(n4205) );
XOR U7010 ( .A(c1402), .B(n4206), .Z(c1403) );
ANDN U7011 ( .B(n4207), .A(n4208), .Z(n4206) );
XOR U7012 ( .A(c1402), .B(b[1402]), .Z(n4207) );
XNOR U7013 ( .A(b[1402]), .B(n4208), .Z(c[1402]) );
XNOR U7014 ( .A(a[1402]), .B(c1402), .Z(n4208) );
XOR U7015 ( .A(c1403), .B(n4209), .Z(c1404) );
ANDN U7016 ( .B(n4210), .A(n4211), .Z(n4209) );
XOR U7017 ( .A(c1403), .B(b[1403]), .Z(n4210) );
XNOR U7018 ( .A(b[1403]), .B(n4211), .Z(c[1403]) );
XNOR U7019 ( .A(a[1403]), .B(c1403), .Z(n4211) );
XOR U7020 ( .A(c1404), .B(n4212), .Z(c1405) );
ANDN U7021 ( .B(n4213), .A(n4214), .Z(n4212) );
XOR U7022 ( .A(c1404), .B(b[1404]), .Z(n4213) );
XNOR U7023 ( .A(b[1404]), .B(n4214), .Z(c[1404]) );
XNOR U7024 ( .A(a[1404]), .B(c1404), .Z(n4214) );
XOR U7025 ( .A(c1405), .B(n4215), .Z(c1406) );
ANDN U7026 ( .B(n4216), .A(n4217), .Z(n4215) );
XOR U7027 ( .A(c1405), .B(b[1405]), .Z(n4216) );
XNOR U7028 ( .A(b[1405]), .B(n4217), .Z(c[1405]) );
XNOR U7029 ( .A(a[1405]), .B(c1405), .Z(n4217) );
XOR U7030 ( .A(c1406), .B(n4218), .Z(c1407) );
ANDN U7031 ( .B(n4219), .A(n4220), .Z(n4218) );
XOR U7032 ( .A(c1406), .B(b[1406]), .Z(n4219) );
XNOR U7033 ( .A(b[1406]), .B(n4220), .Z(c[1406]) );
XNOR U7034 ( .A(a[1406]), .B(c1406), .Z(n4220) );
XOR U7035 ( .A(c1407), .B(n4221), .Z(c1408) );
ANDN U7036 ( .B(n4222), .A(n4223), .Z(n4221) );
XOR U7037 ( .A(c1407), .B(b[1407]), .Z(n4222) );
XNOR U7038 ( .A(b[1407]), .B(n4223), .Z(c[1407]) );
XNOR U7039 ( .A(a[1407]), .B(c1407), .Z(n4223) );
XOR U7040 ( .A(c1408), .B(n4224), .Z(c1409) );
ANDN U7041 ( .B(n4225), .A(n4226), .Z(n4224) );
XOR U7042 ( .A(c1408), .B(b[1408]), .Z(n4225) );
XNOR U7043 ( .A(b[1408]), .B(n4226), .Z(c[1408]) );
XNOR U7044 ( .A(a[1408]), .B(c1408), .Z(n4226) );
XOR U7045 ( .A(c1409), .B(n4227), .Z(c1410) );
ANDN U7046 ( .B(n4228), .A(n4229), .Z(n4227) );
XOR U7047 ( .A(c1409), .B(b[1409]), .Z(n4228) );
XNOR U7048 ( .A(b[1409]), .B(n4229), .Z(c[1409]) );
XNOR U7049 ( .A(a[1409]), .B(c1409), .Z(n4229) );
XOR U7050 ( .A(c1410), .B(n4230), .Z(c1411) );
ANDN U7051 ( .B(n4231), .A(n4232), .Z(n4230) );
XOR U7052 ( .A(c1410), .B(b[1410]), .Z(n4231) );
XNOR U7053 ( .A(b[1410]), .B(n4232), .Z(c[1410]) );
XNOR U7054 ( .A(a[1410]), .B(c1410), .Z(n4232) );
XOR U7055 ( .A(c1411), .B(n4233), .Z(c1412) );
ANDN U7056 ( .B(n4234), .A(n4235), .Z(n4233) );
XOR U7057 ( .A(c1411), .B(b[1411]), .Z(n4234) );
XNOR U7058 ( .A(b[1411]), .B(n4235), .Z(c[1411]) );
XNOR U7059 ( .A(a[1411]), .B(c1411), .Z(n4235) );
XOR U7060 ( .A(c1412), .B(n4236), .Z(c1413) );
ANDN U7061 ( .B(n4237), .A(n4238), .Z(n4236) );
XOR U7062 ( .A(c1412), .B(b[1412]), .Z(n4237) );
XNOR U7063 ( .A(b[1412]), .B(n4238), .Z(c[1412]) );
XNOR U7064 ( .A(a[1412]), .B(c1412), .Z(n4238) );
XOR U7065 ( .A(c1413), .B(n4239), .Z(c1414) );
ANDN U7066 ( .B(n4240), .A(n4241), .Z(n4239) );
XOR U7067 ( .A(c1413), .B(b[1413]), .Z(n4240) );
XNOR U7068 ( .A(b[1413]), .B(n4241), .Z(c[1413]) );
XNOR U7069 ( .A(a[1413]), .B(c1413), .Z(n4241) );
XOR U7070 ( .A(c1414), .B(n4242), .Z(c1415) );
ANDN U7071 ( .B(n4243), .A(n4244), .Z(n4242) );
XOR U7072 ( .A(c1414), .B(b[1414]), .Z(n4243) );
XNOR U7073 ( .A(b[1414]), .B(n4244), .Z(c[1414]) );
XNOR U7074 ( .A(a[1414]), .B(c1414), .Z(n4244) );
XOR U7075 ( .A(c1415), .B(n4245), .Z(c1416) );
ANDN U7076 ( .B(n4246), .A(n4247), .Z(n4245) );
XOR U7077 ( .A(c1415), .B(b[1415]), .Z(n4246) );
XNOR U7078 ( .A(b[1415]), .B(n4247), .Z(c[1415]) );
XNOR U7079 ( .A(a[1415]), .B(c1415), .Z(n4247) );
XOR U7080 ( .A(c1416), .B(n4248), .Z(c1417) );
ANDN U7081 ( .B(n4249), .A(n4250), .Z(n4248) );
XOR U7082 ( .A(c1416), .B(b[1416]), .Z(n4249) );
XNOR U7083 ( .A(b[1416]), .B(n4250), .Z(c[1416]) );
XNOR U7084 ( .A(a[1416]), .B(c1416), .Z(n4250) );
XOR U7085 ( .A(c1417), .B(n4251), .Z(c1418) );
ANDN U7086 ( .B(n4252), .A(n4253), .Z(n4251) );
XOR U7087 ( .A(c1417), .B(b[1417]), .Z(n4252) );
XNOR U7088 ( .A(b[1417]), .B(n4253), .Z(c[1417]) );
XNOR U7089 ( .A(a[1417]), .B(c1417), .Z(n4253) );
XOR U7090 ( .A(c1418), .B(n4254), .Z(c1419) );
ANDN U7091 ( .B(n4255), .A(n4256), .Z(n4254) );
XOR U7092 ( .A(c1418), .B(b[1418]), .Z(n4255) );
XNOR U7093 ( .A(b[1418]), .B(n4256), .Z(c[1418]) );
XNOR U7094 ( .A(a[1418]), .B(c1418), .Z(n4256) );
XOR U7095 ( .A(c1419), .B(n4257), .Z(c1420) );
ANDN U7096 ( .B(n4258), .A(n4259), .Z(n4257) );
XOR U7097 ( .A(c1419), .B(b[1419]), .Z(n4258) );
XNOR U7098 ( .A(b[1419]), .B(n4259), .Z(c[1419]) );
XNOR U7099 ( .A(a[1419]), .B(c1419), .Z(n4259) );
XOR U7100 ( .A(c1420), .B(n4260), .Z(c1421) );
ANDN U7101 ( .B(n4261), .A(n4262), .Z(n4260) );
XOR U7102 ( .A(c1420), .B(b[1420]), .Z(n4261) );
XNOR U7103 ( .A(b[1420]), .B(n4262), .Z(c[1420]) );
XNOR U7104 ( .A(a[1420]), .B(c1420), .Z(n4262) );
XOR U7105 ( .A(c1421), .B(n4263), .Z(c1422) );
ANDN U7106 ( .B(n4264), .A(n4265), .Z(n4263) );
XOR U7107 ( .A(c1421), .B(b[1421]), .Z(n4264) );
XNOR U7108 ( .A(b[1421]), .B(n4265), .Z(c[1421]) );
XNOR U7109 ( .A(a[1421]), .B(c1421), .Z(n4265) );
XOR U7110 ( .A(c1422), .B(n4266), .Z(c1423) );
ANDN U7111 ( .B(n4267), .A(n4268), .Z(n4266) );
XOR U7112 ( .A(c1422), .B(b[1422]), .Z(n4267) );
XNOR U7113 ( .A(b[1422]), .B(n4268), .Z(c[1422]) );
XNOR U7114 ( .A(a[1422]), .B(c1422), .Z(n4268) );
XOR U7115 ( .A(c1423), .B(n4269), .Z(c1424) );
ANDN U7116 ( .B(n4270), .A(n4271), .Z(n4269) );
XOR U7117 ( .A(c1423), .B(b[1423]), .Z(n4270) );
XNOR U7118 ( .A(b[1423]), .B(n4271), .Z(c[1423]) );
XNOR U7119 ( .A(a[1423]), .B(c1423), .Z(n4271) );
XOR U7120 ( .A(c1424), .B(n4272), .Z(c1425) );
ANDN U7121 ( .B(n4273), .A(n4274), .Z(n4272) );
XOR U7122 ( .A(c1424), .B(b[1424]), .Z(n4273) );
XNOR U7123 ( .A(b[1424]), .B(n4274), .Z(c[1424]) );
XNOR U7124 ( .A(a[1424]), .B(c1424), .Z(n4274) );
XOR U7125 ( .A(c1425), .B(n4275), .Z(c1426) );
ANDN U7126 ( .B(n4276), .A(n4277), .Z(n4275) );
XOR U7127 ( .A(c1425), .B(b[1425]), .Z(n4276) );
XNOR U7128 ( .A(b[1425]), .B(n4277), .Z(c[1425]) );
XNOR U7129 ( .A(a[1425]), .B(c1425), .Z(n4277) );
XOR U7130 ( .A(c1426), .B(n4278), .Z(c1427) );
ANDN U7131 ( .B(n4279), .A(n4280), .Z(n4278) );
XOR U7132 ( .A(c1426), .B(b[1426]), .Z(n4279) );
XNOR U7133 ( .A(b[1426]), .B(n4280), .Z(c[1426]) );
XNOR U7134 ( .A(a[1426]), .B(c1426), .Z(n4280) );
XOR U7135 ( .A(c1427), .B(n4281), .Z(c1428) );
ANDN U7136 ( .B(n4282), .A(n4283), .Z(n4281) );
XOR U7137 ( .A(c1427), .B(b[1427]), .Z(n4282) );
XNOR U7138 ( .A(b[1427]), .B(n4283), .Z(c[1427]) );
XNOR U7139 ( .A(a[1427]), .B(c1427), .Z(n4283) );
XOR U7140 ( .A(c1428), .B(n4284), .Z(c1429) );
ANDN U7141 ( .B(n4285), .A(n4286), .Z(n4284) );
XOR U7142 ( .A(c1428), .B(b[1428]), .Z(n4285) );
XNOR U7143 ( .A(b[1428]), .B(n4286), .Z(c[1428]) );
XNOR U7144 ( .A(a[1428]), .B(c1428), .Z(n4286) );
XOR U7145 ( .A(c1429), .B(n4287), .Z(c1430) );
ANDN U7146 ( .B(n4288), .A(n4289), .Z(n4287) );
XOR U7147 ( .A(c1429), .B(b[1429]), .Z(n4288) );
XNOR U7148 ( .A(b[1429]), .B(n4289), .Z(c[1429]) );
XNOR U7149 ( .A(a[1429]), .B(c1429), .Z(n4289) );
XOR U7150 ( .A(c1430), .B(n4290), .Z(c1431) );
ANDN U7151 ( .B(n4291), .A(n4292), .Z(n4290) );
XOR U7152 ( .A(c1430), .B(b[1430]), .Z(n4291) );
XNOR U7153 ( .A(b[1430]), .B(n4292), .Z(c[1430]) );
XNOR U7154 ( .A(a[1430]), .B(c1430), .Z(n4292) );
XOR U7155 ( .A(c1431), .B(n4293), .Z(c1432) );
ANDN U7156 ( .B(n4294), .A(n4295), .Z(n4293) );
XOR U7157 ( .A(c1431), .B(b[1431]), .Z(n4294) );
XNOR U7158 ( .A(b[1431]), .B(n4295), .Z(c[1431]) );
XNOR U7159 ( .A(a[1431]), .B(c1431), .Z(n4295) );
XOR U7160 ( .A(c1432), .B(n4296), .Z(c1433) );
ANDN U7161 ( .B(n4297), .A(n4298), .Z(n4296) );
XOR U7162 ( .A(c1432), .B(b[1432]), .Z(n4297) );
XNOR U7163 ( .A(b[1432]), .B(n4298), .Z(c[1432]) );
XNOR U7164 ( .A(a[1432]), .B(c1432), .Z(n4298) );
XOR U7165 ( .A(c1433), .B(n4299), .Z(c1434) );
ANDN U7166 ( .B(n4300), .A(n4301), .Z(n4299) );
XOR U7167 ( .A(c1433), .B(b[1433]), .Z(n4300) );
XNOR U7168 ( .A(b[1433]), .B(n4301), .Z(c[1433]) );
XNOR U7169 ( .A(a[1433]), .B(c1433), .Z(n4301) );
XOR U7170 ( .A(c1434), .B(n4302), .Z(c1435) );
ANDN U7171 ( .B(n4303), .A(n4304), .Z(n4302) );
XOR U7172 ( .A(c1434), .B(b[1434]), .Z(n4303) );
XNOR U7173 ( .A(b[1434]), .B(n4304), .Z(c[1434]) );
XNOR U7174 ( .A(a[1434]), .B(c1434), .Z(n4304) );
XOR U7175 ( .A(c1435), .B(n4305), .Z(c1436) );
ANDN U7176 ( .B(n4306), .A(n4307), .Z(n4305) );
XOR U7177 ( .A(c1435), .B(b[1435]), .Z(n4306) );
XNOR U7178 ( .A(b[1435]), .B(n4307), .Z(c[1435]) );
XNOR U7179 ( .A(a[1435]), .B(c1435), .Z(n4307) );
XOR U7180 ( .A(c1436), .B(n4308), .Z(c1437) );
ANDN U7181 ( .B(n4309), .A(n4310), .Z(n4308) );
XOR U7182 ( .A(c1436), .B(b[1436]), .Z(n4309) );
XNOR U7183 ( .A(b[1436]), .B(n4310), .Z(c[1436]) );
XNOR U7184 ( .A(a[1436]), .B(c1436), .Z(n4310) );
XOR U7185 ( .A(c1437), .B(n4311), .Z(c1438) );
ANDN U7186 ( .B(n4312), .A(n4313), .Z(n4311) );
XOR U7187 ( .A(c1437), .B(b[1437]), .Z(n4312) );
XNOR U7188 ( .A(b[1437]), .B(n4313), .Z(c[1437]) );
XNOR U7189 ( .A(a[1437]), .B(c1437), .Z(n4313) );
XOR U7190 ( .A(c1438), .B(n4314), .Z(c1439) );
ANDN U7191 ( .B(n4315), .A(n4316), .Z(n4314) );
XOR U7192 ( .A(c1438), .B(b[1438]), .Z(n4315) );
XNOR U7193 ( .A(b[1438]), .B(n4316), .Z(c[1438]) );
XNOR U7194 ( .A(a[1438]), .B(c1438), .Z(n4316) );
XOR U7195 ( .A(c1439), .B(n4317), .Z(c1440) );
ANDN U7196 ( .B(n4318), .A(n4319), .Z(n4317) );
XOR U7197 ( .A(c1439), .B(b[1439]), .Z(n4318) );
XNOR U7198 ( .A(b[1439]), .B(n4319), .Z(c[1439]) );
XNOR U7199 ( .A(a[1439]), .B(c1439), .Z(n4319) );
XOR U7200 ( .A(c1440), .B(n4320), .Z(c1441) );
ANDN U7201 ( .B(n4321), .A(n4322), .Z(n4320) );
XOR U7202 ( .A(c1440), .B(b[1440]), .Z(n4321) );
XNOR U7203 ( .A(b[1440]), .B(n4322), .Z(c[1440]) );
XNOR U7204 ( .A(a[1440]), .B(c1440), .Z(n4322) );
XOR U7205 ( .A(c1441), .B(n4323), .Z(c1442) );
ANDN U7206 ( .B(n4324), .A(n4325), .Z(n4323) );
XOR U7207 ( .A(c1441), .B(b[1441]), .Z(n4324) );
XNOR U7208 ( .A(b[1441]), .B(n4325), .Z(c[1441]) );
XNOR U7209 ( .A(a[1441]), .B(c1441), .Z(n4325) );
XOR U7210 ( .A(c1442), .B(n4326), .Z(c1443) );
ANDN U7211 ( .B(n4327), .A(n4328), .Z(n4326) );
XOR U7212 ( .A(c1442), .B(b[1442]), .Z(n4327) );
XNOR U7213 ( .A(b[1442]), .B(n4328), .Z(c[1442]) );
XNOR U7214 ( .A(a[1442]), .B(c1442), .Z(n4328) );
XOR U7215 ( .A(c1443), .B(n4329), .Z(c1444) );
ANDN U7216 ( .B(n4330), .A(n4331), .Z(n4329) );
XOR U7217 ( .A(c1443), .B(b[1443]), .Z(n4330) );
XNOR U7218 ( .A(b[1443]), .B(n4331), .Z(c[1443]) );
XNOR U7219 ( .A(a[1443]), .B(c1443), .Z(n4331) );
XOR U7220 ( .A(c1444), .B(n4332), .Z(c1445) );
ANDN U7221 ( .B(n4333), .A(n4334), .Z(n4332) );
XOR U7222 ( .A(c1444), .B(b[1444]), .Z(n4333) );
XNOR U7223 ( .A(b[1444]), .B(n4334), .Z(c[1444]) );
XNOR U7224 ( .A(a[1444]), .B(c1444), .Z(n4334) );
XOR U7225 ( .A(c1445), .B(n4335), .Z(c1446) );
ANDN U7226 ( .B(n4336), .A(n4337), .Z(n4335) );
XOR U7227 ( .A(c1445), .B(b[1445]), .Z(n4336) );
XNOR U7228 ( .A(b[1445]), .B(n4337), .Z(c[1445]) );
XNOR U7229 ( .A(a[1445]), .B(c1445), .Z(n4337) );
XOR U7230 ( .A(c1446), .B(n4338), .Z(c1447) );
ANDN U7231 ( .B(n4339), .A(n4340), .Z(n4338) );
XOR U7232 ( .A(c1446), .B(b[1446]), .Z(n4339) );
XNOR U7233 ( .A(b[1446]), .B(n4340), .Z(c[1446]) );
XNOR U7234 ( .A(a[1446]), .B(c1446), .Z(n4340) );
XOR U7235 ( .A(c1447), .B(n4341), .Z(c1448) );
ANDN U7236 ( .B(n4342), .A(n4343), .Z(n4341) );
XOR U7237 ( .A(c1447), .B(b[1447]), .Z(n4342) );
XNOR U7238 ( .A(b[1447]), .B(n4343), .Z(c[1447]) );
XNOR U7239 ( .A(a[1447]), .B(c1447), .Z(n4343) );
XOR U7240 ( .A(c1448), .B(n4344), .Z(c1449) );
ANDN U7241 ( .B(n4345), .A(n4346), .Z(n4344) );
XOR U7242 ( .A(c1448), .B(b[1448]), .Z(n4345) );
XNOR U7243 ( .A(b[1448]), .B(n4346), .Z(c[1448]) );
XNOR U7244 ( .A(a[1448]), .B(c1448), .Z(n4346) );
XOR U7245 ( .A(c1449), .B(n4347), .Z(c1450) );
ANDN U7246 ( .B(n4348), .A(n4349), .Z(n4347) );
XOR U7247 ( .A(c1449), .B(b[1449]), .Z(n4348) );
XNOR U7248 ( .A(b[1449]), .B(n4349), .Z(c[1449]) );
XNOR U7249 ( .A(a[1449]), .B(c1449), .Z(n4349) );
XOR U7250 ( .A(c1450), .B(n4350), .Z(c1451) );
ANDN U7251 ( .B(n4351), .A(n4352), .Z(n4350) );
XOR U7252 ( .A(c1450), .B(b[1450]), .Z(n4351) );
XNOR U7253 ( .A(b[1450]), .B(n4352), .Z(c[1450]) );
XNOR U7254 ( .A(a[1450]), .B(c1450), .Z(n4352) );
XOR U7255 ( .A(c1451), .B(n4353), .Z(c1452) );
ANDN U7256 ( .B(n4354), .A(n4355), .Z(n4353) );
XOR U7257 ( .A(c1451), .B(b[1451]), .Z(n4354) );
XNOR U7258 ( .A(b[1451]), .B(n4355), .Z(c[1451]) );
XNOR U7259 ( .A(a[1451]), .B(c1451), .Z(n4355) );
XOR U7260 ( .A(c1452), .B(n4356), .Z(c1453) );
ANDN U7261 ( .B(n4357), .A(n4358), .Z(n4356) );
XOR U7262 ( .A(c1452), .B(b[1452]), .Z(n4357) );
XNOR U7263 ( .A(b[1452]), .B(n4358), .Z(c[1452]) );
XNOR U7264 ( .A(a[1452]), .B(c1452), .Z(n4358) );
XOR U7265 ( .A(c1453), .B(n4359), .Z(c1454) );
ANDN U7266 ( .B(n4360), .A(n4361), .Z(n4359) );
XOR U7267 ( .A(c1453), .B(b[1453]), .Z(n4360) );
XNOR U7268 ( .A(b[1453]), .B(n4361), .Z(c[1453]) );
XNOR U7269 ( .A(a[1453]), .B(c1453), .Z(n4361) );
XOR U7270 ( .A(c1454), .B(n4362), .Z(c1455) );
ANDN U7271 ( .B(n4363), .A(n4364), .Z(n4362) );
XOR U7272 ( .A(c1454), .B(b[1454]), .Z(n4363) );
XNOR U7273 ( .A(b[1454]), .B(n4364), .Z(c[1454]) );
XNOR U7274 ( .A(a[1454]), .B(c1454), .Z(n4364) );
XOR U7275 ( .A(c1455), .B(n4365), .Z(c1456) );
ANDN U7276 ( .B(n4366), .A(n4367), .Z(n4365) );
XOR U7277 ( .A(c1455), .B(b[1455]), .Z(n4366) );
XNOR U7278 ( .A(b[1455]), .B(n4367), .Z(c[1455]) );
XNOR U7279 ( .A(a[1455]), .B(c1455), .Z(n4367) );
XOR U7280 ( .A(c1456), .B(n4368), .Z(c1457) );
ANDN U7281 ( .B(n4369), .A(n4370), .Z(n4368) );
XOR U7282 ( .A(c1456), .B(b[1456]), .Z(n4369) );
XNOR U7283 ( .A(b[1456]), .B(n4370), .Z(c[1456]) );
XNOR U7284 ( .A(a[1456]), .B(c1456), .Z(n4370) );
XOR U7285 ( .A(c1457), .B(n4371), .Z(c1458) );
ANDN U7286 ( .B(n4372), .A(n4373), .Z(n4371) );
XOR U7287 ( .A(c1457), .B(b[1457]), .Z(n4372) );
XNOR U7288 ( .A(b[1457]), .B(n4373), .Z(c[1457]) );
XNOR U7289 ( .A(a[1457]), .B(c1457), .Z(n4373) );
XOR U7290 ( .A(c1458), .B(n4374), .Z(c1459) );
ANDN U7291 ( .B(n4375), .A(n4376), .Z(n4374) );
XOR U7292 ( .A(c1458), .B(b[1458]), .Z(n4375) );
XNOR U7293 ( .A(b[1458]), .B(n4376), .Z(c[1458]) );
XNOR U7294 ( .A(a[1458]), .B(c1458), .Z(n4376) );
XOR U7295 ( .A(c1459), .B(n4377), .Z(c1460) );
ANDN U7296 ( .B(n4378), .A(n4379), .Z(n4377) );
XOR U7297 ( .A(c1459), .B(b[1459]), .Z(n4378) );
XNOR U7298 ( .A(b[1459]), .B(n4379), .Z(c[1459]) );
XNOR U7299 ( .A(a[1459]), .B(c1459), .Z(n4379) );
XOR U7300 ( .A(c1460), .B(n4380), .Z(c1461) );
ANDN U7301 ( .B(n4381), .A(n4382), .Z(n4380) );
XOR U7302 ( .A(c1460), .B(b[1460]), .Z(n4381) );
XNOR U7303 ( .A(b[1460]), .B(n4382), .Z(c[1460]) );
XNOR U7304 ( .A(a[1460]), .B(c1460), .Z(n4382) );
XOR U7305 ( .A(c1461), .B(n4383), .Z(c1462) );
ANDN U7306 ( .B(n4384), .A(n4385), .Z(n4383) );
XOR U7307 ( .A(c1461), .B(b[1461]), .Z(n4384) );
XNOR U7308 ( .A(b[1461]), .B(n4385), .Z(c[1461]) );
XNOR U7309 ( .A(a[1461]), .B(c1461), .Z(n4385) );
XOR U7310 ( .A(c1462), .B(n4386), .Z(c1463) );
ANDN U7311 ( .B(n4387), .A(n4388), .Z(n4386) );
XOR U7312 ( .A(c1462), .B(b[1462]), .Z(n4387) );
XNOR U7313 ( .A(b[1462]), .B(n4388), .Z(c[1462]) );
XNOR U7314 ( .A(a[1462]), .B(c1462), .Z(n4388) );
XOR U7315 ( .A(c1463), .B(n4389), .Z(c1464) );
ANDN U7316 ( .B(n4390), .A(n4391), .Z(n4389) );
XOR U7317 ( .A(c1463), .B(b[1463]), .Z(n4390) );
XNOR U7318 ( .A(b[1463]), .B(n4391), .Z(c[1463]) );
XNOR U7319 ( .A(a[1463]), .B(c1463), .Z(n4391) );
XOR U7320 ( .A(c1464), .B(n4392), .Z(c1465) );
ANDN U7321 ( .B(n4393), .A(n4394), .Z(n4392) );
XOR U7322 ( .A(c1464), .B(b[1464]), .Z(n4393) );
XNOR U7323 ( .A(b[1464]), .B(n4394), .Z(c[1464]) );
XNOR U7324 ( .A(a[1464]), .B(c1464), .Z(n4394) );
XOR U7325 ( .A(c1465), .B(n4395), .Z(c1466) );
ANDN U7326 ( .B(n4396), .A(n4397), .Z(n4395) );
XOR U7327 ( .A(c1465), .B(b[1465]), .Z(n4396) );
XNOR U7328 ( .A(b[1465]), .B(n4397), .Z(c[1465]) );
XNOR U7329 ( .A(a[1465]), .B(c1465), .Z(n4397) );
XOR U7330 ( .A(c1466), .B(n4398), .Z(c1467) );
ANDN U7331 ( .B(n4399), .A(n4400), .Z(n4398) );
XOR U7332 ( .A(c1466), .B(b[1466]), .Z(n4399) );
XNOR U7333 ( .A(b[1466]), .B(n4400), .Z(c[1466]) );
XNOR U7334 ( .A(a[1466]), .B(c1466), .Z(n4400) );
XOR U7335 ( .A(c1467), .B(n4401), .Z(c1468) );
ANDN U7336 ( .B(n4402), .A(n4403), .Z(n4401) );
XOR U7337 ( .A(c1467), .B(b[1467]), .Z(n4402) );
XNOR U7338 ( .A(b[1467]), .B(n4403), .Z(c[1467]) );
XNOR U7339 ( .A(a[1467]), .B(c1467), .Z(n4403) );
XOR U7340 ( .A(c1468), .B(n4404), .Z(c1469) );
ANDN U7341 ( .B(n4405), .A(n4406), .Z(n4404) );
XOR U7342 ( .A(c1468), .B(b[1468]), .Z(n4405) );
XNOR U7343 ( .A(b[1468]), .B(n4406), .Z(c[1468]) );
XNOR U7344 ( .A(a[1468]), .B(c1468), .Z(n4406) );
XOR U7345 ( .A(c1469), .B(n4407), .Z(c1470) );
ANDN U7346 ( .B(n4408), .A(n4409), .Z(n4407) );
XOR U7347 ( .A(c1469), .B(b[1469]), .Z(n4408) );
XNOR U7348 ( .A(b[1469]), .B(n4409), .Z(c[1469]) );
XNOR U7349 ( .A(a[1469]), .B(c1469), .Z(n4409) );
XOR U7350 ( .A(c1470), .B(n4410), .Z(c1471) );
ANDN U7351 ( .B(n4411), .A(n4412), .Z(n4410) );
XOR U7352 ( .A(c1470), .B(b[1470]), .Z(n4411) );
XNOR U7353 ( .A(b[1470]), .B(n4412), .Z(c[1470]) );
XNOR U7354 ( .A(a[1470]), .B(c1470), .Z(n4412) );
XOR U7355 ( .A(c1471), .B(n4413), .Z(c1472) );
ANDN U7356 ( .B(n4414), .A(n4415), .Z(n4413) );
XOR U7357 ( .A(c1471), .B(b[1471]), .Z(n4414) );
XNOR U7358 ( .A(b[1471]), .B(n4415), .Z(c[1471]) );
XNOR U7359 ( .A(a[1471]), .B(c1471), .Z(n4415) );
XOR U7360 ( .A(c1472), .B(n4416), .Z(c1473) );
ANDN U7361 ( .B(n4417), .A(n4418), .Z(n4416) );
XOR U7362 ( .A(c1472), .B(b[1472]), .Z(n4417) );
XNOR U7363 ( .A(b[1472]), .B(n4418), .Z(c[1472]) );
XNOR U7364 ( .A(a[1472]), .B(c1472), .Z(n4418) );
XOR U7365 ( .A(c1473), .B(n4419), .Z(c1474) );
ANDN U7366 ( .B(n4420), .A(n4421), .Z(n4419) );
XOR U7367 ( .A(c1473), .B(b[1473]), .Z(n4420) );
XNOR U7368 ( .A(b[1473]), .B(n4421), .Z(c[1473]) );
XNOR U7369 ( .A(a[1473]), .B(c1473), .Z(n4421) );
XOR U7370 ( .A(c1474), .B(n4422), .Z(c1475) );
ANDN U7371 ( .B(n4423), .A(n4424), .Z(n4422) );
XOR U7372 ( .A(c1474), .B(b[1474]), .Z(n4423) );
XNOR U7373 ( .A(b[1474]), .B(n4424), .Z(c[1474]) );
XNOR U7374 ( .A(a[1474]), .B(c1474), .Z(n4424) );
XOR U7375 ( .A(c1475), .B(n4425), .Z(c1476) );
ANDN U7376 ( .B(n4426), .A(n4427), .Z(n4425) );
XOR U7377 ( .A(c1475), .B(b[1475]), .Z(n4426) );
XNOR U7378 ( .A(b[1475]), .B(n4427), .Z(c[1475]) );
XNOR U7379 ( .A(a[1475]), .B(c1475), .Z(n4427) );
XOR U7380 ( .A(c1476), .B(n4428), .Z(c1477) );
ANDN U7381 ( .B(n4429), .A(n4430), .Z(n4428) );
XOR U7382 ( .A(c1476), .B(b[1476]), .Z(n4429) );
XNOR U7383 ( .A(b[1476]), .B(n4430), .Z(c[1476]) );
XNOR U7384 ( .A(a[1476]), .B(c1476), .Z(n4430) );
XOR U7385 ( .A(c1477), .B(n4431), .Z(c1478) );
ANDN U7386 ( .B(n4432), .A(n4433), .Z(n4431) );
XOR U7387 ( .A(c1477), .B(b[1477]), .Z(n4432) );
XNOR U7388 ( .A(b[1477]), .B(n4433), .Z(c[1477]) );
XNOR U7389 ( .A(a[1477]), .B(c1477), .Z(n4433) );
XOR U7390 ( .A(c1478), .B(n4434), .Z(c1479) );
ANDN U7391 ( .B(n4435), .A(n4436), .Z(n4434) );
XOR U7392 ( .A(c1478), .B(b[1478]), .Z(n4435) );
XNOR U7393 ( .A(b[1478]), .B(n4436), .Z(c[1478]) );
XNOR U7394 ( .A(a[1478]), .B(c1478), .Z(n4436) );
XOR U7395 ( .A(c1479), .B(n4437), .Z(c1480) );
ANDN U7396 ( .B(n4438), .A(n4439), .Z(n4437) );
XOR U7397 ( .A(c1479), .B(b[1479]), .Z(n4438) );
XNOR U7398 ( .A(b[1479]), .B(n4439), .Z(c[1479]) );
XNOR U7399 ( .A(a[1479]), .B(c1479), .Z(n4439) );
XOR U7400 ( .A(c1480), .B(n4440), .Z(c1481) );
ANDN U7401 ( .B(n4441), .A(n4442), .Z(n4440) );
XOR U7402 ( .A(c1480), .B(b[1480]), .Z(n4441) );
XNOR U7403 ( .A(b[1480]), .B(n4442), .Z(c[1480]) );
XNOR U7404 ( .A(a[1480]), .B(c1480), .Z(n4442) );
XOR U7405 ( .A(c1481), .B(n4443), .Z(c1482) );
ANDN U7406 ( .B(n4444), .A(n4445), .Z(n4443) );
XOR U7407 ( .A(c1481), .B(b[1481]), .Z(n4444) );
XNOR U7408 ( .A(b[1481]), .B(n4445), .Z(c[1481]) );
XNOR U7409 ( .A(a[1481]), .B(c1481), .Z(n4445) );
XOR U7410 ( .A(c1482), .B(n4446), .Z(c1483) );
ANDN U7411 ( .B(n4447), .A(n4448), .Z(n4446) );
XOR U7412 ( .A(c1482), .B(b[1482]), .Z(n4447) );
XNOR U7413 ( .A(b[1482]), .B(n4448), .Z(c[1482]) );
XNOR U7414 ( .A(a[1482]), .B(c1482), .Z(n4448) );
XOR U7415 ( .A(c1483), .B(n4449), .Z(c1484) );
ANDN U7416 ( .B(n4450), .A(n4451), .Z(n4449) );
XOR U7417 ( .A(c1483), .B(b[1483]), .Z(n4450) );
XNOR U7418 ( .A(b[1483]), .B(n4451), .Z(c[1483]) );
XNOR U7419 ( .A(a[1483]), .B(c1483), .Z(n4451) );
XOR U7420 ( .A(c1484), .B(n4452), .Z(c1485) );
ANDN U7421 ( .B(n4453), .A(n4454), .Z(n4452) );
XOR U7422 ( .A(c1484), .B(b[1484]), .Z(n4453) );
XNOR U7423 ( .A(b[1484]), .B(n4454), .Z(c[1484]) );
XNOR U7424 ( .A(a[1484]), .B(c1484), .Z(n4454) );
XOR U7425 ( .A(c1485), .B(n4455), .Z(c1486) );
ANDN U7426 ( .B(n4456), .A(n4457), .Z(n4455) );
XOR U7427 ( .A(c1485), .B(b[1485]), .Z(n4456) );
XNOR U7428 ( .A(b[1485]), .B(n4457), .Z(c[1485]) );
XNOR U7429 ( .A(a[1485]), .B(c1485), .Z(n4457) );
XOR U7430 ( .A(c1486), .B(n4458), .Z(c1487) );
ANDN U7431 ( .B(n4459), .A(n4460), .Z(n4458) );
XOR U7432 ( .A(c1486), .B(b[1486]), .Z(n4459) );
XNOR U7433 ( .A(b[1486]), .B(n4460), .Z(c[1486]) );
XNOR U7434 ( .A(a[1486]), .B(c1486), .Z(n4460) );
XOR U7435 ( .A(c1487), .B(n4461), .Z(c1488) );
ANDN U7436 ( .B(n4462), .A(n4463), .Z(n4461) );
XOR U7437 ( .A(c1487), .B(b[1487]), .Z(n4462) );
XNOR U7438 ( .A(b[1487]), .B(n4463), .Z(c[1487]) );
XNOR U7439 ( .A(a[1487]), .B(c1487), .Z(n4463) );
XOR U7440 ( .A(c1488), .B(n4464), .Z(c1489) );
ANDN U7441 ( .B(n4465), .A(n4466), .Z(n4464) );
XOR U7442 ( .A(c1488), .B(b[1488]), .Z(n4465) );
XNOR U7443 ( .A(b[1488]), .B(n4466), .Z(c[1488]) );
XNOR U7444 ( .A(a[1488]), .B(c1488), .Z(n4466) );
XOR U7445 ( .A(c1489), .B(n4467), .Z(c1490) );
ANDN U7446 ( .B(n4468), .A(n4469), .Z(n4467) );
XOR U7447 ( .A(c1489), .B(b[1489]), .Z(n4468) );
XNOR U7448 ( .A(b[1489]), .B(n4469), .Z(c[1489]) );
XNOR U7449 ( .A(a[1489]), .B(c1489), .Z(n4469) );
XOR U7450 ( .A(c1490), .B(n4470), .Z(c1491) );
ANDN U7451 ( .B(n4471), .A(n4472), .Z(n4470) );
XOR U7452 ( .A(c1490), .B(b[1490]), .Z(n4471) );
XNOR U7453 ( .A(b[1490]), .B(n4472), .Z(c[1490]) );
XNOR U7454 ( .A(a[1490]), .B(c1490), .Z(n4472) );
XOR U7455 ( .A(c1491), .B(n4473), .Z(c1492) );
ANDN U7456 ( .B(n4474), .A(n4475), .Z(n4473) );
XOR U7457 ( .A(c1491), .B(b[1491]), .Z(n4474) );
XNOR U7458 ( .A(b[1491]), .B(n4475), .Z(c[1491]) );
XNOR U7459 ( .A(a[1491]), .B(c1491), .Z(n4475) );
XOR U7460 ( .A(c1492), .B(n4476), .Z(c1493) );
ANDN U7461 ( .B(n4477), .A(n4478), .Z(n4476) );
XOR U7462 ( .A(c1492), .B(b[1492]), .Z(n4477) );
XNOR U7463 ( .A(b[1492]), .B(n4478), .Z(c[1492]) );
XNOR U7464 ( .A(a[1492]), .B(c1492), .Z(n4478) );
XOR U7465 ( .A(c1493), .B(n4479), .Z(c1494) );
ANDN U7466 ( .B(n4480), .A(n4481), .Z(n4479) );
XOR U7467 ( .A(c1493), .B(b[1493]), .Z(n4480) );
XNOR U7468 ( .A(b[1493]), .B(n4481), .Z(c[1493]) );
XNOR U7469 ( .A(a[1493]), .B(c1493), .Z(n4481) );
XOR U7470 ( .A(c1494), .B(n4482), .Z(c1495) );
ANDN U7471 ( .B(n4483), .A(n4484), .Z(n4482) );
XOR U7472 ( .A(c1494), .B(b[1494]), .Z(n4483) );
XNOR U7473 ( .A(b[1494]), .B(n4484), .Z(c[1494]) );
XNOR U7474 ( .A(a[1494]), .B(c1494), .Z(n4484) );
XOR U7475 ( .A(c1495), .B(n4485), .Z(c1496) );
ANDN U7476 ( .B(n4486), .A(n4487), .Z(n4485) );
XOR U7477 ( .A(c1495), .B(b[1495]), .Z(n4486) );
XNOR U7478 ( .A(b[1495]), .B(n4487), .Z(c[1495]) );
XNOR U7479 ( .A(a[1495]), .B(c1495), .Z(n4487) );
XOR U7480 ( .A(c1496), .B(n4488), .Z(c1497) );
ANDN U7481 ( .B(n4489), .A(n4490), .Z(n4488) );
XOR U7482 ( .A(c1496), .B(b[1496]), .Z(n4489) );
XNOR U7483 ( .A(b[1496]), .B(n4490), .Z(c[1496]) );
XNOR U7484 ( .A(a[1496]), .B(c1496), .Z(n4490) );
XOR U7485 ( .A(c1497), .B(n4491), .Z(c1498) );
ANDN U7486 ( .B(n4492), .A(n4493), .Z(n4491) );
XOR U7487 ( .A(c1497), .B(b[1497]), .Z(n4492) );
XNOR U7488 ( .A(b[1497]), .B(n4493), .Z(c[1497]) );
XNOR U7489 ( .A(a[1497]), .B(c1497), .Z(n4493) );
XOR U7490 ( .A(c1498), .B(n4494), .Z(c1499) );
ANDN U7491 ( .B(n4495), .A(n4496), .Z(n4494) );
XOR U7492 ( .A(c1498), .B(b[1498]), .Z(n4495) );
XNOR U7493 ( .A(b[1498]), .B(n4496), .Z(c[1498]) );
XNOR U7494 ( .A(a[1498]), .B(c1498), .Z(n4496) );
XOR U7495 ( .A(c1499), .B(n4497), .Z(c1500) );
ANDN U7496 ( .B(n4498), .A(n4499), .Z(n4497) );
XOR U7497 ( .A(c1499), .B(b[1499]), .Z(n4498) );
XNOR U7498 ( .A(b[1499]), .B(n4499), .Z(c[1499]) );
XNOR U7499 ( .A(a[1499]), .B(c1499), .Z(n4499) );
XOR U7500 ( .A(c1500), .B(n4500), .Z(c1501) );
ANDN U7501 ( .B(n4501), .A(n4502), .Z(n4500) );
XOR U7502 ( .A(c1500), .B(b[1500]), .Z(n4501) );
XNOR U7503 ( .A(b[1500]), .B(n4502), .Z(c[1500]) );
XNOR U7504 ( .A(a[1500]), .B(c1500), .Z(n4502) );
XOR U7505 ( .A(c1501), .B(n4503), .Z(c1502) );
ANDN U7506 ( .B(n4504), .A(n4505), .Z(n4503) );
XOR U7507 ( .A(c1501), .B(b[1501]), .Z(n4504) );
XNOR U7508 ( .A(b[1501]), .B(n4505), .Z(c[1501]) );
XNOR U7509 ( .A(a[1501]), .B(c1501), .Z(n4505) );
XOR U7510 ( .A(c1502), .B(n4506), .Z(c1503) );
ANDN U7511 ( .B(n4507), .A(n4508), .Z(n4506) );
XOR U7512 ( .A(c1502), .B(b[1502]), .Z(n4507) );
XNOR U7513 ( .A(b[1502]), .B(n4508), .Z(c[1502]) );
XNOR U7514 ( .A(a[1502]), .B(c1502), .Z(n4508) );
XOR U7515 ( .A(c1503), .B(n4509), .Z(c1504) );
ANDN U7516 ( .B(n4510), .A(n4511), .Z(n4509) );
XOR U7517 ( .A(c1503), .B(b[1503]), .Z(n4510) );
XNOR U7518 ( .A(b[1503]), .B(n4511), .Z(c[1503]) );
XNOR U7519 ( .A(a[1503]), .B(c1503), .Z(n4511) );
XOR U7520 ( .A(c1504), .B(n4512), .Z(c1505) );
ANDN U7521 ( .B(n4513), .A(n4514), .Z(n4512) );
XOR U7522 ( .A(c1504), .B(b[1504]), .Z(n4513) );
XNOR U7523 ( .A(b[1504]), .B(n4514), .Z(c[1504]) );
XNOR U7524 ( .A(a[1504]), .B(c1504), .Z(n4514) );
XOR U7525 ( .A(c1505), .B(n4515), .Z(c1506) );
ANDN U7526 ( .B(n4516), .A(n4517), .Z(n4515) );
XOR U7527 ( .A(c1505), .B(b[1505]), .Z(n4516) );
XNOR U7528 ( .A(b[1505]), .B(n4517), .Z(c[1505]) );
XNOR U7529 ( .A(a[1505]), .B(c1505), .Z(n4517) );
XOR U7530 ( .A(c1506), .B(n4518), .Z(c1507) );
ANDN U7531 ( .B(n4519), .A(n4520), .Z(n4518) );
XOR U7532 ( .A(c1506), .B(b[1506]), .Z(n4519) );
XNOR U7533 ( .A(b[1506]), .B(n4520), .Z(c[1506]) );
XNOR U7534 ( .A(a[1506]), .B(c1506), .Z(n4520) );
XOR U7535 ( .A(c1507), .B(n4521), .Z(c1508) );
ANDN U7536 ( .B(n4522), .A(n4523), .Z(n4521) );
XOR U7537 ( .A(c1507), .B(b[1507]), .Z(n4522) );
XNOR U7538 ( .A(b[1507]), .B(n4523), .Z(c[1507]) );
XNOR U7539 ( .A(a[1507]), .B(c1507), .Z(n4523) );
XOR U7540 ( .A(c1508), .B(n4524), .Z(c1509) );
ANDN U7541 ( .B(n4525), .A(n4526), .Z(n4524) );
XOR U7542 ( .A(c1508), .B(b[1508]), .Z(n4525) );
XNOR U7543 ( .A(b[1508]), .B(n4526), .Z(c[1508]) );
XNOR U7544 ( .A(a[1508]), .B(c1508), .Z(n4526) );
XOR U7545 ( .A(c1509), .B(n4527), .Z(c1510) );
ANDN U7546 ( .B(n4528), .A(n4529), .Z(n4527) );
XOR U7547 ( .A(c1509), .B(b[1509]), .Z(n4528) );
XNOR U7548 ( .A(b[1509]), .B(n4529), .Z(c[1509]) );
XNOR U7549 ( .A(a[1509]), .B(c1509), .Z(n4529) );
XOR U7550 ( .A(c1510), .B(n4530), .Z(c1511) );
ANDN U7551 ( .B(n4531), .A(n4532), .Z(n4530) );
XOR U7552 ( .A(c1510), .B(b[1510]), .Z(n4531) );
XNOR U7553 ( .A(b[1510]), .B(n4532), .Z(c[1510]) );
XNOR U7554 ( .A(a[1510]), .B(c1510), .Z(n4532) );
XOR U7555 ( .A(c1511), .B(n4533), .Z(c1512) );
ANDN U7556 ( .B(n4534), .A(n4535), .Z(n4533) );
XOR U7557 ( .A(c1511), .B(b[1511]), .Z(n4534) );
XNOR U7558 ( .A(b[1511]), .B(n4535), .Z(c[1511]) );
XNOR U7559 ( .A(a[1511]), .B(c1511), .Z(n4535) );
XOR U7560 ( .A(c1512), .B(n4536), .Z(c1513) );
ANDN U7561 ( .B(n4537), .A(n4538), .Z(n4536) );
XOR U7562 ( .A(c1512), .B(b[1512]), .Z(n4537) );
XNOR U7563 ( .A(b[1512]), .B(n4538), .Z(c[1512]) );
XNOR U7564 ( .A(a[1512]), .B(c1512), .Z(n4538) );
XOR U7565 ( .A(c1513), .B(n4539), .Z(c1514) );
ANDN U7566 ( .B(n4540), .A(n4541), .Z(n4539) );
XOR U7567 ( .A(c1513), .B(b[1513]), .Z(n4540) );
XNOR U7568 ( .A(b[1513]), .B(n4541), .Z(c[1513]) );
XNOR U7569 ( .A(a[1513]), .B(c1513), .Z(n4541) );
XOR U7570 ( .A(c1514), .B(n4542), .Z(c1515) );
ANDN U7571 ( .B(n4543), .A(n4544), .Z(n4542) );
XOR U7572 ( .A(c1514), .B(b[1514]), .Z(n4543) );
XNOR U7573 ( .A(b[1514]), .B(n4544), .Z(c[1514]) );
XNOR U7574 ( .A(a[1514]), .B(c1514), .Z(n4544) );
XOR U7575 ( .A(c1515), .B(n4545), .Z(c1516) );
ANDN U7576 ( .B(n4546), .A(n4547), .Z(n4545) );
XOR U7577 ( .A(c1515), .B(b[1515]), .Z(n4546) );
XNOR U7578 ( .A(b[1515]), .B(n4547), .Z(c[1515]) );
XNOR U7579 ( .A(a[1515]), .B(c1515), .Z(n4547) );
XOR U7580 ( .A(c1516), .B(n4548), .Z(c1517) );
ANDN U7581 ( .B(n4549), .A(n4550), .Z(n4548) );
XOR U7582 ( .A(c1516), .B(b[1516]), .Z(n4549) );
XNOR U7583 ( .A(b[1516]), .B(n4550), .Z(c[1516]) );
XNOR U7584 ( .A(a[1516]), .B(c1516), .Z(n4550) );
XOR U7585 ( .A(c1517), .B(n4551), .Z(c1518) );
ANDN U7586 ( .B(n4552), .A(n4553), .Z(n4551) );
XOR U7587 ( .A(c1517), .B(b[1517]), .Z(n4552) );
XNOR U7588 ( .A(b[1517]), .B(n4553), .Z(c[1517]) );
XNOR U7589 ( .A(a[1517]), .B(c1517), .Z(n4553) );
XOR U7590 ( .A(c1518), .B(n4554), .Z(c1519) );
ANDN U7591 ( .B(n4555), .A(n4556), .Z(n4554) );
XOR U7592 ( .A(c1518), .B(b[1518]), .Z(n4555) );
XNOR U7593 ( .A(b[1518]), .B(n4556), .Z(c[1518]) );
XNOR U7594 ( .A(a[1518]), .B(c1518), .Z(n4556) );
XOR U7595 ( .A(c1519), .B(n4557), .Z(c1520) );
ANDN U7596 ( .B(n4558), .A(n4559), .Z(n4557) );
XOR U7597 ( .A(c1519), .B(b[1519]), .Z(n4558) );
XNOR U7598 ( .A(b[1519]), .B(n4559), .Z(c[1519]) );
XNOR U7599 ( .A(a[1519]), .B(c1519), .Z(n4559) );
XOR U7600 ( .A(c1520), .B(n4560), .Z(c1521) );
ANDN U7601 ( .B(n4561), .A(n4562), .Z(n4560) );
XOR U7602 ( .A(c1520), .B(b[1520]), .Z(n4561) );
XNOR U7603 ( .A(b[1520]), .B(n4562), .Z(c[1520]) );
XNOR U7604 ( .A(a[1520]), .B(c1520), .Z(n4562) );
XOR U7605 ( .A(c1521), .B(n4563), .Z(c1522) );
ANDN U7606 ( .B(n4564), .A(n4565), .Z(n4563) );
XOR U7607 ( .A(c1521), .B(b[1521]), .Z(n4564) );
XNOR U7608 ( .A(b[1521]), .B(n4565), .Z(c[1521]) );
XNOR U7609 ( .A(a[1521]), .B(c1521), .Z(n4565) );
XOR U7610 ( .A(c1522), .B(n4566), .Z(c1523) );
ANDN U7611 ( .B(n4567), .A(n4568), .Z(n4566) );
XOR U7612 ( .A(c1522), .B(b[1522]), .Z(n4567) );
XNOR U7613 ( .A(b[1522]), .B(n4568), .Z(c[1522]) );
XNOR U7614 ( .A(a[1522]), .B(c1522), .Z(n4568) );
XOR U7615 ( .A(c1523), .B(n4569), .Z(c1524) );
ANDN U7616 ( .B(n4570), .A(n4571), .Z(n4569) );
XOR U7617 ( .A(c1523), .B(b[1523]), .Z(n4570) );
XNOR U7618 ( .A(b[1523]), .B(n4571), .Z(c[1523]) );
XNOR U7619 ( .A(a[1523]), .B(c1523), .Z(n4571) );
XOR U7620 ( .A(c1524), .B(n4572), .Z(c1525) );
ANDN U7621 ( .B(n4573), .A(n4574), .Z(n4572) );
XOR U7622 ( .A(c1524), .B(b[1524]), .Z(n4573) );
XNOR U7623 ( .A(b[1524]), .B(n4574), .Z(c[1524]) );
XNOR U7624 ( .A(a[1524]), .B(c1524), .Z(n4574) );
XOR U7625 ( .A(c1525), .B(n4575), .Z(c1526) );
ANDN U7626 ( .B(n4576), .A(n4577), .Z(n4575) );
XOR U7627 ( .A(c1525), .B(b[1525]), .Z(n4576) );
XNOR U7628 ( .A(b[1525]), .B(n4577), .Z(c[1525]) );
XNOR U7629 ( .A(a[1525]), .B(c1525), .Z(n4577) );
XOR U7630 ( .A(c1526), .B(n4578), .Z(c1527) );
ANDN U7631 ( .B(n4579), .A(n4580), .Z(n4578) );
XOR U7632 ( .A(c1526), .B(b[1526]), .Z(n4579) );
XNOR U7633 ( .A(b[1526]), .B(n4580), .Z(c[1526]) );
XNOR U7634 ( .A(a[1526]), .B(c1526), .Z(n4580) );
XOR U7635 ( .A(c1527), .B(n4581), .Z(c1528) );
ANDN U7636 ( .B(n4582), .A(n4583), .Z(n4581) );
XOR U7637 ( .A(c1527), .B(b[1527]), .Z(n4582) );
XNOR U7638 ( .A(b[1527]), .B(n4583), .Z(c[1527]) );
XNOR U7639 ( .A(a[1527]), .B(c1527), .Z(n4583) );
XOR U7640 ( .A(c1528), .B(n4584), .Z(c1529) );
ANDN U7641 ( .B(n4585), .A(n4586), .Z(n4584) );
XOR U7642 ( .A(c1528), .B(b[1528]), .Z(n4585) );
XNOR U7643 ( .A(b[1528]), .B(n4586), .Z(c[1528]) );
XNOR U7644 ( .A(a[1528]), .B(c1528), .Z(n4586) );
XOR U7645 ( .A(c1529), .B(n4587), .Z(c1530) );
ANDN U7646 ( .B(n4588), .A(n4589), .Z(n4587) );
XOR U7647 ( .A(c1529), .B(b[1529]), .Z(n4588) );
XNOR U7648 ( .A(b[1529]), .B(n4589), .Z(c[1529]) );
XNOR U7649 ( .A(a[1529]), .B(c1529), .Z(n4589) );
XOR U7650 ( .A(c1530), .B(n4590), .Z(c1531) );
ANDN U7651 ( .B(n4591), .A(n4592), .Z(n4590) );
XOR U7652 ( .A(c1530), .B(b[1530]), .Z(n4591) );
XNOR U7653 ( .A(b[1530]), .B(n4592), .Z(c[1530]) );
XNOR U7654 ( .A(a[1530]), .B(c1530), .Z(n4592) );
XOR U7655 ( .A(c1531), .B(n4593), .Z(c1532) );
ANDN U7656 ( .B(n4594), .A(n4595), .Z(n4593) );
XOR U7657 ( .A(c1531), .B(b[1531]), .Z(n4594) );
XNOR U7658 ( .A(b[1531]), .B(n4595), .Z(c[1531]) );
XNOR U7659 ( .A(a[1531]), .B(c1531), .Z(n4595) );
XOR U7660 ( .A(c1532), .B(n4596), .Z(c1533) );
ANDN U7661 ( .B(n4597), .A(n4598), .Z(n4596) );
XOR U7662 ( .A(c1532), .B(b[1532]), .Z(n4597) );
XNOR U7663 ( .A(b[1532]), .B(n4598), .Z(c[1532]) );
XNOR U7664 ( .A(a[1532]), .B(c1532), .Z(n4598) );
XOR U7665 ( .A(c1533), .B(n4599), .Z(c1534) );
ANDN U7666 ( .B(n4600), .A(n4601), .Z(n4599) );
XOR U7667 ( .A(c1533), .B(b[1533]), .Z(n4600) );
XNOR U7668 ( .A(b[1533]), .B(n4601), .Z(c[1533]) );
XNOR U7669 ( .A(a[1533]), .B(c1533), .Z(n4601) );
XOR U7670 ( .A(c1534), .B(n4602), .Z(c1535) );
ANDN U7671 ( .B(n4603), .A(n4604), .Z(n4602) );
XOR U7672 ( .A(c1534), .B(b[1534]), .Z(n4603) );
XNOR U7673 ( .A(b[1534]), .B(n4604), .Z(c[1534]) );
XNOR U7674 ( .A(a[1534]), .B(c1534), .Z(n4604) );
XOR U7675 ( .A(c1535), .B(n4605), .Z(c1536) );
ANDN U7676 ( .B(n4606), .A(n4607), .Z(n4605) );
XOR U7677 ( .A(c1535), .B(b[1535]), .Z(n4606) );
XNOR U7678 ( .A(b[1535]), .B(n4607), .Z(c[1535]) );
XNOR U7679 ( .A(a[1535]), .B(c1535), .Z(n4607) );
XOR U7680 ( .A(c1536), .B(n4608), .Z(c1537) );
ANDN U7681 ( .B(n4609), .A(n4610), .Z(n4608) );
XOR U7682 ( .A(c1536), .B(b[1536]), .Z(n4609) );
XNOR U7683 ( .A(b[1536]), .B(n4610), .Z(c[1536]) );
XNOR U7684 ( .A(a[1536]), .B(c1536), .Z(n4610) );
XOR U7685 ( .A(c1537), .B(n4611), .Z(c1538) );
ANDN U7686 ( .B(n4612), .A(n4613), .Z(n4611) );
XOR U7687 ( .A(c1537), .B(b[1537]), .Z(n4612) );
XNOR U7688 ( .A(b[1537]), .B(n4613), .Z(c[1537]) );
XNOR U7689 ( .A(a[1537]), .B(c1537), .Z(n4613) );
XOR U7690 ( .A(c1538), .B(n4614), .Z(c1539) );
ANDN U7691 ( .B(n4615), .A(n4616), .Z(n4614) );
XOR U7692 ( .A(c1538), .B(b[1538]), .Z(n4615) );
XNOR U7693 ( .A(b[1538]), .B(n4616), .Z(c[1538]) );
XNOR U7694 ( .A(a[1538]), .B(c1538), .Z(n4616) );
XOR U7695 ( .A(c1539), .B(n4617), .Z(c1540) );
ANDN U7696 ( .B(n4618), .A(n4619), .Z(n4617) );
XOR U7697 ( .A(c1539), .B(b[1539]), .Z(n4618) );
XNOR U7698 ( .A(b[1539]), .B(n4619), .Z(c[1539]) );
XNOR U7699 ( .A(a[1539]), .B(c1539), .Z(n4619) );
XOR U7700 ( .A(c1540), .B(n4620), .Z(c1541) );
ANDN U7701 ( .B(n4621), .A(n4622), .Z(n4620) );
XOR U7702 ( .A(c1540), .B(b[1540]), .Z(n4621) );
XNOR U7703 ( .A(b[1540]), .B(n4622), .Z(c[1540]) );
XNOR U7704 ( .A(a[1540]), .B(c1540), .Z(n4622) );
XOR U7705 ( .A(c1541), .B(n4623), .Z(c1542) );
ANDN U7706 ( .B(n4624), .A(n4625), .Z(n4623) );
XOR U7707 ( .A(c1541), .B(b[1541]), .Z(n4624) );
XNOR U7708 ( .A(b[1541]), .B(n4625), .Z(c[1541]) );
XNOR U7709 ( .A(a[1541]), .B(c1541), .Z(n4625) );
XOR U7710 ( .A(c1542), .B(n4626), .Z(c1543) );
ANDN U7711 ( .B(n4627), .A(n4628), .Z(n4626) );
XOR U7712 ( .A(c1542), .B(b[1542]), .Z(n4627) );
XNOR U7713 ( .A(b[1542]), .B(n4628), .Z(c[1542]) );
XNOR U7714 ( .A(a[1542]), .B(c1542), .Z(n4628) );
XOR U7715 ( .A(c1543), .B(n4629), .Z(c1544) );
ANDN U7716 ( .B(n4630), .A(n4631), .Z(n4629) );
XOR U7717 ( .A(c1543), .B(b[1543]), .Z(n4630) );
XNOR U7718 ( .A(b[1543]), .B(n4631), .Z(c[1543]) );
XNOR U7719 ( .A(a[1543]), .B(c1543), .Z(n4631) );
XOR U7720 ( .A(c1544), .B(n4632), .Z(c1545) );
ANDN U7721 ( .B(n4633), .A(n4634), .Z(n4632) );
XOR U7722 ( .A(c1544), .B(b[1544]), .Z(n4633) );
XNOR U7723 ( .A(b[1544]), .B(n4634), .Z(c[1544]) );
XNOR U7724 ( .A(a[1544]), .B(c1544), .Z(n4634) );
XOR U7725 ( .A(c1545), .B(n4635), .Z(c1546) );
ANDN U7726 ( .B(n4636), .A(n4637), .Z(n4635) );
XOR U7727 ( .A(c1545), .B(b[1545]), .Z(n4636) );
XNOR U7728 ( .A(b[1545]), .B(n4637), .Z(c[1545]) );
XNOR U7729 ( .A(a[1545]), .B(c1545), .Z(n4637) );
XOR U7730 ( .A(c1546), .B(n4638), .Z(c1547) );
ANDN U7731 ( .B(n4639), .A(n4640), .Z(n4638) );
XOR U7732 ( .A(c1546), .B(b[1546]), .Z(n4639) );
XNOR U7733 ( .A(b[1546]), .B(n4640), .Z(c[1546]) );
XNOR U7734 ( .A(a[1546]), .B(c1546), .Z(n4640) );
XOR U7735 ( .A(c1547), .B(n4641), .Z(c1548) );
ANDN U7736 ( .B(n4642), .A(n4643), .Z(n4641) );
XOR U7737 ( .A(c1547), .B(b[1547]), .Z(n4642) );
XNOR U7738 ( .A(b[1547]), .B(n4643), .Z(c[1547]) );
XNOR U7739 ( .A(a[1547]), .B(c1547), .Z(n4643) );
XOR U7740 ( .A(c1548), .B(n4644), .Z(c1549) );
ANDN U7741 ( .B(n4645), .A(n4646), .Z(n4644) );
XOR U7742 ( .A(c1548), .B(b[1548]), .Z(n4645) );
XNOR U7743 ( .A(b[1548]), .B(n4646), .Z(c[1548]) );
XNOR U7744 ( .A(a[1548]), .B(c1548), .Z(n4646) );
XOR U7745 ( .A(c1549), .B(n4647), .Z(c1550) );
ANDN U7746 ( .B(n4648), .A(n4649), .Z(n4647) );
XOR U7747 ( .A(c1549), .B(b[1549]), .Z(n4648) );
XNOR U7748 ( .A(b[1549]), .B(n4649), .Z(c[1549]) );
XNOR U7749 ( .A(a[1549]), .B(c1549), .Z(n4649) );
XOR U7750 ( .A(c1550), .B(n4650), .Z(c1551) );
ANDN U7751 ( .B(n4651), .A(n4652), .Z(n4650) );
XOR U7752 ( .A(c1550), .B(b[1550]), .Z(n4651) );
XNOR U7753 ( .A(b[1550]), .B(n4652), .Z(c[1550]) );
XNOR U7754 ( .A(a[1550]), .B(c1550), .Z(n4652) );
XOR U7755 ( .A(c1551), .B(n4653), .Z(c1552) );
ANDN U7756 ( .B(n4654), .A(n4655), .Z(n4653) );
XOR U7757 ( .A(c1551), .B(b[1551]), .Z(n4654) );
XNOR U7758 ( .A(b[1551]), .B(n4655), .Z(c[1551]) );
XNOR U7759 ( .A(a[1551]), .B(c1551), .Z(n4655) );
XOR U7760 ( .A(c1552), .B(n4656), .Z(c1553) );
ANDN U7761 ( .B(n4657), .A(n4658), .Z(n4656) );
XOR U7762 ( .A(c1552), .B(b[1552]), .Z(n4657) );
XNOR U7763 ( .A(b[1552]), .B(n4658), .Z(c[1552]) );
XNOR U7764 ( .A(a[1552]), .B(c1552), .Z(n4658) );
XOR U7765 ( .A(c1553), .B(n4659), .Z(c1554) );
ANDN U7766 ( .B(n4660), .A(n4661), .Z(n4659) );
XOR U7767 ( .A(c1553), .B(b[1553]), .Z(n4660) );
XNOR U7768 ( .A(b[1553]), .B(n4661), .Z(c[1553]) );
XNOR U7769 ( .A(a[1553]), .B(c1553), .Z(n4661) );
XOR U7770 ( .A(c1554), .B(n4662), .Z(c1555) );
ANDN U7771 ( .B(n4663), .A(n4664), .Z(n4662) );
XOR U7772 ( .A(c1554), .B(b[1554]), .Z(n4663) );
XNOR U7773 ( .A(b[1554]), .B(n4664), .Z(c[1554]) );
XNOR U7774 ( .A(a[1554]), .B(c1554), .Z(n4664) );
XOR U7775 ( .A(c1555), .B(n4665), .Z(c1556) );
ANDN U7776 ( .B(n4666), .A(n4667), .Z(n4665) );
XOR U7777 ( .A(c1555), .B(b[1555]), .Z(n4666) );
XNOR U7778 ( .A(b[1555]), .B(n4667), .Z(c[1555]) );
XNOR U7779 ( .A(a[1555]), .B(c1555), .Z(n4667) );
XOR U7780 ( .A(c1556), .B(n4668), .Z(c1557) );
ANDN U7781 ( .B(n4669), .A(n4670), .Z(n4668) );
XOR U7782 ( .A(c1556), .B(b[1556]), .Z(n4669) );
XNOR U7783 ( .A(b[1556]), .B(n4670), .Z(c[1556]) );
XNOR U7784 ( .A(a[1556]), .B(c1556), .Z(n4670) );
XOR U7785 ( .A(c1557), .B(n4671), .Z(c1558) );
ANDN U7786 ( .B(n4672), .A(n4673), .Z(n4671) );
XOR U7787 ( .A(c1557), .B(b[1557]), .Z(n4672) );
XNOR U7788 ( .A(b[1557]), .B(n4673), .Z(c[1557]) );
XNOR U7789 ( .A(a[1557]), .B(c1557), .Z(n4673) );
XOR U7790 ( .A(c1558), .B(n4674), .Z(c1559) );
ANDN U7791 ( .B(n4675), .A(n4676), .Z(n4674) );
XOR U7792 ( .A(c1558), .B(b[1558]), .Z(n4675) );
XNOR U7793 ( .A(b[1558]), .B(n4676), .Z(c[1558]) );
XNOR U7794 ( .A(a[1558]), .B(c1558), .Z(n4676) );
XOR U7795 ( .A(c1559), .B(n4677), .Z(c1560) );
ANDN U7796 ( .B(n4678), .A(n4679), .Z(n4677) );
XOR U7797 ( .A(c1559), .B(b[1559]), .Z(n4678) );
XNOR U7798 ( .A(b[1559]), .B(n4679), .Z(c[1559]) );
XNOR U7799 ( .A(a[1559]), .B(c1559), .Z(n4679) );
XOR U7800 ( .A(c1560), .B(n4680), .Z(c1561) );
ANDN U7801 ( .B(n4681), .A(n4682), .Z(n4680) );
XOR U7802 ( .A(c1560), .B(b[1560]), .Z(n4681) );
XNOR U7803 ( .A(b[1560]), .B(n4682), .Z(c[1560]) );
XNOR U7804 ( .A(a[1560]), .B(c1560), .Z(n4682) );
XOR U7805 ( .A(c1561), .B(n4683), .Z(c1562) );
ANDN U7806 ( .B(n4684), .A(n4685), .Z(n4683) );
XOR U7807 ( .A(c1561), .B(b[1561]), .Z(n4684) );
XNOR U7808 ( .A(b[1561]), .B(n4685), .Z(c[1561]) );
XNOR U7809 ( .A(a[1561]), .B(c1561), .Z(n4685) );
XOR U7810 ( .A(c1562), .B(n4686), .Z(c1563) );
ANDN U7811 ( .B(n4687), .A(n4688), .Z(n4686) );
XOR U7812 ( .A(c1562), .B(b[1562]), .Z(n4687) );
XNOR U7813 ( .A(b[1562]), .B(n4688), .Z(c[1562]) );
XNOR U7814 ( .A(a[1562]), .B(c1562), .Z(n4688) );
XOR U7815 ( .A(c1563), .B(n4689), .Z(c1564) );
ANDN U7816 ( .B(n4690), .A(n4691), .Z(n4689) );
XOR U7817 ( .A(c1563), .B(b[1563]), .Z(n4690) );
XNOR U7818 ( .A(b[1563]), .B(n4691), .Z(c[1563]) );
XNOR U7819 ( .A(a[1563]), .B(c1563), .Z(n4691) );
XOR U7820 ( .A(c1564), .B(n4692), .Z(c1565) );
ANDN U7821 ( .B(n4693), .A(n4694), .Z(n4692) );
XOR U7822 ( .A(c1564), .B(b[1564]), .Z(n4693) );
XNOR U7823 ( .A(b[1564]), .B(n4694), .Z(c[1564]) );
XNOR U7824 ( .A(a[1564]), .B(c1564), .Z(n4694) );
XOR U7825 ( .A(c1565), .B(n4695), .Z(c1566) );
ANDN U7826 ( .B(n4696), .A(n4697), .Z(n4695) );
XOR U7827 ( .A(c1565), .B(b[1565]), .Z(n4696) );
XNOR U7828 ( .A(b[1565]), .B(n4697), .Z(c[1565]) );
XNOR U7829 ( .A(a[1565]), .B(c1565), .Z(n4697) );
XOR U7830 ( .A(c1566), .B(n4698), .Z(c1567) );
ANDN U7831 ( .B(n4699), .A(n4700), .Z(n4698) );
XOR U7832 ( .A(c1566), .B(b[1566]), .Z(n4699) );
XNOR U7833 ( .A(b[1566]), .B(n4700), .Z(c[1566]) );
XNOR U7834 ( .A(a[1566]), .B(c1566), .Z(n4700) );
XOR U7835 ( .A(c1567), .B(n4701), .Z(c1568) );
ANDN U7836 ( .B(n4702), .A(n4703), .Z(n4701) );
XOR U7837 ( .A(c1567), .B(b[1567]), .Z(n4702) );
XNOR U7838 ( .A(b[1567]), .B(n4703), .Z(c[1567]) );
XNOR U7839 ( .A(a[1567]), .B(c1567), .Z(n4703) );
XOR U7840 ( .A(c1568), .B(n4704), .Z(c1569) );
ANDN U7841 ( .B(n4705), .A(n4706), .Z(n4704) );
XOR U7842 ( .A(c1568), .B(b[1568]), .Z(n4705) );
XNOR U7843 ( .A(b[1568]), .B(n4706), .Z(c[1568]) );
XNOR U7844 ( .A(a[1568]), .B(c1568), .Z(n4706) );
XOR U7845 ( .A(c1569), .B(n4707), .Z(c1570) );
ANDN U7846 ( .B(n4708), .A(n4709), .Z(n4707) );
XOR U7847 ( .A(c1569), .B(b[1569]), .Z(n4708) );
XNOR U7848 ( .A(b[1569]), .B(n4709), .Z(c[1569]) );
XNOR U7849 ( .A(a[1569]), .B(c1569), .Z(n4709) );
XOR U7850 ( .A(c1570), .B(n4710), .Z(c1571) );
ANDN U7851 ( .B(n4711), .A(n4712), .Z(n4710) );
XOR U7852 ( .A(c1570), .B(b[1570]), .Z(n4711) );
XNOR U7853 ( .A(b[1570]), .B(n4712), .Z(c[1570]) );
XNOR U7854 ( .A(a[1570]), .B(c1570), .Z(n4712) );
XOR U7855 ( .A(c1571), .B(n4713), .Z(c1572) );
ANDN U7856 ( .B(n4714), .A(n4715), .Z(n4713) );
XOR U7857 ( .A(c1571), .B(b[1571]), .Z(n4714) );
XNOR U7858 ( .A(b[1571]), .B(n4715), .Z(c[1571]) );
XNOR U7859 ( .A(a[1571]), .B(c1571), .Z(n4715) );
XOR U7860 ( .A(c1572), .B(n4716), .Z(c1573) );
ANDN U7861 ( .B(n4717), .A(n4718), .Z(n4716) );
XOR U7862 ( .A(c1572), .B(b[1572]), .Z(n4717) );
XNOR U7863 ( .A(b[1572]), .B(n4718), .Z(c[1572]) );
XNOR U7864 ( .A(a[1572]), .B(c1572), .Z(n4718) );
XOR U7865 ( .A(c1573), .B(n4719), .Z(c1574) );
ANDN U7866 ( .B(n4720), .A(n4721), .Z(n4719) );
XOR U7867 ( .A(c1573), .B(b[1573]), .Z(n4720) );
XNOR U7868 ( .A(b[1573]), .B(n4721), .Z(c[1573]) );
XNOR U7869 ( .A(a[1573]), .B(c1573), .Z(n4721) );
XOR U7870 ( .A(c1574), .B(n4722), .Z(c1575) );
ANDN U7871 ( .B(n4723), .A(n4724), .Z(n4722) );
XOR U7872 ( .A(c1574), .B(b[1574]), .Z(n4723) );
XNOR U7873 ( .A(b[1574]), .B(n4724), .Z(c[1574]) );
XNOR U7874 ( .A(a[1574]), .B(c1574), .Z(n4724) );
XOR U7875 ( .A(c1575), .B(n4725), .Z(c1576) );
ANDN U7876 ( .B(n4726), .A(n4727), .Z(n4725) );
XOR U7877 ( .A(c1575), .B(b[1575]), .Z(n4726) );
XNOR U7878 ( .A(b[1575]), .B(n4727), .Z(c[1575]) );
XNOR U7879 ( .A(a[1575]), .B(c1575), .Z(n4727) );
XOR U7880 ( .A(c1576), .B(n4728), .Z(c1577) );
ANDN U7881 ( .B(n4729), .A(n4730), .Z(n4728) );
XOR U7882 ( .A(c1576), .B(b[1576]), .Z(n4729) );
XNOR U7883 ( .A(b[1576]), .B(n4730), .Z(c[1576]) );
XNOR U7884 ( .A(a[1576]), .B(c1576), .Z(n4730) );
XOR U7885 ( .A(c1577), .B(n4731), .Z(c1578) );
ANDN U7886 ( .B(n4732), .A(n4733), .Z(n4731) );
XOR U7887 ( .A(c1577), .B(b[1577]), .Z(n4732) );
XNOR U7888 ( .A(b[1577]), .B(n4733), .Z(c[1577]) );
XNOR U7889 ( .A(a[1577]), .B(c1577), .Z(n4733) );
XOR U7890 ( .A(c1578), .B(n4734), .Z(c1579) );
ANDN U7891 ( .B(n4735), .A(n4736), .Z(n4734) );
XOR U7892 ( .A(c1578), .B(b[1578]), .Z(n4735) );
XNOR U7893 ( .A(b[1578]), .B(n4736), .Z(c[1578]) );
XNOR U7894 ( .A(a[1578]), .B(c1578), .Z(n4736) );
XOR U7895 ( .A(c1579), .B(n4737), .Z(c1580) );
ANDN U7896 ( .B(n4738), .A(n4739), .Z(n4737) );
XOR U7897 ( .A(c1579), .B(b[1579]), .Z(n4738) );
XNOR U7898 ( .A(b[1579]), .B(n4739), .Z(c[1579]) );
XNOR U7899 ( .A(a[1579]), .B(c1579), .Z(n4739) );
XOR U7900 ( .A(c1580), .B(n4740), .Z(c1581) );
ANDN U7901 ( .B(n4741), .A(n4742), .Z(n4740) );
XOR U7902 ( .A(c1580), .B(b[1580]), .Z(n4741) );
XNOR U7903 ( .A(b[1580]), .B(n4742), .Z(c[1580]) );
XNOR U7904 ( .A(a[1580]), .B(c1580), .Z(n4742) );
XOR U7905 ( .A(c1581), .B(n4743), .Z(c1582) );
ANDN U7906 ( .B(n4744), .A(n4745), .Z(n4743) );
XOR U7907 ( .A(c1581), .B(b[1581]), .Z(n4744) );
XNOR U7908 ( .A(b[1581]), .B(n4745), .Z(c[1581]) );
XNOR U7909 ( .A(a[1581]), .B(c1581), .Z(n4745) );
XOR U7910 ( .A(c1582), .B(n4746), .Z(c1583) );
ANDN U7911 ( .B(n4747), .A(n4748), .Z(n4746) );
XOR U7912 ( .A(c1582), .B(b[1582]), .Z(n4747) );
XNOR U7913 ( .A(b[1582]), .B(n4748), .Z(c[1582]) );
XNOR U7914 ( .A(a[1582]), .B(c1582), .Z(n4748) );
XOR U7915 ( .A(c1583), .B(n4749), .Z(c1584) );
ANDN U7916 ( .B(n4750), .A(n4751), .Z(n4749) );
XOR U7917 ( .A(c1583), .B(b[1583]), .Z(n4750) );
XNOR U7918 ( .A(b[1583]), .B(n4751), .Z(c[1583]) );
XNOR U7919 ( .A(a[1583]), .B(c1583), .Z(n4751) );
XOR U7920 ( .A(c1584), .B(n4752), .Z(c1585) );
ANDN U7921 ( .B(n4753), .A(n4754), .Z(n4752) );
XOR U7922 ( .A(c1584), .B(b[1584]), .Z(n4753) );
XNOR U7923 ( .A(b[1584]), .B(n4754), .Z(c[1584]) );
XNOR U7924 ( .A(a[1584]), .B(c1584), .Z(n4754) );
XOR U7925 ( .A(c1585), .B(n4755), .Z(c1586) );
ANDN U7926 ( .B(n4756), .A(n4757), .Z(n4755) );
XOR U7927 ( .A(c1585), .B(b[1585]), .Z(n4756) );
XNOR U7928 ( .A(b[1585]), .B(n4757), .Z(c[1585]) );
XNOR U7929 ( .A(a[1585]), .B(c1585), .Z(n4757) );
XOR U7930 ( .A(c1586), .B(n4758), .Z(c1587) );
ANDN U7931 ( .B(n4759), .A(n4760), .Z(n4758) );
XOR U7932 ( .A(c1586), .B(b[1586]), .Z(n4759) );
XNOR U7933 ( .A(b[1586]), .B(n4760), .Z(c[1586]) );
XNOR U7934 ( .A(a[1586]), .B(c1586), .Z(n4760) );
XOR U7935 ( .A(c1587), .B(n4761), .Z(c1588) );
ANDN U7936 ( .B(n4762), .A(n4763), .Z(n4761) );
XOR U7937 ( .A(c1587), .B(b[1587]), .Z(n4762) );
XNOR U7938 ( .A(b[1587]), .B(n4763), .Z(c[1587]) );
XNOR U7939 ( .A(a[1587]), .B(c1587), .Z(n4763) );
XOR U7940 ( .A(c1588), .B(n4764), .Z(c1589) );
ANDN U7941 ( .B(n4765), .A(n4766), .Z(n4764) );
XOR U7942 ( .A(c1588), .B(b[1588]), .Z(n4765) );
XNOR U7943 ( .A(b[1588]), .B(n4766), .Z(c[1588]) );
XNOR U7944 ( .A(a[1588]), .B(c1588), .Z(n4766) );
XOR U7945 ( .A(c1589), .B(n4767), .Z(c1590) );
ANDN U7946 ( .B(n4768), .A(n4769), .Z(n4767) );
XOR U7947 ( .A(c1589), .B(b[1589]), .Z(n4768) );
XNOR U7948 ( .A(b[1589]), .B(n4769), .Z(c[1589]) );
XNOR U7949 ( .A(a[1589]), .B(c1589), .Z(n4769) );
XOR U7950 ( .A(c1590), .B(n4770), .Z(c1591) );
ANDN U7951 ( .B(n4771), .A(n4772), .Z(n4770) );
XOR U7952 ( .A(c1590), .B(b[1590]), .Z(n4771) );
XNOR U7953 ( .A(b[1590]), .B(n4772), .Z(c[1590]) );
XNOR U7954 ( .A(a[1590]), .B(c1590), .Z(n4772) );
XOR U7955 ( .A(c1591), .B(n4773), .Z(c1592) );
ANDN U7956 ( .B(n4774), .A(n4775), .Z(n4773) );
XOR U7957 ( .A(c1591), .B(b[1591]), .Z(n4774) );
XNOR U7958 ( .A(b[1591]), .B(n4775), .Z(c[1591]) );
XNOR U7959 ( .A(a[1591]), .B(c1591), .Z(n4775) );
XOR U7960 ( .A(c1592), .B(n4776), .Z(c1593) );
ANDN U7961 ( .B(n4777), .A(n4778), .Z(n4776) );
XOR U7962 ( .A(c1592), .B(b[1592]), .Z(n4777) );
XNOR U7963 ( .A(b[1592]), .B(n4778), .Z(c[1592]) );
XNOR U7964 ( .A(a[1592]), .B(c1592), .Z(n4778) );
XOR U7965 ( .A(c1593), .B(n4779), .Z(c1594) );
ANDN U7966 ( .B(n4780), .A(n4781), .Z(n4779) );
XOR U7967 ( .A(c1593), .B(b[1593]), .Z(n4780) );
XNOR U7968 ( .A(b[1593]), .B(n4781), .Z(c[1593]) );
XNOR U7969 ( .A(a[1593]), .B(c1593), .Z(n4781) );
XOR U7970 ( .A(c1594), .B(n4782), .Z(c1595) );
ANDN U7971 ( .B(n4783), .A(n4784), .Z(n4782) );
XOR U7972 ( .A(c1594), .B(b[1594]), .Z(n4783) );
XNOR U7973 ( .A(b[1594]), .B(n4784), .Z(c[1594]) );
XNOR U7974 ( .A(a[1594]), .B(c1594), .Z(n4784) );
XOR U7975 ( .A(c1595), .B(n4785), .Z(c1596) );
ANDN U7976 ( .B(n4786), .A(n4787), .Z(n4785) );
XOR U7977 ( .A(c1595), .B(b[1595]), .Z(n4786) );
XNOR U7978 ( .A(b[1595]), .B(n4787), .Z(c[1595]) );
XNOR U7979 ( .A(a[1595]), .B(c1595), .Z(n4787) );
XOR U7980 ( .A(c1596), .B(n4788), .Z(c1597) );
ANDN U7981 ( .B(n4789), .A(n4790), .Z(n4788) );
XOR U7982 ( .A(c1596), .B(b[1596]), .Z(n4789) );
XNOR U7983 ( .A(b[1596]), .B(n4790), .Z(c[1596]) );
XNOR U7984 ( .A(a[1596]), .B(c1596), .Z(n4790) );
XOR U7985 ( .A(c1597), .B(n4791), .Z(c1598) );
ANDN U7986 ( .B(n4792), .A(n4793), .Z(n4791) );
XOR U7987 ( .A(c1597), .B(b[1597]), .Z(n4792) );
XNOR U7988 ( .A(b[1597]), .B(n4793), .Z(c[1597]) );
XNOR U7989 ( .A(a[1597]), .B(c1597), .Z(n4793) );
XOR U7990 ( .A(c1598), .B(n4794), .Z(c1599) );
ANDN U7991 ( .B(n4795), .A(n4796), .Z(n4794) );
XOR U7992 ( .A(c1598), .B(b[1598]), .Z(n4795) );
XNOR U7993 ( .A(b[1598]), .B(n4796), .Z(c[1598]) );
XNOR U7994 ( .A(a[1598]), .B(c1598), .Z(n4796) );
XOR U7995 ( .A(c1599), .B(n4797), .Z(c1600) );
ANDN U7996 ( .B(n4798), .A(n4799), .Z(n4797) );
XOR U7997 ( .A(c1599), .B(b[1599]), .Z(n4798) );
XNOR U7998 ( .A(b[1599]), .B(n4799), .Z(c[1599]) );
XNOR U7999 ( .A(a[1599]), .B(c1599), .Z(n4799) );
XOR U8000 ( .A(c1600), .B(n4800), .Z(c1601) );
ANDN U8001 ( .B(n4801), .A(n4802), .Z(n4800) );
XOR U8002 ( .A(c1600), .B(b[1600]), .Z(n4801) );
XNOR U8003 ( .A(b[1600]), .B(n4802), .Z(c[1600]) );
XNOR U8004 ( .A(a[1600]), .B(c1600), .Z(n4802) );
XOR U8005 ( .A(c1601), .B(n4803), .Z(c1602) );
ANDN U8006 ( .B(n4804), .A(n4805), .Z(n4803) );
XOR U8007 ( .A(c1601), .B(b[1601]), .Z(n4804) );
XNOR U8008 ( .A(b[1601]), .B(n4805), .Z(c[1601]) );
XNOR U8009 ( .A(a[1601]), .B(c1601), .Z(n4805) );
XOR U8010 ( .A(c1602), .B(n4806), .Z(c1603) );
ANDN U8011 ( .B(n4807), .A(n4808), .Z(n4806) );
XOR U8012 ( .A(c1602), .B(b[1602]), .Z(n4807) );
XNOR U8013 ( .A(b[1602]), .B(n4808), .Z(c[1602]) );
XNOR U8014 ( .A(a[1602]), .B(c1602), .Z(n4808) );
XOR U8015 ( .A(c1603), .B(n4809), .Z(c1604) );
ANDN U8016 ( .B(n4810), .A(n4811), .Z(n4809) );
XOR U8017 ( .A(c1603), .B(b[1603]), .Z(n4810) );
XNOR U8018 ( .A(b[1603]), .B(n4811), .Z(c[1603]) );
XNOR U8019 ( .A(a[1603]), .B(c1603), .Z(n4811) );
XOR U8020 ( .A(c1604), .B(n4812), .Z(c1605) );
ANDN U8021 ( .B(n4813), .A(n4814), .Z(n4812) );
XOR U8022 ( .A(c1604), .B(b[1604]), .Z(n4813) );
XNOR U8023 ( .A(b[1604]), .B(n4814), .Z(c[1604]) );
XNOR U8024 ( .A(a[1604]), .B(c1604), .Z(n4814) );
XOR U8025 ( .A(c1605), .B(n4815), .Z(c1606) );
ANDN U8026 ( .B(n4816), .A(n4817), .Z(n4815) );
XOR U8027 ( .A(c1605), .B(b[1605]), .Z(n4816) );
XNOR U8028 ( .A(b[1605]), .B(n4817), .Z(c[1605]) );
XNOR U8029 ( .A(a[1605]), .B(c1605), .Z(n4817) );
XOR U8030 ( .A(c1606), .B(n4818), .Z(c1607) );
ANDN U8031 ( .B(n4819), .A(n4820), .Z(n4818) );
XOR U8032 ( .A(c1606), .B(b[1606]), .Z(n4819) );
XNOR U8033 ( .A(b[1606]), .B(n4820), .Z(c[1606]) );
XNOR U8034 ( .A(a[1606]), .B(c1606), .Z(n4820) );
XOR U8035 ( .A(c1607), .B(n4821), .Z(c1608) );
ANDN U8036 ( .B(n4822), .A(n4823), .Z(n4821) );
XOR U8037 ( .A(c1607), .B(b[1607]), .Z(n4822) );
XNOR U8038 ( .A(b[1607]), .B(n4823), .Z(c[1607]) );
XNOR U8039 ( .A(a[1607]), .B(c1607), .Z(n4823) );
XOR U8040 ( .A(c1608), .B(n4824), .Z(c1609) );
ANDN U8041 ( .B(n4825), .A(n4826), .Z(n4824) );
XOR U8042 ( .A(c1608), .B(b[1608]), .Z(n4825) );
XNOR U8043 ( .A(b[1608]), .B(n4826), .Z(c[1608]) );
XNOR U8044 ( .A(a[1608]), .B(c1608), .Z(n4826) );
XOR U8045 ( .A(c1609), .B(n4827), .Z(c1610) );
ANDN U8046 ( .B(n4828), .A(n4829), .Z(n4827) );
XOR U8047 ( .A(c1609), .B(b[1609]), .Z(n4828) );
XNOR U8048 ( .A(b[1609]), .B(n4829), .Z(c[1609]) );
XNOR U8049 ( .A(a[1609]), .B(c1609), .Z(n4829) );
XOR U8050 ( .A(c1610), .B(n4830), .Z(c1611) );
ANDN U8051 ( .B(n4831), .A(n4832), .Z(n4830) );
XOR U8052 ( .A(c1610), .B(b[1610]), .Z(n4831) );
XNOR U8053 ( .A(b[1610]), .B(n4832), .Z(c[1610]) );
XNOR U8054 ( .A(a[1610]), .B(c1610), .Z(n4832) );
XOR U8055 ( .A(c1611), .B(n4833), .Z(c1612) );
ANDN U8056 ( .B(n4834), .A(n4835), .Z(n4833) );
XOR U8057 ( .A(c1611), .B(b[1611]), .Z(n4834) );
XNOR U8058 ( .A(b[1611]), .B(n4835), .Z(c[1611]) );
XNOR U8059 ( .A(a[1611]), .B(c1611), .Z(n4835) );
XOR U8060 ( .A(c1612), .B(n4836), .Z(c1613) );
ANDN U8061 ( .B(n4837), .A(n4838), .Z(n4836) );
XOR U8062 ( .A(c1612), .B(b[1612]), .Z(n4837) );
XNOR U8063 ( .A(b[1612]), .B(n4838), .Z(c[1612]) );
XNOR U8064 ( .A(a[1612]), .B(c1612), .Z(n4838) );
XOR U8065 ( .A(c1613), .B(n4839), .Z(c1614) );
ANDN U8066 ( .B(n4840), .A(n4841), .Z(n4839) );
XOR U8067 ( .A(c1613), .B(b[1613]), .Z(n4840) );
XNOR U8068 ( .A(b[1613]), .B(n4841), .Z(c[1613]) );
XNOR U8069 ( .A(a[1613]), .B(c1613), .Z(n4841) );
XOR U8070 ( .A(c1614), .B(n4842), .Z(c1615) );
ANDN U8071 ( .B(n4843), .A(n4844), .Z(n4842) );
XOR U8072 ( .A(c1614), .B(b[1614]), .Z(n4843) );
XNOR U8073 ( .A(b[1614]), .B(n4844), .Z(c[1614]) );
XNOR U8074 ( .A(a[1614]), .B(c1614), .Z(n4844) );
XOR U8075 ( .A(c1615), .B(n4845), .Z(c1616) );
ANDN U8076 ( .B(n4846), .A(n4847), .Z(n4845) );
XOR U8077 ( .A(c1615), .B(b[1615]), .Z(n4846) );
XNOR U8078 ( .A(b[1615]), .B(n4847), .Z(c[1615]) );
XNOR U8079 ( .A(a[1615]), .B(c1615), .Z(n4847) );
XOR U8080 ( .A(c1616), .B(n4848), .Z(c1617) );
ANDN U8081 ( .B(n4849), .A(n4850), .Z(n4848) );
XOR U8082 ( .A(c1616), .B(b[1616]), .Z(n4849) );
XNOR U8083 ( .A(b[1616]), .B(n4850), .Z(c[1616]) );
XNOR U8084 ( .A(a[1616]), .B(c1616), .Z(n4850) );
XOR U8085 ( .A(c1617), .B(n4851), .Z(c1618) );
ANDN U8086 ( .B(n4852), .A(n4853), .Z(n4851) );
XOR U8087 ( .A(c1617), .B(b[1617]), .Z(n4852) );
XNOR U8088 ( .A(b[1617]), .B(n4853), .Z(c[1617]) );
XNOR U8089 ( .A(a[1617]), .B(c1617), .Z(n4853) );
XOR U8090 ( .A(c1618), .B(n4854), .Z(c1619) );
ANDN U8091 ( .B(n4855), .A(n4856), .Z(n4854) );
XOR U8092 ( .A(c1618), .B(b[1618]), .Z(n4855) );
XNOR U8093 ( .A(b[1618]), .B(n4856), .Z(c[1618]) );
XNOR U8094 ( .A(a[1618]), .B(c1618), .Z(n4856) );
XOR U8095 ( .A(c1619), .B(n4857), .Z(c1620) );
ANDN U8096 ( .B(n4858), .A(n4859), .Z(n4857) );
XOR U8097 ( .A(c1619), .B(b[1619]), .Z(n4858) );
XNOR U8098 ( .A(b[1619]), .B(n4859), .Z(c[1619]) );
XNOR U8099 ( .A(a[1619]), .B(c1619), .Z(n4859) );
XOR U8100 ( .A(c1620), .B(n4860), .Z(c1621) );
ANDN U8101 ( .B(n4861), .A(n4862), .Z(n4860) );
XOR U8102 ( .A(c1620), .B(b[1620]), .Z(n4861) );
XNOR U8103 ( .A(b[1620]), .B(n4862), .Z(c[1620]) );
XNOR U8104 ( .A(a[1620]), .B(c1620), .Z(n4862) );
XOR U8105 ( .A(c1621), .B(n4863), .Z(c1622) );
ANDN U8106 ( .B(n4864), .A(n4865), .Z(n4863) );
XOR U8107 ( .A(c1621), .B(b[1621]), .Z(n4864) );
XNOR U8108 ( .A(b[1621]), .B(n4865), .Z(c[1621]) );
XNOR U8109 ( .A(a[1621]), .B(c1621), .Z(n4865) );
XOR U8110 ( .A(c1622), .B(n4866), .Z(c1623) );
ANDN U8111 ( .B(n4867), .A(n4868), .Z(n4866) );
XOR U8112 ( .A(c1622), .B(b[1622]), .Z(n4867) );
XNOR U8113 ( .A(b[1622]), .B(n4868), .Z(c[1622]) );
XNOR U8114 ( .A(a[1622]), .B(c1622), .Z(n4868) );
XOR U8115 ( .A(c1623), .B(n4869), .Z(c1624) );
ANDN U8116 ( .B(n4870), .A(n4871), .Z(n4869) );
XOR U8117 ( .A(c1623), .B(b[1623]), .Z(n4870) );
XNOR U8118 ( .A(b[1623]), .B(n4871), .Z(c[1623]) );
XNOR U8119 ( .A(a[1623]), .B(c1623), .Z(n4871) );
XOR U8120 ( .A(c1624), .B(n4872), .Z(c1625) );
ANDN U8121 ( .B(n4873), .A(n4874), .Z(n4872) );
XOR U8122 ( .A(c1624), .B(b[1624]), .Z(n4873) );
XNOR U8123 ( .A(b[1624]), .B(n4874), .Z(c[1624]) );
XNOR U8124 ( .A(a[1624]), .B(c1624), .Z(n4874) );
XOR U8125 ( .A(c1625), .B(n4875), .Z(c1626) );
ANDN U8126 ( .B(n4876), .A(n4877), .Z(n4875) );
XOR U8127 ( .A(c1625), .B(b[1625]), .Z(n4876) );
XNOR U8128 ( .A(b[1625]), .B(n4877), .Z(c[1625]) );
XNOR U8129 ( .A(a[1625]), .B(c1625), .Z(n4877) );
XOR U8130 ( .A(c1626), .B(n4878), .Z(c1627) );
ANDN U8131 ( .B(n4879), .A(n4880), .Z(n4878) );
XOR U8132 ( .A(c1626), .B(b[1626]), .Z(n4879) );
XNOR U8133 ( .A(b[1626]), .B(n4880), .Z(c[1626]) );
XNOR U8134 ( .A(a[1626]), .B(c1626), .Z(n4880) );
XOR U8135 ( .A(c1627), .B(n4881), .Z(c1628) );
ANDN U8136 ( .B(n4882), .A(n4883), .Z(n4881) );
XOR U8137 ( .A(c1627), .B(b[1627]), .Z(n4882) );
XNOR U8138 ( .A(b[1627]), .B(n4883), .Z(c[1627]) );
XNOR U8139 ( .A(a[1627]), .B(c1627), .Z(n4883) );
XOR U8140 ( .A(c1628), .B(n4884), .Z(c1629) );
ANDN U8141 ( .B(n4885), .A(n4886), .Z(n4884) );
XOR U8142 ( .A(c1628), .B(b[1628]), .Z(n4885) );
XNOR U8143 ( .A(b[1628]), .B(n4886), .Z(c[1628]) );
XNOR U8144 ( .A(a[1628]), .B(c1628), .Z(n4886) );
XOR U8145 ( .A(c1629), .B(n4887), .Z(c1630) );
ANDN U8146 ( .B(n4888), .A(n4889), .Z(n4887) );
XOR U8147 ( .A(c1629), .B(b[1629]), .Z(n4888) );
XNOR U8148 ( .A(b[1629]), .B(n4889), .Z(c[1629]) );
XNOR U8149 ( .A(a[1629]), .B(c1629), .Z(n4889) );
XOR U8150 ( .A(c1630), .B(n4890), .Z(c1631) );
ANDN U8151 ( .B(n4891), .A(n4892), .Z(n4890) );
XOR U8152 ( .A(c1630), .B(b[1630]), .Z(n4891) );
XNOR U8153 ( .A(b[1630]), .B(n4892), .Z(c[1630]) );
XNOR U8154 ( .A(a[1630]), .B(c1630), .Z(n4892) );
XOR U8155 ( .A(c1631), .B(n4893), .Z(c1632) );
ANDN U8156 ( .B(n4894), .A(n4895), .Z(n4893) );
XOR U8157 ( .A(c1631), .B(b[1631]), .Z(n4894) );
XNOR U8158 ( .A(b[1631]), .B(n4895), .Z(c[1631]) );
XNOR U8159 ( .A(a[1631]), .B(c1631), .Z(n4895) );
XOR U8160 ( .A(c1632), .B(n4896), .Z(c1633) );
ANDN U8161 ( .B(n4897), .A(n4898), .Z(n4896) );
XOR U8162 ( .A(c1632), .B(b[1632]), .Z(n4897) );
XNOR U8163 ( .A(b[1632]), .B(n4898), .Z(c[1632]) );
XNOR U8164 ( .A(a[1632]), .B(c1632), .Z(n4898) );
XOR U8165 ( .A(c1633), .B(n4899), .Z(c1634) );
ANDN U8166 ( .B(n4900), .A(n4901), .Z(n4899) );
XOR U8167 ( .A(c1633), .B(b[1633]), .Z(n4900) );
XNOR U8168 ( .A(b[1633]), .B(n4901), .Z(c[1633]) );
XNOR U8169 ( .A(a[1633]), .B(c1633), .Z(n4901) );
XOR U8170 ( .A(c1634), .B(n4902), .Z(c1635) );
ANDN U8171 ( .B(n4903), .A(n4904), .Z(n4902) );
XOR U8172 ( .A(c1634), .B(b[1634]), .Z(n4903) );
XNOR U8173 ( .A(b[1634]), .B(n4904), .Z(c[1634]) );
XNOR U8174 ( .A(a[1634]), .B(c1634), .Z(n4904) );
XOR U8175 ( .A(c1635), .B(n4905), .Z(c1636) );
ANDN U8176 ( .B(n4906), .A(n4907), .Z(n4905) );
XOR U8177 ( .A(c1635), .B(b[1635]), .Z(n4906) );
XNOR U8178 ( .A(b[1635]), .B(n4907), .Z(c[1635]) );
XNOR U8179 ( .A(a[1635]), .B(c1635), .Z(n4907) );
XOR U8180 ( .A(c1636), .B(n4908), .Z(c1637) );
ANDN U8181 ( .B(n4909), .A(n4910), .Z(n4908) );
XOR U8182 ( .A(c1636), .B(b[1636]), .Z(n4909) );
XNOR U8183 ( .A(b[1636]), .B(n4910), .Z(c[1636]) );
XNOR U8184 ( .A(a[1636]), .B(c1636), .Z(n4910) );
XOR U8185 ( .A(c1637), .B(n4911), .Z(c1638) );
ANDN U8186 ( .B(n4912), .A(n4913), .Z(n4911) );
XOR U8187 ( .A(c1637), .B(b[1637]), .Z(n4912) );
XNOR U8188 ( .A(b[1637]), .B(n4913), .Z(c[1637]) );
XNOR U8189 ( .A(a[1637]), .B(c1637), .Z(n4913) );
XOR U8190 ( .A(c1638), .B(n4914), .Z(c1639) );
ANDN U8191 ( .B(n4915), .A(n4916), .Z(n4914) );
XOR U8192 ( .A(c1638), .B(b[1638]), .Z(n4915) );
XNOR U8193 ( .A(b[1638]), .B(n4916), .Z(c[1638]) );
XNOR U8194 ( .A(a[1638]), .B(c1638), .Z(n4916) );
XOR U8195 ( .A(c1639), .B(n4917), .Z(c1640) );
ANDN U8196 ( .B(n4918), .A(n4919), .Z(n4917) );
XOR U8197 ( .A(c1639), .B(b[1639]), .Z(n4918) );
XNOR U8198 ( .A(b[1639]), .B(n4919), .Z(c[1639]) );
XNOR U8199 ( .A(a[1639]), .B(c1639), .Z(n4919) );
XOR U8200 ( .A(c1640), .B(n4920), .Z(c1641) );
ANDN U8201 ( .B(n4921), .A(n4922), .Z(n4920) );
XOR U8202 ( .A(c1640), .B(b[1640]), .Z(n4921) );
XNOR U8203 ( .A(b[1640]), .B(n4922), .Z(c[1640]) );
XNOR U8204 ( .A(a[1640]), .B(c1640), .Z(n4922) );
XOR U8205 ( .A(c1641), .B(n4923), .Z(c1642) );
ANDN U8206 ( .B(n4924), .A(n4925), .Z(n4923) );
XOR U8207 ( .A(c1641), .B(b[1641]), .Z(n4924) );
XNOR U8208 ( .A(b[1641]), .B(n4925), .Z(c[1641]) );
XNOR U8209 ( .A(a[1641]), .B(c1641), .Z(n4925) );
XOR U8210 ( .A(c1642), .B(n4926), .Z(c1643) );
ANDN U8211 ( .B(n4927), .A(n4928), .Z(n4926) );
XOR U8212 ( .A(c1642), .B(b[1642]), .Z(n4927) );
XNOR U8213 ( .A(b[1642]), .B(n4928), .Z(c[1642]) );
XNOR U8214 ( .A(a[1642]), .B(c1642), .Z(n4928) );
XOR U8215 ( .A(c1643), .B(n4929), .Z(c1644) );
ANDN U8216 ( .B(n4930), .A(n4931), .Z(n4929) );
XOR U8217 ( .A(c1643), .B(b[1643]), .Z(n4930) );
XNOR U8218 ( .A(b[1643]), .B(n4931), .Z(c[1643]) );
XNOR U8219 ( .A(a[1643]), .B(c1643), .Z(n4931) );
XOR U8220 ( .A(c1644), .B(n4932), .Z(c1645) );
ANDN U8221 ( .B(n4933), .A(n4934), .Z(n4932) );
XOR U8222 ( .A(c1644), .B(b[1644]), .Z(n4933) );
XNOR U8223 ( .A(b[1644]), .B(n4934), .Z(c[1644]) );
XNOR U8224 ( .A(a[1644]), .B(c1644), .Z(n4934) );
XOR U8225 ( .A(c1645), .B(n4935), .Z(c1646) );
ANDN U8226 ( .B(n4936), .A(n4937), .Z(n4935) );
XOR U8227 ( .A(c1645), .B(b[1645]), .Z(n4936) );
XNOR U8228 ( .A(b[1645]), .B(n4937), .Z(c[1645]) );
XNOR U8229 ( .A(a[1645]), .B(c1645), .Z(n4937) );
XOR U8230 ( .A(c1646), .B(n4938), .Z(c1647) );
ANDN U8231 ( .B(n4939), .A(n4940), .Z(n4938) );
XOR U8232 ( .A(c1646), .B(b[1646]), .Z(n4939) );
XNOR U8233 ( .A(b[1646]), .B(n4940), .Z(c[1646]) );
XNOR U8234 ( .A(a[1646]), .B(c1646), .Z(n4940) );
XOR U8235 ( .A(c1647), .B(n4941), .Z(c1648) );
ANDN U8236 ( .B(n4942), .A(n4943), .Z(n4941) );
XOR U8237 ( .A(c1647), .B(b[1647]), .Z(n4942) );
XNOR U8238 ( .A(b[1647]), .B(n4943), .Z(c[1647]) );
XNOR U8239 ( .A(a[1647]), .B(c1647), .Z(n4943) );
XOR U8240 ( .A(c1648), .B(n4944), .Z(c1649) );
ANDN U8241 ( .B(n4945), .A(n4946), .Z(n4944) );
XOR U8242 ( .A(c1648), .B(b[1648]), .Z(n4945) );
XNOR U8243 ( .A(b[1648]), .B(n4946), .Z(c[1648]) );
XNOR U8244 ( .A(a[1648]), .B(c1648), .Z(n4946) );
XOR U8245 ( .A(c1649), .B(n4947), .Z(c1650) );
ANDN U8246 ( .B(n4948), .A(n4949), .Z(n4947) );
XOR U8247 ( .A(c1649), .B(b[1649]), .Z(n4948) );
XNOR U8248 ( .A(b[1649]), .B(n4949), .Z(c[1649]) );
XNOR U8249 ( .A(a[1649]), .B(c1649), .Z(n4949) );
XOR U8250 ( .A(c1650), .B(n4950), .Z(c1651) );
ANDN U8251 ( .B(n4951), .A(n4952), .Z(n4950) );
XOR U8252 ( .A(c1650), .B(b[1650]), .Z(n4951) );
XNOR U8253 ( .A(b[1650]), .B(n4952), .Z(c[1650]) );
XNOR U8254 ( .A(a[1650]), .B(c1650), .Z(n4952) );
XOR U8255 ( .A(c1651), .B(n4953), .Z(c1652) );
ANDN U8256 ( .B(n4954), .A(n4955), .Z(n4953) );
XOR U8257 ( .A(c1651), .B(b[1651]), .Z(n4954) );
XNOR U8258 ( .A(b[1651]), .B(n4955), .Z(c[1651]) );
XNOR U8259 ( .A(a[1651]), .B(c1651), .Z(n4955) );
XOR U8260 ( .A(c1652), .B(n4956), .Z(c1653) );
ANDN U8261 ( .B(n4957), .A(n4958), .Z(n4956) );
XOR U8262 ( .A(c1652), .B(b[1652]), .Z(n4957) );
XNOR U8263 ( .A(b[1652]), .B(n4958), .Z(c[1652]) );
XNOR U8264 ( .A(a[1652]), .B(c1652), .Z(n4958) );
XOR U8265 ( .A(c1653), .B(n4959), .Z(c1654) );
ANDN U8266 ( .B(n4960), .A(n4961), .Z(n4959) );
XOR U8267 ( .A(c1653), .B(b[1653]), .Z(n4960) );
XNOR U8268 ( .A(b[1653]), .B(n4961), .Z(c[1653]) );
XNOR U8269 ( .A(a[1653]), .B(c1653), .Z(n4961) );
XOR U8270 ( .A(c1654), .B(n4962), .Z(c1655) );
ANDN U8271 ( .B(n4963), .A(n4964), .Z(n4962) );
XOR U8272 ( .A(c1654), .B(b[1654]), .Z(n4963) );
XNOR U8273 ( .A(b[1654]), .B(n4964), .Z(c[1654]) );
XNOR U8274 ( .A(a[1654]), .B(c1654), .Z(n4964) );
XOR U8275 ( .A(c1655), .B(n4965), .Z(c1656) );
ANDN U8276 ( .B(n4966), .A(n4967), .Z(n4965) );
XOR U8277 ( .A(c1655), .B(b[1655]), .Z(n4966) );
XNOR U8278 ( .A(b[1655]), .B(n4967), .Z(c[1655]) );
XNOR U8279 ( .A(a[1655]), .B(c1655), .Z(n4967) );
XOR U8280 ( .A(c1656), .B(n4968), .Z(c1657) );
ANDN U8281 ( .B(n4969), .A(n4970), .Z(n4968) );
XOR U8282 ( .A(c1656), .B(b[1656]), .Z(n4969) );
XNOR U8283 ( .A(b[1656]), .B(n4970), .Z(c[1656]) );
XNOR U8284 ( .A(a[1656]), .B(c1656), .Z(n4970) );
XOR U8285 ( .A(c1657), .B(n4971), .Z(c1658) );
ANDN U8286 ( .B(n4972), .A(n4973), .Z(n4971) );
XOR U8287 ( .A(c1657), .B(b[1657]), .Z(n4972) );
XNOR U8288 ( .A(b[1657]), .B(n4973), .Z(c[1657]) );
XNOR U8289 ( .A(a[1657]), .B(c1657), .Z(n4973) );
XOR U8290 ( .A(c1658), .B(n4974), .Z(c1659) );
ANDN U8291 ( .B(n4975), .A(n4976), .Z(n4974) );
XOR U8292 ( .A(c1658), .B(b[1658]), .Z(n4975) );
XNOR U8293 ( .A(b[1658]), .B(n4976), .Z(c[1658]) );
XNOR U8294 ( .A(a[1658]), .B(c1658), .Z(n4976) );
XOR U8295 ( .A(c1659), .B(n4977), .Z(c1660) );
ANDN U8296 ( .B(n4978), .A(n4979), .Z(n4977) );
XOR U8297 ( .A(c1659), .B(b[1659]), .Z(n4978) );
XNOR U8298 ( .A(b[1659]), .B(n4979), .Z(c[1659]) );
XNOR U8299 ( .A(a[1659]), .B(c1659), .Z(n4979) );
XOR U8300 ( .A(c1660), .B(n4980), .Z(c1661) );
ANDN U8301 ( .B(n4981), .A(n4982), .Z(n4980) );
XOR U8302 ( .A(c1660), .B(b[1660]), .Z(n4981) );
XNOR U8303 ( .A(b[1660]), .B(n4982), .Z(c[1660]) );
XNOR U8304 ( .A(a[1660]), .B(c1660), .Z(n4982) );
XOR U8305 ( .A(c1661), .B(n4983), .Z(c1662) );
ANDN U8306 ( .B(n4984), .A(n4985), .Z(n4983) );
XOR U8307 ( .A(c1661), .B(b[1661]), .Z(n4984) );
XNOR U8308 ( .A(b[1661]), .B(n4985), .Z(c[1661]) );
XNOR U8309 ( .A(a[1661]), .B(c1661), .Z(n4985) );
XOR U8310 ( .A(c1662), .B(n4986), .Z(c1663) );
ANDN U8311 ( .B(n4987), .A(n4988), .Z(n4986) );
XOR U8312 ( .A(c1662), .B(b[1662]), .Z(n4987) );
XNOR U8313 ( .A(b[1662]), .B(n4988), .Z(c[1662]) );
XNOR U8314 ( .A(a[1662]), .B(c1662), .Z(n4988) );
XOR U8315 ( .A(c1663), .B(n4989), .Z(c1664) );
ANDN U8316 ( .B(n4990), .A(n4991), .Z(n4989) );
XOR U8317 ( .A(c1663), .B(b[1663]), .Z(n4990) );
XNOR U8318 ( .A(b[1663]), .B(n4991), .Z(c[1663]) );
XNOR U8319 ( .A(a[1663]), .B(c1663), .Z(n4991) );
XOR U8320 ( .A(c1664), .B(n4992), .Z(c1665) );
ANDN U8321 ( .B(n4993), .A(n4994), .Z(n4992) );
XOR U8322 ( .A(c1664), .B(b[1664]), .Z(n4993) );
XNOR U8323 ( .A(b[1664]), .B(n4994), .Z(c[1664]) );
XNOR U8324 ( .A(a[1664]), .B(c1664), .Z(n4994) );
XOR U8325 ( .A(c1665), .B(n4995), .Z(c1666) );
ANDN U8326 ( .B(n4996), .A(n4997), .Z(n4995) );
XOR U8327 ( .A(c1665), .B(b[1665]), .Z(n4996) );
XNOR U8328 ( .A(b[1665]), .B(n4997), .Z(c[1665]) );
XNOR U8329 ( .A(a[1665]), .B(c1665), .Z(n4997) );
XOR U8330 ( .A(c1666), .B(n4998), .Z(c1667) );
ANDN U8331 ( .B(n4999), .A(n5000), .Z(n4998) );
XOR U8332 ( .A(c1666), .B(b[1666]), .Z(n4999) );
XNOR U8333 ( .A(b[1666]), .B(n5000), .Z(c[1666]) );
XNOR U8334 ( .A(a[1666]), .B(c1666), .Z(n5000) );
XOR U8335 ( .A(c1667), .B(n5001), .Z(c1668) );
ANDN U8336 ( .B(n5002), .A(n5003), .Z(n5001) );
XOR U8337 ( .A(c1667), .B(b[1667]), .Z(n5002) );
XNOR U8338 ( .A(b[1667]), .B(n5003), .Z(c[1667]) );
XNOR U8339 ( .A(a[1667]), .B(c1667), .Z(n5003) );
XOR U8340 ( .A(c1668), .B(n5004), .Z(c1669) );
ANDN U8341 ( .B(n5005), .A(n5006), .Z(n5004) );
XOR U8342 ( .A(c1668), .B(b[1668]), .Z(n5005) );
XNOR U8343 ( .A(b[1668]), .B(n5006), .Z(c[1668]) );
XNOR U8344 ( .A(a[1668]), .B(c1668), .Z(n5006) );
XOR U8345 ( .A(c1669), .B(n5007), .Z(c1670) );
ANDN U8346 ( .B(n5008), .A(n5009), .Z(n5007) );
XOR U8347 ( .A(c1669), .B(b[1669]), .Z(n5008) );
XNOR U8348 ( .A(b[1669]), .B(n5009), .Z(c[1669]) );
XNOR U8349 ( .A(a[1669]), .B(c1669), .Z(n5009) );
XOR U8350 ( .A(c1670), .B(n5010), .Z(c1671) );
ANDN U8351 ( .B(n5011), .A(n5012), .Z(n5010) );
XOR U8352 ( .A(c1670), .B(b[1670]), .Z(n5011) );
XNOR U8353 ( .A(b[1670]), .B(n5012), .Z(c[1670]) );
XNOR U8354 ( .A(a[1670]), .B(c1670), .Z(n5012) );
XOR U8355 ( .A(c1671), .B(n5013), .Z(c1672) );
ANDN U8356 ( .B(n5014), .A(n5015), .Z(n5013) );
XOR U8357 ( .A(c1671), .B(b[1671]), .Z(n5014) );
XNOR U8358 ( .A(b[1671]), .B(n5015), .Z(c[1671]) );
XNOR U8359 ( .A(a[1671]), .B(c1671), .Z(n5015) );
XOR U8360 ( .A(c1672), .B(n5016), .Z(c1673) );
ANDN U8361 ( .B(n5017), .A(n5018), .Z(n5016) );
XOR U8362 ( .A(c1672), .B(b[1672]), .Z(n5017) );
XNOR U8363 ( .A(b[1672]), .B(n5018), .Z(c[1672]) );
XNOR U8364 ( .A(a[1672]), .B(c1672), .Z(n5018) );
XOR U8365 ( .A(c1673), .B(n5019), .Z(c1674) );
ANDN U8366 ( .B(n5020), .A(n5021), .Z(n5019) );
XOR U8367 ( .A(c1673), .B(b[1673]), .Z(n5020) );
XNOR U8368 ( .A(b[1673]), .B(n5021), .Z(c[1673]) );
XNOR U8369 ( .A(a[1673]), .B(c1673), .Z(n5021) );
XOR U8370 ( .A(c1674), .B(n5022), .Z(c1675) );
ANDN U8371 ( .B(n5023), .A(n5024), .Z(n5022) );
XOR U8372 ( .A(c1674), .B(b[1674]), .Z(n5023) );
XNOR U8373 ( .A(b[1674]), .B(n5024), .Z(c[1674]) );
XNOR U8374 ( .A(a[1674]), .B(c1674), .Z(n5024) );
XOR U8375 ( .A(c1675), .B(n5025), .Z(c1676) );
ANDN U8376 ( .B(n5026), .A(n5027), .Z(n5025) );
XOR U8377 ( .A(c1675), .B(b[1675]), .Z(n5026) );
XNOR U8378 ( .A(b[1675]), .B(n5027), .Z(c[1675]) );
XNOR U8379 ( .A(a[1675]), .B(c1675), .Z(n5027) );
XOR U8380 ( .A(c1676), .B(n5028), .Z(c1677) );
ANDN U8381 ( .B(n5029), .A(n5030), .Z(n5028) );
XOR U8382 ( .A(c1676), .B(b[1676]), .Z(n5029) );
XNOR U8383 ( .A(b[1676]), .B(n5030), .Z(c[1676]) );
XNOR U8384 ( .A(a[1676]), .B(c1676), .Z(n5030) );
XOR U8385 ( .A(c1677), .B(n5031), .Z(c1678) );
ANDN U8386 ( .B(n5032), .A(n5033), .Z(n5031) );
XOR U8387 ( .A(c1677), .B(b[1677]), .Z(n5032) );
XNOR U8388 ( .A(b[1677]), .B(n5033), .Z(c[1677]) );
XNOR U8389 ( .A(a[1677]), .B(c1677), .Z(n5033) );
XOR U8390 ( .A(c1678), .B(n5034), .Z(c1679) );
ANDN U8391 ( .B(n5035), .A(n5036), .Z(n5034) );
XOR U8392 ( .A(c1678), .B(b[1678]), .Z(n5035) );
XNOR U8393 ( .A(b[1678]), .B(n5036), .Z(c[1678]) );
XNOR U8394 ( .A(a[1678]), .B(c1678), .Z(n5036) );
XOR U8395 ( .A(c1679), .B(n5037), .Z(c1680) );
ANDN U8396 ( .B(n5038), .A(n5039), .Z(n5037) );
XOR U8397 ( .A(c1679), .B(b[1679]), .Z(n5038) );
XNOR U8398 ( .A(b[1679]), .B(n5039), .Z(c[1679]) );
XNOR U8399 ( .A(a[1679]), .B(c1679), .Z(n5039) );
XOR U8400 ( .A(c1680), .B(n5040), .Z(c1681) );
ANDN U8401 ( .B(n5041), .A(n5042), .Z(n5040) );
XOR U8402 ( .A(c1680), .B(b[1680]), .Z(n5041) );
XNOR U8403 ( .A(b[1680]), .B(n5042), .Z(c[1680]) );
XNOR U8404 ( .A(a[1680]), .B(c1680), .Z(n5042) );
XOR U8405 ( .A(c1681), .B(n5043), .Z(c1682) );
ANDN U8406 ( .B(n5044), .A(n5045), .Z(n5043) );
XOR U8407 ( .A(c1681), .B(b[1681]), .Z(n5044) );
XNOR U8408 ( .A(b[1681]), .B(n5045), .Z(c[1681]) );
XNOR U8409 ( .A(a[1681]), .B(c1681), .Z(n5045) );
XOR U8410 ( .A(c1682), .B(n5046), .Z(c1683) );
ANDN U8411 ( .B(n5047), .A(n5048), .Z(n5046) );
XOR U8412 ( .A(c1682), .B(b[1682]), .Z(n5047) );
XNOR U8413 ( .A(b[1682]), .B(n5048), .Z(c[1682]) );
XNOR U8414 ( .A(a[1682]), .B(c1682), .Z(n5048) );
XOR U8415 ( .A(c1683), .B(n5049), .Z(c1684) );
ANDN U8416 ( .B(n5050), .A(n5051), .Z(n5049) );
XOR U8417 ( .A(c1683), .B(b[1683]), .Z(n5050) );
XNOR U8418 ( .A(b[1683]), .B(n5051), .Z(c[1683]) );
XNOR U8419 ( .A(a[1683]), .B(c1683), .Z(n5051) );
XOR U8420 ( .A(c1684), .B(n5052), .Z(c1685) );
ANDN U8421 ( .B(n5053), .A(n5054), .Z(n5052) );
XOR U8422 ( .A(c1684), .B(b[1684]), .Z(n5053) );
XNOR U8423 ( .A(b[1684]), .B(n5054), .Z(c[1684]) );
XNOR U8424 ( .A(a[1684]), .B(c1684), .Z(n5054) );
XOR U8425 ( .A(c1685), .B(n5055), .Z(c1686) );
ANDN U8426 ( .B(n5056), .A(n5057), .Z(n5055) );
XOR U8427 ( .A(c1685), .B(b[1685]), .Z(n5056) );
XNOR U8428 ( .A(b[1685]), .B(n5057), .Z(c[1685]) );
XNOR U8429 ( .A(a[1685]), .B(c1685), .Z(n5057) );
XOR U8430 ( .A(c1686), .B(n5058), .Z(c1687) );
ANDN U8431 ( .B(n5059), .A(n5060), .Z(n5058) );
XOR U8432 ( .A(c1686), .B(b[1686]), .Z(n5059) );
XNOR U8433 ( .A(b[1686]), .B(n5060), .Z(c[1686]) );
XNOR U8434 ( .A(a[1686]), .B(c1686), .Z(n5060) );
XOR U8435 ( .A(c1687), .B(n5061), .Z(c1688) );
ANDN U8436 ( .B(n5062), .A(n5063), .Z(n5061) );
XOR U8437 ( .A(c1687), .B(b[1687]), .Z(n5062) );
XNOR U8438 ( .A(b[1687]), .B(n5063), .Z(c[1687]) );
XNOR U8439 ( .A(a[1687]), .B(c1687), .Z(n5063) );
XOR U8440 ( .A(c1688), .B(n5064), .Z(c1689) );
ANDN U8441 ( .B(n5065), .A(n5066), .Z(n5064) );
XOR U8442 ( .A(c1688), .B(b[1688]), .Z(n5065) );
XNOR U8443 ( .A(b[1688]), .B(n5066), .Z(c[1688]) );
XNOR U8444 ( .A(a[1688]), .B(c1688), .Z(n5066) );
XOR U8445 ( .A(c1689), .B(n5067), .Z(c1690) );
ANDN U8446 ( .B(n5068), .A(n5069), .Z(n5067) );
XOR U8447 ( .A(c1689), .B(b[1689]), .Z(n5068) );
XNOR U8448 ( .A(b[1689]), .B(n5069), .Z(c[1689]) );
XNOR U8449 ( .A(a[1689]), .B(c1689), .Z(n5069) );
XOR U8450 ( .A(c1690), .B(n5070), .Z(c1691) );
ANDN U8451 ( .B(n5071), .A(n5072), .Z(n5070) );
XOR U8452 ( .A(c1690), .B(b[1690]), .Z(n5071) );
XNOR U8453 ( .A(b[1690]), .B(n5072), .Z(c[1690]) );
XNOR U8454 ( .A(a[1690]), .B(c1690), .Z(n5072) );
XOR U8455 ( .A(c1691), .B(n5073), .Z(c1692) );
ANDN U8456 ( .B(n5074), .A(n5075), .Z(n5073) );
XOR U8457 ( .A(c1691), .B(b[1691]), .Z(n5074) );
XNOR U8458 ( .A(b[1691]), .B(n5075), .Z(c[1691]) );
XNOR U8459 ( .A(a[1691]), .B(c1691), .Z(n5075) );
XOR U8460 ( .A(c1692), .B(n5076), .Z(c1693) );
ANDN U8461 ( .B(n5077), .A(n5078), .Z(n5076) );
XOR U8462 ( .A(c1692), .B(b[1692]), .Z(n5077) );
XNOR U8463 ( .A(b[1692]), .B(n5078), .Z(c[1692]) );
XNOR U8464 ( .A(a[1692]), .B(c1692), .Z(n5078) );
XOR U8465 ( .A(c1693), .B(n5079), .Z(c1694) );
ANDN U8466 ( .B(n5080), .A(n5081), .Z(n5079) );
XOR U8467 ( .A(c1693), .B(b[1693]), .Z(n5080) );
XNOR U8468 ( .A(b[1693]), .B(n5081), .Z(c[1693]) );
XNOR U8469 ( .A(a[1693]), .B(c1693), .Z(n5081) );
XOR U8470 ( .A(c1694), .B(n5082), .Z(c1695) );
ANDN U8471 ( .B(n5083), .A(n5084), .Z(n5082) );
XOR U8472 ( .A(c1694), .B(b[1694]), .Z(n5083) );
XNOR U8473 ( .A(b[1694]), .B(n5084), .Z(c[1694]) );
XNOR U8474 ( .A(a[1694]), .B(c1694), .Z(n5084) );
XOR U8475 ( .A(c1695), .B(n5085), .Z(c1696) );
ANDN U8476 ( .B(n5086), .A(n5087), .Z(n5085) );
XOR U8477 ( .A(c1695), .B(b[1695]), .Z(n5086) );
XNOR U8478 ( .A(b[1695]), .B(n5087), .Z(c[1695]) );
XNOR U8479 ( .A(a[1695]), .B(c1695), .Z(n5087) );
XOR U8480 ( .A(c1696), .B(n5088), .Z(c1697) );
ANDN U8481 ( .B(n5089), .A(n5090), .Z(n5088) );
XOR U8482 ( .A(c1696), .B(b[1696]), .Z(n5089) );
XNOR U8483 ( .A(b[1696]), .B(n5090), .Z(c[1696]) );
XNOR U8484 ( .A(a[1696]), .B(c1696), .Z(n5090) );
XOR U8485 ( .A(c1697), .B(n5091), .Z(c1698) );
ANDN U8486 ( .B(n5092), .A(n5093), .Z(n5091) );
XOR U8487 ( .A(c1697), .B(b[1697]), .Z(n5092) );
XNOR U8488 ( .A(b[1697]), .B(n5093), .Z(c[1697]) );
XNOR U8489 ( .A(a[1697]), .B(c1697), .Z(n5093) );
XOR U8490 ( .A(c1698), .B(n5094), .Z(c1699) );
ANDN U8491 ( .B(n5095), .A(n5096), .Z(n5094) );
XOR U8492 ( .A(c1698), .B(b[1698]), .Z(n5095) );
XNOR U8493 ( .A(b[1698]), .B(n5096), .Z(c[1698]) );
XNOR U8494 ( .A(a[1698]), .B(c1698), .Z(n5096) );
XOR U8495 ( .A(c1699), .B(n5097), .Z(c1700) );
ANDN U8496 ( .B(n5098), .A(n5099), .Z(n5097) );
XOR U8497 ( .A(c1699), .B(b[1699]), .Z(n5098) );
XNOR U8498 ( .A(b[1699]), .B(n5099), .Z(c[1699]) );
XNOR U8499 ( .A(a[1699]), .B(c1699), .Z(n5099) );
XOR U8500 ( .A(c1700), .B(n5100), .Z(c1701) );
ANDN U8501 ( .B(n5101), .A(n5102), .Z(n5100) );
XOR U8502 ( .A(c1700), .B(b[1700]), .Z(n5101) );
XNOR U8503 ( .A(b[1700]), .B(n5102), .Z(c[1700]) );
XNOR U8504 ( .A(a[1700]), .B(c1700), .Z(n5102) );
XOR U8505 ( .A(c1701), .B(n5103), .Z(c1702) );
ANDN U8506 ( .B(n5104), .A(n5105), .Z(n5103) );
XOR U8507 ( .A(c1701), .B(b[1701]), .Z(n5104) );
XNOR U8508 ( .A(b[1701]), .B(n5105), .Z(c[1701]) );
XNOR U8509 ( .A(a[1701]), .B(c1701), .Z(n5105) );
XOR U8510 ( .A(c1702), .B(n5106), .Z(c1703) );
ANDN U8511 ( .B(n5107), .A(n5108), .Z(n5106) );
XOR U8512 ( .A(c1702), .B(b[1702]), .Z(n5107) );
XNOR U8513 ( .A(b[1702]), .B(n5108), .Z(c[1702]) );
XNOR U8514 ( .A(a[1702]), .B(c1702), .Z(n5108) );
XOR U8515 ( .A(c1703), .B(n5109), .Z(c1704) );
ANDN U8516 ( .B(n5110), .A(n5111), .Z(n5109) );
XOR U8517 ( .A(c1703), .B(b[1703]), .Z(n5110) );
XNOR U8518 ( .A(b[1703]), .B(n5111), .Z(c[1703]) );
XNOR U8519 ( .A(a[1703]), .B(c1703), .Z(n5111) );
XOR U8520 ( .A(c1704), .B(n5112), .Z(c1705) );
ANDN U8521 ( .B(n5113), .A(n5114), .Z(n5112) );
XOR U8522 ( .A(c1704), .B(b[1704]), .Z(n5113) );
XNOR U8523 ( .A(b[1704]), .B(n5114), .Z(c[1704]) );
XNOR U8524 ( .A(a[1704]), .B(c1704), .Z(n5114) );
XOR U8525 ( .A(c1705), .B(n5115), .Z(c1706) );
ANDN U8526 ( .B(n5116), .A(n5117), .Z(n5115) );
XOR U8527 ( .A(c1705), .B(b[1705]), .Z(n5116) );
XNOR U8528 ( .A(b[1705]), .B(n5117), .Z(c[1705]) );
XNOR U8529 ( .A(a[1705]), .B(c1705), .Z(n5117) );
XOR U8530 ( .A(c1706), .B(n5118), .Z(c1707) );
ANDN U8531 ( .B(n5119), .A(n5120), .Z(n5118) );
XOR U8532 ( .A(c1706), .B(b[1706]), .Z(n5119) );
XNOR U8533 ( .A(b[1706]), .B(n5120), .Z(c[1706]) );
XNOR U8534 ( .A(a[1706]), .B(c1706), .Z(n5120) );
XOR U8535 ( .A(c1707), .B(n5121), .Z(c1708) );
ANDN U8536 ( .B(n5122), .A(n5123), .Z(n5121) );
XOR U8537 ( .A(c1707), .B(b[1707]), .Z(n5122) );
XNOR U8538 ( .A(b[1707]), .B(n5123), .Z(c[1707]) );
XNOR U8539 ( .A(a[1707]), .B(c1707), .Z(n5123) );
XOR U8540 ( .A(c1708), .B(n5124), .Z(c1709) );
ANDN U8541 ( .B(n5125), .A(n5126), .Z(n5124) );
XOR U8542 ( .A(c1708), .B(b[1708]), .Z(n5125) );
XNOR U8543 ( .A(b[1708]), .B(n5126), .Z(c[1708]) );
XNOR U8544 ( .A(a[1708]), .B(c1708), .Z(n5126) );
XOR U8545 ( .A(c1709), .B(n5127), .Z(c1710) );
ANDN U8546 ( .B(n5128), .A(n5129), .Z(n5127) );
XOR U8547 ( .A(c1709), .B(b[1709]), .Z(n5128) );
XNOR U8548 ( .A(b[1709]), .B(n5129), .Z(c[1709]) );
XNOR U8549 ( .A(a[1709]), .B(c1709), .Z(n5129) );
XOR U8550 ( .A(c1710), .B(n5130), .Z(c1711) );
ANDN U8551 ( .B(n5131), .A(n5132), .Z(n5130) );
XOR U8552 ( .A(c1710), .B(b[1710]), .Z(n5131) );
XNOR U8553 ( .A(b[1710]), .B(n5132), .Z(c[1710]) );
XNOR U8554 ( .A(a[1710]), .B(c1710), .Z(n5132) );
XOR U8555 ( .A(c1711), .B(n5133), .Z(c1712) );
ANDN U8556 ( .B(n5134), .A(n5135), .Z(n5133) );
XOR U8557 ( .A(c1711), .B(b[1711]), .Z(n5134) );
XNOR U8558 ( .A(b[1711]), .B(n5135), .Z(c[1711]) );
XNOR U8559 ( .A(a[1711]), .B(c1711), .Z(n5135) );
XOR U8560 ( .A(c1712), .B(n5136), .Z(c1713) );
ANDN U8561 ( .B(n5137), .A(n5138), .Z(n5136) );
XOR U8562 ( .A(c1712), .B(b[1712]), .Z(n5137) );
XNOR U8563 ( .A(b[1712]), .B(n5138), .Z(c[1712]) );
XNOR U8564 ( .A(a[1712]), .B(c1712), .Z(n5138) );
XOR U8565 ( .A(c1713), .B(n5139), .Z(c1714) );
ANDN U8566 ( .B(n5140), .A(n5141), .Z(n5139) );
XOR U8567 ( .A(c1713), .B(b[1713]), .Z(n5140) );
XNOR U8568 ( .A(b[1713]), .B(n5141), .Z(c[1713]) );
XNOR U8569 ( .A(a[1713]), .B(c1713), .Z(n5141) );
XOR U8570 ( .A(c1714), .B(n5142), .Z(c1715) );
ANDN U8571 ( .B(n5143), .A(n5144), .Z(n5142) );
XOR U8572 ( .A(c1714), .B(b[1714]), .Z(n5143) );
XNOR U8573 ( .A(b[1714]), .B(n5144), .Z(c[1714]) );
XNOR U8574 ( .A(a[1714]), .B(c1714), .Z(n5144) );
XOR U8575 ( .A(c1715), .B(n5145), .Z(c1716) );
ANDN U8576 ( .B(n5146), .A(n5147), .Z(n5145) );
XOR U8577 ( .A(c1715), .B(b[1715]), .Z(n5146) );
XNOR U8578 ( .A(b[1715]), .B(n5147), .Z(c[1715]) );
XNOR U8579 ( .A(a[1715]), .B(c1715), .Z(n5147) );
XOR U8580 ( .A(c1716), .B(n5148), .Z(c1717) );
ANDN U8581 ( .B(n5149), .A(n5150), .Z(n5148) );
XOR U8582 ( .A(c1716), .B(b[1716]), .Z(n5149) );
XNOR U8583 ( .A(b[1716]), .B(n5150), .Z(c[1716]) );
XNOR U8584 ( .A(a[1716]), .B(c1716), .Z(n5150) );
XOR U8585 ( .A(c1717), .B(n5151), .Z(c1718) );
ANDN U8586 ( .B(n5152), .A(n5153), .Z(n5151) );
XOR U8587 ( .A(c1717), .B(b[1717]), .Z(n5152) );
XNOR U8588 ( .A(b[1717]), .B(n5153), .Z(c[1717]) );
XNOR U8589 ( .A(a[1717]), .B(c1717), .Z(n5153) );
XOR U8590 ( .A(c1718), .B(n5154), .Z(c1719) );
ANDN U8591 ( .B(n5155), .A(n5156), .Z(n5154) );
XOR U8592 ( .A(c1718), .B(b[1718]), .Z(n5155) );
XNOR U8593 ( .A(b[1718]), .B(n5156), .Z(c[1718]) );
XNOR U8594 ( .A(a[1718]), .B(c1718), .Z(n5156) );
XOR U8595 ( .A(c1719), .B(n5157), .Z(c1720) );
ANDN U8596 ( .B(n5158), .A(n5159), .Z(n5157) );
XOR U8597 ( .A(c1719), .B(b[1719]), .Z(n5158) );
XNOR U8598 ( .A(b[1719]), .B(n5159), .Z(c[1719]) );
XNOR U8599 ( .A(a[1719]), .B(c1719), .Z(n5159) );
XOR U8600 ( .A(c1720), .B(n5160), .Z(c1721) );
ANDN U8601 ( .B(n5161), .A(n5162), .Z(n5160) );
XOR U8602 ( .A(c1720), .B(b[1720]), .Z(n5161) );
XNOR U8603 ( .A(b[1720]), .B(n5162), .Z(c[1720]) );
XNOR U8604 ( .A(a[1720]), .B(c1720), .Z(n5162) );
XOR U8605 ( .A(c1721), .B(n5163), .Z(c1722) );
ANDN U8606 ( .B(n5164), .A(n5165), .Z(n5163) );
XOR U8607 ( .A(c1721), .B(b[1721]), .Z(n5164) );
XNOR U8608 ( .A(b[1721]), .B(n5165), .Z(c[1721]) );
XNOR U8609 ( .A(a[1721]), .B(c1721), .Z(n5165) );
XOR U8610 ( .A(c1722), .B(n5166), .Z(c1723) );
ANDN U8611 ( .B(n5167), .A(n5168), .Z(n5166) );
XOR U8612 ( .A(c1722), .B(b[1722]), .Z(n5167) );
XNOR U8613 ( .A(b[1722]), .B(n5168), .Z(c[1722]) );
XNOR U8614 ( .A(a[1722]), .B(c1722), .Z(n5168) );
XOR U8615 ( .A(c1723), .B(n5169), .Z(c1724) );
ANDN U8616 ( .B(n5170), .A(n5171), .Z(n5169) );
XOR U8617 ( .A(c1723), .B(b[1723]), .Z(n5170) );
XNOR U8618 ( .A(b[1723]), .B(n5171), .Z(c[1723]) );
XNOR U8619 ( .A(a[1723]), .B(c1723), .Z(n5171) );
XOR U8620 ( .A(c1724), .B(n5172), .Z(c1725) );
ANDN U8621 ( .B(n5173), .A(n5174), .Z(n5172) );
XOR U8622 ( .A(c1724), .B(b[1724]), .Z(n5173) );
XNOR U8623 ( .A(b[1724]), .B(n5174), .Z(c[1724]) );
XNOR U8624 ( .A(a[1724]), .B(c1724), .Z(n5174) );
XOR U8625 ( .A(c1725), .B(n5175), .Z(c1726) );
ANDN U8626 ( .B(n5176), .A(n5177), .Z(n5175) );
XOR U8627 ( .A(c1725), .B(b[1725]), .Z(n5176) );
XNOR U8628 ( .A(b[1725]), .B(n5177), .Z(c[1725]) );
XNOR U8629 ( .A(a[1725]), .B(c1725), .Z(n5177) );
XOR U8630 ( .A(c1726), .B(n5178), .Z(c1727) );
ANDN U8631 ( .B(n5179), .A(n5180), .Z(n5178) );
XOR U8632 ( .A(c1726), .B(b[1726]), .Z(n5179) );
XNOR U8633 ( .A(b[1726]), .B(n5180), .Z(c[1726]) );
XNOR U8634 ( .A(a[1726]), .B(c1726), .Z(n5180) );
XOR U8635 ( .A(c1727), .B(n5181), .Z(c1728) );
ANDN U8636 ( .B(n5182), .A(n5183), .Z(n5181) );
XOR U8637 ( .A(c1727), .B(b[1727]), .Z(n5182) );
XNOR U8638 ( .A(b[1727]), .B(n5183), .Z(c[1727]) );
XNOR U8639 ( .A(a[1727]), .B(c1727), .Z(n5183) );
XOR U8640 ( .A(c1728), .B(n5184), .Z(c1729) );
ANDN U8641 ( .B(n5185), .A(n5186), .Z(n5184) );
XOR U8642 ( .A(c1728), .B(b[1728]), .Z(n5185) );
XNOR U8643 ( .A(b[1728]), .B(n5186), .Z(c[1728]) );
XNOR U8644 ( .A(a[1728]), .B(c1728), .Z(n5186) );
XOR U8645 ( .A(c1729), .B(n5187), .Z(c1730) );
ANDN U8646 ( .B(n5188), .A(n5189), .Z(n5187) );
XOR U8647 ( .A(c1729), .B(b[1729]), .Z(n5188) );
XNOR U8648 ( .A(b[1729]), .B(n5189), .Z(c[1729]) );
XNOR U8649 ( .A(a[1729]), .B(c1729), .Z(n5189) );
XOR U8650 ( .A(c1730), .B(n5190), .Z(c1731) );
ANDN U8651 ( .B(n5191), .A(n5192), .Z(n5190) );
XOR U8652 ( .A(c1730), .B(b[1730]), .Z(n5191) );
XNOR U8653 ( .A(b[1730]), .B(n5192), .Z(c[1730]) );
XNOR U8654 ( .A(a[1730]), .B(c1730), .Z(n5192) );
XOR U8655 ( .A(c1731), .B(n5193), .Z(c1732) );
ANDN U8656 ( .B(n5194), .A(n5195), .Z(n5193) );
XOR U8657 ( .A(c1731), .B(b[1731]), .Z(n5194) );
XNOR U8658 ( .A(b[1731]), .B(n5195), .Z(c[1731]) );
XNOR U8659 ( .A(a[1731]), .B(c1731), .Z(n5195) );
XOR U8660 ( .A(c1732), .B(n5196), .Z(c1733) );
ANDN U8661 ( .B(n5197), .A(n5198), .Z(n5196) );
XOR U8662 ( .A(c1732), .B(b[1732]), .Z(n5197) );
XNOR U8663 ( .A(b[1732]), .B(n5198), .Z(c[1732]) );
XNOR U8664 ( .A(a[1732]), .B(c1732), .Z(n5198) );
XOR U8665 ( .A(c1733), .B(n5199), .Z(c1734) );
ANDN U8666 ( .B(n5200), .A(n5201), .Z(n5199) );
XOR U8667 ( .A(c1733), .B(b[1733]), .Z(n5200) );
XNOR U8668 ( .A(b[1733]), .B(n5201), .Z(c[1733]) );
XNOR U8669 ( .A(a[1733]), .B(c1733), .Z(n5201) );
XOR U8670 ( .A(c1734), .B(n5202), .Z(c1735) );
ANDN U8671 ( .B(n5203), .A(n5204), .Z(n5202) );
XOR U8672 ( .A(c1734), .B(b[1734]), .Z(n5203) );
XNOR U8673 ( .A(b[1734]), .B(n5204), .Z(c[1734]) );
XNOR U8674 ( .A(a[1734]), .B(c1734), .Z(n5204) );
XOR U8675 ( .A(c1735), .B(n5205), .Z(c1736) );
ANDN U8676 ( .B(n5206), .A(n5207), .Z(n5205) );
XOR U8677 ( .A(c1735), .B(b[1735]), .Z(n5206) );
XNOR U8678 ( .A(b[1735]), .B(n5207), .Z(c[1735]) );
XNOR U8679 ( .A(a[1735]), .B(c1735), .Z(n5207) );
XOR U8680 ( .A(c1736), .B(n5208), .Z(c1737) );
ANDN U8681 ( .B(n5209), .A(n5210), .Z(n5208) );
XOR U8682 ( .A(c1736), .B(b[1736]), .Z(n5209) );
XNOR U8683 ( .A(b[1736]), .B(n5210), .Z(c[1736]) );
XNOR U8684 ( .A(a[1736]), .B(c1736), .Z(n5210) );
XOR U8685 ( .A(c1737), .B(n5211), .Z(c1738) );
ANDN U8686 ( .B(n5212), .A(n5213), .Z(n5211) );
XOR U8687 ( .A(c1737), .B(b[1737]), .Z(n5212) );
XNOR U8688 ( .A(b[1737]), .B(n5213), .Z(c[1737]) );
XNOR U8689 ( .A(a[1737]), .B(c1737), .Z(n5213) );
XOR U8690 ( .A(c1738), .B(n5214), .Z(c1739) );
ANDN U8691 ( .B(n5215), .A(n5216), .Z(n5214) );
XOR U8692 ( .A(c1738), .B(b[1738]), .Z(n5215) );
XNOR U8693 ( .A(b[1738]), .B(n5216), .Z(c[1738]) );
XNOR U8694 ( .A(a[1738]), .B(c1738), .Z(n5216) );
XOR U8695 ( .A(c1739), .B(n5217), .Z(c1740) );
ANDN U8696 ( .B(n5218), .A(n5219), .Z(n5217) );
XOR U8697 ( .A(c1739), .B(b[1739]), .Z(n5218) );
XNOR U8698 ( .A(b[1739]), .B(n5219), .Z(c[1739]) );
XNOR U8699 ( .A(a[1739]), .B(c1739), .Z(n5219) );
XOR U8700 ( .A(c1740), .B(n5220), .Z(c1741) );
ANDN U8701 ( .B(n5221), .A(n5222), .Z(n5220) );
XOR U8702 ( .A(c1740), .B(b[1740]), .Z(n5221) );
XNOR U8703 ( .A(b[1740]), .B(n5222), .Z(c[1740]) );
XNOR U8704 ( .A(a[1740]), .B(c1740), .Z(n5222) );
XOR U8705 ( .A(c1741), .B(n5223), .Z(c1742) );
ANDN U8706 ( .B(n5224), .A(n5225), .Z(n5223) );
XOR U8707 ( .A(c1741), .B(b[1741]), .Z(n5224) );
XNOR U8708 ( .A(b[1741]), .B(n5225), .Z(c[1741]) );
XNOR U8709 ( .A(a[1741]), .B(c1741), .Z(n5225) );
XOR U8710 ( .A(c1742), .B(n5226), .Z(c1743) );
ANDN U8711 ( .B(n5227), .A(n5228), .Z(n5226) );
XOR U8712 ( .A(c1742), .B(b[1742]), .Z(n5227) );
XNOR U8713 ( .A(b[1742]), .B(n5228), .Z(c[1742]) );
XNOR U8714 ( .A(a[1742]), .B(c1742), .Z(n5228) );
XOR U8715 ( .A(c1743), .B(n5229), .Z(c1744) );
ANDN U8716 ( .B(n5230), .A(n5231), .Z(n5229) );
XOR U8717 ( .A(c1743), .B(b[1743]), .Z(n5230) );
XNOR U8718 ( .A(b[1743]), .B(n5231), .Z(c[1743]) );
XNOR U8719 ( .A(a[1743]), .B(c1743), .Z(n5231) );
XOR U8720 ( .A(c1744), .B(n5232), .Z(c1745) );
ANDN U8721 ( .B(n5233), .A(n5234), .Z(n5232) );
XOR U8722 ( .A(c1744), .B(b[1744]), .Z(n5233) );
XNOR U8723 ( .A(b[1744]), .B(n5234), .Z(c[1744]) );
XNOR U8724 ( .A(a[1744]), .B(c1744), .Z(n5234) );
XOR U8725 ( .A(c1745), .B(n5235), .Z(c1746) );
ANDN U8726 ( .B(n5236), .A(n5237), .Z(n5235) );
XOR U8727 ( .A(c1745), .B(b[1745]), .Z(n5236) );
XNOR U8728 ( .A(b[1745]), .B(n5237), .Z(c[1745]) );
XNOR U8729 ( .A(a[1745]), .B(c1745), .Z(n5237) );
XOR U8730 ( .A(c1746), .B(n5238), .Z(c1747) );
ANDN U8731 ( .B(n5239), .A(n5240), .Z(n5238) );
XOR U8732 ( .A(c1746), .B(b[1746]), .Z(n5239) );
XNOR U8733 ( .A(b[1746]), .B(n5240), .Z(c[1746]) );
XNOR U8734 ( .A(a[1746]), .B(c1746), .Z(n5240) );
XOR U8735 ( .A(c1747), .B(n5241), .Z(c1748) );
ANDN U8736 ( .B(n5242), .A(n5243), .Z(n5241) );
XOR U8737 ( .A(c1747), .B(b[1747]), .Z(n5242) );
XNOR U8738 ( .A(b[1747]), .B(n5243), .Z(c[1747]) );
XNOR U8739 ( .A(a[1747]), .B(c1747), .Z(n5243) );
XOR U8740 ( .A(c1748), .B(n5244), .Z(c1749) );
ANDN U8741 ( .B(n5245), .A(n5246), .Z(n5244) );
XOR U8742 ( .A(c1748), .B(b[1748]), .Z(n5245) );
XNOR U8743 ( .A(b[1748]), .B(n5246), .Z(c[1748]) );
XNOR U8744 ( .A(a[1748]), .B(c1748), .Z(n5246) );
XOR U8745 ( .A(c1749), .B(n5247), .Z(c1750) );
ANDN U8746 ( .B(n5248), .A(n5249), .Z(n5247) );
XOR U8747 ( .A(c1749), .B(b[1749]), .Z(n5248) );
XNOR U8748 ( .A(b[1749]), .B(n5249), .Z(c[1749]) );
XNOR U8749 ( .A(a[1749]), .B(c1749), .Z(n5249) );
XOR U8750 ( .A(c1750), .B(n5250), .Z(c1751) );
ANDN U8751 ( .B(n5251), .A(n5252), .Z(n5250) );
XOR U8752 ( .A(c1750), .B(b[1750]), .Z(n5251) );
XNOR U8753 ( .A(b[1750]), .B(n5252), .Z(c[1750]) );
XNOR U8754 ( .A(a[1750]), .B(c1750), .Z(n5252) );
XOR U8755 ( .A(c1751), .B(n5253), .Z(c1752) );
ANDN U8756 ( .B(n5254), .A(n5255), .Z(n5253) );
XOR U8757 ( .A(c1751), .B(b[1751]), .Z(n5254) );
XNOR U8758 ( .A(b[1751]), .B(n5255), .Z(c[1751]) );
XNOR U8759 ( .A(a[1751]), .B(c1751), .Z(n5255) );
XOR U8760 ( .A(c1752), .B(n5256), .Z(c1753) );
ANDN U8761 ( .B(n5257), .A(n5258), .Z(n5256) );
XOR U8762 ( .A(c1752), .B(b[1752]), .Z(n5257) );
XNOR U8763 ( .A(b[1752]), .B(n5258), .Z(c[1752]) );
XNOR U8764 ( .A(a[1752]), .B(c1752), .Z(n5258) );
XOR U8765 ( .A(c1753), .B(n5259), .Z(c1754) );
ANDN U8766 ( .B(n5260), .A(n5261), .Z(n5259) );
XOR U8767 ( .A(c1753), .B(b[1753]), .Z(n5260) );
XNOR U8768 ( .A(b[1753]), .B(n5261), .Z(c[1753]) );
XNOR U8769 ( .A(a[1753]), .B(c1753), .Z(n5261) );
XOR U8770 ( .A(c1754), .B(n5262), .Z(c1755) );
ANDN U8771 ( .B(n5263), .A(n5264), .Z(n5262) );
XOR U8772 ( .A(c1754), .B(b[1754]), .Z(n5263) );
XNOR U8773 ( .A(b[1754]), .B(n5264), .Z(c[1754]) );
XNOR U8774 ( .A(a[1754]), .B(c1754), .Z(n5264) );
XOR U8775 ( .A(c1755), .B(n5265), .Z(c1756) );
ANDN U8776 ( .B(n5266), .A(n5267), .Z(n5265) );
XOR U8777 ( .A(c1755), .B(b[1755]), .Z(n5266) );
XNOR U8778 ( .A(b[1755]), .B(n5267), .Z(c[1755]) );
XNOR U8779 ( .A(a[1755]), .B(c1755), .Z(n5267) );
XOR U8780 ( .A(c1756), .B(n5268), .Z(c1757) );
ANDN U8781 ( .B(n5269), .A(n5270), .Z(n5268) );
XOR U8782 ( .A(c1756), .B(b[1756]), .Z(n5269) );
XNOR U8783 ( .A(b[1756]), .B(n5270), .Z(c[1756]) );
XNOR U8784 ( .A(a[1756]), .B(c1756), .Z(n5270) );
XOR U8785 ( .A(c1757), .B(n5271), .Z(c1758) );
ANDN U8786 ( .B(n5272), .A(n5273), .Z(n5271) );
XOR U8787 ( .A(c1757), .B(b[1757]), .Z(n5272) );
XNOR U8788 ( .A(b[1757]), .B(n5273), .Z(c[1757]) );
XNOR U8789 ( .A(a[1757]), .B(c1757), .Z(n5273) );
XOR U8790 ( .A(c1758), .B(n5274), .Z(c1759) );
ANDN U8791 ( .B(n5275), .A(n5276), .Z(n5274) );
XOR U8792 ( .A(c1758), .B(b[1758]), .Z(n5275) );
XNOR U8793 ( .A(b[1758]), .B(n5276), .Z(c[1758]) );
XNOR U8794 ( .A(a[1758]), .B(c1758), .Z(n5276) );
XOR U8795 ( .A(c1759), .B(n5277), .Z(c1760) );
ANDN U8796 ( .B(n5278), .A(n5279), .Z(n5277) );
XOR U8797 ( .A(c1759), .B(b[1759]), .Z(n5278) );
XNOR U8798 ( .A(b[1759]), .B(n5279), .Z(c[1759]) );
XNOR U8799 ( .A(a[1759]), .B(c1759), .Z(n5279) );
XOR U8800 ( .A(c1760), .B(n5280), .Z(c1761) );
ANDN U8801 ( .B(n5281), .A(n5282), .Z(n5280) );
XOR U8802 ( .A(c1760), .B(b[1760]), .Z(n5281) );
XNOR U8803 ( .A(b[1760]), .B(n5282), .Z(c[1760]) );
XNOR U8804 ( .A(a[1760]), .B(c1760), .Z(n5282) );
XOR U8805 ( .A(c1761), .B(n5283), .Z(c1762) );
ANDN U8806 ( .B(n5284), .A(n5285), .Z(n5283) );
XOR U8807 ( .A(c1761), .B(b[1761]), .Z(n5284) );
XNOR U8808 ( .A(b[1761]), .B(n5285), .Z(c[1761]) );
XNOR U8809 ( .A(a[1761]), .B(c1761), .Z(n5285) );
XOR U8810 ( .A(c1762), .B(n5286), .Z(c1763) );
ANDN U8811 ( .B(n5287), .A(n5288), .Z(n5286) );
XOR U8812 ( .A(c1762), .B(b[1762]), .Z(n5287) );
XNOR U8813 ( .A(b[1762]), .B(n5288), .Z(c[1762]) );
XNOR U8814 ( .A(a[1762]), .B(c1762), .Z(n5288) );
XOR U8815 ( .A(c1763), .B(n5289), .Z(c1764) );
ANDN U8816 ( .B(n5290), .A(n5291), .Z(n5289) );
XOR U8817 ( .A(c1763), .B(b[1763]), .Z(n5290) );
XNOR U8818 ( .A(b[1763]), .B(n5291), .Z(c[1763]) );
XNOR U8819 ( .A(a[1763]), .B(c1763), .Z(n5291) );
XOR U8820 ( .A(c1764), .B(n5292), .Z(c1765) );
ANDN U8821 ( .B(n5293), .A(n5294), .Z(n5292) );
XOR U8822 ( .A(c1764), .B(b[1764]), .Z(n5293) );
XNOR U8823 ( .A(b[1764]), .B(n5294), .Z(c[1764]) );
XNOR U8824 ( .A(a[1764]), .B(c1764), .Z(n5294) );
XOR U8825 ( .A(c1765), .B(n5295), .Z(c1766) );
ANDN U8826 ( .B(n5296), .A(n5297), .Z(n5295) );
XOR U8827 ( .A(c1765), .B(b[1765]), .Z(n5296) );
XNOR U8828 ( .A(b[1765]), .B(n5297), .Z(c[1765]) );
XNOR U8829 ( .A(a[1765]), .B(c1765), .Z(n5297) );
XOR U8830 ( .A(c1766), .B(n5298), .Z(c1767) );
ANDN U8831 ( .B(n5299), .A(n5300), .Z(n5298) );
XOR U8832 ( .A(c1766), .B(b[1766]), .Z(n5299) );
XNOR U8833 ( .A(b[1766]), .B(n5300), .Z(c[1766]) );
XNOR U8834 ( .A(a[1766]), .B(c1766), .Z(n5300) );
XOR U8835 ( .A(c1767), .B(n5301), .Z(c1768) );
ANDN U8836 ( .B(n5302), .A(n5303), .Z(n5301) );
XOR U8837 ( .A(c1767), .B(b[1767]), .Z(n5302) );
XNOR U8838 ( .A(b[1767]), .B(n5303), .Z(c[1767]) );
XNOR U8839 ( .A(a[1767]), .B(c1767), .Z(n5303) );
XOR U8840 ( .A(c1768), .B(n5304), .Z(c1769) );
ANDN U8841 ( .B(n5305), .A(n5306), .Z(n5304) );
XOR U8842 ( .A(c1768), .B(b[1768]), .Z(n5305) );
XNOR U8843 ( .A(b[1768]), .B(n5306), .Z(c[1768]) );
XNOR U8844 ( .A(a[1768]), .B(c1768), .Z(n5306) );
XOR U8845 ( .A(c1769), .B(n5307), .Z(c1770) );
ANDN U8846 ( .B(n5308), .A(n5309), .Z(n5307) );
XOR U8847 ( .A(c1769), .B(b[1769]), .Z(n5308) );
XNOR U8848 ( .A(b[1769]), .B(n5309), .Z(c[1769]) );
XNOR U8849 ( .A(a[1769]), .B(c1769), .Z(n5309) );
XOR U8850 ( .A(c1770), .B(n5310), .Z(c1771) );
ANDN U8851 ( .B(n5311), .A(n5312), .Z(n5310) );
XOR U8852 ( .A(c1770), .B(b[1770]), .Z(n5311) );
XNOR U8853 ( .A(b[1770]), .B(n5312), .Z(c[1770]) );
XNOR U8854 ( .A(a[1770]), .B(c1770), .Z(n5312) );
XOR U8855 ( .A(c1771), .B(n5313), .Z(c1772) );
ANDN U8856 ( .B(n5314), .A(n5315), .Z(n5313) );
XOR U8857 ( .A(c1771), .B(b[1771]), .Z(n5314) );
XNOR U8858 ( .A(b[1771]), .B(n5315), .Z(c[1771]) );
XNOR U8859 ( .A(a[1771]), .B(c1771), .Z(n5315) );
XOR U8860 ( .A(c1772), .B(n5316), .Z(c1773) );
ANDN U8861 ( .B(n5317), .A(n5318), .Z(n5316) );
XOR U8862 ( .A(c1772), .B(b[1772]), .Z(n5317) );
XNOR U8863 ( .A(b[1772]), .B(n5318), .Z(c[1772]) );
XNOR U8864 ( .A(a[1772]), .B(c1772), .Z(n5318) );
XOR U8865 ( .A(c1773), .B(n5319), .Z(c1774) );
ANDN U8866 ( .B(n5320), .A(n5321), .Z(n5319) );
XOR U8867 ( .A(c1773), .B(b[1773]), .Z(n5320) );
XNOR U8868 ( .A(b[1773]), .B(n5321), .Z(c[1773]) );
XNOR U8869 ( .A(a[1773]), .B(c1773), .Z(n5321) );
XOR U8870 ( .A(c1774), .B(n5322), .Z(c1775) );
ANDN U8871 ( .B(n5323), .A(n5324), .Z(n5322) );
XOR U8872 ( .A(c1774), .B(b[1774]), .Z(n5323) );
XNOR U8873 ( .A(b[1774]), .B(n5324), .Z(c[1774]) );
XNOR U8874 ( .A(a[1774]), .B(c1774), .Z(n5324) );
XOR U8875 ( .A(c1775), .B(n5325), .Z(c1776) );
ANDN U8876 ( .B(n5326), .A(n5327), .Z(n5325) );
XOR U8877 ( .A(c1775), .B(b[1775]), .Z(n5326) );
XNOR U8878 ( .A(b[1775]), .B(n5327), .Z(c[1775]) );
XNOR U8879 ( .A(a[1775]), .B(c1775), .Z(n5327) );
XOR U8880 ( .A(c1776), .B(n5328), .Z(c1777) );
ANDN U8881 ( .B(n5329), .A(n5330), .Z(n5328) );
XOR U8882 ( .A(c1776), .B(b[1776]), .Z(n5329) );
XNOR U8883 ( .A(b[1776]), .B(n5330), .Z(c[1776]) );
XNOR U8884 ( .A(a[1776]), .B(c1776), .Z(n5330) );
XOR U8885 ( .A(c1777), .B(n5331), .Z(c1778) );
ANDN U8886 ( .B(n5332), .A(n5333), .Z(n5331) );
XOR U8887 ( .A(c1777), .B(b[1777]), .Z(n5332) );
XNOR U8888 ( .A(b[1777]), .B(n5333), .Z(c[1777]) );
XNOR U8889 ( .A(a[1777]), .B(c1777), .Z(n5333) );
XOR U8890 ( .A(c1778), .B(n5334), .Z(c1779) );
ANDN U8891 ( .B(n5335), .A(n5336), .Z(n5334) );
XOR U8892 ( .A(c1778), .B(b[1778]), .Z(n5335) );
XNOR U8893 ( .A(b[1778]), .B(n5336), .Z(c[1778]) );
XNOR U8894 ( .A(a[1778]), .B(c1778), .Z(n5336) );
XOR U8895 ( .A(c1779), .B(n5337), .Z(c1780) );
ANDN U8896 ( .B(n5338), .A(n5339), .Z(n5337) );
XOR U8897 ( .A(c1779), .B(b[1779]), .Z(n5338) );
XNOR U8898 ( .A(b[1779]), .B(n5339), .Z(c[1779]) );
XNOR U8899 ( .A(a[1779]), .B(c1779), .Z(n5339) );
XOR U8900 ( .A(c1780), .B(n5340), .Z(c1781) );
ANDN U8901 ( .B(n5341), .A(n5342), .Z(n5340) );
XOR U8902 ( .A(c1780), .B(b[1780]), .Z(n5341) );
XNOR U8903 ( .A(b[1780]), .B(n5342), .Z(c[1780]) );
XNOR U8904 ( .A(a[1780]), .B(c1780), .Z(n5342) );
XOR U8905 ( .A(c1781), .B(n5343), .Z(c1782) );
ANDN U8906 ( .B(n5344), .A(n5345), .Z(n5343) );
XOR U8907 ( .A(c1781), .B(b[1781]), .Z(n5344) );
XNOR U8908 ( .A(b[1781]), .B(n5345), .Z(c[1781]) );
XNOR U8909 ( .A(a[1781]), .B(c1781), .Z(n5345) );
XOR U8910 ( .A(c1782), .B(n5346), .Z(c1783) );
ANDN U8911 ( .B(n5347), .A(n5348), .Z(n5346) );
XOR U8912 ( .A(c1782), .B(b[1782]), .Z(n5347) );
XNOR U8913 ( .A(b[1782]), .B(n5348), .Z(c[1782]) );
XNOR U8914 ( .A(a[1782]), .B(c1782), .Z(n5348) );
XOR U8915 ( .A(c1783), .B(n5349), .Z(c1784) );
ANDN U8916 ( .B(n5350), .A(n5351), .Z(n5349) );
XOR U8917 ( .A(c1783), .B(b[1783]), .Z(n5350) );
XNOR U8918 ( .A(b[1783]), .B(n5351), .Z(c[1783]) );
XNOR U8919 ( .A(a[1783]), .B(c1783), .Z(n5351) );
XOR U8920 ( .A(c1784), .B(n5352), .Z(c1785) );
ANDN U8921 ( .B(n5353), .A(n5354), .Z(n5352) );
XOR U8922 ( .A(c1784), .B(b[1784]), .Z(n5353) );
XNOR U8923 ( .A(b[1784]), .B(n5354), .Z(c[1784]) );
XNOR U8924 ( .A(a[1784]), .B(c1784), .Z(n5354) );
XOR U8925 ( .A(c1785), .B(n5355), .Z(c1786) );
ANDN U8926 ( .B(n5356), .A(n5357), .Z(n5355) );
XOR U8927 ( .A(c1785), .B(b[1785]), .Z(n5356) );
XNOR U8928 ( .A(b[1785]), .B(n5357), .Z(c[1785]) );
XNOR U8929 ( .A(a[1785]), .B(c1785), .Z(n5357) );
XOR U8930 ( .A(c1786), .B(n5358), .Z(c1787) );
ANDN U8931 ( .B(n5359), .A(n5360), .Z(n5358) );
XOR U8932 ( .A(c1786), .B(b[1786]), .Z(n5359) );
XNOR U8933 ( .A(b[1786]), .B(n5360), .Z(c[1786]) );
XNOR U8934 ( .A(a[1786]), .B(c1786), .Z(n5360) );
XOR U8935 ( .A(c1787), .B(n5361), .Z(c1788) );
ANDN U8936 ( .B(n5362), .A(n5363), .Z(n5361) );
XOR U8937 ( .A(c1787), .B(b[1787]), .Z(n5362) );
XNOR U8938 ( .A(b[1787]), .B(n5363), .Z(c[1787]) );
XNOR U8939 ( .A(a[1787]), .B(c1787), .Z(n5363) );
XOR U8940 ( .A(c1788), .B(n5364), .Z(c1789) );
ANDN U8941 ( .B(n5365), .A(n5366), .Z(n5364) );
XOR U8942 ( .A(c1788), .B(b[1788]), .Z(n5365) );
XNOR U8943 ( .A(b[1788]), .B(n5366), .Z(c[1788]) );
XNOR U8944 ( .A(a[1788]), .B(c1788), .Z(n5366) );
XOR U8945 ( .A(c1789), .B(n5367), .Z(c1790) );
ANDN U8946 ( .B(n5368), .A(n5369), .Z(n5367) );
XOR U8947 ( .A(c1789), .B(b[1789]), .Z(n5368) );
XNOR U8948 ( .A(b[1789]), .B(n5369), .Z(c[1789]) );
XNOR U8949 ( .A(a[1789]), .B(c1789), .Z(n5369) );
XOR U8950 ( .A(c1790), .B(n5370), .Z(c1791) );
ANDN U8951 ( .B(n5371), .A(n5372), .Z(n5370) );
XOR U8952 ( .A(c1790), .B(b[1790]), .Z(n5371) );
XNOR U8953 ( .A(b[1790]), .B(n5372), .Z(c[1790]) );
XNOR U8954 ( .A(a[1790]), .B(c1790), .Z(n5372) );
XOR U8955 ( .A(c1791), .B(n5373), .Z(c1792) );
ANDN U8956 ( .B(n5374), .A(n5375), .Z(n5373) );
XOR U8957 ( .A(c1791), .B(b[1791]), .Z(n5374) );
XNOR U8958 ( .A(b[1791]), .B(n5375), .Z(c[1791]) );
XNOR U8959 ( .A(a[1791]), .B(c1791), .Z(n5375) );
XOR U8960 ( .A(c1792), .B(n5376), .Z(c1793) );
ANDN U8961 ( .B(n5377), .A(n5378), .Z(n5376) );
XOR U8962 ( .A(c1792), .B(b[1792]), .Z(n5377) );
XNOR U8963 ( .A(b[1792]), .B(n5378), .Z(c[1792]) );
XNOR U8964 ( .A(a[1792]), .B(c1792), .Z(n5378) );
XOR U8965 ( .A(c1793), .B(n5379), .Z(c1794) );
ANDN U8966 ( .B(n5380), .A(n5381), .Z(n5379) );
XOR U8967 ( .A(c1793), .B(b[1793]), .Z(n5380) );
XNOR U8968 ( .A(b[1793]), .B(n5381), .Z(c[1793]) );
XNOR U8969 ( .A(a[1793]), .B(c1793), .Z(n5381) );
XOR U8970 ( .A(c1794), .B(n5382), .Z(c1795) );
ANDN U8971 ( .B(n5383), .A(n5384), .Z(n5382) );
XOR U8972 ( .A(c1794), .B(b[1794]), .Z(n5383) );
XNOR U8973 ( .A(b[1794]), .B(n5384), .Z(c[1794]) );
XNOR U8974 ( .A(a[1794]), .B(c1794), .Z(n5384) );
XOR U8975 ( .A(c1795), .B(n5385), .Z(c1796) );
ANDN U8976 ( .B(n5386), .A(n5387), .Z(n5385) );
XOR U8977 ( .A(c1795), .B(b[1795]), .Z(n5386) );
XNOR U8978 ( .A(b[1795]), .B(n5387), .Z(c[1795]) );
XNOR U8979 ( .A(a[1795]), .B(c1795), .Z(n5387) );
XOR U8980 ( .A(c1796), .B(n5388), .Z(c1797) );
ANDN U8981 ( .B(n5389), .A(n5390), .Z(n5388) );
XOR U8982 ( .A(c1796), .B(b[1796]), .Z(n5389) );
XNOR U8983 ( .A(b[1796]), .B(n5390), .Z(c[1796]) );
XNOR U8984 ( .A(a[1796]), .B(c1796), .Z(n5390) );
XOR U8985 ( .A(c1797), .B(n5391), .Z(c1798) );
ANDN U8986 ( .B(n5392), .A(n5393), .Z(n5391) );
XOR U8987 ( .A(c1797), .B(b[1797]), .Z(n5392) );
XNOR U8988 ( .A(b[1797]), .B(n5393), .Z(c[1797]) );
XNOR U8989 ( .A(a[1797]), .B(c1797), .Z(n5393) );
XOR U8990 ( .A(c1798), .B(n5394), .Z(c1799) );
ANDN U8991 ( .B(n5395), .A(n5396), .Z(n5394) );
XOR U8992 ( .A(c1798), .B(b[1798]), .Z(n5395) );
XNOR U8993 ( .A(b[1798]), .B(n5396), .Z(c[1798]) );
XNOR U8994 ( .A(a[1798]), .B(c1798), .Z(n5396) );
XOR U8995 ( .A(c1799), .B(n5397), .Z(c1800) );
ANDN U8996 ( .B(n5398), .A(n5399), .Z(n5397) );
XOR U8997 ( .A(c1799), .B(b[1799]), .Z(n5398) );
XNOR U8998 ( .A(b[1799]), .B(n5399), .Z(c[1799]) );
XNOR U8999 ( .A(a[1799]), .B(c1799), .Z(n5399) );
XOR U9000 ( .A(c1800), .B(n5400), .Z(c1801) );
ANDN U9001 ( .B(n5401), .A(n5402), .Z(n5400) );
XOR U9002 ( .A(c1800), .B(b[1800]), .Z(n5401) );
XNOR U9003 ( .A(b[1800]), .B(n5402), .Z(c[1800]) );
XNOR U9004 ( .A(a[1800]), .B(c1800), .Z(n5402) );
XOR U9005 ( .A(c1801), .B(n5403), .Z(c1802) );
ANDN U9006 ( .B(n5404), .A(n5405), .Z(n5403) );
XOR U9007 ( .A(c1801), .B(b[1801]), .Z(n5404) );
XNOR U9008 ( .A(b[1801]), .B(n5405), .Z(c[1801]) );
XNOR U9009 ( .A(a[1801]), .B(c1801), .Z(n5405) );
XOR U9010 ( .A(c1802), .B(n5406), .Z(c1803) );
ANDN U9011 ( .B(n5407), .A(n5408), .Z(n5406) );
XOR U9012 ( .A(c1802), .B(b[1802]), .Z(n5407) );
XNOR U9013 ( .A(b[1802]), .B(n5408), .Z(c[1802]) );
XNOR U9014 ( .A(a[1802]), .B(c1802), .Z(n5408) );
XOR U9015 ( .A(c1803), .B(n5409), .Z(c1804) );
ANDN U9016 ( .B(n5410), .A(n5411), .Z(n5409) );
XOR U9017 ( .A(c1803), .B(b[1803]), .Z(n5410) );
XNOR U9018 ( .A(b[1803]), .B(n5411), .Z(c[1803]) );
XNOR U9019 ( .A(a[1803]), .B(c1803), .Z(n5411) );
XOR U9020 ( .A(c1804), .B(n5412), .Z(c1805) );
ANDN U9021 ( .B(n5413), .A(n5414), .Z(n5412) );
XOR U9022 ( .A(c1804), .B(b[1804]), .Z(n5413) );
XNOR U9023 ( .A(b[1804]), .B(n5414), .Z(c[1804]) );
XNOR U9024 ( .A(a[1804]), .B(c1804), .Z(n5414) );
XOR U9025 ( .A(c1805), .B(n5415), .Z(c1806) );
ANDN U9026 ( .B(n5416), .A(n5417), .Z(n5415) );
XOR U9027 ( .A(c1805), .B(b[1805]), .Z(n5416) );
XNOR U9028 ( .A(b[1805]), .B(n5417), .Z(c[1805]) );
XNOR U9029 ( .A(a[1805]), .B(c1805), .Z(n5417) );
XOR U9030 ( .A(c1806), .B(n5418), .Z(c1807) );
ANDN U9031 ( .B(n5419), .A(n5420), .Z(n5418) );
XOR U9032 ( .A(c1806), .B(b[1806]), .Z(n5419) );
XNOR U9033 ( .A(b[1806]), .B(n5420), .Z(c[1806]) );
XNOR U9034 ( .A(a[1806]), .B(c1806), .Z(n5420) );
XOR U9035 ( .A(c1807), .B(n5421), .Z(c1808) );
ANDN U9036 ( .B(n5422), .A(n5423), .Z(n5421) );
XOR U9037 ( .A(c1807), .B(b[1807]), .Z(n5422) );
XNOR U9038 ( .A(b[1807]), .B(n5423), .Z(c[1807]) );
XNOR U9039 ( .A(a[1807]), .B(c1807), .Z(n5423) );
XOR U9040 ( .A(c1808), .B(n5424), .Z(c1809) );
ANDN U9041 ( .B(n5425), .A(n5426), .Z(n5424) );
XOR U9042 ( .A(c1808), .B(b[1808]), .Z(n5425) );
XNOR U9043 ( .A(b[1808]), .B(n5426), .Z(c[1808]) );
XNOR U9044 ( .A(a[1808]), .B(c1808), .Z(n5426) );
XOR U9045 ( .A(c1809), .B(n5427), .Z(c1810) );
ANDN U9046 ( .B(n5428), .A(n5429), .Z(n5427) );
XOR U9047 ( .A(c1809), .B(b[1809]), .Z(n5428) );
XNOR U9048 ( .A(b[1809]), .B(n5429), .Z(c[1809]) );
XNOR U9049 ( .A(a[1809]), .B(c1809), .Z(n5429) );
XOR U9050 ( .A(c1810), .B(n5430), .Z(c1811) );
ANDN U9051 ( .B(n5431), .A(n5432), .Z(n5430) );
XOR U9052 ( .A(c1810), .B(b[1810]), .Z(n5431) );
XNOR U9053 ( .A(b[1810]), .B(n5432), .Z(c[1810]) );
XNOR U9054 ( .A(a[1810]), .B(c1810), .Z(n5432) );
XOR U9055 ( .A(c1811), .B(n5433), .Z(c1812) );
ANDN U9056 ( .B(n5434), .A(n5435), .Z(n5433) );
XOR U9057 ( .A(c1811), .B(b[1811]), .Z(n5434) );
XNOR U9058 ( .A(b[1811]), .B(n5435), .Z(c[1811]) );
XNOR U9059 ( .A(a[1811]), .B(c1811), .Z(n5435) );
XOR U9060 ( .A(c1812), .B(n5436), .Z(c1813) );
ANDN U9061 ( .B(n5437), .A(n5438), .Z(n5436) );
XOR U9062 ( .A(c1812), .B(b[1812]), .Z(n5437) );
XNOR U9063 ( .A(b[1812]), .B(n5438), .Z(c[1812]) );
XNOR U9064 ( .A(a[1812]), .B(c1812), .Z(n5438) );
XOR U9065 ( .A(c1813), .B(n5439), .Z(c1814) );
ANDN U9066 ( .B(n5440), .A(n5441), .Z(n5439) );
XOR U9067 ( .A(c1813), .B(b[1813]), .Z(n5440) );
XNOR U9068 ( .A(b[1813]), .B(n5441), .Z(c[1813]) );
XNOR U9069 ( .A(a[1813]), .B(c1813), .Z(n5441) );
XOR U9070 ( .A(c1814), .B(n5442), .Z(c1815) );
ANDN U9071 ( .B(n5443), .A(n5444), .Z(n5442) );
XOR U9072 ( .A(c1814), .B(b[1814]), .Z(n5443) );
XNOR U9073 ( .A(b[1814]), .B(n5444), .Z(c[1814]) );
XNOR U9074 ( .A(a[1814]), .B(c1814), .Z(n5444) );
XOR U9075 ( .A(c1815), .B(n5445), .Z(c1816) );
ANDN U9076 ( .B(n5446), .A(n5447), .Z(n5445) );
XOR U9077 ( .A(c1815), .B(b[1815]), .Z(n5446) );
XNOR U9078 ( .A(b[1815]), .B(n5447), .Z(c[1815]) );
XNOR U9079 ( .A(a[1815]), .B(c1815), .Z(n5447) );
XOR U9080 ( .A(c1816), .B(n5448), .Z(c1817) );
ANDN U9081 ( .B(n5449), .A(n5450), .Z(n5448) );
XOR U9082 ( .A(c1816), .B(b[1816]), .Z(n5449) );
XNOR U9083 ( .A(b[1816]), .B(n5450), .Z(c[1816]) );
XNOR U9084 ( .A(a[1816]), .B(c1816), .Z(n5450) );
XOR U9085 ( .A(c1817), .B(n5451), .Z(c1818) );
ANDN U9086 ( .B(n5452), .A(n5453), .Z(n5451) );
XOR U9087 ( .A(c1817), .B(b[1817]), .Z(n5452) );
XNOR U9088 ( .A(b[1817]), .B(n5453), .Z(c[1817]) );
XNOR U9089 ( .A(a[1817]), .B(c1817), .Z(n5453) );
XOR U9090 ( .A(c1818), .B(n5454), .Z(c1819) );
ANDN U9091 ( .B(n5455), .A(n5456), .Z(n5454) );
XOR U9092 ( .A(c1818), .B(b[1818]), .Z(n5455) );
XNOR U9093 ( .A(b[1818]), .B(n5456), .Z(c[1818]) );
XNOR U9094 ( .A(a[1818]), .B(c1818), .Z(n5456) );
XOR U9095 ( .A(c1819), .B(n5457), .Z(c1820) );
ANDN U9096 ( .B(n5458), .A(n5459), .Z(n5457) );
XOR U9097 ( .A(c1819), .B(b[1819]), .Z(n5458) );
XNOR U9098 ( .A(b[1819]), .B(n5459), .Z(c[1819]) );
XNOR U9099 ( .A(a[1819]), .B(c1819), .Z(n5459) );
XOR U9100 ( .A(c1820), .B(n5460), .Z(c1821) );
ANDN U9101 ( .B(n5461), .A(n5462), .Z(n5460) );
XOR U9102 ( .A(c1820), .B(b[1820]), .Z(n5461) );
XNOR U9103 ( .A(b[1820]), .B(n5462), .Z(c[1820]) );
XNOR U9104 ( .A(a[1820]), .B(c1820), .Z(n5462) );
XOR U9105 ( .A(c1821), .B(n5463), .Z(c1822) );
ANDN U9106 ( .B(n5464), .A(n5465), .Z(n5463) );
XOR U9107 ( .A(c1821), .B(b[1821]), .Z(n5464) );
XNOR U9108 ( .A(b[1821]), .B(n5465), .Z(c[1821]) );
XNOR U9109 ( .A(a[1821]), .B(c1821), .Z(n5465) );
XOR U9110 ( .A(c1822), .B(n5466), .Z(c1823) );
ANDN U9111 ( .B(n5467), .A(n5468), .Z(n5466) );
XOR U9112 ( .A(c1822), .B(b[1822]), .Z(n5467) );
XNOR U9113 ( .A(b[1822]), .B(n5468), .Z(c[1822]) );
XNOR U9114 ( .A(a[1822]), .B(c1822), .Z(n5468) );
XOR U9115 ( .A(c1823), .B(n5469), .Z(c1824) );
ANDN U9116 ( .B(n5470), .A(n5471), .Z(n5469) );
XOR U9117 ( .A(c1823), .B(b[1823]), .Z(n5470) );
XNOR U9118 ( .A(b[1823]), .B(n5471), .Z(c[1823]) );
XNOR U9119 ( .A(a[1823]), .B(c1823), .Z(n5471) );
XOR U9120 ( .A(c1824), .B(n5472), .Z(c1825) );
ANDN U9121 ( .B(n5473), .A(n5474), .Z(n5472) );
XOR U9122 ( .A(c1824), .B(b[1824]), .Z(n5473) );
XNOR U9123 ( .A(b[1824]), .B(n5474), .Z(c[1824]) );
XNOR U9124 ( .A(a[1824]), .B(c1824), .Z(n5474) );
XOR U9125 ( .A(c1825), .B(n5475), .Z(c1826) );
ANDN U9126 ( .B(n5476), .A(n5477), .Z(n5475) );
XOR U9127 ( .A(c1825), .B(b[1825]), .Z(n5476) );
XNOR U9128 ( .A(b[1825]), .B(n5477), .Z(c[1825]) );
XNOR U9129 ( .A(a[1825]), .B(c1825), .Z(n5477) );
XOR U9130 ( .A(c1826), .B(n5478), .Z(c1827) );
ANDN U9131 ( .B(n5479), .A(n5480), .Z(n5478) );
XOR U9132 ( .A(c1826), .B(b[1826]), .Z(n5479) );
XNOR U9133 ( .A(b[1826]), .B(n5480), .Z(c[1826]) );
XNOR U9134 ( .A(a[1826]), .B(c1826), .Z(n5480) );
XOR U9135 ( .A(c1827), .B(n5481), .Z(c1828) );
ANDN U9136 ( .B(n5482), .A(n5483), .Z(n5481) );
XOR U9137 ( .A(c1827), .B(b[1827]), .Z(n5482) );
XNOR U9138 ( .A(b[1827]), .B(n5483), .Z(c[1827]) );
XNOR U9139 ( .A(a[1827]), .B(c1827), .Z(n5483) );
XOR U9140 ( .A(c1828), .B(n5484), .Z(c1829) );
ANDN U9141 ( .B(n5485), .A(n5486), .Z(n5484) );
XOR U9142 ( .A(c1828), .B(b[1828]), .Z(n5485) );
XNOR U9143 ( .A(b[1828]), .B(n5486), .Z(c[1828]) );
XNOR U9144 ( .A(a[1828]), .B(c1828), .Z(n5486) );
XOR U9145 ( .A(c1829), .B(n5487), .Z(c1830) );
ANDN U9146 ( .B(n5488), .A(n5489), .Z(n5487) );
XOR U9147 ( .A(c1829), .B(b[1829]), .Z(n5488) );
XNOR U9148 ( .A(b[1829]), .B(n5489), .Z(c[1829]) );
XNOR U9149 ( .A(a[1829]), .B(c1829), .Z(n5489) );
XOR U9150 ( .A(c1830), .B(n5490), .Z(c1831) );
ANDN U9151 ( .B(n5491), .A(n5492), .Z(n5490) );
XOR U9152 ( .A(c1830), .B(b[1830]), .Z(n5491) );
XNOR U9153 ( .A(b[1830]), .B(n5492), .Z(c[1830]) );
XNOR U9154 ( .A(a[1830]), .B(c1830), .Z(n5492) );
XOR U9155 ( .A(c1831), .B(n5493), .Z(c1832) );
ANDN U9156 ( .B(n5494), .A(n5495), .Z(n5493) );
XOR U9157 ( .A(c1831), .B(b[1831]), .Z(n5494) );
XNOR U9158 ( .A(b[1831]), .B(n5495), .Z(c[1831]) );
XNOR U9159 ( .A(a[1831]), .B(c1831), .Z(n5495) );
XOR U9160 ( .A(c1832), .B(n5496), .Z(c1833) );
ANDN U9161 ( .B(n5497), .A(n5498), .Z(n5496) );
XOR U9162 ( .A(c1832), .B(b[1832]), .Z(n5497) );
XNOR U9163 ( .A(b[1832]), .B(n5498), .Z(c[1832]) );
XNOR U9164 ( .A(a[1832]), .B(c1832), .Z(n5498) );
XOR U9165 ( .A(c1833), .B(n5499), .Z(c1834) );
ANDN U9166 ( .B(n5500), .A(n5501), .Z(n5499) );
XOR U9167 ( .A(c1833), .B(b[1833]), .Z(n5500) );
XNOR U9168 ( .A(b[1833]), .B(n5501), .Z(c[1833]) );
XNOR U9169 ( .A(a[1833]), .B(c1833), .Z(n5501) );
XOR U9170 ( .A(c1834), .B(n5502), .Z(c1835) );
ANDN U9171 ( .B(n5503), .A(n5504), .Z(n5502) );
XOR U9172 ( .A(c1834), .B(b[1834]), .Z(n5503) );
XNOR U9173 ( .A(b[1834]), .B(n5504), .Z(c[1834]) );
XNOR U9174 ( .A(a[1834]), .B(c1834), .Z(n5504) );
XOR U9175 ( .A(c1835), .B(n5505), .Z(c1836) );
ANDN U9176 ( .B(n5506), .A(n5507), .Z(n5505) );
XOR U9177 ( .A(c1835), .B(b[1835]), .Z(n5506) );
XNOR U9178 ( .A(b[1835]), .B(n5507), .Z(c[1835]) );
XNOR U9179 ( .A(a[1835]), .B(c1835), .Z(n5507) );
XOR U9180 ( .A(c1836), .B(n5508), .Z(c1837) );
ANDN U9181 ( .B(n5509), .A(n5510), .Z(n5508) );
XOR U9182 ( .A(c1836), .B(b[1836]), .Z(n5509) );
XNOR U9183 ( .A(b[1836]), .B(n5510), .Z(c[1836]) );
XNOR U9184 ( .A(a[1836]), .B(c1836), .Z(n5510) );
XOR U9185 ( .A(c1837), .B(n5511), .Z(c1838) );
ANDN U9186 ( .B(n5512), .A(n5513), .Z(n5511) );
XOR U9187 ( .A(c1837), .B(b[1837]), .Z(n5512) );
XNOR U9188 ( .A(b[1837]), .B(n5513), .Z(c[1837]) );
XNOR U9189 ( .A(a[1837]), .B(c1837), .Z(n5513) );
XOR U9190 ( .A(c1838), .B(n5514), .Z(c1839) );
ANDN U9191 ( .B(n5515), .A(n5516), .Z(n5514) );
XOR U9192 ( .A(c1838), .B(b[1838]), .Z(n5515) );
XNOR U9193 ( .A(b[1838]), .B(n5516), .Z(c[1838]) );
XNOR U9194 ( .A(a[1838]), .B(c1838), .Z(n5516) );
XOR U9195 ( .A(c1839), .B(n5517), .Z(c1840) );
ANDN U9196 ( .B(n5518), .A(n5519), .Z(n5517) );
XOR U9197 ( .A(c1839), .B(b[1839]), .Z(n5518) );
XNOR U9198 ( .A(b[1839]), .B(n5519), .Z(c[1839]) );
XNOR U9199 ( .A(a[1839]), .B(c1839), .Z(n5519) );
XOR U9200 ( .A(c1840), .B(n5520), .Z(c1841) );
ANDN U9201 ( .B(n5521), .A(n5522), .Z(n5520) );
XOR U9202 ( .A(c1840), .B(b[1840]), .Z(n5521) );
XNOR U9203 ( .A(b[1840]), .B(n5522), .Z(c[1840]) );
XNOR U9204 ( .A(a[1840]), .B(c1840), .Z(n5522) );
XOR U9205 ( .A(c1841), .B(n5523), .Z(c1842) );
ANDN U9206 ( .B(n5524), .A(n5525), .Z(n5523) );
XOR U9207 ( .A(c1841), .B(b[1841]), .Z(n5524) );
XNOR U9208 ( .A(b[1841]), .B(n5525), .Z(c[1841]) );
XNOR U9209 ( .A(a[1841]), .B(c1841), .Z(n5525) );
XOR U9210 ( .A(c1842), .B(n5526), .Z(c1843) );
ANDN U9211 ( .B(n5527), .A(n5528), .Z(n5526) );
XOR U9212 ( .A(c1842), .B(b[1842]), .Z(n5527) );
XNOR U9213 ( .A(b[1842]), .B(n5528), .Z(c[1842]) );
XNOR U9214 ( .A(a[1842]), .B(c1842), .Z(n5528) );
XOR U9215 ( .A(c1843), .B(n5529), .Z(c1844) );
ANDN U9216 ( .B(n5530), .A(n5531), .Z(n5529) );
XOR U9217 ( .A(c1843), .B(b[1843]), .Z(n5530) );
XNOR U9218 ( .A(b[1843]), .B(n5531), .Z(c[1843]) );
XNOR U9219 ( .A(a[1843]), .B(c1843), .Z(n5531) );
XOR U9220 ( .A(c1844), .B(n5532), .Z(c1845) );
ANDN U9221 ( .B(n5533), .A(n5534), .Z(n5532) );
XOR U9222 ( .A(c1844), .B(b[1844]), .Z(n5533) );
XNOR U9223 ( .A(b[1844]), .B(n5534), .Z(c[1844]) );
XNOR U9224 ( .A(a[1844]), .B(c1844), .Z(n5534) );
XOR U9225 ( .A(c1845), .B(n5535), .Z(c1846) );
ANDN U9226 ( .B(n5536), .A(n5537), .Z(n5535) );
XOR U9227 ( .A(c1845), .B(b[1845]), .Z(n5536) );
XNOR U9228 ( .A(b[1845]), .B(n5537), .Z(c[1845]) );
XNOR U9229 ( .A(a[1845]), .B(c1845), .Z(n5537) );
XOR U9230 ( .A(c1846), .B(n5538), .Z(c1847) );
ANDN U9231 ( .B(n5539), .A(n5540), .Z(n5538) );
XOR U9232 ( .A(c1846), .B(b[1846]), .Z(n5539) );
XNOR U9233 ( .A(b[1846]), .B(n5540), .Z(c[1846]) );
XNOR U9234 ( .A(a[1846]), .B(c1846), .Z(n5540) );
XOR U9235 ( .A(c1847), .B(n5541), .Z(c1848) );
ANDN U9236 ( .B(n5542), .A(n5543), .Z(n5541) );
XOR U9237 ( .A(c1847), .B(b[1847]), .Z(n5542) );
XNOR U9238 ( .A(b[1847]), .B(n5543), .Z(c[1847]) );
XNOR U9239 ( .A(a[1847]), .B(c1847), .Z(n5543) );
XOR U9240 ( .A(c1848), .B(n5544), .Z(c1849) );
ANDN U9241 ( .B(n5545), .A(n5546), .Z(n5544) );
XOR U9242 ( .A(c1848), .B(b[1848]), .Z(n5545) );
XNOR U9243 ( .A(b[1848]), .B(n5546), .Z(c[1848]) );
XNOR U9244 ( .A(a[1848]), .B(c1848), .Z(n5546) );
XOR U9245 ( .A(c1849), .B(n5547), .Z(c1850) );
ANDN U9246 ( .B(n5548), .A(n5549), .Z(n5547) );
XOR U9247 ( .A(c1849), .B(b[1849]), .Z(n5548) );
XNOR U9248 ( .A(b[1849]), .B(n5549), .Z(c[1849]) );
XNOR U9249 ( .A(a[1849]), .B(c1849), .Z(n5549) );
XOR U9250 ( .A(c1850), .B(n5550), .Z(c1851) );
ANDN U9251 ( .B(n5551), .A(n5552), .Z(n5550) );
XOR U9252 ( .A(c1850), .B(b[1850]), .Z(n5551) );
XNOR U9253 ( .A(b[1850]), .B(n5552), .Z(c[1850]) );
XNOR U9254 ( .A(a[1850]), .B(c1850), .Z(n5552) );
XOR U9255 ( .A(c1851), .B(n5553), .Z(c1852) );
ANDN U9256 ( .B(n5554), .A(n5555), .Z(n5553) );
XOR U9257 ( .A(c1851), .B(b[1851]), .Z(n5554) );
XNOR U9258 ( .A(b[1851]), .B(n5555), .Z(c[1851]) );
XNOR U9259 ( .A(a[1851]), .B(c1851), .Z(n5555) );
XOR U9260 ( .A(c1852), .B(n5556), .Z(c1853) );
ANDN U9261 ( .B(n5557), .A(n5558), .Z(n5556) );
XOR U9262 ( .A(c1852), .B(b[1852]), .Z(n5557) );
XNOR U9263 ( .A(b[1852]), .B(n5558), .Z(c[1852]) );
XNOR U9264 ( .A(a[1852]), .B(c1852), .Z(n5558) );
XOR U9265 ( .A(c1853), .B(n5559), .Z(c1854) );
ANDN U9266 ( .B(n5560), .A(n5561), .Z(n5559) );
XOR U9267 ( .A(c1853), .B(b[1853]), .Z(n5560) );
XNOR U9268 ( .A(b[1853]), .B(n5561), .Z(c[1853]) );
XNOR U9269 ( .A(a[1853]), .B(c1853), .Z(n5561) );
XOR U9270 ( .A(c1854), .B(n5562), .Z(c1855) );
ANDN U9271 ( .B(n5563), .A(n5564), .Z(n5562) );
XOR U9272 ( .A(c1854), .B(b[1854]), .Z(n5563) );
XNOR U9273 ( .A(b[1854]), .B(n5564), .Z(c[1854]) );
XNOR U9274 ( .A(a[1854]), .B(c1854), .Z(n5564) );
XOR U9275 ( .A(c1855), .B(n5565), .Z(c1856) );
ANDN U9276 ( .B(n5566), .A(n5567), .Z(n5565) );
XOR U9277 ( .A(c1855), .B(b[1855]), .Z(n5566) );
XNOR U9278 ( .A(b[1855]), .B(n5567), .Z(c[1855]) );
XNOR U9279 ( .A(a[1855]), .B(c1855), .Z(n5567) );
XOR U9280 ( .A(c1856), .B(n5568), .Z(c1857) );
ANDN U9281 ( .B(n5569), .A(n5570), .Z(n5568) );
XOR U9282 ( .A(c1856), .B(b[1856]), .Z(n5569) );
XNOR U9283 ( .A(b[1856]), .B(n5570), .Z(c[1856]) );
XNOR U9284 ( .A(a[1856]), .B(c1856), .Z(n5570) );
XOR U9285 ( .A(c1857), .B(n5571), .Z(c1858) );
ANDN U9286 ( .B(n5572), .A(n5573), .Z(n5571) );
XOR U9287 ( .A(c1857), .B(b[1857]), .Z(n5572) );
XNOR U9288 ( .A(b[1857]), .B(n5573), .Z(c[1857]) );
XNOR U9289 ( .A(a[1857]), .B(c1857), .Z(n5573) );
XOR U9290 ( .A(c1858), .B(n5574), .Z(c1859) );
ANDN U9291 ( .B(n5575), .A(n5576), .Z(n5574) );
XOR U9292 ( .A(c1858), .B(b[1858]), .Z(n5575) );
XNOR U9293 ( .A(b[1858]), .B(n5576), .Z(c[1858]) );
XNOR U9294 ( .A(a[1858]), .B(c1858), .Z(n5576) );
XOR U9295 ( .A(c1859), .B(n5577), .Z(c1860) );
ANDN U9296 ( .B(n5578), .A(n5579), .Z(n5577) );
XOR U9297 ( .A(c1859), .B(b[1859]), .Z(n5578) );
XNOR U9298 ( .A(b[1859]), .B(n5579), .Z(c[1859]) );
XNOR U9299 ( .A(a[1859]), .B(c1859), .Z(n5579) );
XOR U9300 ( .A(c1860), .B(n5580), .Z(c1861) );
ANDN U9301 ( .B(n5581), .A(n5582), .Z(n5580) );
XOR U9302 ( .A(c1860), .B(b[1860]), .Z(n5581) );
XNOR U9303 ( .A(b[1860]), .B(n5582), .Z(c[1860]) );
XNOR U9304 ( .A(a[1860]), .B(c1860), .Z(n5582) );
XOR U9305 ( .A(c1861), .B(n5583), .Z(c1862) );
ANDN U9306 ( .B(n5584), .A(n5585), .Z(n5583) );
XOR U9307 ( .A(c1861), .B(b[1861]), .Z(n5584) );
XNOR U9308 ( .A(b[1861]), .B(n5585), .Z(c[1861]) );
XNOR U9309 ( .A(a[1861]), .B(c1861), .Z(n5585) );
XOR U9310 ( .A(c1862), .B(n5586), .Z(c1863) );
ANDN U9311 ( .B(n5587), .A(n5588), .Z(n5586) );
XOR U9312 ( .A(c1862), .B(b[1862]), .Z(n5587) );
XNOR U9313 ( .A(b[1862]), .B(n5588), .Z(c[1862]) );
XNOR U9314 ( .A(a[1862]), .B(c1862), .Z(n5588) );
XOR U9315 ( .A(c1863), .B(n5589), .Z(c1864) );
ANDN U9316 ( .B(n5590), .A(n5591), .Z(n5589) );
XOR U9317 ( .A(c1863), .B(b[1863]), .Z(n5590) );
XNOR U9318 ( .A(b[1863]), .B(n5591), .Z(c[1863]) );
XNOR U9319 ( .A(a[1863]), .B(c1863), .Z(n5591) );
XOR U9320 ( .A(c1864), .B(n5592), .Z(c1865) );
ANDN U9321 ( .B(n5593), .A(n5594), .Z(n5592) );
XOR U9322 ( .A(c1864), .B(b[1864]), .Z(n5593) );
XNOR U9323 ( .A(b[1864]), .B(n5594), .Z(c[1864]) );
XNOR U9324 ( .A(a[1864]), .B(c1864), .Z(n5594) );
XOR U9325 ( .A(c1865), .B(n5595), .Z(c1866) );
ANDN U9326 ( .B(n5596), .A(n5597), .Z(n5595) );
XOR U9327 ( .A(c1865), .B(b[1865]), .Z(n5596) );
XNOR U9328 ( .A(b[1865]), .B(n5597), .Z(c[1865]) );
XNOR U9329 ( .A(a[1865]), .B(c1865), .Z(n5597) );
XOR U9330 ( .A(c1866), .B(n5598), .Z(c1867) );
ANDN U9331 ( .B(n5599), .A(n5600), .Z(n5598) );
XOR U9332 ( .A(c1866), .B(b[1866]), .Z(n5599) );
XNOR U9333 ( .A(b[1866]), .B(n5600), .Z(c[1866]) );
XNOR U9334 ( .A(a[1866]), .B(c1866), .Z(n5600) );
XOR U9335 ( .A(c1867), .B(n5601), .Z(c1868) );
ANDN U9336 ( .B(n5602), .A(n5603), .Z(n5601) );
XOR U9337 ( .A(c1867), .B(b[1867]), .Z(n5602) );
XNOR U9338 ( .A(b[1867]), .B(n5603), .Z(c[1867]) );
XNOR U9339 ( .A(a[1867]), .B(c1867), .Z(n5603) );
XOR U9340 ( .A(c1868), .B(n5604), .Z(c1869) );
ANDN U9341 ( .B(n5605), .A(n5606), .Z(n5604) );
XOR U9342 ( .A(c1868), .B(b[1868]), .Z(n5605) );
XNOR U9343 ( .A(b[1868]), .B(n5606), .Z(c[1868]) );
XNOR U9344 ( .A(a[1868]), .B(c1868), .Z(n5606) );
XOR U9345 ( .A(c1869), .B(n5607), .Z(c1870) );
ANDN U9346 ( .B(n5608), .A(n5609), .Z(n5607) );
XOR U9347 ( .A(c1869), .B(b[1869]), .Z(n5608) );
XNOR U9348 ( .A(b[1869]), .B(n5609), .Z(c[1869]) );
XNOR U9349 ( .A(a[1869]), .B(c1869), .Z(n5609) );
XOR U9350 ( .A(c1870), .B(n5610), .Z(c1871) );
ANDN U9351 ( .B(n5611), .A(n5612), .Z(n5610) );
XOR U9352 ( .A(c1870), .B(b[1870]), .Z(n5611) );
XNOR U9353 ( .A(b[1870]), .B(n5612), .Z(c[1870]) );
XNOR U9354 ( .A(a[1870]), .B(c1870), .Z(n5612) );
XOR U9355 ( .A(c1871), .B(n5613), .Z(c1872) );
ANDN U9356 ( .B(n5614), .A(n5615), .Z(n5613) );
XOR U9357 ( .A(c1871), .B(b[1871]), .Z(n5614) );
XNOR U9358 ( .A(b[1871]), .B(n5615), .Z(c[1871]) );
XNOR U9359 ( .A(a[1871]), .B(c1871), .Z(n5615) );
XOR U9360 ( .A(c1872), .B(n5616), .Z(c1873) );
ANDN U9361 ( .B(n5617), .A(n5618), .Z(n5616) );
XOR U9362 ( .A(c1872), .B(b[1872]), .Z(n5617) );
XNOR U9363 ( .A(b[1872]), .B(n5618), .Z(c[1872]) );
XNOR U9364 ( .A(a[1872]), .B(c1872), .Z(n5618) );
XOR U9365 ( .A(c1873), .B(n5619), .Z(c1874) );
ANDN U9366 ( .B(n5620), .A(n5621), .Z(n5619) );
XOR U9367 ( .A(c1873), .B(b[1873]), .Z(n5620) );
XNOR U9368 ( .A(b[1873]), .B(n5621), .Z(c[1873]) );
XNOR U9369 ( .A(a[1873]), .B(c1873), .Z(n5621) );
XOR U9370 ( .A(c1874), .B(n5622), .Z(c1875) );
ANDN U9371 ( .B(n5623), .A(n5624), .Z(n5622) );
XOR U9372 ( .A(c1874), .B(b[1874]), .Z(n5623) );
XNOR U9373 ( .A(b[1874]), .B(n5624), .Z(c[1874]) );
XNOR U9374 ( .A(a[1874]), .B(c1874), .Z(n5624) );
XOR U9375 ( .A(c1875), .B(n5625), .Z(c1876) );
ANDN U9376 ( .B(n5626), .A(n5627), .Z(n5625) );
XOR U9377 ( .A(c1875), .B(b[1875]), .Z(n5626) );
XNOR U9378 ( .A(b[1875]), .B(n5627), .Z(c[1875]) );
XNOR U9379 ( .A(a[1875]), .B(c1875), .Z(n5627) );
XOR U9380 ( .A(c1876), .B(n5628), .Z(c1877) );
ANDN U9381 ( .B(n5629), .A(n5630), .Z(n5628) );
XOR U9382 ( .A(c1876), .B(b[1876]), .Z(n5629) );
XNOR U9383 ( .A(b[1876]), .B(n5630), .Z(c[1876]) );
XNOR U9384 ( .A(a[1876]), .B(c1876), .Z(n5630) );
XOR U9385 ( .A(c1877), .B(n5631), .Z(c1878) );
ANDN U9386 ( .B(n5632), .A(n5633), .Z(n5631) );
XOR U9387 ( .A(c1877), .B(b[1877]), .Z(n5632) );
XNOR U9388 ( .A(b[1877]), .B(n5633), .Z(c[1877]) );
XNOR U9389 ( .A(a[1877]), .B(c1877), .Z(n5633) );
XOR U9390 ( .A(c1878), .B(n5634), .Z(c1879) );
ANDN U9391 ( .B(n5635), .A(n5636), .Z(n5634) );
XOR U9392 ( .A(c1878), .B(b[1878]), .Z(n5635) );
XNOR U9393 ( .A(b[1878]), .B(n5636), .Z(c[1878]) );
XNOR U9394 ( .A(a[1878]), .B(c1878), .Z(n5636) );
XOR U9395 ( .A(c1879), .B(n5637), .Z(c1880) );
ANDN U9396 ( .B(n5638), .A(n5639), .Z(n5637) );
XOR U9397 ( .A(c1879), .B(b[1879]), .Z(n5638) );
XNOR U9398 ( .A(b[1879]), .B(n5639), .Z(c[1879]) );
XNOR U9399 ( .A(a[1879]), .B(c1879), .Z(n5639) );
XOR U9400 ( .A(c1880), .B(n5640), .Z(c1881) );
ANDN U9401 ( .B(n5641), .A(n5642), .Z(n5640) );
XOR U9402 ( .A(c1880), .B(b[1880]), .Z(n5641) );
XNOR U9403 ( .A(b[1880]), .B(n5642), .Z(c[1880]) );
XNOR U9404 ( .A(a[1880]), .B(c1880), .Z(n5642) );
XOR U9405 ( .A(c1881), .B(n5643), .Z(c1882) );
ANDN U9406 ( .B(n5644), .A(n5645), .Z(n5643) );
XOR U9407 ( .A(c1881), .B(b[1881]), .Z(n5644) );
XNOR U9408 ( .A(b[1881]), .B(n5645), .Z(c[1881]) );
XNOR U9409 ( .A(a[1881]), .B(c1881), .Z(n5645) );
XOR U9410 ( .A(c1882), .B(n5646), .Z(c1883) );
ANDN U9411 ( .B(n5647), .A(n5648), .Z(n5646) );
XOR U9412 ( .A(c1882), .B(b[1882]), .Z(n5647) );
XNOR U9413 ( .A(b[1882]), .B(n5648), .Z(c[1882]) );
XNOR U9414 ( .A(a[1882]), .B(c1882), .Z(n5648) );
XOR U9415 ( .A(c1883), .B(n5649), .Z(c1884) );
ANDN U9416 ( .B(n5650), .A(n5651), .Z(n5649) );
XOR U9417 ( .A(c1883), .B(b[1883]), .Z(n5650) );
XNOR U9418 ( .A(b[1883]), .B(n5651), .Z(c[1883]) );
XNOR U9419 ( .A(a[1883]), .B(c1883), .Z(n5651) );
XOR U9420 ( .A(c1884), .B(n5652), .Z(c1885) );
ANDN U9421 ( .B(n5653), .A(n5654), .Z(n5652) );
XOR U9422 ( .A(c1884), .B(b[1884]), .Z(n5653) );
XNOR U9423 ( .A(b[1884]), .B(n5654), .Z(c[1884]) );
XNOR U9424 ( .A(a[1884]), .B(c1884), .Z(n5654) );
XOR U9425 ( .A(c1885), .B(n5655), .Z(c1886) );
ANDN U9426 ( .B(n5656), .A(n5657), .Z(n5655) );
XOR U9427 ( .A(c1885), .B(b[1885]), .Z(n5656) );
XNOR U9428 ( .A(b[1885]), .B(n5657), .Z(c[1885]) );
XNOR U9429 ( .A(a[1885]), .B(c1885), .Z(n5657) );
XOR U9430 ( .A(c1886), .B(n5658), .Z(c1887) );
ANDN U9431 ( .B(n5659), .A(n5660), .Z(n5658) );
XOR U9432 ( .A(c1886), .B(b[1886]), .Z(n5659) );
XNOR U9433 ( .A(b[1886]), .B(n5660), .Z(c[1886]) );
XNOR U9434 ( .A(a[1886]), .B(c1886), .Z(n5660) );
XOR U9435 ( .A(c1887), .B(n5661), .Z(c1888) );
ANDN U9436 ( .B(n5662), .A(n5663), .Z(n5661) );
XOR U9437 ( .A(c1887), .B(b[1887]), .Z(n5662) );
XNOR U9438 ( .A(b[1887]), .B(n5663), .Z(c[1887]) );
XNOR U9439 ( .A(a[1887]), .B(c1887), .Z(n5663) );
XOR U9440 ( .A(c1888), .B(n5664), .Z(c1889) );
ANDN U9441 ( .B(n5665), .A(n5666), .Z(n5664) );
XOR U9442 ( .A(c1888), .B(b[1888]), .Z(n5665) );
XNOR U9443 ( .A(b[1888]), .B(n5666), .Z(c[1888]) );
XNOR U9444 ( .A(a[1888]), .B(c1888), .Z(n5666) );
XOR U9445 ( .A(c1889), .B(n5667), .Z(c1890) );
ANDN U9446 ( .B(n5668), .A(n5669), .Z(n5667) );
XOR U9447 ( .A(c1889), .B(b[1889]), .Z(n5668) );
XNOR U9448 ( .A(b[1889]), .B(n5669), .Z(c[1889]) );
XNOR U9449 ( .A(a[1889]), .B(c1889), .Z(n5669) );
XOR U9450 ( .A(c1890), .B(n5670), .Z(c1891) );
ANDN U9451 ( .B(n5671), .A(n5672), .Z(n5670) );
XOR U9452 ( .A(c1890), .B(b[1890]), .Z(n5671) );
XNOR U9453 ( .A(b[1890]), .B(n5672), .Z(c[1890]) );
XNOR U9454 ( .A(a[1890]), .B(c1890), .Z(n5672) );
XOR U9455 ( .A(c1891), .B(n5673), .Z(c1892) );
ANDN U9456 ( .B(n5674), .A(n5675), .Z(n5673) );
XOR U9457 ( .A(c1891), .B(b[1891]), .Z(n5674) );
XNOR U9458 ( .A(b[1891]), .B(n5675), .Z(c[1891]) );
XNOR U9459 ( .A(a[1891]), .B(c1891), .Z(n5675) );
XOR U9460 ( .A(c1892), .B(n5676), .Z(c1893) );
ANDN U9461 ( .B(n5677), .A(n5678), .Z(n5676) );
XOR U9462 ( .A(c1892), .B(b[1892]), .Z(n5677) );
XNOR U9463 ( .A(b[1892]), .B(n5678), .Z(c[1892]) );
XNOR U9464 ( .A(a[1892]), .B(c1892), .Z(n5678) );
XOR U9465 ( .A(c1893), .B(n5679), .Z(c1894) );
ANDN U9466 ( .B(n5680), .A(n5681), .Z(n5679) );
XOR U9467 ( .A(c1893), .B(b[1893]), .Z(n5680) );
XNOR U9468 ( .A(b[1893]), .B(n5681), .Z(c[1893]) );
XNOR U9469 ( .A(a[1893]), .B(c1893), .Z(n5681) );
XOR U9470 ( .A(c1894), .B(n5682), .Z(c1895) );
ANDN U9471 ( .B(n5683), .A(n5684), .Z(n5682) );
XOR U9472 ( .A(c1894), .B(b[1894]), .Z(n5683) );
XNOR U9473 ( .A(b[1894]), .B(n5684), .Z(c[1894]) );
XNOR U9474 ( .A(a[1894]), .B(c1894), .Z(n5684) );
XOR U9475 ( .A(c1895), .B(n5685), .Z(c1896) );
ANDN U9476 ( .B(n5686), .A(n5687), .Z(n5685) );
XOR U9477 ( .A(c1895), .B(b[1895]), .Z(n5686) );
XNOR U9478 ( .A(b[1895]), .B(n5687), .Z(c[1895]) );
XNOR U9479 ( .A(a[1895]), .B(c1895), .Z(n5687) );
XOR U9480 ( .A(c1896), .B(n5688), .Z(c1897) );
ANDN U9481 ( .B(n5689), .A(n5690), .Z(n5688) );
XOR U9482 ( .A(c1896), .B(b[1896]), .Z(n5689) );
XNOR U9483 ( .A(b[1896]), .B(n5690), .Z(c[1896]) );
XNOR U9484 ( .A(a[1896]), .B(c1896), .Z(n5690) );
XOR U9485 ( .A(c1897), .B(n5691), .Z(c1898) );
ANDN U9486 ( .B(n5692), .A(n5693), .Z(n5691) );
XOR U9487 ( .A(c1897), .B(b[1897]), .Z(n5692) );
XNOR U9488 ( .A(b[1897]), .B(n5693), .Z(c[1897]) );
XNOR U9489 ( .A(a[1897]), .B(c1897), .Z(n5693) );
XOR U9490 ( .A(c1898), .B(n5694), .Z(c1899) );
ANDN U9491 ( .B(n5695), .A(n5696), .Z(n5694) );
XOR U9492 ( .A(c1898), .B(b[1898]), .Z(n5695) );
XNOR U9493 ( .A(b[1898]), .B(n5696), .Z(c[1898]) );
XNOR U9494 ( .A(a[1898]), .B(c1898), .Z(n5696) );
XOR U9495 ( .A(c1899), .B(n5697), .Z(c1900) );
ANDN U9496 ( .B(n5698), .A(n5699), .Z(n5697) );
XOR U9497 ( .A(c1899), .B(b[1899]), .Z(n5698) );
XNOR U9498 ( .A(b[1899]), .B(n5699), .Z(c[1899]) );
XNOR U9499 ( .A(a[1899]), .B(c1899), .Z(n5699) );
XOR U9500 ( .A(c1900), .B(n5700), .Z(c1901) );
ANDN U9501 ( .B(n5701), .A(n5702), .Z(n5700) );
XOR U9502 ( .A(c1900), .B(b[1900]), .Z(n5701) );
XNOR U9503 ( .A(b[1900]), .B(n5702), .Z(c[1900]) );
XNOR U9504 ( .A(a[1900]), .B(c1900), .Z(n5702) );
XOR U9505 ( .A(c1901), .B(n5703), .Z(c1902) );
ANDN U9506 ( .B(n5704), .A(n5705), .Z(n5703) );
XOR U9507 ( .A(c1901), .B(b[1901]), .Z(n5704) );
XNOR U9508 ( .A(b[1901]), .B(n5705), .Z(c[1901]) );
XNOR U9509 ( .A(a[1901]), .B(c1901), .Z(n5705) );
XOR U9510 ( .A(c1902), .B(n5706), .Z(c1903) );
ANDN U9511 ( .B(n5707), .A(n5708), .Z(n5706) );
XOR U9512 ( .A(c1902), .B(b[1902]), .Z(n5707) );
XNOR U9513 ( .A(b[1902]), .B(n5708), .Z(c[1902]) );
XNOR U9514 ( .A(a[1902]), .B(c1902), .Z(n5708) );
XOR U9515 ( .A(c1903), .B(n5709), .Z(c1904) );
ANDN U9516 ( .B(n5710), .A(n5711), .Z(n5709) );
XOR U9517 ( .A(c1903), .B(b[1903]), .Z(n5710) );
XNOR U9518 ( .A(b[1903]), .B(n5711), .Z(c[1903]) );
XNOR U9519 ( .A(a[1903]), .B(c1903), .Z(n5711) );
XOR U9520 ( .A(c1904), .B(n5712), .Z(c1905) );
ANDN U9521 ( .B(n5713), .A(n5714), .Z(n5712) );
XOR U9522 ( .A(c1904), .B(b[1904]), .Z(n5713) );
XNOR U9523 ( .A(b[1904]), .B(n5714), .Z(c[1904]) );
XNOR U9524 ( .A(a[1904]), .B(c1904), .Z(n5714) );
XOR U9525 ( .A(c1905), .B(n5715), .Z(c1906) );
ANDN U9526 ( .B(n5716), .A(n5717), .Z(n5715) );
XOR U9527 ( .A(c1905), .B(b[1905]), .Z(n5716) );
XNOR U9528 ( .A(b[1905]), .B(n5717), .Z(c[1905]) );
XNOR U9529 ( .A(a[1905]), .B(c1905), .Z(n5717) );
XOR U9530 ( .A(c1906), .B(n5718), .Z(c1907) );
ANDN U9531 ( .B(n5719), .A(n5720), .Z(n5718) );
XOR U9532 ( .A(c1906), .B(b[1906]), .Z(n5719) );
XNOR U9533 ( .A(b[1906]), .B(n5720), .Z(c[1906]) );
XNOR U9534 ( .A(a[1906]), .B(c1906), .Z(n5720) );
XOR U9535 ( .A(c1907), .B(n5721), .Z(c1908) );
ANDN U9536 ( .B(n5722), .A(n5723), .Z(n5721) );
XOR U9537 ( .A(c1907), .B(b[1907]), .Z(n5722) );
XNOR U9538 ( .A(b[1907]), .B(n5723), .Z(c[1907]) );
XNOR U9539 ( .A(a[1907]), .B(c1907), .Z(n5723) );
XOR U9540 ( .A(c1908), .B(n5724), .Z(c1909) );
ANDN U9541 ( .B(n5725), .A(n5726), .Z(n5724) );
XOR U9542 ( .A(c1908), .B(b[1908]), .Z(n5725) );
XNOR U9543 ( .A(b[1908]), .B(n5726), .Z(c[1908]) );
XNOR U9544 ( .A(a[1908]), .B(c1908), .Z(n5726) );
XOR U9545 ( .A(c1909), .B(n5727), .Z(c1910) );
ANDN U9546 ( .B(n5728), .A(n5729), .Z(n5727) );
XOR U9547 ( .A(c1909), .B(b[1909]), .Z(n5728) );
XNOR U9548 ( .A(b[1909]), .B(n5729), .Z(c[1909]) );
XNOR U9549 ( .A(a[1909]), .B(c1909), .Z(n5729) );
XOR U9550 ( .A(c1910), .B(n5730), .Z(c1911) );
ANDN U9551 ( .B(n5731), .A(n5732), .Z(n5730) );
XOR U9552 ( .A(c1910), .B(b[1910]), .Z(n5731) );
XNOR U9553 ( .A(b[1910]), .B(n5732), .Z(c[1910]) );
XNOR U9554 ( .A(a[1910]), .B(c1910), .Z(n5732) );
XOR U9555 ( .A(c1911), .B(n5733), .Z(c1912) );
ANDN U9556 ( .B(n5734), .A(n5735), .Z(n5733) );
XOR U9557 ( .A(c1911), .B(b[1911]), .Z(n5734) );
XNOR U9558 ( .A(b[1911]), .B(n5735), .Z(c[1911]) );
XNOR U9559 ( .A(a[1911]), .B(c1911), .Z(n5735) );
XOR U9560 ( .A(c1912), .B(n5736), .Z(c1913) );
ANDN U9561 ( .B(n5737), .A(n5738), .Z(n5736) );
XOR U9562 ( .A(c1912), .B(b[1912]), .Z(n5737) );
XNOR U9563 ( .A(b[1912]), .B(n5738), .Z(c[1912]) );
XNOR U9564 ( .A(a[1912]), .B(c1912), .Z(n5738) );
XOR U9565 ( .A(c1913), .B(n5739), .Z(c1914) );
ANDN U9566 ( .B(n5740), .A(n5741), .Z(n5739) );
XOR U9567 ( .A(c1913), .B(b[1913]), .Z(n5740) );
XNOR U9568 ( .A(b[1913]), .B(n5741), .Z(c[1913]) );
XNOR U9569 ( .A(a[1913]), .B(c1913), .Z(n5741) );
XOR U9570 ( .A(c1914), .B(n5742), .Z(c1915) );
ANDN U9571 ( .B(n5743), .A(n5744), .Z(n5742) );
XOR U9572 ( .A(c1914), .B(b[1914]), .Z(n5743) );
XNOR U9573 ( .A(b[1914]), .B(n5744), .Z(c[1914]) );
XNOR U9574 ( .A(a[1914]), .B(c1914), .Z(n5744) );
XOR U9575 ( .A(c1915), .B(n5745), .Z(c1916) );
ANDN U9576 ( .B(n5746), .A(n5747), .Z(n5745) );
XOR U9577 ( .A(c1915), .B(b[1915]), .Z(n5746) );
XNOR U9578 ( .A(b[1915]), .B(n5747), .Z(c[1915]) );
XNOR U9579 ( .A(a[1915]), .B(c1915), .Z(n5747) );
XOR U9580 ( .A(c1916), .B(n5748), .Z(c1917) );
ANDN U9581 ( .B(n5749), .A(n5750), .Z(n5748) );
XOR U9582 ( .A(c1916), .B(b[1916]), .Z(n5749) );
XNOR U9583 ( .A(b[1916]), .B(n5750), .Z(c[1916]) );
XNOR U9584 ( .A(a[1916]), .B(c1916), .Z(n5750) );
XOR U9585 ( .A(c1917), .B(n5751), .Z(c1918) );
ANDN U9586 ( .B(n5752), .A(n5753), .Z(n5751) );
XOR U9587 ( .A(c1917), .B(b[1917]), .Z(n5752) );
XNOR U9588 ( .A(b[1917]), .B(n5753), .Z(c[1917]) );
XNOR U9589 ( .A(a[1917]), .B(c1917), .Z(n5753) );
XOR U9590 ( .A(c1918), .B(n5754), .Z(c1919) );
ANDN U9591 ( .B(n5755), .A(n5756), .Z(n5754) );
XOR U9592 ( .A(c1918), .B(b[1918]), .Z(n5755) );
XNOR U9593 ( .A(b[1918]), .B(n5756), .Z(c[1918]) );
XNOR U9594 ( .A(a[1918]), .B(c1918), .Z(n5756) );
XOR U9595 ( .A(c1919), .B(n5757), .Z(c1920) );
ANDN U9596 ( .B(n5758), .A(n5759), .Z(n5757) );
XOR U9597 ( .A(c1919), .B(b[1919]), .Z(n5758) );
XNOR U9598 ( .A(b[1919]), .B(n5759), .Z(c[1919]) );
XNOR U9599 ( .A(a[1919]), .B(c1919), .Z(n5759) );
XOR U9600 ( .A(c1920), .B(n5760), .Z(c1921) );
ANDN U9601 ( .B(n5761), .A(n5762), .Z(n5760) );
XOR U9602 ( .A(c1920), .B(b[1920]), .Z(n5761) );
XNOR U9603 ( .A(b[1920]), .B(n5762), .Z(c[1920]) );
XNOR U9604 ( .A(a[1920]), .B(c1920), .Z(n5762) );
XOR U9605 ( .A(c1921), .B(n5763), .Z(c1922) );
ANDN U9606 ( .B(n5764), .A(n5765), .Z(n5763) );
XOR U9607 ( .A(c1921), .B(b[1921]), .Z(n5764) );
XNOR U9608 ( .A(b[1921]), .B(n5765), .Z(c[1921]) );
XNOR U9609 ( .A(a[1921]), .B(c1921), .Z(n5765) );
XOR U9610 ( .A(c1922), .B(n5766), .Z(c1923) );
ANDN U9611 ( .B(n5767), .A(n5768), .Z(n5766) );
XOR U9612 ( .A(c1922), .B(b[1922]), .Z(n5767) );
XNOR U9613 ( .A(b[1922]), .B(n5768), .Z(c[1922]) );
XNOR U9614 ( .A(a[1922]), .B(c1922), .Z(n5768) );
XOR U9615 ( .A(c1923), .B(n5769), .Z(c1924) );
ANDN U9616 ( .B(n5770), .A(n5771), .Z(n5769) );
XOR U9617 ( .A(c1923), .B(b[1923]), .Z(n5770) );
XNOR U9618 ( .A(b[1923]), .B(n5771), .Z(c[1923]) );
XNOR U9619 ( .A(a[1923]), .B(c1923), .Z(n5771) );
XOR U9620 ( .A(c1924), .B(n5772), .Z(c1925) );
ANDN U9621 ( .B(n5773), .A(n5774), .Z(n5772) );
XOR U9622 ( .A(c1924), .B(b[1924]), .Z(n5773) );
XNOR U9623 ( .A(b[1924]), .B(n5774), .Z(c[1924]) );
XNOR U9624 ( .A(a[1924]), .B(c1924), .Z(n5774) );
XOR U9625 ( .A(c1925), .B(n5775), .Z(c1926) );
ANDN U9626 ( .B(n5776), .A(n5777), .Z(n5775) );
XOR U9627 ( .A(c1925), .B(b[1925]), .Z(n5776) );
XNOR U9628 ( .A(b[1925]), .B(n5777), .Z(c[1925]) );
XNOR U9629 ( .A(a[1925]), .B(c1925), .Z(n5777) );
XOR U9630 ( .A(c1926), .B(n5778), .Z(c1927) );
ANDN U9631 ( .B(n5779), .A(n5780), .Z(n5778) );
XOR U9632 ( .A(c1926), .B(b[1926]), .Z(n5779) );
XNOR U9633 ( .A(b[1926]), .B(n5780), .Z(c[1926]) );
XNOR U9634 ( .A(a[1926]), .B(c1926), .Z(n5780) );
XOR U9635 ( .A(c1927), .B(n5781), .Z(c1928) );
ANDN U9636 ( .B(n5782), .A(n5783), .Z(n5781) );
XOR U9637 ( .A(c1927), .B(b[1927]), .Z(n5782) );
XNOR U9638 ( .A(b[1927]), .B(n5783), .Z(c[1927]) );
XNOR U9639 ( .A(a[1927]), .B(c1927), .Z(n5783) );
XOR U9640 ( .A(c1928), .B(n5784), .Z(c1929) );
ANDN U9641 ( .B(n5785), .A(n5786), .Z(n5784) );
XOR U9642 ( .A(c1928), .B(b[1928]), .Z(n5785) );
XNOR U9643 ( .A(b[1928]), .B(n5786), .Z(c[1928]) );
XNOR U9644 ( .A(a[1928]), .B(c1928), .Z(n5786) );
XOR U9645 ( .A(c1929), .B(n5787), .Z(c1930) );
ANDN U9646 ( .B(n5788), .A(n5789), .Z(n5787) );
XOR U9647 ( .A(c1929), .B(b[1929]), .Z(n5788) );
XNOR U9648 ( .A(b[1929]), .B(n5789), .Z(c[1929]) );
XNOR U9649 ( .A(a[1929]), .B(c1929), .Z(n5789) );
XOR U9650 ( .A(c1930), .B(n5790), .Z(c1931) );
ANDN U9651 ( .B(n5791), .A(n5792), .Z(n5790) );
XOR U9652 ( .A(c1930), .B(b[1930]), .Z(n5791) );
XNOR U9653 ( .A(b[1930]), .B(n5792), .Z(c[1930]) );
XNOR U9654 ( .A(a[1930]), .B(c1930), .Z(n5792) );
XOR U9655 ( .A(c1931), .B(n5793), .Z(c1932) );
ANDN U9656 ( .B(n5794), .A(n5795), .Z(n5793) );
XOR U9657 ( .A(c1931), .B(b[1931]), .Z(n5794) );
XNOR U9658 ( .A(b[1931]), .B(n5795), .Z(c[1931]) );
XNOR U9659 ( .A(a[1931]), .B(c1931), .Z(n5795) );
XOR U9660 ( .A(c1932), .B(n5796), .Z(c1933) );
ANDN U9661 ( .B(n5797), .A(n5798), .Z(n5796) );
XOR U9662 ( .A(c1932), .B(b[1932]), .Z(n5797) );
XNOR U9663 ( .A(b[1932]), .B(n5798), .Z(c[1932]) );
XNOR U9664 ( .A(a[1932]), .B(c1932), .Z(n5798) );
XOR U9665 ( .A(c1933), .B(n5799), .Z(c1934) );
ANDN U9666 ( .B(n5800), .A(n5801), .Z(n5799) );
XOR U9667 ( .A(c1933), .B(b[1933]), .Z(n5800) );
XNOR U9668 ( .A(b[1933]), .B(n5801), .Z(c[1933]) );
XNOR U9669 ( .A(a[1933]), .B(c1933), .Z(n5801) );
XOR U9670 ( .A(c1934), .B(n5802), .Z(c1935) );
ANDN U9671 ( .B(n5803), .A(n5804), .Z(n5802) );
XOR U9672 ( .A(c1934), .B(b[1934]), .Z(n5803) );
XNOR U9673 ( .A(b[1934]), .B(n5804), .Z(c[1934]) );
XNOR U9674 ( .A(a[1934]), .B(c1934), .Z(n5804) );
XOR U9675 ( .A(c1935), .B(n5805), .Z(c1936) );
ANDN U9676 ( .B(n5806), .A(n5807), .Z(n5805) );
XOR U9677 ( .A(c1935), .B(b[1935]), .Z(n5806) );
XNOR U9678 ( .A(b[1935]), .B(n5807), .Z(c[1935]) );
XNOR U9679 ( .A(a[1935]), .B(c1935), .Z(n5807) );
XOR U9680 ( .A(c1936), .B(n5808), .Z(c1937) );
ANDN U9681 ( .B(n5809), .A(n5810), .Z(n5808) );
XOR U9682 ( .A(c1936), .B(b[1936]), .Z(n5809) );
XNOR U9683 ( .A(b[1936]), .B(n5810), .Z(c[1936]) );
XNOR U9684 ( .A(a[1936]), .B(c1936), .Z(n5810) );
XOR U9685 ( .A(c1937), .B(n5811), .Z(c1938) );
ANDN U9686 ( .B(n5812), .A(n5813), .Z(n5811) );
XOR U9687 ( .A(c1937), .B(b[1937]), .Z(n5812) );
XNOR U9688 ( .A(b[1937]), .B(n5813), .Z(c[1937]) );
XNOR U9689 ( .A(a[1937]), .B(c1937), .Z(n5813) );
XOR U9690 ( .A(c1938), .B(n5814), .Z(c1939) );
ANDN U9691 ( .B(n5815), .A(n5816), .Z(n5814) );
XOR U9692 ( .A(c1938), .B(b[1938]), .Z(n5815) );
XNOR U9693 ( .A(b[1938]), .B(n5816), .Z(c[1938]) );
XNOR U9694 ( .A(a[1938]), .B(c1938), .Z(n5816) );
XOR U9695 ( .A(c1939), .B(n5817), .Z(c1940) );
ANDN U9696 ( .B(n5818), .A(n5819), .Z(n5817) );
XOR U9697 ( .A(c1939), .B(b[1939]), .Z(n5818) );
XNOR U9698 ( .A(b[1939]), .B(n5819), .Z(c[1939]) );
XNOR U9699 ( .A(a[1939]), .B(c1939), .Z(n5819) );
XOR U9700 ( .A(c1940), .B(n5820), .Z(c1941) );
ANDN U9701 ( .B(n5821), .A(n5822), .Z(n5820) );
XOR U9702 ( .A(c1940), .B(b[1940]), .Z(n5821) );
XNOR U9703 ( .A(b[1940]), .B(n5822), .Z(c[1940]) );
XNOR U9704 ( .A(a[1940]), .B(c1940), .Z(n5822) );
XOR U9705 ( .A(c1941), .B(n5823), .Z(c1942) );
ANDN U9706 ( .B(n5824), .A(n5825), .Z(n5823) );
XOR U9707 ( .A(c1941), .B(b[1941]), .Z(n5824) );
XNOR U9708 ( .A(b[1941]), .B(n5825), .Z(c[1941]) );
XNOR U9709 ( .A(a[1941]), .B(c1941), .Z(n5825) );
XOR U9710 ( .A(c1942), .B(n5826), .Z(c1943) );
ANDN U9711 ( .B(n5827), .A(n5828), .Z(n5826) );
XOR U9712 ( .A(c1942), .B(b[1942]), .Z(n5827) );
XNOR U9713 ( .A(b[1942]), .B(n5828), .Z(c[1942]) );
XNOR U9714 ( .A(a[1942]), .B(c1942), .Z(n5828) );
XOR U9715 ( .A(c1943), .B(n5829), .Z(c1944) );
ANDN U9716 ( .B(n5830), .A(n5831), .Z(n5829) );
XOR U9717 ( .A(c1943), .B(b[1943]), .Z(n5830) );
XNOR U9718 ( .A(b[1943]), .B(n5831), .Z(c[1943]) );
XNOR U9719 ( .A(a[1943]), .B(c1943), .Z(n5831) );
XOR U9720 ( .A(c1944), .B(n5832), .Z(c1945) );
ANDN U9721 ( .B(n5833), .A(n5834), .Z(n5832) );
XOR U9722 ( .A(c1944), .B(b[1944]), .Z(n5833) );
XNOR U9723 ( .A(b[1944]), .B(n5834), .Z(c[1944]) );
XNOR U9724 ( .A(a[1944]), .B(c1944), .Z(n5834) );
XOR U9725 ( .A(c1945), .B(n5835), .Z(c1946) );
ANDN U9726 ( .B(n5836), .A(n5837), .Z(n5835) );
XOR U9727 ( .A(c1945), .B(b[1945]), .Z(n5836) );
XNOR U9728 ( .A(b[1945]), .B(n5837), .Z(c[1945]) );
XNOR U9729 ( .A(a[1945]), .B(c1945), .Z(n5837) );
XOR U9730 ( .A(c1946), .B(n5838), .Z(c1947) );
ANDN U9731 ( .B(n5839), .A(n5840), .Z(n5838) );
XOR U9732 ( .A(c1946), .B(b[1946]), .Z(n5839) );
XNOR U9733 ( .A(b[1946]), .B(n5840), .Z(c[1946]) );
XNOR U9734 ( .A(a[1946]), .B(c1946), .Z(n5840) );
XOR U9735 ( .A(c1947), .B(n5841), .Z(c1948) );
ANDN U9736 ( .B(n5842), .A(n5843), .Z(n5841) );
XOR U9737 ( .A(c1947), .B(b[1947]), .Z(n5842) );
XNOR U9738 ( .A(b[1947]), .B(n5843), .Z(c[1947]) );
XNOR U9739 ( .A(a[1947]), .B(c1947), .Z(n5843) );
XOR U9740 ( .A(c1948), .B(n5844), .Z(c1949) );
ANDN U9741 ( .B(n5845), .A(n5846), .Z(n5844) );
XOR U9742 ( .A(c1948), .B(b[1948]), .Z(n5845) );
XNOR U9743 ( .A(b[1948]), .B(n5846), .Z(c[1948]) );
XNOR U9744 ( .A(a[1948]), .B(c1948), .Z(n5846) );
XOR U9745 ( .A(c1949), .B(n5847), .Z(c1950) );
ANDN U9746 ( .B(n5848), .A(n5849), .Z(n5847) );
XOR U9747 ( .A(c1949), .B(b[1949]), .Z(n5848) );
XNOR U9748 ( .A(b[1949]), .B(n5849), .Z(c[1949]) );
XNOR U9749 ( .A(a[1949]), .B(c1949), .Z(n5849) );
XOR U9750 ( .A(c1950), .B(n5850), .Z(c1951) );
ANDN U9751 ( .B(n5851), .A(n5852), .Z(n5850) );
XOR U9752 ( .A(c1950), .B(b[1950]), .Z(n5851) );
XNOR U9753 ( .A(b[1950]), .B(n5852), .Z(c[1950]) );
XNOR U9754 ( .A(a[1950]), .B(c1950), .Z(n5852) );
XOR U9755 ( .A(c1951), .B(n5853), .Z(c1952) );
ANDN U9756 ( .B(n5854), .A(n5855), .Z(n5853) );
XOR U9757 ( .A(c1951), .B(b[1951]), .Z(n5854) );
XNOR U9758 ( .A(b[1951]), .B(n5855), .Z(c[1951]) );
XNOR U9759 ( .A(a[1951]), .B(c1951), .Z(n5855) );
XOR U9760 ( .A(c1952), .B(n5856), .Z(c1953) );
ANDN U9761 ( .B(n5857), .A(n5858), .Z(n5856) );
XOR U9762 ( .A(c1952), .B(b[1952]), .Z(n5857) );
XNOR U9763 ( .A(b[1952]), .B(n5858), .Z(c[1952]) );
XNOR U9764 ( .A(a[1952]), .B(c1952), .Z(n5858) );
XOR U9765 ( .A(c1953), .B(n5859), .Z(c1954) );
ANDN U9766 ( .B(n5860), .A(n5861), .Z(n5859) );
XOR U9767 ( .A(c1953), .B(b[1953]), .Z(n5860) );
XNOR U9768 ( .A(b[1953]), .B(n5861), .Z(c[1953]) );
XNOR U9769 ( .A(a[1953]), .B(c1953), .Z(n5861) );
XOR U9770 ( .A(c1954), .B(n5862), .Z(c1955) );
ANDN U9771 ( .B(n5863), .A(n5864), .Z(n5862) );
XOR U9772 ( .A(c1954), .B(b[1954]), .Z(n5863) );
XNOR U9773 ( .A(b[1954]), .B(n5864), .Z(c[1954]) );
XNOR U9774 ( .A(a[1954]), .B(c1954), .Z(n5864) );
XOR U9775 ( .A(c1955), .B(n5865), .Z(c1956) );
ANDN U9776 ( .B(n5866), .A(n5867), .Z(n5865) );
XOR U9777 ( .A(c1955), .B(b[1955]), .Z(n5866) );
XNOR U9778 ( .A(b[1955]), .B(n5867), .Z(c[1955]) );
XNOR U9779 ( .A(a[1955]), .B(c1955), .Z(n5867) );
XOR U9780 ( .A(c1956), .B(n5868), .Z(c1957) );
ANDN U9781 ( .B(n5869), .A(n5870), .Z(n5868) );
XOR U9782 ( .A(c1956), .B(b[1956]), .Z(n5869) );
XNOR U9783 ( .A(b[1956]), .B(n5870), .Z(c[1956]) );
XNOR U9784 ( .A(a[1956]), .B(c1956), .Z(n5870) );
XOR U9785 ( .A(c1957), .B(n5871), .Z(c1958) );
ANDN U9786 ( .B(n5872), .A(n5873), .Z(n5871) );
XOR U9787 ( .A(c1957), .B(b[1957]), .Z(n5872) );
XNOR U9788 ( .A(b[1957]), .B(n5873), .Z(c[1957]) );
XNOR U9789 ( .A(a[1957]), .B(c1957), .Z(n5873) );
XOR U9790 ( .A(c1958), .B(n5874), .Z(c1959) );
ANDN U9791 ( .B(n5875), .A(n5876), .Z(n5874) );
XOR U9792 ( .A(c1958), .B(b[1958]), .Z(n5875) );
XNOR U9793 ( .A(b[1958]), .B(n5876), .Z(c[1958]) );
XNOR U9794 ( .A(a[1958]), .B(c1958), .Z(n5876) );
XOR U9795 ( .A(c1959), .B(n5877), .Z(c1960) );
ANDN U9796 ( .B(n5878), .A(n5879), .Z(n5877) );
XOR U9797 ( .A(c1959), .B(b[1959]), .Z(n5878) );
XNOR U9798 ( .A(b[1959]), .B(n5879), .Z(c[1959]) );
XNOR U9799 ( .A(a[1959]), .B(c1959), .Z(n5879) );
XOR U9800 ( .A(c1960), .B(n5880), .Z(c1961) );
ANDN U9801 ( .B(n5881), .A(n5882), .Z(n5880) );
XOR U9802 ( .A(c1960), .B(b[1960]), .Z(n5881) );
XNOR U9803 ( .A(b[1960]), .B(n5882), .Z(c[1960]) );
XNOR U9804 ( .A(a[1960]), .B(c1960), .Z(n5882) );
XOR U9805 ( .A(c1961), .B(n5883), .Z(c1962) );
ANDN U9806 ( .B(n5884), .A(n5885), .Z(n5883) );
XOR U9807 ( .A(c1961), .B(b[1961]), .Z(n5884) );
XNOR U9808 ( .A(b[1961]), .B(n5885), .Z(c[1961]) );
XNOR U9809 ( .A(a[1961]), .B(c1961), .Z(n5885) );
XOR U9810 ( .A(c1962), .B(n5886), .Z(c1963) );
ANDN U9811 ( .B(n5887), .A(n5888), .Z(n5886) );
XOR U9812 ( .A(c1962), .B(b[1962]), .Z(n5887) );
XNOR U9813 ( .A(b[1962]), .B(n5888), .Z(c[1962]) );
XNOR U9814 ( .A(a[1962]), .B(c1962), .Z(n5888) );
XOR U9815 ( .A(c1963), .B(n5889), .Z(c1964) );
ANDN U9816 ( .B(n5890), .A(n5891), .Z(n5889) );
XOR U9817 ( .A(c1963), .B(b[1963]), .Z(n5890) );
XNOR U9818 ( .A(b[1963]), .B(n5891), .Z(c[1963]) );
XNOR U9819 ( .A(a[1963]), .B(c1963), .Z(n5891) );
XOR U9820 ( .A(c1964), .B(n5892), .Z(c1965) );
ANDN U9821 ( .B(n5893), .A(n5894), .Z(n5892) );
XOR U9822 ( .A(c1964), .B(b[1964]), .Z(n5893) );
XNOR U9823 ( .A(b[1964]), .B(n5894), .Z(c[1964]) );
XNOR U9824 ( .A(a[1964]), .B(c1964), .Z(n5894) );
XOR U9825 ( .A(c1965), .B(n5895), .Z(c1966) );
ANDN U9826 ( .B(n5896), .A(n5897), .Z(n5895) );
XOR U9827 ( .A(c1965), .B(b[1965]), .Z(n5896) );
XNOR U9828 ( .A(b[1965]), .B(n5897), .Z(c[1965]) );
XNOR U9829 ( .A(a[1965]), .B(c1965), .Z(n5897) );
XOR U9830 ( .A(c1966), .B(n5898), .Z(c1967) );
ANDN U9831 ( .B(n5899), .A(n5900), .Z(n5898) );
XOR U9832 ( .A(c1966), .B(b[1966]), .Z(n5899) );
XNOR U9833 ( .A(b[1966]), .B(n5900), .Z(c[1966]) );
XNOR U9834 ( .A(a[1966]), .B(c1966), .Z(n5900) );
XOR U9835 ( .A(c1967), .B(n5901), .Z(c1968) );
ANDN U9836 ( .B(n5902), .A(n5903), .Z(n5901) );
XOR U9837 ( .A(c1967), .B(b[1967]), .Z(n5902) );
XNOR U9838 ( .A(b[1967]), .B(n5903), .Z(c[1967]) );
XNOR U9839 ( .A(a[1967]), .B(c1967), .Z(n5903) );
XOR U9840 ( .A(c1968), .B(n5904), .Z(c1969) );
ANDN U9841 ( .B(n5905), .A(n5906), .Z(n5904) );
XOR U9842 ( .A(c1968), .B(b[1968]), .Z(n5905) );
XNOR U9843 ( .A(b[1968]), .B(n5906), .Z(c[1968]) );
XNOR U9844 ( .A(a[1968]), .B(c1968), .Z(n5906) );
XOR U9845 ( .A(c1969), .B(n5907), .Z(c1970) );
ANDN U9846 ( .B(n5908), .A(n5909), .Z(n5907) );
XOR U9847 ( .A(c1969), .B(b[1969]), .Z(n5908) );
XNOR U9848 ( .A(b[1969]), .B(n5909), .Z(c[1969]) );
XNOR U9849 ( .A(a[1969]), .B(c1969), .Z(n5909) );
XOR U9850 ( .A(c1970), .B(n5910), .Z(c1971) );
ANDN U9851 ( .B(n5911), .A(n5912), .Z(n5910) );
XOR U9852 ( .A(c1970), .B(b[1970]), .Z(n5911) );
XNOR U9853 ( .A(b[1970]), .B(n5912), .Z(c[1970]) );
XNOR U9854 ( .A(a[1970]), .B(c1970), .Z(n5912) );
XOR U9855 ( .A(c1971), .B(n5913), .Z(c1972) );
ANDN U9856 ( .B(n5914), .A(n5915), .Z(n5913) );
XOR U9857 ( .A(c1971), .B(b[1971]), .Z(n5914) );
XNOR U9858 ( .A(b[1971]), .B(n5915), .Z(c[1971]) );
XNOR U9859 ( .A(a[1971]), .B(c1971), .Z(n5915) );
XOR U9860 ( .A(c1972), .B(n5916), .Z(c1973) );
ANDN U9861 ( .B(n5917), .A(n5918), .Z(n5916) );
XOR U9862 ( .A(c1972), .B(b[1972]), .Z(n5917) );
XNOR U9863 ( .A(b[1972]), .B(n5918), .Z(c[1972]) );
XNOR U9864 ( .A(a[1972]), .B(c1972), .Z(n5918) );
XOR U9865 ( .A(c1973), .B(n5919), .Z(c1974) );
ANDN U9866 ( .B(n5920), .A(n5921), .Z(n5919) );
XOR U9867 ( .A(c1973), .B(b[1973]), .Z(n5920) );
XNOR U9868 ( .A(b[1973]), .B(n5921), .Z(c[1973]) );
XNOR U9869 ( .A(a[1973]), .B(c1973), .Z(n5921) );
XOR U9870 ( .A(c1974), .B(n5922), .Z(c1975) );
ANDN U9871 ( .B(n5923), .A(n5924), .Z(n5922) );
XOR U9872 ( .A(c1974), .B(b[1974]), .Z(n5923) );
XNOR U9873 ( .A(b[1974]), .B(n5924), .Z(c[1974]) );
XNOR U9874 ( .A(a[1974]), .B(c1974), .Z(n5924) );
XOR U9875 ( .A(c1975), .B(n5925), .Z(c1976) );
ANDN U9876 ( .B(n5926), .A(n5927), .Z(n5925) );
XOR U9877 ( .A(c1975), .B(b[1975]), .Z(n5926) );
XNOR U9878 ( .A(b[1975]), .B(n5927), .Z(c[1975]) );
XNOR U9879 ( .A(a[1975]), .B(c1975), .Z(n5927) );
XOR U9880 ( .A(c1976), .B(n5928), .Z(c1977) );
ANDN U9881 ( .B(n5929), .A(n5930), .Z(n5928) );
XOR U9882 ( .A(c1976), .B(b[1976]), .Z(n5929) );
XNOR U9883 ( .A(b[1976]), .B(n5930), .Z(c[1976]) );
XNOR U9884 ( .A(a[1976]), .B(c1976), .Z(n5930) );
XOR U9885 ( .A(c1977), .B(n5931), .Z(c1978) );
ANDN U9886 ( .B(n5932), .A(n5933), .Z(n5931) );
XOR U9887 ( .A(c1977), .B(b[1977]), .Z(n5932) );
XNOR U9888 ( .A(b[1977]), .B(n5933), .Z(c[1977]) );
XNOR U9889 ( .A(a[1977]), .B(c1977), .Z(n5933) );
XOR U9890 ( .A(c1978), .B(n5934), .Z(c1979) );
ANDN U9891 ( .B(n5935), .A(n5936), .Z(n5934) );
XOR U9892 ( .A(c1978), .B(b[1978]), .Z(n5935) );
XNOR U9893 ( .A(b[1978]), .B(n5936), .Z(c[1978]) );
XNOR U9894 ( .A(a[1978]), .B(c1978), .Z(n5936) );
XOR U9895 ( .A(c1979), .B(n5937), .Z(c1980) );
ANDN U9896 ( .B(n5938), .A(n5939), .Z(n5937) );
XOR U9897 ( .A(c1979), .B(b[1979]), .Z(n5938) );
XNOR U9898 ( .A(b[1979]), .B(n5939), .Z(c[1979]) );
XNOR U9899 ( .A(a[1979]), .B(c1979), .Z(n5939) );
XOR U9900 ( .A(c1980), .B(n5940), .Z(c1981) );
ANDN U9901 ( .B(n5941), .A(n5942), .Z(n5940) );
XOR U9902 ( .A(c1980), .B(b[1980]), .Z(n5941) );
XNOR U9903 ( .A(b[1980]), .B(n5942), .Z(c[1980]) );
XNOR U9904 ( .A(a[1980]), .B(c1980), .Z(n5942) );
XOR U9905 ( .A(c1981), .B(n5943), .Z(c1982) );
ANDN U9906 ( .B(n5944), .A(n5945), .Z(n5943) );
XOR U9907 ( .A(c1981), .B(b[1981]), .Z(n5944) );
XNOR U9908 ( .A(b[1981]), .B(n5945), .Z(c[1981]) );
XNOR U9909 ( .A(a[1981]), .B(c1981), .Z(n5945) );
XOR U9910 ( .A(c1982), .B(n5946), .Z(c1983) );
ANDN U9911 ( .B(n5947), .A(n5948), .Z(n5946) );
XOR U9912 ( .A(c1982), .B(b[1982]), .Z(n5947) );
XNOR U9913 ( .A(b[1982]), .B(n5948), .Z(c[1982]) );
XNOR U9914 ( .A(a[1982]), .B(c1982), .Z(n5948) );
XOR U9915 ( .A(c1983), .B(n5949), .Z(c1984) );
ANDN U9916 ( .B(n5950), .A(n5951), .Z(n5949) );
XOR U9917 ( .A(c1983), .B(b[1983]), .Z(n5950) );
XNOR U9918 ( .A(b[1983]), .B(n5951), .Z(c[1983]) );
XNOR U9919 ( .A(a[1983]), .B(c1983), .Z(n5951) );
XOR U9920 ( .A(c1984), .B(n5952), .Z(c1985) );
ANDN U9921 ( .B(n5953), .A(n5954), .Z(n5952) );
XOR U9922 ( .A(c1984), .B(b[1984]), .Z(n5953) );
XNOR U9923 ( .A(b[1984]), .B(n5954), .Z(c[1984]) );
XNOR U9924 ( .A(a[1984]), .B(c1984), .Z(n5954) );
XOR U9925 ( .A(c1985), .B(n5955), .Z(c1986) );
ANDN U9926 ( .B(n5956), .A(n5957), .Z(n5955) );
XOR U9927 ( .A(c1985), .B(b[1985]), .Z(n5956) );
XNOR U9928 ( .A(b[1985]), .B(n5957), .Z(c[1985]) );
XNOR U9929 ( .A(a[1985]), .B(c1985), .Z(n5957) );
XOR U9930 ( .A(c1986), .B(n5958), .Z(c1987) );
ANDN U9931 ( .B(n5959), .A(n5960), .Z(n5958) );
XOR U9932 ( .A(c1986), .B(b[1986]), .Z(n5959) );
XNOR U9933 ( .A(b[1986]), .B(n5960), .Z(c[1986]) );
XNOR U9934 ( .A(a[1986]), .B(c1986), .Z(n5960) );
XOR U9935 ( .A(c1987), .B(n5961), .Z(c1988) );
ANDN U9936 ( .B(n5962), .A(n5963), .Z(n5961) );
XOR U9937 ( .A(c1987), .B(b[1987]), .Z(n5962) );
XNOR U9938 ( .A(b[1987]), .B(n5963), .Z(c[1987]) );
XNOR U9939 ( .A(a[1987]), .B(c1987), .Z(n5963) );
XOR U9940 ( .A(c1988), .B(n5964), .Z(c1989) );
ANDN U9941 ( .B(n5965), .A(n5966), .Z(n5964) );
XOR U9942 ( .A(c1988), .B(b[1988]), .Z(n5965) );
XNOR U9943 ( .A(b[1988]), .B(n5966), .Z(c[1988]) );
XNOR U9944 ( .A(a[1988]), .B(c1988), .Z(n5966) );
XOR U9945 ( .A(c1989), .B(n5967), .Z(c1990) );
ANDN U9946 ( .B(n5968), .A(n5969), .Z(n5967) );
XOR U9947 ( .A(c1989), .B(b[1989]), .Z(n5968) );
XNOR U9948 ( .A(b[1989]), .B(n5969), .Z(c[1989]) );
XNOR U9949 ( .A(a[1989]), .B(c1989), .Z(n5969) );
XOR U9950 ( .A(c1990), .B(n5970), .Z(c1991) );
ANDN U9951 ( .B(n5971), .A(n5972), .Z(n5970) );
XOR U9952 ( .A(c1990), .B(b[1990]), .Z(n5971) );
XNOR U9953 ( .A(b[1990]), .B(n5972), .Z(c[1990]) );
XNOR U9954 ( .A(a[1990]), .B(c1990), .Z(n5972) );
XOR U9955 ( .A(c1991), .B(n5973), .Z(c1992) );
ANDN U9956 ( .B(n5974), .A(n5975), .Z(n5973) );
XOR U9957 ( .A(c1991), .B(b[1991]), .Z(n5974) );
XNOR U9958 ( .A(b[1991]), .B(n5975), .Z(c[1991]) );
XNOR U9959 ( .A(a[1991]), .B(c1991), .Z(n5975) );
XOR U9960 ( .A(c1992), .B(n5976), .Z(c1993) );
ANDN U9961 ( .B(n5977), .A(n5978), .Z(n5976) );
XOR U9962 ( .A(c1992), .B(b[1992]), .Z(n5977) );
XNOR U9963 ( .A(b[1992]), .B(n5978), .Z(c[1992]) );
XNOR U9964 ( .A(a[1992]), .B(c1992), .Z(n5978) );
XOR U9965 ( .A(c1993), .B(n5979), .Z(c1994) );
ANDN U9966 ( .B(n5980), .A(n5981), .Z(n5979) );
XOR U9967 ( .A(c1993), .B(b[1993]), .Z(n5980) );
XNOR U9968 ( .A(b[1993]), .B(n5981), .Z(c[1993]) );
XNOR U9969 ( .A(a[1993]), .B(c1993), .Z(n5981) );
XOR U9970 ( .A(c1994), .B(n5982), .Z(c1995) );
ANDN U9971 ( .B(n5983), .A(n5984), .Z(n5982) );
XOR U9972 ( .A(c1994), .B(b[1994]), .Z(n5983) );
XNOR U9973 ( .A(b[1994]), .B(n5984), .Z(c[1994]) );
XNOR U9974 ( .A(a[1994]), .B(c1994), .Z(n5984) );
XOR U9975 ( .A(c1995), .B(n5985), .Z(c1996) );
ANDN U9976 ( .B(n5986), .A(n5987), .Z(n5985) );
XOR U9977 ( .A(c1995), .B(b[1995]), .Z(n5986) );
XNOR U9978 ( .A(b[1995]), .B(n5987), .Z(c[1995]) );
XNOR U9979 ( .A(a[1995]), .B(c1995), .Z(n5987) );
XOR U9980 ( .A(c1996), .B(n5988), .Z(c1997) );
ANDN U9981 ( .B(n5989), .A(n5990), .Z(n5988) );
XOR U9982 ( .A(c1996), .B(b[1996]), .Z(n5989) );
XNOR U9983 ( .A(b[1996]), .B(n5990), .Z(c[1996]) );
XNOR U9984 ( .A(a[1996]), .B(c1996), .Z(n5990) );
XOR U9985 ( .A(c1997), .B(n5991), .Z(c1998) );
ANDN U9986 ( .B(n5992), .A(n5993), .Z(n5991) );
XOR U9987 ( .A(c1997), .B(b[1997]), .Z(n5992) );
XNOR U9988 ( .A(b[1997]), .B(n5993), .Z(c[1997]) );
XNOR U9989 ( .A(a[1997]), .B(c1997), .Z(n5993) );
XOR U9990 ( .A(c1998), .B(n5994), .Z(c1999) );
ANDN U9991 ( .B(n5995), .A(n5996), .Z(n5994) );
XOR U9992 ( .A(c1998), .B(b[1998]), .Z(n5995) );
XNOR U9993 ( .A(b[1998]), .B(n5996), .Z(c[1998]) );
XNOR U9994 ( .A(a[1998]), .B(c1998), .Z(n5996) );
XOR U9995 ( .A(c1999), .B(n5997), .Z(c2000) );
ANDN U9996 ( .B(n5998), .A(n5999), .Z(n5997) );
XOR U9997 ( .A(c1999), .B(b[1999]), .Z(n5998) );
XNOR U9998 ( .A(b[1999]), .B(n5999), .Z(c[1999]) );
XNOR U9999 ( .A(a[1999]), .B(c1999), .Z(n5999) );
XOR U10000 ( .A(c2000), .B(n6000), .Z(c2001) );
ANDN U10001 ( .B(n6001), .A(n6002), .Z(n6000) );
XOR U10002 ( .A(c2000), .B(b[2000]), .Z(n6001) );
XNOR U10003 ( .A(b[2000]), .B(n6002), .Z(c[2000]) );
XNOR U10004 ( .A(a[2000]), .B(c2000), .Z(n6002) );
XOR U10005 ( .A(c2001), .B(n6003), .Z(c2002) );
ANDN U10006 ( .B(n6004), .A(n6005), .Z(n6003) );
XOR U10007 ( .A(c2001), .B(b[2001]), .Z(n6004) );
XNOR U10008 ( .A(b[2001]), .B(n6005), .Z(c[2001]) );
XNOR U10009 ( .A(a[2001]), .B(c2001), .Z(n6005) );
XOR U10010 ( .A(c2002), .B(n6006), .Z(c2003) );
ANDN U10011 ( .B(n6007), .A(n6008), .Z(n6006) );
XOR U10012 ( .A(c2002), .B(b[2002]), .Z(n6007) );
XNOR U10013 ( .A(b[2002]), .B(n6008), .Z(c[2002]) );
XNOR U10014 ( .A(a[2002]), .B(c2002), .Z(n6008) );
XOR U10015 ( .A(c2003), .B(n6009), .Z(c2004) );
ANDN U10016 ( .B(n6010), .A(n6011), .Z(n6009) );
XOR U10017 ( .A(c2003), .B(b[2003]), .Z(n6010) );
XNOR U10018 ( .A(b[2003]), .B(n6011), .Z(c[2003]) );
XNOR U10019 ( .A(a[2003]), .B(c2003), .Z(n6011) );
XOR U10020 ( .A(c2004), .B(n6012), .Z(c2005) );
ANDN U10021 ( .B(n6013), .A(n6014), .Z(n6012) );
XOR U10022 ( .A(c2004), .B(b[2004]), .Z(n6013) );
XNOR U10023 ( .A(b[2004]), .B(n6014), .Z(c[2004]) );
XNOR U10024 ( .A(a[2004]), .B(c2004), .Z(n6014) );
XOR U10025 ( .A(c2005), .B(n6015), .Z(c2006) );
ANDN U10026 ( .B(n6016), .A(n6017), .Z(n6015) );
XOR U10027 ( .A(c2005), .B(b[2005]), .Z(n6016) );
XNOR U10028 ( .A(b[2005]), .B(n6017), .Z(c[2005]) );
XNOR U10029 ( .A(a[2005]), .B(c2005), .Z(n6017) );
XOR U10030 ( .A(c2006), .B(n6018), .Z(c2007) );
ANDN U10031 ( .B(n6019), .A(n6020), .Z(n6018) );
XOR U10032 ( .A(c2006), .B(b[2006]), .Z(n6019) );
XNOR U10033 ( .A(b[2006]), .B(n6020), .Z(c[2006]) );
XNOR U10034 ( .A(a[2006]), .B(c2006), .Z(n6020) );
XOR U10035 ( .A(c2007), .B(n6021), .Z(c2008) );
ANDN U10036 ( .B(n6022), .A(n6023), .Z(n6021) );
XOR U10037 ( .A(c2007), .B(b[2007]), .Z(n6022) );
XNOR U10038 ( .A(b[2007]), .B(n6023), .Z(c[2007]) );
XNOR U10039 ( .A(a[2007]), .B(c2007), .Z(n6023) );
XOR U10040 ( .A(c2008), .B(n6024), .Z(c2009) );
ANDN U10041 ( .B(n6025), .A(n6026), .Z(n6024) );
XOR U10042 ( .A(c2008), .B(b[2008]), .Z(n6025) );
XNOR U10043 ( .A(b[2008]), .B(n6026), .Z(c[2008]) );
XNOR U10044 ( .A(a[2008]), .B(c2008), .Z(n6026) );
XOR U10045 ( .A(c2009), .B(n6027), .Z(c2010) );
ANDN U10046 ( .B(n6028), .A(n6029), .Z(n6027) );
XOR U10047 ( .A(c2009), .B(b[2009]), .Z(n6028) );
XNOR U10048 ( .A(b[2009]), .B(n6029), .Z(c[2009]) );
XNOR U10049 ( .A(a[2009]), .B(c2009), .Z(n6029) );
XOR U10050 ( .A(c2010), .B(n6030), .Z(c2011) );
ANDN U10051 ( .B(n6031), .A(n6032), .Z(n6030) );
XOR U10052 ( .A(c2010), .B(b[2010]), .Z(n6031) );
XNOR U10053 ( .A(b[2010]), .B(n6032), .Z(c[2010]) );
XNOR U10054 ( .A(a[2010]), .B(c2010), .Z(n6032) );
XOR U10055 ( .A(c2011), .B(n6033), .Z(c2012) );
ANDN U10056 ( .B(n6034), .A(n6035), .Z(n6033) );
XOR U10057 ( .A(c2011), .B(b[2011]), .Z(n6034) );
XNOR U10058 ( .A(b[2011]), .B(n6035), .Z(c[2011]) );
XNOR U10059 ( .A(a[2011]), .B(c2011), .Z(n6035) );
XOR U10060 ( .A(c2012), .B(n6036), .Z(c2013) );
ANDN U10061 ( .B(n6037), .A(n6038), .Z(n6036) );
XOR U10062 ( .A(c2012), .B(b[2012]), .Z(n6037) );
XNOR U10063 ( .A(b[2012]), .B(n6038), .Z(c[2012]) );
XNOR U10064 ( .A(a[2012]), .B(c2012), .Z(n6038) );
XOR U10065 ( .A(c2013), .B(n6039), .Z(c2014) );
ANDN U10066 ( .B(n6040), .A(n6041), .Z(n6039) );
XOR U10067 ( .A(c2013), .B(b[2013]), .Z(n6040) );
XNOR U10068 ( .A(b[2013]), .B(n6041), .Z(c[2013]) );
XNOR U10069 ( .A(a[2013]), .B(c2013), .Z(n6041) );
XOR U10070 ( .A(c2014), .B(n6042), .Z(c2015) );
ANDN U10071 ( .B(n6043), .A(n6044), .Z(n6042) );
XOR U10072 ( .A(c2014), .B(b[2014]), .Z(n6043) );
XNOR U10073 ( .A(b[2014]), .B(n6044), .Z(c[2014]) );
XNOR U10074 ( .A(a[2014]), .B(c2014), .Z(n6044) );
XOR U10075 ( .A(c2015), .B(n6045), .Z(c2016) );
ANDN U10076 ( .B(n6046), .A(n6047), .Z(n6045) );
XOR U10077 ( .A(c2015), .B(b[2015]), .Z(n6046) );
XNOR U10078 ( .A(b[2015]), .B(n6047), .Z(c[2015]) );
XNOR U10079 ( .A(a[2015]), .B(c2015), .Z(n6047) );
XOR U10080 ( .A(c2016), .B(n6048), .Z(c2017) );
ANDN U10081 ( .B(n6049), .A(n6050), .Z(n6048) );
XOR U10082 ( .A(c2016), .B(b[2016]), .Z(n6049) );
XNOR U10083 ( .A(b[2016]), .B(n6050), .Z(c[2016]) );
XNOR U10084 ( .A(a[2016]), .B(c2016), .Z(n6050) );
XOR U10085 ( .A(c2017), .B(n6051), .Z(c2018) );
ANDN U10086 ( .B(n6052), .A(n6053), .Z(n6051) );
XOR U10087 ( .A(c2017), .B(b[2017]), .Z(n6052) );
XNOR U10088 ( .A(b[2017]), .B(n6053), .Z(c[2017]) );
XNOR U10089 ( .A(a[2017]), .B(c2017), .Z(n6053) );
XOR U10090 ( .A(c2018), .B(n6054), .Z(c2019) );
ANDN U10091 ( .B(n6055), .A(n6056), .Z(n6054) );
XOR U10092 ( .A(c2018), .B(b[2018]), .Z(n6055) );
XNOR U10093 ( .A(b[2018]), .B(n6056), .Z(c[2018]) );
XNOR U10094 ( .A(a[2018]), .B(c2018), .Z(n6056) );
XOR U10095 ( .A(c2019), .B(n6057), .Z(c2020) );
ANDN U10096 ( .B(n6058), .A(n6059), .Z(n6057) );
XOR U10097 ( .A(c2019), .B(b[2019]), .Z(n6058) );
XNOR U10098 ( .A(b[2019]), .B(n6059), .Z(c[2019]) );
XNOR U10099 ( .A(a[2019]), .B(c2019), .Z(n6059) );
XOR U10100 ( .A(c2020), .B(n6060), .Z(c2021) );
ANDN U10101 ( .B(n6061), .A(n6062), .Z(n6060) );
XOR U10102 ( .A(c2020), .B(b[2020]), .Z(n6061) );
XNOR U10103 ( .A(b[2020]), .B(n6062), .Z(c[2020]) );
XNOR U10104 ( .A(a[2020]), .B(c2020), .Z(n6062) );
XOR U10105 ( .A(c2021), .B(n6063), .Z(c2022) );
ANDN U10106 ( .B(n6064), .A(n6065), .Z(n6063) );
XOR U10107 ( .A(c2021), .B(b[2021]), .Z(n6064) );
XNOR U10108 ( .A(b[2021]), .B(n6065), .Z(c[2021]) );
XNOR U10109 ( .A(a[2021]), .B(c2021), .Z(n6065) );
XOR U10110 ( .A(c2022), .B(n6066), .Z(c2023) );
ANDN U10111 ( .B(n6067), .A(n6068), .Z(n6066) );
XOR U10112 ( .A(c2022), .B(b[2022]), .Z(n6067) );
XNOR U10113 ( .A(b[2022]), .B(n6068), .Z(c[2022]) );
XNOR U10114 ( .A(a[2022]), .B(c2022), .Z(n6068) );
XOR U10115 ( .A(c2023), .B(n6069), .Z(c2024) );
ANDN U10116 ( .B(n6070), .A(n6071), .Z(n6069) );
XOR U10117 ( .A(c2023), .B(b[2023]), .Z(n6070) );
XNOR U10118 ( .A(b[2023]), .B(n6071), .Z(c[2023]) );
XNOR U10119 ( .A(a[2023]), .B(c2023), .Z(n6071) );
XOR U10120 ( .A(c2024), .B(n6072), .Z(c2025) );
ANDN U10121 ( .B(n6073), .A(n6074), .Z(n6072) );
XOR U10122 ( .A(c2024), .B(b[2024]), .Z(n6073) );
XNOR U10123 ( .A(b[2024]), .B(n6074), .Z(c[2024]) );
XNOR U10124 ( .A(a[2024]), .B(c2024), .Z(n6074) );
XOR U10125 ( .A(c2025), .B(n6075), .Z(c2026) );
ANDN U10126 ( .B(n6076), .A(n6077), .Z(n6075) );
XOR U10127 ( .A(c2025), .B(b[2025]), .Z(n6076) );
XNOR U10128 ( .A(b[2025]), .B(n6077), .Z(c[2025]) );
XNOR U10129 ( .A(a[2025]), .B(c2025), .Z(n6077) );
XOR U10130 ( .A(c2026), .B(n6078), .Z(c2027) );
ANDN U10131 ( .B(n6079), .A(n6080), .Z(n6078) );
XOR U10132 ( .A(c2026), .B(b[2026]), .Z(n6079) );
XNOR U10133 ( .A(b[2026]), .B(n6080), .Z(c[2026]) );
XNOR U10134 ( .A(a[2026]), .B(c2026), .Z(n6080) );
XOR U10135 ( .A(c2027), .B(n6081), .Z(c2028) );
ANDN U10136 ( .B(n6082), .A(n6083), .Z(n6081) );
XOR U10137 ( .A(c2027), .B(b[2027]), .Z(n6082) );
XNOR U10138 ( .A(b[2027]), .B(n6083), .Z(c[2027]) );
XNOR U10139 ( .A(a[2027]), .B(c2027), .Z(n6083) );
XOR U10140 ( .A(c2028), .B(n6084), .Z(c2029) );
ANDN U10141 ( .B(n6085), .A(n6086), .Z(n6084) );
XOR U10142 ( .A(c2028), .B(b[2028]), .Z(n6085) );
XNOR U10143 ( .A(b[2028]), .B(n6086), .Z(c[2028]) );
XNOR U10144 ( .A(a[2028]), .B(c2028), .Z(n6086) );
XOR U10145 ( .A(c2029), .B(n6087), .Z(c2030) );
ANDN U10146 ( .B(n6088), .A(n6089), .Z(n6087) );
XOR U10147 ( .A(c2029), .B(b[2029]), .Z(n6088) );
XNOR U10148 ( .A(b[2029]), .B(n6089), .Z(c[2029]) );
XNOR U10149 ( .A(a[2029]), .B(c2029), .Z(n6089) );
XOR U10150 ( .A(c2030), .B(n6090), .Z(c2031) );
ANDN U10151 ( .B(n6091), .A(n6092), .Z(n6090) );
XOR U10152 ( .A(c2030), .B(b[2030]), .Z(n6091) );
XNOR U10153 ( .A(b[2030]), .B(n6092), .Z(c[2030]) );
XNOR U10154 ( .A(a[2030]), .B(c2030), .Z(n6092) );
XOR U10155 ( .A(c2031), .B(n6093), .Z(c2032) );
ANDN U10156 ( .B(n6094), .A(n6095), .Z(n6093) );
XOR U10157 ( .A(c2031), .B(b[2031]), .Z(n6094) );
XNOR U10158 ( .A(b[2031]), .B(n6095), .Z(c[2031]) );
XNOR U10159 ( .A(a[2031]), .B(c2031), .Z(n6095) );
XOR U10160 ( .A(c2032), .B(n6096), .Z(c2033) );
ANDN U10161 ( .B(n6097), .A(n6098), .Z(n6096) );
XOR U10162 ( .A(c2032), .B(b[2032]), .Z(n6097) );
XNOR U10163 ( .A(b[2032]), .B(n6098), .Z(c[2032]) );
XNOR U10164 ( .A(a[2032]), .B(c2032), .Z(n6098) );
XOR U10165 ( .A(c2033), .B(n6099), .Z(c2034) );
ANDN U10166 ( .B(n6100), .A(n6101), .Z(n6099) );
XOR U10167 ( .A(c2033), .B(b[2033]), .Z(n6100) );
XNOR U10168 ( .A(b[2033]), .B(n6101), .Z(c[2033]) );
XNOR U10169 ( .A(a[2033]), .B(c2033), .Z(n6101) );
XOR U10170 ( .A(c2034), .B(n6102), .Z(c2035) );
ANDN U10171 ( .B(n6103), .A(n6104), .Z(n6102) );
XOR U10172 ( .A(c2034), .B(b[2034]), .Z(n6103) );
XNOR U10173 ( .A(b[2034]), .B(n6104), .Z(c[2034]) );
XNOR U10174 ( .A(a[2034]), .B(c2034), .Z(n6104) );
XOR U10175 ( .A(c2035), .B(n6105), .Z(c2036) );
ANDN U10176 ( .B(n6106), .A(n6107), .Z(n6105) );
XOR U10177 ( .A(c2035), .B(b[2035]), .Z(n6106) );
XNOR U10178 ( .A(b[2035]), .B(n6107), .Z(c[2035]) );
XNOR U10179 ( .A(a[2035]), .B(c2035), .Z(n6107) );
XOR U10180 ( .A(c2036), .B(n6108), .Z(c2037) );
ANDN U10181 ( .B(n6109), .A(n6110), .Z(n6108) );
XOR U10182 ( .A(c2036), .B(b[2036]), .Z(n6109) );
XNOR U10183 ( .A(b[2036]), .B(n6110), .Z(c[2036]) );
XNOR U10184 ( .A(a[2036]), .B(c2036), .Z(n6110) );
XOR U10185 ( .A(c2037), .B(n6111), .Z(c2038) );
ANDN U10186 ( .B(n6112), .A(n6113), .Z(n6111) );
XOR U10187 ( .A(c2037), .B(b[2037]), .Z(n6112) );
XNOR U10188 ( .A(b[2037]), .B(n6113), .Z(c[2037]) );
XNOR U10189 ( .A(a[2037]), .B(c2037), .Z(n6113) );
XOR U10190 ( .A(c2038), .B(n6114), .Z(c2039) );
ANDN U10191 ( .B(n6115), .A(n6116), .Z(n6114) );
XOR U10192 ( .A(c2038), .B(b[2038]), .Z(n6115) );
XNOR U10193 ( .A(b[2038]), .B(n6116), .Z(c[2038]) );
XNOR U10194 ( .A(a[2038]), .B(c2038), .Z(n6116) );
XOR U10195 ( .A(c2039), .B(n6117), .Z(c2040) );
ANDN U10196 ( .B(n6118), .A(n6119), .Z(n6117) );
XOR U10197 ( .A(c2039), .B(b[2039]), .Z(n6118) );
XNOR U10198 ( .A(b[2039]), .B(n6119), .Z(c[2039]) );
XNOR U10199 ( .A(a[2039]), .B(c2039), .Z(n6119) );
XOR U10200 ( .A(c2040), .B(n6120), .Z(c2041) );
ANDN U10201 ( .B(n6121), .A(n6122), .Z(n6120) );
XOR U10202 ( .A(c2040), .B(b[2040]), .Z(n6121) );
XNOR U10203 ( .A(b[2040]), .B(n6122), .Z(c[2040]) );
XNOR U10204 ( .A(a[2040]), .B(c2040), .Z(n6122) );
XOR U10205 ( .A(c2041), .B(n6123), .Z(c2042) );
ANDN U10206 ( .B(n6124), .A(n6125), .Z(n6123) );
XOR U10207 ( .A(c2041), .B(b[2041]), .Z(n6124) );
XNOR U10208 ( .A(b[2041]), .B(n6125), .Z(c[2041]) );
XNOR U10209 ( .A(a[2041]), .B(c2041), .Z(n6125) );
XOR U10210 ( .A(c2042), .B(n6126), .Z(c2043) );
ANDN U10211 ( .B(n6127), .A(n6128), .Z(n6126) );
XOR U10212 ( .A(c2042), .B(b[2042]), .Z(n6127) );
XNOR U10213 ( .A(b[2042]), .B(n6128), .Z(c[2042]) );
XNOR U10214 ( .A(a[2042]), .B(c2042), .Z(n6128) );
XOR U10215 ( .A(c2043), .B(n6129), .Z(c2044) );
ANDN U10216 ( .B(n6130), .A(n6131), .Z(n6129) );
XOR U10217 ( .A(c2043), .B(b[2043]), .Z(n6130) );
XNOR U10218 ( .A(b[2043]), .B(n6131), .Z(c[2043]) );
XNOR U10219 ( .A(a[2043]), .B(c2043), .Z(n6131) );
XOR U10220 ( .A(c2044), .B(n6132), .Z(c2045) );
ANDN U10221 ( .B(n6133), .A(n6134), .Z(n6132) );
XOR U10222 ( .A(c2044), .B(b[2044]), .Z(n6133) );
XNOR U10223 ( .A(b[2044]), .B(n6134), .Z(c[2044]) );
XNOR U10224 ( .A(a[2044]), .B(c2044), .Z(n6134) );
XOR U10225 ( .A(c2045), .B(n6135), .Z(c2046) );
ANDN U10226 ( .B(n6136), .A(n6137), .Z(n6135) );
XOR U10227 ( .A(c2045), .B(b[2045]), .Z(n6136) );
XNOR U10228 ( .A(b[2045]), .B(n6137), .Z(c[2045]) );
XNOR U10229 ( .A(a[2045]), .B(c2045), .Z(n6137) );
XOR U10230 ( .A(c2046), .B(n6138), .Z(c2047) );
ANDN U10231 ( .B(n6139), .A(n6140), .Z(n6138) );
XOR U10232 ( .A(c2046), .B(b[2046]), .Z(n6139) );
XNOR U10233 ( .A(b[2046]), .B(n6140), .Z(c[2046]) );
XNOR U10234 ( .A(a[2046]), .B(c2046), .Z(n6140) );
XOR U10235 ( .A(c2047), .B(n6141), .Z(c2048) );
ANDN U10236 ( .B(n6142), .A(n6143), .Z(n6141) );
XOR U10237 ( .A(c2047), .B(b[2047]), .Z(n6142) );
XNOR U10238 ( .A(b[2047]), .B(n6143), .Z(c[2047]) );
XNOR U10239 ( .A(a[2047]), .B(c2047), .Z(n6143) );
XOR U10240 ( .A(c2048), .B(n6144), .Z(c2049) );
ANDN U10241 ( .B(n6145), .A(n6146), .Z(n6144) );
XOR U10242 ( .A(c2048), .B(b[2048]), .Z(n6145) );
XNOR U10243 ( .A(b[2048]), .B(n6146), .Z(c[2048]) );
XNOR U10244 ( .A(a[2048]), .B(c2048), .Z(n6146) );
XOR U10245 ( .A(c2049), .B(n6147), .Z(c2050) );
ANDN U10246 ( .B(n6148), .A(n6149), .Z(n6147) );
XOR U10247 ( .A(c2049), .B(b[2049]), .Z(n6148) );
XNOR U10248 ( .A(b[2049]), .B(n6149), .Z(c[2049]) );
XNOR U10249 ( .A(a[2049]), .B(c2049), .Z(n6149) );
XOR U10250 ( .A(c2050), .B(n6150), .Z(c2051) );
ANDN U10251 ( .B(n6151), .A(n6152), .Z(n6150) );
XOR U10252 ( .A(c2050), .B(b[2050]), .Z(n6151) );
XNOR U10253 ( .A(b[2050]), .B(n6152), .Z(c[2050]) );
XNOR U10254 ( .A(a[2050]), .B(c2050), .Z(n6152) );
XOR U10255 ( .A(c2051), .B(n6153), .Z(c2052) );
ANDN U10256 ( .B(n6154), .A(n6155), .Z(n6153) );
XOR U10257 ( .A(c2051), .B(b[2051]), .Z(n6154) );
XNOR U10258 ( .A(b[2051]), .B(n6155), .Z(c[2051]) );
XNOR U10259 ( .A(a[2051]), .B(c2051), .Z(n6155) );
XOR U10260 ( .A(c2052), .B(n6156), .Z(c2053) );
ANDN U10261 ( .B(n6157), .A(n6158), .Z(n6156) );
XOR U10262 ( .A(c2052), .B(b[2052]), .Z(n6157) );
XNOR U10263 ( .A(b[2052]), .B(n6158), .Z(c[2052]) );
XNOR U10264 ( .A(a[2052]), .B(c2052), .Z(n6158) );
XOR U10265 ( .A(c2053), .B(n6159), .Z(c2054) );
ANDN U10266 ( .B(n6160), .A(n6161), .Z(n6159) );
XOR U10267 ( .A(c2053), .B(b[2053]), .Z(n6160) );
XNOR U10268 ( .A(b[2053]), .B(n6161), .Z(c[2053]) );
XNOR U10269 ( .A(a[2053]), .B(c2053), .Z(n6161) );
XOR U10270 ( .A(c2054), .B(n6162), .Z(c2055) );
ANDN U10271 ( .B(n6163), .A(n6164), .Z(n6162) );
XOR U10272 ( .A(c2054), .B(b[2054]), .Z(n6163) );
XNOR U10273 ( .A(b[2054]), .B(n6164), .Z(c[2054]) );
XNOR U10274 ( .A(a[2054]), .B(c2054), .Z(n6164) );
XOR U10275 ( .A(c2055), .B(n6165), .Z(c2056) );
ANDN U10276 ( .B(n6166), .A(n6167), .Z(n6165) );
XOR U10277 ( .A(c2055), .B(b[2055]), .Z(n6166) );
XNOR U10278 ( .A(b[2055]), .B(n6167), .Z(c[2055]) );
XNOR U10279 ( .A(a[2055]), .B(c2055), .Z(n6167) );
XOR U10280 ( .A(c2056), .B(n6168), .Z(c2057) );
ANDN U10281 ( .B(n6169), .A(n6170), .Z(n6168) );
XOR U10282 ( .A(c2056), .B(b[2056]), .Z(n6169) );
XNOR U10283 ( .A(b[2056]), .B(n6170), .Z(c[2056]) );
XNOR U10284 ( .A(a[2056]), .B(c2056), .Z(n6170) );
XOR U10285 ( .A(c2057), .B(n6171), .Z(c2058) );
ANDN U10286 ( .B(n6172), .A(n6173), .Z(n6171) );
XOR U10287 ( .A(c2057), .B(b[2057]), .Z(n6172) );
XNOR U10288 ( .A(b[2057]), .B(n6173), .Z(c[2057]) );
XNOR U10289 ( .A(a[2057]), .B(c2057), .Z(n6173) );
XOR U10290 ( .A(c2058), .B(n6174), .Z(c2059) );
ANDN U10291 ( .B(n6175), .A(n6176), .Z(n6174) );
XOR U10292 ( .A(c2058), .B(b[2058]), .Z(n6175) );
XNOR U10293 ( .A(b[2058]), .B(n6176), .Z(c[2058]) );
XNOR U10294 ( .A(a[2058]), .B(c2058), .Z(n6176) );
XOR U10295 ( .A(c2059), .B(n6177), .Z(c2060) );
ANDN U10296 ( .B(n6178), .A(n6179), .Z(n6177) );
XOR U10297 ( .A(c2059), .B(b[2059]), .Z(n6178) );
XNOR U10298 ( .A(b[2059]), .B(n6179), .Z(c[2059]) );
XNOR U10299 ( .A(a[2059]), .B(c2059), .Z(n6179) );
XOR U10300 ( .A(c2060), .B(n6180), .Z(c2061) );
ANDN U10301 ( .B(n6181), .A(n6182), .Z(n6180) );
XOR U10302 ( .A(c2060), .B(b[2060]), .Z(n6181) );
XNOR U10303 ( .A(b[2060]), .B(n6182), .Z(c[2060]) );
XNOR U10304 ( .A(a[2060]), .B(c2060), .Z(n6182) );
XOR U10305 ( .A(c2061), .B(n6183), .Z(c2062) );
ANDN U10306 ( .B(n6184), .A(n6185), .Z(n6183) );
XOR U10307 ( .A(c2061), .B(b[2061]), .Z(n6184) );
XNOR U10308 ( .A(b[2061]), .B(n6185), .Z(c[2061]) );
XNOR U10309 ( .A(a[2061]), .B(c2061), .Z(n6185) );
XOR U10310 ( .A(c2062), .B(n6186), .Z(c2063) );
ANDN U10311 ( .B(n6187), .A(n6188), .Z(n6186) );
XOR U10312 ( .A(c2062), .B(b[2062]), .Z(n6187) );
XNOR U10313 ( .A(b[2062]), .B(n6188), .Z(c[2062]) );
XNOR U10314 ( .A(a[2062]), .B(c2062), .Z(n6188) );
XOR U10315 ( .A(c2063), .B(n6189), .Z(c2064) );
ANDN U10316 ( .B(n6190), .A(n6191), .Z(n6189) );
XOR U10317 ( .A(c2063), .B(b[2063]), .Z(n6190) );
XNOR U10318 ( .A(b[2063]), .B(n6191), .Z(c[2063]) );
XNOR U10319 ( .A(a[2063]), .B(c2063), .Z(n6191) );
XOR U10320 ( .A(c2064), .B(n6192), .Z(c2065) );
ANDN U10321 ( .B(n6193), .A(n6194), .Z(n6192) );
XOR U10322 ( .A(c2064), .B(b[2064]), .Z(n6193) );
XNOR U10323 ( .A(b[2064]), .B(n6194), .Z(c[2064]) );
XNOR U10324 ( .A(a[2064]), .B(c2064), .Z(n6194) );
XOR U10325 ( .A(c2065), .B(n6195), .Z(c2066) );
ANDN U10326 ( .B(n6196), .A(n6197), .Z(n6195) );
XOR U10327 ( .A(c2065), .B(b[2065]), .Z(n6196) );
XNOR U10328 ( .A(b[2065]), .B(n6197), .Z(c[2065]) );
XNOR U10329 ( .A(a[2065]), .B(c2065), .Z(n6197) );
XOR U10330 ( .A(c2066), .B(n6198), .Z(c2067) );
ANDN U10331 ( .B(n6199), .A(n6200), .Z(n6198) );
XOR U10332 ( .A(c2066), .B(b[2066]), .Z(n6199) );
XNOR U10333 ( .A(b[2066]), .B(n6200), .Z(c[2066]) );
XNOR U10334 ( .A(a[2066]), .B(c2066), .Z(n6200) );
XOR U10335 ( .A(c2067), .B(n6201), .Z(c2068) );
ANDN U10336 ( .B(n6202), .A(n6203), .Z(n6201) );
XOR U10337 ( .A(c2067), .B(b[2067]), .Z(n6202) );
XNOR U10338 ( .A(b[2067]), .B(n6203), .Z(c[2067]) );
XNOR U10339 ( .A(a[2067]), .B(c2067), .Z(n6203) );
XOR U10340 ( .A(c2068), .B(n6204), .Z(c2069) );
ANDN U10341 ( .B(n6205), .A(n6206), .Z(n6204) );
XOR U10342 ( .A(c2068), .B(b[2068]), .Z(n6205) );
XNOR U10343 ( .A(b[2068]), .B(n6206), .Z(c[2068]) );
XNOR U10344 ( .A(a[2068]), .B(c2068), .Z(n6206) );
XOR U10345 ( .A(c2069), .B(n6207), .Z(c2070) );
ANDN U10346 ( .B(n6208), .A(n6209), .Z(n6207) );
XOR U10347 ( .A(c2069), .B(b[2069]), .Z(n6208) );
XNOR U10348 ( .A(b[2069]), .B(n6209), .Z(c[2069]) );
XNOR U10349 ( .A(a[2069]), .B(c2069), .Z(n6209) );
XOR U10350 ( .A(c2070), .B(n6210), .Z(c2071) );
ANDN U10351 ( .B(n6211), .A(n6212), .Z(n6210) );
XOR U10352 ( .A(c2070), .B(b[2070]), .Z(n6211) );
XNOR U10353 ( .A(b[2070]), .B(n6212), .Z(c[2070]) );
XNOR U10354 ( .A(a[2070]), .B(c2070), .Z(n6212) );
XOR U10355 ( .A(c2071), .B(n6213), .Z(c2072) );
ANDN U10356 ( .B(n6214), .A(n6215), .Z(n6213) );
XOR U10357 ( .A(c2071), .B(b[2071]), .Z(n6214) );
XNOR U10358 ( .A(b[2071]), .B(n6215), .Z(c[2071]) );
XNOR U10359 ( .A(a[2071]), .B(c2071), .Z(n6215) );
XOR U10360 ( .A(c2072), .B(n6216), .Z(c2073) );
ANDN U10361 ( .B(n6217), .A(n6218), .Z(n6216) );
XOR U10362 ( .A(c2072), .B(b[2072]), .Z(n6217) );
XNOR U10363 ( .A(b[2072]), .B(n6218), .Z(c[2072]) );
XNOR U10364 ( .A(a[2072]), .B(c2072), .Z(n6218) );
XOR U10365 ( .A(c2073), .B(n6219), .Z(c2074) );
ANDN U10366 ( .B(n6220), .A(n6221), .Z(n6219) );
XOR U10367 ( .A(c2073), .B(b[2073]), .Z(n6220) );
XNOR U10368 ( .A(b[2073]), .B(n6221), .Z(c[2073]) );
XNOR U10369 ( .A(a[2073]), .B(c2073), .Z(n6221) );
XOR U10370 ( .A(c2074), .B(n6222), .Z(c2075) );
ANDN U10371 ( .B(n6223), .A(n6224), .Z(n6222) );
XOR U10372 ( .A(c2074), .B(b[2074]), .Z(n6223) );
XNOR U10373 ( .A(b[2074]), .B(n6224), .Z(c[2074]) );
XNOR U10374 ( .A(a[2074]), .B(c2074), .Z(n6224) );
XOR U10375 ( .A(c2075), .B(n6225), .Z(c2076) );
ANDN U10376 ( .B(n6226), .A(n6227), .Z(n6225) );
XOR U10377 ( .A(c2075), .B(b[2075]), .Z(n6226) );
XNOR U10378 ( .A(b[2075]), .B(n6227), .Z(c[2075]) );
XNOR U10379 ( .A(a[2075]), .B(c2075), .Z(n6227) );
XOR U10380 ( .A(c2076), .B(n6228), .Z(c2077) );
ANDN U10381 ( .B(n6229), .A(n6230), .Z(n6228) );
XOR U10382 ( .A(c2076), .B(b[2076]), .Z(n6229) );
XNOR U10383 ( .A(b[2076]), .B(n6230), .Z(c[2076]) );
XNOR U10384 ( .A(a[2076]), .B(c2076), .Z(n6230) );
XOR U10385 ( .A(c2077), .B(n6231), .Z(c2078) );
ANDN U10386 ( .B(n6232), .A(n6233), .Z(n6231) );
XOR U10387 ( .A(c2077), .B(b[2077]), .Z(n6232) );
XNOR U10388 ( .A(b[2077]), .B(n6233), .Z(c[2077]) );
XNOR U10389 ( .A(a[2077]), .B(c2077), .Z(n6233) );
XOR U10390 ( .A(c2078), .B(n6234), .Z(c2079) );
ANDN U10391 ( .B(n6235), .A(n6236), .Z(n6234) );
XOR U10392 ( .A(c2078), .B(b[2078]), .Z(n6235) );
XNOR U10393 ( .A(b[2078]), .B(n6236), .Z(c[2078]) );
XNOR U10394 ( .A(a[2078]), .B(c2078), .Z(n6236) );
XOR U10395 ( .A(c2079), .B(n6237), .Z(c2080) );
ANDN U10396 ( .B(n6238), .A(n6239), .Z(n6237) );
XOR U10397 ( .A(c2079), .B(b[2079]), .Z(n6238) );
XNOR U10398 ( .A(b[2079]), .B(n6239), .Z(c[2079]) );
XNOR U10399 ( .A(a[2079]), .B(c2079), .Z(n6239) );
XOR U10400 ( .A(c2080), .B(n6240), .Z(c2081) );
ANDN U10401 ( .B(n6241), .A(n6242), .Z(n6240) );
XOR U10402 ( .A(c2080), .B(b[2080]), .Z(n6241) );
XNOR U10403 ( .A(b[2080]), .B(n6242), .Z(c[2080]) );
XNOR U10404 ( .A(a[2080]), .B(c2080), .Z(n6242) );
XOR U10405 ( .A(c2081), .B(n6243), .Z(c2082) );
ANDN U10406 ( .B(n6244), .A(n6245), .Z(n6243) );
XOR U10407 ( .A(c2081), .B(b[2081]), .Z(n6244) );
XNOR U10408 ( .A(b[2081]), .B(n6245), .Z(c[2081]) );
XNOR U10409 ( .A(a[2081]), .B(c2081), .Z(n6245) );
XOR U10410 ( .A(c2082), .B(n6246), .Z(c2083) );
ANDN U10411 ( .B(n6247), .A(n6248), .Z(n6246) );
XOR U10412 ( .A(c2082), .B(b[2082]), .Z(n6247) );
XNOR U10413 ( .A(b[2082]), .B(n6248), .Z(c[2082]) );
XNOR U10414 ( .A(a[2082]), .B(c2082), .Z(n6248) );
XOR U10415 ( .A(c2083), .B(n6249), .Z(c2084) );
ANDN U10416 ( .B(n6250), .A(n6251), .Z(n6249) );
XOR U10417 ( .A(c2083), .B(b[2083]), .Z(n6250) );
XNOR U10418 ( .A(b[2083]), .B(n6251), .Z(c[2083]) );
XNOR U10419 ( .A(a[2083]), .B(c2083), .Z(n6251) );
XOR U10420 ( .A(c2084), .B(n6252), .Z(c2085) );
ANDN U10421 ( .B(n6253), .A(n6254), .Z(n6252) );
XOR U10422 ( .A(c2084), .B(b[2084]), .Z(n6253) );
XNOR U10423 ( .A(b[2084]), .B(n6254), .Z(c[2084]) );
XNOR U10424 ( .A(a[2084]), .B(c2084), .Z(n6254) );
XOR U10425 ( .A(c2085), .B(n6255), .Z(c2086) );
ANDN U10426 ( .B(n6256), .A(n6257), .Z(n6255) );
XOR U10427 ( .A(c2085), .B(b[2085]), .Z(n6256) );
XNOR U10428 ( .A(b[2085]), .B(n6257), .Z(c[2085]) );
XNOR U10429 ( .A(a[2085]), .B(c2085), .Z(n6257) );
XOR U10430 ( .A(c2086), .B(n6258), .Z(c2087) );
ANDN U10431 ( .B(n6259), .A(n6260), .Z(n6258) );
XOR U10432 ( .A(c2086), .B(b[2086]), .Z(n6259) );
XNOR U10433 ( .A(b[2086]), .B(n6260), .Z(c[2086]) );
XNOR U10434 ( .A(a[2086]), .B(c2086), .Z(n6260) );
XOR U10435 ( .A(c2087), .B(n6261), .Z(c2088) );
ANDN U10436 ( .B(n6262), .A(n6263), .Z(n6261) );
XOR U10437 ( .A(c2087), .B(b[2087]), .Z(n6262) );
XNOR U10438 ( .A(b[2087]), .B(n6263), .Z(c[2087]) );
XNOR U10439 ( .A(a[2087]), .B(c2087), .Z(n6263) );
XOR U10440 ( .A(c2088), .B(n6264), .Z(c2089) );
ANDN U10441 ( .B(n6265), .A(n6266), .Z(n6264) );
XOR U10442 ( .A(c2088), .B(b[2088]), .Z(n6265) );
XNOR U10443 ( .A(b[2088]), .B(n6266), .Z(c[2088]) );
XNOR U10444 ( .A(a[2088]), .B(c2088), .Z(n6266) );
XOR U10445 ( .A(c2089), .B(n6267), .Z(c2090) );
ANDN U10446 ( .B(n6268), .A(n6269), .Z(n6267) );
XOR U10447 ( .A(c2089), .B(b[2089]), .Z(n6268) );
XNOR U10448 ( .A(b[2089]), .B(n6269), .Z(c[2089]) );
XNOR U10449 ( .A(a[2089]), .B(c2089), .Z(n6269) );
XOR U10450 ( .A(c2090), .B(n6270), .Z(c2091) );
ANDN U10451 ( .B(n6271), .A(n6272), .Z(n6270) );
XOR U10452 ( .A(c2090), .B(b[2090]), .Z(n6271) );
XNOR U10453 ( .A(b[2090]), .B(n6272), .Z(c[2090]) );
XNOR U10454 ( .A(a[2090]), .B(c2090), .Z(n6272) );
XOR U10455 ( .A(c2091), .B(n6273), .Z(c2092) );
ANDN U10456 ( .B(n6274), .A(n6275), .Z(n6273) );
XOR U10457 ( .A(c2091), .B(b[2091]), .Z(n6274) );
XNOR U10458 ( .A(b[2091]), .B(n6275), .Z(c[2091]) );
XNOR U10459 ( .A(a[2091]), .B(c2091), .Z(n6275) );
XOR U10460 ( .A(c2092), .B(n6276), .Z(c2093) );
ANDN U10461 ( .B(n6277), .A(n6278), .Z(n6276) );
XOR U10462 ( .A(c2092), .B(b[2092]), .Z(n6277) );
XNOR U10463 ( .A(b[2092]), .B(n6278), .Z(c[2092]) );
XNOR U10464 ( .A(a[2092]), .B(c2092), .Z(n6278) );
XOR U10465 ( .A(c2093), .B(n6279), .Z(c2094) );
ANDN U10466 ( .B(n6280), .A(n6281), .Z(n6279) );
XOR U10467 ( .A(c2093), .B(b[2093]), .Z(n6280) );
XNOR U10468 ( .A(b[2093]), .B(n6281), .Z(c[2093]) );
XNOR U10469 ( .A(a[2093]), .B(c2093), .Z(n6281) );
XOR U10470 ( .A(c2094), .B(n6282), .Z(c2095) );
ANDN U10471 ( .B(n6283), .A(n6284), .Z(n6282) );
XOR U10472 ( .A(c2094), .B(b[2094]), .Z(n6283) );
XNOR U10473 ( .A(b[2094]), .B(n6284), .Z(c[2094]) );
XNOR U10474 ( .A(a[2094]), .B(c2094), .Z(n6284) );
XOR U10475 ( .A(c2095), .B(n6285), .Z(c2096) );
ANDN U10476 ( .B(n6286), .A(n6287), .Z(n6285) );
XOR U10477 ( .A(c2095), .B(b[2095]), .Z(n6286) );
XNOR U10478 ( .A(b[2095]), .B(n6287), .Z(c[2095]) );
XNOR U10479 ( .A(a[2095]), .B(c2095), .Z(n6287) );
XOR U10480 ( .A(c2096), .B(n6288), .Z(c2097) );
ANDN U10481 ( .B(n6289), .A(n6290), .Z(n6288) );
XOR U10482 ( .A(c2096), .B(b[2096]), .Z(n6289) );
XNOR U10483 ( .A(b[2096]), .B(n6290), .Z(c[2096]) );
XNOR U10484 ( .A(a[2096]), .B(c2096), .Z(n6290) );
XOR U10485 ( .A(c2097), .B(n6291), .Z(c2098) );
ANDN U10486 ( .B(n6292), .A(n6293), .Z(n6291) );
XOR U10487 ( .A(c2097), .B(b[2097]), .Z(n6292) );
XNOR U10488 ( .A(b[2097]), .B(n6293), .Z(c[2097]) );
XNOR U10489 ( .A(a[2097]), .B(c2097), .Z(n6293) );
XOR U10490 ( .A(c2098), .B(n6294), .Z(c2099) );
ANDN U10491 ( .B(n6295), .A(n6296), .Z(n6294) );
XOR U10492 ( .A(c2098), .B(b[2098]), .Z(n6295) );
XNOR U10493 ( .A(b[2098]), .B(n6296), .Z(c[2098]) );
XNOR U10494 ( .A(a[2098]), .B(c2098), .Z(n6296) );
XOR U10495 ( .A(c2099), .B(n6297), .Z(c2100) );
ANDN U10496 ( .B(n6298), .A(n6299), .Z(n6297) );
XOR U10497 ( .A(c2099), .B(b[2099]), .Z(n6298) );
XNOR U10498 ( .A(b[2099]), .B(n6299), .Z(c[2099]) );
XNOR U10499 ( .A(a[2099]), .B(c2099), .Z(n6299) );
XOR U10500 ( .A(c2100), .B(n6300), .Z(c2101) );
ANDN U10501 ( .B(n6301), .A(n6302), .Z(n6300) );
XOR U10502 ( .A(c2100), .B(b[2100]), .Z(n6301) );
XNOR U10503 ( .A(b[2100]), .B(n6302), .Z(c[2100]) );
XNOR U10504 ( .A(a[2100]), .B(c2100), .Z(n6302) );
XOR U10505 ( .A(c2101), .B(n6303), .Z(c2102) );
ANDN U10506 ( .B(n6304), .A(n6305), .Z(n6303) );
XOR U10507 ( .A(c2101), .B(b[2101]), .Z(n6304) );
XNOR U10508 ( .A(b[2101]), .B(n6305), .Z(c[2101]) );
XNOR U10509 ( .A(a[2101]), .B(c2101), .Z(n6305) );
XOR U10510 ( .A(c2102), .B(n6306), .Z(c2103) );
ANDN U10511 ( .B(n6307), .A(n6308), .Z(n6306) );
XOR U10512 ( .A(c2102), .B(b[2102]), .Z(n6307) );
XNOR U10513 ( .A(b[2102]), .B(n6308), .Z(c[2102]) );
XNOR U10514 ( .A(a[2102]), .B(c2102), .Z(n6308) );
XOR U10515 ( .A(c2103), .B(n6309), .Z(c2104) );
ANDN U10516 ( .B(n6310), .A(n6311), .Z(n6309) );
XOR U10517 ( .A(c2103), .B(b[2103]), .Z(n6310) );
XNOR U10518 ( .A(b[2103]), .B(n6311), .Z(c[2103]) );
XNOR U10519 ( .A(a[2103]), .B(c2103), .Z(n6311) );
XOR U10520 ( .A(c2104), .B(n6312), .Z(c2105) );
ANDN U10521 ( .B(n6313), .A(n6314), .Z(n6312) );
XOR U10522 ( .A(c2104), .B(b[2104]), .Z(n6313) );
XNOR U10523 ( .A(b[2104]), .B(n6314), .Z(c[2104]) );
XNOR U10524 ( .A(a[2104]), .B(c2104), .Z(n6314) );
XOR U10525 ( .A(c2105), .B(n6315), .Z(c2106) );
ANDN U10526 ( .B(n6316), .A(n6317), .Z(n6315) );
XOR U10527 ( .A(c2105), .B(b[2105]), .Z(n6316) );
XNOR U10528 ( .A(b[2105]), .B(n6317), .Z(c[2105]) );
XNOR U10529 ( .A(a[2105]), .B(c2105), .Z(n6317) );
XOR U10530 ( .A(c2106), .B(n6318), .Z(c2107) );
ANDN U10531 ( .B(n6319), .A(n6320), .Z(n6318) );
XOR U10532 ( .A(c2106), .B(b[2106]), .Z(n6319) );
XNOR U10533 ( .A(b[2106]), .B(n6320), .Z(c[2106]) );
XNOR U10534 ( .A(a[2106]), .B(c2106), .Z(n6320) );
XOR U10535 ( .A(c2107), .B(n6321), .Z(c2108) );
ANDN U10536 ( .B(n6322), .A(n6323), .Z(n6321) );
XOR U10537 ( .A(c2107), .B(b[2107]), .Z(n6322) );
XNOR U10538 ( .A(b[2107]), .B(n6323), .Z(c[2107]) );
XNOR U10539 ( .A(a[2107]), .B(c2107), .Z(n6323) );
XOR U10540 ( .A(c2108), .B(n6324), .Z(c2109) );
ANDN U10541 ( .B(n6325), .A(n6326), .Z(n6324) );
XOR U10542 ( .A(c2108), .B(b[2108]), .Z(n6325) );
XNOR U10543 ( .A(b[2108]), .B(n6326), .Z(c[2108]) );
XNOR U10544 ( .A(a[2108]), .B(c2108), .Z(n6326) );
XOR U10545 ( .A(c2109), .B(n6327), .Z(c2110) );
ANDN U10546 ( .B(n6328), .A(n6329), .Z(n6327) );
XOR U10547 ( .A(c2109), .B(b[2109]), .Z(n6328) );
XNOR U10548 ( .A(b[2109]), .B(n6329), .Z(c[2109]) );
XNOR U10549 ( .A(a[2109]), .B(c2109), .Z(n6329) );
XOR U10550 ( .A(c2110), .B(n6330), .Z(c2111) );
ANDN U10551 ( .B(n6331), .A(n6332), .Z(n6330) );
XOR U10552 ( .A(c2110), .B(b[2110]), .Z(n6331) );
XNOR U10553 ( .A(b[2110]), .B(n6332), .Z(c[2110]) );
XNOR U10554 ( .A(a[2110]), .B(c2110), .Z(n6332) );
XOR U10555 ( .A(c2111), .B(n6333), .Z(c2112) );
ANDN U10556 ( .B(n6334), .A(n6335), .Z(n6333) );
XOR U10557 ( .A(c2111), .B(b[2111]), .Z(n6334) );
XNOR U10558 ( .A(b[2111]), .B(n6335), .Z(c[2111]) );
XNOR U10559 ( .A(a[2111]), .B(c2111), .Z(n6335) );
XOR U10560 ( .A(c2112), .B(n6336), .Z(c2113) );
ANDN U10561 ( .B(n6337), .A(n6338), .Z(n6336) );
XOR U10562 ( .A(c2112), .B(b[2112]), .Z(n6337) );
XNOR U10563 ( .A(b[2112]), .B(n6338), .Z(c[2112]) );
XNOR U10564 ( .A(a[2112]), .B(c2112), .Z(n6338) );
XOR U10565 ( .A(c2113), .B(n6339), .Z(c2114) );
ANDN U10566 ( .B(n6340), .A(n6341), .Z(n6339) );
XOR U10567 ( .A(c2113), .B(b[2113]), .Z(n6340) );
XNOR U10568 ( .A(b[2113]), .B(n6341), .Z(c[2113]) );
XNOR U10569 ( .A(a[2113]), .B(c2113), .Z(n6341) );
XOR U10570 ( .A(c2114), .B(n6342), .Z(c2115) );
ANDN U10571 ( .B(n6343), .A(n6344), .Z(n6342) );
XOR U10572 ( .A(c2114), .B(b[2114]), .Z(n6343) );
XNOR U10573 ( .A(b[2114]), .B(n6344), .Z(c[2114]) );
XNOR U10574 ( .A(a[2114]), .B(c2114), .Z(n6344) );
XOR U10575 ( .A(c2115), .B(n6345), .Z(c2116) );
ANDN U10576 ( .B(n6346), .A(n6347), .Z(n6345) );
XOR U10577 ( .A(c2115), .B(b[2115]), .Z(n6346) );
XNOR U10578 ( .A(b[2115]), .B(n6347), .Z(c[2115]) );
XNOR U10579 ( .A(a[2115]), .B(c2115), .Z(n6347) );
XOR U10580 ( .A(c2116), .B(n6348), .Z(c2117) );
ANDN U10581 ( .B(n6349), .A(n6350), .Z(n6348) );
XOR U10582 ( .A(c2116), .B(b[2116]), .Z(n6349) );
XNOR U10583 ( .A(b[2116]), .B(n6350), .Z(c[2116]) );
XNOR U10584 ( .A(a[2116]), .B(c2116), .Z(n6350) );
XOR U10585 ( .A(c2117), .B(n6351), .Z(c2118) );
ANDN U10586 ( .B(n6352), .A(n6353), .Z(n6351) );
XOR U10587 ( .A(c2117), .B(b[2117]), .Z(n6352) );
XNOR U10588 ( .A(b[2117]), .B(n6353), .Z(c[2117]) );
XNOR U10589 ( .A(a[2117]), .B(c2117), .Z(n6353) );
XOR U10590 ( .A(c2118), .B(n6354), .Z(c2119) );
ANDN U10591 ( .B(n6355), .A(n6356), .Z(n6354) );
XOR U10592 ( .A(c2118), .B(b[2118]), .Z(n6355) );
XNOR U10593 ( .A(b[2118]), .B(n6356), .Z(c[2118]) );
XNOR U10594 ( .A(a[2118]), .B(c2118), .Z(n6356) );
XOR U10595 ( .A(c2119), .B(n6357), .Z(c2120) );
ANDN U10596 ( .B(n6358), .A(n6359), .Z(n6357) );
XOR U10597 ( .A(c2119), .B(b[2119]), .Z(n6358) );
XNOR U10598 ( .A(b[2119]), .B(n6359), .Z(c[2119]) );
XNOR U10599 ( .A(a[2119]), .B(c2119), .Z(n6359) );
XOR U10600 ( .A(c2120), .B(n6360), .Z(c2121) );
ANDN U10601 ( .B(n6361), .A(n6362), .Z(n6360) );
XOR U10602 ( .A(c2120), .B(b[2120]), .Z(n6361) );
XNOR U10603 ( .A(b[2120]), .B(n6362), .Z(c[2120]) );
XNOR U10604 ( .A(a[2120]), .B(c2120), .Z(n6362) );
XOR U10605 ( .A(c2121), .B(n6363), .Z(c2122) );
ANDN U10606 ( .B(n6364), .A(n6365), .Z(n6363) );
XOR U10607 ( .A(c2121), .B(b[2121]), .Z(n6364) );
XNOR U10608 ( .A(b[2121]), .B(n6365), .Z(c[2121]) );
XNOR U10609 ( .A(a[2121]), .B(c2121), .Z(n6365) );
XOR U10610 ( .A(c2122), .B(n6366), .Z(c2123) );
ANDN U10611 ( .B(n6367), .A(n6368), .Z(n6366) );
XOR U10612 ( .A(c2122), .B(b[2122]), .Z(n6367) );
XNOR U10613 ( .A(b[2122]), .B(n6368), .Z(c[2122]) );
XNOR U10614 ( .A(a[2122]), .B(c2122), .Z(n6368) );
XOR U10615 ( .A(c2123), .B(n6369), .Z(c2124) );
ANDN U10616 ( .B(n6370), .A(n6371), .Z(n6369) );
XOR U10617 ( .A(c2123), .B(b[2123]), .Z(n6370) );
XNOR U10618 ( .A(b[2123]), .B(n6371), .Z(c[2123]) );
XNOR U10619 ( .A(a[2123]), .B(c2123), .Z(n6371) );
XOR U10620 ( .A(c2124), .B(n6372), .Z(c2125) );
ANDN U10621 ( .B(n6373), .A(n6374), .Z(n6372) );
XOR U10622 ( .A(c2124), .B(b[2124]), .Z(n6373) );
XNOR U10623 ( .A(b[2124]), .B(n6374), .Z(c[2124]) );
XNOR U10624 ( .A(a[2124]), .B(c2124), .Z(n6374) );
XOR U10625 ( .A(c2125), .B(n6375), .Z(c2126) );
ANDN U10626 ( .B(n6376), .A(n6377), .Z(n6375) );
XOR U10627 ( .A(c2125), .B(b[2125]), .Z(n6376) );
XNOR U10628 ( .A(b[2125]), .B(n6377), .Z(c[2125]) );
XNOR U10629 ( .A(a[2125]), .B(c2125), .Z(n6377) );
XOR U10630 ( .A(c2126), .B(n6378), .Z(c2127) );
ANDN U10631 ( .B(n6379), .A(n6380), .Z(n6378) );
XOR U10632 ( .A(c2126), .B(b[2126]), .Z(n6379) );
XNOR U10633 ( .A(b[2126]), .B(n6380), .Z(c[2126]) );
XNOR U10634 ( .A(a[2126]), .B(c2126), .Z(n6380) );
XOR U10635 ( .A(c2127), .B(n6381), .Z(c2128) );
ANDN U10636 ( .B(n6382), .A(n6383), .Z(n6381) );
XOR U10637 ( .A(c2127), .B(b[2127]), .Z(n6382) );
XNOR U10638 ( .A(b[2127]), .B(n6383), .Z(c[2127]) );
XNOR U10639 ( .A(a[2127]), .B(c2127), .Z(n6383) );
XOR U10640 ( .A(c2128), .B(n6384), .Z(c2129) );
ANDN U10641 ( .B(n6385), .A(n6386), .Z(n6384) );
XOR U10642 ( .A(c2128), .B(b[2128]), .Z(n6385) );
XNOR U10643 ( .A(b[2128]), .B(n6386), .Z(c[2128]) );
XNOR U10644 ( .A(a[2128]), .B(c2128), .Z(n6386) );
XOR U10645 ( .A(c2129), .B(n6387), .Z(c2130) );
ANDN U10646 ( .B(n6388), .A(n6389), .Z(n6387) );
XOR U10647 ( .A(c2129), .B(b[2129]), .Z(n6388) );
XNOR U10648 ( .A(b[2129]), .B(n6389), .Z(c[2129]) );
XNOR U10649 ( .A(a[2129]), .B(c2129), .Z(n6389) );
XOR U10650 ( .A(c2130), .B(n6390), .Z(c2131) );
ANDN U10651 ( .B(n6391), .A(n6392), .Z(n6390) );
XOR U10652 ( .A(c2130), .B(b[2130]), .Z(n6391) );
XNOR U10653 ( .A(b[2130]), .B(n6392), .Z(c[2130]) );
XNOR U10654 ( .A(a[2130]), .B(c2130), .Z(n6392) );
XOR U10655 ( .A(c2131), .B(n6393), .Z(c2132) );
ANDN U10656 ( .B(n6394), .A(n6395), .Z(n6393) );
XOR U10657 ( .A(c2131), .B(b[2131]), .Z(n6394) );
XNOR U10658 ( .A(b[2131]), .B(n6395), .Z(c[2131]) );
XNOR U10659 ( .A(a[2131]), .B(c2131), .Z(n6395) );
XOR U10660 ( .A(c2132), .B(n6396), .Z(c2133) );
ANDN U10661 ( .B(n6397), .A(n6398), .Z(n6396) );
XOR U10662 ( .A(c2132), .B(b[2132]), .Z(n6397) );
XNOR U10663 ( .A(b[2132]), .B(n6398), .Z(c[2132]) );
XNOR U10664 ( .A(a[2132]), .B(c2132), .Z(n6398) );
XOR U10665 ( .A(c2133), .B(n6399), .Z(c2134) );
ANDN U10666 ( .B(n6400), .A(n6401), .Z(n6399) );
XOR U10667 ( .A(c2133), .B(b[2133]), .Z(n6400) );
XNOR U10668 ( .A(b[2133]), .B(n6401), .Z(c[2133]) );
XNOR U10669 ( .A(a[2133]), .B(c2133), .Z(n6401) );
XOR U10670 ( .A(c2134), .B(n6402), .Z(c2135) );
ANDN U10671 ( .B(n6403), .A(n6404), .Z(n6402) );
XOR U10672 ( .A(c2134), .B(b[2134]), .Z(n6403) );
XNOR U10673 ( .A(b[2134]), .B(n6404), .Z(c[2134]) );
XNOR U10674 ( .A(a[2134]), .B(c2134), .Z(n6404) );
XOR U10675 ( .A(c2135), .B(n6405), .Z(c2136) );
ANDN U10676 ( .B(n6406), .A(n6407), .Z(n6405) );
XOR U10677 ( .A(c2135), .B(b[2135]), .Z(n6406) );
XNOR U10678 ( .A(b[2135]), .B(n6407), .Z(c[2135]) );
XNOR U10679 ( .A(a[2135]), .B(c2135), .Z(n6407) );
XOR U10680 ( .A(c2136), .B(n6408), .Z(c2137) );
ANDN U10681 ( .B(n6409), .A(n6410), .Z(n6408) );
XOR U10682 ( .A(c2136), .B(b[2136]), .Z(n6409) );
XNOR U10683 ( .A(b[2136]), .B(n6410), .Z(c[2136]) );
XNOR U10684 ( .A(a[2136]), .B(c2136), .Z(n6410) );
XOR U10685 ( .A(c2137), .B(n6411), .Z(c2138) );
ANDN U10686 ( .B(n6412), .A(n6413), .Z(n6411) );
XOR U10687 ( .A(c2137), .B(b[2137]), .Z(n6412) );
XNOR U10688 ( .A(b[2137]), .B(n6413), .Z(c[2137]) );
XNOR U10689 ( .A(a[2137]), .B(c2137), .Z(n6413) );
XOR U10690 ( .A(c2138), .B(n6414), .Z(c2139) );
ANDN U10691 ( .B(n6415), .A(n6416), .Z(n6414) );
XOR U10692 ( .A(c2138), .B(b[2138]), .Z(n6415) );
XNOR U10693 ( .A(b[2138]), .B(n6416), .Z(c[2138]) );
XNOR U10694 ( .A(a[2138]), .B(c2138), .Z(n6416) );
XOR U10695 ( .A(c2139), .B(n6417), .Z(c2140) );
ANDN U10696 ( .B(n6418), .A(n6419), .Z(n6417) );
XOR U10697 ( .A(c2139), .B(b[2139]), .Z(n6418) );
XNOR U10698 ( .A(b[2139]), .B(n6419), .Z(c[2139]) );
XNOR U10699 ( .A(a[2139]), .B(c2139), .Z(n6419) );
XOR U10700 ( .A(c2140), .B(n6420), .Z(c2141) );
ANDN U10701 ( .B(n6421), .A(n6422), .Z(n6420) );
XOR U10702 ( .A(c2140), .B(b[2140]), .Z(n6421) );
XNOR U10703 ( .A(b[2140]), .B(n6422), .Z(c[2140]) );
XNOR U10704 ( .A(a[2140]), .B(c2140), .Z(n6422) );
XOR U10705 ( .A(c2141), .B(n6423), .Z(c2142) );
ANDN U10706 ( .B(n6424), .A(n6425), .Z(n6423) );
XOR U10707 ( .A(c2141), .B(b[2141]), .Z(n6424) );
XNOR U10708 ( .A(b[2141]), .B(n6425), .Z(c[2141]) );
XNOR U10709 ( .A(a[2141]), .B(c2141), .Z(n6425) );
XOR U10710 ( .A(c2142), .B(n6426), .Z(c2143) );
ANDN U10711 ( .B(n6427), .A(n6428), .Z(n6426) );
XOR U10712 ( .A(c2142), .B(b[2142]), .Z(n6427) );
XNOR U10713 ( .A(b[2142]), .B(n6428), .Z(c[2142]) );
XNOR U10714 ( .A(a[2142]), .B(c2142), .Z(n6428) );
XOR U10715 ( .A(c2143), .B(n6429), .Z(c2144) );
ANDN U10716 ( .B(n6430), .A(n6431), .Z(n6429) );
XOR U10717 ( .A(c2143), .B(b[2143]), .Z(n6430) );
XNOR U10718 ( .A(b[2143]), .B(n6431), .Z(c[2143]) );
XNOR U10719 ( .A(a[2143]), .B(c2143), .Z(n6431) );
XOR U10720 ( .A(c2144), .B(n6432), .Z(c2145) );
ANDN U10721 ( .B(n6433), .A(n6434), .Z(n6432) );
XOR U10722 ( .A(c2144), .B(b[2144]), .Z(n6433) );
XNOR U10723 ( .A(b[2144]), .B(n6434), .Z(c[2144]) );
XNOR U10724 ( .A(a[2144]), .B(c2144), .Z(n6434) );
XOR U10725 ( .A(c2145), .B(n6435), .Z(c2146) );
ANDN U10726 ( .B(n6436), .A(n6437), .Z(n6435) );
XOR U10727 ( .A(c2145), .B(b[2145]), .Z(n6436) );
XNOR U10728 ( .A(b[2145]), .B(n6437), .Z(c[2145]) );
XNOR U10729 ( .A(a[2145]), .B(c2145), .Z(n6437) );
XOR U10730 ( .A(c2146), .B(n6438), .Z(c2147) );
ANDN U10731 ( .B(n6439), .A(n6440), .Z(n6438) );
XOR U10732 ( .A(c2146), .B(b[2146]), .Z(n6439) );
XNOR U10733 ( .A(b[2146]), .B(n6440), .Z(c[2146]) );
XNOR U10734 ( .A(a[2146]), .B(c2146), .Z(n6440) );
XOR U10735 ( .A(c2147), .B(n6441), .Z(c2148) );
ANDN U10736 ( .B(n6442), .A(n6443), .Z(n6441) );
XOR U10737 ( .A(c2147), .B(b[2147]), .Z(n6442) );
XNOR U10738 ( .A(b[2147]), .B(n6443), .Z(c[2147]) );
XNOR U10739 ( .A(a[2147]), .B(c2147), .Z(n6443) );
XOR U10740 ( .A(c2148), .B(n6444), .Z(c2149) );
ANDN U10741 ( .B(n6445), .A(n6446), .Z(n6444) );
XOR U10742 ( .A(c2148), .B(b[2148]), .Z(n6445) );
XNOR U10743 ( .A(b[2148]), .B(n6446), .Z(c[2148]) );
XNOR U10744 ( .A(a[2148]), .B(c2148), .Z(n6446) );
XOR U10745 ( .A(c2149), .B(n6447), .Z(c2150) );
ANDN U10746 ( .B(n6448), .A(n6449), .Z(n6447) );
XOR U10747 ( .A(c2149), .B(b[2149]), .Z(n6448) );
XNOR U10748 ( .A(b[2149]), .B(n6449), .Z(c[2149]) );
XNOR U10749 ( .A(a[2149]), .B(c2149), .Z(n6449) );
XOR U10750 ( .A(c2150), .B(n6450), .Z(c2151) );
ANDN U10751 ( .B(n6451), .A(n6452), .Z(n6450) );
XOR U10752 ( .A(c2150), .B(b[2150]), .Z(n6451) );
XNOR U10753 ( .A(b[2150]), .B(n6452), .Z(c[2150]) );
XNOR U10754 ( .A(a[2150]), .B(c2150), .Z(n6452) );
XOR U10755 ( .A(c2151), .B(n6453), .Z(c2152) );
ANDN U10756 ( .B(n6454), .A(n6455), .Z(n6453) );
XOR U10757 ( .A(c2151), .B(b[2151]), .Z(n6454) );
XNOR U10758 ( .A(b[2151]), .B(n6455), .Z(c[2151]) );
XNOR U10759 ( .A(a[2151]), .B(c2151), .Z(n6455) );
XOR U10760 ( .A(c2152), .B(n6456), .Z(c2153) );
ANDN U10761 ( .B(n6457), .A(n6458), .Z(n6456) );
XOR U10762 ( .A(c2152), .B(b[2152]), .Z(n6457) );
XNOR U10763 ( .A(b[2152]), .B(n6458), .Z(c[2152]) );
XNOR U10764 ( .A(a[2152]), .B(c2152), .Z(n6458) );
XOR U10765 ( .A(c2153), .B(n6459), .Z(c2154) );
ANDN U10766 ( .B(n6460), .A(n6461), .Z(n6459) );
XOR U10767 ( .A(c2153), .B(b[2153]), .Z(n6460) );
XNOR U10768 ( .A(b[2153]), .B(n6461), .Z(c[2153]) );
XNOR U10769 ( .A(a[2153]), .B(c2153), .Z(n6461) );
XOR U10770 ( .A(c2154), .B(n6462), .Z(c2155) );
ANDN U10771 ( .B(n6463), .A(n6464), .Z(n6462) );
XOR U10772 ( .A(c2154), .B(b[2154]), .Z(n6463) );
XNOR U10773 ( .A(b[2154]), .B(n6464), .Z(c[2154]) );
XNOR U10774 ( .A(a[2154]), .B(c2154), .Z(n6464) );
XOR U10775 ( .A(c2155), .B(n6465), .Z(c2156) );
ANDN U10776 ( .B(n6466), .A(n6467), .Z(n6465) );
XOR U10777 ( .A(c2155), .B(b[2155]), .Z(n6466) );
XNOR U10778 ( .A(b[2155]), .B(n6467), .Z(c[2155]) );
XNOR U10779 ( .A(a[2155]), .B(c2155), .Z(n6467) );
XOR U10780 ( .A(c2156), .B(n6468), .Z(c2157) );
ANDN U10781 ( .B(n6469), .A(n6470), .Z(n6468) );
XOR U10782 ( .A(c2156), .B(b[2156]), .Z(n6469) );
XNOR U10783 ( .A(b[2156]), .B(n6470), .Z(c[2156]) );
XNOR U10784 ( .A(a[2156]), .B(c2156), .Z(n6470) );
XOR U10785 ( .A(c2157), .B(n6471), .Z(c2158) );
ANDN U10786 ( .B(n6472), .A(n6473), .Z(n6471) );
XOR U10787 ( .A(c2157), .B(b[2157]), .Z(n6472) );
XNOR U10788 ( .A(b[2157]), .B(n6473), .Z(c[2157]) );
XNOR U10789 ( .A(a[2157]), .B(c2157), .Z(n6473) );
XOR U10790 ( .A(c2158), .B(n6474), .Z(c2159) );
ANDN U10791 ( .B(n6475), .A(n6476), .Z(n6474) );
XOR U10792 ( .A(c2158), .B(b[2158]), .Z(n6475) );
XNOR U10793 ( .A(b[2158]), .B(n6476), .Z(c[2158]) );
XNOR U10794 ( .A(a[2158]), .B(c2158), .Z(n6476) );
XOR U10795 ( .A(c2159), .B(n6477), .Z(c2160) );
ANDN U10796 ( .B(n6478), .A(n6479), .Z(n6477) );
XOR U10797 ( .A(c2159), .B(b[2159]), .Z(n6478) );
XNOR U10798 ( .A(b[2159]), .B(n6479), .Z(c[2159]) );
XNOR U10799 ( .A(a[2159]), .B(c2159), .Z(n6479) );
XOR U10800 ( .A(c2160), .B(n6480), .Z(c2161) );
ANDN U10801 ( .B(n6481), .A(n6482), .Z(n6480) );
XOR U10802 ( .A(c2160), .B(b[2160]), .Z(n6481) );
XNOR U10803 ( .A(b[2160]), .B(n6482), .Z(c[2160]) );
XNOR U10804 ( .A(a[2160]), .B(c2160), .Z(n6482) );
XOR U10805 ( .A(c2161), .B(n6483), .Z(c2162) );
ANDN U10806 ( .B(n6484), .A(n6485), .Z(n6483) );
XOR U10807 ( .A(c2161), .B(b[2161]), .Z(n6484) );
XNOR U10808 ( .A(b[2161]), .B(n6485), .Z(c[2161]) );
XNOR U10809 ( .A(a[2161]), .B(c2161), .Z(n6485) );
XOR U10810 ( .A(c2162), .B(n6486), .Z(c2163) );
ANDN U10811 ( .B(n6487), .A(n6488), .Z(n6486) );
XOR U10812 ( .A(c2162), .B(b[2162]), .Z(n6487) );
XNOR U10813 ( .A(b[2162]), .B(n6488), .Z(c[2162]) );
XNOR U10814 ( .A(a[2162]), .B(c2162), .Z(n6488) );
XOR U10815 ( .A(c2163), .B(n6489), .Z(c2164) );
ANDN U10816 ( .B(n6490), .A(n6491), .Z(n6489) );
XOR U10817 ( .A(c2163), .B(b[2163]), .Z(n6490) );
XNOR U10818 ( .A(b[2163]), .B(n6491), .Z(c[2163]) );
XNOR U10819 ( .A(a[2163]), .B(c2163), .Z(n6491) );
XOR U10820 ( .A(c2164), .B(n6492), .Z(c2165) );
ANDN U10821 ( .B(n6493), .A(n6494), .Z(n6492) );
XOR U10822 ( .A(c2164), .B(b[2164]), .Z(n6493) );
XNOR U10823 ( .A(b[2164]), .B(n6494), .Z(c[2164]) );
XNOR U10824 ( .A(a[2164]), .B(c2164), .Z(n6494) );
XOR U10825 ( .A(c2165), .B(n6495), .Z(c2166) );
ANDN U10826 ( .B(n6496), .A(n6497), .Z(n6495) );
XOR U10827 ( .A(c2165), .B(b[2165]), .Z(n6496) );
XNOR U10828 ( .A(b[2165]), .B(n6497), .Z(c[2165]) );
XNOR U10829 ( .A(a[2165]), .B(c2165), .Z(n6497) );
XOR U10830 ( .A(c2166), .B(n6498), .Z(c2167) );
ANDN U10831 ( .B(n6499), .A(n6500), .Z(n6498) );
XOR U10832 ( .A(c2166), .B(b[2166]), .Z(n6499) );
XNOR U10833 ( .A(b[2166]), .B(n6500), .Z(c[2166]) );
XNOR U10834 ( .A(a[2166]), .B(c2166), .Z(n6500) );
XOR U10835 ( .A(c2167), .B(n6501), .Z(c2168) );
ANDN U10836 ( .B(n6502), .A(n6503), .Z(n6501) );
XOR U10837 ( .A(c2167), .B(b[2167]), .Z(n6502) );
XNOR U10838 ( .A(b[2167]), .B(n6503), .Z(c[2167]) );
XNOR U10839 ( .A(a[2167]), .B(c2167), .Z(n6503) );
XOR U10840 ( .A(c2168), .B(n6504), .Z(c2169) );
ANDN U10841 ( .B(n6505), .A(n6506), .Z(n6504) );
XOR U10842 ( .A(c2168), .B(b[2168]), .Z(n6505) );
XNOR U10843 ( .A(b[2168]), .B(n6506), .Z(c[2168]) );
XNOR U10844 ( .A(a[2168]), .B(c2168), .Z(n6506) );
XOR U10845 ( .A(c2169), .B(n6507), .Z(c2170) );
ANDN U10846 ( .B(n6508), .A(n6509), .Z(n6507) );
XOR U10847 ( .A(c2169), .B(b[2169]), .Z(n6508) );
XNOR U10848 ( .A(b[2169]), .B(n6509), .Z(c[2169]) );
XNOR U10849 ( .A(a[2169]), .B(c2169), .Z(n6509) );
XOR U10850 ( .A(c2170), .B(n6510), .Z(c2171) );
ANDN U10851 ( .B(n6511), .A(n6512), .Z(n6510) );
XOR U10852 ( .A(c2170), .B(b[2170]), .Z(n6511) );
XNOR U10853 ( .A(b[2170]), .B(n6512), .Z(c[2170]) );
XNOR U10854 ( .A(a[2170]), .B(c2170), .Z(n6512) );
XOR U10855 ( .A(c2171), .B(n6513), .Z(c2172) );
ANDN U10856 ( .B(n6514), .A(n6515), .Z(n6513) );
XOR U10857 ( .A(c2171), .B(b[2171]), .Z(n6514) );
XNOR U10858 ( .A(b[2171]), .B(n6515), .Z(c[2171]) );
XNOR U10859 ( .A(a[2171]), .B(c2171), .Z(n6515) );
XOR U10860 ( .A(c2172), .B(n6516), .Z(c2173) );
ANDN U10861 ( .B(n6517), .A(n6518), .Z(n6516) );
XOR U10862 ( .A(c2172), .B(b[2172]), .Z(n6517) );
XNOR U10863 ( .A(b[2172]), .B(n6518), .Z(c[2172]) );
XNOR U10864 ( .A(a[2172]), .B(c2172), .Z(n6518) );
XOR U10865 ( .A(c2173), .B(n6519), .Z(c2174) );
ANDN U10866 ( .B(n6520), .A(n6521), .Z(n6519) );
XOR U10867 ( .A(c2173), .B(b[2173]), .Z(n6520) );
XNOR U10868 ( .A(b[2173]), .B(n6521), .Z(c[2173]) );
XNOR U10869 ( .A(a[2173]), .B(c2173), .Z(n6521) );
XOR U10870 ( .A(c2174), .B(n6522), .Z(c2175) );
ANDN U10871 ( .B(n6523), .A(n6524), .Z(n6522) );
XOR U10872 ( .A(c2174), .B(b[2174]), .Z(n6523) );
XNOR U10873 ( .A(b[2174]), .B(n6524), .Z(c[2174]) );
XNOR U10874 ( .A(a[2174]), .B(c2174), .Z(n6524) );
XOR U10875 ( .A(c2175), .B(n6525), .Z(c2176) );
ANDN U10876 ( .B(n6526), .A(n6527), .Z(n6525) );
XOR U10877 ( .A(c2175), .B(b[2175]), .Z(n6526) );
XNOR U10878 ( .A(b[2175]), .B(n6527), .Z(c[2175]) );
XNOR U10879 ( .A(a[2175]), .B(c2175), .Z(n6527) );
XOR U10880 ( .A(c2176), .B(n6528), .Z(c2177) );
ANDN U10881 ( .B(n6529), .A(n6530), .Z(n6528) );
XOR U10882 ( .A(c2176), .B(b[2176]), .Z(n6529) );
XNOR U10883 ( .A(b[2176]), .B(n6530), .Z(c[2176]) );
XNOR U10884 ( .A(a[2176]), .B(c2176), .Z(n6530) );
XOR U10885 ( .A(c2177), .B(n6531), .Z(c2178) );
ANDN U10886 ( .B(n6532), .A(n6533), .Z(n6531) );
XOR U10887 ( .A(c2177), .B(b[2177]), .Z(n6532) );
XNOR U10888 ( .A(b[2177]), .B(n6533), .Z(c[2177]) );
XNOR U10889 ( .A(a[2177]), .B(c2177), .Z(n6533) );
XOR U10890 ( .A(c2178), .B(n6534), .Z(c2179) );
ANDN U10891 ( .B(n6535), .A(n6536), .Z(n6534) );
XOR U10892 ( .A(c2178), .B(b[2178]), .Z(n6535) );
XNOR U10893 ( .A(b[2178]), .B(n6536), .Z(c[2178]) );
XNOR U10894 ( .A(a[2178]), .B(c2178), .Z(n6536) );
XOR U10895 ( .A(c2179), .B(n6537), .Z(c2180) );
ANDN U10896 ( .B(n6538), .A(n6539), .Z(n6537) );
XOR U10897 ( .A(c2179), .B(b[2179]), .Z(n6538) );
XNOR U10898 ( .A(b[2179]), .B(n6539), .Z(c[2179]) );
XNOR U10899 ( .A(a[2179]), .B(c2179), .Z(n6539) );
XOR U10900 ( .A(c2180), .B(n6540), .Z(c2181) );
ANDN U10901 ( .B(n6541), .A(n6542), .Z(n6540) );
XOR U10902 ( .A(c2180), .B(b[2180]), .Z(n6541) );
XNOR U10903 ( .A(b[2180]), .B(n6542), .Z(c[2180]) );
XNOR U10904 ( .A(a[2180]), .B(c2180), .Z(n6542) );
XOR U10905 ( .A(c2181), .B(n6543), .Z(c2182) );
ANDN U10906 ( .B(n6544), .A(n6545), .Z(n6543) );
XOR U10907 ( .A(c2181), .B(b[2181]), .Z(n6544) );
XNOR U10908 ( .A(b[2181]), .B(n6545), .Z(c[2181]) );
XNOR U10909 ( .A(a[2181]), .B(c2181), .Z(n6545) );
XOR U10910 ( .A(c2182), .B(n6546), .Z(c2183) );
ANDN U10911 ( .B(n6547), .A(n6548), .Z(n6546) );
XOR U10912 ( .A(c2182), .B(b[2182]), .Z(n6547) );
XNOR U10913 ( .A(b[2182]), .B(n6548), .Z(c[2182]) );
XNOR U10914 ( .A(a[2182]), .B(c2182), .Z(n6548) );
XOR U10915 ( .A(c2183), .B(n6549), .Z(c2184) );
ANDN U10916 ( .B(n6550), .A(n6551), .Z(n6549) );
XOR U10917 ( .A(c2183), .B(b[2183]), .Z(n6550) );
XNOR U10918 ( .A(b[2183]), .B(n6551), .Z(c[2183]) );
XNOR U10919 ( .A(a[2183]), .B(c2183), .Z(n6551) );
XOR U10920 ( .A(c2184), .B(n6552), .Z(c2185) );
ANDN U10921 ( .B(n6553), .A(n6554), .Z(n6552) );
XOR U10922 ( .A(c2184), .B(b[2184]), .Z(n6553) );
XNOR U10923 ( .A(b[2184]), .B(n6554), .Z(c[2184]) );
XNOR U10924 ( .A(a[2184]), .B(c2184), .Z(n6554) );
XOR U10925 ( .A(c2185), .B(n6555), .Z(c2186) );
ANDN U10926 ( .B(n6556), .A(n6557), .Z(n6555) );
XOR U10927 ( .A(c2185), .B(b[2185]), .Z(n6556) );
XNOR U10928 ( .A(b[2185]), .B(n6557), .Z(c[2185]) );
XNOR U10929 ( .A(a[2185]), .B(c2185), .Z(n6557) );
XOR U10930 ( .A(c2186), .B(n6558), .Z(c2187) );
ANDN U10931 ( .B(n6559), .A(n6560), .Z(n6558) );
XOR U10932 ( .A(c2186), .B(b[2186]), .Z(n6559) );
XNOR U10933 ( .A(b[2186]), .B(n6560), .Z(c[2186]) );
XNOR U10934 ( .A(a[2186]), .B(c2186), .Z(n6560) );
XOR U10935 ( .A(c2187), .B(n6561), .Z(c2188) );
ANDN U10936 ( .B(n6562), .A(n6563), .Z(n6561) );
XOR U10937 ( .A(c2187), .B(b[2187]), .Z(n6562) );
XNOR U10938 ( .A(b[2187]), .B(n6563), .Z(c[2187]) );
XNOR U10939 ( .A(a[2187]), .B(c2187), .Z(n6563) );
XOR U10940 ( .A(c2188), .B(n6564), .Z(c2189) );
ANDN U10941 ( .B(n6565), .A(n6566), .Z(n6564) );
XOR U10942 ( .A(c2188), .B(b[2188]), .Z(n6565) );
XNOR U10943 ( .A(b[2188]), .B(n6566), .Z(c[2188]) );
XNOR U10944 ( .A(a[2188]), .B(c2188), .Z(n6566) );
XOR U10945 ( .A(c2189), .B(n6567), .Z(c2190) );
ANDN U10946 ( .B(n6568), .A(n6569), .Z(n6567) );
XOR U10947 ( .A(c2189), .B(b[2189]), .Z(n6568) );
XNOR U10948 ( .A(b[2189]), .B(n6569), .Z(c[2189]) );
XNOR U10949 ( .A(a[2189]), .B(c2189), .Z(n6569) );
XOR U10950 ( .A(c2190), .B(n6570), .Z(c2191) );
ANDN U10951 ( .B(n6571), .A(n6572), .Z(n6570) );
XOR U10952 ( .A(c2190), .B(b[2190]), .Z(n6571) );
XNOR U10953 ( .A(b[2190]), .B(n6572), .Z(c[2190]) );
XNOR U10954 ( .A(a[2190]), .B(c2190), .Z(n6572) );
XOR U10955 ( .A(c2191), .B(n6573), .Z(c2192) );
ANDN U10956 ( .B(n6574), .A(n6575), .Z(n6573) );
XOR U10957 ( .A(c2191), .B(b[2191]), .Z(n6574) );
XNOR U10958 ( .A(b[2191]), .B(n6575), .Z(c[2191]) );
XNOR U10959 ( .A(a[2191]), .B(c2191), .Z(n6575) );
XOR U10960 ( .A(c2192), .B(n6576), .Z(c2193) );
ANDN U10961 ( .B(n6577), .A(n6578), .Z(n6576) );
XOR U10962 ( .A(c2192), .B(b[2192]), .Z(n6577) );
XNOR U10963 ( .A(b[2192]), .B(n6578), .Z(c[2192]) );
XNOR U10964 ( .A(a[2192]), .B(c2192), .Z(n6578) );
XOR U10965 ( .A(c2193), .B(n6579), .Z(c2194) );
ANDN U10966 ( .B(n6580), .A(n6581), .Z(n6579) );
XOR U10967 ( .A(c2193), .B(b[2193]), .Z(n6580) );
XNOR U10968 ( .A(b[2193]), .B(n6581), .Z(c[2193]) );
XNOR U10969 ( .A(a[2193]), .B(c2193), .Z(n6581) );
XOR U10970 ( .A(c2194), .B(n6582), .Z(c2195) );
ANDN U10971 ( .B(n6583), .A(n6584), .Z(n6582) );
XOR U10972 ( .A(c2194), .B(b[2194]), .Z(n6583) );
XNOR U10973 ( .A(b[2194]), .B(n6584), .Z(c[2194]) );
XNOR U10974 ( .A(a[2194]), .B(c2194), .Z(n6584) );
XOR U10975 ( .A(c2195), .B(n6585), .Z(c2196) );
ANDN U10976 ( .B(n6586), .A(n6587), .Z(n6585) );
XOR U10977 ( .A(c2195), .B(b[2195]), .Z(n6586) );
XNOR U10978 ( .A(b[2195]), .B(n6587), .Z(c[2195]) );
XNOR U10979 ( .A(a[2195]), .B(c2195), .Z(n6587) );
XOR U10980 ( .A(c2196), .B(n6588), .Z(c2197) );
ANDN U10981 ( .B(n6589), .A(n6590), .Z(n6588) );
XOR U10982 ( .A(c2196), .B(b[2196]), .Z(n6589) );
XNOR U10983 ( .A(b[2196]), .B(n6590), .Z(c[2196]) );
XNOR U10984 ( .A(a[2196]), .B(c2196), .Z(n6590) );
XOR U10985 ( .A(c2197), .B(n6591), .Z(c2198) );
ANDN U10986 ( .B(n6592), .A(n6593), .Z(n6591) );
XOR U10987 ( .A(c2197), .B(b[2197]), .Z(n6592) );
XNOR U10988 ( .A(b[2197]), .B(n6593), .Z(c[2197]) );
XNOR U10989 ( .A(a[2197]), .B(c2197), .Z(n6593) );
XOR U10990 ( .A(c2198), .B(n6594), .Z(c2199) );
ANDN U10991 ( .B(n6595), .A(n6596), .Z(n6594) );
XOR U10992 ( .A(c2198), .B(b[2198]), .Z(n6595) );
XNOR U10993 ( .A(b[2198]), .B(n6596), .Z(c[2198]) );
XNOR U10994 ( .A(a[2198]), .B(c2198), .Z(n6596) );
XOR U10995 ( .A(c2199), .B(n6597), .Z(c2200) );
ANDN U10996 ( .B(n6598), .A(n6599), .Z(n6597) );
XOR U10997 ( .A(c2199), .B(b[2199]), .Z(n6598) );
XNOR U10998 ( .A(b[2199]), .B(n6599), .Z(c[2199]) );
XNOR U10999 ( .A(a[2199]), .B(c2199), .Z(n6599) );
XOR U11000 ( .A(c2200), .B(n6600), .Z(c2201) );
ANDN U11001 ( .B(n6601), .A(n6602), .Z(n6600) );
XOR U11002 ( .A(c2200), .B(b[2200]), .Z(n6601) );
XNOR U11003 ( .A(b[2200]), .B(n6602), .Z(c[2200]) );
XNOR U11004 ( .A(a[2200]), .B(c2200), .Z(n6602) );
XOR U11005 ( .A(c2201), .B(n6603), .Z(c2202) );
ANDN U11006 ( .B(n6604), .A(n6605), .Z(n6603) );
XOR U11007 ( .A(c2201), .B(b[2201]), .Z(n6604) );
XNOR U11008 ( .A(b[2201]), .B(n6605), .Z(c[2201]) );
XNOR U11009 ( .A(a[2201]), .B(c2201), .Z(n6605) );
XOR U11010 ( .A(c2202), .B(n6606), .Z(c2203) );
ANDN U11011 ( .B(n6607), .A(n6608), .Z(n6606) );
XOR U11012 ( .A(c2202), .B(b[2202]), .Z(n6607) );
XNOR U11013 ( .A(b[2202]), .B(n6608), .Z(c[2202]) );
XNOR U11014 ( .A(a[2202]), .B(c2202), .Z(n6608) );
XOR U11015 ( .A(c2203), .B(n6609), .Z(c2204) );
ANDN U11016 ( .B(n6610), .A(n6611), .Z(n6609) );
XOR U11017 ( .A(c2203), .B(b[2203]), .Z(n6610) );
XNOR U11018 ( .A(b[2203]), .B(n6611), .Z(c[2203]) );
XNOR U11019 ( .A(a[2203]), .B(c2203), .Z(n6611) );
XOR U11020 ( .A(c2204), .B(n6612), .Z(c2205) );
ANDN U11021 ( .B(n6613), .A(n6614), .Z(n6612) );
XOR U11022 ( .A(c2204), .B(b[2204]), .Z(n6613) );
XNOR U11023 ( .A(b[2204]), .B(n6614), .Z(c[2204]) );
XNOR U11024 ( .A(a[2204]), .B(c2204), .Z(n6614) );
XOR U11025 ( .A(c2205), .B(n6615), .Z(c2206) );
ANDN U11026 ( .B(n6616), .A(n6617), .Z(n6615) );
XOR U11027 ( .A(c2205), .B(b[2205]), .Z(n6616) );
XNOR U11028 ( .A(b[2205]), .B(n6617), .Z(c[2205]) );
XNOR U11029 ( .A(a[2205]), .B(c2205), .Z(n6617) );
XOR U11030 ( .A(c2206), .B(n6618), .Z(c2207) );
ANDN U11031 ( .B(n6619), .A(n6620), .Z(n6618) );
XOR U11032 ( .A(c2206), .B(b[2206]), .Z(n6619) );
XNOR U11033 ( .A(b[2206]), .B(n6620), .Z(c[2206]) );
XNOR U11034 ( .A(a[2206]), .B(c2206), .Z(n6620) );
XOR U11035 ( .A(c2207), .B(n6621), .Z(c2208) );
ANDN U11036 ( .B(n6622), .A(n6623), .Z(n6621) );
XOR U11037 ( .A(c2207), .B(b[2207]), .Z(n6622) );
XNOR U11038 ( .A(b[2207]), .B(n6623), .Z(c[2207]) );
XNOR U11039 ( .A(a[2207]), .B(c2207), .Z(n6623) );
XOR U11040 ( .A(c2208), .B(n6624), .Z(c2209) );
ANDN U11041 ( .B(n6625), .A(n6626), .Z(n6624) );
XOR U11042 ( .A(c2208), .B(b[2208]), .Z(n6625) );
XNOR U11043 ( .A(b[2208]), .B(n6626), .Z(c[2208]) );
XNOR U11044 ( .A(a[2208]), .B(c2208), .Z(n6626) );
XOR U11045 ( .A(c2209), .B(n6627), .Z(c2210) );
ANDN U11046 ( .B(n6628), .A(n6629), .Z(n6627) );
XOR U11047 ( .A(c2209), .B(b[2209]), .Z(n6628) );
XNOR U11048 ( .A(b[2209]), .B(n6629), .Z(c[2209]) );
XNOR U11049 ( .A(a[2209]), .B(c2209), .Z(n6629) );
XOR U11050 ( .A(c2210), .B(n6630), .Z(c2211) );
ANDN U11051 ( .B(n6631), .A(n6632), .Z(n6630) );
XOR U11052 ( .A(c2210), .B(b[2210]), .Z(n6631) );
XNOR U11053 ( .A(b[2210]), .B(n6632), .Z(c[2210]) );
XNOR U11054 ( .A(a[2210]), .B(c2210), .Z(n6632) );
XOR U11055 ( .A(c2211), .B(n6633), .Z(c2212) );
ANDN U11056 ( .B(n6634), .A(n6635), .Z(n6633) );
XOR U11057 ( .A(c2211), .B(b[2211]), .Z(n6634) );
XNOR U11058 ( .A(b[2211]), .B(n6635), .Z(c[2211]) );
XNOR U11059 ( .A(a[2211]), .B(c2211), .Z(n6635) );
XOR U11060 ( .A(c2212), .B(n6636), .Z(c2213) );
ANDN U11061 ( .B(n6637), .A(n6638), .Z(n6636) );
XOR U11062 ( .A(c2212), .B(b[2212]), .Z(n6637) );
XNOR U11063 ( .A(b[2212]), .B(n6638), .Z(c[2212]) );
XNOR U11064 ( .A(a[2212]), .B(c2212), .Z(n6638) );
XOR U11065 ( .A(c2213), .B(n6639), .Z(c2214) );
ANDN U11066 ( .B(n6640), .A(n6641), .Z(n6639) );
XOR U11067 ( .A(c2213), .B(b[2213]), .Z(n6640) );
XNOR U11068 ( .A(b[2213]), .B(n6641), .Z(c[2213]) );
XNOR U11069 ( .A(a[2213]), .B(c2213), .Z(n6641) );
XOR U11070 ( .A(c2214), .B(n6642), .Z(c2215) );
ANDN U11071 ( .B(n6643), .A(n6644), .Z(n6642) );
XOR U11072 ( .A(c2214), .B(b[2214]), .Z(n6643) );
XNOR U11073 ( .A(b[2214]), .B(n6644), .Z(c[2214]) );
XNOR U11074 ( .A(a[2214]), .B(c2214), .Z(n6644) );
XOR U11075 ( .A(c2215), .B(n6645), .Z(c2216) );
ANDN U11076 ( .B(n6646), .A(n6647), .Z(n6645) );
XOR U11077 ( .A(c2215), .B(b[2215]), .Z(n6646) );
XNOR U11078 ( .A(b[2215]), .B(n6647), .Z(c[2215]) );
XNOR U11079 ( .A(a[2215]), .B(c2215), .Z(n6647) );
XOR U11080 ( .A(c2216), .B(n6648), .Z(c2217) );
ANDN U11081 ( .B(n6649), .A(n6650), .Z(n6648) );
XOR U11082 ( .A(c2216), .B(b[2216]), .Z(n6649) );
XNOR U11083 ( .A(b[2216]), .B(n6650), .Z(c[2216]) );
XNOR U11084 ( .A(a[2216]), .B(c2216), .Z(n6650) );
XOR U11085 ( .A(c2217), .B(n6651), .Z(c2218) );
ANDN U11086 ( .B(n6652), .A(n6653), .Z(n6651) );
XOR U11087 ( .A(c2217), .B(b[2217]), .Z(n6652) );
XNOR U11088 ( .A(b[2217]), .B(n6653), .Z(c[2217]) );
XNOR U11089 ( .A(a[2217]), .B(c2217), .Z(n6653) );
XOR U11090 ( .A(c2218), .B(n6654), .Z(c2219) );
ANDN U11091 ( .B(n6655), .A(n6656), .Z(n6654) );
XOR U11092 ( .A(c2218), .B(b[2218]), .Z(n6655) );
XNOR U11093 ( .A(b[2218]), .B(n6656), .Z(c[2218]) );
XNOR U11094 ( .A(a[2218]), .B(c2218), .Z(n6656) );
XOR U11095 ( .A(c2219), .B(n6657), .Z(c2220) );
ANDN U11096 ( .B(n6658), .A(n6659), .Z(n6657) );
XOR U11097 ( .A(c2219), .B(b[2219]), .Z(n6658) );
XNOR U11098 ( .A(b[2219]), .B(n6659), .Z(c[2219]) );
XNOR U11099 ( .A(a[2219]), .B(c2219), .Z(n6659) );
XOR U11100 ( .A(c2220), .B(n6660), .Z(c2221) );
ANDN U11101 ( .B(n6661), .A(n6662), .Z(n6660) );
XOR U11102 ( .A(c2220), .B(b[2220]), .Z(n6661) );
XNOR U11103 ( .A(b[2220]), .B(n6662), .Z(c[2220]) );
XNOR U11104 ( .A(a[2220]), .B(c2220), .Z(n6662) );
XOR U11105 ( .A(c2221), .B(n6663), .Z(c2222) );
ANDN U11106 ( .B(n6664), .A(n6665), .Z(n6663) );
XOR U11107 ( .A(c2221), .B(b[2221]), .Z(n6664) );
XNOR U11108 ( .A(b[2221]), .B(n6665), .Z(c[2221]) );
XNOR U11109 ( .A(a[2221]), .B(c2221), .Z(n6665) );
XOR U11110 ( .A(c2222), .B(n6666), .Z(c2223) );
ANDN U11111 ( .B(n6667), .A(n6668), .Z(n6666) );
XOR U11112 ( .A(c2222), .B(b[2222]), .Z(n6667) );
XNOR U11113 ( .A(b[2222]), .B(n6668), .Z(c[2222]) );
XNOR U11114 ( .A(a[2222]), .B(c2222), .Z(n6668) );
XOR U11115 ( .A(c2223), .B(n6669), .Z(c2224) );
ANDN U11116 ( .B(n6670), .A(n6671), .Z(n6669) );
XOR U11117 ( .A(c2223), .B(b[2223]), .Z(n6670) );
XNOR U11118 ( .A(b[2223]), .B(n6671), .Z(c[2223]) );
XNOR U11119 ( .A(a[2223]), .B(c2223), .Z(n6671) );
XOR U11120 ( .A(c2224), .B(n6672), .Z(c2225) );
ANDN U11121 ( .B(n6673), .A(n6674), .Z(n6672) );
XOR U11122 ( .A(c2224), .B(b[2224]), .Z(n6673) );
XNOR U11123 ( .A(b[2224]), .B(n6674), .Z(c[2224]) );
XNOR U11124 ( .A(a[2224]), .B(c2224), .Z(n6674) );
XOR U11125 ( .A(c2225), .B(n6675), .Z(c2226) );
ANDN U11126 ( .B(n6676), .A(n6677), .Z(n6675) );
XOR U11127 ( .A(c2225), .B(b[2225]), .Z(n6676) );
XNOR U11128 ( .A(b[2225]), .B(n6677), .Z(c[2225]) );
XNOR U11129 ( .A(a[2225]), .B(c2225), .Z(n6677) );
XOR U11130 ( .A(c2226), .B(n6678), .Z(c2227) );
ANDN U11131 ( .B(n6679), .A(n6680), .Z(n6678) );
XOR U11132 ( .A(c2226), .B(b[2226]), .Z(n6679) );
XNOR U11133 ( .A(b[2226]), .B(n6680), .Z(c[2226]) );
XNOR U11134 ( .A(a[2226]), .B(c2226), .Z(n6680) );
XOR U11135 ( .A(c2227), .B(n6681), .Z(c2228) );
ANDN U11136 ( .B(n6682), .A(n6683), .Z(n6681) );
XOR U11137 ( .A(c2227), .B(b[2227]), .Z(n6682) );
XNOR U11138 ( .A(b[2227]), .B(n6683), .Z(c[2227]) );
XNOR U11139 ( .A(a[2227]), .B(c2227), .Z(n6683) );
XOR U11140 ( .A(c2228), .B(n6684), .Z(c2229) );
ANDN U11141 ( .B(n6685), .A(n6686), .Z(n6684) );
XOR U11142 ( .A(c2228), .B(b[2228]), .Z(n6685) );
XNOR U11143 ( .A(b[2228]), .B(n6686), .Z(c[2228]) );
XNOR U11144 ( .A(a[2228]), .B(c2228), .Z(n6686) );
XOR U11145 ( .A(c2229), .B(n6687), .Z(c2230) );
ANDN U11146 ( .B(n6688), .A(n6689), .Z(n6687) );
XOR U11147 ( .A(c2229), .B(b[2229]), .Z(n6688) );
XNOR U11148 ( .A(b[2229]), .B(n6689), .Z(c[2229]) );
XNOR U11149 ( .A(a[2229]), .B(c2229), .Z(n6689) );
XOR U11150 ( .A(c2230), .B(n6690), .Z(c2231) );
ANDN U11151 ( .B(n6691), .A(n6692), .Z(n6690) );
XOR U11152 ( .A(c2230), .B(b[2230]), .Z(n6691) );
XNOR U11153 ( .A(b[2230]), .B(n6692), .Z(c[2230]) );
XNOR U11154 ( .A(a[2230]), .B(c2230), .Z(n6692) );
XOR U11155 ( .A(c2231), .B(n6693), .Z(c2232) );
ANDN U11156 ( .B(n6694), .A(n6695), .Z(n6693) );
XOR U11157 ( .A(c2231), .B(b[2231]), .Z(n6694) );
XNOR U11158 ( .A(b[2231]), .B(n6695), .Z(c[2231]) );
XNOR U11159 ( .A(a[2231]), .B(c2231), .Z(n6695) );
XOR U11160 ( .A(c2232), .B(n6696), .Z(c2233) );
ANDN U11161 ( .B(n6697), .A(n6698), .Z(n6696) );
XOR U11162 ( .A(c2232), .B(b[2232]), .Z(n6697) );
XNOR U11163 ( .A(b[2232]), .B(n6698), .Z(c[2232]) );
XNOR U11164 ( .A(a[2232]), .B(c2232), .Z(n6698) );
XOR U11165 ( .A(c2233), .B(n6699), .Z(c2234) );
ANDN U11166 ( .B(n6700), .A(n6701), .Z(n6699) );
XOR U11167 ( .A(c2233), .B(b[2233]), .Z(n6700) );
XNOR U11168 ( .A(b[2233]), .B(n6701), .Z(c[2233]) );
XNOR U11169 ( .A(a[2233]), .B(c2233), .Z(n6701) );
XOR U11170 ( .A(c2234), .B(n6702), .Z(c2235) );
ANDN U11171 ( .B(n6703), .A(n6704), .Z(n6702) );
XOR U11172 ( .A(c2234), .B(b[2234]), .Z(n6703) );
XNOR U11173 ( .A(b[2234]), .B(n6704), .Z(c[2234]) );
XNOR U11174 ( .A(a[2234]), .B(c2234), .Z(n6704) );
XOR U11175 ( .A(c2235), .B(n6705), .Z(c2236) );
ANDN U11176 ( .B(n6706), .A(n6707), .Z(n6705) );
XOR U11177 ( .A(c2235), .B(b[2235]), .Z(n6706) );
XNOR U11178 ( .A(b[2235]), .B(n6707), .Z(c[2235]) );
XNOR U11179 ( .A(a[2235]), .B(c2235), .Z(n6707) );
XOR U11180 ( .A(c2236), .B(n6708), .Z(c2237) );
ANDN U11181 ( .B(n6709), .A(n6710), .Z(n6708) );
XOR U11182 ( .A(c2236), .B(b[2236]), .Z(n6709) );
XNOR U11183 ( .A(b[2236]), .B(n6710), .Z(c[2236]) );
XNOR U11184 ( .A(a[2236]), .B(c2236), .Z(n6710) );
XOR U11185 ( .A(c2237), .B(n6711), .Z(c2238) );
ANDN U11186 ( .B(n6712), .A(n6713), .Z(n6711) );
XOR U11187 ( .A(c2237), .B(b[2237]), .Z(n6712) );
XNOR U11188 ( .A(b[2237]), .B(n6713), .Z(c[2237]) );
XNOR U11189 ( .A(a[2237]), .B(c2237), .Z(n6713) );
XOR U11190 ( .A(c2238), .B(n6714), .Z(c2239) );
ANDN U11191 ( .B(n6715), .A(n6716), .Z(n6714) );
XOR U11192 ( .A(c2238), .B(b[2238]), .Z(n6715) );
XNOR U11193 ( .A(b[2238]), .B(n6716), .Z(c[2238]) );
XNOR U11194 ( .A(a[2238]), .B(c2238), .Z(n6716) );
XOR U11195 ( .A(c2239), .B(n6717), .Z(c2240) );
ANDN U11196 ( .B(n6718), .A(n6719), .Z(n6717) );
XOR U11197 ( .A(c2239), .B(b[2239]), .Z(n6718) );
XNOR U11198 ( .A(b[2239]), .B(n6719), .Z(c[2239]) );
XNOR U11199 ( .A(a[2239]), .B(c2239), .Z(n6719) );
XOR U11200 ( .A(c2240), .B(n6720), .Z(c2241) );
ANDN U11201 ( .B(n6721), .A(n6722), .Z(n6720) );
XOR U11202 ( .A(c2240), .B(b[2240]), .Z(n6721) );
XNOR U11203 ( .A(b[2240]), .B(n6722), .Z(c[2240]) );
XNOR U11204 ( .A(a[2240]), .B(c2240), .Z(n6722) );
XOR U11205 ( .A(c2241), .B(n6723), .Z(c2242) );
ANDN U11206 ( .B(n6724), .A(n6725), .Z(n6723) );
XOR U11207 ( .A(c2241), .B(b[2241]), .Z(n6724) );
XNOR U11208 ( .A(b[2241]), .B(n6725), .Z(c[2241]) );
XNOR U11209 ( .A(a[2241]), .B(c2241), .Z(n6725) );
XOR U11210 ( .A(c2242), .B(n6726), .Z(c2243) );
ANDN U11211 ( .B(n6727), .A(n6728), .Z(n6726) );
XOR U11212 ( .A(c2242), .B(b[2242]), .Z(n6727) );
XNOR U11213 ( .A(b[2242]), .B(n6728), .Z(c[2242]) );
XNOR U11214 ( .A(a[2242]), .B(c2242), .Z(n6728) );
XOR U11215 ( .A(c2243), .B(n6729), .Z(c2244) );
ANDN U11216 ( .B(n6730), .A(n6731), .Z(n6729) );
XOR U11217 ( .A(c2243), .B(b[2243]), .Z(n6730) );
XNOR U11218 ( .A(b[2243]), .B(n6731), .Z(c[2243]) );
XNOR U11219 ( .A(a[2243]), .B(c2243), .Z(n6731) );
XOR U11220 ( .A(c2244), .B(n6732), .Z(c2245) );
ANDN U11221 ( .B(n6733), .A(n6734), .Z(n6732) );
XOR U11222 ( .A(c2244), .B(b[2244]), .Z(n6733) );
XNOR U11223 ( .A(b[2244]), .B(n6734), .Z(c[2244]) );
XNOR U11224 ( .A(a[2244]), .B(c2244), .Z(n6734) );
XOR U11225 ( .A(c2245), .B(n6735), .Z(c2246) );
ANDN U11226 ( .B(n6736), .A(n6737), .Z(n6735) );
XOR U11227 ( .A(c2245), .B(b[2245]), .Z(n6736) );
XNOR U11228 ( .A(b[2245]), .B(n6737), .Z(c[2245]) );
XNOR U11229 ( .A(a[2245]), .B(c2245), .Z(n6737) );
XOR U11230 ( .A(c2246), .B(n6738), .Z(c2247) );
ANDN U11231 ( .B(n6739), .A(n6740), .Z(n6738) );
XOR U11232 ( .A(c2246), .B(b[2246]), .Z(n6739) );
XNOR U11233 ( .A(b[2246]), .B(n6740), .Z(c[2246]) );
XNOR U11234 ( .A(a[2246]), .B(c2246), .Z(n6740) );
XOR U11235 ( .A(c2247), .B(n6741), .Z(c2248) );
ANDN U11236 ( .B(n6742), .A(n6743), .Z(n6741) );
XOR U11237 ( .A(c2247), .B(b[2247]), .Z(n6742) );
XNOR U11238 ( .A(b[2247]), .B(n6743), .Z(c[2247]) );
XNOR U11239 ( .A(a[2247]), .B(c2247), .Z(n6743) );
XOR U11240 ( .A(c2248), .B(n6744), .Z(c2249) );
ANDN U11241 ( .B(n6745), .A(n6746), .Z(n6744) );
XOR U11242 ( .A(c2248), .B(b[2248]), .Z(n6745) );
XNOR U11243 ( .A(b[2248]), .B(n6746), .Z(c[2248]) );
XNOR U11244 ( .A(a[2248]), .B(c2248), .Z(n6746) );
XOR U11245 ( .A(c2249), .B(n6747), .Z(c2250) );
ANDN U11246 ( .B(n6748), .A(n6749), .Z(n6747) );
XOR U11247 ( .A(c2249), .B(b[2249]), .Z(n6748) );
XNOR U11248 ( .A(b[2249]), .B(n6749), .Z(c[2249]) );
XNOR U11249 ( .A(a[2249]), .B(c2249), .Z(n6749) );
XOR U11250 ( .A(c2250), .B(n6750), .Z(c2251) );
ANDN U11251 ( .B(n6751), .A(n6752), .Z(n6750) );
XOR U11252 ( .A(c2250), .B(b[2250]), .Z(n6751) );
XNOR U11253 ( .A(b[2250]), .B(n6752), .Z(c[2250]) );
XNOR U11254 ( .A(a[2250]), .B(c2250), .Z(n6752) );
XOR U11255 ( .A(c2251), .B(n6753), .Z(c2252) );
ANDN U11256 ( .B(n6754), .A(n6755), .Z(n6753) );
XOR U11257 ( .A(c2251), .B(b[2251]), .Z(n6754) );
XNOR U11258 ( .A(b[2251]), .B(n6755), .Z(c[2251]) );
XNOR U11259 ( .A(a[2251]), .B(c2251), .Z(n6755) );
XOR U11260 ( .A(c2252), .B(n6756), .Z(c2253) );
ANDN U11261 ( .B(n6757), .A(n6758), .Z(n6756) );
XOR U11262 ( .A(c2252), .B(b[2252]), .Z(n6757) );
XNOR U11263 ( .A(b[2252]), .B(n6758), .Z(c[2252]) );
XNOR U11264 ( .A(a[2252]), .B(c2252), .Z(n6758) );
XOR U11265 ( .A(c2253), .B(n6759), .Z(c2254) );
ANDN U11266 ( .B(n6760), .A(n6761), .Z(n6759) );
XOR U11267 ( .A(c2253), .B(b[2253]), .Z(n6760) );
XNOR U11268 ( .A(b[2253]), .B(n6761), .Z(c[2253]) );
XNOR U11269 ( .A(a[2253]), .B(c2253), .Z(n6761) );
XOR U11270 ( .A(c2254), .B(n6762), .Z(c2255) );
ANDN U11271 ( .B(n6763), .A(n6764), .Z(n6762) );
XOR U11272 ( .A(c2254), .B(b[2254]), .Z(n6763) );
XNOR U11273 ( .A(b[2254]), .B(n6764), .Z(c[2254]) );
XNOR U11274 ( .A(a[2254]), .B(c2254), .Z(n6764) );
XOR U11275 ( .A(c2255), .B(n6765), .Z(c2256) );
ANDN U11276 ( .B(n6766), .A(n6767), .Z(n6765) );
XOR U11277 ( .A(c2255), .B(b[2255]), .Z(n6766) );
XNOR U11278 ( .A(b[2255]), .B(n6767), .Z(c[2255]) );
XNOR U11279 ( .A(a[2255]), .B(c2255), .Z(n6767) );
XOR U11280 ( .A(c2256), .B(n6768), .Z(c2257) );
ANDN U11281 ( .B(n6769), .A(n6770), .Z(n6768) );
XOR U11282 ( .A(c2256), .B(b[2256]), .Z(n6769) );
XNOR U11283 ( .A(b[2256]), .B(n6770), .Z(c[2256]) );
XNOR U11284 ( .A(a[2256]), .B(c2256), .Z(n6770) );
XOR U11285 ( .A(c2257), .B(n6771), .Z(c2258) );
ANDN U11286 ( .B(n6772), .A(n6773), .Z(n6771) );
XOR U11287 ( .A(c2257), .B(b[2257]), .Z(n6772) );
XNOR U11288 ( .A(b[2257]), .B(n6773), .Z(c[2257]) );
XNOR U11289 ( .A(a[2257]), .B(c2257), .Z(n6773) );
XOR U11290 ( .A(c2258), .B(n6774), .Z(c2259) );
ANDN U11291 ( .B(n6775), .A(n6776), .Z(n6774) );
XOR U11292 ( .A(c2258), .B(b[2258]), .Z(n6775) );
XNOR U11293 ( .A(b[2258]), .B(n6776), .Z(c[2258]) );
XNOR U11294 ( .A(a[2258]), .B(c2258), .Z(n6776) );
XOR U11295 ( .A(c2259), .B(n6777), .Z(c2260) );
ANDN U11296 ( .B(n6778), .A(n6779), .Z(n6777) );
XOR U11297 ( .A(c2259), .B(b[2259]), .Z(n6778) );
XNOR U11298 ( .A(b[2259]), .B(n6779), .Z(c[2259]) );
XNOR U11299 ( .A(a[2259]), .B(c2259), .Z(n6779) );
XOR U11300 ( .A(c2260), .B(n6780), .Z(c2261) );
ANDN U11301 ( .B(n6781), .A(n6782), .Z(n6780) );
XOR U11302 ( .A(c2260), .B(b[2260]), .Z(n6781) );
XNOR U11303 ( .A(b[2260]), .B(n6782), .Z(c[2260]) );
XNOR U11304 ( .A(a[2260]), .B(c2260), .Z(n6782) );
XOR U11305 ( .A(c2261), .B(n6783), .Z(c2262) );
ANDN U11306 ( .B(n6784), .A(n6785), .Z(n6783) );
XOR U11307 ( .A(c2261), .B(b[2261]), .Z(n6784) );
XNOR U11308 ( .A(b[2261]), .B(n6785), .Z(c[2261]) );
XNOR U11309 ( .A(a[2261]), .B(c2261), .Z(n6785) );
XOR U11310 ( .A(c2262), .B(n6786), .Z(c2263) );
ANDN U11311 ( .B(n6787), .A(n6788), .Z(n6786) );
XOR U11312 ( .A(c2262), .B(b[2262]), .Z(n6787) );
XNOR U11313 ( .A(b[2262]), .B(n6788), .Z(c[2262]) );
XNOR U11314 ( .A(a[2262]), .B(c2262), .Z(n6788) );
XOR U11315 ( .A(c2263), .B(n6789), .Z(c2264) );
ANDN U11316 ( .B(n6790), .A(n6791), .Z(n6789) );
XOR U11317 ( .A(c2263), .B(b[2263]), .Z(n6790) );
XNOR U11318 ( .A(b[2263]), .B(n6791), .Z(c[2263]) );
XNOR U11319 ( .A(a[2263]), .B(c2263), .Z(n6791) );
XOR U11320 ( .A(c2264), .B(n6792), .Z(c2265) );
ANDN U11321 ( .B(n6793), .A(n6794), .Z(n6792) );
XOR U11322 ( .A(c2264), .B(b[2264]), .Z(n6793) );
XNOR U11323 ( .A(b[2264]), .B(n6794), .Z(c[2264]) );
XNOR U11324 ( .A(a[2264]), .B(c2264), .Z(n6794) );
XOR U11325 ( .A(c2265), .B(n6795), .Z(c2266) );
ANDN U11326 ( .B(n6796), .A(n6797), .Z(n6795) );
XOR U11327 ( .A(c2265), .B(b[2265]), .Z(n6796) );
XNOR U11328 ( .A(b[2265]), .B(n6797), .Z(c[2265]) );
XNOR U11329 ( .A(a[2265]), .B(c2265), .Z(n6797) );
XOR U11330 ( .A(c2266), .B(n6798), .Z(c2267) );
ANDN U11331 ( .B(n6799), .A(n6800), .Z(n6798) );
XOR U11332 ( .A(c2266), .B(b[2266]), .Z(n6799) );
XNOR U11333 ( .A(b[2266]), .B(n6800), .Z(c[2266]) );
XNOR U11334 ( .A(a[2266]), .B(c2266), .Z(n6800) );
XOR U11335 ( .A(c2267), .B(n6801), .Z(c2268) );
ANDN U11336 ( .B(n6802), .A(n6803), .Z(n6801) );
XOR U11337 ( .A(c2267), .B(b[2267]), .Z(n6802) );
XNOR U11338 ( .A(b[2267]), .B(n6803), .Z(c[2267]) );
XNOR U11339 ( .A(a[2267]), .B(c2267), .Z(n6803) );
XOR U11340 ( .A(c2268), .B(n6804), .Z(c2269) );
ANDN U11341 ( .B(n6805), .A(n6806), .Z(n6804) );
XOR U11342 ( .A(c2268), .B(b[2268]), .Z(n6805) );
XNOR U11343 ( .A(b[2268]), .B(n6806), .Z(c[2268]) );
XNOR U11344 ( .A(a[2268]), .B(c2268), .Z(n6806) );
XOR U11345 ( .A(c2269), .B(n6807), .Z(c2270) );
ANDN U11346 ( .B(n6808), .A(n6809), .Z(n6807) );
XOR U11347 ( .A(c2269), .B(b[2269]), .Z(n6808) );
XNOR U11348 ( .A(b[2269]), .B(n6809), .Z(c[2269]) );
XNOR U11349 ( .A(a[2269]), .B(c2269), .Z(n6809) );
XOR U11350 ( .A(c2270), .B(n6810), .Z(c2271) );
ANDN U11351 ( .B(n6811), .A(n6812), .Z(n6810) );
XOR U11352 ( .A(c2270), .B(b[2270]), .Z(n6811) );
XNOR U11353 ( .A(b[2270]), .B(n6812), .Z(c[2270]) );
XNOR U11354 ( .A(a[2270]), .B(c2270), .Z(n6812) );
XOR U11355 ( .A(c2271), .B(n6813), .Z(c2272) );
ANDN U11356 ( .B(n6814), .A(n6815), .Z(n6813) );
XOR U11357 ( .A(c2271), .B(b[2271]), .Z(n6814) );
XNOR U11358 ( .A(b[2271]), .B(n6815), .Z(c[2271]) );
XNOR U11359 ( .A(a[2271]), .B(c2271), .Z(n6815) );
XOR U11360 ( .A(c2272), .B(n6816), .Z(c2273) );
ANDN U11361 ( .B(n6817), .A(n6818), .Z(n6816) );
XOR U11362 ( .A(c2272), .B(b[2272]), .Z(n6817) );
XNOR U11363 ( .A(b[2272]), .B(n6818), .Z(c[2272]) );
XNOR U11364 ( .A(a[2272]), .B(c2272), .Z(n6818) );
XOR U11365 ( .A(c2273), .B(n6819), .Z(c2274) );
ANDN U11366 ( .B(n6820), .A(n6821), .Z(n6819) );
XOR U11367 ( .A(c2273), .B(b[2273]), .Z(n6820) );
XNOR U11368 ( .A(b[2273]), .B(n6821), .Z(c[2273]) );
XNOR U11369 ( .A(a[2273]), .B(c2273), .Z(n6821) );
XOR U11370 ( .A(c2274), .B(n6822), .Z(c2275) );
ANDN U11371 ( .B(n6823), .A(n6824), .Z(n6822) );
XOR U11372 ( .A(c2274), .B(b[2274]), .Z(n6823) );
XNOR U11373 ( .A(b[2274]), .B(n6824), .Z(c[2274]) );
XNOR U11374 ( .A(a[2274]), .B(c2274), .Z(n6824) );
XOR U11375 ( .A(c2275), .B(n6825), .Z(c2276) );
ANDN U11376 ( .B(n6826), .A(n6827), .Z(n6825) );
XOR U11377 ( .A(c2275), .B(b[2275]), .Z(n6826) );
XNOR U11378 ( .A(b[2275]), .B(n6827), .Z(c[2275]) );
XNOR U11379 ( .A(a[2275]), .B(c2275), .Z(n6827) );
XOR U11380 ( .A(c2276), .B(n6828), .Z(c2277) );
ANDN U11381 ( .B(n6829), .A(n6830), .Z(n6828) );
XOR U11382 ( .A(c2276), .B(b[2276]), .Z(n6829) );
XNOR U11383 ( .A(b[2276]), .B(n6830), .Z(c[2276]) );
XNOR U11384 ( .A(a[2276]), .B(c2276), .Z(n6830) );
XOR U11385 ( .A(c2277), .B(n6831), .Z(c2278) );
ANDN U11386 ( .B(n6832), .A(n6833), .Z(n6831) );
XOR U11387 ( .A(c2277), .B(b[2277]), .Z(n6832) );
XNOR U11388 ( .A(b[2277]), .B(n6833), .Z(c[2277]) );
XNOR U11389 ( .A(a[2277]), .B(c2277), .Z(n6833) );
XOR U11390 ( .A(c2278), .B(n6834), .Z(c2279) );
ANDN U11391 ( .B(n6835), .A(n6836), .Z(n6834) );
XOR U11392 ( .A(c2278), .B(b[2278]), .Z(n6835) );
XNOR U11393 ( .A(b[2278]), .B(n6836), .Z(c[2278]) );
XNOR U11394 ( .A(a[2278]), .B(c2278), .Z(n6836) );
XOR U11395 ( .A(c2279), .B(n6837), .Z(c2280) );
ANDN U11396 ( .B(n6838), .A(n6839), .Z(n6837) );
XOR U11397 ( .A(c2279), .B(b[2279]), .Z(n6838) );
XNOR U11398 ( .A(b[2279]), .B(n6839), .Z(c[2279]) );
XNOR U11399 ( .A(a[2279]), .B(c2279), .Z(n6839) );
XOR U11400 ( .A(c2280), .B(n6840), .Z(c2281) );
ANDN U11401 ( .B(n6841), .A(n6842), .Z(n6840) );
XOR U11402 ( .A(c2280), .B(b[2280]), .Z(n6841) );
XNOR U11403 ( .A(b[2280]), .B(n6842), .Z(c[2280]) );
XNOR U11404 ( .A(a[2280]), .B(c2280), .Z(n6842) );
XOR U11405 ( .A(c2281), .B(n6843), .Z(c2282) );
ANDN U11406 ( .B(n6844), .A(n6845), .Z(n6843) );
XOR U11407 ( .A(c2281), .B(b[2281]), .Z(n6844) );
XNOR U11408 ( .A(b[2281]), .B(n6845), .Z(c[2281]) );
XNOR U11409 ( .A(a[2281]), .B(c2281), .Z(n6845) );
XOR U11410 ( .A(c2282), .B(n6846), .Z(c2283) );
ANDN U11411 ( .B(n6847), .A(n6848), .Z(n6846) );
XOR U11412 ( .A(c2282), .B(b[2282]), .Z(n6847) );
XNOR U11413 ( .A(b[2282]), .B(n6848), .Z(c[2282]) );
XNOR U11414 ( .A(a[2282]), .B(c2282), .Z(n6848) );
XOR U11415 ( .A(c2283), .B(n6849), .Z(c2284) );
ANDN U11416 ( .B(n6850), .A(n6851), .Z(n6849) );
XOR U11417 ( .A(c2283), .B(b[2283]), .Z(n6850) );
XNOR U11418 ( .A(b[2283]), .B(n6851), .Z(c[2283]) );
XNOR U11419 ( .A(a[2283]), .B(c2283), .Z(n6851) );
XOR U11420 ( .A(c2284), .B(n6852), .Z(c2285) );
ANDN U11421 ( .B(n6853), .A(n6854), .Z(n6852) );
XOR U11422 ( .A(c2284), .B(b[2284]), .Z(n6853) );
XNOR U11423 ( .A(b[2284]), .B(n6854), .Z(c[2284]) );
XNOR U11424 ( .A(a[2284]), .B(c2284), .Z(n6854) );
XOR U11425 ( .A(c2285), .B(n6855), .Z(c2286) );
ANDN U11426 ( .B(n6856), .A(n6857), .Z(n6855) );
XOR U11427 ( .A(c2285), .B(b[2285]), .Z(n6856) );
XNOR U11428 ( .A(b[2285]), .B(n6857), .Z(c[2285]) );
XNOR U11429 ( .A(a[2285]), .B(c2285), .Z(n6857) );
XOR U11430 ( .A(c2286), .B(n6858), .Z(c2287) );
ANDN U11431 ( .B(n6859), .A(n6860), .Z(n6858) );
XOR U11432 ( .A(c2286), .B(b[2286]), .Z(n6859) );
XNOR U11433 ( .A(b[2286]), .B(n6860), .Z(c[2286]) );
XNOR U11434 ( .A(a[2286]), .B(c2286), .Z(n6860) );
XOR U11435 ( .A(c2287), .B(n6861), .Z(c2288) );
ANDN U11436 ( .B(n6862), .A(n6863), .Z(n6861) );
XOR U11437 ( .A(c2287), .B(b[2287]), .Z(n6862) );
XNOR U11438 ( .A(b[2287]), .B(n6863), .Z(c[2287]) );
XNOR U11439 ( .A(a[2287]), .B(c2287), .Z(n6863) );
XOR U11440 ( .A(c2288), .B(n6864), .Z(c2289) );
ANDN U11441 ( .B(n6865), .A(n6866), .Z(n6864) );
XOR U11442 ( .A(c2288), .B(b[2288]), .Z(n6865) );
XNOR U11443 ( .A(b[2288]), .B(n6866), .Z(c[2288]) );
XNOR U11444 ( .A(a[2288]), .B(c2288), .Z(n6866) );
XOR U11445 ( .A(c2289), .B(n6867), .Z(c2290) );
ANDN U11446 ( .B(n6868), .A(n6869), .Z(n6867) );
XOR U11447 ( .A(c2289), .B(b[2289]), .Z(n6868) );
XNOR U11448 ( .A(b[2289]), .B(n6869), .Z(c[2289]) );
XNOR U11449 ( .A(a[2289]), .B(c2289), .Z(n6869) );
XOR U11450 ( .A(c2290), .B(n6870), .Z(c2291) );
ANDN U11451 ( .B(n6871), .A(n6872), .Z(n6870) );
XOR U11452 ( .A(c2290), .B(b[2290]), .Z(n6871) );
XNOR U11453 ( .A(b[2290]), .B(n6872), .Z(c[2290]) );
XNOR U11454 ( .A(a[2290]), .B(c2290), .Z(n6872) );
XOR U11455 ( .A(c2291), .B(n6873), .Z(c2292) );
ANDN U11456 ( .B(n6874), .A(n6875), .Z(n6873) );
XOR U11457 ( .A(c2291), .B(b[2291]), .Z(n6874) );
XNOR U11458 ( .A(b[2291]), .B(n6875), .Z(c[2291]) );
XNOR U11459 ( .A(a[2291]), .B(c2291), .Z(n6875) );
XOR U11460 ( .A(c2292), .B(n6876), .Z(c2293) );
ANDN U11461 ( .B(n6877), .A(n6878), .Z(n6876) );
XOR U11462 ( .A(c2292), .B(b[2292]), .Z(n6877) );
XNOR U11463 ( .A(b[2292]), .B(n6878), .Z(c[2292]) );
XNOR U11464 ( .A(a[2292]), .B(c2292), .Z(n6878) );
XOR U11465 ( .A(c2293), .B(n6879), .Z(c2294) );
ANDN U11466 ( .B(n6880), .A(n6881), .Z(n6879) );
XOR U11467 ( .A(c2293), .B(b[2293]), .Z(n6880) );
XNOR U11468 ( .A(b[2293]), .B(n6881), .Z(c[2293]) );
XNOR U11469 ( .A(a[2293]), .B(c2293), .Z(n6881) );
XOR U11470 ( .A(c2294), .B(n6882), .Z(c2295) );
ANDN U11471 ( .B(n6883), .A(n6884), .Z(n6882) );
XOR U11472 ( .A(c2294), .B(b[2294]), .Z(n6883) );
XNOR U11473 ( .A(b[2294]), .B(n6884), .Z(c[2294]) );
XNOR U11474 ( .A(a[2294]), .B(c2294), .Z(n6884) );
XOR U11475 ( .A(c2295), .B(n6885), .Z(c2296) );
ANDN U11476 ( .B(n6886), .A(n6887), .Z(n6885) );
XOR U11477 ( .A(c2295), .B(b[2295]), .Z(n6886) );
XNOR U11478 ( .A(b[2295]), .B(n6887), .Z(c[2295]) );
XNOR U11479 ( .A(a[2295]), .B(c2295), .Z(n6887) );
XOR U11480 ( .A(c2296), .B(n6888), .Z(c2297) );
ANDN U11481 ( .B(n6889), .A(n6890), .Z(n6888) );
XOR U11482 ( .A(c2296), .B(b[2296]), .Z(n6889) );
XNOR U11483 ( .A(b[2296]), .B(n6890), .Z(c[2296]) );
XNOR U11484 ( .A(a[2296]), .B(c2296), .Z(n6890) );
XOR U11485 ( .A(c2297), .B(n6891), .Z(c2298) );
ANDN U11486 ( .B(n6892), .A(n6893), .Z(n6891) );
XOR U11487 ( .A(c2297), .B(b[2297]), .Z(n6892) );
XNOR U11488 ( .A(b[2297]), .B(n6893), .Z(c[2297]) );
XNOR U11489 ( .A(a[2297]), .B(c2297), .Z(n6893) );
XOR U11490 ( .A(c2298), .B(n6894), .Z(c2299) );
ANDN U11491 ( .B(n6895), .A(n6896), .Z(n6894) );
XOR U11492 ( .A(c2298), .B(b[2298]), .Z(n6895) );
XNOR U11493 ( .A(b[2298]), .B(n6896), .Z(c[2298]) );
XNOR U11494 ( .A(a[2298]), .B(c2298), .Z(n6896) );
XOR U11495 ( .A(c2299), .B(n6897), .Z(c2300) );
ANDN U11496 ( .B(n6898), .A(n6899), .Z(n6897) );
XOR U11497 ( .A(c2299), .B(b[2299]), .Z(n6898) );
XNOR U11498 ( .A(b[2299]), .B(n6899), .Z(c[2299]) );
XNOR U11499 ( .A(a[2299]), .B(c2299), .Z(n6899) );
XOR U11500 ( .A(c2300), .B(n6900), .Z(c2301) );
ANDN U11501 ( .B(n6901), .A(n6902), .Z(n6900) );
XOR U11502 ( .A(c2300), .B(b[2300]), .Z(n6901) );
XNOR U11503 ( .A(b[2300]), .B(n6902), .Z(c[2300]) );
XNOR U11504 ( .A(a[2300]), .B(c2300), .Z(n6902) );
XOR U11505 ( .A(c2301), .B(n6903), .Z(c2302) );
ANDN U11506 ( .B(n6904), .A(n6905), .Z(n6903) );
XOR U11507 ( .A(c2301), .B(b[2301]), .Z(n6904) );
XNOR U11508 ( .A(b[2301]), .B(n6905), .Z(c[2301]) );
XNOR U11509 ( .A(a[2301]), .B(c2301), .Z(n6905) );
XOR U11510 ( .A(c2302), .B(n6906), .Z(c2303) );
ANDN U11511 ( .B(n6907), .A(n6908), .Z(n6906) );
XOR U11512 ( .A(c2302), .B(b[2302]), .Z(n6907) );
XNOR U11513 ( .A(b[2302]), .B(n6908), .Z(c[2302]) );
XNOR U11514 ( .A(a[2302]), .B(c2302), .Z(n6908) );
XOR U11515 ( .A(c2303), .B(n6909), .Z(c2304) );
ANDN U11516 ( .B(n6910), .A(n6911), .Z(n6909) );
XOR U11517 ( .A(c2303), .B(b[2303]), .Z(n6910) );
XNOR U11518 ( .A(b[2303]), .B(n6911), .Z(c[2303]) );
XNOR U11519 ( .A(a[2303]), .B(c2303), .Z(n6911) );
XOR U11520 ( .A(c2304), .B(n6912), .Z(c2305) );
ANDN U11521 ( .B(n6913), .A(n6914), .Z(n6912) );
XOR U11522 ( .A(c2304), .B(b[2304]), .Z(n6913) );
XNOR U11523 ( .A(b[2304]), .B(n6914), .Z(c[2304]) );
XNOR U11524 ( .A(a[2304]), .B(c2304), .Z(n6914) );
XOR U11525 ( .A(c2305), .B(n6915), .Z(c2306) );
ANDN U11526 ( .B(n6916), .A(n6917), .Z(n6915) );
XOR U11527 ( .A(c2305), .B(b[2305]), .Z(n6916) );
XNOR U11528 ( .A(b[2305]), .B(n6917), .Z(c[2305]) );
XNOR U11529 ( .A(a[2305]), .B(c2305), .Z(n6917) );
XOR U11530 ( .A(c2306), .B(n6918), .Z(c2307) );
ANDN U11531 ( .B(n6919), .A(n6920), .Z(n6918) );
XOR U11532 ( .A(c2306), .B(b[2306]), .Z(n6919) );
XNOR U11533 ( .A(b[2306]), .B(n6920), .Z(c[2306]) );
XNOR U11534 ( .A(a[2306]), .B(c2306), .Z(n6920) );
XOR U11535 ( .A(c2307), .B(n6921), .Z(c2308) );
ANDN U11536 ( .B(n6922), .A(n6923), .Z(n6921) );
XOR U11537 ( .A(c2307), .B(b[2307]), .Z(n6922) );
XNOR U11538 ( .A(b[2307]), .B(n6923), .Z(c[2307]) );
XNOR U11539 ( .A(a[2307]), .B(c2307), .Z(n6923) );
XOR U11540 ( .A(c2308), .B(n6924), .Z(c2309) );
ANDN U11541 ( .B(n6925), .A(n6926), .Z(n6924) );
XOR U11542 ( .A(c2308), .B(b[2308]), .Z(n6925) );
XNOR U11543 ( .A(b[2308]), .B(n6926), .Z(c[2308]) );
XNOR U11544 ( .A(a[2308]), .B(c2308), .Z(n6926) );
XOR U11545 ( .A(c2309), .B(n6927), .Z(c2310) );
ANDN U11546 ( .B(n6928), .A(n6929), .Z(n6927) );
XOR U11547 ( .A(c2309), .B(b[2309]), .Z(n6928) );
XNOR U11548 ( .A(b[2309]), .B(n6929), .Z(c[2309]) );
XNOR U11549 ( .A(a[2309]), .B(c2309), .Z(n6929) );
XOR U11550 ( .A(c2310), .B(n6930), .Z(c2311) );
ANDN U11551 ( .B(n6931), .A(n6932), .Z(n6930) );
XOR U11552 ( .A(c2310), .B(b[2310]), .Z(n6931) );
XNOR U11553 ( .A(b[2310]), .B(n6932), .Z(c[2310]) );
XNOR U11554 ( .A(a[2310]), .B(c2310), .Z(n6932) );
XOR U11555 ( .A(c2311), .B(n6933), .Z(c2312) );
ANDN U11556 ( .B(n6934), .A(n6935), .Z(n6933) );
XOR U11557 ( .A(c2311), .B(b[2311]), .Z(n6934) );
XNOR U11558 ( .A(b[2311]), .B(n6935), .Z(c[2311]) );
XNOR U11559 ( .A(a[2311]), .B(c2311), .Z(n6935) );
XOR U11560 ( .A(c2312), .B(n6936), .Z(c2313) );
ANDN U11561 ( .B(n6937), .A(n6938), .Z(n6936) );
XOR U11562 ( .A(c2312), .B(b[2312]), .Z(n6937) );
XNOR U11563 ( .A(b[2312]), .B(n6938), .Z(c[2312]) );
XNOR U11564 ( .A(a[2312]), .B(c2312), .Z(n6938) );
XOR U11565 ( .A(c2313), .B(n6939), .Z(c2314) );
ANDN U11566 ( .B(n6940), .A(n6941), .Z(n6939) );
XOR U11567 ( .A(c2313), .B(b[2313]), .Z(n6940) );
XNOR U11568 ( .A(b[2313]), .B(n6941), .Z(c[2313]) );
XNOR U11569 ( .A(a[2313]), .B(c2313), .Z(n6941) );
XOR U11570 ( .A(c2314), .B(n6942), .Z(c2315) );
ANDN U11571 ( .B(n6943), .A(n6944), .Z(n6942) );
XOR U11572 ( .A(c2314), .B(b[2314]), .Z(n6943) );
XNOR U11573 ( .A(b[2314]), .B(n6944), .Z(c[2314]) );
XNOR U11574 ( .A(a[2314]), .B(c2314), .Z(n6944) );
XOR U11575 ( .A(c2315), .B(n6945), .Z(c2316) );
ANDN U11576 ( .B(n6946), .A(n6947), .Z(n6945) );
XOR U11577 ( .A(c2315), .B(b[2315]), .Z(n6946) );
XNOR U11578 ( .A(b[2315]), .B(n6947), .Z(c[2315]) );
XNOR U11579 ( .A(a[2315]), .B(c2315), .Z(n6947) );
XOR U11580 ( .A(c2316), .B(n6948), .Z(c2317) );
ANDN U11581 ( .B(n6949), .A(n6950), .Z(n6948) );
XOR U11582 ( .A(c2316), .B(b[2316]), .Z(n6949) );
XNOR U11583 ( .A(b[2316]), .B(n6950), .Z(c[2316]) );
XNOR U11584 ( .A(a[2316]), .B(c2316), .Z(n6950) );
XOR U11585 ( .A(c2317), .B(n6951), .Z(c2318) );
ANDN U11586 ( .B(n6952), .A(n6953), .Z(n6951) );
XOR U11587 ( .A(c2317), .B(b[2317]), .Z(n6952) );
XNOR U11588 ( .A(b[2317]), .B(n6953), .Z(c[2317]) );
XNOR U11589 ( .A(a[2317]), .B(c2317), .Z(n6953) );
XOR U11590 ( .A(c2318), .B(n6954), .Z(c2319) );
ANDN U11591 ( .B(n6955), .A(n6956), .Z(n6954) );
XOR U11592 ( .A(c2318), .B(b[2318]), .Z(n6955) );
XNOR U11593 ( .A(b[2318]), .B(n6956), .Z(c[2318]) );
XNOR U11594 ( .A(a[2318]), .B(c2318), .Z(n6956) );
XOR U11595 ( .A(c2319), .B(n6957), .Z(c2320) );
ANDN U11596 ( .B(n6958), .A(n6959), .Z(n6957) );
XOR U11597 ( .A(c2319), .B(b[2319]), .Z(n6958) );
XNOR U11598 ( .A(b[2319]), .B(n6959), .Z(c[2319]) );
XNOR U11599 ( .A(a[2319]), .B(c2319), .Z(n6959) );
XOR U11600 ( .A(c2320), .B(n6960), .Z(c2321) );
ANDN U11601 ( .B(n6961), .A(n6962), .Z(n6960) );
XOR U11602 ( .A(c2320), .B(b[2320]), .Z(n6961) );
XNOR U11603 ( .A(b[2320]), .B(n6962), .Z(c[2320]) );
XNOR U11604 ( .A(a[2320]), .B(c2320), .Z(n6962) );
XOR U11605 ( .A(c2321), .B(n6963), .Z(c2322) );
ANDN U11606 ( .B(n6964), .A(n6965), .Z(n6963) );
XOR U11607 ( .A(c2321), .B(b[2321]), .Z(n6964) );
XNOR U11608 ( .A(b[2321]), .B(n6965), .Z(c[2321]) );
XNOR U11609 ( .A(a[2321]), .B(c2321), .Z(n6965) );
XOR U11610 ( .A(c2322), .B(n6966), .Z(c2323) );
ANDN U11611 ( .B(n6967), .A(n6968), .Z(n6966) );
XOR U11612 ( .A(c2322), .B(b[2322]), .Z(n6967) );
XNOR U11613 ( .A(b[2322]), .B(n6968), .Z(c[2322]) );
XNOR U11614 ( .A(a[2322]), .B(c2322), .Z(n6968) );
XOR U11615 ( .A(c2323), .B(n6969), .Z(c2324) );
ANDN U11616 ( .B(n6970), .A(n6971), .Z(n6969) );
XOR U11617 ( .A(c2323), .B(b[2323]), .Z(n6970) );
XNOR U11618 ( .A(b[2323]), .B(n6971), .Z(c[2323]) );
XNOR U11619 ( .A(a[2323]), .B(c2323), .Z(n6971) );
XOR U11620 ( .A(c2324), .B(n6972), .Z(c2325) );
ANDN U11621 ( .B(n6973), .A(n6974), .Z(n6972) );
XOR U11622 ( .A(c2324), .B(b[2324]), .Z(n6973) );
XNOR U11623 ( .A(b[2324]), .B(n6974), .Z(c[2324]) );
XNOR U11624 ( .A(a[2324]), .B(c2324), .Z(n6974) );
XOR U11625 ( .A(c2325), .B(n6975), .Z(c2326) );
ANDN U11626 ( .B(n6976), .A(n6977), .Z(n6975) );
XOR U11627 ( .A(c2325), .B(b[2325]), .Z(n6976) );
XNOR U11628 ( .A(b[2325]), .B(n6977), .Z(c[2325]) );
XNOR U11629 ( .A(a[2325]), .B(c2325), .Z(n6977) );
XOR U11630 ( .A(c2326), .B(n6978), .Z(c2327) );
ANDN U11631 ( .B(n6979), .A(n6980), .Z(n6978) );
XOR U11632 ( .A(c2326), .B(b[2326]), .Z(n6979) );
XNOR U11633 ( .A(b[2326]), .B(n6980), .Z(c[2326]) );
XNOR U11634 ( .A(a[2326]), .B(c2326), .Z(n6980) );
XOR U11635 ( .A(c2327), .B(n6981), .Z(c2328) );
ANDN U11636 ( .B(n6982), .A(n6983), .Z(n6981) );
XOR U11637 ( .A(c2327), .B(b[2327]), .Z(n6982) );
XNOR U11638 ( .A(b[2327]), .B(n6983), .Z(c[2327]) );
XNOR U11639 ( .A(a[2327]), .B(c2327), .Z(n6983) );
XOR U11640 ( .A(c2328), .B(n6984), .Z(c2329) );
ANDN U11641 ( .B(n6985), .A(n6986), .Z(n6984) );
XOR U11642 ( .A(c2328), .B(b[2328]), .Z(n6985) );
XNOR U11643 ( .A(b[2328]), .B(n6986), .Z(c[2328]) );
XNOR U11644 ( .A(a[2328]), .B(c2328), .Z(n6986) );
XOR U11645 ( .A(c2329), .B(n6987), .Z(c2330) );
ANDN U11646 ( .B(n6988), .A(n6989), .Z(n6987) );
XOR U11647 ( .A(c2329), .B(b[2329]), .Z(n6988) );
XNOR U11648 ( .A(b[2329]), .B(n6989), .Z(c[2329]) );
XNOR U11649 ( .A(a[2329]), .B(c2329), .Z(n6989) );
XOR U11650 ( .A(c2330), .B(n6990), .Z(c2331) );
ANDN U11651 ( .B(n6991), .A(n6992), .Z(n6990) );
XOR U11652 ( .A(c2330), .B(b[2330]), .Z(n6991) );
XNOR U11653 ( .A(b[2330]), .B(n6992), .Z(c[2330]) );
XNOR U11654 ( .A(a[2330]), .B(c2330), .Z(n6992) );
XOR U11655 ( .A(c2331), .B(n6993), .Z(c2332) );
ANDN U11656 ( .B(n6994), .A(n6995), .Z(n6993) );
XOR U11657 ( .A(c2331), .B(b[2331]), .Z(n6994) );
XNOR U11658 ( .A(b[2331]), .B(n6995), .Z(c[2331]) );
XNOR U11659 ( .A(a[2331]), .B(c2331), .Z(n6995) );
XOR U11660 ( .A(c2332), .B(n6996), .Z(c2333) );
ANDN U11661 ( .B(n6997), .A(n6998), .Z(n6996) );
XOR U11662 ( .A(c2332), .B(b[2332]), .Z(n6997) );
XNOR U11663 ( .A(b[2332]), .B(n6998), .Z(c[2332]) );
XNOR U11664 ( .A(a[2332]), .B(c2332), .Z(n6998) );
XOR U11665 ( .A(c2333), .B(n6999), .Z(c2334) );
ANDN U11666 ( .B(n7000), .A(n7001), .Z(n6999) );
XOR U11667 ( .A(c2333), .B(b[2333]), .Z(n7000) );
XNOR U11668 ( .A(b[2333]), .B(n7001), .Z(c[2333]) );
XNOR U11669 ( .A(a[2333]), .B(c2333), .Z(n7001) );
XOR U11670 ( .A(c2334), .B(n7002), .Z(c2335) );
ANDN U11671 ( .B(n7003), .A(n7004), .Z(n7002) );
XOR U11672 ( .A(c2334), .B(b[2334]), .Z(n7003) );
XNOR U11673 ( .A(b[2334]), .B(n7004), .Z(c[2334]) );
XNOR U11674 ( .A(a[2334]), .B(c2334), .Z(n7004) );
XOR U11675 ( .A(c2335), .B(n7005), .Z(c2336) );
ANDN U11676 ( .B(n7006), .A(n7007), .Z(n7005) );
XOR U11677 ( .A(c2335), .B(b[2335]), .Z(n7006) );
XNOR U11678 ( .A(b[2335]), .B(n7007), .Z(c[2335]) );
XNOR U11679 ( .A(a[2335]), .B(c2335), .Z(n7007) );
XOR U11680 ( .A(c2336), .B(n7008), .Z(c2337) );
ANDN U11681 ( .B(n7009), .A(n7010), .Z(n7008) );
XOR U11682 ( .A(c2336), .B(b[2336]), .Z(n7009) );
XNOR U11683 ( .A(b[2336]), .B(n7010), .Z(c[2336]) );
XNOR U11684 ( .A(a[2336]), .B(c2336), .Z(n7010) );
XOR U11685 ( .A(c2337), .B(n7011), .Z(c2338) );
ANDN U11686 ( .B(n7012), .A(n7013), .Z(n7011) );
XOR U11687 ( .A(c2337), .B(b[2337]), .Z(n7012) );
XNOR U11688 ( .A(b[2337]), .B(n7013), .Z(c[2337]) );
XNOR U11689 ( .A(a[2337]), .B(c2337), .Z(n7013) );
XOR U11690 ( .A(c2338), .B(n7014), .Z(c2339) );
ANDN U11691 ( .B(n7015), .A(n7016), .Z(n7014) );
XOR U11692 ( .A(c2338), .B(b[2338]), .Z(n7015) );
XNOR U11693 ( .A(b[2338]), .B(n7016), .Z(c[2338]) );
XNOR U11694 ( .A(a[2338]), .B(c2338), .Z(n7016) );
XOR U11695 ( .A(c2339), .B(n7017), .Z(c2340) );
ANDN U11696 ( .B(n7018), .A(n7019), .Z(n7017) );
XOR U11697 ( .A(c2339), .B(b[2339]), .Z(n7018) );
XNOR U11698 ( .A(b[2339]), .B(n7019), .Z(c[2339]) );
XNOR U11699 ( .A(a[2339]), .B(c2339), .Z(n7019) );
XOR U11700 ( .A(c2340), .B(n7020), .Z(c2341) );
ANDN U11701 ( .B(n7021), .A(n7022), .Z(n7020) );
XOR U11702 ( .A(c2340), .B(b[2340]), .Z(n7021) );
XNOR U11703 ( .A(b[2340]), .B(n7022), .Z(c[2340]) );
XNOR U11704 ( .A(a[2340]), .B(c2340), .Z(n7022) );
XOR U11705 ( .A(c2341), .B(n7023), .Z(c2342) );
ANDN U11706 ( .B(n7024), .A(n7025), .Z(n7023) );
XOR U11707 ( .A(c2341), .B(b[2341]), .Z(n7024) );
XNOR U11708 ( .A(b[2341]), .B(n7025), .Z(c[2341]) );
XNOR U11709 ( .A(a[2341]), .B(c2341), .Z(n7025) );
XOR U11710 ( .A(c2342), .B(n7026), .Z(c2343) );
ANDN U11711 ( .B(n7027), .A(n7028), .Z(n7026) );
XOR U11712 ( .A(c2342), .B(b[2342]), .Z(n7027) );
XNOR U11713 ( .A(b[2342]), .B(n7028), .Z(c[2342]) );
XNOR U11714 ( .A(a[2342]), .B(c2342), .Z(n7028) );
XOR U11715 ( .A(c2343), .B(n7029), .Z(c2344) );
ANDN U11716 ( .B(n7030), .A(n7031), .Z(n7029) );
XOR U11717 ( .A(c2343), .B(b[2343]), .Z(n7030) );
XNOR U11718 ( .A(b[2343]), .B(n7031), .Z(c[2343]) );
XNOR U11719 ( .A(a[2343]), .B(c2343), .Z(n7031) );
XOR U11720 ( .A(c2344), .B(n7032), .Z(c2345) );
ANDN U11721 ( .B(n7033), .A(n7034), .Z(n7032) );
XOR U11722 ( .A(c2344), .B(b[2344]), .Z(n7033) );
XNOR U11723 ( .A(b[2344]), .B(n7034), .Z(c[2344]) );
XNOR U11724 ( .A(a[2344]), .B(c2344), .Z(n7034) );
XOR U11725 ( .A(c2345), .B(n7035), .Z(c2346) );
ANDN U11726 ( .B(n7036), .A(n7037), .Z(n7035) );
XOR U11727 ( .A(c2345), .B(b[2345]), .Z(n7036) );
XNOR U11728 ( .A(b[2345]), .B(n7037), .Z(c[2345]) );
XNOR U11729 ( .A(a[2345]), .B(c2345), .Z(n7037) );
XOR U11730 ( .A(c2346), .B(n7038), .Z(c2347) );
ANDN U11731 ( .B(n7039), .A(n7040), .Z(n7038) );
XOR U11732 ( .A(c2346), .B(b[2346]), .Z(n7039) );
XNOR U11733 ( .A(b[2346]), .B(n7040), .Z(c[2346]) );
XNOR U11734 ( .A(a[2346]), .B(c2346), .Z(n7040) );
XOR U11735 ( .A(c2347), .B(n7041), .Z(c2348) );
ANDN U11736 ( .B(n7042), .A(n7043), .Z(n7041) );
XOR U11737 ( .A(c2347), .B(b[2347]), .Z(n7042) );
XNOR U11738 ( .A(b[2347]), .B(n7043), .Z(c[2347]) );
XNOR U11739 ( .A(a[2347]), .B(c2347), .Z(n7043) );
XOR U11740 ( .A(c2348), .B(n7044), .Z(c2349) );
ANDN U11741 ( .B(n7045), .A(n7046), .Z(n7044) );
XOR U11742 ( .A(c2348), .B(b[2348]), .Z(n7045) );
XNOR U11743 ( .A(b[2348]), .B(n7046), .Z(c[2348]) );
XNOR U11744 ( .A(a[2348]), .B(c2348), .Z(n7046) );
XOR U11745 ( .A(c2349), .B(n7047), .Z(c2350) );
ANDN U11746 ( .B(n7048), .A(n7049), .Z(n7047) );
XOR U11747 ( .A(c2349), .B(b[2349]), .Z(n7048) );
XNOR U11748 ( .A(b[2349]), .B(n7049), .Z(c[2349]) );
XNOR U11749 ( .A(a[2349]), .B(c2349), .Z(n7049) );
XOR U11750 ( .A(c2350), .B(n7050), .Z(c2351) );
ANDN U11751 ( .B(n7051), .A(n7052), .Z(n7050) );
XOR U11752 ( .A(c2350), .B(b[2350]), .Z(n7051) );
XNOR U11753 ( .A(b[2350]), .B(n7052), .Z(c[2350]) );
XNOR U11754 ( .A(a[2350]), .B(c2350), .Z(n7052) );
XOR U11755 ( .A(c2351), .B(n7053), .Z(c2352) );
ANDN U11756 ( .B(n7054), .A(n7055), .Z(n7053) );
XOR U11757 ( .A(c2351), .B(b[2351]), .Z(n7054) );
XNOR U11758 ( .A(b[2351]), .B(n7055), .Z(c[2351]) );
XNOR U11759 ( .A(a[2351]), .B(c2351), .Z(n7055) );
XOR U11760 ( .A(c2352), .B(n7056), .Z(c2353) );
ANDN U11761 ( .B(n7057), .A(n7058), .Z(n7056) );
XOR U11762 ( .A(c2352), .B(b[2352]), .Z(n7057) );
XNOR U11763 ( .A(b[2352]), .B(n7058), .Z(c[2352]) );
XNOR U11764 ( .A(a[2352]), .B(c2352), .Z(n7058) );
XOR U11765 ( .A(c2353), .B(n7059), .Z(c2354) );
ANDN U11766 ( .B(n7060), .A(n7061), .Z(n7059) );
XOR U11767 ( .A(c2353), .B(b[2353]), .Z(n7060) );
XNOR U11768 ( .A(b[2353]), .B(n7061), .Z(c[2353]) );
XNOR U11769 ( .A(a[2353]), .B(c2353), .Z(n7061) );
XOR U11770 ( .A(c2354), .B(n7062), .Z(c2355) );
ANDN U11771 ( .B(n7063), .A(n7064), .Z(n7062) );
XOR U11772 ( .A(c2354), .B(b[2354]), .Z(n7063) );
XNOR U11773 ( .A(b[2354]), .B(n7064), .Z(c[2354]) );
XNOR U11774 ( .A(a[2354]), .B(c2354), .Z(n7064) );
XOR U11775 ( .A(c2355), .B(n7065), .Z(c2356) );
ANDN U11776 ( .B(n7066), .A(n7067), .Z(n7065) );
XOR U11777 ( .A(c2355), .B(b[2355]), .Z(n7066) );
XNOR U11778 ( .A(b[2355]), .B(n7067), .Z(c[2355]) );
XNOR U11779 ( .A(a[2355]), .B(c2355), .Z(n7067) );
XOR U11780 ( .A(c2356), .B(n7068), .Z(c2357) );
ANDN U11781 ( .B(n7069), .A(n7070), .Z(n7068) );
XOR U11782 ( .A(c2356), .B(b[2356]), .Z(n7069) );
XNOR U11783 ( .A(b[2356]), .B(n7070), .Z(c[2356]) );
XNOR U11784 ( .A(a[2356]), .B(c2356), .Z(n7070) );
XOR U11785 ( .A(c2357), .B(n7071), .Z(c2358) );
ANDN U11786 ( .B(n7072), .A(n7073), .Z(n7071) );
XOR U11787 ( .A(c2357), .B(b[2357]), .Z(n7072) );
XNOR U11788 ( .A(b[2357]), .B(n7073), .Z(c[2357]) );
XNOR U11789 ( .A(a[2357]), .B(c2357), .Z(n7073) );
XOR U11790 ( .A(c2358), .B(n7074), .Z(c2359) );
ANDN U11791 ( .B(n7075), .A(n7076), .Z(n7074) );
XOR U11792 ( .A(c2358), .B(b[2358]), .Z(n7075) );
XNOR U11793 ( .A(b[2358]), .B(n7076), .Z(c[2358]) );
XNOR U11794 ( .A(a[2358]), .B(c2358), .Z(n7076) );
XOR U11795 ( .A(c2359), .B(n7077), .Z(c2360) );
ANDN U11796 ( .B(n7078), .A(n7079), .Z(n7077) );
XOR U11797 ( .A(c2359), .B(b[2359]), .Z(n7078) );
XNOR U11798 ( .A(b[2359]), .B(n7079), .Z(c[2359]) );
XNOR U11799 ( .A(a[2359]), .B(c2359), .Z(n7079) );
XOR U11800 ( .A(c2360), .B(n7080), .Z(c2361) );
ANDN U11801 ( .B(n7081), .A(n7082), .Z(n7080) );
XOR U11802 ( .A(c2360), .B(b[2360]), .Z(n7081) );
XNOR U11803 ( .A(b[2360]), .B(n7082), .Z(c[2360]) );
XNOR U11804 ( .A(a[2360]), .B(c2360), .Z(n7082) );
XOR U11805 ( .A(c2361), .B(n7083), .Z(c2362) );
ANDN U11806 ( .B(n7084), .A(n7085), .Z(n7083) );
XOR U11807 ( .A(c2361), .B(b[2361]), .Z(n7084) );
XNOR U11808 ( .A(b[2361]), .B(n7085), .Z(c[2361]) );
XNOR U11809 ( .A(a[2361]), .B(c2361), .Z(n7085) );
XOR U11810 ( .A(c2362), .B(n7086), .Z(c2363) );
ANDN U11811 ( .B(n7087), .A(n7088), .Z(n7086) );
XOR U11812 ( .A(c2362), .B(b[2362]), .Z(n7087) );
XNOR U11813 ( .A(b[2362]), .B(n7088), .Z(c[2362]) );
XNOR U11814 ( .A(a[2362]), .B(c2362), .Z(n7088) );
XOR U11815 ( .A(c2363), .B(n7089), .Z(c2364) );
ANDN U11816 ( .B(n7090), .A(n7091), .Z(n7089) );
XOR U11817 ( .A(c2363), .B(b[2363]), .Z(n7090) );
XNOR U11818 ( .A(b[2363]), .B(n7091), .Z(c[2363]) );
XNOR U11819 ( .A(a[2363]), .B(c2363), .Z(n7091) );
XOR U11820 ( .A(c2364), .B(n7092), .Z(c2365) );
ANDN U11821 ( .B(n7093), .A(n7094), .Z(n7092) );
XOR U11822 ( .A(c2364), .B(b[2364]), .Z(n7093) );
XNOR U11823 ( .A(b[2364]), .B(n7094), .Z(c[2364]) );
XNOR U11824 ( .A(a[2364]), .B(c2364), .Z(n7094) );
XOR U11825 ( .A(c2365), .B(n7095), .Z(c2366) );
ANDN U11826 ( .B(n7096), .A(n7097), .Z(n7095) );
XOR U11827 ( .A(c2365), .B(b[2365]), .Z(n7096) );
XNOR U11828 ( .A(b[2365]), .B(n7097), .Z(c[2365]) );
XNOR U11829 ( .A(a[2365]), .B(c2365), .Z(n7097) );
XOR U11830 ( .A(c2366), .B(n7098), .Z(c2367) );
ANDN U11831 ( .B(n7099), .A(n7100), .Z(n7098) );
XOR U11832 ( .A(c2366), .B(b[2366]), .Z(n7099) );
XNOR U11833 ( .A(b[2366]), .B(n7100), .Z(c[2366]) );
XNOR U11834 ( .A(a[2366]), .B(c2366), .Z(n7100) );
XOR U11835 ( .A(c2367), .B(n7101), .Z(c2368) );
ANDN U11836 ( .B(n7102), .A(n7103), .Z(n7101) );
XOR U11837 ( .A(c2367), .B(b[2367]), .Z(n7102) );
XNOR U11838 ( .A(b[2367]), .B(n7103), .Z(c[2367]) );
XNOR U11839 ( .A(a[2367]), .B(c2367), .Z(n7103) );
XOR U11840 ( .A(c2368), .B(n7104), .Z(c2369) );
ANDN U11841 ( .B(n7105), .A(n7106), .Z(n7104) );
XOR U11842 ( .A(c2368), .B(b[2368]), .Z(n7105) );
XNOR U11843 ( .A(b[2368]), .B(n7106), .Z(c[2368]) );
XNOR U11844 ( .A(a[2368]), .B(c2368), .Z(n7106) );
XOR U11845 ( .A(c2369), .B(n7107), .Z(c2370) );
ANDN U11846 ( .B(n7108), .A(n7109), .Z(n7107) );
XOR U11847 ( .A(c2369), .B(b[2369]), .Z(n7108) );
XNOR U11848 ( .A(b[2369]), .B(n7109), .Z(c[2369]) );
XNOR U11849 ( .A(a[2369]), .B(c2369), .Z(n7109) );
XOR U11850 ( .A(c2370), .B(n7110), .Z(c2371) );
ANDN U11851 ( .B(n7111), .A(n7112), .Z(n7110) );
XOR U11852 ( .A(c2370), .B(b[2370]), .Z(n7111) );
XNOR U11853 ( .A(b[2370]), .B(n7112), .Z(c[2370]) );
XNOR U11854 ( .A(a[2370]), .B(c2370), .Z(n7112) );
XOR U11855 ( .A(c2371), .B(n7113), .Z(c2372) );
ANDN U11856 ( .B(n7114), .A(n7115), .Z(n7113) );
XOR U11857 ( .A(c2371), .B(b[2371]), .Z(n7114) );
XNOR U11858 ( .A(b[2371]), .B(n7115), .Z(c[2371]) );
XNOR U11859 ( .A(a[2371]), .B(c2371), .Z(n7115) );
XOR U11860 ( .A(c2372), .B(n7116), .Z(c2373) );
ANDN U11861 ( .B(n7117), .A(n7118), .Z(n7116) );
XOR U11862 ( .A(c2372), .B(b[2372]), .Z(n7117) );
XNOR U11863 ( .A(b[2372]), .B(n7118), .Z(c[2372]) );
XNOR U11864 ( .A(a[2372]), .B(c2372), .Z(n7118) );
XOR U11865 ( .A(c2373), .B(n7119), .Z(c2374) );
ANDN U11866 ( .B(n7120), .A(n7121), .Z(n7119) );
XOR U11867 ( .A(c2373), .B(b[2373]), .Z(n7120) );
XNOR U11868 ( .A(b[2373]), .B(n7121), .Z(c[2373]) );
XNOR U11869 ( .A(a[2373]), .B(c2373), .Z(n7121) );
XOR U11870 ( .A(c2374), .B(n7122), .Z(c2375) );
ANDN U11871 ( .B(n7123), .A(n7124), .Z(n7122) );
XOR U11872 ( .A(c2374), .B(b[2374]), .Z(n7123) );
XNOR U11873 ( .A(b[2374]), .B(n7124), .Z(c[2374]) );
XNOR U11874 ( .A(a[2374]), .B(c2374), .Z(n7124) );
XOR U11875 ( .A(c2375), .B(n7125), .Z(c2376) );
ANDN U11876 ( .B(n7126), .A(n7127), .Z(n7125) );
XOR U11877 ( .A(c2375), .B(b[2375]), .Z(n7126) );
XNOR U11878 ( .A(b[2375]), .B(n7127), .Z(c[2375]) );
XNOR U11879 ( .A(a[2375]), .B(c2375), .Z(n7127) );
XOR U11880 ( .A(c2376), .B(n7128), .Z(c2377) );
ANDN U11881 ( .B(n7129), .A(n7130), .Z(n7128) );
XOR U11882 ( .A(c2376), .B(b[2376]), .Z(n7129) );
XNOR U11883 ( .A(b[2376]), .B(n7130), .Z(c[2376]) );
XNOR U11884 ( .A(a[2376]), .B(c2376), .Z(n7130) );
XOR U11885 ( .A(c2377), .B(n7131), .Z(c2378) );
ANDN U11886 ( .B(n7132), .A(n7133), .Z(n7131) );
XOR U11887 ( .A(c2377), .B(b[2377]), .Z(n7132) );
XNOR U11888 ( .A(b[2377]), .B(n7133), .Z(c[2377]) );
XNOR U11889 ( .A(a[2377]), .B(c2377), .Z(n7133) );
XOR U11890 ( .A(c2378), .B(n7134), .Z(c2379) );
ANDN U11891 ( .B(n7135), .A(n7136), .Z(n7134) );
XOR U11892 ( .A(c2378), .B(b[2378]), .Z(n7135) );
XNOR U11893 ( .A(b[2378]), .B(n7136), .Z(c[2378]) );
XNOR U11894 ( .A(a[2378]), .B(c2378), .Z(n7136) );
XOR U11895 ( .A(c2379), .B(n7137), .Z(c2380) );
ANDN U11896 ( .B(n7138), .A(n7139), .Z(n7137) );
XOR U11897 ( .A(c2379), .B(b[2379]), .Z(n7138) );
XNOR U11898 ( .A(b[2379]), .B(n7139), .Z(c[2379]) );
XNOR U11899 ( .A(a[2379]), .B(c2379), .Z(n7139) );
XOR U11900 ( .A(c2380), .B(n7140), .Z(c2381) );
ANDN U11901 ( .B(n7141), .A(n7142), .Z(n7140) );
XOR U11902 ( .A(c2380), .B(b[2380]), .Z(n7141) );
XNOR U11903 ( .A(b[2380]), .B(n7142), .Z(c[2380]) );
XNOR U11904 ( .A(a[2380]), .B(c2380), .Z(n7142) );
XOR U11905 ( .A(c2381), .B(n7143), .Z(c2382) );
ANDN U11906 ( .B(n7144), .A(n7145), .Z(n7143) );
XOR U11907 ( .A(c2381), .B(b[2381]), .Z(n7144) );
XNOR U11908 ( .A(b[2381]), .B(n7145), .Z(c[2381]) );
XNOR U11909 ( .A(a[2381]), .B(c2381), .Z(n7145) );
XOR U11910 ( .A(c2382), .B(n7146), .Z(c2383) );
ANDN U11911 ( .B(n7147), .A(n7148), .Z(n7146) );
XOR U11912 ( .A(c2382), .B(b[2382]), .Z(n7147) );
XNOR U11913 ( .A(b[2382]), .B(n7148), .Z(c[2382]) );
XNOR U11914 ( .A(a[2382]), .B(c2382), .Z(n7148) );
XOR U11915 ( .A(c2383), .B(n7149), .Z(c2384) );
ANDN U11916 ( .B(n7150), .A(n7151), .Z(n7149) );
XOR U11917 ( .A(c2383), .B(b[2383]), .Z(n7150) );
XNOR U11918 ( .A(b[2383]), .B(n7151), .Z(c[2383]) );
XNOR U11919 ( .A(a[2383]), .B(c2383), .Z(n7151) );
XOR U11920 ( .A(c2384), .B(n7152), .Z(c2385) );
ANDN U11921 ( .B(n7153), .A(n7154), .Z(n7152) );
XOR U11922 ( .A(c2384), .B(b[2384]), .Z(n7153) );
XNOR U11923 ( .A(b[2384]), .B(n7154), .Z(c[2384]) );
XNOR U11924 ( .A(a[2384]), .B(c2384), .Z(n7154) );
XOR U11925 ( .A(c2385), .B(n7155), .Z(c2386) );
ANDN U11926 ( .B(n7156), .A(n7157), .Z(n7155) );
XOR U11927 ( .A(c2385), .B(b[2385]), .Z(n7156) );
XNOR U11928 ( .A(b[2385]), .B(n7157), .Z(c[2385]) );
XNOR U11929 ( .A(a[2385]), .B(c2385), .Z(n7157) );
XOR U11930 ( .A(c2386), .B(n7158), .Z(c2387) );
ANDN U11931 ( .B(n7159), .A(n7160), .Z(n7158) );
XOR U11932 ( .A(c2386), .B(b[2386]), .Z(n7159) );
XNOR U11933 ( .A(b[2386]), .B(n7160), .Z(c[2386]) );
XNOR U11934 ( .A(a[2386]), .B(c2386), .Z(n7160) );
XOR U11935 ( .A(c2387), .B(n7161), .Z(c2388) );
ANDN U11936 ( .B(n7162), .A(n7163), .Z(n7161) );
XOR U11937 ( .A(c2387), .B(b[2387]), .Z(n7162) );
XNOR U11938 ( .A(b[2387]), .B(n7163), .Z(c[2387]) );
XNOR U11939 ( .A(a[2387]), .B(c2387), .Z(n7163) );
XOR U11940 ( .A(c2388), .B(n7164), .Z(c2389) );
ANDN U11941 ( .B(n7165), .A(n7166), .Z(n7164) );
XOR U11942 ( .A(c2388), .B(b[2388]), .Z(n7165) );
XNOR U11943 ( .A(b[2388]), .B(n7166), .Z(c[2388]) );
XNOR U11944 ( .A(a[2388]), .B(c2388), .Z(n7166) );
XOR U11945 ( .A(c2389), .B(n7167), .Z(c2390) );
ANDN U11946 ( .B(n7168), .A(n7169), .Z(n7167) );
XOR U11947 ( .A(c2389), .B(b[2389]), .Z(n7168) );
XNOR U11948 ( .A(b[2389]), .B(n7169), .Z(c[2389]) );
XNOR U11949 ( .A(a[2389]), .B(c2389), .Z(n7169) );
XOR U11950 ( .A(c2390), .B(n7170), .Z(c2391) );
ANDN U11951 ( .B(n7171), .A(n7172), .Z(n7170) );
XOR U11952 ( .A(c2390), .B(b[2390]), .Z(n7171) );
XNOR U11953 ( .A(b[2390]), .B(n7172), .Z(c[2390]) );
XNOR U11954 ( .A(a[2390]), .B(c2390), .Z(n7172) );
XOR U11955 ( .A(c2391), .B(n7173), .Z(c2392) );
ANDN U11956 ( .B(n7174), .A(n7175), .Z(n7173) );
XOR U11957 ( .A(c2391), .B(b[2391]), .Z(n7174) );
XNOR U11958 ( .A(b[2391]), .B(n7175), .Z(c[2391]) );
XNOR U11959 ( .A(a[2391]), .B(c2391), .Z(n7175) );
XOR U11960 ( .A(c2392), .B(n7176), .Z(c2393) );
ANDN U11961 ( .B(n7177), .A(n7178), .Z(n7176) );
XOR U11962 ( .A(c2392), .B(b[2392]), .Z(n7177) );
XNOR U11963 ( .A(b[2392]), .B(n7178), .Z(c[2392]) );
XNOR U11964 ( .A(a[2392]), .B(c2392), .Z(n7178) );
XOR U11965 ( .A(c2393), .B(n7179), .Z(c2394) );
ANDN U11966 ( .B(n7180), .A(n7181), .Z(n7179) );
XOR U11967 ( .A(c2393), .B(b[2393]), .Z(n7180) );
XNOR U11968 ( .A(b[2393]), .B(n7181), .Z(c[2393]) );
XNOR U11969 ( .A(a[2393]), .B(c2393), .Z(n7181) );
XOR U11970 ( .A(c2394), .B(n7182), .Z(c2395) );
ANDN U11971 ( .B(n7183), .A(n7184), .Z(n7182) );
XOR U11972 ( .A(c2394), .B(b[2394]), .Z(n7183) );
XNOR U11973 ( .A(b[2394]), .B(n7184), .Z(c[2394]) );
XNOR U11974 ( .A(a[2394]), .B(c2394), .Z(n7184) );
XOR U11975 ( .A(c2395), .B(n7185), .Z(c2396) );
ANDN U11976 ( .B(n7186), .A(n7187), .Z(n7185) );
XOR U11977 ( .A(c2395), .B(b[2395]), .Z(n7186) );
XNOR U11978 ( .A(b[2395]), .B(n7187), .Z(c[2395]) );
XNOR U11979 ( .A(a[2395]), .B(c2395), .Z(n7187) );
XOR U11980 ( .A(c2396), .B(n7188), .Z(c2397) );
ANDN U11981 ( .B(n7189), .A(n7190), .Z(n7188) );
XOR U11982 ( .A(c2396), .B(b[2396]), .Z(n7189) );
XNOR U11983 ( .A(b[2396]), .B(n7190), .Z(c[2396]) );
XNOR U11984 ( .A(a[2396]), .B(c2396), .Z(n7190) );
XOR U11985 ( .A(c2397), .B(n7191), .Z(c2398) );
ANDN U11986 ( .B(n7192), .A(n7193), .Z(n7191) );
XOR U11987 ( .A(c2397), .B(b[2397]), .Z(n7192) );
XNOR U11988 ( .A(b[2397]), .B(n7193), .Z(c[2397]) );
XNOR U11989 ( .A(a[2397]), .B(c2397), .Z(n7193) );
XOR U11990 ( .A(c2398), .B(n7194), .Z(c2399) );
ANDN U11991 ( .B(n7195), .A(n7196), .Z(n7194) );
XOR U11992 ( .A(c2398), .B(b[2398]), .Z(n7195) );
XNOR U11993 ( .A(b[2398]), .B(n7196), .Z(c[2398]) );
XNOR U11994 ( .A(a[2398]), .B(c2398), .Z(n7196) );
XOR U11995 ( .A(c2399), .B(n7197), .Z(c2400) );
ANDN U11996 ( .B(n7198), .A(n7199), .Z(n7197) );
XOR U11997 ( .A(c2399), .B(b[2399]), .Z(n7198) );
XNOR U11998 ( .A(b[2399]), .B(n7199), .Z(c[2399]) );
XNOR U11999 ( .A(a[2399]), .B(c2399), .Z(n7199) );
XOR U12000 ( .A(c2400), .B(n7200), .Z(c2401) );
ANDN U12001 ( .B(n7201), .A(n7202), .Z(n7200) );
XOR U12002 ( .A(c2400), .B(b[2400]), .Z(n7201) );
XNOR U12003 ( .A(b[2400]), .B(n7202), .Z(c[2400]) );
XNOR U12004 ( .A(a[2400]), .B(c2400), .Z(n7202) );
XOR U12005 ( .A(c2401), .B(n7203), .Z(c2402) );
ANDN U12006 ( .B(n7204), .A(n7205), .Z(n7203) );
XOR U12007 ( .A(c2401), .B(b[2401]), .Z(n7204) );
XNOR U12008 ( .A(b[2401]), .B(n7205), .Z(c[2401]) );
XNOR U12009 ( .A(a[2401]), .B(c2401), .Z(n7205) );
XOR U12010 ( .A(c2402), .B(n7206), .Z(c2403) );
ANDN U12011 ( .B(n7207), .A(n7208), .Z(n7206) );
XOR U12012 ( .A(c2402), .B(b[2402]), .Z(n7207) );
XNOR U12013 ( .A(b[2402]), .B(n7208), .Z(c[2402]) );
XNOR U12014 ( .A(a[2402]), .B(c2402), .Z(n7208) );
XOR U12015 ( .A(c2403), .B(n7209), .Z(c2404) );
ANDN U12016 ( .B(n7210), .A(n7211), .Z(n7209) );
XOR U12017 ( .A(c2403), .B(b[2403]), .Z(n7210) );
XNOR U12018 ( .A(b[2403]), .B(n7211), .Z(c[2403]) );
XNOR U12019 ( .A(a[2403]), .B(c2403), .Z(n7211) );
XOR U12020 ( .A(c2404), .B(n7212), .Z(c2405) );
ANDN U12021 ( .B(n7213), .A(n7214), .Z(n7212) );
XOR U12022 ( .A(c2404), .B(b[2404]), .Z(n7213) );
XNOR U12023 ( .A(b[2404]), .B(n7214), .Z(c[2404]) );
XNOR U12024 ( .A(a[2404]), .B(c2404), .Z(n7214) );
XOR U12025 ( .A(c2405), .B(n7215), .Z(c2406) );
ANDN U12026 ( .B(n7216), .A(n7217), .Z(n7215) );
XOR U12027 ( .A(c2405), .B(b[2405]), .Z(n7216) );
XNOR U12028 ( .A(b[2405]), .B(n7217), .Z(c[2405]) );
XNOR U12029 ( .A(a[2405]), .B(c2405), .Z(n7217) );
XOR U12030 ( .A(c2406), .B(n7218), .Z(c2407) );
ANDN U12031 ( .B(n7219), .A(n7220), .Z(n7218) );
XOR U12032 ( .A(c2406), .B(b[2406]), .Z(n7219) );
XNOR U12033 ( .A(b[2406]), .B(n7220), .Z(c[2406]) );
XNOR U12034 ( .A(a[2406]), .B(c2406), .Z(n7220) );
XOR U12035 ( .A(c2407), .B(n7221), .Z(c2408) );
ANDN U12036 ( .B(n7222), .A(n7223), .Z(n7221) );
XOR U12037 ( .A(c2407), .B(b[2407]), .Z(n7222) );
XNOR U12038 ( .A(b[2407]), .B(n7223), .Z(c[2407]) );
XNOR U12039 ( .A(a[2407]), .B(c2407), .Z(n7223) );
XOR U12040 ( .A(c2408), .B(n7224), .Z(c2409) );
ANDN U12041 ( .B(n7225), .A(n7226), .Z(n7224) );
XOR U12042 ( .A(c2408), .B(b[2408]), .Z(n7225) );
XNOR U12043 ( .A(b[2408]), .B(n7226), .Z(c[2408]) );
XNOR U12044 ( .A(a[2408]), .B(c2408), .Z(n7226) );
XOR U12045 ( .A(c2409), .B(n7227), .Z(c2410) );
ANDN U12046 ( .B(n7228), .A(n7229), .Z(n7227) );
XOR U12047 ( .A(c2409), .B(b[2409]), .Z(n7228) );
XNOR U12048 ( .A(b[2409]), .B(n7229), .Z(c[2409]) );
XNOR U12049 ( .A(a[2409]), .B(c2409), .Z(n7229) );
XOR U12050 ( .A(c2410), .B(n7230), .Z(c2411) );
ANDN U12051 ( .B(n7231), .A(n7232), .Z(n7230) );
XOR U12052 ( .A(c2410), .B(b[2410]), .Z(n7231) );
XNOR U12053 ( .A(b[2410]), .B(n7232), .Z(c[2410]) );
XNOR U12054 ( .A(a[2410]), .B(c2410), .Z(n7232) );
XOR U12055 ( .A(c2411), .B(n7233), .Z(c2412) );
ANDN U12056 ( .B(n7234), .A(n7235), .Z(n7233) );
XOR U12057 ( .A(c2411), .B(b[2411]), .Z(n7234) );
XNOR U12058 ( .A(b[2411]), .B(n7235), .Z(c[2411]) );
XNOR U12059 ( .A(a[2411]), .B(c2411), .Z(n7235) );
XOR U12060 ( .A(c2412), .B(n7236), .Z(c2413) );
ANDN U12061 ( .B(n7237), .A(n7238), .Z(n7236) );
XOR U12062 ( .A(c2412), .B(b[2412]), .Z(n7237) );
XNOR U12063 ( .A(b[2412]), .B(n7238), .Z(c[2412]) );
XNOR U12064 ( .A(a[2412]), .B(c2412), .Z(n7238) );
XOR U12065 ( .A(c2413), .B(n7239), .Z(c2414) );
ANDN U12066 ( .B(n7240), .A(n7241), .Z(n7239) );
XOR U12067 ( .A(c2413), .B(b[2413]), .Z(n7240) );
XNOR U12068 ( .A(b[2413]), .B(n7241), .Z(c[2413]) );
XNOR U12069 ( .A(a[2413]), .B(c2413), .Z(n7241) );
XOR U12070 ( .A(c2414), .B(n7242), .Z(c2415) );
ANDN U12071 ( .B(n7243), .A(n7244), .Z(n7242) );
XOR U12072 ( .A(c2414), .B(b[2414]), .Z(n7243) );
XNOR U12073 ( .A(b[2414]), .B(n7244), .Z(c[2414]) );
XNOR U12074 ( .A(a[2414]), .B(c2414), .Z(n7244) );
XOR U12075 ( .A(c2415), .B(n7245), .Z(c2416) );
ANDN U12076 ( .B(n7246), .A(n7247), .Z(n7245) );
XOR U12077 ( .A(c2415), .B(b[2415]), .Z(n7246) );
XNOR U12078 ( .A(b[2415]), .B(n7247), .Z(c[2415]) );
XNOR U12079 ( .A(a[2415]), .B(c2415), .Z(n7247) );
XOR U12080 ( .A(c2416), .B(n7248), .Z(c2417) );
ANDN U12081 ( .B(n7249), .A(n7250), .Z(n7248) );
XOR U12082 ( .A(c2416), .B(b[2416]), .Z(n7249) );
XNOR U12083 ( .A(b[2416]), .B(n7250), .Z(c[2416]) );
XNOR U12084 ( .A(a[2416]), .B(c2416), .Z(n7250) );
XOR U12085 ( .A(c2417), .B(n7251), .Z(c2418) );
ANDN U12086 ( .B(n7252), .A(n7253), .Z(n7251) );
XOR U12087 ( .A(c2417), .B(b[2417]), .Z(n7252) );
XNOR U12088 ( .A(b[2417]), .B(n7253), .Z(c[2417]) );
XNOR U12089 ( .A(a[2417]), .B(c2417), .Z(n7253) );
XOR U12090 ( .A(c2418), .B(n7254), .Z(c2419) );
ANDN U12091 ( .B(n7255), .A(n7256), .Z(n7254) );
XOR U12092 ( .A(c2418), .B(b[2418]), .Z(n7255) );
XNOR U12093 ( .A(b[2418]), .B(n7256), .Z(c[2418]) );
XNOR U12094 ( .A(a[2418]), .B(c2418), .Z(n7256) );
XOR U12095 ( .A(c2419), .B(n7257), .Z(c2420) );
ANDN U12096 ( .B(n7258), .A(n7259), .Z(n7257) );
XOR U12097 ( .A(c2419), .B(b[2419]), .Z(n7258) );
XNOR U12098 ( .A(b[2419]), .B(n7259), .Z(c[2419]) );
XNOR U12099 ( .A(a[2419]), .B(c2419), .Z(n7259) );
XOR U12100 ( .A(c2420), .B(n7260), .Z(c2421) );
ANDN U12101 ( .B(n7261), .A(n7262), .Z(n7260) );
XOR U12102 ( .A(c2420), .B(b[2420]), .Z(n7261) );
XNOR U12103 ( .A(b[2420]), .B(n7262), .Z(c[2420]) );
XNOR U12104 ( .A(a[2420]), .B(c2420), .Z(n7262) );
XOR U12105 ( .A(c2421), .B(n7263), .Z(c2422) );
ANDN U12106 ( .B(n7264), .A(n7265), .Z(n7263) );
XOR U12107 ( .A(c2421), .B(b[2421]), .Z(n7264) );
XNOR U12108 ( .A(b[2421]), .B(n7265), .Z(c[2421]) );
XNOR U12109 ( .A(a[2421]), .B(c2421), .Z(n7265) );
XOR U12110 ( .A(c2422), .B(n7266), .Z(c2423) );
ANDN U12111 ( .B(n7267), .A(n7268), .Z(n7266) );
XOR U12112 ( .A(c2422), .B(b[2422]), .Z(n7267) );
XNOR U12113 ( .A(b[2422]), .B(n7268), .Z(c[2422]) );
XNOR U12114 ( .A(a[2422]), .B(c2422), .Z(n7268) );
XOR U12115 ( .A(c2423), .B(n7269), .Z(c2424) );
ANDN U12116 ( .B(n7270), .A(n7271), .Z(n7269) );
XOR U12117 ( .A(c2423), .B(b[2423]), .Z(n7270) );
XNOR U12118 ( .A(b[2423]), .B(n7271), .Z(c[2423]) );
XNOR U12119 ( .A(a[2423]), .B(c2423), .Z(n7271) );
XOR U12120 ( .A(c2424), .B(n7272), .Z(c2425) );
ANDN U12121 ( .B(n7273), .A(n7274), .Z(n7272) );
XOR U12122 ( .A(c2424), .B(b[2424]), .Z(n7273) );
XNOR U12123 ( .A(b[2424]), .B(n7274), .Z(c[2424]) );
XNOR U12124 ( .A(a[2424]), .B(c2424), .Z(n7274) );
XOR U12125 ( .A(c2425), .B(n7275), .Z(c2426) );
ANDN U12126 ( .B(n7276), .A(n7277), .Z(n7275) );
XOR U12127 ( .A(c2425), .B(b[2425]), .Z(n7276) );
XNOR U12128 ( .A(b[2425]), .B(n7277), .Z(c[2425]) );
XNOR U12129 ( .A(a[2425]), .B(c2425), .Z(n7277) );
XOR U12130 ( .A(c2426), .B(n7278), .Z(c2427) );
ANDN U12131 ( .B(n7279), .A(n7280), .Z(n7278) );
XOR U12132 ( .A(c2426), .B(b[2426]), .Z(n7279) );
XNOR U12133 ( .A(b[2426]), .B(n7280), .Z(c[2426]) );
XNOR U12134 ( .A(a[2426]), .B(c2426), .Z(n7280) );
XOR U12135 ( .A(c2427), .B(n7281), .Z(c2428) );
ANDN U12136 ( .B(n7282), .A(n7283), .Z(n7281) );
XOR U12137 ( .A(c2427), .B(b[2427]), .Z(n7282) );
XNOR U12138 ( .A(b[2427]), .B(n7283), .Z(c[2427]) );
XNOR U12139 ( .A(a[2427]), .B(c2427), .Z(n7283) );
XOR U12140 ( .A(c2428), .B(n7284), .Z(c2429) );
ANDN U12141 ( .B(n7285), .A(n7286), .Z(n7284) );
XOR U12142 ( .A(c2428), .B(b[2428]), .Z(n7285) );
XNOR U12143 ( .A(b[2428]), .B(n7286), .Z(c[2428]) );
XNOR U12144 ( .A(a[2428]), .B(c2428), .Z(n7286) );
XOR U12145 ( .A(c2429), .B(n7287), .Z(c2430) );
ANDN U12146 ( .B(n7288), .A(n7289), .Z(n7287) );
XOR U12147 ( .A(c2429), .B(b[2429]), .Z(n7288) );
XNOR U12148 ( .A(b[2429]), .B(n7289), .Z(c[2429]) );
XNOR U12149 ( .A(a[2429]), .B(c2429), .Z(n7289) );
XOR U12150 ( .A(c2430), .B(n7290), .Z(c2431) );
ANDN U12151 ( .B(n7291), .A(n7292), .Z(n7290) );
XOR U12152 ( .A(c2430), .B(b[2430]), .Z(n7291) );
XNOR U12153 ( .A(b[2430]), .B(n7292), .Z(c[2430]) );
XNOR U12154 ( .A(a[2430]), .B(c2430), .Z(n7292) );
XOR U12155 ( .A(c2431), .B(n7293), .Z(c2432) );
ANDN U12156 ( .B(n7294), .A(n7295), .Z(n7293) );
XOR U12157 ( .A(c2431), .B(b[2431]), .Z(n7294) );
XNOR U12158 ( .A(b[2431]), .B(n7295), .Z(c[2431]) );
XNOR U12159 ( .A(a[2431]), .B(c2431), .Z(n7295) );
XOR U12160 ( .A(c2432), .B(n7296), .Z(c2433) );
ANDN U12161 ( .B(n7297), .A(n7298), .Z(n7296) );
XOR U12162 ( .A(c2432), .B(b[2432]), .Z(n7297) );
XNOR U12163 ( .A(b[2432]), .B(n7298), .Z(c[2432]) );
XNOR U12164 ( .A(a[2432]), .B(c2432), .Z(n7298) );
XOR U12165 ( .A(c2433), .B(n7299), .Z(c2434) );
ANDN U12166 ( .B(n7300), .A(n7301), .Z(n7299) );
XOR U12167 ( .A(c2433), .B(b[2433]), .Z(n7300) );
XNOR U12168 ( .A(b[2433]), .B(n7301), .Z(c[2433]) );
XNOR U12169 ( .A(a[2433]), .B(c2433), .Z(n7301) );
XOR U12170 ( .A(c2434), .B(n7302), .Z(c2435) );
ANDN U12171 ( .B(n7303), .A(n7304), .Z(n7302) );
XOR U12172 ( .A(c2434), .B(b[2434]), .Z(n7303) );
XNOR U12173 ( .A(b[2434]), .B(n7304), .Z(c[2434]) );
XNOR U12174 ( .A(a[2434]), .B(c2434), .Z(n7304) );
XOR U12175 ( .A(c2435), .B(n7305), .Z(c2436) );
ANDN U12176 ( .B(n7306), .A(n7307), .Z(n7305) );
XOR U12177 ( .A(c2435), .B(b[2435]), .Z(n7306) );
XNOR U12178 ( .A(b[2435]), .B(n7307), .Z(c[2435]) );
XNOR U12179 ( .A(a[2435]), .B(c2435), .Z(n7307) );
XOR U12180 ( .A(c2436), .B(n7308), .Z(c2437) );
ANDN U12181 ( .B(n7309), .A(n7310), .Z(n7308) );
XOR U12182 ( .A(c2436), .B(b[2436]), .Z(n7309) );
XNOR U12183 ( .A(b[2436]), .B(n7310), .Z(c[2436]) );
XNOR U12184 ( .A(a[2436]), .B(c2436), .Z(n7310) );
XOR U12185 ( .A(c2437), .B(n7311), .Z(c2438) );
ANDN U12186 ( .B(n7312), .A(n7313), .Z(n7311) );
XOR U12187 ( .A(c2437), .B(b[2437]), .Z(n7312) );
XNOR U12188 ( .A(b[2437]), .B(n7313), .Z(c[2437]) );
XNOR U12189 ( .A(a[2437]), .B(c2437), .Z(n7313) );
XOR U12190 ( .A(c2438), .B(n7314), .Z(c2439) );
ANDN U12191 ( .B(n7315), .A(n7316), .Z(n7314) );
XOR U12192 ( .A(c2438), .B(b[2438]), .Z(n7315) );
XNOR U12193 ( .A(b[2438]), .B(n7316), .Z(c[2438]) );
XNOR U12194 ( .A(a[2438]), .B(c2438), .Z(n7316) );
XOR U12195 ( .A(c2439), .B(n7317), .Z(c2440) );
ANDN U12196 ( .B(n7318), .A(n7319), .Z(n7317) );
XOR U12197 ( .A(c2439), .B(b[2439]), .Z(n7318) );
XNOR U12198 ( .A(b[2439]), .B(n7319), .Z(c[2439]) );
XNOR U12199 ( .A(a[2439]), .B(c2439), .Z(n7319) );
XOR U12200 ( .A(c2440), .B(n7320), .Z(c2441) );
ANDN U12201 ( .B(n7321), .A(n7322), .Z(n7320) );
XOR U12202 ( .A(c2440), .B(b[2440]), .Z(n7321) );
XNOR U12203 ( .A(b[2440]), .B(n7322), .Z(c[2440]) );
XNOR U12204 ( .A(a[2440]), .B(c2440), .Z(n7322) );
XOR U12205 ( .A(c2441), .B(n7323), .Z(c2442) );
ANDN U12206 ( .B(n7324), .A(n7325), .Z(n7323) );
XOR U12207 ( .A(c2441), .B(b[2441]), .Z(n7324) );
XNOR U12208 ( .A(b[2441]), .B(n7325), .Z(c[2441]) );
XNOR U12209 ( .A(a[2441]), .B(c2441), .Z(n7325) );
XOR U12210 ( .A(c2442), .B(n7326), .Z(c2443) );
ANDN U12211 ( .B(n7327), .A(n7328), .Z(n7326) );
XOR U12212 ( .A(c2442), .B(b[2442]), .Z(n7327) );
XNOR U12213 ( .A(b[2442]), .B(n7328), .Z(c[2442]) );
XNOR U12214 ( .A(a[2442]), .B(c2442), .Z(n7328) );
XOR U12215 ( .A(c2443), .B(n7329), .Z(c2444) );
ANDN U12216 ( .B(n7330), .A(n7331), .Z(n7329) );
XOR U12217 ( .A(c2443), .B(b[2443]), .Z(n7330) );
XNOR U12218 ( .A(b[2443]), .B(n7331), .Z(c[2443]) );
XNOR U12219 ( .A(a[2443]), .B(c2443), .Z(n7331) );
XOR U12220 ( .A(c2444), .B(n7332), .Z(c2445) );
ANDN U12221 ( .B(n7333), .A(n7334), .Z(n7332) );
XOR U12222 ( .A(c2444), .B(b[2444]), .Z(n7333) );
XNOR U12223 ( .A(b[2444]), .B(n7334), .Z(c[2444]) );
XNOR U12224 ( .A(a[2444]), .B(c2444), .Z(n7334) );
XOR U12225 ( .A(c2445), .B(n7335), .Z(c2446) );
ANDN U12226 ( .B(n7336), .A(n7337), .Z(n7335) );
XOR U12227 ( .A(c2445), .B(b[2445]), .Z(n7336) );
XNOR U12228 ( .A(b[2445]), .B(n7337), .Z(c[2445]) );
XNOR U12229 ( .A(a[2445]), .B(c2445), .Z(n7337) );
XOR U12230 ( .A(c2446), .B(n7338), .Z(c2447) );
ANDN U12231 ( .B(n7339), .A(n7340), .Z(n7338) );
XOR U12232 ( .A(c2446), .B(b[2446]), .Z(n7339) );
XNOR U12233 ( .A(b[2446]), .B(n7340), .Z(c[2446]) );
XNOR U12234 ( .A(a[2446]), .B(c2446), .Z(n7340) );
XOR U12235 ( .A(c2447), .B(n7341), .Z(c2448) );
ANDN U12236 ( .B(n7342), .A(n7343), .Z(n7341) );
XOR U12237 ( .A(c2447), .B(b[2447]), .Z(n7342) );
XNOR U12238 ( .A(b[2447]), .B(n7343), .Z(c[2447]) );
XNOR U12239 ( .A(a[2447]), .B(c2447), .Z(n7343) );
XOR U12240 ( .A(c2448), .B(n7344), .Z(c2449) );
ANDN U12241 ( .B(n7345), .A(n7346), .Z(n7344) );
XOR U12242 ( .A(c2448), .B(b[2448]), .Z(n7345) );
XNOR U12243 ( .A(b[2448]), .B(n7346), .Z(c[2448]) );
XNOR U12244 ( .A(a[2448]), .B(c2448), .Z(n7346) );
XOR U12245 ( .A(c2449), .B(n7347), .Z(c2450) );
ANDN U12246 ( .B(n7348), .A(n7349), .Z(n7347) );
XOR U12247 ( .A(c2449), .B(b[2449]), .Z(n7348) );
XNOR U12248 ( .A(b[2449]), .B(n7349), .Z(c[2449]) );
XNOR U12249 ( .A(a[2449]), .B(c2449), .Z(n7349) );
XOR U12250 ( .A(c2450), .B(n7350), .Z(c2451) );
ANDN U12251 ( .B(n7351), .A(n7352), .Z(n7350) );
XOR U12252 ( .A(c2450), .B(b[2450]), .Z(n7351) );
XNOR U12253 ( .A(b[2450]), .B(n7352), .Z(c[2450]) );
XNOR U12254 ( .A(a[2450]), .B(c2450), .Z(n7352) );
XOR U12255 ( .A(c2451), .B(n7353), .Z(c2452) );
ANDN U12256 ( .B(n7354), .A(n7355), .Z(n7353) );
XOR U12257 ( .A(c2451), .B(b[2451]), .Z(n7354) );
XNOR U12258 ( .A(b[2451]), .B(n7355), .Z(c[2451]) );
XNOR U12259 ( .A(a[2451]), .B(c2451), .Z(n7355) );
XOR U12260 ( .A(c2452), .B(n7356), .Z(c2453) );
ANDN U12261 ( .B(n7357), .A(n7358), .Z(n7356) );
XOR U12262 ( .A(c2452), .B(b[2452]), .Z(n7357) );
XNOR U12263 ( .A(b[2452]), .B(n7358), .Z(c[2452]) );
XNOR U12264 ( .A(a[2452]), .B(c2452), .Z(n7358) );
XOR U12265 ( .A(c2453), .B(n7359), .Z(c2454) );
ANDN U12266 ( .B(n7360), .A(n7361), .Z(n7359) );
XOR U12267 ( .A(c2453), .B(b[2453]), .Z(n7360) );
XNOR U12268 ( .A(b[2453]), .B(n7361), .Z(c[2453]) );
XNOR U12269 ( .A(a[2453]), .B(c2453), .Z(n7361) );
XOR U12270 ( .A(c2454), .B(n7362), .Z(c2455) );
ANDN U12271 ( .B(n7363), .A(n7364), .Z(n7362) );
XOR U12272 ( .A(c2454), .B(b[2454]), .Z(n7363) );
XNOR U12273 ( .A(b[2454]), .B(n7364), .Z(c[2454]) );
XNOR U12274 ( .A(a[2454]), .B(c2454), .Z(n7364) );
XOR U12275 ( .A(c2455), .B(n7365), .Z(c2456) );
ANDN U12276 ( .B(n7366), .A(n7367), .Z(n7365) );
XOR U12277 ( .A(c2455), .B(b[2455]), .Z(n7366) );
XNOR U12278 ( .A(b[2455]), .B(n7367), .Z(c[2455]) );
XNOR U12279 ( .A(a[2455]), .B(c2455), .Z(n7367) );
XOR U12280 ( .A(c2456), .B(n7368), .Z(c2457) );
ANDN U12281 ( .B(n7369), .A(n7370), .Z(n7368) );
XOR U12282 ( .A(c2456), .B(b[2456]), .Z(n7369) );
XNOR U12283 ( .A(b[2456]), .B(n7370), .Z(c[2456]) );
XNOR U12284 ( .A(a[2456]), .B(c2456), .Z(n7370) );
XOR U12285 ( .A(c2457), .B(n7371), .Z(c2458) );
ANDN U12286 ( .B(n7372), .A(n7373), .Z(n7371) );
XOR U12287 ( .A(c2457), .B(b[2457]), .Z(n7372) );
XNOR U12288 ( .A(b[2457]), .B(n7373), .Z(c[2457]) );
XNOR U12289 ( .A(a[2457]), .B(c2457), .Z(n7373) );
XOR U12290 ( .A(c2458), .B(n7374), .Z(c2459) );
ANDN U12291 ( .B(n7375), .A(n7376), .Z(n7374) );
XOR U12292 ( .A(c2458), .B(b[2458]), .Z(n7375) );
XNOR U12293 ( .A(b[2458]), .B(n7376), .Z(c[2458]) );
XNOR U12294 ( .A(a[2458]), .B(c2458), .Z(n7376) );
XOR U12295 ( .A(c2459), .B(n7377), .Z(c2460) );
ANDN U12296 ( .B(n7378), .A(n7379), .Z(n7377) );
XOR U12297 ( .A(c2459), .B(b[2459]), .Z(n7378) );
XNOR U12298 ( .A(b[2459]), .B(n7379), .Z(c[2459]) );
XNOR U12299 ( .A(a[2459]), .B(c2459), .Z(n7379) );
XOR U12300 ( .A(c2460), .B(n7380), .Z(c2461) );
ANDN U12301 ( .B(n7381), .A(n7382), .Z(n7380) );
XOR U12302 ( .A(c2460), .B(b[2460]), .Z(n7381) );
XNOR U12303 ( .A(b[2460]), .B(n7382), .Z(c[2460]) );
XNOR U12304 ( .A(a[2460]), .B(c2460), .Z(n7382) );
XOR U12305 ( .A(c2461), .B(n7383), .Z(c2462) );
ANDN U12306 ( .B(n7384), .A(n7385), .Z(n7383) );
XOR U12307 ( .A(c2461), .B(b[2461]), .Z(n7384) );
XNOR U12308 ( .A(b[2461]), .B(n7385), .Z(c[2461]) );
XNOR U12309 ( .A(a[2461]), .B(c2461), .Z(n7385) );
XOR U12310 ( .A(c2462), .B(n7386), .Z(c2463) );
ANDN U12311 ( .B(n7387), .A(n7388), .Z(n7386) );
XOR U12312 ( .A(c2462), .B(b[2462]), .Z(n7387) );
XNOR U12313 ( .A(b[2462]), .B(n7388), .Z(c[2462]) );
XNOR U12314 ( .A(a[2462]), .B(c2462), .Z(n7388) );
XOR U12315 ( .A(c2463), .B(n7389), .Z(c2464) );
ANDN U12316 ( .B(n7390), .A(n7391), .Z(n7389) );
XOR U12317 ( .A(c2463), .B(b[2463]), .Z(n7390) );
XNOR U12318 ( .A(b[2463]), .B(n7391), .Z(c[2463]) );
XNOR U12319 ( .A(a[2463]), .B(c2463), .Z(n7391) );
XOR U12320 ( .A(c2464), .B(n7392), .Z(c2465) );
ANDN U12321 ( .B(n7393), .A(n7394), .Z(n7392) );
XOR U12322 ( .A(c2464), .B(b[2464]), .Z(n7393) );
XNOR U12323 ( .A(b[2464]), .B(n7394), .Z(c[2464]) );
XNOR U12324 ( .A(a[2464]), .B(c2464), .Z(n7394) );
XOR U12325 ( .A(c2465), .B(n7395), .Z(c2466) );
ANDN U12326 ( .B(n7396), .A(n7397), .Z(n7395) );
XOR U12327 ( .A(c2465), .B(b[2465]), .Z(n7396) );
XNOR U12328 ( .A(b[2465]), .B(n7397), .Z(c[2465]) );
XNOR U12329 ( .A(a[2465]), .B(c2465), .Z(n7397) );
XOR U12330 ( .A(c2466), .B(n7398), .Z(c2467) );
ANDN U12331 ( .B(n7399), .A(n7400), .Z(n7398) );
XOR U12332 ( .A(c2466), .B(b[2466]), .Z(n7399) );
XNOR U12333 ( .A(b[2466]), .B(n7400), .Z(c[2466]) );
XNOR U12334 ( .A(a[2466]), .B(c2466), .Z(n7400) );
XOR U12335 ( .A(c2467), .B(n7401), .Z(c2468) );
ANDN U12336 ( .B(n7402), .A(n7403), .Z(n7401) );
XOR U12337 ( .A(c2467), .B(b[2467]), .Z(n7402) );
XNOR U12338 ( .A(b[2467]), .B(n7403), .Z(c[2467]) );
XNOR U12339 ( .A(a[2467]), .B(c2467), .Z(n7403) );
XOR U12340 ( .A(c2468), .B(n7404), .Z(c2469) );
ANDN U12341 ( .B(n7405), .A(n7406), .Z(n7404) );
XOR U12342 ( .A(c2468), .B(b[2468]), .Z(n7405) );
XNOR U12343 ( .A(b[2468]), .B(n7406), .Z(c[2468]) );
XNOR U12344 ( .A(a[2468]), .B(c2468), .Z(n7406) );
XOR U12345 ( .A(c2469), .B(n7407), .Z(c2470) );
ANDN U12346 ( .B(n7408), .A(n7409), .Z(n7407) );
XOR U12347 ( .A(c2469), .B(b[2469]), .Z(n7408) );
XNOR U12348 ( .A(b[2469]), .B(n7409), .Z(c[2469]) );
XNOR U12349 ( .A(a[2469]), .B(c2469), .Z(n7409) );
XOR U12350 ( .A(c2470), .B(n7410), .Z(c2471) );
ANDN U12351 ( .B(n7411), .A(n7412), .Z(n7410) );
XOR U12352 ( .A(c2470), .B(b[2470]), .Z(n7411) );
XNOR U12353 ( .A(b[2470]), .B(n7412), .Z(c[2470]) );
XNOR U12354 ( .A(a[2470]), .B(c2470), .Z(n7412) );
XOR U12355 ( .A(c2471), .B(n7413), .Z(c2472) );
ANDN U12356 ( .B(n7414), .A(n7415), .Z(n7413) );
XOR U12357 ( .A(c2471), .B(b[2471]), .Z(n7414) );
XNOR U12358 ( .A(b[2471]), .B(n7415), .Z(c[2471]) );
XNOR U12359 ( .A(a[2471]), .B(c2471), .Z(n7415) );
XOR U12360 ( .A(c2472), .B(n7416), .Z(c2473) );
ANDN U12361 ( .B(n7417), .A(n7418), .Z(n7416) );
XOR U12362 ( .A(c2472), .B(b[2472]), .Z(n7417) );
XNOR U12363 ( .A(b[2472]), .B(n7418), .Z(c[2472]) );
XNOR U12364 ( .A(a[2472]), .B(c2472), .Z(n7418) );
XOR U12365 ( .A(c2473), .B(n7419), .Z(c2474) );
ANDN U12366 ( .B(n7420), .A(n7421), .Z(n7419) );
XOR U12367 ( .A(c2473), .B(b[2473]), .Z(n7420) );
XNOR U12368 ( .A(b[2473]), .B(n7421), .Z(c[2473]) );
XNOR U12369 ( .A(a[2473]), .B(c2473), .Z(n7421) );
XOR U12370 ( .A(c2474), .B(n7422), .Z(c2475) );
ANDN U12371 ( .B(n7423), .A(n7424), .Z(n7422) );
XOR U12372 ( .A(c2474), .B(b[2474]), .Z(n7423) );
XNOR U12373 ( .A(b[2474]), .B(n7424), .Z(c[2474]) );
XNOR U12374 ( .A(a[2474]), .B(c2474), .Z(n7424) );
XOR U12375 ( .A(c2475), .B(n7425), .Z(c2476) );
ANDN U12376 ( .B(n7426), .A(n7427), .Z(n7425) );
XOR U12377 ( .A(c2475), .B(b[2475]), .Z(n7426) );
XNOR U12378 ( .A(b[2475]), .B(n7427), .Z(c[2475]) );
XNOR U12379 ( .A(a[2475]), .B(c2475), .Z(n7427) );
XOR U12380 ( .A(c2476), .B(n7428), .Z(c2477) );
ANDN U12381 ( .B(n7429), .A(n7430), .Z(n7428) );
XOR U12382 ( .A(c2476), .B(b[2476]), .Z(n7429) );
XNOR U12383 ( .A(b[2476]), .B(n7430), .Z(c[2476]) );
XNOR U12384 ( .A(a[2476]), .B(c2476), .Z(n7430) );
XOR U12385 ( .A(c2477), .B(n7431), .Z(c2478) );
ANDN U12386 ( .B(n7432), .A(n7433), .Z(n7431) );
XOR U12387 ( .A(c2477), .B(b[2477]), .Z(n7432) );
XNOR U12388 ( .A(b[2477]), .B(n7433), .Z(c[2477]) );
XNOR U12389 ( .A(a[2477]), .B(c2477), .Z(n7433) );
XOR U12390 ( .A(c2478), .B(n7434), .Z(c2479) );
ANDN U12391 ( .B(n7435), .A(n7436), .Z(n7434) );
XOR U12392 ( .A(c2478), .B(b[2478]), .Z(n7435) );
XNOR U12393 ( .A(b[2478]), .B(n7436), .Z(c[2478]) );
XNOR U12394 ( .A(a[2478]), .B(c2478), .Z(n7436) );
XOR U12395 ( .A(c2479), .B(n7437), .Z(c2480) );
ANDN U12396 ( .B(n7438), .A(n7439), .Z(n7437) );
XOR U12397 ( .A(c2479), .B(b[2479]), .Z(n7438) );
XNOR U12398 ( .A(b[2479]), .B(n7439), .Z(c[2479]) );
XNOR U12399 ( .A(a[2479]), .B(c2479), .Z(n7439) );
XOR U12400 ( .A(c2480), .B(n7440), .Z(c2481) );
ANDN U12401 ( .B(n7441), .A(n7442), .Z(n7440) );
XOR U12402 ( .A(c2480), .B(b[2480]), .Z(n7441) );
XNOR U12403 ( .A(b[2480]), .B(n7442), .Z(c[2480]) );
XNOR U12404 ( .A(a[2480]), .B(c2480), .Z(n7442) );
XOR U12405 ( .A(c2481), .B(n7443), .Z(c2482) );
ANDN U12406 ( .B(n7444), .A(n7445), .Z(n7443) );
XOR U12407 ( .A(c2481), .B(b[2481]), .Z(n7444) );
XNOR U12408 ( .A(b[2481]), .B(n7445), .Z(c[2481]) );
XNOR U12409 ( .A(a[2481]), .B(c2481), .Z(n7445) );
XOR U12410 ( .A(c2482), .B(n7446), .Z(c2483) );
ANDN U12411 ( .B(n7447), .A(n7448), .Z(n7446) );
XOR U12412 ( .A(c2482), .B(b[2482]), .Z(n7447) );
XNOR U12413 ( .A(b[2482]), .B(n7448), .Z(c[2482]) );
XNOR U12414 ( .A(a[2482]), .B(c2482), .Z(n7448) );
XOR U12415 ( .A(c2483), .B(n7449), .Z(c2484) );
ANDN U12416 ( .B(n7450), .A(n7451), .Z(n7449) );
XOR U12417 ( .A(c2483), .B(b[2483]), .Z(n7450) );
XNOR U12418 ( .A(b[2483]), .B(n7451), .Z(c[2483]) );
XNOR U12419 ( .A(a[2483]), .B(c2483), .Z(n7451) );
XOR U12420 ( .A(c2484), .B(n7452), .Z(c2485) );
ANDN U12421 ( .B(n7453), .A(n7454), .Z(n7452) );
XOR U12422 ( .A(c2484), .B(b[2484]), .Z(n7453) );
XNOR U12423 ( .A(b[2484]), .B(n7454), .Z(c[2484]) );
XNOR U12424 ( .A(a[2484]), .B(c2484), .Z(n7454) );
XOR U12425 ( .A(c2485), .B(n7455), .Z(c2486) );
ANDN U12426 ( .B(n7456), .A(n7457), .Z(n7455) );
XOR U12427 ( .A(c2485), .B(b[2485]), .Z(n7456) );
XNOR U12428 ( .A(b[2485]), .B(n7457), .Z(c[2485]) );
XNOR U12429 ( .A(a[2485]), .B(c2485), .Z(n7457) );
XOR U12430 ( .A(c2486), .B(n7458), .Z(c2487) );
ANDN U12431 ( .B(n7459), .A(n7460), .Z(n7458) );
XOR U12432 ( .A(c2486), .B(b[2486]), .Z(n7459) );
XNOR U12433 ( .A(b[2486]), .B(n7460), .Z(c[2486]) );
XNOR U12434 ( .A(a[2486]), .B(c2486), .Z(n7460) );
XOR U12435 ( .A(c2487), .B(n7461), .Z(c2488) );
ANDN U12436 ( .B(n7462), .A(n7463), .Z(n7461) );
XOR U12437 ( .A(c2487), .B(b[2487]), .Z(n7462) );
XNOR U12438 ( .A(b[2487]), .B(n7463), .Z(c[2487]) );
XNOR U12439 ( .A(a[2487]), .B(c2487), .Z(n7463) );
XOR U12440 ( .A(c2488), .B(n7464), .Z(c2489) );
ANDN U12441 ( .B(n7465), .A(n7466), .Z(n7464) );
XOR U12442 ( .A(c2488), .B(b[2488]), .Z(n7465) );
XNOR U12443 ( .A(b[2488]), .B(n7466), .Z(c[2488]) );
XNOR U12444 ( .A(a[2488]), .B(c2488), .Z(n7466) );
XOR U12445 ( .A(c2489), .B(n7467), .Z(c2490) );
ANDN U12446 ( .B(n7468), .A(n7469), .Z(n7467) );
XOR U12447 ( .A(c2489), .B(b[2489]), .Z(n7468) );
XNOR U12448 ( .A(b[2489]), .B(n7469), .Z(c[2489]) );
XNOR U12449 ( .A(a[2489]), .B(c2489), .Z(n7469) );
XOR U12450 ( .A(c2490), .B(n7470), .Z(c2491) );
ANDN U12451 ( .B(n7471), .A(n7472), .Z(n7470) );
XOR U12452 ( .A(c2490), .B(b[2490]), .Z(n7471) );
XNOR U12453 ( .A(b[2490]), .B(n7472), .Z(c[2490]) );
XNOR U12454 ( .A(a[2490]), .B(c2490), .Z(n7472) );
XOR U12455 ( .A(c2491), .B(n7473), .Z(c2492) );
ANDN U12456 ( .B(n7474), .A(n7475), .Z(n7473) );
XOR U12457 ( .A(c2491), .B(b[2491]), .Z(n7474) );
XNOR U12458 ( .A(b[2491]), .B(n7475), .Z(c[2491]) );
XNOR U12459 ( .A(a[2491]), .B(c2491), .Z(n7475) );
XOR U12460 ( .A(c2492), .B(n7476), .Z(c2493) );
ANDN U12461 ( .B(n7477), .A(n7478), .Z(n7476) );
XOR U12462 ( .A(c2492), .B(b[2492]), .Z(n7477) );
XNOR U12463 ( .A(b[2492]), .B(n7478), .Z(c[2492]) );
XNOR U12464 ( .A(a[2492]), .B(c2492), .Z(n7478) );
XOR U12465 ( .A(c2493), .B(n7479), .Z(c2494) );
ANDN U12466 ( .B(n7480), .A(n7481), .Z(n7479) );
XOR U12467 ( .A(c2493), .B(b[2493]), .Z(n7480) );
XNOR U12468 ( .A(b[2493]), .B(n7481), .Z(c[2493]) );
XNOR U12469 ( .A(a[2493]), .B(c2493), .Z(n7481) );
XOR U12470 ( .A(c2494), .B(n7482), .Z(c2495) );
ANDN U12471 ( .B(n7483), .A(n7484), .Z(n7482) );
XOR U12472 ( .A(c2494), .B(b[2494]), .Z(n7483) );
XNOR U12473 ( .A(b[2494]), .B(n7484), .Z(c[2494]) );
XNOR U12474 ( .A(a[2494]), .B(c2494), .Z(n7484) );
XOR U12475 ( .A(c2495), .B(n7485), .Z(c2496) );
ANDN U12476 ( .B(n7486), .A(n7487), .Z(n7485) );
XOR U12477 ( .A(c2495), .B(b[2495]), .Z(n7486) );
XNOR U12478 ( .A(b[2495]), .B(n7487), .Z(c[2495]) );
XNOR U12479 ( .A(a[2495]), .B(c2495), .Z(n7487) );
XOR U12480 ( .A(c2496), .B(n7488), .Z(c2497) );
ANDN U12481 ( .B(n7489), .A(n7490), .Z(n7488) );
XOR U12482 ( .A(c2496), .B(b[2496]), .Z(n7489) );
XNOR U12483 ( .A(b[2496]), .B(n7490), .Z(c[2496]) );
XNOR U12484 ( .A(a[2496]), .B(c2496), .Z(n7490) );
XOR U12485 ( .A(c2497), .B(n7491), .Z(c2498) );
ANDN U12486 ( .B(n7492), .A(n7493), .Z(n7491) );
XOR U12487 ( .A(c2497), .B(b[2497]), .Z(n7492) );
XNOR U12488 ( .A(b[2497]), .B(n7493), .Z(c[2497]) );
XNOR U12489 ( .A(a[2497]), .B(c2497), .Z(n7493) );
XOR U12490 ( .A(c2498), .B(n7494), .Z(c2499) );
ANDN U12491 ( .B(n7495), .A(n7496), .Z(n7494) );
XOR U12492 ( .A(c2498), .B(b[2498]), .Z(n7495) );
XNOR U12493 ( .A(b[2498]), .B(n7496), .Z(c[2498]) );
XNOR U12494 ( .A(a[2498]), .B(c2498), .Z(n7496) );
XOR U12495 ( .A(c2499), .B(n7497), .Z(c2500) );
ANDN U12496 ( .B(n7498), .A(n7499), .Z(n7497) );
XOR U12497 ( .A(c2499), .B(b[2499]), .Z(n7498) );
XNOR U12498 ( .A(b[2499]), .B(n7499), .Z(c[2499]) );
XNOR U12499 ( .A(a[2499]), .B(c2499), .Z(n7499) );
XOR U12500 ( .A(c2500), .B(n7500), .Z(c2501) );
ANDN U12501 ( .B(n7501), .A(n7502), .Z(n7500) );
XOR U12502 ( .A(c2500), .B(b[2500]), .Z(n7501) );
XNOR U12503 ( .A(b[2500]), .B(n7502), .Z(c[2500]) );
XNOR U12504 ( .A(a[2500]), .B(c2500), .Z(n7502) );
XOR U12505 ( .A(c2501), .B(n7503), .Z(c2502) );
ANDN U12506 ( .B(n7504), .A(n7505), .Z(n7503) );
XOR U12507 ( .A(c2501), .B(b[2501]), .Z(n7504) );
XNOR U12508 ( .A(b[2501]), .B(n7505), .Z(c[2501]) );
XNOR U12509 ( .A(a[2501]), .B(c2501), .Z(n7505) );
XOR U12510 ( .A(c2502), .B(n7506), .Z(c2503) );
ANDN U12511 ( .B(n7507), .A(n7508), .Z(n7506) );
XOR U12512 ( .A(c2502), .B(b[2502]), .Z(n7507) );
XNOR U12513 ( .A(b[2502]), .B(n7508), .Z(c[2502]) );
XNOR U12514 ( .A(a[2502]), .B(c2502), .Z(n7508) );
XOR U12515 ( .A(c2503), .B(n7509), .Z(c2504) );
ANDN U12516 ( .B(n7510), .A(n7511), .Z(n7509) );
XOR U12517 ( .A(c2503), .B(b[2503]), .Z(n7510) );
XNOR U12518 ( .A(b[2503]), .B(n7511), .Z(c[2503]) );
XNOR U12519 ( .A(a[2503]), .B(c2503), .Z(n7511) );
XOR U12520 ( .A(c2504), .B(n7512), .Z(c2505) );
ANDN U12521 ( .B(n7513), .A(n7514), .Z(n7512) );
XOR U12522 ( .A(c2504), .B(b[2504]), .Z(n7513) );
XNOR U12523 ( .A(b[2504]), .B(n7514), .Z(c[2504]) );
XNOR U12524 ( .A(a[2504]), .B(c2504), .Z(n7514) );
XOR U12525 ( .A(c2505), .B(n7515), .Z(c2506) );
ANDN U12526 ( .B(n7516), .A(n7517), .Z(n7515) );
XOR U12527 ( .A(c2505), .B(b[2505]), .Z(n7516) );
XNOR U12528 ( .A(b[2505]), .B(n7517), .Z(c[2505]) );
XNOR U12529 ( .A(a[2505]), .B(c2505), .Z(n7517) );
XOR U12530 ( .A(c2506), .B(n7518), .Z(c2507) );
ANDN U12531 ( .B(n7519), .A(n7520), .Z(n7518) );
XOR U12532 ( .A(c2506), .B(b[2506]), .Z(n7519) );
XNOR U12533 ( .A(b[2506]), .B(n7520), .Z(c[2506]) );
XNOR U12534 ( .A(a[2506]), .B(c2506), .Z(n7520) );
XOR U12535 ( .A(c2507), .B(n7521), .Z(c2508) );
ANDN U12536 ( .B(n7522), .A(n7523), .Z(n7521) );
XOR U12537 ( .A(c2507), .B(b[2507]), .Z(n7522) );
XNOR U12538 ( .A(b[2507]), .B(n7523), .Z(c[2507]) );
XNOR U12539 ( .A(a[2507]), .B(c2507), .Z(n7523) );
XOR U12540 ( .A(c2508), .B(n7524), .Z(c2509) );
ANDN U12541 ( .B(n7525), .A(n7526), .Z(n7524) );
XOR U12542 ( .A(c2508), .B(b[2508]), .Z(n7525) );
XNOR U12543 ( .A(b[2508]), .B(n7526), .Z(c[2508]) );
XNOR U12544 ( .A(a[2508]), .B(c2508), .Z(n7526) );
XOR U12545 ( .A(c2509), .B(n7527), .Z(c2510) );
ANDN U12546 ( .B(n7528), .A(n7529), .Z(n7527) );
XOR U12547 ( .A(c2509), .B(b[2509]), .Z(n7528) );
XNOR U12548 ( .A(b[2509]), .B(n7529), .Z(c[2509]) );
XNOR U12549 ( .A(a[2509]), .B(c2509), .Z(n7529) );
XOR U12550 ( .A(c2510), .B(n7530), .Z(c2511) );
ANDN U12551 ( .B(n7531), .A(n7532), .Z(n7530) );
XOR U12552 ( .A(c2510), .B(b[2510]), .Z(n7531) );
XNOR U12553 ( .A(b[2510]), .B(n7532), .Z(c[2510]) );
XNOR U12554 ( .A(a[2510]), .B(c2510), .Z(n7532) );
XOR U12555 ( .A(c2511), .B(n7533), .Z(c2512) );
ANDN U12556 ( .B(n7534), .A(n7535), .Z(n7533) );
XOR U12557 ( .A(c2511), .B(b[2511]), .Z(n7534) );
XNOR U12558 ( .A(b[2511]), .B(n7535), .Z(c[2511]) );
XNOR U12559 ( .A(a[2511]), .B(c2511), .Z(n7535) );
XOR U12560 ( .A(c2512), .B(n7536), .Z(c2513) );
ANDN U12561 ( .B(n7537), .A(n7538), .Z(n7536) );
XOR U12562 ( .A(c2512), .B(b[2512]), .Z(n7537) );
XNOR U12563 ( .A(b[2512]), .B(n7538), .Z(c[2512]) );
XNOR U12564 ( .A(a[2512]), .B(c2512), .Z(n7538) );
XOR U12565 ( .A(c2513), .B(n7539), .Z(c2514) );
ANDN U12566 ( .B(n7540), .A(n7541), .Z(n7539) );
XOR U12567 ( .A(c2513), .B(b[2513]), .Z(n7540) );
XNOR U12568 ( .A(b[2513]), .B(n7541), .Z(c[2513]) );
XNOR U12569 ( .A(a[2513]), .B(c2513), .Z(n7541) );
XOR U12570 ( .A(c2514), .B(n7542), .Z(c2515) );
ANDN U12571 ( .B(n7543), .A(n7544), .Z(n7542) );
XOR U12572 ( .A(c2514), .B(b[2514]), .Z(n7543) );
XNOR U12573 ( .A(b[2514]), .B(n7544), .Z(c[2514]) );
XNOR U12574 ( .A(a[2514]), .B(c2514), .Z(n7544) );
XOR U12575 ( .A(c2515), .B(n7545), .Z(c2516) );
ANDN U12576 ( .B(n7546), .A(n7547), .Z(n7545) );
XOR U12577 ( .A(c2515), .B(b[2515]), .Z(n7546) );
XNOR U12578 ( .A(b[2515]), .B(n7547), .Z(c[2515]) );
XNOR U12579 ( .A(a[2515]), .B(c2515), .Z(n7547) );
XOR U12580 ( .A(c2516), .B(n7548), .Z(c2517) );
ANDN U12581 ( .B(n7549), .A(n7550), .Z(n7548) );
XOR U12582 ( .A(c2516), .B(b[2516]), .Z(n7549) );
XNOR U12583 ( .A(b[2516]), .B(n7550), .Z(c[2516]) );
XNOR U12584 ( .A(a[2516]), .B(c2516), .Z(n7550) );
XOR U12585 ( .A(c2517), .B(n7551), .Z(c2518) );
ANDN U12586 ( .B(n7552), .A(n7553), .Z(n7551) );
XOR U12587 ( .A(c2517), .B(b[2517]), .Z(n7552) );
XNOR U12588 ( .A(b[2517]), .B(n7553), .Z(c[2517]) );
XNOR U12589 ( .A(a[2517]), .B(c2517), .Z(n7553) );
XOR U12590 ( .A(c2518), .B(n7554), .Z(c2519) );
ANDN U12591 ( .B(n7555), .A(n7556), .Z(n7554) );
XOR U12592 ( .A(c2518), .B(b[2518]), .Z(n7555) );
XNOR U12593 ( .A(b[2518]), .B(n7556), .Z(c[2518]) );
XNOR U12594 ( .A(a[2518]), .B(c2518), .Z(n7556) );
XOR U12595 ( .A(c2519), .B(n7557), .Z(c2520) );
ANDN U12596 ( .B(n7558), .A(n7559), .Z(n7557) );
XOR U12597 ( .A(c2519), .B(b[2519]), .Z(n7558) );
XNOR U12598 ( .A(b[2519]), .B(n7559), .Z(c[2519]) );
XNOR U12599 ( .A(a[2519]), .B(c2519), .Z(n7559) );
XOR U12600 ( .A(c2520), .B(n7560), .Z(c2521) );
ANDN U12601 ( .B(n7561), .A(n7562), .Z(n7560) );
XOR U12602 ( .A(c2520), .B(b[2520]), .Z(n7561) );
XNOR U12603 ( .A(b[2520]), .B(n7562), .Z(c[2520]) );
XNOR U12604 ( .A(a[2520]), .B(c2520), .Z(n7562) );
XOR U12605 ( .A(c2521), .B(n7563), .Z(c2522) );
ANDN U12606 ( .B(n7564), .A(n7565), .Z(n7563) );
XOR U12607 ( .A(c2521), .B(b[2521]), .Z(n7564) );
XNOR U12608 ( .A(b[2521]), .B(n7565), .Z(c[2521]) );
XNOR U12609 ( .A(a[2521]), .B(c2521), .Z(n7565) );
XOR U12610 ( .A(c2522), .B(n7566), .Z(c2523) );
ANDN U12611 ( .B(n7567), .A(n7568), .Z(n7566) );
XOR U12612 ( .A(c2522), .B(b[2522]), .Z(n7567) );
XNOR U12613 ( .A(b[2522]), .B(n7568), .Z(c[2522]) );
XNOR U12614 ( .A(a[2522]), .B(c2522), .Z(n7568) );
XOR U12615 ( .A(c2523), .B(n7569), .Z(c2524) );
ANDN U12616 ( .B(n7570), .A(n7571), .Z(n7569) );
XOR U12617 ( .A(c2523), .B(b[2523]), .Z(n7570) );
XNOR U12618 ( .A(b[2523]), .B(n7571), .Z(c[2523]) );
XNOR U12619 ( .A(a[2523]), .B(c2523), .Z(n7571) );
XOR U12620 ( .A(c2524), .B(n7572), .Z(c2525) );
ANDN U12621 ( .B(n7573), .A(n7574), .Z(n7572) );
XOR U12622 ( .A(c2524), .B(b[2524]), .Z(n7573) );
XNOR U12623 ( .A(b[2524]), .B(n7574), .Z(c[2524]) );
XNOR U12624 ( .A(a[2524]), .B(c2524), .Z(n7574) );
XOR U12625 ( .A(c2525), .B(n7575), .Z(c2526) );
ANDN U12626 ( .B(n7576), .A(n7577), .Z(n7575) );
XOR U12627 ( .A(c2525), .B(b[2525]), .Z(n7576) );
XNOR U12628 ( .A(b[2525]), .B(n7577), .Z(c[2525]) );
XNOR U12629 ( .A(a[2525]), .B(c2525), .Z(n7577) );
XOR U12630 ( .A(c2526), .B(n7578), .Z(c2527) );
ANDN U12631 ( .B(n7579), .A(n7580), .Z(n7578) );
XOR U12632 ( .A(c2526), .B(b[2526]), .Z(n7579) );
XNOR U12633 ( .A(b[2526]), .B(n7580), .Z(c[2526]) );
XNOR U12634 ( .A(a[2526]), .B(c2526), .Z(n7580) );
XOR U12635 ( .A(c2527), .B(n7581), .Z(c2528) );
ANDN U12636 ( .B(n7582), .A(n7583), .Z(n7581) );
XOR U12637 ( .A(c2527), .B(b[2527]), .Z(n7582) );
XNOR U12638 ( .A(b[2527]), .B(n7583), .Z(c[2527]) );
XNOR U12639 ( .A(a[2527]), .B(c2527), .Z(n7583) );
XOR U12640 ( .A(c2528), .B(n7584), .Z(c2529) );
ANDN U12641 ( .B(n7585), .A(n7586), .Z(n7584) );
XOR U12642 ( .A(c2528), .B(b[2528]), .Z(n7585) );
XNOR U12643 ( .A(b[2528]), .B(n7586), .Z(c[2528]) );
XNOR U12644 ( .A(a[2528]), .B(c2528), .Z(n7586) );
XOR U12645 ( .A(c2529), .B(n7587), .Z(c2530) );
ANDN U12646 ( .B(n7588), .A(n7589), .Z(n7587) );
XOR U12647 ( .A(c2529), .B(b[2529]), .Z(n7588) );
XNOR U12648 ( .A(b[2529]), .B(n7589), .Z(c[2529]) );
XNOR U12649 ( .A(a[2529]), .B(c2529), .Z(n7589) );
XOR U12650 ( .A(c2530), .B(n7590), .Z(c2531) );
ANDN U12651 ( .B(n7591), .A(n7592), .Z(n7590) );
XOR U12652 ( .A(c2530), .B(b[2530]), .Z(n7591) );
XNOR U12653 ( .A(b[2530]), .B(n7592), .Z(c[2530]) );
XNOR U12654 ( .A(a[2530]), .B(c2530), .Z(n7592) );
XOR U12655 ( .A(c2531), .B(n7593), .Z(c2532) );
ANDN U12656 ( .B(n7594), .A(n7595), .Z(n7593) );
XOR U12657 ( .A(c2531), .B(b[2531]), .Z(n7594) );
XNOR U12658 ( .A(b[2531]), .B(n7595), .Z(c[2531]) );
XNOR U12659 ( .A(a[2531]), .B(c2531), .Z(n7595) );
XOR U12660 ( .A(c2532), .B(n7596), .Z(c2533) );
ANDN U12661 ( .B(n7597), .A(n7598), .Z(n7596) );
XOR U12662 ( .A(c2532), .B(b[2532]), .Z(n7597) );
XNOR U12663 ( .A(b[2532]), .B(n7598), .Z(c[2532]) );
XNOR U12664 ( .A(a[2532]), .B(c2532), .Z(n7598) );
XOR U12665 ( .A(c2533), .B(n7599), .Z(c2534) );
ANDN U12666 ( .B(n7600), .A(n7601), .Z(n7599) );
XOR U12667 ( .A(c2533), .B(b[2533]), .Z(n7600) );
XNOR U12668 ( .A(b[2533]), .B(n7601), .Z(c[2533]) );
XNOR U12669 ( .A(a[2533]), .B(c2533), .Z(n7601) );
XOR U12670 ( .A(c2534), .B(n7602), .Z(c2535) );
ANDN U12671 ( .B(n7603), .A(n7604), .Z(n7602) );
XOR U12672 ( .A(c2534), .B(b[2534]), .Z(n7603) );
XNOR U12673 ( .A(b[2534]), .B(n7604), .Z(c[2534]) );
XNOR U12674 ( .A(a[2534]), .B(c2534), .Z(n7604) );
XOR U12675 ( .A(c2535), .B(n7605), .Z(c2536) );
ANDN U12676 ( .B(n7606), .A(n7607), .Z(n7605) );
XOR U12677 ( .A(c2535), .B(b[2535]), .Z(n7606) );
XNOR U12678 ( .A(b[2535]), .B(n7607), .Z(c[2535]) );
XNOR U12679 ( .A(a[2535]), .B(c2535), .Z(n7607) );
XOR U12680 ( .A(c2536), .B(n7608), .Z(c2537) );
ANDN U12681 ( .B(n7609), .A(n7610), .Z(n7608) );
XOR U12682 ( .A(c2536), .B(b[2536]), .Z(n7609) );
XNOR U12683 ( .A(b[2536]), .B(n7610), .Z(c[2536]) );
XNOR U12684 ( .A(a[2536]), .B(c2536), .Z(n7610) );
XOR U12685 ( .A(c2537), .B(n7611), .Z(c2538) );
ANDN U12686 ( .B(n7612), .A(n7613), .Z(n7611) );
XOR U12687 ( .A(c2537), .B(b[2537]), .Z(n7612) );
XNOR U12688 ( .A(b[2537]), .B(n7613), .Z(c[2537]) );
XNOR U12689 ( .A(a[2537]), .B(c2537), .Z(n7613) );
XOR U12690 ( .A(c2538), .B(n7614), .Z(c2539) );
ANDN U12691 ( .B(n7615), .A(n7616), .Z(n7614) );
XOR U12692 ( .A(c2538), .B(b[2538]), .Z(n7615) );
XNOR U12693 ( .A(b[2538]), .B(n7616), .Z(c[2538]) );
XNOR U12694 ( .A(a[2538]), .B(c2538), .Z(n7616) );
XOR U12695 ( .A(c2539), .B(n7617), .Z(c2540) );
ANDN U12696 ( .B(n7618), .A(n7619), .Z(n7617) );
XOR U12697 ( .A(c2539), .B(b[2539]), .Z(n7618) );
XNOR U12698 ( .A(b[2539]), .B(n7619), .Z(c[2539]) );
XNOR U12699 ( .A(a[2539]), .B(c2539), .Z(n7619) );
XOR U12700 ( .A(c2540), .B(n7620), .Z(c2541) );
ANDN U12701 ( .B(n7621), .A(n7622), .Z(n7620) );
XOR U12702 ( .A(c2540), .B(b[2540]), .Z(n7621) );
XNOR U12703 ( .A(b[2540]), .B(n7622), .Z(c[2540]) );
XNOR U12704 ( .A(a[2540]), .B(c2540), .Z(n7622) );
XOR U12705 ( .A(c2541), .B(n7623), .Z(c2542) );
ANDN U12706 ( .B(n7624), .A(n7625), .Z(n7623) );
XOR U12707 ( .A(c2541), .B(b[2541]), .Z(n7624) );
XNOR U12708 ( .A(b[2541]), .B(n7625), .Z(c[2541]) );
XNOR U12709 ( .A(a[2541]), .B(c2541), .Z(n7625) );
XOR U12710 ( .A(c2542), .B(n7626), .Z(c2543) );
ANDN U12711 ( .B(n7627), .A(n7628), .Z(n7626) );
XOR U12712 ( .A(c2542), .B(b[2542]), .Z(n7627) );
XNOR U12713 ( .A(b[2542]), .B(n7628), .Z(c[2542]) );
XNOR U12714 ( .A(a[2542]), .B(c2542), .Z(n7628) );
XOR U12715 ( .A(c2543), .B(n7629), .Z(c2544) );
ANDN U12716 ( .B(n7630), .A(n7631), .Z(n7629) );
XOR U12717 ( .A(c2543), .B(b[2543]), .Z(n7630) );
XNOR U12718 ( .A(b[2543]), .B(n7631), .Z(c[2543]) );
XNOR U12719 ( .A(a[2543]), .B(c2543), .Z(n7631) );
XOR U12720 ( .A(c2544), .B(n7632), .Z(c2545) );
ANDN U12721 ( .B(n7633), .A(n7634), .Z(n7632) );
XOR U12722 ( .A(c2544), .B(b[2544]), .Z(n7633) );
XNOR U12723 ( .A(b[2544]), .B(n7634), .Z(c[2544]) );
XNOR U12724 ( .A(a[2544]), .B(c2544), .Z(n7634) );
XOR U12725 ( .A(c2545), .B(n7635), .Z(c2546) );
ANDN U12726 ( .B(n7636), .A(n7637), .Z(n7635) );
XOR U12727 ( .A(c2545), .B(b[2545]), .Z(n7636) );
XNOR U12728 ( .A(b[2545]), .B(n7637), .Z(c[2545]) );
XNOR U12729 ( .A(a[2545]), .B(c2545), .Z(n7637) );
XOR U12730 ( .A(c2546), .B(n7638), .Z(c2547) );
ANDN U12731 ( .B(n7639), .A(n7640), .Z(n7638) );
XOR U12732 ( .A(c2546), .B(b[2546]), .Z(n7639) );
XNOR U12733 ( .A(b[2546]), .B(n7640), .Z(c[2546]) );
XNOR U12734 ( .A(a[2546]), .B(c2546), .Z(n7640) );
XOR U12735 ( .A(c2547), .B(n7641), .Z(c2548) );
ANDN U12736 ( .B(n7642), .A(n7643), .Z(n7641) );
XOR U12737 ( .A(c2547), .B(b[2547]), .Z(n7642) );
XNOR U12738 ( .A(b[2547]), .B(n7643), .Z(c[2547]) );
XNOR U12739 ( .A(a[2547]), .B(c2547), .Z(n7643) );
XOR U12740 ( .A(c2548), .B(n7644), .Z(c2549) );
ANDN U12741 ( .B(n7645), .A(n7646), .Z(n7644) );
XOR U12742 ( .A(c2548), .B(b[2548]), .Z(n7645) );
XNOR U12743 ( .A(b[2548]), .B(n7646), .Z(c[2548]) );
XNOR U12744 ( .A(a[2548]), .B(c2548), .Z(n7646) );
XOR U12745 ( .A(c2549), .B(n7647), .Z(c2550) );
ANDN U12746 ( .B(n7648), .A(n7649), .Z(n7647) );
XOR U12747 ( .A(c2549), .B(b[2549]), .Z(n7648) );
XNOR U12748 ( .A(b[2549]), .B(n7649), .Z(c[2549]) );
XNOR U12749 ( .A(a[2549]), .B(c2549), .Z(n7649) );
XOR U12750 ( .A(c2550), .B(n7650), .Z(c2551) );
ANDN U12751 ( .B(n7651), .A(n7652), .Z(n7650) );
XOR U12752 ( .A(c2550), .B(b[2550]), .Z(n7651) );
XNOR U12753 ( .A(b[2550]), .B(n7652), .Z(c[2550]) );
XNOR U12754 ( .A(a[2550]), .B(c2550), .Z(n7652) );
XOR U12755 ( .A(c2551), .B(n7653), .Z(c2552) );
ANDN U12756 ( .B(n7654), .A(n7655), .Z(n7653) );
XOR U12757 ( .A(c2551), .B(b[2551]), .Z(n7654) );
XNOR U12758 ( .A(b[2551]), .B(n7655), .Z(c[2551]) );
XNOR U12759 ( .A(a[2551]), .B(c2551), .Z(n7655) );
XOR U12760 ( .A(c2552), .B(n7656), .Z(c2553) );
ANDN U12761 ( .B(n7657), .A(n7658), .Z(n7656) );
XOR U12762 ( .A(c2552), .B(b[2552]), .Z(n7657) );
XNOR U12763 ( .A(b[2552]), .B(n7658), .Z(c[2552]) );
XNOR U12764 ( .A(a[2552]), .B(c2552), .Z(n7658) );
XOR U12765 ( .A(c2553), .B(n7659), .Z(c2554) );
ANDN U12766 ( .B(n7660), .A(n7661), .Z(n7659) );
XOR U12767 ( .A(c2553), .B(b[2553]), .Z(n7660) );
XNOR U12768 ( .A(b[2553]), .B(n7661), .Z(c[2553]) );
XNOR U12769 ( .A(a[2553]), .B(c2553), .Z(n7661) );
XOR U12770 ( .A(c2554), .B(n7662), .Z(c2555) );
ANDN U12771 ( .B(n7663), .A(n7664), .Z(n7662) );
XOR U12772 ( .A(c2554), .B(b[2554]), .Z(n7663) );
XNOR U12773 ( .A(b[2554]), .B(n7664), .Z(c[2554]) );
XNOR U12774 ( .A(a[2554]), .B(c2554), .Z(n7664) );
XOR U12775 ( .A(c2555), .B(n7665), .Z(c2556) );
ANDN U12776 ( .B(n7666), .A(n7667), .Z(n7665) );
XOR U12777 ( .A(c2555), .B(b[2555]), .Z(n7666) );
XNOR U12778 ( .A(b[2555]), .B(n7667), .Z(c[2555]) );
XNOR U12779 ( .A(a[2555]), .B(c2555), .Z(n7667) );
XOR U12780 ( .A(c2556), .B(n7668), .Z(c2557) );
ANDN U12781 ( .B(n7669), .A(n7670), .Z(n7668) );
XOR U12782 ( .A(c2556), .B(b[2556]), .Z(n7669) );
XNOR U12783 ( .A(b[2556]), .B(n7670), .Z(c[2556]) );
XNOR U12784 ( .A(a[2556]), .B(c2556), .Z(n7670) );
XOR U12785 ( .A(c2557), .B(n7671), .Z(c2558) );
ANDN U12786 ( .B(n7672), .A(n7673), .Z(n7671) );
XOR U12787 ( .A(c2557), .B(b[2557]), .Z(n7672) );
XNOR U12788 ( .A(b[2557]), .B(n7673), .Z(c[2557]) );
XNOR U12789 ( .A(a[2557]), .B(c2557), .Z(n7673) );
XOR U12790 ( .A(c2558), .B(n7674), .Z(c2559) );
ANDN U12791 ( .B(n7675), .A(n7676), .Z(n7674) );
XOR U12792 ( .A(c2558), .B(b[2558]), .Z(n7675) );
XNOR U12793 ( .A(b[2558]), .B(n7676), .Z(c[2558]) );
XNOR U12794 ( .A(a[2558]), .B(c2558), .Z(n7676) );
XOR U12795 ( .A(c2559), .B(n7677), .Z(c2560) );
ANDN U12796 ( .B(n7678), .A(n7679), .Z(n7677) );
XOR U12797 ( .A(c2559), .B(b[2559]), .Z(n7678) );
XNOR U12798 ( .A(b[2559]), .B(n7679), .Z(c[2559]) );
XNOR U12799 ( .A(a[2559]), .B(c2559), .Z(n7679) );
XOR U12800 ( .A(c2560), .B(n7680), .Z(c2561) );
ANDN U12801 ( .B(n7681), .A(n7682), .Z(n7680) );
XOR U12802 ( .A(c2560), .B(b[2560]), .Z(n7681) );
XNOR U12803 ( .A(b[2560]), .B(n7682), .Z(c[2560]) );
XNOR U12804 ( .A(a[2560]), .B(c2560), .Z(n7682) );
XOR U12805 ( .A(c2561), .B(n7683), .Z(c2562) );
ANDN U12806 ( .B(n7684), .A(n7685), .Z(n7683) );
XOR U12807 ( .A(c2561), .B(b[2561]), .Z(n7684) );
XNOR U12808 ( .A(b[2561]), .B(n7685), .Z(c[2561]) );
XNOR U12809 ( .A(a[2561]), .B(c2561), .Z(n7685) );
XOR U12810 ( .A(c2562), .B(n7686), .Z(c2563) );
ANDN U12811 ( .B(n7687), .A(n7688), .Z(n7686) );
XOR U12812 ( .A(c2562), .B(b[2562]), .Z(n7687) );
XNOR U12813 ( .A(b[2562]), .B(n7688), .Z(c[2562]) );
XNOR U12814 ( .A(a[2562]), .B(c2562), .Z(n7688) );
XOR U12815 ( .A(c2563), .B(n7689), .Z(c2564) );
ANDN U12816 ( .B(n7690), .A(n7691), .Z(n7689) );
XOR U12817 ( .A(c2563), .B(b[2563]), .Z(n7690) );
XNOR U12818 ( .A(b[2563]), .B(n7691), .Z(c[2563]) );
XNOR U12819 ( .A(a[2563]), .B(c2563), .Z(n7691) );
XOR U12820 ( .A(c2564), .B(n7692), .Z(c2565) );
ANDN U12821 ( .B(n7693), .A(n7694), .Z(n7692) );
XOR U12822 ( .A(c2564), .B(b[2564]), .Z(n7693) );
XNOR U12823 ( .A(b[2564]), .B(n7694), .Z(c[2564]) );
XNOR U12824 ( .A(a[2564]), .B(c2564), .Z(n7694) );
XOR U12825 ( .A(c2565), .B(n7695), .Z(c2566) );
ANDN U12826 ( .B(n7696), .A(n7697), .Z(n7695) );
XOR U12827 ( .A(c2565), .B(b[2565]), .Z(n7696) );
XNOR U12828 ( .A(b[2565]), .B(n7697), .Z(c[2565]) );
XNOR U12829 ( .A(a[2565]), .B(c2565), .Z(n7697) );
XOR U12830 ( .A(c2566), .B(n7698), .Z(c2567) );
ANDN U12831 ( .B(n7699), .A(n7700), .Z(n7698) );
XOR U12832 ( .A(c2566), .B(b[2566]), .Z(n7699) );
XNOR U12833 ( .A(b[2566]), .B(n7700), .Z(c[2566]) );
XNOR U12834 ( .A(a[2566]), .B(c2566), .Z(n7700) );
XOR U12835 ( .A(c2567), .B(n7701), .Z(c2568) );
ANDN U12836 ( .B(n7702), .A(n7703), .Z(n7701) );
XOR U12837 ( .A(c2567), .B(b[2567]), .Z(n7702) );
XNOR U12838 ( .A(b[2567]), .B(n7703), .Z(c[2567]) );
XNOR U12839 ( .A(a[2567]), .B(c2567), .Z(n7703) );
XOR U12840 ( .A(c2568), .B(n7704), .Z(c2569) );
ANDN U12841 ( .B(n7705), .A(n7706), .Z(n7704) );
XOR U12842 ( .A(c2568), .B(b[2568]), .Z(n7705) );
XNOR U12843 ( .A(b[2568]), .B(n7706), .Z(c[2568]) );
XNOR U12844 ( .A(a[2568]), .B(c2568), .Z(n7706) );
XOR U12845 ( .A(c2569), .B(n7707), .Z(c2570) );
ANDN U12846 ( .B(n7708), .A(n7709), .Z(n7707) );
XOR U12847 ( .A(c2569), .B(b[2569]), .Z(n7708) );
XNOR U12848 ( .A(b[2569]), .B(n7709), .Z(c[2569]) );
XNOR U12849 ( .A(a[2569]), .B(c2569), .Z(n7709) );
XOR U12850 ( .A(c2570), .B(n7710), .Z(c2571) );
ANDN U12851 ( .B(n7711), .A(n7712), .Z(n7710) );
XOR U12852 ( .A(c2570), .B(b[2570]), .Z(n7711) );
XNOR U12853 ( .A(b[2570]), .B(n7712), .Z(c[2570]) );
XNOR U12854 ( .A(a[2570]), .B(c2570), .Z(n7712) );
XOR U12855 ( .A(c2571), .B(n7713), .Z(c2572) );
ANDN U12856 ( .B(n7714), .A(n7715), .Z(n7713) );
XOR U12857 ( .A(c2571), .B(b[2571]), .Z(n7714) );
XNOR U12858 ( .A(b[2571]), .B(n7715), .Z(c[2571]) );
XNOR U12859 ( .A(a[2571]), .B(c2571), .Z(n7715) );
XOR U12860 ( .A(c2572), .B(n7716), .Z(c2573) );
ANDN U12861 ( .B(n7717), .A(n7718), .Z(n7716) );
XOR U12862 ( .A(c2572), .B(b[2572]), .Z(n7717) );
XNOR U12863 ( .A(b[2572]), .B(n7718), .Z(c[2572]) );
XNOR U12864 ( .A(a[2572]), .B(c2572), .Z(n7718) );
XOR U12865 ( .A(c2573), .B(n7719), .Z(c2574) );
ANDN U12866 ( .B(n7720), .A(n7721), .Z(n7719) );
XOR U12867 ( .A(c2573), .B(b[2573]), .Z(n7720) );
XNOR U12868 ( .A(b[2573]), .B(n7721), .Z(c[2573]) );
XNOR U12869 ( .A(a[2573]), .B(c2573), .Z(n7721) );
XOR U12870 ( .A(c2574), .B(n7722), .Z(c2575) );
ANDN U12871 ( .B(n7723), .A(n7724), .Z(n7722) );
XOR U12872 ( .A(c2574), .B(b[2574]), .Z(n7723) );
XNOR U12873 ( .A(b[2574]), .B(n7724), .Z(c[2574]) );
XNOR U12874 ( .A(a[2574]), .B(c2574), .Z(n7724) );
XOR U12875 ( .A(c2575), .B(n7725), .Z(c2576) );
ANDN U12876 ( .B(n7726), .A(n7727), .Z(n7725) );
XOR U12877 ( .A(c2575), .B(b[2575]), .Z(n7726) );
XNOR U12878 ( .A(b[2575]), .B(n7727), .Z(c[2575]) );
XNOR U12879 ( .A(a[2575]), .B(c2575), .Z(n7727) );
XOR U12880 ( .A(c2576), .B(n7728), .Z(c2577) );
ANDN U12881 ( .B(n7729), .A(n7730), .Z(n7728) );
XOR U12882 ( .A(c2576), .B(b[2576]), .Z(n7729) );
XNOR U12883 ( .A(b[2576]), .B(n7730), .Z(c[2576]) );
XNOR U12884 ( .A(a[2576]), .B(c2576), .Z(n7730) );
XOR U12885 ( .A(c2577), .B(n7731), .Z(c2578) );
ANDN U12886 ( .B(n7732), .A(n7733), .Z(n7731) );
XOR U12887 ( .A(c2577), .B(b[2577]), .Z(n7732) );
XNOR U12888 ( .A(b[2577]), .B(n7733), .Z(c[2577]) );
XNOR U12889 ( .A(a[2577]), .B(c2577), .Z(n7733) );
XOR U12890 ( .A(c2578), .B(n7734), .Z(c2579) );
ANDN U12891 ( .B(n7735), .A(n7736), .Z(n7734) );
XOR U12892 ( .A(c2578), .B(b[2578]), .Z(n7735) );
XNOR U12893 ( .A(b[2578]), .B(n7736), .Z(c[2578]) );
XNOR U12894 ( .A(a[2578]), .B(c2578), .Z(n7736) );
XOR U12895 ( .A(c2579), .B(n7737), .Z(c2580) );
ANDN U12896 ( .B(n7738), .A(n7739), .Z(n7737) );
XOR U12897 ( .A(c2579), .B(b[2579]), .Z(n7738) );
XNOR U12898 ( .A(b[2579]), .B(n7739), .Z(c[2579]) );
XNOR U12899 ( .A(a[2579]), .B(c2579), .Z(n7739) );
XOR U12900 ( .A(c2580), .B(n7740), .Z(c2581) );
ANDN U12901 ( .B(n7741), .A(n7742), .Z(n7740) );
XOR U12902 ( .A(c2580), .B(b[2580]), .Z(n7741) );
XNOR U12903 ( .A(b[2580]), .B(n7742), .Z(c[2580]) );
XNOR U12904 ( .A(a[2580]), .B(c2580), .Z(n7742) );
XOR U12905 ( .A(c2581), .B(n7743), .Z(c2582) );
ANDN U12906 ( .B(n7744), .A(n7745), .Z(n7743) );
XOR U12907 ( .A(c2581), .B(b[2581]), .Z(n7744) );
XNOR U12908 ( .A(b[2581]), .B(n7745), .Z(c[2581]) );
XNOR U12909 ( .A(a[2581]), .B(c2581), .Z(n7745) );
XOR U12910 ( .A(c2582), .B(n7746), .Z(c2583) );
ANDN U12911 ( .B(n7747), .A(n7748), .Z(n7746) );
XOR U12912 ( .A(c2582), .B(b[2582]), .Z(n7747) );
XNOR U12913 ( .A(b[2582]), .B(n7748), .Z(c[2582]) );
XNOR U12914 ( .A(a[2582]), .B(c2582), .Z(n7748) );
XOR U12915 ( .A(c2583), .B(n7749), .Z(c2584) );
ANDN U12916 ( .B(n7750), .A(n7751), .Z(n7749) );
XOR U12917 ( .A(c2583), .B(b[2583]), .Z(n7750) );
XNOR U12918 ( .A(b[2583]), .B(n7751), .Z(c[2583]) );
XNOR U12919 ( .A(a[2583]), .B(c2583), .Z(n7751) );
XOR U12920 ( .A(c2584), .B(n7752), .Z(c2585) );
ANDN U12921 ( .B(n7753), .A(n7754), .Z(n7752) );
XOR U12922 ( .A(c2584), .B(b[2584]), .Z(n7753) );
XNOR U12923 ( .A(b[2584]), .B(n7754), .Z(c[2584]) );
XNOR U12924 ( .A(a[2584]), .B(c2584), .Z(n7754) );
XOR U12925 ( .A(c2585), .B(n7755), .Z(c2586) );
ANDN U12926 ( .B(n7756), .A(n7757), .Z(n7755) );
XOR U12927 ( .A(c2585), .B(b[2585]), .Z(n7756) );
XNOR U12928 ( .A(b[2585]), .B(n7757), .Z(c[2585]) );
XNOR U12929 ( .A(a[2585]), .B(c2585), .Z(n7757) );
XOR U12930 ( .A(c2586), .B(n7758), .Z(c2587) );
ANDN U12931 ( .B(n7759), .A(n7760), .Z(n7758) );
XOR U12932 ( .A(c2586), .B(b[2586]), .Z(n7759) );
XNOR U12933 ( .A(b[2586]), .B(n7760), .Z(c[2586]) );
XNOR U12934 ( .A(a[2586]), .B(c2586), .Z(n7760) );
XOR U12935 ( .A(c2587), .B(n7761), .Z(c2588) );
ANDN U12936 ( .B(n7762), .A(n7763), .Z(n7761) );
XOR U12937 ( .A(c2587), .B(b[2587]), .Z(n7762) );
XNOR U12938 ( .A(b[2587]), .B(n7763), .Z(c[2587]) );
XNOR U12939 ( .A(a[2587]), .B(c2587), .Z(n7763) );
XOR U12940 ( .A(c2588), .B(n7764), .Z(c2589) );
ANDN U12941 ( .B(n7765), .A(n7766), .Z(n7764) );
XOR U12942 ( .A(c2588), .B(b[2588]), .Z(n7765) );
XNOR U12943 ( .A(b[2588]), .B(n7766), .Z(c[2588]) );
XNOR U12944 ( .A(a[2588]), .B(c2588), .Z(n7766) );
XOR U12945 ( .A(c2589), .B(n7767), .Z(c2590) );
ANDN U12946 ( .B(n7768), .A(n7769), .Z(n7767) );
XOR U12947 ( .A(c2589), .B(b[2589]), .Z(n7768) );
XNOR U12948 ( .A(b[2589]), .B(n7769), .Z(c[2589]) );
XNOR U12949 ( .A(a[2589]), .B(c2589), .Z(n7769) );
XOR U12950 ( .A(c2590), .B(n7770), .Z(c2591) );
ANDN U12951 ( .B(n7771), .A(n7772), .Z(n7770) );
XOR U12952 ( .A(c2590), .B(b[2590]), .Z(n7771) );
XNOR U12953 ( .A(b[2590]), .B(n7772), .Z(c[2590]) );
XNOR U12954 ( .A(a[2590]), .B(c2590), .Z(n7772) );
XOR U12955 ( .A(c2591), .B(n7773), .Z(c2592) );
ANDN U12956 ( .B(n7774), .A(n7775), .Z(n7773) );
XOR U12957 ( .A(c2591), .B(b[2591]), .Z(n7774) );
XNOR U12958 ( .A(b[2591]), .B(n7775), .Z(c[2591]) );
XNOR U12959 ( .A(a[2591]), .B(c2591), .Z(n7775) );
XOR U12960 ( .A(c2592), .B(n7776), .Z(c2593) );
ANDN U12961 ( .B(n7777), .A(n7778), .Z(n7776) );
XOR U12962 ( .A(c2592), .B(b[2592]), .Z(n7777) );
XNOR U12963 ( .A(b[2592]), .B(n7778), .Z(c[2592]) );
XNOR U12964 ( .A(a[2592]), .B(c2592), .Z(n7778) );
XOR U12965 ( .A(c2593), .B(n7779), .Z(c2594) );
ANDN U12966 ( .B(n7780), .A(n7781), .Z(n7779) );
XOR U12967 ( .A(c2593), .B(b[2593]), .Z(n7780) );
XNOR U12968 ( .A(b[2593]), .B(n7781), .Z(c[2593]) );
XNOR U12969 ( .A(a[2593]), .B(c2593), .Z(n7781) );
XOR U12970 ( .A(c2594), .B(n7782), .Z(c2595) );
ANDN U12971 ( .B(n7783), .A(n7784), .Z(n7782) );
XOR U12972 ( .A(c2594), .B(b[2594]), .Z(n7783) );
XNOR U12973 ( .A(b[2594]), .B(n7784), .Z(c[2594]) );
XNOR U12974 ( .A(a[2594]), .B(c2594), .Z(n7784) );
XOR U12975 ( .A(c2595), .B(n7785), .Z(c2596) );
ANDN U12976 ( .B(n7786), .A(n7787), .Z(n7785) );
XOR U12977 ( .A(c2595), .B(b[2595]), .Z(n7786) );
XNOR U12978 ( .A(b[2595]), .B(n7787), .Z(c[2595]) );
XNOR U12979 ( .A(a[2595]), .B(c2595), .Z(n7787) );
XOR U12980 ( .A(c2596), .B(n7788), .Z(c2597) );
ANDN U12981 ( .B(n7789), .A(n7790), .Z(n7788) );
XOR U12982 ( .A(c2596), .B(b[2596]), .Z(n7789) );
XNOR U12983 ( .A(b[2596]), .B(n7790), .Z(c[2596]) );
XNOR U12984 ( .A(a[2596]), .B(c2596), .Z(n7790) );
XOR U12985 ( .A(c2597), .B(n7791), .Z(c2598) );
ANDN U12986 ( .B(n7792), .A(n7793), .Z(n7791) );
XOR U12987 ( .A(c2597), .B(b[2597]), .Z(n7792) );
XNOR U12988 ( .A(b[2597]), .B(n7793), .Z(c[2597]) );
XNOR U12989 ( .A(a[2597]), .B(c2597), .Z(n7793) );
XOR U12990 ( .A(c2598), .B(n7794), .Z(c2599) );
ANDN U12991 ( .B(n7795), .A(n7796), .Z(n7794) );
XOR U12992 ( .A(c2598), .B(b[2598]), .Z(n7795) );
XNOR U12993 ( .A(b[2598]), .B(n7796), .Z(c[2598]) );
XNOR U12994 ( .A(a[2598]), .B(c2598), .Z(n7796) );
XOR U12995 ( .A(c2599), .B(n7797), .Z(c2600) );
ANDN U12996 ( .B(n7798), .A(n7799), .Z(n7797) );
XOR U12997 ( .A(c2599), .B(b[2599]), .Z(n7798) );
XNOR U12998 ( .A(b[2599]), .B(n7799), .Z(c[2599]) );
XNOR U12999 ( .A(a[2599]), .B(c2599), .Z(n7799) );
XOR U13000 ( .A(c2600), .B(n7800), .Z(c2601) );
ANDN U13001 ( .B(n7801), .A(n7802), .Z(n7800) );
XOR U13002 ( .A(c2600), .B(b[2600]), .Z(n7801) );
XNOR U13003 ( .A(b[2600]), .B(n7802), .Z(c[2600]) );
XNOR U13004 ( .A(a[2600]), .B(c2600), .Z(n7802) );
XOR U13005 ( .A(c2601), .B(n7803), .Z(c2602) );
ANDN U13006 ( .B(n7804), .A(n7805), .Z(n7803) );
XOR U13007 ( .A(c2601), .B(b[2601]), .Z(n7804) );
XNOR U13008 ( .A(b[2601]), .B(n7805), .Z(c[2601]) );
XNOR U13009 ( .A(a[2601]), .B(c2601), .Z(n7805) );
XOR U13010 ( .A(c2602), .B(n7806), .Z(c2603) );
ANDN U13011 ( .B(n7807), .A(n7808), .Z(n7806) );
XOR U13012 ( .A(c2602), .B(b[2602]), .Z(n7807) );
XNOR U13013 ( .A(b[2602]), .B(n7808), .Z(c[2602]) );
XNOR U13014 ( .A(a[2602]), .B(c2602), .Z(n7808) );
XOR U13015 ( .A(c2603), .B(n7809), .Z(c2604) );
ANDN U13016 ( .B(n7810), .A(n7811), .Z(n7809) );
XOR U13017 ( .A(c2603), .B(b[2603]), .Z(n7810) );
XNOR U13018 ( .A(b[2603]), .B(n7811), .Z(c[2603]) );
XNOR U13019 ( .A(a[2603]), .B(c2603), .Z(n7811) );
XOR U13020 ( .A(c2604), .B(n7812), .Z(c2605) );
ANDN U13021 ( .B(n7813), .A(n7814), .Z(n7812) );
XOR U13022 ( .A(c2604), .B(b[2604]), .Z(n7813) );
XNOR U13023 ( .A(b[2604]), .B(n7814), .Z(c[2604]) );
XNOR U13024 ( .A(a[2604]), .B(c2604), .Z(n7814) );
XOR U13025 ( .A(c2605), .B(n7815), .Z(c2606) );
ANDN U13026 ( .B(n7816), .A(n7817), .Z(n7815) );
XOR U13027 ( .A(c2605), .B(b[2605]), .Z(n7816) );
XNOR U13028 ( .A(b[2605]), .B(n7817), .Z(c[2605]) );
XNOR U13029 ( .A(a[2605]), .B(c2605), .Z(n7817) );
XOR U13030 ( .A(c2606), .B(n7818), .Z(c2607) );
ANDN U13031 ( .B(n7819), .A(n7820), .Z(n7818) );
XOR U13032 ( .A(c2606), .B(b[2606]), .Z(n7819) );
XNOR U13033 ( .A(b[2606]), .B(n7820), .Z(c[2606]) );
XNOR U13034 ( .A(a[2606]), .B(c2606), .Z(n7820) );
XOR U13035 ( .A(c2607), .B(n7821), .Z(c2608) );
ANDN U13036 ( .B(n7822), .A(n7823), .Z(n7821) );
XOR U13037 ( .A(c2607), .B(b[2607]), .Z(n7822) );
XNOR U13038 ( .A(b[2607]), .B(n7823), .Z(c[2607]) );
XNOR U13039 ( .A(a[2607]), .B(c2607), .Z(n7823) );
XOR U13040 ( .A(c2608), .B(n7824), .Z(c2609) );
ANDN U13041 ( .B(n7825), .A(n7826), .Z(n7824) );
XOR U13042 ( .A(c2608), .B(b[2608]), .Z(n7825) );
XNOR U13043 ( .A(b[2608]), .B(n7826), .Z(c[2608]) );
XNOR U13044 ( .A(a[2608]), .B(c2608), .Z(n7826) );
XOR U13045 ( .A(c2609), .B(n7827), .Z(c2610) );
ANDN U13046 ( .B(n7828), .A(n7829), .Z(n7827) );
XOR U13047 ( .A(c2609), .B(b[2609]), .Z(n7828) );
XNOR U13048 ( .A(b[2609]), .B(n7829), .Z(c[2609]) );
XNOR U13049 ( .A(a[2609]), .B(c2609), .Z(n7829) );
XOR U13050 ( .A(c2610), .B(n7830), .Z(c2611) );
ANDN U13051 ( .B(n7831), .A(n7832), .Z(n7830) );
XOR U13052 ( .A(c2610), .B(b[2610]), .Z(n7831) );
XNOR U13053 ( .A(b[2610]), .B(n7832), .Z(c[2610]) );
XNOR U13054 ( .A(a[2610]), .B(c2610), .Z(n7832) );
XOR U13055 ( .A(c2611), .B(n7833), .Z(c2612) );
ANDN U13056 ( .B(n7834), .A(n7835), .Z(n7833) );
XOR U13057 ( .A(c2611), .B(b[2611]), .Z(n7834) );
XNOR U13058 ( .A(b[2611]), .B(n7835), .Z(c[2611]) );
XNOR U13059 ( .A(a[2611]), .B(c2611), .Z(n7835) );
XOR U13060 ( .A(c2612), .B(n7836), .Z(c2613) );
ANDN U13061 ( .B(n7837), .A(n7838), .Z(n7836) );
XOR U13062 ( .A(c2612), .B(b[2612]), .Z(n7837) );
XNOR U13063 ( .A(b[2612]), .B(n7838), .Z(c[2612]) );
XNOR U13064 ( .A(a[2612]), .B(c2612), .Z(n7838) );
XOR U13065 ( .A(c2613), .B(n7839), .Z(c2614) );
ANDN U13066 ( .B(n7840), .A(n7841), .Z(n7839) );
XOR U13067 ( .A(c2613), .B(b[2613]), .Z(n7840) );
XNOR U13068 ( .A(b[2613]), .B(n7841), .Z(c[2613]) );
XNOR U13069 ( .A(a[2613]), .B(c2613), .Z(n7841) );
XOR U13070 ( .A(c2614), .B(n7842), .Z(c2615) );
ANDN U13071 ( .B(n7843), .A(n7844), .Z(n7842) );
XOR U13072 ( .A(c2614), .B(b[2614]), .Z(n7843) );
XNOR U13073 ( .A(b[2614]), .B(n7844), .Z(c[2614]) );
XNOR U13074 ( .A(a[2614]), .B(c2614), .Z(n7844) );
XOR U13075 ( .A(c2615), .B(n7845), .Z(c2616) );
ANDN U13076 ( .B(n7846), .A(n7847), .Z(n7845) );
XOR U13077 ( .A(c2615), .B(b[2615]), .Z(n7846) );
XNOR U13078 ( .A(b[2615]), .B(n7847), .Z(c[2615]) );
XNOR U13079 ( .A(a[2615]), .B(c2615), .Z(n7847) );
XOR U13080 ( .A(c2616), .B(n7848), .Z(c2617) );
ANDN U13081 ( .B(n7849), .A(n7850), .Z(n7848) );
XOR U13082 ( .A(c2616), .B(b[2616]), .Z(n7849) );
XNOR U13083 ( .A(b[2616]), .B(n7850), .Z(c[2616]) );
XNOR U13084 ( .A(a[2616]), .B(c2616), .Z(n7850) );
XOR U13085 ( .A(c2617), .B(n7851), .Z(c2618) );
ANDN U13086 ( .B(n7852), .A(n7853), .Z(n7851) );
XOR U13087 ( .A(c2617), .B(b[2617]), .Z(n7852) );
XNOR U13088 ( .A(b[2617]), .B(n7853), .Z(c[2617]) );
XNOR U13089 ( .A(a[2617]), .B(c2617), .Z(n7853) );
XOR U13090 ( .A(c2618), .B(n7854), .Z(c2619) );
ANDN U13091 ( .B(n7855), .A(n7856), .Z(n7854) );
XOR U13092 ( .A(c2618), .B(b[2618]), .Z(n7855) );
XNOR U13093 ( .A(b[2618]), .B(n7856), .Z(c[2618]) );
XNOR U13094 ( .A(a[2618]), .B(c2618), .Z(n7856) );
XOR U13095 ( .A(c2619), .B(n7857), .Z(c2620) );
ANDN U13096 ( .B(n7858), .A(n7859), .Z(n7857) );
XOR U13097 ( .A(c2619), .B(b[2619]), .Z(n7858) );
XNOR U13098 ( .A(b[2619]), .B(n7859), .Z(c[2619]) );
XNOR U13099 ( .A(a[2619]), .B(c2619), .Z(n7859) );
XOR U13100 ( .A(c2620), .B(n7860), .Z(c2621) );
ANDN U13101 ( .B(n7861), .A(n7862), .Z(n7860) );
XOR U13102 ( .A(c2620), .B(b[2620]), .Z(n7861) );
XNOR U13103 ( .A(b[2620]), .B(n7862), .Z(c[2620]) );
XNOR U13104 ( .A(a[2620]), .B(c2620), .Z(n7862) );
XOR U13105 ( .A(c2621), .B(n7863), .Z(c2622) );
ANDN U13106 ( .B(n7864), .A(n7865), .Z(n7863) );
XOR U13107 ( .A(c2621), .B(b[2621]), .Z(n7864) );
XNOR U13108 ( .A(b[2621]), .B(n7865), .Z(c[2621]) );
XNOR U13109 ( .A(a[2621]), .B(c2621), .Z(n7865) );
XOR U13110 ( .A(c2622), .B(n7866), .Z(c2623) );
ANDN U13111 ( .B(n7867), .A(n7868), .Z(n7866) );
XOR U13112 ( .A(c2622), .B(b[2622]), .Z(n7867) );
XNOR U13113 ( .A(b[2622]), .B(n7868), .Z(c[2622]) );
XNOR U13114 ( .A(a[2622]), .B(c2622), .Z(n7868) );
XOR U13115 ( .A(c2623), .B(n7869), .Z(c2624) );
ANDN U13116 ( .B(n7870), .A(n7871), .Z(n7869) );
XOR U13117 ( .A(c2623), .B(b[2623]), .Z(n7870) );
XNOR U13118 ( .A(b[2623]), .B(n7871), .Z(c[2623]) );
XNOR U13119 ( .A(a[2623]), .B(c2623), .Z(n7871) );
XOR U13120 ( .A(c2624), .B(n7872), .Z(c2625) );
ANDN U13121 ( .B(n7873), .A(n7874), .Z(n7872) );
XOR U13122 ( .A(c2624), .B(b[2624]), .Z(n7873) );
XNOR U13123 ( .A(b[2624]), .B(n7874), .Z(c[2624]) );
XNOR U13124 ( .A(a[2624]), .B(c2624), .Z(n7874) );
XOR U13125 ( .A(c2625), .B(n7875), .Z(c2626) );
ANDN U13126 ( .B(n7876), .A(n7877), .Z(n7875) );
XOR U13127 ( .A(c2625), .B(b[2625]), .Z(n7876) );
XNOR U13128 ( .A(b[2625]), .B(n7877), .Z(c[2625]) );
XNOR U13129 ( .A(a[2625]), .B(c2625), .Z(n7877) );
XOR U13130 ( .A(c2626), .B(n7878), .Z(c2627) );
ANDN U13131 ( .B(n7879), .A(n7880), .Z(n7878) );
XOR U13132 ( .A(c2626), .B(b[2626]), .Z(n7879) );
XNOR U13133 ( .A(b[2626]), .B(n7880), .Z(c[2626]) );
XNOR U13134 ( .A(a[2626]), .B(c2626), .Z(n7880) );
XOR U13135 ( .A(c2627), .B(n7881), .Z(c2628) );
ANDN U13136 ( .B(n7882), .A(n7883), .Z(n7881) );
XOR U13137 ( .A(c2627), .B(b[2627]), .Z(n7882) );
XNOR U13138 ( .A(b[2627]), .B(n7883), .Z(c[2627]) );
XNOR U13139 ( .A(a[2627]), .B(c2627), .Z(n7883) );
XOR U13140 ( .A(c2628), .B(n7884), .Z(c2629) );
ANDN U13141 ( .B(n7885), .A(n7886), .Z(n7884) );
XOR U13142 ( .A(c2628), .B(b[2628]), .Z(n7885) );
XNOR U13143 ( .A(b[2628]), .B(n7886), .Z(c[2628]) );
XNOR U13144 ( .A(a[2628]), .B(c2628), .Z(n7886) );
XOR U13145 ( .A(c2629), .B(n7887), .Z(c2630) );
ANDN U13146 ( .B(n7888), .A(n7889), .Z(n7887) );
XOR U13147 ( .A(c2629), .B(b[2629]), .Z(n7888) );
XNOR U13148 ( .A(b[2629]), .B(n7889), .Z(c[2629]) );
XNOR U13149 ( .A(a[2629]), .B(c2629), .Z(n7889) );
XOR U13150 ( .A(c2630), .B(n7890), .Z(c2631) );
ANDN U13151 ( .B(n7891), .A(n7892), .Z(n7890) );
XOR U13152 ( .A(c2630), .B(b[2630]), .Z(n7891) );
XNOR U13153 ( .A(b[2630]), .B(n7892), .Z(c[2630]) );
XNOR U13154 ( .A(a[2630]), .B(c2630), .Z(n7892) );
XOR U13155 ( .A(c2631), .B(n7893), .Z(c2632) );
ANDN U13156 ( .B(n7894), .A(n7895), .Z(n7893) );
XOR U13157 ( .A(c2631), .B(b[2631]), .Z(n7894) );
XNOR U13158 ( .A(b[2631]), .B(n7895), .Z(c[2631]) );
XNOR U13159 ( .A(a[2631]), .B(c2631), .Z(n7895) );
XOR U13160 ( .A(c2632), .B(n7896), .Z(c2633) );
ANDN U13161 ( .B(n7897), .A(n7898), .Z(n7896) );
XOR U13162 ( .A(c2632), .B(b[2632]), .Z(n7897) );
XNOR U13163 ( .A(b[2632]), .B(n7898), .Z(c[2632]) );
XNOR U13164 ( .A(a[2632]), .B(c2632), .Z(n7898) );
XOR U13165 ( .A(c2633), .B(n7899), .Z(c2634) );
ANDN U13166 ( .B(n7900), .A(n7901), .Z(n7899) );
XOR U13167 ( .A(c2633), .B(b[2633]), .Z(n7900) );
XNOR U13168 ( .A(b[2633]), .B(n7901), .Z(c[2633]) );
XNOR U13169 ( .A(a[2633]), .B(c2633), .Z(n7901) );
XOR U13170 ( .A(c2634), .B(n7902), .Z(c2635) );
ANDN U13171 ( .B(n7903), .A(n7904), .Z(n7902) );
XOR U13172 ( .A(c2634), .B(b[2634]), .Z(n7903) );
XNOR U13173 ( .A(b[2634]), .B(n7904), .Z(c[2634]) );
XNOR U13174 ( .A(a[2634]), .B(c2634), .Z(n7904) );
XOR U13175 ( .A(c2635), .B(n7905), .Z(c2636) );
ANDN U13176 ( .B(n7906), .A(n7907), .Z(n7905) );
XOR U13177 ( .A(c2635), .B(b[2635]), .Z(n7906) );
XNOR U13178 ( .A(b[2635]), .B(n7907), .Z(c[2635]) );
XNOR U13179 ( .A(a[2635]), .B(c2635), .Z(n7907) );
XOR U13180 ( .A(c2636), .B(n7908), .Z(c2637) );
ANDN U13181 ( .B(n7909), .A(n7910), .Z(n7908) );
XOR U13182 ( .A(c2636), .B(b[2636]), .Z(n7909) );
XNOR U13183 ( .A(b[2636]), .B(n7910), .Z(c[2636]) );
XNOR U13184 ( .A(a[2636]), .B(c2636), .Z(n7910) );
XOR U13185 ( .A(c2637), .B(n7911), .Z(c2638) );
ANDN U13186 ( .B(n7912), .A(n7913), .Z(n7911) );
XOR U13187 ( .A(c2637), .B(b[2637]), .Z(n7912) );
XNOR U13188 ( .A(b[2637]), .B(n7913), .Z(c[2637]) );
XNOR U13189 ( .A(a[2637]), .B(c2637), .Z(n7913) );
XOR U13190 ( .A(c2638), .B(n7914), .Z(c2639) );
ANDN U13191 ( .B(n7915), .A(n7916), .Z(n7914) );
XOR U13192 ( .A(c2638), .B(b[2638]), .Z(n7915) );
XNOR U13193 ( .A(b[2638]), .B(n7916), .Z(c[2638]) );
XNOR U13194 ( .A(a[2638]), .B(c2638), .Z(n7916) );
XOR U13195 ( .A(c2639), .B(n7917), .Z(c2640) );
ANDN U13196 ( .B(n7918), .A(n7919), .Z(n7917) );
XOR U13197 ( .A(c2639), .B(b[2639]), .Z(n7918) );
XNOR U13198 ( .A(b[2639]), .B(n7919), .Z(c[2639]) );
XNOR U13199 ( .A(a[2639]), .B(c2639), .Z(n7919) );
XOR U13200 ( .A(c2640), .B(n7920), .Z(c2641) );
ANDN U13201 ( .B(n7921), .A(n7922), .Z(n7920) );
XOR U13202 ( .A(c2640), .B(b[2640]), .Z(n7921) );
XNOR U13203 ( .A(b[2640]), .B(n7922), .Z(c[2640]) );
XNOR U13204 ( .A(a[2640]), .B(c2640), .Z(n7922) );
XOR U13205 ( .A(c2641), .B(n7923), .Z(c2642) );
ANDN U13206 ( .B(n7924), .A(n7925), .Z(n7923) );
XOR U13207 ( .A(c2641), .B(b[2641]), .Z(n7924) );
XNOR U13208 ( .A(b[2641]), .B(n7925), .Z(c[2641]) );
XNOR U13209 ( .A(a[2641]), .B(c2641), .Z(n7925) );
XOR U13210 ( .A(c2642), .B(n7926), .Z(c2643) );
ANDN U13211 ( .B(n7927), .A(n7928), .Z(n7926) );
XOR U13212 ( .A(c2642), .B(b[2642]), .Z(n7927) );
XNOR U13213 ( .A(b[2642]), .B(n7928), .Z(c[2642]) );
XNOR U13214 ( .A(a[2642]), .B(c2642), .Z(n7928) );
XOR U13215 ( .A(c2643), .B(n7929), .Z(c2644) );
ANDN U13216 ( .B(n7930), .A(n7931), .Z(n7929) );
XOR U13217 ( .A(c2643), .B(b[2643]), .Z(n7930) );
XNOR U13218 ( .A(b[2643]), .B(n7931), .Z(c[2643]) );
XNOR U13219 ( .A(a[2643]), .B(c2643), .Z(n7931) );
XOR U13220 ( .A(c2644), .B(n7932), .Z(c2645) );
ANDN U13221 ( .B(n7933), .A(n7934), .Z(n7932) );
XOR U13222 ( .A(c2644), .B(b[2644]), .Z(n7933) );
XNOR U13223 ( .A(b[2644]), .B(n7934), .Z(c[2644]) );
XNOR U13224 ( .A(a[2644]), .B(c2644), .Z(n7934) );
XOR U13225 ( .A(c2645), .B(n7935), .Z(c2646) );
ANDN U13226 ( .B(n7936), .A(n7937), .Z(n7935) );
XOR U13227 ( .A(c2645), .B(b[2645]), .Z(n7936) );
XNOR U13228 ( .A(b[2645]), .B(n7937), .Z(c[2645]) );
XNOR U13229 ( .A(a[2645]), .B(c2645), .Z(n7937) );
XOR U13230 ( .A(c2646), .B(n7938), .Z(c2647) );
ANDN U13231 ( .B(n7939), .A(n7940), .Z(n7938) );
XOR U13232 ( .A(c2646), .B(b[2646]), .Z(n7939) );
XNOR U13233 ( .A(b[2646]), .B(n7940), .Z(c[2646]) );
XNOR U13234 ( .A(a[2646]), .B(c2646), .Z(n7940) );
XOR U13235 ( .A(c2647), .B(n7941), .Z(c2648) );
ANDN U13236 ( .B(n7942), .A(n7943), .Z(n7941) );
XOR U13237 ( .A(c2647), .B(b[2647]), .Z(n7942) );
XNOR U13238 ( .A(b[2647]), .B(n7943), .Z(c[2647]) );
XNOR U13239 ( .A(a[2647]), .B(c2647), .Z(n7943) );
XOR U13240 ( .A(c2648), .B(n7944), .Z(c2649) );
ANDN U13241 ( .B(n7945), .A(n7946), .Z(n7944) );
XOR U13242 ( .A(c2648), .B(b[2648]), .Z(n7945) );
XNOR U13243 ( .A(b[2648]), .B(n7946), .Z(c[2648]) );
XNOR U13244 ( .A(a[2648]), .B(c2648), .Z(n7946) );
XOR U13245 ( .A(c2649), .B(n7947), .Z(c2650) );
ANDN U13246 ( .B(n7948), .A(n7949), .Z(n7947) );
XOR U13247 ( .A(c2649), .B(b[2649]), .Z(n7948) );
XNOR U13248 ( .A(b[2649]), .B(n7949), .Z(c[2649]) );
XNOR U13249 ( .A(a[2649]), .B(c2649), .Z(n7949) );
XOR U13250 ( .A(c2650), .B(n7950), .Z(c2651) );
ANDN U13251 ( .B(n7951), .A(n7952), .Z(n7950) );
XOR U13252 ( .A(c2650), .B(b[2650]), .Z(n7951) );
XNOR U13253 ( .A(b[2650]), .B(n7952), .Z(c[2650]) );
XNOR U13254 ( .A(a[2650]), .B(c2650), .Z(n7952) );
XOR U13255 ( .A(c2651), .B(n7953), .Z(c2652) );
ANDN U13256 ( .B(n7954), .A(n7955), .Z(n7953) );
XOR U13257 ( .A(c2651), .B(b[2651]), .Z(n7954) );
XNOR U13258 ( .A(b[2651]), .B(n7955), .Z(c[2651]) );
XNOR U13259 ( .A(a[2651]), .B(c2651), .Z(n7955) );
XOR U13260 ( .A(c2652), .B(n7956), .Z(c2653) );
ANDN U13261 ( .B(n7957), .A(n7958), .Z(n7956) );
XOR U13262 ( .A(c2652), .B(b[2652]), .Z(n7957) );
XNOR U13263 ( .A(b[2652]), .B(n7958), .Z(c[2652]) );
XNOR U13264 ( .A(a[2652]), .B(c2652), .Z(n7958) );
XOR U13265 ( .A(c2653), .B(n7959), .Z(c2654) );
ANDN U13266 ( .B(n7960), .A(n7961), .Z(n7959) );
XOR U13267 ( .A(c2653), .B(b[2653]), .Z(n7960) );
XNOR U13268 ( .A(b[2653]), .B(n7961), .Z(c[2653]) );
XNOR U13269 ( .A(a[2653]), .B(c2653), .Z(n7961) );
XOR U13270 ( .A(c2654), .B(n7962), .Z(c2655) );
ANDN U13271 ( .B(n7963), .A(n7964), .Z(n7962) );
XOR U13272 ( .A(c2654), .B(b[2654]), .Z(n7963) );
XNOR U13273 ( .A(b[2654]), .B(n7964), .Z(c[2654]) );
XNOR U13274 ( .A(a[2654]), .B(c2654), .Z(n7964) );
XOR U13275 ( .A(c2655), .B(n7965), .Z(c2656) );
ANDN U13276 ( .B(n7966), .A(n7967), .Z(n7965) );
XOR U13277 ( .A(c2655), .B(b[2655]), .Z(n7966) );
XNOR U13278 ( .A(b[2655]), .B(n7967), .Z(c[2655]) );
XNOR U13279 ( .A(a[2655]), .B(c2655), .Z(n7967) );
XOR U13280 ( .A(c2656), .B(n7968), .Z(c2657) );
ANDN U13281 ( .B(n7969), .A(n7970), .Z(n7968) );
XOR U13282 ( .A(c2656), .B(b[2656]), .Z(n7969) );
XNOR U13283 ( .A(b[2656]), .B(n7970), .Z(c[2656]) );
XNOR U13284 ( .A(a[2656]), .B(c2656), .Z(n7970) );
XOR U13285 ( .A(c2657), .B(n7971), .Z(c2658) );
ANDN U13286 ( .B(n7972), .A(n7973), .Z(n7971) );
XOR U13287 ( .A(c2657), .B(b[2657]), .Z(n7972) );
XNOR U13288 ( .A(b[2657]), .B(n7973), .Z(c[2657]) );
XNOR U13289 ( .A(a[2657]), .B(c2657), .Z(n7973) );
XOR U13290 ( .A(c2658), .B(n7974), .Z(c2659) );
ANDN U13291 ( .B(n7975), .A(n7976), .Z(n7974) );
XOR U13292 ( .A(c2658), .B(b[2658]), .Z(n7975) );
XNOR U13293 ( .A(b[2658]), .B(n7976), .Z(c[2658]) );
XNOR U13294 ( .A(a[2658]), .B(c2658), .Z(n7976) );
XOR U13295 ( .A(c2659), .B(n7977), .Z(c2660) );
ANDN U13296 ( .B(n7978), .A(n7979), .Z(n7977) );
XOR U13297 ( .A(c2659), .B(b[2659]), .Z(n7978) );
XNOR U13298 ( .A(b[2659]), .B(n7979), .Z(c[2659]) );
XNOR U13299 ( .A(a[2659]), .B(c2659), .Z(n7979) );
XOR U13300 ( .A(c2660), .B(n7980), .Z(c2661) );
ANDN U13301 ( .B(n7981), .A(n7982), .Z(n7980) );
XOR U13302 ( .A(c2660), .B(b[2660]), .Z(n7981) );
XNOR U13303 ( .A(b[2660]), .B(n7982), .Z(c[2660]) );
XNOR U13304 ( .A(a[2660]), .B(c2660), .Z(n7982) );
XOR U13305 ( .A(c2661), .B(n7983), .Z(c2662) );
ANDN U13306 ( .B(n7984), .A(n7985), .Z(n7983) );
XOR U13307 ( .A(c2661), .B(b[2661]), .Z(n7984) );
XNOR U13308 ( .A(b[2661]), .B(n7985), .Z(c[2661]) );
XNOR U13309 ( .A(a[2661]), .B(c2661), .Z(n7985) );
XOR U13310 ( .A(c2662), .B(n7986), .Z(c2663) );
ANDN U13311 ( .B(n7987), .A(n7988), .Z(n7986) );
XOR U13312 ( .A(c2662), .B(b[2662]), .Z(n7987) );
XNOR U13313 ( .A(b[2662]), .B(n7988), .Z(c[2662]) );
XNOR U13314 ( .A(a[2662]), .B(c2662), .Z(n7988) );
XOR U13315 ( .A(c2663), .B(n7989), .Z(c2664) );
ANDN U13316 ( .B(n7990), .A(n7991), .Z(n7989) );
XOR U13317 ( .A(c2663), .B(b[2663]), .Z(n7990) );
XNOR U13318 ( .A(b[2663]), .B(n7991), .Z(c[2663]) );
XNOR U13319 ( .A(a[2663]), .B(c2663), .Z(n7991) );
XOR U13320 ( .A(c2664), .B(n7992), .Z(c2665) );
ANDN U13321 ( .B(n7993), .A(n7994), .Z(n7992) );
XOR U13322 ( .A(c2664), .B(b[2664]), .Z(n7993) );
XNOR U13323 ( .A(b[2664]), .B(n7994), .Z(c[2664]) );
XNOR U13324 ( .A(a[2664]), .B(c2664), .Z(n7994) );
XOR U13325 ( .A(c2665), .B(n7995), .Z(c2666) );
ANDN U13326 ( .B(n7996), .A(n7997), .Z(n7995) );
XOR U13327 ( .A(c2665), .B(b[2665]), .Z(n7996) );
XNOR U13328 ( .A(b[2665]), .B(n7997), .Z(c[2665]) );
XNOR U13329 ( .A(a[2665]), .B(c2665), .Z(n7997) );
XOR U13330 ( .A(c2666), .B(n7998), .Z(c2667) );
ANDN U13331 ( .B(n7999), .A(n8000), .Z(n7998) );
XOR U13332 ( .A(c2666), .B(b[2666]), .Z(n7999) );
XNOR U13333 ( .A(b[2666]), .B(n8000), .Z(c[2666]) );
XNOR U13334 ( .A(a[2666]), .B(c2666), .Z(n8000) );
XOR U13335 ( .A(c2667), .B(n8001), .Z(c2668) );
ANDN U13336 ( .B(n8002), .A(n8003), .Z(n8001) );
XOR U13337 ( .A(c2667), .B(b[2667]), .Z(n8002) );
XNOR U13338 ( .A(b[2667]), .B(n8003), .Z(c[2667]) );
XNOR U13339 ( .A(a[2667]), .B(c2667), .Z(n8003) );
XOR U13340 ( .A(c2668), .B(n8004), .Z(c2669) );
ANDN U13341 ( .B(n8005), .A(n8006), .Z(n8004) );
XOR U13342 ( .A(c2668), .B(b[2668]), .Z(n8005) );
XNOR U13343 ( .A(b[2668]), .B(n8006), .Z(c[2668]) );
XNOR U13344 ( .A(a[2668]), .B(c2668), .Z(n8006) );
XOR U13345 ( .A(c2669), .B(n8007), .Z(c2670) );
ANDN U13346 ( .B(n8008), .A(n8009), .Z(n8007) );
XOR U13347 ( .A(c2669), .B(b[2669]), .Z(n8008) );
XNOR U13348 ( .A(b[2669]), .B(n8009), .Z(c[2669]) );
XNOR U13349 ( .A(a[2669]), .B(c2669), .Z(n8009) );
XOR U13350 ( .A(c2670), .B(n8010), .Z(c2671) );
ANDN U13351 ( .B(n8011), .A(n8012), .Z(n8010) );
XOR U13352 ( .A(c2670), .B(b[2670]), .Z(n8011) );
XNOR U13353 ( .A(b[2670]), .B(n8012), .Z(c[2670]) );
XNOR U13354 ( .A(a[2670]), .B(c2670), .Z(n8012) );
XOR U13355 ( .A(c2671), .B(n8013), .Z(c2672) );
ANDN U13356 ( .B(n8014), .A(n8015), .Z(n8013) );
XOR U13357 ( .A(c2671), .B(b[2671]), .Z(n8014) );
XNOR U13358 ( .A(b[2671]), .B(n8015), .Z(c[2671]) );
XNOR U13359 ( .A(a[2671]), .B(c2671), .Z(n8015) );
XOR U13360 ( .A(c2672), .B(n8016), .Z(c2673) );
ANDN U13361 ( .B(n8017), .A(n8018), .Z(n8016) );
XOR U13362 ( .A(c2672), .B(b[2672]), .Z(n8017) );
XNOR U13363 ( .A(b[2672]), .B(n8018), .Z(c[2672]) );
XNOR U13364 ( .A(a[2672]), .B(c2672), .Z(n8018) );
XOR U13365 ( .A(c2673), .B(n8019), .Z(c2674) );
ANDN U13366 ( .B(n8020), .A(n8021), .Z(n8019) );
XOR U13367 ( .A(c2673), .B(b[2673]), .Z(n8020) );
XNOR U13368 ( .A(b[2673]), .B(n8021), .Z(c[2673]) );
XNOR U13369 ( .A(a[2673]), .B(c2673), .Z(n8021) );
XOR U13370 ( .A(c2674), .B(n8022), .Z(c2675) );
ANDN U13371 ( .B(n8023), .A(n8024), .Z(n8022) );
XOR U13372 ( .A(c2674), .B(b[2674]), .Z(n8023) );
XNOR U13373 ( .A(b[2674]), .B(n8024), .Z(c[2674]) );
XNOR U13374 ( .A(a[2674]), .B(c2674), .Z(n8024) );
XOR U13375 ( .A(c2675), .B(n8025), .Z(c2676) );
ANDN U13376 ( .B(n8026), .A(n8027), .Z(n8025) );
XOR U13377 ( .A(c2675), .B(b[2675]), .Z(n8026) );
XNOR U13378 ( .A(b[2675]), .B(n8027), .Z(c[2675]) );
XNOR U13379 ( .A(a[2675]), .B(c2675), .Z(n8027) );
XOR U13380 ( .A(c2676), .B(n8028), .Z(c2677) );
ANDN U13381 ( .B(n8029), .A(n8030), .Z(n8028) );
XOR U13382 ( .A(c2676), .B(b[2676]), .Z(n8029) );
XNOR U13383 ( .A(b[2676]), .B(n8030), .Z(c[2676]) );
XNOR U13384 ( .A(a[2676]), .B(c2676), .Z(n8030) );
XOR U13385 ( .A(c2677), .B(n8031), .Z(c2678) );
ANDN U13386 ( .B(n8032), .A(n8033), .Z(n8031) );
XOR U13387 ( .A(c2677), .B(b[2677]), .Z(n8032) );
XNOR U13388 ( .A(b[2677]), .B(n8033), .Z(c[2677]) );
XNOR U13389 ( .A(a[2677]), .B(c2677), .Z(n8033) );
XOR U13390 ( .A(c2678), .B(n8034), .Z(c2679) );
ANDN U13391 ( .B(n8035), .A(n8036), .Z(n8034) );
XOR U13392 ( .A(c2678), .B(b[2678]), .Z(n8035) );
XNOR U13393 ( .A(b[2678]), .B(n8036), .Z(c[2678]) );
XNOR U13394 ( .A(a[2678]), .B(c2678), .Z(n8036) );
XOR U13395 ( .A(c2679), .B(n8037), .Z(c2680) );
ANDN U13396 ( .B(n8038), .A(n8039), .Z(n8037) );
XOR U13397 ( .A(c2679), .B(b[2679]), .Z(n8038) );
XNOR U13398 ( .A(b[2679]), .B(n8039), .Z(c[2679]) );
XNOR U13399 ( .A(a[2679]), .B(c2679), .Z(n8039) );
XOR U13400 ( .A(c2680), .B(n8040), .Z(c2681) );
ANDN U13401 ( .B(n8041), .A(n8042), .Z(n8040) );
XOR U13402 ( .A(c2680), .B(b[2680]), .Z(n8041) );
XNOR U13403 ( .A(b[2680]), .B(n8042), .Z(c[2680]) );
XNOR U13404 ( .A(a[2680]), .B(c2680), .Z(n8042) );
XOR U13405 ( .A(c2681), .B(n8043), .Z(c2682) );
ANDN U13406 ( .B(n8044), .A(n8045), .Z(n8043) );
XOR U13407 ( .A(c2681), .B(b[2681]), .Z(n8044) );
XNOR U13408 ( .A(b[2681]), .B(n8045), .Z(c[2681]) );
XNOR U13409 ( .A(a[2681]), .B(c2681), .Z(n8045) );
XOR U13410 ( .A(c2682), .B(n8046), .Z(c2683) );
ANDN U13411 ( .B(n8047), .A(n8048), .Z(n8046) );
XOR U13412 ( .A(c2682), .B(b[2682]), .Z(n8047) );
XNOR U13413 ( .A(b[2682]), .B(n8048), .Z(c[2682]) );
XNOR U13414 ( .A(a[2682]), .B(c2682), .Z(n8048) );
XOR U13415 ( .A(c2683), .B(n8049), .Z(c2684) );
ANDN U13416 ( .B(n8050), .A(n8051), .Z(n8049) );
XOR U13417 ( .A(c2683), .B(b[2683]), .Z(n8050) );
XNOR U13418 ( .A(b[2683]), .B(n8051), .Z(c[2683]) );
XNOR U13419 ( .A(a[2683]), .B(c2683), .Z(n8051) );
XOR U13420 ( .A(c2684), .B(n8052), .Z(c2685) );
ANDN U13421 ( .B(n8053), .A(n8054), .Z(n8052) );
XOR U13422 ( .A(c2684), .B(b[2684]), .Z(n8053) );
XNOR U13423 ( .A(b[2684]), .B(n8054), .Z(c[2684]) );
XNOR U13424 ( .A(a[2684]), .B(c2684), .Z(n8054) );
XOR U13425 ( .A(c2685), .B(n8055), .Z(c2686) );
ANDN U13426 ( .B(n8056), .A(n8057), .Z(n8055) );
XOR U13427 ( .A(c2685), .B(b[2685]), .Z(n8056) );
XNOR U13428 ( .A(b[2685]), .B(n8057), .Z(c[2685]) );
XNOR U13429 ( .A(a[2685]), .B(c2685), .Z(n8057) );
XOR U13430 ( .A(c2686), .B(n8058), .Z(c2687) );
ANDN U13431 ( .B(n8059), .A(n8060), .Z(n8058) );
XOR U13432 ( .A(c2686), .B(b[2686]), .Z(n8059) );
XNOR U13433 ( .A(b[2686]), .B(n8060), .Z(c[2686]) );
XNOR U13434 ( .A(a[2686]), .B(c2686), .Z(n8060) );
XOR U13435 ( .A(c2687), .B(n8061), .Z(c2688) );
ANDN U13436 ( .B(n8062), .A(n8063), .Z(n8061) );
XOR U13437 ( .A(c2687), .B(b[2687]), .Z(n8062) );
XNOR U13438 ( .A(b[2687]), .B(n8063), .Z(c[2687]) );
XNOR U13439 ( .A(a[2687]), .B(c2687), .Z(n8063) );
XOR U13440 ( .A(c2688), .B(n8064), .Z(c2689) );
ANDN U13441 ( .B(n8065), .A(n8066), .Z(n8064) );
XOR U13442 ( .A(c2688), .B(b[2688]), .Z(n8065) );
XNOR U13443 ( .A(b[2688]), .B(n8066), .Z(c[2688]) );
XNOR U13444 ( .A(a[2688]), .B(c2688), .Z(n8066) );
XOR U13445 ( .A(c2689), .B(n8067), .Z(c2690) );
ANDN U13446 ( .B(n8068), .A(n8069), .Z(n8067) );
XOR U13447 ( .A(c2689), .B(b[2689]), .Z(n8068) );
XNOR U13448 ( .A(b[2689]), .B(n8069), .Z(c[2689]) );
XNOR U13449 ( .A(a[2689]), .B(c2689), .Z(n8069) );
XOR U13450 ( .A(c2690), .B(n8070), .Z(c2691) );
ANDN U13451 ( .B(n8071), .A(n8072), .Z(n8070) );
XOR U13452 ( .A(c2690), .B(b[2690]), .Z(n8071) );
XNOR U13453 ( .A(b[2690]), .B(n8072), .Z(c[2690]) );
XNOR U13454 ( .A(a[2690]), .B(c2690), .Z(n8072) );
XOR U13455 ( .A(c2691), .B(n8073), .Z(c2692) );
ANDN U13456 ( .B(n8074), .A(n8075), .Z(n8073) );
XOR U13457 ( .A(c2691), .B(b[2691]), .Z(n8074) );
XNOR U13458 ( .A(b[2691]), .B(n8075), .Z(c[2691]) );
XNOR U13459 ( .A(a[2691]), .B(c2691), .Z(n8075) );
XOR U13460 ( .A(c2692), .B(n8076), .Z(c2693) );
ANDN U13461 ( .B(n8077), .A(n8078), .Z(n8076) );
XOR U13462 ( .A(c2692), .B(b[2692]), .Z(n8077) );
XNOR U13463 ( .A(b[2692]), .B(n8078), .Z(c[2692]) );
XNOR U13464 ( .A(a[2692]), .B(c2692), .Z(n8078) );
XOR U13465 ( .A(c2693), .B(n8079), .Z(c2694) );
ANDN U13466 ( .B(n8080), .A(n8081), .Z(n8079) );
XOR U13467 ( .A(c2693), .B(b[2693]), .Z(n8080) );
XNOR U13468 ( .A(b[2693]), .B(n8081), .Z(c[2693]) );
XNOR U13469 ( .A(a[2693]), .B(c2693), .Z(n8081) );
XOR U13470 ( .A(c2694), .B(n8082), .Z(c2695) );
ANDN U13471 ( .B(n8083), .A(n8084), .Z(n8082) );
XOR U13472 ( .A(c2694), .B(b[2694]), .Z(n8083) );
XNOR U13473 ( .A(b[2694]), .B(n8084), .Z(c[2694]) );
XNOR U13474 ( .A(a[2694]), .B(c2694), .Z(n8084) );
XOR U13475 ( .A(c2695), .B(n8085), .Z(c2696) );
ANDN U13476 ( .B(n8086), .A(n8087), .Z(n8085) );
XOR U13477 ( .A(c2695), .B(b[2695]), .Z(n8086) );
XNOR U13478 ( .A(b[2695]), .B(n8087), .Z(c[2695]) );
XNOR U13479 ( .A(a[2695]), .B(c2695), .Z(n8087) );
XOR U13480 ( .A(c2696), .B(n8088), .Z(c2697) );
ANDN U13481 ( .B(n8089), .A(n8090), .Z(n8088) );
XOR U13482 ( .A(c2696), .B(b[2696]), .Z(n8089) );
XNOR U13483 ( .A(b[2696]), .B(n8090), .Z(c[2696]) );
XNOR U13484 ( .A(a[2696]), .B(c2696), .Z(n8090) );
XOR U13485 ( .A(c2697), .B(n8091), .Z(c2698) );
ANDN U13486 ( .B(n8092), .A(n8093), .Z(n8091) );
XOR U13487 ( .A(c2697), .B(b[2697]), .Z(n8092) );
XNOR U13488 ( .A(b[2697]), .B(n8093), .Z(c[2697]) );
XNOR U13489 ( .A(a[2697]), .B(c2697), .Z(n8093) );
XOR U13490 ( .A(c2698), .B(n8094), .Z(c2699) );
ANDN U13491 ( .B(n8095), .A(n8096), .Z(n8094) );
XOR U13492 ( .A(c2698), .B(b[2698]), .Z(n8095) );
XNOR U13493 ( .A(b[2698]), .B(n8096), .Z(c[2698]) );
XNOR U13494 ( .A(a[2698]), .B(c2698), .Z(n8096) );
XOR U13495 ( .A(c2699), .B(n8097), .Z(c2700) );
ANDN U13496 ( .B(n8098), .A(n8099), .Z(n8097) );
XOR U13497 ( .A(c2699), .B(b[2699]), .Z(n8098) );
XNOR U13498 ( .A(b[2699]), .B(n8099), .Z(c[2699]) );
XNOR U13499 ( .A(a[2699]), .B(c2699), .Z(n8099) );
XOR U13500 ( .A(c2700), .B(n8100), .Z(c2701) );
ANDN U13501 ( .B(n8101), .A(n8102), .Z(n8100) );
XOR U13502 ( .A(c2700), .B(b[2700]), .Z(n8101) );
XNOR U13503 ( .A(b[2700]), .B(n8102), .Z(c[2700]) );
XNOR U13504 ( .A(a[2700]), .B(c2700), .Z(n8102) );
XOR U13505 ( .A(c2701), .B(n8103), .Z(c2702) );
ANDN U13506 ( .B(n8104), .A(n8105), .Z(n8103) );
XOR U13507 ( .A(c2701), .B(b[2701]), .Z(n8104) );
XNOR U13508 ( .A(b[2701]), .B(n8105), .Z(c[2701]) );
XNOR U13509 ( .A(a[2701]), .B(c2701), .Z(n8105) );
XOR U13510 ( .A(c2702), .B(n8106), .Z(c2703) );
ANDN U13511 ( .B(n8107), .A(n8108), .Z(n8106) );
XOR U13512 ( .A(c2702), .B(b[2702]), .Z(n8107) );
XNOR U13513 ( .A(b[2702]), .B(n8108), .Z(c[2702]) );
XNOR U13514 ( .A(a[2702]), .B(c2702), .Z(n8108) );
XOR U13515 ( .A(c2703), .B(n8109), .Z(c2704) );
ANDN U13516 ( .B(n8110), .A(n8111), .Z(n8109) );
XOR U13517 ( .A(c2703), .B(b[2703]), .Z(n8110) );
XNOR U13518 ( .A(b[2703]), .B(n8111), .Z(c[2703]) );
XNOR U13519 ( .A(a[2703]), .B(c2703), .Z(n8111) );
XOR U13520 ( .A(c2704), .B(n8112), .Z(c2705) );
ANDN U13521 ( .B(n8113), .A(n8114), .Z(n8112) );
XOR U13522 ( .A(c2704), .B(b[2704]), .Z(n8113) );
XNOR U13523 ( .A(b[2704]), .B(n8114), .Z(c[2704]) );
XNOR U13524 ( .A(a[2704]), .B(c2704), .Z(n8114) );
XOR U13525 ( .A(c2705), .B(n8115), .Z(c2706) );
ANDN U13526 ( .B(n8116), .A(n8117), .Z(n8115) );
XOR U13527 ( .A(c2705), .B(b[2705]), .Z(n8116) );
XNOR U13528 ( .A(b[2705]), .B(n8117), .Z(c[2705]) );
XNOR U13529 ( .A(a[2705]), .B(c2705), .Z(n8117) );
XOR U13530 ( .A(c2706), .B(n8118), .Z(c2707) );
ANDN U13531 ( .B(n8119), .A(n8120), .Z(n8118) );
XOR U13532 ( .A(c2706), .B(b[2706]), .Z(n8119) );
XNOR U13533 ( .A(b[2706]), .B(n8120), .Z(c[2706]) );
XNOR U13534 ( .A(a[2706]), .B(c2706), .Z(n8120) );
XOR U13535 ( .A(c2707), .B(n8121), .Z(c2708) );
ANDN U13536 ( .B(n8122), .A(n8123), .Z(n8121) );
XOR U13537 ( .A(c2707), .B(b[2707]), .Z(n8122) );
XNOR U13538 ( .A(b[2707]), .B(n8123), .Z(c[2707]) );
XNOR U13539 ( .A(a[2707]), .B(c2707), .Z(n8123) );
XOR U13540 ( .A(c2708), .B(n8124), .Z(c2709) );
ANDN U13541 ( .B(n8125), .A(n8126), .Z(n8124) );
XOR U13542 ( .A(c2708), .B(b[2708]), .Z(n8125) );
XNOR U13543 ( .A(b[2708]), .B(n8126), .Z(c[2708]) );
XNOR U13544 ( .A(a[2708]), .B(c2708), .Z(n8126) );
XOR U13545 ( .A(c2709), .B(n8127), .Z(c2710) );
ANDN U13546 ( .B(n8128), .A(n8129), .Z(n8127) );
XOR U13547 ( .A(c2709), .B(b[2709]), .Z(n8128) );
XNOR U13548 ( .A(b[2709]), .B(n8129), .Z(c[2709]) );
XNOR U13549 ( .A(a[2709]), .B(c2709), .Z(n8129) );
XOR U13550 ( .A(c2710), .B(n8130), .Z(c2711) );
ANDN U13551 ( .B(n8131), .A(n8132), .Z(n8130) );
XOR U13552 ( .A(c2710), .B(b[2710]), .Z(n8131) );
XNOR U13553 ( .A(b[2710]), .B(n8132), .Z(c[2710]) );
XNOR U13554 ( .A(a[2710]), .B(c2710), .Z(n8132) );
XOR U13555 ( .A(c2711), .B(n8133), .Z(c2712) );
ANDN U13556 ( .B(n8134), .A(n8135), .Z(n8133) );
XOR U13557 ( .A(c2711), .B(b[2711]), .Z(n8134) );
XNOR U13558 ( .A(b[2711]), .B(n8135), .Z(c[2711]) );
XNOR U13559 ( .A(a[2711]), .B(c2711), .Z(n8135) );
XOR U13560 ( .A(c2712), .B(n8136), .Z(c2713) );
ANDN U13561 ( .B(n8137), .A(n8138), .Z(n8136) );
XOR U13562 ( .A(c2712), .B(b[2712]), .Z(n8137) );
XNOR U13563 ( .A(b[2712]), .B(n8138), .Z(c[2712]) );
XNOR U13564 ( .A(a[2712]), .B(c2712), .Z(n8138) );
XOR U13565 ( .A(c2713), .B(n8139), .Z(c2714) );
ANDN U13566 ( .B(n8140), .A(n8141), .Z(n8139) );
XOR U13567 ( .A(c2713), .B(b[2713]), .Z(n8140) );
XNOR U13568 ( .A(b[2713]), .B(n8141), .Z(c[2713]) );
XNOR U13569 ( .A(a[2713]), .B(c2713), .Z(n8141) );
XOR U13570 ( .A(c2714), .B(n8142), .Z(c2715) );
ANDN U13571 ( .B(n8143), .A(n8144), .Z(n8142) );
XOR U13572 ( .A(c2714), .B(b[2714]), .Z(n8143) );
XNOR U13573 ( .A(b[2714]), .B(n8144), .Z(c[2714]) );
XNOR U13574 ( .A(a[2714]), .B(c2714), .Z(n8144) );
XOR U13575 ( .A(c2715), .B(n8145), .Z(c2716) );
ANDN U13576 ( .B(n8146), .A(n8147), .Z(n8145) );
XOR U13577 ( .A(c2715), .B(b[2715]), .Z(n8146) );
XNOR U13578 ( .A(b[2715]), .B(n8147), .Z(c[2715]) );
XNOR U13579 ( .A(a[2715]), .B(c2715), .Z(n8147) );
XOR U13580 ( .A(c2716), .B(n8148), .Z(c2717) );
ANDN U13581 ( .B(n8149), .A(n8150), .Z(n8148) );
XOR U13582 ( .A(c2716), .B(b[2716]), .Z(n8149) );
XNOR U13583 ( .A(b[2716]), .B(n8150), .Z(c[2716]) );
XNOR U13584 ( .A(a[2716]), .B(c2716), .Z(n8150) );
XOR U13585 ( .A(c2717), .B(n8151), .Z(c2718) );
ANDN U13586 ( .B(n8152), .A(n8153), .Z(n8151) );
XOR U13587 ( .A(c2717), .B(b[2717]), .Z(n8152) );
XNOR U13588 ( .A(b[2717]), .B(n8153), .Z(c[2717]) );
XNOR U13589 ( .A(a[2717]), .B(c2717), .Z(n8153) );
XOR U13590 ( .A(c2718), .B(n8154), .Z(c2719) );
ANDN U13591 ( .B(n8155), .A(n8156), .Z(n8154) );
XOR U13592 ( .A(c2718), .B(b[2718]), .Z(n8155) );
XNOR U13593 ( .A(b[2718]), .B(n8156), .Z(c[2718]) );
XNOR U13594 ( .A(a[2718]), .B(c2718), .Z(n8156) );
XOR U13595 ( .A(c2719), .B(n8157), .Z(c2720) );
ANDN U13596 ( .B(n8158), .A(n8159), .Z(n8157) );
XOR U13597 ( .A(c2719), .B(b[2719]), .Z(n8158) );
XNOR U13598 ( .A(b[2719]), .B(n8159), .Z(c[2719]) );
XNOR U13599 ( .A(a[2719]), .B(c2719), .Z(n8159) );
XOR U13600 ( .A(c2720), .B(n8160), .Z(c2721) );
ANDN U13601 ( .B(n8161), .A(n8162), .Z(n8160) );
XOR U13602 ( .A(c2720), .B(b[2720]), .Z(n8161) );
XNOR U13603 ( .A(b[2720]), .B(n8162), .Z(c[2720]) );
XNOR U13604 ( .A(a[2720]), .B(c2720), .Z(n8162) );
XOR U13605 ( .A(c2721), .B(n8163), .Z(c2722) );
ANDN U13606 ( .B(n8164), .A(n8165), .Z(n8163) );
XOR U13607 ( .A(c2721), .B(b[2721]), .Z(n8164) );
XNOR U13608 ( .A(b[2721]), .B(n8165), .Z(c[2721]) );
XNOR U13609 ( .A(a[2721]), .B(c2721), .Z(n8165) );
XOR U13610 ( .A(c2722), .B(n8166), .Z(c2723) );
ANDN U13611 ( .B(n8167), .A(n8168), .Z(n8166) );
XOR U13612 ( .A(c2722), .B(b[2722]), .Z(n8167) );
XNOR U13613 ( .A(b[2722]), .B(n8168), .Z(c[2722]) );
XNOR U13614 ( .A(a[2722]), .B(c2722), .Z(n8168) );
XOR U13615 ( .A(c2723), .B(n8169), .Z(c2724) );
ANDN U13616 ( .B(n8170), .A(n8171), .Z(n8169) );
XOR U13617 ( .A(c2723), .B(b[2723]), .Z(n8170) );
XNOR U13618 ( .A(b[2723]), .B(n8171), .Z(c[2723]) );
XNOR U13619 ( .A(a[2723]), .B(c2723), .Z(n8171) );
XOR U13620 ( .A(c2724), .B(n8172), .Z(c2725) );
ANDN U13621 ( .B(n8173), .A(n8174), .Z(n8172) );
XOR U13622 ( .A(c2724), .B(b[2724]), .Z(n8173) );
XNOR U13623 ( .A(b[2724]), .B(n8174), .Z(c[2724]) );
XNOR U13624 ( .A(a[2724]), .B(c2724), .Z(n8174) );
XOR U13625 ( .A(c2725), .B(n8175), .Z(c2726) );
ANDN U13626 ( .B(n8176), .A(n8177), .Z(n8175) );
XOR U13627 ( .A(c2725), .B(b[2725]), .Z(n8176) );
XNOR U13628 ( .A(b[2725]), .B(n8177), .Z(c[2725]) );
XNOR U13629 ( .A(a[2725]), .B(c2725), .Z(n8177) );
XOR U13630 ( .A(c2726), .B(n8178), .Z(c2727) );
ANDN U13631 ( .B(n8179), .A(n8180), .Z(n8178) );
XOR U13632 ( .A(c2726), .B(b[2726]), .Z(n8179) );
XNOR U13633 ( .A(b[2726]), .B(n8180), .Z(c[2726]) );
XNOR U13634 ( .A(a[2726]), .B(c2726), .Z(n8180) );
XOR U13635 ( .A(c2727), .B(n8181), .Z(c2728) );
ANDN U13636 ( .B(n8182), .A(n8183), .Z(n8181) );
XOR U13637 ( .A(c2727), .B(b[2727]), .Z(n8182) );
XNOR U13638 ( .A(b[2727]), .B(n8183), .Z(c[2727]) );
XNOR U13639 ( .A(a[2727]), .B(c2727), .Z(n8183) );
XOR U13640 ( .A(c2728), .B(n8184), .Z(c2729) );
ANDN U13641 ( .B(n8185), .A(n8186), .Z(n8184) );
XOR U13642 ( .A(c2728), .B(b[2728]), .Z(n8185) );
XNOR U13643 ( .A(b[2728]), .B(n8186), .Z(c[2728]) );
XNOR U13644 ( .A(a[2728]), .B(c2728), .Z(n8186) );
XOR U13645 ( .A(c2729), .B(n8187), .Z(c2730) );
ANDN U13646 ( .B(n8188), .A(n8189), .Z(n8187) );
XOR U13647 ( .A(c2729), .B(b[2729]), .Z(n8188) );
XNOR U13648 ( .A(b[2729]), .B(n8189), .Z(c[2729]) );
XNOR U13649 ( .A(a[2729]), .B(c2729), .Z(n8189) );
XOR U13650 ( .A(c2730), .B(n8190), .Z(c2731) );
ANDN U13651 ( .B(n8191), .A(n8192), .Z(n8190) );
XOR U13652 ( .A(c2730), .B(b[2730]), .Z(n8191) );
XNOR U13653 ( .A(b[2730]), .B(n8192), .Z(c[2730]) );
XNOR U13654 ( .A(a[2730]), .B(c2730), .Z(n8192) );
XOR U13655 ( .A(c2731), .B(n8193), .Z(c2732) );
ANDN U13656 ( .B(n8194), .A(n8195), .Z(n8193) );
XOR U13657 ( .A(c2731), .B(b[2731]), .Z(n8194) );
XNOR U13658 ( .A(b[2731]), .B(n8195), .Z(c[2731]) );
XNOR U13659 ( .A(a[2731]), .B(c2731), .Z(n8195) );
XOR U13660 ( .A(c2732), .B(n8196), .Z(c2733) );
ANDN U13661 ( .B(n8197), .A(n8198), .Z(n8196) );
XOR U13662 ( .A(c2732), .B(b[2732]), .Z(n8197) );
XNOR U13663 ( .A(b[2732]), .B(n8198), .Z(c[2732]) );
XNOR U13664 ( .A(a[2732]), .B(c2732), .Z(n8198) );
XOR U13665 ( .A(c2733), .B(n8199), .Z(c2734) );
ANDN U13666 ( .B(n8200), .A(n8201), .Z(n8199) );
XOR U13667 ( .A(c2733), .B(b[2733]), .Z(n8200) );
XNOR U13668 ( .A(b[2733]), .B(n8201), .Z(c[2733]) );
XNOR U13669 ( .A(a[2733]), .B(c2733), .Z(n8201) );
XOR U13670 ( .A(c2734), .B(n8202), .Z(c2735) );
ANDN U13671 ( .B(n8203), .A(n8204), .Z(n8202) );
XOR U13672 ( .A(c2734), .B(b[2734]), .Z(n8203) );
XNOR U13673 ( .A(b[2734]), .B(n8204), .Z(c[2734]) );
XNOR U13674 ( .A(a[2734]), .B(c2734), .Z(n8204) );
XOR U13675 ( .A(c2735), .B(n8205), .Z(c2736) );
ANDN U13676 ( .B(n8206), .A(n8207), .Z(n8205) );
XOR U13677 ( .A(c2735), .B(b[2735]), .Z(n8206) );
XNOR U13678 ( .A(b[2735]), .B(n8207), .Z(c[2735]) );
XNOR U13679 ( .A(a[2735]), .B(c2735), .Z(n8207) );
XOR U13680 ( .A(c2736), .B(n8208), .Z(c2737) );
ANDN U13681 ( .B(n8209), .A(n8210), .Z(n8208) );
XOR U13682 ( .A(c2736), .B(b[2736]), .Z(n8209) );
XNOR U13683 ( .A(b[2736]), .B(n8210), .Z(c[2736]) );
XNOR U13684 ( .A(a[2736]), .B(c2736), .Z(n8210) );
XOR U13685 ( .A(c2737), .B(n8211), .Z(c2738) );
ANDN U13686 ( .B(n8212), .A(n8213), .Z(n8211) );
XOR U13687 ( .A(c2737), .B(b[2737]), .Z(n8212) );
XNOR U13688 ( .A(b[2737]), .B(n8213), .Z(c[2737]) );
XNOR U13689 ( .A(a[2737]), .B(c2737), .Z(n8213) );
XOR U13690 ( .A(c2738), .B(n8214), .Z(c2739) );
ANDN U13691 ( .B(n8215), .A(n8216), .Z(n8214) );
XOR U13692 ( .A(c2738), .B(b[2738]), .Z(n8215) );
XNOR U13693 ( .A(b[2738]), .B(n8216), .Z(c[2738]) );
XNOR U13694 ( .A(a[2738]), .B(c2738), .Z(n8216) );
XOR U13695 ( .A(c2739), .B(n8217), .Z(c2740) );
ANDN U13696 ( .B(n8218), .A(n8219), .Z(n8217) );
XOR U13697 ( .A(c2739), .B(b[2739]), .Z(n8218) );
XNOR U13698 ( .A(b[2739]), .B(n8219), .Z(c[2739]) );
XNOR U13699 ( .A(a[2739]), .B(c2739), .Z(n8219) );
XOR U13700 ( .A(c2740), .B(n8220), .Z(c2741) );
ANDN U13701 ( .B(n8221), .A(n8222), .Z(n8220) );
XOR U13702 ( .A(c2740), .B(b[2740]), .Z(n8221) );
XNOR U13703 ( .A(b[2740]), .B(n8222), .Z(c[2740]) );
XNOR U13704 ( .A(a[2740]), .B(c2740), .Z(n8222) );
XOR U13705 ( .A(c2741), .B(n8223), .Z(c2742) );
ANDN U13706 ( .B(n8224), .A(n8225), .Z(n8223) );
XOR U13707 ( .A(c2741), .B(b[2741]), .Z(n8224) );
XNOR U13708 ( .A(b[2741]), .B(n8225), .Z(c[2741]) );
XNOR U13709 ( .A(a[2741]), .B(c2741), .Z(n8225) );
XOR U13710 ( .A(c2742), .B(n8226), .Z(c2743) );
ANDN U13711 ( .B(n8227), .A(n8228), .Z(n8226) );
XOR U13712 ( .A(c2742), .B(b[2742]), .Z(n8227) );
XNOR U13713 ( .A(b[2742]), .B(n8228), .Z(c[2742]) );
XNOR U13714 ( .A(a[2742]), .B(c2742), .Z(n8228) );
XOR U13715 ( .A(c2743), .B(n8229), .Z(c2744) );
ANDN U13716 ( .B(n8230), .A(n8231), .Z(n8229) );
XOR U13717 ( .A(c2743), .B(b[2743]), .Z(n8230) );
XNOR U13718 ( .A(b[2743]), .B(n8231), .Z(c[2743]) );
XNOR U13719 ( .A(a[2743]), .B(c2743), .Z(n8231) );
XOR U13720 ( .A(c2744), .B(n8232), .Z(c2745) );
ANDN U13721 ( .B(n8233), .A(n8234), .Z(n8232) );
XOR U13722 ( .A(c2744), .B(b[2744]), .Z(n8233) );
XNOR U13723 ( .A(b[2744]), .B(n8234), .Z(c[2744]) );
XNOR U13724 ( .A(a[2744]), .B(c2744), .Z(n8234) );
XOR U13725 ( .A(c2745), .B(n8235), .Z(c2746) );
ANDN U13726 ( .B(n8236), .A(n8237), .Z(n8235) );
XOR U13727 ( .A(c2745), .B(b[2745]), .Z(n8236) );
XNOR U13728 ( .A(b[2745]), .B(n8237), .Z(c[2745]) );
XNOR U13729 ( .A(a[2745]), .B(c2745), .Z(n8237) );
XOR U13730 ( .A(c2746), .B(n8238), .Z(c2747) );
ANDN U13731 ( .B(n8239), .A(n8240), .Z(n8238) );
XOR U13732 ( .A(c2746), .B(b[2746]), .Z(n8239) );
XNOR U13733 ( .A(b[2746]), .B(n8240), .Z(c[2746]) );
XNOR U13734 ( .A(a[2746]), .B(c2746), .Z(n8240) );
XOR U13735 ( .A(c2747), .B(n8241), .Z(c2748) );
ANDN U13736 ( .B(n8242), .A(n8243), .Z(n8241) );
XOR U13737 ( .A(c2747), .B(b[2747]), .Z(n8242) );
XNOR U13738 ( .A(b[2747]), .B(n8243), .Z(c[2747]) );
XNOR U13739 ( .A(a[2747]), .B(c2747), .Z(n8243) );
XOR U13740 ( .A(c2748), .B(n8244), .Z(c2749) );
ANDN U13741 ( .B(n8245), .A(n8246), .Z(n8244) );
XOR U13742 ( .A(c2748), .B(b[2748]), .Z(n8245) );
XNOR U13743 ( .A(b[2748]), .B(n8246), .Z(c[2748]) );
XNOR U13744 ( .A(a[2748]), .B(c2748), .Z(n8246) );
XOR U13745 ( .A(c2749), .B(n8247), .Z(c2750) );
ANDN U13746 ( .B(n8248), .A(n8249), .Z(n8247) );
XOR U13747 ( .A(c2749), .B(b[2749]), .Z(n8248) );
XNOR U13748 ( .A(b[2749]), .B(n8249), .Z(c[2749]) );
XNOR U13749 ( .A(a[2749]), .B(c2749), .Z(n8249) );
XOR U13750 ( .A(c2750), .B(n8250), .Z(c2751) );
ANDN U13751 ( .B(n8251), .A(n8252), .Z(n8250) );
XOR U13752 ( .A(c2750), .B(b[2750]), .Z(n8251) );
XNOR U13753 ( .A(b[2750]), .B(n8252), .Z(c[2750]) );
XNOR U13754 ( .A(a[2750]), .B(c2750), .Z(n8252) );
XOR U13755 ( .A(c2751), .B(n8253), .Z(c2752) );
ANDN U13756 ( .B(n8254), .A(n8255), .Z(n8253) );
XOR U13757 ( .A(c2751), .B(b[2751]), .Z(n8254) );
XNOR U13758 ( .A(b[2751]), .B(n8255), .Z(c[2751]) );
XNOR U13759 ( .A(a[2751]), .B(c2751), .Z(n8255) );
XOR U13760 ( .A(c2752), .B(n8256), .Z(c2753) );
ANDN U13761 ( .B(n8257), .A(n8258), .Z(n8256) );
XOR U13762 ( .A(c2752), .B(b[2752]), .Z(n8257) );
XNOR U13763 ( .A(b[2752]), .B(n8258), .Z(c[2752]) );
XNOR U13764 ( .A(a[2752]), .B(c2752), .Z(n8258) );
XOR U13765 ( .A(c2753), .B(n8259), .Z(c2754) );
ANDN U13766 ( .B(n8260), .A(n8261), .Z(n8259) );
XOR U13767 ( .A(c2753), .B(b[2753]), .Z(n8260) );
XNOR U13768 ( .A(b[2753]), .B(n8261), .Z(c[2753]) );
XNOR U13769 ( .A(a[2753]), .B(c2753), .Z(n8261) );
XOR U13770 ( .A(c2754), .B(n8262), .Z(c2755) );
ANDN U13771 ( .B(n8263), .A(n8264), .Z(n8262) );
XOR U13772 ( .A(c2754), .B(b[2754]), .Z(n8263) );
XNOR U13773 ( .A(b[2754]), .B(n8264), .Z(c[2754]) );
XNOR U13774 ( .A(a[2754]), .B(c2754), .Z(n8264) );
XOR U13775 ( .A(c2755), .B(n8265), .Z(c2756) );
ANDN U13776 ( .B(n8266), .A(n8267), .Z(n8265) );
XOR U13777 ( .A(c2755), .B(b[2755]), .Z(n8266) );
XNOR U13778 ( .A(b[2755]), .B(n8267), .Z(c[2755]) );
XNOR U13779 ( .A(a[2755]), .B(c2755), .Z(n8267) );
XOR U13780 ( .A(c2756), .B(n8268), .Z(c2757) );
ANDN U13781 ( .B(n8269), .A(n8270), .Z(n8268) );
XOR U13782 ( .A(c2756), .B(b[2756]), .Z(n8269) );
XNOR U13783 ( .A(b[2756]), .B(n8270), .Z(c[2756]) );
XNOR U13784 ( .A(a[2756]), .B(c2756), .Z(n8270) );
XOR U13785 ( .A(c2757), .B(n8271), .Z(c2758) );
ANDN U13786 ( .B(n8272), .A(n8273), .Z(n8271) );
XOR U13787 ( .A(c2757), .B(b[2757]), .Z(n8272) );
XNOR U13788 ( .A(b[2757]), .B(n8273), .Z(c[2757]) );
XNOR U13789 ( .A(a[2757]), .B(c2757), .Z(n8273) );
XOR U13790 ( .A(c2758), .B(n8274), .Z(c2759) );
ANDN U13791 ( .B(n8275), .A(n8276), .Z(n8274) );
XOR U13792 ( .A(c2758), .B(b[2758]), .Z(n8275) );
XNOR U13793 ( .A(b[2758]), .B(n8276), .Z(c[2758]) );
XNOR U13794 ( .A(a[2758]), .B(c2758), .Z(n8276) );
XOR U13795 ( .A(c2759), .B(n8277), .Z(c2760) );
ANDN U13796 ( .B(n8278), .A(n8279), .Z(n8277) );
XOR U13797 ( .A(c2759), .B(b[2759]), .Z(n8278) );
XNOR U13798 ( .A(b[2759]), .B(n8279), .Z(c[2759]) );
XNOR U13799 ( .A(a[2759]), .B(c2759), .Z(n8279) );
XOR U13800 ( .A(c2760), .B(n8280), .Z(c2761) );
ANDN U13801 ( .B(n8281), .A(n8282), .Z(n8280) );
XOR U13802 ( .A(c2760), .B(b[2760]), .Z(n8281) );
XNOR U13803 ( .A(b[2760]), .B(n8282), .Z(c[2760]) );
XNOR U13804 ( .A(a[2760]), .B(c2760), .Z(n8282) );
XOR U13805 ( .A(c2761), .B(n8283), .Z(c2762) );
ANDN U13806 ( .B(n8284), .A(n8285), .Z(n8283) );
XOR U13807 ( .A(c2761), .B(b[2761]), .Z(n8284) );
XNOR U13808 ( .A(b[2761]), .B(n8285), .Z(c[2761]) );
XNOR U13809 ( .A(a[2761]), .B(c2761), .Z(n8285) );
XOR U13810 ( .A(c2762), .B(n8286), .Z(c2763) );
ANDN U13811 ( .B(n8287), .A(n8288), .Z(n8286) );
XOR U13812 ( .A(c2762), .B(b[2762]), .Z(n8287) );
XNOR U13813 ( .A(b[2762]), .B(n8288), .Z(c[2762]) );
XNOR U13814 ( .A(a[2762]), .B(c2762), .Z(n8288) );
XOR U13815 ( .A(c2763), .B(n8289), .Z(c2764) );
ANDN U13816 ( .B(n8290), .A(n8291), .Z(n8289) );
XOR U13817 ( .A(c2763), .B(b[2763]), .Z(n8290) );
XNOR U13818 ( .A(b[2763]), .B(n8291), .Z(c[2763]) );
XNOR U13819 ( .A(a[2763]), .B(c2763), .Z(n8291) );
XOR U13820 ( .A(c2764), .B(n8292), .Z(c2765) );
ANDN U13821 ( .B(n8293), .A(n8294), .Z(n8292) );
XOR U13822 ( .A(c2764), .B(b[2764]), .Z(n8293) );
XNOR U13823 ( .A(b[2764]), .B(n8294), .Z(c[2764]) );
XNOR U13824 ( .A(a[2764]), .B(c2764), .Z(n8294) );
XOR U13825 ( .A(c2765), .B(n8295), .Z(c2766) );
ANDN U13826 ( .B(n8296), .A(n8297), .Z(n8295) );
XOR U13827 ( .A(c2765), .B(b[2765]), .Z(n8296) );
XNOR U13828 ( .A(b[2765]), .B(n8297), .Z(c[2765]) );
XNOR U13829 ( .A(a[2765]), .B(c2765), .Z(n8297) );
XOR U13830 ( .A(c2766), .B(n8298), .Z(c2767) );
ANDN U13831 ( .B(n8299), .A(n8300), .Z(n8298) );
XOR U13832 ( .A(c2766), .B(b[2766]), .Z(n8299) );
XNOR U13833 ( .A(b[2766]), .B(n8300), .Z(c[2766]) );
XNOR U13834 ( .A(a[2766]), .B(c2766), .Z(n8300) );
XOR U13835 ( .A(c2767), .B(n8301), .Z(c2768) );
ANDN U13836 ( .B(n8302), .A(n8303), .Z(n8301) );
XOR U13837 ( .A(c2767), .B(b[2767]), .Z(n8302) );
XNOR U13838 ( .A(b[2767]), .B(n8303), .Z(c[2767]) );
XNOR U13839 ( .A(a[2767]), .B(c2767), .Z(n8303) );
XOR U13840 ( .A(c2768), .B(n8304), .Z(c2769) );
ANDN U13841 ( .B(n8305), .A(n8306), .Z(n8304) );
XOR U13842 ( .A(c2768), .B(b[2768]), .Z(n8305) );
XNOR U13843 ( .A(b[2768]), .B(n8306), .Z(c[2768]) );
XNOR U13844 ( .A(a[2768]), .B(c2768), .Z(n8306) );
XOR U13845 ( .A(c2769), .B(n8307), .Z(c2770) );
ANDN U13846 ( .B(n8308), .A(n8309), .Z(n8307) );
XOR U13847 ( .A(c2769), .B(b[2769]), .Z(n8308) );
XNOR U13848 ( .A(b[2769]), .B(n8309), .Z(c[2769]) );
XNOR U13849 ( .A(a[2769]), .B(c2769), .Z(n8309) );
XOR U13850 ( .A(c2770), .B(n8310), .Z(c2771) );
ANDN U13851 ( .B(n8311), .A(n8312), .Z(n8310) );
XOR U13852 ( .A(c2770), .B(b[2770]), .Z(n8311) );
XNOR U13853 ( .A(b[2770]), .B(n8312), .Z(c[2770]) );
XNOR U13854 ( .A(a[2770]), .B(c2770), .Z(n8312) );
XOR U13855 ( .A(c2771), .B(n8313), .Z(c2772) );
ANDN U13856 ( .B(n8314), .A(n8315), .Z(n8313) );
XOR U13857 ( .A(c2771), .B(b[2771]), .Z(n8314) );
XNOR U13858 ( .A(b[2771]), .B(n8315), .Z(c[2771]) );
XNOR U13859 ( .A(a[2771]), .B(c2771), .Z(n8315) );
XOR U13860 ( .A(c2772), .B(n8316), .Z(c2773) );
ANDN U13861 ( .B(n8317), .A(n8318), .Z(n8316) );
XOR U13862 ( .A(c2772), .B(b[2772]), .Z(n8317) );
XNOR U13863 ( .A(b[2772]), .B(n8318), .Z(c[2772]) );
XNOR U13864 ( .A(a[2772]), .B(c2772), .Z(n8318) );
XOR U13865 ( .A(c2773), .B(n8319), .Z(c2774) );
ANDN U13866 ( .B(n8320), .A(n8321), .Z(n8319) );
XOR U13867 ( .A(c2773), .B(b[2773]), .Z(n8320) );
XNOR U13868 ( .A(b[2773]), .B(n8321), .Z(c[2773]) );
XNOR U13869 ( .A(a[2773]), .B(c2773), .Z(n8321) );
XOR U13870 ( .A(c2774), .B(n8322), .Z(c2775) );
ANDN U13871 ( .B(n8323), .A(n8324), .Z(n8322) );
XOR U13872 ( .A(c2774), .B(b[2774]), .Z(n8323) );
XNOR U13873 ( .A(b[2774]), .B(n8324), .Z(c[2774]) );
XNOR U13874 ( .A(a[2774]), .B(c2774), .Z(n8324) );
XOR U13875 ( .A(c2775), .B(n8325), .Z(c2776) );
ANDN U13876 ( .B(n8326), .A(n8327), .Z(n8325) );
XOR U13877 ( .A(c2775), .B(b[2775]), .Z(n8326) );
XNOR U13878 ( .A(b[2775]), .B(n8327), .Z(c[2775]) );
XNOR U13879 ( .A(a[2775]), .B(c2775), .Z(n8327) );
XOR U13880 ( .A(c2776), .B(n8328), .Z(c2777) );
ANDN U13881 ( .B(n8329), .A(n8330), .Z(n8328) );
XOR U13882 ( .A(c2776), .B(b[2776]), .Z(n8329) );
XNOR U13883 ( .A(b[2776]), .B(n8330), .Z(c[2776]) );
XNOR U13884 ( .A(a[2776]), .B(c2776), .Z(n8330) );
XOR U13885 ( .A(c2777), .B(n8331), .Z(c2778) );
ANDN U13886 ( .B(n8332), .A(n8333), .Z(n8331) );
XOR U13887 ( .A(c2777), .B(b[2777]), .Z(n8332) );
XNOR U13888 ( .A(b[2777]), .B(n8333), .Z(c[2777]) );
XNOR U13889 ( .A(a[2777]), .B(c2777), .Z(n8333) );
XOR U13890 ( .A(c2778), .B(n8334), .Z(c2779) );
ANDN U13891 ( .B(n8335), .A(n8336), .Z(n8334) );
XOR U13892 ( .A(c2778), .B(b[2778]), .Z(n8335) );
XNOR U13893 ( .A(b[2778]), .B(n8336), .Z(c[2778]) );
XNOR U13894 ( .A(a[2778]), .B(c2778), .Z(n8336) );
XOR U13895 ( .A(c2779), .B(n8337), .Z(c2780) );
ANDN U13896 ( .B(n8338), .A(n8339), .Z(n8337) );
XOR U13897 ( .A(c2779), .B(b[2779]), .Z(n8338) );
XNOR U13898 ( .A(b[2779]), .B(n8339), .Z(c[2779]) );
XNOR U13899 ( .A(a[2779]), .B(c2779), .Z(n8339) );
XOR U13900 ( .A(c2780), .B(n8340), .Z(c2781) );
ANDN U13901 ( .B(n8341), .A(n8342), .Z(n8340) );
XOR U13902 ( .A(c2780), .B(b[2780]), .Z(n8341) );
XNOR U13903 ( .A(b[2780]), .B(n8342), .Z(c[2780]) );
XNOR U13904 ( .A(a[2780]), .B(c2780), .Z(n8342) );
XOR U13905 ( .A(c2781), .B(n8343), .Z(c2782) );
ANDN U13906 ( .B(n8344), .A(n8345), .Z(n8343) );
XOR U13907 ( .A(c2781), .B(b[2781]), .Z(n8344) );
XNOR U13908 ( .A(b[2781]), .B(n8345), .Z(c[2781]) );
XNOR U13909 ( .A(a[2781]), .B(c2781), .Z(n8345) );
XOR U13910 ( .A(c2782), .B(n8346), .Z(c2783) );
ANDN U13911 ( .B(n8347), .A(n8348), .Z(n8346) );
XOR U13912 ( .A(c2782), .B(b[2782]), .Z(n8347) );
XNOR U13913 ( .A(b[2782]), .B(n8348), .Z(c[2782]) );
XNOR U13914 ( .A(a[2782]), .B(c2782), .Z(n8348) );
XOR U13915 ( .A(c2783), .B(n8349), .Z(c2784) );
ANDN U13916 ( .B(n8350), .A(n8351), .Z(n8349) );
XOR U13917 ( .A(c2783), .B(b[2783]), .Z(n8350) );
XNOR U13918 ( .A(b[2783]), .B(n8351), .Z(c[2783]) );
XNOR U13919 ( .A(a[2783]), .B(c2783), .Z(n8351) );
XOR U13920 ( .A(c2784), .B(n8352), .Z(c2785) );
ANDN U13921 ( .B(n8353), .A(n8354), .Z(n8352) );
XOR U13922 ( .A(c2784), .B(b[2784]), .Z(n8353) );
XNOR U13923 ( .A(b[2784]), .B(n8354), .Z(c[2784]) );
XNOR U13924 ( .A(a[2784]), .B(c2784), .Z(n8354) );
XOR U13925 ( .A(c2785), .B(n8355), .Z(c2786) );
ANDN U13926 ( .B(n8356), .A(n8357), .Z(n8355) );
XOR U13927 ( .A(c2785), .B(b[2785]), .Z(n8356) );
XNOR U13928 ( .A(b[2785]), .B(n8357), .Z(c[2785]) );
XNOR U13929 ( .A(a[2785]), .B(c2785), .Z(n8357) );
XOR U13930 ( .A(c2786), .B(n8358), .Z(c2787) );
ANDN U13931 ( .B(n8359), .A(n8360), .Z(n8358) );
XOR U13932 ( .A(c2786), .B(b[2786]), .Z(n8359) );
XNOR U13933 ( .A(b[2786]), .B(n8360), .Z(c[2786]) );
XNOR U13934 ( .A(a[2786]), .B(c2786), .Z(n8360) );
XOR U13935 ( .A(c2787), .B(n8361), .Z(c2788) );
ANDN U13936 ( .B(n8362), .A(n8363), .Z(n8361) );
XOR U13937 ( .A(c2787), .B(b[2787]), .Z(n8362) );
XNOR U13938 ( .A(b[2787]), .B(n8363), .Z(c[2787]) );
XNOR U13939 ( .A(a[2787]), .B(c2787), .Z(n8363) );
XOR U13940 ( .A(c2788), .B(n8364), .Z(c2789) );
ANDN U13941 ( .B(n8365), .A(n8366), .Z(n8364) );
XOR U13942 ( .A(c2788), .B(b[2788]), .Z(n8365) );
XNOR U13943 ( .A(b[2788]), .B(n8366), .Z(c[2788]) );
XNOR U13944 ( .A(a[2788]), .B(c2788), .Z(n8366) );
XOR U13945 ( .A(c2789), .B(n8367), .Z(c2790) );
ANDN U13946 ( .B(n8368), .A(n8369), .Z(n8367) );
XOR U13947 ( .A(c2789), .B(b[2789]), .Z(n8368) );
XNOR U13948 ( .A(b[2789]), .B(n8369), .Z(c[2789]) );
XNOR U13949 ( .A(a[2789]), .B(c2789), .Z(n8369) );
XOR U13950 ( .A(c2790), .B(n8370), .Z(c2791) );
ANDN U13951 ( .B(n8371), .A(n8372), .Z(n8370) );
XOR U13952 ( .A(c2790), .B(b[2790]), .Z(n8371) );
XNOR U13953 ( .A(b[2790]), .B(n8372), .Z(c[2790]) );
XNOR U13954 ( .A(a[2790]), .B(c2790), .Z(n8372) );
XOR U13955 ( .A(c2791), .B(n8373), .Z(c2792) );
ANDN U13956 ( .B(n8374), .A(n8375), .Z(n8373) );
XOR U13957 ( .A(c2791), .B(b[2791]), .Z(n8374) );
XNOR U13958 ( .A(b[2791]), .B(n8375), .Z(c[2791]) );
XNOR U13959 ( .A(a[2791]), .B(c2791), .Z(n8375) );
XOR U13960 ( .A(c2792), .B(n8376), .Z(c2793) );
ANDN U13961 ( .B(n8377), .A(n8378), .Z(n8376) );
XOR U13962 ( .A(c2792), .B(b[2792]), .Z(n8377) );
XNOR U13963 ( .A(b[2792]), .B(n8378), .Z(c[2792]) );
XNOR U13964 ( .A(a[2792]), .B(c2792), .Z(n8378) );
XOR U13965 ( .A(c2793), .B(n8379), .Z(c2794) );
ANDN U13966 ( .B(n8380), .A(n8381), .Z(n8379) );
XOR U13967 ( .A(c2793), .B(b[2793]), .Z(n8380) );
XNOR U13968 ( .A(b[2793]), .B(n8381), .Z(c[2793]) );
XNOR U13969 ( .A(a[2793]), .B(c2793), .Z(n8381) );
XOR U13970 ( .A(c2794), .B(n8382), .Z(c2795) );
ANDN U13971 ( .B(n8383), .A(n8384), .Z(n8382) );
XOR U13972 ( .A(c2794), .B(b[2794]), .Z(n8383) );
XNOR U13973 ( .A(b[2794]), .B(n8384), .Z(c[2794]) );
XNOR U13974 ( .A(a[2794]), .B(c2794), .Z(n8384) );
XOR U13975 ( .A(c2795), .B(n8385), .Z(c2796) );
ANDN U13976 ( .B(n8386), .A(n8387), .Z(n8385) );
XOR U13977 ( .A(c2795), .B(b[2795]), .Z(n8386) );
XNOR U13978 ( .A(b[2795]), .B(n8387), .Z(c[2795]) );
XNOR U13979 ( .A(a[2795]), .B(c2795), .Z(n8387) );
XOR U13980 ( .A(c2796), .B(n8388), .Z(c2797) );
ANDN U13981 ( .B(n8389), .A(n8390), .Z(n8388) );
XOR U13982 ( .A(c2796), .B(b[2796]), .Z(n8389) );
XNOR U13983 ( .A(b[2796]), .B(n8390), .Z(c[2796]) );
XNOR U13984 ( .A(a[2796]), .B(c2796), .Z(n8390) );
XOR U13985 ( .A(c2797), .B(n8391), .Z(c2798) );
ANDN U13986 ( .B(n8392), .A(n8393), .Z(n8391) );
XOR U13987 ( .A(c2797), .B(b[2797]), .Z(n8392) );
XNOR U13988 ( .A(b[2797]), .B(n8393), .Z(c[2797]) );
XNOR U13989 ( .A(a[2797]), .B(c2797), .Z(n8393) );
XOR U13990 ( .A(c2798), .B(n8394), .Z(c2799) );
ANDN U13991 ( .B(n8395), .A(n8396), .Z(n8394) );
XOR U13992 ( .A(c2798), .B(b[2798]), .Z(n8395) );
XNOR U13993 ( .A(b[2798]), .B(n8396), .Z(c[2798]) );
XNOR U13994 ( .A(a[2798]), .B(c2798), .Z(n8396) );
XOR U13995 ( .A(c2799), .B(n8397), .Z(c2800) );
ANDN U13996 ( .B(n8398), .A(n8399), .Z(n8397) );
XOR U13997 ( .A(c2799), .B(b[2799]), .Z(n8398) );
XNOR U13998 ( .A(b[2799]), .B(n8399), .Z(c[2799]) );
XNOR U13999 ( .A(a[2799]), .B(c2799), .Z(n8399) );
XOR U14000 ( .A(c2800), .B(n8400), .Z(c2801) );
ANDN U14001 ( .B(n8401), .A(n8402), .Z(n8400) );
XOR U14002 ( .A(c2800), .B(b[2800]), .Z(n8401) );
XNOR U14003 ( .A(b[2800]), .B(n8402), .Z(c[2800]) );
XNOR U14004 ( .A(a[2800]), .B(c2800), .Z(n8402) );
XOR U14005 ( .A(c2801), .B(n8403), .Z(c2802) );
ANDN U14006 ( .B(n8404), .A(n8405), .Z(n8403) );
XOR U14007 ( .A(c2801), .B(b[2801]), .Z(n8404) );
XNOR U14008 ( .A(b[2801]), .B(n8405), .Z(c[2801]) );
XNOR U14009 ( .A(a[2801]), .B(c2801), .Z(n8405) );
XOR U14010 ( .A(c2802), .B(n8406), .Z(c2803) );
ANDN U14011 ( .B(n8407), .A(n8408), .Z(n8406) );
XOR U14012 ( .A(c2802), .B(b[2802]), .Z(n8407) );
XNOR U14013 ( .A(b[2802]), .B(n8408), .Z(c[2802]) );
XNOR U14014 ( .A(a[2802]), .B(c2802), .Z(n8408) );
XOR U14015 ( .A(c2803), .B(n8409), .Z(c2804) );
ANDN U14016 ( .B(n8410), .A(n8411), .Z(n8409) );
XOR U14017 ( .A(c2803), .B(b[2803]), .Z(n8410) );
XNOR U14018 ( .A(b[2803]), .B(n8411), .Z(c[2803]) );
XNOR U14019 ( .A(a[2803]), .B(c2803), .Z(n8411) );
XOR U14020 ( .A(c2804), .B(n8412), .Z(c2805) );
ANDN U14021 ( .B(n8413), .A(n8414), .Z(n8412) );
XOR U14022 ( .A(c2804), .B(b[2804]), .Z(n8413) );
XNOR U14023 ( .A(b[2804]), .B(n8414), .Z(c[2804]) );
XNOR U14024 ( .A(a[2804]), .B(c2804), .Z(n8414) );
XOR U14025 ( .A(c2805), .B(n8415), .Z(c2806) );
ANDN U14026 ( .B(n8416), .A(n8417), .Z(n8415) );
XOR U14027 ( .A(c2805), .B(b[2805]), .Z(n8416) );
XNOR U14028 ( .A(b[2805]), .B(n8417), .Z(c[2805]) );
XNOR U14029 ( .A(a[2805]), .B(c2805), .Z(n8417) );
XOR U14030 ( .A(c2806), .B(n8418), .Z(c2807) );
ANDN U14031 ( .B(n8419), .A(n8420), .Z(n8418) );
XOR U14032 ( .A(c2806), .B(b[2806]), .Z(n8419) );
XNOR U14033 ( .A(b[2806]), .B(n8420), .Z(c[2806]) );
XNOR U14034 ( .A(a[2806]), .B(c2806), .Z(n8420) );
XOR U14035 ( .A(c2807), .B(n8421), .Z(c2808) );
ANDN U14036 ( .B(n8422), .A(n8423), .Z(n8421) );
XOR U14037 ( .A(c2807), .B(b[2807]), .Z(n8422) );
XNOR U14038 ( .A(b[2807]), .B(n8423), .Z(c[2807]) );
XNOR U14039 ( .A(a[2807]), .B(c2807), .Z(n8423) );
XOR U14040 ( .A(c2808), .B(n8424), .Z(c2809) );
ANDN U14041 ( .B(n8425), .A(n8426), .Z(n8424) );
XOR U14042 ( .A(c2808), .B(b[2808]), .Z(n8425) );
XNOR U14043 ( .A(b[2808]), .B(n8426), .Z(c[2808]) );
XNOR U14044 ( .A(a[2808]), .B(c2808), .Z(n8426) );
XOR U14045 ( .A(c2809), .B(n8427), .Z(c2810) );
ANDN U14046 ( .B(n8428), .A(n8429), .Z(n8427) );
XOR U14047 ( .A(c2809), .B(b[2809]), .Z(n8428) );
XNOR U14048 ( .A(b[2809]), .B(n8429), .Z(c[2809]) );
XNOR U14049 ( .A(a[2809]), .B(c2809), .Z(n8429) );
XOR U14050 ( .A(c2810), .B(n8430), .Z(c2811) );
ANDN U14051 ( .B(n8431), .A(n8432), .Z(n8430) );
XOR U14052 ( .A(c2810), .B(b[2810]), .Z(n8431) );
XNOR U14053 ( .A(b[2810]), .B(n8432), .Z(c[2810]) );
XNOR U14054 ( .A(a[2810]), .B(c2810), .Z(n8432) );
XOR U14055 ( .A(c2811), .B(n8433), .Z(c2812) );
ANDN U14056 ( .B(n8434), .A(n8435), .Z(n8433) );
XOR U14057 ( .A(c2811), .B(b[2811]), .Z(n8434) );
XNOR U14058 ( .A(b[2811]), .B(n8435), .Z(c[2811]) );
XNOR U14059 ( .A(a[2811]), .B(c2811), .Z(n8435) );
XOR U14060 ( .A(c2812), .B(n8436), .Z(c2813) );
ANDN U14061 ( .B(n8437), .A(n8438), .Z(n8436) );
XOR U14062 ( .A(c2812), .B(b[2812]), .Z(n8437) );
XNOR U14063 ( .A(b[2812]), .B(n8438), .Z(c[2812]) );
XNOR U14064 ( .A(a[2812]), .B(c2812), .Z(n8438) );
XOR U14065 ( .A(c2813), .B(n8439), .Z(c2814) );
ANDN U14066 ( .B(n8440), .A(n8441), .Z(n8439) );
XOR U14067 ( .A(c2813), .B(b[2813]), .Z(n8440) );
XNOR U14068 ( .A(b[2813]), .B(n8441), .Z(c[2813]) );
XNOR U14069 ( .A(a[2813]), .B(c2813), .Z(n8441) );
XOR U14070 ( .A(c2814), .B(n8442), .Z(c2815) );
ANDN U14071 ( .B(n8443), .A(n8444), .Z(n8442) );
XOR U14072 ( .A(c2814), .B(b[2814]), .Z(n8443) );
XNOR U14073 ( .A(b[2814]), .B(n8444), .Z(c[2814]) );
XNOR U14074 ( .A(a[2814]), .B(c2814), .Z(n8444) );
XOR U14075 ( .A(c2815), .B(n8445), .Z(c2816) );
ANDN U14076 ( .B(n8446), .A(n8447), .Z(n8445) );
XOR U14077 ( .A(c2815), .B(b[2815]), .Z(n8446) );
XNOR U14078 ( .A(b[2815]), .B(n8447), .Z(c[2815]) );
XNOR U14079 ( .A(a[2815]), .B(c2815), .Z(n8447) );
XOR U14080 ( .A(c2816), .B(n8448), .Z(c2817) );
ANDN U14081 ( .B(n8449), .A(n8450), .Z(n8448) );
XOR U14082 ( .A(c2816), .B(b[2816]), .Z(n8449) );
XNOR U14083 ( .A(b[2816]), .B(n8450), .Z(c[2816]) );
XNOR U14084 ( .A(a[2816]), .B(c2816), .Z(n8450) );
XOR U14085 ( .A(c2817), .B(n8451), .Z(c2818) );
ANDN U14086 ( .B(n8452), .A(n8453), .Z(n8451) );
XOR U14087 ( .A(c2817), .B(b[2817]), .Z(n8452) );
XNOR U14088 ( .A(b[2817]), .B(n8453), .Z(c[2817]) );
XNOR U14089 ( .A(a[2817]), .B(c2817), .Z(n8453) );
XOR U14090 ( .A(c2818), .B(n8454), .Z(c2819) );
ANDN U14091 ( .B(n8455), .A(n8456), .Z(n8454) );
XOR U14092 ( .A(c2818), .B(b[2818]), .Z(n8455) );
XNOR U14093 ( .A(b[2818]), .B(n8456), .Z(c[2818]) );
XNOR U14094 ( .A(a[2818]), .B(c2818), .Z(n8456) );
XOR U14095 ( .A(c2819), .B(n8457), .Z(c2820) );
ANDN U14096 ( .B(n8458), .A(n8459), .Z(n8457) );
XOR U14097 ( .A(c2819), .B(b[2819]), .Z(n8458) );
XNOR U14098 ( .A(b[2819]), .B(n8459), .Z(c[2819]) );
XNOR U14099 ( .A(a[2819]), .B(c2819), .Z(n8459) );
XOR U14100 ( .A(c2820), .B(n8460), .Z(c2821) );
ANDN U14101 ( .B(n8461), .A(n8462), .Z(n8460) );
XOR U14102 ( .A(c2820), .B(b[2820]), .Z(n8461) );
XNOR U14103 ( .A(b[2820]), .B(n8462), .Z(c[2820]) );
XNOR U14104 ( .A(a[2820]), .B(c2820), .Z(n8462) );
XOR U14105 ( .A(c2821), .B(n8463), .Z(c2822) );
ANDN U14106 ( .B(n8464), .A(n8465), .Z(n8463) );
XOR U14107 ( .A(c2821), .B(b[2821]), .Z(n8464) );
XNOR U14108 ( .A(b[2821]), .B(n8465), .Z(c[2821]) );
XNOR U14109 ( .A(a[2821]), .B(c2821), .Z(n8465) );
XOR U14110 ( .A(c2822), .B(n8466), .Z(c2823) );
ANDN U14111 ( .B(n8467), .A(n8468), .Z(n8466) );
XOR U14112 ( .A(c2822), .B(b[2822]), .Z(n8467) );
XNOR U14113 ( .A(b[2822]), .B(n8468), .Z(c[2822]) );
XNOR U14114 ( .A(a[2822]), .B(c2822), .Z(n8468) );
XOR U14115 ( .A(c2823), .B(n8469), .Z(c2824) );
ANDN U14116 ( .B(n8470), .A(n8471), .Z(n8469) );
XOR U14117 ( .A(c2823), .B(b[2823]), .Z(n8470) );
XNOR U14118 ( .A(b[2823]), .B(n8471), .Z(c[2823]) );
XNOR U14119 ( .A(a[2823]), .B(c2823), .Z(n8471) );
XOR U14120 ( .A(c2824), .B(n8472), .Z(c2825) );
ANDN U14121 ( .B(n8473), .A(n8474), .Z(n8472) );
XOR U14122 ( .A(c2824), .B(b[2824]), .Z(n8473) );
XNOR U14123 ( .A(b[2824]), .B(n8474), .Z(c[2824]) );
XNOR U14124 ( .A(a[2824]), .B(c2824), .Z(n8474) );
XOR U14125 ( .A(c2825), .B(n8475), .Z(c2826) );
ANDN U14126 ( .B(n8476), .A(n8477), .Z(n8475) );
XOR U14127 ( .A(c2825), .B(b[2825]), .Z(n8476) );
XNOR U14128 ( .A(b[2825]), .B(n8477), .Z(c[2825]) );
XNOR U14129 ( .A(a[2825]), .B(c2825), .Z(n8477) );
XOR U14130 ( .A(c2826), .B(n8478), .Z(c2827) );
ANDN U14131 ( .B(n8479), .A(n8480), .Z(n8478) );
XOR U14132 ( .A(c2826), .B(b[2826]), .Z(n8479) );
XNOR U14133 ( .A(b[2826]), .B(n8480), .Z(c[2826]) );
XNOR U14134 ( .A(a[2826]), .B(c2826), .Z(n8480) );
XOR U14135 ( .A(c2827), .B(n8481), .Z(c2828) );
ANDN U14136 ( .B(n8482), .A(n8483), .Z(n8481) );
XOR U14137 ( .A(c2827), .B(b[2827]), .Z(n8482) );
XNOR U14138 ( .A(b[2827]), .B(n8483), .Z(c[2827]) );
XNOR U14139 ( .A(a[2827]), .B(c2827), .Z(n8483) );
XOR U14140 ( .A(c2828), .B(n8484), .Z(c2829) );
ANDN U14141 ( .B(n8485), .A(n8486), .Z(n8484) );
XOR U14142 ( .A(c2828), .B(b[2828]), .Z(n8485) );
XNOR U14143 ( .A(b[2828]), .B(n8486), .Z(c[2828]) );
XNOR U14144 ( .A(a[2828]), .B(c2828), .Z(n8486) );
XOR U14145 ( .A(c2829), .B(n8487), .Z(c2830) );
ANDN U14146 ( .B(n8488), .A(n8489), .Z(n8487) );
XOR U14147 ( .A(c2829), .B(b[2829]), .Z(n8488) );
XNOR U14148 ( .A(b[2829]), .B(n8489), .Z(c[2829]) );
XNOR U14149 ( .A(a[2829]), .B(c2829), .Z(n8489) );
XOR U14150 ( .A(c2830), .B(n8490), .Z(c2831) );
ANDN U14151 ( .B(n8491), .A(n8492), .Z(n8490) );
XOR U14152 ( .A(c2830), .B(b[2830]), .Z(n8491) );
XNOR U14153 ( .A(b[2830]), .B(n8492), .Z(c[2830]) );
XNOR U14154 ( .A(a[2830]), .B(c2830), .Z(n8492) );
XOR U14155 ( .A(c2831), .B(n8493), .Z(c2832) );
ANDN U14156 ( .B(n8494), .A(n8495), .Z(n8493) );
XOR U14157 ( .A(c2831), .B(b[2831]), .Z(n8494) );
XNOR U14158 ( .A(b[2831]), .B(n8495), .Z(c[2831]) );
XNOR U14159 ( .A(a[2831]), .B(c2831), .Z(n8495) );
XOR U14160 ( .A(c2832), .B(n8496), .Z(c2833) );
ANDN U14161 ( .B(n8497), .A(n8498), .Z(n8496) );
XOR U14162 ( .A(c2832), .B(b[2832]), .Z(n8497) );
XNOR U14163 ( .A(b[2832]), .B(n8498), .Z(c[2832]) );
XNOR U14164 ( .A(a[2832]), .B(c2832), .Z(n8498) );
XOR U14165 ( .A(c2833), .B(n8499), .Z(c2834) );
ANDN U14166 ( .B(n8500), .A(n8501), .Z(n8499) );
XOR U14167 ( .A(c2833), .B(b[2833]), .Z(n8500) );
XNOR U14168 ( .A(b[2833]), .B(n8501), .Z(c[2833]) );
XNOR U14169 ( .A(a[2833]), .B(c2833), .Z(n8501) );
XOR U14170 ( .A(c2834), .B(n8502), .Z(c2835) );
ANDN U14171 ( .B(n8503), .A(n8504), .Z(n8502) );
XOR U14172 ( .A(c2834), .B(b[2834]), .Z(n8503) );
XNOR U14173 ( .A(b[2834]), .B(n8504), .Z(c[2834]) );
XNOR U14174 ( .A(a[2834]), .B(c2834), .Z(n8504) );
XOR U14175 ( .A(c2835), .B(n8505), .Z(c2836) );
ANDN U14176 ( .B(n8506), .A(n8507), .Z(n8505) );
XOR U14177 ( .A(c2835), .B(b[2835]), .Z(n8506) );
XNOR U14178 ( .A(b[2835]), .B(n8507), .Z(c[2835]) );
XNOR U14179 ( .A(a[2835]), .B(c2835), .Z(n8507) );
XOR U14180 ( .A(c2836), .B(n8508), .Z(c2837) );
ANDN U14181 ( .B(n8509), .A(n8510), .Z(n8508) );
XOR U14182 ( .A(c2836), .B(b[2836]), .Z(n8509) );
XNOR U14183 ( .A(b[2836]), .B(n8510), .Z(c[2836]) );
XNOR U14184 ( .A(a[2836]), .B(c2836), .Z(n8510) );
XOR U14185 ( .A(c2837), .B(n8511), .Z(c2838) );
ANDN U14186 ( .B(n8512), .A(n8513), .Z(n8511) );
XOR U14187 ( .A(c2837), .B(b[2837]), .Z(n8512) );
XNOR U14188 ( .A(b[2837]), .B(n8513), .Z(c[2837]) );
XNOR U14189 ( .A(a[2837]), .B(c2837), .Z(n8513) );
XOR U14190 ( .A(c2838), .B(n8514), .Z(c2839) );
ANDN U14191 ( .B(n8515), .A(n8516), .Z(n8514) );
XOR U14192 ( .A(c2838), .B(b[2838]), .Z(n8515) );
XNOR U14193 ( .A(b[2838]), .B(n8516), .Z(c[2838]) );
XNOR U14194 ( .A(a[2838]), .B(c2838), .Z(n8516) );
XOR U14195 ( .A(c2839), .B(n8517), .Z(c2840) );
ANDN U14196 ( .B(n8518), .A(n8519), .Z(n8517) );
XOR U14197 ( .A(c2839), .B(b[2839]), .Z(n8518) );
XNOR U14198 ( .A(b[2839]), .B(n8519), .Z(c[2839]) );
XNOR U14199 ( .A(a[2839]), .B(c2839), .Z(n8519) );
XOR U14200 ( .A(c2840), .B(n8520), .Z(c2841) );
ANDN U14201 ( .B(n8521), .A(n8522), .Z(n8520) );
XOR U14202 ( .A(c2840), .B(b[2840]), .Z(n8521) );
XNOR U14203 ( .A(b[2840]), .B(n8522), .Z(c[2840]) );
XNOR U14204 ( .A(a[2840]), .B(c2840), .Z(n8522) );
XOR U14205 ( .A(c2841), .B(n8523), .Z(c2842) );
ANDN U14206 ( .B(n8524), .A(n8525), .Z(n8523) );
XOR U14207 ( .A(c2841), .B(b[2841]), .Z(n8524) );
XNOR U14208 ( .A(b[2841]), .B(n8525), .Z(c[2841]) );
XNOR U14209 ( .A(a[2841]), .B(c2841), .Z(n8525) );
XOR U14210 ( .A(c2842), .B(n8526), .Z(c2843) );
ANDN U14211 ( .B(n8527), .A(n8528), .Z(n8526) );
XOR U14212 ( .A(c2842), .B(b[2842]), .Z(n8527) );
XNOR U14213 ( .A(b[2842]), .B(n8528), .Z(c[2842]) );
XNOR U14214 ( .A(a[2842]), .B(c2842), .Z(n8528) );
XOR U14215 ( .A(c2843), .B(n8529), .Z(c2844) );
ANDN U14216 ( .B(n8530), .A(n8531), .Z(n8529) );
XOR U14217 ( .A(c2843), .B(b[2843]), .Z(n8530) );
XNOR U14218 ( .A(b[2843]), .B(n8531), .Z(c[2843]) );
XNOR U14219 ( .A(a[2843]), .B(c2843), .Z(n8531) );
XOR U14220 ( .A(c2844), .B(n8532), .Z(c2845) );
ANDN U14221 ( .B(n8533), .A(n8534), .Z(n8532) );
XOR U14222 ( .A(c2844), .B(b[2844]), .Z(n8533) );
XNOR U14223 ( .A(b[2844]), .B(n8534), .Z(c[2844]) );
XNOR U14224 ( .A(a[2844]), .B(c2844), .Z(n8534) );
XOR U14225 ( .A(c2845), .B(n8535), .Z(c2846) );
ANDN U14226 ( .B(n8536), .A(n8537), .Z(n8535) );
XOR U14227 ( .A(c2845), .B(b[2845]), .Z(n8536) );
XNOR U14228 ( .A(b[2845]), .B(n8537), .Z(c[2845]) );
XNOR U14229 ( .A(a[2845]), .B(c2845), .Z(n8537) );
XOR U14230 ( .A(c2846), .B(n8538), .Z(c2847) );
ANDN U14231 ( .B(n8539), .A(n8540), .Z(n8538) );
XOR U14232 ( .A(c2846), .B(b[2846]), .Z(n8539) );
XNOR U14233 ( .A(b[2846]), .B(n8540), .Z(c[2846]) );
XNOR U14234 ( .A(a[2846]), .B(c2846), .Z(n8540) );
XOR U14235 ( .A(c2847), .B(n8541), .Z(c2848) );
ANDN U14236 ( .B(n8542), .A(n8543), .Z(n8541) );
XOR U14237 ( .A(c2847), .B(b[2847]), .Z(n8542) );
XNOR U14238 ( .A(b[2847]), .B(n8543), .Z(c[2847]) );
XNOR U14239 ( .A(a[2847]), .B(c2847), .Z(n8543) );
XOR U14240 ( .A(c2848), .B(n8544), .Z(c2849) );
ANDN U14241 ( .B(n8545), .A(n8546), .Z(n8544) );
XOR U14242 ( .A(c2848), .B(b[2848]), .Z(n8545) );
XNOR U14243 ( .A(b[2848]), .B(n8546), .Z(c[2848]) );
XNOR U14244 ( .A(a[2848]), .B(c2848), .Z(n8546) );
XOR U14245 ( .A(c2849), .B(n8547), .Z(c2850) );
ANDN U14246 ( .B(n8548), .A(n8549), .Z(n8547) );
XOR U14247 ( .A(c2849), .B(b[2849]), .Z(n8548) );
XNOR U14248 ( .A(b[2849]), .B(n8549), .Z(c[2849]) );
XNOR U14249 ( .A(a[2849]), .B(c2849), .Z(n8549) );
XOR U14250 ( .A(c2850), .B(n8550), .Z(c2851) );
ANDN U14251 ( .B(n8551), .A(n8552), .Z(n8550) );
XOR U14252 ( .A(c2850), .B(b[2850]), .Z(n8551) );
XNOR U14253 ( .A(b[2850]), .B(n8552), .Z(c[2850]) );
XNOR U14254 ( .A(a[2850]), .B(c2850), .Z(n8552) );
XOR U14255 ( .A(c2851), .B(n8553), .Z(c2852) );
ANDN U14256 ( .B(n8554), .A(n8555), .Z(n8553) );
XOR U14257 ( .A(c2851), .B(b[2851]), .Z(n8554) );
XNOR U14258 ( .A(b[2851]), .B(n8555), .Z(c[2851]) );
XNOR U14259 ( .A(a[2851]), .B(c2851), .Z(n8555) );
XOR U14260 ( .A(c2852), .B(n8556), .Z(c2853) );
ANDN U14261 ( .B(n8557), .A(n8558), .Z(n8556) );
XOR U14262 ( .A(c2852), .B(b[2852]), .Z(n8557) );
XNOR U14263 ( .A(b[2852]), .B(n8558), .Z(c[2852]) );
XNOR U14264 ( .A(a[2852]), .B(c2852), .Z(n8558) );
XOR U14265 ( .A(c2853), .B(n8559), .Z(c2854) );
ANDN U14266 ( .B(n8560), .A(n8561), .Z(n8559) );
XOR U14267 ( .A(c2853), .B(b[2853]), .Z(n8560) );
XNOR U14268 ( .A(b[2853]), .B(n8561), .Z(c[2853]) );
XNOR U14269 ( .A(a[2853]), .B(c2853), .Z(n8561) );
XOR U14270 ( .A(c2854), .B(n8562), .Z(c2855) );
ANDN U14271 ( .B(n8563), .A(n8564), .Z(n8562) );
XOR U14272 ( .A(c2854), .B(b[2854]), .Z(n8563) );
XNOR U14273 ( .A(b[2854]), .B(n8564), .Z(c[2854]) );
XNOR U14274 ( .A(a[2854]), .B(c2854), .Z(n8564) );
XOR U14275 ( .A(c2855), .B(n8565), .Z(c2856) );
ANDN U14276 ( .B(n8566), .A(n8567), .Z(n8565) );
XOR U14277 ( .A(c2855), .B(b[2855]), .Z(n8566) );
XNOR U14278 ( .A(b[2855]), .B(n8567), .Z(c[2855]) );
XNOR U14279 ( .A(a[2855]), .B(c2855), .Z(n8567) );
XOR U14280 ( .A(c2856), .B(n8568), .Z(c2857) );
ANDN U14281 ( .B(n8569), .A(n8570), .Z(n8568) );
XOR U14282 ( .A(c2856), .B(b[2856]), .Z(n8569) );
XNOR U14283 ( .A(b[2856]), .B(n8570), .Z(c[2856]) );
XNOR U14284 ( .A(a[2856]), .B(c2856), .Z(n8570) );
XOR U14285 ( .A(c2857), .B(n8571), .Z(c2858) );
ANDN U14286 ( .B(n8572), .A(n8573), .Z(n8571) );
XOR U14287 ( .A(c2857), .B(b[2857]), .Z(n8572) );
XNOR U14288 ( .A(b[2857]), .B(n8573), .Z(c[2857]) );
XNOR U14289 ( .A(a[2857]), .B(c2857), .Z(n8573) );
XOR U14290 ( .A(c2858), .B(n8574), .Z(c2859) );
ANDN U14291 ( .B(n8575), .A(n8576), .Z(n8574) );
XOR U14292 ( .A(c2858), .B(b[2858]), .Z(n8575) );
XNOR U14293 ( .A(b[2858]), .B(n8576), .Z(c[2858]) );
XNOR U14294 ( .A(a[2858]), .B(c2858), .Z(n8576) );
XOR U14295 ( .A(c2859), .B(n8577), .Z(c2860) );
ANDN U14296 ( .B(n8578), .A(n8579), .Z(n8577) );
XOR U14297 ( .A(c2859), .B(b[2859]), .Z(n8578) );
XNOR U14298 ( .A(b[2859]), .B(n8579), .Z(c[2859]) );
XNOR U14299 ( .A(a[2859]), .B(c2859), .Z(n8579) );
XOR U14300 ( .A(c2860), .B(n8580), .Z(c2861) );
ANDN U14301 ( .B(n8581), .A(n8582), .Z(n8580) );
XOR U14302 ( .A(c2860), .B(b[2860]), .Z(n8581) );
XNOR U14303 ( .A(b[2860]), .B(n8582), .Z(c[2860]) );
XNOR U14304 ( .A(a[2860]), .B(c2860), .Z(n8582) );
XOR U14305 ( .A(c2861), .B(n8583), .Z(c2862) );
ANDN U14306 ( .B(n8584), .A(n8585), .Z(n8583) );
XOR U14307 ( .A(c2861), .B(b[2861]), .Z(n8584) );
XNOR U14308 ( .A(b[2861]), .B(n8585), .Z(c[2861]) );
XNOR U14309 ( .A(a[2861]), .B(c2861), .Z(n8585) );
XOR U14310 ( .A(c2862), .B(n8586), .Z(c2863) );
ANDN U14311 ( .B(n8587), .A(n8588), .Z(n8586) );
XOR U14312 ( .A(c2862), .B(b[2862]), .Z(n8587) );
XNOR U14313 ( .A(b[2862]), .B(n8588), .Z(c[2862]) );
XNOR U14314 ( .A(a[2862]), .B(c2862), .Z(n8588) );
XOR U14315 ( .A(c2863), .B(n8589), .Z(c2864) );
ANDN U14316 ( .B(n8590), .A(n8591), .Z(n8589) );
XOR U14317 ( .A(c2863), .B(b[2863]), .Z(n8590) );
XNOR U14318 ( .A(b[2863]), .B(n8591), .Z(c[2863]) );
XNOR U14319 ( .A(a[2863]), .B(c2863), .Z(n8591) );
XOR U14320 ( .A(c2864), .B(n8592), .Z(c2865) );
ANDN U14321 ( .B(n8593), .A(n8594), .Z(n8592) );
XOR U14322 ( .A(c2864), .B(b[2864]), .Z(n8593) );
XNOR U14323 ( .A(b[2864]), .B(n8594), .Z(c[2864]) );
XNOR U14324 ( .A(a[2864]), .B(c2864), .Z(n8594) );
XOR U14325 ( .A(c2865), .B(n8595), .Z(c2866) );
ANDN U14326 ( .B(n8596), .A(n8597), .Z(n8595) );
XOR U14327 ( .A(c2865), .B(b[2865]), .Z(n8596) );
XNOR U14328 ( .A(b[2865]), .B(n8597), .Z(c[2865]) );
XNOR U14329 ( .A(a[2865]), .B(c2865), .Z(n8597) );
XOR U14330 ( .A(c2866), .B(n8598), .Z(c2867) );
ANDN U14331 ( .B(n8599), .A(n8600), .Z(n8598) );
XOR U14332 ( .A(c2866), .B(b[2866]), .Z(n8599) );
XNOR U14333 ( .A(b[2866]), .B(n8600), .Z(c[2866]) );
XNOR U14334 ( .A(a[2866]), .B(c2866), .Z(n8600) );
XOR U14335 ( .A(c2867), .B(n8601), .Z(c2868) );
ANDN U14336 ( .B(n8602), .A(n8603), .Z(n8601) );
XOR U14337 ( .A(c2867), .B(b[2867]), .Z(n8602) );
XNOR U14338 ( .A(b[2867]), .B(n8603), .Z(c[2867]) );
XNOR U14339 ( .A(a[2867]), .B(c2867), .Z(n8603) );
XOR U14340 ( .A(c2868), .B(n8604), .Z(c2869) );
ANDN U14341 ( .B(n8605), .A(n8606), .Z(n8604) );
XOR U14342 ( .A(c2868), .B(b[2868]), .Z(n8605) );
XNOR U14343 ( .A(b[2868]), .B(n8606), .Z(c[2868]) );
XNOR U14344 ( .A(a[2868]), .B(c2868), .Z(n8606) );
XOR U14345 ( .A(c2869), .B(n8607), .Z(c2870) );
ANDN U14346 ( .B(n8608), .A(n8609), .Z(n8607) );
XOR U14347 ( .A(c2869), .B(b[2869]), .Z(n8608) );
XNOR U14348 ( .A(b[2869]), .B(n8609), .Z(c[2869]) );
XNOR U14349 ( .A(a[2869]), .B(c2869), .Z(n8609) );
XOR U14350 ( .A(c2870), .B(n8610), .Z(c2871) );
ANDN U14351 ( .B(n8611), .A(n8612), .Z(n8610) );
XOR U14352 ( .A(c2870), .B(b[2870]), .Z(n8611) );
XNOR U14353 ( .A(b[2870]), .B(n8612), .Z(c[2870]) );
XNOR U14354 ( .A(a[2870]), .B(c2870), .Z(n8612) );
XOR U14355 ( .A(c2871), .B(n8613), .Z(c2872) );
ANDN U14356 ( .B(n8614), .A(n8615), .Z(n8613) );
XOR U14357 ( .A(c2871), .B(b[2871]), .Z(n8614) );
XNOR U14358 ( .A(b[2871]), .B(n8615), .Z(c[2871]) );
XNOR U14359 ( .A(a[2871]), .B(c2871), .Z(n8615) );
XOR U14360 ( .A(c2872), .B(n8616), .Z(c2873) );
ANDN U14361 ( .B(n8617), .A(n8618), .Z(n8616) );
XOR U14362 ( .A(c2872), .B(b[2872]), .Z(n8617) );
XNOR U14363 ( .A(b[2872]), .B(n8618), .Z(c[2872]) );
XNOR U14364 ( .A(a[2872]), .B(c2872), .Z(n8618) );
XOR U14365 ( .A(c2873), .B(n8619), .Z(c2874) );
ANDN U14366 ( .B(n8620), .A(n8621), .Z(n8619) );
XOR U14367 ( .A(c2873), .B(b[2873]), .Z(n8620) );
XNOR U14368 ( .A(b[2873]), .B(n8621), .Z(c[2873]) );
XNOR U14369 ( .A(a[2873]), .B(c2873), .Z(n8621) );
XOR U14370 ( .A(c2874), .B(n8622), .Z(c2875) );
ANDN U14371 ( .B(n8623), .A(n8624), .Z(n8622) );
XOR U14372 ( .A(c2874), .B(b[2874]), .Z(n8623) );
XNOR U14373 ( .A(b[2874]), .B(n8624), .Z(c[2874]) );
XNOR U14374 ( .A(a[2874]), .B(c2874), .Z(n8624) );
XOR U14375 ( .A(c2875), .B(n8625), .Z(c2876) );
ANDN U14376 ( .B(n8626), .A(n8627), .Z(n8625) );
XOR U14377 ( .A(c2875), .B(b[2875]), .Z(n8626) );
XNOR U14378 ( .A(b[2875]), .B(n8627), .Z(c[2875]) );
XNOR U14379 ( .A(a[2875]), .B(c2875), .Z(n8627) );
XOR U14380 ( .A(c2876), .B(n8628), .Z(c2877) );
ANDN U14381 ( .B(n8629), .A(n8630), .Z(n8628) );
XOR U14382 ( .A(c2876), .B(b[2876]), .Z(n8629) );
XNOR U14383 ( .A(b[2876]), .B(n8630), .Z(c[2876]) );
XNOR U14384 ( .A(a[2876]), .B(c2876), .Z(n8630) );
XOR U14385 ( .A(c2877), .B(n8631), .Z(c2878) );
ANDN U14386 ( .B(n8632), .A(n8633), .Z(n8631) );
XOR U14387 ( .A(c2877), .B(b[2877]), .Z(n8632) );
XNOR U14388 ( .A(b[2877]), .B(n8633), .Z(c[2877]) );
XNOR U14389 ( .A(a[2877]), .B(c2877), .Z(n8633) );
XOR U14390 ( .A(c2878), .B(n8634), .Z(c2879) );
ANDN U14391 ( .B(n8635), .A(n8636), .Z(n8634) );
XOR U14392 ( .A(c2878), .B(b[2878]), .Z(n8635) );
XNOR U14393 ( .A(b[2878]), .B(n8636), .Z(c[2878]) );
XNOR U14394 ( .A(a[2878]), .B(c2878), .Z(n8636) );
XOR U14395 ( .A(c2879), .B(n8637), .Z(c2880) );
ANDN U14396 ( .B(n8638), .A(n8639), .Z(n8637) );
XOR U14397 ( .A(c2879), .B(b[2879]), .Z(n8638) );
XNOR U14398 ( .A(b[2879]), .B(n8639), .Z(c[2879]) );
XNOR U14399 ( .A(a[2879]), .B(c2879), .Z(n8639) );
XOR U14400 ( .A(c2880), .B(n8640), .Z(c2881) );
ANDN U14401 ( .B(n8641), .A(n8642), .Z(n8640) );
XOR U14402 ( .A(c2880), .B(b[2880]), .Z(n8641) );
XNOR U14403 ( .A(b[2880]), .B(n8642), .Z(c[2880]) );
XNOR U14404 ( .A(a[2880]), .B(c2880), .Z(n8642) );
XOR U14405 ( .A(c2881), .B(n8643), .Z(c2882) );
ANDN U14406 ( .B(n8644), .A(n8645), .Z(n8643) );
XOR U14407 ( .A(c2881), .B(b[2881]), .Z(n8644) );
XNOR U14408 ( .A(b[2881]), .B(n8645), .Z(c[2881]) );
XNOR U14409 ( .A(a[2881]), .B(c2881), .Z(n8645) );
XOR U14410 ( .A(c2882), .B(n8646), .Z(c2883) );
ANDN U14411 ( .B(n8647), .A(n8648), .Z(n8646) );
XOR U14412 ( .A(c2882), .B(b[2882]), .Z(n8647) );
XNOR U14413 ( .A(b[2882]), .B(n8648), .Z(c[2882]) );
XNOR U14414 ( .A(a[2882]), .B(c2882), .Z(n8648) );
XOR U14415 ( .A(c2883), .B(n8649), .Z(c2884) );
ANDN U14416 ( .B(n8650), .A(n8651), .Z(n8649) );
XOR U14417 ( .A(c2883), .B(b[2883]), .Z(n8650) );
XNOR U14418 ( .A(b[2883]), .B(n8651), .Z(c[2883]) );
XNOR U14419 ( .A(a[2883]), .B(c2883), .Z(n8651) );
XOR U14420 ( .A(c2884), .B(n8652), .Z(c2885) );
ANDN U14421 ( .B(n8653), .A(n8654), .Z(n8652) );
XOR U14422 ( .A(c2884), .B(b[2884]), .Z(n8653) );
XNOR U14423 ( .A(b[2884]), .B(n8654), .Z(c[2884]) );
XNOR U14424 ( .A(a[2884]), .B(c2884), .Z(n8654) );
XOR U14425 ( .A(c2885), .B(n8655), .Z(c2886) );
ANDN U14426 ( .B(n8656), .A(n8657), .Z(n8655) );
XOR U14427 ( .A(c2885), .B(b[2885]), .Z(n8656) );
XNOR U14428 ( .A(b[2885]), .B(n8657), .Z(c[2885]) );
XNOR U14429 ( .A(a[2885]), .B(c2885), .Z(n8657) );
XOR U14430 ( .A(c2886), .B(n8658), .Z(c2887) );
ANDN U14431 ( .B(n8659), .A(n8660), .Z(n8658) );
XOR U14432 ( .A(c2886), .B(b[2886]), .Z(n8659) );
XNOR U14433 ( .A(b[2886]), .B(n8660), .Z(c[2886]) );
XNOR U14434 ( .A(a[2886]), .B(c2886), .Z(n8660) );
XOR U14435 ( .A(c2887), .B(n8661), .Z(c2888) );
ANDN U14436 ( .B(n8662), .A(n8663), .Z(n8661) );
XOR U14437 ( .A(c2887), .B(b[2887]), .Z(n8662) );
XNOR U14438 ( .A(b[2887]), .B(n8663), .Z(c[2887]) );
XNOR U14439 ( .A(a[2887]), .B(c2887), .Z(n8663) );
XOR U14440 ( .A(c2888), .B(n8664), .Z(c2889) );
ANDN U14441 ( .B(n8665), .A(n8666), .Z(n8664) );
XOR U14442 ( .A(c2888), .B(b[2888]), .Z(n8665) );
XNOR U14443 ( .A(b[2888]), .B(n8666), .Z(c[2888]) );
XNOR U14444 ( .A(a[2888]), .B(c2888), .Z(n8666) );
XOR U14445 ( .A(c2889), .B(n8667), .Z(c2890) );
ANDN U14446 ( .B(n8668), .A(n8669), .Z(n8667) );
XOR U14447 ( .A(c2889), .B(b[2889]), .Z(n8668) );
XNOR U14448 ( .A(b[2889]), .B(n8669), .Z(c[2889]) );
XNOR U14449 ( .A(a[2889]), .B(c2889), .Z(n8669) );
XOR U14450 ( .A(c2890), .B(n8670), .Z(c2891) );
ANDN U14451 ( .B(n8671), .A(n8672), .Z(n8670) );
XOR U14452 ( .A(c2890), .B(b[2890]), .Z(n8671) );
XNOR U14453 ( .A(b[2890]), .B(n8672), .Z(c[2890]) );
XNOR U14454 ( .A(a[2890]), .B(c2890), .Z(n8672) );
XOR U14455 ( .A(c2891), .B(n8673), .Z(c2892) );
ANDN U14456 ( .B(n8674), .A(n8675), .Z(n8673) );
XOR U14457 ( .A(c2891), .B(b[2891]), .Z(n8674) );
XNOR U14458 ( .A(b[2891]), .B(n8675), .Z(c[2891]) );
XNOR U14459 ( .A(a[2891]), .B(c2891), .Z(n8675) );
XOR U14460 ( .A(c2892), .B(n8676), .Z(c2893) );
ANDN U14461 ( .B(n8677), .A(n8678), .Z(n8676) );
XOR U14462 ( .A(c2892), .B(b[2892]), .Z(n8677) );
XNOR U14463 ( .A(b[2892]), .B(n8678), .Z(c[2892]) );
XNOR U14464 ( .A(a[2892]), .B(c2892), .Z(n8678) );
XOR U14465 ( .A(c2893), .B(n8679), .Z(c2894) );
ANDN U14466 ( .B(n8680), .A(n8681), .Z(n8679) );
XOR U14467 ( .A(c2893), .B(b[2893]), .Z(n8680) );
XNOR U14468 ( .A(b[2893]), .B(n8681), .Z(c[2893]) );
XNOR U14469 ( .A(a[2893]), .B(c2893), .Z(n8681) );
XOR U14470 ( .A(c2894), .B(n8682), .Z(c2895) );
ANDN U14471 ( .B(n8683), .A(n8684), .Z(n8682) );
XOR U14472 ( .A(c2894), .B(b[2894]), .Z(n8683) );
XNOR U14473 ( .A(b[2894]), .B(n8684), .Z(c[2894]) );
XNOR U14474 ( .A(a[2894]), .B(c2894), .Z(n8684) );
XOR U14475 ( .A(c2895), .B(n8685), .Z(c2896) );
ANDN U14476 ( .B(n8686), .A(n8687), .Z(n8685) );
XOR U14477 ( .A(c2895), .B(b[2895]), .Z(n8686) );
XNOR U14478 ( .A(b[2895]), .B(n8687), .Z(c[2895]) );
XNOR U14479 ( .A(a[2895]), .B(c2895), .Z(n8687) );
XOR U14480 ( .A(c2896), .B(n8688), .Z(c2897) );
ANDN U14481 ( .B(n8689), .A(n8690), .Z(n8688) );
XOR U14482 ( .A(c2896), .B(b[2896]), .Z(n8689) );
XNOR U14483 ( .A(b[2896]), .B(n8690), .Z(c[2896]) );
XNOR U14484 ( .A(a[2896]), .B(c2896), .Z(n8690) );
XOR U14485 ( .A(c2897), .B(n8691), .Z(c2898) );
ANDN U14486 ( .B(n8692), .A(n8693), .Z(n8691) );
XOR U14487 ( .A(c2897), .B(b[2897]), .Z(n8692) );
XNOR U14488 ( .A(b[2897]), .B(n8693), .Z(c[2897]) );
XNOR U14489 ( .A(a[2897]), .B(c2897), .Z(n8693) );
XOR U14490 ( .A(c2898), .B(n8694), .Z(c2899) );
ANDN U14491 ( .B(n8695), .A(n8696), .Z(n8694) );
XOR U14492 ( .A(c2898), .B(b[2898]), .Z(n8695) );
XNOR U14493 ( .A(b[2898]), .B(n8696), .Z(c[2898]) );
XNOR U14494 ( .A(a[2898]), .B(c2898), .Z(n8696) );
XOR U14495 ( .A(c2899), .B(n8697), .Z(c2900) );
ANDN U14496 ( .B(n8698), .A(n8699), .Z(n8697) );
XOR U14497 ( .A(c2899), .B(b[2899]), .Z(n8698) );
XNOR U14498 ( .A(b[2899]), .B(n8699), .Z(c[2899]) );
XNOR U14499 ( .A(a[2899]), .B(c2899), .Z(n8699) );
XOR U14500 ( .A(c2900), .B(n8700), .Z(c2901) );
ANDN U14501 ( .B(n8701), .A(n8702), .Z(n8700) );
XOR U14502 ( .A(c2900), .B(b[2900]), .Z(n8701) );
XNOR U14503 ( .A(b[2900]), .B(n8702), .Z(c[2900]) );
XNOR U14504 ( .A(a[2900]), .B(c2900), .Z(n8702) );
XOR U14505 ( .A(c2901), .B(n8703), .Z(c2902) );
ANDN U14506 ( .B(n8704), .A(n8705), .Z(n8703) );
XOR U14507 ( .A(c2901), .B(b[2901]), .Z(n8704) );
XNOR U14508 ( .A(b[2901]), .B(n8705), .Z(c[2901]) );
XNOR U14509 ( .A(a[2901]), .B(c2901), .Z(n8705) );
XOR U14510 ( .A(c2902), .B(n8706), .Z(c2903) );
ANDN U14511 ( .B(n8707), .A(n8708), .Z(n8706) );
XOR U14512 ( .A(c2902), .B(b[2902]), .Z(n8707) );
XNOR U14513 ( .A(b[2902]), .B(n8708), .Z(c[2902]) );
XNOR U14514 ( .A(a[2902]), .B(c2902), .Z(n8708) );
XOR U14515 ( .A(c2903), .B(n8709), .Z(c2904) );
ANDN U14516 ( .B(n8710), .A(n8711), .Z(n8709) );
XOR U14517 ( .A(c2903), .B(b[2903]), .Z(n8710) );
XNOR U14518 ( .A(b[2903]), .B(n8711), .Z(c[2903]) );
XNOR U14519 ( .A(a[2903]), .B(c2903), .Z(n8711) );
XOR U14520 ( .A(c2904), .B(n8712), .Z(c2905) );
ANDN U14521 ( .B(n8713), .A(n8714), .Z(n8712) );
XOR U14522 ( .A(c2904), .B(b[2904]), .Z(n8713) );
XNOR U14523 ( .A(b[2904]), .B(n8714), .Z(c[2904]) );
XNOR U14524 ( .A(a[2904]), .B(c2904), .Z(n8714) );
XOR U14525 ( .A(c2905), .B(n8715), .Z(c2906) );
ANDN U14526 ( .B(n8716), .A(n8717), .Z(n8715) );
XOR U14527 ( .A(c2905), .B(b[2905]), .Z(n8716) );
XNOR U14528 ( .A(b[2905]), .B(n8717), .Z(c[2905]) );
XNOR U14529 ( .A(a[2905]), .B(c2905), .Z(n8717) );
XOR U14530 ( .A(c2906), .B(n8718), .Z(c2907) );
ANDN U14531 ( .B(n8719), .A(n8720), .Z(n8718) );
XOR U14532 ( .A(c2906), .B(b[2906]), .Z(n8719) );
XNOR U14533 ( .A(b[2906]), .B(n8720), .Z(c[2906]) );
XNOR U14534 ( .A(a[2906]), .B(c2906), .Z(n8720) );
XOR U14535 ( .A(c2907), .B(n8721), .Z(c2908) );
ANDN U14536 ( .B(n8722), .A(n8723), .Z(n8721) );
XOR U14537 ( .A(c2907), .B(b[2907]), .Z(n8722) );
XNOR U14538 ( .A(b[2907]), .B(n8723), .Z(c[2907]) );
XNOR U14539 ( .A(a[2907]), .B(c2907), .Z(n8723) );
XOR U14540 ( .A(c2908), .B(n8724), .Z(c2909) );
ANDN U14541 ( .B(n8725), .A(n8726), .Z(n8724) );
XOR U14542 ( .A(c2908), .B(b[2908]), .Z(n8725) );
XNOR U14543 ( .A(b[2908]), .B(n8726), .Z(c[2908]) );
XNOR U14544 ( .A(a[2908]), .B(c2908), .Z(n8726) );
XOR U14545 ( .A(c2909), .B(n8727), .Z(c2910) );
ANDN U14546 ( .B(n8728), .A(n8729), .Z(n8727) );
XOR U14547 ( .A(c2909), .B(b[2909]), .Z(n8728) );
XNOR U14548 ( .A(b[2909]), .B(n8729), .Z(c[2909]) );
XNOR U14549 ( .A(a[2909]), .B(c2909), .Z(n8729) );
XOR U14550 ( .A(c2910), .B(n8730), .Z(c2911) );
ANDN U14551 ( .B(n8731), .A(n8732), .Z(n8730) );
XOR U14552 ( .A(c2910), .B(b[2910]), .Z(n8731) );
XNOR U14553 ( .A(b[2910]), .B(n8732), .Z(c[2910]) );
XNOR U14554 ( .A(a[2910]), .B(c2910), .Z(n8732) );
XOR U14555 ( .A(c2911), .B(n8733), .Z(c2912) );
ANDN U14556 ( .B(n8734), .A(n8735), .Z(n8733) );
XOR U14557 ( .A(c2911), .B(b[2911]), .Z(n8734) );
XNOR U14558 ( .A(b[2911]), .B(n8735), .Z(c[2911]) );
XNOR U14559 ( .A(a[2911]), .B(c2911), .Z(n8735) );
XOR U14560 ( .A(c2912), .B(n8736), .Z(c2913) );
ANDN U14561 ( .B(n8737), .A(n8738), .Z(n8736) );
XOR U14562 ( .A(c2912), .B(b[2912]), .Z(n8737) );
XNOR U14563 ( .A(b[2912]), .B(n8738), .Z(c[2912]) );
XNOR U14564 ( .A(a[2912]), .B(c2912), .Z(n8738) );
XOR U14565 ( .A(c2913), .B(n8739), .Z(c2914) );
ANDN U14566 ( .B(n8740), .A(n8741), .Z(n8739) );
XOR U14567 ( .A(c2913), .B(b[2913]), .Z(n8740) );
XNOR U14568 ( .A(b[2913]), .B(n8741), .Z(c[2913]) );
XNOR U14569 ( .A(a[2913]), .B(c2913), .Z(n8741) );
XOR U14570 ( .A(c2914), .B(n8742), .Z(c2915) );
ANDN U14571 ( .B(n8743), .A(n8744), .Z(n8742) );
XOR U14572 ( .A(c2914), .B(b[2914]), .Z(n8743) );
XNOR U14573 ( .A(b[2914]), .B(n8744), .Z(c[2914]) );
XNOR U14574 ( .A(a[2914]), .B(c2914), .Z(n8744) );
XOR U14575 ( .A(c2915), .B(n8745), .Z(c2916) );
ANDN U14576 ( .B(n8746), .A(n8747), .Z(n8745) );
XOR U14577 ( .A(c2915), .B(b[2915]), .Z(n8746) );
XNOR U14578 ( .A(b[2915]), .B(n8747), .Z(c[2915]) );
XNOR U14579 ( .A(a[2915]), .B(c2915), .Z(n8747) );
XOR U14580 ( .A(c2916), .B(n8748), .Z(c2917) );
ANDN U14581 ( .B(n8749), .A(n8750), .Z(n8748) );
XOR U14582 ( .A(c2916), .B(b[2916]), .Z(n8749) );
XNOR U14583 ( .A(b[2916]), .B(n8750), .Z(c[2916]) );
XNOR U14584 ( .A(a[2916]), .B(c2916), .Z(n8750) );
XOR U14585 ( .A(c2917), .B(n8751), .Z(c2918) );
ANDN U14586 ( .B(n8752), .A(n8753), .Z(n8751) );
XOR U14587 ( .A(c2917), .B(b[2917]), .Z(n8752) );
XNOR U14588 ( .A(b[2917]), .B(n8753), .Z(c[2917]) );
XNOR U14589 ( .A(a[2917]), .B(c2917), .Z(n8753) );
XOR U14590 ( .A(c2918), .B(n8754), .Z(c2919) );
ANDN U14591 ( .B(n8755), .A(n8756), .Z(n8754) );
XOR U14592 ( .A(c2918), .B(b[2918]), .Z(n8755) );
XNOR U14593 ( .A(b[2918]), .B(n8756), .Z(c[2918]) );
XNOR U14594 ( .A(a[2918]), .B(c2918), .Z(n8756) );
XOR U14595 ( .A(c2919), .B(n8757), .Z(c2920) );
ANDN U14596 ( .B(n8758), .A(n8759), .Z(n8757) );
XOR U14597 ( .A(c2919), .B(b[2919]), .Z(n8758) );
XNOR U14598 ( .A(b[2919]), .B(n8759), .Z(c[2919]) );
XNOR U14599 ( .A(a[2919]), .B(c2919), .Z(n8759) );
XOR U14600 ( .A(c2920), .B(n8760), .Z(c2921) );
ANDN U14601 ( .B(n8761), .A(n8762), .Z(n8760) );
XOR U14602 ( .A(c2920), .B(b[2920]), .Z(n8761) );
XNOR U14603 ( .A(b[2920]), .B(n8762), .Z(c[2920]) );
XNOR U14604 ( .A(a[2920]), .B(c2920), .Z(n8762) );
XOR U14605 ( .A(c2921), .B(n8763), .Z(c2922) );
ANDN U14606 ( .B(n8764), .A(n8765), .Z(n8763) );
XOR U14607 ( .A(c2921), .B(b[2921]), .Z(n8764) );
XNOR U14608 ( .A(b[2921]), .B(n8765), .Z(c[2921]) );
XNOR U14609 ( .A(a[2921]), .B(c2921), .Z(n8765) );
XOR U14610 ( .A(c2922), .B(n8766), .Z(c2923) );
ANDN U14611 ( .B(n8767), .A(n8768), .Z(n8766) );
XOR U14612 ( .A(c2922), .B(b[2922]), .Z(n8767) );
XNOR U14613 ( .A(b[2922]), .B(n8768), .Z(c[2922]) );
XNOR U14614 ( .A(a[2922]), .B(c2922), .Z(n8768) );
XOR U14615 ( .A(c2923), .B(n8769), .Z(c2924) );
ANDN U14616 ( .B(n8770), .A(n8771), .Z(n8769) );
XOR U14617 ( .A(c2923), .B(b[2923]), .Z(n8770) );
XNOR U14618 ( .A(b[2923]), .B(n8771), .Z(c[2923]) );
XNOR U14619 ( .A(a[2923]), .B(c2923), .Z(n8771) );
XOR U14620 ( .A(c2924), .B(n8772), .Z(c2925) );
ANDN U14621 ( .B(n8773), .A(n8774), .Z(n8772) );
XOR U14622 ( .A(c2924), .B(b[2924]), .Z(n8773) );
XNOR U14623 ( .A(b[2924]), .B(n8774), .Z(c[2924]) );
XNOR U14624 ( .A(a[2924]), .B(c2924), .Z(n8774) );
XOR U14625 ( .A(c2925), .B(n8775), .Z(c2926) );
ANDN U14626 ( .B(n8776), .A(n8777), .Z(n8775) );
XOR U14627 ( .A(c2925), .B(b[2925]), .Z(n8776) );
XNOR U14628 ( .A(b[2925]), .B(n8777), .Z(c[2925]) );
XNOR U14629 ( .A(a[2925]), .B(c2925), .Z(n8777) );
XOR U14630 ( .A(c2926), .B(n8778), .Z(c2927) );
ANDN U14631 ( .B(n8779), .A(n8780), .Z(n8778) );
XOR U14632 ( .A(c2926), .B(b[2926]), .Z(n8779) );
XNOR U14633 ( .A(b[2926]), .B(n8780), .Z(c[2926]) );
XNOR U14634 ( .A(a[2926]), .B(c2926), .Z(n8780) );
XOR U14635 ( .A(c2927), .B(n8781), .Z(c2928) );
ANDN U14636 ( .B(n8782), .A(n8783), .Z(n8781) );
XOR U14637 ( .A(c2927), .B(b[2927]), .Z(n8782) );
XNOR U14638 ( .A(b[2927]), .B(n8783), .Z(c[2927]) );
XNOR U14639 ( .A(a[2927]), .B(c2927), .Z(n8783) );
XOR U14640 ( .A(c2928), .B(n8784), .Z(c2929) );
ANDN U14641 ( .B(n8785), .A(n8786), .Z(n8784) );
XOR U14642 ( .A(c2928), .B(b[2928]), .Z(n8785) );
XNOR U14643 ( .A(b[2928]), .B(n8786), .Z(c[2928]) );
XNOR U14644 ( .A(a[2928]), .B(c2928), .Z(n8786) );
XOR U14645 ( .A(c2929), .B(n8787), .Z(c2930) );
ANDN U14646 ( .B(n8788), .A(n8789), .Z(n8787) );
XOR U14647 ( .A(c2929), .B(b[2929]), .Z(n8788) );
XNOR U14648 ( .A(b[2929]), .B(n8789), .Z(c[2929]) );
XNOR U14649 ( .A(a[2929]), .B(c2929), .Z(n8789) );
XOR U14650 ( .A(c2930), .B(n8790), .Z(c2931) );
ANDN U14651 ( .B(n8791), .A(n8792), .Z(n8790) );
XOR U14652 ( .A(c2930), .B(b[2930]), .Z(n8791) );
XNOR U14653 ( .A(b[2930]), .B(n8792), .Z(c[2930]) );
XNOR U14654 ( .A(a[2930]), .B(c2930), .Z(n8792) );
XOR U14655 ( .A(c2931), .B(n8793), .Z(c2932) );
ANDN U14656 ( .B(n8794), .A(n8795), .Z(n8793) );
XOR U14657 ( .A(c2931), .B(b[2931]), .Z(n8794) );
XNOR U14658 ( .A(b[2931]), .B(n8795), .Z(c[2931]) );
XNOR U14659 ( .A(a[2931]), .B(c2931), .Z(n8795) );
XOR U14660 ( .A(c2932), .B(n8796), .Z(c2933) );
ANDN U14661 ( .B(n8797), .A(n8798), .Z(n8796) );
XOR U14662 ( .A(c2932), .B(b[2932]), .Z(n8797) );
XNOR U14663 ( .A(b[2932]), .B(n8798), .Z(c[2932]) );
XNOR U14664 ( .A(a[2932]), .B(c2932), .Z(n8798) );
XOR U14665 ( .A(c2933), .B(n8799), .Z(c2934) );
ANDN U14666 ( .B(n8800), .A(n8801), .Z(n8799) );
XOR U14667 ( .A(c2933), .B(b[2933]), .Z(n8800) );
XNOR U14668 ( .A(b[2933]), .B(n8801), .Z(c[2933]) );
XNOR U14669 ( .A(a[2933]), .B(c2933), .Z(n8801) );
XOR U14670 ( .A(c2934), .B(n8802), .Z(c2935) );
ANDN U14671 ( .B(n8803), .A(n8804), .Z(n8802) );
XOR U14672 ( .A(c2934), .B(b[2934]), .Z(n8803) );
XNOR U14673 ( .A(b[2934]), .B(n8804), .Z(c[2934]) );
XNOR U14674 ( .A(a[2934]), .B(c2934), .Z(n8804) );
XOR U14675 ( .A(c2935), .B(n8805), .Z(c2936) );
ANDN U14676 ( .B(n8806), .A(n8807), .Z(n8805) );
XOR U14677 ( .A(c2935), .B(b[2935]), .Z(n8806) );
XNOR U14678 ( .A(b[2935]), .B(n8807), .Z(c[2935]) );
XNOR U14679 ( .A(a[2935]), .B(c2935), .Z(n8807) );
XOR U14680 ( .A(c2936), .B(n8808), .Z(c2937) );
ANDN U14681 ( .B(n8809), .A(n8810), .Z(n8808) );
XOR U14682 ( .A(c2936), .B(b[2936]), .Z(n8809) );
XNOR U14683 ( .A(b[2936]), .B(n8810), .Z(c[2936]) );
XNOR U14684 ( .A(a[2936]), .B(c2936), .Z(n8810) );
XOR U14685 ( .A(c2937), .B(n8811), .Z(c2938) );
ANDN U14686 ( .B(n8812), .A(n8813), .Z(n8811) );
XOR U14687 ( .A(c2937), .B(b[2937]), .Z(n8812) );
XNOR U14688 ( .A(b[2937]), .B(n8813), .Z(c[2937]) );
XNOR U14689 ( .A(a[2937]), .B(c2937), .Z(n8813) );
XOR U14690 ( .A(c2938), .B(n8814), .Z(c2939) );
ANDN U14691 ( .B(n8815), .A(n8816), .Z(n8814) );
XOR U14692 ( .A(c2938), .B(b[2938]), .Z(n8815) );
XNOR U14693 ( .A(b[2938]), .B(n8816), .Z(c[2938]) );
XNOR U14694 ( .A(a[2938]), .B(c2938), .Z(n8816) );
XOR U14695 ( .A(c2939), .B(n8817), .Z(c2940) );
ANDN U14696 ( .B(n8818), .A(n8819), .Z(n8817) );
XOR U14697 ( .A(c2939), .B(b[2939]), .Z(n8818) );
XNOR U14698 ( .A(b[2939]), .B(n8819), .Z(c[2939]) );
XNOR U14699 ( .A(a[2939]), .B(c2939), .Z(n8819) );
XOR U14700 ( .A(c2940), .B(n8820), .Z(c2941) );
ANDN U14701 ( .B(n8821), .A(n8822), .Z(n8820) );
XOR U14702 ( .A(c2940), .B(b[2940]), .Z(n8821) );
XNOR U14703 ( .A(b[2940]), .B(n8822), .Z(c[2940]) );
XNOR U14704 ( .A(a[2940]), .B(c2940), .Z(n8822) );
XOR U14705 ( .A(c2941), .B(n8823), .Z(c2942) );
ANDN U14706 ( .B(n8824), .A(n8825), .Z(n8823) );
XOR U14707 ( .A(c2941), .B(b[2941]), .Z(n8824) );
XNOR U14708 ( .A(b[2941]), .B(n8825), .Z(c[2941]) );
XNOR U14709 ( .A(a[2941]), .B(c2941), .Z(n8825) );
XOR U14710 ( .A(c2942), .B(n8826), .Z(c2943) );
ANDN U14711 ( .B(n8827), .A(n8828), .Z(n8826) );
XOR U14712 ( .A(c2942), .B(b[2942]), .Z(n8827) );
XNOR U14713 ( .A(b[2942]), .B(n8828), .Z(c[2942]) );
XNOR U14714 ( .A(a[2942]), .B(c2942), .Z(n8828) );
XOR U14715 ( .A(c2943), .B(n8829), .Z(c2944) );
ANDN U14716 ( .B(n8830), .A(n8831), .Z(n8829) );
XOR U14717 ( .A(c2943), .B(b[2943]), .Z(n8830) );
XNOR U14718 ( .A(b[2943]), .B(n8831), .Z(c[2943]) );
XNOR U14719 ( .A(a[2943]), .B(c2943), .Z(n8831) );
XOR U14720 ( .A(c2944), .B(n8832), .Z(c2945) );
ANDN U14721 ( .B(n8833), .A(n8834), .Z(n8832) );
XOR U14722 ( .A(c2944), .B(b[2944]), .Z(n8833) );
XNOR U14723 ( .A(b[2944]), .B(n8834), .Z(c[2944]) );
XNOR U14724 ( .A(a[2944]), .B(c2944), .Z(n8834) );
XOR U14725 ( .A(c2945), .B(n8835), .Z(c2946) );
ANDN U14726 ( .B(n8836), .A(n8837), .Z(n8835) );
XOR U14727 ( .A(c2945), .B(b[2945]), .Z(n8836) );
XNOR U14728 ( .A(b[2945]), .B(n8837), .Z(c[2945]) );
XNOR U14729 ( .A(a[2945]), .B(c2945), .Z(n8837) );
XOR U14730 ( .A(c2946), .B(n8838), .Z(c2947) );
ANDN U14731 ( .B(n8839), .A(n8840), .Z(n8838) );
XOR U14732 ( .A(c2946), .B(b[2946]), .Z(n8839) );
XNOR U14733 ( .A(b[2946]), .B(n8840), .Z(c[2946]) );
XNOR U14734 ( .A(a[2946]), .B(c2946), .Z(n8840) );
XOR U14735 ( .A(c2947), .B(n8841), .Z(c2948) );
ANDN U14736 ( .B(n8842), .A(n8843), .Z(n8841) );
XOR U14737 ( .A(c2947), .B(b[2947]), .Z(n8842) );
XNOR U14738 ( .A(b[2947]), .B(n8843), .Z(c[2947]) );
XNOR U14739 ( .A(a[2947]), .B(c2947), .Z(n8843) );
XOR U14740 ( .A(c2948), .B(n8844), .Z(c2949) );
ANDN U14741 ( .B(n8845), .A(n8846), .Z(n8844) );
XOR U14742 ( .A(c2948), .B(b[2948]), .Z(n8845) );
XNOR U14743 ( .A(b[2948]), .B(n8846), .Z(c[2948]) );
XNOR U14744 ( .A(a[2948]), .B(c2948), .Z(n8846) );
XOR U14745 ( .A(c2949), .B(n8847), .Z(c2950) );
ANDN U14746 ( .B(n8848), .A(n8849), .Z(n8847) );
XOR U14747 ( .A(c2949), .B(b[2949]), .Z(n8848) );
XNOR U14748 ( .A(b[2949]), .B(n8849), .Z(c[2949]) );
XNOR U14749 ( .A(a[2949]), .B(c2949), .Z(n8849) );
XOR U14750 ( .A(c2950), .B(n8850), .Z(c2951) );
ANDN U14751 ( .B(n8851), .A(n8852), .Z(n8850) );
XOR U14752 ( .A(c2950), .B(b[2950]), .Z(n8851) );
XNOR U14753 ( .A(b[2950]), .B(n8852), .Z(c[2950]) );
XNOR U14754 ( .A(a[2950]), .B(c2950), .Z(n8852) );
XOR U14755 ( .A(c2951), .B(n8853), .Z(c2952) );
ANDN U14756 ( .B(n8854), .A(n8855), .Z(n8853) );
XOR U14757 ( .A(c2951), .B(b[2951]), .Z(n8854) );
XNOR U14758 ( .A(b[2951]), .B(n8855), .Z(c[2951]) );
XNOR U14759 ( .A(a[2951]), .B(c2951), .Z(n8855) );
XOR U14760 ( .A(c2952), .B(n8856), .Z(c2953) );
ANDN U14761 ( .B(n8857), .A(n8858), .Z(n8856) );
XOR U14762 ( .A(c2952), .B(b[2952]), .Z(n8857) );
XNOR U14763 ( .A(b[2952]), .B(n8858), .Z(c[2952]) );
XNOR U14764 ( .A(a[2952]), .B(c2952), .Z(n8858) );
XOR U14765 ( .A(c2953), .B(n8859), .Z(c2954) );
ANDN U14766 ( .B(n8860), .A(n8861), .Z(n8859) );
XOR U14767 ( .A(c2953), .B(b[2953]), .Z(n8860) );
XNOR U14768 ( .A(b[2953]), .B(n8861), .Z(c[2953]) );
XNOR U14769 ( .A(a[2953]), .B(c2953), .Z(n8861) );
XOR U14770 ( .A(c2954), .B(n8862), .Z(c2955) );
ANDN U14771 ( .B(n8863), .A(n8864), .Z(n8862) );
XOR U14772 ( .A(c2954), .B(b[2954]), .Z(n8863) );
XNOR U14773 ( .A(b[2954]), .B(n8864), .Z(c[2954]) );
XNOR U14774 ( .A(a[2954]), .B(c2954), .Z(n8864) );
XOR U14775 ( .A(c2955), .B(n8865), .Z(c2956) );
ANDN U14776 ( .B(n8866), .A(n8867), .Z(n8865) );
XOR U14777 ( .A(c2955), .B(b[2955]), .Z(n8866) );
XNOR U14778 ( .A(b[2955]), .B(n8867), .Z(c[2955]) );
XNOR U14779 ( .A(a[2955]), .B(c2955), .Z(n8867) );
XOR U14780 ( .A(c2956), .B(n8868), .Z(c2957) );
ANDN U14781 ( .B(n8869), .A(n8870), .Z(n8868) );
XOR U14782 ( .A(c2956), .B(b[2956]), .Z(n8869) );
XNOR U14783 ( .A(b[2956]), .B(n8870), .Z(c[2956]) );
XNOR U14784 ( .A(a[2956]), .B(c2956), .Z(n8870) );
XOR U14785 ( .A(c2957), .B(n8871), .Z(c2958) );
ANDN U14786 ( .B(n8872), .A(n8873), .Z(n8871) );
XOR U14787 ( .A(c2957), .B(b[2957]), .Z(n8872) );
XNOR U14788 ( .A(b[2957]), .B(n8873), .Z(c[2957]) );
XNOR U14789 ( .A(a[2957]), .B(c2957), .Z(n8873) );
XOR U14790 ( .A(c2958), .B(n8874), .Z(c2959) );
ANDN U14791 ( .B(n8875), .A(n8876), .Z(n8874) );
XOR U14792 ( .A(c2958), .B(b[2958]), .Z(n8875) );
XNOR U14793 ( .A(b[2958]), .B(n8876), .Z(c[2958]) );
XNOR U14794 ( .A(a[2958]), .B(c2958), .Z(n8876) );
XOR U14795 ( .A(c2959), .B(n8877), .Z(c2960) );
ANDN U14796 ( .B(n8878), .A(n8879), .Z(n8877) );
XOR U14797 ( .A(c2959), .B(b[2959]), .Z(n8878) );
XNOR U14798 ( .A(b[2959]), .B(n8879), .Z(c[2959]) );
XNOR U14799 ( .A(a[2959]), .B(c2959), .Z(n8879) );
XOR U14800 ( .A(c2960), .B(n8880), .Z(c2961) );
ANDN U14801 ( .B(n8881), .A(n8882), .Z(n8880) );
XOR U14802 ( .A(c2960), .B(b[2960]), .Z(n8881) );
XNOR U14803 ( .A(b[2960]), .B(n8882), .Z(c[2960]) );
XNOR U14804 ( .A(a[2960]), .B(c2960), .Z(n8882) );
XOR U14805 ( .A(c2961), .B(n8883), .Z(c2962) );
ANDN U14806 ( .B(n8884), .A(n8885), .Z(n8883) );
XOR U14807 ( .A(c2961), .B(b[2961]), .Z(n8884) );
XNOR U14808 ( .A(b[2961]), .B(n8885), .Z(c[2961]) );
XNOR U14809 ( .A(a[2961]), .B(c2961), .Z(n8885) );
XOR U14810 ( .A(c2962), .B(n8886), .Z(c2963) );
ANDN U14811 ( .B(n8887), .A(n8888), .Z(n8886) );
XOR U14812 ( .A(c2962), .B(b[2962]), .Z(n8887) );
XNOR U14813 ( .A(b[2962]), .B(n8888), .Z(c[2962]) );
XNOR U14814 ( .A(a[2962]), .B(c2962), .Z(n8888) );
XOR U14815 ( .A(c2963), .B(n8889), .Z(c2964) );
ANDN U14816 ( .B(n8890), .A(n8891), .Z(n8889) );
XOR U14817 ( .A(c2963), .B(b[2963]), .Z(n8890) );
XNOR U14818 ( .A(b[2963]), .B(n8891), .Z(c[2963]) );
XNOR U14819 ( .A(a[2963]), .B(c2963), .Z(n8891) );
XOR U14820 ( .A(c2964), .B(n8892), .Z(c2965) );
ANDN U14821 ( .B(n8893), .A(n8894), .Z(n8892) );
XOR U14822 ( .A(c2964), .B(b[2964]), .Z(n8893) );
XNOR U14823 ( .A(b[2964]), .B(n8894), .Z(c[2964]) );
XNOR U14824 ( .A(a[2964]), .B(c2964), .Z(n8894) );
XOR U14825 ( .A(c2965), .B(n8895), .Z(c2966) );
ANDN U14826 ( .B(n8896), .A(n8897), .Z(n8895) );
XOR U14827 ( .A(c2965), .B(b[2965]), .Z(n8896) );
XNOR U14828 ( .A(b[2965]), .B(n8897), .Z(c[2965]) );
XNOR U14829 ( .A(a[2965]), .B(c2965), .Z(n8897) );
XOR U14830 ( .A(c2966), .B(n8898), .Z(c2967) );
ANDN U14831 ( .B(n8899), .A(n8900), .Z(n8898) );
XOR U14832 ( .A(c2966), .B(b[2966]), .Z(n8899) );
XNOR U14833 ( .A(b[2966]), .B(n8900), .Z(c[2966]) );
XNOR U14834 ( .A(a[2966]), .B(c2966), .Z(n8900) );
XOR U14835 ( .A(c2967), .B(n8901), .Z(c2968) );
ANDN U14836 ( .B(n8902), .A(n8903), .Z(n8901) );
XOR U14837 ( .A(c2967), .B(b[2967]), .Z(n8902) );
XNOR U14838 ( .A(b[2967]), .B(n8903), .Z(c[2967]) );
XNOR U14839 ( .A(a[2967]), .B(c2967), .Z(n8903) );
XOR U14840 ( .A(c2968), .B(n8904), .Z(c2969) );
ANDN U14841 ( .B(n8905), .A(n8906), .Z(n8904) );
XOR U14842 ( .A(c2968), .B(b[2968]), .Z(n8905) );
XNOR U14843 ( .A(b[2968]), .B(n8906), .Z(c[2968]) );
XNOR U14844 ( .A(a[2968]), .B(c2968), .Z(n8906) );
XOR U14845 ( .A(c2969), .B(n8907), .Z(c2970) );
ANDN U14846 ( .B(n8908), .A(n8909), .Z(n8907) );
XOR U14847 ( .A(c2969), .B(b[2969]), .Z(n8908) );
XNOR U14848 ( .A(b[2969]), .B(n8909), .Z(c[2969]) );
XNOR U14849 ( .A(a[2969]), .B(c2969), .Z(n8909) );
XOR U14850 ( .A(c2970), .B(n8910), .Z(c2971) );
ANDN U14851 ( .B(n8911), .A(n8912), .Z(n8910) );
XOR U14852 ( .A(c2970), .B(b[2970]), .Z(n8911) );
XNOR U14853 ( .A(b[2970]), .B(n8912), .Z(c[2970]) );
XNOR U14854 ( .A(a[2970]), .B(c2970), .Z(n8912) );
XOR U14855 ( .A(c2971), .B(n8913), .Z(c2972) );
ANDN U14856 ( .B(n8914), .A(n8915), .Z(n8913) );
XOR U14857 ( .A(c2971), .B(b[2971]), .Z(n8914) );
XNOR U14858 ( .A(b[2971]), .B(n8915), .Z(c[2971]) );
XNOR U14859 ( .A(a[2971]), .B(c2971), .Z(n8915) );
XOR U14860 ( .A(c2972), .B(n8916), .Z(c2973) );
ANDN U14861 ( .B(n8917), .A(n8918), .Z(n8916) );
XOR U14862 ( .A(c2972), .B(b[2972]), .Z(n8917) );
XNOR U14863 ( .A(b[2972]), .B(n8918), .Z(c[2972]) );
XNOR U14864 ( .A(a[2972]), .B(c2972), .Z(n8918) );
XOR U14865 ( .A(c2973), .B(n8919), .Z(c2974) );
ANDN U14866 ( .B(n8920), .A(n8921), .Z(n8919) );
XOR U14867 ( .A(c2973), .B(b[2973]), .Z(n8920) );
XNOR U14868 ( .A(b[2973]), .B(n8921), .Z(c[2973]) );
XNOR U14869 ( .A(a[2973]), .B(c2973), .Z(n8921) );
XOR U14870 ( .A(c2974), .B(n8922), .Z(c2975) );
ANDN U14871 ( .B(n8923), .A(n8924), .Z(n8922) );
XOR U14872 ( .A(c2974), .B(b[2974]), .Z(n8923) );
XNOR U14873 ( .A(b[2974]), .B(n8924), .Z(c[2974]) );
XNOR U14874 ( .A(a[2974]), .B(c2974), .Z(n8924) );
XOR U14875 ( .A(c2975), .B(n8925), .Z(c2976) );
ANDN U14876 ( .B(n8926), .A(n8927), .Z(n8925) );
XOR U14877 ( .A(c2975), .B(b[2975]), .Z(n8926) );
XNOR U14878 ( .A(b[2975]), .B(n8927), .Z(c[2975]) );
XNOR U14879 ( .A(a[2975]), .B(c2975), .Z(n8927) );
XOR U14880 ( .A(c2976), .B(n8928), .Z(c2977) );
ANDN U14881 ( .B(n8929), .A(n8930), .Z(n8928) );
XOR U14882 ( .A(c2976), .B(b[2976]), .Z(n8929) );
XNOR U14883 ( .A(b[2976]), .B(n8930), .Z(c[2976]) );
XNOR U14884 ( .A(a[2976]), .B(c2976), .Z(n8930) );
XOR U14885 ( .A(c2977), .B(n8931), .Z(c2978) );
ANDN U14886 ( .B(n8932), .A(n8933), .Z(n8931) );
XOR U14887 ( .A(c2977), .B(b[2977]), .Z(n8932) );
XNOR U14888 ( .A(b[2977]), .B(n8933), .Z(c[2977]) );
XNOR U14889 ( .A(a[2977]), .B(c2977), .Z(n8933) );
XOR U14890 ( .A(c2978), .B(n8934), .Z(c2979) );
ANDN U14891 ( .B(n8935), .A(n8936), .Z(n8934) );
XOR U14892 ( .A(c2978), .B(b[2978]), .Z(n8935) );
XNOR U14893 ( .A(b[2978]), .B(n8936), .Z(c[2978]) );
XNOR U14894 ( .A(a[2978]), .B(c2978), .Z(n8936) );
XOR U14895 ( .A(c2979), .B(n8937), .Z(c2980) );
ANDN U14896 ( .B(n8938), .A(n8939), .Z(n8937) );
XOR U14897 ( .A(c2979), .B(b[2979]), .Z(n8938) );
XNOR U14898 ( .A(b[2979]), .B(n8939), .Z(c[2979]) );
XNOR U14899 ( .A(a[2979]), .B(c2979), .Z(n8939) );
XOR U14900 ( .A(c2980), .B(n8940), .Z(c2981) );
ANDN U14901 ( .B(n8941), .A(n8942), .Z(n8940) );
XOR U14902 ( .A(c2980), .B(b[2980]), .Z(n8941) );
XNOR U14903 ( .A(b[2980]), .B(n8942), .Z(c[2980]) );
XNOR U14904 ( .A(a[2980]), .B(c2980), .Z(n8942) );
XOR U14905 ( .A(c2981), .B(n8943), .Z(c2982) );
ANDN U14906 ( .B(n8944), .A(n8945), .Z(n8943) );
XOR U14907 ( .A(c2981), .B(b[2981]), .Z(n8944) );
XNOR U14908 ( .A(b[2981]), .B(n8945), .Z(c[2981]) );
XNOR U14909 ( .A(a[2981]), .B(c2981), .Z(n8945) );
XOR U14910 ( .A(c2982), .B(n8946), .Z(c2983) );
ANDN U14911 ( .B(n8947), .A(n8948), .Z(n8946) );
XOR U14912 ( .A(c2982), .B(b[2982]), .Z(n8947) );
XNOR U14913 ( .A(b[2982]), .B(n8948), .Z(c[2982]) );
XNOR U14914 ( .A(a[2982]), .B(c2982), .Z(n8948) );
XOR U14915 ( .A(c2983), .B(n8949), .Z(c2984) );
ANDN U14916 ( .B(n8950), .A(n8951), .Z(n8949) );
XOR U14917 ( .A(c2983), .B(b[2983]), .Z(n8950) );
XNOR U14918 ( .A(b[2983]), .B(n8951), .Z(c[2983]) );
XNOR U14919 ( .A(a[2983]), .B(c2983), .Z(n8951) );
XOR U14920 ( .A(c2984), .B(n8952), .Z(c2985) );
ANDN U14921 ( .B(n8953), .A(n8954), .Z(n8952) );
XOR U14922 ( .A(c2984), .B(b[2984]), .Z(n8953) );
XNOR U14923 ( .A(b[2984]), .B(n8954), .Z(c[2984]) );
XNOR U14924 ( .A(a[2984]), .B(c2984), .Z(n8954) );
XOR U14925 ( .A(c2985), .B(n8955), .Z(c2986) );
ANDN U14926 ( .B(n8956), .A(n8957), .Z(n8955) );
XOR U14927 ( .A(c2985), .B(b[2985]), .Z(n8956) );
XNOR U14928 ( .A(b[2985]), .B(n8957), .Z(c[2985]) );
XNOR U14929 ( .A(a[2985]), .B(c2985), .Z(n8957) );
XOR U14930 ( .A(c2986), .B(n8958), .Z(c2987) );
ANDN U14931 ( .B(n8959), .A(n8960), .Z(n8958) );
XOR U14932 ( .A(c2986), .B(b[2986]), .Z(n8959) );
XNOR U14933 ( .A(b[2986]), .B(n8960), .Z(c[2986]) );
XNOR U14934 ( .A(a[2986]), .B(c2986), .Z(n8960) );
XOR U14935 ( .A(c2987), .B(n8961), .Z(c2988) );
ANDN U14936 ( .B(n8962), .A(n8963), .Z(n8961) );
XOR U14937 ( .A(c2987), .B(b[2987]), .Z(n8962) );
XNOR U14938 ( .A(b[2987]), .B(n8963), .Z(c[2987]) );
XNOR U14939 ( .A(a[2987]), .B(c2987), .Z(n8963) );
XOR U14940 ( .A(c2988), .B(n8964), .Z(c2989) );
ANDN U14941 ( .B(n8965), .A(n8966), .Z(n8964) );
XOR U14942 ( .A(c2988), .B(b[2988]), .Z(n8965) );
XNOR U14943 ( .A(b[2988]), .B(n8966), .Z(c[2988]) );
XNOR U14944 ( .A(a[2988]), .B(c2988), .Z(n8966) );
XOR U14945 ( .A(c2989), .B(n8967), .Z(c2990) );
ANDN U14946 ( .B(n8968), .A(n8969), .Z(n8967) );
XOR U14947 ( .A(c2989), .B(b[2989]), .Z(n8968) );
XNOR U14948 ( .A(b[2989]), .B(n8969), .Z(c[2989]) );
XNOR U14949 ( .A(a[2989]), .B(c2989), .Z(n8969) );
XOR U14950 ( .A(c2990), .B(n8970), .Z(c2991) );
ANDN U14951 ( .B(n8971), .A(n8972), .Z(n8970) );
XOR U14952 ( .A(c2990), .B(b[2990]), .Z(n8971) );
XNOR U14953 ( .A(b[2990]), .B(n8972), .Z(c[2990]) );
XNOR U14954 ( .A(a[2990]), .B(c2990), .Z(n8972) );
XOR U14955 ( .A(c2991), .B(n8973), .Z(c2992) );
ANDN U14956 ( .B(n8974), .A(n8975), .Z(n8973) );
XOR U14957 ( .A(c2991), .B(b[2991]), .Z(n8974) );
XNOR U14958 ( .A(b[2991]), .B(n8975), .Z(c[2991]) );
XNOR U14959 ( .A(a[2991]), .B(c2991), .Z(n8975) );
XOR U14960 ( .A(c2992), .B(n8976), .Z(c2993) );
ANDN U14961 ( .B(n8977), .A(n8978), .Z(n8976) );
XOR U14962 ( .A(c2992), .B(b[2992]), .Z(n8977) );
XNOR U14963 ( .A(b[2992]), .B(n8978), .Z(c[2992]) );
XNOR U14964 ( .A(a[2992]), .B(c2992), .Z(n8978) );
XOR U14965 ( .A(c2993), .B(n8979), .Z(c2994) );
ANDN U14966 ( .B(n8980), .A(n8981), .Z(n8979) );
XOR U14967 ( .A(c2993), .B(b[2993]), .Z(n8980) );
XNOR U14968 ( .A(b[2993]), .B(n8981), .Z(c[2993]) );
XNOR U14969 ( .A(a[2993]), .B(c2993), .Z(n8981) );
XOR U14970 ( .A(c2994), .B(n8982), .Z(c2995) );
ANDN U14971 ( .B(n8983), .A(n8984), .Z(n8982) );
XOR U14972 ( .A(c2994), .B(b[2994]), .Z(n8983) );
XNOR U14973 ( .A(b[2994]), .B(n8984), .Z(c[2994]) );
XNOR U14974 ( .A(a[2994]), .B(c2994), .Z(n8984) );
XOR U14975 ( .A(c2995), .B(n8985), .Z(c2996) );
ANDN U14976 ( .B(n8986), .A(n8987), .Z(n8985) );
XOR U14977 ( .A(c2995), .B(b[2995]), .Z(n8986) );
XNOR U14978 ( .A(b[2995]), .B(n8987), .Z(c[2995]) );
XNOR U14979 ( .A(a[2995]), .B(c2995), .Z(n8987) );
XOR U14980 ( .A(c2996), .B(n8988), .Z(c2997) );
ANDN U14981 ( .B(n8989), .A(n8990), .Z(n8988) );
XOR U14982 ( .A(c2996), .B(b[2996]), .Z(n8989) );
XNOR U14983 ( .A(b[2996]), .B(n8990), .Z(c[2996]) );
XNOR U14984 ( .A(a[2996]), .B(c2996), .Z(n8990) );
XOR U14985 ( .A(c2997), .B(n8991), .Z(c2998) );
ANDN U14986 ( .B(n8992), .A(n8993), .Z(n8991) );
XOR U14987 ( .A(c2997), .B(b[2997]), .Z(n8992) );
XNOR U14988 ( .A(b[2997]), .B(n8993), .Z(c[2997]) );
XNOR U14989 ( .A(a[2997]), .B(c2997), .Z(n8993) );
XOR U14990 ( .A(c2998), .B(n8994), .Z(c2999) );
ANDN U14991 ( .B(n8995), .A(n8996), .Z(n8994) );
XOR U14992 ( .A(c2998), .B(b[2998]), .Z(n8995) );
XNOR U14993 ( .A(b[2998]), .B(n8996), .Z(c[2998]) );
XNOR U14994 ( .A(a[2998]), .B(c2998), .Z(n8996) );
XOR U14995 ( .A(c2999), .B(n8997), .Z(c3000) );
ANDN U14996 ( .B(n8998), .A(n8999), .Z(n8997) );
XOR U14997 ( .A(c2999), .B(b[2999]), .Z(n8998) );
XNOR U14998 ( .A(b[2999]), .B(n8999), .Z(c[2999]) );
XNOR U14999 ( .A(a[2999]), .B(c2999), .Z(n8999) );
XOR U15000 ( .A(c3000), .B(n9000), .Z(c3001) );
ANDN U15001 ( .B(n9001), .A(n9002), .Z(n9000) );
XOR U15002 ( .A(c3000), .B(b[3000]), .Z(n9001) );
XNOR U15003 ( .A(b[3000]), .B(n9002), .Z(c[3000]) );
XNOR U15004 ( .A(a[3000]), .B(c3000), .Z(n9002) );
XOR U15005 ( .A(c3001), .B(n9003), .Z(c3002) );
ANDN U15006 ( .B(n9004), .A(n9005), .Z(n9003) );
XOR U15007 ( .A(c3001), .B(b[3001]), .Z(n9004) );
XNOR U15008 ( .A(b[3001]), .B(n9005), .Z(c[3001]) );
XNOR U15009 ( .A(a[3001]), .B(c3001), .Z(n9005) );
XOR U15010 ( .A(c3002), .B(n9006), .Z(c3003) );
ANDN U15011 ( .B(n9007), .A(n9008), .Z(n9006) );
XOR U15012 ( .A(c3002), .B(b[3002]), .Z(n9007) );
XNOR U15013 ( .A(b[3002]), .B(n9008), .Z(c[3002]) );
XNOR U15014 ( .A(a[3002]), .B(c3002), .Z(n9008) );
XOR U15015 ( .A(c3003), .B(n9009), .Z(c3004) );
ANDN U15016 ( .B(n9010), .A(n9011), .Z(n9009) );
XOR U15017 ( .A(c3003), .B(b[3003]), .Z(n9010) );
XNOR U15018 ( .A(b[3003]), .B(n9011), .Z(c[3003]) );
XNOR U15019 ( .A(a[3003]), .B(c3003), .Z(n9011) );
XOR U15020 ( .A(c3004), .B(n9012), .Z(c3005) );
ANDN U15021 ( .B(n9013), .A(n9014), .Z(n9012) );
XOR U15022 ( .A(c3004), .B(b[3004]), .Z(n9013) );
XNOR U15023 ( .A(b[3004]), .B(n9014), .Z(c[3004]) );
XNOR U15024 ( .A(a[3004]), .B(c3004), .Z(n9014) );
XOR U15025 ( .A(c3005), .B(n9015), .Z(c3006) );
ANDN U15026 ( .B(n9016), .A(n9017), .Z(n9015) );
XOR U15027 ( .A(c3005), .B(b[3005]), .Z(n9016) );
XNOR U15028 ( .A(b[3005]), .B(n9017), .Z(c[3005]) );
XNOR U15029 ( .A(a[3005]), .B(c3005), .Z(n9017) );
XOR U15030 ( .A(c3006), .B(n9018), .Z(c3007) );
ANDN U15031 ( .B(n9019), .A(n9020), .Z(n9018) );
XOR U15032 ( .A(c3006), .B(b[3006]), .Z(n9019) );
XNOR U15033 ( .A(b[3006]), .B(n9020), .Z(c[3006]) );
XNOR U15034 ( .A(a[3006]), .B(c3006), .Z(n9020) );
XOR U15035 ( .A(c3007), .B(n9021), .Z(c3008) );
ANDN U15036 ( .B(n9022), .A(n9023), .Z(n9021) );
XOR U15037 ( .A(c3007), .B(b[3007]), .Z(n9022) );
XNOR U15038 ( .A(b[3007]), .B(n9023), .Z(c[3007]) );
XNOR U15039 ( .A(a[3007]), .B(c3007), .Z(n9023) );
XOR U15040 ( .A(c3008), .B(n9024), .Z(c3009) );
ANDN U15041 ( .B(n9025), .A(n9026), .Z(n9024) );
XOR U15042 ( .A(c3008), .B(b[3008]), .Z(n9025) );
XNOR U15043 ( .A(b[3008]), .B(n9026), .Z(c[3008]) );
XNOR U15044 ( .A(a[3008]), .B(c3008), .Z(n9026) );
XOR U15045 ( .A(c3009), .B(n9027), .Z(c3010) );
ANDN U15046 ( .B(n9028), .A(n9029), .Z(n9027) );
XOR U15047 ( .A(c3009), .B(b[3009]), .Z(n9028) );
XNOR U15048 ( .A(b[3009]), .B(n9029), .Z(c[3009]) );
XNOR U15049 ( .A(a[3009]), .B(c3009), .Z(n9029) );
XOR U15050 ( .A(c3010), .B(n9030), .Z(c3011) );
ANDN U15051 ( .B(n9031), .A(n9032), .Z(n9030) );
XOR U15052 ( .A(c3010), .B(b[3010]), .Z(n9031) );
XNOR U15053 ( .A(b[3010]), .B(n9032), .Z(c[3010]) );
XNOR U15054 ( .A(a[3010]), .B(c3010), .Z(n9032) );
XOR U15055 ( .A(c3011), .B(n9033), .Z(c3012) );
ANDN U15056 ( .B(n9034), .A(n9035), .Z(n9033) );
XOR U15057 ( .A(c3011), .B(b[3011]), .Z(n9034) );
XNOR U15058 ( .A(b[3011]), .B(n9035), .Z(c[3011]) );
XNOR U15059 ( .A(a[3011]), .B(c3011), .Z(n9035) );
XOR U15060 ( .A(c3012), .B(n9036), .Z(c3013) );
ANDN U15061 ( .B(n9037), .A(n9038), .Z(n9036) );
XOR U15062 ( .A(c3012), .B(b[3012]), .Z(n9037) );
XNOR U15063 ( .A(b[3012]), .B(n9038), .Z(c[3012]) );
XNOR U15064 ( .A(a[3012]), .B(c3012), .Z(n9038) );
XOR U15065 ( .A(c3013), .B(n9039), .Z(c3014) );
ANDN U15066 ( .B(n9040), .A(n9041), .Z(n9039) );
XOR U15067 ( .A(c3013), .B(b[3013]), .Z(n9040) );
XNOR U15068 ( .A(b[3013]), .B(n9041), .Z(c[3013]) );
XNOR U15069 ( .A(a[3013]), .B(c3013), .Z(n9041) );
XOR U15070 ( .A(c3014), .B(n9042), .Z(c3015) );
ANDN U15071 ( .B(n9043), .A(n9044), .Z(n9042) );
XOR U15072 ( .A(c3014), .B(b[3014]), .Z(n9043) );
XNOR U15073 ( .A(b[3014]), .B(n9044), .Z(c[3014]) );
XNOR U15074 ( .A(a[3014]), .B(c3014), .Z(n9044) );
XOR U15075 ( .A(c3015), .B(n9045), .Z(c3016) );
ANDN U15076 ( .B(n9046), .A(n9047), .Z(n9045) );
XOR U15077 ( .A(c3015), .B(b[3015]), .Z(n9046) );
XNOR U15078 ( .A(b[3015]), .B(n9047), .Z(c[3015]) );
XNOR U15079 ( .A(a[3015]), .B(c3015), .Z(n9047) );
XOR U15080 ( .A(c3016), .B(n9048), .Z(c3017) );
ANDN U15081 ( .B(n9049), .A(n9050), .Z(n9048) );
XOR U15082 ( .A(c3016), .B(b[3016]), .Z(n9049) );
XNOR U15083 ( .A(b[3016]), .B(n9050), .Z(c[3016]) );
XNOR U15084 ( .A(a[3016]), .B(c3016), .Z(n9050) );
XOR U15085 ( .A(c3017), .B(n9051), .Z(c3018) );
ANDN U15086 ( .B(n9052), .A(n9053), .Z(n9051) );
XOR U15087 ( .A(c3017), .B(b[3017]), .Z(n9052) );
XNOR U15088 ( .A(b[3017]), .B(n9053), .Z(c[3017]) );
XNOR U15089 ( .A(a[3017]), .B(c3017), .Z(n9053) );
XOR U15090 ( .A(c3018), .B(n9054), .Z(c3019) );
ANDN U15091 ( .B(n9055), .A(n9056), .Z(n9054) );
XOR U15092 ( .A(c3018), .B(b[3018]), .Z(n9055) );
XNOR U15093 ( .A(b[3018]), .B(n9056), .Z(c[3018]) );
XNOR U15094 ( .A(a[3018]), .B(c3018), .Z(n9056) );
XOR U15095 ( .A(c3019), .B(n9057), .Z(c3020) );
ANDN U15096 ( .B(n9058), .A(n9059), .Z(n9057) );
XOR U15097 ( .A(c3019), .B(b[3019]), .Z(n9058) );
XNOR U15098 ( .A(b[3019]), .B(n9059), .Z(c[3019]) );
XNOR U15099 ( .A(a[3019]), .B(c3019), .Z(n9059) );
XOR U15100 ( .A(c3020), .B(n9060), .Z(c3021) );
ANDN U15101 ( .B(n9061), .A(n9062), .Z(n9060) );
XOR U15102 ( .A(c3020), .B(b[3020]), .Z(n9061) );
XNOR U15103 ( .A(b[3020]), .B(n9062), .Z(c[3020]) );
XNOR U15104 ( .A(a[3020]), .B(c3020), .Z(n9062) );
XOR U15105 ( .A(c3021), .B(n9063), .Z(c3022) );
ANDN U15106 ( .B(n9064), .A(n9065), .Z(n9063) );
XOR U15107 ( .A(c3021), .B(b[3021]), .Z(n9064) );
XNOR U15108 ( .A(b[3021]), .B(n9065), .Z(c[3021]) );
XNOR U15109 ( .A(a[3021]), .B(c3021), .Z(n9065) );
XOR U15110 ( .A(c3022), .B(n9066), .Z(c3023) );
ANDN U15111 ( .B(n9067), .A(n9068), .Z(n9066) );
XOR U15112 ( .A(c3022), .B(b[3022]), .Z(n9067) );
XNOR U15113 ( .A(b[3022]), .B(n9068), .Z(c[3022]) );
XNOR U15114 ( .A(a[3022]), .B(c3022), .Z(n9068) );
XOR U15115 ( .A(c3023), .B(n9069), .Z(c3024) );
ANDN U15116 ( .B(n9070), .A(n9071), .Z(n9069) );
XOR U15117 ( .A(c3023), .B(b[3023]), .Z(n9070) );
XNOR U15118 ( .A(b[3023]), .B(n9071), .Z(c[3023]) );
XNOR U15119 ( .A(a[3023]), .B(c3023), .Z(n9071) );
XOR U15120 ( .A(c3024), .B(n9072), .Z(c3025) );
ANDN U15121 ( .B(n9073), .A(n9074), .Z(n9072) );
XOR U15122 ( .A(c3024), .B(b[3024]), .Z(n9073) );
XNOR U15123 ( .A(b[3024]), .B(n9074), .Z(c[3024]) );
XNOR U15124 ( .A(a[3024]), .B(c3024), .Z(n9074) );
XOR U15125 ( .A(c3025), .B(n9075), .Z(c3026) );
ANDN U15126 ( .B(n9076), .A(n9077), .Z(n9075) );
XOR U15127 ( .A(c3025), .B(b[3025]), .Z(n9076) );
XNOR U15128 ( .A(b[3025]), .B(n9077), .Z(c[3025]) );
XNOR U15129 ( .A(a[3025]), .B(c3025), .Z(n9077) );
XOR U15130 ( .A(c3026), .B(n9078), .Z(c3027) );
ANDN U15131 ( .B(n9079), .A(n9080), .Z(n9078) );
XOR U15132 ( .A(c3026), .B(b[3026]), .Z(n9079) );
XNOR U15133 ( .A(b[3026]), .B(n9080), .Z(c[3026]) );
XNOR U15134 ( .A(a[3026]), .B(c3026), .Z(n9080) );
XOR U15135 ( .A(c3027), .B(n9081), .Z(c3028) );
ANDN U15136 ( .B(n9082), .A(n9083), .Z(n9081) );
XOR U15137 ( .A(c3027), .B(b[3027]), .Z(n9082) );
XNOR U15138 ( .A(b[3027]), .B(n9083), .Z(c[3027]) );
XNOR U15139 ( .A(a[3027]), .B(c3027), .Z(n9083) );
XOR U15140 ( .A(c3028), .B(n9084), .Z(c3029) );
ANDN U15141 ( .B(n9085), .A(n9086), .Z(n9084) );
XOR U15142 ( .A(c3028), .B(b[3028]), .Z(n9085) );
XNOR U15143 ( .A(b[3028]), .B(n9086), .Z(c[3028]) );
XNOR U15144 ( .A(a[3028]), .B(c3028), .Z(n9086) );
XOR U15145 ( .A(c3029), .B(n9087), .Z(c3030) );
ANDN U15146 ( .B(n9088), .A(n9089), .Z(n9087) );
XOR U15147 ( .A(c3029), .B(b[3029]), .Z(n9088) );
XNOR U15148 ( .A(b[3029]), .B(n9089), .Z(c[3029]) );
XNOR U15149 ( .A(a[3029]), .B(c3029), .Z(n9089) );
XOR U15150 ( .A(c3030), .B(n9090), .Z(c3031) );
ANDN U15151 ( .B(n9091), .A(n9092), .Z(n9090) );
XOR U15152 ( .A(c3030), .B(b[3030]), .Z(n9091) );
XNOR U15153 ( .A(b[3030]), .B(n9092), .Z(c[3030]) );
XNOR U15154 ( .A(a[3030]), .B(c3030), .Z(n9092) );
XOR U15155 ( .A(c3031), .B(n9093), .Z(c3032) );
ANDN U15156 ( .B(n9094), .A(n9095), .Z(n9093) );
XOR U15157 ( .A(c3031), .B(b[3031]), .Z(n9094) );
XNOR U15158 ( .A(b[3031]), .B(n9095), .Z(c[3031]) );
XNOR U15159 ( .A(a[3031]), .B(c3031), .Z(n9095) );
XOR U15160 ( .A(c3032), .B(n9096), .Z(c3033) );
ANDN U15161 ( .B(n9097), .A(n9098), .Z(n9096) );
XOR U15162 ( .A(c3032), .B(b[3032]), .Z(n9097) );
XNOR U15163 ( .A(b[3032]), .B(n9098), .Z(c[3032]) );
XNOR U15164 ( .A(a[3032]), .B(c3032), .Z(n9098) );
XOR U15165 ( .A(c3033), .B(n9099), .Z(c3034) );
ANDN U15166 ( .B(n9100), .A(n9101), .Z(n9099) );
XOR U15167 ( .A(c3033), .B(b[3033]), .Z(n9100) );
XNOR U15168 ( .A(b[3033]), .B(n9101), .Z(c[3033]) );
XNOR U15169 ( .A(a[3033]), .B(c3033), .Z(n9101) );
XOR U15170 ( .A(c3034), .B(n9102), .Z(c3035) );
ANDN U15171 ( .B(n9103), .A(n9104), .Z(n9102) );
XOR U15172 ( .A(c3034), .B(b[3034]), .Z(n9103) );
XNOR U15173 ( .A(b[3034]), .B(n9104), .Z(c[3034]) );
XNOR U15174 ( .A(a[3034]), .B(c3034), .Z(n9104) );
XOR U15175 ( .A(c3035), .B(n9105), .Z(c3036) );
ANDN U15176 ( .B(n9106), .A(n9107), .Z(n9105) );
XOR U15177 ( .A(c3035), .B(b[3035]), .Z(n9106) );
XNOR U15178 ( .A(b[3035]), .B(n9107), .Z(c[3035]) );
XNOR U15179 ( .A(a[3035]), .B(c3035), .Z(n9107) );
XOR U15180 ( .A(c3036), .B(n9108), .Z(c3037) );
ANDN U15181 ( .B(n9109), .A(n9110), .Z(n9108) );
XOR U15182 ( .A(c3036), .B(b[3036]), .Z(n9109) );
XNOR U15183 ( .A(b[3036]), .B(n9110), .Z(c[3036]) );
XNOR U15184 ( .A(a[3036]), .B(c3036), .Z(n9110) );
XOR U15185 ( .A(c3037), .B(n9111), .Z(c3038) );
ANDN U15186 ( .B(n9112), .A(n9113), .Z(n9111) );
XOR U15187 ( .A(c3037), .B(b[3037]), .Z(n9112) );
XNOR U15188 ( .A(b[3037]), .B(n9113), .Z(c[3037]) );
XNOR U15189 ( .A(a[3037]), .B(c3037), .Z(n9113) );
XOR U15190 ( .A(c3038), .B(n9114), .Z(c3039) );
ANDN U15191 ( .B(n9115), .A(n9116), .Z(n9114) );
XOR U15192 ( .A(c3038), .B(b[3038]), .Z(n9115) );
XNOR U15193 ( .A(b[3038]), .B(n9116), .Z(c[3038]) );
XNOR U15194 ( .A(a[3038]), .B(c3038), .Z(n9116) );
XOR U15195 ( .A(c3039), .B(n9117), .Z(c3040) );
ANDN U15196 ( .B(n9118), .A(n9119), .Z(n9117) );
XOR U15197 ( .A(c3039), .B(b[3039]), .Z(n9118) );
XNOR U15198 ( .A(b[3039]), .B(n9119), .Z(c[3039]) );
XNOR U15199 ( .A(a[3039]), .B(c3039), .Z(n9119) );
XOR U15200 ( .A(c3040), .B(n9120), .Z(c3041) );
ANDN U15201 ( .B(n9121), .A(n9122), .Z(n9120) );
XOR U15202 ( .A(c3040), .B(b[3040]), .Z(n9121) );
XNOR U15203 ( .A(b[3040]), .B(n9122), .Z(c[3040]) );
XNOR U15204 ( .A(a[3040]), .B(c3040), .Z(n9122) );
XOR U15205 ( .A(c3041), .B(n9123), .Z(c3042) );
ANDN U15206 ( .B(n9124), .A(n9125), .Z(n9123) );
XOR U15207 ( .A(c3041), .B(b[3041]), .Z(n9124) );
XNOR U15208 ( .A(b[3041]), .B(n9125), .Z(c[3041]) );
XNOR U15209 ( .A(a[3041]), .B(c3041), .Z(n9125) );
XOR U15210 ( .A(c3042), .B(n9126), .Z(c3043) );
ANDN U15211 ( .B(n9127), .A(n9128), .Z(n9126) );
XOR U15212 ( .A(c3042), .B(b[3042]), .Z(n9127) );
XNOR U15213 ( .A(b[3042]), .B(n9128), .Z(c[3042]) );
XNOR U15214 ( .A(a[3042]), .B(c3042), .Z(n9128) );
XOR U15215 ( .A(c3043), .B(n9129), .Z(c3044) );
ANDN U15216 ( .B(n9130), .A(n9131), .Z(n9129) );
XOR U15217 ( .A(c3043), .B(b[3043]), .Z(n9130) );
XNOR U15218 ( .A(b[3043]), .B(n9131), .Z(c[3043]) );
XNOR U15219 ( .A(a[3043]), .B(c3043), .Z(n9131) );
XOR U15220 ( .A(c3044), .B(n9132), .Z(c3045) );
ANDN U15221 ( .B(n9133), .A(n9134), .Z(n9132) );
XOR U15222 ( .A(c3044), .B(b[3044]), .Z(n9133) );
XNOR U15223 ( .A(b[3044]), .B(n9134), .Z(c[3044]) );
XNOR U15224 ( .A(a[3044]), .B(c3044), .Z(n9134) );
XOR U15225 ( .A(c3045), .B(n9135), .Z(c3046) );
ANDN U15226 ( .B(n9136), .A(n9137), .Z(n9135) );
XOR U15227 ( .A(c3045), .B(b[3045]), .Z(n9136) );
XNOR U15228 ( .A(b[3045]), .B(n9137), .Z(c[3045]) );
XNOR U15229 ( .A(a[3045]), .B(c3045), .Z(n9137) );
XOR U15230 ( .A(c3046), .B(n9138), .Z(c3047) );
ANDN U15231 ( .B(n9139), .A(n9140), .Z(n9138) );
XOR U15232 ( .A(c3046), .B(b[3046]), .Z(n9139) );
XNOR U15233 ( .A(b[3046]), .B(n9140), .Z(c[3046]) );
XNOR U15234 ( .A(a[3046]), .B(c3046), .Z(n9140) );
XOR U15235 ( .A(c3047), .B(n9141), .Z(c3048) );
ANDN U15236 ( .B(n9142), .A(n9143), .Z(n9141) );
XOR U15237 ( .A(c3047), .B(b[3047]), .Z(n9142) );
XNOR U15238 ( .A(b[3047]), .B(n9143), .Z(c[3047]) );
XNOR U15239 ( .A(a[3047]), .B(c3047), .Z(n9143) );
XOR U15240 ( .A(c3048), .B(n9144), .Z(c3049) );
ANDN U15241 ( .B(n9145), .A(n9146), .Z(n9144) );
XOR U15242 ( .A(c3048), .B(b[3048]), .Z(n9145) );
XNOR U15243 ( .A(b[3048]), .B(n9146), .Z(c[3048]) );
XNOR U15244 ( .A(a[3048]), .B(c3048), .Z(n9146) );
XOR U15245 ( .A(c3049), .B(n9147), .Z(c3050) );
ANDN U15246 ( .B(n9148), .A(n9149), .Z(n9147) );
XOR U15247 ( .A(c3049), .B(b[3049]), .Z(n9148) );
XNOR U15248 ( .A(b[3049]), .B(n9149), .Z(c[3049]) );
XNOR U15249 ( .A(a[3049]), .B(c3049), .Z(n9149) );
XOR U15250 ( .A(c3050), .B(n9150), .Z(c3051) );
ANDN U15251 ( .B(n9151), .A(n9152), .Z(n9150) );
XOR U15252 ( .A(c3050), .B(b[3050]), .Z(n9151) );
XNOR U15253 ( .A(b[3050]), .B(n9152), .Z(c[3050]) );
XNOR U15254 ( .A(a[3050]), .B(c3050), .Z(n9152) );
XOR U15255 ( .A(c3051), .B(n9153), .Z(c3052) );
ANDN U15256 ( .B(n9154), .A(n9155), .Z(n9153) );
XOR U15257 ( .A(c3051), .B(b[3051]), .Z(n9154) );
XNOR U15258 ( .A(b[3051]), .B(n9155), .Z(c[3051]) );
XNOR U15259 ( .A(a[3051]), .B(c3051), .Z(n9155) );
XOR U15260 ( .A(c3052), .B(n9156), .Z(c3053) );
ANDN U15261 ( .B(n9157), .A(n9158), .Z(n9156) );
XOR U15262 ( .A(c3052), .B(b[3052]), .Z(n9157) );
XNOR U15263 ( .A(b[3052]), .B(n9158), .Z(c[3052]) );
XNOR U15264 ( .A(a[3052]), .B(c3052), .Z(n9158) );
XOR U15265 ( .A(c3053), .B(n9159), .Z(c3054) );
ANDN U15266 ( .B(n9160), .A(n9161), .Z(n9159) );
XOR U15267 ( .A(c3053), .B(b[3053]), .Z(n9160) );
XNOR U15268 ( .A(b[3053]), .B(n9161), .Z(c[3053]) );
XNOR U15269 ( .A(a[3053]), .B(c3053), .Z(n9161) );
XOR U15270 ( .A(c3054), .B(n9162), .Z(c3055) );
ANDN U15271 ( .B(n9163), .A(n9164), .Z(n9162) );
XOR U15272 ( .A(c3054), .B(b[3054]), .Z(n9163) );
XNOR U15273 ( .A(b[3054]), .B(n9164), .Z(c[3054]) );
XNOR U15274 ( .A(a[3054]), .B(c3054), .Z(n9164) );
XOR U15275 ( .A(c3055), .B(n9165), .Z(c3056) );
ANDN U15276 ( .B(n9166), .A(n9167), .Z(n9165) );
XOR U15277 ( .A(c3055), .B(b[3055]), .Z(n9166) );
XNOR U15278 ( .A(b[3055]), .B(n9167), .Z(c[3055]) );
XNOR U15279 ( .A(a[3055]), .B(c3055), .Z(n9167) );
XOR U15280 ( .A(c3056), .B(n9168), .Z(c3057) );
ANDN U15281 ( .B(n9169), .A(n9170), .Z(n9168) );
XOR U15282 ( .A(c3056), .B(b[3056]), .Z(n9169) );
XNOR U15283 ( .A(b[3056]), .B(n9170), .Z(c[3056]) );
XNOR U15284 ( .A(a[3056]), .B(c3056), .Z(n9170) );
XOR U15285 ( .A(c3057), .B(n9171), .Z(c3058) );
ANDN U15286 ( .B(n9172), .A(n9173), .Z(n9171) );
XOR U15287 ( .A(c3057), .B(b[3057]), .Z(n9172) );
XNOR U15288 ( .A(b[3057]), .B(n9173), .Z(c[3057]) );
XNOR U15289 ( .A(a[3057]), .B(c3057), .Z(n9173) );
XOR U15290 ( .A(c3058), .B(n9174), .Z(c3059) );
ANDN U15291 ( .B(n9175), .A(n9176), .Z(n9174) );
XOR U15292 ( .A(c3058), .B(b[3058]), .Z(n9175) );
XNOR U15293 ( .A(b[3058]), .B(n9176), .Z(c[3058]) );
XNOR U15294 ( .A(a[3058]), .B(c3058), .Z(n9176) );
XOR U15295 ( .A(c3059), .B(n9177), .Z(c3060) );
ANDN U15296 ( .B(n9178), .A(n9179), .Z(n9177) );
XOR U15297 ( .A(c3059), .B(b[3059]), .Z(n9178) );
XNOR U15298 ( .A(b[3059]), .B(n9179), .Z(c[3059]) );
XNOR U15299 ( .A(a[3059]), .B(c3059), .Z(n9179) );
XOR U15300 ( .A(c3060), .B(n9180), .Z(c3061) );
ANDN U15301 ( .B(n9181), .A(n9182), .Z(n9180) );
XOR U15302 ( .A(c3060), .B(b[3060]), .Z(n9181) );
XNOR U15303 ( .A(b[3060]), .B(n9182), .Z(c[3060]) );
XNOR U15304 ( .A(a[3060]), .B(c3060), .Z(n9182) );
XOR U15305 ( .A(c3061), .B(n9183), .Z(c3062) );
ANDN U15306 ( .B(n9184), .A(n9185), .Z(n9183) );
XOR U15307 ( .A(c3061), .B(b[3061]), .Z(n9184) );
XNOR U15308 ( .A(b[3061]), .B(n9185), .Z(c[3061]) );
XNOR U15309 ( .A(a[3061]), .B(c3061), .Z(n9185) );
XOR U15310 ( .A(c3062), .B(n9186), .Z(c3063) );
ANDN U15311 ( .B(n9187), .A(n9188), .Z(n9186) );
XOR U15312 ( .A(c3062), .B(b[3062]), .Z(n9187) );
XNOR U15313 ( .A(b[3062]), .B(n9188), .Z(c[3062]) );
XNOR U15314 ( .A(a[3062]), .B(c3062), .Z(n9188) );
XOR U15315 ( .A(c3063), .B(n9189), .Z(c3064) );
ANDN U15316 ( .B(n9190), .A(n9191), .Z(n9189) );
XOR U15317 ( .A(c3063), .B(b[3063]), .Z(n9190) );
XNOR U15318 ( .A(b[3063]), .B(n9191), .Z(c[3063]) );
XNOR U15319 ( .A(a[3063]), .B(c3063), .Z(n9191) );
XOR U15320 ( .A(c3064), .B(n9192), .Z(c3065) );
ANDN U15321 ( .B(n9193), .A(n9194), .Z(n9192) );
XOR U15322 ( .A(c3064), .B(b[3064]), .Z(n9193) );
XNOR U15323 ( .A(b[3064]), .B(n9194), .Z(c[3064]) );
XNOR U15324 ( .A(a[3064]), .B(c3064), .Z(n9194) );
XOR U15325 ( .A(c3065), .B(n9195), .Z(c3066) );
ANDN U15326 ( .B(n9196), .A(n9197), .Z(n9195) );
XOR U15327 ( .A(c3065), .B(b[3065]), .Z(n9196) );
XNOR U15328 ( .A(b[3065]), .B(n9197), .Z(c[3065]) );
XNOR U15329 ( .A(a[3065]), .B(c3065), .Z(n9197) );
XOR U15330 ( .A(c3066), .B(n9198), .Z(c3067) );
ANDN U15331 ( .B(n9199), .A(n9200), .Z(n9198) );
XOR U15332 ( .A(c3066), .B(b[3066]), .Z(n9199) );
XNOR U15333 ( .A(b[3066]), .B(n9200), .Z(c[3066]) );
XNOR U15334 ( .A(a[3066]), .B(c3066), .Z(n9200) );
XOR U15335 ( .A(c3067), .B(n9201), .Z(c3068) );
ANDN U15336 ( .B(n9202), .A(n9203), .Z(n9201) );
XOR U15337 ( .A(c3067), .B(b[3067]), .Z(n9202) );
XNOR U15338 ( .A(b[3067]), .B(n9203), .Z(c[3067]) );
XNOR U15339 ( .A(a[3067]), .B(c3067), .Z(n9203) );
XOR U15340 ( .A(c3068), .B(n9204), .Z(c3069) );
ANDN U15341 ( .B(n9205), .A(n9206), .Z(n9204) );
XOR U15342 ( .A(c3068), .B(b[3068]), .Z(n9205) );
XNOR U15343 ( .A(b[3068]), .B(n9206), .Z(c[3068]) );
XNOR U15344 ( .A(a[3068]), .B(c3068), .Z(n9206) );
XOR U15345 ( .A(c3069), .B(n9207), .Z(c3070) );
ANDN U15346 ( .B(n9208), .A(n9209), .Z(n9207) );
XOR U15347 ( .A(c3069), .B(b[3069]), .Z(n9208) );
XNOR U15348 ( .A(b[3069]), .B(n9209), .Z(c[3069]) );
XNOR U15349 ( .A(a[3069]), .B(c3069), .Z(n9209) );
XOR U15350 ( .A(c3070), .B(n9210), .Z(c3071) );
ANDN U15351 ( .B(n9211), .A(n9212), .Z(n9210) );
XOR U15352 ( .A(c3070), .B(b[3070]), .Z(n9211) );
XNOR U15353 ( .A(b[3070]), .B(n9212), .Z(c[3070]) );
XNOR U15354 ( .A(a[3070]), .B(c3070), .Z(n9212) );
XOR U15355 ( .A(c3071), .B(n9213), .Z(c3072) );
ANDN U15356 ( .B(n9214), .A(n9215), .Z(n9213) );
XOR U15357 ( .A(c3071), .B(b[3071]), .Z(n9214) );
XNOR U15358 ( .A(b[3071]), .B(n9215), .Z(c[3071]) );
XNOR U15359 ( .A(a[3071]), .B(c3071), .Z(n9215) );
XOR U15360 ( .A(c3072), .B(n9216), .Z(c3073) );
ANDN U15361 ( .B(n9217), .A(n9218), .Z(n9216) );
XOR U15362 ( .A(c3072), .B(b[3072]), .Z(n9217) );
XNOR U15363 ( .A(b[3072]), .B(n9218), .Z(c[3072]) );
XNOR U15364 ( .A(a[3072]), .B(c3072), .Z(n9218) );
XOR U15365 ( .A(c3073), .B(n9219), .Z(c3074) );
ANDN U15366 ( .B(n9220), .A(n9221), .Z(n9219) );
XOR U15367 ( .A(c3073), .B(b[3073]), .Z(n9220) );
XNOR U15368 ( .A(b[3073]), .B(n9221), .Z(c[3073]) );
XNOR U15369 ( .A(a[3073]), .B(c3073), .Z(n9221) );
XOR U15370 ( .A(c3074), .B(n9222), .Z(c3075) );
ANDN U15371 ( .B(n9223), .A(n9224), .Z(n9222) );
XOR U15372 ( .A(c3074), .B(b[3074]), .Z(n9223) );
XNOR U15373 ( .A(b[3074]), .B(n9224), .Z(c[3074]) );
XNOR U15374 ( .A(a[3074]), .B(c3074), .Z(n9224) );
XOR U15375 ( .A(c3075), .B(n9225), .Z(c3076) );
ANDN U15376 ( .B(n9226), .A(n9227), .Z(n9225) );
XOR U15377 ( .A(c3075), .B(b[3075]), .Z(n9226) );
XNOR U15378 ( .A(b[3075]), .B(n9227), .Z(c[3075]) );
XNOR U15379 ( .A(a[3075]), .B(c3075), .Z(n9227) );
XOR U15380 ( .A(c3076), .B(n9228), .Z(c3077) );
ANDN U15381 ( .B(n9229), .A(n9230), .Z(n9228) );
XOR U15382 ( .A(c3076), .B(b[3076]), .Z(n9229) );
XNOR U15383 ( .A(b[3076]), .B(n9230), .Z(c[3076]) );
XNOR U15384 ( .A(a[3076]), .B(c3076), .Z(n9230) );
XOR U15385 ( .A(c3077), .B(n9231), .Z(c3078) );
ANDN U15386 ( .B(n9232), .A(n9233), .Z(n9231) );
XOR U15387 ( .A(c3077), .B(b[3077]), .Z(n9232) );
XNOR U15388 ( .A(b[3077]), .B(n9233), .Z(c[3077]) );
XNOR U15389 ( .A(a[3077]), .B(c3077), .Z(n9233) );
XOR U15390 ( .A(c3078), .B(n9234), .Z(c3079) );
ANDN U15391 ( .B(n9235), .A(n9236), .Z(n9234) );
XOR U15392 ( .A(c3078), .B(b[3078]), .Z(n9235) );
XNOR U15393 ( .A(b[3078]), .B(n9236), .Z(c[3078]) );
XNOR U15394 ( .A(a[3078]), .B(c3078), .Z(n9236) );
XOR U15395 ( .A(c3079), .B(n9237), .Z(c3080) );
ANDN U15396 ( .B(n9238), .A(n9239), .Z(n9237) );
XOR U15397 ( .A(c3079), .B(b[3079]), .Z(n9238) );
XNOR U15398 ( .A(b[3079]), .B(n9239), .Z(c[3079]) );
XNOR U15399 ( .A(a[3079]), .B(c3079), .Z(n9239) );
XOR U15400 ( .A(c3080), .B(n9240), .Z(c3081) );
ANDN U15401 ( .B(n9241), .A(n9242), .Z(n9240) );
XOR U15402 ( .A(c3080), .B(b[3080]), .Z(n9241) );
XNOR U15403 ( .A(b[3080]), .B(n9242), .Z(c[3080]) );
XNOR U15404 ( .A(a[3080]), .B(c3080), .Z(n9242) );
XOR U15405 ( .A(c3081), .B(n9243), .Z(c3082) );
ANDN U15406 ( .B(n9244), .A(n9245), .Z(n9243) );
XOR U15407 ( .A(c3081), .B(b[3081]), .Z(n9244) );
XNOR U15408 ( .A(b[3081]), .B(n9245), .Z(c[3081]) );
XNOR U15409 ( .A(a[3081]), .B(c3081), .Z(n9245) );
XOR U15410 ( .A(c3082), .B(n9246), .Z(c3083) );
ANDN U15411 ( .B(n9247), .A(n9248), .Z(n9246) );
XOR U15412 ( .A(c3082), .B(b[3082]), .Z(n9247) );
XNOR U15413 ( .A(b[3082]), .B(n9248), .Z(c[3082]) );
XNOR U15414 ( .A(a[3082]), .B(c3082), .Z(n9248) );
XOR U15415 ( .A(c3083), .B(n9249), .Z(c3084) );
ANDN U15416 ( .B(n9250), .A(n9251), .Z(n9249) );
XOR U15417 ( .A(c3083), .B(b[3083]), .Z(n9250) );
XNOR U15418 ( .A(b[3083]), .B(n9251), .Z(c[3083]) );
XNOR U15419 ( .A(a[3083]), .B(c3083), .Z(n9251) );
XOR U15420 ( .A(c3084), .B(n9252), .Z(c3085) );
ANDN U15421 ( .B(n9253), .A(n9254), .Z(n9252) );
XOR U15422 ( .A(c3084), .B(b[3084]), .Z(n9253) );
XNOR U15423 ( .A(b[3084]), .B(n9254), .Z(c[3084]) );
XNOR U15424 ( .A(a[3084]), .B(c3084), .Z(n9254) );
XOR U15425 ( .A(c3085), .B(n9255), .Z(c3086) );
ANDN U15426 ( .B(n9256), .A(n9257), .Z(n9255) );
XOR U15427 ( .A(c3085), .B(b[3085]), .Z(n9256) );
XNOR U15428 ( .A(b[3085]), .B(n9257), .Z(c[3085]) );
XNOR U15429 ( .A(a[3085]), .B(c3085), .Z(n9257) );
XOR U15430 ( .A(c3086), .B(n9258), .Z(c3087) );
ANDN U15431 ( .B(n9259), .A(n9260), .Z(n9258) );
XOR U15432 ( .A(c3086), .B(b[3086]), .Z(n9259) );
XNOR U15433 ( .A(b[3086]), .B(n9260), .Z(c[3086]) );
XNOR U15434 ( .A(a[3086]), .B(c3086), .Z(n9260) );
XOR U15435 ( .A(c3087), .B(n9261), .Z(c3088) );
ANDN U15436 ( .B(n9262), .A(n9263), .Z(n9261) );
XOR U15437 ( .A(c3087), .B(b[3087]), .Z(n9262) );
XNOR U15438 ( .A(b[3087]), .B(n9263), .Z(c[3087]) );
XNOR U15439 ( .A(a[3087]), .B(c3087), .Z(n9263) );
XOR U15440 ( .A(c3088), .B(n9264), .Z(c3089) );
ANDN U15441 ( .B(n9265), .A(n9266), .Z(n9264) );
XOR U15442 ( .A(c3088), .B(b[3088]), .Z(n9265) );
XNOR U15443 ( .A(b[3088]), .B(n9266), .Z(c[3088]) );
XNOR U15444 ( .A(a[3088]), .B(c3088), .Z(n9266) );
XOR U15445 ( .A(c3089), .B(n9267), .Z(c3090) );
ANDN U15446 ( .B(n9268), .A(n9269), .Z(n9267) );
XOR U15447 ( .A(c3089), .B(b[3089]), .Z(n9268) );
XNOR U15448 ( .A(b[3089]), .B(n9269), .Z(c[3089]) );
XNOR U15449 ( .A(a[3089]), .B(c3089), .Z(n9269) );
XOR U15450 ( .A(c3090), .B(n9270), .Z(c3091) );
ANDN U15451 ( .B(n9271), .A(n9272), .Z(n9270) );
XOR U15452 ( .A(c3090), .B(b[3090]), .Z(n9271) );
XNOR U15453 ( .A(b[3090]), .B(n9272), .Z(c[3090]) );
XNOR U15454 ( .A(a[3090]), .B(c3090), .Z(n9272) );
XOR U15455 ( .A(c3091), .B(n9273), .Z(c3092) );
ANDN U15456 ( .B(n9274), .A(n9275), .Z(n9273) );
XOR U15457 ( .A(c3091), .B(b[3091]), .Z(n9274) );
XNOR U15458 ( .A(b[3091]), .B(n9275), .Z(c[3091]) );
XNOR U15459 ( .A(a[3091]), .B(c3091), .Z(n9275) );
XOR U15460 ( .A(c3092), .B(n9276), .Z(c3093) );
ANDN U15461 ( .B(n9277), .A(n9278), .Z(n9276) );
XOR U15462 ( .A(c3092), .B(b[3092]), .Z(n9277) );
XNOR U15463 ( .A(b[3092]), .B(n9278), .Z(c[3092]) );
XNOR U15464 ( .A(a[3092]), .B(c3092), .Z(n9278) );
XOR U15465 ( .A(c3093), .B(n9279), .Z(c3094) );
ANDN U15466 ( .B(n9280), .A(n9281), .Z(n9279) );
XOR U15467 ( .A(c3093), .B(b[3093]), .Z(n9280) );
XNOR U15468 ( .A(b[3093]), .B(n9281), .Z(c[3093]) );
XNOR U15469 ( .A(a[3093]), .B(c3093), .Z(n9281) );
XOR U15470 ( .A(c3094), .B(n9282), .Z(c3095) );
ANDN U15471 ( .B(n9283), .A(n9284), .Z(n9282) );
XOR U15472 ( .A(c3094), .B(b[3094]), .Z(n9283) );
XNOR U15473 ( .A(b[3094]), .B(n9284), .Z(c[3094]) );
XNOR U15474 ( .A(a[3094]), .B(c3094), .Z(n9284) );
XOR U15475 ( .A(c3095), .B(n9285), .Z(c3096) );
ANDN U15476 ( .B(n9286), .A(n9287), .Z(n9285) );
XOR U15477 ( .A(c3095), .B(b[3095]), .Z(n9286) );
XNOR U15478 ( .A(b[3095]), .B(n9287), .Z(c[3095]) );
XNOR U15479 ( .A(a[3095]), .B(c3095), .Z(n9287) );
XOR U15480 ( .A(c3096), .B(n9288), .Z(c3097) );
ANDN U15481 ( .B(n9289), .A(n9290), .Z(n9288) );
XOR U15482 ( .A(c3096), .B(b[3096]), .Z(n9289) );
XNOR U15483 ( .A(b[3096]), .B(n9290), .Z(c[3096]) );
XNOR U15484 ( .A(a[3096]), .B(c3096), .Z(n9290) );
XOR U15485 ( .A(c3097), .B(n9291), .Z(c3098) );
ANDN U15486 ( .B(n9292), .A(n9293), .Z(n9291) );
XOR U15487 ( .A(c3097), .B(b[3097]), .Z(n9292) );
XNOR U15488 ( .A(b[3097]), .B(n9293), .Z(c[3097]) );
XNOR U15489 ( .A(a[3097]), .B(c3097), .Z(n9293) );
XOR U15490 ( .A(c3098), .B(n9294), .Z(c3099) );
ANDN U15491 ( .B(n9295), .A(n9296), .Z(n9294) );
XOR U15492 ( .A(c3098), .B(b[3098]), .Z(n9295) );
XNOR U15493 ( .A(b[3098]), .B(n9296), .Z(c[3098]) );
XNOR U15494 ( .A(a[3098]), .B(c3098), .Z(n9296) );
XOR U15495 ( .A(c3099), .B(n9297), .Z(c3100) );
ANDN U15496 ( .B(n9298), .A(n9299), .Z(n9297) );
XOR U15497 ( .A(c3099), .B(b[3099]), .Z(n9298) );
XNOR U15498 ( .A(b[3099]), .B(n9299), .Z(c[3099]) );
XNOR U15499 ( .A(a[3099]), .B(c3099), .Z(n9299) );
XOR U15500 ( .A(c3100), .B(n9300), .Z(c3101) );
ANDN U15501 ( .B(n9301), .A(n9302), .Z(n9300) );
XOR U15502 ( .A(c3100), .B(b[3100]), .Z(n9301) );
XNOR U15503 ( .A(b[3100]), .B(n9302), .Z(c[3100]) );
XNOR U15504 ( .A(a[3100]), .B(c3100), .Z(n9302) );
XOR U15505 ( .A(c3101), .B(n9303), .Z(c3102) );
ANDN U15506 ( .B(n9304), .A(n9305), .Z(n9303) );
XOR U15507 ( .A(c3101), .B(b[3101]), .Z(n9304) );
XNOR U15508 ( .A(b[3101]), .B(n9305), .Z(c[3101]) );
XNOR U15509 ( .A(a[3101]), .B(c3101), .Z(n9305) );
XOR U15510 ( .A(c3102), .B(n9306), .Z(c3103) );
ANDN U15511 ( .B(n9307), .A(n9308), .Z(n9306) );
XOR U15512 ( .A(c3102), .B(b[3102]), .Z(n9307) );
XNOR U15513 ( .A(b[3102]), .B(n9308), .Z(c[3102]) );
XNOR U15514 ( .A(a[3102]), .B(c3102), .Z(n9308) );
XOR U15515 ( .A(c3103), .B(n9309), .Z(c3104) );
ANDN U15516 ( .B(n9310), .A(n9311), .Z(n9309) );
XOR U15517 ( .A(c3103), .B(b[3103]), .Z(n9310) );
XNOR U15518 ( .A(b[3103]), .B(n9311), .Z(c[3103]) );
XNOR U15519 ( .A(a[3103]), .B(c3103), .Z(n9311) );
XOR U15520 ( .A(c3104), .B(n9312), .Z(c3105) );
ANDN U15521 ( .B(n9313), .A(n9314), .Z(n9312) );
XOR U15522 ( .A(c3104), .B(b[3104]), .Z(n9313) );
XNOR U15523 ( .A(b[3104]), .B(n9314), .Z(c[3104]) );
XNOR U15524 ( .A(a[3104]), .B(c3104), .Z(n9314) );
XOR U15525 ( .A(c3105), .B(n9315), .Z(c3106) );
ANDN U15526 ( .B(n9316), .A(n9317), .Z(n9315) );
XOR U15527 ( .A(c3105), .B(b[3105]), .Z(n9316) );
XNOR U15528 ( .A(b[3105]), .B(n9317), .Z(c[3105]) );
XNOR U15529 ( .A(a[3105]), .B(c3105), .Z(n9317) );
XOR U15530 ( .A(c3106), .B(n9318), .Z(c3107) );
ANDN U15531 ( .B(n9319), .A(n9320), .Z(n9318) );
XOR U15532 ( .A(c3106), .B(b[3106]), .Z(n9319) );
XNOR U15533 ( .A(b[3106]), .B(n9320), .Z(c[3106]) );
XNOR U15534 ( .A(a[3106]), .B(c3106), .Z(n9320) );
XOR U15535 ( .A(c3107), .B(n9321), .Z(c3108) );
ANDN U15536 ( .B(n9322), .A(n9323), .Z(n9321) );
XOR U15537 ( .A(c3107), .B(b[3107]), .Z(n9322) );
XNOR U15538 ( .A(b[3107]), .B(n9323), .Z(c[3107]) );
XNOR U15539 ( .A(a[3107]), .B(c3107), .Z(n9323) );
XOR U15540 ( .A(c3108), .B(n9324), .Z(c3109) );
ANDN U15541 ( .B(n9325), .A(n9326), .Z(n9324) );
XOR U15542 ( .A(c3108), .B(b[3108]), .Z(n9325) );
XNOR U15543 ( .A(b[3108]), .B(n9326), .Z(c[3108]) );
XNOR U15544 ( .A(a[3108]), .B(c3108), .Z(n9326) );
XOR U15545 ( .A(c3109), .B(n9327), .Z(c3110) );
ANDN U15546 ( .B(n9328), .A(n9329), .Z(n9327) );
XOR U15547 ( .A(c3109), .B(b[3109]), .Z(n9328) );
XNOR U15548 ( .A(b[3109]), .B(n9329), .Z(c[3109]) );
XNOR U15549 ( .A(a[3109]), .B(c3109), .Z(n9329) );
XOR U15550 ( .A(c3110), .B(n9330), .Z(c3111) );
ANDN U15551 ( .B(n9331), .A(n9332), .Z(n9330) );
XOR U15552 ( .A(c3110), .B(b[3110]), .Z(n9331) );
XNOR U15553 ( .A(b[3110]), .B(n9332), .Z(c[3110]) );
XNOR U15554 ( .A(a[3110]), .B(c3110), .Z(n9332) );
XOR U15555 ( .A(c3111), .B(n9333), .Z(c3112) );
ANDN U15556 ( .B(n9334), .A(n9335), .Z(n9333) );
XOR U15557 ( .A(c3111), .B(b[3111]), .Z(n9334) );
XNOR U15558 ( .A(b[3111]), .B(n9335), .Z(c[3111]) );
XNOR U15559 ( .A(a[3111]), .B(c3111), .Z(n9335) );
XOR U15560 ( .A(c3112), .B(n9336), .Z(c3113) );
ANDN U15561 ( .B(n9337), .A(n9338), .Z(n9336) );
XOR U15562 ( .A(c3112), .B(b[3112]), .Z(n9337) );
XNOR U15563 ( .A(b[3112]), .B(n9338), .Z(c[3112]) );
XNOR U15564 ( .A(a[3112]), .B(c3112), .Z(n9338) );
XOR U15565 ( .A(c3113), .B(n9339), .Z(c3114) );
ANDN U15566 ( .B(n9340), .A(n9341), .Z(n9339) );
XOR U15567 ( .A(c3113), .B(b[3113]), .Z(n9340) );
XNOR U15568 ( .A(b[3113]), .B(n9341), .Z(c[3113]) );
XNOR U15569 ( .A(a[3113]), .B(c3113), .Z(n9341) );
XOR U15570 ( .A(c3114), .B(n9342), .Z(c3115) );
ANDN U15571 ( .B(n9343), .A(n9344), .Z(n9342) );
XOR U15572 ( .A(c3114), .B(b[3114]), .Z(n9343) );
XNOR U15573 ( .A(b[3114]), .B(n9344), .Z(c[3114]) );
XNOR U15574 ( .A(a[3114]), .B(c3114), .Z(n9344) );
XOR U15575 ( .A(c3115), .B(n9345), .Z(c3116) );
ANDN U15576 ( .B(n9346), .A(n9347), .Z(n9345) );
XOR U15577 ( .A(c3115), .B(b[3115]), .Z(n9346) );
XNOR U15578 ( .A(b[3115]), .B(n9347), .Z(c[3115]) );
XNOR U15579 ( .A(a[3115]), .B(c3115), .Z(n9347) );
XOR U15580 ( .A(c3116), .B(n9348), .Z(c3117) );
ANDN U15581 ( .B(n9349), .A(n9350), .Z(n9348) );
XOR U15582 ( .A(c3116), .B(b[3116]), .Z(n9349) );
XNOR U15583 ( .A(b[3116]), .B(n9350), .Z(c[3116]) );
XNOR U15584 ( .A(a[3116]), .B(c3116), .Z(n9350) );
XOR U15585 ( .A(c3117), .B(n9351), .Z(c3118) );
ANDN U15586 ( .B(n9352), .A(n9353), .Z(n9351) );
XOR U15587 ( .A(c3117), .B(b[3117]), .Z(n9352) );
XNOR U15588 ( .A(b[3117]), .B(n9353), .Z(c[3117]) );
XNOR U15589 ( .A(a[3117]), .B(c3117), .Z(n9353) );
XOR U15590 ( .A(c3118), .B(n9354), .Z(c3119) );
ANDN U15591 ( .B(n9355), .A(n9356), .Z(n9354) );
XOR U15592 ( .A(c3118), .B(b[3118]), .Z(n9355) );
XNOR U15593 ( .A(b[3118]), .B(n9356), .Z(c[3118]) );
XNOR U15594 ( .A(a[3118]), .B(c3118), .Z(n9356) );
XOR U15595 ( .A(c3119), .B(n9357), .Z(c3120) );
ANDN U15596 ( .B(n9358), .A(n9359), .Z(n9357) );
XOR U15597 ( .A(c3119), .B(b[3119]), .Z(n9358) );
XNOR U15598 ( .A(b[3119]), .B(n9359), .Z(c[3119]) );
XNOR U15599 ( .A(a[3119]), .B(c3119), .Z(n9359) );
XOR U15600 ( .A(c3120), .B(n9360), .Z(c3121) );
ANDN U15601 ( .B(n9361), .A(n9362), .Z(n9360) );
XOR U15602 ( .A(c3120), .B(b[3120]), .Z(n9361) );
XNOR U15603 ( .A(b[3120]), .B(n9362), .Z(c[3120]) );
XNOR U15604 ( .A(a[3120]), .B(c3120), .Z(n9362) );
XOR U15605 ( .A(c3121), .B(n9363), .Z(c3122) );
ANDN U15606 ( .B(n9364), .A(n9365), .Z(n9363) );
XOR U15607 ( .A(c3121), .B(b[3121]), .Z(n9364) );
XNOR U15608 ( .A(b[3121]), .B(n9365), .Z(c[3121]) );
XNOR U15609 ( .A(a[3121]), .B(c3121), .Z(n9365) );
XOR U15610 ( .A(c3122), .B(n9366), .Z(c3123) );
ANDN U15611 ( .B(n9367), .A(n9368), .Z(n9366) );
XOR U15612 ( .A(c3122), .B(b[3122]), .Z(n9367) );
XNOR U15613 ( .A(b[3122]), .B(n9368), .Z(c[3122]) );
XNOR U15614 ( .A(a[3122]), .B(c3122), .Z(n9368) );
XOR U15615 ( .A(c3123), .B(n9369), .Z(c3124) );
ANDN U15616 ( .B(n9370), .A(n9371), .Z(n9369) );
XOR U15617 ( .A(c3123), .B(b[3123]), .Z(n9370) );
XNOR U15618 ( .A(b[3123]), .B(n9371), .Z(c[3123]) );
XNOR U15619 ( .A(a[3123]), .B(c3123), .Z(n9371) );
XOR U15620 ( .A(c3124), .B(n9372), .Z(c3125) );
ANDN U15621 ( .B(n9373), .A(n9374), .Z(n9372) );
XOR U15622 ( .A(c3124), .B(b[3124]), .Z(n9373) );
XNOR U15623 ( .A(b[3124]), .B(n9374), .Z(c[3124]) );
XNOR U15624 ( .A(a[3124]), .B(c3124), .Z(n9374) );
XOR U15625 ( .A(c3125), .B(n9375), .Z(c3126) );
ANDN U15626 ( .B(n9376), .A(n9377), .Z(n9375) );
XOR U15627 ( .A(c3125), .B(b[3125]), .Z(n9376) );
XNOR U15628 ( .A(b[3125]), .B(n9377), .Z(c[3125]) );
XNOR U15629 ( .A(a[3125]), .B(c3125), .Z(n9377) );
XOR U15630 ( .A(c3126), .B(n9378), .Z(c3127) );
ANDN U15631 ( .B(n9379), .A(n9380), .Z(n9378) );
XOR U15632 ( .A(c3126), .B(b[3126]), .Z(n9379) );
XNOR U15633 ( .A(b[3126]), .B(n9380), .Z(c[3126]) );
XNOR U15634 ( .A(a[3126]), .B(c3126), .Z(n9380) );
XOR U15635 ( .A(c3127), .B(n9381), .Z(c3128) );
ANDN U15636 ( .B(n9382), .A(n9383), .Z(n9381) );
XOR U15637 ( .A(c3127), .B(b[3127]), .Z(n9382) );
XNOR U15638 ( .A(b[3127]), .B(n9383), .Z(c[3127]) );
XNOR U15639 ( .A(a[3127]), .B(c3127), .Z(n9383) );
XOR U15640 ( .A(c3128), .B(n9384), .Z(c3129) );
ANDN U15641 ( .B(n9385), .A(n9386), .Z(n9384) );
XOR U15642 ( .A(c3128), .B(b[3128]), .Z(n9385) );
XNOR U15643 ( .A(b[3128]), .B(n9386), .Z(c[3128]) );
XNOR U15644 ( .A(a[3128]), .B(c3128), .Z(n9386) );
XOR U15645 ( .A(c3129), .B(n9387), .Z(c3130) );
ANDN U15646 ( .B(n9388), .A(n9389), .Z(n9387) );
XOR U15647 ( .A(c3129), .B(b[3129]), .Z(n9388) );
XNOR U15648 ( .A(b[3129]), .B(n9389), .Z(c[3129]) );
XNOR U15649 ( .A(a[3129]), .B(c3129), .Z(n9389) );
XOR U15650 ( .A(c3130), .B(n9390), .Z(c3131) );
ANDN U15651 ( .B(n9391), .A(n9392), .Z(n9390) );
XOR U15652 ( .A(c3130), .B(b[3130]), .Z(n9391) );
XNOR U15653 ( .A(b[3130]), .B(n9392), .Z(c[3130]) );
XNOR U15654 ( .A(a[3130]), .B(c3130), .Z(n9392) );
XOR U15655 ( .A(c3131), .B(n9393), .Z(c3132) );
ANDN U15656 ( .B(n9394), .A(n9395), .Z(n9393) );
XOR U15657 ( .A(c3131), .B(b[3131]), .Z(n9394) );
XNOR U15658 ( .A(b[3131]), .B(n9395), .Z(c[3131]) );
XNOR U15659 ( .A(a[3131]), .B(c3131), .Z(n9395) );
XOR U15660 ( .A(c3132), .B(n9396), .Z(c3133) );
ANDN U15661 ( .B(n9397), .A(n9398), .Z(n9396) );
XOR U15662 ( .A(c3132), .B(b[3132]), .Z(n9397) );
XNOR U15663 ( .A(b[3132]), .B(n9398), .Z(c[3132]) );
XNOR U15664 ( .A(a[3132]), .B(c3132), .Z(n9398) );
XOR U15665 ( .A(c3133), .B(n9399), .Z(c3134) );
ANDN U15666 ( .B(n9400), .A(n9401), .Z(n9399) );
XOR U15667 ( .A(c3133), .B(b[3133]), .Z(n9400) );
XNOR U15668 ( .A(b[3133]), .B(n9401), .Z(c[3133]) );
XNOR U15669 ( .A(a[3133]), .B(c3133), .Z(n9401) );
XOR U15670 ( .A(c3134), .B(n9402), .Z(c3135) );
ANDN U15671 ( .B(n9403), .A(n9404), .Z(n9402) );
XOR U15672 ( .A(c3134), .B(b[3134]), .Z(n9403) );
XNOR U15673 ( .A(b[3134]), .B(n9404), .Z(c[3134]) );
XNOR U15674 ( .A(a[3134]), .B(c3134), .Z(n9404) );
XOR U15675 ( .A(c3135), .B(n9405), .Z(c3136) );
ANDN U15676 ( .B(n9406), .A(n9407), .Z(n9405) );
XOR U15677 ( .A(c3135), .B(b[3135]), .Z(n9406) );
XNOR U15678 ( .A(b[3135]), .B(n9407), .Z(c[3135]) );
XNOR U15679 ( .A(a[3135]), .B(c3135), .Z(n9407) );
XOR U15680 ( .A(c3136), .B(n9408), .Z(c3137) );
ANDN U15681 ( .B(n9409), .A(n9410), .Z(n9408) );
XOR U15682 ( .A(c3136), .B(b[3136]), .Z(n9409) );
XNOR U15683 ( .A(b[3136]), .B(n9410), .Z(c[3136]) );
XNOR U15684 ( .A(a[3136]), .B(c3136), .Z(n9410) );
XOR U15685 ( .A(c3137), .B(n9411), .Z(c3138) );
ANDN U15686 ( .B(n9412), .A(n9413), .Z(n9411) );
XOR U15687 ( .A(c3137), .B(b[3137]), .Z(n9412) );
XNOR U15688 ( .A(b[3137]), .B(n9413), .Z(c[3137]) );
XNOR U15689 ( .A(a[3137]), .B(c3137), .Z(n9413) );
XOR U15690 ( .A(c3138), .B(n9414), .Z(c3139) );
ANDN U15691 ( .B(n9415), .A(n9416), .Z(n9414) );
XOR U15692 ( .A(c3138), .B(b[3138]), .Z(n9415) );
XNOR U15693 ( .A(b[3138]), .B(n9416), .Z(c[3138]) );
XNOR U15694 ( .A(a[3138]), .B(c3138), .Z(n9416) );
XOR U15695 ( .A(c3139), .B(n9417), .Z(c3140) );
ANDN U15696 ( .B(n9418), .A(n9419), .Z(n9417) );
XOR U15697 ( .A(c3139), .B(b[3139]), .Z(n9418) );
XNOR U15698 ( .A(b[3139]), .B(n9419), .Z(c[3139]) );
XNOR U15699 ( .A(a[3139]), .B(c3139), .Z(n9419) );
XOR U15700 ( .A(c3140), .B(n9420), .Z(c3141) );
ANDN U15701 ( .B(n9421), .A(n9422), .Z(n9420) );
XOR U15702 ( .A(c3140), .B(b[3140]), .Z(n9421) );
XNOR U15703 ( .A(b[3140]), .B(n9422), .Z(c[3140]) );
XNOR U15704 ( .A(a[3140]), .B(c3140), .Z(n9422) );
XOR U15705 ( .A(c3141), .B(n9423), .Z(c3142) );
ANDN U15706 ( .B(n9424), .A(n9425), .Z(n9423) );
XOR U15707 ( .A(c3141), .B(b[3141]), .Z(n9424) );
XNOR U15708 ( .A(b[3141]), .B(n9425), .Z(c[3141]) );
XNOR U15709 ( .A(a[3141]), .B(c3141), .Z(n9425) );
XOR U15710 ( .A(c3142), .B(n9426), .Z(c3143) );
ANDN U15711 ( .B(n9427), .A(n9428), .Z(n9426) );
XOR U15712 ( .A(c3142), .B(b[3142]), .Z(n9427) );
XNOR U15713 ( .A(b[3142]), .B(n9428), .Z(c[3142]) );
XNOR U15714 ( .A(a[3142]), .B(c3142), .Z(n9428) );
XOR U15715 ( .A(c3143), .B(n9429), .Z(c3144) );
ANDN U15716 ( .B(n9430), .A(n9431), .Z(n9429) );
XOR U15717 ( .A(c3143), .B(b[3143]), .Z(n9430) );
XNOR U15718 ( .A(b[3143]), .B(n9431), .Z(c[3143]) );
XNOR U15719 ( .A(a[3143]), .B(c3143), .Z(n9431) );
XOR U15720 ( .A(c3144), .B(n9432), .Z(c3145) );
ANDN U15721 ( .B(n9433), .A(n9434), .Z(n9432) );
XOR U15722 ( .A(c3144), .B(b[3144]), .Z(n9433) );
XNOR U15723 ( .A(b[3144]), .B(n9434), .Z(c[3144]) );
XNOR U15724 ( .A(a[3144]), .B(c3144), .Z(n9434) );
XOR U15725 ( .A(c3145), .B(n9435), .Z(c3146) );
ANDN U15726 ( .B(n9436), .A(n9437), .Z(n9435) );
XOR U15727 ( .A(c3145), .B(b[3145]), .Z(n9436) );
XNOR U15728 ( .A(b[3145]), .B(n9437), .Z(c[3145]) );
XNOR U15729 ( .A(a[3145]), .B(c3145), .Z(n9437) );
XOR U15730 ( .A(c3146), .B(n9438), .Z(c3147) );
ANDN U15731 ( .B(n9439), .A(n9440), .Z(n9438) );
XOR U15732 ( .A(c3146), .B(b[3146]), .Z(n9439) );
XNOR U15733 ( .A(b[3146]), .B(n9440), .Z(c[3146]) );
XNOR U15734 ( .A(a[3146]), .B(c3146), .Z(n9440) );
XOR U15735 ( .A(c3147), .B(n9441), .Z(c3148) );
ANDN U15736 ( .B(n9442), .A(n9443), .Z(n9441) );
XOR U15737 ( .A(c3147), .B(b[3147]), .Z(n9442) );
XNOR U15738 ( .A(b[3147]), .B(n9443), .Z(c[3147]) );
XNOR U15739 ( .A(a[3147]), .B(c3147), .Z(n9443) );
XOR U15740 ( .A(c3148), .B(n9444), .Z(c3149) );
ANDN U15741 ( .B(n9445), .A(n9446), .Z(n9444) );
XOR U15742 ( .A(c3148), .B(b[3148]), .Z(n9445) );
XNOR U15743 ( .A(b[3148]), .B(n9446), .Z(c[3148]) );
XNOR U15744 ( .A(a[3148]), .B(c3148), .Z(n9446) );
XOR U15745 ( .A(c3149), .B(n9447), .Z(c3150) );
ANDN U15746 ( .B(n9448), .A(n9449), .Z(n9447) );
XOR U15747 ( .A(c3149), .B(b[3149]), .Z(n9448) );
XNOR U15748 ( .A(b[3149]), .B(n9449), .Z(c[3149]) );
XNOR U15749 ( .A(a[3149]), .B(c3149), .Z(n9449) );
XOR U15750 ( .A(c3150), .B(n9450), .Z(c3151) );
ANDN U15751 ( .B(n9451), .A(n9452), .Z(n9450) );
XOR U15752 ( .A(c3150), .B(b[3150]), .Z(n9451) );
XNOR U15753 ( .A(b[3150]), .B(n9452), .Z(c[3150]) );
XNOR U15754 ( .A(a[3150]), .B(c3150), .Z(n9452) );
XOR U15755 ( .A(c3151), .B(n9453), .Z(c3152) );
ANDN U15756 ( .B(n9454), .A(n9455), .Z(n9453) );
XOR U15757 ( .A(c3151), .B(b[3151]), .Z(n9454) );
XNOR U15758 ( .A(b[3151]), .B(n9455), .Z(c[3151]) );
XNOR U15759 ( .A(a[3151]), .B(c3151), .Z(n9455) );
XOR U15760 ( .A(c3152), .B(n9456), .Z(c3153) );
ANDN U15761 ( .B(n9457), .A(n9458), .Z(n9456) );
XOR U15762 ( .A(c3152), .B(b[3152]), .Z(n9457) );
XNOR U15763 ( .A(b[3152]), .B(n9458), .Z(c[3152]) );
XNOR U15764 ( .A(a[3152]), .B(c3152), .Z(n9458) );
XOR U15765 ( .A(c3153), .B(n9459), .Z(c3154) );
ANDN U15766 ( .B(n9460), .A(n9461), .Z(n9459) );
XOR U15767 ( .A(c3153), .B(b[3153]), .Z(n9460) );
XNOR U15768 ( .A(b[3153]), .B(n9461), .Z(c[3153]) );
XNOR U15769 ( .A(a[3153]), .B(c3153), .Z(n9461) );
XOR U15770 ( .A(c3154), .B(n9462), .Z(c3155) );
ANDN U15771 ( .B(n9463), .A(n9464), .Z(n9462) );
XOR U15772 ( .A(c3154), .B(b[3154]), .Z(n9463) );
XNOR U15773 ( .A(b[3154]), .B(n9464), .Z(c[3154]) );
XNOR U15774 ( .A(a[3154]), .B(c3154), .Z(n9464) );
XOR U15775 ( .A(c3155), .B(n9465), .Z(c3156) );
ANDN U15776 ( .B(n9466), .A(n9467), .Z(n9465) );
XOR U15777 ( .A(c3155), .B(b[3155]), .Z(n9466) );
XNOR U15778 ( .A(b[3155]), .B(n9467), .Z(c[3155]) );
XNOR U15779 ( .A(a[3155]), .B(c3155), .Z(n9467) );
XOR U15780 ( .A(c3156), .B(n9468), .Z(c3157) );
ANDN U15781 ( .B(n9469), .A(n9470), .Z(n9468) );
XOR U15782 ( .A(c3156), .B(b[3156]), .Z(n9469) );
XNOR U15783 ( .A(b[3156]), .B(n9470), .Z(c[3156]) );
XNOR U15784 ( .A(a[3156]), .B(c3156), .Z(n9470) );
XOR U15785 ( .A(c3157), .B(n9471), .Z(c3158) );
ANDN U15786 ( .B(n9472), .A(n9473), .Z(n9471) );
XOR U15787 ( .A(c3157), .B(b[3157]), .Z(n9472) );
XNOR U15788 ( .A(b[3157]), .B(n9473), .Z(c[3157]) );
XNOR U15789 ( .A(a[3157]), .B(c3157), .Z(n9473) );
XOR U15790 ( .A(c3158), .B(n9474), .Z(c3159) );
ANDN U15791 ( .B(n9475), .A(n9476), .Z(n9474) );
XOR U15792 ( .A(c3158), .B(b[3158]), .Z(n9475) );
XNOR U15793 ( .A(b[3158]), .B(n9476), .Z(c[3158]) );
XNOR U15794 ( .A(a[3158]), .B(c3158), .Z(n9476) );
XOR U15795 ( .A(c3159), .B(n9477), .Z(c3160) );
ANDN U15796 ( .B(n9478), .A(n9479), .Z(n9477) );
XOR U15797 ( .A(c3159), .B(b[3159]), .Z(n9478) );
XNOR U15798 ( .A(b[3159]), .B(n9479), .Z(c[3159]) );
XNOR U15799 ( .A(a[3159]), .B(c3159), .Z(n9479) );
XOR U15800 ( .A(c3160), .B(n9480), .Z(c3161) );
ANDN U15801 ( .B(n9481), .A(n9482), .Z(n9480) );
XOR U15802 ( .A(c3160), .B(b[3160]), .Z(n9481) );
XNOR U15803 ( .A(b[3160]), .B(n9482), .Z(c[3160]) );
XNOR U15804 ( .A(a[3160]), .B(c3160), .Z(n9482) );
XOR U15805 ( .A(c3161), .B(n9483), .Z(c3162) );
ANDN U15806 ( .B(n9484), .A(n9485), .Z(n9483) );
XOR U15807 ( .A(c3161), .B(b[3161]), .Z(n9484) );
XNOR U15808 ( .A(b[3161]), .B(n9485), .Z(c[3161]) );
XNOR U15809 ( .A(a[3161]), .B(c3161), .Z(n9485) );
XOR U15810 ( .A(c3162), .B(n9486), .Z(c3163) );
ANDN U15811 ( .B(n9487), .A(n9488), .Z(n9486) );
XOR U15812 ( .A(c3162), .B(b[3162]), .Z(n9487) );
XNOR U15813 ( .A(b[3162]), .B(n9488), .Z(c[3162]) );
XNOR U15814 ( .A(a[3162]), .B(c3162), .Z(n9488) );
XOR U15815 ( .A(c3163), .B(n9489), .Z(c3164) );
ANDN U15816 ( .B(n9490), .A(n9491), .Z(n9489) );
XOR U15817 ( .A(c3163), .B(b[3163]), .Z(n9490) );
XNOR U15818 ( .A(b[3163]), .B(n9491), .Z(c[3163]) );
XNOR U15819 ( .A(a[3163]), .B(c3163), .Z(n9491) );
XOR U15820 ( .A(c3164), .B(n9492), .Z(c3165) );
ANDN U15821 ( .B(n9493), .A(n9494), .Z(n9492) );
XOR U15822 ( .A(c3164), .B(b[3164]), .Z(n9493) );
XNOR U15823 ( .A(b[3164]), .B(n9494), .Z(c[3164]) );
XNOR U15824 ( .A(a[3164]), .B(c3164), .Z(n9494) );
XOR U15825 ( .A(c3165), .B(n9495), .Z(c3166) );
ANDN U15826 ( .B(n9496), .A(n9497), .Z(n9495) );
XOR U15827 ( .A(c3165), .B(b[3165]), .Z(n9496) );
XNOR U15828 ( .A(b[3165]), .B(n9497), .Z(c[3165]) );
XNOR U15829 ( .A(a[3165]), .B(c3165), .Z(n9497) );
XOR U15830 ( .A(c3166), .B(n9498), .Z(c3167) );
ANDN U15831 ( .B(n9499), .A(n9500), .Z(n9498) );
XOR U15832 ( .A(c3166), .B(b[3166]), .Z(n9499) );
XNOR U15833 ( .A(b[3166]), .B(n9500), .Z(c[3166]) );
XNOR U15834 ( .A(a[3166]), .B(c3166), .Z(n9500) );
XOR U15835 ( .A(c3167), .B(n9501), .Z(c3168) );
ANDN U15836 ( .B(n9502), .A(n9503), .Z(n9501) );
XOR U15837 ( .A(c3167), .B(b[3167]), .Z(n9502) );
XNOR U15838 ( .A(b[3167]), .B(n9503), .Z(c[3167]) );
XNOR U15839 ( .A(a[3167]), .B(c3167), .Z(n9503) );
XOR U15840 ( .A(c3168), .B(n9504), .Z(c3169) );
ANDN U15841 ( .B(n9505), .A(n9506), .Z(n9504) );
XOR U15842 ( .A(c3168), .B(b[3168]), .Z(n9505) );
XNOR U15843 ( .A(b[3168]), .B(n9506), .Z(c[3168]) );
XNOR U15844 ( .A(a[3168]), .B(c3168), .Z(n9506) );
XOR U15845 ( .A(c3169), .B(n9507), .Z(c3170) );
ANDN U15846 ( .B(n9508), .A(n9509), .Z(n9507) );
XOR U15847 ( .A(c3169), .B(b[3169]), .Z(n9508) );
XNOR U15848 ( .A(b[3169]), .B(n9509), .Z(c[3169]) );
XNOR U15849 ( .A(a[3169]), .B(c3169), .Z(n9509) );
XOR U15850 ( .A(c3170), .B(n9510), .Z(c3171) );
ANDN U15851 ( .B(n9511), .A(n9512), .Z(n9510) );
XOR U15852 ( .A(c3170), .B(b[3170]), .Z(n9511) );
XNOR U15853 ( .A(b[3170]), .B(n9512), .Z(c[3170]) );
XNOR U15854 ( .A(a[3170]), .B(c3170), .Z(n9512) );
XOR U15855 ( .A(c3171), .B(n9513), .Z(c3172) );
ANDN U15856 ( .B(n9514), .A(n9515), .Z(n9513) );
XOR U15857 ( .A(c3171), .B(b[3171]), .Z(n9514) );
XNOR U15858 ( .A(b[3171]), .B(n9515), .Z(c[3171]) );
XNOR U15859 ( .A(a[3171]), .B(c3171), .Z(n9515) );
XOR U15860 ( .A(c3172), .B(n9516), .Z(c3173) );
ANDN U15861 ( .B(n9517), .A(n9518), .Z(n9516) );
XOR U15862 ( .A(c3172), .B(b[3172]), .Z(n9517) );
XNOR U15863 ( .A(b[3172]), .B(n9518), .Z(c[3172]) );
XNOR U15864 ( .A(a[3172]), .B(c3172), .Z(n9518) );
XOR U15865 ( .A(c3173), .B(n9519), .Z(c3174) );
ANDN U15866 ( .B(n9520), .A(n9521), .Z(n9519) );
XOR U15867 ( .A(c3173), .B(b[3173]), .Z(n9520) );
XNOR U15868 ( .A(b[3173]), .B(n9521), .Z(c[3173]) );
XNOR U15869 ( .A(a[3173]), .B(c3173), .Z(n9521) );
XOR U15870 ( .A(c3174), .B(n9522), .Z(c3175) );
ANDN U15871 ( .B(n9523), .A(n9524), .Z(n9522) );
XOR U15872 ( .A(c3174), .B(b[3174]), .Z(n9523) );
XNOR U15873 ( .A(b[3174]), .B(n9524), .Z(c[3174]) );
XNOR U15874 ( .A(a[3174]), .B(c3174), .Z(n9524) );
XOR U15875 ( .A(c3175), .B(n9525), .Z(c3176) );
ANDN U15876 ( .B(n9526), .A(n9527), .Z(n9525) );
XOR U15877 ( .A(c3175), .B(b[3175]), .Z(n9526) );
XNOR U15878 ( .A(b[3175]), .B(n9527), .Z(c[3175]) );
XNOR U15879 ( .A(a[3175]), .B(c3175), .Z(n9527) );
XOR U15880 ( .A(c3176), .B(n9528), .Z(c3177) );
ANDN U15881 ( .B(n9529), .A(n9530), .Z(n9528) );
XOR U15882 ( .A(c3176), .B(b[3176]), .Z(n9529) );
XNOR U15883 ( .A(b[3176]), .B(n9530), .Z(c[3176]) );
XNOR U15884 ( .A(a[3176]), .B(c3176), .Z(n9530) );
XOR U15885 ( .A(c3177), .B(n9531), .Z(c3178) );
ANDN U15886 ( .B(n9532), .A(n9533), .Z(n9531) );
XOR U15887 ( .A(c3177), .B(b[3177]), .Z(n9532) );
XNOR U15888 ( .A(b[3177]), .B(n9533), .Z(c[3177]) );
XNOR U15889 ( .A(a[3177]), .B(c3177), .Z(n9533) );
XOR U15890 ( .A(c3178), .B(n9534), .Z(c3179) );
ANDN U15891 ( .B(n9535), .A(n9536), .Z(n9534) );
XOR U15892 ( .A(c3178), .B(b[3178]), .Z(n9535) );
XNOR U15893 ( .A(b[3178]), .B(n9536), .Z(c[3178]) );
XNOR U15894 ( .A(a[3178]), .B(c3178), .Z(n9536) );
XOR U15895 ( .A(c3179), .B(n9537), .Z(c3180) );
ANDN U15896 ( .B(n9538), .A(n9539), .Z(n9537) );
XOR U15897 ( .A(c3179), .B(b[3179]), .Z(n9538) );
XNOR U15898 ( .A(b[3179]), .B(n9539), .Z(c[3179]) );
XNOR U15899 ( .A(a[3179]), .B(c3179), .Z(n9539) );
XOR U15900 ( .A(c3180), .B(n9540), .Z(c3181) );
ANDN U15901 ( .B(n9541), .A(n9542), .Z(n9540) );
XOR U15902 ( .A(c3180), .B(b[3180]), .Z(n9541) );
XNOR U15903 ( .A(b[3180]), .B(n9542), .Z(c[3180]) );
XNOR U15904 ( .A(a[3180]), .B(c3180), .Z(n9542) );
XOR U15905 ( .A(c3181), .B(n9543), .Z(c3182) );
ANDN U15906 ( .B(n9544), .A(n9545), .Z(n9543) );
XOR U15907 ( .A(c3181), .B(b[3181]), .Z(n9544) );
XNOR U15908 ( .A(b[3181]), .B(n9545), .Z(c[3181]) );
XNOR U15909 ( .A(a[3181]), .B(c3181), .Z(n9545) );
XOR U15910 ( .A(c3182), .B(n9546), .Z(c3183) );
ANDN U15911 ( .B(n9547), .A(n9548), .Z(n9546) );
XOR U15912 ( .A(c3182), .B(b[3182]), .Z(n9547) );
XNOR U15913 ( .A(b[3182]), .B(n9548), .Z(c[3182]) );
XNOR U15914 ( .A(a[3182]), .B(c3182), .Z(n9548) );
XOR U15915 ( .A(c3183), .B(n9549), .Z(c3184) );
ANDN U15916 ( .B(n9550), .A(n9551), .Z(n9549) );
XOR U15917 ( .A(c3183), .B(b[3183]), .Z(n9550) );
XNOR U15918 ( .A(b[3183]), .B(n9551), .Z(c[3183]) );
XNOR U15919 ( .A(a[3183]), .B(c3183), .Z(n9551) );
XOR U15920 ( .A(c3184), .B(n9552), .Z(c3185) );
ANDN U15921 ( .B(n9553), .A(n9554), .Z(n9552) );
XOR U15922 ( .A(c3184), .B(b[3184]), .Z(n9553) );
XNOR U15923 ( .A(b[3184]), .B(n9554), .Z(c[3184]) );
XNOR U15924 ( .A(a[3184]), .B(c3184), .Z(n9554) );
XOR U15925 ( .A(c3185), .B(n9555), .Z(c3186) );
ANDN U15926 ( .B(n9556), .A(n9557), .Z(n9555) );
XOR U15927 ( .A(c3185), .B(b[3185]), .Z(n9556) );
XNOR U15928 ( .A(b[3185]), .B(n9557), .Z(c[3185]) );
XNOR U15929 ( .A(a[3185]), .B(c3185), .Z(n9557) );
XOR U15930 ( .A(c3186), .B(n9558), .Z(c3187) );
ANDN U15931 ( .B(n9559), .A(n9560), .Z(n9558) );
XOR U15932 ( .A(c3186), .B(b[3186]), .Z(n9559) );
XNOR U15933 ( .A(b[3186]), .B(n9560), .Z(c[3186]) );
XNOR U15934 ( .A(a[3186]), .B(c3186), .Z(n9560) );
XOR U15935 ( .A(c3187), .B(n9561), .Z(c3188) );
ANDN U15936 ( .B(n9562), .A(n9563), .Z(n9561) );
XOR U15937 ( .A(c3187), .B(b[3187]), .Z(n9562) );
XNOR U15938 ( .A(b[3187]), .B(n9563), .Z(c[3187]) );
XNOR U15939 ( .A(a[3187]), .B(c3187), .Z(n9563) );
XOR U15940 ( .A(c3188), .B(n9564), .Z(c3189) );
ANDN U15941 ( .B(n9565), .A(n9566), .Z(n9564) );
XOR U15942 ( .A(c3188), .B(b[3188]), .Z(n9565) );
XNOR U15943 ( .A(b[3188]), .B(n9566), .Z(c[3188]) );
XNOR U15944 ( .A(a[3188]), .B(c3188), .Z(n9566) );
XOR U15945 ( .A(c3189), .B(n9567), .Z(c3190) );
ANDN U15946 ( .B(n9568), .A(n9569), .Z(n9567) );
XOR U15947 ( .A(c3189), .B(b[3189]), .Z(n9568) );
XNOR U15948 ( .A(b[3189]), .B(n9569), .Z(c[3189]) );
XNOR U15949 ( .A(a[3189]), .B(c3189), .Z(n9569) );
XOR U15950 ( .A(c3190), .B(n9570), .Z(c3191) );
ANDN U15951 ( .B(n9571), .A(n9572), .Z(n9570) );
XOR U15952 ( .A(c3190), .B(b[3190]), .Z(n9571) );
XNOR U15953 ( .A(b[3190]), .B(n9572), .Z(c[3190]) );
XNOR U15954 ( .A(a[3190]), .B(c3190), .Z(n9572) );
XOR U15955 ( .A(c3191), .B(n9573), .Z(c3192) );
ANDN U15956 ( .B(n9574), .A(n9575), .Z(n9573) );
XOR U15957 ( .A(c3191), .B(b[3191]), .Z(n9574) );
XNOR U15958 ( .A(b[3191]), .B(n9575), .Z(c[3191]) );
XNOR U15959 ( .A(a[3191]), .B(c3191), .Z(n9575) );
XOR U15960 ( .A(c3192), .B(n9576), .Z(c3193) );
ANDN U15961 ( .B(n9577), .A(n9578), .Z(n9576) );
XOR U15962 ( .A(c3192), .B(b[3192]), .Z(n9577) );
XNOR U15963 ( .A(b[3192]), .B(n9578), .Z(c[3192]) );
XNOR U15964 ( .A(a[3192]), .B(c3192), .Z(n9578) );
XOR U15965 ( .A(c3193), .B(n9579), .Z(c3194) );
ANDN U15966 ( .B(n9580), .A(n9581), .Z(n9579) );
XOR U15967 ( .A(c3193), .B(b[3193]), .Z(n9580) );
XNOR U15968 ( .A(b[3193]), .B(n9581), .Z(c[3193]) );
XNOR U15969 ( .A(a[3193]), .B(c3193), .Z(n9581) );
XOR U15970 ( .A(c3194), .B(n9582), .Z(c3195) );
ANDN U15971 ( .B(n9583), .A(n9584), .Z(n9582) );
XOR U15972 ( .A(c3194), .B(b[3194]), .Z(n9583) );
XNOR U15973 ( .A(b[3194]), .B(n9584), .Z(c[3194]) );
XNOR U15974 ( .A(a[3194]), .B(c3194), .Z(n9584) );
XOR U15975 ( .A(c3195), .B(n9585), .Z(c3196) );
ANDN U15976 ( .B(n9586), .A(n9587), .Z(n9585) );
XOR U15977 ( .A(c3195), .B(b[3195]), .Z(n9586) );
XNOR U15978 ( .A(b[3195]), .B(n9587), .Z(c[3195]) );
XNOR U15979 ( .A(a[3195]), .B(c3195), .Z(n9587) );
XOR U15980 ( .A(c3196), .B(n9588), .Z(c3197) );
ANDN U15981 ( .B(n9589), .A(n9590), .Z(n9588) );
XOR U15982 ( .A(c3196), .B(b[3196]), .Z(n9589) );
XNOR U15983 ( .A(b[3196]), .B(n9590), .Z(c[3196]) );
XNOR U15984 ( .A(a[3196]), .B(c3196), .Z(n9590) );
XOR U15985 ( .A(c3197), .B(n9591), .Z(c3198) );
ANDN U15986 ( .B(n9592), .A(n9593), .Z(n9591) );
XOR U15987 ( .A(c3197), .B(b[3197]), .Z(n9592) );
XNOR U15988 ( .A(b[3197]), .B(n9593), .Z(c[3197]) );
XNOR U15989 ( .A(a[3197]), .B(c3197), .Z(n9593) );
XOR U15990 ( .A(c3198), .B(n9594), .Z(c3199) );
ANDN U15991 ( .B(n9595), .A(n9596), .Z(n9594) );
XOR U15992 ( .A(c3198), .B(b[3198]), .Z(n9595) );
XNOR U15993 ( .A(b[3198]), .B(n9596), .Z(c[3198]) );
XNOR U15994 ( .A(a[3198]), .B(c3198), .Z(n9596) );
XOR U15995 ( .A(c3199), .B(n9597), .Z(c3200) );
ANDN U15996 ( .B(n9598), .A(n9599), .Z(n9597) );
XOR U15997 ( .A(c3199), .B(b[3199]), .Z(n9598) );
XNOR U15998 ( .A(b[3199]), .B(n9599), .Z(c[3199]) );
XNOR U15999 ( .A(a[3199]), .B(c3199), .Z(n9599) );
XOR U16000 ( .A(c3200), .B(n9600), .Z(c3201) );
ANDN U16001 ( .B(n9601), .A(n9602), .Z(n9600) );
XOR U16002 ( .A(c3200), .B(b[3200]), .Z(n9601) );
XNOR U16003 ( .A(b[3200]), .B(n9602), .Z(c[3200]) );
XNOR U16004 ( .A(a[3200]), .B(c3200), .Z(n9602) );
XOR U16005 ( .A(c3201), .B(n9603), .Z(c3202) );
ANDN U16006 ( .B(n9604), .A(n9605), .Z(n9603) );
XOR U16007 ( .A(c3201), .B(b[3201]), .Z(n9604) );
XNOR U16008 ( .A(b[3201]), .B(n9605), .Z(c[3201]) );
XNOR U16009 ( .A(a[3201]), .B(c3201), .Z(n9605) );
XOR U16010 ( .A(c3202), .B(n9606), .Z(c3203) );
ANDN U16011 ( .B(n9607), .A(n9608), .Z(n9606) );
XOR U16012 ( .A(c3202), .B(b[3202]), .Z(n9607) );
XNOR U16013 ( .A(b[3202]), .B(n9608), .Z(c[3202]) );
XNOR U16014 ( .A(a[3202]), .B(c3202), .Z(n9608) );
XOR U16015 ( .A(c3203), .B(n9609), .Z(c3204) );
ANDN U16016 ( .B(n9610), .A(n9611), .Z(n9609) );
XOR U16017 ( .A(c3203), .B(b[3203]), .Z(n9610) );
XNOR U16018 ( .A(b[3203]), .B(n9611), .Z(c[3203]) );
XNOR U16019 ( .A(a[3203]), .B(c3203), .Z(n9611) );
XOR U16020 ( .A(c3204), .B(n9612), .Z(c3205) );
ANDN U16021 ( .B(n9613), .A(n9614), .Z(n9612) );
XOR U16022 ( .A(c3204), .B(b[3204]), .Z(n9613) );
XNOR U16023 ( .A(b[3204]), .B(n9614), .Z(c[3204]) );
XNOR U16024 ( .A(a[3204]), .B(c3204), .Z(n9614) );
XOR U16025 ( .A(c3205), .B(n9615), .Z(c3206) );
ANDN U16026 ( .B(n9616), .A(n9617), .Z(n9615) );
XOR U16027 ( .A(c3205), .B(b[3205]), .Z(n9616) );
XNOR U16028 ( .A(b[3205]), .B(n9617), .Z(c[3205]) );
XNOR U16029 ( .A(a[3205]), .B(c3205), .Z(n9617) );
XOR U16030 ( .A(c3206), .B(n9618), .Z(c3207) );
ANDN U16031 ( .B(n9619), .A(n9620), .Z(n9618) );
XOR U16032 ( .A(c3206), .B(b[3206]), .Z(n9619) );
XNOR U16033 ( .A(b[3206]), .B(n9620), .Z(c[3206]) );
XNOR U16034 ( .A(a[3206]), .B(c3206), .Z(n9620) );
XOR U16035 ( .A(c3207), .B(n9621), .Z(c3208) );
ANDN U16036 ( .B(n9622), .A(n9623), .Z(n9621) );
XOR U16037 ( .A(c3207), .B(b[3207]), .Z(n9622) );
XNOR U16038 ( .A(b[3207]), .B(n9623), .Z(c[3207]) );
XNOR U16039 ( .A(a[3207]), .B(c3207), .Z(n9623) );
XOR U16040 ( .A(c3208), .B(n9624), .Z(c3209) );
ANDN U16041 ( .B(n9625), .A(n9626), .Z(n9624) );
XOR U16042 ( .A(c3208), .B(b[3208]), .Z(n9625) );
XNOR U16043 ( .A(b[3208]), .B(n9626), .Z(c[3208]) );
XNOR U16044 ( .A(a[3208]), .B(c3208), .Z(n9626) );
XOR U16045 ( .A(c3209), .B(n9627), .Z(c3210) );
ANDN U16046 ( .B(n9628), .A(n9629), .Z(n9627) );
XOR U16047 ( .A(c3209), .B(b[3209]), .Z(n9628) );
XNOR U16048 ( .A(b[3209]), .B(n9629), .Z(c[3209]) );
XNOR U16049 ( .A(a[3209]), .B(c3209), .Z(n9629) );
XOR U16050 ( .A(c3210), .B(n9630), .Z(c3211) );
ANDN U16051 ( .B(n9631), .A(n9632), .Z(n9630) );
XOR U16052 ( .A(c3210), .B(b[3210]), .Z(n9631) );
XNOR U16053 ( .A(b[3210]), .B(n9632), .Z(c[3210]) );
XNOR U16054 ( .A(a[3210]), .B(c3210), .Z(n9632) );
XOR U16055 ( .A(c3211), .B(n9633), .Z(c3212) );
ANDN U16056 ( .B(n9634), .A(n9635), .Z(n9633) );
XOR U16057 ( .A(c3211), .B(b[3211]), .Z(n9634) );
XNOR U16058 ( .A(b[3211]), .B(n9635), .Z(c[3211]) );
XNOR U16059 ( .A(a[3211]), .B(c3211), .Z(n9635) );
XOR U16060 ( .A(c3212), .B(n9636), .Z(c3213) );
ANDN U16061 ( .B(n9637), .A(n9638), .Z(n9636) );
XOR U16062 ( .A(c3212), .B(b[3212]), .Z(n9637) );
XNOR U16063 ( .A(b[3212]), .B(n9638), .Z(c[3212]) );
XNOR U16064 ( .A(a[3212]), .B(c3212), .Z(n9638) );
XOR U16065 ( .A(c3213), .B(n9639), .Z(c3214) );
ANDN U16066 ( .B(n9640), .A(n9641), .Z(n9639) );
XOR U16067 ( .A(c3213), .B(b[3213]), .Z(n9640) );
XNOR U16068 ( .A(b[3213]), .B(n9641), .Z(c[3213]) );
XNOR U16069 ( .A(a[3213]), .B(c3213), .Z(n9641) );
XOR U16070 ( .A(c3214), .B(n9642), .Z(c3215) );
ANDN U16071 ( .B(n9643), .A(n9644), .Z(n9642) );
XOR U16072 ( .A(c3214), .B(b[3214]), .Z(n9643) );
XNOR U16073 ( .A(b[3214]), .B(n9644), .Z(c[3214]) );
XNOR U16074 ( .A(a[3214]), .B(c3214), .Z(n9644) );
XOR U16075 ( .A(c3215), .B(n9645), .Z(c3216) );
ANDN U16076 ( .B(n9646), .A(n9647), .Z(n9645) );
XOR U16077 ( .A(c3215), .B(b[3215]), .Z(n9646) );
XNOR U16078 ( .A(b[3215]), .B(n9647), .Z(c[3215]) );
XNOR U16079 ( .A(a[3215]), .B(c3215), .Z(n9647) );
XOR U16080 ( .A(c3216), .B(n9648), .Z(c3217) );
ANDN U16081 ( .B(n9649), .A(n9650), .Z(n9648) );
XOR U16082 ( .A(c3216), .B(b[3216]), .Z(n9649) );
XNOR U16083 ( .A(b[3216]), .B(n9650), .Z(c[3216]) );
XNOR U16084 ( .A(a[3216]), .B(c3216), .Z(n9650) );
XOR U16085 ( .A(c3217), .B(n9651), .Z(c3218) );
ANDN U16086 ( .B(n9652), .A(n9653), .Z(n9651) );
XOR U16087 ( .A(c3217), .B(b[3217]), .Z(n9652) );
XNOR U16088 ( .A(b[3217]), .B(n9653), .Z(c[3217]) );
XNOR U16089 ( .A(a[3217]), .B(c3217), .Z(n9653) );
XOR U16090 ( .A(c3218), .B(n9654), .Z(c3219) );
ANDN U16091 ( .B(n9655), .A(n9656), .Z(n9654) );
XOR U16092 ( .A(c3218), .B(b[3218]), .Z(n9655) );
XNOR U16093 ( .A(b[3218]), .B(n9656), .Z(c[3218]) );
XNOR U16094 ( .A(a[3218]), .B(c3218), .Z(n9656) );
XOR U16095 ( .A(c3219), .B(n9657), .Z(c3220) );
ANDN U16096 ( .B(n9658), .A(n9659), .Z(n9657) );
XOR U16097 ( .A(c3219), .B(b[3219]), .Z(n9658) );
XNOR U16098 ( .A(b[3219]), .B(n9659), .Z(c[3219]) );
XNOR U16099 ( .A(a[3219]), .B(c3219), .Z(n9659) );
XOR U16100 ( .A(c3220), .B(n9660), .Z(c3221) );
ANDN U16101 ( .B(n9661), .A(n9662), .Z(n9660) );
XOR U16102 ( .A(c3220), .B(b[3220]), .Z(n9661) );
XNOR U16103 ( .A(b[3220]), .B(n9662), .Z(c[3220]) );
XNOR U16104 ( .A(a[3220]), .B(c3220), .Z(n9662) );
XOR U16105 ( .A(c3221), .B(n9663), .Z(c3222) );
ANDN U16106 ( .B(n9664), .A(n9665), .Z(n9663) );
XOR U16107 ( .A(c3221), .B(b[3221]), .Z(n9664) );
XNOR U16108 ( .A(b[3221]), .B(n9665), .Z(c[3221]) );
XNOR U16109 ( .A(a[3221]), .B(c3221), .Z(n9665) );
XOR U16110 ( .A(c3222), .B(n9666), .Z(c3223) );
ANDN U16111 ( .B(n9667), .A(n9668), .Z(n9666) );
XOR U16112 ( .A(c3222), .B(b[3222]), .Z(n9667) );
XNOR U16113 ( .A(b[3222]), .B(n9668), .Z(c[3222]) );
XNOR U16114 ( .A(a[3222]), .B(c3222), .Z(n9668) );
XOR U16115 ( .A(c3223), .B(n9669), .Z(c3224) );
ANDN U16116 ( .B(n9670), .A(n9671), .Z(n9669) );
XOR U16117 ( .A(c3223), .B(b[3223]), .Z(n9670) );
XNOR U16118 ( .A(b[3223]), .B(n9671), .Z(c[3223]) );
XNOR U16119 ( .A(a[3223]), .B(c3223), .Z(n9671) );
XOR U16120 ( .A(c3224), .B(n9672), .Z(c3225) );
ANDN U16121 ( .B(n9673), .A(n9674), .Z(n9672) );
XOR U16122 ( .A(c3224), .B(b[3224]), .Z(n9673) );
XNOR U16123 ( .A(b[3224]), .B(n9674), .Z(c[3224]) );
XNOR U16124 ( .A(a[3224]), .B(c3224), .Z(n9674) );
XOR U16125 ( .A(c3225), .B(n9675), .Z(c3226) );
ANDN U16126 ( .B(n9676), .A(n9677), .Z(n9675) );
XOR U16127 ( .A(c3225), .B(b[3225]), .Z(n9676) );
XNOR U16128 ( .A(b[3225]), .B(n9677), .Z(c[3225]) );
XNOR U16129 ( .A(a[3225]), .B(c3225), .Z(n9677) );
XOR U16130 ( .A(c3226), .B(n9678), .Z(c3227) );
ANDN U16131 ( .B(n9679), .A(n9680), .Z(n9678) );
XOR U16132 ( .A(c3226), .B(b[3226]), .Z(n9679) );
XNOR U16133 ( .A(b[3226]), .B(n9680), .Z(c[3226]) );
XNOR U16134 ( .A(a[3226]), .B(c3226), .Z(n9680) );
XOR U16135 ( .A(c3227), .B(n9681), .Z(c3228) );
ANDN U16136 ( .B(n9682), .A(n9683), .Z(n9681) );
XOR U16137 ( .A(c3227), .B(b[3227]), .Z(n9682) );
XNOR U16138 ( .A(b[3227]), .B(n9683), .Z(c[3227]) );
XNOR U16139 ( .A(a[3227]), .B(c3227), .Z(n9683) );
XOR U16140 ( .A(c3228), .B(n9684), .Z(c3229) );
ANDN U16141 ( .B(n9685), .A(n9686), .Z(n9684) );
XOR U16142 ( .A(c3228), .B(b[3228]), .Z(n9685) );
XNOR U16143 ( .A(b[3228]), .B(n9686), .Z(c[3228]) );
XNOR U16144 ( .A(a[3228]), .B(c3228), .Z(n9686) );
XOR U16145 ( .A(c3229), .B(n9687), .Z(c3230) );
ANDN U16146 ( .B(n9688), .A(n9689), .Z(n9687) );
XOR U16147 ( .A(c3229), .B(b[3229]), .Z(n9688) );
XNOR U16148 ( .A(b[3229]), .B(n9689), .Z(c[3229]) );
XNOR U16149 ( .A(a[3229]), .B(c3229), .Z(n9689) );
XOR U16150 ( .A(c3230), .B(n9690), .Z(c3231) );
ANDN U16151 ( .B(n9691), .A(n9692), .Z(n9690) );
XOR U16152 ( .A(c3230), .B(b[3230]), .Z(n9691) );
XNOR U16153 ( .A(b[3230]), .B(n9692), .Z(c[3230]) );
XNOR U16154 ( .A(a[3230]), .B(c3230), .Z(n9692) );
XOR U16155 ( .A(c3231), .B(n9693), .Z(c3232) );
ANDN U16156 ( .B(n9694), .A(n9695), .Z(n9693) );
XOR U16157 ( .A(c3231), .B(b[3231]), .Z(n9694) );
XNOR U16158 ( .A(b[3231]), .B(n9695), .Z(c[3231]) );
XNOR U16159 ( .A(a[3231]), .B(c3231), .Z(n9695) );
XOR U16160 ( .A(c3232), .B(n9696), .Z(c3233) );
ANDN U16161 ( .B(n9697), .A(n9698), .Z(n9696) );
XOR U16162 ( .A(c3232), .B(b[3232]), .Z(n9697) );
XNOR U16163 ( .A(b[3232]), .B(n9698), .Z(c[3232]) );
XNOR U16164 ( .A(a[3232]), .B(c3232), .Z(n9698) );
XOR U16165 ( .A(c3233), .B(n9699), .Z(c3234) );
ANDN U16166 ( .B(n9700), .A(n9701), .Z(n9699) );
XOR U16167 ( .A(c3233), .B(b[3233]), .Z(n9700) );
XNOR U16168 ( .A(b[3233]), .B(n9701), .Z(c[3233]) );
XNOR U16169 ( .A(a[3233]), .B(c3233), .Z(n9701) );
XOR U16170 ( .A(c3234), .B(n9702), .Z(c3235) );
ANDN U16171 ( .B(n9703), .A(n9704), .Z(n9702) );
XOR U16172 ( .A(c3234), .B(b[3234]), .Z(n9703) );
XNOR U16173 ( .A(b[3234]), .B(n9704), .Z(c[3234]) );
XNOR U16174 ( .A(a[3234]), .B(c3234), .Z(n9704) );
XOR U16175 ( .A(c3235), .B(n9705), .Z(c3236) );
ANDN U16176 ( .B(n9706), .A(n9707), .Z(n9705) );
XOR U16177 ( .A(c3235), .B(b[3235]), .Z(n9706) );
XNOR U16178 ( .A(b[3235]), .B(n9707), .Z(c[3235]) );
XNOR U16179 ( .A(a[3235]), .B(c3235), .Z(n9707) );
XOR U16180 ( .A(c3236), .B(n9708), .Z(c3237) );
ANDN U16181 ( .B(n9709), .A(n9710), .Z(n9708) );
XOR U16182 ( .A(c3236), .B(b[3236]), .Z(n9709) );
XNOR U16183 ( .A(b[3236]), .B(n9710), .Z(c[3236]) );
XNOR U16184 ( .A(a[3236]), .B(c3236), .Z(n9710) );
XOR U16185 ( .A(c3237), .B(n9711), .Z(c3238) );
ANDN U16186 ( .B(n9712), .A(n9713), .Z(n9711) );
XOR U16187 ( .A(c3237), .B(b[3237]), .Z(n9712) );
XNOR U16188 ( .A(b[3237]), .B(n9713), .Z(c[3237]) );
XNOR U16189 ( .A(a[3237]), .B(c3237), .Z(n9713) );
XOR U16190 ( .A(c3238), .B(n9714), .Z(c3239) );
ANDN U16191 ( .B(n9715), .A(n9716), .Z(n9714) );
XOR U16192 ( .A(c3238), .B(b[3238]), .Z(n9715) );
XNOR U16193 ( .A(b[3238]), .B(n9716), .Z(c[3238]) );
XNOR U16194 ( .A(a[3238]), .B(c3238), .Z(n9716) );
XOR U16195 ( .A(c3239), .B(n9717), .Z(c3240) );
ANDN U16196 ( .B(n9718), .A(n9719), .Z(n9717) );
XOR U16197 ( .A(c3239), .B(b[3239]), .Z(n9718) );
XNOR U16198 ( .A(b[3239]), .B(n9719), .Z(c[3239]) );
XNOR U16199 ( .A(a[3239]), .B(c3239), .Z(n9719) );
XOR U16200 ( .A(c3240), .B(n9720), .Z(c3241) );
ANDN U16201 ( .B(n9721), .A(n9722), .Z(n9720) );
XOR U16202 ( .A(c3240), .B(b[3240]), .Z(n9721) );
XNOR U16203 ( .A(b[3240]), .B(n9722), .Z(c[3240]) );
XNOR U16204 ( .A(a[3240]), .B(c3240), .Z(n9722) );
XOR U16205 ( .A(c3241), .B(n9723), .Z(c3242) );
ANDN U16206 ( .B(n9724), .A(n9725), .Z(n9723) );
XOR U16207 ( .A(c3241), .B(b[3241]), .Z(n9724) );
XNOR U16208 ( .A(b[3241]), .B(n9725), .Z(c[3241]) );
XNOR U16209 ( .A(a[3241]), .B(c3241), .Z(n9725) );
XOR U16210 ( .A(c3242), .B(n9726), .Z(c3243) );
ANDN U16211 ( .B(n9727), .A(n9728), .Z(n9726) );
XOR U16212 ( .A(c3242), .B(b[3242]), .Z(n9727) );
XNOR U16213 ( .A(b[3242]), .B(n9728), .Z(c[3242]) );
XNOR U16214 ( .A(a[3242]), .B(c3242), .Z(n9728) );
XOR U16215 ( .A(c3243), .B(n9729), .Z(c3244) );
ANDN U16216 ( .B(n9730), .A(n9731), .Z(n9729) );
XOR U16217 ( .A(c3243), .B(b[3243]), .Z(n9730) );
XNOR U16218 ( .A(b[3243]), .B(n9731), .Z(c[3243]) );
XNOR U16219 ( .A(a[3243]), .B(c3243), .Z(n9731) );
XOR U16220 ( .A(c3244), .B(n9732), .Z(c3245) );
ANDN U16221 ( .B(n9733), .A(n9734), .Z(n9732) );
XOR U16222 ( .A(c3244), .B(b[3244]), .Z(n9733) );
XNOR U16223 ( .A(b[3244]), .B(n9734), .Z(c[3244]) );
XNOR U16224 ( .A(a[3244]), .B(c3244), .Z(n9734) );
XOR U16225 ( .A(c3245), .B(n9735), .Z(c3246) );
ANDN U16226 ( .B(n9736), .A(n9737), .Z(n9735) );
XOR U16227 ( .A(c3245), .B(b[3245]), .Z(n9736) );
XNOR U16228 ( .A(b[3245]), .B(n9737), .Z(c[3245]) );
XNOR U16229 ( .A(a[3245]), .B(c3245), .Z(n9737) );
XOR U16230 ( .A(c3246), .B(n9738), .Z(c3247) );
ANDN U16231 ( .B(n9739), .A(n9740), .Z(n9738) );
XOR U16232 ( .A(c3246), .B(b[3246]), .Z(n9739) );
XNOR U16233 ( .A(b[3246]), .B(n9740), .Z(c[3246]) );
XNOR U16234 ( .A(a[3246]), .B(c3246), .Z(n9740) );
XOR U16235 ( .A(c3247), .B(n9741), .Z(c3248) );
ANDN U16236 ( .B(n9742), .A(n9743), .Z(n9741) );
XOR U16237 ( .A(c3247), .B(b[3247]), .Z(n9742) );
XNOR U16238 ( .A(b[3247]), .B(n9743), .Z(c[3247]) );
XNOR U16239 ( .A(a[3247]), .B(c3247), .Z(n9743) );
XOR U16240 ( .A(c3248), .B(n9744), .Z(c3249) );
ANDN U16241 ( .B(n9745), .A(n9746), .Z(n9744) );
XOR U16242 ( .A(c3248), .B(b[3248]), .Z(n9745) );
XNOR U16243 ( .A(b[3248]), .B(n9746), .Z(c[3248]) );
XNOR U16244 ( .A(a[3248]), .B(c3248), .Z(n9746) );
XOR U16245 ( .A(c3249), .B(n9747), .Z(c3250) );
ANDN U16246 ( .B(n9748), .A(n9749), .Z(n9747) );
XOR U16247 ( .A(c3249), .B(b[3249]), .Z(n9748) );
XNOR U16248 ( .A(b[3249]), .B(n9749), .Z(c[3249]) );
XNOR U16249 ( .A(a[3249]), .B(c3249), .Z(n9749) );
XOR U16250 ( .A(c3250), .B(n9750), .Z(c3251) );
ANDN U16251 ( .B(n9751), .A(n9752), .Z(n9750) );
XOR U16252 ( .A(c3250), .B(b[3250]), .Z(n9751) );
XNOR U16253 ( .A(b[3250]), .B(n9752), .Z(c[3250]) );
XNOR U16254 ( .A(a[3250]), .B(c3250), .Z(n9752) );
XOR U16255 ( .A(c3251), .B(n9753), .Z(c3252) );
ANDN U16256 ( .B(n9754), .A(n9755), .Z(n9753) );
XOR U16257 ( .A(c3251), .B(b[3251]), .Z(n9754) );
XNOR U16258 ( .A(b[3251]), .B(n9755), .Z(c[3251]) );
XNOR U16259 ( .A(a[3251]), .B(c3251), .Z(n9755) );
XOR U16260 ( .A(c3252), .B(n9756), .Z(c3253) );
ANDN U16261 ( .B(n9757), .A(n9758), .Z(n9756) );
XOR U16262 ( .A(c3252), .B(b[3252]), .Z(n9757) );
XNOR U16263 ( .A(b[3252]), .B(n9758), .Z(c[3252]) );
XNOR U16264 ( .A(a[3252]), .B(c3252), .Z(n9758) );
XOR U16265 ( .A(c3253), .B(n9759), .Z(c3254) );
ANDN U16266 ( .B(n9760), .A(n9761), .Z(n9759) );
XOR U16267 ( .A(c3253), .B(b[3253]), .Z(n9760) );
XNOR U16268 ( .A(b[3253]), .B(n9761), .Z(c[3253]) );
XNOR U16269 ( .A(a[3253]), .B(c3253), .Z(n9761) );
XOR U16270 ( .A(c3254), .B(n9762), .Z(c3255) );
ANDN U16271 ( .B(n9763), .A(n9764), .Z(n9762) );
XOR U16272 ( .A(c3254), .B(b[3254]), .Z(n9763) );
XNOR U16273 ( .A(b[3254]), .B(n9764), .Z(c[3254]) );
XNOR U16274 ( .A(a[3254]), .B(c3254), .Z(n9764) );
XOR U16275 ( .A(c3255), .B(n9765), .Z(c3256) );
ANDN U16276 ( .B(n9766), .A(n9767), .Z(n9765) );
XOR U16277 ( .A(c3255), .B(b[3255]), .Z(n9766) );
XNOR U16278 ( .A(b[3255]), .B(n9767), .Z(c[3255]) );
XNOR U16279 ( .A(a[3255]), .B(c3255), .Z(n9767) );
XOR U16280 ( .A(c3256), .B(n9768), .Z(c3257) );
ANDN U16281 ( .B(n9769), .A(n9770), .Z(n9768) );
XOR U16282 ( .A(c3256), .B(b[3256]), .Z(n9769) );
XNOR U16283 ( .A(b[3256]), .B(n9770), .Z(c[3256]) );
XNOR U16284 ( .A(a[3256]), .B(c3256), .Z(n9770) );
XOR U16285 ( .A(c3257), .B(n9771), .Z(c3258) );
ANDN U16286 ( .B(n9772), .A(n9773), .Z(n9771) );
XOR U16287 ( .A(c3257), .B(b[3257]), .Z(n9772) );
XNOR U16288 ( .A(b[3257]), .B(n9773), .Z(c[3257]) );
XNOR U16289 ( .A(a[3257]), .B(c3257), .Z(n9773) );
XOR U16290 ( .A(c3258), .B(n9774), .Z(c3259) );
ANDN U16291 ( .B(n9775), .A(n9776), .Z(n9774) );
XOR U16292 ( .A(c3258), .B(b[3258]), .Z(n9775) );
XNOR U16293 ( .A(b[3258]), .B(n9776), .Z(c[3258]) );
XNOR U16294 ( .A(a[3258]), .B(c3258), .Z(n9776) );
XOR U16295 ( .A(c3259), .B(n9777), .Z(c3260) );
ANDN U16296 ( .B(n9778), .A(n9779), .Z(n9777) );
XOR U16297 ( .A(c3259), .B(b[3259]), .Z(n9778) );
XNOR U16298 ( .A(b[3259]), .B(n9779), .Z(c[3259]) );
XNOR U16299 ( .A(a[3259]), .B(c3259), .Z(n9779) );
XOR U16300 ( .A(c3260), .B(n9780), .Z(c3261) );
ANDN U16301 ( .B(n9781), .A(n9782), .Z(n9780) );
XOR U16302 ( .A(c3260), .B(b[3260]), .Z(n9781) );
XNOR U16303 ( .A(b[3260]), .B(n9782), .Z(c[3260]) );
XNOR U16304 ( .A(a[3260]), .B(c3260), .Z(n9782) );
XOR U16305 ( .A(c3261), .B(n9783), .Z(c3262) );
ANDN U16306 ( .B(n9784), .A(n9785), .Z(n9783) );
XOR U16307 ( .A(c3261), .B(b[3261]), .Z(n9784) );
XNOR U16308 ( .A(b[3261]), .B(n9785), .Z(c[3261]) );
XNOR U16309 ( .A(a[3261]), .B(c3261), .Z(n9785) );
XOR U16310 ( .A(c3262), .B(n9786), .Z(c3263) );
ANDN U16311 ( .B(n9787), .A(n9788), .Z(n9786) );
XOR U16312 ( .A(c3262), .B(b[3262]), .Z(n9787) );
XNOR U16313 ( .A(b[3262]), .B(n9788), .Z(c[3262]) );
XNOR U16314 ( .A(a[3262]), .B(c3262), .Z(n9788) );
XOR U16315 ( .A(c3263), .B(n9789), .Z(c3264) );
ANDN U16316 ( .B(n9790), .A(n9791), .Z(n9789) );
XOR U16317 ( .A(c3263), .B(b[3263]), .Z(n9790) );
XNOR U16318 ( .A(b[3263]), .B(n9791), .Z(c[3263]) );
XNOR U16319 ( .A(a[3263]), .B(c3263), .Z(n9791) );
XOR U16320 ( .A(c3264), .B(n9792), .Z(c3265) );
ANDN U16321 ( .B(n9793), .A(n9794), .Z(n9792) );
XOR U16322 ( .A(c3264), .B(b[3264]), .Z(n9793) );
XNOR U16323 ( .A(b[3264]), .B(n9794), .Z(c[3264]) );
XNOR U16324 ( .A(a[3264]), .B(c3264), .Z(n9794) );
XOR U16325 ( .A(c3265), .B(n9795), .Z(c3266) );
ANDN U16326 ( .B(n9796), .A(n9797), .Z(n9795) );
XOR U16327 ( .A(c3265), .B(b[3265]), .Z(n9796) );
XNOR U16328 ( .A(b[3265]), .B(n9797), .Z(c[3265]) );
XNOR U16329 ( .A(a[3265]), .B(c3265), .Z(n9797) );
XOR U16330 ( .A(c3266), .B(n9798), .Z(c3267) );
ANDN U16331 ( .B(n9799), .A(n9800), .Z(n9798) );
XOR U16332 ( .A(c3266), .B(b[3266]), .Z(n9799) );
XNOR U16333 ( .A(b[3266]), .B(n9800), .Z(c[3266]) );
XNOR U16334 ( .A(a[3266]), .B(c3266), .Z(n9800) );
XOR U16335 ( .A(c3267), .B(n9801), .Z(c3268) );
ANDN U16336 ( .B(n9802), .A(n9803), .Z(n9801) );
XOR U16337 ( .A(c3267), .B(b[3267]), .Z(n9802) );
XNOR U16338 ( .A(b[3267]), .B(n9803), .Z(c[3267]) );
XNOR U16339 ( .A(a[3267]), .B(c3267), .Z(n9803) );
XOR U16340 ( .A(c3268), .B(n9804), .Z(c3269) );
ANDN U16341 ( .B(n9805), .A(n9806), .Z(n9804) );
XOR U16342 ( .A(c3268), .B(b[3268]), .Z(n9805) );
XNOR U16343 ( .A(b[3268]), .B(n9806), .Z(c[3268]) );
XNOR U16344 ( .A(a[3268]), .B(c3268), .Z(n9806) );
XOR U16345 ( .A(c3269), .B(n9807), .Z(c3270) );
ANDN U16346 ( .B(n9808), .A(n9809), .Z(n9807) );
XOR U16347 ( .A(c3269), .B(b[3269]), .Z(n9808) );
XNOR U16348 ( .A(b[3269]), .B(n9809), .Z(c[3269]) );
XNOR U16349 ( .A(a[3269]), .B(c3269), .Z(n9809) );
XOR U16350 ( .A(c3270), .B(n9810), .Z(c3271) );
ANDN U16351 ( .B(n9811), .A(n9812), .Z(n9810) );
XOR U16352 ( .A(c3270), .B(b[3270]), .Z(n9811) );
XNOR U16353 ( .A(b[3270]), .B(n9812), .Z(c[3270]) );
XNOR U16354 ( .A(a[3270]), .B(c3270), .Z(n9812) );
XOR U16355 ( .A(c3271), .B(n9813), .Z(c3272) );
ANDN U16356 ( .B(n9814), .A(n9815), .Z(n9813) );
XOR U16357 ( .A(c3271), .B(b[3271]), .Z(n9814) );
XNOR U16358 ( .A(b[3271]), .B(n9815), .Z(c[3271]) );
XNOR U16359 ( .A(a[3271]), .B(c3271), .Z(n9815) );
XOR U16360 ( .A(c3272), .B(n9816), .Z(c3273) );
ANDN U16361 ( .B(n9817), .A(n9818), .Z(n9816) );
XOR U16362 ( .A(c3272), .B(b[3272]), .Z(n9817) );
XNOR U16363 ( .A(b[3272]), .B(n9818), .Z(c[3272]) );
XNOR U16364 ( .A(a[3272]), .B(c3272), .Z(n9818) );
XOR U16365 ( .A(c3273), .B(n9819), .Z(c3274) );
ANDN U16366 ( .B(n9820), .A(n9821), .Z(n9819) );
XOR U16367 ( .A(c3273), .B(b[3273]), .Z(n9820) );
XNOR U16368 ( .A(b[3273]), .B(n9821), .Z(c[3273]) );
XNOR U16369 ( .A(a[3273]), .B(c3273), .Z(n9821) );
XOR U16370 ( .A(c3274), .B(n9822), .Z(c3275) );
ANDN U16371 ( .B(n9823), .A(n9824), .Z(n9822) );
XOR U16372 ( .A(c3274), .B(b[3274]), .Z(n9823) );
XNOR U16373 ( .A(b[3274]), .B(n9824), .Z(c[3274]) );
XNOR U16374 ( .A(a[3274]), .B(c3274), .Z(n9824) );
XOR U16375 ( .A(c3275), .B(n9825), .Z(c3276) );
ANDN U16376 ( .B(n9826), .A(n9827), .Z(n9825) );
XOR U16377 ( .A(c3275), .B(b[3275]), .Z(n9826) );
XNOR U16378 ( .A(b[3275]), .B(n9827), .Z(c[3275]) );
XNOR U16379 ( .A(a[3275]), .B(c3275), .Z(n9827) );
XOR U16380 ( .A(c3276), .B(n9828), .Z(c3277) );
ANDN U16381 ( .B(n9829), .A(n9830), .Z(n9828) );
XOR U16382 ( .A(c3276), .B(b[3276]), .Z(n9829) );
XNOR U16383 ( .A(b[3276]), .B(n9830), .Z(c[3276]) );
XNOR U16384 ( .A(a[3276]), .B(c3276), .Z(n9830) );
XOR U16385 ( .A(c3277), .B(n9831), .Z(c3278) );
ANDN U16386 ( .B(n9832), .A(n9833), .Z(n9831) );
XOR U16387 ( .A(c3277), .B(b[3277]), .Z(n9832) );
XNOR U16388 ( .A(b[3277]), .B(n9833), .Z(c[3277]) );
XNOR U16389 ( .A(a[3277]), .B(c3277), .Z(n9833) );
XOR U16390 ( .A(c3278), .B(n9834), .Z(c3279) );
ANDN U16391 ( .B(n9835), .A(n9836), .Z(n9834) );
XOR U16392 ( .A(c3278), .B(b[3278]), .Z(n9835) );
XNOR U16393 ( .A(b[3278]), .B(n9836), .Z(c[3278]) );
XNOR U16394 ( .A(a[3278]), .B(c3278), .Z(n9836) );
XOR U16395 ( .A(c3279), .B(n9837), .Z(c3280) );
ANDN U16396 ( .B(n9838), .A(n9839), .Z(n9837) );
XOR U16397 ( .A(c3279), .B(b[3279]), .Z(n9838) );
XNOR U16398 ( .A(b[3279]), .B(n9839), .Z(c[3279]) );
XNOR U16399 ( .A(a[3279]), .B(c3279), .Z(n9839) );
XOR U16400 ( .A(c3280), .B(n9840), .Z(c3281) );
ANDN U16401 ( .B(n9841), .A(n9842), .Z(n9840) );
XOR U16402 ( .A(c3280), .B(b[3280]), .Z(n9841) );
XNOR U16403 ( .A(b[3280]), .B(n9842), .Z(c[3280]) );
XNOR U16404 ( .A(a[3280]), .B(c3280), .Z(n9842) );
XOR U16405 ( .A(c3281), .B(n9843), .Z(c3282) );
ANDN U16406 ( .B(n9844), .A(n9845), .Z(n9843) );
XOR U16407 ( .A(c3281), .B(b[3281]), .Z(n9844) );
XNOR U16408 ( .A(b[3281]), .B(n9845), .Z(c[3281]) );
XNOR U16409 ( .A(a[3281]), .B(c3281), .Z(n9845) );
XOR U16410 ( .A(c3282), .B(n9846), .Z(c3283) );
ANDN U16411 ( .B(n9847), .A(n9848), .Z(n9846) );
XOR U16412 ( .A(c3282), .B(b[3282]), .Z(n9847) );
XNOR U16413 ( .A(b[3282]), .B(n9848), .Z(c[3282]) );
XNOR U16414 ( .A(a[3282]), .B(c3282), .Z(n9848) );
XOR U16415 ( .A(c3283), .B(n9849), .Z(c3284) );
ANDN U16416 ( .B(n9850), .A(n9851), .Z(n9849) );
XOR U16417 ( .A(c3283), .B(b[3283]), .Z(n9850) );
XNOR U16418 ( .A(b[3283]), .B(n9851), .Z(c[3283]) );
XNOR U16419 ( .A(a[3283]), .B(c3283), .Z(n9851) );
XOR U16420 ( .A(c3284), .B(n9852), .Z(c3285) );
ANDN U16421 ( .B(n9853), .A(n9854), .Z(n9852) );
XOR U16422 ( .A(c3284), .B(b[3284]), .Z(n9853) );
XNOR U16423 ( .A(b[3284]), .B(n9854), .Z(c[3284]) );
XNOR U16424 ( .A(a[3284]), .B(c3284), .Z(n9854) );
XOR U16425 ( .A(c3285), .B(n9855), .Z(c3286) );
ANDN U16426 ( .B(n9856), .A(n9857), .Z(n9855) );
XOR U16427 ( .A(c3285), .B(b[3285]), .Z(n9856) );
XNOR U16428 ( .A(b[3285]), .B(n9857), .Z(c[3285]) );
XNOR U16429 ( .A(a[3285]), .B(c3285), .Z(n9857) );
XOR U16430 ( .A(c3286), .B(n9858), .Z(c3287) );
ANDN U16431 ( .B(n9859), .A(n9860), .Z(n9858) );
XOR U16432 ( .A(c3286), .B(b[3286]), .Z(n9859) );
XNOR U16433 ( .A(b[3286]), .B(n9860), .Z(c[3286]) );
XNOR U16434 ( .A(a[3286]), .B(c3286), .Z(n9860) );
XOR U16435 ( .A(c3287), .B(n9861), .Z(c3288) );
ANDN U16436 ( .B(n9862), .A(n9863), .Z(n9861) );
XOR U16437 ( .A(c3287), .B(b[3287]), .Z(n9862) );
XNOR U16438 ( .A(b[3287]), .B(n9863), .Z(c[3287]) );
XNOR U16439 ( .A(a[3287]), .B(c3287), .Z(n9863) );
XOR U16440 ( .A(c3288), .B(n9864), .Z(c3289) );
ANDN U16441 ( .B(n9865), .A(n9866), .Z(n9864) );
XOR U16442 ( .A(c3288), .B(b[3288]), .Z(n9865) );
XNOR U16443 ( .A(b[3288]), .B(n9866), .Z(c[3288]) );
XNOR U16444 ( .A(a[3288]), .B(c3288), .Z(n9866) );
XOR U16445 ( .A(c3289), .B(n9867), .Z(c3290) );
ANDN U16446 ( .B(n9868), .A(n9869), .Z(n9867) );
XOR U16447 ( .A(c3289), .B(b[3289]), .Z(n9868) );
XNOR U16448 ( .A(b[3289]), .B(n9869), .Z(c[3289]) );
XNOR U16449 ( .A(a[3289]), .B(c3289), .Z(n9869) );
XOR U16450 ( .A(c3290), .B(n9870), .Z(c3291) );
ANDN U16451 ( .B(n9871), .A(n9872), .Z(n9870) );
XOR U16452 ( .A(c3290), .B(b[3290]), .Z(n9871) );
XNOR U16453 ( .A(b[3290]), .B(n9872), .Z(c[3290]) );
XNOR U16454 ( .A(a[3290]), .B(c3290), .Z(n9872) );
XOR U16455 ( .A(c3291), .B(n9873), .Z(c3292) );
ANDN U16456 ( .B(n9874), .A(n9875), .Z(n9873) );
XOR U16457 ( .A(c3291), .B(b[3291]), .Z(n9874) );
XNOR U16458 ( .A(b[3291]), .B(n9875), .Z(c[3291]) );
XNOR U16459 ( .A(a[3291]), .B(c3291), .Z(n9875) );
XOR U16460 ( .A(c3292), .B(n9876), .Z(c3293) );
ANDN U16461 ( .B(n9877), .A(n9878), .Z(n9876) );
XOR U16462 ( .A(c3292), .B(b[3292]), .Z(n9877) );
XNOR U16463 ( .A(b[3292]), .B(n9878), .Z(c[3292]) );
XNOR U16464 ( .A(a[3292]), .B(c3292), .Z(n9878) );
XOR U16465 ( .A(c3293), .B(n9879), .Z(c3294) );
ANDN U16466 ( .B(n9880), .A(n9881), .Z(n9879) );
XOR U16467 ( .A(c3293), .B(b[3293]), .Z(n9880) );
XNOR U16468 ( .A(b[3293]), .B(n9881), .Z(c[3293]) );
XNOR U16469 ( .A(a[3293]), .B(c3293), .Z(n9881) );
XOR U16470 ( .A(c3294), .B(n9882), .Z(c3295) );
ANDN U16471 ( .B(n9883), .A(n9884), .Z(n9882) );
XOR U16472 ( .A(c3294), .B(b[3294]), .Z(n9883) );
XNOR U16473 ( .A(b[3294]), .B(n9884), .Z(c[3294]) );
XNOR U16474 ( .A(a[3294]), .B(c3294), .Z(n9884) );
XOR U16475 ( .A(c3295), .B(n9885), .Z(c3296) );
ANDN U16476 ( .B(n9886), .A(n9887), .Z(n9885) );
XOR U16477 ( .A(c3295), .B(b[3295]), .Z(n9886) );
XNOR U16478 ( .A(b[3295]), .B(n9887), .Z(c[3295]) );
XNOR U16479 ( .A(a[3295]), .B(c3295), .Z(n9887) );
XOR U16480 ( .A(c3296), .B(n9888), .Z(c3297) );
ANDN U16481 ( .B(n9889), .A(n9890), .Z(n9888) );
XOR U16482 ( .A(c3296), .B(b[3296]), .Z(n9889) );
XNOR U16483 ( .A(b[3296]), .B(n9890), .Z(c[3296]) );
XNOR U16484 ( .A(a[3296]), .B(c3296), .Z(n9890) );
XOR U16485 ( .A(c3297), .B(n9891), .Z(c3298) );
ANDN U16486 ( .B(n9892), .A(n9893), .Z(n9891) );
XOR U16487 ( .A(c3297), .B(b[3297]), .Z(n9892) );
XNOR U16488 ( .A(b[3297]), .B(n9893), .Z(c[3297]) );
XNOR U16489 ( .A(a[3297]), .B(c3297), .Z(n9893) );
XOR U16490 ( .A(c3298), .B(n9894), .Z(c3299) );
ANDN U16491 ( .B(n9895), .A(n9896), .Z(n9894) );
XOR U16492 ( .A(c3298), .B(b[3298]), .Z(n9895) );
XNOR U16493 ( .A(b[3298]), .B(n9896), .Z(c[3298]) );
XNOR U16494 ( .A(a[3298]), .B(c3298), .Z(n9896) );
XOR U16495 ( .A(c3299), .B(n9897), .Z(c3300) );
ANDN U16496 ( .B(n9898), .A(n9899), .Z(n9897) );
XOR U16497 ( .A(c3299), .B(b[3299]), .Z(n9898) );
XNOR U16498 ( .A(b[3299]), .B(n9899), .Z(c[3299]) );
XNOR U16499 ( .A(a[3299]), .B(c3299), .Z(n9899) );
XOR U16500 ( .A(c3300), .B(n9900), .Z(c3301) );
ANDN U16501 ( .B(n9901), .A(n9902), .Z(n9900) );
XOR U16502 ( .A(c3300), .B(b[3300]), .Z(n9901) );
XNOR U16503 ( .A(b[3300]), .B(n9902), .Z(c[3300]) );
XNOR U16504 ( .A(a[3300]), .B(c3300), .Z(n9902) );
XOR U16505 ( .A(c3301), .B(n9903), .Z(c3302) );
ANDN U16506 ( .B(n9904), .A(n9905), .Z(n9903) );
XOR U16507 ( .A(c3301), .B(b[3301]), .Z(n9904) );
XNOR U16508 ( .A(b[3301]), .B(n9905), .Z(c[3301]) );
XNOR U16509 ( .A(a[3301]), .B(c3301), .Z(n9905) );
XOR U16510 ( .A(c3302), .B(n9906), .Z(c3303) );
ANDN U16511 ( .B(n9907), .A(n9908), .Z(n9906) );
XOR U16512 ( .A(c3302), .B(b[3302]), .Z(n9907) );
XNOR U16513 ( .A(b[3302]), .B(n9908), .Z(c[3302]) );
XNOR U16514 ( .A(a[3302]), .B(c3302), .Z(n9908) );
XOR U16515 ( .A(c3303), .B(n9909), .Z(c3304) );
ANDN U16516 ( .B(n9910), .A(n9911), .Z(n9909) );
XOR U16517 ( .A(c3303), .B(b[3303]), .Z(n9910) );
XNOR U16518 ( .A(b[3303]), .B(n9911), .Z(c[3303]) );
XNOR U16519 ( .A(a[3303]), .B(c3303), .Z(n9911) );
XOR U16520 ( .A(c3304), .B(n9912), .Z(c3305) );
ANDN U16521 ( .B(n9913), .A(n9914), .Z(n9912) );
XOR U16522 ( .A(c3304), .B(b[3304]), .Z(n9913) );
XNOR U16523 ( .A(b[3304]), .B(n9914), .Z(c[3304]) );
XNOR U16524 ( .A(a[3304]), .B(c3304), .Z(n9914) );
XOR U16525 ( .A(c3305), .B(n9915), .Z(c3306) );
ANDN U16526 ( .B(n9916), .A(n9917), .Z(n9915) );
XOR U16527 ( .A(c3305), .B(b[3305]), .Z(n9916) );
XNOR U16528 ( .A(b[3305]), .B(n9917), .Z(c[3305]) );
XNOR U16529 ( .A(a[3305]), .B(c3305), .Z(n9917) );
XOR U16530 ( .A(c3306), .B(n9918), .Z(c3307) );
ANDN U16531 ( .B(n9919), .A(n9920), .Z(n9918) );
XOR U16532 ( .A(c3306), .B(b[3306]), .Z(n9919) );
XNOR U16533 ( .A(b[3306]), .B(n9920), .Z(c[3306]) );
XNOR U16534 ( .A(a[3306]), .B(c3306), .Z(n9920) );
XOR U16535 ( .A(c3307), .B(n9921), .Z(c3308) );
ANDN U16536 ( .B(n9922), .A(n9923), .Z(n9921) );
XOR U16537 ( .A(c3307), .B(b[3307]), .Z(n9922) );
XNOR U16538 ( .A(b[3307]), .B(n9923), .Z(c[3307]) );
XNOR U16539 ( .A(a[3307]), .B(c3307), .Z(n9923) );
XOR U16540 ( .A(c3308), .B(n9924), .Z(c3309) );
ANDN U16541 ( .B(n9925), .A(n9926), .Z(n9924) );
XOR U16542 ( .A(c3308), .B(b[3308]), .Z(n9925) );
XNOR U16543 ( .A(b[3308]), .B(n9926), .Z(c[3308]) );
XNOR U16544 ( .A(a[3308]), .B(c3308), .Z(n9926) );
XOR U16545 ( .A(c3309), .B(n9927), .Z(c3310) );
ANDN U16546 ( .B(n9928), .A(n9929), .Z(n9927) );
XOR U16547 ( .A(c3309), .B(b[3309]), .Z(n9928) );
XNOR U16548 ( .A(b[3309]), .B(n9929), .Z(c[3309]) );
XNOR U16549 ( .A(a[3309]), .B(c3309), .Z(n9929) );
XOR U16550 ( .A(c3310), .B(n9930), .Z(c3311) );
ANDN U16551 ( .B(n9931), .A(n9932), .Z(n9930) );
XOR U16552 ( .A(c3310), .B(b[3310]), .Z(n9931) );
XNOR U16553 ( .A(b[3310]), .B(n9932), .Z(c[3310]) );
XNOR U16554 ( .A(a[3310]), .B(c3310), .Z(n9932) );
XOR U16555 ( .A(c3311), .B(n9933), .Z(c3312) );
ANDN U16556 ( .B(n9934), .A(n9935), .Z(n9933) );
XOR U16557 ( .A(c3311), .B(b[3311]), .Z(n9934) );
XNOR U16558 ( .A(b[3311]), .B(n9935), .Z(c[3311]) );
XNOR U16559 ( .A(a[3311]), .B(c3311), .Z(n9935) );
XOR U16560 ( .A(c3312), .B(n9936), .Z(c3313) );
ANDN U16561 ( .B(n9937), .A(n9938), .Z(n9936) );
XOR U16562 ( .A(c3312), .B(b[3312]), .Z(n9937) );
XNOR U16563 ( .A(b[3312]), .B(n9938), .Z(c[3312]) );
XNOR U16564 ( .A(a[3312]), .B(c3312), .Z(n9938) );
XOR U16565 ( .A(c3313), .B(n9939), .Z(c3314) );
ANDN U16566 ( .B(n9940), .A(n9941), .Z(n9939) );
XOR U16567 ( .A(c3313), .B(b[3313]), .Z(n9940) );
XNOR U16568 ( .A(b[3313]), .B(n9941), .Z(c[3313]) );
XNOR U16569 ( .A(a[3313]), .B(c3313), .Z(n9941) );
XOR U16570 ( .A(c3314), .B(n9942), .Z(c3315) );
ANDN U16571 ( .B(n9943), .A(n9944), .Z(n9942) );
XOR U16572 ( .A(c3314), .B(b[3314]), .Z(n9943) );
XNOR U16573 ( .A(b[3314]), .B(n9944), .Z(c[3314]) );
XNOR U16574 ( .A(a[3314]), .B(c3314), .Z(n9944) );
XOR U16575 ( .A(c3315), .B(n9945), .Z(c3316) );
ANDN U16576 ( .B(n9946), .A(n9947), .Z(n9945) );
XOR U16577 ( .A(c3315), .B(b[3315]), .Z(n9946) );
XNOR U16578 ( .A(b[3315]), .B(n9947), .Z(c[3315]) );
XNOR U16579 ( .A(a[3315]), .B(c3315), .Z(n9947) );
XOR U16580 ( .A(c3316), .B(n9948), .Z(c3317) );
ANDN U16581 ( .B(n9949), .A(n9950), .Z(n9948) );
XOR U16582 ( .A(c3316), .B(b[3316]), .Z(n9949) );
XNOR U16583 ( .A(b[3316]), .B(n9950), .Z(c[3316]) );
XNOR U16584 ( .A(a[3316]), .B(c3316), .Z(n9950) );
XOR U16585 ( .A(c3317), .B(n9951), .Z(c3318) );
ANDN U16586 ( .B(n9952), .A(n9953), .Z(n9951) );
XOR U16587 ( .A(c3317), .B(b[3317]), .Z(n9952) );
XNOR U16588 ( .A(b[3317]), .B(n9953), .Z(c[3317]) );
XNOR U16589 ( .A(a[3317]), .B(c3317), .Z(n9953) );
XOR U16590 ( .A(c3318), .B(n9954), .Z(c3319) );
ANDN U16591 ( .B(n9955), .A(n9956), .Z(n9954) );
XOR U16592 ( .A(c3318), .B(b[3318]), .Z(n9955) );
XNOR U16593 ( .A(b[3318]), .B(n9956), .Z(c[3318]) );
XNOR U16594 ( .A(a[3318]), .B(c3318), .Z(n9956) );
XOR U16595 ( .A(c3319), .B(n9957), .Z(c3320) );
ANDN U16596 ( .B(n9958), .A(n9959), .Z(n9957) );
XOR U16597 ( .A(c3319), .B(b[3319]), .Z(n9958) );
XNOR U16598 ( .A(b[3319]), .B(n9959), .Z(c[3319]) );
XNOR U16599 ( .A(a[3319]), .B(c3319), .Z(n9959) );
XOR U16600 ( .A(c3320), .B(n9960), .Z(c3321) );
ANDN U16601 ( .B(n9961), .A(n9962), .Z(n9960) );
XOR U16602 ( .A(c3320), .B(b[3320]), .Z(n9961) );
XNOR U16603 ( .A(b[3320]), .B(n9962), .Z(c[3320]) );
XNOR U16604 ( .A(a[3320]), .B(c3320), .Z(n9962) );
XOR U16605 ( .A(c3321), .B(n9963), .Z(c3322) );
ANDN U16606 ( .B(n9964), .A(n9965), .Z(n9963) );
XOR U16607 ( .A(c3321), .B(b[3321]), .Z(n9964) );
XNOR U16608 ( .A(b[3321]), .B(n9965), .Z(c[3321]) );
XNOR U16609 ( .A(a[3321]), .B(c3321), .Z(n9965) );
XOR U16610 ( .A(c3322), .B(n9966), .Z(c3323) );
ANDN U16611 ( .B(n9967), .A(n9968), .Z(n9966) );
XOR U16612 ( .A(c3322), .B(b[3322]), .Z(n9967) );
XNOR U16613 ( .A(b[3322]), .B(n9968), .Z(c[3322]) );
XNOR U16614 ( .A(a[3322]), .B(c3322), .Z(n9968) );
XOR U16615 ( .A(c3323), .B(n9969), .Z(c3324) );
ANDN U16616 ( .B(n9970), .A(n9971), .Z(n9969) );
XOR U16617 ( .A(c3323), .B(b[3323]), .Z(n9970) );
XNOR U16618 ( .A(b[3323]), .B(n9971), .Z(c[3323]) );
XNOR U16619 ( .A(a[3323]), .B(c3323), .Z(n9971) );
XOR U16620 ( .A(c3324), .B(n9972), .Z(c3325) );
ANDN U16621 ( .B(n9973), .A(n9974), .Z(n9972) );
XOR U16622 ( .A(c3324), .B(b[3324]), .Z(n9973) );
XNOR U16623 ( .A(b[3324]), .B(n9974), .Z(c[3324]) );
XNOR U16624 ( .A(a[3324]), .B(c3324), .Z(n9974) );
XOR U16625 ( .A(c3325), .B(n9975), .Z(c3326) );
ANDN U16626 ( .B(n9976), .A(n9977), .Z(n9975) );
XOR U16627 ( .A(c3325), .B(b[3325]), .Z(n9976) );
XNOR U16628 ( .A(b[3325]), .B(n9977), .Z(c[3325]) );
XNOR U16629 ( .A(a[3325]), .B(c3325), .Z(n9977) );
XOR U16630 ( .A(c3326), .B(n9978), .Z(c3327) );
ANDN U16631 ( .B(n9979), .A(n9980), .Z(n9978) );
XOR U16632 ( .A(c3326), .B(b[3326]), .Z(n9979) );
XNOR U16633 ( .A(b[3326]), .B(n9980), .Z(c[3326]) );
XNOR U16634 ( .A(a[3326]), .B(c3326), .Z(n9980) );
XOR U16635 ( .A(c3327), .B(n9981), .Z(c3328) );
ANDN U16636 ( .B(n9982), .A(n9983), .Z(n9981) );
XOR U16637 ( .A(c3327), .B(b[3327]), .Z(n9982) );
XNOR U16638 ( .A(b[3327]), .B(n9983), .Z(c[3327]) );
XNOR U16639 ( .A(a[3327]), .B(c3327), .Z(n9983) );
XOR U16640 ( .A(c3328), .B(n9984), .Z(c3329) );
ANDN U16641 ( .B(n9985), .A(n9986), .Z(n9984) );
XOR U16642 ( .A(c3328), .B(b[3328]), .Z(n9985) );
XNOR U16643 ( .A(b[3328]), .B(n9986), .Z(c[3328]) );
XNOR U16644 ( .A(a[3328]), .B(c3328), .Z(n9986) );
XOR U16645 ( .A(c3329), .B(n9987), .Z(c3330) );
ANDN U16646 ( .B(n9988), .A(n9989), .Z(n9987) );
XOR U16647 ( .A(c3329), .B(b[3329]), .Z(n9988) );
XNOR U16648 ( .A(b[3329]), .B(n9989), .Z(c[3329]) );
XNOR U16649 ( .A(a[3329]), .B(c3329), .Z(n9989) );
XOR U16650 ( .A(c3330), .B(n9990), .Z(c3331) );
ANDN U16651 ( .B(n9991), .A(n9992), .Z(n9990) );
XOR U16652 ( .A(c3330), .B(b[3330]), .Z(n9991) );
XNOR U16653 ( .A(b[3330]), .B(n9992), .Z(c[3330]) );
XNOR U16654 ( .A(a[3330]), .B(c3330), .Z(n9992) );
XOR U16655 ( .A(c3331), .B(n9993), .Z(c3332) );
ANDN U16656 ( .B(n9994), .A(n9995), .Z(n9993) );
XOR U16657 ( .A(c3331), .B(b[3331]), .Z(n9994) );
XNOR U16658 ( .A(b[3331]), .B(n9995), .Z(c[3331]) );
XNOR U16659 ( .A(a[3331]), .B(c3331), .Z(n9995) );
XOR U16660 ( .A(c3332), .B(n9996), .Z(c3333) );
ANDN U16661 ( .B(n9997), .A(n9998), .Z(n9996) );
XOR U16662 ( .A(c3332), .B(b[3332]), .Z(n9997) );
XNOR U16663 ( .A(b[3332]), .B(n9998), .Z(c[3332]) );
XNOR U16664 ( .A(a[3332]), .B(c3332), .Z(n9998) );
XOR U16665 ( .A(c3333), .B(n9999), .Z(c3334) );
ANDN U16666 ( .B(n10000), .A(n10001), .Z(n9999) );
XOR U16667 ( .A(c3333), .B(b[3333]), .Z(n10000) );
XNOR U16668 ( .A(b[3333]), .B(n10001), .Z(c[3333]) );
XNOR U16669 ( .A(a[3333]), .B(c3333), .Z(n10001) );
XOR U16670 ( .A(c3334), .B(n10002), .Z(c3335) );
ANDN U16671 ( .B(n10003), .A(n10004), .Z(n10002) );
XOR U16672 ( .A(c3334), .B(b[3334]), .Z(n10003) );
XNOR U16673 ( .A(b[3334]), .B(n10004), .Z(c[3334]) );
XNOR U16674 ( .A(a[3334]), .B(c3334), .Z(n10004) );
XOR U16675 ( .A(c3335), .B(n10005), .Z(c3336) );
ANDN U16676 ( .B(n10006), .A(n10007), .Z(n10005) );
XOR U16677 ( .A(c3335), .B(b[3335]), .Z(n10006) );
XNOR U16678 ( .A(b[3335]), .B(n10007), .Z(c[3335]) );
XNOR U16679 ( .A(a[3335]), .B(c3335), .Z(n10007) );
XOR U16680 ( .A(c3336), .B(n10008), .Z(c3337) );
ANDN U16681 ( .B(n10009), .A(n10010), .Z(n10008) );
XOR U16682 ( .A(c3336), .B(b[3336]), .Z(n10009) );
XNOR U16683 ( .A(b[3336]), .B(n10010), .Z(c[3336]) );
XNOR U16684 ( .A(a[3336]), .B(c3336), .Z(n10010) );
XOR U16685 ( .A(c3337), .B(n10011), .Z(c3338) );
ANDN U16686 ( .B(n10012), .A(n10013), .Z(n10011) );
XOR U16687 ( .A(c3337), .B(b[3337]), .Z(n10012) );
XNOR U16688 ( .A(b[3337]), .B(n10013), .Z(c[3337]) );
XNOR U16689 ( .A(a[3337]), .B(c3337), .Z(n10013) );
XOR U16690 ( .A(c3338), .B(n10014), .Z(c3339) );
ANDN U16691 ( .B(n10015), .A(n10016), .Z(n10014) );
XOR U16692 ( .A(c3338), .B(b[3338]), .Z(n10015) );
XNOR U16693 ( .A(b[3338]), .B(n10016), .Z(c[3338]) );
XNOR U16694 ( .A(a[3338]), .B(c3338), .Z(n10016) );
XOR U16695 ( .A(c3339), .B(n10017), .Z(c3340) );
ANDN U16696 ( .B(n10018), .A(n10019), .Z(n10017) );
XOR U16697 ( .A(c3339), .B(b[3339]), .Z(n10018) );
XNOR U16698 ( .A(b[3339]), .B(n10019), .Z(c[3339]) );
XNOR U16699 ( .A(a[3339]), .B(c3339), .Z(n10019) );
XOR U16700 ( .A(c3340), .B(n10020), .Z(c3341) );
ANDN U16701 ( .B(n10021), .A(n10022), .Z(n10020) );
XOR U16702 ( .A(c3340), .B(b[3340]), .Z(n10021) );
XNOR U16703 ( .A(b[3340]), .B(n10022), .Z(c[3340]) );
XNOR U16704 ( .A(a[3340]), .B(c3340), .Z(n10022) );
XOR U16705 ( .A(c3341), .B(n10023), .Z(c3342) );
ANDN U16706 ( .B(n10024), .A(n10025), .Z(n10023) );
XOR U16707 ( .A(c3341), .B(b[3341]), .Z(n10024) );
XNOR U16708 ( .A(b[3341]), .B(n10025), .Z(c[3341]) );
XNOR U16709 ( .A(a[3341]), .B(c3341), .Z(n10025) );
XOR U16710 ( .A(c3342), .B(n10026), .Z(c3343) );
ANDN U16711 ( .B(n10027), .A(n10028), .Z(n10026) );
XOR U16712 ( .A(c3342), .B(b[3342]), .Z(n10027) );
XNOR U16713 ( .A(b[3342]), .B(n10028), .Z(c[3342]) );
XNOR U16714 ( .A(a[3342]), .B(c3342), .Z(n10028) );
XOR U16715 ( .A(c3343), .B(n10029), .Z(c3344) );
ANDN U16716 ( .B(n10030), .A(n10031), .Z(n10029) );
XOR U16717 ( .A(c3343), .B(b[3343]), .Z(n10030) );
XNOR U16718 ( .A(b[3343]), .B(n10031), .Z(c[3343]) );
XNOR U16719 ( .A(a[3343]), .B(c3343), .Z(n10031) );
XOR U16720 ( .A(c3344), .B(n10032), .Z(c3345) );
ANDN U16721 ( .B(n10033), .A(n10034), .Z(n10032) );
XOR U16722 ( .A(c3344), .B(b[3344]), .Z(n10033) );
XNOR U16723 ( .A(b[3344]), .B(n10034), .Z(c[3344]) );
XNOR U16724 ( .A(a[3344]), .B(c3344), .Z(n10034) );
XOR U16725 ( .A(c3345), .B(n10035), .Z(c3346) );
ANDN U16726 ( .B(n10036), .A(n10037), .Z(n10035) );
XOR U16727 ( .A(c3345), .B(b[3345]), .Z(n10036) );
XNOR U16728 ( .A(b[3345]), .B(n10037), .Z(c[3345]) );
XNOR U16729 ( .A(a[3345]), .B(c3345), .Z(n10037) );
XOR U16730 ( .A(c3346), .B(n10038), .Z(c3347) );
ANDN U16731 ( .B(n10039), .A(n10040), .Z(n10038) );
XOR U16732 ( .A(c3346), .B(b[3346]), .Z(n10039) );
XNOR U16733 ( .A(b[3346]), .B(n10040), .Z(c[3346]) );
XNOR U16734 ( .A(a[3346]), .B(c3346), .Z(n10040) );
XOR U16735 ( .A(c3347), .B(n10041), .Z(c3348) );
ANDN U16736 ( .B(n10042), .A(n10043), .Z(n10041) );
XOR U16737 ( .A(c3347), .B(b[3347]), .Z(n10042) );
XNOR U16738 ( .A(b[3347]), .B(n10043), .Z(c[3347]) );
XNOR U16739 ( .A(a[3347]), .B(c3347), .Z(n10043) );
XOR U16740 ( .A(c3348), .B(n10044), .Z(c3349) );
ANDN U16741 ( .B(n10045), .A(n10046), .Z(n10044) );
XOR U16742 ( .A(c3348), .B(b[3348]), .Z(n10045) );
XNOR U16743 ( .A(b[3348]), .B(n10046), .Z(c[3348]) );
XNOR U16744 ( .A(a[3348]), .B(c3348), .Z(n10046) );
XOR U16745 ( .A(c3349), .B(n10047), .Z(c3350) );
ANDN U16746 ( .B(n10048), .A(n10049), .Z(n10047) );
XOR U16747 ( .A(c3349), .B(b[3349]), .Z(n10048) );
XNOR U16748 ( .A(b[3349]), .B(n10049), .Z(c[3349]) );
XNOR U16749 ( .A(a[3349]), .B(c3349), .Z(n10049) );
XOR U16750 ( .A(c3350), .B(n10050), .Z(c3351) );
ANDN U16751 ( .B(n10051), .A(n10052), .Z(n10050) );
XOR U16752 ( .A(c3350), .B(b[3350]), .Z(n10051) );
XNOR U16753 ( .A(b[3350]), .B(n10052), .Z(c[3350]) );
XNOR U16754 ( .A(a[3350]), .B(c3350), .Z(n10052) );
XOR U16755 ( .A(c3351), .B(n10053), .Z(c3352) );
ANDN U16756 ( .B(n10054), .A(n10055), .Z(n10053) );
XOR U16757 ( .A(c3351), .B(b[3351]), .Z(n10054) );
XNOR U16758 ( .A(b[3351]), .B(n10055), .Z(c[3351]) );
XNOR U16759 ( .A(a[3351]), .B(c3351), .Z(n10055) );
XOR U16760 ( .A(c3352), .B(n10056), .Z(c3353) );
ANDN U16761 ( .B(n10057), .A(n10058), .Z(n10056) );
XOR U16762 ( .A(c3352), .B(b[3352]), .Z(n10057) );
XNOR U16763 ( .A(b[3352]), .B(n10058), .Z(c[3352]) );
XNOR U16764 ( .A(a[3352]), .B(c3352), .Z(n10058) );
XOR U16765 ( .A(c3353), .B(n10059), .Z(c3354) );
ANDN U16766 ( .B(n10060), .A(n10061), .Z(n10059) );
XOR U16767 ( .A(c3353), .B(b[3353]), .Z(n10060) );
XNOR U16768 ( .A(b[3353]), .B(n10061), .Z(c[3353]) );
XNOR U16769 ( .A(a[3353]), .B(c3353), .Z(n10061) );
XOR U16770 ( .A(c3354), .B(n10062), .Z(c3355) );
ANDN U16771 ( .B(n10063), .A(n10064), .Z(n10062) );
XOR U16772 ( .A(c3354), .B(b[3354]), .Z(n10063) );
XNOR U16773 ( .A(b[3354]), .B(n10064), .Z(c[3354]) );
XNOR U16774 ( .A(a[3354]), .B(c3354), .Z(n10064) );
XOR U16775 ( .A(c3355), .B(n10065), .Z(c3356) );
ANDN U16776 ( .B(n10066), .A(n10067), .Z(n10065) );
XOR U16777 ( .A(c3355), .B(b[3355]), .Z(n10066) );
XNOR U16778 ( .A(b[3355]), .B(n10067), .Z(c[3355]) );
XNOR U16779 ( .A(a[3355]), .B(c3355), .Z(n10067) );
XOR U16780 ( .A(c3356), .B(n10068), .Z(c3357) );
ANDN U16781 ( .B(n10069), .A(n10070), .Z(n10068) );
XOR U16782 ( .A(c3356), .B(b[3356]), .Z(n10069) );
XNOR U16783 ( .A(b[3356]), .B(n10070), .Z(c[3356]) );
XNOR U16784 ( .A(a[3356]), .B(c3356), .Z(n10070) );
XOR U16785 ( .A(c3357), .B(n10071), .Z(c3358) );
ANDN U16786 ( .B(n10072), .A(n10073), .Z(n10071) );
XOR U16787 ( .A(c3357), .B(b[3357]), .Z(n10072) );
XNOR U16788 ( .A(b[3357]), .B(n10073), .Z(c[3357]) );
XNOR U16789 ( .A(a[3357]), .B(c3357), .Z(n10073) );
XOR U16790 ( .A(c3358), .B(n10074), .Z(c3359) );
ANDN U16791 ( .B(n10075), .A(n10076), .Z(n10074) );
XOR U16792 ( .A(c3358), .B(b[3358]), .Z(n10075) );
XNOR U16793 ( .A(b[3358]), .B(n10076), .Z(c[3358]) );
XNOR U16794 ( .A(a[3358]), .B(c3358), .Z(n10076) );
XOR U16795 ( .A(c3359), .B(n10077), .Z(c3360) );
ANDN U16796 ( .B(n10078), .A(n10079), .Z(n10077) );
XOR U16797 ( .A(c3359), .B(b[3359]), .Z(n10078) );
XNOR U16798 ( .A(b[3359]), .B(n10079), .Z(c[3359]) );
XNOR U16799 ( .A(a[3359]), .B(c3359), .Z(n10079) );
XOR U16800 ( .A(c3360), .B(n10080), .Z(c3361) );
ANDN U16801 ( .B(n10081), .A(n10082), .Z(n10080) );
XOR U16802 ( .A(c3360), .B(b[3360]), .Z(n10081) );
XNOR U16803 ( .A(b[3360]), .B(n10082), .Z(c[3360]) );
XNOR U16804 ( .A(a[3360]), .B(c3360), .Z(n10082) );
XOR U16805 ( .A(c3361), .B(n10083), .Z(c3362) );
ANDN U16806 ( .B(n10084), .A(n10085), .Z(n10083) );
XOR U16807 ( .A(c3361), .B(b[3361]), .Z(n10084) );
XNOR U16808 ( .A(b[3361]), .B(n10085), .Z(c[3361]) );
XNOR U16809 ( .A(a[3361]), .B(c3361), .Z(n10085) );
XOR U16810 ( .A(c3362), .B(n10086), .Z(c3363) );
ANDN U16811 ( .B(n10087), .A(n10088), .Z(n10086) );
XOR U16812 ( .A(c3362), .B(b[3362]), .Z(n10087) );
XNOR U16813 ( .A(b[3362]), .B(n10088), .Z(c[3362]) );
XNOR U16814 ( .A(a[3362]), .B(c3362), .Z(n10088) );
XOR U16815 ( .A(c3363), .B(n10089), .Z(c3364) );
ANDN U16816 ( .B(n10090), .A(n10091), .Z(n10089) );
XOR U16817 ( .A(c3363), .B(b[3363]), .Z(n10090) );
XNOR U16818 ( .A(b[3363]), .B(n10091), .Z(c[3363]) );
XNOR U16819 ( .A(a[3363]), .B(c3363), .Z(n10091) );
XOR U16820 ( .A(c3364), .B(n10092), .Z(c3365) );
ANDN U16821 ( .B(n10093), .A(n10094), .Z(n10092) );
XOR U16822 ( .A(c3364), .B(b[3364]), .Z(n10093) );
XNOR U16823 ( .A(b[3364]), .B(n10094), .Z(c[3364]) );
XNOR U16824 ( .A(a[3364]), .B(c3364), .Z(n10094) );
XOR U16825 ( .A(c3365), .B(n10095), .Z(c3366) );
ANDN U16826 ( .B(n10096), .A(n10097), .Z(n10095) );
XOR U16827 ( .A(c3365), .B(b[3365]), .Z(n10096) );
XNOR U16828 ( .A(b[3365]), .B(n10097), .Z(c[3365]) );
XNOR U16829 ( .A(a[3365]), .B(c3365), .Z(n10097) );
XOR U16830 ( .A(c3366), .B(n10098), .Z(c3367) );
ANDN U16831 ( .B(n10099), .A(n10100), .Z(n10098) );
XOR U16832 ( .A(c3366), .B(b[3366]), .Z(n10099) );
XNOR U16833 ( .A(b[3366]), .B(n10100), .Z(c[3366]) );
XNOR U16834 ( .A(a[3366]), .B(c3366), .Z(n10100) );
XOR U16835 ( .A(c3367), .B(n10101), .Z(c3368) );
ANDN U16836 ( .B(n10102), .A(n10103), .Z(n10101) );
XOR U16837 ( .A(c3367), .B(b[3367]), .Z(n10102) );
XNOR U16838 ( .A(b[3367]), .B(n10103), .Z(c[3367]) );
XNOR U16839 ( .A(a[3367]), .B(c3367), .Z(n10103) );
XOR U16840 ( .A(c3368), .B(n10104), .Z(c3369) );
ANDN U16841 ( .B(n10105), .A(n10106), .Z(n10104) );
XOR U16842 ( .A(c3368), .B(b[3368]), .Z(n10105) );
XNOR U16843 ( .A(b[3368]), .B(n10106), .Z(c[3368]) );
XNOR U16844 ( .A(a[3368]), .B(c3368), .Z(n10106) );
XOR U16845 ( .A(c3369), .B(n10107), .Z(c3370) );
ANDN U16846 ( .B(n10108), .A(n10109), .Z(n10107) );
XOR U16847 ( .A(c3369), .B(b[3369]), .Z(n10108) );
XNOR U16848 ( .A(b[3369]), .B(n10109), .Z(c[3369]) );
XNOR U16849 ( .A(a[3369]), .B(c3369), .Z(n10109) );
XOR U16850 ( .A(c3370), .B(n10110), .Z(c3371) );
ANDN U16851 ( .B(n10111), .A(n10112), .Z(n10110) );
XOR U16852 ( .A(c3370), .B(b[3370]), .Z(n10111) );
XNOR U16853 ( .A(b[3370]), .B(n10112), .Z(c[3370]) );
XNOR U16854 ( .A(a[3370]), .B(c3370), .Z(n10112) );
XOR U16855 ( .A(c3371), .B(n10113), .Z(c3372) );
ANDN U16856 ( .B(n10114), .A(n10115), .Z(n10113) );
XOR U16857 ( .A(c3371), .B(b[3371]), .Z(n10114) );
XNOR U16858 ( .A(b[3371]), .B(n10115), .Z(c[3371]) );
XNOR U16859 ( .A(a[3371]), .B(c3371), .Z(n10115) );
XOR U16860 ( .A(c3372), .B(n10116), .Z(c3373) );
ANDN U16861 ( .B(n10117), .A(n10118), .Z(n10116) );
XOR U16862 ( .A(c3372), .B(b[3372]), .Z(n10117) );
XNOR U16863 ( .A(b[3372]), .B(n10118), .Z(c[3372]) );
XNOR U16864 ( .A(a[3372]), .B(c3372), .Z(n10118) );
XOR U16865 ( .A(c3373), .B(n10119), .Z(c3374) );
ANDN U16866 ( .B(n10120), .A(n10121), .Z(n10119) );
XOR U16867 ( .A(c3373), .B(b[3373]), .Z(n10120) );
XNOR U16868 ( .A(b[3373]), .B(n10121), .Z(c[3373]) );
XNOR U16869 ( .A(a[3373]), .B(c3373), .Z(n10121) );
XOR U16870 ( .A(c3374), .B(n10122), .Z(c3375) );
ANDN U16871 ( .B(n10123), .A(n10124), .Z(n10122) );
XOR U16872 ( .A(c3374), .B(b[3374]), .Z(n10123) );
XNOR U16873 ( .A(b[3374]), .B(n10124), .Z(c[3374]) );
XNOR U16874 ( .A(a[3374]), .B(c3374), .Z(n10124) );
XOR U16875 ( .A(c3375), .B(n10125), .Z(c3376) );
ANDN U16876 ( .B(n10126), .A(n10127), .Z(n10125) );
XOR U16877 ( .A(c3375), .B(b[3375]), .Z(n10126) );
XNOR U16878 ( .A(b[3375]), .B(n10127), .Z(c[3375]) );
XNOR U16879 ( .A(a[3375]), .B(c3375), .Z(n10127) );
XOR U16880 ( .A(c3376), .B(n10128), .Z(c3377) );
ANDN U16881 ( .B(n10129), .A(n10130), .Z(n10128) );
XOR U16882 ( .A(c3376), .B(b[3376]), .Z(n10129) );
XNOR U16883 ( .A(b[3376]), .B(n10130), .Z(c[3376]) );
XNOR U16884 ( .A(a[3376]), .B(c3376), .Z(n10130) );
XOR U16885 ( .A(c3377), .B(n10131), .Z(c3378) );
ANDN U16886 ( .B(n10132), .A(n10133), .Z(n10131) );
XOR U16887 ( .A(c3377), .B(b[3377]), .Z(n10132) );
XNOR U16888 ( .A(b[3377]), .B(n10133), .Z(c[3377]) );
XNOR U16889 ( .A(a[3377]), .B(c3377), .Z(n10133) );
XOR U16890 ( .A(c3378), .B(n10134), .Z(c3379) );
ANDN U16891 ( .B(n10135), .A(n10136), .Z(n10134) );
XOR U16892 ( .A(c3378), .B(b[3378]), .Z(n10135) );
XNOR U16893 ( .A(b[3378]), .B(n10136), .Z(c[3378]) );
XNOR U16894 ( .A(a[3378]), .B(c3378), .Z(n10136) );
XOR U16895 ( .A(c3379), .B(n10137), .Z(c3380) );
ANDN U16896 ( .B(n10138), .A(n10139), .Z(n10137) );
XOR U16897 ( .A(c3379), .B(b[3379]), .Z(n10138) );
XNOR U16898 ( .A(b[3379]), .B(n10139), .Z(c[3379]) );
XNOR U16899 ( .A(a[3379]), .B(c3379), .Z(n10139) );
XOR U16900 ( .A(c3380), .B(n10140), .Z(c3381) );
ANDN U16901 ( .B(n10141), .A(n10142), .Z(n10140) );
XOR U16902 ( .A(c3380), .B(b[3380]), .Z(n10141) );
XNOR U16903 ( .A(b[3380]), .B(n10142), .Z(c[3380]) );
XNOR U16904 ( .A(a[3380]), .B(c3380), .Z(n10142) );
XOR U16905 ( .A(c3381), .B(n10143), .Z(c3382) );
ANDN U16906 ( .B(n10144), .A(n10145), .Z(n10143) );
XOR U16907 ( .A(c3381), .B(b[3381]), .Z(n10144) );
XNOR U16908 ( .A(b[3381]), .B(n10145), .Z(c[3381]) );
XNOR U16909 ( .A(a[3381]), .B(c3381), .Z(n10145) );
XOR U16910 ( .A(c3382), .B(n10146), .Z(c3383) );
ANDN U16911 ( .B(n10147), .A(n10148), .Z(n10146) );
XOR U16912 ( .A(c3382), .B(b[3382]), .Z(n10147) );
XNOR U16913 ( .A(b[3382]), .B(n10148), .Z(c[3382]) );
XNOR U16914 ( .A(a[3382]), .B(c3382), .Z(n10148) );
XOR U16915 ( .A(c3383), .B(n10149), .Z(c3384) );
ANDN U16916 ( .B(n10150), .A(n10151), .Z(n10149) );
XOR U16917 ( .A(c3383), .B(b[3383]), .Z(n10150) );
XNOR U16918 ( .A(b[3383]), .B(n10151), .Z(c[3383]) );
XNOR U16919 ( .A(a[3383]), .B(c3383), .Z(n10151) );
XOR U16920 ( .A(c3384), .B(n10152), .Z(c3385) );
ANDN U16921 ( .B(n10153), .A(n10154), .Z(n10152) );
XOR U16922 ( .A(c3384), .B(b[3384]), .Z(n10153) );
XNOR U16923 ( .A(b[3384]), .B(n10154), .Z(c[3384]) );
XNOR U16924 ( .A(a[3384]), .B(c3384), .Z(n10154) );
XOR U16925 ( .A(c3385), .B(n10155), .Z(c3386) );
ANDN U16926 ( .B(n10156), .A(n10157), .Z(n10155) );
XOR U16927 ( .A(c3385), .B(b[3385]), .Z(n10156) );
XNOR U16928 ( .A(b[3385]), .B(n10157), .Z(c[3385]) );
XNOR U16929 ( .A(a[3385]), .B(c3385), .Z(n10157) );
XOR U16930 ( .A(c3386), .B(n10158), .Z(c3387) );
ANDN U16931 ( .B(n10159), .A(n10160), .Z(n10158) );
XOR U16932 ( .A(c3386), .B(b[3386]), .Z(n10159) );
XNOR U16933 ( .A(b[3386]), .B(n10160), .Z(c[3386]) );
XNOR U16934 ( .A(a[3386]), .B(c3386), .Z(n10160) );
XOR U16935 ( .A(c3387), .B(n10161), .Z(c3388) );
ANDN U16936 ( .B(n10162), .A(n10163), .Z(n10161) );
XOR U16937 ( .A(c3387), .B(b[3387]), .Z(n10162) );
XNOR U16938 ( .A(b[3387]), .B(n10163), .Z(c[3387]) );
XNOR U16939 ( .A(a[3387]), .B(c3387), .Z(n10163) );
XOR U16940 ( .A(c3388), .B(n10164), .Z(c3389) );
ANDN U16941 ( .B(n10165), .A(n10166), .Z(n10164) );
XOR U16942 ( .A(c3388), .B(b[3388]), .Z(n10165) );
XNOR U16943 ( .A(b[3388]), .B(n10166), .Z(c[3388]) );
XNOR U16944 ( .A(a[3388]), .B(c3388), .Z(n10166) );
XOR U16945 ( .A(c3389), .B(n10167), .Z(c3390) );
ANDN U16946 ( .B(n10168), .A(n10169), .Z(n10167) );
XOR U16947 ( .A(c3389), .B(b[3389]), .Z(n10168) );
XNOR U16948 ( .A(b[3389]), .B(n10169), .Z(c[3389]) );
XNOR U16949 ( .A(a[3389]), .B(c3389), .Z(n10169) );
XOR U16950 ( .A(c3390), .B(n10170), .Z(c3391) );
ANDN U16951 ( .B(n10171), .A(n10172), .Z(n10170) );
XOR U16952 ( .A(c3390), .B(b[3390]), .Z(n10171) );
XNOR U16953 ( .A(b[3390]), .B(n10172), .Z(c[3390]) );
XNOR U16954 ( .A(a[3390]), .B(c3390), .Z(n10172) );
XOR U16955 ( .A(c3391), .B(n10173), .Z(c3392) );
ANDN U16956 ( .B(n10174), .A(n10175), .Z(n10173) );
XOR U16957 ( .A(c3391), .B(b[3391]), .Z(n10174) );
XNOR U16958 ( .A(b[3391]), .B(n10175), .Z(c[3391]) );
XNOR U16959 ( .A(a[3391]), .B(c3391), .Z(n10175) );
XOR U16960 ( .A(c3392), .B(n10176), .Z(c3393) );
ANDN U16961 ( .B(n10177), .A(n10178), .Z(n10176) );
XOR U16962 ( .A(c3392), .B(b[3392]), .Z(n10177) );
XNOR U16963 ( .A(b[3392]), .B(n10178), .Z(c[3392]) );
XNOR U16964 ( .A(a[3392]), .B(c3392), .Z(n10178) );
XOR U16965 ( .A(c3393), .B(n10179), .Z(c3394) );
ANDN U16966 ( .B(n10180), .A(n10181), .Z(n10179) );
XOR U16967 ( .A(c3393), .B(b[3393]), .Z(n10180) );
XNOR U16968 ( .A(b[3393]), .B(n10181), .Z(c[3393]) );
XNOR U16969 ( .A(a[3393]), .B(c3393), .Z(n10181) );
XOR U16970 ( .A(c3394), .B(n10182), .Z(c3395) );
ANDN U16971 ( .B(n10183), .A(n10184), .Z(n10182) );
XOR U16972 ( .A(c3394), .B(b[3394]), .Z(n10183) );
XNOR U16973 ( .A(b[3394]), .B(n10184), .Z(c[3394]) );
XNOR U16974 ( .A(a[3394]), .B(c3394), .Z(n10184) );
XOR U16975 ( .A(c3395), .B(n10185), .Z(c3396) );
ANDN U16976 ( .B(n10186), .A(n10187), .Z(n10185) );
XOR U16977 ( .A(c3395), .B(b[3395]), .Z(n10186) );
XNOR U16978 ( .A(b[3395]), .B(n10187), .Z(c[3395]) );
XNOR U16979 ( .A(a[3395]), .B(c3395), .Z(n10187) );
XOR U16980 ( .A(c3396), .B(n10188), .Z(c3397) );
ANDN U16981 ( .B(n10189), .A(n10190), .Z(n10188) );
XOR U16982 ( .A(c3396), .B(b[3396]), .Z(n10189) );
XNOR U16983 ( .A(b[3396]), .B(n10190), .Z(c[3396]) );
XNOR U16984 ( .A(a[3396]), .B(c3396), .Z(n10190) );
XOR U16985 ( .A(c3397), .B(n10191), .Z(c3398) );
ANDN U16986 ( .B(n10192), .A(n10193), .Z(n10191) );
XOR U16987 ( .A(c3397), .B(b[3397]), .Z(n10192) );
XNOR U16988 ( .A(b[3397]), .B(n10193), .Z(c[3397]) );
XNOR U16989 ( .A(a[3397]), .B(c3397), .Z(n10193) );
XOR U16990 ( .A(c3398), .B(n10194), .Z(c3399) );
ANDN U16991 ( .B(n10195), .A(n10196), .Z(n10194) );
XOR U16992 ( .A(c3398), .B(b[3398]), .Z(n10195) );
XNOR U16993 ( .A(b[3398]), .B(n10196), .Z(c[3398]) );
XNOR U16994 ( .A(a[3398]), .B(c3398), .Z(n10196) );
XOR U16995 ( .A(c3399), .B(n10197), .Z(c3400) );
ANDN U16996 ( .B(n10198), .A(n10199), .Z(n10197) );
XOR U16997 ( .A(c3399), .B(b[3399]), .Z(n10198) );
XNOR U16998 ( .A(b[3399]), .B(n10199), .Z(c[3399]) );
XNOR U16999 ( .A(a[3399]), .B(c3399), .Z(n10199) );
XOR U17000 ( .A(c3400), .B(n10200), .Z(c3401) );
ANDN U17001 ( .B(n10201), .A(n10202), .Z(n10200) );
XOR U17002 ( .A(c3400), .B(b[3400]), .Z(n10201) );
XNOR U17003 ( .A(b[3400]), .B(n10202), .Z(c[3400]) );
XNOR U17004 ( .A(a[3400]), .B(c3400), .Z(n10202) );
XOR U17005 ( .A(c3401), .B(n10203), .Z(c3402) );
ANDN U17006 ( .B(n10204), .A(n10205), .Z(n10203) );
XOR U17007 ( .A(c3401), .B(b[3401]), .Z(n10204) );
XNOR U17008 ( .A(b[3401]), .B(n10205), .Z(c[3401]) );
XNOR U17009 ( .A(a[3401]), .B(c3401), .Z(n10205) );
XOR U17010 ( .A(c3402), .B(n10206), .Z(c3403) );
ANDN U17011 ( .B(n10207), .A(n10208), .Z(n10206) );
XOR U17012 ( .A(c3402), .B(b[3402]), .Z(n10207) );
XNOR U17013 ( .A(b[3402]), .B(n10208), .Z(c[3402]) );
XNOR U17014 ( .A(a[3402]), .B(c3402), .Z(n10208) );
XOR U17015 ( .A(c3403), .B(n10209), .Z(c3404) );
ANDN U17016 ( .B(n10210), .A(n10211), .Z(n10209) );
XOR U17017 ( .A(c3403), .B(b[3403]), .Z(n10210) );
XNOR U17018 ( .A(b[3403]), .B(n10211), .Z(c[3403]) );
XNOR U17019 ( .A(a[3403]), .B(c3403), .Z(n10211) );
XOR U17020 ( .A(c3404), .B(n10212), .Z(c3405) );
ANDN U17021 ( .B(n10213), .A(n10214), .Z(n10212) );
XOR U17022 ( .A(c3404), .B(b[3404]), .Z(n10213) );
XNOR U17023 ( .A(b[3404]), .B(n10214), .Z(c[3404]) );
XNOR U17024 ( .A(a[3404]), .B(c3404), .Z(n10214) );
XOR U17025 ( .A(c3405), .B(n10215), .Z(c3406) );
ANDN U17026 ( .B(n10216), .A(n10217), .Z(n10215) );
XOR U17027 ( .A(c3405), .B(b[3405]), .Z(n10216) );
XNOR U17028 ( .A(b[3405]), .B(n10217), .Z(c[3405]) );
XNOR U17029 ( .A(a[3405]), .B(c3405), .Z(n10217) );
XOR U17030 ( .A(c3406), .B(n10218), .Z(c3407) );
ANDN U17031 ( .B(n10219), .A(n10220), .Z(n10218) );
XOR U17032 ( .A(c3406), .B(b[3406]), .Z(n10219) );
XNOR U17033 ( .A(b[3406]), .B(n10220), .Z(c[3406]) );
XNOR U17034 ( .A(a[3406]), .B(c3406), .Z(n10220) );
XOR U17035 ( .A(c3407), .B(n10221), .Z(c3408) );
ANDN U17036 ( .B(n10222), .A(n10223), .Z(n10221) );
XOR U17037 ( .A(c3407), .B(b[3407]), .Z(n10222) );
XNOR U17038 ( .A(b[3407]), .B(n10223), .Z(c[3407]) );
XNOR U17039 ( .A(a[3407]), .B(c3407), .Z(n10223) );
XOR U17040 ( .A(c3408), .B(n10224), .Z(c3409) );
ANDN U17041 ( .B(n10225), .A(n10226), .Z(n10224) );
XOR U17042 ( .A(c3408), .B(b[3408]), .Z(n10225) );
XNOR U17043 ( .A(b[3408]), .B(n10226), .Z(c[3408]) );
XNOR U17044 ( .A(a[3408]), .B(c3408), .Z(n10226) );
XOR U17045 ( .A(c3409), .B(n10227), .Z(c3410) );
ANDN U17046 ( .B(n10228), .A(n10229), .Z(n10227) );
XOR U17047 ( .A(c3409), .B(b[3409]), .Z(n10228) );
XNOR U17048 ( .A(b[3409]), .B(n10229), .Z(c[3409]) );
XNOR U17049 ( .A(a[3409]), .B(c3409), .Z(n10229) );
XOR U17050 ( .A(c3410), .B(n10230), .Z(c3411) );
ANDN U17051 ( .B(n10231), .A(n10232), .Z(n10230) );
XOR U17052 ( .A(c3410), .B(b[3410]), .Z(n10231) );
XNOR U17053 ( .A(b[3410]), .B(n10232), .Z(c[3410]) );
XNOR U17054 ( .A(a[3410]), .B(c3410), .Z(n10232) );
XOR U17055 ( .A(c3411), .B(n10233), .Z(c3412) );
ANDN U17056 ( .B(n10234), .A(n10235), .Z(n10233) );
XOR U17057 ( .A(c3411), .B(b[3411]), .Z(n10234) );
XNOR U17058 ( .A(b[3411]), .B(n10235), .Z(c[3411]) );
XNOR U17059 ( .A(a[3411]), .B(c3411), .Z(n10235) );
XOR U17060 ( .A(c3412), .B(n10236), .Z(c3413) );
ANDN U17061 ( .B(n10237), .A(n10238), .Z(n10236) );
XOR U17062 ( .A(c3412), .B(b[3412]), .Z(n10237) );
XNOR U17063 ( .A(b[3412]), .B(n10238), .Z(c[3412]) );
XNOR U17064 ( .A(a[3412]), .B(c3412), .Z(n10238) );
XOR U17065 ( .A(c3413), .B(n10239), .Z(c3414) );
ANDN U17066 ( .B(n10240), .A(n10241), .Z(n10239) );
XOR U17067 ( .A(c3413), .B(b[3413]), .Z(n10240) );
XNOR U17068 ( .A(b[3413]), .B(n10241), .Z(c[3413]) );
XNOR U17069 ( .A(a[3413]), .B(c3413), .Z(n10241) );
XOR U17070 ( .A(c3414), .B(n10242), .Z(c3415) );
ANDN U17071 ( .B(n10243), .A(n10244), .Z(n10242) );
XOR U17072 ( .A(c3414), .B(b[3414]), .Z(n10243) );
XNOR U17073 ( .A(b[3414]), .B(n10244), .Z(c[3414]) );
XNOR U17074 ( .A(a[3414]), .B(c3414), .Z(n10244) );
XOR U17075 ( .A(c3415), .B(n10245), .Z(c3416) );
ANDN U17076 ( .B(n10246), .A(n10247), .Z(n10245) );
XOR U17077 ( .A(c3415), .B(b[3415]), .Z(n10246) );
XNOR U17078 ( .A(b[3415]), .B(n10247), .Z(c[3415]) );
XNOR U17079 ( .A(a[3415]), .B(c3415), .Z(n10247) );
XOR U17080 ( .A(c3416), .B(n10248), .Z(c3417) );
ANDN U17081 ( .B(n10249), .A(n10250), .Z(n10248) );
XOR U17082 ( .A(c3416), .B(b[3416]), .Z(n10249) );
XNOR U17083 ( .A(b[3416]), .B(n10250), .Z(c[3416]) );
XNOR U17084 ( .A(a[3416]), .B(c3416), .Z(n10250) );
XOR U17085 ( .A(c3417), .B(n10251), .Z(c3418) );
ANDN U17086 ( .B(n10252), .A(n10253), .Z(n10251) );
XOR U17087 ( .A(c3417), .B(b[3417]), .Z(n10252) );
XNOR U17088 ( .A(b[3417]), .B(n10253), .Z(c[3417]) );
XNOR U17089 ( .A(a[3417]), .B(c3417), .Z(n10253) );
XOR U17090 ( .A(c3418), .B(n10254), .Z(c3419) );
ANDN U17091 ( .B(n10255), .A(n10256), .Z(n10254) );
XOR U17092 ( .A(c3418), .B(b[3418]), .Z(n10255) );
XNOR U17093 ( .A(b[3418]), .B(n10256), .Z(c[3418]) );
XNOR U17094 ( .A(a[3418]), .B(c3418), .Z(n10256) );
XOR U17095 ( .A(c3419), .B(n10257), .Z(c3420) );
ANDN U17096 ( .B(n10258), .A(n10259), .Z(n10257) );
XOR U17097 ( .A(c3419), .B(b[3419]), .Z(n10258) );
XNOR U17098 ( .A(b[3419]), .B(n10259), .Z(c[3419]) );
XNOR U17099 ( .A(a[3419]), .B(c3419), .Z(n10259) );
XOR U17100 ( .A(c3420), .B(n10260), .Z(c3421) );
ANDN U17101 ( .B(n10261), .A(n10262), .Z(n10260) );
XOR U17102 ( .A(c3420), .B(b[3420]), .Z(n10261) );
XNOR U17103 ( .A(b[3420]), .B(n10262), .Z(c[3420]) );
XNOR U17104 ( .A(a[3420]), .B(c3420), .Z(n10262) );
XOR U17105 ( .A(c3421), .B(n10263), .Z(c3422) );
ANDN U17106 ( .B(n10264), .A(n10265), .Z(n10263) );
XOR U17107 ( .A(c3421), .B(b[3421]), .Z(n10264) );
XNOR U17108 ( .A(b[3421]), .B(n10265), .Z(c[3421]) );
XNOR U17109 ( .A(a[3421]), .B(c3421), .Z(n10265) );
XOR U17110 ( .A(c3422), .B(n10266), .Z(c3423) );
ANDN U17111 ( .B(n10267), .A(n10268), .Z(n10266) );
XOR U17112 ( .A(c3422), .B(b[3422]), .Z(n10267) );
XNOR U17113 ( .A(b[3422]), .B(n10268), .Z(c[3422]) );
XNOR U17114 ( .A(a[3422]), .B(c3422), .Z(n10268) );
XOR U17115 ( .A(c3423), .B(n10269), .Z(c3424) );
ANDN U17116 ( .B(n10270), .A(n10271), .Z(n10269) );
XOR U17117 ( .A(c3423), .B(b[3423]), .Z(n10270) );
XNOR U17118 ( .A(b[3423]), .B(n10271), .Z(c[3423]) );
XNOR U17119 ( .A(a[3423]), .B(c3423), .Z(n10271) );
XOR U17120 ( .A(c3424), .B(n10272), .Z(c3425) );
ANDN U17121 ( .B(n10273), .A(n10274), .Z(n10272) );
XOR U17122 ( .A(c3424), .B(b[3424]), .Z(n10273) );
XNOR U17123 ( .A(b[3424]), .B(n10274), .Z(c[3424]) );
XNOR U17124 ( .A(a[3424]), .B(c3424), .Z(n10274) );
XOR U17125 ( .A(c3425), .B(n10275), .Z(c3426) );
ANDN U17126 ( .B(n10276), .A(n10277), .Z(n10275) );
XOR U17127 ( .A(c3425), .B(b[3425]), .Z(n10276) );
XNOR U17128 ( .A(b[3425]), .B(n10277), .Z(c[3425]) );
XNOR U17129 ( .A(a[3425]), .B(c3425), .Z(n10277) );
XOR U17130 ( .A(c3426), .B(n10278), .Z(c3427) );
ANDN U17131 ( .B(n10279), .A(n10280), .Z(n10278) );
XOR U17132 ( .A(c3426), .B(b[3426]), .Z(n10279) );
XNOR U17133 ( .A(b[3426]), .B(n10280), .Z(c[3426]) );
XNOR U17134 ( .A(a[3426]), .B(c3426), .Z(n10280) );
XOR U17135 ( .A(c3427), .B(n10281), .Z(c3428) );
ANDN U17136 ( .B(n10282), .A(n10283), .Z(n10281) );
XOR U17137 ( .A(c3427), .B(b[3427]), .Z(n10282) );
XNOR U17138 ( .A(b[3427]), .B(n10283), .Z(c[3427]) );
XNOR U17139 ( .A(a[3427]), .B(c3427), .Z(n10283) );
XOR U17140 ( .A(c3428), .B(n10284), .Z(c3429) );
ANDN U17141 ( .B(n10285), .A(n10286), .Z(n10284) );
XOR U17142 ( .A(c3428), .B(b[3428]), .Z(n10285) );
XNOR U17143 ( .A(b[3428]), .B(n10286), .Z(c[3428]) );
XNOR U17144 ( .A(a[3428]), .B(c3428), .Z(n10286) );
XOR U17145 ( .A(c3429), .B(n10287), .Z(c3430) );
ANDN U17146 ( .B(n10288), .A(n10289), .Z(n10287) );
XOR U17147 ( .A(c3429), .B(b[3429]), .Z(n10288) );
XNOR U17148 ( .A(b[3429]), .B(n10289), .Z(c[3429]) );
XNOR U17149 ( .A(a[3429]), .B(c3429), .Z(n10289) );
XOR U17150 ( .A(c3430), .B(n10290), .Z(c3431) );
ANDN U17151 ( .B(n10291), .A(n10292), .Z(n10290) );
XOR U17152 ( .A(c3430), .B(b[3430]), .Z(n10291) );
XNOR U17153 ( .A(b[3430]), .B(n10292), .Z(c[3430]) );
XNOR U17154 ( .A(a[3430]), .B(c3430), .Z(n10292) );
XOR U17155 ( .A(c3431), .B(n10293), .Z(c3432) );
ANDN U17156 ( .B(n10294), .A(n10295), .Z(n10293) );
XOR U17157 ( .A(c3431), .B(b[3431]), .Z(n10294) );
XNOR U17158 ( .A(b[3431]), .B(n10295), .Z(c[3431]) );
XNOR U17159 ( .A(a[3431]), .B(c3431), .Z(n10295) );
XOR U17160 ( .A(c3432), .B(n10296), .Z(c3433) );
ANDN U17161 ( .B(n10297), .A(n10298), .Z(n10296) );
XOR U17162 ( .A(c3432), .B(b[3432]), .Z(n10297) );
XNOR U17163 ( .A(b[3432]), .B(n10298), .Z(c[3432]) );
XNOR U17164 ( .A(a[3432]), .B(c3432), .Z(n10298) );
XOR U17165 ( .A(c3433), .B(n10299), .Z(c3434) );
ANDN U17166 ( .B(n10300), .A(n10301), .Z(n10299) );
XOR U17167 ( .A(c3433), .B(b[3433]), .Z(n10300) );
XNOR U17168 ( .A(b[3433]), .B(n10301), .Z(c[3433]) );
XNOR U17169 ( .A(a[3433]), .B(c3433), .Z(n10301) );
XOR U17170 ( .A(c3434), .B(n10302), .Z(c3435) );
ANDN U17171 ( .B(n10303), .A(n10304), .Z(n10302) );
XOR U17172 ( .A(c3434), .B(b[3434]), .Z(n10303) );
XNOR U17173 ( .A(b[3434]), .B(n10304), .Z(c[3434]) );
XNOR U17174 ( .A(a[3434]), .B(c3434), .Z(n10304) );
XOR U17175 ( .A(c3435), .B(n10305), .Z(c3436) );
ANDN U17176 ( .B(n10306), .A(n10307), .Z(n10305) );
XOR U17177 ( .A(c3435), .B(b[3435]), .Z(n10306) );
XNOR U17178 ( .A(b[3435]), .B(n10307), .Z(c[3435]) );
XNOR U17179 ( .A(a[3435]), .B(c3435), .Z(n10307) );
XOR U17180 ( .A(c3436), .B(n10308), .Z(c3437) );
ANDN U17181 ( .B(n10309), .A(n10310), .Z(n10308) );
XOR U17182 ( .A(c3436), .B(b[3436]), .Z(n10309) );
XNOR U17183 ( .A(b[3436]), .B(n10310), .Z(c[3436]) );
XNOR U17184 ( .A(a[3436]), .B(c3436), .Z(n10310) );
XOR U17185 ( .A(c3437), .B(n10311), .Z(c3438) );
ANDN U17186 ( .B(n10312), .A(n10313), .Z(n10311) );
XOR U17187 ( .A(c3437), .B(b[3437]), .Z(n10312) );
XNOR U17188 ( .A(b[3437]), .B(n10313), .Z(c[3437]) );
XNOR U17189 ( .A(a[3437]), .B(c3437), .Z(n10313) );
XOR U17190 ( .A(c3438), .B(n10314), .Z(c3439) );
ANDN U17191 ( .B(n10315), .A(n10316), .Z(n10314) );
XOR U17192 ( .A(c3438), .B(b[3438]), .Z(n10315) );
XNOR U17193 ( .A(b[3438]), .B(n10316), .Z(c[3438]) );
XNOR U17194 ( .A(a[3438]), .B(c3438), .Z(n10316) );
XOR U17195 ( .A(c3439), .B(n10317), .Z(c3440) );
ANDN U17196 ( .B(n10318), .A(n10319), .Z(n10317) );
XOR U17197 ( .A(c3439), .B(b[3439]), .Z(n10318) );
XNOR U17198 ( .A(b[3439]), .B(n10319), .Z(c[3439]) );
XNOR U17199 ( .A(a[3439]), .B(c3439), .Z(n10319) );
XOR U17200 ( .A(c3440), .B(n10320), .Z(c3441) );
ANDN U17201 ( .B(n10321), .A(n10322), .Z(n10320) );
XOR U17202 ( .A(c3440), .B(b[3440]), .Z(n10321) );
XNOR U17203 ( .A(b[3440]), .B(n10322), .Z(c[3440]) );
XNOR U17204 ( .A(a[3440]), .B(c3440), .Z(n10322) );
XOR U17205 ( .A(c3441), .B(n10323), .Z(c3442) );
ANDN U17206 ( .B(n10324), .A(n10325), .Z(n10323) );
XOR U17207 ( .A(c3441), .B(b[3441]), .Z(n10324) );
XNOR U17208 ( .A(b[3441]), .B(n10325), .Z(c[3441]) );
XNOR U17209 ( .A(a[3441]), .B(c3441), .Z(n10325) );
XOR U17210 ( .A(c3442), .B(n10326), .Z(c3443) );
ANDN U17211 ( .B(n10327), .A(n10328), .Z(n10326) );
XOR U17212 ( .A(c3442), .B(b[3442]), .Z(n10327) );
XNOR U17213 ( .A(b[3442]), .B(n10328), .Z(c[3442]) );
XNOR U17214 ( .A(a[3442]), .B(c3442), .Z(n10328) );
XOR U17215 ( .A(c3443), .B(n10329), .Z(c3444) );
ANDN U17216 ( .B(n10330), .A(n10331), .Z(n10329) );
XOR U17217 ( .A(c3443), .B(b[3443]), .Z(n10330) );
XNOR U17218 ( .A(b[3443]), .B(n10331), .Z(c[3443]) );
XNOR U17219 ( .A(a[3443]), .B(c3443), .Z(n10331) );
XOR U17220 ( .A(c3444), .B(n10332), .Z(c3445) );
ANDN U17221 ( .B(n10333), .A(n10334), .Z(n10332) );
XOR U17222 ( .A(c3444), .B(b[3444]), .Z(n10333) );
XNOR U17223 ( .A(b[3444]), .B(n10334), .Z(c[3444]) );
XNOR U17224 ( .A(a[3444]), .B(c3444), .Z(n10334) );
XOR U17225 ( .A(c3445), .B(n10335), .Z(c3446) );
ANDN U17226 ( .B(n10336), .A(n10337), .Z(n10335) );
XOR U17227 ( .A(c3445), .B(b[3445]), .Z(n10336) );
XNOR U17228 ( .A(b[3445]), .B(n10337), .Z(c[3445]) );
XNOR U17229 ( .A(a[3445]), .B(c3445), .Z(n10337) );
XOR U17230 ( .A(c3446), .B(n10338), .Z(c3447) );
ANDN U17231 ( .B(n10339), .A(n10340), .Z(n10338) );
XOR U17232 ( .A(c3446), .B(b[3446]), .Z(n10339) );
XNOR U17233 ( .A(b[3446]), .B(n10340), .Z(c[3446]) );
XNOR U17234 ( .A(a[3446]), .B(c3446), .Z(n10340) );
XOR U17235 ( .A(c3447), .B(n10341), .Z(c3448) );
ANDN U17236 ( .B(n10342), .A(n10343), .Z(n10341) );
XOR U17237 ( .A(c3447), .B(b[3447]), .Z(n10342) );
XNOR U17238 ( .A(b[3447]), .B(n10343), .Z(c[3447]) );
XNOR U17239 ( .A(a[3447]), .B(c3447), .Z(n10343) );
XOR U17240 ( .A(c3448), .B(n10344), .Z(c3449) );
ANDN U17241 ( .B(n10345), .A(n10346), .Z(n10344) );
XOR U17242 ( .A(c3448), .B(b[3448]), .Z(n10345) );
XNOR U17243 ( .A(b[3448]), .B(n10346), .Z(c[3448]) );
XNOR U17244 ( .A(a[3448]), .B(c3448), .Z(n10346) );
XOR U17245 ( .A(c3449), .B(n10347), .Z(c3450) );
ANDN U17246 ( .B(n10348), .A(n10349), .Z(n10347) );
XOR U17247 ( .A(c3449), .B(b[3449]), .Z(n10348) );
XNOR U17248 ( .A(b[3449]), .B(n10349), .Z(c[3449]) );
XNOR U17249 ( .A(a[3449]), .B(c3449), .Z(n10349) );
XOR U17250 ( .A(c3450), .B(n10350), .Z(c3451) );
ANDN U17251 ( .B(n10351), .A(n10352), .Z(n10350) );
XOR U17252 ( .A(c3450), .B(b[3450]), .Z(n10351) );
XNOR U17253 ( .A(b[3450]), .B(n10352), .Z(c[3450]) );
XNOR U17254 ( .A(a[3450]), .B(c3450), .Z(n10352) );
XOR U17255 ( .A(c3451), .B(n10353), .Z(c3452) );
ANDN U17256 ( .B(n10354), .A(n10355), .Z(n10353) );
XOR U17257 ( .A(c3451), .B(b[3451]), .Z(n10354) );
XNOR U17258 ( .A(b[3451]), .B(n10355), .Z(c[3451]) );
XNOR U17259 ( .A(a[3451]), .B(c3451), .Z(n10355) );
XOR U17260 ( .A(c3452), .B(n10356), .Z(c3453) );
ANDN U17261 ( .B(n10357), .A(n10358), .Z(n10356) );
XOR U17262 ( .A(c3452), .B(b[3452]), .Z(n10357) );
XNOR U17263 ( .A(b[3452]), .B(n10358), .Z(c[3452]) );
XNOR U17264 ( .A(a[3452]), .B(c3452), .Z(n10358) );
XOR U17265 ( .A(c3453), .B(n10359), .Z(c3454) );
ANDN U17266 ( .B(n10360), .A(n10361), .Z(n10359) );
XOR U17267 ( .A(c3453), .B(b[3453]), .Z(n10360) );
XNOR U17268 ( .A(b[3453]), .B(n10361), .Z(c[3453]) );
XNOR U17269 ( .A(a[3453]), .B(c3453), .Z(n10361) );
XOR U17270 ( .A(c3454), .B(n10362), .Z(c3455) );
ANDN U17271 ( .B(n10363), .A(n10364), .Z(n10362) );
XOR U17272 ( .A(c3454), .B(b[3454]), .Z(n10363) );
XNOR U17273 ( .A(b[3454]), .B(n10364), .Z(c[3454]) );
XNOR U17274 ( .A(a[3454]), .B(c3454), .Z(n10364) );
XOR U17275 ( .A(c3455), .B(n10365), .Z(c3456) );
ANDN U17276 ( .B(n10366), .A(n10367), .Z(n10365) );
XOR U17277 ( .A(c3455), .B(b[3455]), .Z(n10366) );
XNOR U17278 ( .A(b[3455]), .B(n10367), .Z(c[3455]) );
XNOR U17279 ( .A(a[3455]), .B(c3455), .Z(n10367) );
XOR U17280 ( .A(c3456), .B(n10368), .Z(c3457) );
ANDN U17281 ( .B(n10369), .A(n10370), .Z(n10368) );
XOR U17282 ( .A(c3456), .B(b[3456]), .Z(n10369) );
XNOR U17283 ( .A(b[3456]), .B(n10370), .Z(c[3456]) );
XNOR U17284 ( .A(a[3456]), .B(c3456), .Z(n10370) );
XOR U17285 ( .A(c3457), .B(n10371), .Z(c3458) );
ANDN U17286 ( .B(n10372), .A(n10373), .Z(n10371) );
XOR U17287 ( .A(c3457), .B(b[3457]), .Z(n10372) );
XNOR U17288 ( .A(b[3457]), .B(n10373), .Z(c[3457]) );
XNOR U17289 ( .A(a[3457]), .B(c3457), .Z(n10373) );
XOR U17290 ( .A(c3458), .B(n10374), .Z(c3459) );
ANDN U17291 ( .B(n10375), .A(n10376), .Z(n10374) );
XOR U17292 ( .A(c3458), .B(b[3458]), .Z(n10375) );
XNOR U17293 ( .A(b[3458]), .B(n10376), .Z(c[3458]) );
XNOR U17294 ( .A(a[3458]), .B(c3458), .Z(n10376) );
XOR U17295 ( .A(c3459), .B(n10377), .Z(c3460) );
ANDN U17296 ( .B(n10378), .A(n10379), .Z(n10377) );
XOR U17297 ( .A(c3459), .B(b[3459]), .Z(n10378) );
XNOR U17298 ( .A(b[3459]), .B(n10379), .Z(c[3459]) );
XNOR U17299 ( .A(a[3459]), .B(c3459), .Z(n10379) );
XOR U17300 ( .A(c3460), .B(n10380), .Z(c3461) );
ANDN U17301 ( .B(n10381), .A(n10382), .Z(n10380) );
XOR U17302 ( .A(c3460), .B(b[3460]), .Z(n10381) );
XNOR U17303 ( .A(b[3460]), .B(n10382), .Z(c[3460]) );
XNOR U17304 ( .A(a[3460]), .B(c3460), .Z(n10382) );
XOR U17305 ( .A(c3461), .B(n10383), .Z(c3462) );
ANDN U17306 ( .B(n10384), .A(n10385), .Z(n10383) );
XOR U17307 ( .A(c3461), .B(b[3461]), .Z(n10384) );
XNOR U17308 ( .A(b[3461]), .B(n10385), .Z(c[3461]) );
XNOR U17309 ( .A(a[3461]), .B(c3461), .Z(n10385) );
XOR U17310 ( .A(c3462), .B(n10386), .Z(c3463) );
ANDN U17311 ( .B(n10387), .A(n10388), .Z(n10386) );
XOR U17312 ( .A(c3462), .B(b[3462]), .Z(n10387) );
XNOR U17313 ( .A(b[3462]), .B(n10388), .Z(c[3462]) );
XNOR U17314 ( .A(a[3462]), .B(c3462), .Z(n10388) );
XOR U17315 ( .A(c3463), .B(n10389), .Z(c3464) );
ANDN U17316 ( .B(n10390), .A(n10391), .Z(n10389) );
XOR U17317 ( .A(c3463), .B(b[3463]), .Z(n10390) );
XNOR U17318 ( .A(b[3463]), .B(n10391), .Z(c[3463]) );
XNOR U17319 ( .A(a[3463]), .B(c3463), .Z(n10391) );
XOR U17320 ( .A(c3464), .B(n10392), .Z(c3465) );
ANDN U17321 ( .B(n10393), .A(n10394), .Z(n10392) );
XOR U17322 ( .A(c3464), .B(b[3464]), .Z(n10393) );
XNOR U17323 ( .A(b[3464]), .B(n10394), .Z(c[3464]) );
XNOR U17324 ( .A(a[3464]), .B(c3464), .Z(n10394) );
XOR U17325 ( .A(c3465), .B(n10395), .Z(c3466) );
ANDN U17326 ( .B(n10396), .A(n10397), .Z(n10395) );
XOR U17327 ( .A(c3465), .B(b[3465]), .Z(n10396) );
XNOR U17328 ( .A(b[3465]), .B(n10397), .Z(c[3465]) );
XNOR U17329 ( .A(a[3465]), .B(c3465), .Z(n10397) );
XOR U17330 ( .A(c3466), .B(n10398), .Z(c3467) );
ANDN U17331 ( .B(n10399), .A(n10400), .Z(n10398) );
XOR U17332 ( .A(c3466), .B(b[3466]), .Z(n10399) );
XNOR U17333 ( .A(b[3466]), .B(n10400), .Z(c[3466]) );
XNOR U17334 ( .A(a[3466]), .B(c3466), .Z(n10400) );
XOR U17335 ( .A(c3467), .B(n10401), .Z(c3468) );
ANDN U17336 ( .B(n10402), .A(n10403), .Z(n10401) );
XOR U17337 ( .A(c3467), .B(b[3467]), .Z(n10402) );
XNOR U17338 ( .A(b[3467]), .B(n10403), .Z(c[3467]) );
XNOR U17339 ( .A(a[3467]), .B(c3467), .Z(n10403) );
XOR U17340 ( .A(c3468), .B(n10404), .Z(c3469) );
ANDN U17341 ( .B(n10405), .A(n10406), .Z(n10404) );
XOR U17342 ( .A(c3468), .B(b[3468]), .Z(n10405) );
XNOR U17343 ( .A(b[3468]), .B(n10406), .Z(c[3468]) );
XNOR U17344 ( .A(a[3468]), .B(c3468), .Z(n10406) );
XOR U17345 ( .A(c3469), .B(n10407), .Z(c3470) );
ANDN U17346 ( .B(n10408), .A(n10409), .Z(n10407) );
XOR U17347 ( .A(c3469), .B(b[3469]), .Z(n10408) );
XNOR U17348 ( .A(b[3469]), .B(n10409), .Z(c[3469]) );
XNOR U17349 ( .A(a[3469]), .B(c3469), .Z(n10409) );
XOR U17350 ( .A(c3470), .B(n10410), .Z(c3471) );
ANDN U17351 ( .B(n10411), .A(n10412), .Z(n10410) );
XOR U17352 ( .A(c3470), .B(b[3470]), .Z(n10411) );
XNOR U17353 ( .A(b[3470]), .B(n10412), .Z(c[3470]) );
XNOR U17354 ( .A(a[3470]), .B(c3470), .Z(n10412) );
XOR U17355 ( .A(c3471), .B(n10413), .Z(c3472) );
ANDN U17356 ( .B(n10414), .A(n10415), .Z(n10413) );
XOR U17357 ( .A(c3471), .B(b[3471]), .Z(n10414) );
XNOR U17358 ( .A(b[3471]), .B(n10415), .Z(c[3471]) );
XNOR U17359 ( .A(a[3471]), .B(c3471), .Z(n10415) );
XOR U17360 ( .A(c3472), .B(n10416), .Z(c3473) );
ANDN U17361 ( .B(n10417), .A(n10418), .Z(n10416) );
XOR U17362 ( .A(c3472), .B(b[3472]), .Z(n10417) );
XNOR U17363 ( .A(b[3472]), .B(n10418), .Z(c[3472]) );
XNOR U17364 ( .A(a[3472]), .B(c3472), .Z(n10418) );
XOR U17365 ( .A(c3473), .B(n10419), .Z(c3474) );
ANDN U17366 ( .B(n10420), .A(n10421), .Z(n10419) );
XOR U17367 ( .A(c3473), .B(b[3473]), .Z(n10420) );
XNOR U17368 ( .A(b[3473]), .B(n10421), .Z(c[3473]) );
XNOR U17369 ( .A(a[3473]), .B(c3473), .Z(n10421) );
XOR U17370 ( .A(c3474), .B(n10422), .Z(c3475) );
ANDN U17371 ( .B(n10423), .A(n10424), .Z(n10422) );
XOR U17372 ( .A(c3474), .B(b[3474]), .Z(n10423) );
XNOR U17373 ( .A(b[3474]), .B(n10424), .Z(c[3474]) );
XNOR U17374 ( .A(a[3474]), .B(c3474), .Z(n10424) );
XOR U17375 ( .A(c3475), .B(n10425), .Z(c3476) );
ANDN U17376 ( .B(n10426), .A(n10427), .Z(n10425) );
XOR U17377 ( .A(c3475), .B(b[3475]), .Z(n10426) );
XNOR U17378 ( .A(b[3475]), .B(n10427), .Z(c[3475]) );
XNOR U17379 ( .A(a[3475]), .B(c3475), .Z(n10427) );
XOR U17380 ( .A(c3476), .B(n10428), .Z(c3477) );
ANDN U17381 ( .B(n10429), .A(n10430), .Z(n10428) );
XOR U17382 ( .A(c3476), .B(b[3476]), .Z(n10429) );
XNOR U17383 ( .A(b[3476]), .B(n10430), .Z(c[3476]) );
XNOR U17384 ( .A(a[3476]), .B(c3476), .Z(n10430) );
XOR U17385 ( .A(c3477), .B(n10431), .Z(c3478) );
ANDN U17386 ( .B(n10432), .A(n10433), .Z(n10431) );
XOR U17387 ( .A(c3477), .B(b[3477]), .Z(n10432) );
XNOR U17388 ( .A(b[3477]), .B(n10433), .Z(c[3477]) );
XNOR U17389 ( .A(a[3477]), .B(c3477), .Z(n10433) );
XOR U17390 ( .A(c3478), .B(n10434), .Z(c3479) );
ANDN U17391 ( .B(n10435), .A(n10436), .Z(n10434) );
XOR U17392 ( .A(c3478), .B(b[3478]), .Z(n10435) );
XNOR U17393 ( .A(b[3478]), .B(n10436), .Z(c[3478]) );
XNOR U17394 ( .A(a[3478]), .B(c3478), .Z(n10436) );
XOR U17395 ( .A(c3479), .B(n10437), .Z(c3480) );
ANDN U17396 ( .B(n10438), .A(n10439), .Z(n10437) );
XOR U17397 ( .A(c3479), .B(b[3479]), .Z(n10438) );
XNOR U17398 ( .A(b[3479]), .B(n10439), .Z(c[3479]) );
XNOR U17399 ( .A(a[3479]), .B(c3479), .Z(n10439) );
XOR U17400 ( .A(c3480), .B(n10440), .Z(c3481) );
ANDN U17401 ( .B(n10441), .A(n10442), .Z(n10440) );
XOR U17402 ( .A(c3480), .B(b[3480]), .Z(n10441) );
XNOR U17403 ( .A(b[3480]), .B(n10442), .Z(c[3480]) );
XNOR U17404 ( .A(a[3480]), .B(c3480), .Z(n10442) );
XOR U17405 ( .A(c3481), .B(n10443), .Z(c3482) );
ANDN U17406 ( .B(n10444), .A(n10445), .Z(n10443) );
XOR U17407 ( .A(c3481), .B(b[3481]), .Z(n10444) );
XNOR U17408 ( .A(b[3481]), .B(n10445), .Z(c[3481]) );
XNOR U17409 ( .A(a[3481]), .B(c3481), .Z(n10445) );
XOR U17410 ( .A(c3482), .B(n10446), .Z(c3483) );
ANDN U17411 ( .B(n10447), .A(n10448), .Z(n10446) );
XOR U17412 ( .A(c3482), .B(b[3482]), .Z(n10447) );
XNOR U17413 ( .A(b[3482]), .B(n10448), .Z(c[3482]) );
XNOR U17414 ( .A(a[3482]), .B(c3482), .Z(n10448) );
XOR U17415 ( .A(c3483), .B(n10449), .Z(c3484) );
ANDN U17416 ( .B(n10450), .A(n10451), .Z(n10449) );
XOR U17417 ( .A(c3483), .B(b[3483]), .Z(n10450) );
XNOR U17418 ( .A(b[3483]), .B(n10451), .Z(c[3483]) );
XNOR U17419 ( .A(a[3483]), .B(c3483), .Z(n10451) );
XOR U17420 ( .A(c3484), .B(n10452), .Z(c3485) );
ANDN U17421 ( .B(n10453), .A(n10454), .Z(n10452) );
XOR U17422 ( .A(c3484), .B(b[3484]), .Z(n10453) );
XNOR U17423 ( .A(b[3484]), .B(n10454), .Z(c[3484]) );
XNOR U17424 ( .A(a[3484]), .B(c3484), .Z(n10454) );
XOR U17425 ( .A(c3485), .B(n10455), .Z(c3486) );
ANDN U17426 ( .B(n10456), .A(n10457), .Z(n10455) );
XOR U17427 ( .A(c3485), .B(b[3485]), .Z(n10456) );
XNOR U17428 ( .A(b[3485]), .B(n10457), .Z(c[3485]) );
XNOR U17429 ( .A(a[3485]), .B(c3485), .Z(n10457) );
XOR U17430 ( .A(c3486), .B(n10458), .Z(c3487) );
ANDN U17431 ( .B(n10459), .A(n10460), .Z(n10458) );
XOR U17432 ( .A(c3486), .B(b[3486]), .Z(n10459) );
XNOR U17433 ( .A(b[3486]), .B(n10460), .Z(c[3486]) );
XNOR U17434 ( .A(a[3486]), .B(c3486), .Z(n10460) );
XOR U17435 ( .A(c3487), .B(n10461), .Z(c3488) );
ANDN U17436 ( .B(n10462), .A(n10463), .Z(n10461) );
XOR U17437 ( .A(c3487), .B(b[3487]), .Z(n10462) );
XNOR U17438 ( .A(b[3487]), .B(n10463), .Z(c[3487]) );
XNOR U17439 ( .A(a[3487]), .B(c3487), .Z(n10463) );
XOR U17440 ( .A(c3488), .B(n10464), .Z(c3489) );
ANDN U17441 ( .B(n10465), .A(n10466), .Z(n10464) );
XOR U17442 ( .A(c3488), .B(b[3488]), .Z(n10465) );
XNOR U17443 ( .A(b[3488]), .B(n10466), .Z(c[3488]) );
XNOR U17444 ( .A(a[3488]), .B(c3488), .Z(n10466) );
XOR U17445 ( .A(c3489), .B(n10467), .Z(c3490) );
ANDN U17446 ( .B(n10468), .A(n10469), .Z(n10467) );
XOR U17447 ( .A(c3489), .B(b[3489]), .Z(n10468) );
XNOR U17448 ( .A(b[3489]), .B(n10469), .Z(c[3489]) );
XNOR U17449 ( .A(a[3489]), .B(c3489), .Z(n10469) );
XOR U17450 ( .A(c3490), .B(n10470), .Z(c3491) );
ANDN U17451 ( .B(n10471), .A(n10472), .Z(n10470) );
XOR U17452 ( .A(c3490), .B(b[3490]), .Z(n10471) );
XNOR U17453 ( .A(b[3490]), .B(n10472), .Z(c[3490]) );
XNOR U17454 ( .A(a[3490]), .B(c3490), .Z(n10472) );
XOR U17455 ( .A(c3491), .B(n10473), .Z(c3492) );
ANDN U17456 ( .B(n10474), .A(n10475), .Z(n10473) );
XOR U17457 ( .A(c3491), .B(b[3491]), .Z(n10474) );
XNOR U17458 ( .A(b[3491]), .B(n10475), .Z(c[3491]) );
XNOR U17459 ( .A(a[3491]), .B(c3491), .Z(n10475) );
XOR U17460 ( .A(c3492), .B(n10476), .Z(c3493) );
ANDN U17461 ( .B(n10477), .A(n10478), .Z(n10476) );
XOR U17462 ( .A(c3492), .B(b[3492]), .Z(n10477) );
XNOR U17463 ( .A(b[3492]), .B(n10478), .Z(c[3492]) );
XNOR U17464 ( .A(a[3492]), .B(c3492), .Z(n10478) );
XOR U17465 ( .A(c3493), .B(n10479), .Z(c3494) );
ANDN U17466 ( .B(n10480), .A(n10481), .Z(n10479) );
XOR U17467 ( .A(c3493), .B(b[3493]), .Z(n10480) );
XNOR U17468 ( .A(b[3493]), .B(n10481), .Z(c[3493]) );
XNOR U17469 ( .A(a[3493]), .B(c3493), .Z(n10481) );
XOR U17470 ( .A(c3494), .B(n10482), .Z(c3495) );
ANDN U17471 ( .B(n10483), .A(n10484), .Z(n10482) );
XOR U17472 ( .A(c3494), .B(b[3494]), .Z(n10483) );
XNOR U17473 ( .A(b[3494]), .B(n10484), .Z(c[3494]) );
XNOR U17474 ( .A(a[3494]), .B(c3494), .Z(n10484) );
XOR U17475 ( .A(c3495), .B(n10485), .Z(c3496) );
ANDN U17476 ( .B(n10486), .A(n10487), .Z(n10485) );
XOR U17477 ( .A(c3495), .B(b[3495]), .Z(n10486) );
XNOR U17478 ( .A(b[3495]), .B(n10487), .Z(c[3495]) );
XNOR U17479 ( .A(a[3495]), .B(c3495), .Z(n10487) );
XOR U17480 ( .A(c3496), .B(n10488), .Z(c3497) );
ANDN U17481 ( .B(n10489), .A(n10490), .Z(n10488) );
XOR U17482 ( .A(c3496), .B(b[3496]), .Z(n10489) );
XNOR U17483 ( .A(b[3496]), .B(n10490), .Z(c[3496]) );
XNOR U17484 ( .A(a[3496]), .B(c3496), .Z(n10490) );
XOR U17485 ( .A(c3497), .B(n10491), .Z(c3498) );
ANDN U17486 ( .B(n10492), .A(n10493), .Z(n10491) );
XOR U17487 ( .A(c3497), .B(b[3497]), .Z(n10492) );
XNOR U17488 ( .A(b[3497]), .B(n10493), .Z(c[3497]) );
XNOR U17489 ( .A(a[3497]), .B(c3497), .Z(n10493) );
XOR U17490 ( .A(c3498), .B(n10494), .Z(c3499) );
ANDN U17491 ( .B(n10495), .A(n10496), .Z(n10494) );
XOR U17492 ( .A(c3498), .B(b[3498]), .Z(n10495) );
XNOR U17493 ( .A(b[3498]), .B(n10496), .Z(c[3498]) );
XNOR U17494 ( .A(a[3498]), .B(c3498), .Z(n10496) );
XOR U17495 ( .A(c3499), .B(n10497), .Z(c3500) );
ANDN U17496 ( .B(n10498), .A(n10499), .Z(n10497) );
XOR U17497 ( .A(c3499), .B(b[3499]), .Z(n10498) );
XNOR U17498 ( .A(b[3499]), .B(n10499), .Z(c[3499]) );
XNOR U17499 ( .A(a[3499]), .B(c3499), .Z(n10499) );
XOR U17500 ( .A(c3500), .B(n10500), .Z(c3501) );
ANDN U17501 ( .B(n10501), .A(n10502), .Z(n10500) );
XOR U17502 ( .A(c3500), .B(b[3500]), .Z(n10501) );
XNOR U17503 ( .A(b[3500]), .B(n10502), .Z(c[3500]) );
XNOR U17504 ( .A(a[3500]), .B(c3500), .Z(n10502) );
XOR U17505 ( .A(c3501), .B(n10503), .Z(c3502) );
ANDN U17506 ( .B(n10504), .A(n10505), .Z(n10503) );
XOR U17507 ( .A(c3501), .B(b[3501]), .Z(n10504) );
XNOR U17508 ( .A(b[3501]), .B(n10505), .Z(c[3501]) );
XNOR U17509 ( .A(a[3501]), .B(c3501), .Z(n10505) );
XOR U17510 ( .A(c3502), .B(n10506), .Z(c3503) );
ANDN U17511 ( .B(n10507), .A(n10508), .Z(n10506) );
XOR U17512 ( .A(c3502), .B(b[3502]), .Z(n10507) );
XNOR U17513 ( .A(b[3502]), .B(n10508), .Z(c[3502]) );
XNOR U17514 ( .A(a[3502]), .B(c3502), .Z(n10508) );
XOR U17515 ( .A(c3503), .B(n10509), .Z(c3504) );
ANDN U17516 ( .B(n10510), .A(n10511), .Z(n10509) );
XOR U17517 ( .A(c3503), .B(b[3503]), .Z(n10510) );
XNOR U17518 ( .A(b[3503]), .B(n10511), .Z(c[3503]) );
XNOR U17519 ( .A(a[3503]), .B(c3503), .Z(n10511) );
XOR U17520 ( .A(c3504), .B(n10512), .Z(c3505) );
ANDN U17521 ( .B(n10513), .A(n10514), .Z(n10512) );
XOR U17522 ( .A(c3504), .B(b[3504]), .Z(n10513) );
XNOR U17523 ( .A(b[3504]), .B(n10514), .Z(c[3504]) );
XNOR U17524 ( .A(a[3504]), .B(c3504), .Z(n10514) );
XOR U17525 ( .A(c3505), .B(n10515), .Z(c3506) );
ANDN U17526 ( .B(n10516), .A(n10517), .Z(n10515) );
XOR U17527 ( .A(c3505), .B(b[3505]), .Z(n10516) );
XNOR U17528 ( .A(b[3505]), .B(n10517), .Z(c[3505]) );
XNOR U17529 ( .A(a[3505]), .B(c3505), .Z(n10517) );
XOR U17530 ( .A(c3506), .B(n10518), .Z(c3507) );
ANDN U17531 ( .B(n10519), .A(n10520), .Z(n10518) );
XOR U17532 ( .A(c3506), .B(b[3506]), .Z(n10519) );
XNOR U17533 ( .A(b[3506]), .B(n10520), .Z(c[3506]) );
XNOR U17534 ( .A(a[3506]), .B(c3506), .Z(n10520) );
XOR U17535 ( .A(c3507), .B(n10521), .Z(c3508) );
ANDN U17536 ( .B(n10522), .A(n10523), .Z(n10521) );
XOR U17537 ( .A(c3507), .B(b[3507]), .Z(n10522) );
XNOR U17538 ( .A(b[3507]), .B(n10523), .Z(c[3507]) );
XNOR U17539 ( .A(a[3507]), .B(c3507), .Z(n10523) );
XOR U17540 ( .A(c3508), .B(n10524), .Z(c3509) );
ANDN U17541 ( .B(n10525), .A(n10526), .Z(n10524) );
XOR U17542 ( .A(c3508), .B(b[3508]), .Z(n10525) );
XNOR U17543 ( .A(b[3508]), .B(n10526), .Z(c[3508]) );
XNOR U17544 ( .A(a[3508]), .B(c3508), .Z(n10526) );
XOR U17545 ( .A(c3509), .B(n10527), .Z(c3510) );
ANDN U17546 ( .B(n10528), .A(n10529), .Z(n10527) );
XOR U17547 ( .A(c3509), .B(b[3509]), .Z(n10528) );
XNOR U17548 ( .A(b[3509]), .B(n10529), .Z(c[3509]) );
XNOR U17549 ( .A(a[3509]), .B(c3509), .Z(n10529) );
XOR U17550 ( .A(c3510), .B(n10530), .Z(c3511) );
ANDN U17551 ( .B(n10531), .A(n10532), .Z(n10530) );
XOR U17552 ( .A(c3510), .B(b[3510]), .Z(n10531) );
XNOR U17553 ( .A(b[3510]), .B(n10532), .Z(c[3510]) );
XNOR U17554 ( .A(a[3510]), .B(c3510), .Z(n10532) );
XOR U17555 ( .A(c3511), .B(n10533), .Z(c3512) );
ANDN U17556 ( .B(n10534), .A(n10535), .Z(n10533) );
XOR U17557 ( .A(c3511), .B(b[3511]), .Z(n10534) );
XNOR U17558 ( .A(b[3511]), .B(n10535), .Z(c[3511]) );
XNOR U17559 ( .A(a[3511]), .B(c3511), .Z(n10535) );
XOR U17560 ( .A(c3512), .B(n10536), .Z(c3513) );
ANDN U17561 ( .B(n10537), .A(n10538), .Z(n10536) );
XOR U17562 ( .A(c3512), .B(b[3512]), .Z(n10537) );
XNOR U17563 ( .A(b[3512]), .B(n10538), .Z(c[3512]) );
XNOR U17564 ( .A(a[3512]), .B(c3512), .Z(n10538) );
XOR U17565 ( .A(c3513), .B(n10539), .Z(c3514) );
ANDN U17566 ( .B(n10540), .A(n10541), .Z(n10539) );
XOR U17567 ( .A(c3513), .B(b[3513]), .Z(n10540) );
XNOR U17568 ( .A(b[3513]), .B(n10541), .Z(c[3513]) );
XNOR U17569 ( .A(a[3513]), .B(c3513), .Z(n10541) );
XOR U17570 ( .A(c3514), .B(n10542), .Z(c3515) );
ANDN U17571 ( .B(n10543), .A(n10544), .Z(n10542) );
XOR U17572 ( .A(c3514), .B(b[3514]), .Z(n10543) );
XNOR U17573 ( .A(b[3514]), .B(n10544), .Z(c[3514]) );
XNOR U17574 ( .A(a[3514]), .B(c3514), .Z(n10544) );
XOR U17575 ( .A(c3515), .B(n10545), .Z(c3516) );
ANDN U17576 ( .B(n10546), .A(n10547), .Z(n10545) );
XOR U17577 ( .A(c3515), .B(b[3515]), .Z(n10546) );
XNOR U17578 ( .A(b[3515]), .B(n10547), .Z(c[3515]) );
XNOR U17579 ( .A(a[3515]), .B(c3515), .Z(n10547) );
XOR U17580 ( .A(c3516), .B(n10548), .Z(c3517) );
ANDN U17581 ( .B(n10549), .A(n10550), .Z(n10548) );
XOR U17582 ( .A(c3516), .B(b[3516]), .Z(n10549) );
XNOR U17583 ( .A(b[3516]), .B(n10550), .Z(c[3516]) );
XNOR U17584 ( .A(a[3516]), .B(c3516), .Z(n10550) );
XOR U17585 ( .A(c3517), .B(n10551), .Z(c3518) );
ANDN U17586 ( .B(n10552), .A(n10553), .Z(n10551) );
XOR U17587 ( .A(c3517), .B(b[3517]), .Z(n10552) );
XNOR U17588 ( .A(b[3517]), .B(n10553), .Z(c[3517]) );
XNOR U17589 ( .A(a[3517]), .B(c3517), .Z(n10553) );
XOR U17590 ( .A(c3518), .B(n10554), .Z(c3519) );
ANDN U17591 ( .B(n10555), .A(n10556), .Z(n10554) );
XOR U17592 ( .A(c3518), .B(b[3518]), .Z(n10555) );
XNOR U17593 ( .A(b[3518]), .B(n10556), .Z(c[3518]) );
XNOR U17594 ( .A(a[3518]), .B(c3518), .Z(n10556) );
XOR U17595 ( .A(c3519), .B(n10557), .Z(c3520) );
ANDN U17596 ( .B(n10558), .A(n10559), .Z(n10557) );
XOR U17597 ( .A(c3519), .B(b[3519]), .Z(n10558) );
XNOR U17598 ( .A(b[3519]), .B(n10559), .Z(c[3519]) );
XNOR U17599 ( .A(a[3519]), .B(c3519), .Z(n10559) );
XOR U17600 ( .A(c3520), .B(n10560), .Z(c3521) );
ANDN U17601 ( .B(n10561), .A(n10562), .Z(n10560) );
XOR U17602 ( .A(c3520), .B(b[3520]), .Z(n10561) );
XNOR U17603 ( .A(b[3520]), .B(n10562), .Z(c[3520]) );
XNOR U17604 ( .A(a[3520]), .B(c3520), .Z(n10562) );
XOR U17605 ( .A(c3521), .B(n10563), .Z(c3522) );
ANDN U17606 ( .B(n10564), .A(n10565), .Z(n10563) );
XOR U17607 ( .A(c3521), .B(b[3521]), .Z(n10564) );
XNOR U17608 ( .A(b[3521]), .B(n10565), .Z(c[3521]) );
XNOR U17609 ( .A(a[3521]), .B(c3521), .Z(n10565) );
XOR U17610 ( .A(c3522), .B(n10566), .Z(c3523) );
ANDN U17611 ( .B(n10567), .A(n10568), .Z(n10566) );
XOR U17612 ( .A(c3522), .B(b[3522]), .Z(n10567) );
XNOR U17613 ( .A(b[3522]), .B(n10568), .Z(c[3522]) );
XNOR U17614 ( .A(a[3522]), .B(c3522), .Z(n10568) );
XOR U17615 ( .A(c3523), .B(n10569), .Z(c3524) );
ANDN U17616 ( .B(n10570), .A(n10571), .Z(n10569) );
XOR U17617 ( .A(c3523), .B(b[3523]), .Z(n10570) );
XNOR U17618 ( .A(b[3523]), .B(n10571), .Z(c[3523]) );
XNOR U17619 ( .A(a[3523]), .B(c3523), .Z(n10571) );
XOR U17620 ( .A(c3524), .B(n10572), .Z(c3525) );
ANDN U17621 ( .B(n10573), .A(n10574), .Z(n10572) );
XOR U17622 ( .A(c3524), .B(b[3524]), .Z(n10573) );
XNOR U17623 ( .A(b[3524]), .B(n10574), .Z(c[3524]) );
XNOR U17624 ( .A(a[3524]), .B(c3524), .Z(n10574) );
XOR U17625 ( .A(c3525), .B(n10575), .Z(c3526) );
ANDN U17626 ( .B(n10576), .A(n10577), .Z(n10575) );
XOR U17627 ( .A(c3525), .B(b[3525]), .Z(n10576) );
XNOR U17628 ( .A(b[3525]), .B(n10577), .Z(c[3525]) );
XNOR U17629 ( .A(a[3525]), .B(c3525), .Z(n10577) );
XOR U17630 ( .A(c3526), .B(n10578), .Z(c3527) );
ANDN U17631 ( .B(n10579), .A(n10580), .Z(n10578) );
XOR U17632 ( .A(c3526), .B(b[3526]), .Z(n10579) );
XNOR U17633 ( .A(b[3526]), .B(n10580), .Z(c[3526]) );
XNOR U17634 ( .A(a[3526]), .B(c3526), .Z(n10580) );
XOR U17635 ( .A(c3527), .B(n10581), .Z(c3528) );
ANDN U17636 ( .B(n10582), .A(n10583), .Z(n10581) );
XOR U17637 ( .A(c3527), .B(b[3527]), .Z(n10582) );
XNOR U17638 ( .A(b[3527]), .B(n10583), .Z(c[3527]) );
XNOR U17639 ( .A(a[3527]), .B(c3527), .Z(n10583) );
XOR U17640 ( .A(c3528), .B(n10584), .Z(c3529) );
ANDN U17641 ( .B(n10585), .A(n10586), .Z(n10584) );
XOR U17642 ( .A(c3528), .B(b[3528]), .Z(n10585) );
XNOR U17643 ( .A(b[3528]), .B(n10586), .Z(c[3528]) );
XNOR U17644 ( .A(a[3528]), .B(c3528), .Z(n10586) );
XOR U17645 ( .A(c3529), .B(n10587), .Z(c3530) );
ANDN U17646 ( .B(n10588), .A(n10589), .Z(n10587) );
XOR U17647 ( .A(c3529), .B(b[3529]), .Z(n10588) );
XNOR U17648 ( .A(b[3529]), .B(n10589), .Z(c[3529]) );
XNOR U17649 ( .A(a[3529]), .B(c3529), .Z(n10589) );
XOR U17650 ( .A(c3530), .B(n10590), .Z(c3531) );
ANDN U17651 ( .B(n10591), .A(n10592), .Z(n10590) );
XOR U17652 ( .A(c3530), .B(b[3530]), .Z(n10591) );
XNOR U17653 ( .A(b[3530]), .B(n10592), .Z(c[3530]) );
XNOR U17654 ( .A(a[3530]), .B(c3530), .Z(n10592) );
XOR U17655 ( .A(c3531), .B(n10593), .Z(c3532) );
ANDN U17656 ( .B(n10594), .A(n10595), .Z(n10593) );
XOR U17657 ( .A(c3531), .B(b[3531]), .Z(n10594) );
XNOR U17658 ( .A(b[3531]), .B(n10595), .Z(c[3531]) );
XNOR U17659 ( .A(a[3531]), .B(c3531), .Z(n10595) );
XOR U17660 ( .A(c3532), .B(n10596), .Z(c3533) );
ANDN U17661 ( .B(n10597), .A(n10598), .Z(n10596) );
XOR U17662 ( .A(c3532), .B(b[3532]), .Z(n10597) );
XNOR U17663 ( .A(b[3532]), .B(n10598), .Z(c[3532]) );
XNOR U17664 ( .A(a[3532]), .B(c3532), .Z(n10598) );
XOR U17665 ( .A(c3533), .B(n10599), .Z(c3534) );
ANDN U17666 ( .B(n10600), .A(n10601), .Z(n10599) );
XOR U17667 ( .A(c3533), .B(b[3533]), .Z(n10600) );
XNOR U17668 ( .A(b[3533]), .B(n10601), .Z(c[3533]) );
XNOR U17669 ( .A(a[3533]), .B(c3533), .Z(n10601) );
XOR U17670 ( .A(c3534), .B(n10602), .Z(c3535) );
ANDN U17671 ( .B(n10603), .A(n10604), .Z(n10602) );
XOR U17672 ( .A(c3534), .B(b[3534]), .Z(n10603) );
XNOR U17673 ( .A(b[3534]), .B(n10604), .Z(c[3534]) );
XNOR U17674 ( .A(a[3534]), .B(c3534), .Z(n10604) );
XOR U17675 ( .A(c3535), .B(n10605), .Z(c3536) );
ANDN U17676 ( .B(n10606), .A(n10607), .Z(n10605) );
XOR U17677 ( .A(c3535), .B(b[3535]), .Z(n10606) );
XNOR U17678 ( .A(b[3535]), .B(n10607), .Z(c[3535]) );
XNOR U17679 ( .A(a[3535]), .B(c3535), .Z(n10607) );
XOR U17680 ( .A(c3536), .B(n10608), .Z(c3537) );
ANDN U17681 ( .B(n10609), .A(n10610), .Z(n10608) );
XOR U17682 ( .A(c3536), .B(b[3536]), .Z(n10609) );
XNOR U17683 ( .A(b[3536]), .B(n10610), .Z(c[3536]) );
XNOR U17684 ( .A(a[3536]), .B(c3536), .Z(n10610) );
XOR U17685 ( .A(c3537), .B(n10611), .Z(c3538) );
ANDN U17686 ( .B(n10612), .A(n10613), .Z(n10611) );
XOR U17687 ( .A(c3537), .B(b[3537]), .Z(n10612) );
XNOR U17688 ( .A(b[3537]), .B(n10613), .Z(c[3537]) );
XNOR U17689 ( .A(a[3537]), .B(c3537), .Z(n10613) );
XOR U17690 ( .A(c3538), .B(n10614), .Z(c3539) );
ANDN U17691 ( .B(n10615), .A(n10616), .Z(n10614) );
XOR U17692 ( .A(c3538), .B(b[3538]), .Z(n10615) );
XNOR U17693 ( .A(b[3538]), .B(n10616), .Z(c[3538]) );
XNOR U17694 ( .A(a[3538]), .B(c3538), .Z(n10616) );
XOR U17695 ( .A(c3539), .B(n10617), .Z(c3540) );
ANDN U17696 ( .B(n10618), .A(n10619), .Z(n10617) );
XOR U17697 ( .A(c3539), .B(b[3539]), .Z(n10618) );
XNOR U17698 ( .A(b[3539]), .B(n10619), .Z(c[3539]) );
XNOR U17699 ( .A(a[3539]), .B(c3539), .Z(n10619) );
XOR U17700 ( .A(c3540), .B(n10620), .Z(c3541) );
ANDN U17701 ( .B(n10621), .A(n10622), .Z(n10620) );
XOR U17702 ( .A(c3540), .B(b[3540]), .Z(n10621) );
XNOR U17703 ( .A(b[3540]), .B(n10622), .Z(c[3540]) );
XNOR U17704 ( .A(a[3540]), .B(c3540), .Z(n10622) );
XOR U17705 ( .A(c3541), .B(n10623), .Z(c3542) );
ANDN U17706 ( .B(n10624), .A(n10625), .Z(n10623) );
XOR U17707 ( .A(c3541), .B(b[3541]), .Z(n10624) );
XNOR U17708 ( .A(b[3541]), .B(n10625), .Z(c[3541]) );
XNOR U17709 ( .A(a[3541]), .B(c3541), .Z(n10625) );
XOR U17710 ( .A(c3542), .B(n10626), .Z(c3543) );
ANDN U17711 ( .B(n10627), .A(n10628), .Z(n10626) );
XOR U17712 ( .A(c3542), .B(b[3542]), .Z(n10627) );
XNOR U17713 ( .A(b[3542]), .B(n10628), .Z(c[3542]) );
XNOR U17714 ( .A(a[3542]), .B(c3542), .Z(n10628) );
XOR U17715 ( .A(c3543), .B(n10629), .Z(c3544) );
ANDN U17716 ( .B(n10630), .A(n10631), .Z(n10629) );
XOR U17717 ( .A(c3543), .B(b[3543]), .Z(n10630) );
XNOR U17718 ( .A(b[3543]), .B(n10631), .Z(c[3543]) );
XNOR U17719 ( .A(a[3543]), .B(c3543), .Z(n10631) );
XOR U17720 ( .A(c3544), .B(n10632), .Z(c3545) );
ANDN U17721 ( .B(n10633), .A(n10634), .Z(n10632) );
XOR U17722 ( .A(c3544), .B(b[3544]), .Z(n10633) );
XNOR U17723 ( .A(b[3544]), .B(n10634), .Z(c[3544]) );
XNOR U17724 ( .A(a[3544]), .B(c3544), .Z(n10634) );
XOR U17725 ( .A(c3545), .B(n10635), .Z(c3546) );
ANDN U17726 ( .B(n10636), .A(n10637), .Z(n10635) );
XOR U17727 ( .A(c3545), .B(b[3545]), .Z(n10636) );
XNOR U17728 ( .A(b[3545]), .B(n10637), .Z(c[3545]) );
XNOR U17729 ( .A(a[3545]), .B(c3545), .Z(n10637) );
XOR U17730 ( .A(c3546), .B(n10638), .Z(c3547) );
ANDN U17731 ( .B(n10639), .A(n10640), .Z(n10638) );
XOR U17732 ( .A(c3546), .B(b[3546]), .Z(n10639) );
XNOR U17733 ( .A(b[3546]), .B(n10640), .Z(c[3546]) );
XNOR U17734 ( .A(a[3546]), .B(c3546), .Z(n10640) );
XOR U17735 ( .A(c3547), .B(n10641), .Z(c3548) );
ANDN U17736 ( .B(n10642), .A(n10643), .Z(n10641) );
XOR U17737 ( .A(c3547), .B(b[3547]), .Z(n10642) );
XNOR U17738 ( .A(b[3547]), .B(n10643), .Z(c[3547]) );
XNOR U17739 ( .A(a[3547]), .B(c3547), .Z(n10643) );
XOR U17740 ( .A(c3548), .B(n10644), .Z(c3549) );
ANDN U17741 ( .B(n10645), .A(n10646), .Z(n10644) );
XOR U17742 ( .A(c3548), .B(b[3548]), .Z(n10645) );
XNOR U17743 ( .A(b[3548]), .B(n10646), .Z(c[3548]) );
XNOR U17744 ( .A(a[3548]), .B(c3548), .Z(n10646) );
XOR U17745 ( .A(c3549), .B(n10647), .Z(c3550) );
ANDN U17746 ( .B(n10648), .A(n10649), .Z(n10647) );
XOR U17747 ( .A(c3549), .B(b[3549]), .Z(n10648) );
XNOR U17748 ( .A(b[3549]), .B(n10649), .Z(c[3549]) );
XNOR U17749 ( .A(a[3549]), .B(c3549), .Z(n10649) );
XOR U17750 ( .A(c3550), .B(n10650), .Z(c3551) );
ANDN U17751 ( .B(n10651), .A(n10652), .Z(n10650) );
XOR U17752 ( .A(c3550), .B(b[3550]), .Z(n10651) );
XNOR U17753 ( .A(b[3550]), .B(n10652), .Z(c[3550]) );
XNOR U17754 ( .A(a[3550]), .B(c3550), .Z(n10652) );
XOR U17755 ( .A(c3551), .B(n10653), .Z(c3552) );
ANDN U17756 ( .B(n10654), .A(n10655), .Z(n10653) );
XOR U17757 ( .A(c3551), .B(b[3551]), .Z(n10654) );
XNOR U17758 ( .A(b[3551]), .B(n10655), .Z(c[3551]) );
XNOR U17759 ( .A(a[3551]), .B(c3551), .Z(n10655) );
XOR U17760 ( .A(c3552), .B(n10656), .Z(c3553) );
ANDN U17761 ( .B(n10657), .A(n10658), .Z(n10656) );
XOR U17762 ( .A(c3552), .B(b[3552]), .Z(n10657) );
XNOR U17763 ( .A(b[3552]), .B(n10658), .Z(c[3552]) );
XNOR U17764 ( .A(a[3552]), .B(c3552), .Z(n10658) );
XOR U17765 ( .A(c3553), .B(n10659), .Z(c3554) );
ANDN U17766 ( .B(n10660), .A(n10661), .Z(n10659) );
XOR U17767 ( .A(c3553), .B(b[3553]), .Z(n10660) );
XNOR U17768 ( .A(b[3553]), .B(n10661), .Z(c[3553]) );
XNOR U17769 ( .A(a[3553]), .B(c3553), .Z(n10661) );
XOR U17770 ( .A(c3554), .B(n10662), .Z(c3555) );
ANDN U17771 ( .B(n10663), .A(n10664), .Z(n10662) );
XOR U17772 ( .A(c3554), .B(b[3554]), .Z(n10663) );
XNOR U17773 ( .A(b[3554]), .B(n10664), .Z(c[3554]) );
XNOR U17774 ( .A(a[3554]), .B(c3554), .Z(n10664) );
XOR U17775 ( .A(c3555), .B(n10665), .Z(c3556) );
ANDN U17776 ( .B(n10666), .A(n10667), .Z(n10665) );
XOR U17777 ( .A(c3555), .B(b[3555]), .Z(n10666) );
XNOR U17778 ( .A(b[3555]), .B(n10667), .Z(c[3555]) );
XNOR U17779 ( .A(a[3555]), .B(c3555), .Z(n10667) );
XOR U17780 ( .A(c3556), .B(n10668), .Z(c3557) );
ANDN U17781 ( .B(n10669), .A(n10670), .Z(n10668) );
XOR U17782 ( .A(c3556), .B(b[3556]), .Z(n10669) );
XNOR U17783 ( .A(b[3556]), .B(n10670), .Z(c[3556]) );
XNOR U17784 ( .A(a[3556]), .B(c3556), .Z(n10670) );
XOR U17785 ( .A(c3557), .B(n10671), .Z(c3558) );
ANDN U17786 ( .B(n10672), .A(n10673), .Z(n10671) );
XOR U17787 ( .A(c3557), .B(b[3557]), .Z(n10672) );
XNOR U17788 ( .A(b[3557]), .B(n10673), .Z(c[3557]) );
XNOR U17789 ( .A(a[3557]), .B(c3557), .Z(n10673) );
XOR U17790 ( .A(c3558), .B(n10674), .Z(c3559) );
ANDN U17791 ( .B(n10675), .A(n10676), .Z(n10674) );
XOR U17792 ( .A(c3558), .B(b[3558]), .Z(n10675) );
XNOR U17793 ( .A(b[3558]), .B(n10676), .Z(c[3558]) );
XNOR U17794 ( .A(a[3558]), .B(c3558), .Z(n10676) );
XOR U17795 ( .A(c3559), .B(n10677), .Z(c3560) );
ANDN U17796 ( .B(n10678), .A(n10679), .Z(n10677) );
XOR U17797 ( .A(c3559), .B(b[3559]), .Z(n10678) );
XNOR U17798 ( .A(b[3559]), .B(n10679), .Z(c[3559]) );
XNOR U17799 ( .A(a[3559]), .B(c3559), .Z(n10679) );
XOR U17800 ( .A(c3560), .B(n10680), .Z(c3561) );
ANDN U17801 ( .B(n10681), .A(n10682), .Z(n10680) );
XOR U17802 ( .A(c3560), .B(b[3560]), .Z(n10681) );
XNOR U17803 ( .A(b[3560]), .B(n10682), .Z(c[3560]) );
XNOR U17804 ( .A(a[3560]), .B(c3560), .Z(n10682) );
XOR U17805 ( .A(c3561), .B(n10683), .Z(c3562) );
ANDN U17806 ( .B(n10684), .A(n10685), .Z(n10683) );
XOR U17807 ( .A(c3561), .B(b[3561]), .Z(n10684) );
XNOR U17808 ( .A(b[3561]), .B(n10685), .Z(c[3561]) );
XNOR U17809 ( .A(a[3561]), .B(c3561), .Z(n10685) );
XOR U17810 ( .A(c3562), .B(n10686), .Z(c3563) );
ANDN U17811 ( .B(n10687), .A(n10688), .Z(n10686) );
XOR U17812 ( .A(c3562), .B(b[3562]), .Z(n10687) );
XNOR U17813 ( .A(b[3562]), .B(n10688), .Z(c[3562]) );
XNOR U17814 ( .A(a[3562]), .B(c3562), .Z(n10688) );
XOR U17815 ( .A(c3563), .B(n10689), .Z(c3564) );
ANDN U17816 ( .B(n10690), .A(n10691), .Z(n10689) );
XOR U17817 ( .A(c3563), .B(b[3563]), .Z(n10690) );
XNOR U17818 ( .A(b[3563]), .B(n10691), .Z(c[3563]) );
XNOR U17819 ( .A(a[3563]), .B(c3563), .Z(n10691) );
XOR U17820 ( .A(c3564), .B(n10692), .Z(c3565) );
ANDN U17821 ( .B(n10693), .A(n10694), .Z(n10692) );
XOR U17822 ( .A(c3564), .B(b[3564]), .Z(n10693) );
XNOR U17823 ( .A(b[3564]), .B(n10694), .Z(c[3564]) );
XNOR U17824 ( .A(a[3564]), .B(c3564), .Z(n10694) );
XOR U17825 ( .A(c3565), .B(n10695), .Z(c3566) );
ANDN U17826 ( .B(n10696), .A(n10697), .Z(n10695) );
XOR U17827 ( .A(c3565), .B(b[3565]), .Z(n10696) );
XNOR U17828 ( .A(b[3565]), .B(n10697), .Z(c[3565]) );
XNOR U17829 ( .A(a[3565]), .B(c3565), .Z(n10697) );
XOR U17830 ( .A(c3566), .B(n10698), .Z(c3567) );
ANDN U17831 ( .B(n10699), .A(n10700), .Z(n10698) );
XOR U17832 ( .A(c3566), .B(b[3566]), .Z(n10699) );
XNOR U17833 ( .A(b[3566]), .B(n10700), .Z(c[3566]) );
XNOR U17834 ( .A(a[3566]), .B(c3566), .Z(n10700) );
XOR U17835 ( .A(c3567), .B(n10701), .Z(c3568) );
ANDN U17836 ( .B(n10702), .A(n10703), .Z(n10701) );
XOR U17837 ( .A(c3567), .B(b[3567]), .Z(n10702) );
XNOR U17838 ( .A(b[3567]), .B(n10703), .Z(c[3567]) );
XNOR U17839 ( .A(a[3567]), .B(c3567), .Z(n10703) );
XOR U17840 ( .A(c3568), .B(n10704), .Z(c3569) );
ANDN U17841 ( .B(n10705), .A(n10706), .Z(n10704) );
XOR U17842 ( .A(c3568), .B(b[3568]), .Z(n10705) );
XNOR U17843 ( .A(b[3568]), .B(n10706), .Z(c[3568]) );
XNOR U17844 ( .A(a[3568]), .B(c3568), .Z(n10706) );
XOR U17845 ( .A(c3569), .B(n10707), .Z(c3570) );
ANDN U17846 ( .B(n10708), .A(n10709), .Z(n10707) );
XOR U17847 ( .A(c3569), .B(b[3569]), .Z(n10708) );
XNOR U17848 ( .A(b[3569]), .B(n10709), .Z(c[3569]) );
XNOR U17849 ( .A(a[3569]), .B(c3569), .Z(n10709) );
XOR U17850 ( .A(c3570), .B(n10710), .Z(c3571) );
ANDN U17851 ( .B(n10711), .A(n10712), .Z(n10710) );
XOR U17852 ( .A(c3570), .B(b[3570]), .Z(n10711) );
XNOR U17853 ( .A(b[3570]), .B(n10712), .Z(c[3570]) );
XNOR U17854 ( .A(a[3570]), .B(c3570), .Z(n10712) );
XOR U17855 ( .A(c3571), .B(n10713), .Z(c3572) );
ANDN U17856 ( .B(n10714), .A(n10715), .Z(n10713) );
XOR U17857 ( .A(c3571), .B(b[3571]), .Z(n10714) );
XNOR U17858 ( .A(b[3571]), .B(n10715), .Z(c[3571]) );
XNOR U17859 ( .A(a[3571]), .B(c3571), .Z(n10715) );
XOR U17860 ( .A(c3572), .B(n10716), .Z(c3573) );
ANDN U17861 ( .B(n10717), .A(n10718), .Z(n10716) );
XOR U17862 ( .A(c3572), .B(b[3572]), .Z(n10717) );
XNOR U17863 ( .A(b[3572]), .B(n10718), .Z(c[3572]) );
XNOR U17864 ( .A(a[3572]), .B(c3572), .Z(n10718) );
XOR U17865 ( .A(c3573), .B(n10719), .Z(c3574) );
ANDN U17866 ( .B(n10720), .A(n10721), .Z(n10719) );
XOR U17867 ( .A(c3573), .B(b[3573]), .Z(n10720) );
XNOR U17868 ( .A(b[3573]), .B(n10721), .Z(c[3573]) );
XNOR U17869 ( .A(a[3573]), .B(c3573), .Z(n10721) );
XOR U17870 ( .A(c3574), .B(n10722), .Z(c3575) );
ANDN U17871 ( .B(n10723), .A(n10724), .Z(n10722) );
XOR U17872 ( .A(c3574), .B(b[3574]), .Z(n10723) );
XNOR U17873 ( .A(b[3574]), .B(n10724), .Z(c[3574]) );
XNOR U17874 ( .A(a[3574]), .B(c3574), .Z(n10724) );
XOR U17875 ( .A(c3575), .B(n10725), .Z(c3576) );
ANDN U17876 ( .B(n10726), .A(n10727), .Z(n10725) );
XOR U17877 ( .A(c3575), .B(b[3575]), .Z(n10726) );
XNOR U17878 ( .A(b[3575]), .B(n10727), .Z(c[3575]) );
XNOR U17879 ( .A(a[3575]), .B(c3575), .Z(n10727) );
XOR U17880 ( .A(c3576), .B(n10728), .Z(c3577) );
ANDN U17881 ( .B(n10729), .A(n10730), .Z(n10728) );
XOR U17882 ( .A(c3576), .B(b[3576]), .Z(n10729) );
XNOR U17883 ( .A(b[3576]), .B(n10730), .Z(c[3576]) );
XNOR U17884 ( .A(a[3576]), .B(c3576), .Z(n10730) );
XOR U17885 ( .A(c3577), .B(n10731), .Z(c3578) );
ANDN U17886 ( .B(n10732), .A(n10733), .Z(n10731) );
XOR U17887 ( .A(c3577), .B(b[3577]), .Z(n10732) );
XNOR U17888 ( .A(b[3577]), .B(n10733), .Z(c[3577]) );
XNOR U17889 ( .A(a[3577]), .B(c3577), .Z(n10733) );
XOR U17890 ( .A(c3578), .B(n10734), .Z(c3579) );
ANDN U17891 ( .B(n10735), .A(n10736), .Z(n10734) );
XOR U17892 ( .A(c3578), .B(b[3578]), .Z(n10735) );
XNOR U17893 ( .A(b[3578]), .B(n10736), .Z(c[3578]) );
XNOR U17894 ( .A(a[3578]), .B(c3578), .Z(n10736) );
XOR U17895 ( .A(c3579), .B(n10737), .Z(c3580) );
ANDN U17896 ( .B(n10738), .A(n10739), .Z(n10737) );
XOR U17897 ( .A(c3579), .B(b[3579]), .Z(n10738) );
XNOR U17898 ( .A(b[3579]), .B(n10739), .Z(c[3579]) );
XNOR U17899 ( .A(a[3579]), .B(c3579), .Z(n10739) );
XOR U17900 ( .A(c3580), .B(n10740), .Z(c3581) );
ANDN U17901 ( .B(n10741), .A(n10742), .Z(n10740) );
XOR U17902 ( .A(c3580), .B(b[3580]), .Z(n10741) );
XNOR U17903 ( .A(b[3580]), .B(n10742), .Z(c[3580]) );
XNOR U17904 ( .A(a[3580]), .B(c3580), .Z(n10742) );
XOR U17905 ( .A(c3581), .B(n10743), .Z(c3582) );
ANDN U17906 ( .B(n10744), .A(n10745), .Z(n10743) );
XOR U17907 ( .A(c3581), .B(b[3581]), .Z(n10744) );
XNOR U17908 ( .A(b[3581]), .B(n10745), .Z(c[3581]) );
XNOR U17909 ( .A(a[3581]), .B(c3581), .Z(n10745) );
XOR U17910 ( .A(c3582), .B(n10746), .Z(c3583) );
ANDN U17911 ( .B(n10747), .A(n10748), .Z(n10746) );
XOR U17912 ( .A(c3582), .B(b[3582]), .Z(n10747) );
XNOR U17913 ( .A(b[3582]), .B(n10748), .Z(c[3582]) );
XNOR U17914 ( .A(a[3582]), .B(c3582), .Z(n10748) );
XOR U17915 ( .A(c3583), .B(n10749), .Z(c3584) );
ANDN U17916 ( .B(n10750), .A(n10751), .Z(n10749) );
XOR U17917 ( .A(c3583), .B(b[3583]), .Z(n10750) );
XNOR U17918 ( .A(b[3583]), .B(n10751), .Z(c[3583]) );
XNOR U17919 ( .A(a[3583]), .B(c3583), .Z(n10751) );
XOR U17920 ( .A(c3584), .B(n10752), .Z(c3585) );
ANDN U17921 ( .B(n10753), .A(n10754), .Z(n10752) );
XOR U17922 ( .A(c3584), .B(b[3584]), .Z(n10753) );
XNOR U17923 ( .A(b[3584]), .B(n10754), .Z(c[3584]) );
XNOR U17924 ( .A(a[3584]), .B(c3584), .Z(n10754) );
XOR U17925 ( .A(c3585), .B(n10755), .Z(c3586) );
ANDN U17926 ( .B(n10756), .A(n10757), .Z(n10755) );
XOR U17927 ( .A(c3585), .B(b[3585]), .Z(n10756) );
XNOR U17928 ( .A(b[3585]), .B(n10757), .Z(c[3585]) );
XNOR U17929 ( .A(a[3585]), .B(c3585), .Z(n10757) );
XOR U17930 ( .A(c3586), .B(n10758), .Z(c3587) );
ANDN U17931 ( .B(n10759), .A(n10760), .Z(n10758) );
XOR U17932 ( .A(c3586), .B(b[3586]), .Z(n10759) );
XNOR U17933 ( .A(b[3586]), .B(n10760), .Z(c[3586]) );
XNOR U17934 ( .A(a[3586]), .B(c3586), .Z(n10760) );
XOR U17935 ( .A(c3587), .B(n10761), .Z(c3588) );
ANDN U17936 ( .B(n10762), .A(n10763), .Z(n10761) );
XOR U17937 ( .A(c3587), .B(b[3587]), .Z(n10762) );
XNOR U17938 ( .A(b[3587]), .B(n10763), .Z(c[3587]) );
XNOR U17939 ( .A(a[3587]), .B(c3587), .Z(n10763) );
XOR U17940 ( .A(c3588), .B(n10764), .Z(c3589) );
ANDN U17941 ( .B(n10765), .A(n10766), .Z(n10764) );
XOR U17942 ( .A(c3588), .B(b[3588]), .Z(n10765) );
XNOR U17943 ( .A(b[3588]), .B(n10766), .Z(c[3588]) );
XNOR U17944 ( .A(a[3588]), .B(c3588), .Z(n10766) );
XOR U17945 ( .A(c3589), .B(n10767), .Z(c3590) );
ANDN U17946 ( .B(n10768), .A(n10769), .Z(n10767) );
XOR U17947 ( .A(c3589), .B(b[3589]), .Z(n10768) );
XNOR U17948 ( .A(b[3589]), .B(n10769), .Z(c[3589]) );
XNOR U17949 ( .A(a[3589]), .B(c3589), .Z(n10769) );
XOR U17950 ( .A(c3590), .B(n10770), .Z(c3591) );
ANDN U17951 ( .B(n10771), .A(n10772), .Z(n10770) );
XOR U17952 ( .A(c3590), .B(b[3590]), .Z(n10771) );
XNOR U17953 ( .A(b[3590]), .B(n10772), .Z(c[3590]) );
XNOR U17954 ( .A(a[3590]), .B(c3590), .Z(n10772) );
XOR U17955 ( .A(c3591), .B(n10773), .Z(c3592) );
ANDN U17956 ( .B(n10774), .A(n10775), .Z(n10773) );
XOR U17957 ( .A(c3591), .B(b[3591]), .Z(n10774) );
XNOR U17958 ( .A(b[3591]), .B(n10775), .Z(c[3591]) );
XNOR U17959 ( .A(a[3591]), .B(c3591), .Z(n10775) );
XOR U17960 ( .A(c3592), .B(n10776), .Z(c3593) );
ANDN U17961 ( .B(n10777), .A(n10778), .Z(n10776) );
XOR U17962 ( .A(c3592), .B(b[3592]), .Z(n10777) );
XNOR U17963 ( .A(b[3592]), .B(n10778), .Z(c[3592]) );
XNOR U17964 ( .A(a[3592]), .B(c3592), .Z(n10778) );
XOR U17965 ( .A(c3593), .B(n10779), .Z(c3594) );
ANDN U17966 ( .B(n10780), .A(n10781), .Z(n10779) );
XOR U17967 ( .A(c3593), .B(b[3593]), .Z(n10780) );
XNOR U17968 ( .A(b[3593]), .B(n10781), .Z(c[3593]) );
XNOR U17969 ( .A(a[3593]), .B(c3593), .Z(n10781) );
XOR U17970 ( .A(c3594), .B(n10782), .Z(c3595) );
ANDN U17971 ( .B(n10783), .A(n10784), .Z(n10782) );
XOR U17972 ( .A(c3594), .B(b[3594]), .Z(n10783) );
XNOR U17973 ( .A(b[3594]), .B(n10784), .Z(c[3594]) );
XNOR U17974 ( .A(a[3594]), .B(c3594), .Z(n10784) );
XOR U17975 ( .A(c3595), .B(n10785), .Z(c3596) );
ANDN U17976 ( .B(n10786), .A(n10787), .Z(n10785) );
XOR U17977 ( .A(c3595), .B(b[3595]), .Z(n10786) );
XNOR U17978 ( .A(b[3595]), .B(n10787), .Z(c[3595]) );
XNOR U17979 ( .A(a[3595]), .B(c3595), .Z(n10787) );
XOR U17980 ( .A(c3596), .B(n10788), .Z(c3597) );
ANDN U17981 ( .B(n10789), .A(n10790), .Z(n10788) );
XOR U17982 ( .A(c3596), .B(b[3596]), .Z(n10789) );
XNOR U17983 ( .A(b[3596]), .B(n10790), .Z(c[3596]) );
XNOR U17984 ( .A(a[3596]), .B(c3596), .Z(n10790) );
XOR U17985 ( .A(c3597), .B(n10791), .Z(c3598) );
ANDN U17986 ( .B(n10792), .A(n10793), .Z(n10791) );
XOR U17987 ( .A(c3597), .B(b[3597]), .Z(n10792) );
XNOR U17988 ( .A(b[3597]), .B(n10793), .Z(c[3597]) );
XNOR U17989 ( .A(a[3597]), .B(c3597), .Z(n10793) );
XOR U17990 ( .A(c3598), .B(n10794), .Z(c3599) );
ANDN U17991 ( .B(n10795), .A(n10796), .Z(n10794) );
XOR U17992 ( .A(c3598), .B(b[3598]), .Z(n10795) );
XNOR U17993 ( .A(b[3598]), .B(n10796), .Z(c[3598]) );
XNOR U17994 ( .A(a[3598]), .B(c3598), .Z(n10796) );
XOR U17995 ( .A(c3599), .B(n10797), .Z(c3600) );
ANDN U17996 ( .B(n10798), .A(n10799), .Z(n10797) );
XOR U17997 ( .A(c3599), .B(b[3599]), .Z(n10798) );
XNOR U17998 ( .A(b[3599]), .B(n10799), .Z(c[3599]) );
XNOR U17999 ( .A(a[3599]), .B(c3599), .Z(n10799) );
XOR U18000 ( .A(c3600), .B(n10800), .Z(c3601) );
ANDN U18001 ( .B(n10801), .A(n10802), .Z(n10800) );
XOR U18002 ( .A(c3600), .B(b[3600]), .Z(n10801) );
XNOR U18003 ( .A(b[3600]), .B(n10802), .Z(c[3600]) );
XNOR U18004 ( .A(a[3600]), .B(c3600), .Z(n10802) );
XOR U18005 ( .A(c3601), .B(n10803), .Z(c3602) );
ANDN U18006 ( .B(n10804), .A(n10805), .Z(n10803) );
XOR U18007 ( .A(c3601), .B(b[3601]), .Z(n10804) );
XNOR U18008 ( .A(b[3601]), .B(n10805), .Z(c[3601]) );
XNOR U18009 ( .A(a[3601]), .B(c3601), .Z(n10805) );
XOR U18010 ( .A(c3602), .B(n10806), .Z(c3603) );
ANDN U18011 ( .B(n10807), .A(n10808), .Z(n10806) );
XOR U18012 ( .A(c3602), .B(b[3602]), .Z(n10807) );
XNOR U18013 ( .A(b[3602]), .B(n10808), .Z(c[3602]) );
XNOR U18014 ( .A(a[3602]), .B(c3602), .Z(n10808) );
XOR U18015 ( .A(c3603), .B(n10809), .Z(c3604) );
ANDN U18016 ( .B(n10810), .A(n10811), .Z(n10809) );
XOR U18017 ( .A(c3603), .B(b[3603]), .Z(n10810) );
XNOR U18018 ( .A(b[3603]), .B(n10811), .Z(c[3603]) );
XNOR U18019 ( .A(a[3603]), .B(c3603), .Z(n10811) );
XOR U18020 ( .A(c3604), .B(n10812), .Z(c3605) );
ANDN U18021 ( .B(n10813), .A(n10814), .Z(n10812) );
XOR U18022 ( .A(c3604), .B(b[3604]), .Z(n10813) );
XNOR U18023 ( .A(b[3604]), .B(n10814), .Z(c[3604]) );
XNOR U18024 ( .A(a[3604]), .B(c3604), .Z(n10814) );
XOR U18025 ( .A(c3605), .B(n10815), .Z(c3606) );
ANDN U18026 ( .B(n10816), .A(n10817), .Z(n10815) );
XOR U18027 ( .A(c3605), .B(b[3605]), .Z(n10816) );
XNOR U18028 ( .A(b[3605]), .B(n10817), .Z(c[3605]) );
XNOR U18029 ( .A(a[3605]), .B(c3605), .Z(n10817) );
XOR U18030 ( .A(c3606), .B(n10818), .Z(c3607) );
ANDN U18031 ( .B(n10819), .A(n10820), .Z(n10818) );
XOR U18032 ( .A(c3606), .B(b[3606]), .Z(n10819) );
XNOR U18033 ( .A(b[3606]), .B(n10820), .Z(c[3606]) );
XNOR U18034 ( .A(a[3606]), .B(c3606), .Z(n10820) );
XOR U18035 ( .A(c3607), .B(n10821), .Z(c3608) );
ANDN U18036 ( .B(n10822), .A(n10823), .Z(n10821) );
XOR U18037 ( .A(c3607), .B(b[3607]), .Z(n10822) );
XNOR U18038 ( .A(b[3607]), .B(n10823), .Z(c[3607]) );
XNOR U18039 ( .A(a[3607]), .B(c3607), .Z(n10823) );
XOR U18040 ( .A(c3608), .B(n10824), .Z(c3609) );
ANDN U18041 ( .B(n10825), .A(n10826), .Z(n10824) );
XOR U18042 ( .A(c3608), .B(b[3608]), .Z(n10825) );
XNOR U18043 ( .A(b[3608]), .B(n10826), .Z(c[3608]) );
XNOR U18044 ( .A(a[3608]), .B(c3608), .Z(n10826) );
XOR U18045 ( .A(c3609), .B(n10827), .Z(c3610) );
ANDN U18046 ( .B(n10828), .A(n10829), .Z(n10827) );
XOR U18047 ( .A(c3609), .B(b[3609]), .Z(n10828) );
XNOR U18048 ( .A(b[3609]), .B(n10829), .Z(c[3609]) );
XNOR U18049 ( .A(a[3609]), .B(c3609), .Z(n10829) );
XOR U18050 ( .A(c3610), .B(n10830), .Z(c3611) );
ANDN U18051 ( .B(n10831), .A(n10832), .Z(n10830) );
XOR U18052 ( .A(c3610), .B(b[3610]), .Z(n10831) );
XNOR U18053 ( .A(b[3610]), .B(n10832), .Z(c[3610]) );
XNOR U18054 ( .A(a[3610]), .B(c3610), .Z(n10832) );
XOR U18055 ( .A(c3611), .B(n10833), .Z(c3612) );
ANDN U18056 ( .B(n10834), .A(n10835), .Z(n10833) );
XOR U18057 ( .A(c3611), .B(b[3611]), .Z(n10834) );
XNOR U18058 ( .A(b[3611]), .B(n10835), .Z(c[3611]) );
XNOR U18059 ( .A(a[3611]), .B(c3611), .Z(n10835) );
XOR U18060 ( .A(c3612), .B(n10836), .Z(c3613) );
ANDN U18061 ( .B(n10837), .A(n10838), .Z(n10836) );
XOR U18062 ( .A(c3612), .B(b[3612]), .Z(n10837) );
XNOR U18063 ( .A(b[3612]), .B(n10838), .Z(c[3612]) );
XNOR U18064 ( .A(a[3612]), .B(c3612), .Z(n10838) );
XOR U18065 ( .A(c3613), .B(n10839), .Z(c3614) );
ANDN U18066 ( .B(n10840), .A(n10841), .Z(n10839) );
XOR U18067 ( .A(c3613), .B(b[3613]), .Z(n10840) );
XNOR U18068 ( .A(b[3613]), .B(n10841), .Z(c[3613]) );
XNOR U18069 ( .A(a[3613]), .B(c3613), .Z(n10841) );
XOR U18070 ( .A(c3614), .B(n10842), .Z(c3615) );
ANDN U18071 ( .B(n10843), .A(n10844), .Z(n10842) );
XOR U18072 ( .A(c3614), .B(b[3614]), .Z(n10843) );
XNOR U18073 ( .A(b[3614]), .B(n10844), .Z(c[3614]) );
XNOR U18074 ( .A(a[3614]), .B(c3614), .Z(n10844) );
XOR U18075 ( .A(c3615), .B(n10845), .Z(c3616) );
ANDN U18076 ( .B(n10846), .A(n10847), .Z(n10845) );
XOR U18077 ( .A(c3615), .B(b[3615]), .Z(n10846) );
XNOR U18078 ( .A(b[3615]), .B(n10847), .Z(c[3615]) );
XNOR U18079 ( .A(a[3615]), .B(c3615), .Z(n10847) );
XOR U18080 ( .A(c3616), .B(n10848), .Z(c3617) );
ANDN U18081 ( .B(n10849), .A(n10850), .Z(n10848) );
XOR U18082 ( .A(c3616), .B(b[3616]), .Z(n10849) );
XNOR U18083 ( .A(b[3616]), .B(n10850), .Z(c[3616]) );
XNOR U18084 ( .A(a[3616]), .B(c3616), .Z(n10850) );
XOR U18085 ( .A(c3617), .B(n10851), .Z(c3618) );
ANDN U18086 ( .B(n10852), .A(n10853), .Z(n10851) );
XOR U18087 ( .A(c3617), .B(b[3617]), .Z(n10852) );
XNOR U18088 ( .A(b[3617]), .B(n10853), .Z(c[3617]) );
XNOR U18089 ( .A(a[3617]), .B(c3617), .Z(n10853) );
XOR U18090 ( .A(c3618), .B(n10854), .Z(c3619) );
ANDN U18091 ( .B(n10855), .A(n10856), .Z(n10854) );
XOR U18092 ( .A(c3618), .B(b[3618]), .Z(n10855) );
XNOR U18093 ( .A(b[3618]), .B(n10856), .Z(c[3618]) );
XNOR U18094 ( .A(a[3618]), .B(c3618), .Z(n10856) );
XOR U18095 ( .A(c3619), .B(n10857), .Z(c3620) );
ANDN U18096 ( .B(n10858), .A(n10859), .Z(n10857) );
XOR U18097 ( .A(c3619), .B(b[3619]), .Z(n10858) );
XNOR U18098 ( .A(b[3619]), .B(n10859), .Z(c[3619]) );
XNOR U18099 ( .A(a[3619]), .B(c3619), .Z(n10859) );
XOR U18100 ( .A(c3620), .B(n10860), .Z(c3621) );
ANDN U18101 ( .B(n10861), .A(n10862), .Z(n10860) );
XOR U18102 ( .A(c3620), .B(b[3620]), .Z(n10861) );
XNOR U18103 ( .A(b[3620]), .B(n10862), .Z(c[3620]) );
XNOR U18104 ( .A(a[3620]), .B(c3620), .Z(n10862) );
XOR U18105 ( .A(c3621), .B(n10863), .Z(c3622) );
ANDN U18106 ( .B(n10864), .A(n10865), .Z(n10863) );
XOR U18107 ( .A(c3621), .B(b[3621]), .Z(n10864) );
XNOR U18108 ( .A(b[3621]), .B(n10865), .Z(c[3621]) );
XNOR U18109 ( .A(a[3621]), .B(c3621), .Z(n10865) );
XOR U18110 ( .A(c3622), .B(n10866), .Z(c3623) );
ANDN U18111 ( .B(n10867), .A(n10868), .Z(n10866) );
XOR U18112 ( .A(c3622), .B(b[3622]), .Z(n10867) );
XNOR U18113 ( .A(b[3622]), .B(n10868), .Z(c[3622]) );
XNOR U18114 ( .A(a[3622]), .B(c3622), .Z(n10868) );
XOR U18115 ( .A(c3623), .B(n10869), .Z(c3624) );
ANDN U18116 ( .B(n10870), .A(n10871), .Z(n10869) );
XOR U18117 ( .A(c3623), .B(b[3623]), .Z(n10870) );
XNOR U18118 ( .A(b[3623]), .B(n10871), .Z(c[3623]) );
XNOR U18119 ( .A(a[3623]), .B(c3623), .Z(n10871) );
XOR U18120 ( .A(c3624), .B(n10872), .Z(c3625) );
ANDN U18121 ( .B(n10873), .A(n10874), .Z(n10872) );
XOR U18122 ( .A(c3624), .B(b[3624]), .Z(n10873) );
XNOR U18123 ( .A(b[3624]), .B(n10874), .Z(c[3624]) );
XNOR U18124 ( .A(a[3624]), .B(c3624), .Z(n10874) );
XOR U18125 ( .A(c3625), .B(n10875), .Z(c3626) );
ANDN U18126 ( .B(n10876), .A(n10877), .Z(n10875) );
XOR U18127 ( .A(c3625), .B(b[3625]), .Z(n10876) );
XNOR U18128 ( .A(b[3625]), .B(n10877), .Z(c[3625]) );
XNOR U18129 ( .A(a[3625]), .B(c3625), .Z(n10877) );
XOR U18130 ( .A(c3626), .B(n10878), .Z(c3627) );
ANDN U18131 ( .B(n10879), .A(n10880), .Z(n10878) );
XOR U18132 ( .A(c3626), .B(b[3626]), .Z(n10879) );
XNOR U18133 ( .A(b[3626]), .B(n10880), .Z(c[3626]) );
XNOR U18134 ( .A(a[3626]), .B(c3626), .Z(n10880) );
XOR U18135 ( .A(c3627), .B(n10881), .Z(c3628) );
ANDN U18136 ( .B(n10882), .A(n10883), .Z(n10881) );
XOR U18137 ( .A(c3627), .B(b[3627]), .Z(n10882) );
XNOR U18138 ( .A(b[3627]), .B(n10883), .Z(c[3627]) );
XNOR U18139 ( .A(a[3627]), .B(c3627), .Z(n10883) );
XOR U18140 ( .A(c3628), .B(n10884), .Z(c3629) );
ANDN U18141 ( .B(n10885), .A(n10886), .Z(n10884) );
XOR U18142 ( .A(c3628), .B(b[3628]), .Z(n10885) );
XNOR U18143 ( .A(b[3628]), .B(n10886), .Z(c[3628]) );
XNOR U18144 ( .A(a[3628]), .B(c3628), .Z(n10886) );
XOR U18145 ( .A(c3629), .B(n10887), .Z(c3630) );
ANDN U18146 ( .B(n10888), .A(n10889), .Z(n10887) );
XOR U18147 ( .A(c3629), .B(b[3629]), .Z(n10888) );
XNOR U18148 ( .A(b[3629]), .B(n10889), .Z(c[3629]) );
XNOR U18149 ( .A(a[3629]), .B(c3629), .Z(n10889) );
XOR U18150 ( .A(c3630), .B(n10890), .Z(c3631) );
ANDN U18151 ( .B(n10891), .A(n10892), .Z(n10890) );
XOR U18152 ( .A(c3630), .B(b[3630]), .Z(n10891) );
XNOR U18153 ( .A(b[3630]), .B(n10892), .Z(c[3630]) );
XNOR U18154 ( .A(a[3630]), .B(c3630), .Z(n10892) );
XOR U18155 ( .A(c3631), .B(n10893), .Z(c3632) );
ANDN U18156 ( .B(n10894), .A(n10895), .Z(n10893) );
XOR U18157 ( .A(c3631), .B(b[3631]), .Z(n10894) );
XNOR U18158 ( .A(b[3631]), .B(n10895), .Z(c[3631]) );
XNOR U18159 ( .A(a[3631]), .B(c3631), .Z(n10895) );
XOR U18160 ( .A(c3632), .B(n10896), .Z(c3633) );
ANDN U18161 ( .B(n10897), .A(n10898), .Z(n10896) );
XOR U18162 ( .A(c3632), .B(b[3632]), .Z(n10897) );
XNOR U18163 ( .A(b[3632]), .B(n10898), .Z(c[3632]) );
XNOR U18164 ( .A(a[3632]), .B(c3632), .Z(n10898) );
XOR U18165 ( .A(c3633), .B(n10899), .Z(c3634) );
ANDN U18166 ( .B(n10900), .A(n10901), .Z(n10899) );
XOR U18167 ( .A(c3633), .B(b[3633]), .Z(n10900) );
XNOR U18168 ( .A(b[3633]), .B(n10901), .Z(c[3633]) );
XNOR U18169 ( .A(a[3633]), .B(c3633), .Z(n10901) );
XOR U18170 ( .A(c3634), .B(n10902), .Z(c3635) );
ANDN U18171 ( .B(n10903), .A(n10904), .Z(n10902) );
XOR U18172 ( .A(c3634), .B(b[3634]), .Z(n10903) );
XNOR U18173 ( .A(b[3634]), .B(n10904), .Z(c[3634]) );
XNOR U18174 ( .A(a[3634]), .B(c3634), .Z(n10904) );
XOR U18175 ( .A(c3635), .B(n10905), .Z(c3636) );
ANDN U18176 ( .B(n10906), .A(n10907), .Z(n10905) );
XOR U18177 ( .A(c3635), .B(b[3635]), .Z(n10906) );
XNOR U18178 ( .A(b[3635]), .B(n10907), .Z(c[3635]) );
XNOR U18179 ( .A(a[3635]), .B(c3635), .Z(n10907) );
XOR U18180 ( .A(c3636), .B(n10908), .Z(c3637) );
ANDN U18181 ( .B(n10909), .A(n10910), .Z(n10908) );
XOR U18182 ( .A(c3636), .B(b[3636]), .Z(n10909) );
XNOR U18183 ( .A(b[3636]), .B(n10910), .Z(c[3636]) );
XNOR U18184 ( .A(a[3636]), .B(c3636), .Z(n10910) );
XOR U18185 ( .A(c3637), .B(n10911), .Z(c3638) );
ANDN U18186 ( .B(n10912), .A(n10913), .Z(n10911) );
XOR U18187 ( .A(c3637), .B(b[3637]), .Z(n10912) );
XNOR U18188 ( .A(b[3637]), .B(n10913), .Z(c[3637]) );
XNOR U18189 ( .A(a[3637]), .B(c3637), .Z(n10913) );
XOR U18190 ( .A(c3638), .B(n10914), .Z(c3639) );
ANDN U18191 ( .B(n10915), .A(n10916), .Z(n10914) );
XOR U18192 ( .A(c3638), .B(b[3638]), .Z(n10915) );
XNOR U18193 ( .A(b[3638]), .B(n10916), .Z(c[3638]) );
XNOR U18194 ( .A(a[3638]), .B(c3638), .Z(n10916) );
XOR U18195 ( .A(c3639), .B(n10917), .Z(c3640) );
ANDN U18196 ( .B(n10918), .A(n10919), .Z(n10917) );
XOR U18197 ( .A(c3639), .B(b[3639]), .Z(n10918) );
XNOR U18198 ( .A(b[3639]), .B(n10919), .Z(c[3639]) );
XNOR U18199 ( .A(a[3639]), .B(c3639), .Z(n10919) );
XOR U18200 ( .A(c3640), .B(n10920), .Z(c3641) );
ANDN U18201 ( .B(n10921), .A(n10922), .Z(n10920) );
XOR U18202 ( .A(c3640), .B(b[3640]), .Z(n10921) );
XNOR U18203 ( .A(b[3640]), .B(n10922), .Z(c[3640]) );
XNOR U18204 ( .A(a[3640]), .B(c3640), .Z(n10922) );
XOR U18205 ( .A(c3641), .B(n10923), .Z(c3642) );
ANDN U18206 ( .B(n10924), .A(n10925), .Z(n10923) );
XOR U18207 ( .A(c3641), .B(b[3641]), .Z(n10924) );
XNOR U18208 ( .A(b[3641]), .B(n10925), .Z(c[3641]) );
XNOR U18209 ( .A(a[3641]), .B(c3641), .Z(n10925) );
XOR U18210 ( .A(c3642), .B(n10926), .Z(c3643) );
ANDN U18211 ( .B(n10927), .A(n10928), .Z(n10926) );
XOR U18212 ( .A(c3642), .B(b[3642]), .Z(n10927) );
XNOR U18213 ( .A(b[3642]), .B(n10928), .Z(c[3642]) );
XNOR U18214 ( .A(a[3642]), .B(c3642), .Z(n10928) );
XOR U18215 ( .A(c3643), .B(n10929), .Z(c3644) );
ANDN U18216 ( .B(n10930), .A(n10931), .Z(n10929) );
XOR U18217 ( .A(c3643), .B(b[3643]), .Z(n10930) );
XNOR U18218 ( .A(b[3643]), .B(n10931), .Z(c[3643]) );
XNOR U18219 ( .A(a[3643]), .B(c3643), .Z(n10931) );
XOR U18220 ( .A(c3644), .B(n10932), .Z(c3645) );
ANDN U18221 ( .B(n10933), .A(n10934), .Z(n10932) );
XOR U18222 ( .A(c3644), .B(b[3644]), .Z(n10933) );
XNOR U18223 ( .A(b[3644]), .B(n10934), .Z(c[3644]) );
XNOR U18224 ( .A(a[3644]), .B(c3644), .Z(n10934) );
XOR U18225 ( .A(c3645), .B(n10935), .Z(c3646) );
ANDN U18226 ( .B(n10936), .A(n10937), .Z(n10935) );
XOR U18227 ( .A(c3645), .B(b[3645]), .Z(n10936) );
XNOR U18228 ( .A(b[3645]), .B(n10937), .Z(c[3645]) );
XNOR U18229 ( .A(a[3645]), .B(c3645), .Z(n10937) );
XOR U18230 ( .A(c3646), .B(n10938), .Z(c3647) );
ANDN U18231 ( .B(n10939), .A(n10940), .Z(n10938) );
XOR U18232 ( .A(c3646), .B(b[3646]), .Z(n10939) );
XNOR U18233 ( .A(b[3646]), .B(n10940), .Z(c[3646]) );
XNOR U18234 ( .A(a[3646]), .B(c3646), .Z(n10940) );
XOR U18235 ( .A(c3647), .B(n10941), .Z(c3648) );
ANDN U18236 ( .B(n10942), .A(n10943), .Z(n10941) );
XOR U18237 ( .A(c3647), .B(b[3647]), .Z(n10942) );
XNOR U18238 ( .A(b[3647]), .B(n10943), .Z(c[3647]) );
XNOR U18239 ( .A(a[3647]), .B(c3647), .Z(n10943) );
XOR U18240 ( .A(c3648), .B(n10944), .Z(c3649) );
ANDN U18241 ( .B(n10945), .A(n10946), .Z(n10944) );
XOR U18242 ( .A(c3648), .B(b[3648]), .Z(n10945) );
XNOR U18243 ( .A(b[3648]), .B(n10946), .Z(c[3648]) );
XNOR U18244 ( .A(a[3648]), .B(c3648), .Z(n10946) );
XOR U18245 ( .A(c3649), .B(n10947), .Z(c3650) );
ANDN U18246 ( .B(n10948), .A(n10949), .Z(n10947) );
XOR U18247 ( .A(c3649), .B(b[3649]), .Z(n10948) );
XNOR U18248 ( .A(b[3649]), .B(n10949), .Z(c[3649]) );
XNOR U18249 ( .A(a[3649]), .B(c3649), .Z(n10949) );
XOR U18250 ( .A(c3650), .B(n10950), .Z(c3651) );
ANDN U18251 ( .B(n10951), .A(n10952), .Z(n10950) );
XOR U18252 ( .A(c3650), .B(b[3650]), .Z(n10951) );
XNOR U18253 ( .A(b[3650]), .B(n10952), .Z(c[3650]) );
XNOR U18254 ( .A(a[3650]), .B(c3650), .Z(n10952) );
XOR U18255 ( .A(c3651), .B(n10953), .Z(c3652) );
ANDN U18256 ( .B(n10954), .A(n10955), .Z(n10953) );
XOR U18257 ( .A(c3651), .B(b[3651]), .Z(n10954) );
XNOR U18258 ( .A(b[3651]), .B(n10955), .Z(c[3651]) );
XNOR U18259 ( .A(a[3651]), .B(c3651), .Z(n10955) );
XOR U18260 ( .A(c3652), .B(n10956), .Z(c3653) );
ANDN U18261 ( .B(n10957), .A(n10958), .Z(n10956) );
XOR U18262 ( .A(c3652), .B(b[3652]), .Z(n10957) );
XNOR U18263 ( .A(b[3652]), .B(n10958), .Z(c[3652]) );
XNOR U18264 ( .A(a[3652]), .B(c3652), .Z(n10958) );
XOR U18265 ( .A(c3653), .B(n10959), .Z(c3654) );
ANDN U18266 ( .B(n10960), .A(n10961), .Z(n10959) );
XOR U18267 ( .A(c3653), .B(b[3653]), .Z(n10960) );
XNOR U18268 ( .A(b[3653]), .B(n10961), .Z(c[3653]) );
XNOR U18269 ( .A(a[3653]), .B(c3653), .Z(n10961) );
XOR U18270 ( .A(c3654), .B(n10962), .Z(c3655) );
ANDN U18271 ( .B(n10963), .A(n10964), .Z(n10962) );
XOR U18272 ( .A(c3654), .B(b[3654]), .Z(n10963) );
XNOR U18273 ( .A(b[3654]), .B(n10964), .Z(c[3654]) );
XNOR U18274 ( .A(a[3654]), .B(c3654), .Z(n10964) );
XOR U18275 ( .A(c3655), .B(n10965), .Z(c3656) );
ANDN U18276 ( .B(n10966), .A(n10967), .Z(n10965) );
XOR U18277 ( .A(c3655), .B(b[3655]), .Z(n10966) );
XNOR U18278 ( .A(b[3655]), .B(n10967), .Z(c[3655]) );
XNOR U18279 ( .A(a[3655]), .B(c3655), .Z(n10967) );
XOR U18280 ( .A(c3656), .B(n10968), .Z(c3657) );
ANDN U18281 ( .B(n10969), .A(n10970), .Z(n10968) );
XOR U18282 ( .A(c3656), .B(b[3656]), .Z(n10969) );
XNOR U18283 ( .A(b[3656]), .B(n10970), .Z(c[3656]) );
XNOR U18284 ( .A(a[3656]), .B(c3656), .Z(n10970) );
XOR U18285 ( .A(c3657), .B(n10971), .Z(c3658) );
ANDN U18286 ( .B(n10972), .A(n10973), .Z(n10971) );
XOR U18287 ( .A(c3657), .B(b[3657]), .Z(n10972) );
XNOR U18288 ( .A(b[3657]), .B(n10973), .Z(c[3657]) );
XNOR U18289 ( .A(a[3657]), .B(c3657), .Z(n10973) );
XOR U18290 ( .A(c3658), .B(n10974), .Z(c3659) );
ANDN U18291 ( .B(n10975), .A(n10976), .Z(n10974) );
XOR U18292 ( .A(c3658), .B(b[3658]), .Z(n10975) );
XNOR U18293 ( .A(b[3658]), .B(n10976), .Z(c[3658]) );
XNOR U18294 ( .A(a[3658]), .B(c3658), .Z(n10976) );
XOR U18295 ( .A(c3659), .B(n10977), .Z(c3660) );
ANDN U18296 ( .B(n10978), .A(n10979), .Z(n10977) );
XOR U18297 ( .A(c3659), .B(b[3659]), .Z(n10978) );
XNOR U18298 ( .A(b[3659]), .B(n10979), .Z(c[3659]) );
XNOR U18299 ( .A(a[3659]), .B(c3659), .Z(n10979) );
XOR U18300 ( .A(c3660), .B(n10980), .Z(c3661) );
ANDN U18301 ( .B(n10981), .A(n10982), .Z(n10980) );
XOR U18302 ( .A(c3660), .B(b[3660]), .Z(n10981) );
XNOR U18303 ( .A(b[3660]), .B(n10982), .Z(c[3660]) );
XNOR U18304 ( .A(a[3660]), .B(c3660), .Z(n10982) );
XOR U18305 ( .A(c3661), .B(n10983), .Z(c3662) );
ANDN U18306 ( .B(n10984), .A(n10985), .Z(n10983) );
XOR U18307 ( .A(c3661), .B(b[3661]), .Z(n10984) );
XNOR U18308 ( .A(b[3661]), .B(n10985), .Z(c[3661]) );
XNOR U18309 ( .A(a[3661]), .B(c3661), .Z(n10985) );
XOR U18310 ( .A(c3662), .B(n10986), .Z(c3663) );
ANDN U18311 ( .B(n10987), .A(n10988), .Z(n10986) );
XOR U18312 ( .A(c3662), .B(b[3662]), .Z(n10987) );
XNOR U18313 ( .A(b[3662]), .B(n10988), .Z(c[3662]) );
XNOR U18314 ( .A(a[3662]), .B(c3662), .Z(n10988) );
XOR U18315 ( .A(c3663), .B(n10989), .Z(c3664) );
ANDN U18316 ( .B(n10990), .A(n10991), .Z(n10989) );
XOR U18317 ( .A(c3663), .B(b[3663]), .Z(n10990) );
XNOR U18318 ( .A(b[3663]), .B(n10991), .Z(c[3663]) );
XNOR U18319 ( .A(a[3663]), .B(c3663), .Z(n10991) );
XOR U18320 ( .A(c3664), .B(n10992), .Z(c3665) );
ANDN U18321 ( .B(n10993), .A(n10994), .Z(n10992) );
XOR U18322 ( .A(c3664), .B(b[3664]), .Z(n10993) );
XNOR U18323 ( .A(b[3664]), .B(n10994), .Z(c[3664]) );
XNOR U18324 ( .A(a[3664]), .B(c3664), .Z(n10994) );
XOR U18325 ( .A(c3665), .B(n10995), .Z(c3666) );
ANDN U18326 ( .B(n10996), .A(n10997), .Z(n10995) );
XOR U18327 ( .A(c3665), .B(b[3665]), .Z(n10996) );
XNOR U18328 ( .A(b[3665]), .B(n10997), .Z(c[3665]) );
XNOR U18329 ( .A(a[3665]), .B(c3665), .Z(n10997) );
XOR U18330 ( .A(c3666), .B(n10998), .Z(c3667) );
ANDN U18331 ( .B(n10999), .A(n11000), .Z(n10998) );
XOR U18332 ( .A(c3666), .B(b[3666]), .Z(n10999) );
XNOR U18333 ( .A(b[3666]), .B(n11000), .Z(c[3666]) );
XNOR U18334 ( .A(a[3666]), .B(c3666), .Z(n11000) );
XOR U18335 ( .A(c3667), .B(n11001), .Z(c3668) );
ANDN U18336 ( .B(n11002), .A(n11003), .Z(n11001) );
XOR U18337 ( .A(c3667), .B(b[3667]), .Z(n11002) );
XNOR U18338 ( .A(b[3667]), .B(n11003), .Z(c[3667]) );
XNOR U18339 ( .A(a[3667]), .B(c3667), .Z(n11003) );
XOR U18340 ( .A(c3668), .B(n11004), .Z(c3669) );
ANDN U18341 ( .B(n11005), .A(n11006), .Z(n11004) );
XOR U18342 ( .A(c3668), .B(b[3668]), .Z(n11005) );
XNOR U18343 ( .A(b[3668]), .B(n11006), .Z(c[3668]) );
XNOR U18344 ( .A(a[3668]), .B(c3668), .Z(n11006) );
XOR U18345 ( .A(c3669), .B(n11007), .Z(c3670) );
ANDN U18346 ( .B(n11008), .A(n11009), .Z(n11007) );
XOR U18347 ( .A(c3669), .B(b[3669]), .Z(n11008) );
XNOR U18348 ( .A(b[3669]), .B(n11009), .Z(c[3669]) );
XNOR U18349 ( .A(a[3669]), .B(c3669), .Z(n11009) );
XOR U18350 ( .A(c3670), .B(n11010), .Z(c3671) );
ANDN U18351 ( .B(n11011), .A(n11012), .Z(n11010) );
XOR U18352 ( .A(c3670), .B(b[3670]), .Z(n11011) );
XNOR U18353 ( .A(b[3670]), .B(n11012), .Z(c[3670]) );
XNOR U18354 ( .A(a[3670]), .B(c3670), .Z(n11012) );
XOR U18355 ( .A(c3671), .B(n11013), .Z(c3672) );
ANDN U18356 ( .B(n11014), .A(n11015), .Z(n11013) );
XOR U18357 ( .A(c3671), .B(b[3671]), .Z(n11014) );
XNOR U18358 ( .A(b[3671]), .B(n11015), .Z(c[3671]) );
XNOR U18359 ( .A(a[3671]), .B(c3671), .Z(n11015) );
XOR U18360 ( .A(c3672), .B(n11016), .Z(c3673) );
ANDN U18361 ( .B(n11017), .A(n11018), .Z(n11016) );
XOR U18362 ( .A(c3672), .B(b[3672]), .Z(n11017) );
XNOR U18363 ( .A(b[3672]), .B(n11018), .Z(c[3672]) );
XNOR U18364 ( .A(a[3672]), .B(c3672), .Z(n11018) );
XOR U18365 ( .A(c3673), .B(n11019), .Z(c3674) );
ANDN U18366 ( .B(n11020), .A(n11021), .Z(n11019) );
XOR U18367 ( .A(c3673), .B(b[3673]), .Z(n11020) );
XNOR U18368 ( .A(b[3673]), .B(n11021), .Z(c[3673]) );
XNOR U18369 ( .A(a[3673]), .B(c3673), .Z(n11021) );
XOR U18370 ( .A(c3674), .B(n11022), .Z(c3675) );
ANDN U18371 ( .B(n11023), .A(n11024), .Z(n11022) );
XOR U18372 ( .A(c3674), .B(b[3674]), .Z(n11023) );
XNOR U18373 ( .A(b[3674]), .B(n11024), .Z(c[3674]) );
XNOR U18374 ( .A(a[3674]), .B(c3674), .Z(n11024) );
XOR U18375 ( .A(c3675), .B(n11025), .Z(c3676) );
ANDN U18376 ( .B(n11026), .A(n11027), .Z(n11025) );
XOR U18377 ( .A(c3675), .B(b[3675]), .Z(n11026) );
XNOR U18378 ( .A(b[3675]), .B(n11027), .Z(c[3675]) );
XNOR U18379 ( .A(a[3675]), .B(c3675), .Z(n11027) );
XOR U18380 ( .A(c3676), .B(n11028), .Z(c3677) );
ANDN U18381 ( .B(n11029), .A(n11030), .Z(n11028) );
XOR U18382 ( .A(c3676), .B(b[3676]), .Z(n11029) );
XNOR U18383 ( .A(b[3676]), .B(n11030), .Z(c[3676]) );
XNOR U18384 ( .A(a[3676]), .B(c3676), .Z(n11030) );
XOR U18385 ( .A(c3677), .B(n11031), .Z(c3678) );
ANDN U18386 ( .B(n11032), .A(n11033), .Z(n11031) );
XOR U18387 ( .A(c3677), .B(b[3677]), .Z(n11032) );
XNOR U18388 ( .A(b[3677]), .B(n11033), .Z(c[3677]) );
XNOR U18389 ( .A(a[3677]), .B(c3677), .Z(n11033) );
XOR U18390 ( .A(c3678), .B(n11034), .Z(c3679) );
ANDN U18391 ( .B(n11035), .A(n11036), .Z(n11034) );
XOR U18392 ( .A(c3678), .B(b[3678]), .Z(n11035) );
XNOR U18393 ( .A(b[3678]), .B(n11036), .Z(c[3678]) );
XNOR U18394 ( .A(a[3678]), .B(c3678), .Z(n11036) );
XOR U18395 ( .A(c3679), .B(n11037), .Z(c3680) );
ANDN U18396 ( .B(n11038), .A(n11039), .Z(n11037) );
XOR U18397 ( .A(c3679), .B(b[3679]), .Z(n11038) );
XNOR U18398 ( .A(b[3679]), .B(n11039), .Z(c[3679]) );
XNOR U18399 ( .A(a[3679]), .B(c3679), .Z(n11039) );
XOR U18400 ( .A(c3680), .B(n11040), .Z(c3681) );
ANDN U18401 ( .B(n11041), .A(n11042), .Z(n11040) );
XOR U18402 ( .A(c3680), .B(b[3680]), .Z(n11041) );
XNOR U18403 ( .A(b[3680]), .B(n11042), .Z(c[3680]) );
XNOR U18404 ( .A(a[3680]), .B(c3680), .Z(n11042) );
XOR U18405 ( .A(c3681), .B(n11043), .Z(c3682) );
ANDN U18406 ( .B(n11044), .A(n11045), .Z(n11043) );
XOR U18407 ( .A(c3681), .B(b[3681]), .Z(n11044) );
XNOR U18408 ( .A(b[3681]), .B(n11045), .Z(c[3681]) );
XNOR U18409 ( .A(a[3681]), .B(c3681), .Z(n11045) );
XOR U18410 ( .A(c3682), .B(n11046), .Z(c3683) );
ANDN U18411 ( .B(n11047), .A(n11048), .Z(n11046) );
XOR U18412 ( .A(c3682), .B(b[3682]), .Z(n11047) );
XNOR U18413 ( .A(b[3682]), .B(n11048), .Z(c[3682]) );
XNOR U18414 ( .A(a[3682]), .B(c3682), .Z(n11048) );
XOR U18415 ( .A(c3683), .B(n11049), .Z(c3684) );
ANDN U18416 ( .B(n11050), .A(n11051), .Z(n11049) );
XOR U18417 ( .A(c3683), .B(b[3683]), .Z(n11050) );
XNOR U18418 ( .A(b[3683]), .B(n11051), .Z(c[3683]) );
XNOR U18419 ( .A(a[3683]), .B(c3683), .Z(n11051) );
XOR U18420 ( .A(c3684), .B(n11052), .Z(c3685) );
ANDN U18421 ( .B(n11053), .A(n11054), .Z(n11052) );
XOR U18422 ( .A(c3684), .B(b[3684]), .Z(n11053) );
XNOR U18423 ( .A(b[3684]), .B(n11054), .Z(c[3684]) );
XNOR U18424 ( .A(a[3684]), .B(c3684), .Z(n11054) );
XOR U18425 ( .A(c3685), .B(n11055), .Z(c3686) );
ANDN U18426 ( .B(n11056), .A(n11057), .Z(n11055) );
XOR U18427 ( .A(c3685), .B(b[3685]), .Z(n11056) );
XNOR U18428 ( .A(b[3685]), .B(n11057), .Z(c[3685]) );
XNOR U18429 ( .A(a[3685]), .B(c3685), .Z(n11057) );
XOR U18430 ( .A(c3686), .B(n11058), .Z(c3687) );
ANDN U18431 ( .B(n11059), .A(n11060), .Z(n11058) );
XOR U18432 ( .A(c3686), .B(b[3686]), .Z(n11059) );
XNOR U18433 ( .A(b[3686]), .B(n11060), .Z(c[3686]) );
XNOR U18434 ( .A(a[3686]), .B(c3686), .Z(n11060) );
XOR U18435 ( .A(c3687), .B(n11061), .Z(c3688) );
ANDN U18436 ( .B(n11062), .A(n11063), .Z(n11061) );
XOR U18437 ( .A(c3687), .B(b[3687]), .Z(n11062) );
XNOR U18438 ( .A(b[3687]), .B(n11063), .Z(c[3687]) );
XNOR U18439 ( .A(a[3687]), .B(c3687), .Z(n11063) );
XOR U18440 ( .A(c3688), .B(n11064), .Z(c3689) );
ANDN U18441 ( .B(n11065), .A(n11066), .Z(n11064) );
XOR U18442 ( .A(c3688), .B(b[3688]), .Z(n11065) );
XNOR U18443 ( .A(b[3688]), .B(n11066), .Z(c[3688]) );
XNOR U18444 ( .A(a[3688]), .B(c3688), .Z(n11066) );
XOR U18445 ( .A(c3689), .B(n11067), .Z(c3690) );
ANDN U18446 ( .B(n11068), .A(n11069), .Z(n11067) );
XOR U18447 ( .A(c3689), .B(b[3689]), .Z(n11068) );
XNOR U18448 ( .A(b[3689]), .B(n11069), .Z(c[3689]) );
XNOR U18449 ( .A(a[3689]), .B(c3689), .Z(n11069) );
XOR U18450 ( .A(c3690), .B(n11070), .Z(c3691) );
ANDN U18451 ( .B(n11071), .A(n11072), .Z(n11070) );
XOR U18452 ( .A(c3690), .B(b[3690]), .Z(n11071) );
XNOR U18453 ( .A(b[3690]), .B(n11072), .Z(c[3690]) );
XNOR U18454 ( .A(a[3690]), .B(c3690), .Z(n11072) );
XOR U18455 ( .A(c3691), .B(n11073), .Z(c3692) );
ANDN U18456 ( .B(n11074), .A(n11075), .Z(n11073) );
XOR U18457 ( .A(c3691), .B(b[3691]), .Z(n11074) );
XNOR U18458 ( .A(b[3691]), .B(n11075), .Z(c[3691]) );
XNOR U18459 ( .A(a[3691]), .B(c3691), .Z(n11075) );
XOR U18460 ( .A(c3692), .B(n11076), .Z(c3693) );
ANDN U18461 ( .B(n11077), .A(n11078), .Z(n11076) );
XOR U18462 ( .A(c3692), .B(b[3692]), .Z(n11077) );
XNOR U18463 ( .A(b[3692]), .B(n11078), .Z(c[3692]) );
XNOR U18464 ( .A(a[3692]), .B(c3692), .Z(n11078) );
XOR U18465 ( .A(c3693), .B(n11079), .Z(c3694) );
ANDN U18466 ( .B(n11080), .A(n11081), .Z(n11079) );
XOR U18467 ( .A(c3693), .B(b[3693]), .Z(n11080) );
XNOR U18468 ( .A(b[3693]), .B(n11081), .Z(c[3693]) );
XNOR U18469 ( .A(a[3693]), .B(c3693), .Z(n11081) );
XOR U18470 ( .A(c3694), .B(n11082), .Z(c3695) );
ANDN U18471 ( .B(n11083), .A(n11084), .Z(n11082) );
XOR U18472 ( .A(c3694), .B(b[3694]), .Z(n11083) );
XNOR U18473 ( .A(b[3694]), .B(n11084), .Z(c[3694]) );
XNOR U18474 ( .A(a[3694]), .B(c3694), .Z(n11084) );
XOR U18475 ( .A(c3695), .B(n11085), .Z(c3696) );
ANDN U18476 ( .B(n11086), .A(n11087), .Z(n11085) );
XOR U18477 ( .A(c3695), .B(b[3695]), .Z(n11086) );
XNOR U18478 ( .A(b[3695]), .B(n11087), .Z(c[3695]) );
XNOR U18479 ( .A(a[3695]), .B(c3695), .Z(n11087) );
XOR U18480 ( .A(c3696), .B(n11088), .Z(c3697) );
ANDN U18481 ( .B(n11089), .A(n11090), .Z(n11088) );
XOR U18482 ( .A(c3696), .B(b[3696]), .Z(n11089) );
XNOR U18483 ( .A(b[3696]), .B(n11090), .Z(c[3696]) );
XNOR U18484 ( .A(a[3696]), .B(c3696), .Z(n11090) );
XOR U18485 ( .A(c3697), .B(n11091), .Z(c3698) );
ANDN U18486 ( .B(n11092), .A(n11093), .Z(n11091) );
XOR U18487 ( .A(c3697), .B(b[3697]), .Z(n11092) );
XNOR U18488 ( .A(b[3697]), .B(n11093), .Z(c[3697]) );
XNOR U18489 ( .A(a[3697]), .B(c3697), .Z(n11093) );
XOR U18490 ( .A(c3698), .B(n11094), .Z(c3699) );
ANDN U18491 ( .B(n11095), .A(n11096), .Z(n11094) );
XOR U18492 ( .A(c3698), .B(b[3698]), .Z(n11095) );
XNOR U18493 ( .A(b[3698]), .B(n11096), .Z(c[3698]) );
XNOR U18494 ( .A(a[3698]), .B(c3698), .Z(n11096) );
XOR U18495 ( .A(c3699), .B(n11097), .Z(c3700) );
ANDN U18496 ( .B(n11098), .A(n11099), .Z(n11097) );
XOR U18497 ( .A(c3699), .B(b[3699]), .Z(n11098) );
XNOR U18498 ( .A(b[3699]), .B(n11099), .Z(c[3699]) );
XNOR U18499 ( .A(a[3699]), .B(c3699), .Z(n11099) );
XOR U18500 ( .A(c3700), .B(n11100), .Z(c3701) );
ANDN U18501 ( .B(n11101), .A(n11102), .Z(n11100) );
XOR U18502 ( .A(c3700), .B(b[3700]), .Z(n11101) );
XNOR U18503 ( .A(b[3700]), .B(n11102), .Z(c[3700]) );
XNOR U18504 ( .A(a[3700]), .B(c3700), .Z(n11102) );
XOR U18505 ( .A(c3701), .B(n11103), .Z(c3702) );
ANDN U18506 ( .B(n11104), .A(n11105), .Z(n11103) );
XOR U18507 ( .A(c3701), .B(b[3701]), .Z(n11104) );
XNOR U18508 ( .A(b[3701]), .B(n11105), .Z(c[3701]) );
XNOR U18509 ( .A(a[3701]), .B(c3701), .Z(n11105) );
XOR U18510 ( .A(c3702), .B(n11106), .Z(c3703) );
ANDN U18511 ( .B(n11107), .A(n11108), .Z(n11106) );
XOR U18512 ( .A(c3702), .B(b[3702]), .Z(n11107) );
XNOR U18513 ( .A(b[3702]), .B(n11108), .Z(c[3702]) );
XNOR U18514 ( .A(a[3702]), .B(c3702), .Z(n11108) );
XOR U18515 ( .A(c3703), .B(n11109), .Z(c3704) );
ANDN U18516 ( .B(n11110), .A(n11111), .Z(n11109) );
XOR U18517 ( .A(c3703), .B(b[3703]), .Z(n11110) );
XNOR U18518 ( .A(b[3703]), .B(n11111), .Z(c[3703]) );
XNOR U18519 ( .A(a[3703]), .B(c3703), .Z(n11111) );
XOR U18520 ( .A(c3704), .B(n11112), .Z(c3705) );
ANDN U18521 ( .B(n11113), .A(n11114), .Z(n11112) );
XOR U18522 ( .A(c3704), .B(b[3704]), .Z(n11113) );
XNOR U18523 ( .A(b[3704]), .B(n11114), .Z(c[3704]) );
XNOR U18524 ( .A(a[3704]), .B(c3704), .Z(n11114) );
XOR U18525 ( .A(c3705), .B(n11115), .Z(c3706) );
ANDN U18526 ( .B(n11116), .A(n11117), .Z(n11115) );
XOR U18527 ( .A(c3705), .B(b[3705]), .Z(n11116) );
XNOR U18528 ( .A(b[3705]), .B(n11117), .Z(c[3705]) );
XNOR U18529 ( .A(a[3705]), .B(c3705), .Z(n11117) );
XOR U18530 ( .A(c3706), .B(n11118), .Z(c3707) );
ANDN U18531 ( .B(n11119), .A(n11120), .Z(n11118) );
XOR U18532 ( .A(c3706), .B(b[3706]), .Z(n11119) );
XNOR U18533 ( .A(b[3706]), .B(n11120), .Z(c[3706]) );
XNOR U18534 ( .A(a[3706]), .B(c3706), .Z(n11120) );
XOR U18535 ( .A(c3707), .B(n11121), .Z(c3708) );
ANDN U18536 ( .B(n11122), .A(n11123), .Z(n11121) );
XOR U18537 ( .A(c3707), .B(b[3707]), .Z(n11122) );
XNOR U18538 ( .A(b[3707]), .B(n11123), .Z(c[3707]) );
XNOR U18539 ( .A(a[3707]), .B(c3707), .Z(n11123) );
XOR U18540 ( .A(c3708), .B(n11124), .Z(c3709) );
ANDN U18541 ( .B(n11125), .A(n11126), .Z(n11124) );
XOR U18542 ( .A(c3708), .B(b[3708]), .Z(n11125) );
XNOR U18543 ( .A(b[3708]), .B(n11126), .Z(c[3708]) );
XNOR U18544 ( .A(a[3708]), .B(c3708), .Z(n11126) );
XOR U18545 ( .A(c3709), .B(n11127), .Z(c3710) );
ANDN U18546 ( .B(n11128), .A(n11129), .Z(n11127) );
XOR U18547 ( .A(c3709), .B(b[3709]), .Z(n11128) );
XNOR U18548 ( .A(b[3709]), .B(n11129), .Z(c[3709]) );
XNOR U18549 ( .A(a[3709]), .B(c3709), .Z(n11129) );
XOR U18550 ( .A(c3710), .B(n11130), .Z(c3711) );
ANDN U18551 ( .B(n11131), .A(n11132), .Z(n11130) );
XOR U18552 ( .A(c3710), .B(b[3710]), .Z(n11131) );
XNOR U18553 ( .A(b[3710]), .B(n11132), .Z(c[3710]) );
XNOR U18554 ( .A(a[3710]), .B(c3710), .Z(n11132) );
XOR U18555 ( .A(c3711), .B(n11133), .Z(c3712) );
ANDN U18556 ( .B(n11134), .A(n11135), .Z(n11133) );
XOR U18557 ( .A(c3711), .B(b[3711]), .Z(n11134) );
XNOR U18558 ( .A(b[3711]), .B(n11135), .Z(c[3711]) );
XNOR U18559 ( .A(a[3711]), .B(c3711), .Z(n11135) );
XOR U18560 ( .A(c3712), .B(n11136), .Z(c3713) );
ANDN U18561 ( .B(n11137), .A(n11138), .Z(n11136) );
XOR U18562 ( .A(c3712), .B(b[3712]), .Z(n11137) );
XNOR U18563 ( .A(b[3712]), .B(n11138), .Z(c[3712]) );
XNOR U18564 ( .A(a[3712]), .B(c3712), .Z(n11138) );
XOR U18565 ( .A(c3713), .B(n11139), .Z(c3714) );
ANDN U18566 ( .B(n11140), .A(n11141), .Z(n11139) );
XOR U18567 ( .A(c3713), .B(b[3713]), .Z(n11140) );
XNOR U18568 ( .A(b[3713]), .B(n11141), .Z(c[3713]) );
XNOR U18569 ( .A(a[3713]), .B(c3713), .Z(n11141) );
XOR U18570 ( .A(c3714), .B(n11142), .Z(c3715) );
ANDN U18571 ( .B(n11143), .A(n11144), .Z(n11142) );
XOR U18572 ( .A(c3714), .B(b[3714]), .Z(n11143) );
XNOR U18573 ( .A(b[3714]), .B(n11144), .Z(c[3714]) );
XNOR U18574 ( .A(a[3714]), .B(c3714), .Z(n11144) );
XOR U18575 ( .A(c3715), .B(n11145), .Z(c3716) );
ANDN U18576 ( .B(n11146), .A(n11147), .Z(n11145) );
XOR U18577 ( .A(c3715), .B(b[3715]), .Z(n11146) );
XNOR U18578 ( .A(b[3715]), .B(n11147), .Z(c[3715]) );
XNOR U18579 ( .A(a[3715]), .B(c3715), .Z(n11147) );
XOR U18580 ( .A(c3716), .B(n11148), .Z(c3717) );
ANDN U18581 ( .B(n11149), .A(n11150), .Z(n11148) );
XOR U18582 ( .A(c3716), .B(b[3716]), .Z(n11149) );
XNOR U18583 ( .A(b[3716]), .B(n11150), .Z(c[3716]) );
XNOR U18584 ( .A(a[3716]), .B(c3716), .Z(n11150) );
XOR U18585 ( .A(c3717), .B(n11151), .Z(c3718) );
ANDN U18586 ( .B(n11152), .A(n11153), .Z(n11151) );
XOR U18587 ( .A(c3717), .B(b[3717]), .Z(n11152) );
XNOR U18588 ( .A(b[3717]), .B(n11153), .Z(c[3717]) );
XNOR U18589 ( .A(a[3717]), .B(c3717), .Z(n11153) );
XOR U18590 ( .A(c3718), .B(n11154), .Z(c3719) );
ANDN U18591 ( .B(n11155), .A(n11156), .Z(n11154) );
XOR U18592 ( .A(c3718), .B(b[3718]), .Z(n11155) );
XNOR U18593 ( .A(b[3718]), .B(n11156), .Z(c[3718]) );
XNOR U18594 ( .A(a[3718]), .B(c3718), .Z(n11156) );
XOR U18595 ( .A(c3719), .B(n11157), .Z(c3720) );
ANDN U18596 ( .B(n11158), .A(n11159), .Z(n11157) );
XOR U18597 ( .A(c3719), .B(b[3719]), .Z(n11158) );
XNOR U18598 ( .A(b[3719]), .B(n11159), .Z(c[3719]) );
XNOR U18599 ( .A(a[3719]), .B(c3719), .Z(n11159) );
XOR U18600 ( .A(c3720), .B(n11160), .Z(c3721) );
ANDN U18601 ( .B(n11161), .A(n11162), .Z(n11160) );
XOR U18602 ( .A(c3720), .B(b[3720]), .Z(n11161) );
XNOR U18603 ( .A(b[3720]), .B(n11162), .Z(c[3720]) );
XNOR U18604 ( .A(a[3720]), .B(c3720), .Z(n11162) );
XOR U18605 ( .A(c3721), .B(n11163), .Z(c3722) );
ANDN U18606 ( .B(n11164), .A(n11165), .Z(n11163) );
XOR U18607 ( .A(c3721), .B(b[3721]), .Z(n11164) );
XNOR U18608 ( .A(b[3721]), .B(n11165), .Z(c[3721]) );
XNOR U18609 ( .A(a[3721]), .B(c3721), .Z(n11165) );
XOR U18610 ( .A(c3722), .B(n11166), .Z(c3723) );
ANDN U18611 ( .B(n11167), .A(n11168), .Z(n11166) );
XOR U18612 ( .A(c3722), .B(b[3722]), .Z(n11167) );
XNOR U18613 ( .A(b[3722]), .B(n11168), .Z(c[3722]) );
XNOR U18614 ( .A(a[3722]), .B(c3722), .Z(n11168) );
XOR U18615 ( .A(c3723), .B(n11169), .Z(c3724) );
ANDN U18616 ( .B(n11170), .A(n11171), .Z(n11169) );
XOR U18617 ( .A(c3723), .B(b[3723]), .Z(n11170) );
XNOR U18618 ( .A(b[3723]), .B(n11171), .Z(c[3723]) );
XNOR U18619 ( .A(a[3723]), .B(c3723), .Z(n11171) );
XOR U18620 ( .A(c3724), .B(n11172), .Z(c3725) );
ANDN U18621 ( .B(n11173), .A(n11174), .Z(n11172) );
XOR U18622 ( .A(c3724), .B(b[3724]), .Z(n11173) );
XNOR U18623 ( .A(b[3724]), .B(n11174), .Z(c[3724]) );
XNOR U18624 ( .A(a[3724]), .B(c3724), .Z(n11174) );
XOR U18625 ( .A(c3725), .B(n11175), .Z(c3726) );
ANDN U18626 ( .B(n11176), .A(n11177), .Z(n11175) );
XOR U18627 ( .A(c3725), .B(b[3725]), .Z(n11176) );
XNOR U18628 ( .A(b[3725]), .B(n11177), .Z(c[3725]) );
XNOR U18629 ( .A(a[3725]), .B(c3725), .Z(n11177) );
XOR U18630 ( .A(c3726), .B(n11178), .Z(c3727) );
ANDN U18631 ( .B(n11179), .A(n11180), .Z(n11178) );
XOR U18632 ( .A(c3726), .B(b[3726]), .Z(n11179) );
XNOR U18633 ( .A(b[3726]), .B(n11180), .Z(c[3726]) );
XNOR U18634 ( .A(a[3726]), .B(c3726), .Z(n11180) );
XOR U18635 ( .A(c3727), .B(n11181), .Z(c3728) );
ANDN U18636 ( .B(n11182), .A(n11183), .Z(n11181) );
XOR U18637 ( .A(c3727), .B(b[3727]), .Z(n11182) );
XNOR U18638 ( .A(b[3727]), .B(n11183), .Z(c[3727]) );
XNOR U18639 ( .A(a[3727]), .B(c3727), .Z(n11183) );
XOR U18640 ( .A(c3728), .B(n11184), .Z(c3729) );
ANDN U18641 ( .B(n11185), .A(n11186), .Z(n11184) );
XOR U18642 ( .A(c3728), .B(b[3728]), .Z(n11185) );
XNOR U18643 ( .A(b[3728]), .B(n11186), .Z(c[3728]) );
XNOR U18644 ( .A(a[3728]), .B(c3728), .Z(n11186) );
XOR U18645 ( .A(c3729), .B(n11187), .Z(c3730) );
ANDN U18646 ( .B(n11188), .A(n11189), .Z(n11187) );
XOR U18647 ( .A(c3729), .B(b[3729]), .Z(n11188) );
XNOR U18648 ( .A(b[3729]), .B(n11189), .Z(c[3729]) );
XNOR U18649 ( .A(a[3729]), .B(c3729), .Z(n11189) );
XOR U18650 ( .A(c3730), .B(n11190), .Z(c3731) );
ANDN U18651 ( .B(n11191), .A(n11192), .Z(n11190) );
XOR U18652 ( .A(c3730), .B(b[3730]), .Z(n11191) );
XNOR U18653 ( .A(b[3730]), .B(n11192), .Z(c[3730]) );
XNOR U18654 ( .A(a[3730]), .B(c3730), .Z(n11192) );
XOR U18655 ( .A(c3731), .B(n11193), .Z(c3732) );
ANDN U18656 ( .B(n11194), .A(n11195), .Z(n11193) );
XOR U18657 ( .A(c3731), .B(b[3731]), .Z(n11194) );
XNOR U18658 ( .A(b[3731]), .B(n11195), .Z(c[3731]) );
XNOR U18659 ( .A(a[3731]), .B(c3731), .Z(n11195) );
XOR U18660 ( .A(c3732), .B(n11196), .Z(c3733) );
ANDN U18661 ( .B(n11197), .A(n11198), .Z(n11196) );
XOR U18662 ( .A(c3732), .B(b[3732]), .Z(n11197) );
XNOR U18663 ( .A(b[3732]), .B(n11198), .Z(c[3732]) );
XNOR U18664 ( .A(a[3732]), .B(c3732), .Z(n11198) );
XOR U18665 ( .A(c3733), .B(n11199), .Z(c3734) );
ANDN U18666 ( .B(n11200), .A(n11201), .Z(n11199) );
XOR U18667 ( .A(c3733), .B(b[3733]), .Z(n11200) );
XNOR U18668 ( .A(b[3733]), .B(n11201), .Z(c[3733]) );
XNOR U18669 ( .A(a[3733]), .B(c3733), .Z(n11201) );
XOR U18670 ( .A(c3734), .B(n11202), .Z(c3735) );
ANDN U18671 ( .B(n11203), .A(n11204), .Z(n11202) );
XOR U18672 ( .A(c3734), .B(b[3734]), .Z(n11203) );
XNOR U18673 ( .A(b[3734]), .B(n11204), .Z(c[3734]) );
XNOR U18674 ( .A(a[3734]), .B(c3734), .Z(n11204) );
XOR U18675 ( .A(c3735), .B(n11205), .Z(c3736) );
ANDN U18676 ( .B(n11206), .A(n11207), .Z(n11205) );
XOR U18677 ( .A(c3735), .B(b[3735]), .Z(n11206) );
XNOR U18678 ( .A(b[3735]), .B(n11207), .Z(c[3735]) );
XNOR U18679 ( .A(a[3735]), .B(c3735), .Z(n11207) );
XOR U18680 ( .A(c3736), .B(n11208), .Z(c3737) );
ANDN U18681 ( .B(n11209), .A(n11210), .Z(n11208) );
XOR U18682 ( .A(c3736), .B(b[3736]), .Z(n11209) );
XNOR U18683 ( .A(b[3736]), .B(n11210), .Z(c[3736]) );
XNOR U18684 ( .A(a[3736]), .B(c3736), .Z(n11210) );
XOR U18685 ( .A(c3737), .B(n11211), .Z(c3738) );
ANDN U18686 ( .B(n11212), .A(n11213), .Z(n11211) );
XOR U18687 ( .A(c3737), .B(b[3737]), .Z(n11212) );
XNOR U18688 ( .A(b[3737]), .B(n11213), .Z(c[3737]) );
XNOR U18689 ( .A(a[3737]), .B(c3737), .Z(n11213) );
XOR U18690 ( .A(c3738), .B(n11214), .Z(c3739) );
ANDN U18691 ( .B(n11215), .A(n11216), .Z(n11214) );
XOR U18692 ( .A(c3738), .B(b[3738]), .Z(n11215) );
XNOR U18693 ( .A(b[3738]), .B(n11216), .Z(c[3738]) );
XNOR U18694 ( .A(a[3738]), .B(c3738), .Z(n11216) );
XOR U18695 ( .A(c3739), .B(n11217), .Z(c3740) );
ANDN U18696 ( .B(n11218), .A(n11219), .Z(n11217) );
XOR U18697 ( .A(c3739), .B(b[3739]), .Z(n11218) );
XNOR U18698 ( .A(b[3739]), .B(n11219), .Z(c[3739]) );
XNOR U18699 ( .A(a[3739]), .B(c3739), .Z(n11219) );
XOR U18700 ( .A(c3740), .B(n11220), .Z(c3741) );
ANDN U18701 ( .B(n11221), .A(n11222), .Z(n11220) );
XOR U18702 ( .A(c3740), .B(b[3740]), .Z(n11221) );
XNOR U18703 ( .A(b[3740]), .B(n11222), .Z(c[3740]) );
XNOR U18704 ( .A(a[3740]), .B(c3740), .Z(n11222) );
XOR U18705 ( .A(c3741), .B(n11223), .Z(c3742) );
ANDN U18706 ( .B(n11224), .A(n11225), .Z(n11223) );
XOR U18707 ( .A(c3741), .B(b[3741]), .Z(n11224) );
XNOR U18708 ( .A(b[3741]), .B(n11225), .Z(c[3741]) );
XNOR U18709 ( .A(a[3741]), .B(c3741), .Z(n11225) );
XOR U18710 ( .A(c3742), .B(n11226), .Z(c3743) );
ANDN U18711 ( .B(n11227), .A(n11228), .Z(n11226) );
XOR U18712 ( .A(c3742), .B(b[3742]), .Z(n11227) );
XNOR U18713 ( .A(b[3742]), .B(n11228), .Z(c[3742]) );
XNOR U18714 ( .A(a[3742]), .B(c3742), .Z(n11228) );
XOR U18715 ( .A(c3743), .B(n11229), .Z(c3744) );
ANDN U18716 ( .B(n11230), .A(n11231), .Z(n11229) );
XOR U18717 ( .A(c3743), .B(b[3743]), .Z(n11230) );
XNOR U18718 ( .A(b[3743]), .B(n11231), .Z(c[3743]) );
XNOR U18719 ( .A(a[3743]), .B(c3743), .Z(n11231) );
XOR U18720 ( .A(c3744), .B(n11232), .Z(c3745) );
ANDN U18721 ( .B(n11233), .A(n11234), .Z(n11232) );
XOR U18722 ( .A(c3744), .B(b[3744]), .Z(n11233) );
XNOR U18723 ( .A(b[3744]), .B(n11234), .Z(c[3744]) );
XNOR U18724 ( .A(a[3744]), .B(c3744), .Z(n11234) );
XOR U18725 ( .A(c3745), .B(n11235), .Z(c3746) );
ANDN U18726 ( .B(n11236), .A(n11237), .Z(n11235) );
XOR U18727 ( .A(c3745), .B(b[3745]), .Z(n11236) );
XNOR U18728 ( .A(b[3745]), .B(n11237), .Z(c[3745]) );
XNOR U18729 ( .A(a[3745]), .B(c3745), .Z(n11237) );
XOR U18730 ( .A(c3746), .B(n11238), .Z(c3747) );
ANDN U18731 ( .B(n11239), .A(n11240), .Z(n11238) );
XOR U18732 ( .A(c3746), .B(b[3746]), .Z(n11239) );
XNOR U18733 ( .A(b[3746]), .B(n11240), .Z(c[3746]) );
XNOR U18734 ( .A(a[3746]), .B(c3746), .Z(n11240) );
XOR U18735 ( .A(c3747), .B(n11241), .Z(c3748) );
ANDN U18736 ( .B(n11242), .A(n11243), .Z(n11241) );
XOR U18737 ( .A(c3747), .B(b[3747]), .Z(n11242) );
XNOR U18738 ( .A(b[3747]), .B(n11243), .Z(c[3747]) );
XNOR U18739 ( .A(a[3747]), .B(c3747), .Z(n11243) );
XOR U18740 ( .A(c3748), .B(n11244), .Z(c3749) );
ANDN U18741 ( .B(n11245), .A(n11246), .Z(n11244) );
XOR U18742 ( .A(c3748), .B(b[3748]), .Z(n11245) );
XNOR U18743 ( .A(b[3748]), .B(n11246), .Z(c[3748]) );
XNOR U18744 ( .A(a[3748]), .B(c3748), .Z(n11246) );
XOR U18745 ( .A(c3749), .B(n11247), .Z(c3750) );
ANDN U18746 ( .B(n11248), .A(n11249), .Z(n11247) );
XOR U18747 ( .A(c3749), .B(b[3749]), .Z(n11248) );
XNOR U18748 ( .A(b[3749]), .B(n11249), .Z(c[3749]) );
XNOR U18749 ( .A(a[3749]), .B(c3749), .Z(n11249) );
XOR U18750 ( .A(c3750), .B(n11250), .Z(c3751) );
ANDN U18751 ( .B(n11251), .A(n11252), .Z(n11250) );
XOR U18752 ( .A(c3750), .B(b[3750]), .Z(n11251) );
XNOR U18753 ( .A(b[3750]), .B(n11252), .Z(c[3750]) );
XNOR U18754 ( .A(a[3750]), .B(c3750), .Z(n11252) );
XOR U18755 ( .A(c3751), .B(n11253), .Z(c3752) );
ANDN U18756 ( .B(n11254), .A(n11255), .Z(n11253) );
XOR U18757 ( .A(c3751), .B(b[3751]), .Z(n11254) );
XNOR U18758 ( .A(b[3751]), .B(n11255), .Z(c[3751]) );
XNOR U18759 ( .A(a[3751]), .B(c3751), .Z(n11255) );
XOR U18760 ( .A(c3752), .B(n11256), .Z(c3753) );
ANDN U18761 ( .B(n11257), .A(n11258), .Z(n11256) );
XOR U18762 ( .A(c3752), .B(b[3752]), .Z(n11257) );
XNOR U18763 ( .A(b[3752]), .B(n11258), .Z(c[3752]) );
XNOR U18764 ( .A(a[3752]), .B(c3752), .Z(n11258) );
XOR U18765 ( .A(c3753), .B(n11259), .Z(c3754) );
ANDN U18766 ( .B(n11260), .A(n11261), .Z(n11259) );
XOR U18767 ( .A(c3753), .B(b[3753]), .Z(n11260) );
XNOR U18768 ( .A(b[3753]), .B(n11261), .Z(c[3753]) );
XNOR U18769 ( .A(a[3753]), .B(c3753), .Z(n11261) );
XOR U18770 ( .A(c3754), .B(n11262), .Z(c3755) );
ANDN U18771 ( .B(n11263), .A(n11264), .Z(n11262) );
XOR U18772 ( .A(c3754), .B(b[3754]), .Z(n11263) );
XNOR U18773 ( .A(b[3754]), .B(n11264), .Z(c[3754]) );
XNOR U18774 ( .A(a[3754]), .B(c3754), .Z(n11264) );
XOR U18775 ( .A(c3755), .B(n11265), .Z(c3756) );
ANDN U18776 ( .B(n11266), .A(n11267), .Z(n11265) );
XOR U18777 ( .A(c3755), .B(b[3755]), .Z(n11266) );
XNOR U18778 ( .A(b[3755]), .B(n11267), .Z(c[3755]) );
XNOR U18779 ( .A(a[3755]), .B(c3755), .Z(n11267) );
XOR U18780 ( .A(c3756), .B(n11268), .Z(c3757) );
ANDN U18781 ( .B(n11269), .A(n11270), .Z(n11268) );
XOR U18782 ( .A(c3756), .B(b[3756]), .Z(n11269) );
XNOR U18783 ( .A(b[3756]), .B(n11270), .Z(c[3756]) );
XNOR U18784 ( .A(a[3756]), .B(c3756), .Z(n11270) );
XOR U18785 ( .A(c3757), .B(n11271), .Z(c3758) );
ANDN U18786 ( .B(n11272), .A(n11273), .Z(n11271) );
XOR U18787 ( .A(c3757), .B(b[3757]), .Z(n11272) );
XNOR U18788 ( .A(b[3757]), .B(n11273), .Z(c[3757]) );
XNOR U18789 ( .A(a[3757]), .B(c3757), .Z(n11273) );
XOR U18790 ( .A(c3758), .B(n11274), .Z(c3759) );
ANDN U18791 ( .B(n11275), .A(n11276), .Z(n11274) );
XOR U18792 ( .A(c3758), .B(b[3758]), .Z(n11275) );
XNOR U18793 ( .A(b[3758]), .B(n11276), .Z(c[3758]) );
XNOR U18794 ( .A(a[3758]), .B(c3758), .Z(n11276) );
XOR U18795 ( .A(c3759), .B(n11277), .Z(c3760) );
ANDN U18796 ( .B(n11278), .A(n11279), .Z(n11277) );
XOR U18797 ( .A(c3759), .B(b[3759]), .Z(n11278) );
XNOR U18798 ( .A(b[3759]), .B(n11279), .Z(c[3759]) );
XNOR U18799 ( .A(a[3759]), .B(c3759), .Z(n11279) );
XOR U18800 ( .A(c3760), .B(n11280), .Z(c3761) );
ANDN U18801 ( .B(n11281), .A(n11282), .Z(n11280) );
XOR U18802 ( .A(c3760), .B(b[3760]), .Z(n11281) );
XNOR U18803 ( .A(b[3760]), .B(n11282), .Z(c[3760]) );
XNOR U18804 ( .A(a[3760]), .B(c3760), .Z(n11282) );
XOR U18805 ( .A(c3761), .B(n11283), .Z(c3762) );
ANDN U18806 ( .B(n11284), .A(n11285), .Z(n11283) );
XOR U18807 ( .A(c3761), .B(b[3761]), .Z(n11284) );
XNOR U18808 ( .A(b[3761]), .B(n11285), .Z(c[3761]) );
XNOR U18809 ( .A(a[3761]), .B(c3761), .Z(n11285) );
XOR U18810 ( .A(c3762), .B(n11286), .Z(c3763) );
ANDN U18811 ( .B(n11287), .A(n11288), .Z(n11286) );
XOR U18812 ( .A(c3762), .B(b[3762]), .Z(n11287) );
XNOR U18813 ( .A(b[3762]), .B(n11288), .Z(c[3762]) );
XNOR U18814 ( .A(a[3762]), .B(c3762), .Z(n11288) );
XOR U18815 ( .A(c3763), .B(n11289), .Z(c3764) );
ANDN U18816 ( .B(n11290), .A(n11291), .Z(n11289) );
XOR U18817 ( .A(c3763), .B(b[3763]), .Z(n11290) );
XNOR U18818 ( .A(b[3763]), .B(n11291), .Z(c[3763]) );
XNOR U18819 ( .A(a[3763]), .B(c3763), .Z(n11291) );
XOR U18820 ( .A(c3764), .B(n11292), .Z(c3765) );
ANDN U18821 ( .B(n11293), .A(n11294), .Z(n11292) );
XOR U18822 ( .A(c3764), .B(b[3764]), .Z(n11293) );
XNOR U18823 ( .A(b[3764]), .B(n11294), .Z(c[3764]) );
XNOR U18824 ( .A(a[3764]), .B(c3764), .Z(n11294) );
XOR U18825 ( .A(c3765), .B(n11295), .Z(c3766) );
ANDN U18826 ( .B(n11296), .A(n11297), .Z(n11295) );
XOR U18827 ( .A(c3765), .B(b[3765]), .Z(n11296) );
XNOR U18828 ( .A(b[3765]), .B(n11297), .Z(c[3765]) );
XNOR U18829 ( .A(a[3765]), .B(c3765), .Z(n11297) );
XOR U18830 ( .A(c3766), .B(n11298), .Z(c3767) );
ANDN U18831 ( .B(n11299), .A(n11300), .Z(n11298) );
XOR U18832 ( .A(c3766), .B(b[3766]), .Z(n11299) );
XNOR U18833 ( .A(b[3766]), .B(n11300), .Z(c[3766]) );
XNOR U18834 ( .A(a[3766]), .B(c3766), .Z(n11300) );
XOR U18835 ( .A(c3767), .B(n11301), .Z(c3768) );
ANDN U18836 ( .B(n11302), .A(n11303), .Z(n11301) );
XOR U18837 ( .A(c3767), .B(b[3767]), .Z(n11302) );
XNOR U18838 ( .A(b[3767]), .B(n11303), .Z(c[3767]) );
XNOR U18839 ( .A(a[3767]), .B(c3767), .Z(n11303) );
XOR U18840 ( .A(c3768), .B(n11304), .Z(c3769) );
ANDN U18841 ( .B(n11305), .A(n11306), .Z(n11304) );
XOR U18842 ( .A(c3768), .B(b[3768]), .Z(n11305) );
XNOR U18843 ( .A(b[3768]), .B(n11306), .Z(c[3768]) );
XNOR U18844 ( .A(a[3768]), .B(c3768), .Z(n11306) );
XOR U18845 ( .A(c3769), .B(n11307), .Z(c3770) );
ANDN U18846 ( .B(n11308), .A(n11309), .Z(n11307) );
XOR U18847 ( .A(c3769), .B(b[3769]), .Z(n11308) );
XNOR U18848 ( .A(b[3769]), .B(n11309), .Z(c[3769]) );
XNOR U18849 ( .A(a[3769]), .B(c3769), .Z(n11309) );
XOR U18850 ( .A(c3770), .B(n11310), .Z(c3771) );
ANDN U18851 ( .B(n11311), .A(n11312), .Z(n11310) );
XOR U18852 ( .A(c3770), .B(b[3770]), .Z(n11311) );
XNOR U18853 ( .A(b[3770]), .B(n11312), .Z(c[3770]) );
XNOR U18854 ( .A(a[3770]), .B(c3770), .Z(n11312) );
XOR U18855 ( .A(c3771), .B(n11313), .Z(c3772) );
ANDN U18856 ( .B(n11314), .A(n11315), .Z(n11313) );
XOR U18857 ( .A(c3771), .B(b[3771]), .Z(n11314) );
XNOR U18858 ( .A(b[3771]), .B(n11315), .Z(c[3771]) );
XNOR U18859 ( .A(a[3771]), .B(c3771), .Z(n11315) );
XOR U18860 ( .A(c3772), .B(n11316), .Z(c3773) );
ANDN U18861 ( .B(n11317), .A(n11318), .Z(n11316) );
XOR U18862 ( .A(c3772), .B(b[3772]), .Z(n11317) );
XNOR U18863 ( .A(b[3772]), .B(n11318), .Z(c[3772]) );
XNOR U18864 ( .A(a[3772]), .B(c3772), .Z(n11318) );
XOR U18865 ( .A(c3773), .B(n11319), .Z(c3774) );
ANDN U18866 ( .B(n11320), .A(n11321), .Z(n11319) );
XOR U18867 ( .A(c3773), .B(b[3773]), .Z(n11320) );
XNOR U18868 ( .A(b[3773]), .B(n11321), .Z(c[3773]) );
XNOR U18869 ( .A(a[3773]), .B(c3773), .Z(n11321) );
XOR U18870 ( .A(c3774), .B(n11322), .Z(c3775) );
ANDN U18871 ( .B(n11323), .A(n11324), .Z(n11322) );
XOR U18872 ( .A(c3774), .B(b[3774]), .Z(n11323) );
XNOR U18873 ( .A(b[3774]), .B(n11324), .Z(c[3774]) );
XNOR U18874 ( .A(a[3774]), .B(c3774), .Z(n11324) );
XOR U18875 ( .A(c3775), .B(n11325), .Z(c3776) );
ANDN U18876 ( .B(n11326), .A(n11327), .Z(n11325) );
XOR U18877 ( .A(c3775), .B(b[3775]), .Z(n11326) );
XNOR U18878 ( .A(b[3775]), .B(n11327), .Z(c[3775]) );
XNOR U18879 ( .A(a[3775]), .B(c3775), .Z(n11327) );
XOR U18880 ( .A(c3776), .B(n11328), .Z(c3777) );
ANDN U18881 ( .B(n11329), .A(n11330), .Z(n11328) );
XOR U18882 ( .A(c3776), .B(b[3776]), .Z(n11329) );
XNOR U18883 ( .A(b[3776]), .B(n11330), .Z(c[3776]) );
XNOR U18884 ( .A(a[3776]), .B(c3776), .Z(n11330) );
XOR U18885 ( .A(c3777), .B(n11331), .Z(c3778) );
ANDN U18886 ( .B(n11332), .A(n11333), .Z(n11331) );
XOR U18887 ( .A(c3777), .B(b[3777]), .Z(n11332) );
XNOR U18888 ( .A(b[3777]), .B(n11333), .Z(c[3777]) );
XNOR U18889 ( .A(a[3777]), .B(c3777), .Z(n11333) );
XOR U18890 ( .A(c3778), .B(n11334), .Z(c3779) );
ANDN U18891 ( .B(n11335), .A(n11336), .Z(n11334) );
XOR U18892 ( .A(c3778), .B(b[3778]), .Z(n11335) );
XNOR U18893 ( .A(b[3778]), .B(n11336), .Z(c[3778]) );
XNOR U18894 ( .A(a[3778]), .B(c3778), .Z(n11336) );
XOR U18895 ( .A(c3779), .B(n11337), .Z(c3780) );
ANDN U18896 ( .B(n11338), .A(n11339), .Z(n11337) );
XOR U18897 ( .A(c3779), .B(b[3779]), .Z(n11338) );
XNOR U18898 ( .A(b[3779]), .B(n11339), .Z(c[3779]) );
XNOR U18899 ( .A(a[3779]), .B(c3779), .Z(n11339) );
XOR U18900 ( .A(c3780), .B(n11340), .Z(c3781) );
ANDN U18901 ( .B(n11341), .A(n11342), .Z(n11340) );
XOR U18902 ( .A(c3780), .B(b[3780]), .Z(n11341) );
XNOR U18903 ( .A(b[3780]), .B(n11342), .Z(c[3780]) );
XNOR U18904 ( .A(a[3780]), .B(c3780), .Z(n11342) );
XOR U18905 ( .A(c3781), .B(n11343), .Z(c3782) );
ANDN U18906 ( .B(n11344), .A(n11345), .Z(n11343) );
XOR U18907 ( .A(c3781), .B(b[3781]), .Z(n11344) );
XNOR U18908 ( .A(b[3781]), .B(n11345), .Z(c[3781]) );
XNOR U18909 ( .A(a[3781]), .B(c3781), .Z(n11345) );
XOR U18910 ( .A(c3782), .B(n11346), .Z(c3783) );
ANDN U18911 ( .B(n11347), .A(n11348), .Z(n11346) );
XOR U18912 ( .A(c3782), .B(b[3782]), .Z(n11347) );
XNOR U18913 ( .A(b[3782]), .B(n11348), .Z(c[3782]) );
XNOR U18914 ( .A(a[3782]), .B(c3782), .Z(n11348) );
XOR U18915 ( .A(c3783), .B(n11349), .Z(c3784) );
ANDN U18916 ( .B(n11350), .A(n11351), .Z(n11349) );
XOR U18917 ( .A(c3783), .B(b[3783]), .Z(n11350) );
XNOR U18918 ( .A(b[3783]), .B(n11351), .Z(c[3783]) );
XNOR U18919 ( .A(a[3783]), .B(c3783), .Z(n11351) );
XOR U18920 ( .A(c3784), .B(n11352), .Z(c3785) );
ANDN U18921 ( .B(n11353), .A(n11354), .Z(n11352) );
XOR U18922 ( .A(c3784), .B(b[3784]), .Z(n11353) );
XNOR U18923 ( .A(b[3784]), .B(n11354), .Z(c[3784]) );
XNOR U18924 ( .A(a[3784]), .B(c3784), .Z(n11354) );
XOR U18925 ( .A(c3785), .B(n11355), .Z(c3786) );
ANDN U18926 ( .B(n11356), .A(n11357), .Z(n11355) );
XOR U18927 ( .A(c3785), .B(b[3785]), .Z(n11356) );
XNOR U18928 ( .A(b[3785]), .B(n11357), .Z(c[3785]) );
XNOR U18929 ( .A(a[3785]), .B(c3785), .Z(n11357) );
XOR U18930 ( .A(c3786), .B(n11358), .Z(c3787) );
ANDN U18931 ( .B(n11359), .A(n11360), .Z(n11358) );
XOR U18932 ( .A(c3786), .B(b[3786]), .Z(n11359) );
XNOR U18933 ( .A(b[3786]), .B(n11360), .Z(c[3786]) );
XNOR U18934 ( .A(a[3786]), .B(c3786), .Z(n11360) );
XOR U18935 ( .A(c3787), .B(n11361), .Z(c3788) );
ANDN U18936 ( .B(n11362), .A(n11363), .Z(n11361) );
XOR U18937 ( .A(c3787), .B(b[3787]), .Z(n11362) );
XNOR U18938 ( .A(b[3787]), .B(n11363), .Z(c[3787]) );
XNOR U18939 ( .A(a[3787]), .B(c3787), .Z(n11363) );
XOR U18940 ( .A(c3788), .B(n11364), .Z(c3789) );
ANDN U18941 ( .B(n11365), .A(n11366), .Z(n11364) );
XOR U18942 ( .A(c3788), .B(b[3788]), .Z(n11365) );
XNOR U18943 ( .A(b[3788]), .B(n11366), .Z(c[3788]) );
XNOR U18944 ( .A(a[3788]), .B(c3788), .Z(n11366) );
XOR U18945 ( .A(c3789), .B(n11367), .Z(c3790) );
ANDN U18946 ( .B(n11368), .A(n11369), .Z(n11367) );
XOR U18947 ( .A(c3789), .B(b[3789]), .Z(n11368) );
XNOR U18948 ( .A(b[3789]), .B(n11369), .Z(c[3789]) );
XNOR U18949 ( .A(a[3789]), .B(c3789), .Z(n11369) );
XOR U18950 ( .A(c3790), .B(n11370), .Z(c3791) );
ANDN U18951 ( .B(n11371), .A(n11372), .Z(n11370) );
XOR U18952 ( .A(c3790), .B(b[3790]), .Z(n11371) );
XNOR U18953 ( .A(b[3790]), .B(n11372), .Z(c[3790]) );
XNOR U18954 ( .A(a[3790]), .B(c3790), .Z(n11372) );
XOR U18955 ( .A(c3791), .B(n11373), .Z(c3792) );
ANDN U18956 ( .B(n11374), .A(n11375), .Z(n11373) );
XOR U18957 ( .A(c3791), .B(b[3791]), .Z(n11374) );
XNOR U18958 ( .A(b[3791]), .B(n11375), .Z(c[3791]) );
XNOR U18959 ( .A(a[3791]), .B(c3791), .Z(n11375) );
XOR U18960 ( .A(c3792), .B(n11376), .Z(c3793) );
ANDN U18961 ( .B(n11377), .A(n11378), .Z(n11376) );
XOR U18962 ( .A(c3792), .B(b[3792]), .Z(n11377) );
XNOR U18963 ( .A(b[3792]), .B(n11378), .Z(c[3792]) );
XNOR U18964 ( .A(a[3792]), .B(c3792), .Z(n11378) );
XOR U18965 ( .A(c3793), .B(n11379), .Z(c3794) );
ANDN U18966 ( .B(n11380), .A(n11381), .Z(n11379) );
XOR U18967 ( .A(c3793), .B(b[3793]), .Z(n11380) );
XNOR U18968 ( .A(b[3793]), .B(n11381), .Z(c[3793]) );
XNOR U18969 ( .A(a[3793]), .B(c3793), .Z(n11381) );
XOR U18970 ( .A(c3794), .B(n11382), .Z(c3795) );
ANDN U18971 ( .B(n11383), .A(n11384), .Z(n11382) );
XOR U18972 ( .A(c3794), .B(b[3794]), .Z(n11383) );
XNOR U18973 ( .A(b[3794]), .B(n11384), .Z(c[3794]) );
XNOR U18974 ( .A(a[3794]), .B(c3794), .Z(n11384) );
XOR U18975 ( .A(c3795), .B(n11385), .Z(c3796) );
ANDN U18976 ( .B(n11386), .A(n11387), .Z(n11385) );
XOR U18977 ( .A(c3795), .B(b[3795]), .Z(n11386) );
XNOR U18978 ( .A(b[3795]), .B(n11387), .Z(c[3795]) );
XNOR U18979 ( .A(a[3795]), .B(c3795), .Z(n11387) );
XOR U18980 ( .A(c3796), .B(n11388), .Z(c3797) );
ANDN U18981 ( .B(n11389), .A(n11390), .Z(n11388) );
XOR U18982 ( .A(c3796), .B(b[3796]), .Z(n11389) );
XNOR U18983 ( .A(b[3796]), .B(n11390), .Z(c[3796]) );
XNOR U18984 ( .A(a[3796]), .B(c3796), .Z(n11390) );
XOR U18985 ( .A(c3797), .B(n11391), .Z(c3798) );
ANDN U18986 ( .B(n11392), .A(n11393), .Z(n11391) );
XOR U18987 ( .A(c3797), .B(b[3797]), .Z(n11392) );
XNOR U18988 ( .A(b[3797]), .B(n11393), .Z(c[3797]) );
XNOR U18989 ( .A(a[3797]), .B(c3797), .Z(n11393) );
XOR U18990 ( .A(c3798), .B(n11394), .Z(c3799) );
ANDN U18991 ( .B(n11395), .A(n11396), .Z(n11394) );
XOR U18992 ( .A(c3798), .B(b[3798]), .Z(n11395) );
XNOR U18993 ( .A(b[3798]), .B(n11396), .Z(c[3798]) );
XNOR U18994 ( .A(a[3798]), .B(c3798), .Z(n11396) );
XOR U18995 ( .A(c3799), .B(n11397), .Z(c3800) );
ANDN U18996 ( .B(n11398), .A(n11399), .Z(n11397) );
XOR U18997 ( .A(c3799), .B(b[3799]), .Z(n11398) );
XNOR U18998 ( .A(b[3799]), .B(n11399), .Z(c[3799]) );
XNOR U18999 ( .A(a[3799]), .B(c3799), .Z(n11399) );
XOR U19000 ( .A(c3800), .B(n11400), .Z(c3801) );
ANDN U19001 ( .B(n11401), .A(n11402), .Z(n11400) );
XOR U19002 ( .A(c3800), .B(b[3800]), .Z(n11401) );
XNOR U19003 ( .A(b[3800]), .B(n11402), .Z(c[3800]) );
XNOR U19004 ( .A(a[3800]), .B(c3800), .Z(n11402) );
XOR U19005 ( .A(c3801), .B(n11403), .Z(c3802) );
ANDN U19006 ( .B(n11404), .A(n11405), .Z(n11403) );
XOR U19007 ( .A(c3801), .B(b[3801]), .Z(n11404) );
XNOR U19008 ( .A(b[3801]), .B(n11405), .Z(c[3801]) );
XNOR U19009 ( .A(a[3801]), .B(c3801), .Z(n11405) );
XOR U19010 ( .A(c3802), .B(n11406), .Z(c3803) );
ANDN U19011 ( .B(n11407), .A(n11408), .Z(n11406) );
XOR U19012 ( .A(c3802), .B(b[3802]), .Z(n11407) );
XNOR U19013 ( .A(b[3802]), .B(n11408), .Z(c[3802]) );
XNOR U19014 ( .A(a[3802]), .B(c3802), .Z(n11408) );
XOR U19015 ( .A(c3803), .B(n11409), .Z(c3804) );
ANDN U19016 ( .B(n11410), .A(n11411), .Z(n11409) );
XOR U19017 ( .A(c3803), .B(b[3803]), .Z(n11410) );
XNOR U19018 ( .A(b[3803]), .B(n11411), .Z(c[3803]) );
XNOR U19019 ( .A(a[3803]), .B(c3803), .Z(n11411) );
XOR U19020 ( .A(c3804), .B(n11412), .Z(c3805) );
ANDN U19021 ( .B(n11413), .A(n11414), .Z(n11412) );
XOR U19022 ( .A(c3804), .B(b[3804]), .Z(n11413) );
XNOR U19023 ( .A(b[3804]), .B(n11414), .Z(c[3804]) );
XNOR U19024 ( .A(a[3804]), .B(c3804), .Z(n11414) );
XOR U19025 ( .A(c3805), .B(n11415), .Z(c3806) );
ANDN U19026 ( .B(n11416), .A(n11417), .Z(n11415) );
XOR U19027 ( .A(c3805), .B(b[3805]), .Z(n11416) );
XNOR U19028 ( .A(b[3805]), .B(n11417), .Z(c[3805]) );
XNOR U19029 ( .A(a[3805]), .B(c3805), .Z(n11417) );
XOR U19030 ( .A(c3806), .B(n11418), .Z(c3807) );
ANDN U19031 ( .B(n11419), .A(n11420), .Z(n11418) );
XOR U19032 ( .A(c3806), .B(b[3806]), .Z(n11419) );
XNOR U19033 ( .A(b[3806]), .B(n11420), .Z(c[3806]) );
XNOR U19034 ( .A(a[3806]), .B(c3806), .Z(n11420) );
XOR U19035 ( .A(c3807), .B(n11421), .Z(c3808) );
ANDN U19036 ( .B(n11422), .A(n11423), .Z(n11421) );
XOR U19037 ( .A(c3807), .B(b[3807]), .Z(n11422) );
XNOR U19038 ( .A(b[3807]), .B(n11423), .Z(c[3807]) );
XNOR U19039 ( .A(a[3807]), .B(c3807), .Z(n11423) );
XOR U19040 ( .A(c3808), .B(n11424), .Z(c3809) );
ANDN U19041 ( .B(n11425), .A(n11426), .Z(n11424) );
XOR U19042 ( .A(c3808), .B(b[3808]), .Z(n11425) );
XNOR U19043 ( .A(b[3808]), .B(n11426), .Z(c[3808]) );
XNOR U19044 ( .A(a[3808]), .B(c3808), .Z(n11426) );
XOR U19045 ( .A(c3809), .B(n11427), .Z(c3810) );
ANDN U19046 ( .B(n11428), .A(n11429), .Z(n11427) );
XOR U19047 ( .A(c3809), .B(b[3809]), .Z(n11428) );
XNOR U19048 ( .A(b[3809]), .B(n11429), .Z(c[3809]) );
XNOR U19049 ( .A(a[3809]), .B(c3809), .Z(n11429) );
XOR U19050 ( .A(c3810), .B(n11430), .Z(c3811) );
ANDN U19051 ( .B(n11431), .A(n11432), .Z(n11430) );
XOR U19052 ( .A(c3810), .B(b[3810]), .Z(n11431) );
XNOR U19053 ( .A(b[3810]), .B(n11432), .Z(c[3810]) );
XNOR U19054 ( .A(a[3810]), .B(c3810), .Z(n11432) );
XOR U19055 ( .A(c3811), .B(n11433), .Z(c3812) );
ANDN U19056 ( .B(n11434), .A(n11435), .Z(n11433) );
XOR U19057 ( .A(c3811), .B(b[3811]), .Z(n11434) );
XNOR U19058 ( .A(b[3811]), .B(n11435), .Z(c[3811]) );
XNOR U19059 ( .A(a[3811]), .B(c3811), .Z(n11435) );
XOR U19060 ( .A(c3812), .B(n11436), .Z(c3813) );
ANDN U19061 ( .B(n11437), .A(n11438), .Z(n11436) );
XOR U19062 ( .A(c3812), .B(b[3812]), .Z(n11437) );
XNOR U19063 ( .A(b[3812]), .B(n11438), .Z(c[3812]) );
XNOR U19064 ( .A(a[3812]), .B(c3812), .Z(n11438) );
XOR U19065 ( .A(c3813), .B(n11439), .Z(c3814) );
ANDN U19066 ( .B(n11440), .A(n11441), .Z(n11439) );
XOR U19067 ( .A(c3813), .B(b[3813]), .Z(n11440) );
XNOR U19068 ( .A(b[3813]), .B(n11441), .Z(c[3813]) );
XNOR U19069 ( .A(a[3813]), .B(c3813), .Z(n11441) );
XOR U19070 ( .A(c3814), .B(n11442), .Z(c3815) );
ANDN U19071 ( .B(n11443), .A(n11444), .Z(n11442) );
XOR U19072 ( .A(c3814), .B(b[3814]), .Z(n11443) );
XNOR U19073 ( .A(b[3814]), .B(n11444), .Z(c[3814]) );
XNOR U19074 ( .A(a[3814]), .B(c3814), .Z(n11444) );
XOR U19075 ( .A(c3815), .B(n11445), .Z(c3816) );
ANDN U19076 ( .B(n11446), .A(n11447), .Z(n11445) );
XOR U19077 ( .A(c3815), .B(b[3815]), .Z(n11446) );
XNOR U19078 ( .A(b[3815]), .B(n11447), .Z(c[3815]) );
XNOR U19079 ( .A(a[3815]), .B(c3815), .Z(n11447) );
XOR U19080 ( .A(c3816), .B(n11448), .Z(c3817) );
ANDN U19081 ( .B(n11449), .A(n11450), .Z(n11448) );
XOR U19082 ( .A(c3816), .B(b[3816]), .Z(n11449) );
XNOR U19083 ( .A(b[3816]), .B(n11450), .Z(c[3816]) );
XNOR U19084 ( .A(a[3816]), .B(c3816), .Z(n11450) );
XOR U19085 ( .A(c3817), .B(n11451), .Z(c3818) );
ANDN U19086 ( .B(n11452), .A(n11453), .Z(n11451) );
XOR U19087 ( .A(c3817), .B(b[3817]), .Z(n11452) );
XNOR U19088 ( .A(b[3817]), .B(n11453), .Z(c[3817]) );
XNOR U19089 ( .A(a[3817]), .B(c3817), .Z(n11453) );
XOR U19090 ( .A(c3818), .B(n11454), .Z(c3819) );
ANDN U19091 ( .B(n11455), .A(n11456), .Z(n11454) );
XOR U19092 ( .A(c3818), .B(b[3818]), .Z(n11455) );
XNOR U19093 ( .A(b[3818]), .B(n11456), .Z(c[3818]) );
XNOR U19094 ( .A(a[3818]), .B(c3818), .Z(n11456) );
XOR U19095 ( .A(c3819), .B(n11457), .Z(c3820) );
ANDN U19096 ( .B(n11458), .A(n11459), .Z(n11457) );
XOR U19097 ( .A(c3819), .B(b[3819]), .Z(n11458) );
XNOR U19098 ( .A(b[3819]), .B(n11459), .Z(c[3819]) );
XNOR U19099 ( .A(a[3819]), .B(c3819), .Z(n11459) );
XOR U19100 ( .A(c3820), .B(n11460), .Z(c3821) );
ANDN U19101 ( .B(n11461), .A(n11462), .Z(n11460) );
XOR U19102 ( .A(c3820), .B(b[3820]), .Z(n11461) );
XNOR U19103 ( .A(b[3820]), .B(n11462), .Z(c[3820]) );
XNOR U19104 ( .A(a[3820]), .B(c3820), .Z(n11462) );
XOR U19105 ( .A(c3821), .B(n11463), .Z(c3822) );
ANDN U19106 ( .B(n11464), .A(n11465), .Z(n11463) );
XOR U19107 ( .A(c3821), .B(b[3821]), .Z(n11464) );
XNOR U19108 ( .A(b[3821]), .B(n11465), .Z(c[3821]) );
XNOR U19109 ( .A(a[3821]), .B(c3821), .Z(n11465) );
XOR U19110 ( .A(c3822), .B(n11466), .Z(c3823) );
ANDN U19111 ( .B(n11467), .A(n11468), .Z(n11466) );
XOR U19112 ( .A(c3822), .B(b[3822]), .Z(n11467) );
XNOR U19113 ( .A(b[3822]), .B(n11468), .Z(c[3822]) );
XNOR U19114 ( .A(a[3822]), .B(c3822), .Z(n11468) );
XOR U19115 ( .A(c3823), .B(n11469), .Z(c3824) );
ANDN U19116 ( .B(n11470), .A(n11471), .Z(n11469) );
XOR U19117 ( .A(c3823), .B(b[3823]), .Z(n11470) );
XNOR U19118 ( .A(b[3823]), .B(n11471), .Z(c[3823]) );
XNOR U19119 ( .A(a[3823]), .B(c3823), .Z(n11471) );
XOR U19120 ( .A(c3824), .B(n11472), .Z(c3825) );
ANDN U19121 ( .B(n11473), .A(n11474), .Z(n11472) );
XOR U19122 ( .A(c3824), .B(b[3824]), .Z(n11473) );
XNOR U19123 ( .A(b[3824]), .B(n11474), .Z(c[3824]) );
XNOR U19124 ( .A(a[3824]), .B(c3824), .Z(n11474) );
XOR U19125 ( .A(c3825), .B(n11475), .Z(c3826) );
ANDN U19126 ( .B(n11476), .A(n11477), .Z(n11475) );
XOR U19127 ( .A(c3825), .B(b[3825]), .Z(n11476) );
XNOR U19128 ( .A(b[3825]), .B(n11477), .Z(c[3825]) );
XNOR U19129 ( .A(a[3825]), .B(c3825), .Z(n11477) );
XOR U19130 ( .A(c3826), .B(n11478), .Z(c3827) );
ANDN U19131 ( .B(n11479), .A(n11480), .Z(n11478) );
XOR U19132 ( .A(c3826), .B(b[3826]), .Z(n11479) );
XNOR U19133 ( .A(b[3826]), .B(n11480), .Z(c[3826]) );
XNOR U19134 ( .A(a[3826]), .B(c3826), .Z(n11480) );
XOR U19135 ( .A(c3827), .B(n11481), .Z(c3828) );
ANDN U19136 ( .B(n11482), .A(n11483), .Z(n11481) );
XOR U19137 ( .A(c3827), .B(b[3827]), .Z(n11482) );
XNOR U19138 ( .A(b[3827]), .B(n11483), .Z(c[3827]) );
XNOR U19139 ( .A(a[3827]), .B(c3827), .Z(n11483) );
XOR U19140 ( .A(c3828), .B(n11484), .Z(c3829) );
ANDN U19141 ( .B(n11485), .A(n11486), .Z(n11484) );
XOR U19142 ( .A(c3828), .B(b[3828]), .Z(n11485) );
XNOR U19143 ( .A(b[3828]), .B(n11486), .Z(c[3828]) );
XNOR U19144 ( .A(a[3828]), .B(c3828), .Z(n11486) );
XOR U19145 ( .A(c3829), .B(n11487), .Z(c3830) );
ANDN U19146 ( .B(n11488), .A(n11489), .Z(n11487) );
XOR U19147 ( .A(c3829), .B(b[3829]), .Z(n11488) );
XNOR U19148 ( .A(b[3829]), .B(n11489), .Z(c[3829]) );
XNOR U19149 ( .A(a[3829]), .B(c3829), .Z(n11489) );
XOR U19150 ( .A(c3830), .B(n11490), .Z(c3831) );
ANDN U19151 ( .B(n11491), .A(n11492), .Z(n11490) );
XOR U19152 ( .A(c3830), .B(b[3830]), .Z(n11491) );
XNOR U19153 ( .A(b[3830]), .B(n11492), .Z(c[3830]) );
XNOR U19154 ( .A(a[3830]), .B(c3830), .Z(n11492) );
XOR U19155 ( .A(c3831), .B(n11493), .Z(c3832) );
ANDN U19156 ( .B(n11494), .A(n11495), .Z(n11493) );
XOR U19157 ( .A(c3831), .B(b[3831]), .Z(n11494) );
XNOR U19158 ( .A(b[3831]), .B(n11495), .Z(c[3831]) );
XNOR U19159 ( .A(a[3831]), .B(c3831), .Z(n11495) );
XOR U19160 ( .A(c3832), .B(n11496), .Z(c3833) );
ANDN U19161 ( .B(n11497), .A(n11498), .Z(n11496) );
XOR U19162 ( .A(c3832), .B(b[3832]), .Z(n11497) );
XNOR U19163 ( .A(b[3832]), .B(n11498), .Z(c[3832]) );
XNOR U19164 ( .A(a[3832]), .B(c3832), .Z(n11498) );
XOR U19165 ( .A(c3833), .B(n11499), .Z(c3834) );
ANDN U19166 ( .B(n11500), .A(n11501), .Z(n11499) );
XOR U19167 ( .A(c3833), .B(b[3833]), .Z(n11500) );
XNOR U19168 ( .A(b[3833]), .B(n11501), .Z(c[3833]) );
XNOR U19169 ( .A(a[3833]), .B(c3833), .Z(n11501) );
XOR U19170 ( .A(c3834), .B(n11502), .Z(c3835) );
ANDN U19171 ( .B(n11503), .A(n11504), .Z(n11502) );
XOR U19172 ( .A(c3834), .B(b[3834]), .Z(n11503) );
XNOR U19173 ( .A(b[3834]), .B(n11504), .Z(c[3834]) );
XNOR U19174 ( .A(a[3834]), .B(c3834), .Z(n11504) );
XOR U19175 ( .A(c3835), .B(n11505), .Z(c3836) );
ANDN U19176 ( .B(n11506), .A(n11507), .Z(n11505) );
XOR U19177 ( .A(c3835), .B(b[3835]), .Z(n11506) );
XNOR U19178 ( .A(b[3835]), .B(n11507), .Z(c[3835]) );
XNOR U19179 ( .A(a[3835]), .B(c3835), .Z(n11507) );
XOR U19180 ( .A(c3836), .B(n11508), .Z(c3837) );
ANDN U19181 ( .B(n11509), .A(n11510), .Z(n11508) );
XOR U19182 ( .A(c3836), .B(b[3836]), .Z(n11509) );
XNOR U19183 ( .A(b[3836]), .B(n11510), .Z(c[3836]) );
XNOR U19184 ( .A(a[3836]), .B(c3836), .Z(n11510) );
XOR U19185 ( .A(c3837), .B(n11511), .Z(c3838) );
ANDN U19186 ( .B(n11512), .A(n11513), .Z(n11511) );
XOR U19187 ( .A(c3837), .B(b[3837]), .Z(n11512) );
XNOR U19188 ( .A(b[3837]), .B(n11513), .Z(c[3837]) );
XNOR U19189 ( .A(a[3837]), .B(c3837), .Z(n11513) );
XOR U19190 ( .A(c3838), .B(n11514), .Z(c3839) );
ANDN U19191 ( .B(n11515), .A(n11516), .Z(n11514) );
XOR U19192 ( .A(c3838), .B(b[3838]), .Z(n11515) );
XNOR U19193 ( .A(b[3838]), .B(n11516), .Z(c[3838]) );
XNOR U19194 ( .A(a[3838]), .B(c3838), .Z(n11516) );
XOR U19195 ( .A(c3839), .B(n11517), .Z(c3840) );
ANDN U19196 ( .B(n11518), .A(n11519), .Z(n11517) );
XOR U19197 ( .A(c3839), .B(b[3839]), .Z(n11518) );
XNOR U19198 ( .A(b[3839]), .B(n11519), .Z(c[3839]) );
XNOR U19199 ( .A(a[3839]), .B(c3839), .Z(n11519) );
XOR U19200 ( .A(c3840), .B(n11520), .Z(c3841) );
ANDN U19201 ( .B(n11521), .A(n11522), .Z(n11520) );
XOR U19202 ( .A(c3840), .B(b[3840]), .Z(n11521) );
XNOR U19203 ( .A(b[3840]), .B(n11522), .Z(c[3840]) );
XNOR U19204 ( .A(a[3840]), .B(c3840), .Z(n11522) );
XOR U19205 ( .A(c3841), .B(n11523), .Z(c3842) );
ANDN U19206 ( .B(n11524), .A(n11525), .Z(n11523) );
XOR U19207 ( .A(c3841), .B(b[3841]), .Z(n11524) );
XNOR U19208 ( .A(b[3841]), .B(n11525), .Z(c[3841]) );
XNOR U19209 ( .A(a[3841]), .B(c3841), .Z(n11525) );
XOR U19210 ( .A(c3842), .B(n11526), .Z(c3843) );
ANDN U19211 ( .B(n11527), .A(n11528), .Z(n11526) );
XOR U19212 ( .A(c3842), .B(b[3842]), .Z(n11527) );
XNOR U19213 ( .A(b[3842]), .B(n11528), .Z(c[3842]) );
XNOR U19214 ( .A(a[3842]), .B(c3842), .Z(n11528) );
XOR U19215 ( .A(c3843), .B(n11529), .Z(c3844) );
ANDN U19216 ( .B(n11530), .A(n11531), .Z(n11529) );
XOR U19217 ( .A(c3843), .B(b[3843]), .Z(n11530) );
XNOR U19218 ( .A(b[3843]), .B(n11531), .Z(c[3843]) );
XNOR U19219 ( .A(a[3843]), .B(c3843), .Z(n11531) );
XOR U19220 ( .A(c3844), .B(n11532), .Z(c3845) );
ANDN U19221 ( .B(n11533), .A(n11534), .Z(n11532) );
XOR U19222 ( .A(c3844), .B(b[3844]), .Z(n11533) );
XNOR U19223 ( .A(b[3844]), .B(n11534), .Z(c[3844]) );
XNOR U19224 ( .A(a[3844]), .B(c3844), .Z(n11534) );
XOR U19225 ( .A(c3845), .B(n11535), .Z(c3846) );
ANDN U19226 ( .B(n11536), .A(n11537), .Z(n11535) );
XOR U19227 ( .A(c3845), .B(b[3845]), .Z(n11536) );
XNOR U19228 ( .A(b[3845]), .B(n11537), .Z(c[3845]) );
XNOR U19229 ( .A(a[3845]), .B(c3845), .Z(n11537) );
XOR U19230 ( .A(c3846), .B(n11538), .Z(c3847) );
ANDN U19231 ( .B(n11539), .A(n11540), .Z(n11538) );
XOR U19232 ( .A(c3846), .B(b[3846]), .Z(n11539) );
XNOR U19233 ( .A(b[3846]), .B(n11540), .Z(c[3846]) );
XNOR U19234 ( .A(a[3846]), .B(c3846), .Z(n11540) );
XOR U19235 ( .A(c3847), .B(n11541), .Z(c3848) );
ANDN U19236 ( .B(n11542), .A(n11543), .Z(n11541) );
XOR U19237 ( .A(c3847), .B(b[3847]), .Z(n11542) );
XNOR U19238 ( .A(b[3847]), .B(n11543), .Z(c[3847]) );
XNOR U19239 ( .A(a[3847]), .B(c3847), .Z(n11543) );
XOR U19240 ( .A(c3848), .B(n11544), .Z(c3849) );
ANDN U19241 ( .B(n11545), .A(n11546), .Z(n11544) );
XOR U19242 ( .A(c3848), .B(b[3848]), .Z(n11545) );
XNOR U19243 ( .A(b[3848]), .B(n11546), .Z(c[3848]) );
XNOR U19244 ( .A(a[3848]), .B(c3848), .Z(n11546) );
XOR U19245 ( .A(c3849), .B(n11547), .Z(c3850) );
ANDN U19246 ( .B(n11548), .A(n11549), .Z(n11547) );
XOR U19247 ( .A(c3849), .B(b[3849]), .Z(n11548) );
XNOR U19248 ( .A(b[3849]), .B(n11549), .Z(c[3849]) );
XNOR U19249 ( .A(a[3849]), .B(c3849), .Z(n11549) );
XOR U19250 ( .A(c3850), .B(n11550), .Z(c3851) );
ANDN U19251 ( .B(n11551), .A(n11552), .Z(n11550) );
XOR U19252 ( .A(c3850), .B(b[3850]), .Z(n11551) );
XNOR U19253 ( .A(b[3850]), .B(n11552), .Z(c[3850]) );
XNOR U19254 ( .A(a[3850]), .B(c3850), .Z(n11552) );
XOR U19255 ( .A(c3851), .B(n11553), .Z(c3852) );
ANDN U19256 ( .B(n11554), .A(n11555), .Z(n11553) );
XOR U19257 ( .A(c3851), .B(b[3851]), .Z(n11554) );
XNOR U19258 ( .A(b[3851]), .B(n11555), .Z(c[3851]) );
XNOR U19259 ( .A(a[3851]), .B(c3851), .Z(n11555) );
XOR U19260 ( .A(c3852), .B(n11556), .Z(c3853) );
ANDN U19261 ( .B(n11557), .A(n11558), .Z(n11556) );
XOR U19262 ( .A(c3852), .B(b[3852]), .Z(n11557) );
XNOR U19263 ( .A(b[3852]), .B(n11558), .Z(c[3852]) );
XNOR U19264 ( .A(a[3852]), .B(c3852), .Z(n11558) );
XOR U19265 ( .A(c3853), .B(n11559), .Z(c3854) );
ANDN U19266 ( .B(n11560), .A(n11561), .Z(n11559) );
XOR U19267 ( .A(c3853), .B(b[3853]), .Z(n11560) );
XNOR U19268 ( .A(b[3853]), .B(n11561), .Z(c[3853]) );
XNOR U19269 ( .A(a[3853]), .B(c3853), .Z(n11561) );
XOR U19270 ( .A(c3854), .B(n11562), .Z(c3855) );
ANDN U19271 ( .B(n11563), .A(n11564), .Z(n11562) );
XOR U19272 ( .A(c3854), .B(b[3854]), .Z(n11563) );
XNOR U19273 ( .A(b[3854]), .B(n11564), .Z(c[3854]) );
XNOR U19274 ( .A(a[3854]), .B(c3854), .Z(n11564) );
XOR U19275 ( .A(c3855), .B(n11565), .Z(c3856) );
ANDN U19276 ( .B(n11566), .A(n11567), .Z(n11565) );
XOR U19277 ( .A(c3855), .B(b[3855]), .Z(n11566) );
XNOR U19278 ( .A(b[3855]), .B(n11567), .Z(c[3855]) );
XNOR U19279 ( .A(a[3855]), .B(c3855), .Z(n11567) );
XOR U19280 ( .A(c3856), .B(n11568), .Z(c3857) );
ANDN U19281 ( .B(n11569), .A(n11570), .Z(n11568) );
XOR U19282 ( .A(c3856), .B(b[3856]), .Z(n11569) );
XNOR U19283 ( .A(b[3856]), .B(n11570), .Z(c[3856]) );
XNOR U19284 ( .A(a[3856]), .B(c3856), .Z(n11570) );
XOR U19285 ( .A(c3857), .B(n11571), .Z(c3858) );
ANDN U19286 ( .B(n11572), .A(n11573), .Z(n11571) );
XOR U19287 ( .A(c3857), .B(b[3857]), .Z(n11572) );
XNOR U19288 ( .A(b[3857]), .B(n11573), .Z(c[3857]) );
XNOR U19289 ( .A(a[3857]), .B(c3857), .Z(n11573) );
XOR U19290 ( .A(c3858), .B(n11574), .Z(c3859) );
ANDN U19291 ( .B(n11575), .A(n11576), .Z(n11574) );
XOR U19292 ( .A(c3858), .B(b[3858]), .Z(n11575) );
XNOR U19293 ( .A(b[3858]), .B(n11576), .Z(c[3858]) );
XNOR U19294 ( .A(a[3858]), .B(c3858), .Z(n11576) );
XOR U19295 ( .A(c3859), .B(n11577), .Z(c3860) );
ANDN U19296 ( .B(n11578), .A(n11579), .Z(n11577) );
XOR U19297 ( .A(c3859), .B(b[3859]), .Z(n11578) );
XNOR U19298 ( .A(b[3859]), .B(n11579), .Z(c[3859]) );
XNOR U19299 ( .A(a[3859]), .B(c3859), .Z(n11579) );
XOR U19300 ( .A(c3860), .B(n11580), .Z(c3861) );
ANDN U19301 ( .B(n11581), .A(n11582), .Z(n11580) );
XOR U19302 ( .A(c3860), .B(b[3860]), .Z(n11581) );
XNOR U19303 ( .A(b[3860]), .B(n11582), .Z(c[3860]) );
XNOR U19304 ( .A(a[3860]), .B(c3860), .Z(n11582) );
XOR U19305 ( .A(c3861), .B(n11583), .Z(c3862) );
ANDN U19306 ( .B(n11584), .A(n11585), .Z(n11583) );
XOR U19307 ( .A(c3861), .B(b[3861]), .Z(n11584) );
XNOR U19308 ( .A(b[3861]), .B(n11585), .Z(c[3861]) );
XNOR U19309 ( .A(a[3861]), .B(c3861), .Z(n11585) );
XOR U19310 ( .A(c3862), .B(n11586), .Z(c3863) );
ANDN U19311 ( .B(n11587), .A(n11588), .Z(n11586) );
XOR U19312 ( .A(c3862), .B(b[3862]), .Z(n11587) );
XNOR U19313 ( .A(b[3862]), .B(n11588), .Z(c[3862]) );
XNOR U19314 ( .A(a[3862]), .B(c3862), .Z(n11588) );
XOR U19315 ( .A(c3863), .B(n11589), .Z(c3864) );
ANDN U19316 ( .B(n11590), .A(n11591), .Z(n11589) );
XOR U19317 ( .A(c3863), .B(b[3863]), .Z(n11590) );
XNOR U19318 ( .A(b[3863]), .B(n11591), .Z(c[3863]) );
XNOR U19319 ( .A(a[3863]), .B(c3863), .Z(n11591) );
XOR U19320 ( .A(c3864), .B(n11592), .Z(c3865) );
ANDN U19321 ( .B(n11593), .A(n11594), .Z(n11592) );
XOR U19322 ( .A(c3864), .B(b[3864]), .Z(n11593) );
XNOR U19323 ( .A(b[3864]), .B(n11594), .Z(c[3864]) );
XNOR U19324 ( .A(a[3864]), .B(c3864), .Z(n11594) );
XOR U19325 ( .A(c3865), .B(n11595), .Z(c3866) );
ANDN U19326 ( .B(n11596), .A(n11597), .Z(n11595) );
XOR U19327 ( .A(c3865), .B(b[3865]), .Z(n11596) );
XNOR U19328 ( .A(b[3865]), .B(n11597), .Z(c[3865]) );
XNOR U19329 ( .A(a[3865]), .B(c3865), .Z(n11597) );
XOR U19330 ( .A(c3866), .B(n11598), .Z(c3867) );
ANDN U19331 ( .B(n11599), .A(n11600), .Z(n11598) );
XOR U19332 ( .A(c3866), .B(b[3866]), .Z(n11599) );
XNOR U19333 ( .A(b[3866]), .B(n11600), .Z(c[3866]) );
XNOR U19334 ( .A(a[3866]), .B(c3866), .Z(n11600) );
XOR U19335 ( .A(c3867), .B(n11601), .Z(c3868) );
ANDN U19336 ( .B(n11602), .A(n11603), .Z(n11601) );
XOR U19337 ( .A(c3867), .B(b[3867]), .Z(n11602) );
XNOR U19338 ( .A(b[3867]), .B(n11603), .Z(c[3867]) );
XNOR U19339 ( .A(a[3867]), .B(c3867), .Z(n11603) );
XOR U19340 ( .A(c3868), .B(n11604), .Z(c3869) );
ANDN U19341 ( .B(n11605), .A(n11606), .Z(n11604) );
XOR U19342 ( .A(c3868), .B(b[3868]), .Z(n11605) );
XNOR U19343 ( .A(b[3868]), .B(n11606), .Z(c[3868]) );
XNOR U19344 ( .A(a[3868]), .B(c3868), .Z(n11606) );
XOR U19345 ( .A(c3869), .B(n11607), .Z(c3870) );
ANDN U19346 ( .B(n11608), .A(n11609), .Z(n11607) );
XOR U19347 ( .A(c3869), .B(b[3869]), .Z(n11608) );
XNOR U19348 ( .A(b[3869]), .B(n11609), .Z(c[3869]) );
XNOR U19349 ( .A(a[3869]), .B(c3869), .Z(n11609) );
XOR U19350 ( .A(c3870), .B(n11610), .Z(c3871) );
ANDN U19351 ( .B(n11611), .A(n11612), .Z(n11610) );
XOR U19352 ( .A(c3870), .B(b[3870]), .Z(n11611) );
XNOR U19353 ( .A(b[3870]), .B(n11612), .Z(c[3870]) );
XNOR U19354 ( .A(a[3870]), .B(c3870), .Z(n11612) );
XOR U19355 ( .A(c3871), .B(n11613), .Z(c3872) );
ANDN U19356 ( .B(n11614), .A(n11615), .Z(n11613) );
XOR U19357 ( .A(c3871), .B(b[3871]), .Z(n11614) );
XNOR U19358 ( .A(b[3871]), .B(n11615), .Z(c[3871]) );
XNOR U19359 ( .A(a[3871]), .B(c3871), .Z(n11615) );
XOR U19360 ( .A(c3872), .B(n11616), .Z(c3873) );
ANDN U19361 ( .B(n11617), .A(n11618), .Z(n11616) );
XOR U19362 ( .A(c3872), .B(b[3872]), .Z(n11617) );
XNOR U19363 ( .A(b[3872]), .B(n11618), .Z(c[3872]) );
XNOR U19364 ( .A(a[3872]), .B(c3872), .Z(n11618) );
XOR U19365 ( .A(c3873), .B(n11619), .Z(c3874) );
ANDN U19366 ( .B(n11620), .A(n11621), .Z(n11619) );
XOR U19367 ( .A(c3873), .B(b[3873]), .Z(n11620) );
XNOR U19368 ( .A(b[3873]), .B(n11621), .Z(c[3873]) );
XNOR U19369 ( .A(a[3873]), .B(c3873), .Z(n11621) );
XOR U19370 ( .A(c3874), .B(n11622), .Z(c3875) );
ANDN U19371 ( .B(n11623), .A(n11624), .Z(n11622) );
XOR U19372 ( .A(c3874), .B(b[3874]), .Z(n11623) );
XNOR U19373 ( .A(b[3874]), .B(n11624), .Z(c[3874]) );
XNOR U19374 ( .A(a[3874]), .B(c3874), .Z(n11624) );
XOR U19375 ( .A(c3875), .B(n11625), .Z(c3876) );
ANDN U19376 ( .B(n11626), .A(n11627), .Z(n11625) );
XOR U19377 ( .A(c3875), .B(b[3875]), .Z(n11626) );
XNOR U19378 ( .A(b[3875]), .B(n11627), .Z(c[3875]) );
XNOR U19379 ( .A(a[3875]), .B(c3875), .Z(n11627) );
XOR U19380 ( .A(c3876), .B(n11628), .Z(c3877) );
ANDN U19381 ( .B(n11629), .A(n11630), .Z(n11628) );
XOR U19382 ( .A(c3876), .B(b[3876]), .Z(n11629) );
XNOR U19383 ( .A(b[3876]), .B(n11630), .Z(c[3876]) );
XNOR U19384 ( .A(a[3876]), .B(c3876), .Z(n11630) );
XOR U19385 ( .A(c3877), .B(n11631), .Z(c3878) );
ANDN U19386 ( .B(n11632), .A(n11633), .Z(n11631) );
XOR U19387 ( .A(c3877), .B(b[3877]), .Z(n11632) );
XNOR U19388 ( .A(b[3877]), .B(n11633), .Z(c[3877]) );
XNOR U19389 ( .A(a[3877]), .B(c3877), .Z(n11633) );
XOR U19390 ( .A(c3878), .B(n11634), .Z(c3879) );
ANDN U19391 ( .B(n11635), .A(n11636), .Z(n11634) );
XOR U19392 ( .A(c3878), .B(b[3878]), .Z(n11635) );
XNOR U19393 ( .A(b[3878]), .B(n11636), .Z(c[3878]) );
XNOR U19394 ( .A(a[3878]), .B(c3878), .Z(n11636) );
XOR U19395 ( .A(c3879), .B(n11637), .Z(c3880) );
ANDN U19396 ( .B(n11638), .A(n11639), .Z(n11637) );
XOR U19397 ( .A(c3879), .B(b[3879]), .Z(n11638) );
XNOR U19398 ( .A(b[3879]), .B(n11639), .Z(c[3879]) );
XNOR U19399 ( .A(a[3879]), .B(c3879), .Z(n11639) );
XOR U19400 ( .A(c3880), .B(n11640), .Z(c3881) );
ANDN U19401 ( .B(n11641), .A(n11642), .Z(n11640) );
XOR U19402 ( .A(c3880), .B(b[3880]), .Z(n11641) );
XNOR U19403 ( .A(b[3880]), .B(n11642), .Z(c[3880]) );
XNOR U19404 ( .A(a[3880]), .B(c3880), .Z(n11642) );
XOR U19405 ( .A(c3881), .B(n11643), .Z(c3882) );
ANDN U19406 ( .B(n11644), .A(n11645), .Z(n11643) );
XOR U19407 ( .A(c3881), .B(b[3881]), .Z(n11644) );
XNOR U19408 ( .A(b[3881]), .B(n11645), .Z(c[3881]) );
XNOR U19409 ( .A(a[3881]), .B(c3881), .Z(n11645) );
XOR U19410 ( .A(c3882), .B(n11646), .Z(c3883) );
ANDN U19411 ( .B(n11647), .A(n11648), .Z(n11646) );
XOR U19412 ( .A(c3882), .B(b[3882]), .Z(n11647) );
XNOR U19413 ( .A(b[3882]), .B(n11648), .Z(c[3882]) );
XNOR U19414 ( .A(a[3882]), .B(c3882), .Z(n11648) );
XOR U19415 ( .A(c3883), .B(n11649), .Z(c3884) );
ANDN U19416 ( .B(n11650), .A(n11651), .Z(n11649) );
XOR U19417 ( .A(c3883), .B(b[3883]), .Z(n11650) );
XNOR U19418 ( .A(b[3883]), .B(n11651), .Z(c[3883]) );
XNOR U19419 ( .A(a[3883]), .B(c3883), .Z(n11651) );
XOR U19420 ( .A(c3884), .B(n11652), .Z(c3885) );
ANDN U19421 ( .B(n11653), .A(n11654), .Z(n11652) );
XOR U19422 ( .A(c3884), .B(b[3884]), .Z(n11653) );
XNOR U19423 ( .A(b[3884]), .B(n11654), .Z(c[3884]) );
XNOR U19424 ( .A(a[3884]), .B(c3884), .Z(n11654) );
XOR U19425 ( .A(c3885), .B(n11655), .Z(c3886) );
ANDN U19426 ( .B(n11656), .A(n11657), .Z(n11655) );
XOR U19427 ( .A(c3885), .B(b[3885]), .Z(n11656) );
XNOR U19428 ( .A(b[3885]), .B(n11657), .Z(c[3885]) );
XNOR U19429 ( .A(a[3885]), .B(c3885), .Z(n11657) );
XOR U19430 ( .A(c3886), .B(n11658), .Z(c3887) );
ANDN U19431 ( .B(n11659), .A(n11660), .Z(n11658) );
XOR U19432 ( .A(c3886), .B(b[3886]), .Z(n11659) );
XNOR U19433 ( .A(b[3886]), .B(n11660), .Z(c[3886]) );
XNOR U19434 ( .A(a[3886]), .B(c3886), .Z(n11660) );
XOR U19435 ( .A(c3887), .B(n11661), .Z(c3888) );
ANDN U19436 ( .B(n11662), .A(n11663), .Z(n11661) );
XOR U19437 ( .A(c3887), .B(b[3887]), .Z(n11662) );
XNOR U19438 ( .A(b[3887]), .B(n11663), .Z(c[3887]) );
XNOR U19439 ( .A(a[3887]), .B(c3887), .Z(n11663) );
XOR U19440 ( .A(c3888), .B(n11664), .Z(c3889) );
ANDN U19441 ( .B(n11665), .A(n11666), .Z(n11664) );
XOR U19442 ( .A(c3888), .B(b[3888]), .Z(n11665) );
XNOR U19443 ( .A(b[3888]), .B(n11666), .Z(c[3888]) );
XNOR U19444 ( .A(a[3888]), .B(c3888), .Z(n11666) );
XOR U19445 ( .A(c3889), .B(n11667), .Z(c3890) );
ANDN U19446 ( .B(n11668), .A(n11669), .Z(n11667) );
XOR U19447 ( .A(c3889), .B(b[3889]), .Z(n11668) );
XNOR U19448 ( .A(b[3889]), .B(n11669), .Z(c[3889]) );
XNOR U19449 ( .A(a[3889]), .B(c3889), .Z(n11669) );
XOR U19450 ( .A(c3890), .B(n11670), .Z(c3891) );
ANDN U19451 ( .B(n11671), .A(n11672), .Z(n11670) );
XOR U19452 ( .A(c3890), .B(b[3890]), .Z(n11671) );
XNOR U19453 ( .A(b[3890]), .B(n11672), .Z(c[3890]) );
XNOR U19454 ( .A(a[3890]), .B(c3890), .Z(n11672) );
XOR U19455 ( .A(c3891), .B(n11673), .Z(c3892) );
ANDN U19456 ( .B(n11674), .A(n11675), .Z(n11673) );
XOR U19457 ( .A(c3891), .B(b[3891]), .Z(n11674) );
XNOR U19458 ( .A(b[3891]), .B(n11675), .Z(c[3891]) );
XNOR U19459 ( .A(a[3891]), .B(c3891), .Z(n11675) );
XOR U19460 ( .A(c3892), .B(n11676), .Z(c3893) );
ANDN U19461 ( .B(n11677), .A(n11678), .Z(n11676) );
XOR U19462 ( .A(c3892), .B(b[3892]), .Z(n11677) );
XNOR U19463 ( .A(b[3892]), .B(n11678), .Z(c[3892]) );
XNOR U19464 ( .A(a[3892]), .B(c3892), .Z(n11678) );
XOR U19465 ( .A(c3893), .B(n11679), .Z(c3894) );
ANDN U19466 ( .B(n11680), .A(n11681), .Z(n11679) );
XOR U19467 ( .A(c3893), .B(b[3893]), .Z(n11680) );
XNOR U19468 ( .A(b[3893]), .B(n11681), .Z(c[3893]) );
XNOR U19469 ( .A(a[3893]), .B(c3893), .Z(n11681) );
XOR U19470 ( .A(c3894), .B(n11682), .Z(c3895) );
ANDN U19471 ( .B(n11683), .A(n11684), .Z(n11682) );
XOR U19472 ( .A(c3894), .B(b[3894]), .Z(n11683) );
XNOR U19473 ( .A(b[3894]), .B(n11684), .Z(c[3894]) );
XNOR U19474 ( .A(a[3894]), .B(c3894), .Z(n11684) );
XOR U19475 ( .A(c3895), .B(n11685), .Z(c3896) );
ANDN U19476 ( .B(n11686), .A(n11687), .Z(n11685) );
XOR U19477 ( .A(c3895), .B(b[3895]), .Z(n11686) );
XNOR U19478 ( .A(b[3895]), .B(n11687), .Z(c[3895]) );
XNOR U19479 ( .A(a[3895]), .B(c3895), .Z(n11687) );
XOR U19480 ( .A(c3896), .B(n11688), .Z(c3897) );
ANDN U19481 ( .B(n11689), .A(n11690), .Z(n11688) );
XOR U19482 ( .A(c3896), .B(b[3896]), .Z(n11689) );
XNOR U19483 ( .A(b[3896]), .B(n11690), .Z(c[3896]) );
XNOR U19484 ( .A(a[3896]), .B(c3896), .Z(n11690) );
XOR U19485 ( .A(c3897), .B(n11691), .Z(c3898) );
ANDN U19486 ( .B(n11692), .A(n11693), .Z(n11691) );
XOR U19487 ( .A(c3897), .B(b[3897]), .Z(n11692) );
XNOR U19488 ( .A(b[3897]), .B(n11693), .Z(c[3897]) );
XNOR U19489 ( .A(a[3897]), .B(c3897), .Z(n11693) );
XOR U19490 ( .A(c3898), .B(n11694), .Z(c3899) );
ANDN U19491 ( .B(n11695), .A(n11696), .Z(n11694) );
XOR U19492 ( .A(c3898), .B(b[3898]), .Z(n11695) );
XNOR U19493 ( .A(b[3898]), .B(n11696), .Z(c[3898]) );
XNOR U19494 ( .A(a[3898]), .B(c3898), .Z(n11696) );
XOR U19495 ( .A(c3899), .B(n11697), .Z(c3900) );
ANDN U19496 ( .B(n11698), .A(n11699), .Z(n11697) );
XOR U19497 ( .A(c3899), .B(b[3899]), .Z(n11698) );
XNOR U19498 ( .A(b[3899]), .B(n11699), .Z(c[3899]) );
XNOR U19499 ( .A(a[3899]), .B(c3899), .Z(n11699) );
XOR U19500 ( .A(c3900), .B(n11700), .Z(c3901) );
ANDN U19501 ( .B(n11701), .A(n11702), .Z(n11700) );
XOR U19502 ( .A(c3900), .B(b[3900]), .Z(n11701) );
XNOR U19503 ( .A(b[3900]), .B(n11702), .Z(c[3900]) );
XNOR U19504 ( .A(a[3900]), .B(c3900), .Z(n11702) );
XOR U19505 ( .A(c3901), .B(n11703), .Z(c3902) );
ANDN U19506 ( .B(n11704), .A(n11705), .Z(n11703) );
XOR U19507 ( .A(c3901), .B(b[3901]), .Z(n11704) );
XNOR U19508 ( .A(b[3901]), .B(n11705), .Z(c[3901]) );
XNOR U19509 ( .A(a[3901]), .B(c3901), .Z(n11705) );
XOR U19510 ( .A(c3902), .B(n11706), .Z(c3903) );
ANDN U19511 ( .B(n11707), .A(n11708), .Z(n11706) );
XOR U19512 ( .A(c3902), .B(b[3902]), .Z(n11707) );
XNOR U19513 ( .A(b[3902]), .B(n11708), .Z(c[3902]) );
XNOR U19514 ( .A(a[3902]), .B(c3902), .Z(n11708) );
XOR U19515 ( .A(c3903), .B(n11709), .Z(c3904) );
ANDN U19516 ( .B(n11710), .A(n11711), .Z(n11709) );
XOR U19517 ( .A(c3903), .B(b[3903]), .Z(n11710) );
XNOR U19518 ( .A(b[3903]), .B(n11711), .Z(c[3903]) );
XNOR U19519 ( .A(a[3903]), .B(c3903), .Z(n11711) );
XOR U19520 ( .A(c3904), .B(n11712), .Z(c3905) );
ANDN U19521 ( .B(n11713), .A(n11714), .Z(n11712) );
XOR U19522 ( .A(c3904), .B(b[3904]), .Z(n11713) );
XNOR U19523 ( .A(b[3904]), .B(n11714), .Z(c[3904]) );
XNOR U19524 ( .A(a[3904]), .B(c3904), .Z(n11714) );
XOR U19525 ( .A(c3905), .B(n11715), .Z(c3906) );
ANDN U19526 ( .B(n11716), .A(n11717), .Z(n11715) );
XOR U19527 ( .A(c3905), .B(b[3905]), .Z(n11716) );
XNOR U19528 ( .A(b[3905]), .B(n11717), .Z(c[3905]) );
XNOR U19529 ( .A(a[3905]), .B(c3905), .Z(n11717) );
XOR U19530 ( .A(c3906), .B(n11718), .Z(c3907) );
ANDN U19531 ( .B(n11719), .A(n11720), .Z(n11718) );
XOR U19532 ( .A(c3906), .B(b[3906]), .Z(n11719) );
XNOR U19533 ( .A(b[3906]), .B(n11720), .Z(c[3906]) );
XNOR U19534 ( .A(a[3906]), .B(c3906), .Z(n11720) );
XOR U19535 ( .A(c3907), .B(n11721), .Z(c3908) );
ANDN U19536 ( .B(n11722), .A(n11723), .Z(n11721) );
XOR U19537 ( .A(c3907), .B(b[3907]), .Z(n11722) );
XNOR U19538 ( .A(b[3907]), .B(n11723), .Z(c[3907]) );
XNOR U19539 ( .A(a[3907]), .B(c3907), .Z(n11723) );
XOR U19540 ( .A(c3908), .B(n11724), .Z(c3909) );
ANDN U19541 ( .B(n11725), .A(n11726), .Z(n11724) );
XOR U19542 ( .A(c3908), .B(b[3908]), .Z(n11725) );
XNOR U19543 ( .A(b[3908]), .B(n11726), .Z(c[3908]) );
XNOR U19544 ( .A(a[3908]), .B(c3908), .Z(n11726) );
XOR U19545 ( .A(c3909), .B(n11727), .Z(c3910) );
ANDN U19546 ( .B(n11728), .A(n11729), .Z(n11727) );
XOR U19547 ( .A(c3909), .B(b[3909]), .Z(n11728) );
XNOR U19548 ( .A(b[3909]), .B(n11729), .Z(c[3909]) );
XNOR U19549 ( .A(a[3909]), .B(c3909), .Z(n11729) );
XOR U19550 ( .A(c3910), .B(n11730), .Z(c3911) );
ANDN U19551 ( .B(n11731), .A(n11732), .Z(n11730) );
XOR U19552 ( .A(c3910), .B(b[3910]), .Z(n11731) );
XNOR U19553 ( .A(b[3910]), .B(n11732), .Z(c[3910]) );
XNOR U19554 ( .A(a[3910]), .B(c3910), .Z(n11732) );
XOR U19555 ( .A(c3911), .B(n11733), .Z(c3912) );
ANDN U19556 ( .B(n11734), .A(n11735), .Z(n11733) );
XOR U19557 ( .A(c3911), .B(b[3911]), .Z(n11734) );
XNOR U19558 ( .A(b[3911]), .B(n11735), .Z(c[3911]) );
XNOR U19559 ( .A(a[3911]), .B(c3911), .Z(n11735) );
XOR U19560 ( .A(c3912), .B(n11736), .Z(c3913) );
ANDN U19561 ( .B(n11737), .A(n11738), .Z(n11736) );
XOR U19562 ( .A(c3912), .B(b[3912]), .Z(n11737) );
XNOR U19563 ( .A(b[3912]), .B(n11738), .Z(c[3912]) );
XNOR U19564 ( .A(a[3912]), .B(c3912), .Z(n11738) );
XOR U19565 ( .A(c3913), .B(n11739), .Z(c3914) );
ANDN U19566 ( .B(n11740), .A(n11741), .Z(n11739) );
XOR U19567 ( .A(c3913), .B(b[3913]), .Z(n11740) );
XNOR U19568 ( .A(b[3913]), .B(n11741), .Z(c[3913]) );
XNOR U19569 ( .A(a[3913]), .B(c3913), .Z(n11741) );
XOR U19570 ( .A(c3914), .B(n11742), .Z(c3915) );
ANDN U19571 ( .B(n11743), .A(n11744), .Z(n11742) );
XOR U19572 ( .A(c3914), .B(b[3914]), .Z(n11743) );
XNOR U19573 ( .A(b[3914]), .B(n11744), .Z(c[3914]) );
XNOR U19574 ( .A(a[3914]), .B(c3914), .Z(n11744) );
XOR U19575 ( .A(c3915), .B(n11745), .Z(c3916) );
ANDN U19576 ( .B(n11746), .A(n11747), .Z(n11745) );
XOR U19577 ( .A(c3915), .B(b[3915]), .Z(n11746) );
XNOR U19578 ( .A(b[3915]), .B(n11747), .Z(c[3915]) );
XNOR U19579 ( .A(a[3915]), .B(c3915), .Z(n11747) );
XOR U19580 ( .A(c3916), .B(n11748), .Z(c3917) );
ANDN U19581 ( .B(n11749), .A(n11750), .Z(n11748) );
XOR U19582 ( .A(c3916), .B(b[3916]), .Z(n11749) );
XNOR U19583 ( .A(b[3916]), .B(n11750), .Z(c[3916]) );
XNOR U19584 ( .A(a[3916]), .B(c3916), .Z(n11750) );
XOR U19585 ( .A(c3917), .B(n11751), .Z(c3918) );
ANDN U19586 ( .B(n11752), .A(n11753), .Z(n11751) );
XOR U19587 ( .A(c3917), .B(b[3917]), .Z(n11752) );
XNOR U19588 ( .A(b[3917]), .B(n11753), .Z(c[3917]) );
XNOR U19589 ( .A(a[3917]), .B(c3917), .Z(n11753) );
XOR U19590 ( .A(c3918), .B(n11754), .Z(c3919) );
ANDN U19591 ( .B(n11755), .A(n11756), .Z(n11754) );
XOR U19592 ( .A(c3918), .B(b[3918]), .Z(n11755) );
XNOR U19593 ( .A(b[3918]), .B(n11756), .Z(c[3918]) );
XNOR U19594 ( .A(a[3918]), .B(c3918), .Z(n11756) );
XOR U19595 ( .A(c3919), .B(n11757), .Z(c3920) );
ANDN U19596 ( .B(n11758), .A(n11759), .Z(n11757) );
XOR U19597 ( .A(c3919), .B(b[3919]), .Z(n11758) );
XNOR U19598 ( .A(b[3919]), .B(n11759), .Z(c[3919]) );
XNOR U19599 ( .A(a[3919]), .B(c3919), .Z(n11759) );
XOR U19600 ( .A(c3920), .B(n11760), .Z(c3921) );
ANDN U19601 ( .B(n11761), .A(n11762), .Z(n11760) );
XOR U19602 ( .A(c3920), .B(b[3920]), .Z(n11761) );
XNOR U19603 ( .A(b[3920]), .B(n11762), .Z(c[3920]) );
XNOR U19604 ( .A(a[3920]), .B(c3920), .Z(n11762) );
XOR U19605 ( .A(c3921), .B(n11763), .Z(c3922) );
ANDN U19606 ( .B(n11764), .A(n11765), .Z(n11763) );
XOR U19607 ( .A(c3921), .B(b[3921]), .Z(n11764) );
XNOR U19608 ( .A(b[3921]), .B(n11765), .Z(c[3921]) );
XNOR U19609 ( .A(a[3921]), .B(c3921), .Z(n11765) );
XOR U19610 ( .A(c3922), .B(n11766), .Z(c3923) );
ANDN U19611 ( .B(n11767), .A(n11768), .Z(n11766) );
XOR U19612 ( .A(c3922), .B(b[3922]), .Z(n11767) );
XNOR U19613 ( .A(b[3922]), .B(n11768), .Z(c[3922]) );
XNOR U19614 ( .A(a[3922]), .B(c3922), .Z(n11768) );
XOR U19615 ( .A(c3923), .B(n11769), .Z(c3924) );
ANDN U19616 ( .B(n11770), .A(n11771), .Z(n11769) );
XOR U19617 ( .A(c3923), .B(b[3923]), .Z(n11770) );
XNOR U19618 ( .A(b[3923]), .B(n11771), .Z(c[3923]) );
XNOR U19619 ( .A(a[3923]), .B(c3923), .Z(n11771) );
XOR U19620 ( .A(c3924), .B(n11772), .Z(c3925) );
ANDN U19621 ( .B(n11773), .A(n11774), .Z(n11772) );
XOR U19622 ( .A(c3924), .B(b[3924]), .Z(n11773) );
XNOR U19623 ( .A(b[3924]), .B(n11774), .Z(c[3924]) );
XNOR U19624 ( .A(a[3924]), .B(c3924), .Z(n11774) );
XOR U19625 ( .A(c3925), .B(n11775), .Z(c3926) );
ANDN U19626 ( .B(n11776), .A(n11777), .Z(n11775) );
XOR U19627 ( .A(c3925), .B(b[3925]), .Z(n11776) );
XNOR U19628 ( .A(b[3925]), .B(n11777), .Z(c[3925]) );
XNOR U19629 ( .A(a[3925]), .B(c3925), .Z(n11777) );
XOR U19630 ( .A(c3926), .B(n11778), .Z(c3927) );
ANDN U19631 ( .B(n11779), .A(n11780), .Z(n11778) );
XOR U19632 ( .A(c3926), .B(b[3926]), .Z(n11779) );
XNOR U19633 ( .A(b[3926]), .B(n11780), .Z(c[3926]) );
XNOR U19634 ( .A(a[3926]), .B(c3926), .Z(n11780) );
XOR U19635 ( .A(c3927), .B(n11781), .Z(c3928) );
ANDN U19636 ( .B(n11782), .A(n11783), .Z(n11781) );
XOR U19637 ( .A(c3927), .B(b[3927]), .Z(n11782) );
XNOR U19638 ( .A(b[3927]), .B(n11783), .Z(c[3927]) );
XNOR U19639 ( .A(a[3927]), .B(c3927), .Z(n11783) );
XOR U19640 ( .A(c3928), .B(n11784), .Z(c3929) );
ANDN U19641 ( .B(n11785), .A(n11786), .Z(n11784) );
XOR U19642 ( .A(c3928), .B(b[3928]), .Z(n11785) );
XNOR U19643 ( .A(b[3928]), .B(n11786), .Z(c[3928]) );
XNOR U19644 ( .A(a[3928]), .B(c3928), .Z(n11786) );
XOR U19645 ( .A(c3929), .B(n11787), .Z(c3930) );
ANDN U19646 ( .B(n11788), .A(n11789), .Z(n11787) );
XOR U19647 ( .A(c3929), .B(b[3929]), .Z(n11788) );
XNOR U19648 ( .A(b[3929]), .B(n11789), .Z(c[3929]) );
XNOR U19649 ( .A(a[3929]), .B(c3929), .Z(n11789) );
XOR U19650 ( .A(c3930), .B(n11790), .Z(c3931) );
ANDN U19651 ( .B(n11791), .A(n11792), .Z(n11790) );
XOR U19652 ( .A(c3930), .B(b[3930]), .Z(n11791) );
XNOR U19653 ( .A(b[3930]), .B(n11792), .Z(c[3930]) );
XNOR U19654 ( .A(a[3930]), .B(c3930), .Z(n11792) );
XOR U19655 ( .A(c3931), .B(n11793), .Z(c3932) );
ANDN U19656 ( .B(n11794), .A(n11795), .Z(n11793) );
XOR U19657 ( .A(c3931), .B(b[3931]), .Z(n11794) );
XNOR U19658 ( .A(b[3931]), .B(n11795), .Z(c[3931]) );
XNOR U19659 ( .A(a[3931]), .B(c3931), .Z(n11795) );
XOR U19660 ( .A(c3932), .B(n11796), .Z(c3933) );
ANDN U19661 ( .B(n11797), .A(n11798), .Z(n11796) );
XOR U19662 ( .A(c3932), .B(b[3932]), .Z(n11797) );
XNOR U19663 ( .A(b[3932]), .B(n11798), .Z(c[3932]) );
XNOR U19664 ( .A(a[3932]), .B(c3932), .Z(n11798) );
XOR U19665 ( .A(c3933), .B(n11799), .Z(c3934) );
ANDN U19666 ( .B(n11800), .A(n11801), .Z(n11799) );
XOR U19667 ( .A(c3933), .B(b[3933]), .Z(n11800) );
XNOR U19668 ( .A(b[3933]), .B(n11801), .Z(c[3933]) );
XNOR U19669 ( .A(a[3933]), .B(c3933), .Z(n11801) );
XOR U19670 ( .A(c3934), .B(n11802), .Z(c3935) );
ANDN U19671 ( .B(n11803), .A(n11804), .Z(n11802) );
XOR U19672 ( .A(c3934), .B(b[3934]), .Z(n11803) );
XNOR U19673 ( .A(b[3934]), .B(n11804), .Z(c[3934]) );
XNOR U19674 ( .A(a[3934]), .B(c3934), .Z(n11804) );
XOR U19675 ( .A(c3935), .B(n11805), .Z(c3936) );
ANDN U19676 ( .B(n11806), .A(n11807), .Z(n11805) );
XOR U19677 ( .A(c3935), .B(b[3935]), .Z(n11806) );
XNOR U19678 ( .A(b[3935]), .B(n11807), .Z(c[3935]) );
XNOR U19679 ( .A(a[3935]), .B(c3935), .Z(n11807) );
XOR U19680 ( .A(c3936), .B(n11808), .Z(c3937) );
ANDN U19681 ( .B(n11809), .A(n11810), .Z(n11808) );
XOR U19682 ( .A(c3936), .B(b[3936]), .Z(n11809) );
XNOR U19683 ( .A(b[3936]), .B(n11810), .Z(c[3936]) );
XNOR U19684 ( .A(a[3936]), .B(c3936), .Z(n11810) );
XOR U19685 ( .A(c3937), .B(n11811), .Z(c3938) );
ANDN U19686 ( .B(n11812), .A(n11813), .Z(n11811) );
XOR U19687 ( .A(c3937), .B(b[3937]), .Z(n11812) );
XNOR U19688 ( .A(b[3937]), .B(n11813), .Z(c[3937]) );
XNOR U19689 ( .A(a[3937]), .B(c3937), .Z(n11813) );
XOR U19690 ( .A(c3938), .B(n11814), .Z(c3939) );
ANDN U19691 ( .B(n11815), .A(n11816), .Z(n11814) );
XOR U19692 ( .A(c3938), .B(b[3938]), .Z(n11815) );
XNOR U19693 ( .A(b[3938]), .B(n11816), .Z(c[3938]) );
XNOR U19694 ( .A(a[3938]), .B(c3938), .Z(n11816) );
XOR U19695 ( .A(c3939), .B(n11817), .Z(c3940) );
ANDN U19696 ( .B(n11818), .A(n11819), .Z(n11817) );
XOR U19697 ( .A(c3939), .B(b[3939]), .Z(n11818) );
XNOR U19698 ( .A(b[3939]), .B(n11819), .Z(c[3939]) );
XNOR U19699 ( .A(a[3939]), .B(c3939), .Z(n11819) );
XOR U19700 ( .A(c3940), .B(n11820), .Z(c3941) );
ANDN U19701 ( .B(n11821), .A(n11822), .Z(n11820) );
XOR U19702 ( .A(c3940), .B(b[3940]), .Z(n11821) );
XNOR U19703 ( .A(b[3940]), .B(n11822), .Z(c[3940]) );
XNOR U19704 ( .A(a[3940]), .B(c3940), .Z(n11822) );
XOR U19705 ( .A(c3941), .B(n11823), .Z(c3942) );
ANDN U19706 ( .B(n11824), .A(n11825), .Z(n11823) );
XOR U19707 ( .A(c3941), .B(b[3941]), .Z(n11824) );
XNOR U19708 ( .A(b[3941]), .B(n11825), .Z(c[3941]) );
XNOR U19709 ( .A(a[3941]), .B(c3941), .Z(n11825) );
XOR U19710 ( .A(c3942), .B(n11826), .Z(c3943) );
ANDN U19711 ( .B(n11827), .A(n11828), .Z(n11826) );
XOR U19712 ( .A(c3942), .B(b[3942]), .Z(n11827) );
XNOR U19713 ( .A(b[3942]), .B(n11828), .Z(c[3942]) );
XNOR U19714 ( .A(a[3942]), .B(c3942), .Z(n11828) );
XOR U19715 ( .A(c3943), .B(n11829), .Z(c3944) );
ANDN U19716 ( .B(n11830), .A(n11831), .Z(n11829) );
XOR U19717 ( .A(c3943), .B(b[3943]), .Z(n11830) );
XNOR U19718 ( .A(b[3943]), .B(n11831), .Z(c[3943]) );
XNOR U19719 ( .A(a[3943]), .B(c3943), .Z(n11831) );
XOR U19720 ( .A(c3944), .B(n11832), .Z(c3945) );
ANDN U19721 ( .B(n11833), .A(n11834), .Z(n11832) );
XOR U19722 ( .A(c3944), .B(b[3944]), .Z(n11833) );
XNOR U19723 ( .A(b[3944]), .B(n11834), .Z(c[3944]) );
XNOR U19724 ( .A(a[3944]), .B(c3944), .Z(n11834) );
XOR U19725 ( .A(c3945), .B(n11835), .Z(c3946) );
ANDN U19726 ( .B(n11836), .A(n11837), .Z(n11835) );
XOR U19727 ( .A(c3945), .B(b[3945]), .Z(n11836) );
XNOR U19728 ( .A(b[3945]), .B(n11837), .Z(c[3945]) );
XNOR U19729 ( .A(a[3945]), .B(c3945), .Z(n11837) );
XOR U19730 ( .A(c3946), .B(n11838), .Z(c3947) );
ANDN U19731 ( .B(n11839), .A(n11840), .Z(n11838) );
XOR U19732 ( .A(c3946), .B(b[3946]), .Z(n11839) );
XNOR U19733 ( .A(b[3946]), .B(n11840), .Z(c[3946]) );
XNOR U19734 ( .A(a[3946]), .B(c3946), .Z(n11840) );
XOR U19735 ( .A(c3947), .B(n11841), .Z(c3948) );
ANDN U19736 ( .B(n11842), .A(n11843), .Z(n11841) );
XOR U19737 ( .A(c3947), .B(b[3947]), .Z(n11842) );
XNOR U19738 ( .A(b[3947]), .B(n11843), .Z(c[3947]) );
XNOR U19739 ( .A(a[3947]), .B(c3947), .Z(n11843) );
XOR U19740 ( .A(c3948), .B(n11844), .Z(c3949) );
ANDN U19741 ( .B(n11845), .A(n11846), .Z(n11844) );
XOR U19742 ( .A(c3948), .B(b[3948]), .Z(n11845) );
XNOR U19743 ( .A(b[3948]), .B(n11846), .Z(c[3948]) );
XNOR U19744 ( .A(a[3948]), .B(c3948), .Z(n11846) );
XOR U19745 ( .A(c3949), .B(n11847), .Z(c3950) );
ANDN U19746 ( .B(n11848), .A(n11849), .Z(n11847) );
XOR U19747 ( .A(c3949), .B(b[3949]), .Z(n11848) );
XNOR U19748 ( .A(b[3949]), .B(n11849), .Z(c[3949]) );
XNOR U19749 ( .A(a[3949]), .B(c3949), .Z(n11849) );
XOR U19750 ( .A(c3950), .B(n11850), .Z(c3951) );
ANDN U19751 ( .B(n11851), .A(n11852), .Z(n11850) );
XOR U19752 ( .A(c3950), .B(b[3950]), .Z(n11851) );
XNOR U19753 ( .A(b[3950]), .B(n11852), .Z(c[3950]) );
XNOR U19754 ( .A(a[3950]), .B(c3950), .Z(n11852) );
XOR U19755 ( .A(c3951), .B(n11853), .Z(c3952) );
ANDN U19756 ( .B(n11854), .A(n11855), .Z(n11853) );
XOR U19757 ( .A(c3951), .B(b[3951]), .Z(n11854) );
XNOR U19758 ( .A(b[3951]), .B(n11855), .Z(c[3951]) );
XNOR U19759 ( .A(a[3951]), .B(c3951), .Z(n11855) );
XOR U19760 ( .A(c3952), .B(n11856), .Z(c3953) );
ANDN U19761 ( .B(n11857), .A(n11858), .Z(n11856) );
XOR U19762 ( .A(c3952), .B(b[3952]), .Z(n11857) );
XNOR U19763 ( .A(b[3952]), .B(n11858), .Z(c[3952]) );
XNOR U19764 ( .A(a[3952]), .B(c3952), .Z(n11858) );
XOR U19765 ( .A(c3953), .B(n11859), .Z(c3954) );
ANDN U19766 ( .B(n11860), .A(n11861), .Z(n11859) );
XOR U19767 ( .A(c3953), .B(b[3953]), .Z(n11860) );
XNOR U19768 ( .A(b[3953]), .B(n11861), .Z(c[3953]) );
XNOR U19769 ( .A(a[3953]), .B(c3953), .Z(n11861) );
XOR U19770 ( .A(c3954), .B(n11862), .Z(c3955) );
ANDN U19771 ( .B(n11863), .A(n11864), .Z(n11862) );
XOR U19772 ( .A(c3954), .B(b[3954]), .Z(n11863) );
XNOR U19773 ( .A(b[3954]), .B(n11864), .Z(c[3954]) );
XNOR U19774 ( .A(a[3954]), .B(c3954), .Z(n11864) );
XOR U19775 ( .A(c3955), .B(n11865), .Z(c3956) );
ANDN U19776 ( .B(n11866), .A(n11867), .Z(n11865) );
XOR U19777 ( .A(c3955), .B(b[3955]), .Z(n11866) );
XNOR U19778 ( .A(b[3955]), .B(n11867), .Z(c[3955]) );
XNOR U19779 ( .A(a[3955]), .B(c3955), .Z(n11867) );
XOR U19780 ( .A(c3956), .B(n11868), .Z(c3957) );
ANDN U19781 ( .B(n11869), .A(n11870), .Z(n11868) );
XOR U19782 ( .A(c3956), .B(b[3956]), .Z(n11869) );
XNOR U19783 ( .A(b[3956]), .B(n11870), .Z(c[3956]) );
XNOR U19784 ( .A(a[3956]), .B(c3956), .Z(n11870) );
XOR U19785 ( .A(c3957), .B(n11871), .Z(c3958) );
ANDN U19786 ( .B(n11872), .A(n11873), .Z(n11871) );
XOR U19787 ( .A(c3957), .B(b[3957]), .Z(n11872) );
XNOR U19788 ( .A(b[3957]), .B(n11873), .Z(c[3957]) );
XNOR U19789 ( .A(a[3957]), .B(c3957), .Z(n11873) );
XOR U19790 ( .A(c3958), .B(n11874), .Z(c3959) );
ANDN U19791 ( .B(n11875), .A(n11876), .Z(n11874) );
XOR U19792 ( .A(c3958), .B(b[3958]), .Z(n11875) );
XNOR U19793 ( .A(b[3958]), .B(n11876), .Z(c[3958]) );
XNOR U19794 ( .A(a[3958]), .B(c3958), .Z(n11876) );
XOR U19795 ( .A(c3959), .B(n11877), .Z(c3960) );
ANDN U19796 ( .B(n11878), .A(n11879), .Z(n11877) );
XOR U19797 ( .A(c3959), .B(b[3959]), .Z(n11878) );
XNOR U19798 ( .A(b[3959]), .B(n11879), .Z(c[3959]) );
XNOR U19799 ( .A(a[3959]), .B(c3959), .Z(n11879) );
XOR U19800 ( .A(c3960), .B(n11880), .Z(c3961) );
ANDN U19801 ( .B(n11881), .A(n11882), .Z(n11880) );
XOR U19802 ( .A(c3960), .B(b[3960]), .Z(n11881) );
XNOR U19803 ( .A(b[3960]), .B(n11882), .Z(c[3960]) );
XNOR U19804 ( .A(a[3960]), .B(c3960), .Z(n11882) );
XOR U19805 ( .A(c3961), .B(n11883), .Z(c3962) );
ANDN U19806 ( .B(n11884), .A(n11885), .Z(n11883) );
XOR U19807 ( .A(c3961), .B(b[3961]), .Z(n11884) );
XNOR U19808 ( .A(b[3961]), .B(n11885), .Z(c[3961]) );
XNOR U19809 ( .A(a[3961]), .B(c3961), .Z(n11885) );
XOR U19810 ( .A(c3962), .B(n11886), .Z(c3963) );
ANDN U19811 ( .B(n11887), .A(n11888), .Z(n11886) );
XOR U19812 ( .A(c3962), .B(b[3962]), .Z(n11887) );
XNOR U19813 ( .A(b[3962]), .B(n11888), .Z(c[3962]) );
XNOR U19814 ( .A(a[3962]), .B(c3962), .Z(n11888) );
XOR U19815 ( .A(c3963), .B(n11889), .Z(c3964) );
ANDN U19816 ( .B(n11890), .A(n11891), .Z(n11889) );
XOR U19817 ( .A(c3963), .B(b[3963]), .Z(n11890) );
XNOR U19818 ( .A(b[3963]), .B(n11891), .Z(c[3963]) );
XNOR U19819 ( .A(a[3963]), .B(c3963), .Z(n11891) );
XOR U19820 ( .A(c3964), .B(n11892), .Z(c3965) );
ANDN U19821 ( .B(n11893), .A(n11894), .Z(n11892) );
XOR U19822 ( .A(c3964), .B(b[3964]), .Z(n11893) );
XNOR U19823 ( .A(b[3964]), .B(n11894), .Z(c[3964]) );
XNOR U19824 ( .A(a[3964]), .B(c3964), .Z(n11894) );
XOR U19825 ( .A(c3965), .B(n11895), .Z(c3966) );
ANDN U19826 ( .B(n11896), .A(n11897), .Z(n11895) );
XOR U19827 ( .A(c3965), .B(b[3965]), .Z(n11896) );
XNOR U19828 ( .A(b[3965]), .B(n11897), .Z(c[3965]) );
XNOR U19829 ( .A(a[3965]), .B(c3965), .Z(n11897) );
XOR U19830 ( .A(c3966), .B(n11898), .Z(c3967) );
ANDN U19831 ( .B(n11899), .A(n11900), .Z(n11898) );
XOR U19832 ( .A(c3966), .B(b[3966]), .Z(n11899) );
XNOR U19833 ( .A(b[3966]), .B(n11900), .Z(c[3966]) );
XNOR U19834 ( .A(a[3966]), .B(c3966), .Z(n11900) );
XOR U19835 ( .A(c3967), .B(n11901), .Z(c3968) );
ANDN U19836 ( .B(n11902), .A(n11903), .Z(n11901) );
XOR U19837 ( .A(c3967), .B(b[3967]), .Z(n11902) );
XNOR U19838 ( .A(b[3967]), .B(n11903), .Z(c[3967]) );
XNOR U19839 ( .A(a[3967]), .B(c3967), .Z(n11903) );
XOR U19840 ( .A(c3968), .B(n11904), .Z(c3969) );
ANDN U19841 ( .B(n11905), .A(n11906), .Z(n11904) );
XOR U19842 ( .A(c3968), .B(b[3968]), .Z(n11905) );
XNOR U19843 ( .A(b[3968]), .B(n11906), .Z(c[3968]) );
XNOR U19844 ( .A(a[3968]), .B(c3968), .Z(n11906) );
XOR U19845 ( .A(c3969), .B(n11907), .Z(c3970) );
ANDN U19846 ( .B(n11908), .A(n11909), .Z(n11907) );
XOR U19847 ( .A(c3969), .B(b[3969]), .Z(n11908) );
XNOR U19848 ( .A(b[3969]), .B(n11909), .Z(c[3969]) );
XNOR U19849 ( .A(a[3969]), .B(c3969), .Z(n11909) );
XOR U19850 ( .A(c3970), .B(n11910), .Z(c3971) );
ANDN U19851 ( .B(n11911), .A(n11912), .Z(n11910) );
XOR U19852 ( .A(c3970), .B(b[3970]), .Z(n11911) );
XNOR U19853 ( .A(b[3970]), .B(n11912), .Z(c[3970]) );
XNOR U19854 ( .A(a[3970]), .B(c3970), .Z(n11912) );
XOR U19855 ( .A(c3971), .B(n11913), .Z(c3972) );
ANDN U19856 ( .B(n11914), .A(n11915), .Z(n11913) );
XOR U19857 ( .A(c3971), .B(b[3971]), .Z(n11914) );
XNOR U19858 ( .A(b[3971]), .B(n11915), .Z(c[3971]) );
XNOR U19859 ( .A(a[3971]), .B(c3971), .Z(n11915) );
XOR U19860 ( .A(c3972), .B(n11916), .Z(c3973) );
ANDN U19861 ( .B(n11917), .A(n11918), .Z(n11916) );
XOR U19862 ( .A(c3972), .B(b[3972]), .Z(n11917) );
XNOR U19863 ( .A(b[3972]), .B(n11918), .Z(c[3972]) );
XNOR U19864 ( .A(a[3972]), .B(c3972), .Z(n11918) );
XOR U19865 ( .A(c3973), .B(n11919), .Z(c3974) );
ANDN U19866 ( .B(n11920), .A(n11921), .Z(n11919) );
XOR U19867 ( .A(c3973), .B(b[3973]), .Z(n11920) );
XNOR U19868 ( .A(b[3973]), .B(n11921), .Z(c[3973]) );
XNOR U19869 ( .A(a[3973]), .B(c3973), .Z(n11921) );
XOR U19870 ( .A(c3974), .B(n11922), .Z(c3975) );
ANDN U19871 ( .B(n11923), .A(n11924), .Z(n11922) );
XOR U19872 ( .A(c3974), .B(b[3974]), .Z(n11923) );
XNOR U19873 ( .A(b[3974]), .B(n11924), .Z(c[3974]) );
XNOR U19874 ( .A(a[3974]), .B(c3974), .Z(n11924) );
XOR U19875 ( .A(c3975), .B(n11925), .Z(c3976) );
ANDN U19876 ( .B(n11926), .A(n11927), .Z(n11925) );
XOR U19877 ( .A(c3975), .B(b[3975]), .Z(n11926) );
XNOR U19878 ( .A(b[3975]), .B(n11927), .Z(c[3975]) );
XNOR U19879 ( .A(a[3975]), .B(c3975), .Z(n11927) );
XOR U19880 ( .A(c3976), .B(n11928), .Z(c3977) );
ANDN U19881 ( .B(n11929), .A(n11930), .Z(n11928) );
XOR U19882 ( .A(c3976), .B(b[3976]), .Z(n11929) );
XNOR U19883 ( .A(b[3976]), .B(n11930), .Z(c[3976]) );
XNOR U19884 ( .A(a[3976]), .B(c3976), .Z(n11930) );
XOR U19885 ( .A(c3977), .B(n11931), .Z(c3978) );
ANDN U19886 ( .B(n11932), .A(n11933), .Z(n11931) );
XOR U19887 ( .A(c3977), .B(b[3977]), .Z(n11932) );
XNOR U19888 ( .A(b[3977]), .B(n11933), .Z(c[3977]) );
XNOR U19889 ( .A(a[3977]), .B(c3977), .Z(n11933) );
XOR U19890 ( .A(c3978), .B(n11934), .Z(c3979) );
ANDN U19891 ( .B(n11935), .A(n11936), .Z(n11934) );
XOR U19892 ( .A(c3978), .B(b[3978]), .Z(n11935) );
XNOR U19893 ( .A(b[3978]), .B(n11936), .Z(c[3978]) );
XNOR U19894 ( .A(a[3978]), .B(c3978), .Z(n11936) );
XOR U19895 ( .A(c3979), .B(n11937), .Z(c3980) );
ANDN U19896 ( .B(n11938), .A(n11939), .Z(n11937) );
XOR U19897 ( .A(c3979), .B(b[3979]), .Z(n11938) );
XNOR U19898 ( .A(b[3979]), .B(n11939), .Z(c[3979]) );
XNOR U19899 ( .A(a[3979]), .B(c3979), .Z(n11939) );
XOR U19900 ( .A(c3980), .B(n11940), .Z(c3981) );
ANDN U19901 ( .B(n11941), .A(n11942), .Z(n11940) );
XOR U19902 ( .A(c3980), .B(b[3980]), .Z(n11941) );
XNOR U19903 ( .A(b[3980]), .B(n11942), .Z(c[3980]) );
XNOR U19904 ( .A(a[3980]), .B(c3980), .Z(n11942) );
XOR U19905 ( .A(c3981), .B(n11943), .Z(c3982) );
ANDN U19906 ( .B(n11944), .A(n11945), .Z(n11943) );
XOR U19907 ( .A(c3981), .B(b[3981]), .Z(n11944) );
XNOR U19908 ( .A(b[3981]), .B(n11945), .Z(c[3981]) );
XNOR U19909 ( .A(a[3981]), .B(c3981), .Z(n11945) );
XOR U19910 ( .A(c3982), .B(n11946), .Z(c3983) );
ANDN U19911 ( .B(n11947), .A(n11948), .Z(n11946) );
XOR U19912 ( .A(c3982), .B(b[3982]), .Z(n11947) );
XNOR U19913 ( .A(b[3982]), .B(n11948), .Z(c[3982]) );
XNOR U19914 ( .A(a[3982]), .B(c3982), .Z(n11948) );
XOR U19915 ( .A(c3983), .B(n11949), .Z(c3984) );
ANDN U19916 ( .B(n11950), .A(n11951), .Z(n11949) );
XOR U19917 ( .A(c3983), .B(b[3983]), .Z(n11950) );
XNOR U19918 ( .A(b[3983]), .B(n11951), .Z(c[3983]) );
XNOR U19919 ( .A(a[3983]), .B(c3983), .Z(n11951) );
XOR U19920 ( .A(c3984), .B(n11952), .Z(c3985) );
ANDN U19921 ( .B(n11953), .A(n11954), .Z(n11952) );
XOR U19922 ( .A(c3984), .B(b[3984]), .Z(n11953) );
XNOR U19923 ( .A(b[3984]), .B(n11954), .Z(c[3984]) );
XNOR U19924 ( .A(a[3984]), .B(c3984), .Z(n11954) );
XOR U19925 ( .A(c3985), .B(n11955), .Z(c3986) );
ANDN U19926 ( .B(n11956), .A(n11957), .Z(n11955) );
XOR U19927 ( .A(c3985), .B(b[3985]), .Z(n11956) );
XNOR U19928 ( .A(b[3985]), .B(n11957), .Z(c[3985]) );
XNOR U19929 ( .A(a[3985]), .B(c3985), .Z(n11957) );
XOR U19930 ( .A(c3986), .B(n11958), .Z(c3987) );
ANDN U19931 ( .B(n11959), .A(n11960), .Z(n11958) );
XOR U19932 ( .A(c3986), .B(b[3986]), .Z(n11959) );
XNOR U19933 ( .A(b[3986]), .B(n11960), .Z(c[3986]) );
XNOR U19934 ( .A(a[3986]), .B(c3986), .Z(n11960) );
XOR U19935 ( .A(c3987), .B(n11961), .Z(c3988) );
ANDN U19936 ( .B(n11962), .A(n11963), .Z(n11961) );
XOR U19937 ( .A(c3987), .B(b[3987]), .Z(n11962) );
XNOR U19938 ( .A(b[3987]), .B(n11963), .Z(c[3987]) );
XNOR U19939 ( .A(a[3987]), .B(c3987), .Z(n11963) );
XOR U19940 ( .A(c3988), .B(n11964), .Z(c3989) );
ANDN U19941 ( .B(n11965), .A(n11966), .Z(n11964) );
XOR U19942 ( .A(c3988), .B(b[3988]), .Z(n11965) );
XNOR U19943 ( .A(b[3988]), .B(n11966), .Z(c[3988]) );
XNOR U19944 ( .A(a[3988]), .B(c3988), .Z(n11966) );
XOR U19945 ( .A(c3989), .B(n11967), .Z(c3990) );
ANDN U19946 ( .B(n11968), .A(n11969), .Z(n11967) );
XOR U19947 ( .A(c3989), .B(b[3989]), .Z(n11968) );
XNOR U19948 ( .A(b[3989]), .B(n11969), .Z(c[3989]) );
XNOR U19949 ( .A(a[3989]), .B(c3989), .Z(n11969) );
XOR U19950 ( .A(c3990), .B(n11970), .Z(c3991) );
ANDN U19951 ( .B(n11971), .A(n11972), .Z(n11970) );
XOR U19952 ( .A(c3990), .B(b[3990]), .Z(n11971) );
XNOR U19953 ( .A(b[3990]), .B(n11972), .Z(c[3990]) );
XNOR U19954 ( .A(a[3990]), .B(c3990), .Z(n11972) );
XOR U19955 ( .A(c3991), .B(n11973), .Z(c3992) );
ANDN U19956 ( .B(n11974), .A(n11975), .Z(n11973) );
XOR U19957 ( .A(c3991), .B(b[3991]), .Z(n11974) );
XNOR U19958 ( .A(b[3991]), .B(n11975), .Z(c[3991]) );
XNOR U19959 ( .A(a[3991]), .B(c3991), .Z(n11975) );
XOR U19960 ( .A(c3992), .B(n11976), .Z(c3993) );
ANDN U19961 ( .B(n11977), .A(n11978), .Z(n11976) );
XOR U19962 ( .A(c3992), .B(b[3992]), .Z(n11977) );
XNOR U19963 ( .A(b[3992]), .B(n11978), .Z(c[3992]) );
XNOR U19964 ( .A(a[3992]), .B(c3992), .Z(n11978) );
XOR U19965 ( .A(c3993), .B(n11979), .Z(c3994) );
ANDN U19966 ( .B(n11980), .A(n11981), .Z(n11979) );
XOR U19967 ( .A(c3993), .B(b[3993]), .Z(n11980) );
XNOR U19968 ( .A(b[3993]), .B(n11981), .Z(c[3993]) );
XNOR U19969 ( .A(a[3993]), .B(c3993), .Z(n11981) );
XOR U19970 ( .A(c3994), .B(n11982), .Z(c3995) );
ANDN U19971 ( .B(n11983), .A(n11984), .Z(n11982) );
XOR U19972 ( .A(c3994), .B(b[3994]), .Z(n11983) );
XNOR U19973 ( .A(b[3994]), .B(n11984), .Z(c[3994]) );
XNOR U19974 ( .A(a[3994]), .B(c3994), .Z(n11984) );
XOR U19975 ( .A(c3995), .B(n11985), .Z(c3996) );
ANDN U19976 ( .B(n11986), .A(n11987), .Z(n11985) );
XOR U19977 ( .A(c3995), .B(b[3995]), .Z(n11986) );
XNOR U19978 ( .A(b[3995]), .B(n11987), .Z(c[3995]) );
XNOR U19979 ( .A(a[3995]), .B(c3995), .Z(n11987) );
XOR U19980 ( .A(c3996), .B(n11988), .Z(c3997) );
ANDN U19981 ( .B(n11989), .A(n11990), .Z(n11988) );
XOR U19982 ( .A(c3996), .B(b[3996]), .Z(n11989) );
XNOR U19983 ( .A(b[3996]), .B(n11990), .Z(c[3996]) );
XNOR U19984 ( .A(a[3996]), .B(c3996), .Z(n11990) );
XOR U19985 ( .A(c3997), .B(n11991), .Z(c3998) );
ANDN U19986 ( .B(n11992), .A(n11993), .Z(n11991) );
XOR U19987 ( .A(c3997), .B(b[3997]), .Z(n11992) );
XNOR U19988 ( .A(b[3997]), .B(n11993), .Z(c[3997]) );
XNOR U19989 ( .A(a[3997]), .B(c3997), .Z(n11993) );
XOR U19990 ( .A(c3998), .B(n11994), .Z(c3999) );
ANDN U19991 ( .B(n11995), .A(n11996), .Z(n11994) );
XOR U19992 ( .A(c3998), .B(b[3998]), .Z(n11995) );
XNOR U19993 ( .A(b[3998]), .B(n11996), .Z(c[3998]) );
XNOR U19994 ( .A(a[3998]), .B(c3998), .Z(n11996) );
XOR U19995 ( .A(c3999), .B(n11997), .Z(c4000) );
ANDN U19996 ( .B(n11998), .A(n11999), .Z(n11997) );
XOR U19997 ( .A(c3999), .B(b[3999]), .Z(n11998) );
XNOR U19998 ( .A(b[3999]), .B(n11999), .Z(c[3999]) );
XNOR U19999 ( .A(a[3999]), .B(c3999), .Z(n11999) );
XOR U20000 ( .A(c4000), .B(n12000), .Z(c4001) );
ANDN U20001 ( .B(n12001), .A(n12002), .Z(n12000) );
XOR U20002 ( .A(c4000), .B(b[4000]), .Z(n12001) );
XNOR U20003 ( .A(b[4000]), .B(n12002), .Z(c[4000]) );
XNOR U20004 ( .A(a[4000]), .B(c4000), .Z(n12002) );
XOR U20005 ( .A(c4001), .B(n12003), .Z(c4002) );
ANDN U20006 ( .B(n12004), .A(n12005), .Z(n12003) );
XOR U20007 ( .A(c4001), .B(b[4001]), .Z(n12004) );
XNOR U20008 ( .A(b[4001]), .B(n12005), .Z(c[4001]) );
XNOR U20009 ( .A(a[4001]), .B(c4001), .Z(n12005) );
XOR U20010 ( .A(c4002), .B(n12006), .Z(c4003) );
ANDN U20011 ( .B(n12007), .A(n12008), .Z(n12006) );
XOR U20012 ( .A(c4002), .B(b[4002]), .Z(n12007) );
XNOR U20013 ( .A(b[4002]), .B(n12008), .Z(c[4002]) );
XNOR U20014 ( .A(a[4002]), .B(c4002), .Z(n12008) );
XOR U20015 ( .A(c4003), .B(n12009), .Z(c4004) );
ANDN U20016 ( .B(n12010), .A(n12011), .Z(n12009) );
XOR U20017 ( .A(c4003), .B(b[4003]), .Z(n12010) );
XNOR U20018 ( .A(b[4003]), .B(n12011), .Z(c[4003]) );
XNOR U20019 ( .A(a[4003]), .B(c4003), .Z(n12011) );
XOR U20020 ( .A(c4004), .B(n12012), .Z(c4005) );
ANDN U20021 ( .B(n12013), .A(n12014), .Z(n12012) );
XOR U20022 ( .A(c4004), .B(b[4004]), .Z(n12013) );
XNOR U20023 ( .A(b[4004]), .B(n12014), .Z(c[4004]) );
XNOR U20024 ( .A(a[4004]), .B(c4004), .Z(n12014) );
XOR U20025 ( .A(c4005), .B(n12015), .Z(c4006) );
ANDN U20026 ( .B(n12016), .A(n12017), .Z(n12015) );
XOR U20027 ( .A(c4005), .B(b[4005]), .Z(n12016) );
XNOR U20028 ( .A(b[4005]), .B(n12017), .Z(c[4005]) );
XNOR U20029 ( .A(a[4005]), .B(c4005), .Z(n12017) );
XOR U20030 ( .A(c4006), .B(n12018), .Z(c4007) );
ANDN U20031 ( .B(n12019), .A(n12020), .Z(n12018) );
XOR U20032 ( .A(c4006), .B(b[4006]), .Z(n12019) );
XNOR U20033 ( .A(b[4006]), .B(n12020), .Z(c[4006]) );
XNOR U20034 ( .A(a[4006]), .B(c4006), .Z(n12020) );
XOR U20035 ( .A(c4007), .B(n12021), .Z(c4008) );
ANDN U20036 ( .B(n12022), .A(n12023), .Z(n12021) );
XOR U20037 ( .A(c4007), .B(b[4007]), .Z(n12022) );
XNOR U20038 ( .A(b[4007]), .B(n12023), .Z(c[4007]) );
XNOR U20039 ( .A(a[4007]), .B(c4007), .Z(n12023) );
XOR U20040 ( .A(c4008), .B(n12024), .Z(c4009) );
ANDN U20041 ( .B(n12025), .A(n12026), .Z(n12024) );
XOR U20042 ( .A(c4008), .B(b[4008]), .Z(n12025) );
XNOR U20043 ( .A(b[4008]), .B(n12026), .Z(c[4008]) );
XNOR U20044 ( .A(a[4008]), .B(c4008), .Z(n12026) );
XOR U20045 ( .A(c4009), .B(n12027), .Z(c4010) );
ANDN U20046 ( .B(n12028), .A(n12029), .Z(n12027) );
XOR U20047 ( .A(c4009), .B(b[4009]), .Z(n12028) );
XNOR U20048 ( .A(b[4009]), .B(n12029), .Z(c[4009]) );
XNOR U20049 ( .A(a[4009]), .B(c4009), .Z(n12029) );
XOR U20050 ( .A(c4010), .B(n12030), .Z(c4011) );
ANDN U20051 ( .B(n12031), .A(n12032), .Z(n12030) );
XOR U20052 ( .A(c4010), .B(b[4010]), .Z(n12031) );
XNOR U20053 ( .A(b[4010]), .B(n12032), .Z(c[4010]) );
XNOR U20054 ( .A(a[4010]), .B(c4010), .Z(n12032) );
XOR U20055 ( .A(c4011), .B(n12033), .Z(c4012) );
ANDN U20056 ( .B(n12034), .A(n12035), .Z(n12033) );
XOR U20057 ( .A(c4011), .B(b[4011]), .Z(n12034) );
XNOR U20058 ( .A(b[4011]), .B(n12035), .Z(c[4011]) );
XNOR U20059 ( .A(a[4011]), .B(c4011), .Z(n12035) );
XOR U20060 ( .A(c4012), .B(n12036), .Z(c4013) );
ANDN U20061 ( .B(n12037), .A(n12038), .Z(n12036) );
XOR U20062 ( .A(c4012), .B(b[4012]), .Z(n12037) );
XNOR U20063 ( .A(b[4012]), .B(n12038), .Z(c[4012]) );
XNOR U20064 ( .A(a[4012]), .B(c4012), .Z(n12038) );
XOR U20065 ( .A(c4013), .B(n12039), .Z(c4014) );
ANDN U20066 ( .B(n12040), .A(n12041), .Z(n12039) );
XOR U20067 ( .A(c4013), .B(b[4013]), .Z(n12040) );
XNOR U20068 ( .A(b[4013]), .B(n12041), .Z(c[4013]) );
XNOR U20069 ( .A(a[4013]), .B(c4013), .Z(n12041) );
XOR U20070 ( .A(c4014), .B(n12042), .Z(c4015) );
ANDN U20071 ( .B(n12043), .A(n12044), .Z(n12042) );
XOR U20072 ( .A(c4014), .B(b[4014]), .Z(n12043) );
XNOR U20073 ( .A(b[4014]), .B(n12044), .Z(c[4014]) );
XNOR U20074 ( .A(a[4014]), .B(c4014), .Z(n12044) );
XOR U20075 ( .A(c4015), .B(n12045), .Z(c4016) );
ANDN U20076 ( .B(n12046), .A(n12047), .Z(n12045) );
XOR U20077 ( .A(c4015), .B(b[4015]), .Z(n12046) );
XNOR U20078 ( .A(b[4015]), .B(n12047), .Z(c[4015]) );
XNOR U20079 ( .A(a[4015]), .B(c4015), .Z(n12047) );
XOR U20080 ( .A(c4016), .B(n12048), .Z(c4017) );
ANDN U20081 ( .B(n12049), .A(n12050), .Z(n12048) );
XOR U20082 ( .A(c4016), .B(b[4016]), .Z(n12049) );
XNOR U20083 ( .A(b[4016]), .B(n12050), .Z(c[4016]) );
XNOR U20084 ( .A(a[4016]), .B(c4016), .Z(n12050) );
XOR U20085 ( .A(c4017), .B(n12051), .Z(c4018) );
ANDN U20086 ( .B(n12052), .A(n12053), .Z(n12051) );
XOR U20087 ( .A(c4017), .B(b[4017]), .Z(n12052) );
XNOR U20088 ( .A(b[4017]), .B(n12053), .Z(c[4017]) );
XNOR U20089 ( .A(a[4017]), .B(c4017), .Z(n12053) );
XOR U20090 ( .A(c4018), .B(n12054), .Z(c4019) );
ANDN U20091 ( .B(n12055), .A(n12056), .Z(n12054) );
XOR U20092 ( .A(c4018), .B(b[4018]), .Z(n12055) );
XNOR U20093 ( .A(b[4018]), .B(n12056), .Z(c[4018]) );
XNOR U20094 ( .A(a[4018]), .B(c4018), .Z(n12056) );
XOR U20095 ( .A(c4019), .B(n12057), .Z(c4020) );
ANDN U20096 ( .B(n12058), .A(n12059), .Z(n12057) );
XOR U20097 ( .A(c4019), .B(b[4019]), .Z(n12058) );
XNOR U20098 ( .A(b[4019]), .B(n12059), .Z(c[4019]) );
XNOR U20099 ( .A(a[4019]), .B(c4019), .Z(n12059) );
XOR U20100 ( .A(c4020), .B(n12060), .Z(c4021) );
ANDN U20101 ( .B(n12061), .A(n12062), .Z(n12060) );
XOR U20102 ( .A(c4020), .B(b[4020]), .Z(n12061) );
XNOR U20103 ( .A(b[4020]), .B(n12062), .Z(c[4020]) );
XNOR U20104 ( .A(a[4020]), .B(c4020), .Z(n12062) );
XOR U20105 ( .A(c4021), .B(n12063), .Z(c4022) );
ANDN U20106 ( .B(n12064), .A(n12065), .Z(n12063) );
XOR U20107 ( .A(c4021), .B(b[4021]), .Z(n12064) );
XNOR U20108 ( .A(b[4021]), .B(n12065), .Z(c[4021]) );
XNOR U20109 ( .A(a[4021]), .B(c4021), .Z(n12065) );
XOR U20110 ( .A(c4022), .B(n12066), .Z(c4023) );
ANDN U20111 ( .B(n12067), .A(n12068), .Z(n12066) );
XOR U20112 ( .A(c4022), .B(b[4022]), .Z(n12067) );
XNOR U20113 ( .A(b[4022]), .B(n12068), .Z(c[4022]) );
XNOR U20114 ( .A(a[4022]), .B(c4022), .Z(n12068) );
XOR U20115 ( .A(c4023), .B(n12069), .Z(c4024) );
ANDN U20116 ( .B(n12070), .A(n12071), .Z(n12069) );
XOR U20117 ( .A(c4023), .B(b[4023]), .Z(n12070) );
XNOR U20118 ( .A(b[4023]), .B(n12071), .Z(c[4023]) );
XNOR U20119 ( .A(a[4023]), .B(c4023), .Z(n12071) );
XOR U20120 ( .A(c4024), .B(n12072), .Z(c4025) );
ANDN U20121 ( .B(n12073), .A(n12074), .Z(n12072) );
XOR U20122 ( .A(c4024), .B(b[4024]), .Z(n12073) );
XNOR U20123 ( .A(b[4024]), .B(n12074), .Z(c[4024]) );
XNOR U20124 ( .A(a[4024]), .B(c4024), .Z(n12074) );
XOR U20125 ( .A(c4025), .B(n12075), .Z(c4026) );
ANDN U20126 ( .B(n12076), .A(n12077), .Z(n12075) );
XOR U20127 ( .A(c4025), .B(b[4025]), .Z(n12076) );
XNOR U20128 ( .A(b[4025]), .B(n12077), .Z(c[4025]) );
XNOR U20129 ( .A(a[4025]), .B(c4025), .Z(n12077) );
XOR U20130 ( .A(c4026), .B(n12078), .Z(c4027) );
ANDN U20131 ( .B(n12079), .A(n12080), .Z(n12078) );
XOR U20132 ( .A(c4026), .B(b[4026]), .Z(n12079) );
XNOR U20133 ( .A(b[4026]), .B(n12080), .Z(c[4026]) );
XNOR U20134 ( .A(a[4026]), .B(c4026), .Z(n12080) );
XOR U20135 ( .A(c4027), .B(n12081), .Z(c4028) );
ANDN U20136 ( .B(n12082), .A(n12083), .Z(n12081) );
XOR U20137 ( .A(c4027), .B(b[4027]), .Z(n12082) );
XNOR U20138 ( .A(b[4027]), .B(n12083), .Z(c[4027]) );
XNOR U20139 ( .A(a[4027]), .B(c4027), .Z(n12083) );
XOR U20140 ( .A(c4028), .B(n12084), .Z(c4029) );
ANDN U20141 ( .B(n12085), .A(n12086), .Z(n12084) );
XOR U20142 ( .A(c4028), .B(b[4028]), .Z(n12085) );
XNOR U20143 ( .A(b[4028]), .B(n12086), .Z(c[4028]) );
XNOR U20144 ( .A(a[4028]), .B(c4028), .Z(n12086) );
XOR U20145 ( .A(c4029), .B(n12087), .Z(c4030) );
ANDN U20146 ( .B(n12088), .A(n12089), .Z(n12087) );
XOR U20147 ( .A(c4029), .B(b[4029]), .Z(n12088) );
XNOR U20148 ( .A(b[4029]), .B(n12089), .Z(c[4029]) );
XNOR U20149 ( .A(a[4029]), .B(c4029), .Z(n12089) );
XOR U20150 ( .A(c4030), .B(n12090), .Z(c4031) );
ANDN U20151 ( .B(n12091), .A(n12092), .Z(n12090) );
XOR U20152 ( .A(c4030), .B(b[4030]), .Z(n12091) );
XNOR U20153 ( .A(b[4030]), .B(n12092), .Z(c[4030]) );
XNOR U20154 ( .A(a[4030]), .B(c4030), .Z(n12092) );
XOR U20155 ( .A(c4031), .B(n12093), .Z(c4032) );
ANDN U20156 ( .B(n12094), .A(n12095), .Z(n12093) );
XOR U20157 ( .A(c4031), .B(b[4031]), .Z(n12094) );
XNOR U20158 ( .A(b[4031]), .B(n12095), .Z(c[4031]) );
XNOR U20159 ( .A(a[4031]), .B(c4031), .Z(n12095) );
XOR U20160 ( .A(c4032), .B(n12096), .Z(c4033) );
ANDN U20161 ( .B(n12097), .A(n12098), .Z(n12096) );
XOR U20162 ( .A(c4032), .B(b[4032]), .Z(n12097) );
XNOR U20163 ( .A(b[4032]), .B(n12098), .Z(c[4032]) );
XNOR U20164 ( .A(a[4032]), .B(c4032), .Z(n12098) );
XOR U20165 ( .A(c4033), .B(n12099), .Z(c4034) );
ANDN U20166 ( .B(n12100), .A(n12101), .Z(n12099) );
XOR U20167 ( .A(c4033), .B(b[4033]), .Z(n12100) );
XNOR U20168 ( .A(b[4033]), .B(n12101), .Z(c[4033]) );
XNOR U20169 ( .A(a[4033]), .B(c4033), .Z(n12101) );
XOR U20170 ( .A(c4034), .B(n12102), .Z(c4035) );
ANDN U20171 ( .B(n12103), .A(n12104), .Z(n12102) );
XOR U20172 ( .A(c4034), .B(b[4034]), .Z(n12103) );
XNOR U20173 ( .A(b[4034]), .B(n12104), .Z(c[4034]) );
XNOR U20174 ( .A(a[4034]), .B(c4034), .Z(n12104) );
XOR U20175 ( .A(c4035), .B(n12105), .Z(c4036) );
ANDN U20176 ( .B(n12106), .A(n12107), .Z(n12105) );
XOR U20177 ( .A(c4035), .B(b[4035]), .Z(n12106) );
XNOR U20178 ( .A(b[4035]), .B(n12107), .Z(c[4035]) );
XNOR U20179 ( .A(a[4035]), .B(c4035), .Z(n12107) );
XOR U20180 ( .A(c4036), .B(n12108), .Z(c4037) );
ANDN U20181 ( .B(n12109), .A(n12110), .Z(n12108) );
XOR U20182 ( .A(c4036), .B(b[4036]), .Z(n12109) );
XNOR U20183 ( .A(b[4036]), .B(n12110), .Z(c[4036]) );
XNOR U20184 ( .A(a[4036]), .B(c4036), .Z(n12110) );
XOR U20185 ( .A(c4037), .B(n12111), .Z(c4038) );
ANDN U20186 ( .B(n12112), .A(n12113), .Z(n12111) );
XOR U20187 ( .A(c4037), .B(b[4037]), .Z(n12112) );
XNOR U20188 ( .A(b[4037]), .B(n12113), .Z(c[4037]) );
XNOR U20189 ( .A(a[4037]), .B(c4037), .Z(n12113) );
XOR U20190 ( .A(c4038), .B(n12114), .Z(c4039) );
ANDN U20191 ( .B(n12115), .A(n12116), .Z(n12114) );
XOR U20192 ( .A(c4038), .B(b[4038]), .Z(n12115) );
XNOR U20193 ( .A(b[4038]), .B(n12116), .Z(c[4038]) );
XNOR U20194 ( .A(a[4038]), .B(c4038), .Z(n12116) );
XOR U20195 ( .A(c4039), .B(n12117), .Z(c4040) );
ANDN U20196 ( .B(n12118), .A(n12119), .Z(n12117) );
XOR U20197 ( .A(c4039), .B(b[4039]), .Z(n12118) );
XNOR U20198 ( .A(b[4039]), .B(n12119), .Z(c[4039]) );
XNOR U20199 ( .A(a[4039]), .B(c4039), .Z(n12119) );
XOR U20200 ( .A(c4040), .B(n12120), .Z(c4041) );
ANDN U20201 ( .B(n12121), .A(n12122), .Z(n12120) );
XOR U20202 ( .A(c4040), .B(b[4040]), .Z(n12121) );
XNOR U20203 ( .A(b[4040]), .B(n12122), .Z(c[4040]) );
XNOR U20204 ( .A(a[4040]), .B(c4040), .Z(n12122) );
XOR U20205 ( .A(c4041), .B(n12123), .Z(c4042) );
ANDN U20206 ( .B(n12124), .A(n12125), .Z(n12123) );
XOR U20207 ( .A(c4041), .B(b[4041]), .Z(n12124) );
XNOR U20208 ( .A(b[4041]), .B(n12125), .Z(c[4041]) );
XNOR U20209 ( .A(a[4041]), .B(c4041), .Z(n12125) );
XOR U20210 ( .A(c4042), .B(n12126), .Z(c4043) );
ANDN U20211 ( .B(n12127), .A(n12128), .Z(n12126) );
XOR U20212 ( .A(c4042), .B(b[4042]), .Z(n12127) );
XNOR U20213 ( .A(b[4042]), .B(n12128), .Z(c[4042]) );
XNOR U20214 ( .A(a[4042]), .B(c4042), .Z(n12128) );
XOR U20215 ( .A(c4043), .B(n12129), .Z(c4044) );
ANDN U20216 ( .B(n12130), .A(n12131), .Z(n12129) );
XOR U20217 ( .A(c4043), .B(b[4043]), .Z(n12130) );
XNOR U20218 ( .A(b[4043]), .B(n12131), .Z(c[4043]) );
XNOR U20219 ( .A(a[4043]), .B(c4043), .Z(n12131) );
XOR U20220 ( .A(c4044), .B(n12132), .Z(c4045) );
ANDN U20221 ( .B(n12133), .A(n12134), .Z(n12132) );
XOR U20222 ( .A(c4044), .B(b[4044]), .Z(n12133) );
XNOR U20223 ( .A(b[4044]), .B(n12134), .Z(c[4044]) );
XNOR U20224 ( .A(a[4044]), .B(c4044), .Z(n12134) );
XOR U20225 ( .A(c4045), .B(n12135), .Z(c4046) );
ANDN U20226 ( .B(n12136), .A(n12137), .Z(n12135) );
XOR U20227 ( .A(c4045), .B(b[4045]), .Z(n12136) );
XNOR U20228 ( .A(b[4045]), .B(n12137), .Z(c[4045]) );
XNOR U20229 ( .A(a[4045]), .B(c4045), .Z(n12137) );
XOR U20230 ( .A(c4046), .B(n12138), .Z(c4047) );
ANDN U20231 ( .B(n12139), .A(n12140), .Z(n12138) );
XOR U20232 ( .A(c4046), .B(b[4046]), .Z(n12139) );
XNOR U20233 ( .A(b[4046]), .B(n12140), .Z(c[4046]) );
XNOR U20234 ( .A(a[4046]), .B(c4046), .Z(n12140) );
XOR U20235 ( .A(c4047), .B(n12141), .Z(c4048) );
ANDN U20236 ( .B(n12142), .A(n12143), .Z(n12141) );
XOR U20237 ( .A(c4047), .B(b[4047]), .Z(n12142) );
XNOR U20238 ( .A(b[4047]), .B(n12143), .Z(c[4047]) );
XNOR U20239 ( .A(a[4047]), .B(c4047), .Z(n12143) );
XOR U20240 ( .A(c4048), .B(n12144), .Z(c4049) );
ANDN U20241 ( .B(n12145), .A(n12146), .Z(n12144) );
XOR U20242 ( .A(c4048), .B(b[4048]), .Z(n12145) );
XNOR U20243 ( .A(b[4048]), .B(n12146), .Z(c[4048]) );
XNOR U20244 ( .A(a[4048]), .B(c4048), .Z(n12146) );
XOR U20245 ( .A(c4049), .B(n12147), .Z(c4050) );
ANDN U20246 ( .B(n12148), .A(n12149), .Z(n12147) );
XOR U20247 ( .A(c4049), .B(b[4049]), .Z(n12148) );
XNOR U20248 ( .A(b[4049]), .B(n12149), .Z(c[4049]) );
XNOR U20249 ( .A(a[4049]), .B(c4049), .Z(n12149) );
XOR U20250 ( .A(c4050), .B(n12150), .Z(c4051) );
ANDN U20251 ( .B(n12151), .A(n12152), .Z(n12150) );
XOR U20252 ( .A(c4050), .B(b[4050]), .Z(n12151) );
XNOR U20253 ( .A(b[4050]), .B(n12152), .Z(c[4050]) );
XNOR U20254 ( .A(a[4050]), .B(c4050), .Z(n12152) );
XOR U20255 ( .A(c4051), .B(n12153), .Z(c4052) );
ANDN U20256 ( .B(n12154), .A(n12155), .Z(n12153) );
XOR U20257 ( .A(c4051), .B(b[4051]), .Z(n12154) );
XNOR U20258 ( .A(b[4051]), .B(n12155), .Z(c[4051]) );
XNOR U20259 ( .A(a[4051]), .B(c4051), .Z(n12155) );
XOR U20260 ( .A(c4052), .B(n12156), .Z(c4053) );
ANDN U20261 ( .B(n12157), .A(n12158), .Z(n12156) );
XOR U20262 ( .A(c4052), .B(b[4052]), .Z(n12157) );
XNOR U20263 ( .A(b[4052]), .B(n12158), .Z(c[4052]) );
XNOR U20264 ( .A(a[4052]), .B(c4052), .Z(n12158) );
XOR U20265 ( .A(c4053), .B(n12159), .Z(c4054) );
ANDN U20266 ( .B(n12160), .A(n12161), .Z(n12159) );
XOR U20267 ( .A(c4053), .B(b[4053]), .Z(n12160) );
XNOR U20268 ( .A(b[4053]), .B(n12161), .Z(c[4053]) );
XNOR U20269 ( .A(a[4053]), .B(c4053), .Z(n12161) );
XOR U20270 ( .A(c4054), .B(n12162), .Z(c4055) );
ANDN U20271 ( .B(n12163), .A(n12164), .Z(n12162) );
XOR U20272 ( .A(c4054), .B(b[4054]), .Z(n12163) );
XNOR U20273 ( .A(b[4054]), .B(n12164), .Z(c[4054]) );
XNOR U20274 ( .A(a[4054]), .B(c4054), .Z(n12164) );
XOR U20275 ( .A(c4055), .B(n12165), .Z(c4056) );
ANDN U20276 ( .B(n12166), .A(n12167), .Z(n12165) );
XOR U20277 ( .A(c4055), .B(b[4055]), .Z(n12166) );
XNOR U20278 ( .A(b[4055]), .B(n12167), .Z(c[4055]) );
XNOR U20279 ( .A(a[4055]), .B(c4055), .Z(n12167) );
XOR U20280 ( .A(c4056), .B(n12168), .Z(c4057) );
ANDN U20281 ( .B(n12169), .A(n12170), .Z(n12168) );
XOR U20282 ( .A(c4056), .B(b[4056]), .Z(n12169) );
XNOR U20283 ( .A(b[4056]), .B(n12170), .Z(c[4056]) );
XNOR U20284 ( .A(a[4056]), .B(c4056), .Z(n12170) );
XOR U20285 ( .A(c4057), .B(n12171), .Z(c4058) );
ANDN U20286 ( .B(n12172), .A(n12173), .Z(n12171) );
XOR U20287 ( .A(c4057), .B(b[4057]), .Z(n12172) );
XNOR U20288 ( .A(b[4057]), .B(n12173), .Z(c[4057]) );
XNOR U20289 ( .A(a[4057]), .B(c4057), .Z(n12173) );
XOR U20290 ( .A(c4058), .B(n12174), .Z(c4059) );
ANDN U20291 ( .B(n12175), .A(n12176), .Z(n12174) );
XOR U20292 ( .A(c4058), .B(b[4058]), .Z(n12175) );
XNOR U20293 ( .A(b[4058]), .B(n12176), .Z(c[4058]) );
XNOR U20294 ( .A(a[4058]), .B(c4058), .Z(n12176) );
XOR U20295 ( .A(c4059), .B(n12177), .Z(c4060) );
ANDN U20296 ( .B(n12178), .A(n12179), .Z(n12177) );
XOR U20297 ( .A(c4059), .B(b[4059]), .Z(n12178) );
XNOR U20298 ( .A(b[4059]), .B(n12179), .Z(c[4059]) );
XNOR U20299 ( .A(a[4059]), .B(c4059), .Z(n12179) );
XOR U20300 ( .A(c4060), .B(n12180), .Z(c4061) );
ANDN U20301 ( .B(n12181), .A(n12182), .Z(n12180) );
XOR U20302 ( .A(c4060), .B(b[4060]), .Z(n12181) );
XNOR U20303 ( .A(b[4060]), .B(n12182), .Z(c[4060]) );
XNOR U20304 ( .A(a[4060]), .B(c4060), .Z(n12182) );
XOR U20305 ( .A(c4061), .B(n12183), .Z(c4062) );
ANDN U20306 ( .B(n12184), .A(n12185), .Z(n12183) );
XOR U20307 ( .A(c4061), .B(b[4061]), .Z(n12184) );
XNOR U20308 ( .A(b[4061]), .B(n12185), .Z(c[4061]) );
XNOR U20309 ( .A(a[4061]), .B(c4061), .Z(n12185) );
XOR U20310 ( .A(c4062), .B(n12186), .Z(c4063) );
ANDN U20311 ( .B(n12187), .A(n12188), .Z(n12186) );
XOR U20312 ( .A(c4062), .B(b[4062]), .Z(n12187) );
XNOR U20313 ( .A(b[4062]), .B(n12188), .Z(c[4062]) );
XNOR U20314 ( .A(a[4062]), .B(c4062), .Z(n12188) );
XOR U20315 ( .A(c4063), .B(n12189), .Z(c4064) );
ANDN U20316 ( .B(n12190), .A(n12191), .Z(n12189) );
XOR U20317 ( .A(c4063), .B(b[4063]), .Z(n12190) );
XNOR U20318 ( .A(b[4063]), .B(n12191), .Z(c[4063]) );
XNOR U20319 ( .A(a[4063]), .B(c4063), .Z(n12191) );
XOR U20320 ( .A(c4064), .B(n12192), .Z(c4065) );
ANDN U20321 ( .B(n12193), .A(n12194), .Z(n12192) );
XOR U20322 ( .A(c4064), .B(b[4064]), .Z(n12193) );
XNOR U20323 ( .A(b[4064]), .B(n12194), .Z(c[4064]) );
XNOR U20324 ( .A(a[4064]), .B(c4064), .Z(n12194) );
XOR U20325 ( .A(c4065), .B(n12195), .Z(c4066) );
ANDN U20326 ( .B(n12196), .A(n12197), .Z(n12195) );
XOR U20327 ( .A(c4065), .B(b[4065]), .Z(n12196) );
XNOR U20328 ( .A(b[4065]), .B(n12197), .Z(c[4065]) );
XNOR U20329 ( .A(a[4065]), .B(c4065), .Z(n12197) );
XOR U20330 ( .A(c4066), .B(n12198), .Z(c4067) );
ANDN U20331 ( .B(n12199), .A(n12200), .Z(n12198) );
XOR U20332 ( .A(c4066), .B(b[4066]), .Z(n12199) );
XNOR U20333 ( .A(b[4066]), .B(n12200), .Z(c[4066]) );
XNOR U20334 ( .A(a[4066]), .B(c4066), .Z(n12200) );
XOR U20335 ( .A(c4067), .B(n12201), .Z(c4068) );
ANDN U20336 ( .B(n12202), .A(n12203), .Z(n12201) );
XOR U20337 ( .A(c4067), .B(b[4067]), .Z(n12202) );
XNOR U20338 ( .A(b[4067]), .B(n12203), .Z(c[4067]) );
XNOR U20339 ( .A(a[4067]), .B(c4067), .Z(n12203) );
XOR U20340 ( .A(c4068), .B(n12204), .Z(c4069) );
ANDN U20341 ( .B(n12205), .A(n12206), .Z(n12204) );
XOR U20342 ( .A(c4068), .B(b[4068]), .Z(n12205) );
XNOR U20343 ( .A(b[4068]), .B(n12206), .Z(c[4068]) );
XNOR U20344 ( .A(a[4068]), .B(c4068), .Z(n12206) );
XOR U20345 ( .A(c4069), .B(n12207), .Z(c4070) );
ANDN U20346 ( .B(n12208), .A(n12209), .Z(n12207) );
XOR U20347 ( .A(c4069), .B(b[4069]), .Z(n12208) );
XNOR U20348 ( .A(b[4069]), .B(n12209), .Z(c[4069]) );
XNOR U20349 ( .A(a[4069]), .B(c4069), .Z(n12209) );
XOR U20350 ( .A(c4070), .B(n12210), .Z(c4071) );
ANDN U20351 ( .B(n12211), .A(n12212), .Z(n12210) );
XOR U20352 ( .A(c4070), .B(b[4070]), .Z(n12211) );
XNOR U20353 ( .A(b[4070]), .B(n12212), .Z(c[4070]) );
XNOR U20354 ( .A(a[4070]), .B(c4070), .Z(n12212) );
XOR U20355 ( .A(c4071), .B(n12213), .Z(c4072) );
ANDN U20356 ( .B(n12214), .A(n12215), .Z(n12213) );
XOR U20357 ( .A(c4071), .B(b[4071]), .Z(n12214) );
XNOR U20358 ( .A(b[4071]), .B(n12215), .Z(c[4071]) );
XNOR U20359 ( .A(a[4071]), .B(c4071), .Z(n12215) );
XOR U20360 ( .A(c4072), .B(n12216), .Z(c4073) );
ANDN U20361 ( .B(n12217), .A(n12218), .Z(n12216) );
XOR U20362 ( .A(c4072), .B(b[4072]), .Z(n12217) );
XNOR U20363 ( .A(b[4072]), .B(n12218), .Z(c[4072]) );
XNOR U20364 ( .A(a[4072]), .B(c4072), .Z(n12218) );
XOR U20365 ( .A(c4073), .B(n12219), .Z(c4074) );
ANDN U20366 ( .B(n12220), .A(n12221), .Z(n12219) );
XOR U20367 ( .A(c4073), .B(b[4073]), .Z(n12220) );
XNOR U20368 ( .A(b[4073]), .B(n12221), .Z(c[4073]) );
XNOR U20369 ( .A(a[4073]), .B(c4073), .Z(n12221) );
XOR U20370 ( .A(c4074), .B(n12222), .Z(c4075) );
ANDN U20371 ( .B(n12223), .A(n12224), .Z(n12222) );
XOR U20372 ( .A(c4074), .B(b[4074]), .Z(n12223) );
XNOR U20373 ( .A(b[4074]), .B(n12224), .Z(c[4074]) );
XNOR U20374 ( .A(a[4074]), .B(c4074), .Z(n12224) );
XOR U20375 ( .A(c4075), .B(n12225), .Z(c4076) );
ANDN U20376 ( .B(n12226), .A(n12227), .Z(n12225) );
XOR U20377 ( .A(c4075), .B(b[4075]), .Z(n12226) );
XNOR U20378 ( .A(b[4075]), .B(n12227), .Z(c[4075]) );
XNOR U20379 ( .A(a[4075]), .B(c4075), .Z(n12227) );
XOR U20380 ( .A(c4076), .B(n12228), .Z(c4077) );
ANDN U20381 ( .B(n12229), .A(n12230), .Z(n12228) );
XOR U20382 ( .A(c4076), .B(b[4076]), .Z(n12229) );
XNOR U20383 ( .A(b[4076]), .B(n12230), .Z(c[4076]) );
XNOR U20384 ( .A(a[4076]), .B(c4076), .Z(n12230) );
XOR U20385 ( .A(c4077), .B(n12231), .Z(c4078) );
ANDN U20386 ( .B(n12232), .A(n12233), .Z(n12231) );
XOR U20387 ( .A(c4077), .B(b[4077]), .Z(n12232) );
XNOR U20388 ( .A(b[4077]), .B(n12233), .Z(c[4077]) );
XNOR U20389 ( .A(a[4077]), .B(c4077), .Z(n12233) );
XOR U20390 ( .A(c4078), .B(n12234), .Z(c4079) );
ANDN U20391 ( .B(n12235), .A(n12236), .Z(n12234) );
XOR U20392 ( .A(c4078), .B(b[4078]), .Z(n12235) );
XNOR U20393 ( .A(b[4078]), .B(n12236), .Z(c[4078]) );
XNOR U20394 ( .A(a[4078]), .B(c4078), .Z(n12236) );
XOR U20395 ( .A(c4079), .B(n12237), .Z(c4080) );
ANDN U20396 ( .B(n12238), .A(n12239), .Z(n12237) );
XOR U20397 ( .A(c4079), .B(b[4079]), .Z(n12238) );
XNOR U20398 ( .A(b[4079]), .B(n12239), .Z(c[4079]) );
XNOR U20399 ( .A(a[4079]), .B(c4079), .Z(n12239) );
XOR U20400 ( .A(c4080), .B(n12240), .Z(c4081) );
ANDN U20401 ( .B(n12241), .A(n12242), .Z(n12240) );
XOR U20402 ( .A(c4080), .B(b[4080]), .Z(n12241) );
XNOR U20403 ( .A(b[4080]), .B(n12242), .Z(c[4080]) );
XNOR U20404 ( .A(a[4080]), .B(c4080), .Z(n12242) );
XOR U20405 ( .A(c4081), .B(n12243), .Z(c4082) );
ANDN U20406 ( .B(n12244), .A(n12245), .Z(n12243) );
XOR U20407 ( .A(c4081), .B(b[4081]), .Z(n12244) );
XNOR U20408 ( .A(b[4081]), .B(n12245), .Z(c[4081]) );
XNOR U20409 ( .A(a[4081]), .B(c4081), .Z(n12245) );
XOR U20410 ( .A(c4082), .B(n12246), .Z(c4083) );
ANDN U20411 ( .B(n12247), .A(n12248), .Z(n12246) );
XOR U20412 ( .A(c4082), .B(b[4082]), .Z(n12247) );
XNOR U20413 ( .A(b[4082]), .B(n12248), .Z(c[4082]) );
XNOR U20414 ( .A(a[4082]), .B(c4082), .Z(n12248) );
XOR U20415 ( .A(c4083), .B(n12249), .Z(c4084) );
ANDN U20416 ( .B(n12250), .A(n12251), .Z(n12249) );
XOR U20417 ( .A(c4083), .B(b[4083]), .Z(n12250) );
XNOR U20418 ( .A(b[4083]), .B(n12251), .Z(c[4083]) );
XNOR U20419 ( .A(a[4083]), .B(c4083), .Z(n12251) );
XOR U20420 ( .A(c4084), .B(n12252), .Z(c4085) );
ANDN U20421 ( .B(n12253), .A(n12254), .Z(n12252) );
XOR U20422 ( .A(c4084), .B(b[4084]), .Z(n12253) );
XNOR U20423 ( .A(b[4084]), .B(n12254), .Z(c[4084]) );
XNOR U20424 ( .A(a[4084]), .B(c4084), .Z(n12254) );
XOR U20425 ( .A(c4085), .B(n12255), .Z(c4086) );
ANDN U20426 ( .B(n12256), .A(n12257), .Z(n12255) );
XOR U20427 ( .A(c4085), .B(b[4085]), .Z(n12256) );
XNOR U20428 ( .A(b[4085]), .B(n12257), .Z(c[4085]) );
XNOR U20429 ( .A(a[4085]), .B(c4085), .Z(n12257) );
XOR U20430 ( .A(c4086), .B(n12258), .Z(c4087) );
ANDN U20431 ( .B(n12259), .A(n12260), .Z(n12258) );
XOR U20432 ( .A(c4086), .B(b[4086]), .Z(n12259) );
XNOR U20433 ( .A(b[4086]), .B(n12260), .Z(c[4086]) );
XNOR U20434 ( .A(a[4086]), .B(c4086), .Z(n12260) );
XOR U20435 ( .A(c4087), .B(n12261), .Z(c4088) );
ANDN U20436 ( .B(n12262), .A(n12263), .Z(n12261) );
XOR U20437 ( .A(c4087), .B(b[4087]), .Z(n12262) );
XNOR U20438 ( .A(b[4087]), .B(n12263), .Z(c[4087]) );
XNOR U20439 ( .A(a[4087]), .B(c4087), .Z(n12263) );
XOR U20440 ( .A(c4088), .B(n12264), .Z(c4089) );
ANDN U20441 ( .B(n12265), .A(n12266), .Z(n12264) );
XOR U20442 ( .A(c4088), .B(b[4088]), .Z(n12265) );
XNOR U20443 ( .A(b[4088]), .B(n12266), .Z(c[4088]) );
XNOR U20444 ( .A(a[4088]), .B(c4088), .Z(n12266) );
XOR U20445 ( .A(c4089), .B(n12267), .Z(c4090) );
ANDN U20446 ( .B(n12268), .A(n12269), .Z(n12267) );
XOR U20447 ( .A(c4089), .B(b[4089]), .Z(n12268) );
XNOR U20448 ( .A(b[4089]), .B(n12269), .Z(c[4089]) );
XNOR U20449 ( .A(a[4089]), .B(c4089), .Z(n12269) );
XOR U20450 ( .A(c4090), .B(n12270), .Z(c4091) );
ANDN U20451 ( .B(n12271), .A(n12272), .Z(n12270) );
XOR U20452 ( .A(c4090), .B(b[4090]), .Z(n12271) );
XNOR U20453 ( .A(b[4090]), .B(n12272), .Z(c[4090]) );
XNOR U20454 ( .A(a[4090]), .B(c4090), .Z(n12272) );
XOR U20455 ( .A(c4091), .B(n12273), .Z(c4092) );
ANDN U20456 ( .B(n12274), .A(n12275), .Z(n12273) );
XOR U20457 ( .A(c4091), .B(b[4091]), .Z(n12274) );
XNOR U20458 ( .A(b[4091]), .B(n12275), .Z(c[4091]) );
XNOR U20459 ( .A(a[4091]), .B(c4091), .Z(n12275) );
XOR U20460 ( .A(c4092), .B(n12276), .Z(c4093) );
ANDN U20461 ( .B(n12277), .A(n12278), .Z(n12276) );
XOR U20462 ( .A(c4092), .B(b[4092]), .Z(n12277) );
XNOR U20463 ( .A(b[4092]), .B(n12278), .Z(c[4092]) );
XNOR U20464 ( .A(a[4092]), .B(c4092), .Z(n12278) );
XOR U20465 ( .A(c4093), .B(n12279), .Z(c4094) );
ANDN U20466 ( .B(n12280), .A(n12281), .Z(n12279) );
XOR U20467 ( .A(c4093), .B(b[4093]), .Z(n12280) );
XNOR U20468 ( .A(b[4093]), .B(n12281), .Z(c[4093]) );
XNOR U20469 ( .A(a[4093]), .B(c4093), .Z(n12281) );
XOR U20470 ( .A(c4094), .B(n12282), .Z(c4095) );
ANDN U20471 ( .B(n12283), .A(n12284), .Z(n12282) );
XOR U20472 ( .A(c4094), .B(b[4094]), .Z(n12283) );
XNOR U20473 ( .A(b[4094]), .B(n12284), .Z(c[4094]) );
XNOR U20474 ( .A(a[4094]), .B(c4094), .Z(n12284) );
XOR U20475 ( .A(c4095), .B(n12285), .Z(c4096) );
ANDN U20476 ( .B(n12286), .A(n12287), .Z(n12285) );
XOR U20477 ( .A(c4095), .B(b[4095]), .Z(n12286) );
XNOR U20478 ( .A(b[4095]), .B(n12287), .Z(c[4095]) );
XNOR U20479 ( .A(a[4095]), .B(c4095), .Z(n12287) );
XOR U20480 ( .A(c4096), .B(n12288), .Z(c4097) );
ANDN U20481 ( .B(n12289), .A(n12290), .Z(n12288) );
XOR U20482 ( .A(c4096), .B(b[4096]), .Z(n12289) );
XNOR U20483 ( .A(b[4096]), .B(n12290), .Z(c[4096]) );
XNOR U20484 ( .A(a[4096]), .B(c4096), .Z(n12290) );
XOR U20485 ( .A(c4097), .B(n12291), .Z(c4098) );
ANDN U20486 ( .B(n12292), .A(n12293), .Z(n12291) );
XOR U20487 ( .A(c4097), .B(b[4097]), .Z(n12292) );
XNOR U20488 ( .A(b[4097]), .B(n12293), .Z(c[4097]) );
XNOR U20489 ( .A(a[4097]), .B(c4097), .Z(n12293) );
XOR U20490 ( .A(c4098), .B(n12294), .Z(c4099) );
ANDN U20491 ( .B(n12295), .A(n12296), .Z(n12294) );
XOR U20492 ( .A(c4098), .B(b[4098]), .Z(n12295) );
XNOR U20493 ( .A(b[4098]), .B(n12296), .Z(c[4098]) );
XNOR U20494 ( .A(a[4098]), .B(c4098), .Z(n12296) );
XOR U20495 ( .A(c4099), .B(n12297), .Z(c4100) );
ANDN U20496 ( .B(n12298), .A(n12299), .Z(n12297) );
XOR U20497 ( .A(c4099), .B(b[4099]), .Z(n12298) );
XNOR U20498 ( .A(b[4099]), .B(n12299), .Z(c[4099]) );
XNOR U20499 ( .A(a[4099]), .B(c4099), .Z(n12299) );
XOR U20500 ( .A(c4100), .B(n12300), .Z(c4101) );
ANDN U20501 ( .B(n12301), .A(n12302), .Z(n12300) );
XOR U20502 ( .A(c4100), .B(b[4100]), .Z(n12301) );
XNOR U20503 ( .A(b[4100]), .B(n12302), .Z(c[4100]) );
XNOR U20504 ( .A(a[4100]), .B(c4100), .Z(n12302) );
XOR U20505 ( .A(c4101), .B(n12303), .Z(c4102) );
ANDN U20506 ( .B(n12304), .A(n12305), .Z(n12303) );
XOR U20507 ( .A(c4101), .B(b[4101]), .Z(n12304) );
XNOR U20508 ( .A(b[4101]), .B(n12305), .Z(c[4101]) );
XNOR U20509 ( .A(a[4101]), .B(c4101), .Z(n12305) );
XOR U20510 ( .A(c4102), .B(n12306), .Z(c4103) );
ANDN U20511 ( .B(n12307), .A(n12308), .Z(n12306) );
XOR U20512 ( .A(c4102), .B(b[4102]), .Z(n12307) );
XNOR U20513 ( .A(b[4102]), .B(n12308), .Z(c[4102]) );
XNOR U20514 ( .A(a[4102]), .B(c4102), .Z(n12308) );
XOR U20515 ( .A(c4103), .B(n12309), .Z(c4104) );
ANDN U20516 ( .B(n12310), .A(n12311), .Z(n12309) );
XOR U20517 ( .A(c4103), .B(b[4103]), .Z(n12310) );
XNOR U20518 ( .A(b[4103]), .B(n12311), .Z(c[4103]) );
XNOR U20519 ( .A(a[4103]), .B(c4103), .Z(n12311) );
XOR U20520 ( .A(c4104), .B(n12312), .Z(c4105) );
ANDN U20521 ( .B(n12313), .A(n12314), .Z(n12312) );
XOR U20522 ( .A(c4104), .B(b[4104]), .Z(n12313) );
XNOR U20523 ( .A(b[4104]), .B(n12314), .Z(c[4104]) );
XNOR U20524 ( .A(a[4104]), .B(c4104), .Z(n12314) );
XOR U20525 ( .A(c4105), .B(n12315), .Z(c4106) );
ANDN U20526 ( .B(n12316), .A(n12317), .Z(n12315) );
XOR U20527 ( .A(c4105), .B(b[4105]), .Z(n12316) );
XNOR U20528 ( .A(b[4105]), .B(n12317), .Z(c[4105]) );
XNOR U20529 ( .A(a[4105]), .B(c4105), .Z(n12317) );
XOR U20530 ( .A(c4106), .B(n12318), .Z(c4107) );
ANDN U20531 ( .B(n12319), .A(n12320), .Z(n12318) );
XOR U20532 ( .A(c4106), .B(b[4106]), .Z(n12319) );
XNOR U20533 ( .A(b[4106]), .B(n12320), .Z(c[4106]) );
XNOR U20534 ( .A(a[4106]), .B(c4106), .Z(n12320) );
XOR U20535 ( .A(c4107), .B(n12321), .Z(c4108) );
ANDN U20536 ( .B(n12322), .A(n12323), .Z(n12321) );
XOR U20537 ( .A(c4107), .B(b[4107]), .Z(n12322) );
XNOR U20538 ( .A(b[4107]), .B(n12323), .Z(c[4107]) );
XNOR U20539 ( .A(a[4107]), .B(c4107), .Z(n12323) );
XOR U20540 ( .A(c4108), .B(n12324), .Z(c4109) );
ANDN U20541 ( .B(n12325), .A(n12326), .Z(n12324) );
XOR U20542 ( .A(c4108), .B(b[4108]), .Z(n12325) );
XNOR U20543 ( .A(b[4108]), .B(n12326), .Z(c[4108]) );
XNOR U20544 ( .A(a[4108]), .B(c4108), .Z(n12326) );
XOR U20545 ( .A(c4109), .B(n12327), .Z(c4110) );
ANDN U20546 ( .B(n12328), .A(n12329), .Z(n12327) );
XOR U20547 ( .A(c4109), .B(b[4109]), .Z(n12328) );
XNOR U20548 ( .A(b[4109]), .B(n12329), .Z(c[4109]) );
XNOR U20549 ( .A(a[4109]), .B(c4109), .Z(n12329) );
XOR U20550 ( .A(c4110), .B(n12330), .Z(c4111) );
ANDN U20551 ( .B(n12331), .A(n12332), .Z(n12330) );
XOR U20552 ( .A(c4110), .B(b[4110]), .Z(n12331) );
XNOR U20553 ( .A(b[4110]), .B(n12332), .Z(c[4110]) );
XNOR U20554 ( .A(a[4110]), .B(c4110), .Z(n12332) );
XOR U20555 ( .A(c4111), .B(n12333), .Z(c4112) );
ANDN U20556 ( .B(n12334), .A(n12335), .Z(n12333) );
XOR U20557 ( .A(c4111), .B(b[4111]), .Z(n12334) );
XNOR U20558 ( .A(b[4111]), .B(n12335), .Z(c[4111]) );
XNOR U20559 ( .A(a[4111]), .B(c4111), .Z(n12335) );
XOR U20560 ( .A(c4112), .B(n12336), .Z(c4113) );
ANDN U20561 ( .B(n12337), .A(n12338), .Z(n12336) );
XOR U20562 ( .A(c4112), .B(b[4112]), .Z(n12337) );
XNOR U20563 ( .A(b[4112]), .B(n12338), .Z(c[4112]) );
XNOR U20564 ( .A(a[4112]), .B(c4112), .Z(n12338) );
XOR U20565 ( .A(c4113), .B(n12339), .Z(c4114) );
ANDN U20566 ( .B(n12340), .A(n12341), .Z(n12339) );
XOR U20567 ( .A(c4113), .B(b[4113]), .Z(n12340) );
XNOR U20568 ( .A(b[4113]), .B(n12341), .Z(c[4113]) );
XNOR U20569 ( .A(a[4113]), .B(c4113), .Z(n12341) );
XOR U20570 ( .A(c4114), .B(n12342), .Z(c4115) );
ANDN U20571 ( .B(n12343), .A(n12344), .Z(n12342) );
XOR U20572 ( .A(c4114), .B(b[4114]), .Z(n12343) );
XNOR U20573 ( .A(b[4114]), .B(n12344), .Z(c[4114]) );
XNOR U20574 ( .A(a[4114]), .B(c4114), .Z(n12344) );
XOR U20575 ( .A(c4115), .B(n12345), .Z(c4116) );
ANDN U20576 ( .B(n12346), .A(n12347), .Z(n12345) );
XOR U20577 ( .A(c4115), .B(b[4115]), .Z(n12346) );
XNOR U20578 ( .A(b[4115]), .B(n12347), .Z(c[4115]) );
XNOR U20579 ( .A(a[4115]), .B(c4115), .Z(n12347) );
XOR U20580 ( .A(c4116), .B(n12348), .Z(c4117) );
ANDN U20581 ( .B(n12349), .A(n12350), .Z(n12348) );
XOR U20582 ( .A(c4116), .B(b[4116]), .Z(n12349) );
XNOR U20583 ( .A(b[4116]), .B(n12350), .Z(c[4116]) );
XNOR U20584 ( .A(a[4116]), .B(c4116), .Z(n12350) );
XOR U20585 ( .A(c4117), .B(n12351), .Z(c4118) );
ANDN U20586 ( .B(n12352), .A(n12353), .Z(n12351) );
XOR U20587 ( .A(c4117), .B(b[4117]), .Z(n12352) );
XNOR U20588 ( .A(b[4117]), .B(n12353), .Z(c[4117]) );
XNOR U20589 ( .A(a[4117]), .B(c4117), .Z(n12353) );
XOR U20590 ( .A(c4118), .B(n12354), .Z(c4119) );
ANDN U20591 ( .B(n12355), .A(n12356), .Z(n12354) );
XOR U20592 ( .A(c4118), .B(b[4118]), .Z(n12355) );
XNOR U20593 ( .A(b[4118]), .B(n12356), .Z(c[4118]) );
XNOR U20594 ( .A(a[4118]), .B(c4118), .Z(n12356) );
XOR U20595 ( .A(c4119), .B(n12357), .Z(c4120) );
ANDN U20596 ( .B(n12358), .A(n12359), .Z(n12357) );
XOR U20597 ( .A(c4119), .B(b[4119]), .Z(n12358) );
XNOR U20598 ( .A(b[4119]), .B(n12359), .Z(c[4119]) );
XNOR U20599 ( .A(a[4119]), .B(c4119), .Z(n12359) );
XOR U20600 ( .A(c4120), .B(n12360), .Z(c4121) );
ANDN U20601 ( .B(n12361), .A(n12362), .Z(n12360) );
XOR U20602 ( .A(c4120), .B(b[4120]), .Z(n12361) );
XNOR U20603 ( .A(b[4120]), .B(n12362), .Z(c[4120]) );
XNOR U20604 ( .A(a[4120]), .B(c4120), .Z(n12362) );
XOR U20605 ( .A(c4121), .B(n12363), .Z(c4122) );
ANDN U20606 ( .B(n12364), .A(n12365), .Z(n12363) );
XOR U20607 ( .A(c4121), .B(b[4121]), .Z(n12364) );
XNOR U20608 ( .A(b[4121]), .B(n12365), .Z(c[4121]) );
XNOR U20609 ( .A(a[4121]), .B(c4121), .Z(n12365) );
XOR U20610 ( .A(c4122), .B(n12366), .Z(c4123) );
ANDN U20611 ( .B(n12367), .A(n12368), .Z(n12366) );
XOR U20612 ( .A(c4122), .B(b[4122]), .Z(n12367) );
XNOR U20613 ( .A(b[4122]), .B(n12368), .Z(c[4122]) );
XNOR U20614 ( .A(a[4122]), .B(c4122), .Z(n12368) );
XOR U20615 ( .A(c4123), .B(n12369), .Z(c4124) );
ANDN U20616 ( .B(n12370), .A(n12371), .Z(n12369) );
XOR U20617 ( .A(c4123), .B(b[4123]), .Z(n12370) );
XNOR U20618 ( .A(b[4123]), .B(n12371), .Z(c[4123]) );
XNOR U20619 ( .A(a[4123]), .B(c4123), .Z(n12371) );
XOR U20620 ( .A(c4124), .B(n12372), .Z(c4125) );
ANDN U20621 ( .B(n12373), .A(n12374), .Z(n12372) );
XOR U20622 ( .A(c4124), .B(b[4124]), .Z(n12373) );
XNOR U20623 ( .A(b[4124]), .B(n12374), .Z(c[4124]) );
XNOR U20624 ( .A(a[4124]), .B(c4124), .Z(n12374) );
XOR U20625 ( .A(c4125), .B(n12375), .Z(c4126) );
ANDN U20626 ( .B(n12376), .A(n12377), .Z(n12375) );
XOR U20627 ( .A(c4125), .B(b[4125]), .Z(n12376) );
XNOR U20628 ( .A(b[4125]), .B(n12377), .Z(c[4125]) );
XNOR U20629 ( .A(a[4125]), .B(c4125), .Z(n12377) );
XOR U20630 ( .A(c4126), .B(n12378), .Z(c4127) );
ANDN U20631 ( .B(n12379), .A(n12380), .Z(n12378) );
XOR U20632 ( .A(c4126), .B(b[4126]), .Z(n12379) );
XNOR U20633 ( .A(b[4126]), .B(n12380), .Z(c[4126]) );
XNOR U20634 ( .A(a[4126]), .B(c4126), .Z(n12380) );
XOR U20635 ( .A(c4127), .B(n12381), .Z(c4128) );
ANDN U20636 ( .B(n12382), .A(n12383), .Z(n12381) );
XOR U20637 ( .A(c4127), .B(b[4127]), .Z(n12382) );
XNOR U20638 ( .A(b[4127]), .B(n12383), .Z(c[4127]) );
XNOR U20639 ( .A(a[4127]), .B(c4127), .Z(n12383) );
XOR U20640 ( .A(c4128), .B(n12384), .Z(c4129) );
ANDN U20641 ( .B(n12385), .A(n12386), .Z(n12384) );
XOR U20642 ( .A(c4128), .B(b[4128]), .Z(n12385) );
XNOR U20643 ( .A(b[4128]), .B(n12386), .Z(c[4128]) );
XNOR U20644 ( .A(a[4128]), .B(c4128), .Z(n12386) );
XOR U20645 ( .A(c4129), .B(n12387), .Z(c4130) );
ANDN U20646 ( .B(n12388), .A(n12389), .Z(n12387) );
XOR U20647 ( .A(c4129), .B(b[4129]), .Z(n12388) );
XNOR U20648 ( .A(b[4129]), .B(n12389), .Z(c[4129]) );
XNOR U20649 ( .A(a[4129]), .B(c4129), .Z(n12389) );
XOR U20650 ( .A(c4130), .B(n12390), .Z(c4131) );
ANDN U20651 ( .B(n12391), .A(n12392), .Z(n12390) );
XOR U20652 ( .A(c4130), .B(b[4130]), .Z(n12391) );
XNOR U20653 ( .A(b[4130]), .B(n12392), .Z(c[4130]) );
XNOR U20654 ( .A(a[4130]), .B(c4130), .Z(n12392) );
XOR U20655 ( .A(c4131), .B(n12393), .Z(c4132) );
ANDN U20656 ( .B(n12394), .A(n12395), .Z(n12393) );
XOR U20657 ( .A(c4131), .B(b[4131]), .Z(n12394) );
XNOR U20658 ( .A(b[4131]), .B(n12395), .Z(c[4131]) );
XNOR U20659 ( .A(a[4131]), .B(c4131), .Z(n12395) );
XOR U20660 ( .A(c4132), .B(n12396), .Z(c4133) );
ANDN U20661 ( .B(n12397), .A(n12398), .Z(n12396) );
XOR U20662 ( .A(c4132), .B(b[4132]), .Z(n12397) );
XNOR U20663 ( .A(b[4132]), .B(n12398), .Z(c[4132]) );
XNOR U20664 ( .A(a[4132]), .B(c4132), .Z(n12398) );
XOR U20665 ( .A(c4133), .B(n12399), .Z(c4134) );
ANDN U20666 ( .B(n12400), .A(n12401), .Z(n12399) );
XOR U20667 ( .A(c4133), .B(b[4133]), .Z(n12400) );
XNOR U20668 ( .A(b[4133]), .B(n12401), .Z(c[4133]) );
XNOR U20669 ( .A(a[4133]), .B(c4133), .Z(n12401) );
XOR U20670 ( .A(c4134), .B(n12402), .Z(c4135) );
ANDN U20671 ( .B(n12403), .A(n12404), .Z(n12402) );
XOR U20672 ( .A(c4134), .B(b[4134]), .Z(n12403) );
XNOR U20673 ( .A(b[4134]), .B(n12404), .Z(c[4134]) );
XNOR U20674 ( .A(a[4134]), .B(c4134), .Z(n12404) );
XOR U20675 ( .A(c4135), .B(n12405), .Z(c4136) );
ANDN U20676 ( .B(n12406), .A(n12407), .Z(n12405) );
XOR U20677 ( .A(c4135), .B(b[4135]), .Z(n12406) );
XNOR U20678 ( .A(b[4135]), .B(n12407), .Z(c[4135]) );
XNOR U20679 ( .A(a[4135]), .B(c4135), .Z(n12407) );
XOR U20680 ( .A(c4136), .B(n12408), .Z(c4137) );
ANDN U20681 ( .B(n12409), .A(n12410), .Z(n12408) );
XOR U20682 ( .A(c4136), .B(b[4136]), .Z(n12409) );
XNOR U20683 ( .A(b[4136]), .B(n12410), .Z(c[4136]) );
XNOR U20684 ( .A(a[4136]), .B(c4136), .Z(n12410) );
XOR U20685 ( .A(c4137), .B(n12411), .Z(c4138) );
ANDN U20686 ( .B(n12412), .A(n12413), .Z(n12411) );
XOR U20687 ( .A(c4137), .B(b[4137]), .Z(n12412) );
XNOR U20688 ( .A(b[4137]), .B(n12413), .Z(c[4137]) );
XNOR U20689 ( .A(a[4137]), .B(c4137), .Z(n12413) );
XOR U20690 ( .A(c4138), .B(n12414), .Z(c4139) );
ANDN U20691 ( .B(n12415), .A(n12416), .Z(n12414) );
XOR U20692 ( .A(c4138), .B(b[4138]), .Z(n12415) );
XNOR U20693 ( .A(b[4138]), .B(n12416), .Z(c[4138]) );
XNOR U20694 ( .A(a[4138]), .B(c4138), .Z(n12416) );
XOR U20695 ( .A(c4139), .B(n12417), .Z(c4140) );
ANDN U20696 ( .B(n12418), .A(n12419), .Z(n12417) );
XOR U20697 ( .A(c4139), .B(b[4139]), .Z(n12418) );
XNOR U20698 ( .A(b[4139]), .B(n12419), .Z(c[4139]) );
XNOR U20699 ( .A(a[4139]), .B(c4139), .Z(n12419) );
XOR U20700 ( .A(c4140), .B(n12420), .Z(c4141) );
ANDN U20701 ( .B(n12421), .A(n12422), .Z(n12420) );
XOR U20702 ( .A(c4140), .B(b[4140]), .Z(n12421) );
XNOR U20703 ( .A(b[4140]), .B(n12422), .Z(c[4140]) );
XNOR U20704 ( .A(a[4140]), .B(c4140), .Z(n12422) );
XOR U20705 ( .A(c4141), .B(n12423), .Z(c4142) );
ANDN U20706 ( .B(n12424), .A(n12425), .Z(n12423) );
XOR U20707 ( .A(c4141), .B(b[4141]), .Z(n12424) );
XNOR U20708 ( .A(b[4141]), .B(n12425), .Z(c[4141]) );
XNOR U20709 ( .A(a[4141]), .B(c4141), .Z(n12425) );
XOR U20710 ( .A(c4142), .B(n12426), .Z(c4143) );
ANDN U20711 ( .B(n12427), .A(n12428), .Z(n12426) );
XOR U20712 ( .A(c4142), .B(b[4142]), .Z(n12427) );
XNOR U20713 ( .A(b[4142]), .B(n12428), .Z(c[4142]) );
XNOR U20714 ( .A(a[4142]), .B(c4142), .Z(n12428) );
XOR U20715 ( .A(c4143), .B(n12429), .Z(c4144) );
ANDN U20716 ( .B(n12430), .A(n12431), .Z(n12429) );
XOR U20717 ( .A(c4143), .B(b[4143]), .Z(n12430) );
XNOR U20718 ( .A(b[4143]), .B(n12431), .Z(c[4143]) );
XNOR U20719 ( .A(a[4143]), .B(c4143), .Z(n12431) );
XOR U20720 ( .A(c4144), .B(n12432), .Z(c4145) );
ANDN U20721 ( .B(n12433), .A(n12434), .Z(n12432) );
XOR U20722 ( .A(c4144), .B(b[4144]), .Z(n12433) );
XNOR U20723 ( .A(b[4144]), .B(n12434), .Z(c[4144]) );
XNOR U20724 ( .A(a[4144]), .B(c4144), .Z(n12434) );
XOR U20725 ( .A(c4145), .B(n12435), .Z(c4146) );
ANDN U20726 ( .B(n12436), .A(n12437), .Z(n12435) );
XOR U20727 ( .A(c4145), .B(b[4145]), .Z(n12436) );
XNOR U20728 ( .A(b[4145]), .B(n12437), .Z(c[4145]) );
XNOR U20729 ( .A(a[4145]), .B(c4145), .Z(n12437) );
XOR U20730 ( .A(c4146), .B(n12438), .Z(c4147) );
ANDN U20731 ( .B(n12439), .A(n12440), .Z(n12438) );
XOR U20732 ( .A(c4146), .B(b[4146]), .Z(n12439) );
XNOR U20733 ( .A(b[4146]), .B(n12440), .Z(c[4146]) );
XNOR U20734 ( .A(a[4146]), .B(c4146), .Z(n12440) );
XOR U20735 ( .A(c4147), .B(n12441), .Z(c4148) );
ANDN U20736 ( .B(n12442), .A(n12443), .Z(n12441) );
XOR U20737 ( .A(c4147), .B(b[4147]), .Z(n12442) );
XNOR U20738 ( .A(b[4147]), .B(n12443), .Z(c[4147]) );
XNOR U20739 ( .A(a[4147]), .B(c4147), .Z(n12443) );
XOR U20740 ( .A(c4148), .B(n12444), .Z(c4149) );
ANDN U20741 ( .B(n12445), .A(n12446), .Z(n12444) );
XOR U20742 ( .A(c4148), .B(b[4148]), .Z(n12445) );
XNOR U20743 ( .A(b[4148]), .B(n12446), .Z(c[4148]) );
XNOR U20744 ( .A(a[4148]), .B(c4148), .Z(n12446) );
XOR U20745 ( .A(c4149), .B(n12447), .Z(c4150) );
ANDN U20746 ( .B(n12448), .A(n12449), .Z(n12447) );
XOR U20747 ( .A(c4149), .B(b[4149]), .Z(n12448) );
XNOR U20748 ( .A(b[4149]), .B(n12449), .Z(c[4149]) );
XNOR U20749 ( .A(a[4149]), .B(c4149), .Z(n12449) );
XOR U20750 ( .A(c4150), .B(n12450), .Z(c4151) );
ANDN U20751 ( .B(n12451), .A(n12452), .Z(n12450) );
XOR U20752 ( .A(c4150), .B(b[4150]), .Z(n12451) );
XNOR U20753 ( .A(b[4150]), .B(n12452), .Z(c[4150]) );
XNOR U20754 ( .A(a[4150]), .B(c4150), .Z(n12452) );
XOR U20755 ( .A(c4151), .B(n12453), .Z(c4152) );
ANDN U20756 ( .B(n12454), .A(n12455), .Z(n12453) );
XOR U20757 ( .A(c4151), .B(b[4151]), .Z(n12454) );
XNOR U20758 ( .A(b[4151]), .B(n12455), .Z(c[4151]) );
XNOR U20759 ( .A(a[4151]), .B(c4151), .Z(n12455) );
XOR U20760 ( .A(c4152), .B(n12456), .Z(c4153) );
ANDN U20761 ( .B(n12457), .A(n12458), .Z(n12456) );
XOR U20762 ( .A(c4152), .B(b[4152]), .Z(n12457) );
XNOR U20763 ( .A(b[4152]), .B(n12458), .Z(c[4152]) );
XNOR U20764 ( .A(a[4152]), .B(c4152), .Z(n12458) );
XOR U20765 ( .A(c4153), .B(n12459), .Z(c4154) );
ANDN U20766 ( .B(n12460), .A(n12461), .Z(n12459) );
XOR U20767 ( .A(c4153), .B(b[4153]), .Z(n12460) );
XNOR U20768 ( .A(b[4153]), .B(n12461), .Z(c[4153]) );
XNOR U20769 ( .A(a[4153]), .B(c4153), .Z(n12461) );
XOR U20770 ( .A(c4154), .B(n12462), .Z(c4155) );
ANDN U20771 ( .B(n12463), .A(n12464), .Z(n12462) );
XOR U20772 ( .A(c4154), .B(b[4154]), .Z(n12463) );
XNOR U20773 ( .A(b[4154]), .B(n12464), .Z(c[4154]) );
XNOR U20774 ( .A(a[4154]), .B(c4154), .Z(n12464) );
XOR U20775 ( .A(c4155), .B(n12465), .Z(c4156) );
ANDN U20776 ( .B(n12466), .A(n12467), .Z(n12465) );
XOR U20777 ( .A(c4155), .B(b[4155]), .Z(n12466) );
XNOR U20778 ( .A(b[4155]), .B(n12467), .Z(c[4155]) );
XNOR U20779 ( .A(a[4155]), .B(c4155), .Z(n12467) );
XOR U20780 ( .A(c4156), .B(n12468), .Z(c4157) );
ANDN U20781 ( .B(n12469), .A(n12470), .Z(n12468) );
XOR U20782 ( .A(c4156), .B(b[4156]), .Z(n12469) );
XNOR U20783 ( .A(b[4156]), .B(n12470), .Z(c[4156]) );
XNOR U20784 ( .A(a[4156]), .B(c4156), .Z(n12470) );
XOR U20785 ( .A(c4157), .B(n12471), .Z(c4158) );
ANDN U20786 ( .B(n12472), .A(n12473), .Z(n12471) );
XOR U20787 ( .A(c4157), .B(b[4157]), .Z(n12472) );
XNOR U20788 ( .A(b[4157]), .B(n12473), .Z(c[4157]) );
XNOR U20789 ( .A(a[4157]), .B(c4157), .Z(n12473) );
XOR U20790 ( .A(c4158), .B(n12474), .Z(c4159) );
ANDN U20791 ( .B(n12475), .A(n12476), .Z(n12474) );
XOR U20792 ( .A(c4158), .B(b[4158]), .Z(n12475) );
XNOR U20793 ( .A(b[4158]), .B(n12476), .Z(c[4158]) );
XNOR U20794 ( .A(a[4158]), .B(c4158), .Z(n12476) );
XOR U20795 ( .A(c4159), .B(n12477), .Z(c4160) );
ANDN U20796 ( .B(n12478), .A(n12479), .Z(n12477) );
XOR U20797 ( .A(c4159), .B(b[4159]), .Z(n12478) );
XNOR U20798 ( .A(b[4159]), .B(n12479), .Z(c[4159]) );
XNOR U20799 ( .A(a[4159]), .B(c4159), .Z(n12479) );
XOR U20800 ( .A(c4160), .B(n12480), .Z(c4161) );
ANDN U20801 ( .B(n12481), .A(n12482), .Z(n12480) );
XOR U20802 ( .A(c4160), .B(b[4160]), .Z(n12481) );
XNOR U20803 ( .A(b[4160]), .B(n12482), .Z(c[4160]) );
XNOR U20804 ( .A(a[4160]), .B(c4160), .Z(n12482) );
XOR U20805 ( .A(c4161), .B(n12483), .Z(c4162) );
ANDN U20806 ( .B(n12484), .A(n12485), .Z(n12483) );
XOR U20807 ( .A(c4161), .B(b[4161]), .Z(n12484) );
XNOR U20808 ( .A(b[4161]), .B(n12485), .Z(c[4161]) );
XNOR U20809 ( .A(a[4161]), .B(c4161), .Z(n12485) );
XOR U20810 ( .A(c4162), .B(n12486), .Z(c4163) );
ANDN U20811 ( .B(n12487), .A(n12488), .Z(n12486) );
XOR U20812 ( .A(c4162), .B(b[4162]), .Z(n12487) );
XNOR U20813 ( .A(b[4162]), .B(n12488), .Z(c[4162]) );
XNOR U20814 ( .A(a[4162]), .B(c4162), .Z(n12488) );
XOR U20815 ( .A(c4163), .B(n12489), .Z(c4164) );
ANDN U20816 ( .B(n12490), .A(n12491), .Z(n12489) );
XOR U20817 ( .A(c4163), .B(b[4163]), .Z(n12490) );
XNOR U20818 ( .A(b[4163]), .B(n12491), .Z(c[4163]) );
XNOR U20819 ( .A(a[4163]), .B(c4163), .Z(n12491) );
XOR U20820 ( .A(c4164), .B(n12492), .Z(c4165) );
ANDN U20821 ( .B(n12493), .A(n12494), .Z(n12492) );
XOR U20822 ( .A(c4164), .B(b[4164]), .Z(n12493) );
XNOR U20823 ( .A(b[4164]), .B(n12494), .Z(c[4164]) );
XNOR U20824 ( .A(a[4164]), .B(c4164), .Z(n12494) );
XOR U20825 ( .A(c4165), .B(n12495), .Z(c4166) );
ANDN U20826 ( .B(n12496), .A(n12497), .Z(n12495) );
XOR U20827 ( .A(c4165), .B(b[4165]), .Z(n12496) );
XNOR U20828 ( .A(b[4165]), .B(n12497), .Z(c[4165]) );
XNOR U20829 ( .A(a[4165]), .B(c4165), .Z(n12497) );
XOR U20830 ( .A(c4166), .B(n12498), .Z(c4167) );
ANDN U20831 ( .B(n12499), .A(n12500), .Z(n12498) );
XOR U20832 ( .A(c4166), .B(b[4166]), .Z(n12499) );
XNOR U20833 ( .A(b[4166]), .B(n12500), .Z(c[4166]) );
XNOR U20834 ( .A(a[4166]), .B(c4166), .Z(n12500) );
XOR U20835 ( .A(c4167), .B(n12501), .Z(c4168) );
ANDN U20836 ( .B(n12502), .A(n12503), .Z(n12501) );
XOR U20837 ( .A(c4167), .B(b[4167]), .Z(n12502) );
XNOR U20838 ( .A(b[4167]), .B(n12503), .Z(c[4167]) );
XNOR U20839 ( .A(a[4167]), .B(c4167), .Z(n12503) );
XOR U20840 ( .A(c4168), .B(n12504), .Z(c4169) );
ANDN U20841 ( .B(n12505), .A(n12506), .Z(n12504) );
XOR U20842 ( .A(c4168), .B(b[4168]), .Z(n12505) );
XNOR U20843 ( .A(b[4168]), .B(n12506), .Z(c[4168]) );
XNOR U20844 ( .A(a[4168]), .B(c4168), .Z(n12506) );
XOR U20845 ( .A(c4169), .B(n12507), .Z(c4170) );
ANDN U20846 ( .B(n12508), .A(n12509), .Z(n12507) );
XOR U20847 ( .A(c4169), .B(b[4169]), .Z(n12508) );
XNOR U20848 ( .A(b[4169]), .B(n12509), .Z(c[4169]) );
XNOR U20849 ( .A(a[4169]), .B(c4169), .Z(n12509) );
XOR U20850 ( .A(c4170), .B(n12510), .Z(c4171) );
ANDN U20851 ( .B(n12511), .A(n12512), .Z(n12510) );
XOR U20852 ( .A(c4170), .B(b[4170]), .Z(n12511) );
XNOR U20853 ( .A(b[4170]), .B(n12512), .Z(c[4170]) );
XNOR U20854 ( .A(a[4170]), .B(c4170), .Z(n12512) );
XOR U20855 ( .A(c4171), .B(n12513), .Z(c4172) );
ANDN U20856 ( .B(n12514), .A(n12515), .Z(n12513) );
XOR U20857 ( .A(c4171), .B(b[4171]), .Z(n12514) );
XNOR U20858 ( .A(b[4171]), .B(n12515), .Z(c[4171]) );
XNOR U20859 ( .A(a[4171]), .B(c4171), .Z(n12515) );
XOR U20860 ( .A(c4172), .B(n12516), .Z(c4173) );
ANDN U20861 ( .B(n12517), .A(n12518), .Z(n12516) );
XOR U20862 ( .A(c4172), .B(b[4172]), .Z(n12517) );
XNOR U20863 ( .A(b[4172]), .B(n12518), .Z(c[4172]) );
XNOR U20864 ( .A(a[4172]), .B(c4172), .Z(n12518) );
XOR U20865 ( .A(c4173), .B(n12519), .Z(c4174) );
ANDN U20866 ( .B(n12520), .A(n12521), .Z(n12519) );
XOR U20867 ( .A(c4173), .B(b[4173]), .Z(n12520) );
XNOR U20868 ( .A(b[4173]), .B(n12521), .Z(c[4173]) );
XNOR U20869 ( .A(a[4173]), .B(c4173), .Z(n12521) );
XOR U20870 ( .A(c4174), .B(n12522), .Z(c4175) );
ANDN U20871 ( .B(n12523), .A(n12524), .Z(n12522) );
XOR U20872 ( .A(c4174), .B(b[4174]), .Z(n12523) );
XNOR U20873 ( .A(b[4174]), .B(n12524), .Z(c[4174]) );
XNOR U20874 ( .A(a[4174]), .B(c4174), .Z(n12524) );
XOR U20875 ( .A(c4175), .B(n12525), .Z(c4176) );
ANDN U20876 ( .B(n12526), .A(n12527), .Z(n12525) );
XOR U20877 ( .A(c4175), .B(b[4175]), .Z(n12526) );
XNOR U20878 ( .A(b[4175]), .B(n12527), .Z(c[4175]) );
XNOR U20879 ( .A(a[4175]), .B(c4175), .Z(n12527) );
XOR U20880 ( .A(c4176), .B(n12528), .Z(c4177) );
ANDN U20881 ( .B(n12529), .A(n12530), .Z(n12528) );
XOR U20882 ( .A(c4176), .B(b[4176]), .Z(n12529) );
XNOR U20883 ( .A(b[4176]), .B(n12530), .Z(c[4176]) );
XNOR U20884 ( .A(a[4176]), .B(c4176), .Z(n12530) );
XOR U20885 ( .A(c4177), .B(n12531), .Z(c4178) );
ANDN U20886 ( .B(n12532), .A(n12533), .Z(n12531) );
XOR U20887 ( .A(c4177), .B(b[4177]), .Z(n12532) );
XNOR U20888 ( .A(b[4177]), .B(n12533), .Z(c[4177]) );
XNOR U20889 ( .A(a[4177]), .B(c4177), .Z(n12533) );
XOR U20890 ( .A(c4178), .B(n12534), .Z(c4179) );
ANDN U20891 ( .B(n12535), .A(n12536), .Z(n12534) );
XOR U20892 ( .A(c4178), .B(b[4178]), .Z(n12535) );
XNOR U20893 ( .A(b[4178]), .B(n12536), .Z(c[4178]) );
XNOR U20894 ( .A(a[4178]), .B(c4178), .Z(n12536) );
XOR U20895 ( .A(c4179), .B(n12537), .Z(c4180) );
ANDN U20896 ( .B(n12538), .A(n12539), .Z(n12537) );
XOR U20897 ( .A(c4179), .B(b[4179]), .Z(n12538) );
XNOR U20898 ( .A(b[4179]), .B(n12539), .Z(c[4179]) );
XNOR U20899 ( .A(a[4179]), .B(c4179), .Z(n12539) );
XOR U20900 ( .A(c4180), .B(n12540), .Z(c4181) );
ANDN U20901 ( .B(n12541), .A(n12542), .Z(n12540) );
XOR U20902 ( .A(c4180), .B(b[4180]), .Z(n12541) );
XNOR U20903 ( .A(b[4180]), .B(n12542), .Z(c[4180]) );
XNOR U20904 ( .A(a[4180]), .B(c4180), .Z(n12542) );
XOR U20905 ( .A(c4181), .B(n12543), .Z(c4182) );
ANDN U20906 ( .B(n12544), .A(n12545), .Z(n12543) );
XOR U20907 ( .A(c4181), .B(b[4181]), .Z(n12544) );
XNOR U20908 ( .A(b[4181]), .B(n12545), .Z(c[4181]) );
XNOR U20909 ( .A(a[4181]), .B(c4181), .Z(n12545) );
XOR U20910 ( .A(c4182), .B(n12546), .Z(c4183) );
ANDN U20911 ( .B(n12547), .A(n12548), .Z(n12546) );
XOR U20912 ( .A(c4182), .B(b[4182]), .Z(n12547) );
XNOR U20913 ( .A(b[4182]), .B(n12548), .Z(c[4182]) );
XNOR U20914 ( .A(a[4182]), .B(c4182), .Z(n12548) );
XOR U20915 ( .A(c4183), .B(n12549), .Z(c4184) );
ANDN U20916 ( .B(n12550), .A(n12551), .Z(n12549) );
XOR U20917 ( .A(c4183), .B(b[4183]), .Z(n12550) );
XNOR U20918 ( .A(b[4183]), .B(n12551), .Z(c[4183]) );
XNOR U20919 ( .A(a[4183]), .B(c4183), .Z(n12551) );
XOR U20920 ( .A(c4184), .B(n12552), .Z(c4185) );
ANDN U20921 ( .B(n12553), .A(n12554), .Z(n12552) );
XOR U20922 ( .A(c4184), .B(b[4184]), .Z(n12553) );
XNOR U20923 ( .A(b[4184]), .B(n12554), .Z(c[4184]) );
XNOR U20924 ( .A(a[4184]), .B(c4184), .Z(n12554) );
XOR U20925 ( .A(c4185), .B(n12555), .Z(c4186) );
ANDN U20926 ( .B(n12556), .A(n12557), .Z(n12555) );
XOR U20927 ( .A(c4185), .B(b[4185]), .Z(n12556) );
XNOR U20928 ( .A(b[4185]), .B(n12557), .Z(c[4185]) );
XNOR U20929 ( .A(a[4185]), .B(c4185), .Z(n12557) );
XOR U20930 ( .A(c4186), .B(n12558), .Z(c4187) );
ANDN U20931 ( .B(n12559), .A(n12560), .Z(n12558) );
XOR U20932 ( .A(c4186), .B(b[4186]), .Z(n12559) );
XNOR U20933 ( .A(b[4186]), .B(n12560), .Z(c[4186]) );
XNOR U20934 ( .A(a[4186]), .B(c4186), .Z(n12560) );
XOR U20935 ( .A(c4187), .B(n12561), .Z(c4188) );
ANDN U20936 ( .B(n12562), .A(n12563), .Z(n12561) );
XOR U20937 ( .A(c4187), .B(b[4187]), .Z(n12562) );
XNOR U20938 ( .A(b[4187]), .B(n12563), .Z(c[4187]) );
XNOR U20939 ( .A(a[4187]), .B(c4187), .Z(n12563) );
XOR U20940 ( .A(c4188), .B(n12564), .Z(c4189) );
ANDN U20941 ( .B(n12565), .A(n12566), .Z(n12564) );
XOR U20942 ( .A(c4188), .B(b[4188]), .Z(n12565) );
XNOR U20943 ( .A(b[4188]), .B(n12566), .Z(c[4188]) );
XNOR U20944 ( .A(a[4188]), .B(c4188), .Z(n12566) );
XOR U20945 ( .A(c4189), .B(n12567), .Z(c4190) );
ANDN U20946 ( .B(n12568), .A(n12569), .Z(n12567) );
XOR U20947 ( .A(c4189), .B(b[4189]), .Z(n12568) );
XNOR U20948 ( .A(b[4189]), .B(n12569), .Z(c[4189]) );
XNOR U20949 ( .A(a[4189]), .B(c4189), .Z(n12569) );
XOR U20950 ( .A(c4190), .B(n12570), .Z(c4191) );
ANDN U20951 ( .B(n12571), .A(n12572), .Z(n12570) );
XOR U20952 ( .A(c4190), .B(b[4190]), .Z(n12571) );
XNOR U20953 ( .A(b[4190]), .B(n12572), .Z(c[4190]) );
XNOR U20954 ( .A(a[4190]), .B(c4190), .Z(n12572) );
XOR U20955 ( .A(c4191), .B(n12573), .Z(c4192) );
ANDN U20956 ( .B(n12574), .A(n12575), .Z(n12573) );
XOR U20957 ( .A(c4191), .B(b[4191]), .Z(n12574) );
XNOR U20958 ( .A(b[4191]), .B(n12575), .Z(c[4191]) );
XNOR U20959 ( .A(a[4191]), .B(c4191), .Z(n12575) );
XOR U20960 ( .A(c4192), .B(n12576), .Z(c4193) );
ANDN U20961 ( .B(n12577), .A(n12578), .Z(n12576) );
XOR U20962 ( .A(c4192), .B(b[4192]), .Z(n12577) );
XNOR U20963 ( .A(b[4192]), .B(n12578), .Z(c[4192]) );
XNOR U20964 ( .A(a[4192]), .B(c4192), .Z(n12578) );
XOR U20965 ( .A(c4193), .B(n12579), .Z(c4194) );
ANDN U20966 ( .B(n12580), .A(n12581), .Z(n12579) );
XOR U20967 ( .A(c4193), .B(b[4193]), .Z(n12580) );
XNOR U20968 ( .A(b[4193]), .B(n12581), .Z(c[4193]) );
XNOR U20969 ( .A(a[4193]), .B(c4193), .Z(n12581) );
XOR U20970 ( .A(c4194), .B(n12582), .Z(c4195) );
ANDN U20971 ( .B(n12583), .A(n12584), .Z(n12582) );
XOR U20972 ( .A(c4194), .B(b[4194]), .Z(n12583) );
XNOR U20973 ( .A(b[4194]), .B(n12584), .Z(c[4194]) );
XNOR U20974 ( .A(a[4194]), .B(c4194), .Z(n12584) );
XOR U20975 ( .A(c4195), .B(n12585), .Z(c4196) );
ANDN U20976 ( .B(n12586), .A(n12587), .Z(n12585) );
XOR U20977 ( .A(c4195), .B(b[4195]), .Z(n12586) );
XNOR U20978 ( .A(b[4195]), .B(n12587), .Z(c[4195]) );
XNOR U20979 ( .A(a[4195]), .B(c4195), .Z(n12587) );
XOR U20980 ( .A(c4196), .B(n12588), .Z(c4197) );
ANDN U20981 ( .B(n12589), .A(n12590), .Z(n12588) );
XOR U20982 ( .A(c4196), .B(b[4196]), .Z(n12589) );
XNOR U20983 ( .A(b[4196]), .B(n12590), .Z(c[4196]) );
XNOR U20984 ( .A(a[4196]), .B(c4196), .Z(n12590) );
XOR U20985 ( .A(c4197), .B(n12591), .Z(c4198) );
ANDN U20986 ( .B(n12592), .A(n12593), .Z(n12591) );
XOR U20987 ( .A(c4197), .B(b[4197]), .Z(n12592) );
XNOR U20988 ( .A(b[4197]), .B(n12593), .Z(c[4197]) );
XNOR U20989 ( .A(a[4197]), .B(c4197), .Z(n12593) );
XOR U20990 ( .A(c4198), .B(n12594), .Z(c4199) );
ANDN U20991 ( .B(n12595), .A(n12596), .Z(n12594) );
XOR U20992 ( .A(c4198), .B(b[4198]), .Z(n12595) );
XNOR U20993 ( .A(b[4198]), .B(n12596), .Z(c[4198]) );
XNOR U20994 ( .A(a[4198]), .B(c4198), .Z(n12596) );
XOR U20995 ( .A(c4199), .B(n12597), .Z(c4200) );
ANDN U20996 ( .B(n12598), .A(n12599), .Z(n12597) );
XOR U20997 ( .A(c4199), .B(b[4199]), .Z(n12598) );
XNOR U20998 ( .A(b[4199]), .B(n12599), .Z(c[4199]) );
XNOR U20999 ( .A(a[4199]), .B(c4199), .Z(n12599) );
XOR U21000 ( .A(c4200), .B(n12600), .Z(c4201) );
ANDN U21001 ( .B(n12601), .A(n12602), .Z(n12600) );
XOR U21002 ( .A(c4200), .B(b[4200]), .Z(n12601) );
XNOR U21003 ( .A(b[4200]), .B(n12602), .Z(c[4200]) );
XNOR U21004 ( .A(a[4200]), .B(c4200), .Z(n12602) );
XOR U21005 ( .A(c4201), .B(n12603), .Z(c4202) );
ANDN U21006 ( .B(n12604), .A(n12605), .Z(n12603) );
XOR U21007 ( .A(c4201), .B(b[4201]), .Z(n12604) );
XNOR U21008 ( .A(b[4201]), .B(n12605), .Z(c[4201]) );
XNOR U21009 ( .A(a[4201]), .B(c4201), .Z(n12605) );
XOR U21010 ( .A(c4202), .B(n12606), .Z(c4203) );
ANDN U21011 ( .B(n12607), .A(n12608), .Z(n12606) );
XOR U21012 ( .A(c4202), .B(b[4202]), .Z(n12607) );
XNOR U21013 ( .A(b[4202]), .B(n12608), .Z(c[4202]) );
XNOR U21014 ( .A(a[4202]), .B(c4202), .Z(n12608) );
XOR U21015 ( .A(c4203), .B(n12609), .Z(c4204) );
ANDN U21016 ( .B(n12610), .A(n12611), .Z(n12609) );
XOR U21017 ( .A(c4203), .B(b[4203]), .Z(n12610) );
XNOR U21018 ( .A(b[4203]), .B(n12611), .Z(c[4203]) );
XNOR U21019 ( .A(a[4203]), .B(c4203), .Z(n12611) );
XOR U21020 ( .A(c4204), .B(n12612), .Z(c4205) );
ANDN U21021 ( .B(n12613), .A(n12614), .Z(n12612) );
XOR U21022 ( .A(c4204), .B(b[4204]), .Z(n12613) );
XNOR U21023 ( .A(b[4204]), .B(n12614), .Z(c[4204]) );
XNOR U21024 ( .A(a[4204]), .B(c4204), .Z(n12614) );
XOR U21025 ( .A(c4205), .B(n12615), .Z(c4206) );
ANDN U21026 ( .B(n12616), .A(n12617), .Z(n12615) );
XOR U21027 ( .A(c4205), .B(b[4205]), .Z(n12616) );
XNOR U21028 ( .A(b[4205]), .B(n12617), .Z(c[4205]) );
XNOR U21029 ( .A(a[4205]), .B(c4205), .Z(n12617) );
XOR U21030 ( .A(c4206), .B(n12618), .Z(c4207) );
ANDN U21031 ( .B(n12619), .A(n12620), .Z(n12618) );
XOR U21032 ( .A(c4206), .B(b[4206]), .Z(n12619) );
XNOR U21033 ( .A(b[4206]), .B(n12620), .Z(c[4206]) );
XNOR U21034 ( .A(a[4206]), .B(c4206), .Z(n12620) );
XOR U21035 ( .A(c4207), .B(n12621), .Z(c4208) );
ANDN U21036 ( .B(n12622), .A(n12623), .Z(n12621) );
XOR U21037 ( .A(c4207), .B(b[4207]), .Z(n12622) );
XNOR U21038 ( .A(b[4207]), .B(n12623), .Z(c[4207]) );
XNOR U21039 ( .A(a[4207]), .B(c4207), .Z(n12623) );
XOR U21040 ( .A(c4208), .B(n12624), .Z(c4209) );
ANDN U21041 ( .B(n12625), .A(n12626), .Z(n12624) );
XOR U21042 ( .A(c4208), .B(b[4208]), .Z(n12625) );
XNOR U21043 ( .A(b[4208]), .B(n12626), .Z(c[4208]) );
XNOR U21044 ( .A(a[4208]), .B(c4208), .Z(n12626) );
XOR U21045 ( .A(c4209), .B(n12627), .Z(c4210) );
ANDN U21046 ( .B(n12628), .A(n12629), .Z(n12627) );
XOR U21047 ( .A(c4209), .B(b[4209]), .Z(n12628) );
XNOR U21048 ( .A(b[4209]), .B(n12629), .Z(c[4209]) );
XNOR U21049 ( .A(a[4209]), .B(c4209), .Z(n12629) );
XOR U21050 ( .A(c4210), .B(n12630), .Z(c4211) );
ANDN U21051 ( .B(n12631), .A(n12632), .Z(n12630) );
XOR U21052 ( .A(c4210), .B(b[4210]), .Z(n12631) );
XNOR U21053 ( .A(b[4210]), .B(n12632), .Z(c[4210]) );
XNOR U21054 ( .A(a[4210]), .B(c4210), .Z(n12632) );
XOR U21055 ( .A(c4211), .B(n12633), .Z(c4212) );
ANDN U21056 ( .B(n12634), .A(n12635), .Z(n12633) );
XOR U21057 ( .A(c4211), .B(b[4211]), .Z(n12634) );
XNOR U21058 ( .A(b[4211]), .B(n12635), .Z(c[4211]) );
XNOR U21059 ( .A(a[4211]), .B(c4211), .Z(n12635) );
XOR U21060 ( .A(c4212), .B(n12636), .Z(c4213) );
ANDN U21061 ( .B(n12637), .A(n12638), .Z(n12636) );
XOR U21062 ( .A(c4212), .B(b[4212]), .Z(n12637) );
XNOR U21063 ( .A(b[4212]), .B(n12638), .Z(c[4212]) );
XNOR U21064 ( .A(a[4212]), .B(c4212), .Z(n12638) );
XOR U21065 ( .A(c4213), .B(n12639), .Z(c4214) );
ANDN U21066 ( .B(n12640), .A(n12641), .Z(n12639) );
XOR U21067 ( .A(c4213), .B(b[4213]), .Z(n12640) );
XNOR U21068 ( .A(b[4213]), .B(n12641), .Z(c[4213]) );
XNOR U21069 ( .A(a[4213]), .B(c4213), .Z(n12641) );
XOR U21070 ( .A(c4214), .B(n12642), .Z(c4215) );
ANDN U21071 ( .B(n12643), .A(n12644), .Z(n12642) );
XOR U21072 ( .A(c4214), .B(b[4214]), .Z(n12643) );
XNOR U21073 ( .A(b[4214]), .B(n12644), .Z(c[4214]) );
XNOR U21074 ( .A(a[4214]), .B(c4214), .Z(n12644) );
XOR U21075 ( .A(c4215), .B(n12645), .Z(c4216) );
ANDN U21076 ( .B(n12646), .A(n12647), .Z(n12645) );
XOR U21077 ( .A(c4215), .B(b[4215]), .Z(n12646) );
XNOR U21078 ( .A(b[4215]), .B(n12647), .Z(c[4215]) );
XNOR U21079 ( .A(a[4215]), .B(c4215), .Z(n12647) );
XOR U21080 ( .A(c4216), .B(n12648), .Z(c4217) );
ANDN U21081 ( .B(n12649), .A(n12650), .Z(n12648) );
XOR U21082 ( .A(c4216), .B(b[4216]), .Z(n12649) );
XNOR U21083 ( .A(b[4216]), .B(n12650), .Z(c[4216]) );
XNOR U21084 ( .A(a[4216]), .B(c4216), .Z(n12650) );
XOR U21085 ( .A(c4217), .B(n12651), .Z(c4218) );
ANDN U21086 ( .B(n12652), .A(n12653), .Z(n12651) );
XOR U21087 ( .A(c4217), .B(b[4217]), .Z(n12652) );
XNOR U21088 ( .A(b[4217]), .B(n12653), .Z(c[4217]) );
XNOR U21089 ( .A(a[4217]), .B(c4217), .Z(n12653) );
XOR U21090 ( .A(c4218), .B(n12654), .Z(c4219) );
ANDN U21091 ( .B(n12655), .A(n12656), .Z(n12654) );
XOR U21092 ( .A(c4218), .B(b[4218]), .Z(n12655) );
XNOR U21093 ( .A(b[4218]), .B(n12656), .Z(c[4218]) );
XNOR U21094 ( .A(a[4218]), .B(c4218), .Z(n12656) );
XOR U21095 ( .A(c4219), .B(n12657), .Z(c4220) );
ANDN U21096 ( .B(n12658), .A(n12659), .Z(n12657) );
XOR U21097 ( .A(c4219), .B(b[4219]), .Z(n12658) );
XNOR U21098 ( .A(b[4219]), .B(n12659), .Z(c[4219]) );
XNOR U21099 ( .A(a[4219]), .B(c4219), .Z(n12659) );
XOR U21100 ( .A(c4220), .B(n12660), .Z(c4221) );
ANDN U21101 ( .B(n12661), .A(n12662), .Z(n12660) );
XOR U21102 ( .A(c4220), .B(b[4220]), .Z(n12661) );
XNOR U21103 ( .A(b[4220]), .B(n12662), .Z(c[4220]) );
XNOR U21104 ( .A(a[4220]), .B(c4220), .Z(n12662) );
XOR U21105 ( .A(c4221), .B(n12663), .Z(c4222) );
ANDN U21106 ( .B(n12664), .A(n12665), .Z(n12663) );
XOR U21107 ( .A(c4221), .B(b[4221]), .Z(n12664) );
XNOR U21108 ( .A(b[4221]), .B(n12665), .Z(c[4221]) );
XNOR U21109 ( .A(a[4221]), .B(c4221), .Z(n12665) );
XOR U21110 ( .A(c4222), .B(n12666), .Z(c4223) );
ANDN U21111 ( .B(n12667), .A(n12668), .Z(n12666) );
XOR U21112 ( .A(c4222), .B(b[4222]), .Z(n12667) );
XNOR U21113 ( .A(b[4222]), .B(n12668), .Z(c[4222]) );
XNOR U21114 ( .A(a[4222]), .B(c4222), .Z(n12668) );
XOR U21115 ( .A(c4223), .B(n12669), .Z(c4224) );
ANDN U21116 ( .B(n12670), .A(n12671), .Z(n12669) );
XOR U21117 ( .A(c4223), .B(b[4223]), .Z(n12670) );
XNOR U21118 ( .A(b[4223]), .B(n12671), .Z(c[4223]) );
XNOR U21119 ( .A(a[4223]), .B(c4223), .Z(n12671) );
XOR U21120 ( .A(c4224), .B(n12672), .Z(c4225) );
ANDN U21121 ( .B(n12673), .A(n12674), .Z(n12672) );
XOR U21122 ( .A(c4224), .B(b[4224]), .Z(n12673) );
XNOR U21123 ( .A(b[4224]), .B(n12674), .Z(c[4224]) );
XNOR U21124 ( .A(a[4224]), .B(c4224), .Z(n12674) );
XOR U21125 ( .A(c4225), .B(n12675), .Z(c4226) );
ANDN U21126 ( .B(n12676), .A(n12677), .Z(n12675) );
XOR U21127 ( .A(c4225), .B(b[4225]), .Z(n12676) );
XNOR U21128 ( .A(b[4225]), .B(n12677), .Z(c[4225]) );
XNOR U21129 ( .A(a[4225]), .B(c4225), .Z(n12677) );
XOR U21130 ( .A(c4226), .B(n12678), .Z(c4227) );
ANDN U21131 ( .B(n12679), .A(n12680), .Z(n12678) );
XOR U21132 ( .A(c4226), .B(b[4226]), .Z(n12679) );
XNOR U21133 ( .A(b[4226]), .B(n12680), .Z(c[4226]) );
XNOR U21134 ( .A(a[4226]), .B(c4226), .Z(n12680) );
XOR U21135 ( .A(c4227), .B(n12681), .Z(c4228) );
ANDN U21136 ( .B(n12682), .A(n12683), .Z(n12681) );
XOR U21137 ( .A(c4227), .B(b[4227]), .Z(n12682) );
XNOR U21138 ( .A(b[4227]), .B(n12683), .Z(c[4227]) );
XNOR U21139 ( .A(a[4227]), .B(c4227), .Z(n12683) );
XOR U21140 ( .A(c4228), .B(n12684), .Z(c4229) );
ANDN U21141 ( .B(n12685), .A(n12686), .Z(n12684) );
XOR U21142 ( .A(c4228), .B(b[4228]), .Z(n12685) );
XNOR U21143 ( .A(b[4228]), .B(n12686), .Z(c[4228]) );
XNOR U21144 ( .A(a[4228]), .B(c4228), .Z(n12686) );
XOR U21145 ( .A(c4229), .B(n12687), .Z(c4230) );
ANDN U21146 ( .B(n12688), .A(n12689), .Z(n12687) );
XOR U21147 ( .A(c4229), .B(b[4229]), .Z(n12688) );
XNOR U21148 ( .A(b[4229]), .B(n12689), .Z(c[4229]) );
XNOR U21149 ( .A(a[4229]), .B(c4229), .Z(n12689) );
XOR U21150 ( .A(c4230), .B(n12690), .Z(c4231) );
ANDN U21151 ( .B(n12691), .A(n12692), .Z(n12690) );
XOR U21152 ( .A(c4230), .B(b[4230]), .Z(n12691) );
XNOR U21153 ( .A(b[4230]), .B(n12692), .Z(c[4230]) );
XNOR U21154 ( .A(a[4230]), .B(c4230), .Z(n12692) );
XOR U21155 ( .A(c4231), .B(n12693), .Z(c4232) );
ANDN U21156 ( .B(n12694), .A(n12695), .Z(n12693) );
XOR U21157 ( .A(c4231), .B(b[4231]), .Z(n12694) );
XNOR U21158 ( .A(b[4231]), .B(n12695), .Z(c[4231]) );
XNOR U21159 ( .A(a[4231]), .B(c4231), .Z(n12695) );
XOR U21160 ( .A(c4232), .B(n12696), .Z(c4233) );
ANDN U21161 ( .B(n12697), .A(n12698), .Z(n12696) );
XOR U21162 ( .A(c4232), .B(b[4232]), .Z(n12697) );
XNOR U21163 ( .A(b[4232]), .B(n12698), .Z(c[4232]) );
XNOR U21164 ( .A(a[4232]), .B(c4232), .Z(n12698) );
XOR U21165 ( .A(c4233), .B(n12699), .Z(c4234) );
ANDN U21166 ( .B(n12700), .A(n12701), .Z(n12699) );
XOR U21167 ( .A(c4233), .B(b[4233]), .Z(n12700) );
XNOR U21168 ( .A(b[4233]), .B(n12701), .Z(c[4233]) );
XNOR U21169 ( .A(a[4233]), .B(c4233), .Z(n12701) );
XOR U21170 ( .A(c4234), .B(n12702), .Z(c4235) );
ANDN U21171 ( .B(n12703), .A(n12704), .Z(n12702) );
XOR U21172 ( .A(c4234), .B(b[4234]), .Z(n12703) );
XNOR U21173 ( .A(b[4234]), .B(n12704), .Z(c[4234]) );
XNOR U21174 ( .A(a[4234]), .B(c4234), .Z(n12704) );
XOR U21175 ( .A(c4235), .B(n12705), .Z(c4236) );
ANDN U21176 ( .B(n12706), .A(n12707), .Z(n12705) );
XOR U21177 ( .A(c4235), .B(b[4235]), .Z(n12706) );
XNOR U21178 ( .A(b[4235]), .B(n12707), .Z(c[4235]) );
XNOR U21179 ( .A(a[4235]), .B(c4235), .Z(n12707) );
XOR U21180 ( .A(c4236), .B(n12708), .Z(c4237) );
ANDN U21181 ( .B(n12709), .A(n12710), .Z(n12708) );
XOR U21182 ( .A(c4236), .B(b[4236]), .Z(n12709) );
XNOR U21183 ( .A(b[4236]), .B(n12710), .Z(c[4236]) );
XNOR U21184 ( .A(a[4236]), .B(c4236), .Z(n12710) );
XOR U21185 ( .A(c4237), .B(n12711), .Z(c4238) );
ANDN U21186 ( .B(n12712), .A(n12713), .Z(n12711) );
XOR U21187 ( .A(c4237), .B(b[4237]), .Z(n12712) );
XNOR U21188 ( .A(b[4237]), .B(n12713), .Z(c[4237]) );
XNOR U21189 ( .A(a[4237]), .B(c4237), .Z(n12713) );
XOR U21190 ( .A(c4238), .B(n12714), .Z(c4239) );
ANDN U21191 ( .B(n12715), .A(n12716), .Z(n12714) );
XOR U21192 ( .A(c4238), .B(b[4238]), .Z(n12715) );
XNOR U21193 ( .A(b[4238]), .B(n12716), .Z(c[4238]) );
XNOR U21194 ( .A(a[4238]), .B(c4238), .Z(n12716) );
XOR U21195 ( .A(c4239), .B(n12717), .Z(c4240) );
ANDN U21196 ( .B(n12718), .A(n12719), .Z(n12717) );
XOR U21197 ( .A(c4239), .B(b[4239]), .Z(n12718) );
XNOR U21198 ( .A(b[4239]), .B(n12719), .Z(c[4239]) );
XNOR U21199 ( .A(a[4239]), .B(c4239), .Z(n12719) );
XOR U21200 ( .A(c4240), .B(n12720), .Z(c4241) );
ANDN U21201 ( .B(n12721), .A(n12722), .Z(n12720) );
XOR U21202 ( .A(c4240), .B(b[4240]), .Z(n12721) );
XNOR U21203 ( .A(b[4240]), .B(n12722), .Z(c[4240]) );
XNOR U21204 ( .A(a[4240]), .B(c4240), .Z(n12722) );
XOR U21205 ( .A(c4241), .B(n12723), .Z(c4242) );
ANDN U21206 ( .B(n12724), .A(n12725), .Z(n12723) );
XOR U21207 ( .A(c4241), .B(b[4241]), .Z(n12724) );
XNOR U21208 ( .A(b[4241]), .B(n12725), .Z(c[4241]) );
XNOR U21209 ( .A(a[4241]), .B(c4241), .Z(n12725) );
XOR U21210 ( .A(c4242), .B(n12726), .Z(c4243) );
ANDN U21211 ( .B(n12727), .A(n12728), .Z(n12726) );
XOR U21212 ( .A(c4242), .B(b[4242]), .Z(n12727) );
XNOR U21213 ( .A(b[4242]), .B(n12728), .Z(c[4242]) );
XNOR U21214 ( .A(a[4242]), .B(c4242), .Z(n12728) );
XOR U21215 ( .A(c4243), .B(n12729), .Z(c4244) );
ANDN U21216 ( .B(n12730), .A(n12731), .Z(n12729) );
XOR U21217 ( .A(c4243), .B(b[4243]), .Z(n12730) );
XNOR U21218 ( .A(b[4243]), .B(n12731), .Z(c[4243]) );
XNOR U21219 ( .A(a[4243]), .B(c4243), .Z(n12731) );
XOR U21220 ( .A(c4244), .B(n12732), .Z(c4245) );
ANDN U21221 ( .B(n12733), .A(n12734), .Z(n12732) );
XOR U21222 ( .A(c4244), .B(b[4244]), .Z(n12733) );
XNOR U21223 ( .A(b[4244]), .B(n12734), .Z(c[4244]) );
XNOR U21224 ( .A(a[4244]), .B(c4244), .Z(n12734) );
XOR U21225 ( .A(c4245), .B(n12735), .Z(c4246) );
ANDN U21226 ( .B(n12736), .A(n12737), .Z(n12735) );
XOR U21227 ( .A(c4245), .B(b[4245]), .Z(n12736) );
XNOR U21228 ( .A(b[4245]), .B(n12737), .Z(c[4245]) );
XNOR U21229 ( .A(a[4245]), .B(c4245), .Z(n12737) );
XOR U21230 ( .A(c4246), .B(n12738), .Z(c4247) );
ANDN U21231 ( .B(n12739), .A(n12740), .Z(n12738) );
XOR U21232 ( .A(c4246), .B(b[4246]), .Z(n12739) );
XNOR U21233 ( .A(b[4246]), .B(n12740), .Z(c[4246]) );
XNOR U21234 ( .A(a[4246]), .B(c4246), .Z(n12740) );
XOR U21235 ( .A(c4247), .B(n12741), .Z(c4248) );
ANDN U21236 ( .B(n12742), .A(n12743), .Z(n12741) );
XOR U21237 ( .A(c4247), .B(b[4247]), .Z(n12742) );
XNOR U21238 ( .A(b[4247]), .B(n12743), .Z(c[4247]) );
XNOR U21239 ( .A(a[4247]), .B(c4247), .Z(n12743) );
XOR U21240 ( .A(c4248), .B(n12744), .Z(c4249) );
ANDN U21241 ( .B(n12745), .A(n12746), .Z(n12744) );
XOR U21242 ( .A(c4248), .B(b[4248]), .Z(n12745) );
XNOR U21243 ( .A(b[4248]), .B(n12746), .Z(c[4248]) );
XNOR U21244 ( .A(a[4248]), .B(c4248), .Z(n12746) );
XOR U21245 ( .A(c4249), .B(n12747), .Z(c4250) );
ANDN U21246 ( .B(n12748), .A(n12749), .Z(n12747) );
XOR U21247 ( .A(c4249), .B(b[4249]), .Z(n12748) );
XNOR U21248 ( .A(b[4249]), .B(n12749), .Z(c[4249]) );
XNOR U21249 ( .A(a[4249]), .B(c4249), .Z(n12749) );
XOR U21250 ( .A(c4250), .B(n12750), .Z(c4251) );
ANDN U21251 ( .B(n12751), .A(n12752), .Z(n12750) );
XOR U21252 ( .A(c4250), .B(b[4250]), .Z(n12751) );
XNOR U21253 ( .A(b[4250]), .B(n12752), .Z(c[4250]) );
XNOR U21254 ( .A(a[4250]), .B(c4250), .Z(n12752) );
XOR U21255 ( .A(c4251), .B(n12753), .Z(c4252) );
ANDN U21256 ( .B(n12754), .A(n12755), .Z(n12753) );
XOR U21257 ( .A(c4251), .B(b[4251]), .Z(n12754) );
XNOR U21258 ( .A(b[4251]), .B(n12755), .Z(c[4251]) );
XNOR U21259 ( .A(a[4251]), .B(c4251), .Z(n12755) );
XOR U21260 ( .A(c4252), .B(n12756), .Z(c4253) );
ANDN U21261 ( .B(n12757), .A(n12758), .Z(n12756) );
XOR U21262 ( .A(c4252), .B(b[4252]), .Z(n12757) );
XNOR U21263 ( .A(b[4252]), .B(n12758), .Z(c[4252]) );
XNOR U21264 ( .A(a[4252]), .B(c4252), .Z(n12758) );
XOR U21265 ( .A(c4253), .B(n12759), .Z(c4254) );
ANDN U21266 ( .B(n12760), .A(n12761), .Z(n12759) );
XOR U21267 ( .A(c4253), .B(b[4253]), .Z(n12760) );
XNOR U21268 ( .A(b[4253]), .B(n12761), .Z(c[4253]) );
XNOR U21269 ( .A(a[4253]), .B(c4253), .Z(n12761) );
XOR U21270 ( .A(c4254), .B(n12762), .Z(c4255) );
ANDN U21271 ( .B(n12763), .A(n12764), .Z(n12762) );
XOR U21272 ( .A(c4254), .B(b[4254]), .Z(n12763) );
XNOR U21273 ( .A(b[4254]), .B(n12764), .Z(c[4254]) );
XNOR U21274 ( .A(a[4254]), .B(c4254), .Z(n12764) );
XOR U21275 ( .A(c4255), .B(n12765), .Z(c4256) );
ANDN U21276 ( .B(n12766), .A(n12767), .Z(n12765) );
XOR U21277 ( .A(c4255), .B(b[4255]), .Z(n12766) );
XNOR U21278 ( .A(b[4255]), .B(n12767), .Z(c[4255]) );
XNOR U21279 ( .A(a[4255]), .B(c4255), .Z(n12767) );
XOR U21280 ( .A(c4256), .B(n12768), .Z(c4257) );
ANDN U21281 ( .B(n12769), .A(n12770), .Z(n12768) );
XOR U21282 ( .A(c4256), .B(b[4256]), .Z(n12769) );
XNOR U21283 ( .A(b[4256]), .B(n12770), .Z(c[4256]) );
XNOR U21284 ( .A(a[4256]), .B(c4256), .Z(n12770) );
XOR U21285 ( .A(c4257), .B(n12771), .Z(c4258) );
ANDN U21286 ( .B(n12772), .A(n12773), .Z(n12771) );
XOR U21287 ( .A(c4257), .B(b[4257]), .Z(n12772) );
XNOR U21288 ( .A(b[4257]), .B(n12773), .Z(c[4257]) );
XNOR U21289 ( .A(a[4257]), .B(c4257), .Z(n12773) );
XOR U21290 ( .A(c4258), .B(n12774), .Z(c4259) );
ANDN U21291 ( .B(n12775), .A(n12776), .Z(n12774) );
XOR U21292 ( .A(c4258), .B(b[4258]), .Z(n12775) );
XNOR U21293 ( .A(b[4258]), .B(n12776), .Z(c[4258]) );
XNOR U21294 ( .A(a[4258]), .B(c4258), .Z(n12776) );
XOR U21295 ( .A(c4259), .B(n12777), .Z(c4260) );
ANDN U21296 ( .B(n12778), .A(n12779), .Z(n12777) );
XOR U21297 ( .A(c4259), .B(b[4259]), .Z(n12778) );
XNOR U21298 ( .A(b[4259]), .B(n12779), .Z(c[4259]) );
XNOR U21299 ( .A(a[4259]), .B(c4259), .Z(n12779) );
XOR U21300 ( .A(c4260), .B(n12780), .Z(c4261) );
ANDN U21301 ( .B(n12781), .A(n12782), .Z(n12780) );
XOR U21302 ( .A(c4260), .B(b[4260]), .Z(n12781) );
XNOR U21303 ( .A(b[4260]), .B(n12782), .Z(c[4260]) );
XNOR U21304 ( .A(a[4260]), .B(c4260), .Z(n12782) );
XOR U21305 ( .A(c4261), .B(n12783), .Z(c4262) );
ANDN U21306 ( .B(n12784), .A(n12785), .Z(n12783) );
XOR U21307 ( .A(c4261), .B(b[4261]), .Z(n12784) );
XNOR U21308 ( .A(b[4261]), .B(n12785), .Z(c[4261]) );
XNOR U21309 ( .A(a[4261]), .B(c4261), .Z(n12785) );
XOR U21310 ( .A(c4262), .B(n12786), .Z(c4263) );
ANDN U21311 ( .B(n12787), .A(n12788), .Z(n12786) );
XOR U21312 ( .A(c4262), .B(b[4262]), .Z(n12787) );
XNOR U21313 ( .A(b[4262]), .B(n12788), .Z(c[4262]) );
XNOR U21314 ( .A(a[4262]), .B(c4262), .Z(n12788) );
XOR U21315 ( .A(c4263), .B(n12789), .Z(c4264) );
ANDN U21316 ( .B(n12790), .A(n12791), .Z(n12789) );
XOR U21317 ( .A(c4263), .B(b[4263]), .Z(n12790) );
XNOR U21318 ( .A(b[4263]), .B(n12791), .Z(c[4263]) );
XNOR U21319 ( .A(a[4263]), .B(c4263), .Z(n12791) );
XOR U21320 ( .A(c4264), .B(n12792), .Z(c4265) );
ANDN U21321 ( .B(n12793), .A(n12794), .Z(n12792) );
XOR U21322 ( .A(c4264), .B(b[4264]), .Z(n12793) );
XNOR U21323 ( .A(b[4264]), .B(n12794), .Z(c[4264]) );
XNOR U21324 ( .A(a[4264]), .B(c4264), .Z(n12794) );
XOR U21325 ( .A(c4265), .B(n12795), .Z(c4266) );
ANDN U21326 ( .B(n12796), .A(n12797), .Z(n12795) );
XOR U21327 ( .A(c4265), .B(b[4265]), .Z(n12796) );
XNOR U21328 ( .A(b[4265]), .B(n12797), .Z(c[4265]) );
XNOR U21329 ( .A(a[4265]), .B(c4265), .Z(n12797) );
XOR U21330 ( .A(c4266), .B(n12798), .Z(c4267) );
ANDN U21331 ( .B(n12799), .A(n12800), .Z(n12798) );
XOR U21332 ( .A(c4266), .B(b[4266]), .Z(n12799) );
XNOR U21333 ( .A(b[4266]), .B(n12800), .Z(c[4266]) );
XNOR U21334 ( .A(a[4266]), .B(c4266), .Z(n12800) );
XOR U21335 ( .A(c4267), .B(n12801), .Z(c4268) );
ANDN U21336 ( .B(n12802), .A(n12803), .Z(n12801) );
XOR U21337 ( .A(c4267), .B(b[4267]), .Z(n12802) );
XNOR U21338 ( .A(b[4267]), .B(n12803), .Z(c[4267]) );
XNOR U21339 ( .A(a[4267]), .B(c4267), .Z(n12803) );
XOR U21340 ( .A(c4268), .B(n12804), .Z(c4269) );
ANDN U21341 ( .B(n12805), .A(n12806), .Z(n12804) );
XOR U21342 ( .A(c4268), .B(b[4268]), .Z(n12805) );
XNOR U21343 ( .A(b[4268]), .B(n12806), .Z(c[4268]) );
XNOR U21344 ( .A(a[4268]), .B(c4268), .Z(n12806) );
XOR U21345 ( .A(c4269), .B(n12807), .Z(c4270) );
ANDN U21346 ( .B(n12808), .A(n12809), .Z(n12807) );
XOR U21347 ( .A(c4269), .B(b[4269]), .Z(n12808) );
XNOR U21348 ( .A(b[4269]), .B(n12809), .Z(c[4269]) );
XNOR U21349 ( .A(a[4269]), .B(c4269), .Z(n12809) );
XOR U21350 ( .A(c4270), .B(n12810), .Z(c4271) );
ANDN U21351 ( .B(n12811), .A(n12812), .Z(n12810) );
XOR U21352 ( .A(c4270), .B(b[4270]), .Z(n12811) );
XNOR U21353 ( .A(b[4270]), .B(n12812), .Z(c[4270]) );
XNOR U21354 ( .A(a[4270]), .B(c4270), .Z(n12812) );
XOR U21355 ( .A(c4271), .B(n12813), .Z(c4272) );
ANDN U21356 ( .B(n12814), .A(n12815), .Z(n12813) );
XOR U21357 ( .A(c4271), .B(b[4271]), .Z(n12814) );
XNOR U21358 ( .A(b[4271]), .B(n12815), .Z(c[4271]) );
XNOR U21359 ( .A(a[4271]), .B(c4271), .Z(n12815) );
XOR U21360 ( .A(c4272), .B(n12816), .Z(c4273) );
ANDN U21361 ( .B(n12817), .A(n12818), .Z(n12816) );
XOR U21362 ( .A(c4272), .B(b[4272]), .Z(n12817) );
XNOR U21363 ( .A(b[4272]), .B(n12818), .Z(c[4272]) );
XNOR U21364 ( .A(a[4272]), .B(c4272), .Z(n12818) );
XOR U21365 ( .A(c4273), .B(n12819), .Z(c4274) );
ANDN U21366 ( .B(n12820), .A(n12821), .Z(n12819) );
XOR U21367 ( .A(c4273), .B(b[4273]), .Z(n12820) );
XNOR U21368 ( .A(b[4273]), .B(n12821), .Z(c[4273]) );
XNOR U21369 ( .A(a[4273]), .B(c4273), .Z(n12821) );
XOR U21370 ( .A(c4274), .B(n12822), .Z(c4275) );
ANDN U21371 ( .B(n12823), .A(n12824), .Z(n12822) );
XOR U21372 ( .A(c4274), .B(b[4274]), .Z(n12823) );
XNOR U21373 ( .A(b[4274]), .B(n12824), .Z(c[4274]) );
XNOR U21374 ( .A(a[4274]), .B(c4274), .Z(n12824) );
XOR U21375 ( .A(c4275), .B(n12825), .Z(c4276) );
ANDN U21376 ( .B(n12826), .A(n12827), .Z(n12825) );
XOR U21377 ( .A(c4275), .B(b[4275]), .Z(n12826) );
XNOR U21378 ( .A(b[4275]), .B(n12827), .Z(c[4275]) );
XNOR U21379 ( .A(a[4275]), .B(c4275), .Z(n12827) );
XOR U21380 ( .A(c4276), .B(n12828), .Z(c4277) );
ANDN U21381 ( .B(n12829), .A(n12830), .Z(n12828) );
XOR U21382 ( .A(c4276), .B(b[4276]), .Z(n12829) );
XNOR U21383 ( .A(b[4276]), .B(n12830), .Z(c[4276]) );
XNOR U21384 ( .A(a[4276]), .B(c4276), .Z(n12830) );
XOR U21385 ( .A(c4277), .B(n12831), .Z(c4278) );
ANDN U21386 ( .B(n12832), .A(n12833), .Z(n12831) );
XOR U21387 ( .A(c4277), .B(b[4277]), .Z(n12832) );
XNOR U21388 ( .A(b[4277]), .B(n12833), .Z(c[4277]) );
XNOR U21389 ( .A(a[4277]), .B(c4277), .Z(n12833) );
XOR U21390 ( .A(c4278), .B(n12834), .Z(c4279) );
ANDN U21391 ( .B(n12835), .A(n12836), .Z(n12834) );
XOR U21392 ( .A(c4278), .B(b[4278]), .Z(n12835) );
XNOR U21393 ( .A(b[4278]), .B(n12836), .Z(c[4278]) );
XNOR U21394 ( .A(a[4278]), .B(c4278), .Z(n12836) );
XOR U21395 ( .A(c4279), .B(n12837), .Z(c4280) );
ANDN U21396 ( .B(n12838), .A(n12839), .Z(n12837) );
XOR U21397 ( .A(c4279), .B(b[4279]), .Z(n12838) );
XNOR U21398 ( .A(b[4279]), .B(n12839), .Z(c[4279]) );
XNOR U21399 ( .A(a[4279]), .B(c4279), .Z(n12839) );
XOR U21400 ( .A(c4280), .B(n12840), .Z(c4281) );
ANDN U21401 ( .B(n12841), .A(n12842), .Z(n12840) );
XOR U21402 ( .A(c4280), .B(b[4280]), .Z(n12841) );
XNOR U21403 ( .A(b[4280]), .B(n12842), .Z(c[4280]) );
XNOR U21404 ( .A(a[4280]), .B(c4280), .Z(n12842) );
XOR U21405 ( .A(c4281), .B(n12843), .Z(c4282) );
ANDN U21406 ( .B(n12844), .A(n12845), .Z(n12843) );
XOR U21407 ( .A(c4281), .B(b[4281]), .Z(n12844) );
XNOR U21408 ( .A(b[4281]), .B(n12845), .Z(c[4281]) );
XNOR U21409 ( .A(a[4281]), .B(c4281), .Z(n12845) );
XOR U21410 ( .A(c4282), .B(n12846), .Z(c4283) );
ANDN U21411 ( .B(n12847), .A(n12848), .Z(n12846) );
XOR U21412 ( .A(c4282), .B(b[4282]), .Z(n12847) );
XNOR U21413 ( .A(b[4282]), .B(n12848), .Z(c[4282]) );
XNOR U21414 ( .A(a[4282]), .B(c4282), .Z(n12848) );
XOR U21415 ( .A(c4283), .B(n12849), .Z(c4284) );
ANDN U21416 ( .B(n12850), .A(n12851), .Z(n12849) );
XOR U21417 ( .A(c4283), .B(b[4283]), .Z(n12850) );
XNOR U21418 ( .A(b[4283]), .B(n12851), .Z(c[4283]) );
XNOR U21419 ( .A(a[4283]), .B(c4283), .Z(n12851) );
XOR U21420 ( .A(c4284), .B(n12852), .Z(c4285) );
ANDN U21421 ( .B(n12853), .A(n12854), .Z(n12852) );
XOR U21422 ( .A(c4284), .B(b[4284]), .Z(n12853) );
XNOR U21423 ( .A(b[4284]), .B(n12854), .Z(c[4284]) );
XNOR U21424 ( .A(a[4284]), .B(c4284), .Z(n12854) );
XOR U21425 ( .A(c4285), .B(n12855), .Z(c4286) );
ANDN U21426 ( .B(n12856), .A(n12857), .Z(n12855) );
XOR U21427 ( .A(c4285), .B(b[4285]), .Z(n12856) );
XNOR U21428 ( .A(b[4285]), .B(n12857), .Z(c[4285]) );
XNOR U21429 ( .A(a[4285]), .B(c4285), .Z(n12857) );
XOR U21430 ( .A(c4286), .B(n12858), .Z(c4287) );
ANDN U21431 ( .B(n12859), .A(n12860), .Z(n12858) );
XOR U21432 ( .A(c4286), .B(b[4286]), .Z(n12859) );
XNOR U21433 ( .A(b[4286]), .B(n12860), .Z(c[4286]) );
XNOR U21434 ( .A(a[4286]), .B(c4286), .Z(n12860) );
XOR U21435 ( .A(c4287), .B(n12861), .Z(c4288) );
ANDN U21436 ( .B(n12862), .A(n12863), .Z(n12861) );
XOR U21437 ( .A(c4287), .B(b[4287]), .Z(n12862) );
XNOR U21438 ( .A(b[4287]), .B(n12863), .Z(c[4287]) );
XNOR U21439 ( .A(a[4287]), .B(c4287), .Z(n12863) );
XOR U21440 ( .A(c4288), .B(n12864), .Z(c4289) );
ANDN U21441 ( .B(n12865), .A(n12866), .Z(n12864) );
XOR U21442 ( .A(c4288), .B(b[4288]), .Z(n12865) );
XNOR U21443 ( .A(b[4288]), .B(n12866), .Z(c[4288]) );
XNOR U21444 ( .A(a[4288]), .B(c4288), .Z(n12866) );
XOR U21445 ( .A(c4289), .B(n12867), .Z(c4290) );
ANDN U21446 ( .B(n12868), .A(n12869), .Z(n12867) );
XOR U21447 ( .A(c4289), .B(b[4289]), .Z(n12868) );
XNOR U21448 ( .A(b[4289]), .B(n12869), .Z(c[4289]) );
XNOR U21449 ( .A(a[4289]), .B(c4289), .Z(n12869) );
XOR U21450 ( .A(c4290), .B(n12870), .Z(c4291) );
ANDN U21451 ( .B(n12871), .A(n12872), .Z(n12870) );
XOR U21452 ( .A(c4290), .B(b[4290]), .Z(n12871) );
XNOR U21453 ( .A(b[4290]), .B(n12872), .Z(c[4290]) );
XNOR U21454 ( .A(a[4290]), .B(c4290), .Z(n12872) );
XOR U21455 ( .A(c4291), .B(n12873), .Z(c4292) );
ANDN U21456 ( .B(n12874), .A(n12875), .Z(n12873) );
XOR U21457 ( .A(c4291), .B(b[4291]), .Z(n12874) );
XNOR U21458 ( .A(b[4291]), .B(n12875), .Z(c[4291]) );
XNOR U21459 ( .A(a[4291]), .B(c4291), .Z(n12875) );
XOR U21460 ( .A(c4292), .B(n12876), .Z(c4293) );
ANDN U21461 ( .B(n12877), .A(n12878), .Z(n12876) );
XOR U21462 ( .A(c4292), .B(b[4292]), .Z(n12877) );
XNOR U21463 ( .A(b[4292]), .B(n12878), .Z(c[4292]) );
XNOR U21464 ( .A(a[4292]), .B(c4292), .Z(n12878) );
XOR U21465 ( .A(c4293), .B(n12879), .Z(c4294) );
ANDN U21466 ( .B(n12880), .A(n12881), .Z(n12879) );
XOR U21467 ( .A(c4293), .B(b[4293]), .Z(n12880) );
XNOR U21468 ( .A(b[4293]), .B(n12881), .Z(c[4293]) );
XNOR U21469 ( .A(a[4293]), .B(c4293), .Z(n12881) );
XOR U21470 ( .A(c4294), .B(n12882), .Z(c4295) );
ANDN U21471 ( .B(n12883), .A(n12884), .Z(n12882) );
XOR U21472 ( .A(c4294), .B(b[4294]), .Z(n12883) );
XNOR U21473 ( .A(b[4294]), .B(n12884), .Z(c[4294]) );
XNOR U21474 ( .A(a[4294]), .B(c4294), .Z(n12884) );
XOR U21475 ( .A(c4295), .B(n12885), .Z(c4296) );
ANDN U21476 ( .B(n12886), .A(n12887), .Z(n12885) );
XOR U21477 ( .A(c4295), .B(b[4295]), .Z(n12886) );
XNOR U21478 ( .A(b[4295]), .B(n12887), .Z(c[4295]) );
XNOR U21479 ( .A(a[4295]), .B(c4295), .Z(n12887) );
XOR U21480 ( .A(c4296), .B(n12888), .Z(c4297) );
ANDN U21481 ( .B(n12889), .A(n12890), .Z(n12888) );
XOR U21482 ( .A(c4296), .B(b[4296]), .Z(n12889) );
XNOR U21483 ( .A(b[4296]), .B(n12890), .Z(c[4296]) );
XNOR U21484 ( .A(a[4296]), .B(c4296), .Z(n12890) );
XOR U21485 ( .A(c4297), .B(n12891), .Z(c4298) );
ANDN U21486 ( .B(n12892), .A(n12893), .Z(n12891) );
XOR U21487 ( .A(c4297), .B(b[4297]), .Z(n12892) );
XNOR U21488 ( .A(b[4297]), .B(n12893), .Z(c[4297]) );
XNOR U21489 ( .A(a[4297]), .B(c4297), .Z(n12893) );
XOR U21490 ( .A(c4298), .B(n12894), .Z(c4299) );
ANDN U21491 ( .B(n12895), .A(n12896), .Z(n12894) );
XOR U21492 ( .A(c4298), .B(b[4298]), .Z(n12895) );
XNOR U21493 ( .A(b[4298]), .B(n12896), .Z(c[4298]) );
XNOR U21494 ( .A(a[4298]), .B(c4298), .Z(n12896) );
XOR U21495 ( .A(c4299), .B(n12897), .Z(c4300) );
ANDN U21496 ( .B(n12898), .A(n12899), .Z(n12897) );
XOR U21497 ( .A(c4299), .B(b[4299]), .Z(n12898) );
XNOR U21498 ( .A(b[4299]), .B(n12899), .Z(c[4299]) );
XNOR U21499 ( .A(a[4299]), .B(c4299), .Z(n12899) );
XOR U21500 ( .A(c4300), .B(n12900), .Z(c4301) );
ANDN U21501 ( .B(n12901), .A(n12902), .Z(n12900) );
XOR U21502 ( .A(c4300), .B(b[4300]), .Z(n12901) );
XNOR U21503 ( .A(b[4300]), .B(n12902), .Z(c[4300]) );
XNOR U21504 ( .A(a[4300]), .B(c4300), .Z(n12902) );
XOR U21505 ( .A(c4301), .B(n12903), .Z(c4302) );
ANDN U21506 ( .B(n12904), .A(n12905), .Z(n12903) );
XOR U21507 ( .A(c4301), .B(b[4301]), .Z(n12904) );
XNOR U21508 ( .A(b[4301]), .B(n12905), .Z(c[4301]) );
XNOR U21509 ( .A(a[4301]), .B(c4301), .Z(n12905) );
XOR U21510 ( .A(c4302), .B(n12906), .Z(c4303) );
ANDN U21511 ( .B(n12907), .A(n12908), .Z(n12906) );
XOR U21512 ( .A(c4302), .B(b[4302]), .Z(n12907) );
XNOR U21513 ( .A(b[4302]), .B(n12908), .Z(c[4302]) );
XNOR U21514 ( .A(a[4302]), .B(c4302), .Z(n12908) );
XOR U21515 ( .A(c4303), .B(n12909), .Z(c4304) );
ANDN U21516 ( .B(n12910), .A(n12911), .Z(n12909) );
XOR U21517 ( .A(c4303), .B(b[4303]), .Z(n12910) );
XNOR U21518 ( .A(b[4303]), .B(n12911), .Z(c[4303]) );
XNOR U21519 ( .A(a[4303]), .B(c4303), .Z(n12911) );
XOR U21520 ( .A(c4304), .B(n12912), .Z(c4305) );
ANDN U21521 ( .B(n12913), .A(n12914), .Z(n12912) );
XOR U21522 ( .A(c4304), .B(b[4304]), .Z(n12913) );
XNOR U21523 ( .A(b[4304]), .B(n12914), .Z(c[4304]) );
XNOR U21524 ( .A(a[4304]), .B(c4304), .Z(n12914) );
XOR U21525 ( .A(c4305), .B(n12915), .Z(c4306) );
ANDN U21526 ( .B(n12916), .A(n12917), .Z(n12915) );
XOR U21527 ( .A(c4305), .B(b[4305]), .Z(n12916) );
XNOR U21528 ( .A(b[4305]), .B(n12917), .Z(c[4305]) );
XNOR U21529 ( .A(a[4305]), .B(c4305), .Z(n12917) );
XOR U21530 ( .A(c4306), .B(n12918), .Z(c4307) );
ANDN U21531 ( .B(n12919), .A(n12920), .Z(n12918) );
XOR U21532 ( .A(c4306), .B(b[4306]), .Z(n12919) );
XNOR U21533 ( .A(b[4306]), .B(n12920), .Z(c[4306]) );
XNOR U21534 ( .A(a[4306]), .B(c4306), .Z(n12920) );
XOR U21535 ( .A(c4307), .B(n12921), .Z(c4308) );
ANDN U21536 ( .B(n12922), .A(n12923), .Z(n12921) );
XOR U21537 ( .A(c4307), .B(b[4307]), .Z(n12922) );
XNOR U21538 ( .A(b[4307]), .B(n12923), .Z(c[4307]) );
XNOR U21539 ( .A(a[4307]), .B(c4307), .Z(n12923) );
XOR U21540 ( .A(c4308), .B(n12924), .Z(c4309) );
ANDN U21541 ( .B(n12925), .A(n12926), .Z(n12924) );
XOR U21542 ( .A(c4308), .B(b[4308]), .Z(n12925) );
XNOR U21543 ( .A(b[4308]), .B(n12926), .Z(c[4308]) );
XNOR U21544 ( .A(a[4308]), .B(c4308), .Z(n12926) );
XOR U21545 ( .A(c4309), .B(n12927), .Z(c4310) );
ANDN U21546 ( .B(n12928), .A(n12929), .Z(n12927) );
XOR U21547 ( .A(c4309), .B(b[4309]), .Z(n12928) );
XNOR U21548 ( .A(b[4309]), .B(n12929), .Z(c[4309]) );
XNOR U21549 ( .A(a[4309]), .B(c4309), .Z(n12929) );
XOR U21550 ( .A(c4310), .B(n12930), .Z(c4311) );
ANDN U21551 ( .B(n12931), .A(n12932), .Z(n12930) );
XOR U21552 ( .A(c4310), .B(b[4310]), .Z(n12931) );
XNOR U21553 ( .A(b[4310]), .B(n12932), .Z(c[4310]) );
XNOR U21554 ( .A(a[4310]), .B(c4310), .Z(n12932) );
XOR U21555 ( .A(c4311), .B(n12933), .Z(c4312) );
ANDN U21556 ( .B(n12934), .A(n12935), .Z(n12933) );
XOR U21557 ( .A(c4311), .B(b[4311]), .Z(n12934) );
XNOR U21558 ( .A(b[4311]), .B(n12935), .Z(c[4311]) );
XNOR U21559 ( .A(a[4311]), .B(c4311), .Z(n12935) );
XOR U21560 ( .A(c4312), .B(n12936), .Z(c4313) );
ANDN U21561 ( .B(n12937), .A(n12938), .Z(n12936) );
XOR U21562 ( .A(c4312), .B(b[4312]), .Z(n12937) );
XNOR U21563 ( .A(b[4312]), .B(n12938), .Z(c[4312]) );
XNOR U21564 ( .A(a[4312]), .B(c4312), .Z(n12938) );
XOR U21565 ( .A(c4313), .B(n12939), .Z(c4314) );
ANDN U21566 ( .B(n12940), .A(n12941), .Z(n12939) );
XOR U21567 ( .A(c4313), .B(b[4313]), .Z(n12940) );
XNOR U21568 ( .A(b[4313]), .B(n12941), .Z(c[4313]) );
XNOR U21569 ( .A(a[4313]), .B(c4313), .Z(n12941) );
XOR U21570 ( .A(c4314), .B(n12942), .Z(c4315) );
ANDN U21571 ( .B(n12943), .A(n12944), .Z(n12942) );
XOR U21572 ( .A(c4314), .B(b[4314]), .Z(n12943) );
XNOR U21573 ( .A(b[4314]), .B(n12944), .Z(c[4314]) );
XNOR U21574 ( .A(a[4314]), .B(c4314), .Z(n12944) );
XOR U21575 ( .A(c4315), .B(n12945), .Z(c4316) );
ANDN U21576 ( .B(n12946), .A(n12947), .Z(n12945) );
XOR U21577 ( .A(c4315), .B(b[4315]), .Z(n12946) );
XNOR U21578 ( .A(b[4315]), .B(n12947), .Z(c[4315]) );
XNOR U21579 ( .A(a[4315]), .B(c4315), .Z(n12947) );
XOR U21580 ( .A(c4316), .B(n12948), .Z(c4317) );
ANDN U21581 ( .B(n12949), .A(n12950), .Z(n12948) );
XOR U21582 ( .A(c4316), .B(b[4316]), .Z(n12949) );
XNOR U21583 ( .A(b[4316]), .B(n12950), .Z(c[4316]) );
XNOR U21584 ( .A(a[4316]), .B(c4316), .Z(n12950) );
XOR U21585 ( .A(c4317), .B(n12951), .Z(c4318) );
ANDN U21586 ( .B(n12952), .A(n12953), .Z(n12951) );
XOR U21587 ( .A(c4317), .B(b[4317]), .Z(n12952) );
XNOR U21588 ( .A(b[4317]), .B(n12953), .Z(c[4317]) );
XNOR U21589 ( .A(a[4317]), .B(c4317), .Z(n12953) );
XOR U21590 ( .A(c4318), .B(n12954), .Z(c4319) );
ANDN U21591 ( .B(n12955), .A(n12956), .Z(n12954) );
XOR U21592 ( .A(c4318), .B(b[4318]), .Z(n12955) );
XNOR U21593 ( .A(b[4318]), .B(n12956), .Z(c[4318]) );
XNOR U21594 ( .A(a[4318]), .B(c4318), .Z(n12956) );
XOR U21595 ( .A(c4319), .B(n12957), .Z(c4320) );
ANDN U21596 ( .B(n12958), .A(n12959), .Z(n12957) );
XOR U21597 ( .A(c4319), .B(b[4319]), .Z(n12958) );
XNOR U21598 ( .A(b[4319]), .B(n12959), .Z(c[4319]) );
XNOR U21599 ( .A(a[4319]), .B(c4319), .Z(n12959) );
XOR U21600 ( .A(c4320), .B(n12960), .Z(c4321) );
ANDN U21601 ( .B(n12961), .A(n12962), .Z(n12960) );
XOR U21602 ( .A(c4320), .B(b[4320]), .Z(n12961) );
XNOR U21603 ( .A(b[4320]), .B(n12962), .Z(c[4320]) );
XNOR U21604 ( .A(a[4320]), .B(c4320), .Z(n12962) );
XOR U21605 ( .A(c4321), .B(n12963), .Z(c4322) );
ANDN U21606 ( .B(n12964), .A(n12965), .Z(n12963) );
XOR U21607 ( .A(c4321), .B(b[4321]), .Z(n12964) );
XNOR U21608 ( .A(b[4321]), .B(n12965), .Z(c[4321]) );
XNOR U21609 ( .A(a[4321]), .B(c4321), .Z(n12965) );
XOR U21610 ( .A(c4322), .B(n12966), .Z(c4323) );
ANDN U21611 ( .B(n12967), .A(n12968), .Z(n12966) );
XOR U21612 ( .A(c4322), .B(b[4322]), .Z(n12967) );
XNOR U21613 ( .A(b[4322]), .B(n12968), .Z(c[4322]) );
XNOR U21614 ( .A(a[4322]), .B(c4322), .Z(n12968) );
XOR U21615 ( .A(c4323), .B(n12969), .Z(c4324) );
ANDN U21616 ( .B(n12970), .A(n12971), .Z(n12969) );
XOR U21617 ( .A(c4323), .B(b[4323]), .Z(n12970) );
XNOR U21618 ( .A(b[4323]), .B(n12971), .Z(c[4323]) );
XNOR U21619 ( .A(a[4323]), .B(c4323), .Z(n12971) );
XOR U21620 ( .A(c4324), .B(n12972), .Z(c4325) );
ANDN U21621 ( .B(n12973), .A(n12974), .Z(n12972) );
XOR U21622 ( .A(c4324), .B(b[4324]), .Z(n12973) );
XNOR U21623 ( .A(b[4324]), .B(n12974), .Z(c[4324]) );
XNOR U21624 ( .A(a[4324]), .B(c4324), .Z(n12974) );
XOR U21625 ( .A(c4325), .B(n12975), .Z(c4326) );
ANDN U21626 ( .B(n12976), .A(n12977), .Z(n12975) );
XOR U21627 ( .A(c4325), .B(b[4325]), .Z(n12976) );
XNOR U21628 ( .A(b[4325]), .B(n12977), .Z(c[4325]) );
XNOR U21629 ( .A(a[4325]), .B(c4325), .Z(n12977) );
XOR U21630 ( .A(c4326), .B(n12978), .Z(c4327) );
ANDN U21631 ( .B(n12979), .A(n12980), .Z(n12978) );
XOR U21632 ( .A(c4326), .B(b[4326]), .Z(n12979) );
XNOR U21633 ( .A(b[4326]), .B(n12980), .Z(c[4326]) );
XNOR U21634 ( .A(a[4326]), .B(c4326), .Z(n12980) );
XOR U21635 ( .A(c4327), .B(n12981), .Z(c4328) );
ANDN U21636 ( .B(n12982), .A(n12983), .Z(n12981) );
XOR U21637 ( .A(c4327), .B(b[4327]), .Z(n12982) );
XNOR U21638 ( .A(b[4327]), .B(n12983), .Z(c[4327]) );
XNOR U21639 ( .A(a[4327]), .B(c4327), .Z(n12983) );
XOR U21640 ( .A(c4328), .B(n12984), .Z(c4329) );
ANDN U21641 ( .B(n12985), .A(n12986), .Z(n12984) );
XOR U21642 ( .A(c4328), .B(b[4328]), .Z(n12985) );
XNOR U21643 ( .A(b[4328]), .B(n12986), .Z(c[4328]) );
XNOR U21644 ( .A(a[4328]), .B(c4328), .Z(n12986) );
XOR U21645 ( .A(c4329), .B(n12987), .Z(c4330) );
ANDN U21646 ( .B(n12988), .A(n12989), .Z(n12987) );
XOR U21647 ( .A(c4329), .B(b[4329]), .Z(n12988) );
XNOR U21648 ( .A(b[4329]), .B(n12989), .Z(c[4329]) );
XNOR U21649 ( .A(a[4329]), .B(c4329), .Z(n12989) );
XOR U21650 ( .A(c4330), .B(n12990), .Z(c4331) );
ANDN U21651 ( .B(n12991), .A(n12992), .Z(n12990) );
XOR U21652 ( .A(c4330), .B(b[4330]), .Z(n12991) );
XNOR U21653 ( .A(b[4330]), .B(n12992), .Z(c[4330]) );
XNOR U21654 ( .A(a[4330]), .B(c4330), .Z(n12992) );
XOR U21655 ( .A(c4331), .B(n12993), .Z(c4332) );
ANDN U21656 ( .B(n12994), .A(n12995), .Z(n12993) );
XOR U21657 ( .A(c4331), .B(b[4331]), .Z(n12994) );
XNOR U21658 ( .A(b[4331]), .B(n12995), .Z(c[4331]) );
XNOR U21659 ( .A(a[4331]), .B(c4331), .Z(n12995) );
XOR U21660 ( .A(c4332), .B(n12996), .Z(c4333) );
ANDN U21661 ( .B(n12997), .A(n12998), .Z(n12996) );
XOR U21662 ( .A(c4332), .B(b[4332]), .Z(n12997) );
XNOR U21663 ( .A(b[4332]), .B(n12998), .Z(c[4332]) );
XNOR U21664 ( .A(a[4332]), .B(c4332), .Z(n12998) );
XOR U21665 ( .A(c4333), .B(n12999), .Z(c4334) );
ANDN U21666 ( .B(n13000), .A(n13001), .Z(n12999) );
XOR U21667 ( .A(c4333), .B(b[4333]), .Z(n13000) );
XNOR U21668 ( .A(b[4333]), .B(n13001), .Z(c[4333]) );
XNOR U21669 ( .A(a[4333]), .B(c4333), .Z(n13001) );
XOR U21670 ( .A(c4334), .B(n13002), .Z(c4335) );
ANDN U21671 ( .B(n13003), .A(n13004), .Z(n13002) );
XOR U21672 ( .A(c4334), .B(b[4334]), .Z(n13003) );
XNOR U21673 ( .A(b[4334]), .B(n13004), .Z(c[4334]) );
XNOR U21674 ( .A(a[4334]), .B(c4334), .Z(n13004) );
XOR U21675 ( .A(c4335), .B(n13005), .Z(c4336) );
ANDN U21676 ( .B(n13006), .A(n13007), .Z(n13005) );
XOR U21677 ( .A(c4335), .B(b[4335]), .Z(n13006) );
XNOR U21678 ( .A(b[4335]), .B(n13007), .Z(c[4335]) );
XNOR U21679 ( .A(a[4335]), .B(c4335), .Z(n13007) );
XOR U21680 ( .A(c4336), .B(n13008), .Z(c4337) );
ANDN U21681 ( .B(n13009), .A(n13010), .Z(n13008) );
XOR U21682 ( .A(c4336), .B(b[4336]), .Z(n13009) );
XNOR U21683 ( .A(b[4336]), .B(n13010), .Z(c[4336]) );
XNOR U21684 ( .A(a[4336]), .B(c4336), .Z(n13010) );
XOR U21685 ( .A(c4337), .B(n13011), .Z(c4338) );
ANDN U21686 ( .B(n13012), .A(n13013), .Z(n13011) );
XOR U21687 ( .A(c4337), .B(b[4337]), .Z(n13012) );
XNOR U21688 ( .A(b[4337]), .B(n13013), .Z(c[4337]) );
XNOR U21689 ( .A(a[4337]), .B(c4337), .Z(n13013) );
XOR U21690 ( .A(c4338), .B(n13014), .Z(c4339) );
ANDN U21691 ( .B(n13015), .A(n13016), .Z(n13014) );
XOR U21692 ( .A(c4338), .B(b[4338]), .Z(n13015) );
XNOR U21693 ( .A(b[4338]), .B(n13016), .Z(c[4338]) );
XNOR U21694 ( .A(a[4338]), .B(c4338), .Z(n13016) );
XOR U21695 ( .A(c4339), .B(n13017), .Z(c4340) );
ANDN U21696 ( .B(n13018), .A(n13019), .Z(n13017) );
XOR U21697 ( .A(c4339), .B(b[4339]), .Z(n13018) );
XNOR U21698 ( .A(b[4339]), .B(n13019), .Z(c[4339]) );
XNOR U21699 ( .A(a[4339]), .B(c4339), .Z(n13019) );
XOR U21700 ( .A(c4340), .B(n13020), .Z(c4341) );
ANDN U21701 ( .B(n13021), .A(n13022), .Z(n13020) );
XOR U21702 ( .A(c4340), .B(b[4340]), .Z(n13021) );
XNOR U21703 ( .A(b[4340]), .B(n13022), .Z(c[4340]) );
XNOR U21704 ( .A(a[4340]), .B(c4340), .Z(n13022) );
XOR U21705 ( .A(c4341), .B(n13023), .Z(c4342) );
ANDN U21706 ( .B(n13024), .A(n13025), .Z(n13023) );
XOR U21707 ( .A(c4341), .B(b[4341]), .Z(n13024) );
XNOR U21708 ( .A(b[4341]), .B(n13025), .Z(c[4341]) );
XNOR U21709 ( .A(a[4341]), .B(c4341), .Z(n13025) );
XOR U21710 ( .A(c4342), .B(n13026), .Z(c4343) );
ANDN U21711 ( .B(n13027), .A(n13028), .Z(n13026) );
XOR U21712 ( .A(c4342), .B(b[4342]), .Z(n13027) );
XNOR U21713 ( .A(b[4342]), .B(n13028), .Z(c[4342]) );
XNOR U21714 ( .A(a[4342]), .B(c4342), .Z(n13028) );
XOR U21715 ( .A(c4343), .B(n13029), .Z(c4344) );
ANDN U21716 ( .B(n13030), .A(n13031), .Z(n13029) );
XOR U21717 ( .A(c4343), .B(b[4343]), .Z(n13030) );
XNOR U21718 ( .A(b[4343]), .B(n13031), .Z(c[4343]) );
XNOR U21719 ( .A(a[4343]), .B(c4343), .Z(n13031) );
XOR U21720 ( .A(c4344), .B(n13032), .Z(c4345) );
ANDN U21721 ( .B(n13033), .A(n13034), .Z(n13032) );
XOR U21722 ( .A(c4344), .B(b[4344]), .Z(n13033) );
XNOR U21723 ( .A(b[4344]), .B(n13034), .Z(c[4344]) );
XNOR U21724 ( .A(a[4344]), .B(c4344), .Z(n13034) );
XOR U21725 ( .A(c4345), .B(n13035), .Z(c4346) );
ANDN U21726 ( .B(n13036), .A(n13037), .Z(n13035) );
XOR U21727 ( .A(c4345), .B(b[4345]), .Z(n13036) );
XNOR U21728 ( .A(b[4345]), .B(n13037), .Z(c[4345]) );
XNOR U21729 ( .A(a[4345]), .B(c4345), .Z(n13037) );
XOR U21730 ( .A(c4346), .B(n13038), .Z(c4347) );
ANDN U21731 ( .B(n13039), .A(n13040), .Z(n13038) );
XOR U21732 ( .A(c4346), .B(b[4346]), .Z(n13039) );
XNOR U21733 ( .A(b[4346]), .B(n13040), .Z(c[4346]) );
XNOR U21734 ( .A(a[4346]), .B(c4346), .Z(n13040) );
XOR U21735 ( .A(c4347), .B(n13041), .Z(c4348) );
ANDN U21736 ( .B(n13042), .A(n13043), .Z(n13041) );
XOR U21737 ( .A(c4347), .B(b[4347]), .Z(n13042) );
XNOR U21738 ( .A(b[4347]), .B(n13043), .Z(c[4347]) );
XNOR U21739 ( .A(a[4347]), .B(c4347), .Z(n13043) );
XOR U21740 ( .A(c4348), .B(n13044), .Z(c4349) );
ANDN U21741 ( .B(n13045), .A(n13046), .Z(n13044) );
XOR U21742 ( .A(c4348), .B(b[4348]), .Z(n13045) );
XNOR U21743 ( .A(b[4348]), .B(n13046), .Z(c[4348]) );
XNOR U21744 ( .A(a[4348]), .B(c4348), .Z(n13046) );
XOR U21745 ( .A(c4349), .B(n13047), .Z(c4350) );
ANDN U21746 ( .B(n13048), .A(n13049), .Z(n13047) );
XOR U21747 ( .A(c4349), .B(b[4349]), .Z(n13048) );
XNOR U21748 ( .A(b[4349]), .B(n13049), .Z(c[4349]) );
XNOR U21749 ( .A(a[4349]), .B(c4349), .Z(n13049) );
XOR U21750 ( .A(c4350), .B(n13050), .Z(c4351) );
ANDN U21751 ( .B(n13051), .A(n13052), .Z(n13050) );
XOR U21752 ( .A(c4350), .B(b[4350]), .Z(n13051) );
XNOR U21753 ( .A(b[4350]), .B(n13052), .Z(c[4350]) );
XNOR U21754 ( .A(a[4350]), .B(c4350), .Z(n13052) );
XOR U21755 ( .A(c4351), .B(n13053), .Z(c4352) );
ANDN U21756 ( .B(n13054), .A(n13055), .Z(n13053) );
XOR U21757 ( .A(c4351), .B(b[4351]), .Z(n13054) );
XNOR U21758 ( .A(b[4351]), .B(n13055), .Z(c[4351]) );
XNOR U21759 ( .A(a[4351]), .B(c4351), .Z(n13055) );
XOR U21760 ( .A(c4352), .B(n13056), .Z(c4353) );
ANDN U21761 ( .B(n13057), .A(n13058), .Z(n13056) );
XOR U21762 ( .A(c4352), .B(b[4352]), .Z(n13057) );
XNOR U21763 ( .A(b[4352]), .B(n13058), .Z(c[4352]) );
XNOR U21764 ( .A(a[4352]), .B(c4352), .Z(n13058) );
XOR U21765 ( .A(c4353), .B(n13059), .Z(c4354) );
ANDN U21766 ( .B(n13060), .A(n13061), .Z(n13059) );
XOR U21767 ( .A(c4353), .B(b[4353]), .Z(n13060) );
XNOR U21768 ( .A(b[4353]), .B(n13061), .Z(c[4353]) );
XNOR U21769 ( .A(a[4353]), .B(c4353), .Z(n13061) );
XOR U21770 ( .A(c4354), .B(n13062), .Z(c4355) );
ANDN U21771 ( .B(n13063), .A(n13064), .Z(n13062) );
XOR U21772 ( .A(c4354), .B(b[4354]), .Z(n13063) );
XNOR U21773 ( .A(b[4354]), .B(n13064), .Z(c[4354]) );
XNOR U21774 ( .A(a[4354]), .B(c4354), .Z(n13064) );
XOR U21775 ( .A(c4355), .B(n13065), .Z(c4356) );
ANDN U21776 ( .B(n13066), .A(n13067), .Z(n13065) );
XOR U21777 ( .A(c4355), .B(b[4355]), .Z(n13066) );
XNOR U21778 ( .A(b[4355]), .B(n13067), .Z(c[4355]) );
XNOR U21779 ( .A(a[4355]), .B(c4355), .Z(n13067) );
XOR U21780 ( .A(c4356), .B(n13068), .Z(c4357) );
ANDN U21781 ( .B(n13069), .A(n13070), .Z(n13068) );
XOR U21782 ( .A(c4356), .B(b[4356]), .Z(n13069) );
XNOR U21783 ( .A(b[4356]), .B(n13070), .Z(c[4356]) );
XNOR U21784 ( .A(a[4356]), .B(c4356), .Z(n13070) );
XOR U21785 ( .A(c4357), .B(n13071), .Z(c4358) );
ANDN U21786 ( .B(n13072), .A(n13073), .Z(n13071) );
XOR U21787 ( .A(c4357), .B(b[4357]), .Z(n13072) );
XNOR U21788 ( .A(b[4357]), .B(n13073), .Z(c[4357]) );
XNOR U21789 ( .A(a[4357]), .B(c4357), .Z(n13073) );
XOR U21790 ( .A(c4358), .B(n13074), .Z(c4359) );
ANDN U21791 ( .B(n13075), .A(n13076), .Z(n13074) );
XOR U21792 ( .A(c4358), .B(b[4358]), .Z(n13075) );
XNOR U21793 ( .A(b[4358]), .B(n13076), .Z(c[4358]) );
XNOR U21794 ( .A(a[4358]), .B(c4358), .Z(n13076) );
XOR U21795 ( .A(c4359), .B(n13077), .Z(c4360) );
ANDN U21796 ( .B(n13078), .A(n13079), .Z(n13077) );
XOR U21797 ( .A(c4359), .B(b[4359]), .Z(n13078) );
XNOR U21798 ( .A(b[4359]), .B(n13079), .Z(c[4359]) );
XNOR U21799 ( .A(a[4359]), .B(c4359), .Z(n13079) );
XOR U21800 ( .A(c4360), .B(n13080), .Z(c4361) );
ANDN U21801 ( .B(n13081), .A(n13082), .Z(n13080) );
XOR U21802 ( .A(c4360), .B(b[4360]), .Z(n13081) );
XNOR U21803 ( .A(b[4360]), .B(n13082), .Z(c[4360]) );
XNOR U21804 ( .A(a[4360]), .B(c4360), .Z(n13082) );
XOR U21805 ( .A(c4361), .B(n13083), .Z(c4362) );
ANDN U21806 ( .B(n13084), .A(n13085), .Z(n13083) );
XOR U21807 ( .A(c4361), .B(b[4361]), .Z(n13084) );
XNOR U21808 ( .A(b[4361]), .B(n13085), .Z(c[4361]) );
XNOR U21809 ( .A(a[4361]), .B(c4361), .Z(n13085) );
XOR U21810 ( .A(c4362), .B(n13086), .Z(c4363) );
ANDN U21811 ( .B(n13087), .A(n13088), .Z(n13086) );
XOR U21812 ( .A(c4362), .B(b[4362]), .Z(n13087) );
XNOR U21813 ( .A(b[4362]), .B(n13088), .Z(c[4362]) );
XNOR U21814 ( .A(a[4362]), .B(c4362), .Z(n13088) );
XOR U21815 ( .A(c4363), .B(n13089), .Z(c4364) );
ANDN U21816 ( .B(n13090), .A(n13091), .Z(n13089) );
XOR U21817 ( .A(c4363), .B(b[4363]), .Z(n13090) );
XNOR U21818 ( .A(b[4363]), .B(n13091), .Z(c[4363]) );
XNOR U21819 ( .A(a[4363]), .B(c4363), .Z(n13091) );
XOR U21820 ( .A(c4364), .B(n13092), .Z(c4365) );
ANDN U21821 ( .B(n13093), .A(n13094), .Z(n13092) );
XOR U21822 ( .A(c4364), .B(b[4364]), .Z(n13093) );
XNOR U21823 ( .A(b[4364]), .B(n13094), .Z(c[4364]) );
XNOR U21824 ( .A(a[4364]), .B(c4364), .Z(n13094) );
XOR U21825 ( .A(c4365), .B(n13095), .Z(c4366) );
ANDN U21826 ( .B(n13096), .A(n13097), .Z(n13095) );
XOR U21827 ( .A(c4365), .B(b[4365]), .Z(n13096) );
XNOR U21828 ( .A(b[4365]), .B(n13097), .Z(c[4365]) );
XNOR U21829 ( .A(a[4365]), .B(c4365), .Z(n13097) );
XOR U21830 ( .A(c4366), .B(n13098), .Z(c4367) );
ANDN U21831 ( .B(n13099), .A(n13100), .Z(n13098) );
XOR U21832 ( .A(c4366), .B(b[4366]), .Z(n13099) );
XNOR U21833 ( .A(b[4366]), .B(n13100), .Z(c[4366]) );
XNOR U21834 ( .A(a[4366]), .B(c4366), .Z(n13100) );
XOR U21835 ( .A(c4367), .B(n13101), .Z(c4368) );
ANDN U21836 ( .B(n13102), .A(n13103), .Z(n13101) );
XOR U21837 ( .A(c4367), .B(b[4367]), .Z(n13102) );
XNOR U21838 ( .A(b[4367]), .B(n13103), .Z(c[4367]) );
XNOR U21839 ( .A(a[4367]), .B(c4367), .Z(n13103) );
XOR U21840 ( .A(c4368), .B(n13104), .Z(c4369) );
ANDN U21841 ( .B(n13105), .A(n13106), .Z(n13104) );
XOR U21842 ( .A(c4368), .B(b[4368]), .Z(n13105) );
XNOR U21843 ( .A(b[4368]), .B(n13106), .Z(c[4368]) );
XNOR U21844 ( .A(a[4368]), .B(c4368), .Z(n13106) );
XOR U21845 ( .A(c4369), .B(n13107), .Z(c4370) );
ANDN U21846 ( .B(n13108), .A(n13109), .Z(n13107) );
XOR U21847 ( .A(c4369), .B(b[4369]), .Z(n13108) );
XNOR U21848 ( .A(b[4369]), .B(n13109), .Z(c[4369]) );
XNOR U21849 ( .A(a[4369]), .B(c4369), .Z(n13109) );
XOR U21850 ( .A(c4370), .B(n13110), .Z(c4371) );
ANDN U21851 ( .B(n13111), .A(n13112), .Z(n13110) );
XOR U21852 ( .A(c4370), .B(b[4370]), .Z(n13111) );
XNOR U21853 ( .A(b[4370]), .B(n13112), .Z(c[4370]) );
XNOR U21854 ( .A(a[4370]), .B(c4370), .Z(n13112) );
XOR U21855 ( .A(c4371), .B(n13113), .Z(c4372) );
ANDN U21856 ( .B(n13114), .A(n13115), .Z(n13113) );
XOR U21857 ( .A(c4371), .B(b[4371]), .Z(n13114) );
XNOR U21858 ( .A(b[4371]), .B(n13115), .Z(c[4371]) );
XNOR U21859 ( .A(a[4371]), .B(c4371), .Z(n13115) );
XOR U21860 ( .A(c4372), .B(n13116), .Z(c4373) );
ANDN U21861 ( .B(n13117), .A(n13118), .Z(n13116) );
XOR U21862 ( .A(c4372), .B(b[4372]), .Z(n13117) );
XNOR U21863 ( .A(b[4372]), .B(n13118), .Z(c[4372]) );
XNOR U21864 ( .A(a[4372]), .B(c4372), .Z(n13118) );
XOR U21865 ( .A(c4373), .B(n13119), .Z(c4374) );
ANDN U21866 ( .B(n13120), .A(n13121), .Z(n13119) );
XOR U21867 ( .A(c4373), .B(b[4373]), .Z(n13120) );
XNOR U21868 ( .A(b[4373]), .B(n13121), .Z(c[4373]) );
XNOR U21869 ( .A(a[4373]), .B(c4373), .Z(n13121) );
XOR U21870 ( .A(c4374), .B(n13122), .Z(c4375) );
ANDN U21871 ( .B(n13123), .A(n13124), .Z(n13122) );
XOR U21872 ( .A(c4374), .B(b[4374]), .Z(n13123) );
XNOR U21873 ( .A(b[4374]), .B(n13124), .Z(c[4374]) );
XNOR U21874 ( .A(a[4374]), .B(c4374), .Z(n13124) );
XOR U21875 ( .A(c4375), .B(n13125), .Z(c4376) );
ANDN U21876 ( .B(n13126), .A(n13127), .Z(n13125) );
XOR U21877 ( .A(c4375), .B(b[4375]), .Z(n13126) );
XNOR U21878 ( .A(b[4375]), .B(n13127), .Z(c[4375]) );
XNOR U21879 ( .A(a[4375]), .B(c4375), .Z(n13127) );
XOR U21880 ( .A(c4376), .B(n13128), .Z(c4377) );
ANDN U21881 ( .B(n13129), .A(n13130), .Z(n13128) );
XOR U21882 ( .A(c4376), .B(b[4376]), .Z(n13129) );
XNOR U21883 ( .A(b[4376]), .B(n13130), .Z(c[4376]) );
XNOR U21884 ( .A(a[4376]), .B(c4376), .Z(n13130) );
XOR U21885 ( .A(c4377), .B(n13131), .Z(c4378) );
ANDN U21886 ( .B(n13132), .A(n13133), .Z(n13131) );
XOR U21887 ( .A(c4377), .B(b[4377]), .Z(n13132) );
XNOR U21888 ( .A(b[4377]), .B(n13133), .Z(c[4377]) );
XNOR U21889 ( .A(a[4377]), .B(c4377), .Z(n13133) );
XOR U21890 ( .A(c4378), .B(n13134), .Z(c4379) );
ANDN U21891 ( .B(n13135), .A(n13136), .Z(n13134) );
XOR U21892 ( .A(c4378), .B(b[4378]), .Z(n13135) );
XNOR U21893 ( .A(b[4378]), .B(n13136), .Z(c[4378]) );
XNOR U21894 ( .A(a[4378]), .B(c4378), .Z(n13136) );
XOR U21895 ( .A(c4379), .B(n13137), .Z(c4380) );
ANDN U21896 ( .B(n13138), .A(n13139), .Z(n13137) );
XOR U21897 ( .A(c4379), .B(b[4379]), .Z(n13138) );
XNOR U21898 ( .A(b[4379]), .B(n13139), .Z(c[4379]) );
XNOR U21899 ( .A(a[4379]), .B(c4379), .Z(n13139) );
XOR U21900 ( .A(c4380), .B(n13140), .Z(c4381) );
ANDN U21901 ( .B(n13141), .A(n13142), .Z(n13140) );
XOR U21902 ( .A(c4380), .B(b[4380]), .Z(n13141) );
XNOR U21903 ( .A(b[4380]), .B(n13142), .Z(c[4380]) );
XNOR U21904 ( .A(a[4380]), .B(c4380), .Z(n13142) );
XOR U21905 ( .A(c4381), .B(n13143), .Z(c4382) );
ANDN U21906 ( .B(n13144), .A(n13145), .Z(n13143) );
XOR U21907 ( .A(c4381), .B(b[4381]), .Z(n13144) );
XNOR U21908 ( .A(b[4381]), .B(n13145), .Z(c[4381]) );
XNOR U21909 ( .A(a[4381]), .B(c4381), .Z(n13145) );
XOR U21910 ( .A(c4382), .B(n13146), .Z(c4383) );
ANDN U21911 ( .B(n13147), .A(n13148), .Z(n13146) );
XOR U21912 ( .A(c4382), .B(b[4382]), .Z(n13147) );
XNOR U21913 ( .A(b[4382]), .B(n13148), .Z(c[4382]) );
XNOR U21914 ( .A(a[4382]), .B(c4382), .Z(n13148) );
XOR U21915 ( .A(c4383), .B(n13149), .Z(c4384) );
ANDN U21916 ( .B(n13150), .A(n13151), .Z(n13149) );
XOR U21917 ( .A(c4383), .B(b[4383]), .Z(n13150) );
XNOR U21918 ( .A(b[4383]), .B(n13151), .Z(c[4383]) );
XNOR U21919 ( .A(a[4383]), .B(c4383), .Z(n13151) );
XOR U21920 ( .A(c4384), .B(n13152), .Z(c4385) );
ANDN U21921 ( .B(n13153), .A(n13154), .Z(n13152) );
XOR U21922 ( .A(c4384), .B(b[4384]), .Z(n13153) );
XNOR U21923 ( .A(b[4384]), .B(n13154), .Z(c[4384]) );
XNOR U21924 ( .A(a[4384]), .B(c4384), .Z(n13154) );
XOR U21925 ( .A(c4385), .B(n13155), .Z(c4386) );
ANDN U21926 ( .B(n13156), .A(n13157), .Z(n13155) );
XOR U21927 ( .A(c4385), .B(b[4385]), .Z(n13156) );
XNOR U21928 ( .A(b[4385]), .B(n13157), .Z(c[4385]) );
XNOR U21929 ( .A(a[4385]), .B(c4385), .Z(n13157) );
XOR U21930 ( .A(c4386), .B(n13158), .Z(c4387) );
ANDN U21931 ( .B(n13159), .A(n13160), .Z(n13158) );
XOR U21932 ( .A(c4386), .B(b[4386]), .Z(n13159) );
XNOR U21933 ( .A(b[4386]), .B(n13160), .Z(c[4386]) );
XNOR U21934 ( .A(a[4386]), .B(c4386), .Z(n13160) );
XOR U21935 ( .A(c4387), .B(n13161), .Z(c4388) );
ANDN U21936 ( .B(n13162), .A(n13163), .Z(n13161) );
XOR U21937 ( .A(c4387), .B(b[4387]), .Z(n13162) );
XNOR U21938 ( .A(b[4387]), .B(n13163), .Z(c[4387]) );
XNOR U21939 ( .A(a[4387]), .B(c4387), .Z(n13163) );
XOR U21940 ( .A(c4388), .B(n13164), .Z(c4389) );
ANDN U21941 ( .B(n13165), .A(n13166), .Z(n13164) );
XOR U21942 ( .A(c4388), .B(b[4388]), .Z(n13165) );
XNOR U21943 ( .A(b[4388]), .B(n13166), .Z(c[4388]) );
XNOR U21944 ( .A(a[4388]), .B(c4388), .Z(n13166) );
XOR U21945 ( .A(c4389), .B(n13167), .Z(c4390) );
ANDN U21946 ( .B(n13168), .A(n13169), .Z(n13167) );
XOR U21947 ( .A(c4389), .B(b[4389]), .Z(n13168) );
XNOR U21948 ( .A(b[4389]), .B(n13169), .Z(c[4389]) );
XNOR U21949 ( .A(a[4389]), .B(c4389), .Z(n13169) );
XOR U21950 ( .A(c4390), .B(n13170), .Z(c4391) );
ANDN U21951 ( .B(n13171), .A(n13172), .Z(n13170) );
XOR U21952 ( .A(c4390), .B(b[4390]), .Z(n13171) );
XNOR U21953 ( .A(b[4390]), .B(n13172), .Z(c[4390]) );
XNOR U21954 ( .A(a[4390]), .B(c4390), .Z(n13172) );
XOR U21955 ( .A(c4391), .B(n13173), .Z(c4392) );
ANDN U21956 ( .B(n13174), .A(n13175), .Z(n13173) );
XOR U21957 ( .A(c4391), .B(b[4391]), .Z(n13174) );
XNOR U21958 ( .A(b[4391]), .B(n13175), .Z(c[4391]) );
XNOR U21959 ( .A(a[4391]), .B(c4391), .Z(n13175) );
XOR U21960 ( .A(c4392), .B(n13176), .Z(c4393) );
ANDN U21961 ( .B(n13177), .A(n13178), .Z(n13176) );
XOR U21962 ( .A(c4392), .B(b[4392]), .Z(n13177) );
XNOR U21963 ( .A(b[4392]), .B(n13178), .Z(c[4392]) );
XNOR U21964 ( .A(a[4392]), .B(c4392), .Z(n13178) );
XOR U21965 ( .A(c4393), .B(n13179), .Z(c4394) );
ANDN U21966 ( .B(n13180), .A(n13181), .Z(n13179) );
XOR U21967 ( .A(c4393), .B(b[4393]), .Z(n13180) );
XNOR U21968 ( .A(b[4393]), .B(n13181), .Z(c[4393]) );
XNOR U21969 ( .A(a[4393]), .B(c4393), .Z(n13181) );
XOR U21970 ( .A(c4394), .B(n13182), .Z(c4395) );
ANDN U21971 ( .B(n13183), .A(n13184), .Z(n13182) );
XOR U21972 ( .A(c4394), .B(b[4394]), .Z(n13183) );
XNOR U21973 ( .A(b[4394]), .B(n13184), .Z(c[4394]) );
XNOR U21974 ( .A(a[4394]), .B(c4394), .Z(n13184) );
XOR U21975 ( .A(c4395), .B(n13185), .Z(c4396) );
ANDN U21976 ( .B(n13186), .A(n13187), .Z(n13185) );
XOR U21977 ( .A(c4395), .B(b[4395]), .Z(n13186) );
XNOR U21978 ( .A(b[4395]), .B(n13187), .Z(c[4395]) );
XNOR U21979 ( .A(a[4395]), .B(c4395), .Z(n13187) );
XOR U21980 ( .A(c4396), .B(n13188), .Z(c4397) );
ANDN U21981 ( .B(n13189), .A(n13190), .Z(n13188) );
XOR U21982 ( .A(c4396), .B(b[4396]), .Z(n13189) );
XNOR U21983 ( .A(b[4396]), .B(n13190), .Z(c[4396]) );
XNOR U21984 ( .A(a[4396]), .B(c4396), .Z(n13190) );
XOR U21985 ( .A(c4397), .B(n13191), .Z(c4398) );
ANDN U21986 ( .B(n13192), .A(n13193), .Z(n13191) );
XOR U21987 ( .A(c4397), .B(b[4397]), .Z(n13192) );
XNOR U21988 ( .A(b[4397]), .B(n13193), .Z(c[4397]) );
XNOR U21989 ( .A(a[4397]), .B(c4397), .Z(n13193) );
XOR U21990 ( .A(c4398), .B(n13194), .Z(c4399) );
ANDN U21991 ( .B(n13195), .A(n13196), .Z(n13194) );
XOR U21992 ( .A(c4398), .B(b[4398]), .Z(n13195) );
XNOR U21993 ( .A(b[4398]), .B(n13196), .Z(c[4398]) );
XNOR U21994 ( .A(a[4398]), .B(c4398), .Z(n13196) );
XOR U21995 ( .A(c4399), .B(n13197), .Z(c4400) );
ANDN U21996 ( .B(n13198), .A(n13199), .Z(n13197) );
XOR U21997 ( .A(c4399), .B(b[4399]), .Z(n13198) );
XNOR U21998 ( .A(b[4399]), .B(n13199), .Z(c[4399]) );
XNOR U21999 ( .A(a[4399]), .B(c4399), .Z(n13199) );
XOR U22000 ( .A(c4400), .B(n13200), .Z(c4401) );
ANDN U22001 ( .B(n13201), .A(n13202), .Z(n13200) );
XOR U22002 ( .A(c4400), .B(b[4400]), .Z(n13201) );
XNOR U22003 ( .A(b[4400]), .B(n13202), .Z(c[4400]) );
XNOR U22004 ( .A(a[4400]), .B(c4400), .Z(n13202) );
XOR U22005 ( .A(c4401), .B(n13203), .Z(c4402) );
ANDN U22006 ( .B(n13204), .A(n13205), .Z(n13203) );
XOR U22007 ( .A(c4401), .B(b[4401]), .Z(n13204) );
XNOR U22008 ( .A(b[4401]), .B(n13205), .Z(c[4401]) );
XNOR U22009 ( .A(a[4401]), .B(c4401), .Z(n13205) );
XOR U22010 ( .A(c4402), .B(n13206), .Z(c4403) );
ANDN U22011 ( .B(n13207), .A(n13208), .Z(n13206) );
XOR U22012 ( .A(c4402), .B(b[4402]), .Z(n13207) );
XNOR U22013 ( .A(b[4402]), .B(n13208), .Z(c[4402]) );
XNOR U22014 ( .A(a[4402]), .B(c4402), .Z(n13208) );
XOR U22015 ( .A(c4403), .B(n13209), .Z(c4404) );
ANDN U22016 ( .B(n13210), .A(n13211), .Z(n13209) );
XOR U22017 ( .A(c4403), .B(b[4403]), .Z(n13210) );
XNOR U22018 ( .A(b[4403]), .B(n13211), .Z(c[4403]) );
XNOR U22019 ( .A(a[4403]), .B(c4403), .Z(n13211) );
XOR U22020 ( .A(c4404), .B(n13212), .Z(c4405) );
ANDN U22021 ( .B(n13213), .A(n13214), .Z(n13212) );
XOR U22022 ( .A(c4404), .B(b[4404]), .Z(n13213) );
XNOR U22023 ( .A(b[4404]), .B(n13214), .Z(c[4404]) );
XNOR U22024 ( .A(a[4404]), .B(c4404), .Z(n13214) );
XOR U22025 ( .A(c4405), .B(n13215), .Z(c4406) );
ANDN U22026 ( .B(n13216), .A(n13217), .Z(n13215) );
XOR U22027 ( .A(c4405), .B(b[4405]), .Z(n13216) );
XNOR U22028 ( .A(b[4405]), .B(n13217), .Z(c[4405]) );
XNOR U22029 ( .A(a[4405]), .B(c4405), .Z(n13217) );
XOR U22030 ( .A(c4406), .B(n13218), .Z(c4407) );
ANDN U22031 ( .B(n13219), .A(n13220), .Z(n13218) );
XOR U22032 ( .A(c4406), .B(b[4406]), .Z(n13219) );
XNOR U22033 ( .A(b[4406]), .B(n13220), .Z(c[4406]) );
XNOR U22034 ( .A(a[4406]), .B(c4406), .Z(n13220) );
XOR U22035 ( .A(c4407), .B(n13221), .Z(c4408) );
ANDN U22036 ( .B(n13222), .A(n13223), .Z(n13221) );
XOR U22037 ( .A(c4407), .B(b[4407]), .Z(n13222) );
XNOR U22038 ( .A(b[4407]), .B(n13223), .Z(c[4407]) );
XNOR U22039 ( .A(a[4407]), .B(c4407), .Z(n13223) );
XOR U22040 ( .A(c4408), .B(n13224), .Z(c4409) );
ANDN U22041 ( .B(n13225), .A(n13226), .Z(n13224) );
XOR U22042 ( .A(c4408), .B(b[4408]), .Z(n13225) );
XNOR U22043 ( .A(b[4408]), .B(n13226), .Z(c[4408]) );
XNOR U22044 ( .A(a[4408]), .B(c4408), .Z(n13226) );
XOR U22045 ( .A(c4409), .B(n13227), .Z(c4410) );
ANDN U22046 ( .B(n13228), .A(n13229), .Z(n13227) );
XOR U22047 ( .A(c4409), .B(b[4409]), .Z(n13228) );
XNOR U22048 ( .A(b[4409]), .B(n13229), .Z(c[4409]) );
XNOR U22049 ( .A(a[4409]), .B(c4409), .Z(n13229) );
XOR U22050 ( .A(c4410), .B(n13230), .Z(c4411) );
ANDN U22051 ( .B(n13231), .A(n13232), .Z(n13230) );
XOR U22052 ( .A(c4410), .B(b[4410]), .Z(n13231) );
XNOR U22053 ( .A(b[4410]), .B(n13232), .Z(c[4410]) );
XNOR U22054 ( .A(a[4410]), .B(c4410), .Z(n13232) );
XOR U22055 ( .A(c4411), .B(n13233), .Z(c4412) );
ANDN U22056 ( .B(n13234), .A(n13235), .Z(n13233) );
XOR U22057 ( .A(c4411), .B(b[4411]), .Z(n13234) );
XNOR U22058 ( .A(b[4411]), .B(n13235), .Z(c[4411]) );
XNOR U22059 ( .A(a[4411]), .B(c4411), .Z(n13235) );
XOR U22060 ( .A(c4412), .B(n13236), .Z(c4413) );
ANDN U22061 ( .B(n13237), .A(n13238), .Z(n13236) );
XOR U22062 ( .A(c4412), .B(b[4412]), .Z(n13237) );
XNOR U22063 ( .A(b[4412]), .B(n13238), .Z(c[4412]) );
XNOR U22064 ( .A(a[4412]), .B(c4412), .Z(n13238) );
XOR U22065 ( .A(c4413), .B(n13239), .Z(c4414) );
ANDN U22066 ( .B(n13240), .A(n13241), .Z(n13239) );
XOR U22067 ( .A(c4413), .B(b[4413]), .Z(n13240) );
XNOR U22068 ( .A(b[4413]), .B(n13241), .Z(c[4413]) );
XNOR U22069 ( .A(a[4413]), .B(c4413), .Z(n13241) );
XOR U22070 ( .A(c4414), .B(n13242), .Z(c4415) );
ANDN U22071 ( .B(n13243), .A(n13244), .Z(n13242) );
XOR U22072 ( .A(c4414), .B(b[4414]), .Z(n13243) );
XNOR U22073 ( .A(b[4414]), .B(n13244), .Z(c[4414]) );
XNOR U22074 ( .A(a[4414]), .B(c4414), .Z(n13244) );
XOR U22075 ( .A(c4415), .B(n13245), .Z(c4416) );
ANDN U22076 ( .B(n13246), .A(n13247), .Z(n13245) );
XOR U22077 ( .A(c4415), .B(b[4415]), .Z(n13246) );
XNOR U22078 ( .A(b[4415]), .B(n13247), .Z(c[4415]) );
XNOR U22079 ( .A(a[4415]), .B(c4415), .Z(n13247) );
XOR U22080 ( .A(c4416), .B(n13248), .Z(c4417) );
ANDN U22081 ( .B(n13249), .A(n13250), .Z(n13248) );
XOR U22082 ( .A(c4416), .B(b[4416]), .Z(n13249) );
XNOR U22083 ( .A(b[4416]), .B(n13250), .Z(c[4416]) );
XNOR U22084 ( .A(a[4416]), .B(c4416), .Z(n13250) );
XOR U22085 ( .A(c4417), .B(n13251), .Z(c4418) );
ANDN U22086 ( .B(n13252), .A(n13253), .Z(n13251) );
XOR U22087 ( .A(c4417), .B(b[4417]), .Z(n13252) );
XNOR U22088 ( .A(b[4417]), .B(n13253), .Z(c[4417]) );
XNOR U22089 ( .A(a[4417]), .B(c4417), .Z(n13253) );
XOR U22090 ( .A(c4418), .B(n13254), .Z(c4419) );
ANDN U22091 ( .B(n13255), .A(n13256), .Z(n13254) );
XOR U22092 ( .A(c4418), .B(b[4418]), .Z(n13255) );
XNOR U22093 ( .A(b[4418]), .B(n13256), .Z(c[4418]) );
XNOR U22094 ( .A(a[4418]), .B(c4418), .Z(n13256) );
XOR U22095 ( .A(c4419), .B(n13257), .Z(c4420) );
ANDN U22096 ( .B(n13258), .A(n13259), .Z(n13257) );
XOR U22097 ( .A(c4419), .B(b[4419]), .Z(n13258) );
XNOR U22098 ( .A(b[4419]), .B(n13259), .Z(c[4419]) );
XNOR U22099 ( .A(a[4419]), .B(c4419), .Z(n13259) );
XOR U22100 ( .A(c4420), .B(n13260), .Z(c4421) );
ANDN U22101 ( .B(n13261), .A(n13262), .Z(n13260) );
XOR U22102 ( .A(c4420), .B(b[4420]), .Z(n13261) );
XNOR U22103 ( .A(b[4420]), .B(n13262), .Z(c[4420]) );
XNOR U22104 ( .A(a[4420]), .B(c4420), .Z(n13262) );
XOR U22105 ( .A(c4421), .B(n13263), .Z(c4422) );
ANDN U22106 ( .B(n13264), .A(n13265), .Z(n13263) );
XOR U22107 ( .A(c4421), .B(b[4421]), .Z(n13264) );
XNOR U22108 ( .A(b[4421]), .B(n13265), .Z(c[4421]) );
XNOR U22109 ( .A(a[4421]), .B(c4421), .Z(n13265) );
XOR U22110 ( .A(c4422), .B(n13266), .Z(c4423) );
ANDN U22111 ( .B(n13267), .A(n13268), .Z(n13266) );
XOR U22112 ( .A(c4422), .B(b[4422]), .Z(n13267) );
XNOR U22113 ( .A(b[4422]), .B(n13268), .Z(c[4422]) );
XNOR U22114 ( .A(a[4422]), .B(c4422), .Z(n13268) );
XOR U22115 ( .A(c4423), .B(n13269), .Z(c4424) );
ANDN U22116 ( .B(n13270), .A(n13271), .Z(n13269) );
XOR U22117 ( .A(c4423), .B(b[4423]), .Z(n13270) );
XNOR U22118 ( .A(b[4423]), .B(n13271), .Z(c[4423]) );
XNOR U22119 ( .A(a[4423]), .B(c4423), .Z(n13271) );
XOR U22120 ( .A(c4424), .B(n13272), .Z(c4425) );
ANDN U22121 ( .B(n13273), .A(n13274), .Z(n13272) );
XOR U22122 ( .A(c4424), .B(b[4424]), .Z(n13273) );
XNOR U22123 ( .A(b[4424]), .B(n13274), .Z(c[4424]) );
XNOR U22124 ( .A(a[4424]), .B(c4424), .Z(n13274) );
XOR U22125 ( .A(c4425), .B(n13275), .Z(c4426) );
ANDN U22126 ( .B(n13276), .A(n13277), .Z(n13275) );
XOR U22127 ( .A(c4425), .B(b[4425]), .Z(n13276) );
XNOR U22128 ( .A(b[4425]), .B(n13277), .Z(c[4425]) );
XNOR U22129 ( .A(a[4425]), .B(c4425), .Z(n13277) );
XOR U22130 ( .A(c4426), .B(n13278), .Z(c4427) );
ANDN U22131 ( .B(n13279), .A(n13280), .Z(n13278) );
XOR U22132 ( .A(c4426), .B(b[4426]), .Z(n13279) );
XNOR U22133 ( .A(b[4426]), .B(n13280), .Z(c[4426]) );
XNOR U22134 ( .A(a[4426]), .B(c4426), .Z(n13280) );
XOR U22135 ( .A(c4427), .B(n13281), .Z(c4428) );
ANDN U22136 ( .B(n13282), .A(n13283), .Z(n13281) );
XOR U22137 ( .A(c4427), .B(b[4427]), .Z(n13282) );
XNOR U22138 ( .A(b[4427]), .B(n13283), .Z(c[4427]) );
XNOR U22139 ( .A(a[4427]), .B(c4427), .Z(n13283) );
XOR U22140 ( .A(c4428), .B(n13284), .Z(c4429) );
ANDN U22141 ( .B(n13285), .A(n13286), .Z(n13284) );
XOR U22142 ( .A(c4428), .B(b[4428]), .Z(n13285) );
XNOR U22143 ( .A(b[4428]), .B(n13286), .Z(c[4428]) );
XNOR U22144 ( .A(a[4428]), .B(c4428), .Z(n13286) );
XOR U22145 ( .A(c4429), .B(n13287), .Z(c4430) );
ANDN U22146 ( .B(n13288), .A(n13289), .Z(n13287) );
XOR U22147 ( .A(c4429), .B(b[4429]), .Z(n13288) );
XNOR U22148 ( .A(b[4429]), .B(n13289), .Z(c[4429]) );
XNOR U22149 ( .A(a[4429]), .B(c4429), .Z(n13289) );
XOR U22150 ( .A(c4430), .B(n13290), .Z(c4431) );
ANDN U22151 ( .B(n13291), .A(n13292), .Z(n13290) );
XOR U22152 ( .A(c4430), .B(b[4430]), .Z(n13291) );
XNOR U22153 ( .A(b[4430]), .B(n13292), .Z(c[4430]) );
XNOR U22154 ( .A(a[4430]), .B(c4430), .Z(n13292) );
XOR U22155 ( .A(c4431), .B(n13293), .Z(c4432) );
ANDN U22156 ( .B(n13294), .A(n13295), .Z(n13293) );
XOR U22157 ( .A(c4431), .B(b[4431]), .Z(n13294) );
XNOR U22158 ( .A(b[4431]), .B(n13295), .Z(c[4431]) );
XNOR U22159 ( .A(a[4431]), .B(c4431), .Z(n13295) );
XOR U22160 ( .A(c4432), .B(n13296), .Z(c4433) );
ANDN U22161 ( .B(n13297), .A(n13298), .Z(n13296) );
XOR U22162 ( .A(c4432), .B(b[4432]), .Z(n13297) );
XNOR U22163 ( .A(b[4432]), .B(n13298), .Z(c[4432]) );
XNOR U22164 ( .A(a[4432]), .B(c4432), .Z(n13298) );
XOR U22165 ( .A(c4433), .B(n13299), .Z(c4434) );
ANDN U22166 ( .B(n13300), .A(n13301), .Z(n13299) );
XOR U22167 ( .A(c4433), .B(b[4433]), .Z(n13300) );
XNOR U22168 ( .A(b[4433]), .B(n13301), .Z(c[4433]) );
XNOR U22169 ( .A(a[4433]), .B(c4433), .Z(n13301) );
XOR U22170 ( .A(c4434), .B(n13302), .Z(c4435) );
ANDN U22171 ( .B(n13303), .A(n13304), .Z(n13302) );
XOR U22172 ( .A(c4434), .B(b[4434]), .Z(n13303) );
XNOR U22173 ( .A(b[4434]), .B(n13304), .Z(c[4434]) );
XNOR U22174 ( .A(a[4434]), .B(c4434), .Z(n13304) );
XOR U22175 ( .A(c4435), .B(n13305), .Z(c4436) );
ANDN U22176 ( .B(n13306), .A(n13307), .Z(n13305) );
XOR U22177 ( .A(c4435), .B(b[4435]), .Z(n13306) );
XNOR U22178 ( .A(b[4435]), .B(n13307), .Z(c[4435]) );
XNOR U22179 ( .A(a[4435]), .B(c4435), .Z(n13307) );
XOR U22180 ( .A(c4436), .B(n13308), .Z(c4437) );
ANDN U22181 ( .B(n13309), .A(n13310), .Z(n13308) );
XOR U22182 ( .A(c4436), .B(b[4436]), .Z(n13309) );
XNOR U22183 ( .A(b[4436]), .B(n13310), .Z(c[4436]) );
XNOR U22184 ( .A(a[4436]), .B(c4436), .Z(n13310) );
XOR U22185 ( .A(c4437), .B(n13311), .Z(c4438) );
ANDN U22186 ( .B(n13312), .A(n13313), .Z(n13311) );
XOR U22187 ( .A(c4437), .B(b[4437]), .Z(n13312) );
XNOR U22188 ( .A(b[4437]), .B(n13313), .Z(c[4437]) );
XNOR U22189 ( .A(a[4437]), .B(c4437), .Z(n13313) );
XOR U22190 ( .A(c4438), .B(n13314), .Z(c4439) );
ANDN U22191 ( .B(n13315), .A(n13316), .Z(n13314) );
XOR U22192 ( .A(c4438), .B(b[4438]), .Z(n13315) );
XNOR U22193 ( .A(b[4438]), .B(n13316), .Z(c[4438]) );
XNOR U22194 ( .A(a[4438]), .B(c4438), .Z(n13316) );
XOR U22195 ( .A(c4439), .B(n13317), .Z(c4440) );
ANDN U22196 ( .B(n13318), .A(n13319), .Z(n13317) );
XOR U22197 ( .A(c4439), .B(b[4439]), .Z(n13318) );
XNOR U22198 ( .A(b[4439]), .B(n13319), .Z(c[4439]) );
XNOR U22199 ( .A(a[4439]), .B(c4439), .Z(n13319) );
XOR U22200 ( .A(c4440), .B(n13320), .Z(c4441) );
ANDN U22201 ( .B(n13321), .A(n13322), .Z(n13320) );
XOR U22202 ( .A(c4440), .B(b[4440]), .Z(n13321) );
XNOR U22203 ( .A(b[4440]), .B(n13322), .Z(c[4440]) );
XNOR U22204 ( .A(a[4440]), .B(c4440), .Z(n13322) );
XOR U22205 ( .A(c4441), .B(n13323), .Z(c4442) );
ANDN U22206 ( .B(n13324), .A(n13325), .Z(n13323) );
XOR U22207 ( .A(c4441), .B(b[4441]), .Z(n13324) );
XNOR U22208 ( .A(b[4441]), .B(n13325), .Z(c[4441]) );
XNOR U22209 ( .A(a[4441]), .B(c4441), .Z(n13325) );
XOR U22210 ( .A(c4442), .B(n13326), .Z(c4443) );
ANDN U22211 ( .B(n13327), .A(n13328), .Z(n13326) );
XOR U22212 ( .A(c4442), .B(b[4442]), .Z(n13327) );
XNOR U22213 ( .A(b[4442]), .B(n13328), .Z(c[4442]) );
XNOR U22214 ( .A(a[4442]), .B(c4442), .Z(n13328) );
XOR U22215 ( .A(c4443), .B(n13329), .Z(c4444) );
ANDN U22216 ( .B(n13330), .A(n13331), .Z(n13329) );
XOR U22217 ( .A(c4443), .B(b[4443]), .Z(n13330) );
XNOR U22218 ( .A(b[4443]), .B(n13331), .Z(c[4443]) );
XNOR U22219 ( .A(a[4443]), .B(c4443), .Z(n13331) );
XOR U22220 ( .A(c4444), .B(n13332), .Z(c4445) );
ANDN U22221 ( .B(n13333), .A(n13334), .Z(n13332) );
XOR U22222 ( .A(c4444), .B(b[4444]), .Z(n13333) );
XNOR U22223 ( .A(b[4444]), .B(n13334), .Z(c[4444]) );
XNOR U22224 ( .A(a[4444]), .B(c4444), .Z(n13334) );
XOR U22225 ( .A(c4445), .B(n13335), .Z(c4446) );
ANDN U22226 ( .B(n13336), .A(n13337), .Z(n13335) );
XOR U22227 ( .A(c4445), .B(b[4445]), .Z(n13336) );
XNOR U22228 ( .A(b[4445]), .B(n13337), .Z(c[4445]) );
XNOR U22229 ( .A(a[4445]), .B(c4445), .Z(n13337) );
XOR U22230 ( .A(c4446), .B(n13338), .Z(c4447) );
ANDN U22231 ( .B(n13339), .A(n13340), .Z(n13338) );
XOR U22232 ( .A(c4446), .B(b[4446]), .Z(n13339) );
XNOR U22233 ( .A(b[4446]), .B(n13340), .Z(c[4446]) );
XNOR U22234 ( .A(a[4446]), .B(c4446), .Z(n13340) );
XOR U22235 ( .A(c4447), .B(n13341), .Z(c4448) );
ANDN U22236 ( .B(n13342), .A(n13343), .Z(n13341) );
XOR U22237 ( .A(c4447), .B(b[4447]), .Z(n13342) );
XNOR U22238 ( .A(b[4447]), .B(n13343), .Z(c[4447]) );
XNOR U22239 ( .A(a[4447]), .B(c4447), .Z(n13343) );
XOR U22240 ( .A(c4448), .B(n13344), .Z(c4449) );
ANDN U22241 ( .B(n13345), .A(n13346), .Z(n13344) );
XOR U22242 ( .A(c4448), .B(b[4448]), .Z(n13345) );
XNOR U22243 ( .A(b[4448]), .B(n13346), .Z(c[4448]) );
XNOR U22244 ( .A(a[4448]), .B(c4448), .Z(n13346) );
XOR U22245 ( .A(c4449), .B(n13347), .Z(c4450) );
ANDN U22246 ( .B(n13348), .A(n13349), .Z(n13347) );
XOR U22247 ( .A(c4449), .B(b[4449]), .Z(n13348) );
XNOR U22248 ( .A(b[4449]), .B(n13349), .Z(c[4449]) );
XNOR U22249 ( .A(a[4449]), .B(c4449), .Z(n13349) );
XOR U22250 ( .A(c4450), .B(n13350), .Z(c4451) );
ANDN U22251 ( .B(n13351), .A(n13352), .Z(n13350) );
XOR U22252 ( .A(c4450), .B(b[4450]), .Z(n13351) );
XNOR U22253 ( .A(b[4450]), .B(n13352), .Z(c[4450]) );
XNOR U22254 ( .A(a[4450]), .B(c4450), .Z(n13352) );
XOR U22255 ( .A(c4451), .B(n13353), .Z(c4452) );
ANDN U22256 ( .B(n13354), .A(n13355), .Z(n13353) );
XOR U22257 ( .A(c4451), .B(b[4451]), .Z(n13354) );
XNOR U22258 ( .A(b[4451]), .B(n13355), .Z(c[4451]) );
XNOR U22259 ( .A(a[4451]), .B(c4451), .Z(n13355) );
XOR U22260 ( .A(c4452), .B(n13356), .Z(c4453) );
ANDN U22261 ( .B(n13357), .A(n13358), .Z(n13356) );
XOR U22262 ( .A(c4452), .B(b[4452]), .Z(n13357) );
XNOR U22263 ( .A(b[4452]), .B(n13358), .Z(c[4452]) );
XNOR U22264 ( .A(a[4452]), .B(c4452), .Z(n13358) );
XOR U22265 ( .A(c4453), .B(n13359), .Z(c4454) );
ANDN U22266 ( .B(n13360), .A(n13361), .Z(n13359) );
XOR U22267 ( .A(c4453), .B(b[4453]), .Z(n13360) );
XNOR U22268 ( .A(b[4453]), .B(n13361), .Z(c[4453]) );
XNOR U22269 ( .A(a[4453]), .B(c4453), .Z(n13361) );
XOR U22270 ( .A(c4454), .B(n13362), .Z(c4455) );
ANDN U22271 ( .B(n13363), .A(n13364), .Z(n13362) );
XOR U22272 ( .A(c4454), .B(b[4454]), .Z(n13363) );
XNOR U22273 ( .A(b[4454]), .B(n13364), .Z(c[4454]) );
XNOR U22274 ( .A(a[4454]), .B(c4454), .Z(n13364) );
XOR U22275 ( .A(c4455), .B(n13365), .Z(c4456) );
ANDN U22276 ( .B(n13366), .A(n13367), .Z(n13365) );
XOR U22277 ( .A(c4455), .B(b[4455]), .Z(n13366) );
XNOR U22278 ( .A(b[4455]), .B(n13367), .Z(c[4455]) );
XNOR U22279 ( .A(a[4455]), .B(c4455), .Z(n13367) );
XOR U22280 ( .A(c4456), .B(n13368), .Z(c4457) );
ANDN U22281 ( .B(n13369), .A(n13370), .Z(n13368) );
XOR U22282 ( .A(c4456), .B(b[4456]), .Z(n13369) );
XNOR U22283 ( .A(b[4456]), .B(n13370), .Z(c[4456]) );
XNOR U22284 ( .A(a[4456]), .B(c4456), .Z(n13370) );
XOR U22285 ( .A(c4457), .B(n13371), .Z(c4458) );
ANDN U22286 ( .B(n13372), .A(n13373), .Z(n13371) );
XOR U22287 ( .A(c4457), .B(b[4457]), .Z(n13372) );
XNOR U22288 ( .A(b[4457]), .B(n13373), .Z(c[4457]) );
XNOR U22289 ( .A(a[4457]), .B(c4457), .Z(n13373) );
XOR U22290 ( .A(c4458), .B(n13374), .Z(c4459) );
ANDN U22291 ( .B(n13375), .A(n13376), .Z(n13374) );
XOR U22292 ( .A(c4458), .B(b[4458]), .Z(n13375) );
XNOR U22293 ( .A(b[4458]), .B(n13376), .Z(c[4458]) );
XNOR U22294 ( .A(a[4458]), .B(c4458), .Z(n13376) );
XOR U22295 ( .A(c4459), .B(n13377), .Z(c4460) );
ANDN U22296 ( .B(n13378), .A(n13379), .Z(n13377) );
XOR U22297 ( .A(c4459), .B(b[4459]), .Z(n13378) );
XNOR U22298 ( .A(b[4459]), .B(n13379), .Z(c[4459]) );
XNOR U22299 ( .A(a[4459]), .B(c4459), .Z(n13379) );
XOR U22300 ( .A(c4460), .B(n13380), .Z(c4461) );
ANDN U22301 ( .B(n13381), .A(n13382), .Z(n13380) );
XOR U22302 ( .A(c4460), .B(b[4460]), .Z(n13381) );
XNOR U22303 ( .A(b[4460]), .B(n13382), .Z(c[4460]) );
XNOR U22304 ( .A(a[4460]), .B(c4460), .Z(n13382) );
XOR U22305 ( .A(c4461), .B(n13383), .Z(c4462) );
ANDN U22306 ( .B(n13384), .A(n13385), .Z(n13383) );
XOR U22307 ( .A(c4461), .B(b[4461]), .Z(n13384) );
XNOR U22308 ( .A(b[4461]), .B(n13385), .Z(c[4461]) );
XNOR U22309 ( .A(a[4461]), .B(c4461), .Z(n13385) );
XOR U22310 ( .A(c4462), .B(n13386), .Z(c4463) );
ANDN U22311 ( .B(n13387), .A(n13388), .Z(n13386) );
XOR U22312 ( .A(c4462), .B(b[4462]), .Z(n13387) );
XNOR U22313 ( .A(b[4462]), .B(n13388), .Z(c[4462]) );
XNOR U22314 ( .A(a[4462]), .B(c4462), .Z(n13388) );
XOR U22315 ( .A(c4463), .B(n13389), .Z(c4464) );
ANDN U22316 ( .B(n13390), .A(n13391), .Z(n13389) );
XOR U22317 ( .A(c4463), .B(b[4463]), .Z(n13390) );
XNOR U22318 ( .A(b[4463]), .B(n13391), .Z(c[4463]) );
XNOR U22319 ( .A(a[4463]), .B(c4463), .Z(n13391) );
XOR U22320 ( .A(c4464), .B(n13392), .Z(c4465) );
ANDN U22321 ( .B(n13393), .A(n13394), .Z(n13392) );
XOR U22322 ( .A(c4464), .B(b[4464]), .Z(n13393) );
XNOR U22323 ( .A(b[4464]), .B(n13394), .Z(c[4464]) );
XNOR U22324 ( .A(a[4464]), .B(c4464), .Z(n13394) );
XOR U22325 ( .A(c4465), .B(n13395), .Z(c4466) );
ANDN U22326 ( .B(n13396), .A(n13397), .Z(n13395) );
XOR U22327 ( .A(c4465), .B(b[4465]), .Z(n13396) );
XNOR U22328 ( .A(b[4465]), .B(n13397), .Z(c[4465]) );
XNOR U22329 ( .A(a[4465]), .B(c4465), .Z(n13397) );
XOR U22330 ( .A(c4466), .B(n13398), .Z(c4467) );
ANDN U22331 ( .B(n13399), .A(n13400), .Z(n13398) );
XOR U22332 ( .A(c4466), .B(b[4466]), .Z(n13399) );
XNOR U22333 ( .A(b[4466]), .B(n13400), .Z(c[4466]) );
XNOR U22334 ( .A(a[4466]), .B(c4466), .Z(n13400) );
XOR U22335 ( .A(c4467), .B(n13401), .Z(c4468) );
ANDN U22336 ( .B(n13402), .A(n13403), .Z(n13401) );
XOR U22337 ( .A(c4467), .B(b[4467]), .Z(n13402) );
XNOR U22338 ( .A(b[4467]), .B(n13403), .Z(c[4467]) );
XNOR U22339 ( .A(a[4467]), .B(c4467), .Z(n13403) );
XOR U22340 ( .A(c4468), .B(n13404), .Z(c4469) );
ANDN U22341 ( .B(n13405), .A(n13406), .Z(n13404) );
XOR U22342 ( .A(c4468), .B(b[4468]), .Z(n13405) );
XNOR U22343 ( .A(b[4468]), .B(n13406), .Z(c[4468]) );
XNOR U22344 ( .A(a[4468]), .B(c4468), .Z(n13406) );
XOR U22345 ( .A(c4469), .B(n13407), .Z(c4470) );
ANDN U22346 ( .B(n13408), .A(n13409), .Z(n13407) );
XOR U22347 ( .A(c4469), .B(b[4469]), .Z(n13408) );
XNOR U22348 ( .A(b[4469]), .B(n13409), .Z(c[4469]) );
XNOR U22349 ( .A(a[4469]), .B(c4469), .Z(n13409) );
XOR U22350 ( .A(c4470), .B(n13410), .Z(c4471) );
ANDN U22351 ( .B(n13411), .A(n13412), .Z(n13410) );
XOR U22352 ( .A(c4470), .B(b[4470]), .Z(n13411) );
XNOR U22353 ( .A(b[4470]), .B(n13412), .Z(c[4470]) );
XNOR U22354 ( .A(a[4470]), .B(c4470), .Z(n13412) );
XOR U22355 ( .A(c4471), .B(n13413), .Z(c4472) );
ANDN U22356 ( .B(n13414), .A(n13415), .Z(n13413) );
XOR U22357 ( .A(c4471), .B(b[4471]), .Z(n13414) );
XNOR U22358 ( .A(b[4471]), .B(n13415), .Z(c[4471]) );
XNOR U22359 ( .A(a[4471]), .B(c4471), .Z(n13415) );
XOR U22360 ( .A(c4472), .B(n13416), .Z(c4473) );
ANDN U22361 ( .B(n13417), .A(n13418), .Z(n13416) );
XOR U22362 ( .A(c4472), .B(b[4472]), .Z(n13417) );
XNOR U22363 ( .A(b[4472]), .B(n13418), .Z(c[4472]) );
XNOR U22364 ( .A(a[4472]), .B(c4472), .Z(n13418) );
XOR U22365 ( .A(c4473), .B(n13419), .Z(c4474) );
ANDN U22366 ( .B(n13420), .A(n13421), .Z(n13419) );
XOR U22367 ( .A(c4473), .B(b[4473]), .Z(n13420) );
XNOR U22368 ( .A(b[4473]), .B(n13421), .Z(c[4473]) );
XNOR U22369 ( .A(a[4473]), .B(c4473), .Z(n13421) );
XOR U22370 ( .A(c4474), .B(n13422), .Z(c4475) );
ANDN U22371 ( .B(n13423), .A(n13424), .Z(n13422) );
XOR U22372 ( .A(c4474), .B(b[4474]), .Z(n13423) );
XNOR U22373 ( .A(b[4474]), .B(n13424), .Z(c[4474]) );
XNOR U22374 ( .A(a[4474]), .B(c4474), .Z(n13424) );
XOR U22375 ( .A(c4475), .B(n13425), .Z(c4476) );
ANDN U22376 ( .B(n13426), .A(n13427), .Z(n13425) );
XOR U22377 ( .A(c4475), .B(b[4475]), .Z(n13426) );
XNOR U22378 ( .A(b[4475]), .B(n13427), .Z(c[4475]) );
XNOR U22379 ( .A(a[4475]), .B(c4475), .Z(n13427) );
XOR U22380 ( .A(c4476), .B(n13428), .Z(c4477) );
ANDN U22381 ( .B(n13429), .A(n13430), .Z(n13428) );
XOR U22382 ( .A(c4476), .B(b[4476]), .Z(n13429) );
XNOR U22383 ( .A(b[4476]), .B(n13430), .Z(c[4476]) );
XNOR U22384 ( .A(a[4476]), .B(c4476), .Z(n13430) );
XOR U22385 ( .A(c4477), .B(n13431), .Z(c4478) );
ANDN U22386 ( .B(n13432), .A(n13433), .Z(n13431) );
XOR U22387 ( .A(c4477), .B(b[4477]), .Z(n13432) );
XNOR U22388 ( .A(b[4477]), .B(n13433), .Z(c[4477]) );
XNOR U22389 ( .A(a[4477]), .B(c4477), .Z(n13433) );
XOR U22390 ( .A(c4478), .B(n13434), .Z(c4479) );
ANDN U22391 ( .B(n13435), .A(n13436), .Z(n13434) );
XOR U22392 ( .A(c4478), .B(b[4478]), .Z(n13435) );
XNOR U22393 ( .A(b[4478]), .B(n13436), .Z(c[4478]) );
XNOR U22394 ( .A(a[4478]), .B(c4478), .Z(n13436) );
XOR U22395 ( .A(c4479), .B(n13437), .Z(c4480) );
ANDN U22396 ( .B(n13438), .A(n13439), .Z(n13437) );
XOR U22397 ( .A(c4479), .B(b[4479]), .Z(n13438) );
XNOR U22398 ( .A(b[4479]), .B(n13439), .Z(c[4479]) );
XNOR U22399 ( .A(a[4479]), .B(c4479), .Z(n13439) );
XOR U22400 ( .A(c4480), .B(n13440), .Z(c4481) );
ANDN U22401 ( .B(n13441), .A(n13442), .Z(n13440) );
XOR U22402 ( .A(c4480), .B(b[4480]), .Z(n13441) );
XNOR U22403 ( .A(b[4480]), .B(n13442), .Z(c[4480]) );
XNOR U22404 ( .A(a[4480]), .B(c4480), .Z(n13442) );
XOR U22405 ( .A(c4481), .B(n13443), .Z(c4482) );
ANDN U22406 ( .B(n13444), .A(n13445), .Z(n13443) );
XOR U22407 ( .A(c4481), .B(b[4481]), .Z(n13444) );
XNOR U22408 ( .A(b[4481]), .B(n13445), .Z(c[4481]) );
XNOR U22409 ( .A(a[4481]), .B(c4481), .Z(n13445) );
XOR U22410 ( .A(c4482), .B(n13446), .Z(c4483) );
ANDN U22411 ( .B(n13447), .A(n13448), .Z(n13446) );
XOR U22412 ( .A(c4482), .B(b[4482]), .Z(n13447) );
XNOR U22413 ( .A(b[4482]), .B(n13448), .Z(c[4482]) );
XNOR U22414 ( .A(a[4482]), .B(c4482), .Z(n13448) );
XOR U22415 ( .A(c4483), .B(n13449), .Z(c4484) );
ANDN U22416 ( .B(n13450), .A(n13451), .Z(n13449) );
XOR U22417 ( .A(c4483), .B(b[4483]), .Z(n13450) );
XNOR U22418 ( .A(b[4483]), .B(n13451), .Z(c[4483]) );
XNOR U22419 ( .A(a[4483]), .B(c4483), .Z(n13451) );
XOR U22420 ( .A(c4484), .B(n13452), .Z(c4485) );
ANDN U22421 ( .B(n13453), .A(n13454), .Z(n13452) );
XOR U22422 ( .A(c4484), .B(b[4484]), .Z(n13453) );
XNOR U22423 ( .A(b[4484]), .B(n13454), .Z(c[4484]) );
XNOR U22424 ( .A(a[4484]), .B(c4484), .Z(n13454) );
XOR U22425 ( .A(c4485), .B(n13455), .Z(c4486) );
ANDN U22426 ( .B(n13456), .A(n13457), .Z(n13455) );
XOR U22427 ( .A(c4485), .B(b[4485]), .Z(n13456) );
XNOR U22428 ( .A(b[4485]), .B(n13457), .Z(c[4485]) );
XNOR U22429 ( .A(a[4485]), .B(c4485), .Z(n13457) );
XOR U22430 ( .A(c4486), .B(n13458), .Z(c4487) );
ANDN U22431 ( .B(n13459), .A(n13460), .Z(n13458) );
XOR U22432 ( .A(c4486), .B(b[4486]), .Z(n13459) );
XNOR U22433 ( .A(b[4486]), .B(n13460), .Z(c[4486]) );
XNOR U22434 ( .A(a[4486]), .B(c4486), .Z(n13460) );
XOR U22435 ( .A(c4487), .B(n13461), .Z(c4488) );
ANDN U22436 ( .B(n13462), .A(n13463), .Z(n13461) );
XOR U22437 ( .A(c4487), .B(b[4487]), .Z(n13462) );
XNOR U22438 ( .A(b[4487]), .B(n13463), .Z(c[4487]) );
XNOR U22439 ( .A(a[4487]), .B(c4487), .Z(n13463) );
XOR U22440 ( .A(c4488), .B(n13464), .Z(c4489) );
ANDN U22441 ( .B(n13465), .A(n13466), .Z(n13464) );
XOR U22442 ( .A(c4488), .B(b[4488]), .Z(n13465) );
XNOR U22443 ( .A(b[4488]), .B(n13466), .Z(c[4488]) );
XNOR U22444 ( .A(a[4488]), .B(c4488), .Z(n13466) );
XOR U22445 ( .A(c4489), .B(n13467), .Z(c4490) );
ANDN U22446 ( .B(n13468), .A(n13469), .Z(n13467) );
XOR U22447 ( .A(c4489), .B(b[4489]), .Z(n13468) );
XNOR U22448 ( .A(b[4489]), .B(n13469), .Z(c[4489]) );
XNOR U22449 ( .A(a[4489]), .B(c4489), .Z(n13469) );
XOR U22450 ( .A(c4490), .B(n13470), .Z(c4491) );
ANDN U22451 ( .B(n13471), .A(n13472), .Z(n13470) );
XOR U22452 ( .A(c4490), .B(b[4490]), .Z(n13471) );
XNOR U22453 ( .A(b[4490]), .B(n13472), .Z(c[4490]) );
XNOR U22454 ( .A(a[4490]), .B(c4490), .Z(n13472) );
XOR U22455 ( .A(c4491), .B(n13473), .Z(c4492) );
ANDN U22456 ( .B(n13474), .A(n13475), .Z(n13473) );
XOR U22457 ( .A(c4491), .B(b[4491]), .Z(n13474) );
XNOR U22458 ( .A(b[4491]), .B(n13475), .Z(c[4491]) );
XNOR U22459 ( .A(a[4491]), .B(c4491), .Z(n13475) );
XOR U22460 ( .A(c4492), .B(n13476), .Z(c4493) );
ANDN U22461 ( .B(n13477), .A(n13478), .Z(n13476) );
XOR U22462 ( .A(c4492), .B(b[4492]), .Z(n13477) );
XNOR U22463 ( .A(b[4492]), .B(n13478), .Z(c[4492]) );
XNOR U22464 ( .A(a[4492]), .B(c4492), .Z(n13478) );
XOR U22465 ( .A(c4493), .B(n13479), .Z(c4494) );
ANDN U22466 ( .B(n13480), .A(n13481), .Z(n13479) );
XOR U22467 ( .A(c4493), .B(b[4493]), .Z(n13480) );
XNOR U22468 ( .A(b[4493]), .B(n13481), .Z(c[4493]) );
XNOR U22469 ( .A(a[4493]), .B(c4493), .Z(n13481) );
XOR U22470 ( .A(c4494), .B(n13482), .Z(c4495) );
ANDN U22471 ( .B(n13483), .A(n13484), .Z(n13482) );
XOR U22472 ( .A(c4494), .B(b[4494]), .Z(n13483) );
XNOR U22473 ( .A(b[4494]), .B(n13484), .Z(c[4494]) );
XNOR U22474 ( .A(a[4494]), .B(c4494), .Z(n13484) );
XOR U22475 ( .A(c4495), .B(n13485), .Z(c4496) );
ANDN U22476 ( .B(n13486), .A(n13487), .Z(n13485) );
XOR U22477 ( .A(c4495), .B(b[4495]), .Z(n13486) );
XNOR U22478 ( .A(b[4495]), .B(n13487), .Z(c[4495]) );
XNOR U22479 ( .A(a[4495]), .B(c4495), .Z(n13487) );
XOR U22480 ( .A(c4496), .B(n13488), .Z(c4497) );
ANDN U22481 ( .B(n13489), .A(n13490), .Z(n13488) );
XOR U22482 ( .A(c4496), .B(b[4496]), .Z(n13489) );
XNOR U22483 ( .A(b[4496]), .B(n13490), .Z(c[4496]) );
XNOR U22484 ( .A(a[4496]), .B(c4496), .Z(n13490) );
XOR U22485 ( .A(c4497), .B(n13491), .Z(c4498) );
ANDN U22486 ( .B(n13492), .A(n13493), .Z(n13491) );
XOR U22487 ( .A(c4497), .B(b[4497]), .Z(n13492) );
XNOR U22488 ( .A(b[4497]), .B(n13493), .Z(c[4497]) );
XNOR U22489 ( .A(a[4497]), .B(c4497), .Z(n13493) );
XOR U22490 ( .A(c4498), .B(n13494), .Z(c4499) );
ANDN U22491 ( .B(n13495), .A(n13496), .Z(n13494) );
XOR U22492 ( .A(c4498), .B(b[4498]), .Z(n13495) );
XNOR U22493 ( .A(b[4498]), .B(n13496), .Z(c[4498]) );
XNOR U22494 ( .A(a[4498]), .B(c4498), .Z(n13496) );
XOR U22495 ( .A(c4499), .B(n13497), .Z(c4500) );
ANDN U22496 ( .B(n13498), .A(n13499), .Z(n13497) );
XOR U22497 ( .A(c4499), .B(b[4499]), .Z(n13498) );
XNOR U22498 ( .A(b[4499]), .B(n13499), .Z(c[4499]) );
XNOR U22499 ( .A(a[4499]), .B(c4499), .Z(n13499) );
XOR U22500 ( .A(c4500), .B(n13500), .Z(c4501) );
ANDN U22501 ( .B(n13501), .A(n13502), .Z(n13500) );
XOR U22502 ( .A(c4500), .B(b[4500]), .Z(n13501) );
XNOR U22503 ( .A(b[4500]), .B(n13502), .Z(c[4500]) );
XNOR U22504 ( .A(a[4500]), .B(c4500), .Z(n13502) );
XOR U22505 ( .A(c4501), .B(n13503), .Z(c4502) );
ANDN U22506 ( .B(n13504), .A(n13505), .Z(n13503) );
XOR U22507 ( .A(c4501), .B(b[4501]), .Z(n13504) );
XNOR U22508 ( .A(b[4501]), .B(n13505), .Z(c[4501]) );
XNOR U22509 ( .A(a[4501]), .B(c4501), .Z(n13505) );
XOR U22510 ( .A(c4502), .B(n13506), .Z(c4503) );
ANDN U22511 ( .B(n13507), .A(n13508), .Z(n13506) );
XOR U22512 ( .A(c4502), .B(b[4502]), .Z(n13507) );
XNOR U22513 ( .A(b[4502]), .B(n13508), .Z(c[4502]) );
XNOR U22514 ( .A(a[4502]), .B(c4502), .Z(n13508) );
XOR U22515 ( .A(c4503), .B(n13509), .Z(c4504) );
ANDN U22516 ( .B(n13510), .A(n13511), .Z(n13509) );
XOR U22517 ( .A(c4503), .B(b[4503]), .Z(n13510) );
XNOR U22518 ( .A(b[4503]), .B(n13511), .Z(c[4503]) );
XNOR U22519 ( .A(a[4503]), .B(c4503), .Z(n13511) );
XOR U22520 ( .A(c4504), .B(n13512), .Z(c4505) );
ANDN U22521 ( .B(n13513), .A(n13514), .Z(n13512) );
XOR U22522 ( .A(c4504), .B(b[4504]), .Z(n13513) );
XNOR U22523 ( .A(b[4504]), .B(n13514), .Z(c[4504]) );
XNOR U22524 ( .A(a[4504]), .B(c4504), .Z(n13514) );
XOR U22525 ( .A(c4505), .B(n13515), .Z(c4506) );
ANDN U22526 ( .B(n13516), .A(n13517), .Z(n13515) );
XOR U22527 ( .A(c4505), .B(b[4505]), .Z(n13516) );
XNOR U22528 ( .A(b[4505]), .B(n13517), .Z(c[4505]) );
XNOR U22529 ( .A(a[4505]), .B(c4505), .Z(n13517) );
XOR U22530 ( .A(c4506), .B(n13518), .Z(c4507) );
ANDN U22531 ( .B(n13519), .A(n13520), .Z(n13518) );
XOR U22532 ( .A(c4506), .B(b[4506]), .Z(n13519) );
XNOR U22533 ( .A(b[4506]), .B(n13520), .Z(c[4506]) );
XNOR U22534 ( .A(a[4506]), .B(c4506), .Z(n13520) );
XOR U22535 ( .A(c4507), .B(n13521), .Z(c4508) );
ANDN U22536 ( .B(n13522), .A(n13523), .Z(n13521) );
XOR U22537 ( .A(c4507), .B(b[4507]), .Z(n13522) );
XNOR U22538 ( .A(b[4507]), .B(n13523), .Z(c[4507]) );
XNOR U22539 ( .A(a[4507]), .B(c4507), .Z(n13523) );
XOR U22540 ( .A(c4508), .B(n13524), .Z(c4509) );
ANDN U22541 ( .B(n13525), .A(n13526), .Z(n13524) );
XOR U22542 ( .A(c4508), .B(b[4508]), .Z(n13525) );
XNOR U22543 ( .A(b[4508]), .B(n13526), .Z(c[4508]) );
XNOR U22544 ( .A(a[4508]), .B(c4508), .Z(n13526) );
XOR U22545 ( .A(c4509), .B(n13527), .Z(c4510) );
ANDN U22546 ( .B(n13528), .A(n13529), .Z(n13527) );
XOR U22547 ( .A(c4509), .B(b[4509]), .Z(n13528) );
XNOR U22548 ( .A(b[4509]), .B(n13529), .Z(c[4509]) );
XNOR U22549 ( .A(a[4509]), .B(c4509), .Z(n13529) );
XOR U22550 ( .A(c4510), .B(n13530), .Z(c4511) );
ANDN U22551 ( .B(n13531), .A(n13532), .Z(n13530) );
XOR U22552 ( .A(c4510), .B(b[4510]), .Z(n13531) );
XNOR U22553 ( .A(b[4510]), .B(n13532), .Z(c[4510]) );
XNOR U22554 ( .A(a[4510]), .B(c4510), .Z(n13532) );
XOR U22555 ( .A(c4511), .B(n13533), .Z(c4512) );
ANDN U22556 ( .B(n13534), .A(n13535), .Z(n13533) );
XOR U22557 ( .A(c4511), .B(b[4511]), .Z(n13534) );
XNOR U22558 ( .A(b[4511]), .B(n13535), .Z(c[4511]) );
XNOR U22559 ( .A(a[4511]), .B(c4511), .Z(n13535) );
XOR U22560 ( .A(c4512), .B(n13536), .Z(c4513) );
ANDN U22561 ( .B(n13537), .A(n13538), .Z(n13536) );
XOR U22562 ( .A(c4512), .B(b[4512]), .Z(n13537) );
XNOR U22563 ( .A(b[4512]), .B(n13538), .Z(c[4512]) );
XNOR U22564 ( .A(a[4512]), .B(c4512), .Z(n13538) );
XOR U22565 ( .A(c4513), .B(n13539), .Z(c4514) );
ANDN U22566 ( .B(n13540), .A(n13541), .Z(n13539) );
XOR U22567 ( .A(c4513), .B(b[4513]), .Z(n13540) );
XNOR U22568 ( .A(b[4513]), .B(n13541), .Z(c[4513]) );
XNOR U22569 ( .A(a[4513]), .B(c4513), .Z(n13541) );
XOR U22570 ( .A(c4514), .B(n13542), .Z(c4515) );
ANDN U22571 ( .B(n13543), .A(n13544), .Z(n13542) );
XOR U22572 ( .A(c4514), .B(b[4514]), .Z(n13543) );
XNOR U22573 ( .A(b[4514]), .B(n13544), .Z(c[4514]) );
XNOR U22574 ( .A(a[4514]), .B(c4514), .Z(n13544) );
XOR U22575 ( .A(c4515), .B(n13545), .Z(c4516) );
ANDN U22576 ( .B(n13546), .A(n13547), .Z(n13545) );
XOR U22577 ( .A(c4515), .B(b[4515]), .Z(n13546) );
XNOR U22578 ( .A(b[4515]), .B(n13547), .Z(c[4515]) );
XNOR U22579 ( .A(a[4515]), .B(c4515), .Z(n13547) );
XOR U22580 ( .A(c4516), .B(n13548), .Z(c4517) );
ANDN U22581 ( .B(n13549), .A(n13550), .Z(n13548) );
XOR U22582 ( .A(c4516), .B(b[4516]), .Z(n13549) );
XNOR U22583 ( .A(b[4516]), .B(n13550), .Z(c[4516]) );
XNOR U22584 ( .A(a[4516]), .B(c4516), .Z(n13550) );
XOR U22585 ( .A(c4517), .B(n13551), .Z(c4518) );
ANDN U22586 ( .B(n13552), .A(n13553), .Z(n13551) );
XOR U22587 ( .A(c4517), .B(b[4517]), .Z(n13552) );
XNOR U22588 ( .A(b[4517]), .B(n13553), .Z(c[4517]) );
XNOR U22589 ( .A(a[4517]), .B(c4517), .Z(n13553) );
XOR U22590 ( .A(c4518), .B(n13554), .Z(c4519) );
ANDN U22591 ( .B(n13555), .A(n13556), .Z(n13554) );
XOR U22592 ( .A(c4518), .B(b[4518]), .Z(n13555) );
XNOR U22593 ( .A(b[4518]), .B(n13556), .Z(c[4518]) );
XNOR U22594 ( .A(a[4518]), .B(c4518), .Z(n13556) );
XOR U22595 ( .A(c4519), .B(n13557), .Z(c4520) );
ANDN U22596 ( .B(n13558), .A(n13559), .Z(n13557) );
XOR U22597 ( .A(c4519), .B(b[4519]), .Z(n13558) );
XNOR U22598 ( .A(b[4519]), .B(n13559), .Z(c[4519]) );
XNOR U22599 ( .A(a[4519]), .B(c4519), .Z(n13559) );
XOR U22600 ( .A(c4520), .B(n13560), .Z(c4521) );
ANDN U22601 ( .B(n13561), .A(n13562), .Z(n13560) );
XOR U22602 ( .A(c4520), .B(b[4520]), .Z(n13561) );
XNOR U22603 ( .A(b[4520]), .B(n13562), .Z(c[4520]) );
XNOR U22604 ( .A(a[4520]), .B(c4520), .Z(n13562) );
XOR U22605 ( .A(c4521), .B(n13563), .Z(c4522) );
ANDN U22606 ( .B(n13564), .A(n13565), .Z(n13563) );
XOR U22607 ( .A(c4521), .B(b[4521]), .Z(n13564) );
XNOR U22608 ( .A(b[4521]), .B(n13565), .Z(c[4521]) );
XNOR U22609 ( .A(a[4521]), .B(c4521), .Z(n13565) );
XOR U22610 ( .A(c4522), .B(n13566), .Z(c4523) );
ANDN U22611 ( .B(n13567), .A(n13568), .Z(n13566) );
XOR U22612 ( .A(c4522), .B(b[4522]), .Z(n13567) );
XNOR U22613 ( .A(b[4522]), .B(n13568), .Z(c[4522]) );
XNOR U22614 ( .A(a[4522]), .B(c4522), .Z(n13568) );
XOR U22615 ( .A(c4523), .B(n13569), .Z(c4524) );
ANDN U22616 ( .B(n13570), .A(n13571), .Z(n13569) );
XOR U22617 ( .A(c4523), .B(b[4523]), .Z(n13570) );
XNOR U22618 ( .A(b[4523]), .B(n13571), .Z(c[4523]) );
XNOR U22619 ( .A(a[4523]), .B(c4523), .Z(n13571) );
XOR U22620 ( .A(c4524), .B(n13572), .Z(c4525) );
ANDN U22621 ( .B(n13573), .A(n13574), .Z(n13572) );
XOR U22622 ( .A(c4524), .B(b[4524]), .Z(n13573) );
XNOR U22623 ( .A(b[4524]), .B(n13574), .Z(c[4524]) );
XNOR U22624 ( .A(a[4524]), .B(c4524), .Z(n13574) );
XOR U22625 ( .A(c4525), .B(n13575), .Z(c4526) );
ANDN U22626 ( .B(n13576), .A(n13577), .Z(n13575) );
XOR U22627 ( .A(c4525), .B(b[4525]), .Z(n13576) );
XNOR U22628 ( .A(b[4525]), .B(n13577), .Z(c[4525]) );
XNOR U22629 ( .A(a[4525]), .B(c4525), .Z(n13577) );
XOR U22630 ( .A(c4526), .B(n13578), .Z(c4527) );
ANDN U22631 ( .B(n13579), .A(n13580), .Z(n13578) );
XOR U22632 ( .A(c4526), .B(b[4526]), .Z(n13579) );
XNOR U22633 ( .A(b[4526]), .B(n13580), .Z(c[4526]) );
XNOR U22634 ( .A(a[4526]), .B(c4526), .Z(n13580) );
XOR U22635 ( .A(c4527), .B(n13581), .Z(c4528) );
ANDN U22636 ( .B(n13582), .A(n13583), .Z(n13581) );
XOR U22637 ( .A(c4527), .B(b[4527]), .Z(n13582) );
XNOR U22638 ( .A(b[4527]), .B(n13583), .Z(c[4527]) );
XNOR U22639 ( .A(a[4527]), .B(c4527), .Z(n13583) );
XOR U22640 ( .A(c4528), .B(n13584), .Z(c4529) );
ANDN U22641 ( .B(n13585), .A(n13586), .Z(n13584) );
XOR U22642 ( .A(c4528), .B(b[4528]), .Z(n13585) );
XNOR U22643 ( .A(b[4528]), .B(n13586), .Z(c[4528]) );
XNOR U22644 ( .A(a[4528]), .B(c4528), .Z(n13586) );
XOR U22645 ( .A(c4529), .B(n13587), .Z(c4530) );
ANDN U22646 ( .B(n13588), .A(n13589), .Z(n13587) );
XOR U22647 ( .A(c4529), .B(b[4529]), .Z(n13588) );
XNOR U22648 ( .A(b[4529]), .B(n13589), .Z(c[4529]) );
XNOR U22649 ( .A(a[4529]), .B(c4529), .Z(n13589) );
XOR U22650 ( .A(c4530), .B(n13590), .Z(c4531) );
ANDN U22651 ( .B(n13591), .A(n13592), .Z(n13590) );
XOR U22652 ( .A(c4530), .B(b[4530]), .Z(n13591) );
XNOR U22653 ( .A(b[4530]), .B(n13592), .Z(c[4530]) );
XNOR U22654 ( .A(a[4530]), .B(c4530), .Z(n13592) );
XOR U22655 ( .A(c4531), .B(n13593), .Z(c4532) );
ANDN U22656 ( .B(n13594), .A(n13595), .Z(n13593) );
XOR U22657 ( .A(c4531), .B(b[4531]), .Z(n13594) );
XNOR U22658 ( .A(b[4531]), .B(n13595), .Z(c[4531]) );
XNOR U22659 ( .A(a[4531]), .B(c4531), .Z(n13595) );
XOR U22660 ( .A(c4532), .B(n13596), .Z(c4533) );
ANDN U22661 ( .B(n13597), .A(n13598), .Z(n13596) );
XOR U22662 ( .A(c4532), .B(b[4532]), .Z(n13597) );
XNOR U22663 ( .A(b[4532]), .B(n13598), .Z(c[4532]) );
XNOR U22664 ( .A(a[4532]), .B(c4532), .Z(n13598) );
XOR U22665 ( .A(c4533), .B(n13599), .Z(c4534) );
ANDN U22666 ( .B(n13600), .A(n13601), .Z(n13599) );
XOR U22667 ( .A(c4533), .B(b[4533]), .Z(n13600) );
XNOR U22668 ( .A(b[4533]), .B(n13601), .Z(c[4533]) );
XNOR U22669 ( .A(a[4533]), .B(c4533), .Z(n13601) );
XOR U22670 ( .A(c4534), .B(n13602), .Z(c4535) );
ANDN U22671 ( .B(n13603), .A(n13604), .Z(n13602) );
XOR U22672 ( .A(c4534), .B(b[4534]), .Z(n13603) );
XNOR U22673 ( .A(b[4534]), .B(n13604), .Z(c[4534]) );
XNOR U22674 ( .A(a[4534]), .B(c4534), .Z(n13604) );
XOR U22675 ( .A(c4535), .B(n13605), .Z(c4536) );
ANDN U22676 ( .B(n13606), .A(n13607), .Z(n13605) );
XOR U22677 ( .A(c4535), .B(b[4535]), .Z(n13606) );
XNOR U22678 ( .A(b[4535]), .B(n13607), .Z(c[4535]) );
XNOR U22679 ( .A(a[4535]), .B(c4535), .Z(n13607) );
XOR U22680 ( .A(c4536), .B(n13608), .Z(c4537) );
ANDN U22681 ( .B(n13609), .A(n13610), .Z(n13608) );
XOR U22682 ( .A(c4536), .B(b[4536]), .Z(n13609) );
XNOR U22683 ( .A(b[4536]), .B(n13610), .Z(c[4536]) );
XNOR U22684 ( .A(a[4536]), .B(c4536), .Z(n13610) );
XOR U22685 ( .A(c4537), .B(n13611), .Z(c4538) );
ANDN U22686 ( .B(n13612), .A(n13613), .Z(n13611) );
XOR U22687 ( .A(c4537), .B(b[4537]), .Z(n13612) );
XNOR U22688 ( .A(b[4537]), .B(n13613), .Z(c[4537]) );
XNOR U22689 ( .A(a[4537]), .B(c4537), .Z(n13613) );
XOR U22690 ( .A(c4538), .B(n13614), .Z(c4539) );
ANDN U22691 ( .B(n13615), .A(n13616), .Z(n13614) );
XOR U22692 ( .A(c4538), .B(b[4538]), .Z(n13615) );
XNOR U22693 ( .A(b[4538]), .B(n13616), .Z(c[4538]) );
XNOR U22694 ( .A(a[4538]), .B(c4538), .Z(n13616) );
XOR U22695 ( .A(c4539), .B(n13617), .Z(c4540) );
ANDN U22696 ( .B(n13618), .A(n13619), .Z(n13617) );
XOR U22697 ( .A(c4539), .B(b[4539]), .Z(n13618) );
XNOR U22698 ( .A(b[4539]), .B(n13619), .Z(c[4539]) );
XNOR U22699 ( .A(a[4539]), .B(c4539), .Z(n13619) );
XOR U22700 ( .A(c4540), .B(n13620), .Z(c4541) );
ANDN U22701 ( .B(n13621), .A(n13622), .Z(n13620) );
XOR U22702 ( .A(c4540), .B(b[4540]), .Z(n13621) );
XNOR U22703 ( .A(b[4540]), .B(n13622), .Z(c[4540]) );
XNOR U22704 ( .A(a[4540]), .B(c4540), .Z(n13622) );
XOR U22705 ( .A(c4541), .B(n13623), .Z(c4542) );
ANDN U22706 ( .B(n13624), .A(n13625), .Z(n13623) );
XOR U22707 ( .A(c4541), .B(b[4541]), .Z(n13624) );
XNOR U22708 ( .A(b[4541]), .B(n13625), .Z(c[4541]) );
XNOR U22709 ( .A(a[4541]), .B(c4541), .Z(n13625) );
XOR U22710 ( .A(c4542), .B(n13626), .Z(c4543) );
ANDN U22711 ( .B(n13627), .A(n13628), .Z(n13626) );
XOR U22712 ( .A(c4542), .B(b[4542]), .Z(n13627) );
XNOR U22713 ( .A(b[4542]), .B(n13628), .Z(c[4542]) );
XNOR U22714 ( .A(a[4542]), .B(c4542), .Z(n13628) );
XOR U22715 ( .A(c4543), .B(n13629), .Z(c4544) );
ANDN U22716 ( .B(n13630), .A(n13631), .Z(n13629) );
XOR U22717 ( .A(c4543), .B(b[4543]), .Z(n13630) );
XNOR U22718 ( .A(b[4543]), .B(n13631), .Z(c[4543]) );
XNOR U22719 ( .A(a[4543]), .B(c4543), .Z(n13631) );
XOR U22720 ( .A(c4544), .B(n13632), .Z(c4545) );
ANDN U22721 ( .B(n13633), .A(n13634), .Z(n13632) );
XOR U22722 ( .A(c4544), .B(b[4544]), .Z(n13633) );
XNOR U22723 ( .A(b[4544]), .B(n13634), .Z(c[4544]) );
XNOR U22724 ( .A(a[4544]), .B(c4544), .Z(n13634) );
XOR U22725 ( .A(c4545), .B(n13635), .Z(c4546) );
ANDN U22726 ( .B(n13636), .A(n13637), .Z(n13635) );
XOR U22727 ( .A(c4545), .B(b[4545]), .Z(n13636) );
XNOR U22728 ( .A(b[4545]), .B(n13637), .Z(c[4545]) );
XNOR U22729 ( .A(a[4545]), .B(c4545), .Z(n13637) );
XOR U22730 ( .A(c4546), .B(n13638), .Z(c4547) );
ANDN U22731 ( .B(n13639), .A(n13640), .Z(n13638) );
XOR U22732 ( .A(c4546), .B(b[4546]), .Z(n13639) );
XNOR U22733 ( .A(b[4546]), .B(n13640), .Z(c[4546]) );
XNOR U22734 ( .A(a[4546]), .B(c4546), .Z(n13640) );
XOR U22735 ( .A(c4547), .B(n13641), .Z(c4548) );
ANDN U22736 ( .B(n13642), .A(n13643), .Z(n13641) );
XOR U22737 ( .A(c4547), .B(b[4547]), .Z(n13642) );
XNOR U22738 ( .A(b[4547]), .B(n13643), .Z(c[4547]) );
XNOR U22739 ( .A(a[4547]), .B(c4547), .Z(n13643) );
XOR U22740 ( .A(c4548), .B(n13644), .Z(c4549) );
ANDN U22741 ( .B(n13645), .A(n13646), .Z(n13644) );
XOR U22742 ( .A(c4548), .B(b[4548]), .Z(n13645) );
XNOR U22743 ( .A(b[4548]), .B(n13646), .Z(c[4548]) );
XNOR U22744 ( .A(a[4548]), .B(c4548), .Z(n13646) );
XOR U22745 ( .A(c4549), .B(n13647), .Z(c4550) );
ANDN U22746 ( .B(n13648), .A(n13649), .Z(n13647) );
XOR U22747 ( .A(c4549), .B(b[4549]), .Z(n13648) );
XNOR U22748 ( .A(b[4549]), .B(n13649), .Z(c[4549]) );
XNOR U22749 ( .A(a[4549]), .B(c4549), .Z(n13649) );
XOR U22750 ( .A(c4550), .B(n13650), .Z(c4551) );
ANDN U22751 ( .B(n13651), .A(n13652), .Z(n13650) );
XOR U22752 ( .A(c4550), .B(b[4550]), .Z(n13651) );
XNOR U22753 ( .A(b[4550]), .B(n13652), .Z(c[4550]) );
XNOR U22754 ( .A(a[4550]), .B(c4550), .Z(n13652) );
XOR U22755 ( .A(c4551), .B(n13653), .Z(c4552) );
ANDN U22756 ( .B(n13654), .A(n13655), .Z(n13653) );
XOR U22757 ( .A(c4551), .B(b[4551]), .Z(n13654) );
XNOR U22758 ( .A(b[4551]), .B(n13655), .Z(c[4551]) );
XNOR U22759 ( .A(a[4551]), .B(c4551), .Z(n13655) );
XOR U22760 ( .A(c4552), .B(n13656), .Z(c4553) );
ANDN U22761 ( .B(n13657), .A(n13658), .Z(n13656) );
XOR U22762 ( .A(c4552), .B(b[4552]), .Z(n13657) );
XNOR U22763 ( .A(b[4552]), .B(n13658), .Z(c[4552]) );
XNOR U22764 ( .A(a[4552]), .B(c4552), .Z(n13658) );
XOR U22765 ( .A(c4553), .B(n13659), .Z(c4554) );
ANDN U22766 ( .B(n13660), .A(n13661), .Z(n13659) );
XOR U22767 ( .A(c4553), .B(b[4553]), .Z(n13660) );
XNOR U22768 ( .A(b[4553]), .B(n13661), .Z(c[4553]) );
XNOR U22769 ( .A(a[4553]), .B(c4553), .Z(n13661) );
XOR U22770 ( .A(c4554), .B(n13662), .Z(c4555) );
ANDN U22771 ( .B(n13663), .A(n13664), .Z(n13662) );
XOR U22772 ( .A(c4554), .B(b[4554]), .Z(n13663) );
XNOR U22773 ( .A(b[4554]), .B(n13664), .Z(c[4554]) );
XNOR U22774 ( .A(a[4554]), .B(c4554), .Z(n13664) );
XOR U22775 ( .A(c4555), .B(n13665), .Z(c4556) );
ANDN U22776 ( .B(n13666), .A(n13667), .Z(n13665) );
XOR U22777 ( .A(c4555), .B(b[4555]), .Z(n13666) );
XNOR U22778 ( .A(b[4555]), .B(n13667), .Z(c[4555]) );
XNOR U22779 ( .A(a[4555]), .B(c4555), .Z(n13667) );
XOR U22780 ( .A(c4556), .B(n13668), .Z(c4557) );
ANDN U22781 ( .B(n13669), .A(n13670), .Z(n13668) );
XOR U22782 ( .A(c4556), .B(b[4556]), .Z(n13669) );
XNOR U22783 ( .A(b[4556]), .B(n13670), .Z(c[4556]) );
XNOR U22784 ( .A(a[4556]), .B(c4556), .Z(n13670) );
XOR U22785 ( .A(c4557), .B(n13671), .Z(c4558) );
ANDN U22786 ( .B(n13672), .A(n13673), .Z(n13671) );
XOR U22787 ( .A(c4557), .B(b[4557]), .Z(n13672) );
XNOR U22788 ( .A(b[4557]), .B(n13673), .Z(c[4557]) );
XNOR U22789 ( .A(a[4557]), .B(c4557), .Z(n13673) );
XOR U22790 ( .A(c4558), .B(n13674), .Z(c4559) );
ANDN U22791 ( .B(n13675), .A(n13676), .Z(n13674) );
XOR U22792 ( .A(c4558), .B(b[4558]), .Z(n13675) );
XNOR U22793 ( .A(b[4558]), .B(n13676), .Z(c[4558]) );
XNOR U22794 ( .A(a[4558]), .B(c4558), .Z(n13676) );
XOR U22795 ( .A(c4559), .B(n13677), .Z(c4560) );
ANDN U22796 ( .B(n13678), .A(n13679), .Z(n13677) );
XOR U22797 ( .A(c4559), .B(b[4559]), .Z(n13678) );
XNOR U22798 ( .A(b[4559]), .B(n13679), .Z(c[4559]) );
XNOR U22799 ( .A(a[4559]), .B(c4559), .Z(n13679) );
XOR U22800 ( .A(c4560), .B(n13680), .Z(c4561) );
ANDN U22801 ( .B(n13681), .A(n13682), .Z(n13680) );
XOR U22802 ( .A(c4560), .B(b[4560]), .Z(n13681) );
XNOR U22803 ( .A(b[4560]), .B(n13682), .Z(c[4560]) );
XNOR U22804 ( .A(a[4560]), .B(c4560), .Z(n13682) );
XOR U22805 ( .A(c4561), .B(n13683), .Z(c4562) );
ANDN U22806 ( .B(n13684), .A(n13685), .Z(n13683) );
XOR U22807 ( .A(c4561), .B(b[4561]), .Z(n13684) );
XNOR U22808 ( .A(b[4561]), .B(n13685), .Z(c[4561]) );
XNOR U22809 ( .A(a[4561]), .B(c4561), .Z(n13685) );
XOR U22810 ( .A(c4562), .B(n13686), .Z(c4563) );
ANDN U22811 ( .B(n13687), .A(n13688), .Z(n13686) );
XOR U22812 ( .A(c4562), .B(b[4562]), .Z(n13687) );
XNOR U22813 ( .A(b[4562]), .B(n13688), .Z(c[4562]) );
XNOR U22814 ( .A(a[4562]), .B(c4562), .Z(n13688) );
XOR U22815 ( .A(c4563), .B(n13689), .Z(c4564) );
ANDN U22816 ( .B(n13690), .A(n13691), .Z(n13689) );
XOR U22817 ( .A(c4563), .B(b[4563]), .Z(n13690) );
XNOR U22818 ( .A(b[4563]), .B(n13691), .Z(c[4563]) );
XNOR U22819 ( .A(a[4563]), .B(c4563), .Z(n13691) );
XOR U22820 ( .A(c4564), .B(n13692), .Z(c4565) );
ANDN U22821 ( .B(n13693), .A(n13694), .Z(n13692) );
XOR U22822 ( .A(c4564), .B(b[4564]), .Z(n13693) );
XNOR U22823 ( .A(b[4564]), .B(n13694), .Z(c[4564]) );
XNOR U22824 ( .A(a[4564]), .B(c4564), .Z(n13694) );
XOR U22825 ( .A(c4565), .B(n13695), .Z(c4566) );
ANDN U22826 ( .B(n13696), .A(n13697), .Z(n13695) );
XOR U22827 ( .A(c4565), .B(b[4565]), .Z(n13696) );
XNOR U22828 ( .A(b[4565]), .B(n13697), .Z(c[4565]) );
XNOR U22829 ( .A(a[4565]), .B(c4565), .Z(n13697) );
XOR U22830 ( .A(c4566), .B(n13698), .Z(c4567) );
ANDN U22831 ( .B(n13699), .A(n13700), .Z(n13698) );
XOR U22832 ( .A(c4566), .B(b[4566]), .Z(n13699) );
XNOR U22833 ( .A(b[4566]), .B(n13700), .Z(c[4566]) );
XNOR U22834 ( .A(a[4566]), .B(c4566), .Z(n13700) );
XOR U22835 ( .A(c4567), .B(n13701), .Z(c4568) );
ANDN U22836 ( .B(n13702), .A(n13703), .Z(n13701) );
XOR U22837 ( .A(c4567), .B(b[4567]), .Z(n13702) );
XNOR U22838 ( .A(b[4567]), .B(n13703), .Z(c[4567]) );
XNOR U22839 ( .A(a[4567]), .B(c4567), .Z(n13703) );
XOR U22840 ( .A(c4568), .B(n13704), .Z(c4569) );
ANDN U22841 ( .B(n13705), .A(n13706), .Z(n13704) );
XOR U22842 ( .A(c4568), .B(b[4568]), .Z(n13705) );
XNOR U22843 ( .A(b[4568]), .B(n13706), .Z(c[4568]) );
XNOR U22844 ( .A(a[4568]), .B(c4568), .Z(n13706) );
XOR U22845 ( .A(c4569), .B(n13707), .Z(c4570) );
ANDN U22846 ( .B(n13708), .A(n13709), .Z(n13707) );
XOR U22847 ( .A(c4569), .B(b[4569]), .Z(n13708) );
XNOR U22848 ( .A(b[4569]), .B(n13709), .Z(c[4569]) );
XNOR U22849 ( .A(a[4569]), .B(c4569), .Z(n13709) );
XOR U22850 ( .A(c4570), .B(n13710), .Z(c4571) );
ANDN U22851 ( .B(n13711), .A(n13712), .Z(n13710) );
XOR U22852 ( .A(c4570), .B(b[4570]), .Z(n13711) );
XNOR U22853 ( .A(b[4570]), .B(n13712), .Z(c[4570]) );
XNOR U22854 ( .A(a[4570]), .B(c4570), .Z(n13712) );
XOR U22855 ( .A(c4571), .B(n13713), .Z(c4572) );
ANDN U22856 ( .B(n13714), .A(n13715), .Z(n13713) );
XOR U22857 ( .A(c4571), .B(b[4571]), .Z(n13714) );
XNOR U22858 ( .A(b[4571]), .B(n13715), .Z(c[4571]) );
XNOR U22859 ( .A(a[4571]), .B(c4571), .Z(n13715) );
XOR U22860 ( .A(c4572), .B(n13716), .Z(c4573) );
ANDN U22861 ( .B(n13717), .A(n13718), .Z(n13716) );
XOR U22862 ( .A(c4572), .B(b[4572]), .Z(n13717) );
XNOR U22863 ( .A(b[4572]), .B(n13718), .Z(c[4572]) );
XNOR U22864 ( .A(a[4572]), .B(c4572), .Z(n13718) );
XOR U22865 ( .A(c4573), .B(n13719), .Z(c4574) );
ANDN U22866 ( .B(n13720), .A(n13721), .Z(n13719) );
XOR U22867 ( .A(c4573), .B(b[4573]), .Z(n13720) );
XNOR U22868 ( .A(b[4573]), .B(n13721), .Z(c[4573]) );
XNOR U22869 ( .A(a[4573]), .B(c4573), .Z(n13721) );
XOR U22870 ( .A(c4574), .B(n13722), .Z(c4575) );
ANDN U22871 ( .B(n13723), .A(n13724), .Z(n13722) );
XOR U22872 ( .A(c4574), .B(b[4574]), .Z(n13723) );
XNOR U22873 ( .A(b[4574]), .B(n13724), .Z(c[4574]) );
XNOR U22874 ( .A(a[4574]), .B(c4574), .Z(n13724) );
XOR U22875 ( .A(c4575), .B(n13725), .Z(c4576) );
ANDN U22876 ( .B(n13726), .A(n13727), .Z(n13725) );
XOR U22877 ( .A(c4575), .B(b[4575]), .Z(n13726) );
XNOR U22878 ( .A(b[4575]), .B(n13727), .Z(c[4575]) );
XNOR U22879 ( .A(a[4575]), .B(c4575), .Z(n13727) );
XOR U22880 ( .A(c4576), .B(n13728), .Z(c4577) );
ANDN U22881 ( .B(n13729), .A(n13730), .Z(n13728) );
XOR U22882 ( .A(c4576), .B(b[4576]), .Z(n13729) );
XNOR U22883 ( .A(b[4576]), .B(n13730), .Z(c[4576]) );
XNOR U22884 ( .A(a[4576]), .B(c4576), .Z(n13730) );
XOR U22885 ( .A(c4577), .B(n13731), .Z(c4578) );
ANDN U22886 ( .B(n13732), .A(n13733), .Z(n13731) );
XOR U22887 ( .A(c4577), .B(b[4577]), .Z(n13732) );
XNOR U22888 ( .A(b[4577]), .B(n13733), .Z(c[4577]) );
XNOR U22889 ( .A(a[4577]), .B(c4577), .Z(n13733) );
XOR U22890 ( .A(c4578), .B(n13734), .Z(c4579) );
ANDN U22891 ( .B(n13735), .A(n13736), .Z(n13734) );
XOR U22892 ( .A(c4578), .B(b[4578]), .Z(n13735) );
XNOR U22893 ( .A(b[4578]), .B(n13736), .Z(c[4578]) );
XNOR U22894 ( .A(a[4578]), .B(c4578), .Z(n13736) );
XOR U22895 ( .A(c4579), .B(n13737), .Z(c4580) );
ANDN U22896 ( .B(n13738), .A(n13739), .Z(n13737) );
XOR U22897 ( .A(c4579), .B(b[4579]), .Z(n13738) );
XNOR U22898 ( .A(b[4579]), .B(n13739), .Z(c[4579]) );
XNOR U22899 ( .A(a[4579]), .B(c4579), .Z(n13739) );
XOR U22900 ( .A(c4580), .B(n13740), .Z(c4581) );
ANDN U22901 ( .B(n13741), .A(n13742), .Z(n13740) );
XOR U22902 ( .A(c4580), .B(b[4580]), .Z(n13741) );
XNOR U22903 ( .A(b[4580]), .B(n13742), .Z(c[4580]) );
XNOR U22904 ( .A(a[4580]), .B(c4580), .Z(n13742) );
XOR U22905 ( .A(c4581), .B(n13743), .Z(c4582) );
ANDN U22906 ( .B(n13744), .A(n13745), .Z(n13743) );
XOR U22907 ( .A(c4581), .B(b[4581]), .Z(n13744) );
XNOR U22908 ( .A(b[4581]), .B(n13745), .Z(c[4581]) );
XNOR U22909 ( .A(a[4581]), .B(c4581), .Z(n13745) );
XOR U22910 ( .A(c4582), .B(n13746), .Z(c4583) );
ANDN U22911 ( .B(n13747), .A(n13748), .Z(n13746) );
XOR U22912 ( .A(c4582), .B(b[4582]), .Z(n13747) );
XNOR U22913 ( .A(b[4582]), .B(n13748), .Z(c[4582]) );
XNOR U22914 ( .A(a[4582]), .B(c4582), .Z(n13748) );
XOR U22915 ( .A(c4583), .B(n13749), .Z(c4584) );
ANDN U22916 ( .B(n13750), .A(n13751), .Z(n13749) );
XOR U22917 ( .A(c4583), .B(b[4583]), .Z(n13750) );
XNOR U22918 ( .A(b[4583]), .B(n13751), .Z(c[4583]) );
XNOR U22919 ( .A(a[4583]), .B(c4583), .Z(n13751) );
XOR U22920 ( .A(c4584), .B(n13752), .Z(c4585) );
ANDN U22921 ( .B(n13753), .A(n13754), .Z(n13752) );
XOR U22922 ( .A(c4584), .B(b[4584]), .Z(n13753) );
XNOR U22923 ( .A(b[4584]), .B(n13754), .Z(c[4584]) );
XNOR U22924 ( .A(a[4584]), .B(c4584), .Z(n13754) );
XOR U22925 ( .A(c4585), .B(n13755), .Z(c4586) );
ANDN U22926 ( .B(n13756), .A(n13757), .Z(n13755) );
XOR U22927 ( .A(c4585), .B(b[4585]), .Z(n13756) );
XNOR U22928 ( .A(b[4585]), .B(n13757), .Z(c[4585]) );
XNOR U22929 ( .A(a[4585]), .B(c4585), .Z(n13757) );
XOR U22930 ( .A(c4586), .B(n13758), .Z(c4587) );
ANDN U22931 ( .B(n13759), .A(n13760), .Z(n13758) );
XOR U22932 ( .A(c4586), .B(b[4586]), .Z(n13759) );
XNOR U22933 ( .A(b[4586]), .B(n13760), .Z(c[4586]) );
XNOR U22934 ( .A(a[4586]), .B(c4586), .Z(n13760) );
XOR U22935 ( .A(c4587), .B(n13761), .Z(c4588) );
ANDN U22936 ( .B(n13762), .A(n13763), .Z(n13761) );
XOR U22937 ( .A(c4587), .B(b[4587]), .Z(n13762) );
XNOR U22938 ( .A(b[4587]), .B(n13763), .Z(c[4587]) );
XNOR U22939 ( .A(a[4587]), .B(c4587), .Z(n13763) );
XOR U22940 ( .A(c4588), .B(n13764), .Z(c4589) );
ANDN U22941 ( .B(n13765), .A(n13766), .Z(n13764) );
XOR U22942 ( .A(c4588), .B(b[4588]), .Z(n13765) );
XNOR U22943 ( .A(b[4588]), .B(n13766), .Z(c[4588]) );
XNOR U22944 ( .A(a[4588]), .B(c4588), .Z(n13766) );
XOR U22945 ( .A(c4589), .B(n13767), .Z(c4590) );
ANDN U22946 ( .B(n13768), .A(n13769), .Z(n13767) );
XOR U22947 ( .A(c4589), .B(b[4589]), .Z(n13768) );
XNOR U22948 ( .A(b[4589]), .B(n13769), .Z(c[4589]) );
XNOR U22949 ( .A(a[4589]), .B(c4589), .Z(n13769) );
XOR U22950 ( .A(c4590), .B(n13770), .Z(c4591) );
ANDN U22951 ( .B(n13771), .A(n13772), .Z(n13770) );
XOR U22952 ( .A(c4590), .B(b[4590]), .Z(n13771) );
XNOR U22953 ( .A(b[4590]), .B(n13772), .Z(c[4590]) );
XNOR U22954 ( .A(a[4590]), .B(c4590), .Z(n13772) );
XOR U22955 ( .A(c4591), .B(n13773), .Z(c4592) );
ANDN U22956 ( .B(n13774), .A(n13775), .Z(n13773) );
XOR U22957 ( .A(c4591), .B(b[4591]), .Z(n13774) );
XNOR U22958 ( .A(b[4591]), .B(n13775), .Z(c[4591]) );
XNOR U22959 ( .A(a[4591]), .B(c4591), .Z(n13775) );
XOR U22960 ( .A(c4592), .B(n13776), .Z(c4593) );
ANDN U22961 ( .B(n13777), .A(n13778), .Z(n13776) );
XOR U22962 ( .A(c4592), .B(b[4592]), .Z(n13777) );
XNOR U22963 ( .A(b[4592]), .B(n13778), .Z(c[4592]) );
XNOR U22964 ( .A(a[4592]), .B(c4592), .Z(n13778) );
XOR U22965 ( .A(c4593), .B(n13779), .Z(c4594) );
ANDN U22966 ( .B(n13780), .A(n13781), .Z(n13779) );
XOR U22967 ( .A(c4593), .B(b[4593]), .Z(n13780) );
XNOR U22968 ( .A(b[4593]), .B(n13781), .Z(c[4593]) );
XNOR U22969 ( .A(a[4593]), .B(c4593), .Z(n13781) );
XOR U22970 ( .A(c4594), .B(n13782), .Z(c4595) );
ANDN U22971 ( .B(n13783), .A(n13784), .Z(n13782) );
XOR U22972 ( .A(c4594), .B(b[4594]), .Z(n13783) );
XNOR U22973 ( .A(b[4594]), .B(n13784), .Z(c[4594]) );
XNOR U22974 ( .A(a[4594]), .B(c4594), .Z(n13784) );
XOR U22975 ( .A(c4595), .B(n13785), .Z(c4596) );
ANDN U22976 ( .B(n13786), .A(n13787), .Z(n13785) );
XOR U22977 ( .A(c4595), .B(b[4595]), .Z(n13786) );
XNOR U22978 ( .A(b[4595]), .B(n13787), .Z(c[4595]) );
XNOR U22979 ( .A(a[4595]), .B(c4595), .Z(n13787) );
XOR U22980 ( .A(c4596), .B(n13788), .Z(c4597) );
ANDN U22981 ( .B(n13789), .A(n13790), .Z(n13788) );
XOR U22982 ( .A(c4596), .B(b[4596]), .Z(n13789) );
XNOR U22983 ( .A(b[4596]), .B(n13790), .Z(c[4596]) );
XNOR U22984 ( .A(a[4596]), .B(c4596), .Z(n13790) );
XOR U22985 ( .A(c4597), .B(n13791), .Z(c4598) );
ANDN U22986 ( .B(n13792), .A(n13793), .Z(n13791) );
XOR U22987 ( .A(c4597), .B(b[4597]), .Z(n13792) );
XNOR U22988 ( .A(b[4597]), .B(n13793), .Z(c[4597]) );
XNOR U22989 ( .A(a[4597]), .B(c4597), .Z(n13793) );
XOR U22990 ( .A(c4598), .B(n13794), .Z(c4599) );
ANDN U22991 ( .B(n13795), .A(n13796), .Z(n13794) );
XOR U22992 ( .A(c4598), .B(b[4598]), .Z(n13795) );
XNOR U22993 ( .A(b[4598]), .B(n13796), .Z(c[4598]) );
XNOR U22994 ( .A(a[4598]), .B(c4598), .Z(n13796) );
XOR U22995 ( .A(c4599), .B(n13797), .Z(c4600) );
ANDN U22996 ( .B(n13798), .A(n13799), .Z(n13797) );
XOR U22997 ( .A(c4599), .B(b[4599]), .Z(n13798) );
XNOR U22998 ( .A(b[4599]), .B(n13799), .Z(c[4599]) );
XNOR U22999 ( .A(a[4599]), .B(c4599), .Z(n13799) );
XOR U23000 ( .A(c4600), .B(n13800), .Z(c4601) );
ANDN U23001 ( .B(n13801), .A(n13802), .Z(n13800) );
XOR U23002 ( .A(c4600), .B(b[4600]), .Z(n13801) );
XNOR U23003 ( .A(b[4600]), .B(n13802), .Z(c[4600]) );
XNOR U23004 ( .A(a[4600]), .B(c4600), .Z(n13802) );
XOR U23005 ( .A(c4601), .B(n13803), .Z(c4602) );
ANDN U23006 ( .B(n13804), .A(n13805), .Z(n13803) );
XOR U23007 ( .A(c4601), .B(b[4601]), .Z(n13804) );
XNOR U23008 ( .A(b[4601]), .B(n13805), .Z(c[4601]) );
XNOR U23009 ( .A(a[4601]), .B(c4601), .Z(n13805) );
XOR U23010 ( .A(c4602), .B(n13806), .Z(c4603) );
ANDN U23011 ( .B(n13807), .A(n13808), .Z(n13806) );
XOR U23012 ( .A(c4602), .B(b[4602]), .Z(n13807) );
XNOR U23013 ( .A(b[4602]), .B(n13808), .Z(c[4602]) );
XNOR U23014 ( .A(a[4602]), .B(c4602), .Z(n13808) );
XOR U23015 ( .A(c4603), .B(n13809), .Z(c4604) );
ANDN U23016 ( .B(n13810), .A(n13811), .Z(n13809) );
XOR U23017 ( .A(c4603), .B(b[4603]), .Z(n13810) );
XNOR U23018 ( .A(b[4603]), .B(n13811), .Z(c[4603]) );
XNOR U23019 ( .A(a[4603]), .B(c4603), .Z(n13811) );
XOR U23020 ( .A(c4604), .B(n13812), .Z(c4605) );
ANDN U23021 ( .B(n13813), .A(n13814), .Z(n13812) );
XOR U23022 ( .A(c4604), .B(b[4604]), .Z(n13813) );
XNOR U23023 ( .A(b[4604]), .B(n13814), .Z(c[4604]) );
XNOR U23024 ( .A(a[4604]), .B(c4604), .Z(n13814) );
XOR U23025 ( .A(c4605), .B(n13815), .Z(c4606) );
ANDN U23026 ( .B(n13816), .A(n13817), .Z(n13815) );
XOR U23027 ( .A(c4605), .B(b[4605]), .Z(n13816) );
XNOR U23028 ( .A(b[4605]), .B(n13817), .Z(c[4605]) );
XNOR U23029 ( .A(a[4605]), .B(c4605), .Z(n13817) );
XOR U23030 ( .A(c4606), .B(n13818), .Z(c4607) );
ANDN U23031 ( .B(n13819), .A(n13820), .Z(n13818) );
XOR U23032 ( .A(c4606), .B(b[4606]), .Z(n13819) );
XNOR U23033 ( .A(b[4606]), .B(n13820), .Z(c[4606]) );
XNOR U23034 ( .A(a[4606]), .B(c4606), .Z(n13820) );
XOR U23035 ( .A(c4607), .B(n13821), .Z(c4608) );
ANDN U23036 ( .B(n13822), .A(n13823), .Z(n13821) );
XOR U23037 ( .A(c4607), .B(b[4607]), .Z(n13822) );
XNOR U23038 ( .A(b[4607]), .B(n13823), .Z(c[4607]) );
XNOR U23039 ( .A(a[4607]), .B(c4607), .Z(n13823) );
XOR U23040 ( .A(c4608), .B(n13824), .Z(c4609) );
ANDN U23041 ( .B(n13825), .A(n13826), .Z(n13824) );
XOR U23042 ( .A(c4608), .B(b[4608]), .Z(n13825) );
XNOR U23043 ( .A(b[4608]), .B(n13826), .Z(c[4608]) );
XNOR U23044 ( .A(a[4608]), .B(c4608), .Z(n13826) );
XOR U23045 ( .A(c4609), .B(n13827), .Z(c4610) );
ANDN U23046 ( .B(n13828), .A(n13829), .Z(n13827) );
XOR U23047 ( .A(c4609), .B(b[4609]), .Z(n13828) );
XNOR U23048 ( .A(b[4609]), .B(n13829), .Z(c[4609]) );
XNOR U23049 ( .A(a[4609]), .B(c4609), .Z(n13829) );
XOR U23050 ( .A(c4610), .B(n13830), .Z(c4611) );
ANDN U23051 ( .B(n13831), .A(n13832), .Z(n13830) );
XOR U23052 ( .A(c4610), .B(b[4610]), .Z(n13831) );
XNOR U23053 ( .A(b[4610]), .B(n13832), .Z(c[4610]) );
XNOR U23054 ( .A(a[4610]), .B(c4610), .Z(n13832) );
XOR U23055 ( .A(c4611), .B(n13833), .Z(c4612) );
ANDN U23056 ( .B(n13834), .A(n13835), .Z(n13833) );
XOR U23057 ( .A(c4611), .B(b[4611]), .Z(n13834) );
XNOR U23058 ( .A(b[4611]), .B(n13835), .Z(c[4611]) );
XNOR U23059 ( .A(a[4611]), .B(c4611), .Z(n13835) );
XOR U23060 ( .A(c4612), .B(n13836), .Z(c4613) );
ANDN U23061 ( .B(n13837), .A(n13838), .Z(n13836) );
XOR U23062 ( .A(c4612), .B(b[4612]), .Z(n13837) );
XNOR U23063 ( .A(b[4612]), .B(n13838), .Z(c[4612]) );
XNOR U23064 ( .A(a[4612]), .B(c4612), .Z(n13838) );
XOR U23065 ( .A(c4613), .B(n13839), .Z(c4614) );
ANDN U23066 ( .B(n13840), .A(n13841), .Z(n13839) );
XOR U23067 ( .A(c4613), .B(b[4613]), .Z(n13840) );
XNOR U23068 ( .A(b[4613]), .B(n13841), .Z(c[4613]) );
XNOR U23069 ( .A(a[4613]), .B(c4613), .Z(n13841) );
XOR U23070 ( .A(c4614), .B(n13842), .Z(c4615) );
ANDN U23071 ( .B(n13843), .A(n13844), .Z(n13842) );
XOR U23072 ( .A(c4614), .B(b[4614]), .Z(n13843) );
XNOR U23073 ( .A(b[4614]), .B(n13844), .Z(c[4614]) );
XNOR U23074 ( .A(a[4614]), .B(c4614), .Z(n13844) );
XOR U23075 ( .A(c4615), .B(n13845), .Z(c4616) );
ANDN U23076 ( .B(n13846), .A(n13847), .Z(n13845) );
XOR U23077 ( .A(c4615), .B(b[4615]), .Z(n13846) );
XNOR U23078 ( .A(b[4615]), .B(n13847), .Z(c[4615]) );
XNOR U23079 ( .A(a[4615]), .B(c4615), .Z(n13847) );
XOR U23080 ( .A(c4616), .B(n13848), .Z(c4617) );
ANDN U23081 ( .B(n13849), .A(n13850), .Z(n13848) );
XOR U23082 ( .A(c4616), .B(b[4616]), .Z(n13849) );
XNOR U23083 ( .A(b[4616]), .B(n13850), .Z(c[4616]) );
XNOR U23084 ( .A(a[4616]), .B(c4616), .Z(n13850) );
XOR U23085 ( .A(c4617), .B(n13851), .Z(c4618) );
ANDN U23086 ( .B(n13852), .A(n13853), .Z(n13851) );
XOR U23087 ( .A(c4617), .B(b[4617]), .Z(n13852) );
XNOR U23088 ( .A(b[4617]), .B(n13853), .Z(c[4617]) );
XNOR U23089 ( .A(a[4617]), .B(c4617), .Z(n13853) );
XOR U23090 ( .A(c4618), .B(n13854), .Z(c4619) );
ANDN U23091 ( .B(n13855), .A(n13856), .Z(n13854) );
XOR U23092 ( .A(c4618), .B(b[4618]), .Z(n13855) );
XNOR U23093 ( .A(b[4618]), .B(n13856), .Z(c[4618]) );
XNOR U23094 ( .A(a[4618]), .B(c4618), .Z(n13856) );
XOR U23095 ( .A(c4619), .B(n13857), .Z(c4620) );
ANDN U23096 ( .B(n13858), .A(n13859), .Z(n13857) );
XOR U23097 ( .A(c4619), .B(b[4619]), .Z(n13858) );
XNOR U23098 ( .A(b[4619]), .B(n13859), .Z(c[4619]) );
XNOR U23099 ( .A(a[4619]), .B(c4619), .Z(n13859) );
XOR U23100 ( .A(c4620), .B(n13860), .Z(c4621) );
ANDN U23101 ( .B(n13861), .A(n13862), .Z(n13860) );
XOR U23102 ( .A(c4620), .B(b[4620]), .Z(n13861) );
XNOR U23103 ( .A(b[4620]), .B(n13862), .Z(c[4620]) );
XNOR U23104 ( .A(a[4620]), .B(c4620), .Z(n13862) );
XOR U23105 ( .A(c4621), .B(n13863), .Z(c4622) );
ANDN U23106 ( .B(n13864), .A(n13865), .Z(n13863) );
XOR U23107 ( .A(c4621), .B(b[4621]), .Z(n13864) );
XNOR U23108 ( .A(b[4621]), .B(n13865), .Z(c[4621]) );
XNOR U23109 ( .A(a[4621]), .B(c4621), .Z(n13865) );
XOR U23110 ( .A(c4622), .B(n13866), .Z(c4623) );
ANDN U23111 ( .B(n13867), .A(n13868), .Z(n13866) );
XOR U23112 ( .A(c4622), .B(b[4622]), .Z(n13867) );
XNOR U23113 ( .A(b[4622]), .B(n13868), .Z(c[4622]) );
XNOR U23114 ( .A(a[4622]), .B(c4622), .Z(n13868) );
XOR U23115 ( .A(c4623), .B(n13869), .Z(c4624) );
ANDN U23116 ( .B(n13870), .A(n13871), .Z(n13869) );
XOR U23117 ( .A(c4623), .B(b[4623]), .Z(n13870) );
XNOR U23118 ( .A(b[4623]), .B(n13871), .Z(c[4623]) );
XNOR U23119 ( .A(a[4623]), .B(c4623), .Z(n13871) );
XOR U23120 ( .A(c4624), .B(n13872), .Z(c4625) );
ANDN U23121 ( .B(n13873), .A(n13874), .Z(n13872) );
XOR U23122 ( .A(c4624), .B(b[4624]), .Z(n13873) );
XNOR U23123 ( .A(b[4624]), .B(n13874), .Z(c[4624]) );
XNOR U23124 ( .A(a[4624]), .B(c4624), .Z(n13874) );
XOR U23125 ( .A(c4625), .B(n13875), .Z(c4626) );
ANDN U23126 ( .B(n13876), .A(n13877), .Z(n13875) );
XOR U23127 ( .A(c4625), .B(b[4625]), .Z(n13876) );
XNOR U23128 ( .A(b[4625]), .B(n13877), .Z(c[4625]) );
XNOR U23129 ( .A(a[4625]), .B(c4625), .Z(n13877) );
XOR U23130 ( .A(c4626), .B(n13878), .Z(c4627) );
ANDN U23131 ( .B(n13879), .A(n13880), .Z(n13878) );
XOR U23132 ( .A(c4626), .B(b[4626]), .Z(n13879) );
XNOR U23133 ( .A(b[4626]), .B(n13880), .Z(c[4626]) );
XNOR U23134 ( .A(a[4626]), .B(c4626), .Z(n13880) );
XOR U23135 ( .A(c4627), .B(n13881), .Z(c4628) );
ANDN U23136 ( .B(n13882), .A(n13883), .Z(n13881) );
XOR U23137 ( .A(c4627), .B(b[4627]), .Z(n13882) );
XNOR U23138 ( .A(b[4627]), .B(n13883), .Z(c[4627]) );
XNOR U23139 ( .A(a[4627]), .B(c4627), .Z(n13883) );
XOR U23140 ( .A(c4628), .B(n13884), .Z(c4629) );
ANDN U23141 ( .B(n13885), .A(n13886), .Z(n13884) );
XOR U23142 ( .A(c4628), .B(b[4628]), .Z(n13885) );
XNOR U23143 ( .A(b[4628]), .B(n13886), .Z(c[4628]) );
XNOR U23144 ( .A(a[4628]), .B(c4628), .Z(n13886) );
XOR U23145 ( .A(c4629), .B(n13887), .Z(c4630) );
ANDN U23146 ( .B(n13888), .A(n13889), .Z(n13887) );
XOR U23147 ( .A(c4629), .B(b[4629]), .Z(n13888) );
XNOR U23148 ( .A(b[4629]), .B(n13889), .Z(c[4629]) );
XNOR U23149 ( .A(a[4629]), .B(c4629), .Z(n13889) );
XOR U23150 ( .A(c4630), .B(n13890), .Z(c4631) );
ANDN U23151 ( .B(n13891), .A(n13892), .Z(n13890) );
XOR U23152 ( .A(c4630), .B(b[4630]), .Z(n13891) );
XNOR U23153 ( .A(b[4630]), .B(n13892), .Z(c[4630]) );
XNOR U23154 ( .A(a[4630]), .B(c4630), .Z(n13892) );
XOR U23155 ( .A(c4631), .B(n13893), .Z(c4632) );
ANDN U23156 ( .B(n13894), .A(n13895), .Z(n13893) );
XOR U23157 ( .A(c4631), .B(b[4631]), .Z(n13894) );
XNOR U23158 ( .A(b[4631]), .B(n13895), .Z(c[4631]) );
XNOR U23159 ( .A(a[4631]), .B(c4631), .Z(n13895) );
XOR U23160 ( .A(c4632), .B(n13896), .Z(c4633) );
ANDN U23161 ( .B(n13897), .A(n13898), .Z(n13896) );
XOR U23162 ( .A(c4632), .B(b[4632]), .Z(n13897) );
XNOR U23163 ( .A(b[4632]), .B(n13898), .Z(c[4632]) );
XNOR U23164 ( .A(a[4632]), .B(c4632), .Z(n13898) );
XOR U23165 ( .A(c4633), .B(n13899), .Z(c4634) );
ANDN U23166 ( .B(n13900), .A(n13901), .Z(n13899) );
XOR U23167 ( .A(c4633), .B(b[4633]), .Z(n13900) );
XNOR U23168 ( .A(b[4633]), .B(n13901), .Z(c[4633]) );
XNOR U23169 ( .A(a[4633]), .B(c4633), .Z(n13901) );
XOR U23170 ( .A(c4634), .B(n13902), .Z(c4635) );
ANDN U23171 ( .B(n13903), .A(n13904), .Z(n13902) );
XOR U23172 ( .A(c4634), .B(b[4634]), .Z(n13903) );
XNOR U23173 ( .A(b[4634]), .B(n13904), .Z(c[4634]) );
XNOR U23174 ( .A(a[4634]), .B(c4634), .Z(n13904) );
XOR U23175 ( .A(c4635), .B(n13905), .Z(c4636) );
ANDN U23176 ( .B(n13906), .A(n13907), .Z(n13905) );
XOR U23177 ( .A(c4635), .B(b[4635]), .Z(n13906) );
XNOR U23178 ( .A(b[4635]), .B(n13907), .Z(c[4635]) );
XNOR U23179 ( .A(a[4635]), .B(c4635), .Z(n13907) );
XOR U23180 ( .A(c4636), .B(n13908), .Z(c4637) );
ANDN U23181 ( .B(n13909), .A(n13910), .Z(n13908) );
XOR U23182 ( .A(c4636), .B(b[4636]), .Z(n13909) );
XNOR U23183 ( .A(b[4636]), .B(n13910), .Z(c[4636]) );
XNOR U23184 ( .A(a[4636]), .B(c4636), .Z(n13910) );
XOR U23185 ( .A(c4637), .B(n13911), .Z(c4638) );
ANDN U23186 ( .B(n13912), .A(n13913), .Z(n13911) );
XOR U23187 ( .A(c4637), .B(b[4637]), .Z(n13912) );
XNOR U23188 ( .A(b[4637]), .B(n13913), .Z(c[4637]) );
XNOR U23189 ( .A(a[4637]), .B(c4637), .Z(n13913) );
XOR U23190 ( .A(c4638), .B(n13914), .Z(c4639) );
ANDN U23191 ( .B(n13915), .A(n13916), .Z(n13914) );
XOR U23192 ( .A(c4638), .B(b[4638]), .Z(n13915) );
XNOR U23193 ( .A(b[4638]), .B(n13916), .Z(c[4638]) );
XNOR U23194 ( .A(a[4638]), .B(c4638), .Z(n13916) );
XOR U23195 ( .A(c4639), .B(n13917), .Z(c4640) );
ANDN U23196 ( .B(n13918), .A(n13919), .Z(n13917) );
XOR U23197 ( .A(c4639), .B(b[4639]), .Z(n13918) );
XNOR U23198 ( .A(b[4639]), .B(n13919), .Z(c[4639]) );
XNOR U23199 ( .A(a[4639]), .B(c4639), .Z(n13919) );
XOR U23200 ( .A(c4640), .B(n13920), .Z(c4641) );
ANDN U23201 ( .B(n13921), .A(n13922), .Z(n13920) );
XOR U23202 ( .A(c4640), .B(b[4640]), .Z(n13921) );
XNOR U23203 ( .A(b[4640]), .B(n13922), .Z(c[4640]) );
XNOR U23204 ( .A(a[4640]), .B(c4640), .Z(n13922) );
XOR U23205 ( .A(c4641), .B(n13923), .Z(c4642) );
ANDN U23206 ( .B(n13924), .A(n13925), .Z(n13923) );
XOR U23207 ( .A(c4641), .B(b[4641]), .Z(n13924) );
XNOR U23208 ( .A(b[4641]), .B(n13925), .Z(c[4641]) );
XNOR U23209 ( .A(a[4641]), .B(c4641), .Z(n13925) );
XOR U23210 ( .A(c4642), .B(n13926), .Z(c4643) );
ANDN U23211 ( .B(n13927), .A(n13928), .Z(n13926) );
XOR U23212 ( .A(c4642), .B(b[4642]), .Z(n13927) );
XNOR U23213 ( .A(b[4642]), .B(n13928), .Z(c[4642]) );
XNOR U23214 ( .A(a[4642]), .B(c4642), .Z(n13928) );
XOR U23215 ( .A(c4643), .B(n13929), .Z(c4644) );
ANDN U23216 ( .B(n13930), .A(n13931), .Z(n13929) );
XOR U23217 ( .A(c4643), .B(b[4643]), .Z(n13930) );
XNOR U23218 ( .A(b[4643]), .B(n13931), .Z(c[4643]) );
XNOR U23219 ( .A(a[4643]), .B(c4643), .Z(n13931) );
XOR U23220 ( .A(c4644), .B(n13932), .Z(c4645) );
ANDN U23221 ( .B(n13933), .A(n13934), .Z(n13932) );
XOR U23222 ( .A(c4644), .B(b[4644]), .Z(n13933) );
XNOR U23223 ( .A(b[4644]), .B(n13934), .Z(c[4644]) );
XNOR U23224 ( .A(a[4644]), .B(c4644), .Z(n13934) );
XOR U23225 ( .A(c4645), .B(n13935), .Z(c4646) );
ANDN U23226 ( .B(n13936), .A(n13937), .Z(n13935) );
XOR U23227 ( .A(c4645), .B(b[4645]), .Z(n13936) );
XNOR U23228 ( .A(b[4645]), .B(n13937), .Z(c[4645]) );
XNOR U23229 ( .A(a[4645]), .B(c4645), .Z(n13937) );
XOR U23230 ( .A(c4646), .B(n13938), .Z(c4647) );
ANDN U23231 ( .B(n13939), .A(n13940), .Z(n13938) );
XOR U23232 ( .A(c4646), .B(b[4646]), .Z(n13939) );
XNOR U23233 ( .A(b[4646]), .B(n13940), .Z(c[4646]) );
XNOR U23234 ( .A(a[4646]), .B(c4646), .Z(n13940) );
XOR U23235 ( .A(c4647), .B(n13941), .Z(c4648) );
ANDN U23236 ( .B(n13942), .A(n13943), .Z(n13941) );
XOR U23237 ( .A(c4647), .B(b[4647]), .Z(n13942) );
XNOR U23238 ( .A(b[4647]), .B(n13943), .Z(c[4647]) );
XNOR U23239 ( .A(a[4647]), .B(c4647), .Z(n13943) );
XOR U23240 ( .A(c4648), .B(n13944), .Z(c4649) );
ANDN U23241 ( .B(n13945), .A(n13946), .Z(n13944) );
XOR U23242 ( .A(c4648), .B(b[4648]), .Z(n13945) );
XNOR U23243 ( .A(b[4648]), .B(n13946), .Z(c[4648]) );
XNOR U23244 ( .A(a[4648]), .B(c4648), .Z(n13946) );
XOR U23245 ( .A(c4649), .B(n13947), .Z(c4650) );
ANDN U23246 ( .B(n13948), .A(n13949), .Z(n13947) );
XOR U23247 ( .A(c4649), .B(b[4649]), .Z(n13948) );
XNOR U23248 ( .A(b[4649]), .B(n13949), .Z(c[4649]) );
XNOR U23249 ( .A(a[4649]), .B(c4649), .Z(n13949) );
XOR U23250 ( .A(c4650), .B(n13950), .Z(c4651) );
ANDN U23251 ( .B(n13951), .A(n13952), .Z(n13950) );
XOR U23252 ( .A(c4650), .B(b[4650]), .Z(n13951) );
XNOR U23253 ( .A(b[4650]), .B(n13952), .Z(c[4650]) );
XNOR U23254 ( .A(a[4650]), .B(c4650), .Z(n13952) );
XOR U23255 ( .A(c4651), .B(n13953), .Z(c4652) );
ANDN U23256 ( .B(n13954), .A(n13955), .Z(n13953) );
XOR U23257 ( .A(c4651), .B(b[4651]), .Z(n13954) );
XNOR U23258 ( .A(b[4651]), .B(n13955), .Z(c[4651]) );
XNOR U23259 ( .A(a[4651]), .B(c4651), .Z(n13955) );
XOR U23260 ( .A(c4652), .B(n13956), .Z(c4653) );
ANDN U23261 ( .B(n13957), .A(n13958), .Z(n13956) );
XOR U23262 ( .A(c4652), .B(b[4652]), .Z(n13957) );
XNOR U23263 ( .A(b[4652]), .B(n13958), .Z(c[4652]) );
XNOR U23264 ( .A(a[4652]), .B(c4652), .Z(n13958) );
XOR U23265 ( .A(c4653), .B(n13959), .Z(c4654) );
ANDN U23266 ( .B(n13960), .A(n13961), .Z(n13959) );
XOR U23267 ( .A(c4653), .B(b[4653]), .Z(n13960) );
XNOR U23268 ( .A(b[4653]), .B(n13961), .Z(c[4653]) );
XNOR U23269 ( .A(a[4653]), .B(c4653), .Z(n13961) );
XOR U23270 ( .A(c4654), .B(n13962), .Z(c4655) );
ANDN U23271 ( .B(n13963), .A(n13964), .Z(n13962) );
XOR U23272 ( .A(c4654), .B(b[4654]), .Z(n13963) );
XNOR U23273 ( .A(b[4654]), .B(n13964), .Z(c[4654]) );
XNOR U23274 ( .A(a[4654]), .B(c4654), .Z(n13964) );
XOR U23275 ( .A(c4655), .B(n13965), .Z(c4656) );
ANDN U23276 ( .B(n13966), .A(n13967), .Z(n13965) );
XOR U23277 ( .A(c4655), .B(b[4655]), .Z(n13966) );
XNOR U23278 ( .A(b[4655]), .B(n13967), .Z(c[4655]) );
XNOR U23279 ( .A(a[4655]), .B(c4655), .Z(n13967) );
XOR U23280 ( .A(c4656), .B(n13968), .Z(c4657) );
ANDN U23281 ( .B(n13969), .A(n13970), .Z(n13968) );
XOR U23282 ( .A(c4656), .B(b[4656]), .Z(n13969) );
XNOR U23283 ( .A(b[4656]), .B(n13970), .Z(c[4656]) );
XNOR U23284 ( .A(a[4656]), .B(c4656), .Z(n13970) );
XOR U23285 ( .A(c4657), .B(n13971), .Z(c4658) );
ANDN U23286 ( .B(n13972), .A(n13973), .Z(n13971) );
XOR U23287 ( .A(c4657), .B(b[4657]), .Z(n13972) );
XNOR U23288 ( .A(b[4657]), .B(n13973), .Z(c[4657]) );
XNOR U23289 ( .A(a[4657]), .B(c4657), .Z(n13973) );
XOR U23290 ( .A(c4658), .B(n13974), .Z(c4659) );
ANDN U23291 ( .B(n13975), .A(n13976), .Z(n13974) );
XOR U23292 ( .A(c4658), .B(b[4658]), .Z(n13975) );
XNOR U23293 ( .A(b[4658]), .B(n13976), .Z(c[4658]) );
XNOR U23294 ( .A(a[4658]), .B(c4658), .Z(n13976) );
XOR U23295 ( .A(c4659), .B(n13977), .Z(c4660) );
ANDN U23296 ( .B(n13978), .A(n13979), .Z(n13977) );
XOR U23297 ( .A(c4659), .B(b[4659]), .Z(n13978) );
XNOR U23298 ( .A(b[4659]), .B(n13979), .Z(c[4659]) );
XNOR U23299 ( .A(a[4659]), .B(c4659), .Z(n13979) );
XOR U23300 ( .A(c4660), .B(n13980), .Z(c4661) );
ANDN U23301 ( .B(n13981), .A(n13982), .Z(n13980) );
XOR U23302 ( .A(c4660), .B(b[4660]), .Z(n13981) );
XNOR U23303 ( .A(b[4660]), .B(n13982), .Z(c[4660]) );
XNOR U23304 ( .A(a[4660]), .B(c4660), .Z(n13982) );
XOR U23305 ( .A(c4661), .B(n13983), .Z(c4662) );
ANDN U23306 ( .B(n13984), .A(n13985), .Z(n13983) );
XOR U23307 ( .A(c4661), .B(b[4661]), .Z(n13984) );
XNOR U23308 ( .A(b[4661]), .B(n13985), .Z(c[4661]) );
XNOR U23309 ( .A(a[4661]), .B(c4661), .Z(n13985) );
XOR U23310 ( .A(c4662), .B(n13986), .Z(c4663) );
ANDN U23311 ( .B(n13987), .A(n13988), .Z(n13986) );
XOR U23312 ( .A(c4662), .B(b[4662]), .Z(n13987) );
XNOR U23313 ( .A(b[4662]), .B(n13988), .Z(c[4662]) );
XNOR U23314 ( .A(a[4662]), .B(c4662), .Z(n13988) );
XOR U23315 ( .A(c4663), .B(n13989), .Z(c4664) );
ANDN U23316 ( .B(n13990), .A(n13991), .Z(n13989) );
XOR U23317 ( .A(c4663), .B(b[4663]), .Z(n13990) );
XNOR U23318 ( .A(b[4663]), .B(n13991), .Z(c[4663]) );
XNOR U23319 ( .A(a[4663]), .B(c4663), .Z(n13991) );
XOR U23320 ( .A(c4664), .B(n13992), .Z(c4665) );
ANDN U23321 ( .B(n13993), .A(n13994), .Z(n13992) );
XOR U23322 ( .A(c4664), .B(b[4664]), .Z(n13993) );
XNOR U23323 ( .A(b[4664]), .B(n13994), .Z(c[4664]) );
XNOR U23324 ( .A(a[4664]), .B(c4664), .Z(n13994) );
XOR U23325 ( .A(c4665), .B(n13995), .Z(c4666) );
ANDN U23326 ( .B(n13996), .A(n13997), .Z(n13995) );
XOR U23327 ( .A(c4665), .B(b[4665]), .Z(n13996) );
XNOR U23328 ( .A(b[4665]), .B(n13997), .Z(c[4665]) );
XNOR U23329 ( .A(a[4665]), .B(c4665), .Z(n13997) );
XOR U23330 ( .A(c4666), .B(n13998), .Z(c4667) );
ANDN U23331 ( .B(n13999), .A(n14000), .Z(n13998) );
XOR U23332 ( .A(c4666), .B(b[4666]), .Z(n13999) );
XNOR U23333 ( .A(b[4666]), .B(n14000), .Z(c[4666]) );
XNOR U23334 ( .A(a[4666]), .B(c4666), .Z(n14000) );
XOR U23335 ( .A(c4667), .B(n14001), .Z(c4668) );
ANDN U23336 ( .B(n14002), .A(n14003), .Z(n14001) );
XOR U23337 ( .A(c4667), .B(b[4667]), .Z(n14002) );
XNOR U23338 ( .A(b[4667]), .B(n14003), .Z(c[4667]) );
XNOR U23339 ( .A(a[4667]), .B(c4667), .Z(n14003) );
XOR U23340 ( .A(c4668), .B(n14004), .Z(c4669) );
ANDN U23341 ( .B(n14005), .A(n14006), .Z(n14004) );
XOR U23342 ( .A(c4668), .B(b[4668]), .Z(n14005) );
XNOR U23343 ( .A(b[4668]), .B(n14006), .Z(c[4668]) );
XNOR U23344 ( .A(a[4668]), .B(c4668), .Z(n14006) );
XOR U23345 ( .A(c4669), .B(n14007), .Z(c4670) );
ANDN U23346 ( .B(n14008), .A(n14009), .Z(n14007) );
XOR U23347 ( .A(c4669), .B(b[4669]), .Z(n14008) );
XNOR U23348 ( .A(b[4669]), .B(n14009), .Z(c[4669]) );
XNOR U23349 ( .A(a[4669]), .B(c4669), .Z(n14009) );
XOR U23350 ( .A(c4670), .B(n14010), .Z(c4671) );
ANDN U23351 ( .B(n14011), .A(n14012), .Z(n14010) );
XOR U23352 ( .A(c4670), .B(b[4670]), .Z(n14011) );
XNOR U23353 ( .A(b[4670]), .B(n14012), .Z(c[4670]) );
XNOR U23354 ( .A(a[4670]), .B(c4670), .Z(n14012) );
XOR U23355 ( .A(c4671), .B(n14013), .Z(c4672) );
ANDN U23356 ( .B(n14014), .A(n14015), .Z(n14013) );
XOR U23357 ( .A(c4671), .B(b[4671]), .Z(n14014) );
XNOR U23358 ( .A(b[4671]), .B(n14015), .Z(c[4671]) );
XNOR U23359 ( .A(a[4671]), .B(c4671), .Z(n14015) );
XOR U23360 ( .A(c4672), .B(n14016), .Z(c4673) );
ANDN U23361 ( .B(n14017), .A(n14018), .Z(n14016) );
XOR U23362 ( .A(c4672), .B(b[4672]), .Z(n14017) );
XNOR U23363 ( .A(b[4672]), .B(n14018), .Z(c[4672]) );
XNOR U23364 ( .A(a[4672]), .B(c4672), .Z(n14018) );
XOR U23365 ( .A(c4673), .B(n14019), .Z(c4674) );
ANDN U23366 ( .B(n14020), .A(n14021), .Z(n14019) );
XOR U23367 ( .A(c4673), .B(b[4673]), .Z(n14020) );
XNOR U23368 ( .A(b[4673]), .B(n14021), .Z(c[4673]) );
XNOR U23369 ( .A(a[4673]), .B(c4673), .Z(n14021) );
XOR U23370 ( .A(c4674), .B(n14022), .Z(c4675) );
ANDN U23371 ( .B(n14023), .A(n14024), .Z(n14022) );
XOR U23372 ( .A(c4674), .B(b[4674]), .Z(n14023) );
XNOR U23373 ( .A(b[4674]), .B(n14024), .Z(c[4674]) );
XNOR U23374 ( .A(a[4674]), .B(c4674), .Z(n14024) );
XOR U23375 ( .A(c4675), .B(n14025), .Z(c4676) );
ANDN U23376 ( .B(n14026), .A(n14027), .Z(n14025) );
XOR U23377 ( .A(c4675), .B(b[4675]), .Z(n14026) );
XNOR U23378 ( .A(b[4675]), .B(n14027), .Z(c[4675]) );
XNOR U23379 ( .A(a[4675]), .B(c4675), .Z(n14027) );
XOR U23380 ( .A(c4676), .B(n14028), .Z(c4677) );
ANDN U23381 ( .B(n14029), .A(n14030), .Z(n14028) );
XOR U23382 ( .A(c4676), .B(b[4676]), .Z(n14029) );
XNOR U23383 ( .A(b[4676]), .B(n14030), .Z(c[4676]) );
XNOR U23384 ( .A(a[4676]), .B(c4676), .Z(n14030) );
XOR U23385 ( .A(c4677), .B(n14031), .Z(c4678) );
ANDN U23386 ( .B(n14032), .A(n14033), .Z(n14031) );
XOR U23387 ( .A(c4677), .B(b[4677]), .Z(n14032) );
XNOR U23388 ( .A(b[4677]), .B(n14033), .Z(c[4677]) );
XNOR U23389 ( .A(a[4677]), .B(c4677), .Z(n14033) );
XOR U23390 ( .A(c4678), .B(n14034), .Z(c4679) );
ANDN U23391 ( .B(n14035), .A(n14036), .Z(n14034) );
XOR U23392 ( .A(c4678), .B(b[4678]), .Z(n14035) );
XNOR U23393 ( .A(b[4678]), .B(n14036), .Z(c[4678]) );
XNOR U23394 ( .A(a[4678]), .B(c4678), .Z(n14036) );
XOR U23395 ( .A(c4679), .B(n14037), .Z(c4680) );
ANDN U23396 ( .B(n14038), .A(n14039), .Z(n14037) );
XOR U23397 ( .A(c4679), .B(b[4679]), .Z(n14038) );
XNOR U23398 ( .A(b[4679]), .B(n14039), .Z(c[4679]) );
XNOR U23399 ( .A(a[4679]), .B(c4679), .Z(n14039) );
XOR U23400 ( .A(c4680), .B(n14040), .Z(c4681) );
ANDN U23401 ( .B(n14041), .A(n14042), .Z(n14040) );
XOR U23402 ( .A(c4680), .B(b[4680]), .Z(n14041) );
XNOR U23403 ( .A(b[4680]), .B(n14042), .Z(c[4680]) );
XNOR U23404 ( .A(a[4680]), .B(c4680), .Z(n14042) );
XOR U23405 ( .A(c4681), .B(n14043), .Z(c4682) );
ANDN U23406 ( .B(n14044), .A(n14045), .Z(n14043) );
XOR U23407 ( .A(c4681), .B(b[4681]), .Z(n14044) );
XNOR U23408 ( .A(b[4681]), .B(n14045), .Z(c[4681]) );
XNOR U23409 ( .A(a[4681]), .B(c4681), .Z(n14045) );
XOR U23410 ( .A(c4682), .B(n14046), .Z(c4683) );
ANDN U23411 ( .B(n14047), .A(n14048), .Z(n14046) );
XOR U23412 ( .A(c4682), .B(b[4682]), .Z(n14047) );
XNOR U23413 ( .A(b[4682]), .B(n14048), .Z(c[4682]) );
XNOR U23414 ( .A(a[4682]), .B(c4682), .Z(n14048) );
XOR U23415 ( .A(c4683), .B(n14049), .Z(c4684) );
ANDN U23416 ( .B(n14050), .A(n14051), .Z(n14049) );
XOR U23417 ( .A(c4683), .B(b[4683]), .Z(n14050) );
XNOR U23418 ( .A(b[4683]), .B(n14051), .Z(c[4683]) );
XNOR U23419 ( .A(a[4683]), .B(c4683), .Z(n14051) );
XOR U23420 ( .A(c4684), .B(n14052), .Z(c4685) );
ANDN U23421 ( .B(n14053), .A(n14054), .Z(n14052) );
XOR U23422 ( .A(c4684), .B(b[4684]), .Z(n14053) );
XNOR U23423 ( .A(b[4684]), .B(n14054), .Z(c[4684]) );
XNOR U23424 ( .A(a[4684]), .B(c4684), .Z(n14054) );
XOR U23425 ( .A(c4685), .B(n14055), .Z(c4686) );
ANDN U23426 ( .B(n14056), .A(n14057), .Z(n14055) );
XOR U23427 ( .A(c4685), .B(b[4685]), .Z(n14056) );
XNOR U23428 ( .A(b[4685]), .B(n14057), .Z(c[4685]) );
XNOR U23429 ( .A(a[4685]), .B(c4685), .Z(n14057) );
XOR U23430 ( .A(c4686), .B(n14058), .Z(c4687) );
ANDN U23431 ( .B(n14059), .A(n14060), .Z(n14058) );
XOR U23432 ( .A(c4686), .B(b[4686]), .Z(n14059) );
XNOR U23433 ( .A(b[4686]), .B(n14060), .Z(c[4686]) );
XNOR U23434 ( .A(a[4686]), .B(c4686), .Z(n14060) );
XOR U23435 ( .A(c4687), .B(n14061), .Z(c4688) );
ANDN U23436 ( .B(n14062), .A(n14063), .Z(n14061) );
XOR U23437 ( .A(c4687), .B(b[4687]), .Z(n14062) );
XNOR U23438 ( .A(b[4687]), .B(n14063), .Z(c[4687]) );
XNOR U23439 ( .A(a[4687]), .B(c4687), .Z(n14063) );
XOR U23440 ( .A(c4688), .B(n14064), .Z(c4689) );
ANDN U23441 ( .B(n14065), .A(n14066), .Z(n14064) );
XOR U23442 ( .A(c4688), .B(b[4688]), .Z(n14065) );
XNOR U23443 ( .A(b[4688]), .B(n14066), .Z(c[4688]) );
XNOR U23444 ( .A(a[4688]), .B(c4688), .Z(n14066) );
XOR U23445 ( .A(c4689), .B(n14067), .Z(c4690) );
ANDN U23446 ( .B(n14068), .A(n14069), .Z(n14067) );
XOR U23447 ( .A(c4689), .B(b[4689]), .Z(n14068) );
XNOR U23448 ( .A(b[4689]), .B(n14069), .Z(c[4689]) );
XNOR U23449 ( .A(a[4689]), .B(c4689), .Z(n14069) );
XOR U23450 ( .A(c4690), .B(n14070), .Z(c4691) );
ANDN U23451 ( .B(n14071), .A(n14072), .Z(n14070) );
XOR U23452 ( .A(c4690), .B(b[4690]), .Z(n14071) );
XNOR U23453 ( .A(b[4690]), .B(n14072), .Z(c[4690]) );
XNOR U23454 ( .A(a[4690]), .B(c4690), .Z(n14072) );
XOR U23455 ( .A(c4691), .B(n14073), .Z(c4692) );
ANDN U23456 ( .B(n14074), .A(n14075), .Z(n14073) );
XOR U23457 ( .A(c4691), .B(b[4691]), .Z(n14074) );
XNOR U23458 ( .A(b[4691]), .B(n14075), .Z(c[4691]) );
XNOR U23459 ( .A(a[4691]), .B(c4691), .Z(n14075) );
XOR U23460 ( .A(c4692), .B(n14076), .Z(c4693) );
ANDN U23461 ( .B(n14077), .A(n14078), .Z(n14076) );
XOR U23462 ( .A(c4692), .B(b[4692]), .Z(n14077) );
XNOR U23463 ( .A(b[4692]), .B(n14078), .Z(c[4692]) );
XNOR U23464 ( .A(a[4692]), .B(c4692), .Z(n14078) );
XOR U23465 ( .A(c4693), .B(n14079), .Z(c4694) );
ANDN U23466 ( .B(n14080), .A(n14081), .Z(n14079) );
XOR U23467 ( .A(c4693), .B(b[4693]), .Z(n14080) );
XNOR U23468 ( .A(b[4693]), .B(n14081), .Z(c[4693]) );
XNOR U23469 ( .A(a[4693]), .B(c4693), .Z(n14081) );
XOR U23470 ( .A(c4694), .B(n14082), .Z(c4695) );
ANDN U23471 ( .B(n14083), .A(n14084), .Z(n14082) );
XOR U23472 ( .A(c4694), .B(b[4694]), .Z(n14083) );
XNOR U23473 ( .A(b[4694]), .B(n14084), .Z(c[4694]) );
XNOR U23474 ( .A(a[4694]), .B(c4694), .Z(n14084) );
XOR U23475 ( .A(c4695), .B(n14085), .Z(c4696) );
ANDN U23476 ( .B(n14086), .A(n14087), .Z(n14085) );
XOR U23477 ( .A(c4695), .B(b[4695]), .Z(n14086) );
XNOR U23478 ( .A(b[4695]), .B(n14087), .Z(c[4695]) );
XNOR U23479 ( .A(a[4695]), .B(c4695), .Z(n14087) );
XOR U23480 ( .A(c4696), .B(n14088), .Z(c4697) );
ANDN U23481 ( .B(n14089), .A(n14090), .Z(n14088) );
XOR U23482 ( .A(c4696), .B(b[4696]), .Z(n14089) );
XNOR U23483 ( .A(b[4696]), .B(n14090), .Z(c[4696]) );
XNOR U23484 ( .A(a[4696]), .B(c4696), .Z(n14090) );
XOR U23485 ( .A(c4697), .B(n14091), .Z(c4698) );
ANDN U23486 ( .B(n14092), .A(n14093), .Z(n14091) );
XOR U23487 ( .A(c4697), .B(b[4697]), .Z(n14092) );
XNOR U23488 ( .A(b[4697]), .B(n14093), .Z(c[4697]) );
XNOR U23489 ( .A(a[4697]), .B(c4697), .Z(n14093) );
XOR U23490 ( .A(c4698), .B(n14094), .Z(c4699) );
ANDN U23491 ( .B(n14095), .A(n14096), .Z(n14094) );
XOR U23492 ( .A(c4698), .B(b[4698]), .Z(n14095) );
XNOR U23493 ( .A(b[4698]), .B(n14096), .Z(c[4698]) );
XNOR U23494 ( .A(a[4698]), .B(c4698), .Z(n14096) );
XOR U23495 ( .A(c4699), .B(n14097), .Z(c4700) );
ANDN U23496 ( .B(n14098), .A(n14099), .Z(n14097) );
XOR U23497 ( .A(c4699), .B(b[4699]), .Z(n14098) );
XNOR U23498 ( .A(b[4699]), .B(n14099), .Z(c[4699]) );
XNOR U23499 ( .A(a[4699]), .B(c4699), .Z(n14099) );
XOR U23500 ( .A(c4700), .B(n14100), .Z(c4701) );
ANDN U23501 ( .B(n14101), .A(n14102), .Z(n14100) );
XOR U23502 ( .A(c4700), .B(b[4700]), .Z(n14101) );
XNOR U23503 ( .A(b[4700]), .B(n14102), .Z(c[4700]) );
XNOR U23504 ( .A(a[4700]), .B(c4700), .Z(n14102) );
XOR U23505 ( .A(c4701), .B(n14103), .Z(c4702) );
ANDN U23506 ( .B(n14104), .A(n14105), .Z(n14103) );
XOR U23507 ( .A(c4701), .B(b[4701]), .Z(n14104) );
XNOR U23508 ( .A(b[4701]), .B(n14105), .Z(c[4701]) );
XNOR U23509 ( .A(a[4701]), .B(c4701), .Z(n14105) );
XOR U23510 ( .A(c4702), .B(n14106), .Z(c4703) );
ANDN U23511 ( .B(n14107), .A(n14108), .Z(n14106) );
XOR U23512 ( .A(c4702), .B(b[4702]), .Z(n14107) );
XNOR U23513 ( .A(b[4702]), .B(n14108), .Z(c[4702]) );
XNOR U23514 ( .A(a[4702]), .B(c4702), .Z(n14108) );
XOR U23515 ( .A(c4703), .B(n14109), .Z(c4704) );
ANDN U23516 ( .B(n14110), .A(n14111), .Z(n14109) );
XOR U23517 ( .A(c4703), .B(b[4703]), .Z(n14110) );
XNOR U23518 ( .A(b[4703]), .B(n14111), .Z(c[4703]) );
XNOR U23519 ( .A(a[4703]), .B(c4703), .Z(n14111) );
XOR U23520 ( .A(c4704), .B(n14112), .Z(c4705) );
ANDN U23521 ( .B(n14113), .A(n14114), .Z(n14112) );
XOR U23522 ( .A(c4704), .B(b[4704]), .Z(n14113) );
XNOR U23523 ( .A(b[4704]), .B(n14114), .Z(c[4704]) );
XNOR U23524 ( .A(a[4704]), .B(c4704), .Z(n14114) );
XOR U23525 ( .A(c4705), .B(n14115), .Z(c4706) );
ANDN U23526 ( .B(n14116), .A(n14117), .Z(n14115) );
XOR U23527 ( .A(c4705), .B(b[4705]), .Z(n14116) );
XNOR U23528 ( .A(b[4705]), .B(n14117), .Z(c[4705]) );
XNOR U23529 ( .A(a[4705]), .B(c4705), .Z(n14117) );
XOR U23530 ( .A(c4706), .B(n14118), .Z(c4707) );
ANDN U23531 ( .B(n14119), .A(n14120), .Z(n14118) );
XOR U23532 ( .A(c4706), .B(b[4706]), .Z(n14119) );
XNOR U23533 ( .A(b[4706]), .B(n14120), .Z(c[4706]) );
XNOR U23534 ( .A(a[4706]), .B(c4706), .Z(n14120) );
XOR U23535 ( .A(c4707), .B(n14121), .Z(c4708) );
ANDN U23536 ( .B(n14122), .A(n14123), .Z(n14121) );
XOR U23537 ( .A(c4707), .B(b[4707]), .Z(n14122) );
XNOR U23538 ( .A(b[4707]), .B(n14123), .Z(c[4707]) );
XNOR U23539 ( .A(a[4707]), .B(c4707), .Z(n14123) );
XOR U23540 ( .A(c4708), .B(n14124), .Z(c4709) );
ANDN U23541 ( .B(n14125), .A(n14126), .Z(n14124) );
XOR U23542 ( .A(c4708), .B(b[4708]), .Z(n14125) );
XNOR U23543 ( .A(b[4708]), .B(n14126), .Z(c[4708]) );
XNOR U23544 ( .A(a[4708]), .B(c4708), .Z(n14126) );
XOR U23545 ( .A(c4709), .B(n14127), .Z(c4710) );
ANDN U23546 ( .B(n14128), .A(n14129), .Z(n14127) );
XOR U23547 ( .A(c4709), .B(b[4709]), .Z(n14128) );
XNOR U23548 ( .A(b[4709]), .B(n14129), .Z(c[4709]) );
XNOR U23549 ( .A(a[4709]), .B(c4709), .Z(n14129) );
XOR U23550 ( .A(c4710), .B(n14130), .Z(c4711) );
ANDN U23551 ( .B(n14131), .A(n14132), .Z(n14130) );
XOR U23552 ( .A(c4710), .B(b[4710]), .Z(n14131) );
XNOR U23553 ( .A(b[4710]), .B(n14132), .Z(c[4710]) );
XNOR U23554 ( .A(a[4710]), .B(c4710), .Z(n14132) );
XOR U23555 ( .A(c4711), .B(n14133), .Z(c4712) );
ANDN U23556 ( .B(n14134), .A(n14135), .Z(n14133) );
XOR U23557 ( .A(c4711), .B(b[4711]), .Z(n14134) );
XNOR U23558 ( .A(b[4711]), .B(n14135), .Z(c[4711]) );
XNOR U23559 ( .A(a[4711]), .B(c4711), .Z(n14135) );
XOR U23560 ( .A(c4712), .B(n14136), .Z(c4713) );
ANDN U23561 ( .B(n14137), .A(n14138), .Z(n14136) );
XOR U23562 ( .A(c4712), .B(b[4712]), .Z(n14137) );
XNOR U23563 ( .A(b[4712]), .B(n14138), .Z(c[4712]) );
XNOR U23564 ( .A(a[4712]), .B(c4712), .Z(n14138) );
XOR U23565 ( .A(c4713), .B(n14139), .Z(c4714) );
ANDN U23566 ( .B(n14140), .A(n14141), .Z(n14139) );
XOR U23567 ( .A(c4713), .B(b[4713]), .Z(n14140) );
XNOR U23568 ( .A(b[4713]), .B(n14141), .Z(c[4713]) );
XNOR U23569 ( .A(a[4713]), .B(c4713), .Z(n14141) );
XOR U23570 ( .A(c4714), .B(n14142), .Z(c4715) );
ANDN U23571 ( .B(n14143), .A(n14144), .Z(n14142) );
XOR U23572 ( .A(c4714), .B(b[4714]), .Z(n14143) );
XNOR U23573 ( .A(b[4714]), .B(n14144), .Z(c[4714]) );
XNOR U23574 ( .A(a[4714]), .B(c4714), .Z(n14144) );
XOR U23575 ( .A(c4715), .B(n14145), .Z(c4716) );
ANDN U23576 ( .B(n14146), .A(n14147), .Z(n14145) );
XOR U23577 ( .A(c4715), .B(b[4715]), .Z(n14146) );
XNOR U23578 ( .A(b[4715]), .B(n14147), .Z(c[4715]) );
XNOR U23579 ( .A(a[4715]), .B(c4715), .Z(n14147) );
XOR U23580 ( .A(c4716), .B(n14148), .Z(c4717) );
ANDN U23581 ( .B(n14149), .A(n14150), .Z(n14148) );
XOR U23582 ( .A(c4716), .B(b[4716]), .Z(n14149) );
XNOR U23583 ( .A(b[4716]), .B(n14150), .Z(c[4716]) );
XNOR U23584 ( .A(a[4716]), .B(c4716), .Z(n14150) );
XOR U23585 ( .A(c4717), .B(n14151), .Z(c4718) );
ANDN U23586 ( .B(n14152), .A(n14153), .Z(n14151) );
XOR U23587 ( .A(c4717), .B(b[4717]), .Z(n14152) );
XNOR U23588 ( .A(b[4717]), .B(n14153), .Z(c[4717]) );
XNOR U23589 ( .A(a[4717]), .B(c4717), .Z(n14153) );
XOR U23590 ( .A(c4718), .B(n14154), .Z(c4719) );
ANDN U23591 ( .B(n14155), .A(n14156), .Z(n14154) );
XOR U23592 ( .A(c4718), .B(b[4718]), .Z(n14155) );
XNOR U23593 ( .A(b[4718]), .B(n14156), .Z(c[4718]) );
XNOR U23594 ( .A(a[4718]), .B(c4718), .Z(n14156) );
XOR U23595 ( .A(c4719), .B(n14157), .Z(c4720) );
ANDN U23596 ( .B(n14158), .A(n14159), .Z(n14157) );
XOR U23597 ( .A(c4719), .B(b[4719]), .Z(n14158) );
XNOR U23598 ( .A(b[4719]), .B(n14159), .Z(c[4719]) );
XNOR U23599 ( .A(a[4719]), .B(c4719), .Z(n14159) );
XOR U23600 ( .A(c4720), .B(n14160), .Z(c4721) );
ANDN U23601 ( .B(n14161), .A(n14162), .Z(n14160) );
XOR U23602 ( .A(c4720), .B(b[4720]), .Z(n14161) );
XNOR U23603 ( .A(b[4720]), .B(n14162), .Z(c[4720]) );
XNOR U23604 ( .A(a[4720]), .B(c4720), .Z(n14162) );
XOR U23605 ( .A(c4721), .B(n14163), .Z(c4722) );
ANDN U23606 ( .B(n14164), .A(n14165), .Z(n14163) );
XOR U23607 ( .A(c4721), .B(b[4721]), .Z(n14164) );
XNOR U23608 ( .A(b[4721]), .B(n14165), .Z(c[4721]) );
XNOR U23609 ( .A(a[4721]), .B(c4721), .Z(n14165) );
XOR U23610 ( .A(c4722), .B(n14166), .Z(c4723) );
ANDN U23611 ( .B(n14167), .A(n14168), .Z(n14166) );
XOR U23612 ( .A(c4722), .B(b[4722]), .Z(n14167) );
XNOR U23613 ( .A(b[4722]), .B(n14168), .Z(c[4722]) );
XNOR U23614 ( .A(a[4722]), .B(c4722), .Z(n14168) );
XOR U23615 ( .A(c4723), .B(n14169), .Z(c4724) );
ANDN U23616 ( .B(n14170), .A(n14171), .Z(n14169) );
XOR U23617 ( .A(c4723), .B(b[4723]), .Z(n14170) );
XNOR U23618 ( .A(b[4723]), .B(n14171), .Z(c[4723]) );
XNOR U23619 ( .A(a[4723]), .B(c4723), .Z(n14171) );
XOR U23620 ( .A(c4724), .B(n14172), .Z(c4725) );
ANDN U23621 ( .B(n14173), .A(n14174), .Z(n14172) );
XOR U23622 ( .A(c4724), .B(b[4724]), .Z(n14173) );
XNOR U23623 ( .A(b[4724]), .B(n14174), .Z(c[4724]) );
XNOR U23624 ( .A(a[4724]), .B(c4724), .Z(n14174) );
XOR U23625 ( .A(c4725), .B(n14175), .Z(c4726) );
ANDN U23626 ( .B(n14176), .A(n14177), .Z(n14175) );
XOR U23627 ( .A(c4725), .B(b[4725]), .Z(n14176) );
XNOR U23628 ( .A(b[4725]), .B(n14177), .Z(c[4725]) );
XNOR U23629 ( .A(a[4725]), .B(c4725), .Z(n14177) );
XOR U23630 ( .A(c4726), .B(n14178), .Z(c4727) );
ANDN U23631 ( .B(n14179), .A(n14180), .Z(n14178) );
XOR U23632 ( .A(c4726), .B(b[4726]), .Z(n14179) );
XNOR U23633 ( .A(b[4726]), .B(n14180), .Z(c[4726]) );
XNOR U23634 ( .A(a[4726]), .B(c4726), .Z(n14180) );
XOR U23635 ( .A(c4727), .B(n14181), .Z(c4728) );
ANDN U23636 ( .B(n14182), .A(n14183), .Z(n14181) );
XOR U23637 ( .A(c4727), .B(b[4727]), .Z(n14182) );
XNOR U23638 ( .A(b[4727]), .B(n14183), .Z(c[4727]) );
XNOR U23639 ( .A(a[4727]), .B(c4727), .Z(n14183) );
XOR U23640 ( .A(c4728), .B(n14184), .Z(c4729) );
ANDN U23641 ( .B(n14185), .A(n14186), .Z(n14184) );
XOR U23642 ( .A(c4728), .B(b[4728]), .Z(n14185) );
XNOR U23643 ( .A(b[4728]), .B(n14186), .Z(c[4728]) );
XNOR U23644 ( .A(a[4728]), .B(c4728), .Z(n14186) );
XOR U23645 ( .A(c4729), .B(n14187), .Z(c4730) );
ANDN U23646 ( .B(n14188), .A(n14189), .Z(n14187) );
XOR U23647 ( .A(c4729), .B(b[4729]), .Z(n14188) );
XNOR U23648 ( .A(b[4729]), .B(n14189), .Z(c[4729]) );
XNOR U23649 ( .A(a[4729]), .B(c4729), .Z(n14189) );
XOR U23650 ( .A(c4730), .B(n14190), .Z(c4731) );
ANDN U23651 ( .B(n14191), .A(n14192), .Z(n14190) );
XOR U23652 ( .A(c4730), .B(b[4730]), .Z(n14191) );
XNOR U23653 ( .A(b[4730]), .B(n14192), .Z(c[4730]) );
XNOR U23654 ( .A(a[4730]), .B(c4730), .Z(n14192) );
XOR U23655 ( .A(c4731), .B(n14193), .Z(c4732) );
ANDN U23656 ( .B(n14194), .A(n14195), .Z(n14193) );
XOR U23657 ( .A(c4731), .B(b[4731]), .Z(n14194) );
XNOR U23658 ( .A(b[4731]), .B(n14195), .Z(c[4731]) );
XNOR U23659 ( .A(a[4731]), .B(c4731), .Z(n14195) );
XOR U23660 ( .A(c4732), .B(n14196), .Z(c4733) );
ANDN U23661 ( .B(n14197), .A(n14198), .Z(n14196) );
XOR U23662 ( .A(c4732), .B(b[4732]), .Z(n14197) );
XNOR U23663 ( .A(b[4732]), .B(n14198), .Z(c[4732]) );
XNOR U23664 ( .A(a[4732]), .B(c4732), .Z(n14198) );
XOR U23665 ( .A(c4733), .B(n14199), .Z(c4734) );
ANDN U23666 ( .B(n14200), .A(n14201), .Z(n14199) );
XOR U23667 ( .A(c4733), .B(b[4733]), .Z(n14200) );
XNOR U23668 ( .A(b[4733]), .B(n14201), .Z(c[4733]) );
XNOR U23669 ( .A(a[4733]), .B(c4733), .Z(n14201) );
XOR U23670 ( .A(c4734), .B(n14202), .Z(c4735) );
ANDN U23671 ( .B(n14203), .A(n14204), .Z(n14202) );
XOR U23672 ( .A(c4734), .B(b[4734]), .Z(n14203) );
XNOR U23673 ( .A(b[4734]), .B(n14204), .Z(c[4734]) );
XNOR U23674 ( .A(a[4734]), .B(c4734), .Z(n14204) );
XOR U23675 ( .A(c4735), .B(n14205), .Z(c4736) );
ANDN U23676 ( .B(n14206), .A(n14207), .Z(n14205) );
XOR U23677 ( .A(c4735), .B(b[4735]), .Z(n14206) );
XNOR U23678 ( .A(b[4735]), .B(n14207), .Z(c[4735]) );
XNOR U23679 ( .A(a[4735]), .B(c4735), .Z(n14207) );
XOR U23680 ( .A(c4736), .B(n14208), .Z(c4737) );
ANDN U23681 ( .B(n14209), .A(n14210), .Z(n14208) );
XOR U23682 ( .A(c4736), .B(b[4736]), .Z(n14209) );
XNOR U23683 ( .A(b[4736]), .B(n14210), .Z(c[4736]) );
XNOR U23684 ( .A(a[4736]), .B(c4736), .Z(n14210) );
XOR U23685 ( .A(c4737), .B(n14211), .Z(c4738) );
ANDN U23686 ( .B(n14212), .A(n14213), .Z(n14211) );
XOR U23687 ( .A(c4737), .B(b[4737]), .Z(n14212) );
XNOR U23688 ( .A(b[4737]), .B(n14213), .Z(c[4737]) );
XNOR U23689 ( .A(a[4737]), .B(c4737), .Z(n14213) );
XOR U23690 ( .A(c4738), .B(n14214), .Z(c4739) );
ANDN U23691 ( .B(n14215), .A(n14216), .Z(n14214) );
XOR U23692 ( .A(c4738), .B(b[4738]), .Z(n14215) );
XNOR U23693 ( .A(b[4738]), .B(n14216), .Z(c[4738]) );
XNOR U23694 ( .A(a[4738]), .B(c4738), .Z(n14216) );
XOR U23695 ( .A(c4739), .B(n14217), .Z(c4740) );
ANDN U23696 ( .B(n14218), .A(n14219), .Z(n14217) );
XOR U23697 ( .A(c4739), .B(b[4739]), .Z(n14218) );
XNOR U23698 ( .A(b[4739]), .B(n14219), .Z(c[4739]) );
XNOR U23699 ( .A(a[4739]), .B(c4739), .Z(n14219) );
XOR U23700 ( .A(c4740), .B(n14220), .Z(c4741) );
ANDN U23701 ( .B(n14221), .A(n14222), .Z(n14220) );
XOR U23702 ( .A(c4740), .B(b[4740]), .Z(n14221) );
XNOR U23703 ( .A(b[4740]), .B(n14222), .Z(c[4740]) );
XNOR U23704 ( .A(a[4740]), .B(c4740), .Z(n14222) );
XOR U23705 ( .A(c4741), .B(n14223), .Z(c4742) );
ANDN U23706 ( .B(n14224), .A(n14225), .Z(n14223) );
XOR U23707 ( .A(c4741), .B(b[4741]), .Z(n14224) );
XNOR U23708 ( .A(b[4741]), .B(n14225), .Z(c[4741]) );
XNOR U23709 ( .A(a[4741]), .B(c4741), .Z(n14225) );
XOR U23710 ( .A(c4742), .B(n14226), .Z(c4743) );
ANDN U23711 ( .B(n14227), .A(n14228), .Z(n14226) );
XOR U23712 ( .A(c4742), .B(b[4742]), .Z(n14227) );
XNOR U23713 ( .A(b[4742]), .B(n14228), .Z(c[4742]) );
XNOR U23714 ( .A(a[4742]), .B(c4742), .Z(n14228) );
XOR U23715 ( .A(c4743), .B(n14229), .Z(c4744) );
ANDN U23716 ( .B(n14230), .A(n14231), .Z(n14229) );
XOR U23717 ( .A(c4743), .B(b[4743]), .Z(n14230) );
XNOR U23718 ( .A(b[4743]), .B(n14231), .Z(c[4743]) );
XNOR U23719 ( .A(a[4743]), .B(c4743), .Z(n14231) );
XOR U23720 ( .A(c4744), .B(n14232), .Z(c4745) );
ANDN U23721 ( .B(n14233), .A(n14234), .Z(n14232) );
XOR U23722 ( .A(c4744), .B(b[4744]), .Z(n14233) );
XNOR U23723 ( .A(b[4744]), .B(n14234), .Z(c[4744]) );
XNOR U23724 ( .A(a[4744]), .B(c4744), .Z(n14234) );
XOR U23725 ( .A(c4745), .B(n14235), .Z(c4746) );
ANDN U23726 ( .B(n14236), .A(n14237), .Z(n14235) );
XOR U23727 ( .A(c4745), .B(b[4745]), .Z(n14236) );
XNOR U23728 ( .A(b[4745]), .B(n14237), .Z(c[4745]) );
XNOR U23729 ( .A(a[4745]), .B(c4745), .Z(n14237) );
XOR U23730 ( .A(c4746), .B(n14238), .Z(c4747) );
ANDN U23731 ( .B(n14239), .A(n14240), .Z(n14238) );
XOR U23732 ( .A(c4746), .B(b[4746]), .Z(n14239) );
XNOR U23733 ( .A(b[4746]), .B(n14240), .Z(c[4746]) );
XNOR U23734 ( .A(a[4746]), .B(c4746), .Z(n14240) );
XOR U23735 ( .A(c4747), .B(n14241), .Z(c4748) );
ANDN U23736 ( .B(n14242), .A(n14243), .Z(n14241) );
XOR U23737 ( .A(c4747), .B(b[4747]), .Z(n14242) );
XNOR U23738 ( .A(b[4747]), .B(n14243), .Z(c[4747]) );
XNOR U23739 ( .A(a[4747]), .B(c4747), .Z(n14243) );
XOR U23740 ( .A(c4748), .B(n14244), .Z(c4749) );
ANDN U23741 ( .B(n14245), .A(n14246), .Z(n14244) );
XOR U23742 ( .A(c4748), .B(b[4748]), .Z(n14245) );
XNOR U23743 ( .A(b[4748]), .B(n14246), .Z(c[4748]) );
XNOR U23744 ( .A(a[4748]), .B(c4748), .Z(n14246) );
XOR U23745 ( .A(c4749), .B(n14247), .Z(c4750) );
ANDN U23746 ( .B(n14248), .A(n14249), .Z(n14247) );
XOR U23747 ( .A(c4749), .B(b[4749]), .Z(n14248) );
XNOR U23748 ( .A(b[4749]), .B(n14249), .Z(c[4749]) );
XNOR U23749 ( .A(a[4749]), .B(c4749), .Z(n14249) );
XOR U23750 ( .A(c4750), .B(n14250), .Z(c4751) );
ANDN U23751 ( .B(n14251), .A(n14252), .Z(n14250) );
XOR U23752 ( .A(c4750), .B(b[4750]), .Z(n14251) );
XNOR U23753 ( .A(b[4750]), .B(n14252), .Z(c[4750]) );
XNOR U23754 ( .A(a[4750]), .B(c4750), .Z(n14252) );
XOR U23755 ( .A(c4751), .B(n14253), .Z(c4752) );
ANDN U23756 ( .B(n14254), .A(n14255), .Z(n14253) );
XOR U23757 ( .A(c4751), .B(b[4751]), .Z(n14254) );
XNOR U23758 ( .A(b[4751]), .B(n14255), .Z(c[4751]) );
XNOR U23759 ( .A(a[4751]), .B(c4751), .Z(n14255) );
XOR U23760 ( .A(c4752), .B(n14256), .Z(c4753) );
ANDN U23761 ( .B(n14257), .A(n14258), .Z(n14256) );
XOR U23762 ( .A(c4752), .B(b[4752]), .Z(n14257) );
XNOR U23763 ( .A(b[4752]), .B(n14258), .Z(c[4752]) );
XNOR U23764 ( .A(a[4752]), .B(c4752), .Z(n14258) );
XOR U23765 ( .A(c4753), .B(n14259), .Z(c4754) );
ANDN U23766 ( .B(n14260), .A(n14261), .Z(n14259) );
XOR U23767 ( .A(c4753), .B(b[4753]), .Z(n14260) );
XNOR U23768 ( .A(b[4753]), .B(n14261), .Z(c[4753]) );
XNOR U23769 ( .A(a[4753]), .B(c4753), .Z(n14261) );
XOR U23770 ( .A(c4754), .B(n14262), .Z(c4755) );
ANDN U23771 ( .B(n14263), .A(n14264), .Z(n14262) );
XOR U23772 ( .A(c4754), .B(b[4754]), .Z(n14263) );
XNOR U23773 ( .A(b[4754]), .B(n14264), .Z(c[4754]) );
XNOR U23774 ( .A(a[4754]), .B(c4754), .Z(n14264) );
XOR U23775 ( .A(c4755), .B(n14265), .Z(c4756) );
ANDN U23776 ( .B(n14266), .A(n14267), .Z(n14265) );
XOR U23777 ( .A(c4755), .B(b[4755]), .Z(n14266) );
XNOR U23778 ( .A(b[4755]), .B(n14267), .Z(c[4755]) );
XNOR U23779 ( .A(a[4755]), .B(c4755), .Z(n14267) );
XOR U23780 ( .A(c4756), .B(n14268), .Z(c4757) );
ANDN U23781 ( .B(n14269), .A(n14270), .Z(n14268) );
XOR U23782 ( .A(c4756), .B(b[4756]), .Z(n14269) );
XNOR U23783 ( .A(b[4756]), .B(n14270), .Z(c[4756]) );
XNOR U23784 ( .A(a[4756]), .B(c4756), .Z(n14270) );
XOR U23785 ( .A(c4757), .B(n14271), .Z(c4758) );
ANDN U23786 ( .B(n14272), .A(n14273), .Z(n14271) );
XOR U23787 ( .A(c4757), .B(b[4757]), .Z(n14272) );
XNOR U23788 ( .A(b[4757]), .B(n14273), .Z(c[4757]) );
XNOR U23789 ( .A(a[4757]), .B(c4757), .Z(n14273) );
XOR U23790 ( .A(c4758), .B(n14274), .Z(c4759) );
ANDN U23791 ( .B(n14275), .A(n14276), .Z(n14274) );
XOR U23792 ( .A(c4758), .B(b[4758]), .Z(n14275) );
XNOR U23793 ( .A(b[4758]), .B(n14276), .Z(c[4758]) );
XNOR U23794 ( .A(a[4758]), .B(c4758), .Z(n14276) );
XOR U23795 ( .A(c4759), .B(n14277), .Z(c4760) );
ANDN U23796 ( .B(n14278), .A(n14279), .Z(n14277) );
XOR U23797 ( .A(c4759), .B(b[4759]), .Z(n14278) );
XNOR U23798 ( .A(b[4759]), .B(n14279), .Z(c[4759]) );
XNOR U23799 ( .A(a[4759]), .B(c4759), .Z(n14279) );
XOR U23800 ( .A(c4760), .B(n14280), .Z(c4761) );
ANDN U23801 ( .B(n14281), .A(n14282), .Z(n14280) );
XOR U23802 ( .A(c4760), .B(b[4760]), .Z(n14281) );
XNOR U23803 ( .A(b[4760]), .B(n14282), .Z(c[4760]) );
XNOR U23804 ( .A(a[4760]), .B(c4760), .Z(n14282) );
XOR U23805 ( .A(c4761), .B(n14283), .Z(c4762) );
ANDN U23806 ( .B(n14284), .A(n14285), .Z(n14283) );
XOR U23807 ( .A(c4761), .B(b[4761]), .Z(n14284) );
XNOR U23808 ( .A(b[4761]), .B(n14285), .Z(c[4761]) );
XNOR U23809 ( .A(a[4761]), .B(c4761), .Z(n14285) );
XOR U23810 ( .A(c4762), .B(n14286), .Z(c4763) );
ANDN U23811 ( .B(n14287), .A(n14288), .Z(n14286) );
XOR U23812 ( .A(c4762), .B(b[4762]), .Z(n14287) );
XNOR U23813 ( .A(b[4762]), .B(n14288), .Z(c[4762]) );
XNOR U23814 ( .A(a[4762]), .B(c4762), .Z(n14288) );
XOR U23815 ( .A(c4763), .B(n14289), .Z(c4764) );
ANDN U23816 ( .B(n14290), .A(n14291), .Z(n14289) );
XOR U23817 ( .A(c4763), .B(b[4763]), .Z(n14290) );
XNOR U23818 ( .A(b[4763]), .B(n14291), .Z(c[4763]) );
XNOR U23819 ( .A(a[4763]), .B(c4763), .Z(n14291) );
XOR U23820 ( .A(c4764), .B(n14292), .Z(c4765) );
ANDN U23821 ( .B(n14293), .A(n14294), .Z(n14292) );
XOR U23822 ( .A(c4764), .B(b[4764]), .Z(n14293) );
XNOR U23823 ( .A(b[4764]), .B(n14294), .Z(c[4764]) );
XNOR U23824 ( .A(a[4764]), .B(c4764), .Z(n14294) );
XOR U23825 ( .A(c4765), .B(n14295), .Z(c4766) );
ANDN U23826 ( .B(n14296), .A(n14297), .Z(n14295) );
XOR U23827 ( .A(c4765), .B(b[4765]), .Z(n14296) );
XNOR U23828 ( .A(b[4765]), .B(n14297), .Z(c[4765]) );
XNOR U23829 ( .A(a[4765]), .B(c4765), .Z(n14297) );
XOR U23830 ( .A(c4766), .B(n14298), .Z(c4767) );
ANDN U23831 ( .B(n14299), .A(n14300), .Z(n14298) );
XOR U23832 ( .A(c4766), .B(b[4766]), .Z(n14299) );
XNOR U23833 ( .A(b[4766]), .B(n14300), .Z(c[4766]) );
XNOR U23834 ( .A(a[4766]), .B(c4766), .Z(n14300) );
XOR U23835 ( .A(c4767), .B(n14301), .Z(c4768) );
ANDN U23836 ( .B(n14302), .A(n14303), .Z(n14301) );
XOR U23837 ( .A(c4767), .B(b[4767]), .Z(n14302) );
XNOR U23838 ( .A(b[4767]), .B(n14303), .Z(c[4767]) );
XNOR U23839 ( .A(a[4767]), .B(c4767), .Z(n14303) );
XOR U23840 ( .A(c4768), .B(n14304), .Z(c4769) );
ANDN U23841 ( .B(n14305), .A(n14306), .Z(n14304) );
XOR U23842 ( .A(c4768), .B(b[4768]), .Z(n14305) );
XNOR U23843 ( .A(b[4768]), .B(n14306), .Z(c[4768]) );
XNOR U23844 ( .A(a[4768]), .B(c4768), .Z(n14306) );
XOR U23845 ( .A(c4769), .B(n14307), .Z(c4770) );
ANDN U23846 ( .B(n14308), .A(n14309), .Z(n14307) );
XOR U23847 ( .A(c4769), .B(b[4769]), .Z(n14308) );
XNOR U23848 ( .A(b[4769]), .B(n14309), .Z(c[4769]) );
XNOR U23849 ( .A(a[4769]), .B(c4769), .Z(n14309) );
XOR U23850 ( .A(c4770), .B(n14310), .Z(c4771) );
ANDN U23851 ( .B(n14311), .A(n14312), .Z(n14310) );
XOR U23852 ( .A(c4770), .B(b[4770]), .Z(n14311) );
XNOR U23853 ( .A(b[4770]), .B(n14312), .Z(c[4770]) );
XNOR U23854 ( .A(a[4770]), .B(c4770), .Z(n14312) );
XOR U23855 ( .A(c4771), .B(n14313), .Z(c4772) );
ANDN U23856 ( .B(n14314), .A(n14315), .Z(n14313) );
XOR U23857 ( .A(c4771), .B(b[4771]), .Z(n14314) );
XNOR U23858 ( .A(b[4771]), .B(n14315), .Z(c[4771]) );
XNOR U23859 ( .A(a[4771]), .B(c4771), .Z(n14315) );
XOR U23860 ( .A(c4772), .B(n14316), .Z(c4773) );
ANDN U23861 ( .B(n14317), .A(n14318), .Z(n14316) );
XOR U23862 ( .A(c4772), .B(b[4772]), .Z(n14317) );
XNOR U23863 ( .A(b[4772]), .B(n14318), .Z(c[4772]) );
XNOR U23864 ( .A(a[4772]), .B(c4772), .Z(n14318) );
XOR U23865 ( .A(c4773), .B(n14319), .Z(c4774) );
ANDN U23866 ( .B(n14320), .A(n14321), .Z(n14319) );
XOR U23867 ( .A(c4773), .B(b[4773]), .Z(n14320) );
XNOR U23868 ( .A(b[4773]), .B(n14321), .Z(c[4773]) );
XNOR U23869 ( .A(a[4773]), .B(c4773), .Z(n14321) );
XOR U23870 ( .A(c4774), .B(n14322), .Z(c4775) );
ANDN U23871 ( .B(n14323), .A(n14324), .Z(n14322) );
XOR U23872 ( .A(c4774), .B(b[4774]), .Z(n14323) );
XNOR U23873 ( .A(b[4774]), .B(n14324), .Z(c[4774]) );
XNOR U23874 ( .A(a[4774]), .B(c4774), .Z(n14324) );
XOR U23875 ( .A(c4775), .B(n14325), .Z(c4776) );
ANDN U23876 ( .B(n14326), .A(n14327), .Z(n14325) );
XOR U23877 ( .A(c4775), .B(b[4775]), .Z(n14326) );
XNOR U23878 ( .A(b[4775]), .B(n14327), .Z(c[4775]) );
XNOR U23879 ( .A(a[4775]), .B(c4775), .Z(n14327) );
XOR U23880 ( .A(c4776), .B(n14328), .Z(c4777) );
ANDN U23881 ( .B(n14329), .A(n14330), .Z(n14328) );
XOR U23882 ( .A(c4776), .B(b[4776]), .Z(n14329) );
XNOR U23883 ( .A(b[4776]), .B(n14330), .Z(c[4776]) );
XNOR U23884 ( .A(a[4776]), .B(c4776), .Z(n14330) );
XOR U23885 ( .A(c4777), .B(n14331), .Z(c4778) );
ANDN U23886 ( .B(n14332), .A(n14333), .Z(n14331) );
XOR U23887 ( .A(c4777), .B(b[4777]), .Z(n14332) );
XNOR U23888 ( .A(b[4777]), .B(n14333), .Z(c[4777]) );
XNOR U23889 ( .A(a[4777]), .B(c4777), .Z(n14333) );
XOR U23890 ( .A(c4778), .B(n14334), .Z(c4779) );
ANDN U23891 ( .B(n14335), .A(n14336), .Z(n14334) );
XOR U23892 ( .A(c4778), .B(b[4778]), .Z(n14335) );
XNOR U23893 ( .A(b[4778]), .B(n14336), .Z(c[4778]) );
XNOR U23894 ( .A(a[4778]), .B(c4778), .Z(n14336) );
XOR U23895 ( .A(c4779), .B(n14337), .Z(c4780) );
ANDN U23896 ( .B(n14338), .A(n14339), .Z(n14337) );
XOR U23897 ( .A(c4779), .B(b[4779]), .Z(n14338) );
XNOR U23898 ( .A(b[4779]), .B(n14339), .Z(c[4779]) );
XNOR U23899 ( .A(a[4779]), .B(c4779), .Z(n14339) );
XOR U23900 ( .A(c4780), .B(n14340), .Z(c4781) );
ANDN U23901 ( .B(n14341), .A(n14342), .Z(n14340) );
XOR U23902 ( .A(c4780), .B(b[4780]), .Z(n14341) );
XNOR U23903 ( .A(b[4780]), .B(n14342), .Z(c[4780]) );
XNOR U23904 ( .A(a[4780]), .B(c4780), .Z(n14342) );
XOR U23905 ( .A(c4781), .B(n14343), .Z(c4782) );
ANDN U23906 ( .B(n14344), .A(n14345), .Z(n14343) );
XOR U23907 ( .A(c4781), .B(b[4781]), .Z(n14344) );
XNOR U23908 ( .A(b[4781]), .B(n14345), .Z(c[4781]) );
XNOR U23909 ( .A(a[4781]), .B(c4781), .Z(n14345) );
XOR U23910 ( .A(c4782), .B(n14346), .Z(c4783) );
ANDN U23911 ( .B(n14347), .A(n14348), .Z(n14346) );
XOR U23912 ( .A(c4782), .B(b[4782]), .Z(n14347) );
XNOR U23913 ( .A(b[4782]), .B(n14348), .Z(c[4782]) );
XNOR U23914 ( .A(a[4782]), .B(c4782), .Z(n14348) );
XOR U23915 ( .A(c4783), .B(n14349), .Z(c4784) );
ANDN U23916 ( .B(n14350), .A(n14351), .Z(n14349) );
XOR U23917 ( .A(c4783), .B(b[4783]), .Z(n14350) );
XNOR U23918 ( .A(b[4783]), .B(n14351), .Z(c[4783]) );
XNOR U23919 ( .A(a[4783]), .B(c4783), .Z(n14351) );
XOR U23920 ( .A(c4784), .B(n14352), .Z(c4785) );
ANDN U23921 ( .B(n14353), .A(n14354), .Z(n14352) );
XOR U23922 ( .A(c4784), .B(b[4784]), .Z(n14353) );
XNOR U23923 ( .A(b[4784]), .B(n14354), .Z(c[4784]) );
XNOR U23924 ( .A(a[4784]), .B(c4784), .Z(n14354) );
XOR U23925 ( .A(c4785), .B(n14355), .Z(c4786) );
ANDN U23926 ( .B(n14356), .A(n14357), .Z(n14355) );
XOR U23927 ( .A(c4785), .B(b[4785]), .Z(n14356) );
XNOR U23928 ( .A(b[4785]), .B(n14357), .Z(c[4785]) );
XNOR U23929 ( .A(a[4785]), .B(c4785), .Z(n14357) );
XOR U23930 ( .A(c4786), .B(n14358), .Z(c4787) );
ANDN U23931 ( .B(n14359), .A(n14360), .Z(n14358) );
XOR U23932 ( .A(c4786), .B(b[4786]), .Z(n14359) );
XNOR U23933 ( .A(b[4786]), .B(n14360), .Z(c[4786]) );
XNOR U23934 ( .A(a[4786]), .B(c4786), .Z(n14360) );
XOR U23935 ( .A(c4787), .B(n14361), .Z(c4788) );
ANDN U23936 ( .B(n14362), .A(n14363), .Z(n14361) );
XOR U23937 ( .A(c4787), .B(b[4787]), .Z(n14362) );
XNOR U23938 ( .A(b[4787]), .B(n14363), .Z(c[4787]) );
XNOR U23939 ( .A(a[4787]), .B(c4787), .Z(n14363) );
XOR U23940 ( .A(c4788), .B(n14364), .Z(c4789) );
ANDN U23941 ( .B(n14365), .A(n14366), .Z(n14364) );
XOR U23942 ( .A(c4788), .B(b[4788]), .Z(n14365) );
XNOR U23943 ( .A(b[4788]), .B(n14366), .Z(c[4788]) );
XNOR U23944 ( .A(a[4788]), .B(c4788), .Z(n14366) );
XOR U23945 ( .A(c4789), .B(n14367), .Z(c4790) );
ANDN U23946 ( .B(n14368), .A(n14369), .Z(n14367) );
XOR U23947 ( .A(c4789), .B(b[4789]), .Z(n14368) );
XNOR U23948 ( .A(b[4789]), .B(n14369), .Z(c[4789]) );
XNOR U23949 ( .A(a[4789]), .B(c4789), .Z(n14369) );
XOR U23950 ( .A(c4790), .B(n14370), .Z(c4791) );
ANDN U23951 ( .B(n14371), .A(n14372), .Z(n14370) );
XOR U23952 ( .A(c4790), .B(b[4790]), .Z(n14371) );
XNOR U23953 ( .A(b[4790]), .B(n14372), .Z(c[4790]) );
XNOR U23954 ( .A(a[4790]), .B(c4790), .Z(n14372) );
XOR U23955 ( .A(c4791), .B(n14373), .Z(c4792) );
ANDN U23956 ( .B(n14374), .A(n14375), .Z(n14373) );
XOR U23957 ( .A(c4791), .B(b[4791]), .Z(n14374) );
XNOR U23958 ( .A(b[4791]), .B(n14375), .Z(c[4791]) );
XNOR U23959 ( .A(a[4791]), .B(c4791), .Z(n14375) );
XOR U23960 ( .A(c4792), .B(n14376), .Z(c4793) );
ANDN U23961 ( .B(n14377), .A(n14378), .Z(n14376) );
XOR U23962 ( .A(c4792), .B(b[4792]), .Z(n14377) );
XNOR U23963 ( .A(b[4792]), .B(n14378), .Z(c[4792]) );
XNOR U23964 ( .A(a[4792]), .B(c4792), .Z(n14378) );
XOR U23965 ( .A(c4793), .B(n14379), .Z(c4794) );
ANDN U23966 ( .B(n14380), .A(n14381), .Z(n14379) );
XOR U23967 ( .A(c4793), .B(b[4793]), .Z(n14380) );
XNOR U23968 ( .A(b[4793]), .B(n14381), .Z(c[4793]) );
XNOR U23969 ( .A(a[4793]), .B(c4793), .Z(n14381) );
XOR U23970 ( .A(c4794), .B(n14382), .Z(c4795) );
ANDN U23971 ( .B(n14383), .A(n14384), .Z(n14382) );
XOR U23972 ( .A(c4794), .B(b[4794]), .Z(n14383) );
XNOR U23973 ( .A(b[4794]), .B(n14384), .Z(c[4794]) );
XNOR U23974 ( .A(a[4794]), .B(c4794), .Z(n14384) );
XOR U23975 ( .A(c4795), .B(n14385), .Z(c4796) );
ANDN U23976 ( .B(n14386), .A(n14387), .Z(n14385) );
XOR U23977 ( .A(c4795), .B(b[4795]), .Z(n14386) );
XNOR U23978 ( .A(b[4795]), .B(n14387), .Z(c[4795]) );
XNOR U23979 ( .A(a[4795]), .B(c4795), .Z(n14387) );
XOR U23980 ( .A(c4796), .B(n14388), .Z(c4797) );
ANDN U23981 ( .B(n14389), .A(n14390), .Z(n14388) );
XOR U23982 ( .A(c4796), .B(b[4796]), .Z(n14389) );
XNOR U23983 ( .A(b[4796]), .B(n14390), .Z(c[4796]) );
XNOR U23984 ( .A(a[4796]), .B(c4796), .Z(n14390) );
XOR U23985 ( .A(c4797), .B(n14391), .Z(c4798) );
ANDN U23986 ( .B(n14392), .A(n14393), .Z(n14391) );
XOR U23987 ( .A(c4797), .B(b[4797]), .Z(n14392) );
XNOR U23988 ( .A(b[4797]), .B(n14393), .Z(c[4797]) );
XNOR U23989 ( .A(a[4797]), .B(c4797), .Z(n14393) );
XOR U23990 ( .A(c4798), .B(n14394), .Z(c4799) );
ANDN U23991 ( .B(n14395), .A(n14396), .Z(n14394) );
XOR U23992 ( .A(c4798), .B(b[4798]), .Z(n14395) );
XNOR U23993 ( .A(b[4798]), .B(n14396), .Z(c[4798]) );
XNOR U23994 ( .A(a[4798]), .B(c4798), .Z(n14396) );
XOR U23995 ( .A(c4799), .B(n14397), .Z(c4800) );
ANDN U23996 ( .B(n14398), .A(n14399), .Z(n14397) );
XOR U23997 ( .A(c4799), .B(b[4799]), .Z(n14398) );
XNOR U23998 ( .A(b[4799]), .B(n14399), .Z(c[4799]) );
XNOR U23999 ( .A(a[4799]), .B(c4799), .Z(n14399) );
XOR U24000 ( .A(c4800), .B(n14400), .Z(c4801) );
ANDN U24001 ( .B(n14401), .A(n14402), .Z(n14400) );
XOR U24002 ( .A(c4800), .B(b[4800]), .Z(n14401) );
XNOR U24003 ( .A(b[4800]), .B(n14402), .Z(c[4800]) );
XNOR U24004 ( .A(a[4800]), .B(c4800), .Z(n14402) );
XOR U24005 ( .A(c4801), .B(n14403), .Z(c4802) );
ANDN U24006 ( .B(n14404), .A(n14405), .Z(n14403) );
XOR U24007 ( .A(c4801), .B(b[4801]), .Z(n14404) );
XNOR U24008 ( .A(b[4801]), .B(n14405), .Z(c[4801]) );
XNOR U24009 ( .A(a[4801]), .B(c4801), .Z(n14405) );
XOR U24010 ( .A(c4802), .B(n14406), .Z(c4803) );
ANDN U24011 ( .B(n14407), .A(n14408), .Z(n14406) );
XOR U24012 ( .A(c4802), .B(b[4802]), .Z(n14407) );
XNOR U24013 ( .A(b[4802]), .B(n14408), .Z(c[4802]) );
XNOR U24014 ( .A(a[4802]), .B(c4802), .Z(n14408) );
XOR U24015 ( .A(c4803), .B(n14409), .Z(c4804) );
ANDN U24016 ( .B(n14410), .A(n14411), .Z(n14409) );
XOR U24017 ( .A(c4803), .B(b[4803]), .Z(n14410) );
XNOR U24018 ( .A(b[4803]), .B(n14411), .Z(c[4803]) );
XNOR U24019 ( .A(a[4803]), .B(c4803), .Z(n14411) );
XOR U24020 ( .A(c4804), .B(n14412), .Z(c4805) );
ANDN U24021 ( .B(n14413), .A(n14414), .Z(n14412) );
XOR U24022 ( .A(c4804), .B(b[4804]), .Z(n14413) );
XNOR U24023 ( .A(b[4804]), .B(n14414), .Z(c[4804]) );
XNOR U24024 ( .A(a[4804]), .B(c4804), .Z(n14414) );
XOR U24025 ( .A(c4805), .B(n14415), .Z(c4806) );
ANDN U24026 ( .B(n14416), .A(n14417), .Z(n14415) );
XOR U24027 ( .A(c4805), .B(b[4805]), .Z(n14416) );
XNOR U24028 ( .A(b[4805]), .B(n14417), .Z(c[4805]) );
XNOR U24029 ( .A(a[4805]), .B(c4805), .Z(n14417) );
XOR U24030 ( .A(c4806), .B(n14418), .Z(c4807) );
ANDN U24031 ( .B(n14419), .A(n14420), .Z(n14418) );
XOR U24032 ( .A(c4806), .B(b[4806]), .Z(n14419) );
XNOR U24033 ( .A(b[4806]), .B(n14420), .Z(c[4806]) );
XNOR U24034 ( .A(a[4806]), .B(c4806), .Z(n14420) );
XOR U24035 ( .A(c4807), .B(n14421), .Z(c4808) );
ANDN U24036 ( .B(n14422), .A(n14423), .Z(n14421) );
XOR U24037 ( .A(c4807), .B(b[4807]), .Z(n14422) );
XNOR U24038 ( .A(b[4807]), .B(n14423), .Z(c[4807]) );
XNOR U24039 ( .A(a[4807]), .B(c4807), .Z(n14423) );
XOR U24040 ( .A(c4808), .B(n14424), .Z(c4809) );
ANDN U24041 ( .B(n14425), .A(n14426), .Z(n14424) );
XOR U24042 ( .A(c4808), .B(b[4808]), .Z(n14425) );
XNOR U24043 ( .A(b[4808]), .B(n14426), .Z(c[4808]) );
XNOR U24044 ( .A(a[4808]), .B(c4808), .Z(n14426) );
XOR U24045 ( .A(c4809), .B(n14427), .Z(c4810) );
ANDN U24046 ( .B(n14428), .A(n14429), .Z(n14427) );
XOR U24047 ( .A(c4809), .B(b[4809]), .Z(n14428) );
XNOR U24048 ( .A(b[4809]), .B(n14429), .Z(c[4809]) );
XNOR U24049 ( .A(a[4809]), .B(c4809), .Z(n14429) );
XOR U24050 ( .A(c4810), .B(n14430), .Z(c4811) );
ANDN U24051 ( .B(n14431), .A(n14432), .Z(n14430) );
XOR U24052 ( .A(c4810), .B(b[4810]), .Z(n14431) );
XNOR U24053 ( .A(b[4810]), .B(n14432), .Z(c[4810]) );
XNOR U24054 ( .A(a[4810]), .B(c4810), .Z(n14432) );
XOR U24055 ( .A(c4811), .B(n14433), .Z(c4812) );
ANDN U24056 ( .B(n14434), .A(n14435), .Z(n14433) );
XOR U24057 ( .A(c4811), .B(b[4811]), .Z(n14434) );
XNOR U24058 ( .A(b[4811]), .B(n14435), .Z(c[4811]) );
XNOR U24059 ( .A(a[4811]), .B(c4811), .Z(n14435) );
XOR U24060 ( .A(c4812), .B(n14436), .Z(c4813) );
ANDN U24061 ( .B(n14437), .A(n14438), .Z(n14436) );
XOR U24062 ( .A(c4812), .B(b[4812]), .Z(n14437) );
XNOR U24063 ( .A(b[4812]), .B(n14438), .Z(c[4812]) );
XNOR U24064 ( .A(a[4812]), .B(c4812), .Z(n14438) );
XOR U24065 ( .A(c4813), .B(n14439), .Z(c4814) );
ANDN U24066 ( .B(n14440), .A(n14441), .Z(n14439) );
XOR U24067 ( .A(c4813), .B(b[4813]), .Z(n14440) );
XNOR U24068 ( .A(b[4813]), .B(n14441), .Z(c[4813]) );
XNOR U24069 ( .A(a[4813]), .B(c4813), .Z(n14441) );
XOR U24070 ( .A(c4814), .B(n14442), .Z(c4815) );
ANDN U24071 ( .B(n14443), .A(n14444), .Z(n14442) );
XOR U24072 ( .A(c4814), .B(b[4814]), .Z(n14443) );
XNOR U24073 ( .A(b[4814]), .B(n14444), .Z(c[4814]) );
XNOR U24074 ( .A(a[4814]), .B(c4814), .Z(n14444) );
XOR U24075 ( .A(c4815), .B(n14445), .Z(c4816) );
ANDN U24076 ( .B(n14446), .A(n14447), .Z(n14445) );
XOR U24077 ( .A(c4815), .B(b[4815]), .Z(n14446) );
XNOR U24078 ( .A(b[4815]), .B(n14447), .Z(c[4815]) );
XNOR U24079 ( .A(a[4815]), .B(c4815), .Z(n14447) );
XOR U24080 ( .A(c4816), .B(n14448), .Z(c4817) );
ANDN U24081 ( .B(n14449), .A(n14450), .Z(n14448) );
XOR U24082 ( .A(c4816), .B(b[4816]), .Z(n14449) );
XNOR U24083 ( .A(b[4816]), .B(n14450), .Z(c[4816]) );
XNOR U24084 ( .A(a[4816]), .B(c4816), .Z(n14450) );
XOR U24085 ( .A(c4817), .B(n14451), .Z(c4818) );
ANDN U24086 ( .B(n14452), .A(n14453), .Z(n14451) );
XOR U24087 ( .A(c4817), .B(b[4817]), .Z(n14452) );
XNOR U24088 ( .A(b[4817]), .B(n14453), .Z(c[4817]) );
XNOR U24089 ( .A(a[4817]), .B(c4817), .Z(n14453) );
XOR U24090 ( .A(c4818), .B(n14454), .Z(c4819) );
ANDN U24091 ( .B(n14455), .A(n14456), .Z(n14454) );
XOR U24092 ( .A(c4818), .B(b[4818]), .Z(n14455) );
XNOR U24093 ( .A(b[4818]), .B(n14456), .Z(c[4818]) );
XNOR U24094 ( .A(a[4818]), .B(c4818), .Z(n14456) );
XOR U24095 ( .A(c4819), .B(n14457), .Z(c4820) );
ANDN U24096 ( .B(n14458), .A(n14459), .Z(n14457) );
XOR U24097 ( .A(c4819), .B(b[4819]), .Z(n14458) );
XNOR U24098 ( .A(b[4819]), .B(n14459), .Z(c[4819]) );
XNOR U24099 ( .A(a[4819]), .B(c4819), .Z(n14459) );
XOR U24100 ( .A(c4820), .B(n14460), .Z(c4821) );
ANDN U24101 ( .B(n14461), .A(n14462), .Z(n14460) );
XOR U24102 ( .A(c4820), .B(b[4820]), .Z(n14461) );
XNOR U24103 ( .A(b[4820]), .B(n14462), .Z(c[4820]) );
XNOR U24104 ( .A(a[4820]), .B(c4820), .Z(n14462) );
XOR U24105 ( .A(c4821), .B(n14463), .Z(c4822) );
ANDN U24106 ( .B(n14464), .A(n14465), .Z(n14463) );
XOR U24107 ( .A(c4821), .B(b[4821]), .Z(n14464) );
XNOR U24108 ( .A(b[4821]), .B(n14465), .Z(c[4821]) );
XNOR U24109 ( .A(a[4821]), .B(c4821), .Z(n14465) );
XOR U24110 ( .A(c4822), .B(n14466), .Z(c4823) );
ANDN U24111 ( .B(n14467), .A(n14468), .Z(n14466) );
XOR U24112 ( .A(c4822), .B(b[4822]), .Z(n14467) );
XNOR U24113 ( .A(b[4822]), .B(n14468), .Z(c[4822]) );
XNOR U24114 ( .A(a[4822]), .B(c4822), .Z(n14468) );
XOR U24115 ( .A(c4823), .B(n14469), .Z(c4824) );
ANDN U24116 ( .B(n14470), .A(n14471), .Z(n14469) );
XOR U24117 ( .A(c4823), .B(b[4823]), .Z(n14470) );
XNOR U24118 ( .A(b[4823]), .B(n14471), .Z(c[4823]) );
XNOR U24119 ( .A(a[4823]), .B(c4823), .Z(n14471) );
XOR U24120 ( .A(c4824), .B(n14472), .Z(c4825) );
ANDN U24121 ( .B(n14473), .A(n14474), .Z(n14472) );
XOR U24122 ( .A(c4824), .B(b[4824]), .Z(n14473) );
XNOR U24123 ( .A(b[4824]), .B(n14474), .Z(c[4824]) );
XNOR U24124 ( .A(a[4824]), .B(c4824), .Z(n14474) );
XOR U24125 ( .A(c4825), .B(n14475), .Z(c4826) );
ANDN U24126 ( .B(n14476), .A(n14477), .Z(n14475) );
XOR U24127 ( .A(c4825), .B(b[4825]), .Z(n14476) );
XNOR U24128 ( .A(b[4825]), .B(n14477), .Z(c[4825]) );
XNOR U24129 ( .A(a[4825]), .B(c4825), .Z(n14477) );
XOR U24130 ( .A(c4826), .B(n14478), .Z(c4827) );
ANDN U24131 ( .B(n14479), .A(n14480), .Z(n14478) );
XOR U24132 ( .A(c4826), .B(b[4826]), .Z(n14479) );
XNOR U24133 ( .A(b[4826]), .B(n14480), .Z(c[4826]) );
XNOR U24134 ( .A(a[4826]), .B(c4826), .Z(n14480) );
XOR U24135 ( .A(c4827), .B(n14481), .Z(c4828) );
ANDN U24136 ( .B(n14482), .A(n14483), .Z(n14481) );
XOR U24137 ( .A(c4827), .B(b[4827]), .Z(n14482) );
XNOR U24138 ( .A(b[4827]), .B(n14483), .Z(c[4827]) );
XNOR U24139 ( .A(a[4827]), .B(c4827), .Z(n14483) );
XOR U24140 ( .A(c4828), .B(n14484), .Z(c4829) );
ANDN U24141 ( .B(n14485), .A(n14486), .Z(n14484) );
XOR U24142 ( .A(c4828), .B(b[4828]), .Z(n14485) );
XNOR U24143 ( .A(b[4828]), .B(n14486), .Z(c[4828]) );
XNOR U24144 ( .A(a[4828]), .B(c4828), .Z(n14486) );
XOR U24145 ( .A(c4829), .B(n14487), .Z(c4830) );
ANDN U24146 ( .B(n14488), .A(n14489), .Z(n14487) );
XOR U24147 ( .A(c4829), .B(b[4829]), .Z(n14488) );
XNOR U24148 ( .A(b[4829]), .B(n14489), .Z(c[4829]) );
XNOR U24149 ( .A(a[4829]), .B(c4829), .Z(n14489) );
XOR U24150 ( .A(c4830), .B(n14490), .Z(c4831) );
ANDN U24151 ( .B(n14491), .A(n14492), .Z(n14490) );
XOR U24152 ( .A(c4830), .B(b[4830]), .Z(n14491) );
XNOR U24153 ( .A(b[4830]), .B(n14492), .Z(c[4830]) );
XNOR U24154 ( .A(a[4830]), .B(c4830), .Z(n14492) );
XOR U24155 ( .A(c4831), .B(n14493), .Z(c4832) );
ANDN U24156 ( .B(n14494), .A(n14495), .Z(n14493) );
XOR U24157 ( .A(c4831), .B(b[4831]), .Z(n14494) );
XNOR U24158 ( .A(b[4831]), .B(n14495), .Z(c[4831]) );
XNOR U24159 ( .A(a[4831]), .B(c4831), .Z(n14495) );
XOR U24160 ( .A(c4832), .B(n14496), .Z(c4833) );
ANDN U24161 ( .B(n14497), .A(n14498), .Z(n14496) );
XOR U24162 ( .A(c4832), .B(b[4832]), .Z(n14497) );
XNOR U24163 ( .A(b[4832]), .B(n14498), .Z(c[4832]) );
XNOR U24164 ( .A(a[4832]), .B(c4832), .Z(n14498) );
XOR U24165 ( .A(c4833), .B(n14499), .Z(c4834) );
ANDN U24166 ( .B(n14500), .A(n14501), .Z(n14499) );
XOR U24167 ( .A(c4833), .B(b[4833]), .Z(n14500) );
XNOR U24168 ( .A(b[4833]), .B(n14501), .Z(c[4833]) );
XNOR U24169 ( .A(a[4833]), .B(c4833), .Z(n14501) );
XOR U24170 ( .A(c4834), .B(n14502), .Z(c4835) );
ANDN U24171 ( .B(n14503), .A(n14504), .Z(n14502) );
XOR U24172 ( .A(c4834), .B(b[4834]), .Z(n14503) );
XNOR U24173 ( .A(b[4834]), .B(n14504), .Z(c[4834]) );
XNOR U24174 ( .A(a[4834]), .B(c4834), .Z(n14504) );
XOR U24175 ( .A(c4835), .B(n14505), .Z(c4836) );
ANDN U24176 ( .B(n14506), .A(n14507), .Z(n14505) );
XOR U24177 ( .A(c4835), .B(b[4835]), .Z(n14506) );
XNOR U24178 ( .A(b[4835]), .B(n14507), .Z(c[4835]) );
XNOR U24179 ( .A(a[4835]), .B(c4835), .Z(n14507) );
XOR U24180 ( .A(c4836), .B(n14508), .Z(c4837) );
ANDN U24181 ( .B(n14509), .A(n14510), .Z(n14508) );
XOR U24182 ( .A(c4836), .B(b[4836]), .Z(n14509) );
XNOR U24183 ( .A(b[4836]), .B(n14510), .Z(c[4836]) );
XNOR U24184 ( .A(a[4836]), .B(c4836), .Z(n14510) );
XOR U24185 ( .A(c4837), .B(n14511), .Z(c4838) );
ANDN U24186 ( .B(n14512), .A(n14513), .Z(n14511) );
XOR U24187 ( .A(c4837), .B(b[4837]), .Z(n14512) );
XNOR U24188 ( .A(b[4837]), .B(n14513), .Z(c[4837]) );
XNOR U24189 ( .A(a[4837]), .B(c4837), .Z(n14513) );
XOR U24190 ( .A(c4838), .B(n14514), .Z(c4839) );
ANDN U24191 ( .B(n14515), .A(n14516), .Z(n14514) );
XOR U24192 ( .A(c4838), .B(b[4838]), .Z(n14515) );
XNOR U24193 ( .A(b[4838]), .B(n14516), .Z(c[4838]) );
XNOR U24194 ( .A(a[4838]), .B(c4838), .Z(n14516) );
XOR U24195 ( .A(c4839), .B(n14517), .Z(c4840) );
ANDN U24196 ( .B(n14518), .A(n14519), .Z(n14517) );
XOR U24197 ( .A(c4839), .B(b[4839]), .Z(n14518) );
XNOR U24198 ( .A(b[4839]), .B(n14519), .Z(c[4839]) );
XNOR U24199 ( .A(a[4839]), .B(c4839), .Z(n14519) );
XOR U24200 ( .A(c4840), .B(n14520), .Z(c4841) );
ANDN U24201 ( .B(n14521), .A(n14522), .Z(n14520) );
XOR U24202 ( .A(c4840), .B(b[4840]), .Z(n14521) );
XNOR U24203 ( .A(b[4840]), .B(n14522), .Z(c[4840]) );
XNOR U24204 ( .A(a[4840]), .B(c4840), .Z(n14522) );
XOR U24205 ( .A(c4841), .B(n14523), .Z(c4842) );
ANDN U24206 ( .B(n14524), .A(n14525), .Z(n14523) );
XOR U24207 ( .A(c4841), .B(b[4841]), .Z(n14524) );
XNOR U24208 ( .A(b[4841]), .B(n14525), .Z(c[4841]) );
XNOR U24209 ( .A(a[4841]), .B(c4841), .Z(n14525) );
XOR U24210 ( .A(c4842), .B(n14526), .Z(c4843) );
ANDN U24211 ( .B(n14527), .A(n14528), .Z(n14526) );
XOR U24212 ( .A(c4842), .B(b[4842]), .Z(n14527) );
XNOR U24213 ( .A(b[4842]), .B(n14528), .Z(c[4842]) );
XNOR U24214 ( .A(a[4842]), .B(c4842), .Z(n14528) );
XOR U24215 ( .A(c4843), .B(n14529), .Z(c4844) );
ANDN U24216 ( .B(n14530), .A(n14531), .Z(n14529) );
XOR U24217 ( .A(c4843), .B(b[4843]), .Z(n14530) );
XNOR U24218 ( .A(b[4843]), .B(n14531), .Z(c[4843]) );
XNOR U24219 ( .A(a[4843]), .B(c4843), .Z(n14531) );
XOR U24220 ( .A(c4844), .B(n14532), .Z(c4845) );
ANDN U24221 ( .B(n14533), .A(n14534), .Z(n14532) );
XOR U24222 ( .A(c4844), .B(b[4844]), .Z(n14533) );
XNOR U24223 ( .A(b[4844]), .B(n14534), .Z(c[4844]) );
XNOR U24224 ( .A(a[4844]), .B(c4844), .Z(n14534) );
XOR U24225 ( .A(c4845), .B(n14535), .Z(c4846) );
ANDN U24226 ( .B(n14536), .A(n14537), .Z(n14535) );
XOR U24227 ( .A(c4845), .B(b[4845]), .Z(n14536) );
XNOR U24228 ( .A(b[4845]), .B(n14537), .Z(c[4845]) );
XNOR U24229 ( .A(a[4845]), .B(c4845), .Z(n14537) );
XOR U24230 ( .A(c4846), .B(n14538), .Z(c4847) );
ANDN U24231 ( .B(n14539), .A(n14540), .Z(n14538) );
XOR U24232 ( .A(c4846), .B(b[4846]), .Z(n14539) );
XNOR U24233 ( .A(b[4846]), .B(n14540), .Z(c[4846]) );
XNOR U24234 ( .A(a[4846]), .B(c4846), .Z(n14540) );
XOR U24235 ( .A(c4847), .B(n14541), .Z(c4848) );
ANDN U24236 ( .B(n14542), .A(n14543), .Z(n14541) );
XOR U24237 ( .A(c4847), .B(b[4847]), .Z(n14542) );
XNOR U24238 ( .A(b[4847]), .B(n14543), .Z(c[4847]) );
XNOR U24239 ( .A(a[4847]), .B(c4847), .Z(n14543) );
XOR U24240 ( .A(c4848), .B(n14544), .Z(c4849) );
ANDN U24241 ( .B(n14545), .A(n14546), .Z(n14544) );
XOR U24242 ( .A(c4848), .B(b[4848]), .Z(n14545) );
XNOR U24243 ( .A(b[4848]), .B(n14546), .Z(c[4848]) );
XNOR U24244 ( .A(a[4848]), .B(c4848), .Z(n14546) );
XOR U24245 ( .A(c4849), .B(n14547), .Z(c4850) );
ANDN U24246 ( .B(n14548), .A(n14549), .Z(n14547) );
XOR U24247 ( .A(c4849), .B(b[4849]), .Z(n14548) );
XNOR U24248 ( .A(b[4849]), .B(n14549), .Z(c[4849]) );
XNOR U24249 ( .A(a[4849]), .B(c4849), .Z(n14549) );
XOR U24250 ( .A(c4850), .B(n14550), .Z(c4851) );
ANDN U24251 ( .B(n14551), .A(n14552), .Z(n14550) );
XOR U24252 ( .A(c4850), .B(b[4850]), .Z(n14551) );
XNOR U24253 ( .A(b[4850]), .B(n14552), .Z(c[4850]) );
XNOR U24254 ( .A(a[4850]), .B(c4850), .Z(n14552) );
XOR U24255 ( .A(c4851), .B(n14553), .Z(c4852) );
ANDN U24256 ( .B(n14554), .A(n14555), .Z(n14553) );
XOR U24257 ( .A(c4851), .B(b[4851]), .Z(n14554) );
XNOR U24258 ( .A(b[4851]), .B(n14555), .Z(c[4851]) );
XNOR U24259 ( .A(a[4851]), .B(c4851), .Z(n14555) );
XOR U24260 ( .A(c4852), .B(n14556), .Z(c4853) );
ANDN U24261 ( .B(n14557), .A(n14558), .Z(n14556) );
XOR U24262 ( .A(c4852), .B(b[4852]), .Z(n14557) );
XNOR U24263 ( .A(b[4852]), .B(n14558), .Z(c[4852]) );
XNOR U24264 ( .A(a[4852]), .B(c4852), .Z(n14558) );
XOR U24265 ( .A(c4853), .B(n14559), .Z(c4854) );
ANDN U24266 ( .B(n14560), .A(n14561), .Z(n14559) );
XOR U24267 ( .A(c4853), .B(b[4853]), .Z(n14560) );
XNOR U24268 ( .A(b[4853]), .B(n14561), .Z(c[4853]) );
XNOR U24269 ( .A(a[4853]), .B(c4853), .Z(n14561) );
XOR U24270 ( .A(c4854), .B(n14562), .Z(c4855) );
ANDN U24271 ( .B(n14563), .A(n14564), .Z(n14562) );
XOR U24272 ( .A(c4854), .B(b[4854]), .Z(n14563) );
XNOR U24273 ( .A(b[4854]), .B(n14564), .Z(c[4854]) );
XNOR U24274 ( .A(a[4854]), .B(c4854), .Z(n14564) );
XOR U24275 ( .A(c4855), .B(n14565), .Z(c4856) );
ANDN U24276 ( .B(n14566), .A(n14567), .Z(n14565) );
XOR U24277 ( .A(c4855), .B(b[4855]), .Z(n14566) );
XNOR U24278 ( .A(b[4855]), .B(n14567), .Z(c[4855]) );
XNOR U24279 ( .A(a[4855]), .B(c4855), .Z(n14567) );
XOR U24280 ( .A(c4856), .B(n14568), .Z(c4857) );
ANDN U24281 ( .B(n14569), .A(n14570), .Z(n14568) );
XOR U24282 ( .A(c4856), .B(b[4856]), .Z(n14569) );
XNOR U24283 ( .A(b[4856]), .B(n14570), .Z(c[4856]) );
XNOR U24284 ( .A(a[4856]), .B(c4856), .Z(n14570) );
XOR U24285 ( .A(c4857), .B(n14571), .Z(c4858) );
ANDN U24286 ( .B(n14572), .A(n14573), .Z(n14571) );
XOR U24287 ( .A(c4857), .B(b[4857]), .Z(n14572) );
XNOR U24288 ( .A(b[4857]), .B(n14573), .Z(c[4857]) );
XNOR U24289 ( .A(a[4857]), .B(c4857), .Z(n14573) );
XOR U24290 ( .A(c4858), .B(n14574), .Z(c4859) );
ANDN U24291 ( .B(n14575), .A(n14576), .Z(n14574) );
XOR U24292 ( .A(c4858), .B(b[4858]), .Z(n14575) );
XNOR U24293 ( .A(b[4858]), .B(n14576), .Z(c[4858]) );
XNOR U24294 ( .A(a[4858]), .B(c4858), .Z(n14576) );
XOR U24295 ( .A(c4859), .B(n14577), .Z(c4860) );
ANDN U24296 ( .B(n14578), .A(n14579), .Z(n14577) );
XOR U24297 ( .A(c4859), .B(b[4859]), .Z(n14578) );
XNOR U24298 ( .A(b[4859]), .B(n14579), .Z(c[4859]) );
XNOR U24299 ( .A(a[4859]), .B(c4859), .Z(n14579) );
XOR U24300 ( .A(c4860), .B(n14580), .Z(c4861) );
ANDN U24301 ( .B(n14581), .A(n14582), .Z(n14580) );
XOR U24302 ( .A(c4860), .B(b[4860]), .Z(n14581) );
XNOR U24303 ( .A(b[4860]), .B(n14582), .Z(c[4860]) );
XNOR U24304 ( .A(a[4860]), .B(c4860), .Z(n14582) );
XOR U24305 ( .A(c4861), .B(n14583), .Z(c4862) );
ANDN U24306 ( .B(n14584), .A(n14585), .Z(n14583) );
XOR U24307 ( .A(c4861), .B(b[4861]), .Z(n14584) );
XNOR U24308 ( .A(b[4861]), .B(n14585), .Z(c[4861]) );
XNOR U24309 ( .A(a[4861]), .B(c4861), .Z(n14585) );
XOR U24310 ( .A(c4862), .B(n14586), .Z(c4863) );
ANDN U24311 ( .B(n14587), .A(n14588), .Z(n14586) );
XOR U24312 ( .A(c4862), .B(b[4862]), .Z(n14587) );
XNOR U24313 ( .A(b[4862]), .B(n14588), .Z(c[4862]) );
XNOR U24314 ( .A(a[4862]), .B(c4862), .Z(n14588) );
XOR U24315 ( .A(c4863), .B(n14589), .Z(c4864) );
ANDN U24316 ( .B(n14590), .A(n14591), .Z(n14589) );
XOR U24317 ( .A(c4863), .B(b[4863]), .Z(n14590) );
XNOR U24318 ( .A(b[4863]), .B(n14591), .Z(c[4863]) );
XNOR U24319 ( .A(a[4863]), .B(c4863), .Z(n14591) );
XOR U24320 ( .A(c4864), .B(n14592), .Z(c4865) );
ANDN U24321 ( .B(n14593), .A(n14594), .Z(n14592) );
XOR U24322 ( .A(c4864), .B(b[4864]), .Z(n14593) );
XNOR U24323 ( .A(b[4864]), .B(n14594), .Z(c[4864]) );
XNOR U24324 ( .A(a[4864]), .B(c4864), .Z(n14594) );
XOR U24325 ( .A(c4865), .B(n14595), .Z(c4866) );
ANDN U24326 ( .B(n14596), .A(n14597), .Z(n14595) );
XOR U24327 ( .A(c4865), .B(b[4865]), .Z(n14596) );
XNOR U24328 ( .A(b[4865]), .B(n14597), .Z(c[4865]) );
XNOR U24329 ( .A(a[4865]), .B(c4865), .Z(n14597) );
XOR U24330 ( .A(c4866), .B(n14598), .Z(c4867) );
ANDN U24331 ( .B(n14599), .A(n14600), .Z(n14598) );
XOR U24332 ( .A(c4866), .B(b[4866]), .Z(n14599) );
XNOR U24333 ( .A(b[4866]), .B(n14600), .Z(c[4866]) );
XNOR U24334 ( .A(a[4866]), .B(c4866), .Z(n14600) );
XOR U24335 ( .A(c4867), .B(n14601), .Z(c4868) );
ANDN U24336 ( .B(n14602), .A(n14603), .Z(n14601) );
XOR U24337 ( .A(c4867), .B(b[4867]), .Z(n14602) );
XNOR U24338 ( .A(b[4867]), .B(n14603), .Z(c[4867]) );
XNOR U24339 ( .A(a[4867]), .B(c4867), .Z(n14603) );
XOR U24340 ( .A(c4868), .B(n14604), .Z(c4869) );
ANDN U24341 ( .B(n14605), .A(n14606), .Z(n14604) );
XOR U24342 ( .A(c4868), .B(b[4868]), .Z(n14605) );
XNOR U24343 ( .A(b[4868]), .B(n14606), .Z(c[4868]) );
XNOR U24344 ( .A(a[4868]), .B(c4868), .Z(n14606) );
XOR U24345 ( .A(c4869), .B(n14607), .Z(c4870) );
ANDN U24346 ( .B(n14608), .A(n14609), .Z(n14607) );
XOR U24347 ( .A(c4869), .B(b[4869]), .Z(n14608) );
XNOR U24348 ( .A(b[4869]), .B(n14609), .Z(c[4869]) );
XNOR U24349 ( .A(a[4869]), .B(c4869), .Z(n14609) );
XOR U24350 ( .A(c4870), .B(n14610), .Z(c4871) );
ANDN U24351 ( .B(n14611), .A(n14612), .Z(n14610) );
XOR U24352 ( .A(c4870), .B(b[4870]), .Z(n14611) );
XNOR U24353 ( .A(b[4870]), .B(n14612), .Z(c[4870]) );
XNOR U24354 ( .A(a[4870]), .B(c4870), .Z(n14612) );
XOR U24355 ( .A(c4871), .B(n14613), .Z(c4872) );
ANDN U24356 ( .B(n14614), .A(n14615), .Z(n14613) );
XOR U24357 ( .A(c4871), .B(b[4871]), .Z(n14614) );
XNOR U24358 ( .A(b[4871]), .B(n14615), .Z(c[4871]) );
XNOR U24359 ( .A(a[4871]), .B(c4871), .Z(n14615) );
XOR U24360 ( .A(c4872), .B(n14616), .Z(c4873) );
ANDN U24361 ( .B(n14617), .A(n14618), .Z(n14616) );
XOR U24362 ( .A(c4872), .B(b[4872]), .Z(n14617) );
XNOR U24363 ( .A(b[4872]), .B(n14618), .Z(c[4872]) );
XNOR U24364 ( .A(a[4872]), .B(c4872), .Z(n14618) );
XOR U24365 ( .A(c4873), .B(n14619), .Z(c4874) );
ANDN U24366 ( .B(n14620), .A(n14621), .Z(n14619) );
XOR U24367 ( .A(c4873), .B(b[4873]), .Z(n14620) );
XNOR U24368 ( .A(b[4873]), .B(n14621), .Z(c[4873]) );
XNOR U24369 ( .A(a[4873]), .B(c4873), .Z(n14621) );
XOR U24370 ( .A(c4874), .B(n14622), .Z(c4875) );
ANDN U24371 ( .B(n14623), .A(n14624), .Z(n14622) );
XOR U24372 ( .A(c4874), .B(b[4874]), .Z(n14623) );
XNOR U24373 ( .A(b[4874]), .B(n14624), .Z(c[4874]) );
XNOR U24374 ( .A(a[4874]), .B(c4874), .Z(n14624) );
XOR U24375 ( .A(c4875), .B(n14625), .Z(c4876) );
ANDN U24376 ( .B(n14626), .A(n14627), .Z(n14625) );
XOR U24377 ( .A(c4875), .B(b[4875]), .Z(n14626) );
XNOR U24378 ( .A(b[4875]), .B(n14627), .Z(c[4875]) );
XNOR U24379 ( .A(a[4875]), .B(c4875), .Z(n14627) );
XOR U24380 ( .A(c4876), .B(n14628), .Z(c4877) );
ANDN U24381 ( .B(n14629), .A(n14630), .Z(n14628) );
XOR U24382 ( .A(c4876), .B(b[4876]), .Z(n14629) );
XNOR U24383 ( .A(b[4876]), .B(n14630), .Z(c[4876]) );
XNOR U24384 ( .A(a[4876]), .B(c4876), .Z(n14630) );
XOR U24385 ( .A(c4877), .B(n14631), .Z(c4878) );
ANDN U24386 ( .B(n14632), .A(n14633), .Z(n14631) );
XOR U24387 ( .A(c4877), .B(b[4877]), .Z(n14632) );
XNOR U24388 ( .A(b[4877]), .B(n14633), .Z(c[4877]) );
XNOR U24389 ( .A(a[4877]), .B(c4877), .Z(n14633) );
XOR U24390 ( .A(c4878), .B(n14634), .Z(c4879) );
ANDN U24391 ( .B(n14635), .A(n14636), .Z(n14634) );
XOR U24392 ( .A(c4878), .B(b[4878]), .Z(n14635) );
XNOR U24393 ( .A(b[4878]), .B(n14636), .Z(c[4878]) );
XNOR U24394 ( .A(a[4878]), .B(c4878), .Z(n14636) );
XOR U24395 ( .A(c4879), .B(n14637), .Z(c4880) );
ANDN U24396 ( .B(n14638), .A(n14639), .Z(n14637) );
XOR U24397 ( .A(c4879), .B(b[4879]), .Z(n14638) );
XNOR U24398 ( .A(b[4879]), .B(n14639), .Z(c[4879]) );
XNOR U24399 ( .A(a[4879]), .B(c4879), .Z(n14639) );
XOR U24400 ( .A(c4880), .B(n14640), .Z(c4881) );
ANDN U24401 ( .B(n14641), .A(n14642), .Z(n14640) );
XOR U24402 ( .A(c4880), .B(b[4880]), .Z(n14641) );
XNOR U24403 ( .A(b[4880]), .B(n14642), .Z(c[4880]) );
XNOR U24404 ( .A(a[4880]), .B(c4880), .Z(n14642) );
XOR U24405 ( .A(c4881), .B(n14643), .Z(c4882) );
ANDN U24406 ( .B(n14644), .A(n14645), .Z(n14643) );
XOR U24407 ( .A(c4881), .B(b[4881]), .Z(n14644) );
XNOR U24408 ( .A(b[4881]), .B(n14645), .Z(c[4881]) );
XNOR U24409 ( .A(a[4881]), .B(c4881), .Z(n14645) );
XOR U24410 ( .A(c4882), .B(n14646), .Z(c4883) );
ANDN U24411 ( .B(n14647), .A(n14648), .Z(n14646) );
XOR U24412 ( .A(c4882), .B(b[4882]), .Z(n14647) );
XNOR U24413 ( .A(b[4882]), .B(n14648), .Z(c[4882]) );
XNOR U24414 ( .A(a[4882]), .B(c4882), .Z(n14648) );
XOR U24415 ( .A(c4883), .B(n14649), .Z(c4884) );
ANDN U24416 ( .B(n14650), .A(n14651), .Z(n14649) );
XOR U24417 ( .A(c4883), .B(b[4883]), .Z(n14650) );
XNOR U24418 ( .A(b[4883]), .B(n14651), .Z(c[4883]) );
XNOR U24419 ( .A(a[4883]), .B(c4883), .Z(n14651) );
XOR U24420 ( .A(c4884), .B(n14652), .Z(c4885) );
ANDN U24421 ( .B(n14653), .A(n14654), .Z(n14652) );
XOR U24422 ( .A(c4884), .B(b[4884]), .Z(n14653) );
XNOR U24423 ( .A(b[4884]), .B(n14654), .Z(c[4884]) );
XNOR U24424 ( .A(a[4884]), .B(c4884), .Z(n14654) );
XOR U24425 ( .A(c4885), .B(n14655), .Z(c4886) );
ANDN U24426 ( .B(n14656), .A(n14657), .Z(n14655) );
XOR U24427 ( .A(c4885), .B(b[4885]), .Z(n14656) );
XNOR U24428 ( .A(b[4885]), .B(n14657), .Z(c[4885]) );
XNOR U24429 ( .A(a[4885]), .B(c4885), .Z(n14657) );
XOR U24430 ( .A(c4886), .B(n14658), .Z(c4887) );
ANDN U24431 ( .B(n14659), .A(n14660), .Z(n14658) );
XOR U24432 ( .A(c4886), .B(b[4886]), .Z(n14659) );
XNOR U24433 ( .A(b[4886]), .B(n14660), .Z(c[4886]) );
XNOR U24434 ( .A(a[4886]), .B(c4886), .Z(n14660) );
XOR U24435 ( .A(c4887), .B(n14661), .Z(c4888) );
ANDN U24436 ( .B(n14662), .A(n14663), .Z(n14661) );
XOR U24437 ( .A(c4887), .B(b[4887]), .Z(n14662) );
XNOR U24438 ( .A(b[4887]), .B(n14663), .Z(c[4887]) );
XNOR U24439 ( .A(a[4887]), .B(c4887), .Z(n14663) );
XOR U24440 ( .A(c4888), .B(n14664), .Z(c4889) );
ANDN U24441 ( .B(n14665), .A(n14666), .Z(n14664) );
XOR U24442 ( .A(c4888), .B(b[4888]), .Z(n14665) );
XNOR U24443 ( .A(b[4888]), .B(n14666), .Z(c[4888]) );
XNOR U24444 ( .A(a[4888]), .B(c4888), .Z(n14666) );
XOR U24445 ( .A(c4889), .B(n14667), .Z(c4890) );
ANDN U24446 ( .B(n14668), .A(n14669), .Z(n14667) );
XOR U24447 ( .A(c4889), .B(b[4889]), .Z(n14668) );
XNOR U24448 ( .A(b[4889]), .B(n14669), .Z(c[4889]) );
XNOR U24449 ( .A(a[4889]), .B(c4889), .Z(n14669) );
XOR U24450 ( .A(c4890), .B(n14670), .Z(c4891) );
ANDN U24451 ( .B(n14671), .A(n14672), .Z(n14670) );
XOR U24452 ( .A(c4890), .B(b[4890]), .Z(n14671) );
XNOR U24453 ( .A(b[4890]), .B(n14672), .Z(c[4890]) );
XNOR U24454 ( .A(a[4890]), .B(c4890), .Z(n14672) );
XOR U24455 ( .A(c4891), .B(n14673), .Z(c4892) );
ANDN U24456 ( .B(n14674), .A(n14675), .Z(n14673) );
XOR U24457 ( .A(c4891), .B(b[4891]), .Z(n14674) );
XNOR U24458 ( .A(b[4891]), .B(n14675), .Z(c[4891]) );
XNOR U24459 ( .A(a[4891]), .B(c4891), .Z(n14675) );
XOR U24460 ( .A(c4892), .B(n14676), .Z(c4893) );
ANDN U24461 ( .B(n14677), .A(n14678), .Z(n14676) );
XOR U24462 ( .A(c4892), .B(b[4892]), .Z(n14677) );
XNOR U24463 ( .A(b[4892]), .B(n14678), .Z(c[4892]) );
XNOR U24464 ( .A(a[4892]), .B(c4892), .Z(n14678) );
XOR U24465 ( .A(c4893), .B(n14679), .Z(c4894) );
ANDN U24466 ( .B(n14680), .A(n14681), .Z(n14679) );
XOR U24467 ( .A(c4893), .B(b[4893]), .Z(n14680) );
XNOR U24468 ( .A(b[4893]), .B(n14681), .Z(c[4893]) );
XNOR U24469 ( .A(a[4893]), .B(c4893), .Z(n14681) );
XOR U24470 ( .A(c4894), .B(n14682), .Z(c4895) );
ANDN U24471 ( .B(n14683), .A(n14684), .Z(n14682) );
XOR U24472 ( .A(c4894), .B(b[4894]), .Z(n14683) );
XNOR U24473 ( .A(b[4894]), .B(n14684), .Z(c[4894]) );
XNOR U24474 ( .A(a[4894]), .B(c4894), .Z(n14684) );
XOR U24475 ( .A(c4895), .B(n14685), .Z(c4896) );
ANDN U24476 ( .B(n14686), .A(n14687), .Z(n14685) );
XOR U24477 ( .A(c4895), .B(b[4895]), .Z(n14686) );
XNOR U24478 ( .A(b[4895]), .B(n14687), .Z(c[4895]) );
XNOR U24479 ( .A(a[4895]), .B(c4895), .Z(n14687) );
XOR U24480 ( .A(c4896), .B(n14688), .Z(c4897) );
ANDN U24481 ( .B(n14689), .A(n14690), .Z(n14688) );
XOR U24482 ( .A(c4896), .B(b[4896]), .Z(n14689) );
XNOR U24483 ( .A(b[4896]), .B(n14690), .Z(c[4896]) );
XNOR U24484 ( .A(a[4896]), .B(c4896), .Z(n14690) );
XOR U24485 ( .A(c4897), .B(n14691), .Z(c4898) );
ANDN U24486 ( .B(n14692), .A(n14693), .Z(n14691) );
XOR U24487 ( .A(c4897), .B(b[4897]), .Z(n14692) );
XNOR U24488 ( .A(b[4897]), .B(n14693), .Z(c[4897]) );
XNOR U24489 ( .A(a[4897]), .B(c4897), .Z(n14693) );
XOR U24490 ( .A(c4898), .B(n14694), .Z(c4899) );
ANDN U24491 ( .B(n14695), .A(n14696), .Z(n14694) );
XOR U24492 ( .A(c4898), .B(b[4898]), .Z(n14695) );
XNOR U24493 ( .A(b[4898]), .B(n14696), .Z(c[4898]) );
XNOR U24494 ( .A(a[4898]), .B(c4898), .Z(n14696) );
XOR U24495 ( .A(c4899), .B(n14697), .Z(c4900) );
ANDN U24496 ( .B(n14698), .A(n14699), .Z(n14697) );
XOR U24497 ( .A(c4899), .B(b[4899]), .Z(n14698) );
XNOR U24498 ( .A(b[4899]), .B(n14699), .Z(c[4899]) );
XNOR U24499 ( .A(a[4899]), .B(c4899), .Z(n14699) );
XOR U24500 ( .A(c4900), .B(n14700), .Z(c4901) );
ANDN U24501 ( .B(n14701), .A(n14702), .Z(n14700) );
XOR U24502 ( .A(c4900), .B(b[4900]), .Z(n14701) );
XNOR U24503 ( .A(b[4900]), .B(n14702), .Z(c[4900]) );
XNOR U24504 ( .A(a[4900]), .B(c4900), .Z(n14702) );
XOR U24505 ( .A(c4901), .B(n14703), .Z(c4902) );
ANDN U24506 ( .B(n14704), .A(n14705), .Z(n14703) );
XOR U24507 ( .A(c4901), .B(b[4901]), .Z(n14704) );
XNOR U24508 ( .A(b[4901]), .B(n14705), .Z(c[4901]) );
XNOR U24509 ( .A(a[4901]), .B(c4901), .Z(n14705) );
XOR U24510 ( .A(c4902), .B(n14706), .Z(c4903) );
ANDN U24511 ( .B(n14707), .A(n14708), .Z(n14706) );
XOR U24512 ( .A(c4902), .B(b[4902]), .Z(n14707) );
XNOR U24513 ( .A(b[4902]), .B(n14708), .Z(c[4902]) );
XNOR U24514 ( .A(a[4902]), .B(c4902), .Z(n14708) );
XOR U24515 ( .A(c4903), .B(n14709), .Z(c4904) );
ANDN U24516 ( .B(n14710), .A(n14711), .Z(n14709) );
XOR U24517 ( .A(c4903), .B(b[4903]), .Z(n14710) );
XNOR U24518 ( .A(b[4903]), .B(n14711), .Z(c[4903]) );
XNOR U24519 ( .A(a[4903]), .B(c4903), .Z(n14711) );
XOR U24520 ( .A(c4904), .B(n14712), .Z(c4905) );
ANDN U24521 ( .B(n14713), .A(n14714), .Z(n14712) );
XOR U24522 ( .A(c4904), .B(b[4904]), .Z(n14713) );
XNOR U24523 ( .A(b[4904]), .B(n14714), .Z(c[4904]) );
XNOR U24524 ( .A(a[4904]), .B(c4904), .Z(n14714) );
XOR U24525 ( .A(c4905), .B(n14715), .Z(c4906) );
ANDN U24526 ( .B(n14716), .A(n14717), .Z(n14715) );
XOR U24527 ( .A(c4905), .B(b[4905]), .Z(n14716) );
XNOR U24528 ( .A(b[4905]), .B(n14717), .Z(c[4905]) );
XNOR U24529 ( .A(a[4905]), .B(c4905), .Z(n14717) );
XOR U24530 ( .A(c4906), .B(n14718), .Z(c4907) );
ANDN U24531 ( .B(n14719), .A(n14720), .Z(n14718) );
XOR U24532 ( .A(c4906), .B(b[4906]), .Z(n14719) );
XNOR U24533 ( .A(b[4906]), .B(n14720), .Z(c[4906]) );
XNOR U24534 ( .A(a[4906]), .B(c4906), .Z(n14720) );
XOR U24535 ( .A(c4907), .B(n14721), .Z(c4908) );
ANDN U24536 ( .B(n14722), .A(n14723), .Z(n14721) );
XOR U24537 ( .A(c4907), .B(b[4907]), .Z(n14722) );
XNOR U24538 ( .A(b[4907]), .B(n14723), .Z(c[4907]) );
XNOR U24539 ( .A(a[4907]), .B(c4907), .Z(n14723) );
XOR U24540 ( .A(c4908), .B(n14724), .Z(c4909) );
ANDN U24541 ( .B(n14725), .A(n14726), .Z(n14724) );
XOR U24542 ( .A(c4908), .B(b[4908]), .Z(n14725) );
XNOR U24543 ( .A(b[4908]), .B(n14726), .Z(c[4908]) );
XNOR U24544 ( .A(a[4908]), .B(c4908), .Z(n14726) );
XOR U24545 ( .A(c4909), .B(n14727), .Z(c4910) );
ANDN U24546 ( .B(n14728), .A(n14729), .Z(n14727) );
XOR U24547 ( .A(c4909), .B(b[4909]), .Z(n14728) );
XNOR U24548 ( .A(b[4909]), .B(n14729), .Z(c[4909]) );
XNOR U24549 ( .A(a[4909]), .B(c4909), .Z(n14729) );
XOR U24550 ( .A(c4910), .B(n14730), .Z(c4911) );
ANDN U24551 ( .B(n14731), .A(n14732), .Z(n14730) );
XOR U24552 ( .A(c4910), .B(b[4910]), .Z(n14731) );
XNOR U24553 ( .A(b[4910]), .B(n14732), .Z(c[4910]) );
XNOR U24554 ( .A(a[4910]), .B(c4910), .Z(n14732) );
XOR U24555 ( .A(c4911), .B(n14733), .Z(c4912) );
ANDN U24556 ( .B(n14734), .A(n14735), .Z(n14733) );
XOR U24557 ( .A(c4911), .B(b[4911]), .Z(n14734) );
XNOR U24558 ( .A(b[4911]), .B(n14735), .Z(c[4911]) );
XNOR U24559 ( .A(a[4911]), .B(c4911), .Z(n14735) );
XOR U24560 ( .A(c4912), .B(n14736), .Z(c4913) );
ANDN U24561 ( .B(n14737), .A(n14738), .Z(n14736) );
XOR U24562 ( .A(c4912), .B(b[4912]), .Z(n14737) );
XNOR U24563 ( .A(b[4912]), .B(n14738), .Z(c[4912]) );
XNOR U24564 ( .A(a[4912]), .B(c4912), .Z(n14738) );
XOR U24565 ( .A(c4913), .B(n14739), .Z(c4914) );
ANDN U24566 ( .B(n14740), .A(n14741), .Z(n14739) );
XOR U24567 ( .A(c4913), .B(b[4913]), .Z(n14740) );
XNOR U24568 ( .A(b[4913]), .B(n14741), .Z(c[4913]) );
XNOR U24569 ( .A(a[4913]), .B(c4913), .Z(n14741) );
XOR U24570 ( .A(c4914), .B(n14742), .Z(c4915) );
ANDN U24571 ( .B(n14743), .A(n14744), .Z(n14742) );
XOR U24572 ( .A(c4914), .B(b[4914]), .Z(n14743) );
XNOR U24573 ( .A(b[4914]), .B(n14744), .Z(c[4914]) );
XNOR U24574 ( .A(a[4914]), .B(c4914), .Z(n14744) );
XOR U24575 ( .A(c4915), .B(n14745), .Z(c4916) );
ANDN U24576 ( .B(n14746), .A(n14747), .Z(n14745) );
XOR U24577 ( .A(c4915), .B(b[4915]), .Z(n14746) );
XNOR U24578 ( .A(b[4915]), .B(n14747), .Z(c[4915]) );
XNOR U24579 ( .A(a[4915]), .B(c4915), .Z(n14747) );
XOR U24580 ( .A(c4916), .B(n14748), .Z(c4917) );
ANDN U24581 ( .B(n14749), .A(n14750), .Z(n14748) );
XOR U24582 ( .A(c4916), .B(b[4916]), .Z(n14749) );
XNOR U24583 ( .A(b[4916]), .B(n14750), .Z(c[4916]) );
XNOR U24584 ( .A(a[4916]), .B(c4916), .Z(n14750) );
XOR U24585 ( .A(c4917), .B(n14751), .Z(c4918) );
ANDN U24586 ( .B(n14752), .A(n14753), .Z(n14751) );
XOR U24587 ( .A(c4917), .B(b[4917]), .Z(n14752) );
XNOR U24588 ( .A(b[4917]), .B(n14753), .Z(c[4917]) );
XNOR U24589 ( .A(a[4917]), .B(c4917), .Z(n14753) );
XOR U24590 ( .A(c4918), .B(n14754), .Z(c4919) );
ANDN U24591 ( .B(n14755), .A(n14756), .Z(n14754) );
XOR U24592 ( .A(c4918), .B(b[4918]), .Z(n14755) );
XNOR U24593 ( .A(b[4918]), .B(n14756), .Z(c[4918]) );
XNOR U24594 ( .A(a[4918]), .B(c4918), .Z(n14756) );
XOR U24595 ( .A(c4919), .B(n14757), .Z(c4920) );
ANDN U24596 ( .B(n14758), .A(n14759), .Z(n14757) );
XOR U24597 ( .A(c4919), .B(b[4919]), .Z(n14758) );
XNOR U24598 ( .A(b[4919]), .B(n14759), .Z(c[4919]) );
XNOR U24599 ( .A(a[4919]), .B(c4919), .Z(n14759) );
XOR U24600 ( .A(c4920), .B(n14760), .Z(c4921) );
ANDN U24601 ( .B(n14761), .A(n14762), .Z(n14760) );
XOR U24602 ( .A(c4920), .B(b[4920]), .Z(n14761) );
XNOR U24603 ( .A(b[4920]), .B(n14762), .Z(c[4920]) );
XNOR U24604 ( .A(a[4920]), .B(c4920), .Z(n14762) );
XOR U24605 ( .A(c4921), .B(n14763), .Z(c4922) );
ANDN U24606 ( .B(n14764), .A(n14765), .Z(n14763) );
XOR U24607 ( .A(c4921), .B(b[4921]), .Z(n14764) );
XNOR U24608 ( .A(b[4921]), .B(n14765), .Z(c[4921]) );
XNOR U24609 ( .A(a[4921]), .B(c4921), .Z(n14765) );
XOR U24610 ( .A(c4922), .B(n14766), .Z(c4923) );
ANDN U24611 ( .B(n14767), .A(n14768), .Z(n14766) );
XOR U24612 ( .A(c4922), .B(b[4922]), .Z(n14767) );
XNOR U24613 ( .A(b[4922]), .B(n14768), .Z(c[4922]) );
XNOR U24614 ( .A(a[4922]), .B(c4922), .Z(n14768) );
XOR U24615 ( .A(c4923), .B(n14769), .Z(c4924) );
ANDN U24616 ( .B(n14770), .A(n14771), .Z(n14769) );
XOR U24617 ( .A(c4923), .B(b[4923]), .Z(n14770) );
XNOR U24618 ( .A(b[4923]), .B(n14771), .Z(c[4923]) );
XNOR U24619 ( .A(a[4923]), .B(c4923), .Z(n14771) );
XOR U24620 ( .A(c4924), .B(n14772), .Z(c4925) );
ANDN U24621 ( .B(n14773), .A(n14774), .Z(n14772) );
XOR U24622 ( .A(c4924), .B(b[4924]), .Z(n14773) );
XNOR U24623 ( .A(b[4924]), .B(n14774), .Z(c[4924]) );
XNOR U24624 ( .A(a[4924]), .B(c4924), .Z(n14774) );
XOR U24625 ( .A(c4925), .B(n14775), .Z(c4926) );
ANDN U24626 ( .B(n14776), .A(n14777), .Z(n14775) );
XOR U24627 ( .A(c4925), .B(b[4925]), .Z(n14776) );
XNOR U24628 ( .A(b[4925]), .B(n14777), .Z(c[4925]) );
XNOR U24629 ( .A(a[4925]), .B(c4925), .Z(n14777) );
XOR U24630 ( .A(c4926), .B(n14778), .Z(c4927) );
ANDN U24631 ( .B(n14779), .A(n14780), .Z(n14778) );
XOR U24632 ( .A(c4926), .B(b[4926]), .Z(n14779) );
XNOR U24633 ( .A(b[4926]), .B(n14780), .Z(c[4926]) );
XNOR U24634 ( .A(a[4926]), .B(c4926), .Z(n14780) );
XOR U24635 ( .A(c4927), .B(n14781), .Z(c4928) );
ANDN U24636 ( .B(n14782), .A(n14783), .Z(n14781) );
XOR U24637 ( .A(c4927), .B(b[4927]), .Z(n14782) );
XNOR U24638 ( .A(b[4927]), .B(n14783), .Z(c[4927]) );
XNOR U24639 ( .A(a[4927]), .B(c4927), .Z(n14783) );
XOR U24640 ( .A(c4928), .B(n14784), .Z(c4929) );
ANDN U24641 ( .B(n14785), .A(n14786), .Z(n14784) );
XOR U24642 ( .A(c4928), .B(b[4928]), .Z(n14785) );
XNOR U24643 ( .A(b[4928]), .B(n14786), .Z(c[4928]) );
XNOR U24644 ( .A(a[4928]), .B(c4928), .Z(n14786) );
XOR U24645 ( .A(c4929), .B(n14787), .Z(c4930) );
ANDN U24646 ( .B(n14788), .A(n14789), .Z(n14787) );
XOR U24647 ( .A(c4929), .B(b[4929]), .Z(n14788) );
XNOR U24648 ( .A(b[4929]), .B(n14789), .Z(c[4929]) );
XNOR U24649 ( .A(a[4929]), .B(c4929), .Z(n14789) );
XOR U24650 ( .A(c4930), .B(n14790), .Z(c4931) );
ANDN U24651 ( .B(n14791), .A(n14792), .Z(n14790) );
XOR U24652 ( .A(c4930), .B(b[4930]), .Z(n14791) );
XNOR U24653 ( .A(b[4930]), .B(n14792), .Z(c[4930]) );
XNOR U24654 ( .A(a[4930]), .B(c4930), .Z(n14792) );
XOR U24655 ( .A(c4931), .B(n14793), .Z(c4932) );
ANDN U24656 ( .B(n14794), .A(n14795), .Z(n14793) );
XOR U24657 ( .A(c4931), .B(b[4931]), .Z(n14794) );
XNOR U24658 ( .A(b[4931]), .B(n14795), .Z(c[4931]) );
XNOR U24659 ( .A(a[4931]), .B(c4931), .Z(n14795) );
XOR U24660 ( .A(c4932), .B(n14796), .Z(c4933) );
ANDN U24661 ( .B(n14797), .A(n14798), .Z(n14796) );
XOR U24662 ( .A(c4932), .B(b[4932]), .Z(n14797) );
XNOR U24663 ( .A(b[4932]), .B(n14798), .Z(c[4932]) );
XNOR U24664 ( .A(a[4932]), .B(c4932), .Z(n14798) );
XOR U24665 ( .A(c4933), .B(n14799), .Z(c4934) );
ANDN U24666 ( .B(n14800), .A(n14801), .Z(n14799) );
XOR U24667 ( .A(c4933), .B(b[4933]), .Z(n14800) );
XNOR U24668 ( .A(b[4933]), .B(n14801), .Z(c[4933]) );
XNOR U24669 ( .A(a[4933]), .B(c4933), .Z(n14801) );
XOR U24670 ( .A(c4934), .B(n14802), .Z(c4935) );
ANDN U24671 ( .B(n14803), .A(n14804), .Z(n14802) );
XOR U24672 ( .A(c4934), .B(b[4934]), .Z(n14803) );
XNOR U24673 ( .A(b[4934]), .B(n14804), .Z(c[4934]) );
XNOR U24674 ( .A(a[4934]), .B(c4934), .Z(n14804) );
XOR U24675 ( .A(c4935), .B(n14805), .Z(c4936) );
ANDN U24676 ( .B(n14806), .A(n14807), .Z(n14805) );
XOR U24677 ( .A(c4935), .B(b[4935]), .Z(n14806) );
XNOR U24678 ( .A(b[4935]), .B(n14807), .Z(c[4935]) );
XNOR U24679 ( .A(a[4935]), .B(c4935), .Z(n14807) );
XOR U24680 ( .A(c4936), .B(n14808), .Z(c4937) );
ANDN U24681 ( .B(n14809), .A(n14810), .Z(n14808) );
XOR U24682 ( .A(c4936), .B(b[4936]), .Z(n14809) );
XNOR U24683 ( .A(b[4936]), .B(n14810), .Z(c[4936]) );
XNOR U24684 ( .A(a[4936]), .B(c4936), .Z(n14810) );
XOR U24685 ( .A(c4937), .B(n14811), .Z(c4938) );
ANDN U24686 ( .B(n14812), .A(n14813), .Z(n14811) );
XOR U24687 ( .A(c4937), .B(b[4937]), .Z(n14812) );
XNOR U24688 ( .A(b[4937]), .B(n14813), .Z(c[4937]) );
XNOR U24689 ( .A(a[4937]), .B(c4937), .Z(n14813) );
XOR U24690 ( .A(c4938), .B(n14814), .Z(c4939) );
ANDN U24691 ( .B(n14815), .A(n14816), .Z(n14814) );
XOR U24692 ( .A(c4938), .B(b[4938]), .Z(n14815) );
XNOR U24693 ( .A(b[4938]), .B(n14816), .Z(c[4938]) );
XNOR U24694 ( .A(a[4938]), .B(c4938), .Z(n14816) );
XOR U24695 ( .A(c4939), .B(n14817), .Z(c4940) );
ANDN U24696 ( .B(n14818), .A(n14819), .Z(n14817) );
XOR U24697 ( .A(c4939), .B(b[4939]), .Z(n14818) );
XNOR U24698 ( .A(b[4939]), .B(n14819), .Z(c[4939]) );
XNOR U24699 ( .A(a[4939]), .B(c4939), .Z(n14819) );
XOR U24700 ( .A(c4940), .B(n14820), .Z(c4941) );
ANDN U24701 ( .B(n14821), .A(n14822), .Z(n14820) );
XOR U24702 ( .A(c4940), .B(b[4940]), .Z(n14821) );
XNOR U24703 ( .A(b[4940]), .B(n14822), .Z(c[4940]) );
XNOR U24704 ( .A(a[4940]), .B(c4940), .Z(n14822) );
XOR U24705 ( .A(c4941), .B(n14823), .Z(c4942) );
ANDN U24706 ( .B(n14824), .A(n14825), .Z(n14823) );
XOR U24707 ( .A(c4941), .B(b[4941]), .Z(n14824) );
XNOR U24708 ( .A(b[4941]), .B(n14825), .Z(c[4941]) );
XNOR U24709 ( .A(a[4941]), .B(c4941), .Z(n14825) );
XOR U24710 ( .A(c4942), .B(n14826), .Z(c4943) );
ANDN U24711 ( .B(n14827), .A(n14828), .Z(n14826) );
XOR U24712 ( .A(c4942), .B(b[4942]), .Z(n14827) );
XNOR U24713 ( .A(b[4942]), .B(n14828), .Z(c[4942]) );
XNOR U24714 ( .A(a[4942]), .B(c4942), .Z(n14828) );
XOR U24715 ( .A(c4943), .B(n14829), .Z(c4944) );
ANDN U24716 ( .B(n14830), .A(n14831), .Z(n14829) );
XOR U24717 ( .A(c4943), .B(b[4943]), .Z(n14830) );
XNOR U24718 ( .A(b[4943]), .B(n14831), .Z(c[4943]) );
XNOR U24719 ( .A(a[4943]), .B(c4943), .Z(n14831) );
XOR U24720 ( .A(c4944), .B(n14832), .Z(c4945) );
ANDN U24721 ( .B(n14833), .A(n14834), .Z(n14832) );
XOR U24722 ( .A(c4944), .B(b[4944]), .Z(n14833) );
XNOR U24723 ( .A(b[4944]), .B(n14834), .Z(c[4944]) );
XNOR U24724 ( .A(a[4944]), .B(c4944), .Z(n14834) );
XOR U24725 ( .A(c4945), .B(n14835), .Z(c4946) );
ANDN U24726 ( .B(n14836), .A(n14837), .Z(n14835) );
XOR U24727 ( .A(c4945), .B(b[4945]), .Z(n14836) );
XNOR U24728 ( .A(b[4945]), .B(n14837), .Z(c[4945]) );
XNOR U24729 ( .A(a[4945]), .B(c4945), .Z(n14837) );
XOR U24730 ( .A(c4946), .B(n14838), .Z(c4947) );
ANDN U24731 ( .B(n14839), .A(n14840), .Z(n14838) );
XOR U24732 ( .A(c4946), .B(b[4946]), .Z(n14839) );
XNOR U24733 ( .A(b[4946]), .B(n14840), .Z(c[4946]) );
XNOR U24734 ( .A(a[4946]), .B(c4946), .Z(n14840) );
XOR U24735 ( .A(c4947), .B(n14841), .Z(c4948) );
ANDN U24736 ( .B(n14842), .A(n14843), .Z(n14841) );
XOR U24737 ( .A(c4947), .B(b[4947]), .Z(n14842) );
XNOR U24738 ( .A(b[4947]), .B(n14843), .Z(c[4947]) );
XNOR U24739 ( .A(a[4947]), .B(c4947), .Z(n14843) );
XOR U24740 ( .A(c4948), .B(n14844), .Z(c4949) );
ANDN U24741 ( .B(n14845), .A(n14846), .Z(n14844) );
XOR U24742 ( .A(c4948), .B(b[4948]), .Z(n14845) );
XNOR U24743 ( .A(b[4948]), .B(n14846), .Z(c[4948]) );
XNOR U24744 ( .A(a[4948]), .B(c4948), .Z(n14846) );
XOR U24745 ( .A(c4949), .B(n14847), .Z(c4950) );
ANDN U24746 ( .B(n14848), .A(n14849), .Z(n14847) );
XOR U24747 ( .A(c4949), .B(b[4949]), .Z(n14848) );
XNOR U24748 ( .A(b[4949]), .B(n14849), .Z(c[4949]) );
XNOR U24749 ( .A(a[4949]), .B(c4949), .Z(n14849) );
XOR U24750 ( .A(c4950), .B(n14850), .Z(c4951) );
ANDN U24751 ( .B(n14851), .A(n14852), .Z(n14850) );
XOR U24752 ( .A(c4950), .B(b[4950]), .Z(n14851) );
XNOR U24753 ( .A(b[4950]), .B(n14852), .Z(c[4950]) );
XNOR U24754 ( .A(a[4950]), .B(c4950), .Z(n14852) );
XOR U24755 ( .A(c4951), .B(n14853), .Z(c4952) );
ANDN U24756 ( .B(n14854), .A(n14855), .Z(n14853) );
XOR U24757 ( .A(c4951), .B(b[4951]), .Z(n14854) );
XNOR U24758 ( .A(b[4951]), .B(n14855), .Z(c[4951]) );
XNOR U24759 ( .A(a[4951]), .B(c4951), .Z(n14855) );
XOR U24760 ( .A(c4952), .B(n14856), .Z(c4953) );
ANDN U24761 ( .B(n14857), .A(n14858), .Z(n14856) );
XOR U24762 ( .A(c4952), .B(b[4952]), .Z(n14857) );
XNOR U24763 ( .A(b[4952]), .B(n14858), .Z(c[4952]) );
XNOR U24764 ( .A(a[4952]), .B(c4952), .Z(n14858) );
XOR U24765 ( .A(c4953), .B(n14859), .Z(c4954) );
ANDN U24766 ( .B(n14860), .A(n14861), .Z(n14859) );
XOR U24767 ( .A(c4953), .B(b[4953]), .Z(n14860) );
XNOR U24768 ( .A(b[4953]), .B(n14861), .Z(c[4953]) );
XNOR U24769 ( .A(a[4953]), .B(c4953), .Z(n14861) );
XOR U24770 ( .A(c4954), .B(n14862), .Z(c4955) );
ANDN U24771 ( .B(n14863), .A(n14864), .Z(n14862) );
XOR U24772 ( .A(c4954), .B(b[4954]), .Z(n14863) );
XNOR U24773 ( .A(b[4954]), .B(n14864), .Z(c[4954]) );
XNOR U24774 ( .A(a[4954]), .B(c4954), .Z(n14864) );
XOR U24775 ( .A(c4955), .B(n14865), .Z(c4956) );
ANDN U24776 ( .B(n14866), .A(n14867), .Z(n14865) );
XOR U24777 ( .A(c4955), .B(b[4955]), .Z(n14866) );
XNOR U24778 ( .A(b[4955]), .B(n14867), .Z(c[4955]) );
XNOR U24779 ( .A(a[4955]), .B(c4955), .Z(n14867) );
XOR U24780 ( .A(c4956), .B(n14868), .Z(c4957) );
ANDN U24781 ( .B(n14869), .A(n14870), .Z(n14868) );
XOR U24782 ( .A(c4956), .B(b[4956]), .Z(n14869) );
XNOR U24783 ( .A(b[4956]), .B(n14870), .Z(c[4956]) );
XNOR U24784 ( .A(a[4956]), .B(c4956), .Z(n14870) );
XOR U24785 ( .A(c4957), .B(n14871), .Z(c4958) );
ANDN U24786 ( .B(n14872), .A(n14873), .Z(n14871) );
XOR U24787 ( .A(c4957), .B(b[4957]), .Z(n14872) );
XNOR U24788 ( .A(b[4957]), .B(n14873), .Z(c[4957]) );
XNOR U24789 ( .A(a[4957]), .B(c4957), .Z(n14873) );
XOR U24790 ( .A(c4958), .B(n14874), .Z(c4959) );
ANDN U24791 ( .B(n14875), .A(n14876), .Z(n14874) );
XOR U24792 ( .A(c4958), .B(b[4958]), .Z(n14875) );
XNOR U24793 ( .A(b[4958]), .B(n14876), .Z(c[4958]) );
XNOR U24794 ( .A(a[4958]), .B(c4958), .Z(n14876) );
XOR U24795 ( .A(c4959), .B(n14877), .Z(c4960) );
ANDN U24796 ( .B(n14878), .A(n14879), .Z(n14877) );
XOR U24797 ( .A(c4959), .B(b[4959]), .Z(n14878) );
XNOR U24798 ( .A(b[4959]), .B(n14879), .Z(c[4959]) );
XNOR U24799 ( .A(a[4959]), .B(c4959), .Z(n14879) );
XOR U24800 ( .A(c4960), .B(n14880), .Z(c4961) );
ANDN U24801 ( .B(n14881), .A(n14882), .Z(n14880) );
XOR U24802 ( .A(c4960), .B(b[4960]), .Z(n14881) );
XNOR U24803 ( .A(b[4960]), .B(n14882), .Z(c[4960]) );
XNOR U24804 ( .A(a[4960]), .B(c4960), .Z(n14882) );
XOR U24805 ( .A(c4961), .B(n14883), .Z(c4962) );
ANDN U24806 ( .B(n14884), .A(n14885), .Z(n14883) );
XOR U24807 ( .A(c4961), .B(b[4961]), .Z(n14884) );
XNOR U24808 ( .A(b[4961]), .B(n14885), .Z(c[4961]) );
XNOR U24809 ( .A(a[4961]), .B(c4961), .Z(n14885) );
XOR U24810 ( .A(c4962), .B(n14886), .Z(c4963) );
ANDN U24811 ( .B(n14887), .A(n14888), .Z(n14886) );
XOR U24812 ( .A(c4962), .B(b[4962]), .Z(n14887) );
XNOR U24813 ( .A(b[4962]), .B(n14888), .Z(c[4962]) );
XNOR U24814 ( .A(a[4962]), .B(c4962), .Z(n14888) );
XOR U24815 ( .A(c4963), .B(n14889), .Z(c4964) );
ANDN U24816 ( .B(n14890), .A(n14891), .Z(n14889) );
XOR U24817 ( .A(c4963), .B(b[4963]), .Z(n14890) );
XNOR U24818 ( .A(b[4963]), .B(n14891), .Z(c[4963]) );
XNOR U24819 ( .A(a[4963]), .B(c4963), .Z(n14891) );
XOR U24820 ( .A(c4964), .B(n14892), .Z(c4965) );
ANDN U24821 ( .B(n14893), .A(n14894), .Z(n14892) );
XOR U24822 ( .A(c4964), .B(b[4964]), .Z(n14893) );
XNOR U24823 ( .A(b[4964]), .B(n14894), .Z(c[4964]) );
XNOR U24824 ( .A(a[4964]), .B(c4964), .Z(n14894) );
XOR U24825 ( .A(c4965), .B(n14895), .Z(c4966) );
ANDN U24826 ( .B(n14896), .A(n14897), .Z(n14895) );
XOR U24827 ( .A(c4965), .B(b[4965]), .Z(n14896) );
XNOR U24828 ( .A(b[4965]), .B(n14897), .Z(c[4965]) );
XNOR U24829 ( .A(a[4965]), .B(c4965), .Z(n14897) );
XOR U24830 ( .A(c4966), .B(n14898), .Z(c4967) );
ANDN U24831 ( .B(n14899), .A(n14900), .Z(n14898) );
XOR U24832 ( .A(c4966), .B(b[4966]), .Z(n14899) );
XNOR U24833 ( .A(b[4966]), .B(n14900), .Z(c[4966]) );
XNOR U24834 ( .A(a[4966]), .B(c4966), .Z(n14900) );
XOR U24835 ( .A(c4967), .B(n14901), .Z(c4968) );
ANDN U24836 ( .B(n14902), .A(n14903), .Z(n14901) );
XOR U24837 ( .A(c4967), .B(b[4967]), .Z(n14902) );
XNOR U24838 ( .A(b[4967]), .B(n14903), .Z(c[4967]) );
XNOR U24839 ( .A(a[4967]), .B(c4967), .Z(n14903) );
XOR U24840 ( .A(c4968), .B(n14904), .Z(c4969) );
ANDN U24841 ( .B(n14905), .A(n14906), .Z(n14904) );
XOR U24842 ( .A(c4968), .B(b[4968]), .Z(n14905) );
XNOR U24843 ( .A(b[4968]), .B(n14906), .Z(c[4968]) );
XNOR U24844 ( .A(a[4968]), .B(c4968), .Z(n14906) );
XOR U24845 ( .A(c4969), .B(n14907), .Z(c4970) );
ANDN U24846 ( .B(n14908), .A(n14909), .Z(n14907) );
XOR U24847 ( .A(c4969), .B(b[4969]), .Z(n14908) );
XNOR U24848 ( .A(b[4969]), .B(n14909), .Z(c[4969]) );
XNOR U24849 ( .A(a[4969]), .B(c4969), .Z(n14909) );
XOR U24850 ( .A(c4970), .B(n14910), .Z(c4971) );
ANDN U24851 ( .B(n14911), .A(n14912), .Z(n14910) );
XOR U24852 ( .A(c4970), .B(b[4970]), .Z(n14911) );
XNOR U24853 ( .A(b[4970]), .B(n14912), .Z(c[4970]) );
XNOR U24854 ( .A(a[4970]), .B(c4970), .Z(n14912) );
XOR U24855 ( .A(c4971), .B(n14913), .Z(c4972) );
ANDN U24856 ( .B(n14914), .A(n14915), .Z(n14913) );
XOR U24857 ( .A(c4971), .B(b[4971]), .Z(n14914) );
XNOR U24858 ( .A(b[4971]), .B(n14915), .Z(c[4971]) );
XNOR U24859 ( .A(a[4971]), .B(c4971), .Z(n14915) );
XOR U24860 ( .A(c4972), .B(n14916), .Z(c4973) );
ANDN U24861 ( .B(n14917), .A(n14918), .Z(n14916) );
XOR U24862 ( .A(c4972), .B(b[4972]), .Z(n14917) );
XNOR U24863 ( .A(b[4972]), .B(n14918), .Z(c[4972]) );
XNOR U24864 ( .A(a[4972]), .B(c4972), .Z(n14918) );
XOR U24865 ( .A(c4973), .B(n14919), .Z(c4974) );
ANDN U24866 ( .B(n14920), .A(n14921), .Z(n14919) );
XOR U24867 ( .A(c4973), .B(b[4973]), .Z(n14920) );
XNOR U24868 ( .A(b[4973]), .B(n14921), .Z(c[4973]) );
XNOR U24869 ( .A(a[4973]), .B(c4973), .Z(n14921) );
XOR U24870 ( .A(c4974), .B(n14922), .Z(c4975) );
ANDN U24871 ( .B(n14923), .A(n14924), .Z(n14922) );
XOR U24872 ( .A(c4974), .B(b[4974]), .Z(n14923) );
XNOR U24873 ( .A(b[4974]), .B(n14924), .Z(c[4974]) );
XNOR U24874 ( .A(a[4974]), .B(c4974), .Z(n14924) );
XOR U24875 ( .A(c4975), .B(n14925), .Z(c4976) );
ANDN U24876 ( .B(n14926), .A(n14927), .Z(n14925) );
XOR U24877 ( .A(c4975), .B(b[4975]), .Z(n14926) );
XNOR U24878 ( .A(b[4975]), .B(n14927), .Z(c[4975]) );
XNOR U24879 ( .A(a[4975]), .B(c4975), .Z(n14927) );
XOR U24880 ( .A(c4976), .B(n14928), .Z(c4977) );
ANDN U24881 ( .B(n14929), .A(n14930), .Z(n14928) );
XOR U24882 ( .A(c4976), .B(b[4976]), .Z(n14929) );
XNOR U24883 ( .A(b[4976]), .B(n14930), .Z(c[4976]) );
XNOR U24884 ( .A(a[4976]), .B(c4976), .Z(n14930) );
XOR U24885 ( .A(c4977), .B(n14931), .Z(c4978) );
ANDN U24886 ( .B(n14932), .A(n14933), .Z(n14931) );
XOR U24887 ( .A(c4977), .B(b[4977]), .Z(n14932) );
XNOR U24888 ( .A(b[4977]), .B(n14933), .Z(c[4977]) );
XNOR U24889 ( .A(a[4977]), .B(c4977), .Z(n14933) );
XOR U24890 ( .A(c4978), .B(n14934), .Z(c4979) );
ANDN U24891 ( .B(n14935), .A(n14936), .Z(n14934) );
XOR U24892 ( .A(c4978), .B(b[4978]), .Z(n14935) );
XNOR U24893 ( .A(b[4978]), .B(n14936), .Z(c[4978]) );
XNOR U24894 ( .A(a[4978]), .B(c4978), .Z(n14936) );
XOR U24895 ( .A(c4979), .B(n14937), .Z(c4980) );
ANDN U24896 ( .B(n14938), .A(n14939), .Z(n14937) );
XOR U24897 ( .A(c4979), .B(b[4979]), .Z(n14938) );
XNOR U24898 ( .A(b[4979]), .B(n14939), .Z(c[4979]) );
XNOR U24899 ( .A(a[4979]), .B(c4979), .Z(n14939) );
XOR U24900 ( .A(c4980), .B(n14940), .Z(c4981) );
ANDN U24901 ( .B(n14941), .A(n14942), .Z(n14940) );
XOR U24902 ( .A(c4980), .B(b[4980]), .Z(n14941) );
XNOR U24903 ( .A(b[4980]), .B(n14942), .Z(c[4980]) );
XNOR U24904 ( .A(a[4980]), .B(c4980), .Z(n14942) );
XOR U24905 ( .A(c4981), .B(n14943), .Z(c4982) );
ANDN U24906 ( .B(n14944), .A(n14945), .Z(n14943) );
XOR U24907 ( .A(c4981), .B(b[4981]), .Z(n14944) );
XNOR U24908 ( .A(b[4981]), .B(n14945), .Z(c[4981]) );
XNOR U24909 ( .A(a[4981]), .B(c4981), .Z(n14945) );
XOR U24910 ( .A(c4982), .B(n14946), .Z(c4983) );
ANDN U24911 ( .B(n14947), .A(n14948), .Z(n14946) );
XOR U24912 ( .A(c4982), .B(b[4982]), .Z(n14947) );
XNOR U24913 ( .A(b[4982]), .B(n14948), .Z(c[4982]) );
XNOR U24914 ( .A(a[4982]), .B(c4982), .Z(n14948) );
XOR U24915 ( .A(c4983), .B(n14949), .Z(c4984) );
ANDN U24916 ( .B(n14950), .A(n14951), .Z(n14949) );
XOR U24917 ( .A(c4983), .B(b[4983]), .Z(n14950) );
XNOR U24918 ( .A(b[4983]), .B(n14951), .Z(c[4983]) );
XNOR U24919 ( .A(a[4983]), .B(c4983), .Z(n14951) );
XOR U24920 ( .A(c4984), .B(n14952), .Z(c4985) );
ANDN U24921 ( .B(n14953), .A(n14954), .Z(n14952) );
XOR U24922 ( .A(c4984), .B(b[4984]), .Z(n14953) );
XNOR U24923 ( .A(b[4984]), .B(n14954), .Z(c[4984]) );
XNOR U24924 ( .A(a[4984]), .B(c4984), .Z(n14954) );
XOR U24925 ( .A(c4985), .B(n14955), .Z(c4986) );
ANDN U24926 ( .B(n14956), .A(n14957), .Z(n14955) );
XOR U24927 ( .A(c4985), .B(b[4985]), .Z(n14956) );
XNOR U24928 ( .A(b[4985]), .B(n14957), .Z(c[4985]) );
XNOR U24929 ( .A(a[4985]), .B(c4985), .Z(n14957) );
XOR U24930 ( .A(c4986), .B(n14958), .Z(c4987) );
ANDN U24931 ( .B(n14959), .A(n14960), .Z(n14958) );
XOR U24932 ( .A(c4986), .B(b[4986]), .Z(n14959) );
XNOR U24933 ( .A(b[4986]), .B(n14960), .Z(c[4986]) );
XNOR U24934 ( .A(a[4986]), .B(c4986), .Z(n14960) );
XOR U24935 ( .A(c4987), .B(n14961), .Z(c4988) );
ANDN U24936 ( .B(n14962), .A(n14963), .Z(n14961) );
XOR U24937 ( .A(c4987), .B(b[4987]), .Z(n14962) );
XNOR U24938 ( .A(b[4987]), .B(n14963), .Z(c[4987]) );
XNOR U24939 ( .A(a[4987]), .B(c4987), .Z(n14963) );
XOR U24940 ( .A(c4988), .B(n14964), .Z(c4989) );
ANDN U24941 ( .B(n14965), .A(n14966), .Z(n14964) );
XOR U24942 ( .A(c4988), .B(b[4988]), .Z(n14965) );
XNOR U24943 ( .A(b[4988]), .B(n14966), .Z(c[4988]) );
XNOR U24944 ( .A(a[4988]), .B(c4988), .Z(n14966) );
XOR U24945 ( .A(c4989), .B(n14967), .Z(c4990) );
ANDN U24946 ( .B(n14968), .A(n14969), .Z(n14967) );
XOR U24947 ( .A(c4989), .B(b[4989]), .Z(n14968) );
XNOR U24948 ( .A(b[4989]), .B(n14969), .Z(c[4989]) );
XNOR U24949 ( .A(a[4989]), .B(c4989), .Z(n14969) );
XOR U24950 ( .A(c4990), .B(n14970), .Z(c4991) );
ANDN U24951 ( .B(n14971), .A(n14972), .Z(n14970) );
XOR U24952 ( .A(c4990), .B(b[4990]), .Z(n14971) );
XNOR U24953 ( .A(b[4990]), .B(n14972), .Z(c[4990]) );
XNOR U24954 ( .A(a[4990]), .B(c4990), .Z(n14972) );
XOR U24955 ( .A(c4991), .B(n14973), .Z(c4992) );
ANDN U24956 ( .B(n14974), .A(n14975), .Z(n14973) );
XOR U24957 ( .A(c4991), .B(b[4991]), .Z(n14974) );
XNOR U24958 ( .A(b[4991]), .B(n14975), .Z(c[4991]) );
XNOR U24959 ( .A(a[4991]), .B(c4991), .Z(n14975) );
XOR U24960 ( .A(c4992), .B(n14976), .Z(c4993) );
ANDN U24961 ( .B(n14977), .A(n14978), .Z(n14976) );
XOR U24962 ( .A(c4992), .B(b[4992]), .Z(n14977) );
XNOR U24963 ( .A(b[4992]), .B(n14978), .Z(c[4992]) );
XNOR U24964 ( .A(a[4992]), .B(c4992), .Z(n14978) );
XOR U24965 ( .A(c4993), .B(n14979), .Z(c4994) );
ANDN U24966 ( .B(n14980), .A(n14981), .Z(n14979) );
XOR U24967 ( .A(c4993), .B(b[4993]), .Z(n14980) );
XNOR U24968 ( .A(b[4993]), .B(n14981), .Z(c[4993]) );
XNOR U24969 ( .A(a[4993]), .B(c4993), .Z(n14981) );
XOR U24970 ( .A(c4994), .B(n14982), .Z(c4995) );
ANDN U24971 ( .B(n14983), .A(n14984), .Z(n14982) );
XOR U24972 ( .A(c4994), .B(b[4994]), .Z(n14983) );
XNOR U24973 ( .A(b[4994]), .B(n14984), .Z(c[4994]) );
XNOR U24974 ( .A(a[4994]), .B(c4994), .Z(n14984) );
XOR U24975 ( .A(c4995), .B(n14985), .Z(c4996) );
ANDN U24976 ( .B(n14986), .A(n14987), .Z(n14985) );
XOR U24977 ( .A(c4995), .B(b[4995]), .Z(n14986) );
XNOR U24978 ( .A(b[4995]), .B(n14987), .Z(c[4995]) );
XNOR U24979 ( .A(a[4995]), .B(c4995), .Z(n14987) );
XOR U24980 ( .A(c4996), .B(n14988), .Z(c4997) );
ANDN U24981 ( .B(n14989), .A(n14990), .Z(n14988) );
XOR U24982 ( .A(c4996), .B(b[4996]), .Z(n14989) );
XNOR U24983 ( .A(b[4996]), .B(n14990), .Z(c[4996]) );
XNOR U24984 ( .A(a[4996]), .B(c4996), .Z(n14990) );
XOR U24985 ( .A(c4997), .B(n14991), .Z(c4998) );
ANDN U24986 ( .B(n14992), .A(n14993), .Z(n14991) );
XOR U24987 ( .A(c4997), .B(b[4997]), .Z(n14992) );
XNOR U24988 ( .A(b[4997]), .B(n14993), .Z(c[4997]) );
XNOR U24989 ( .A(a[4997]), .B(c4997), .Z(n14993) );
XOR U24990 ( .A(c4998), .B(n14994), .Z(c4999) );
ANDN U24991 ( .B(n14995), .A(n14996), .Z(n14994) );
XOR U24992 ( .A(c4998), .B(b[4998]), .Z(n14995) );
XNOR U24993 ( .A(b[4998]), .B(n14996), .Z(c[4998]) );
XNOR U24994 ( .A(a[4998]), .B(c4998), .Z(n14996) );
XOR U24995 ( .A(c4999), .B(n14997), .Z(c5000) );
ANDN U24996 ( .B(n14998), .A(n14999), .Z(n14997) );
XOR U24997 ( .A(c4999), .B(b[4999]), .Z(n14998) );
XNOR U24998 ( .A(b[4999]), .B(n14999), .Z(c[4999]) );
XNOR U24999 ( .A(a[4999]), .B(c4999), .Z(n14999) );
XOR U25000 ( .A(c5000), .B(n15000), .Z(c5001) );
ANDN U25001 ( .B(n15001), .A(n15002), .Z(n15000) );
XOR U25002 ( .A(c5000), .B(b[5000]), .Z(n15001) );
XNOR U25003 ( .A(b[5000]), .B(n15002), .Z(c[5000]) );
XNOR U25004 ( .A(a[5000]), .B(c5000), .Z(n15002) );
XOR U25005 ( .A(c5001), .B(n15003), .Z(c5002) );
ANDN U25006 ( .B(n15004), .A(n15005), .Z(n15003) );
XOR U25007 ( .A(c5001), .B(b[5001]), .Z(n15004) );
XNOR U25008 ( .A(b[5001]), .B(n15005), .Z(c[5001]) );
XNOR U25009 ( .A(a[5001]), .B(c5001), .Z(n15005) );
XOR U25010 ( .A(c5002), .B(n15006), .Z(c5003) );
ANDN U25011 ( .B(n15007), .A(n15008), .Z(n15006) );
XOR U25012 ( .A(c5002), .B(b[5002]), .Z(n15007) );
XNOR U25013 ( .A(b[5002]), .B(n15008), .Z(c[5002]) );
XNOR U25014 ( .A(a[5002]), .B(c5002), .Z(n15008) );
XOR U25015 ( .A(c5003), .B(n15009), .Z(c5004) );
ANDN U25016 ( .B(n15010), .A(n15011), .Z(n15009) );
XOR U25017 ( .A(c5003), .B(b[5003]), .Z(n15010) );
XNOR U25018 ( .A(b[5003]), .B(n15011), .Z(c[5003]) );
XNOR U25019 ( .A(a[5003]), .B(c5003), .Z(n15011) );
XOR U25020 ( .A(c5004), .B(n15012), .Z(c5005) );
ANDN U25021 ( .B(n15013), .A(n15014), .Z(n15012) );
XOR U25022 ( .A(c5004), .B(b[5004]), .Z(n15013) );
XNOR U25023 ( .A(b[5004]), .B(n15014), .Z(c[5004]) );
XNOR U25024 ( .A(a[5004]), .B(c5004), .Z(n15014) );
XOR U25025 ( .A(c5005), .B(n15015), .Z(c5006) );
ANDN U25026 ( .B(n15016), .A(n15017), .Z(n15015) );
XOR U25027 ( .A(c5005), .B(b[5005]), .Z(n15016) );
XNOR U25028 ( .A(b[5005]), .B(n15017), .Z(c[5005]) );
XNOR U25029 ( .A(a[5005]), .B(c5005), .Z(n15017) );
XOR U25030 ( .A(c5006), .B(n15018), .Z(c5007) );
ANDN U25031 ( .B(n15019), .A(n15020), .Z(n15018) );
XOR U25032 ( .A(c5006), .B(b[5006]), .Z(n15019) );
XNOR U25033 ( .A(b[5006]), .B(n15020), .Z(c[5006]) );
XNOR U25034 ( .A(a[5006]), .B(c5006), .Z(n15020) );
XOR U25035 ( .A(c5007), .B(n15021), .Z(c5008) );
ANDN U25036 ( .B(n15022), .A(n15023), .Z(n15021) );
XOR U25037 ( .A(c5007), .B(b[5007]), .Z(n15022) );
XNOR U25038 ( .A(b[5007]), .B(n15023), .Z(c[5007]) );
XNOR U25039 ( .A(a[5007]), .B(c5007), .Z(n15023) );
XOR U25040 ( .A(c5008), .B(n15024), .Z(c5009) );
ANDN U25041 ( .B(n15025), .A(n15026), .Z(n15024) );
XOR U25042 ( .A(c5008), .B(b[5008]), .Z(n15025) );
XNOR U25043 ( .A(b[5008]), .B(n15026), .Z(c[5008]) );
XNOR U25044 ( .A(a[5008]), .B(c5008), .Z(n15026) );
XOR U25045 ( .A(c5009), .B(n15027), .Z(c5010) );
ANDN U25046 ( .B(n15028), .A(n15029), .Z(n15027) );
XOR U25047 ( .A(c5009), .B(b[5009]), .Z(n15028) );
XNOR U25048 ( .A(b[5009]), .B(n15029), .Z(c[5009]) );
XNOR U25049 ( .A(a[5009]), .B(c5009), .Z(n15029) );
XOR U25050 ( .A(c5010), .B(n15030), .Z(c5011) );
ANDN U25051 ( .B(n15031), .A(n15032), .Z(n15030) );
XOR U25052 ( .A(c5010), .B(b[5010]), .Z(n15031) );
XNOR U25053 ( .A(b[5010]), .B(n15032), .Z(c[5010]) );
XNOR U25054 ( .A(a[5010]), .B(c5010), .Z(n15032) );
XOR U25055 ( .A(c5011), .B(n15033), .Z(c5012) );
ANDN U25056 ( .B(n15034), .A(n15035), .Z(n15033) );
XOR U25057 ( .A(c5011), .B(b[5011]), .Z(n15034) );
XNOR U25058 ( .A(b[5011]), .B(n15035), .Z(c[5011]) );
XNOR U25059 ( .A(a[5011]), .B(c5011), .Z(n15035) );
XOR U25060 ( .A(c5012), .B(n15036), .Z(c5013) );
ANDN U25061 ( .B(n15037), .A(n15038), .Z(n15036) );
XOR U25062 ( .A(c5012), .B(b[5012]), .Z(n15037) );
XNOR U25063 ( .A(b[5012]), .B(n15038), .Z(c[5012]) );
XNOR U25064 ( .A(a[5012]), .B(c5012), .Z(n15038) );
XOR U25065 ( .A(c5013), .B(n15039), .Z(c5014) );
ANDN U25066 ( .B(n15040), .A(n15041), .Z(n15039) );
XOR U25067 ( .A(c5013), .B(b[5013]), .Z(n15040) );
XNOR U25068 ( .A(b[5013]), .B(n15041), .Z(c[5013]) );
XNOR U25069 ( .A(a[5013]), .B(c5013), .Z(n15041) );
XOR U25070 ( .A(c5014), .B(n15042), .Z(c5015) );
ANDN U25071 ( .B(n15043), .A(n15044), .Z(n15042) );
XOR U25072 ( .A(c5014), .B(b[5014]), .Z(n15043) );
XNOR U25073 ( .A(b[5014]), .B(n15044), .Z(c[5014]) );
XNOR U25074 ( .A(a[5014]), .B(c5014), .Z(n15044) );
XOR U25075 ( .A(c5015), .B(n15045), .Z(c5016) );
ANDN U25076 ( .B(n15046), .A(n15047), .Z(n15045) );
XOR U25077 ( .A(c5015), .B(b[5015]), .Z(n15046) );
XNOR U25078 ( .A(b[5015]), .B(n15047), .Z(c[5015]) );
XNOR U25079 ( .A(a[5015]), .B(c5015), .Z(n15047) );
XOR U25080 ( .A(c5016), .B(n15048), .Z(c5017) );
ANDN U25081 ( .B(n15049), .A(n15050), .Z(n15048) );
XOR U25082 ( .A(c5016), .B(b[5016]), .Z(n15049) );
XNOR U25083 ( .A(b[5016]), .B(n15050), .Z(c[5016]) );
XNOR U25084 ( .A(a[5016]), .B(c5016), .Z(n15050) );
XOR U25085 ( .A(c5017), .B(n15051), .Z(c5018) );
ANDN U25086 ( .B(n15052), .A(n15053), .Z(n15051) );
XOR U25087 ( .A(c5017), .B(b[5017]), .Z(n15052) );
XNOR U25088 ( .A(b[5017]), .B(n15053), .Z(c[5017]) );
XNOR U25089 ( .A(a[5017]), .B(c5017), .Z(n15053) );
XOR U25090 ( .A(c5018), .B(n15054), .Z(c5019) );
ANDN U25091 ( .B(n15055), .A(n15056), .Z(n15054) );
XOR U25092 ( .A(c5018), .B(b[5018]), .Z(n15055) );
XNOR U25093 ( .A(b[5018]), .B(n15056), .Z(c[5018]) );
XNOR U25094 ( .A(a[5018]), .B(c5018), .Z(n15056) );
XOR U25095 ( .A(c5019), .B(n15057), .Z(c5020) );
ANDN U25096 ( .B(n15058), .A(n15059), .Z(n15057) );
XOR U25097 ( .A(c5019), .B(b[5019]), .Z(n15058) );
XNOR U25098 ( .A(b[5019]), .B(n15059), .Z(c[5019]) );
XNOR U25099 ( .A(a[5019]), .B(c5019), .Z(n15059) );
XOR U25100 ( .A(c5020), .B(n15060), .Z(c5021) );
ANDN U25101 ( .B(n15061), .A(n15062), .Z(n15060) );
XOR U25102 ( .A(c5020), .B(b[5020]), .Z(n15061) );
XNOR U25103 ( .A(b[5020]), .B(n15062), .Z(c[5020]) );
XNOR U25104 ( .A(a[5020]), .B(c5020), .Z(n15062) );
XOR U25105 ( .A(c5021), .B(n15063), .Z(c5022) );
ANDN U25106 ( .B(n15064), .A(n15065), .Z(n15063) );
XOR U25107 ( .A(c5021), .B(b[5021]), .Z(n15064) );
XNOR U25108 ( .A(b[5021]), .B(n15065), .Z(c[5021]) );
XNOR U25109 ( .A(a[5021]), .B(c5021), .Z(n15065) );
XOR U25110 ( .A(c5022), .B(n15066), .Z(c5023) );
ANDN U25111 ( .B(n15067), .A(n15068), .Z(n15066) );
XOR U25112 ( .A(c5022), .B(b[5022]), .Z(n15067) );
XNOR U25113 ( .A(b[5022]), .B(n15068), .Z(c[5022]) );
XNOR U25114 ( .A(a[5022]), .B(c5022), .Z(n15068) );
XOR U25115 ( .A(c5023), .B(n15069), .Z(c5024) );
ANDN U25116 ( .B(n15070), .A(n15071), .Z(n15069) );
XOR U25117 ( .A(c5023), .B(b[5023]), .Z(n15070) );
XNOR U25118 ( .A(b[5023]), .B(n15071), .Z(c[5023]) );
XNOR U25119 ( .A(a[5023]), .B(c5023), .Z(n15071) );
XOR U25120 ( .A(c5024), .B(n15072), .Z(c5025) );
ANDN U25121 ( .B(n15073), .A(n15074), .Z(n15072) );
XOR U25122 ( .A(c5024), .B(b[5024]), .Z(n15073) );
XNOR U25123 ( .A(b[5024]), .B(n15074), .Z(c[5024]) );
XNOR U25124 ( .A(a[5024]), .B(c5024), .Z(n15074) );
XOR U25125 ( .A(c5025), .B(n15075), .Z(c5026) );
ANDN U25126 ( .B(n15076), .A(n15077), .Z(n15075) );
XOR U25127 ( .A(c5025), .B(b[5025]), .Z(n15076) );
XNOR U25128 ( .A(b[5025]), .B(n15077), .Z(c[5025]) );
XNOR U25129 ( .A(a[5025]), .B(c5025), .Z(n15077) );
XOR U25130 ( .A(c5026), .B(n15078), .Z(c5027) );
ANDN U25131 ( .B(n15079), .A(n15080), .Z(n15078) );
XOR U25132 ( .A(c5026), .B(b[5026]), .Z(n15079) );
XNOR U25133 ( .A(b[5026]), .B(n15080), .Z(c[5026]) );
XNOR U25134 ( .A(a[5026]), .B(c5026), .Z(n15080) );
XOR U25135 ( .A(c5027), .B(n15081), .Z(c5028) );
ANDN U25136 ( .B(n15082), .A(n15083), .Z(n15081) );
XOR U25137 ( .A(c5027), .B(b[5027]), .Z(n15082) );
XNOR U25138 ( .A(b[5027]), .B(n15083), .Z(c[5027]) );
XNOR U25139 ( .A(a[5027]), .B(c5027), .Z(n15083) );
XOR U25140 ( .A(c5028), .B(n15084), .Z(c5029) );
ANDN U25141 ( .B(n15085), .A(n15086), .Z(n15084) );
XOR U25142 ( .A(c5028), .B(b[5028]), .Z(n15085) );
XNOR U25143 ( .A(b[5028]), .B(n15086), .Z(c[5028]) );
XNOR U25144 ( .A(a[5028]), .B(c5028), .Z(n15086) );
XOR U25145 ( .A(c5029), .B(n15087), .Z(c5030) );
ANDN U25146 ( .B(n15088), .A(n15089), .Z(n15087) );
XOR U25147 ( .A(c5029), .B(b[5029]), .Z(n15088) );
XNOR U25148 ( .A(b[5029]), .B(n15089), .Z(c[5029]) );
XNOR U25149 ( .A(a[5029]), .B(c5029), .Z(n15089) );
XOR U25150 ( .A(c5030), .B(n15090), .Z(c5031) );
ANDN U25151 ( .B(n15091), .A(n15092), .Z(n15090) );
XOR U25152 ( .A(c5030), .B(b[5030]), .Z(n15091) );
XNOR U25153 ( .A(b[5030]), .B(n15092), .Z(c[5030]) );
XNOR U25154 ( .A(a[5030]), .B(c5030), .Z(n15092) );
XOR U25155 ( .A(c5031), .B(n15093), .Z(c5032) );
ANDN U25156 ( .B(n15094), .A(n15095), .Z(n15093) );
XOR U25157 ( .A(c5031), .B(b[5031]), .Z(n15094) );
XNOR U25158 ( .A(b[5031]), .B(n15095), .Z(c[5031]) );
XNOR U25159 ( .A(a[5031]), .B(c5031), .Z(n15095) );
XOR U25160 ( .A(c5032), .B(n15096), .Z(c5033) );
ANDN U25161 ( .B(n15097), .A(n15098), .Z(n15096) );
XOR U25162 ( .A(c5032), .B(b[5032]), .Z(n15097) );
XNOR U25163 ( .A(b[5032]), .B(n15098), .Z(c[5032]) );
XNOR U25164 ( .A(a[5032]), .B(c5032), .Z(n15098) );
XOR U25165 ( .A(c5033), .B(n15099), .Z(c5034) );
ANDN U25166 ( .B(n15100), .A(n15101), .Z(n15099) );
XOR U25167 ( .A(c5033), .B(b[5033]), .Z(n15100) );
XNOR U25168 ( .A(b[5033]), .B(n15101), .Z(c[5033]) );
XNOR U25169 ( .A(a[5033]), .B(c5033), .Z(n15101) );
XOR U25170 ( .A(c5034), .B(n15102), .Z(c5035) );
ANDN U25171 ( .B(n15103), .A(n15104), .Z(n15102) );
XOR U25172 ( .A(c5034), .B(b[5034]), .Z(n15103) );
XNOR U25173 ( .A(b[5034]), .B(n15104), .Z(c[5034]) );
XNOR U25174 ( .A(a[5034]), .B(c5034), .Z(n15104) );
XOR U25175 ( .A(c5035), .B(n15105), .Z(c5036) );
ANDN U25176 ( .B(n15106), .A(n15107), .Z(n15105) );
XOR U25177 ( .A(c5035), .B(b[5035]), .Z(n15106) );
XNOR U25178 ( .A(b[5035]), .B(n15107), .Z(c[5035]) );
XNOR U25179 ( .A(a[5035]), .B(c5035), .Z(n15107) );
XOR U25180 ( .A(c5036), .B(n15108), .Z(c5037) );
ANDN U25181 ( .B(n15109), .A(n15110), .Z(n15108) );
XOR U25182 ( .A(c5036), .B(b[5036]), .Z(n15109) );
XNOR U25183 ( .A(b[5036]), .B(n15110), .Z(c[5036]) );
XNOR U25184 ( .A(a[5036]), .B(c5036), .Z(n15110) );
XOR U25185 ( .A(c5037), .B(n15111), .Z(c5038) );
ANDN U25186 ( .B(n15112), .A(n15113), .Z(n15111) );
XOR U25187 ( .A(c5037), .B(b[5037]), .Z(n15112) );
XNOR U25188 ( .A(b[5037]), .B(n15113), .Z(c[5037]) );
XNOR U25189 ( .A(a[5037]), .B(c5037), .Z(n15113) );
XOR U25190 ( .A(c5038), .B(n15114), .Z(c5039) );
ANDN U25191 ( .B(n15115), .A(n15116), .Z(n15114) );
XOR U25192 ( .A(c5038), .B(b[5038]), .Z(n15115) );
XNOR U25193 ( .A(b[5038]), .B(n15116), .Z(c[5038]) );
XNOR U25194 ( .A(a[5038]), .B(c5038), .Z(n15116) );
XOR U25195 ( .A(c5039), .B(n15117), .Z(c5040) );
ANDN U25196 ( .B(n15118), .A(n15119), .Z(n15117) );
XOR U25197 ( .A(c5039), .B(b[5039]), .Z(n15118) );
XNOR U25198 ( .A(b[5039]), .B(n15119), .Z(c[5039]) );
XNOR U25199 ( .A(a[5039]), .B(c5039), .Z(n15119) );
XOR U25200 ( .A(c5040), .B(n15120), .Z(c5041) );
ANDN U25201 ( .B(n15121), .A(n15122), .Z(n15120) );
XOR U25202 ( .A(c5040), .B(b[5040]), .Z(n15121) );
XNOR U25203 ( .A(b[5040]), .B(n15122), .Z(c[5040]) );
XNOR U25204 ( .A(a[5040]), .B(c5040), .Z(n15122) );
XOR U25205 ( .A(c5041), .B(n15123), .Z(c5042) );
ANDN U25206 ( .B(n15124), .A(n15125), .Z(n15123) );
XOR U25207 ( .A(c5041), .B(b[5041]), .Z(n15124) );
XNOR U25208 ( .A(b[5041]), .B(n15125), .Z(c[5041]) );
XNOR U25209 ( .A(a[5041]), .B(c5041), .Z(n15125) );
XOR U25210 ( .A(c5042), .B(n15126), .Z(c5043) );
ANDN U25211 ( .B(n15127), .A(n15128), .Z(n15126) );
XOR U25212 ( .A(c5042), .B(b[5042]), .Z(n15127) );
XNOR U25213 ( .A(b[5042]), .B(n15128), .Z(c[5042]) );
XNOR U25214 ( .A(a[5042]), .B(c5042), .Z(n15128) );
XOR U25215 ( .A(c5043), .B(n15129), .Z(c5044) );
ANDN U25216 ( .B(n15130), .A(n15131), .Z(n15129) );
XOR U25217 ( .A(c5043), .B(b[5043]), .Z(n15130) );
XNOR U25218 ( .A(b[5043]), .B(n15131), .Z(c[5043]) );
XNOR U25219 ( .A(a[5043]), .B(c5043), .Z(n15131) );
XOR U25220 ( .A(c5044), .B(n15132), .Z(c5045) );
ANDN U25221 ( .B(n15133), .A(n15134), .Z(n15132) );
XOR U25222 ( .A(c5044), .B(b[5044]), .Z(n15133) );
XNOR U25223 ( .A(b[5044]), .B(n15134), .Z(c[5044]) );
XNOR U25224 ( .A(a[5044]), .B(c5044), .Z(n15134) );
XOR U25225 ( .A(c5045), .B(n15135), .Z(c5046) );
ANDN U25226 ( .B(n15136), .A(n15137), .Z(n15135) );
XOR U25227 ( .A(c5045), .B(b[5045]), .Z(n15136) );
XNOR U25228 ( .A(b[5045]), .B(n15137), .Z(c[5045]) );
XNOR U25229 ( .A(a[5045]), .B(c5045), .Z(n15137) );
XOR U25230 ( .A(c5046), .B(n15138), .Z(c5047) );
ANDN U25231 ( .B(n15139), .A(n15140), .Z(n15138) );
XOR U25232 ( .A(c5046), .B(b[5046]), .Z(n15139) );
XNOR U25233 ( .A(b[5046]), .B(n15140), .Z(c[5046]) );
XNOR U25234 ( .A(a[5046]), .B(c5046), .Z(n15140) );
XOR U25235 ( .A(c5047), .B(n15141), .Z(c5048) );
ANDN U25236 ( .B(n15142), .A(n15143), .Z(n15141) );
XOR U25237 ( .A(c5047), .B(b[5047]), .Z(n15142) );
XNOR U25238 ( .A(b[5047]), .B(n15143), .Z(c[5047]) );
XNOR U25239 ( .A(a[5047]), .B(c5047), .Z(n15143) );
XOR U25240 ( .A(c5048), .B(n15144), .Z(c5049) );
ANDN U25241 ( .B(n15145), .A(n15146), .Z(n15144) );
XOR U25242 ( .A(c5048), .B(b[5048]), .Z(n15145) );
XNOR U25243 ( .A(b[5048]), .B(n15146), .Z(c[5048]) );
XNOR U25244 ( .A(a[5048]), .B(c5048), .Z(n15146) );
XOR U25245 ( .A(c5049), .B(n15147), .Z(c5050) );
ANDN U25246 ( .B(n15148), .A(n15149), .Z(n15147) );
XOR U25247 ( .A(c5049), .B(b[5049]), .Z(n15148) );
XNOR U25248 ( .A(b[5049]), .B(n15149), .Z(c[5049]) );
XNOR U25249 ( .A(a[5049]), .B(c5049), .Z(n15149) );
XOR U25250 ( .A(c5050), .B(n15150), .Z(c5051) );
ANDN U25251 ( .B(n15151), .A(n15152), .Z(n15150) );
XOR U25252 ( .A(c5050), .B(b[5050]), .Z(n15151) );
XNOR U25253 ( .A(b[5050]), .B(n15152), .Z(c[5050]) );
XNOR U25254 ( .A(a[5050]), .B(c5050), .Z(n15152) );
XOR U25255 ( .A(c5051), .B(n15153), .Z(c5052) );
ANDN U25256 ( .B(n15154), .A(n15155), .Z(n15153) );
XOR U25257 ( .A(c5051), .B(b[5051]), .Z(n15154) );
XNOR U25258 ( .A(b[5051]), .B(n15155), .Z(c[5051]) );
XNOR U25259 ( .A(a[5051]), .B(c5051), .Z(n15155) );
XOR U25260 ( .A(c5052), .B(n15156), .Z(c5053) );
ANDN U25261 ( .B(n15157), .A(n15158), .Z(n15156) );
XOR U25262 ( .A(c5052), .B(b[5052]), .Z(n15157) );
XNOR U25263 ( .A(b[5052]), .B(n15158), .Z(c[5052]) );
XNOR U25264 ( .A(a[5052]), .B(c5052), .Z(n15158) );
XOR U25265 ( .A(c5053), .B(n15159), .Z(c5054) );
ANDN U25266 ( .B(n15160), .A(n15161), .Z(n15159) );
XOR U25267 ( .A(c5053), .B(b[5053]), .Z(n15160) );
XNOR U25268 ( .A(b[5053]), .B(n15161), .Z(c[5053]) );
XNOR U25269 ( .A(a[5053]), .B(c5053), .Z(n15161) );
XOR U25270 ( .A(c5054), .B(n15162), .Z(c5055) );
ANDN U25271 ( .B(n15163), .A(n15164), .Z(n15162) );
XOR U25272 ( .A(c5054), .B(b[5054]), .Z(n15163) );
XNOR U25273 ( .A(b[5054]), .B(n15164), .Z(c[5054]) );
XNOR U25274 ( .A(a[5054]), .B(c5054), .Z(n15164) );
XOR U25275 ( .A(c5055), .B(n15165), .Z(c5056) );
ANDN U25276 ( .B(n15166), .A(n15167), .Z(n15165) );
XOR U25277 ( .A(c5055), .B(b[5055]), .Z(n15166) );
XNOR U25278 ( .A(b[5055]), .B(n15167), .Z(c[5055]) );
XNOR U25279 ( .A(a[5055]), .B(c5055), .Z(n15167) );
XOR U25280 ( .A(c5056), .B(n15168), .Z(c5057) );
ANDN U25281 ( .B(n15169), .A(n15170), .Z(n15168) );
XOR U25282 ( .A(c5056), .B(b[5056]), .Z(n15169) );
XNOR U25283 ( .A(b[5056]), .B(n15170), .Z(c[5056]) );
XNOR U25284 ( .A(a[5056]), .B(c5056), .Z(n15170) );
XOR U25285 ( .A(c5057), .B(n15171), .Z(c5058) );
ANDN U25286 ( .B(n15172), .A(n15173), .Z(n15171) );
XOR U25287 ( .A(c5057), .B(b[5057]), .Z(n15172) );
XNOR U25288 ( .A(b[5057]), .B(n15173), .Z(c[5057]) );
XNOR U25289 ( .A(a[5057]), .B(c5057), .Z(n15173) );
XOR U25290 ( .A(c5058), .B(n15174), .Z(c5059) );
ANDN U25291 ( .B(n15175), .A(n15176), .Z(n15174) );
XOR U25292 ( .A(c5058), .B(b[5058]), .Z(n15175) );
XNOR U25293 ( .A(b[5058]), .B(n15176), .Z(c[5058]) );
XNOR U25294 ( .A(a[5058]), .B(c5058), .Z(n15176) );
XOR U25295 ( .A(c5059), .B(n15177), .Z(c5060) );
ANDN U25296 ( .B(n15178), .A(n15179), .Z(n15177) );
XOR U25297 ( .A(c5059), .B(b[5059]), .Z(n15178) );
XNOR U25298 ( .A(b[5059]), .B(n15179), .Z(c[5059]) );
XNOR U25299 ( .A(a[5059]), .B(c5059), .Z(n15179) );
XOR U25300 ( .A(c5060), .B(n15180), .Z(c5061) );
ANDN U25301 ( .B(n15181), .A(n15182), .Z(n15180) );
XOR U25302 ( .A(c5060), .B(b[5060]), .Z(n15181) );
XNOR U25303 ( .A(b[5060]), .B(n15182), .Z(c[5060]) );
XNOR U25304 ( .A(a[5060]), .B(c5060), .Z(n15182) );
XOR U25305 ( .A(c5061), .B(n15183), .Z(c5062) );
ANDN U25306 ( .B(n15184), .A(n15185), .Z(n15183) );
XOR U25307 ( .A(c5061), .B(b[5061]), .Z(n15184) );
XNOR U25308 ( .A(b[5061]), .B(n15185), .Z(c[5061]) );
XNOR U25309 ( .A(a[5061]), .B(c5061), .Z(n15185) );
XOR U25310 ( .A(c5062), .B(n15186), .Z(c5063) );
ANDN U25311 ( .B(n15187), .A(n15188), .Z(n15186) );
XOR U25312 ( .A(c5062), .B(b[5062]), .Z(n15187) );
XNOR U25313 ( .A(b[5062]), .B(n15188), .Z(c[5062]) );
XNOR U25314 ( .A(a[5062]), .B(c5062), .Z(n15188) );
XOR U25315 ( .A(c5063), .B(n15189), .Z(c5064) );
ANDN U25316 ( .B(n15190), .A(n15191), .Z(n15189) );
XOR U25317 ( .A(c5063), .B(b[5063]), .Z(n15190) );
XNOR U25318 ( .A(b[5063]), .B(n15191), .Z(c[5063]) );
XNOR U25319 ( .A(a[5063]), .B(c5063), .Z(n15191) );
XOR U25320 ( .A(c5064), .B(n15192), .Z(c5065) );
ANDN U25321 ( .B(n15193), .A(n15194), .Z(n15192) );
XOR U25322 ( .A(c5064), .B(b[5064]), .Z(n15193) );
XNOR U25323 ( .A(b[5064]), .B(n15194), .Z(c[5064]) );
XNOR U25324 ( .A(a[5064]), .B(c5064), .Z(n15194) );
XOR U25325 ( .A(c5065), .B(n15195), .Z(c5066) );
ANDN U25326 ( .B(n15196), .A(n15197), .Z(n15195) );
XOR U25327 ( .A(c5065), .B(b[5065]), .Z(n15196) );
XNOR U25328 ( .A(b[5065]), .B(n15197), .Z(c[5065]) );
XNOR U25329 ( .A(a[5065]), .B(c5065), .Z(n15197) );
XOR U25330 ( .A(c5066), .B(n15198), .Z(c5067) );
ANDN U25331 ( .B(n15199), .A(n15200), .Z(n15198) );
XOR U25332 ( .A(c5066), .B(b[5066]), .Z(n15199) );
XNOR U25333 ( .A(b[5066]), .B(n15200), .Z(c[5066]) );
XNOR U25334 ( .A(a[5066]), .B(c5066), .Z(n15200) );
XOR U25335 ( .A(c5067), .B(n15201), .Z(c5068) );
ANDN U25336 ( .B(n15202), .A(n15203), .Z(n15201) );
XOR U25337 ( .A(c5067), .B(b[5067]), .Z(n15202) );
XNOR U25338 ( .A(b[5067]), .B(n15203), .Z(c[5067]) );
XNOR U25339 ( .A(a[5067]), .B(c5067), .Z(n15203) );
XOR U25340 ( .A(c5068), .B(n15204), .Z(c5069) );
ANDN U25341 ( .B(n15205), .A(n15206), .Z(n15204) );
XOR U25342 ( .A(c5068), .B(b[5068]), .Z(n15205) );
XNOR U25343 ( .A(b[5068]), .B(n15206), .Z(c[5068]) );
XNOR U25344 ( .A(a[5068]), .B(c5068), .Z(n15206) );
XOR U25345 ( .A(c5069), .B(n15207), .Z(c5070) );
ANDN U25346 ( .B(n15208), .A(n15209), .Z(n15207) );
XOR U25347 ( .A(c5069), .B(b[5069]), .Z(n15208) );
XNOR U25348 ( .A(b[5069]), .B(n15209), .Z(c[5069]) );
XNOR U25349 ( .A(a[5069]), .B(c5069), .Z(n15209) );
XOR U25350 ( .A(c5070), .B(n15210), .Z(c5071) );
ANDN U25351 ( .B(n15211), .A(n15212), .Z(n15210) );
XOR U25352 ( .A(c5070), .B(b[5070]), .Z(n15211) );
XNOR U25353 ( .A(b[5070]), .B(n15212), .Z(c[5070]) );
XNOR U25354 ( .A(a[5070]), .B(c5070), .Z(n15212) );
XOR U25355 ( .A(c5071), .B(n15213), .Z(c5072) );
ANDN U25356 ( .B(n15214), .A(n15215), .Z(n15213) );
XOR U25357 ( .A(c5071), .B(b[5071]), .Z(n15214) );
XNOR U25358 ( .A(b[5071]), .B(n15215), .Z(c[5071]) );
XNOR U25359 ( .A(a[5071]), .B(c5071), .Z(n15215) );
XOR U25360 ( .A(c5072), .B(n15216), .Z(c5073) );
ANDN U25361 ( .B(n15217), .A(n15218), .Z(n15216) );
XOR U25362 ( .A(c5072), .B(b[5072]), .Z(n15217) );
XNOR U25363 ( .A(b[5072]), .B(n15218), .Z(c[5072]) );
XNOR U25364 ( .A(a[5072]), .B(c5072), .Z(n15218) );
XOR U25365 ( .A(c5073), .B(n15219), .Z(c5074) );
ANDN U25366 ( .B(n15220), .A(n15221), .Z(n15219) );
XOR U25367 ( .A(c5073), .B(b[5073]), .Z(n15220) );
XNOR U25368 ( .A(b[5073]), .B(n15221), .Z(c[5073]) );
XNOR U25369 ( .A(a[5073]), .B(c5073), .Z(n15221) );
XOR U25370 ( .A(c5074), .B(n15222), .Z(c5075) );
ANDN U25371 ( .B(n15223), .A(n15224), .Z(n15222) );
XOR U25372 ( .A(c5074), .B(b[5074]), .Z(n15223) );
XNOR U25373 ( .A(b[5074]), .B(n15224), .Z(c[5074]) );
XNOR U25374 ( .A(a[5074]), .B(c5074), .Z(n15224) );
XOR U25375 ( .A(c5075), .B(n15225), .Z(c5076) );
ANDN U25376 ( .B(n15226), .A(n15227), .Z(n15225) );
XOR U25377 ( .A(c5075), .B(b[5075]), .Z(n15226) );
XNOR U25378 ( .A(b[5075]), .B(n15227), .Z(c[5075]) );
XNOR U25379 ( .A(a[5075]), .B(c5075), .Z(n15227) );
XOR U25380 ( .A(c5076), .B(n15228), .Z(c5077) );
ANDN U25381 ( .B(n15229), .A(n15230), .Z(n15228) );
XOR U25382 ( .A(c5076), .B(b[5076]), .Z(n15229) );
XNOR U25383 ( .A(b[5076]), .B(n15230), .Z(c[5076]) );
XNOR U25384 ( .A(a[5076]), .B(c5076), .Z(n15230) );
XOR U25385 ( .A(c5077), .B(n15231), .Z(c5078) );
ANDN U25386 ( .B(n15232), .A(n15233), .Z(n15231) );
XOR U25387 ( .A(c5077), .B(b[5077]), .Z(n15232) );
XNOR U25388 ( .A(b[5077]), .B(n15233), .Z(c[5077]) );
XNOR U25389 ( .A(a[5077]), .B(c5077), .Z(n15233) );
XOR U25390 ( .A(c5078), .B(n15234), .Z(c5079) );
ANDN U25391 ( .B(n15235), .A(n15236), .Z(n15234) );
XOR U25392 ( .A(c5078), .B(b[5078]), .Z(n15235) );
XNOR U25393 ( .A(b[5078]), .B(n15236), .Z(c[5078]) );
XNOR U25394 ( .A(a[5078]), .B(c5078), .Z(n15236) );
XOR U25395 ( .A(c5079), .B(n15237), .Z(c5080) );
ANDN U25396 ( .B(n15238), .A(n15239), .Z(n15237) );
XOR U25397 ( .A(c5079), .B(b[5079]), .Z(n15238) );
XNOR U25398 ( .A(b[5079]), .B(n15239), .Z(c[5079]) );
XNOR U25399 ( .A(a[5079]), .B(c5079), .Z(n15239) );
XOR U25400 ( .A(c5080), .B(n15240), .Z(c5081) );
ANDN U25401 ( .B(n15241), .A(n15242), .Z(n15240) );
XOR U25402 ( .A(c5080), .B(b[5080]), .Z(n15241) );
XNOR U25403 ( .A(b[5080]), .B(n15242), .Z(c[5080]) );
XNOR U25404 ( .A(a[5080]), .B(c5080), .Z(n15242) );
XOR U25405 ( .A(c5081), .B(n15243), .Z(c5082) );
ANDN U25406 ( .B(n15244), .A(n15245), .Z(n15243) );
XOR U25407 ( .A(c5081), .B(b[5081]), .Z(n15244) );
XNOR U25408 ( .A(b[5081]), .B(n15245), .Z(c[5081]) );
XNOR U25409 ( .A(a[5081]), .B(c5081), .Z(n15245) );
XOR U25410 ( .A(c5082), .B(n15246), .Z(c5083) );
ANDN U25411 ( .B(n15247), .A(n15248), .Z(n15246) );
XOR U25412 ( .A(c5082), .B(b[5082]), .Z(n15247) );
XNOR U25413 ( .A(b[5082]), .B(n15248), .Z(c[5082]) );
XNOR U25414 ( .A(a[5082]), .B(c5082), .Z(n15248) );
XOR U25415 ( .A(c5083), .B(n15249), .Z(c5084) );
ANDN U25416 ( .B(n15250), .A(n15251), .Z(n15249) );
XOR U25417 ( .A(c5083), .B(b[5083]), .Z(n15250) );
XNOR U25418 ( .A(b[5083]), .B(n15251), .Z(c[5083]) );
XNOR U25419 ( .A(a[5083]), .B(c5083), .Z(n15251) );
XOR U25420 ( .A(c5084), .B(n15252), .Z(c5085) );
ANDN U25421 ( .B(n15253), .A(n15254), .Z(n15252) );
XOR U25422 ( .A(c5084), .B(b[5084]), .Z(n15253) );
XNOR U25423 ( .A(b[5084]), .B(n15254), .Z(c[5084]) );
XNOR U25424 ( .A(a[5084]), .B(c5084), .Z(n15254) );
XOR U25425 ( .A(c5085), .B(n15255), .Z(c5086) );
ANDN U25426 ( .B(n15256), .A(n15257), .Z(n15255) );
XOR U25427 ( .A(c5085), .B(b[5085]), .Z(n15256) );
XNOR U25428 ( .A(b[5085]), .B(n15257), .Z(c[5085]) );
XNOR U25429 ( .A(a[5085]), .B(c5085), .Z(n15257) );
XOR U25430 ( .A(c5086), .B(n15258), .Z(c5087) );
ANDN U25431 ( .B(n15259), .A(n15260), .Z(n15258) );
XOR U25432 ( .A(c5086), .B(b[5086]), .Z(n15259) );
XNOR U25433 ( .A(b[5086]), .B(n15260), .Z(c[5086]) );
XNOR U25434 ( .A(a[5086]), .B(c5086), .Z(n15260) );
XOR U25435 ( .A(c5087), .B(n15261), .Z(c5088) );
ANDN U25436 ( .B(n15262), .A(n15263), .Z(n15261) );
XOR U25437 ( .A(c5087), .B(b[5087]), .Z(n15262) );
XNOR U25438 ( .A(b[5087]), .B(n15263), .Z(c[5087]) );
XNOR U25439 ( .A(a[5087]), .B(c5087), .Z(n15263) );
XOR U25440 ( .A(c5088), .B(n15264), .Z(c5089) );
ANDN U25441 ( .B(n15265), .A(n15266), .Z(n15264) );
XOR U25442 ( .A(c5088), .B(b[5088]), .Z(n15265) );
XNOR U25443 ( .A(b[5088]), .B(n15266), .Z(c[5088]) );
XNOR U25444 ( .A(a[5088]), .B(c5088), .Z(n15266) );
XOR U25445 ( .A(c5089), .B(n15267), .Z(c5090) );
ANDN U25446 ( .B(n15268), .A(n15269), .Z(n15267) );
XOR U25447 ( .A(c5089), .B(b[5089]), .Z(n15268) );
XNOR U25448 ( .A(b[5089]), .B(n15269), .Z(c[5089]) );
XNOR U25449 ( .A(a[5089]), .B(c5089), .Z(n15269) );
XOR U25450 ( .A(c5090), .B(n15270), .Z(c5091) );
ANDN U25451 ( .B(n15271), .A(n15272), .Z(n15270) );
XOR U25452 ( .A(c5090), .B(b[5090]), .Z(n15271) );
XNOR U25453 ( .A(b[5090]), .B(n15272), .Z(c[5090]) );
XNOR U25454 ( .A(a[5090]), .B(c5090), .Z(n15272) );
XOR U25455 ( .A(c5091), .B(n15273), .Z(c5092) );
ANDN U25456 ( .B(n15274), .A(n15275), .Z(n15273) );
XOR U25457 ( .A(c5091), .B(b[5091]), .Z(n15274) );
XNOR U25458 ( .A(b[5091]), .B(n15275), .Z(c[5091]) );
XNOR U25459 ( .A(a[5091]), .B(c5091), .Z(n15275) );
XOR U25460 ( .A(c5092), .B(n15276), .Z(c5093) );
ANDN U25461 ( .B(n15277), .A(n15278), .Z(n15276) );
XOR U25462 ( .A(c5092), .B(b[5092]), .Z(n15277) );
XNOR U25463 ( .A(b[5092]), .B(n15278), .Z(c[5092]) );
XNOR U25464 ( .A(a[5092]), .B(c5092), .Z(n15278) );
XOR U25465 ( .A(c5093), .B(n15279), .Z(c5094) );
ANDN U25466 ( .B(n15280), .A(n15281), .Z(n15279) );
XOR U25467 ( .A(c5093), .B(b[5093]), .Z(n15280) );
XNOR U25468 ( .A(b[5093]), .B(n15281), .Z(c[5093]) );
XNOR U25469 ( .A(a[5093]), .B(c5093), .Z(n15281) );
XOR U25470 ( .A(c5094), .B(n15282), .Z(c5095) );
ANDN U25471 ( .B(n15283), .A(n15284), .Z(n15282) );
XOR U25472 ( .A(c5094), .B(b[5094]), .Z(n15283) );
XNOR U25473 ( .A(b[5094]), .B(n15284), .Z(c[5094]) );
XNOR U25474 ( .A(a[5094]), .B(c5094), .Z(n15284) );
XOR U25475 ( .A(c5095), .B(n15285), .Z(c5096) );
ANDN U25476 ( .B(n15286), .A(n15287), .Z(n15285) );
XOR U25477 ( .A(c5095), .B(b[5095]), .Z(n15286) );
XNOR U25478 ( .A(b[5095]), .B(n15287), .Z(c[5095]) );
XNOR U25479 ( .A(a[5095]), .B(c5095), .Z(n15287) );
XOR U25480 ( .A(c5096), .B(n15288), .Z(c5097) );
ANDN U25481 ( .B(n15289), .A(n15290), .Z(n15288) );
XOR U25482 ( .A(c5096), .B(b[5096]), .Z(n15289) );
XNOR U25483 ( .A(b[5096]), .B(n15290), .Z(c[5096]) );
XNOR U25484 ( .A(a[5096]), .B(c5096), .Z(n15290) );
XOR U25485 ( .A(c5097), .B(n15291), .Z(c5098) );
ANDN U25486 ( .B(n15292), .A(n15293), .Z(n15291) );
XOR U25487 ( .A(c5097), .B(b[5097]), .Z(n15292) );
XNOR U25488 ( .A(b[5097]), .B(n15293), .Z(c[5097]) );
XNOR U25489 ( .A(a[5097]), .B(c5097), .Z(n15293) );
XOR U25490 ( .A(c5098), .B(n15294), .Z(c5099) );
ANDN U25491 ( .B(n15295), .A(n15296), .Z(n15294) );
XOR U25492 ( .A(c5098), .B(b[5098]), .Z(n15295) );
XNOR U25493 ( .A(b[5098]), .B(n15296), .Z(c[5098]) );
XNOR U25494 ( .A(a[5098]), .B(c5098), .Z(n15296) );
XOR U25495 ( .A(c5099), .B(n15297), .Z(c5100) );
ANDN U25496 ( .B(n15298), .A(n15299), .Z(n15297) );
XOR U25497 ( .A(c5099), .B(b[5099]), .Z(n15298) );
XNOR U25498 ( .A(b[5099]), .B(n15299), .Z(c[5099]) );
XNOR U25499 ( .A(a[5099]), .B(c5099), .Z(n15299) );
XOR U25500 ( .A(c5100), .B(n15300), .Z(c5101) );
ANDN U25501 ( .B(n15301), .A(n15302), .Z(n15300) );
XOR U25502 ( .A(c5100), .B(b[5100]), .Z(n15301) );
XNOR U25503 ( .A(b[5100]), .B(n15302), .Z(c[5100]) );
XNOR U25504 ( .A(a[5100]), .B(c5100), .Z(n15302) );
XOR U25505 ( .A(c5101), .B(n15303), .Z(c5102) );
ANDN U25506 ( .B(n15304), .A(n15305), .Z(n15303) );
XOR U25507 ( .A(c5101), .B(b[5101]), .Z(n15304) );
XNOR U25508 ( .A(b[5101]), .B(n15305), .Z(c[5101]) );
XNOR U25509 ( .A(a[5101]), .B(c5101), .Z(n15305) );
XOR U25510 ( .A(c5102), .B(n15306), .Z(c5103) );
ANDN U25511 ( .B(n15307), .A(n15308), .Z(n15306) );
XOR U25512 ( .A(c5102), .B(b[5102]), .Z(n15307) );
XNOR U25513 ( .A(b[5102]), .B(n15308), .Z(c[5102]) );
XNOR U25514 ( .A(a[5102]), .B(c5102), .Z(n15308) );
XOR U25515 ( .A(c5103), .B(n15309), .Z(c5104) );
ANDN U25516 ( .B(n15310), .A(n15311), .Z(n15309) );
XOR U25517 ( .A(c5103), .B(b[5103]), .Z(n15310) );
XNOR U25518 ( .A(b[5103]), .B(n15311), .Z(c[5103]) );
XNOR U25519 ( .A(a[5103]), .B(c5103), .Z(n15311) );
XOR U25520 ( .A(c5104), .B(n15312), .Z(c5105) );
ANDN U25521 ( .B(n15313), .A(n15314), .Z(n15312) );
XOR U25522 ( .A(c5104), .B(b[5104]), .Z(n15313) );
XNOR U25523 ( .A(b[5104]), .B(n15314), .Z(c[5104]) );
XNOR U25524 ( .A(a[5104]), .B(c5104), .Z(n15314) );
XOR U25525 ( .A(c5105), .B(n15315), .Z(c5106) );
ANDN U25526 ( .B(n15316), .A(n15317), .Z(n15315) );
XOR U25527 ( .A(c5105), .B(b[5105]), .Z(n15316) );
XNOR U25528 ( .A(b[5105]), .B(n15317), .Z(c[5105]) );
XNOR U25529 ( .A(a[5105]), .B(c5105), .Z(n15317) );
XOR U25530 ( .A(c5106), .B(n15318), .Z(c5107) );
ANDN U25531 ( .B(n15319), .A(n15320), .Z(n15318) );
XOR U25532 ( .A(c5106), .B(b[5106]), .Z(n15319) );
XNOR U25533 ( .A(b[5106]), .B(n15320), .Z(c[5106]) );
XNOR U25534 ( .A(a[5106]), .B(c5106), .Z(n15320) );
XOR U25535 ( .A(c5107), .B(n15321), .Z(c5108) );
ANDN U25536 ( .B(n15322), .A(n15323), .Z(n15321) );
XOR U25537 ( .A(c5107), .B(b[5107]), .Z(n15322) );
XNOR U25538 ( .A(b[5107]), .B(n15323), .Z(c[5107]) );
XNOR U25539 ( .A(a[5107]), .B(c5107), .Z(n15323) );
XOR U25540 ( .A(c5108), .B(n15324), .Z(c5109) );
ANDN U25541 ( .B(n15325), .A(n15326), .Z(n15324) );
XOR U25542 ( .A(c5108), .B(b[5108]), .Z(n15325) );
XNOR U25543 ( .A(b[5108]), .B(n15326), .Z(c[5108]) );
XNOR U25544 ( .A(a[5108]), .B(c5108), .Z(n15326) );
XOR U25545 ( .A(c5109), .B(n15327), .Z(c5110) );
ANDN U25546 ( .B(n15328), .A(n15329), .Z(n15327) );
XOR U25547 ( .A(c5109), .B(b[5109]), .Z(n15328) );
XNOR U25548 ( .A(b[5109]), .B(n15329), .Z(c[5109]) );
XNOR U25549 ( .A(a[5109]), .B(c5109), .Z(n15329) );
XOR U25550 ( .A(c5110), .B(n15330), .Z(c5111) );
ANDN U25551 ( .B(n15331), .A(n15332), .Z(n15330) );
XOR U25552 ( .A(c5110), .B(b[5110]), .Z(n15331) );
XNOR U25553 ( .A(b[5110]), .B(n15332), .Z(c[5110]) );
XNOR U25554 ( .A(a[5110]), .B(c5110), .Z(n15332) );
XOR U25555 ( .A(c5111), .B(n15333), .Z(c5112) );
ANDN U25556 ( .B(n15334), .A(n15335), .Z(n15333) );
XOR U25557 ( .A(c5111), .B(b[5111]), .Z(n15334) );
XNOR U25558 ( .A(b[5111]), .B(n15335), .Z(c[5111]) );
XNOR U25559 ( .A(a[5111]), .B(c5111), .Z(n15335) );
XOR U25560 ( .A(c5112), .B(n15336), .Z(c5113) );
ANDN U25561 ( .B(n15337), .A(n15338), .Z(n15336) );
XOR U25562 ( .A(c5112), .B(b[5112]), .Z(n15337) );
XNOR U25563 ( .A(b[5112]), .B(n15338), .Z(c[5112]) );
XNOR U25564 ( .A(a[5112]), .B(c5112), .Z(n15338) );
XOR U25565 ( .A(c5113), .B(n15339), .Z(c5114) );
ANDN U25566 ( .B(n15340), .A(n15341), .Z(n15339) );
XOR U25567 ( .A(c5113), .B(b[5113]), .Z(n15340) );
XNOR U25568 ( .A(b[5113]), .B(n15341), .Z(c[5113]) );
XNOR U25569 ( .A(a[5113]), .B(c5113), .Z(n15341) );
XOR U25570 ( .A(c5114), .B(n15342), .Z(c5115) );
ANDN U25571 ( .B(n15343), .A(n15344), .Z(n15342) );
XOR U25572 ( .A(c5114), .B(b[5114]), .Z(n15343) );
XNOR U25573 ( .A(b[5114]), .B(n15344), .Z(c[5114]) );
XNOR U25574 ( .A(a[5114]), .B(c5114), .Z(n15344) );
XOR U25575 ( .A(c5115), .B(n15345), .Z(c5116) );
ANDN U25576 ( .B(n15346), .A(n15347), .Z(n15345) );
XOR U25577 ( .A(c5115), .B(b[5115]), .Z(n15346) );
XNOR U25578 ( .A(b[5115]), .B(n15347), .Z(c[5115]) );
XNOR U25579 ( .A(a[5115]), .B(c5115), .Z(n15347) );
XOR U25580 ( .A(c5116), .B(n15348), .Z(c5117) );
ANDN U25581 ( .B(n15349), .A(n15350), .Z(n15348) );
XOR U25582 ( .A(c5116), .B(b[5116]), .Z(n15349) );
XNOR U25583 ( .A(b[5116]), .B(n15350), .Z(c[5116]) );
XNOR U25584 ( .A(a[5116]), .B(c5116), .Z(n15350) );
XOR U25585 ( .A(c5117), .B(n15351), .Z(c5118) );
ANDN U25586 ( .B(n15352), .A(n15353), .Z(n15351) );
XOR U25587 ( .A(c5117), .B(b[5117]), .Z(n15352) );
XNOR U25588 ( .A(b[5117]), .B(n15353), .Z(c[5117]) );
XNOR U25589 ( .A(a[5117]), .B(c5117), .Z(n15353) );
XOR U25590 ( .A(c5118), .B(n15354), .Z(c5119) );
ANDN U25591 ( .B(n15355), .A(n15356), .Z(n15354) );
XOR U25592 ( .A(c5118), .B(b[5118]), .Z(n15355) );
XNOR U25593 ( .A(b[5118]), .B(n15356), .Z(c[5118]) );
XNOR U25594 ( .A(a[5118]), .B(c5118), .Z(n15356) );
XOR U25595 ( .A(c5119), .B(n15357), .Z(c5120) );
ANDN U25596 ( .B(n15358), .A(n15359), .Z(n15357) );
XOR U25597 ( .A(c5119), .B(b[5119]), .Z(n15358) );
XNOR U25598 ( .A(b[5119]), .B(n15359), .Z(c[5119]) );
XNOR U25599 ( .A(a[5119]), .B(c5119), .Z(n15359) );
XOR U25600 ( .A(c5120), .B(n15360), .Z(c5121) );
ANDN U25601 ( .B(n15361), .A(n15362), .Z(n15360) );
XOR U25602 ( .A(c5120), .B(b[5120]), .Z(n15361) );
XNOR U25603 ( .A(b[5120]), .B(n15362), .Z(c[5120]) );
XNOR U25604 ( .A(a[5120]), .B(c5120), .Z(n15362) );
XOR U25605 ( .A(c5121), .B(n15363), .Z(c5122) );
ANDN U25606 ( .B(n15364), .A(n15365), .Z(n15363) );
XOR U25607 ( .A(c5121), .B(b[5121]), .Z(n15364) );
XNOR U25608 ( .A(b[5121]), .B(n15365), .Z(c[5121]) );
XNOR U25609 ( .A(a[5121]), .B(c5121), .Z(n15365) );
XOR U25610 ( .A(c5122), .B(n15366), .Z(c5123) );
ANDN U25611 ( .B(n15367), .A(n15368), .Z(n15366) );
XOR U25612 ( .A(c5122), .B(b[5122]), .Z(n15367) );
XNOR U25613 ( .A(b[5122]), .B(n15368), .Z(c[5122]) );
XNOR U25614 ( .A(a[5122]), .B(c5122), .Z(n15368) );
XOR U25615 ( .A(c5123), .B(n15369), .Z(c5124) );
ANDN U25616 ( .B(n15370), .A(n15371), .Z(n15369) );
XOR U25617 ( .A(c5123), .B(b[5123]), .Z(n15370) );
XNOR U25618 ( .A(b[5123]), .B(n15371), .Z(c[5123]) );
XNOR U25619 ( .A(a[5123]), .B(c5123), .Z(n15371) );
XOR U25620 ( .A(c5124), .B(n15372), .Z(c5125) );
ANDN U25621 ( .B(n15373), .A(n15374), .Z(n15372) );
XOR U25622 ( .A(c5124), .B(b[5124]), .Z(n15373) );
XNOR U25623 ( .A(b[5124]), .B(n15374), .Z(c[5124]) );
XNOR U25624 ( .A(a[5124]), .B(c5124), .Z(n15374) );
XOR U25625 ( .A(c5125), .B(n15375), .Z(c5126) );
ANDN U25626 ( .B(n15376), .A(n15377), .Z(n15375) );
XOR U25627 ( .A(c5125), .B(b[5125]), .Z(n15376) );
XNOR U25628 ( .A(b[5125]), .B(n15377), .Z(c[5125]) );
XNOR U25629 ( .A(a[5125]), .B(c5125), .Z(n15377) );
XOR U25630 ( .A(c5126), .B(n15378), .Z(c5127) );
ANDN U25631 ( .B(n15379), .A(n15380), .Z(n15378) );
XOR U25632 ( .A(c5126), .B(b[5126]), .Z(n15379) );
XNOR U25633 ( .A(b[5126]), .B(n15380), .Z(c[5126]) );
XNOR U25634 ( .A(a[5126]), .B(c5126), .Z(n15380) );
XOR U25635 ( .A(c5127), .B(n15381), .Z(c5128) );
ANDN U25636 ( .B(n15382), .A(n15383), .Z(n15381) );
XOR U25637 ( .A(c5127), .B(b[5127]), .Z(n15382) );
XNOR U25638 ( .A(b[5127]), .B(n15383), .Z(c[5127]) );
XNOR U25639 ( .A(a[5127]), .B(c5127), .Z(n15383) );
XOR U25640 ( .A(c5128), .B(n15384), .Z(c5129) );
ANDN U25641 ( .B(n15385), .A(n15386), .Z(n15384) );
XOR U25642 ( .A(c5128), .B(b[5128]), .Z(n15385) );
XNOR U25643 ( .A(b[5128]), .B(n15386), .Z(c[5128]) );
XNOR U25644 ( .A(a[5128]), .B(c5128), .Z(n15386) );
XOR U25645 ( .A(c5129), .B(n15387), .Z(c5130) );
ANDN U25646 ( .B(n15388), .A(n15389), .Z(n15387) );
XOR U25647 ( .A(c5129), .B(b[5129]), .Z(n15388) );
XNOR U25648 ( .A(b[5129]), .B(n15389), .Z(c[5129]) );
XNOR U25649 ( .A(a[5129]), .B(c5129), .Z(n15389) );
XOR U25650 ( .A(c5130), .B(n15390), .Z(c5131) );
ANDN U25651 ( .B(n15391), .A(n15392), .Z(n15390) );
XOR U25652 ( .A(c5130), .B(b[5130]), .Z(n15391) );
XNOR U25653 ( .A(b[5130]), .B(n15392), .Z(c[5130]) );
XNOR U25654 ( .A(a[5130]), .B(c5130), .Z(n15392) );
XOR U25655 ( .A(c5131), .B(n15393), .Z(c5132) );
ANDN U25656 ( .B(n15394), .A(n15395), .Z(n15393) );
XOR U25657 ( .A(c5131), .B(b[5131]), .Z(n15394) );
XNOR U25658 ( .A(b[5131]), .B(n15395), .Z(c[5131]) );
XNOR U25659 ( .A(a[5131]), .B(c5131), .Z(n15395) );
XOR U25660 ( .A(c5132), .B(n15396), .Z(c5133) );
ANDN U25661 ( .B(n15397), .A(n15398), .Z(n15396) );
XOR U25662 ( .A(c5132), .B(b[5132]), .Z(n15397) );
XNOR U25663 ( .A(b[5132]), .B(n15398), .Z(c[5132]) );
XNOR U25664 ( .A(a[5132]), .B(c5132), .Z(n15398) );
XOR U25665 ( .A(c5133), .B(n15399), .Z(c5134) );
ANDN U25666 ( .B(n15400), .A(n15401), .Z(n15399) );
XOR U25667 ( .A(c5133), .B(b[5133]), .Z(n15400) );
XNOR U25668 ( .A(b[5133]), .B(n15401), .Z(c[5133]) );
XNOR U25669 ( .A(a[5133]), .B(c5133), .Z(n15401) );
XOR U25670 ( .A(c5134), .B(n15402), .Z(c5135) );
ANDN U25671 ( .B(n15403), .A(n15404), .Z(n15402) );
XOR U25672 ( .A(c5134), .B(b[5134]), .Z(n15403) );
XNOR U25673 ( .A(b[5134]), .B(n15404), .Z(c[5134]) );
XNOR U25674 ( .A(a[5134]), .B(c5134), .Z(n15404) );
XOR U25675 ( .A(c5135), .B(n15405), .Z(c5136) );
ANDN U25676 ( .B(n15406), .A(n15407), .Z(n15405) );
XOR U25677 ( .A(c5135), .B(b[5135]), .Z(n15406) );
XNOR U25678 ( .A(b[5135]), .B(n15407), .Z(c[5135]) );
XNOR U25679 ( .A(a[5135]), .B(c5135), .Z(n15407) );
XOR U25680 ( .A(c5136), .B(n15408), .Z(c5137) );
ANDN U25681 ( .B(n15409), .A(n15410), .Z(n15408) );
XOR U25682 ( .A(c5136), .B(b[5136]), .Z(n15409) );
XNOR U25683 ( .A(b[5136]), .B(n15410), .Z(c[5136]) );
XNOR U25684 ( .A(a[5136]), .B(c5136), .Z(n15410) );
XOR U25685 ( .A(c5137), .B(n15411), .Z(c5138) );
ANDN U25686 ( .B(n15412), .A(n15413), .Z(n15411) );
XOR U25687 ( .A(c5137), .B(b[5137]), .Z(n15412) );
XNOR U25688 ( .A(b[5137]), .B(n15413), .Z(c[5137]) );
XNOR U25689 ( .A(a[5137]), .B(c5137), .Z(n15413) );
XOR U25690 ( .A(c5138), .B(n15414), .Z(c5139) );
ANDN U25691 ( .B(n15415), .A(n15416), .Z(n15414) );
XOR U25692 ( .A(c5138), .B(b[5138]), .Z(n15415) );
XNOR U25693 ( .A(b[5138]), .B(n15416), .Z(c[5138]) );
XNOR U25694 ( .A(a[5138]), .B(c5138), .Z(n15416) );
XOR U25695 ( .A(c5139), .B(n15417), .Z(c5140) );
ANDN U25696 ( .B(n15418), .A(n15419), .Z(n15417) );
XOR U25697 ( .A(c5139), .B(b[5139]), .Z(n15418) );
XNOR U25698 ( .A(b[5139]), .B(n15419), .Z(c[5139]) );
XNOR U25699 ( .A(a[5139]), .B(c5139), .Z(n15419) );
XOR U25700 ( .A(c5140), .B(n15420), .Z(c5141) );
ANDN U25701 ( .B(n15421), .A(n15422), .Z(n15420) );
XOR U25702 ( .A(c5140), .B(b[5140]), .Z(n15421) );
XNOR U25703 ( .A(b[5140]), .B(n15422), .Z(c[5140]) );
XNOR U25704 ( .A(a[5140]), .B(c5140), .Z(n15422) );
XOR U25705 ( .A(c5141), .B(n15423), .Z(c5142) );
ANDN U25706 ( .B(n15424), .A(n15425), .Z(n15423) );
XOR U25707 ( .A(c5141), .B(b[5141]), .Z(n15424) );
XNOR U25708 ( .A(b[5141]), .B(n15425), .Z(c[5141]) );
XNOR U25709 ( .A(a[5141]), .B(c5141), .Z(n15425) );
XOR U25710 ( .A(c5142), .B(n15426), .Z(c5143) );
ANDN U25711 ( .B(n15427), .A(n15428), .Z(n15426) );
XOR U25712 ( .A(c5142), .B(b[5142]), .Z(n15427) );
XNOR U25713 ( .A(b[5142]), .B(n15428), .Z(c[5142]) );
XNOR U25714 ( .A(a[5142]), .B(c5142), .Z(n15428) );
XOR U25715 ( .A(c5143), .B(n15429), .Z(c5144) );
ANDN U25716 ( .B(n15430), .A(n15431), .Z(n15429) );
XOR U25717 ( .A(c5143), .B(b[5143]), .Z(n15430) );
XNOR U25718 ( .A(b[5143]), .B(n15431), .Z(c[5143]) );
XNOR U25719 ( .A(a[5143]), .B(c5143), .Z(n15431) );
XOR U25720 ( .A(c5144), .B(n15432), .Z(c5145) );
ANDN U25721 ( .B(n15433), .A(n15434), .Z(n15432) );
XOR U25722 ( .A(c5144), .B(b[5144]), .Z(n15433) );
XNOR U25723 ( .A(b[5144]), .B(n15434), .Z(c[5144]) );
XNOR U25724 ( .A(a[5144]), .B(c5144), .Z(n15434) );
XOR U25725 ( .A(c5145), .B(n15435), .Z(c5146) );
ANDN U25726 ( .B(n15436), .A(n15437), .Z(n15435) );
XOR U25727 ( .A(c5145), .B(b[5145]), .Z(n15436) );
XNOR U25728 ( .A(b[5145]), .B(n15437), .Z(c[5145]) );
XNOR U25729 ( .A(a[5145]), .B(c5145), .Z(n15437) );
XOR U25730 ( .A(c5146), .B(n15438), .Z(c5147) );
ANDN U25731 ( .B(n15439), .A(n15440), .Z(n15438) );
XOR U25732 ( .A(c5146), .B(b[5146]), .Z(n15439) );
XNOR U25733 ( .A(b[5146]), .B(n15440), .Z(c[5146]) );
XNOR U25734 ( .A(a[5146]), .B(c5146), .Z(n15440) );
XOR U25735 ( .A(c5147), .B(n15441), .Z(c5148) );
ANDN U25736 ( .B(n15442), .A(n15443), .Z(n15441) );
XOR U25737 ( .A(c5147), .B(b[5147]), .Z(n15442) );
XNOR U25738 ( .A(b[5147]), .B(n15443), .Z(c[5147]) );
XNOR U25739 ( .A(a[5147]), .B(c5147), .Z(n15443) );
XOR U25740 ( .A(c5148), .B(n15444), .Z(c5149) );
ANDN U25741 ( .B(n15445), .A(n15446), .Z(n15444) );
XOR U25742 ( .A(c5148), .B(b[5148]), .Z(n15445) );
XNOR U25743 ( .A(b[5148]), .B(n15446), .Z(c[5148]) );
XNOR U25744 ( .A(a[5148]), .B(c5148), .Z(n15446) );
XOR U25745 ( .A(c5149), .B(n15447), .Z(c5150) );
ANDN U25746 ( .B(n15448), .A(n15449), .Z(n15447) );
XOR U25747 ( .A(c5149), .B(b[5149]), .Z(n15448) );
XNOR U25748 ( .A(b[5149]), .B(n15449), .Z(c[5149]) );
XNOR U25749 ( .A(a[5149]), .B(c5149), .Z(n15449) );
XOR U25750 ( .A(c5150), .B(n15450), .Z(c5151) );
ANDN U25751 ( .B(n15451), .A(n15452), .Z(n15450) );
XOR U25752 ( .A(c5150), .B(b[5150]), .Z(n15451) );
XNOR U25753 ( .A(b[5150]), .B(n15452), .Z(c[5150]) );
XNOR U25754 ( .A(a[5150]), .B(c5150), .Z(n15452) );
XOR U25755 ( .A(c5151), .B(n15453), .Z(c5152) );
ANDN U25756 ( .B(n15454), .A(n15455), .Z(n15453) );
XOR U25757 ( .A(c5151), .B(b[5151]), .Z(n15454) );
XNOR U25758 ( .A(b[5151]), .B(n15455), .Z(c[5151]) );
XNOR U25759 ( .A(a[5151]), .B(c5151), .Z(n15455) );
XOR U25760 ( .A(c5152), .B(n15456), .Z(c5153) );
ANDN U25761 ( .B(n15457), .A(n15458), .Z(n15456) );
XOR U25762 ( .A(c5152), .B(b[5152]), .Z(n15457) );
XNOR U25763 ( .A(b[5152]), .B(n15458), .Z(c[5152]) );
XNOR U25764 ( .A(a[5152]), .B(c5152), .Z(n15458) );
XOR U25765 ( .A(c5153), .B(n15459), .Z(c5154) );
ANDN U25766 ( .B(n15460), .A(n15461), .Z(n15459) );
XOR U25767 ( .A(c5153), .B(b[5153]), .Z(n15460) );
XNOR U25768 ( .A(b[5153]), .B(n15461), .Z(c[5153]) );
XNOR U25769 ( .A(a[5153]), .B(c5153), .Z(n15461) );
XOR U25770 ( .A(c5154), .B(n15462), .Z(c5155) );
ANDN U25771 ( .B(n15463), .A(n15464), .Z(n15462) );
XOR U25772 ( .A(c5154), .B(b[5154]), .Z(n15463) );
XNOR U25773 ( .A(b[5154]), .B(n15464), .Z(c[5154]) );
XNOR U25774 ( .A(a[5154]), .B(c5154), .Z(n15464) );
XOR U25775 ( .A(c5155), .B(n15465), .Z(c5156) );
ANDN U25776 ( .B(n15466), .A(n15467), .Z(n15465) );
XOR U25777 ( .A(c5155), .B(b[5155]), .Z(n15466) );
XNOR U25778 ( .A(b[5155]), .B(n15467), .Z(c[5155]) );
XNOR U25779 ( .A(a[5155]), .B(c5155), .Z(n15467) );
XOR U25780 ( .A(c5156), .B(n15468), .Z(c5157) );
ANDN U25781 ( .B(n15469), .A(n15470), .Z(n15468) );
XOR U25782 ( .A(c5156), .B(b[5156]), .Z(n15469) );
XNOR U25783 ( .A(b[5156]), .B(n15470), .Z(c[5156]) );
XNOR U25784 ( .A(a[5156]), .B(c5156), .Z(n15470) );
XOR U25785 ( .A(c5157), .B(n15471), .Z(c5158) );
ANDN U25786 ( .B(n15472), .A(n15473), .Z(n15471) );
XOR U25787 ( .A(c5157), .B(b[5157]), .Z(n15472) );
XNOR U25788 ( .A(b[5157]), .B(n15473), .Z(c[5157]) );
XNOR U25789 ( .A(a[5157]), .B(c5157), .Z(n15473) );
XOR U25790 ( .A(c5158), .B(n15474), .Z(c5159) );
ANDN U25791 ( .B(n15475), .A(n15476), .Z(n15474) );
XOR U25792 ( .A(c5158), .B(b[5158]), .Z(n15475) );
XNOR U25793 ( .A(b[5158]), .B(n15476), .Z(c[5158]) );
XNOR U25794 ( .A(a[5158]), .B(c5158), .Z(n15476) );
XOR U25795 ( .A(c5159), .B(n15477), .Z(c5160) );
ANDN U25796 ( .B(n15478), .A(n15479), .Z(n15477) );
XOR U25797 ( .A(c5159), .B(b[5159]), .Z(n15478) );
XNOR U25798 ( .A(b[5159]), .B(n15479), .Z(c[5159]) );
XNOR U25799 ( .A(a[5159]), .B(c5159), .Z(n15479) );
XOR U25800 ( .A(c5160), .B(n15480), .Z(c5161) );
ANDN U25801 ( .B(n15481), .A(n15482), .Z(n15480) );
XOR U25802 ( .A(c5160), .B(b[5160]), .Z(n15481) );
XNOR U25803 ( .A(b[5160]), .B(n15482), .Z(c[5160]) );
XNOR U25804 ( .A(a[5160]), .B(c5160), .Z(n15482) );
XOR U25805 ( .A(c5161), .B(n15483), .Z(c5162) );
ANDN U25806 ( .B(n15484), .A(n15485), .Z(n15483) );
XOR U25807 ( .A(c5161), .B(b[5161]), .Z(n15484) );
XNOR U25808 ( .A(b[5161]), .B(n15485), .Z(c[5161]) );
XNOR U25809 ( .A(a[5161]), .B(c5161), .Z(n15485) );
XOR U25810 ( .A(c5162), .B(n15486), .Z(c5163) );
ANDN U25811 ( .B(n15487), .A(n15488), .Z(n15486) );
XOR U25812 ( .A(c5162), .B(b[5162]), .Z(n15487) );
XNOR U25813 ( .A(b[5162]), .B(n15488), .Z(c[5162]) );
XNOR U25814 ( .A(a[5162]), .B(c5162), .Z(n15488) );
XOR U25815 ( .A(c5163), .B(n15489), .Z(c5164) );
ANDN U25816 ( .B(n15490), .A(n15491), .Z(n15489) );
XOR U25817 ( .A(c5163), .B(b[5163]), .Z(n15490) );
XNOR U25818 ( .A(b[5163]), .B(n15491), .Z(c[5163]) );
XNOR U25819 ( .A(a[5163]), .B(c5163), .Z(n15491) );
XOR U25820 ( .A(c5164), .B(n15492), .Z(c5165) );
ANDN U25821 ( .B(n15493), .A(n15494), .Z(n15492) );
XOR U25822 ( .A(c5164), .B(b[5164]), .Z(n15493) );
XNOR U25823 ( .A(b[5164]), .B(n15494), .Z(c[5164]) );
XNOR U25824 ( .A(a[5164]), .B(c5164), .Z(n15494) );
XOR U25825 ( .A(c5165), .B(n15495), .Z(c5166) );
ANDN U25826 ( .B(n15496), .A(n15497), .Z(n15495) );
XOR U25827 ( .A(c5165), .B(b[5165]), .Z(n15496) );
XNOR U25828 ( .A(b[5165]), .B(n15497), .Z(c[5165]) );
XNOR U25829 ( .A(a[5165]), .B(c5165), .Z(n15497) );
XOR U25830 ( .A(c5166), .B(n15498), .Z(c5167) );
ANDN U25831 ( .B(n15499), .A(n15500), .Z(n15498) );
XOR U25832 ( .A(c5166), .B(b[5166]), .Z(n15499) );
XNOR U25833 ( .A(b[5166]), .B(n15500), .Z(c[5166]) );
XNOR U25834 ( .A(a[5166]), .B(c5166), .Z(n15500) );
XOR U25835 ( .A(c5167), .B(n15501), .Z(c5168) );
ANDN U25836 ( .B(n15502), .A(n15503), .Z(n15501) );
XOR U25837 ( .A(c5167), .B(b[5167]), .Z(n15502) );
XNOR U25838 ( .A(b[5167]), .B(n15503), .Z(c[5167]) );
XNOR U25839 ( .A(a[5167]), .B(c5167), .Z(n15503) );
XOR U25840 ( .A(c5168), .B(n15504), .Z(c5169) );
ANDN U25841 ( .B(n15505), .A(n15506), .Z(n15504) );
XOR U25842 ( .A(c5168), .B(b[5168]), .Z(n15505) );
XNOR U25843 ( .A(b[5168]), .B(n15506), .Z(c[5168]) );
XNOR U25844 ( .A(a[5168]), .B(c5168), .Z(n15506) );
XOR U25845 ( .A(c5169), .B(n15507), .Z(c5170) );
ANDN U25846 ( .B(n15508), .A(n15509), .Z(n15507) );
XOR U25847 ( .A(c5169), .B(b[5169]), .Z(n15508) );
XNOR U25848 ( .A(b[5169]), .B(n15509), .Z(c[5169]) );
XNOR U25849 ( .A(a[5169]), .B(c5169), .Z(n15509) );
XOR U25850 ( .A(c5170), .B(n15510), .Z(c5171) );
ANDN U25851 ( .B(n15511), .A(n15512), .Z(n15510) );
XOR U25852 ( .A(c5170), .B(b[5170]), .Z(n15511) );
XNOR U25853 ( .A(b[5170]), .B(n15512), .Z(c[5170]) );
XNOR U25854 ( .A(a[5170]), .B(c5170), .Z(n15512) );
XOR U25855 ( .A(c5171), .B(n15513), .Z(c5172) );
ANDN U25856 ( .B(n15514), .A(n15515), .Z(n15513) );
XOR U25857 ( .A(c5171), .B(b[5171]), .Z(n15514) );
XNOR U25858 ( .A(b[5171]), .B(n15515), .Z(c[5171]) );
XNOR U25859 ( .A(a[5171]), .B(c5171), .Z(n15515) );
XOR U25860 ( .A(c5172), .B(n15516), .Z(c5173) );
ANDN U25861 ( .B(n15517), .A(n15518), .Z(n15516) );
XOR U25862 ( .A(c5172), .B(b[5172]), .Z(n15517) );
XNOR U25863 ( .A(b[5172]), .B(n15518), .Z(c[5172]) );
XNOR U25864 ( .A(a[5172]), .B(c5172), .Z(n15518) );
XOR U25865 ( .A(c5173), .B(n15519), .Z(c5174) );
ANDN U25866 ( .B(n15520), .A(n15521), .Z(n15519) );
XOR U25867 ( .A(c5173), .B(b[5173]), .Z(n15520) );
XNOR U25868 ( .A(b[5173]), .B(n15521), .Z(c[5173]) );
XNOR U25869 ( .A(a[5173]), .B(c5173), .Z(n15521) );
XOR U25870 ( .A(c5174), .B(n15522), .Z(c5175) );
ANDN U25871 ( .B(n15523), .A(n15524), .Z(n15522) );
XOR U25872 ( .A(c5174), .B(b[5174]), .Z(n15523) );
XNOR U25873 ( .A(b[5174]), .B(n15524), .Z(c[5174]) );
XNOR U25874 ( .A(a[5174]), .B(c5174), .Z(n15524) );
XOR U25875 ( .A(c5175), .B(n15525), .Z(c5176) );
ANDN U25876 ( .B(n15526), .A(n15527), .Z(n15525) );
XOR U25877 ( .A(c5175), .B(b[5175]), .Z(n15526) );
XNOR U25878 ( .A(b[5175]), .B(n15527), .Z(c[5175]) );
XNOR U25879 ( .A(a[5175]), .B(c5175), .Z(n15527) );
XOR U25880 ( .A(c5176), .B(n15528), .Z(c5177) );
ANDN U25881 ( .B(n15529), .A(n15530), .Z(n15528) );
XOR U25882 ( .A(c5176), .B(b[5176]), .Z(n15529) );
XNOR U25883 ( .A(b[5176]), .B(n15530), .Z(c[5176]) );
XNOR U25884 ( .A(a[5176]), .B(c5176), .Z(n15530) );
XOR U25885 ( .A(c5177), .B(n15531), .Z(c5178) );
ANDN U25886 ( .B(n15532), .A(n15533), .Z(n15531) );
XOR U25887 ( .A(c5177), .B(b[5177]), .Z(n15532) );
XNOR U25888 ( .A(b[5177]), .B(n15533), .Z(c[5177]) );
XNOR U25889 ( .A(a[5177]), .B(c5177), .Z(n15533) );
XOR U25890 ( .A(c5178), .B(n15534), .Z(c5179) );
ANDN U25891 ( .B(n15535), .A(n15536), .Z(n15534) );
XOR U25892 ( .A(c5178), .B(b[5178]), .Z(n15535) );
XNOR U25893 ( .A(b[5178]), .B(n15536), .Z(c[5178]) );
XNOR U25894 ( .A(a[5178]), .B(c5178), .Z(n15536) );
XOR U25895 ( .A(c5179), .B(n15537), .Z(c5180) );
ANDN U25896 ( .B(n15538), .A(n15539), .Z(n15537) );
XOR U25897 ( .A(c5179), .B(b[5179]), .Z(n15538) );
XNOR U25898 ( .A(b[5179]), .B(n15539), .Z(c[5179]) );
XNOR U25899 ( .A(a[5179]), .B(c5179), .Z(n15539) );
XOR U25900 ( .A(c5180), .B(n15540), .Z(c5181) );
ANDN U25901 ( .B(n15541), .A(n15542), .Z(n15540) );
XOR U25902 ( .A(c5180), .B(b[5180]), .Z(n15541) );
XNOR U25903 ( .A(b[5180]), .B(n15542), .Z(c[5180]) );
XNOR U25904 ( .A(a[5180]), .B(c5180), .Z(n15542) );
XOR U25905 ( .A(c5181), .B(n15543), .Z(c5182) );
ANDN U25906 ( .B(n15544), .A(n15545), .Z(n15543) );
XOR U25907 ( .A(c5181), .B(b[5181]), .Z(n15544) );
XNOR U25908 ( .A(b[5181]), .B(n15545), .Z(c[5181]) );
XNOR U25909 ( .A(a[5181]), .B(c5181), .Z(n15545) );
XOR U25910 ( .A(c5182), .B(n15546), .Z(c5183) );
ANDN U25911 ( .B(n15547), .A(n15548), .Z(n15546) );
XOR U25912 ( .A(c5182), .B(b[5182]), .Z(n15547) );
XNOR U25913 ( .A(b[5182]), .B(n15548), .Z(c[5182]) );
XNOR U25914 ( .A(a[5182]), .B(c5182), .Z(n15548) );
XOR U25915 ( .A(c5183), .B(n15549), .Z(c5184) );
ANDN U25916 ( .B(n15550), .A(n15551), .Z(n15549) );
XOR U25917 ( .A(c5183), .B(b[5183]), .Z(n15550) );
XNOR U25918 ( .A(b[5183]), .B(n15551), .Z(c[5183]) );
XNOR U25919 ( .A(a[5183]), .B(c5183), .Z(n15551) );
XOR U25920 ( .A(c5184), .B(n15552), .Z(c5185) );
ANDN U25921 ( .B(n15553), .A(n15554), .Z(n15552) );
XOR U25922 ( .A(c5184), .B(b[5184]), .Z(n15553) );
XNOR U25923 ( .A(b[5184]), .B(n15554), .Z(c[5184]) );
XNOR U25924 ( .A(a[5184]), .B(c5184), .Z(n15554) );
XOR U25925 ( .A(c5185), .B(n15555), .Z(c5186) );
ANDN U25926 ( .B(n15556), .A(n15557), .Z(n15555) );
XOR U25927 ( .A(c5185), .B(b[5185]), .Z(n15556) );
XNOR U25928 ( .A(b[5185]), .B(n15557), .Z(c[5185]) );
XNOR U25929 ( .A(a[5185]), .B(c5185), .Z(n15557) );
XOR U25930 ( .A(c5186), .B(n15558), .Z(c5187) );
ANDN U25931 ( .B(n15559), .A(n15560), .Z(n15558) );
XOR U25932 ( .A(c5186), .B(b[5186]), .Z(n15559) );
XNOR U25933 ( .A(b[5186]), .B(n15560), .Z(c[5186]) );
XNOR U25934 ( .A(a[5186]), .B(c5186), .Z(n15560) );
XOR U25935 ( .A(c5187), .B(n15561), .Z(c5188) );
ANDN U25936 ( .B(n15562), .A(n15563), .Z(n15561) );
XOR U25937 ( .A(c5187), .B(b[5187]), .Z(n15562) );
XNOR U25938 ( .A(b[5187]), .B(n15563), .Z(c[5187]) );
XNOR U25939 ( .A(a[5187]), .B(c5187), .Z(n15563) );
XOR U25940 ( .A(c5188), .B(n15564), .Z(c5189) );
ANDN U25941 ( .B(n15565), .A(n15566), .Z(n15564) );
XOR U25942 ( .A(c5188), .B(b[5188]), .Z(n15565) );
XNOR U25943 ( .A(b[5188]), .B(n15566), .Z(c[5188]) );
XNOR U25944 ( .A(a[5188]), .B(c5188), .Z(n15566) );
XOR U25945 ( .A(c5189), .B(n15567), .Z(c5190) );
ANDN U25946 ( .B(n15568), .A(n15569), .Z(n15567) );
XOR U25947 ( .A(c5189), .B(b[5189]), .Z(n15568) );
XNOR U25948 ( .A(b[5189]), .B(n15569), .Z(c[5189]) );
XNOR U25949 ( .A(a[5189]), .B(c5189), .Z(n15569) );
XOR U25950 ( .A(c5190), .B(n15570), .Z(c5191) );
ANDN U25951 ( .B(n15571), .A(n15572), .Z(n15570) );
XOR U25952 ( .A(c5190), .B(b[5190]), .Z(n15571) );
XNOR U25953 ( .A(b[5190]), .B(n15572), .Z(c[5190]) );
XNOR U25954 ( .A(a[5190]), .B(c5190), .Z(n15572) );
XOR U25955 ( .A(c5191), .B(n15573), .Z(c5192) );
ANDN U25956 ( .B(n15574), .A(n15575), .Z(n15573) );
XOR U25957 ( .A(c5191), .B(b[5191]), .Z(n15574) );
XNOR U25958 ( .A(b[5191]), .B(n15575), .Z(c[5191]) );
XNOR U25959 ( .A(a[5191]), .B(c5191), .Z(n15575) );
XOR U25960 ( .A(c5192), .B(n15576), .Z(c5193) );
ANDN U25961 ( .B(n15577), .A(n15578), .Z(n15576) );
XOR U25962 ( .A(c5192), .B(b[5192]), .Z(n15577) );
XNOR U25963 ( .A(b[5192]), .B(n15578), .Z(c[5192]) );
XNOR U25964 ( .A(a[5192]), .B(c5192), .Z(n15578) );
XOR U25965 ( .A(c5193), .B(n15579), .Z(c5194) );
ANDN U25966 ( .B(n15580), .A(n15581), .Z(n15579) );
XOR U25967 ( .A(c5193), .B(b[5193]), .Z(n15580) );
XNOR U25968 ( .A(b[5193]), .B(n15581), .Z(c[5193]) );
XNOR U25969 ( .A(a[5193]), .B(c5193), .Z(n15581) );
XOR U25970 ( .A(c5194), .B(n15582), .Z(c5195) );
ANDN U25971 ( .B(n15583), .A(n15584), .Z(n15582) );
XOR U25972 ( .A(c5194), .B(b[5194]), .Z(n15583) );
XNOR U25973 ( .A(b[5194]), .B(n15584), .Z(c[5194]) );
XNOR U25974 ( .A(a[5194]), .B(c5194), .Z(n15584) );
XOR U25975 ( .A(c5195), .B(n15585), .Z(c5196) );
ANDN U25976 ( .B(n15586), .A(n15587), .Z(n15585) );
XOR U25977 ( .A(c5195), .B(b[5195]), .Z(n15586) );
XNOR U25978 ( .A(b[5195]), .B(n15587), .Z(c[5195]) );
XNOR U25979 ( .A(a[5195]), .B(c5195), .Z(n15587) );
XOR U25980 ( .A(c5196), .B(n15588), .Z(c5197) );
ANDN U25981 ( .B(n15589), .A(n15590), .Z(n15588) );
XOR U25982 ( .A(c5196), .B(b[5196]), .Z(n15589) );
XNOR U25983 ( .A(b[5196]), .B(n15590), .Z(c[5196]) );
XNOR U25984 ( .A(a[5196]), .B(c5196), .Z(n15590) );
XOR U25985 ( .A(c5197), .B(n15591), .Z(c5198) );
ANDN U25986 ( .B(n15592), .A(n15593), .Z(n15591) );
XOR U25987 ( .A(c5197), .B(b[5197]), .Z(n15592) );
XNOR U25988 ( .A(b[5197]), .B(n15593), .Z(c[5197]) );
XNOR U25989 ( .A(a[5197]), .B(c5197), .Z(n15593) );
XOR U25990 ( .A(c5198), .B(n15594), .Z(c5199) );
ANDN U25991 ( .B(n15595), .A(n15596), .Z(n15594) );
XOR U25992 ( .A(c5198), .B(b[5198]), .Z(n15595) );
XNOR U25993 ( .A(b[5198]), .B(n15596), .Z(c[5198]) );
XNOR U25994 ( .A(a[5198]), .B(c5198), .Z(n15596) );
XOR U25995 ( .A(c5199), .B(n15597), .Z(c5200) );
ANDN U25996 ( .B(n15598), .A(n15599), .Z(n15597) );
XOR U25997 ( .A(c5199), .B(b[5199]), .Z(n15598) );
XNOR U25998 ( .A(b[5199]), .B(n15599), .Z(c[5199]) );
XNOR U25999 ( .A(a[5199]), .B(c5199), .Z(n15599) );
XOR U26000 ( .A(c5200), .B(n15600), .Z(c5201) );
ANDN U26001 ( .B(n15601), .A(n15602), .Z(n15600) );
XOR U26002 ( .A(c5200), .B(b[5200]), .Z(n15601) );
XNOR U26003 ( .A(b[5200]), .B(n15602), .Z(c[5200]) );
XNOR U26004 ( .A(a[5200]), .B(c5200), .Z(n15602) );
XOR U26005 ( .A(c5201), .B(n15603), .Z(c5202) );
ANDN U26006 ( .B(n15604), .A(n15605), .Z(n15603) );
XOR U26007 ( .A(c5201), .B(b[5201]), .Z(n15604) );
XNOR U26008 ( .A(b[5201]), .B(n15605), .Z(c[5201]) );
XNOR U26009 ( .A(a[5201]), .B(c5201), .Z(n15605) );
XOR U26010 ( .A(c5202), .B(n15606), .Z(c5203) );
ANDN U26011 ( .B(n15607), .A(n15608), .Z(n15606) );
XOR U26012 ( .A(c5202), .B(b[5202]), .Z(n15607) );
XNOR U26013 ( .A(b[5202]), .B(n15608), .Z(c[5202]) );
XNOR U26014 ( .A(a[5202]), .B(c5202), .Z(n15608) );
XOR U26015 ( .A(c5203), .B(n15609), .Z(c5204) );
ANDN U26016 ( .B(n15610), .A(n15611), .Z(n15609) );
XOR U26017 ( .A(c5203), .B(b[5203]), .Z(n15610) );
XNOR U26018 ( .A(b[5203]), .B(n15611), .Z(c[5203]) );
XNOR U26019 ( .A(a[5203]), .B(c5203), .Z(n15611) );
XOR U26020 ( .A(c5204), .B(n15612), .Z(c5205) );
ANDN U26021 ( .B(n15613), .A(n15614), .Z(n15612) );
XOR U26022 ( .A(c5204), .B(b[5204]), .Z(n15613) );
XNOR U26023 ( .A(b[5204]), .B(n15614), .Z(c[5204]) );
XNOR U26024 ( .A(a[5204]), .B(c5204), .Z(n15614) );
XOR U26025 ( .A(c5205), .B(n15615), .Z(c5206) );
ANDN U26026 ( .B(n15616), .A(n15617), .Z(n15615) );
XOR U26027 ( .A(c5205), .B(b[5205]), .Z(n15616) );
XNOR U26028 ( .A(b[5205]), .B(n15617), .Z(c[5205]) );
XNOR U26029 ( .A(a[5205]), .B(c5205), .Z(n15617) );
XOR U26030 ( .A(c5206), .B(n15618), .Z(c5207) );
ANDN U26031 ( .B(n15619), .A(n15620), .Z(n15618) );
XOR U26032 ( .A(c5206), .B(b[5206]), .Z(n15619) );
XNOR U26033 ( .A(b[5206]), .B(n15620), .Z(c[5206]) );
XNOR U26034 ( .A(a[5206]), .B(c5206), .Z(n15620) );
XOR U26035 ( .A(c5207), .B(n15621), .Z(c5208) );
ANDN U26036 ( .B(n15622), .A(n15623), .Z(n15621) );
XOR U26037 ( .A(c5207), .B(b[5207]), .Z(n15622) );
XNOR U26038 ( .A(b[5207]), .B(n15623), .Z(c[5207]) );
XNOR U26039 ( .A(a[5207]), .B(c5207), .Z(n15623) );
XOR U26040 ( .A(c5208), .B(n15624), .Z(c5209) );
ANDN U26041 ( .B(n15625), .A(n15626), .Z(n15624) );
XOR U26042 ( .A(c5208), .B(b[5208]), .Z(n15625) );
XNOR U26043 ( .A(b[5208]), .B(n15626), .Z(c[5208]) );
XNOR U26044 ( .A(a[5208]), .B(c5208), .Z(n15626) );
XOR U26045 ( .A(c5209), .B(n15627), .Z(c5210) );
ANDN U26046 ( .B(n15628), .A(n15629), .Z(n15627) );
XOR U26047 ( .A(c5209), .B(b[5209]), .Z(n15628) );
XNOR U26048 ( .A(b[5209]), .B(n15629), .Z(c[5209]) );
XNOR U26049 ( .A(a[5209]), .B(c5209), .Z(n15629) );
XOR U26050 ( .A(c5210), .B(n15630), .Z(c5211) );
ANDN U26051 ( .B(n15631), .A(n15632), .Z(n15630) );
XOR U26052 ( .A(c5210), .B(b[5210]), .Z(n15631) );
XNOR U26053 ( .A(b[5210]), .B(n15632), .Z(c[5210]) );
XNOR U26054 ( .A(a[5210]), .B(c5210), .Z(n15632) );
XOR U26055 ( .A(c5211), .B(n15633), .Z(c5212) );
ANDN U26056 ( .B(n15634), .A(n15635), .Z(n15633) );
XOR U26057 ( .A(c5211), .B(b[5211]), .Z(n15634) );
XNOR U26058 ( .A(b[5211]), .B(n15635), .Z(c[5211]) );
XNOR U26059 ( .A(a[5211]), .B(c5211), .Z(n15635) );
XOR U26060 ( .A(c5212), .B(n15636), .Z(c5213) );
ANDN U26061 ( .B(n15637), .A(n15638), .Z(n15636) );
XOR U26062 ( .A(c5212), .B(b[5212]), .Z(n15637) );
XNOR U26063 ( .A(b[5212]), .B(n15638), .Z(c[5212]) );
XNOR U26064 ( .A(a[5212]), .B(c5212), .Z(n15638) );
XOR U26065 ( .A(c5213), .B(n15639), .Z(c5214) );
ANDN U26066 ( .B(n15640), .A(n15641), .Z(n15639) );
XOR U26067 ( .A(c5213), .B(b[5213]), .Z(n15640) );
XNOR U26068 ( .A(b[5213]), .B(n15641), .Z(c[5213]) );
XNOR U26069 ( .A(a[5213]), .B(c5213), .Z(n15641) );
XOR U26070 ( .A(c5214), .B(n15642), .Z(c5215) );
ANDN U26071 ( .B(n15643), .A(n15644), .Z(n15642) );
XOR U26072 ( .A(c5214), .B(b[5214]), .Z(n15643) );
XNOR U26073 ( .A(b[5214]), .B(n15644), .Z(c[5214]) );
XNOR U26074 ( .A(a[5214]), .B(c5214), .Z(n15644) );
XOR U26075 ( .A(c5215), .B(n15645), .Z(c5216) );
ANDN U26076 ( .B(n15646), .A(n15647), .Z(n15645) );
XOR U26077 ( .A(c5215), .B(b[5215]), .Z(n15646) );
XNOR U26078 ( .A(b[5215]), .B(n15647), .Z(c[5215]) );
XNOR U26079 ( .A(a[5215]), .B(c5215), .Z(n15647) );
XOR U26080 ( .A(c5216), .B(n15648), .Z(c5217) );
ANDN U26081 ( .B(n15649), .A(n15650), .Z(n15648) );
XOR U26082 ( .A(c5216), .B(b[5216]), .Z(n15649) );
XNOR U26083 ( .A(b[5216]), .B(n15650), .Z(c[5216]) );
XNOR U26084 ( .A(a[5216]), .B(c5216), .Z(n15650) );
XOR U26085 ( .A(c5217), .B(n15651), .Z(c5218) );
ANDN U26086 ( .B(n15652), .A(n15653), .Z(n15651) );
XOR U26087 ( .A(c5217), .B(b[5217]), .Z(n15652) );
XNOR U26088 ( .A(b[5217]), .B(n15653), .Z(c[5217]) );
XNOR U26089 ( .A(a[5217]), .B(c5217), .Z(n15653) );
XOR U26090 ( .A(c5218), .B(n15654), .Z(c5219) );
ANDN U26091 ( .B(n15655), .A(n15656), .Z(n15654) );
XOR U26092 ( .A(c5218), .B(b[5218]), .Z(n15655) );
XNOR U26093 ( .A(b[5218]), .B(n15656), .Z(c[5218]) );
XNOR U26094 ( .A(a[5218]), .B(c5218), .Z(n15656) );
XOR U26095 ( .A(c5219), .B(n15657), .Z(c5220) );
ANDN U26096 ( .B(n15658), .A(n15659), .Z(n15657) );
XOR U26097 ( .A(c5219), .B(b[5219]), .Z(n15658) );
XNOR U26098 ( .A(b[5219]), .B(n15659), .Z(c[5219]) );
XNOR U26099 ( .A(a[5219]), .B(c5219), .Z(n15659) );
XOR U26100 ( .A(c5220), .B(n15660), .Z(c5221) );
ANDN U26101 ( .B(n15661), .A(n15662), .Z(n15660) );
XOR U26102 ( .A(c5220), .B(b[5220]), .Z(n15661) );
XNOR U26103 ( .A(b[5220]), .B(n15662), .Z(c[5220]) );
XNOR U26104 ( .A(a[5220]), .B(c5220), .Z(n15662) );
XOR U26105 ( .A(c5221), .B(n15663), .Z(c5222) );
ANDN U26106 ( .B(n15664), .A(n15665), .Z(n15663) );
XOR U26107 ( .A(c5221), .B(b[5221]), .Z(n15664) );
XNOR U26108 ( .A(b[5221]), .B(n15665), .Z(c[5221]) );
XNOR U26109 ( .A(a[5221]), .B(c5221), .Z(n15665) );
XOR U26110 ( .A(c5222), .B(n15666), .Z(c5223) );
ANDN U26111 ( .B(n15667), .A(n15668), .Z(n15666) );
XOR U26112 ( .A(c5222), .B(b[5222]), .Z(n15667) );
XNOR U26113 ( .A(b[5222]), .B(n15668), .Z(c[5222]) );
XNOR U26114 ( .A(a[5222]), .B(c5222), .Z(n15668) );
XOR U26115 ( .A(c5223), .B(n15669), .Z(c5224) );
ANDN U26116 ( .B(n15670), .A(n15671), .Z(n15669) );
XOR U26117 ( .A(c5223), .B(b[5223]), .Z(n15670) );
XNOR U26118 ( .A(b[5223]), .B(n15671), .Z(c[5223]) );
XNOR U26119 ( .A(a[5223]), .B(c5223), .Z(n15671) );
XOR U26120 ( .A(c5224), .B(n15672), .Z(c5225) );
ANDN U26121 ( .B(n15673), .A(n15674), .Z(n15672) );
XOR U26122 ( .A(c5224), .B(b[5224]), .Z(n15673) );
XNOR U26123 ( .A(b[5224]), .B(n15674), .Z(c[5224]) );
XNOR U26124 ( .A(a[5224]), .B(c5224), .Z(n15674) );
XOR U26125 ( .A(c5225), .B(n15675), .Z(c5226) );
ANDN U26126 ( .B(n15676), .A(n15677), .Z(n15675) );
XOR U26127 ( .A(c5225), .B(b[5225]), .Z(n15676) );
XNOR U26128 ( .A(b[5225]), .B(n15677), .Z(c[5225]) );
XNOR U26129 ( .A(a[5225]), .B(c5225), .Z(n15677) );
XOR U26130 ( .A(c5226), .B(n15678), .Z(c5227) );
ANDN U26131 ( .B(n15679), .A(n15680), .Z(n15678) );
XOR U26132 ( .A(c5226), .B(b[5226]), .Z(n15679) );
XNOR U26133 ( .A(b[5226]), .B(n15680), .Z(c[5226]) );
XNOR U26134 ( .A(a[5226]), .B(c5226), .Z(n15680) );
XOR U26135 ( .A(c5227), .B(n15681), .Z(c5228) );
ANDN U26136 ( .B(n15682), .A(n15683), .Z(n15681) );
XOR U26137 ( .A(c5227), .B(b[5227]), .Z(n15682) );
XNOR U26138 ( .A(b[5227]), .B(n15683), .Z(c[5227]) );
XNOR U26139 ( .A(a[5227]), .B(c5227), .Z(n15683) );
XOR U26140 ( .A(c5228), .B(n15684), .Z(c5229) );
ANDN U26141 ( .B(n15685), .A(n15686), .Z(n15684) );
XOR U26142 ( .A(c5228), .B(b[5228]), .Z(n15685) );
XNOR U26143 ( .A(b[5228]), .B(n15686), .Z(c[5228]) );
XNOR U26144 ( .A(a[5228]), .B(c5228), .Z(n15686) );
XOR U26145 ( .A(c5229), .B(n15687), .Z(c5230) );
ANDN U26146 ( .B(n15688), .A(n15689), .Z(n15687) );
XOR U26147 ( .A(c5229), .B(b[5229]), .Z(n15688) );
XNOR U26148 ( .A(b[5229]), .B(n15689), .Z(c[5229]) );
XNOR U26149 ( .A(a[5229]), .B(c5229), .Z(n15689) );
XOR U26150 ( .A(c5230), .B(n15690), .Z(c5231) );
ANDN U26151 ( .B(n15691), .A(n15692), .Z(n15690) );
XOR U26152 ( .A(c5230), .B(b[5230]), .Z(n15691) );
XNOR U26153 ( .A(b[5230]), .B(n15692), .Z(c[5230]) );
XNOR U26154 ( .A(a[5230]), .B(c5230), .Z(n15692) );
XOR U26155 ( .A(c5231), .B(n15693), .Z(c5232) );
ANDN U26156 ( .B(n15694), .A(n15695), .Z(n15693) );
XOR U26157 ( .A(c5231), .B(b[5231]), .Z(n15694) );
XNOR U26158 ( .A(b[5231]), .B(n15695), .Z(c[5231]) );
XNOR U26159 ( .A(a[5231]), .B(c5231), .Z(n15695) );
XOR U26160 ( .A(c5232), .B(n15696), .Z(c5233) );
ANDN U26161 ( .B(n15697), .A(n15698), .Z(n15696) );
XOR U26162 ( .A(c5232), .B(b[5232]), .Z(n15697) );
XNOR U26163 ( .A(b[5232]), .B(n15698), .Z(c[5232]) );
XNOR U26164 ( .A(a[5232]), .B(c5232), .Z(n15698) );
XOR U26165 ( .A(c5233), .B(n15699), .Z(c5234) );
ANDN U26166 ( .B(n15700), .A(n15701), .Z(n15699) );
XOR U26167 ( .A(c5233), .B(b[5233]), .Z(n15700) );
XNOR U26168 ( .A(b[5233]), .B(n15701), .Z(c[5233]) );
XNOR U26169 ( .A(a[5233]), .B(c5233), .Z(n15701) );
XOR U26170 ( .A(c5234), .B(n15702), .Z(c5235) );
ANDN U26171 ( .B(n15703), .A(n15704), .Z(n15702) );
XOR U26172 ( .A(c5234), .B(b[5234]), .Z(n15703) );
XNOR U26173 ( .A(b[5234]), .B(n15704), .Z(c[5234]) );
XNOR U26174 ( .A(a[5234]), .B(c5234), .Z(n15704) );
XOR U26175 ( .A(c5235), .B(n15705), .Z(c5236) );
ANDN U26176 ( .B(n15706), .A(n15707), .Z(n15705) );
XOR U26177 ( .A(c5235), .B(b[5235]), .Z(n15706) );
XNOR U26178 ( .A(b[5235]), .B(n15707), .Z(c[5235]) );
XNOR U26179 ( .A(a[5235]), .B(c5235), .Z(n15707) );
XOR U26180 ( .A(c5236), .B(n15708), .Z(c5237) );
ANDN U26181 ( .B(n15709), .A(n15710), .Z(n15708) );
XOR U26182 ( .A(c5236), .B(b[5236]), .Z(n15709) );
XNOR U26183 ( .A(b[5236]), .B(n15710), .Z(c[5236]) );
XNOR U26184 ( .A(a[5236]), .B(c5236), .Z(n15710) );
XOR U26185 ( .A(c5237), .B(n15711), .Z(c5238) );
ANDN U26186 ( .B(n15712), .A(n15713), .Z(n15711) );
XOR U26187 ( .A(c5237), .B(b[5237]), .Z(n15712) );
XNOR U26188 ( .A(b[5237]), .B(n15713), .Z(c[5237]) );
XNOR U26189 ( .A(a[5237]), .B(c5237), .Z(n15713) );
XOR U26190 ( .A(c5238), .B(n15714), .Z(c5239) );
ANDN U26191 ( .B(n15715), .A(n15716), .Z(n15714) );
XOR U26192 ( .A(c5238), .B(b[5238]), .Z(n15715) );
XNOR U26193 ( .A(b[5238]), .B(n15716), .Z(c[5238]) );
XNOR U26194 ( .A(a[5238]), .B(c5238), .Z(n15716) );
XOR U26195 ( .A(c5239), .B(n15717), .Z(c5240) );
ANDN U26196 ( .B(n15718), .A(n15719), .Z(n15717) );
XOR U26197 ( .A(c5239), .B(b[5239]), .Z(n15718) );
XNOR U26198 ( .A(b[5239]), .B(n15719), .Z(c[5239]) );
XNOR U26199 ( .A(a[5239]), .B(c5239), .Z(n15719) );
XOR U26200 ( .A(c5240), .B(n15720), .Z(c5241) );
ANDN U26201 ( .B(n15721), .A(n15722), .Z(n15720) );
XOR U26202 ( .A(c5240), .B(b[5240]), .Z(n15721) );
XNOR U26203 ( .A(b[5240]), .B(n15722), .Z(c[5240]) );
XNOR U26204 ( .A(a[5240]), .B(c5240), .Z(n15722) );
XOR U26205 ( .A(c5241), .B(n15723), .Z(c5242) );
ANDN U26206 ( .B(n15724), .A(n15725), .Z(n15723) );
XOR U26207 ( .A(c5241), .B(b[5241]), .Z(n15724) );
XNOR U26208 ( .A(b[5241]), .B(n15725), .Z(c[5241]) );
XNOR U26209 ( .A(a[5241]), .B(c5241), .Z(n15725) );
XOR U26210 ( .A(c5242), .B(n15726), .Z(c5243) );
ANDN U26211 ( .B(n15727), .A(n15728), .Z(n15726) );
XOR U26212 ( .A(c5242), .B(b[5242]), .Z(n15727) );
XNOR U26213 ( .A(b[5242]), .B(n15728), .Z(c[5242]) );
XNOR U26214 ( .A(a[5242]), .B(c5242), .Z(n15728) );
XOR U26215 ( .A(c5243), .B(n15729), .Z(c5244) );
ANDN U26216 ( .B(n15730), .A(n15731), .Z(n15729) );
XOR U26217 ( .A(c5243), .B(b[5243]), .Z(n15730) );
XNOR U26218 ( .A(b[5243]), .B(n15731), .Z(c[5243]) );
XNOR U26219 ( .A(a[5243]), .B(c5243), .Z(n15731) );
XOR U26220 ( .A(c5244), .B(n15732), .Z(c5245) );
ANDN U26221 ( .B(n15733), .A(n15734), .Z(n15732) );
XOR U26222 ( .A(c5244), .B(b[5244]), .Z(n15733) );
XNOR U26223 ( .A(b[5244]), .B(n15734), .Z(c[5244]) );
XNOR U26224 ( .A(a[5244]), .B(c5244), .Z(n15734) );
XOR U26225 ( .A(c5245), .B(n15735), .Z(c5246) );
ANDN U26226 ( .B(n15736), .A(n15737), .Z(n15735) );
XOR U26227 ( .A(c5245), .B(b[5245]), .Z(n15736) );
XNOR U26228 ( .A(b[5245]), .B(n15737), .Z(c[5245]) );
XNOR U26229 ( .A(a[5245]), .B(c5245), .Z(n15737) );
XOR U26230 ( .A(c5246), .B(n15738), .Z(c5247) );
ANDN U26231 ( .B(n15739), .A(n15740), .Z(n15738) );
XOR U26232 ( .A(c5246), .B(b[5246]), .Z(n15739) );
XNOR U26233 ( .A(b[5246]), .B(n15740), .Z(c[5246]) );
XNOR U26234 ( .A(a[5246]), .B(c5246), .Z(n15740) );
XOR U26235 ( .A(c5247), .B(n15741), .Z(c5248) );
ANDN U26236 ( .B(n15742), .A(n15743), .Z(n15741) );
XOR U26237 ( .A(c5247), .B(b[5247]), .Z(n15742) );
XNOR U26238 ( .A(b[5247]), .B(n15743), .Z(c[5247]) );
XNOR U26239 ( .A(a[5247]), .B(c5247), .Z(n15743) );
XOR U26240 ( .A(c5248), .B(n15744), .Z(c5249) );
ANDN U26241 ( .B(n15745), .A(n15746), .Z(n15744) );
XOR U26242 ( .A(c5248), .B(b[5248]), .Z(n15745) );
XNOR U26243 ( .A(b[5248]), .B(n15746), .Z(c[5248]) );
XNOR U26244 ( .A(a[5248]), .B(c5248), .Z(n15746) );
XOR U26245 ( .A(c5249), .B(n15747), .Z(c5250) );
ANDN U26246 ( .B(n15748), .A(n15749), .Z(n15747) );
XOR U26247 ( .A(c5249), .B(b[5249]), .Z(n15748) );
XNOR U26248 ( .A(b[5249]), .B(n15749), .Z(c[5249]) );
XNOR U26249 ( .A(a[5249]), .B(c5249), .Z(n15749) );
XOR U26250 ( .A(c5250), .B(n15750), .Z(c5251) );
ANDN U26251 ( .B(n15751), .A(n15752), .Z(n15750) );
XOR U26252 ( .A(c5250), .B(b[5250]), .Z(n15751) );
XNOR U26253 ( .A(b[5250]), .B(n15752), .Z(c[5250]) );
XNOR U26254 ( .A(a[5250]), .B(c5250), .Z(n15752) );
XOR U26255 ( .A(c5251), .B(n15753), .Z(c5252) );
ANDN U26256 ( .B(n15754), .A(n15755), .Z(n15753) );
XOR U26257 ( .A(c5251), .B(b[5251]), .Z(n15754) );
XNOR U26258 ( .A(b[5251]), .B(n15755), .Z(c[5251]) );
XNOR U26259 ( .A(a[5251]), .B(c5251), .Z(n15755) );
XOR U26260 ( .A(c5252), .B(n15756), .Z(c5253) );
ANDN U26261 ( .B(n15757), .A(n15758), .Z(n15756) );
XOR U26262 ( .A(c5252), .B(b[5252]), .Z(n15757) );
XNOR U26263 ( .A(b[5252]), .B(n15758), .Z(c[5252]) );
XNOR U26264 ( .A(a[5252]), .B(c5252), .Z(n15758) );
XOR U26265 ( .A(c5253), .B(n15759), .Z(c5254) );
ANDN U26266 ( .B(n15760), .A(n15761), .Z(n15759) );
XOR U26267 ( .A(c5253), .B(b[5253]), .Z(n15760) );
XNOR U26268 ( .A(b[5253]), .B(n15761), .Z(c[5253]) );
XNOR U26269 ( .A(a[5253]), .B(c5253), .Z(n15761) );
XOR U26270 ( .A(c5254), .B(n15762), .Z(c5255) );
ANDN U26271 ( .B(n15763), .A(n15764), .Z(n15762) );
XOR U26272 ( .A(c5254), .B(b[5254]), .Z(n15763) );
XNOR U26273 ( .A(b[5254]), .B(n15764), .Z(c[5254]) );
XNOR U26274 ( .A(a[5254]), .B(c5254), .Z(n15764) );
XOR U26275 ( .A(c5255), .B(n15765), .Z(c5256) );
ANDN U26276 ( .B(n15766), .A(n15767), .Z(n15765) );
XOR U26277 ( .A(c5255), .B(b[5255]), .Z(n15766) );
XNOR U26278 ( .A(b[5255]), .B(n15767), .Z(c[5255]) );
XNOR U26279 ( .A(a[5255]), .B(c5255), .Z(n15767) );
XOR U26280 ( .A(c5256), .B(n15768), .Z(c5257) );
ANDN U26281 ( .B(n15769), .A(n15770), .Z(n15768) );
XOR U26282 ( .A(c5256), .B(b[5256]), .Z(n15769) );
XNOR U26283 ( .A(b[5256]), .B(n15770), .Z(c[5256]) );
XNOR U26284 ( .A(a[5256]), .B(c5256), .Z(n15770) );
XOR U26285 ( .A(c5257), .B(n15771), .Z(c5258) );
ANDN U26286 ( .B(n15772), .A(n15773), .Z(n15771) );
XOR U26287 ( .A(c5257), .B(b[5257]), .Z(n15772) );
XNOR U26288 ( .A(b[5257]), .B(n15773), .Z(c[5257]) );
XNOR U26289 ( .A(a[5257]), .B(c5257), .Z(n15773) );
XOR U26290 ( .A(c5258), .B(n15774), .Z(c5259) );
ANDN U26291 ( .B(n15775), .A(n15776), .Z(n15774) );
XOR U26292 ( .A(c5258), .B(b[5258]), .Z(n15775) );
XNOR U26293 ( .A(b[5258]), .B(n15776), .Z(c[5258]) );
XNOR U26294 ( .A(a[5258]), .B(c5258), .Z(n15776) );
XOR U26295 ( .A(c5259), .B(n15777), .Z(c5260) );
ANDN U26296 ( .B(n15778), .A(n15779), .Z(n15777) );
XOR U26297 ( .A(c5259), .B(b[5259]), .Z(n15778) );
XNOR U26298 ( .A(b[5259]), .B(n15779), .Z(c[5259]) );
XNOR U26299 ( .A(a[5259]), .B(c5259), .Z(n15779) );
XOR U26300 ( .A(c5260), .B(n15780), .Z(c5261) );
ANDN U26301 ( .B(n15781), .A(n15782), .Z(n15780) );
XOR U26302 ( .A(c5260), .B(b[5260]), .Z(n15781) );
XNOR U26303 ( .A(b[5260]), .B(n15782), .Z(c[5260]) );
XNOR U26304 ( .A(a[5260]), .B(c5260), .Z(n15782) );
XOR U26305 ( .A(c5261), .B(n15783), .Z(c5262) );
ANDN U26306 ( .B(n15784), .A(n15785), .Z(n15783) );
XOR U26307 ( .A(c5261), .B(b[5261]), .Z(n15784) );
XNOR U26308 ( .A(b[5261]), .B(n15785), .Z(c[5261]) );
XNOR U26309 ( .A(a[5261]), .B(c5261), .Z(n15785) );
XOR U26310 ( .A(c5262), .B(n15786), .Z(c5263) );
ANDN U26311 ( .B(n15787), .A(n15788), .Z(n15786) );
XOR U26312 ( .A(c5262), .B(b[5262]), .Z(n15787) );
XNOR U26313 ( .A(b[5262]), .B(n15788), .Z(c[5262]) );
XNOR U26314 ( .A(a[5262]), .B(c5262), .Z(n15788) );
XOR U26315 ( .A(c5263), .B(n15789), .Z(c5264) );
ANDN U26316 ( .B(n15790), .A(n15791), .Z(n15789) );
XOR U26317 ( .A(c5263), .B(b[5263]), .Z(n15790) );
XNOR U26318 ( .A(b[5263]), .B(n15791), .Z(c[5263]) );
XNOR U26319 ( .A(a[5263]), .B(c5263), .Z(n15791) );
XOR U26320 ( .A(c5264), .B(n15792), .Z(c5265) );
ANDN U26321 ( .B(n15793), .A(n15794), .Z(n15792) );
XOR U26322 ( .A(c5264), .B(b[5264]), .Z(n15793) );
XNOR U26323 ( .A(b[5264]), .B(n15794), .Z(c[5264]) );
XNOR U26324 ( .A(a[5264]), .B(c5264), .Z(n15794) );
XOR U26325 ( .A(c5265), .B(n15795), .Z(c5266) );
ANDN U26326 ( .B(n15796), .A(n15797), .Z(n15795) );
XOR U26327 ( .A(c5265), .B(b[5265]), .Z(n15796) );
XNOR U26328 ( .A(b[5265]), .B(n15797), .Z(c[5265]) );
XNOR U26329 ( .A(a[5265]), .B(c5265), .Z(n15797) );
XOR U26330 ( .A(c5266), .B(n15798), .Z(c5267) );
ANDN U26331 ( .B(n15799), .A(n15800), .Z(n15798) );
XOR U26332 ( .A(c5266), .B(b[5266]), .Z(n15799) );
XNOR U26333 ( .A(b[5266]), .B(n15800), .Z(c[5266]) );
XNOR U26334 ( .A(a[5266]), .B(c5266), .Z(n15800) );
XOR U26335 ( .A(c5267), .B(n15801), .Z(c5268) );
ANDN U26336 ( .B(n15802), .A(n15803), .Z(n15801) );
XOR U26337 ( .A(c5267), .B(b[5267]), .Z(n15802) );
XNOR U26338 ( .A(b[5267]), .B(n15803), .Z(c[5267]) );
XNOR U26339 ( .A(a[5267]), .B(c5267), .Z(n15803) );
XOR U26340 ( .A(c5268), .B(n15804), .Z(c5269) );
ANDN U26341 ( .B(n15805), .A(n15806), .Z(n15804) );
XOR U26342 ( .A(c5268), .B(b[5268]), .Z(n15805) );
XNOR U26343 ( .A(b[5268]), .B(n15806), .Z(c[5268]) );
XNOR U26344 ( .A(a[5268]), .B(c5268), .Z(n15806) );
XOR U26345 ( .A(c5269), .B(n15807), .Z(c5270) );
ANDN U26346 ( .B(n15808), .A(n15809), .Z(n15807) );
XOR U26347 ( .A(c5269), .B(b[5269]), .Z(n15808) );
XNOR U26348 ( .A(b[5269]), .B(n15809), .Z(c[5269]) );
XNOR U26349 ( .A(a[5269]), .B(c5269), .Z(n15809) );
XOR U26350 ( .A(c5270), .B(n15810), .Z(c5271) );
ANDN U26351 ( .B(n15811), .A(n15812), .Z(n15810) );
XOR U26352 ( .A(c5270), .B(b[5270]), .Z(n15811) );
XNOR U26353 ( .A(b[5270]), .B(n15812), .Z(c[5270]) );
XNOR U26354 ( .A(a[5270]), .B(c5270), .Z(n15812) );
XOR U26355 ( .A(c5271), .B(n15813), .Z(c5272) );
ANDN U26356 ( .B(n15814), .A(n15815), .Z(n15813) );
XOR U26357 ( .A(c5271), .B(b[5271]), .Z(n15814) );
XNOR U26358 ( .A(b[5271]), .B(n15815), .Z(c[5271]) );
XNOR U26359 ( .A(a[5271]), .B(c5271), .Z(n15815) );
XOR U26360 ( .A(c5272), .B(n15816), .Z(c5273) );
ANDN U26361 ( .B(n15817), .A(n15818), .Z(n15816) );
XOR U26362 ( .A(c5272), .B(b[5272]), .Z(n15817) );
XNOR U26363 ( .A(b[5272]), .B(n15818), .Z(c[5272]) );
XNOR U26364 ( .A(a[5272]), .B(c5272), .Z(n15818) );
XOR U26365 ( .A(c5273), .B(n15819), .Z(c5274) );
ANDN U26366 ( .B(n15820), .A(n15821), .Z(n15819) );
XOR U26367 ( .A(c5273), .B(b[5273]), .Z(n15820) );
XNOR U26368 ( .A(b[5273]), .B(n15821), .Z(c[5273]) );
XNOR U26369 ( .A(a[5273]), .B(c5273), .Z(n15821) );
XOR U26370 ( .A(c5274), .B(n15822), .Z(c5275) );
ANDN U26371 ( .B(n15823), .A(n15824), .Z(n15822) );
XOR U26372 ( .A(c5274), .B(b[5274]), .Z(n15823) );
XNOR U26373 ( .A(b[5274]), .B(n15824), .Z(c[5274]) );
XNOR U26374 ( .A(a[5274]), .B(c5274), .Z(n15824) );
XOR U26375 ( .A(c5275), .B(n15825), .Z(c5276) );
ANDN U26376 ( .B(n15826), .A(n15827), .Z(n15825) );
XOR U26377 ( .A(c5275), .B(b[5275]), .Z(n15826) );
XNOR U26378 ( .A(b[5275]), .B(n15827), .Z(c[5275]) );
XNOR U26379 ( .A(a[5275]), .B(c5275), .Z(n15827) );
XOR U26380 ( .A(c5276), .B(n15828), .Z(c5277) );
ANDN U26381 ( .B(n15829), .A(n15830), .Z(n15828) );
XOR U26382 ( .A(c5276), .B(b[5276]), .Z(n15829) );
XNOR U26383 ( .A(b[5276]), .B(n15830), .Z(c[5276]) );
XNOR U26384 ( .A(a[5276]), .B(c5276), .Z(n15830) );
XOR U26385 ( .A(c5277), .B(n15831), .Z(c5278) );
ANDN U26386 ( .B(n15832), .A(n15833), .Z(n15831) );
XOR U26387 ( .A(c5277), .B(b[5277]), .Z(n15832) );
XNOR U26388 ( .A(b[5277]), .B(n15833), .Z(c[5277]) );
XNOR U26389 ( .A(a[5277]), .B(c5277), .Z(n15833) );
XOR U26390 ( .A(c5278), .B(n15834), .Z(c5279) );
ANDN U26391 ( .B(n15835), .A(n15836), .Z(n15834) );
XOR U26392 ( .A(c5278), .B(b[5278]), .Z(n15835) );
XNOR U26393 ( .A(b[5278]), .B(n15836), .Z(c[5278]) );
XNOR U26394 ( .A(a[5278]), .B(c5278), .Z(n15836) );
XOR U26395 ( .A(c5279), .B(n15837), .Z(c5280) );
ANDN U26396 ( .B(n15838), .A(n15839), .Z(n15837) );
XOR U26397 ( .A(c5279), .B(b[5279]), .Z(n15838) );
XNOR U26398 ( .A(b[5279]), .B(n15839), .Z(c[5279]) );
XNOR U26399 ( .A(a[5279]), .B(c5279), .Z(n15839) );
XOR U26400 ( .A(c5280), .B(n15840), .Z(c5281) );
ANDN U26401 ( .B(n15841), .A(n15842), .Z(n15840) );
XOR U26402 ( .A(c5280), .B(b[5280]), .Z(n15841) );
XNOR U26403 ( .A(b[5280]), .B(n15842), .Z(c[5280]) );
XNOR U26404 ( .A(a[5280]), .B(c5280), .Z(n15842) );
XOR U26405 ( .A(c5281), .B(n15843), .Z(c5282) );
ANDN U26406 ( .B(n15844), .A(n15845), .Z(n15843) );
XOR U26407 ( .A(c5281), .B(b[5281]), .Z(n15844) );
XNOR U26408 ( .A(b[5281]), .B(n15845), .Z(c[5281]) );
XNOR U26409 ( .A(a[5281]), .B(c5281), .Z(n15845) );
XOR U26410 ( .A(c5282), .B(n15846), .Z(c5283) );
ANDN U26411 ( .B(n15847), .A(n15848), .Z(n15846) );
XOR U26412 ( .A(c5282), .B(b[5282]), .Z(n15847) );
XNOR U26413 ( .A(b[5282]), .B(n15848), .Z(c[5282]) );
XNOR U26414 ( .A(a[5282]), .B(c5282), .Z(n15848) );
XOR U26415 ( .A(c5283), .B(n15849), .Z(c5284) );
ANDN U26416 ( .B(n15850), .A(n15851), .Z(n15849) );
XOR U26417 ( .A(c5283), .B(b[5283]), .Z(n15850) );
XNOR U26418 ( .A(b[5283]), .B(n15851), .Z(c[5283]) );
XNOR U26419 ( .A(a[5283]), .B(c5283), .Z(n15851) );
XOR U26420 ( .A(c5284), .B(n15852), .Z(c5285) );
ANDN U26421 ( .B(n15853), .A(n15854), .Z(n15852) );
XOR U26422 ( .A(c5284), .B(b[5284]), .Z(n15853) );
XNOR U26423 ( .A(b[5284]), .B(n15854), .Z(c[5284]) );
XNOR U26424 ( .A(a[5284]), .B(c5284), .Z(n15854) );
XOR U26425 ( .A(c5285), .B(n15855), .Z(c5286) );
ANDN U26426 ( .B(n15856), .A(n15857), .Z(n15855) );
XOR U26427 ( .A(c5285), .B(b[5285]), .Z(n15856) );
XNOR U26428 ( .A(b[5285]), .B(n15857), .Z(c[5285]) );
XNOR U26429 ( .A(a[5285]), .B(c5285), .Z(n15857) );
XOR U26430 ( .A(c5286), .B(n15858), .Z(c5287) );
ANDN U26431 ( .B(n15859), .A(n15860), .Z(n15858) );
XOR U26432 ( .A(c5286), .B(b[5286]), .Z(n15859) );
XNOR U26433 ( .A(b[5286]), .B(n15860), .Z(c[5286]) );
XNOR U26434 ( .A(a[5286]), .B(c5286), .Z(n15860) );
XOR U26435 ( .A(c5287), .B(n15861), .Z(c5288) );
ANDN U26436 ( .B(n15862), .A(n15863), .Z(n15861) );
XOR U26437 ( .A(c5287), .B(b[5287]), .Z(n15862) );
XNOR U26438 ( .A(b[5287]), .B(n15863), .Z(c[5287]) );
XNOR U26439 ( .A(a[5287]), .B(c5287), .Z(n15863) );
XOR U26440 ( .A(c5288), .B(n15864), .Z(c5289) );
ANDN U26441 ( .B(n15865), .A(n15866), .Z(n15864) );
XOR U26442 ( .A(c5288), .B(b[5288]), .Z(n15865) );
XNOR U26443 ( .A(b[5288]), .B(n15866), .Z(c[5288]) );
XNOR U26444 ( .A(a[5288]), .B(c5288), .Z(n15866) );
XOR U26445 ( .A(c5289), .B(n15867), .Z(c5290) );
ANDN U26446 ( .B(n15868), .A(n15869), .Z(n15867) );
XOR U26447 ( .A(c5289), .B(b[5289]), .Z(n15868) );
XNOR U26448 ( .A(b[5289]), .B(n15869), .Z(c[5289]) );
XNOR U26449 ( .A(a[5289]), .B(c5289), .Z(n15869) );
XOR U26450 ( .A(c5290), .B(n15870), .Z(c5291) );
ANDN U26451 ( .B(n15871), .A(n15872), .Z(n15870) );
XOR U26452 ( .A(c5290), .B(b[5290]), .Z(n15871) );
XNOR U26453 ( .A(b[5290]), .B(n15872), .Z(c[5290]) );
XNOR U26454 ( .A(a[5290]), .B(c5290), .Z(n15872) );
XOR U26455 ( .A(c5291), .B(n15873), .Z(c5292) );
ANDN U26456 ( .B(n15874), .A(n15875), .Z(n15873) );
XOR U26457 ( .A(c5291), .B(b[5291]), .Z(n15874) );
XNOR U26458 ( .A(b[5291]), .B(n15875), .Z(c[5291]) );
XNOR U26459 ( .A(a[5291]), .B(c5291), .Z(n15875) );
XOR U26460 ( .A(c5292), .B(n15876), .Z(c5293) );
ANDN U26461 ( .B(n15877), .A(n15878), .Z(n15876) );
XOR U26462 ( .A(c5292), .B(b[5292]), .Z(n15877) );
XNOR U26463 ( .A(b[5292]), .B(n15878), .Z(c[5292]) );
XNOR U26464 ( .A(a[5292]), .B(c5292), .Z(n15878) );
XOR U26465 ( .A(c5293), .B(n15879), .Z(c5294) );
ANDN U26466 ( .B(n15880), .A(n15881), .Z(n15879) );
XOR U26467 ( .A(c5293), .B(b[5293]), .Z(n15880) );
XNOR U26468 ( .A(b[5293]), .B(n15881), .Z(c[5293]) );
XNOR U26469 ( .A(a[5293]), .B(c5293), .Z(n15881) );
XOR U26470 ( .A(c5294), .B(n15882), .Z(c5295) );
ANDN U26471 ( .B(n15883), .A(n15884), .Z(n15882) );
XOR U26472 ( .A(c5294), .B(b[5294]), .Z(n15883) );
XNOR U26473 ( .A(b[5294]), .B(n15884), .Z(c[5294]) );
XNOR U26474 ( .A(a[5294]), .B(c5294), .Z(n15884) );
XOR U26475 ( .A(c5295), .B(n15885), .Z(c5296) );
ANDN U26476 ( .B(n15886), .A(n15887), .Z(n15885) );
XOR U26477 ( .A(c5295), .B(b[5295]), .Z(n15886) );
XNOR U26478 ( .A(b[5295]), .B(n15887), .Z(c[5295]) );
XNOR U26479 ( .A(a[5295]), .B(c5295), .Z(n15887) );
XOR U26480 ( .A(c5296), .B(n15888), .Z(c5297) );
ANDN U26481 ( .B(n15889), .A(n15890), .Z(n15888) );
XOR U26482 ( .A(c5296), .B(b[5296]), .Z(n15889) );
XNOR U26483 ( .A(b[5296]), .B(n15890), .Z(c[5296]) );
XNOR U26484 ( .A(a[5296]), .B(c5296), .Z(n15890) );
XOR U26485 ( .A(c5297), .B(n15891), .Z(c5298) );
ANDN U26486 ( .B(n15892), .A(n15893), .Z(n15891) );
XOR U26487 ( .A(c5297), .B(b[5297]), .Z(n15892) );
XNOR U26488 ( .A(b[5297]), .B(n15893), .Z(c[5297]) );
XNOR U26489 ( .A(a[5297]), .B(c5297), .Z(n15893) );
XOR U26490 ( .A(c5298), .B(n15894), .Z(c5299) );
ANDN U26491 ( .B(n15895), .A(n15896), .Z(n15894) );
XOR U26492 ( .A(c5298), .B(b[5298]), .Z(n15895) );
XNOR U26493 ( .A(b[5298]), .B(n15896), .Z(c[5298]) );
XNOR U26494 ( .A(a[5298]), .B(c5298), .Z(n15896) );
XOR U26495 ( .A(c5299), .B(n15897), .Z(c5300) );
ANDN U26496 ( .B(n15898), .A(n15899), .Z(n15897) );
XOR U26497 ( .A(c5299), .B(b[5299]), .Z(n15898) );
XNOR U26498 ( .A(b[5299]), .B(n15899), .Z(c[5299]) );
XNOR U26499 ( .A(a[5299]), .B(c5299), .Z(n15899) );
XOR U26500 ( .A(c5300), .B(n15900), .Z(c5301) );
ANDN U26501 ( .B(n15901), .A(n15902), .Z(n15900) );
XOR U26502 ( .A(c5300), .B(b[5300]), .Z(n15901) );
XNOR U26503 ( .A(b[5300]), .B(n15902), .Z(c[5300]) );
XNOR U26504 ( .A(a[5300]), .B(c5300), .Z(n15902) );
XOR U26505 ( .A(c5301), .B(n15903), .Z(c5302) );
ANDN U26506 ( .B(n15904), .A(n15905), .Z(n15903) );
XOR U26507 ( .A(c5301), .B(b[5301]), .Z(n15904) );
XNOR U26508 ( .A(b[5301]), .B(n15905), .Z(c[5301]) );
XNOR U26509 ( .A(a[5301]), .B(c5301), .Z(n15905) );
XOR U26510 ( .A(c5302), .B(n15906), .Z(c5303) );
ANDN U26511 ( .B(n15907), .A(n15908), .Z(n15906) );
XOR U26512 ( .A(c5302), .B(b[5302]), .Z(n15907) );
XNOR U26513 ( .A(b[5302]), .B(n15908), .Z(c[5302]) );
XNOR U26514 ( .A(a[5302]), .B(c5302), .Z(n15908) );
XOR U26515 ( .A(c5303), .B(n15909), .Z(c5304) );
ANDN U26516 ( .B(n15910), .A(n15911), .Z(n15909) );
XOR U26517 ( .A(c5303), .B(b[5303]), .Z(n15910) );
XNOR U26518 ( .A(b[5303]), .B(n15911), .Z(c[5303]) );
XNOR U26519 ( .A(a[5303]), .B(c5303), .Z(n15911) );
XOR U26520 ( .A(c5304), .B(n15912), .Z(c5305) );
ANDN U26521 ( .B(n15913), .A(n15914), .Z(n15912) );
XOR U26522 ( .A(c5304), .B(b[5304]), .Z(n15913) );
XNOR U26523 ( .A(b[5304]), .B(n15914), .Z(c[5304]) );
XNOR U26524 ( .A(a[5304]), .B(c5304), .Z(n15914) );
XOR U26525 ( .A(c5305), .B(n15915), .Z(c5306) );
ANDN U26526 ( .B(n15916), .A(n15917), .Z(n15915) );
XOR U26527 ( .A(c5305), .B(b[5305]), .Z(n15916) );
XNOR U26528 ( .A(b[5305]), .B(n15917), .Z(c[5305]) );
XNOR U26529 ( .A(a[5305]), .B(c5305), .Z(n15917) );
XOR U26530 ( .A(c5306), .B(n15918), .Z(c5307) );
ANDN U26531 ( .B(n15919), .A(n15920), .Z(n15918) );
XOR U26532 ( .A(c5306), .B(b[5306]), .Z(n15919) );
XNOR U26533 ( .A(b[5306]), .B(n15920), .Z(c[5306]) );
XNOR U26534 ( .A(a[5306]), .B(c5306), .Z(n15920) );
XOR U26535 ( .A(c5307), .B(n15921), .Z(c5308) );
ANDN U26536 ( .B(n15922), .A(n15923), .Z(n15921) );
XOR U26537 ( .A(c5307), .B(b[5307]), .Z(n15922) );
XNOR U26538 ( .A(b[5307]), .B(n15923), .Z(c[5307]) );
XNOR U26539 ( .A(a[5307]), .B(c5307), .Z(n15923) );
XOR U26540 ( .A(c5308), .B(n15924), .Z(c5309) );
ANDN U26541 ( .B(n15925), .A(n15926), .Z(n15924) );
XOR U26542 ( .A(c5308), .B(b[5308]), .Z(n15925) );
XNOR U26543 ( .A(b[5308]), .B(n15926), .Z(c[5308]) );
XNOR U26544 ( .A(a[5308]), .B(c5308), .Z(n15926) );
XOR U26545 ( .A(c5309), .B(n15927), .Z(c5310) );
ANDN U26546 ( .B(n15928), .A(n15929), .Z(n15927) );
XOR U26547 ( .A(c5309), .B(b[5309]), .Z(n15928) );
XNOR U26548 ( .A(b[5309]), .B(n15929), .Z(c[5309]) );
XNOR U26549 ( .A(a[5309]), .B(c5309), .Z(n15929) );
XOR U26550 ( .A(c5310), .B(n15930), .Z(c5311) );
ANDN U26551 ( .B(n15931), .A(n15932), .Z(n15930) );
XOR U26552 ( .A(c5310), .B(b[5310]), .Z(n15931) );
XNOR U26553 ( .A(b[5310]), .B(n15932), .Z(c[5310]) );
XNOR U26554 ( .A(a[5310]), .B(c5310), .Z(n15932) );
XOR U26555 ( .A(c5311), .B(n15933), .Z(c5312) );
ANDN U26556 ( .B(n15934), .A(n15935), .Z(n15933) );
XOR U26557 ( .A(c5311), .B(b[5311]), .Z(n15934) );
XNOR U26558 ( .A(b[5311]), .B(n15935), .Z(c[5311]) );
XNOR U26559 ( .A(a[5311]), .B(c5311), .Z(n15935) );
XOR U26560 ( .A(c5312), .B(n15936), .Z(c5313) );
ANDN U26561 ( .B(n15937), .A(n15938), .Z(n15936) );
XOR U26562 ( .A(c5312), .B(b[5312]), .Z(n15937) );
XNOR U26563 ( .A(b[5312]), .B(n15938), .Z(c[5312]) );
XNOR U26564 ( .A(a[5312]), .B(c5312), .Z(n15938) );
XOR U26565 ( .A(c5313), .B(n15939), .Z(c5314) );
ANDN U26566 ( .B(n15940), .A(n15941), .Z(n15939) );
XOR U26567 ( .A(c5313), .B(b[5313]), .Z(n15940) );
XNOR U26568 ( .A(b[5313]), .B(n15941), .Z(c[5313]) );
XNOR U26569 ( .A(a[5313]), .B(c5313), .Z(n15941) );
XOR U26570 ( .A(c5314), .B(n15942), .Z(c5315) );
ANDN U26571 ( .B(n15943), .A(n15944), .Z(n15942) );
XOR U26572 ( .A(c5314), .B(b[5314]), .Z(n15943) );
XNOR U26573 ( .A(b[5314]), .B(n15944), .Z(c[5314]) );
XNOR U26574 ( .A(a[5314]), .B(c5314), .Z(n15944) );
XOR U26575 ( .A(c5315), .B(n15945), .Z(c5316) );
ANDN U26576 ( .B(n15946), .A(n15947), .Z(n15945) );
XOR U26577 ( .A(c5315), .B(b[5315]), .Z(n15946) );
XNOR U26578 ( .A(b[5315]), .B(n15947), .Z(c[5315]) );
XNOR U26579 ( .A(a[5315]), .B(c5315), .Z(n15947) );
XOR U26580 ( .A(c5316), .B(n15948), .Z(c5317) );
ANDN U26581 ( .B(n15949), .A(n15950), .Z(n15948) );
XOR U26582 ( .A(c5316), .B(b[5316]), .Z(n15949) );
XNOR U26583 ( .A(b[5316]), .B(n15950), .Z(c[5316]) );
XNOR U26584 ( .A(a[5316]), .B(c5316), .Z(n15950) );
XOR U26585 ( .A(c5317), .B(n15951), .Z(c5318) );
ANDN U26586 ( .B(n15952), .A(n15953), .Z(n15951) );
XOR U26587 ( .A(c5317), .B(b[5317]), .Z(n15952) );
XNOR U26588 ( .A(b[5317]), .B(n15953), .Z(c[5317]) );
XNOR U26589 ( .A(a[5317]), .B(c5317), .Z(n15953) );
XOR U26590 ( .A(c5318), .B(n15954), .Z(c5319) );
ANDN U26591 ( .B(n15955), .A(n15956), .Z(n15954) );
XOR U26592 ( .A(c5318), .B(b[5318]), .Z(n15955) );
XNOR U26593 ( .A(b[5318]), .B(n15956), .Z(c[5318]) );
XNOR U26594 ( .A(a[5318]), .B(c5318), .Z(n15956) );
XOR U26595 ( .A(c5319), .B(n15957), .Z(c5320) );
ANDN U26596 ( .B(n15958), .A(n15959), .Z(n15957) );
XOR U26597 ( .A(c5319), .B(b[5319]), .Z(n15958) );
XNOR U26598 ( .A(b[5319]), .B(n15959), .Z(c[5319]) );
XNOR U26599 ( .A(a[5319]), .B(c5319), .Z(n15959) );
XOR U26600 ( .A(c5320), .B(n15960), .Z(c5321) );
ANDN U26601 ( .B(n15961), .A(n15962), .Z(n15960) );
XOR U26602 ( .A(c5320), .B(b[5320]), .Z(n15961) );
XNOR U26603 ( .A(b[5320]), .B(n15962), .Z(c[5320]) );
XNOR U26604 ( .A(a[5320]), .B(c5320), .Z(n15962) );
XOR U26605 ( .A(c5321), .B(n15963), .Z(c5322) );
ANDN U26606 ( .B(n15964), .A(n15965), .Z(n15963) );
XOR U26607 ( .A(c5321), .B(b[5321]), .Z(n15964) );
XNOR U26608 ( .A(b[5321]), .B(n15965), .Z(c[5321]) );
XNOR U26609 ( .A(a[5321]), .B(c5321), .Z(n15965) );
XOR U26610 ( .A(c5322), .B(n15966), .Z(c5323) );
ANDN U26611 ( .B(n15967), .A(n15968), .Z(n15966) );
XOR U26612 ( .A(c5322), .B(b[5322]), .Z(n15967) );
XNOR U26613 ( .A(b[5322]), .B(n15968), .Z(c[5322]) );
XNOR U26614 ( .A(a[5322]), .B(c5322), .Z(n15968) );
XOR U26615 ( .A(c5323), .B(n15969), .Z(c5324) );
ANDN U26616 ( .B(n15970), .A(n15971), .Z(n15969) );
XOR U26617 ( .A(c5323), .B(b[5323]), .Z(n15970) );
XNOR U26618 ( .A(b[5323]), .B(n15971), .Z(c[5323]) );
XNOR U26619 ( .A(a[5323]), .B(c5323), .Z(n15971) );
XOR U26620 ( .A(c5324), .B(n15972), .Z(c5325) );
ANDN U26621 ( .B(n15973), .A(n15974), .Z(n15972) );
XOR U26622 ( .A(c5324), .B(b[5324]), .Z(n15973) );
XNOR U26623 ( .A(b[5324]), .B(n15974), .Z(c[5324]) );
XNOR U26624 ( .A(a[5324]), .B(c5324), .Z(n15974) );
XOR U26625 ( .A(c5325), .B(n15975), .Z(c5326) );
ANDN U26626 ( .B(n15976), .A(n15977), .Z(n15975) );
XOR U26627 ( .A(c5325), .B(b[5325]), .Z(n15976) );
XNOR U26628 ( .A(b[5325]), .B(n15977), .Z(c[5325]) );
XNOR U26629 ( .A(a[5325]), .B(c5325), .Z(n15977) );
XOR U26630 ( .A(c5326), .B(n15978), .Z(c5327) );
ANDN U26631 ( .B(n15979), .A(n15980), .Z(n15978) );
XOR U26632 ( .A(c5326), .B(b[5326]), .Z(n15979) );
XNOR U26633 ( .A(b[5326]), .B(n15980), .Z(c[5326]) );
XNOR U26634 ( .A(a[5326]), .B(c5326), .Z(n15980) );
XOR U26635 ( .A(c5327), .B(n15981), .Z(c5328) );
ANDN U26636 ( .B(n15982), .A(n15983), .Z(n15981) );
XOR U26637 ( .A(c5327), .B(b[5327]), .Z(n15982) );
XNOR U26638 ( .A(b[5327]), .B(n15983), .Z(c[5327]) );
XNOR U26639 ( .A(a[5327]), .B(c5327), .Z(n15983) );
XOR U26640 ( .A(c5328), .B(n15984), .Z(c5329) );
ANDN U26641 ( .B(n15985), .A(n15986), .Z(n15984) );
XOR U26642 ( .A(c5328), .B(b[5328]), .Z(n15985) );
XNOR U26643 ( .A(b[5328]), .B(n15986), .Z(c[5328]) );
XNOR U26644 ( .A(a[5328]), .B(c5328), .Z(n15986) );
XOR U26645 ( .A(c5329), .B(n15987), .Z(c5330) );
ANDN U26646 ( .B(n15988), .A(n15989), .Z(n15987) );
XOR U26647 ( .A(c5329), .B(b[5329]), .Z(n15988) );
XNOR U26648 ( .A(b[5329]), .B(n15989), .Z(c[5329]) );
XNOR U26649 ( .A(a[5329]), .B(c5329), .Z(n15989) );
XOR U26650 ( .A(c5330), .B(n15990), .Z(c5331) );
ANDN U26651 ( .B(n15991), .A(n15992), .Z(n15990) );
XOR U26652 ( .A(c5330), .B(b[5330]), .Z(n15991) );
XNOR U26653 ( .A(b[5330]), .B(n15992), .Z(c[5330]) );
XNOR U26654 ( .A(a[5330]), .B(c5330), .Z(n15992) );
XOR U26655 ( .A(c5331), .B(n15993), .Z(c5332) );
ANDN U26656 ( .B(n15994), .A(n15995), .Z(n15993) );
XOR U26657 ( .A(c5331), .B(b[5331]), .Z(n15994) );
XNOR U26658 ( .A(b[5331]), .B(n15995), .Z(c[5331]) );
XNOR U26659 ( .A(a[5331]), .B(c5331), .Z(n15995) );
XOR U26660 ( .A(c5332), .B(n15996), .Z(c5333) );
ANDN U26661 ( .B(n15997), .A(n15998), .Z(n15996) );
XOR U26662 ( .A(c5332), .B(b[5332]), .Z(n15997) );
XNOR U26663 ( .A(b[5332]), .B(n15998), .Z(c[5332]) );
XNOR U26664 ( .A(a[5332]), .B(c5332), .Z(n15998) );
XOR U26665 ( .A(c5333), .B(n15999), .Z(c5334) );
ANDN U26666 ( .B(n16000), .A(n16001), .Z(n15999) );
XOR U26667 ( .A(c5333), .B(b[5333]), .Z(n16000) );
XNOR U26668 ( .A(b[5333]), .B(n16001), .Z(c[5333]) );
XNOR U26669 ( .A(a[5333]), .B(c5333), .Z(n16001) );
XOR U26670 ( .A(c5334), .B(n16002), .Z(c5335) );
ANDN U26671 ( .B(n16003), .A(n16004), .Z(n16002) );
XOR U26672 ( .A(c5334), .B(b[5334]), .Z(n16003) );
XNOR U26673 ( .A(b[5334]), .B(n16004), .Z(c[5334]) );
XNOR U26674 ( .A(a[5334]), .B(c5334), .Z(n16004) );
XOR U26675 ( .A(c5335), .B(n16005), .Z(c5336) );
ANDN U26676 ( .B(n16006), .A(n16007), .Z(n16005) );
XOR U26677 ( .A(c5335), .B(b[5335]), .Z(n16006) );
XNOR U26678 ( .A(b[5335]), .B(n16007), .Z(c[5335]) );
XNOR U26679 ( .A(a[5335]), .B(c5335), .Z(n16007) );
XOR U26680 ( .A(c5336), .B(n16008), .Z(c5337) );
ANDN U26681 ( .B(n16009), .A(n16010), .Z(n16008) );
XOR U26682 ( .A(c5336), .B(b[5336]), .Z(n16009) );
XNOR U26683 ( .A(b[5336]), .B(n16010), .Z(c[5336]) );
XNOR U26684 ( .A(a[5336]), .B(c5336), .Z(n16010) );
XOR U26685 ( .A(c5337), .B(n16011), .Z(c5338) );
ANDN U26686 ( .B(n16012), .A(n16013), .Z(n16011) );
XOR U26687 ( .A(c5337), .B(b[5337]), .Z(n16012) );
XNOR U26688 ( .A(b[5337]), .B(n16013), .Z(c[5337]) );
XNOR U26689 ( .A(a[5337]), .B(c5337), .Z(n16013) );
XOR U26690 ( .A(c5338), .B(n16014), .Z(c5339) );
ANDN U26691 ( .B(n16015), .A(n16016), .Z(n16014) );
XOR U26692 ( .A(c5338), .B(b[5338]), .Z(n16015) );
XNOR U26693 ( .A(b[5338]), .B(n16016), .Z(c[5338]) );
XNOR U26694 ( .A(a[5338]), .B(c5338), .Z(n16016) );
XOR U26695 ( .A(c5339), .B(n16017), .Z(c5340) );
ANDN U26696 ( .B(n16018), .A(n16019), .Z(n16017) );
XOR U26697 ( .A(c5339), .B(b[5339]), .Z(n16018) );
XNOR U26698 ( .A(b[5339]), .B(n16019), .Z(c[5339]) );
XNOR U26699 ( .A(a[5339]), .B(c5339), .Z(n16019) );
XOR U26700 ( .A(c5340), .B(n16020), .Z(c5341) );
ANDN U26701 ( .B(n16021), .A(n16022), .Z(n16020) );
XOR U26702 ( .A(c5340), .B(b[5340]), .Z(n16021) );
XNOR U26703 ( .A(b[5340]), .B(n16022), .Z(c[5340]) );
XNOR U26704 ( .A(a[5340]), .B(c5340), .Z(n16022) );
XOR U26705 ( .A(c5341), .B(n16023), .Z(c5342) );
ANDN U26706 ( .B(n16024), .A(n16025), .Z(n16023) );
XOR U26707 ( .A(c5341), .B(b[5341]), .Z(n16024) );
XNOR U26708 ( .A(b[5341]), .B(n16025), .Z(c[5341]) );
XNOR U26709 ( .A(a[5341]), .B(c5341), .Z(n16025) );
XOR U26710 ( .A(c5342), .B(n16026), .Z(c5343) );
ANDN U26711 ( .B(n16027), .A(n16028), .Z(n16026) );
XOR U26712 ( .A(c5342), .B(b[5342]), .Z(n16027) );
XNOR U26713 ( .A(b[5342]), .B(n16028), .Z(c[5342]) );
XNOR U26714 ( .A(a[5342]), .B(c5342), .Z(n16028) );
XOR U26715 ( .A(c5343), .B(n16029), .Z(c5344) );
ANDN U26716 ( .B(n16030), .A(n16031), .Z(n16029) );
XOR U26717 ( .A(c5343), .B(b[5343]), .Z(n16030) );
XNOR U26718 ( .A(b[5343]), .B(n16031), .Z(c[5343]) );
XNOR U26719 ( .A(a[5343]), .B(c5343), .Z(n16031) );
XOR U26720 ( .A(c5344), .B(n16032), .Z(c5345) );
ANDN U26721 ( .B(n16033), .A(n16034), .Z(n16032) );
XOR U26722 ( .A(c5344), .B(b[5344]), .Z(n16033) );
XNOR U26723 ( .A(b[5344]), .B(n16034), .Z(c[5344]) );
XNOR U26724 ( .A(a[5344]), .B(c5344), .Z(n16034) );
XOR U26725 ( .A(c5345), .B(n16035), .Z(c5346) );
ANDN U26726 ( .B(n16036), .A(n16037), .Z(n16035) );
XOR U26727 ( .A(c5345), .B(b[5345]), .Z(n16036) );
XNOR U26728 ( .A(b[5345]), .B(n16037), .Z(c[5345]) );
XNOR U26729 ( .A(a[5345]), .B(c5345), .Z(n16037) );
XOR U26730 ( .A(c5346), .B(n16038), .Z(c5347) );
ANDN U26731 ( .B(n16039), .A(n16040), .Z(n16038) );
XOR U26732 ( .A(c5346), .B(b[5346]), .Z(n16039) );
XNOR U26733 ( .A(b[5346]), .B(n16040), .Z(c[5346]) );
XNOR U26734 ( .A(a[5346]), .B(c5346), .Z(n16040) );
XOR U26735 ( .A(c5347), .B(n16041), .Z(c5348) );
ANDN U26736 ( .B(n16042), .A(n16043), .Z(n16041) );
XOR U26737 ( .A(c5347), .B(b[5347]), .Z(n16042) );
XNOR U26738 ( .A(b[5347]), .B(n16043), .Z(c[5347]) );
XNOR U26739 ( .A(a[5347]), .B(c5347), .Z(n16043) );
XOR U26740 ( .A(c5348), .B(n16044), .Z(c5349) );
ANDN U26741 ( .B(n16045), .A(n16046), .Z(n16044) );
XOR U26742 ( .A(c5348), .B(b[5348]), .Z(n16045) );
XNOR U26743 ( .A(b[5348]), .B(n16046), .Z(c[5348]) );
XNOR U26744 ( .A(a[5348]), .B(c5348), .Z(n16046) );
XOR U26745 ( .A(c5349), .B(n16047), .Z(c5350) );
ANDN U26746 ( .B(n16048), .A(n16049), .Z(n16047) );
XOR U26747 ( .A(c5349), .B(b[5349]), .Z(n16048) );
XNOR U26748 ( .A(b[5349]), .B(n16049), .Z(c[5349]) );
XNOR U26749 ( .A(a[5349]), .B(c5349), .Z(n16049) );
XOR U26750 ( .A(c5350), .B(n16050), .Z(c5351) );
ANDN U26751 ( .B(n16051), .A(n16052), .Z(n16050) );
XOR U26752 ( .A(c5350), .B(b[5350]), .Z(n16051) );
XNOR U26753 ( .A(b[5350]), .B(n16052), .Z(c[5350]) );
XNOR U26754 ( .A(a[5350]), .B(c5350), .Z(n16052) );
XOR U26755 ( .A(c5351), .B(n16053), .Z(c5352) );
ANDN U26756 ( .B(n16054), .A(n16055), .Z(n16053) );
XOR U26757 ( .A(c5351), .B(b[5351]), .Z(n16054) );
XNOR U26758 ( .A(b[5351]), .B(n16055), .Z(c[5351]) );
XNOR U26759 ( .A(a[5351]), .B(c5351), .Z(n16055) );
XOR U26760 ( .A(c5352), .B(n16056), .Z(c5353) );
ANDN U26761 ( .B(n16057), .A(n16058), .Z(n16056) );
XOR U26762 ( .A(c5352), .B(b[5352]), .Z(n16057) );
XNOR U26763 ( .A(b[5352]), .B(n16058), .Z(c[5352]) );
XNOR U26764 ( .A(a[5352]), .B(c5352), .Z(n16058) );
XOR U26765 ( .A(c5353), .B(n16059), .Z(c5354) );
ANDN U26766 ( .B(n16060), .A(n16061), .Z(n16059) );
XOR U26767 ( .A(c5353), .B(b[5353]), .Z(n16060) );
XNOR U26768 ( .A(b[5353]), .B(n16061), .Z(c[5353]) );
XNOR U26769 ( .A(a[5353]), .B(c5353), .Z(n16061) );
XOR U26770 ( .A(c5354), .B(n16062), .Z(c5355) );
ANDN U26771 ( .B(n16063), .A(n16064), .Z(n16062) );
XOR U26772 ( .A(c5354), .B(b[5354]), .Z(n16063) );
XNOR U26773 ( .A(b[5354]), .B(n16064), .Z(c[5354]) );
XNOR U26774 ( .A(a[5354]), .B(c5354), .Z(n16064) );
XOR U26775 ( .A(c5355), .B(n16065), .Z(c5356) );
ANDN U26776 ( .B(n16066), .A(n16067), .Z(n16065) );
XOR U26777 ( .A(c5355), .B(b[5355]), .Z(n16066) );
XNOR U26778 ( .A(b[5355]), .B(n16067), .Z(c[5355]) );
XNOR U26779 ( .A(a[5355]), .B(c5355), .Z(n16067) );
XOR U26780 ( .A(c5356), .B(n16068), .Z(c5357) );
ANDN U26781 ( .B(n16069), .A(n16070), .Z(n16068) );
XOR U26782 ( .A(c5356), .B(b[5356]), .Z(n16069) );
XNOR U26783 ( .A(b[5356]), .B(n16070), .Z(c[5356]) );
XNOR U26784 ( .A(a[5356]), .B(c5356), .Z(n16070) );
XOR U26785 ( .A(c5357), .B(n16071), .Z(c5358) );
ANDN U26786 ( .B(n16072), .A(n16073), .Z(n16071) );
XOR U26787 ( .A(c5357), .B(b[5357]), .Z(n16072) );
XNOR U26788 ( .A(b[5357]), .B(n16073), .Z(c[5357]) );
XNOR U26789 ( .A(a[5357]), .B(c5357), .Z(n16073) );
XOR U26790 ( .A(c5358), .B(n16074), .Z(c5359) );
ANDN U26791 ( .B(n16075), .A(n16076), .Z(n16074) );
XOR U26792 ( .A(c5358), .B(b[5358]), .Z(n16075) );
XNOR U26793 ( .A(b[5358]), .B(n16076), .Z(c[5358]) );
XNOR U26794 ( .A(a[5358]), .B(c5358), .Z(n16076) );
XOR U26795 ( .A(c5359), .B(n16077), .Z(c5360) );
ANDN U26796 ( .B(n16078), .A(n16079), .Z(n16077) );
XOR U26797 ( .A(c5359), .B(b[5359]), .Z(n16078) );
XNOR U26798 ( .A(b[5359]), .B(n16079), .Z(c[5359]) );
XNOR U26799 ( .A(a[5359]), .B(c5359), .Z(n16079) );
XOR U26800 ( .A(c5360), .B(n16080), .Z(c5361) );
ANDN U26801 ( .B(n16081), .A(n16082), .Z(n16080) );
XOR U26802 ( .A(c5360), .B(b[5360]), .Z(n16081) );
XNOR U26803 ( .A(b[5360]), .B(n16082), .Z(c[5360]) );
XNOR U26804 ( .A(a[5360]), .B(c5360), .Z(n16082) );
XOR U26805 ( .A(c5361), .B(n16083), .Z(c5362) );
ANDN U26806 ( .B(n16084), .A(n16085), .Z(n16083) );
XOR U26807 ( .A(c5361), .B(b[5361]), .Z(n16084) );
XNOR U26808 ( .A(b[5361]), .B(n16085), .Z(c[5361]) );
XNOR U26809 ( .A(a[5361]), .B(c5361), .Z(n16085) );
XOR U26810 ( .A(c5362), .B(n16086), .Z(c5363) );
ANDN U26811 ( .B(n16087), .A(n16088), .Z(n16086) );
XOR U26812 ( .A(c5362), .B(b[5362]), .Z(n16087) );
XNOR U26813 ( .A(b[5362]), .B(n16088), .Z(c[5362]) );
XNOR U26814 ( .A(a[5362]), .B(c5362), .Z(n16088) );
XOR U26815 ( .A(c5363), .B(n16089), .Z(c5364) );
ANDN U26816 ( .B(n16090), .A(n16091), .Z(n16089) );
XOR U26817 ( .A(c5363), .B(b[5363]), .Z(n16090) );
XNOR U26818 ( .A(b[5363]), .B(n16091), .Z(c[5363]) );
XNOR U26819 ( .A(a[5363]), .B(c5363), .Z(n16091) );
XOR U26820 ( .A(c5364), .B(n16092), .Z(c5365) );
ANDN U26821 ( .B(n16093), .A(n16094), .Z(n16092) );
XOR U26822 ( .A(c5364), .B(b[5364]), .Z(n16093) );
XNOR U26823 ( .A(b[5364]), .B(n16094), .Z(c[5364]) );
XNOR U26824 ( .A(a[5364]), .B(c5364), .Z(n16094) );
XOR U26825 ( .A(c5365), .B(n16095), .Z(c5366) );
ANDN U26826 ( .B(n16096), .A(n16097), .Z(n16095) );
XOR U26827 ( .A(c5365), .B(b[5365]), .Z(n16096) );
XNOR U26828 ( .A(b[5365]), .B(n16097), .Z(c[5365]) );
XNOR U26829 ( .A(a[5365]), .B(c5365), .Z(n16097) );
XOR U26830 ( .A(c5366), .B(n16098), .Z(c5367) );
ANDN U26831 ( .B(n16099), .A(n16100), .Z(n16098) );
XOR U26832 ( .A(c5366), .B(b[5366]), .Z(n16099) );
XNOR U26833 ( .A(b[5366]), .B(n16100), .Z(c[5366]) );
XNOR U26834 ( .A(a[5366]), .B(c5366), .Z(n16100) );
XOR U26835 ( .A(c5367), .B(n16101), .Z(c5368) );
ANDN U26836 ( .B(n16102), .A(n16103), .Z(n16101) );
XOR U26837 ( .A(c5367), .B(b[5367]), .Z(n16102) );
XNOR U26838 ( .A(b[5367]), .B(n16103), .Z(c[5367]) );
XNOR U26839 ( .A(a[5367]), .B(c5367), .Z(n16103) );
XOR U26840 ( .A(c5368), .B(n16104), .Z(c5369) );
ANDN U26841 ( .B(n16105), .A(n16106), .Z(n16104) );
XOR U26842 ( .A(c5368), .B(b[5368]), .Z(n16105) );
XNOR U26843 ( .A(b[5368]), .B(n16106), .Z(c[5368]) );
XNOR U26844 ( .A(a[5368]), .B(c5368), .Z(n16106) );
XOR U26845 ( .A(c5369), .B(n16107), .Z(c5370) );
ANDN U26846 ( .B(n16108), .A(n16109), .Z(n16107) );
XOR U26847 ( .A(c5369), .B(b[5369]), .Z(n16108) );
XNOR U26848 ( .A(b[5369]), .B(n16109), .Z(c[5369]) );
XNOR U26849 ( .A(a[5369]), .B(c5369), .Z(n16109) );
XOR U26850 ( .A(c5370), .B(n16110), .Z(c5371) );
ANDN U26851 ( .B(n16111), .A(n16112), .Z(n16110) );
XOR U26852 ( .A(c5370), .B(b[5370]), .Z(n16111) );
XNOR U26853 ( .A(b[5370]), .B(n16112), .Z(c[5370]) );
XNOR U26854 ( .A(a[5370]), .B(c5370), .Z(n16112) );
XOR U26855 ( .A(c5371), .B(n16113), .Z(c5372) );
ANDN U26856 ( .B(n16114), .A(n16115), .Z(n16113) );
XOR U26857 ( .A(c5371), .B(b[5371]), .Z(n16114) );
XNOR U26858 ( .A(b[5371]), .B(n16115), .Z(c[5371]) );
XNOR U26859 ( .A(a[5371]), .B(c5371), .Z(n16115) );
XOR U26860 ( .A(c5372), .B(n16116), .Z(c5373) );
ANDN U26861 ( .B(n16117), .A(n16118), .Z(n16116) );
XOR U26862 ( .A(c5372), .B(b[5372]), .Z(n16117) );
XNOR U26863 ( .A(b[5372]), .B(n16118), .Z(c[5372]) );
XNOR U26864 ( .A(a[5372]), .B(c5372), .Z(n16118) );
XOR U26865 ( .A(c5373), .B(n16119), .Z(c5374) );
ANDN U26866 ( .B(n16120), .A(n16121), .Z(n16119) );
XOR U26867 ( .A(c5373), .B(b[5373]), .Z(n16120) );
XNOR U26868 ( .A(b[5373]), .B(n16121), .Z(c[5373]) );
XNOR U26869 ( .A(a[5373]), .B(c5373), .Z(n16121) );
XOR U26870 ( .A(c5374), .B(n16122), .Z(c5375) );
ANDN U26871 ( .B(n16123), .A(n16124), .Z(n16122) );
XOR U26872 ( .A(c5374), .B(b[5374]), .Z(n16123) );
XNOR U26873 ( .A(b[5374]), .B(n16124), .Z(c[5374]) );
XNOR U26874 ( .A(a[5374]), .B(c5374), .Z(n16124) );
XOR U26875 ( .A(c5375), .B(n16125), .Z(c5376) );
ANDN U26876 ( .B(n16126), .A(n16127), .Z(n16125) );
XOR U26877 ( .A(c5375), .B(b[5375]), .Z(n16126) );
XNOR U26878 ( .A(b[5375]), .B(n16127), .Z(c[5375]) );
XNOR U26879 ( .A(a[5375]), .B(c5375), .Z(n16127) );
XOR U26880 ( .A(c5376), .B(n16128), .Z(c5377) );
ANDN U26881 ( .B(n16129), .A(n16130), .Z(n16128) );
XOR U26882 ( .A(c5376), .B(b[5376]), .Z(n16129) );
XNOR U26883 ( .A(b[5376]), .B(n16130), .Z(c[5376]) );
XNOR U26884 ( .A(a[5376]), .B(c5376), .Z(n16130) );
XOR U26885 ( .A(c5377), .B(n16131), .Z(c5378) );
ANDN U26886 ( .B(n16132), .A(n16133), .Z(n16131) );
XOR U26887 ( .A(c5377), .B(b[5377]), .Z(n16132) );
XNOR U26888 ( .A(b[5377]), .B(n16133), .Z(c[5377]) );
XNOR U26889 ( .A(a[5377]), .B(c5377), .Z(n16133) );
XOR U26890 ( .A(c5378), .B(n16134), .Z(c5379) );
ANDN U26891 ( .B(n16135), .A(n16136), .Z(n16134) );
XOR U26892 ( .A(c5378), .B(b[5378]), .Z(n16135) );
XNOR U26893 ( .A(b[5378]), .B(n16136), .Z(c[5378]) );
XNOR U26894 ( .A(a[5378]), .B(c5378), .Z(n16136) );
XOR U26895 ( .A(c5379), .B(n16137), .Z(c5380) );
ANDN U26896 ( .B(n16138), .A(n16139), .Z(n16137) );
XOR U26897 ( .A(c5379), .B(b[5379]), .Z(n16138) );
XNOR U26898 ( .A(b[5379]), .B(n16139), .Z(c[5379]) );
XNOR U26899 ( .A(a[5379]), .B(c5379), .Z(n16139) );
XOR U26900 ( .A(c5380), .B(n16140), .Z(c5381) );
ANDN U26901 ( .B(n16141), .A(n16142), .Z(n16140) );
XOR U26902 ( .A(c5380), .B(b[5380]), .Z(n16141) );
XNOR U26903 ( .A(b[5380]), .B(n16142), .Z(c[5380]) );
XNOR U26904 ( .A(a[5380]), .B(c5380), .Z(n16142) );
XOR U26905 ( .A(c5381), .B(n16143), .Z(c5382) );
ANDN U26906 ( .B(n16144), .A(n16145), .Z(n16143) );
XOR U26907 ( .A(c5381), .B(b[5381]), .Z(n16144) );
XNOR U26908 ( .A(b[5381]), .B(n16145), .Z(c[5381]) );
XNOR U26909 ( .A(a[5381]), .B(c5381), .Z(n16145) );
XOR U26910 ( .A(c5382), .B(n16146), .Z(c5383) );
ANDN U26911 ( .B(n16147), .A(n16148), .Z(n16146) );
XOR U26912 ( .A(c5382), .B(b[5382]), .Z(n16147) );
XNOR U26913 ( .A(b[5382]), .B(n16148), .Z(c[5382]) );
XNOR U26914 ( .A(a[5382]), .B(c5382), .Z(n16148) );
XOR U26915 ( .A(c5383), .B(n16149), .Z(c5384) );
ANDN U26916 ( .B(n16150), .A(n16151), .Z(n16149) );
XOR U26917 ( .A(c5383), .B(b[5383]), .Z(n16150) );
XNOR U26918 ( .A(b[5383]), .B(n16151), .Z(c[5383]) );
XNOR U26919 ( .A(a[5383]), .B(c5383), .Z(n16151) );
XOR U26920 ( .A(c5384), .B(n16152), .Z(c5385) );
ANDN U26921 ( .B(n16153), .A(n16154), .Z(n16152) );
XOR U26922 ( .A(c5384), .B(b[5384]), .Z(n16153) );
XNOR U26923 ( .A(b[5384]), .B(n16154), .Z(c[5384]) );
XNOR U26924 ( .A(a[5384]), .B(c5384), .Z(n16154) );
XOR U26925 ( .A(c5385), .B(n16155), .Z(c5386) );
ANDN U26926 ( .B(n16156), .A(n16157), .Z(n16155) );
XOR U26927 ( .A(c5385), .B(b[5385]), .Z(n16156) );
XNOR U26928 ( .A(b[5385]), .B(n16157), .Z(c[5385]) );
XNOR U26929 ( .A(a[5385]), .B(c5385), .Z(n16157) );
XOR U26930 ( .A(c5386), .B(n16158), .Z(c5387) );
ANDN U26931 ( .B(n16159), .A(n16160), .Z(n16158) );
XOR U26932 ( .A(c5386), .B(b[5386]), .Z(n16159) );
XNOR U26933 ( .A(b[5386]), .B(n16160), .Z(c[5386]) );
XNOR U26934 ( .A(a[5386]), .B(c5386), .Z(n16160) );
XOR U26935 ( .A(c5387), .B(n16161), .Z(c5388) );
ANDN U26936 ( .B(n16162), .A(n16163), .Z(n16161) );
XOR U26937 ( .A(c5387), .B(b[5387]), .Z(n16162) );
XNOR U26938 ( .A(b[5387]), .B(n16163), .Z(c[5387]) );
XNOR U26939 ( .A(a[5387]), .B(c5387), .Z(n16163) );
XOR U26940 ( .A(c5388), .B(n16164), .Z(c5389) );
ANDN U26941 ( .B(n16165), .A(n16166), .Z(n16164) );
XOR U26942 ( .A(c5388), .B(b[5388]), .Z(n16165) );
XNOR U26943 ( .A(b[5388]), .B(n16166), .Z(c[5388]) );
XNOR U26944 ( .A(a[5388]), .B(c5388), .Z(n16166) );
XOR U26945 ( .A(c5389), .B(n16167), .Z(c5390) );
ANDN U26946 ( .B(n16168), .A(n16169), .Z(n16167) );
XOR U26947 ( .A(c5389), .B(b[5389]), .Z(n16168) );
XNOR U26948 ( .A(b[5389]), .B(n16169), .Z(c[5389]) );
XNOR U26949 ( .A(a[5389]), .B(c5389), .Z(n16169) );
XOR U26950 ( .A(c5390), .B(n16170), .Z(c5391) );
ANDN U26951 ( .B(n16171), .A(n16172), .Z(n16170) );
XOR U26952 ( .A(c5390), .B(b[5390]), .Z(n16171) );
XNOR U26953 ( .A(b[5390]), .B(n16172), .Z(c[5390]) );
XNOR U26954 ( .A(a[5390]), .B(c5390), .Z(n16172) );
XOR U26955 ( .A(c5391), .B(n16173), .Z(c5392) );
ANDN U26956 ( .B(n16174), .A(n16175), .Z(n16173) );
XOR U26957 ( .A(c5391), .B(b[5391]), .Z(n16174) );
XNOR U26958 ( .A(b[5391]), .B(n16175), .Z(c[5391]) );
XNOR U26959 ( .A(a[5391]), .B(c5391), .Z(n16175) );
XOR U26960 ( .A(c5392), .B(n16176), .Z(c5393) );
ANDN U26961 ( .B(n16177), .A(n16178), .Z(n16176) );
XOR U26962 ( .A(c5392), .B(b[5392]), .Z(n16177) );
XNOR U26963 ( .A(b[5392]), .B(n16178), .Z(c[5392]) );
XNOR U26964 ( .A(a[5392]), .B(c5392), .Z(n16178) );
XOR U26965 ( .A(c5393), .B(n16179), .Z(c5394) );
ANDN U26966 ( .B(n16180), .A(n16181), .Z(n16179) );
XOR U26967 ( .A(c5393), .B(b[5393]), .Z(n16180) );
XNOR U26968 ( .A(b[5393]), .B(n16181), .Z(c[5393]) );
XNOR U26969 ( .A(a[5393]), .B(c5393), .Z(n16181) );
XOR U26970 ( .A(c5394), .B(n16182), .Z(c5395) );
ANDN U26971 ( .B(n16183), .A(n16184), .Z(n16182) );
XOR U26972 ( .A(c5394), .B(b[5394]), .Z(n16183) );
XNOR U26973 ( .A(b[5394]), .B(n16184), .Z(c[5394]) );
XNOR U26974 ( .A(a[5394]), .B(c5394), .Z(n16184) );
XOR U26975 ( .A(c5395), .B(n16185), .Z(c5396) );
ANDN U26976 ( .B(n16186), .A(n16187), .Z(n16185) );
XOR U26977 ( .A(c5395), .B(b[5395]), .Z(n16186) );
XNOR U26978 ( .A(b[5395]), .B(n16187), .Z(c[5395]) );
XNOR U26979 ( .A(a[5395]), .B(c5395), .Z(n16187) );
XOR U26980 ( .A(c5396), .B(n16188), .Z(c5397) );
ANDN U26981 ( .B(n16189), .A(n16190), .Z(n16188) );
XOR U26982 ( .A(c5396), .B(b[5396]), .Z(n16189) );
XNOR U26983 ( .A(b[5396]), .B(n16190), .Z(c[5396]) );
XNOR U26984 ( .A(a[5396]), .B(c5396), .Z(n16190) );
XOR U26985 ( .A(c5397), .B(n16191), .Z(c5398) );
ANDN U26986 ( .B(n16192), .A(n16193), .Z(n16191) );
XOR U26987 ( .A(c5397), .B(b[5397]), .Z(n16192) );
XNOR U26988 ( .A(b[5397]), .B(n16193), .Z(c[5397]) );
XNOR U26989 ( .A(a[5397]), .B(c5397), .Z(n16193) );
XOR U26990 ( .A(c5398), .B(n16194), .Z(c5399) );
ANDN U26991 ( .B(n16195), .A(n16196), .Z(n16194) );
XOR U26992 ( .A(c5398), .B(b[5398]), .Z(n16195) );
XNOR U26993 ( .A(b[5398]), .B(n16196), .Z(c[5398]) );
XNOR U26994 ( .A(a[5398]), .B(c5398), .Z(n16196) );
XOR U26995 ( .A(c5399), .B(n16197), .Z(c5400) );
ANDN U26996 ( .B(n16198), .A(n16199), .Z(n16197) );
XOR U26997 ( .A(c5399), .B(b[5399]), .Z(n16198) );
XNOR U26998 ( .A(b[5399]), .B(n16199), .Z(c[5399]) );
XNOR U26999 ( .A(a[5399]), .B(c5399), .Z(n16199) );
XOR U27000 ( .A(c5400), .B(n16200), .Z(c5401) );
ANDN U27001 ( .B(n16201), .A(n16202), .Z(n16200) );
XOR U27002 ( .A(c5400), .B(b[5400]), .Z(n16201) );
XNOR U27003 ( .A(b[5400]), .B(n16202), .Z(c[5400]) );
XNOR U27004 ( .A(a[5400]), .B(c5400), .Z(n16202) );
XOR U27005 ( .A(c5401), .B(n16203), .Z(c5402) );
ANDN U27006 ( .B(n16204), .A(n16205), .Z(n16203) );
XOR U27007 ( .A(c5401), .B(b[5401]), .Z(n16204) );
XNOR U27008 ( .A(b[5401]), .B(n16205), .Z(c[5401]) );
XNOR U27009 ( .A(a[5401]), .B(c5401), .Z(n16205) );
XOR U27010 ( .A(c5402), .B(n16206), .Z(c5403) );
ANDN U27011 ( .B(n16207), .A(n16208), .Z(n16206) );
XOR U27012 ( .A(c5402), .B(b[5402]), .Z(n16207) );
XNOR U27013 ( .A(b[5402]), .B(n16208), .Z(c[5402]) );
XNOR U27014 ( .A(a[5402]), .B(c5402), .Z(n16208) );
XOR U27015 ( .A(c5403), .B(n16209), .Z(c5404) );
ANDN U27016 ( .B(n16210), .A(n16211), .Z(n16209) );
XOR U27017 ( .A(c5403), .B(b[5403]), .Z(n16210) );
XNOR U27018 ( .A(b[5403]), .B(n16211), .Z(c[5403]) );
XNOR U27019 ( .A(a[5403]), .B(c5403), .Z(n16211) );
XOR U27020 ( .A(c5404), .B(n16212), .Z(c5405) );
ANDN U27021 ( .B(n16213), .A(n16214), .Z(n16212) );
XOR U27022 ( .A(c5404), .B(b[5404]), .Z(n16213) );
XNOR U27023 ( .A(b[5404]), .B(n16214), .Z(c[5404]) );
XNOR U27024 ( .A(a[5404]), .B(c5404), .Z(n16214) );
XOR U27025 ( .A(c5405), .B(n16215), .Z(c5406) );
ANDN U27026 ( .B(n16216), .A(n16217), .Z(n16215) );
XOR U27027 ( .A(c5405), .B(b[5405]), .Z(n16216) );
XNOR U27028 ( .A(b[5405]), .B(n16217), .Z(c[5405]) );
XNOR U27029 ( .A(a[5405]), .B(c5405), .Z(n16217) );
XOR U27030 ( .A(c5406), .B(n16218), .Z(c5407) );
ANDN U27031 ( .B(n16219), .A(n16220), .Z(n16218) );
XOR U27032 ( .A(c5406), .B(b[5406]), .Z(n16219) );
XNOR U27033 ( .A(b[5406]), .B(n16220), .Z(c[5406]) );
XNOR U27034 ( .A(a[5406]), .B(c5406), .Z(n16220) );
XOR U27035 ( .A(c5407), .B(n16221), .Z(c5408) );
ANDN U27036 ( .B(n16222), .A(n16223), .Z(n16221) );
XOR U27037 ( .A(c5407), .B(b[5407]), .Z(n16222) );
XNOR U27038 ( .A(b[5407]), .B(n16223), .Z(c[5407]) );
XNOR U27039 ( .A(a[5407]), .B(c5407), .Z(n16223) );
XOR U27040 ( .A(c5408), .B(n16224), .Z(c5409) );
ANDN U27041 ( .B(n16225), .A(n16226), .Z(n16224) );
XOR U27042 ( .A(c5408), .B(b[5408]), .Z(n16225) );
XNOR U27043 ( .A(b[5408]), .B(n16226), .Z(c[5408]) );
XNOR U27044 ( .A(a[5408]), .B(c5408), .Z(n16226) );
XOR U27045 ( .A(c5409), .B(n16227), .Z(c5410) );
ANDN U27046 ( .B(n16228), .A(n16229), .Z(n16227) );
XOR U27047 ( .A(c5409), .B(b[5409]), .Z(n16228) );
XNOR U27048 ( .A(b[5409]), .B(n16229), .Z(c[5409]) );
XNOR U27049 ( .A(a[5409]), .B(c5409), .Z(n16229) );
XOR U27050 ( .A(c5410), .B(n16230), .Z(c5411) );
ANDN U27051 ( .B(n16231), .A(n16232), .Z(n16230) );
XOR U27052 ( .A(c5410), .B(b[5410]), .Z(n16231) );
XNOR U27053 ( .A(b[5410]), .B(n16232), .Z(c[5410]) );
XNOR U27054 ( .A(a[5410]), .B(c5410), .Z(n16232) );
XOR U27055 ( .A(c5411), .B(n16233), .Z(c5412) );
ANDN U27056 ( .B(n16234), .A(n16235), .Z(n16233) );
XOR U27057 ( .A(c5411), .B(b[5411]), .Z(n16234) );
XNOR U27058 ( .A(b[5411]), .B(n16235), .Z(c[5411]) );
XNOR U27059 ( .A(a[5411]), .B(c5411), .Z(n16235) );
XOR U27060 ( .A(c5412), .B(n16236), .Z(c5413) );
ANDN U27061 ( .B(n16237), .A(n16238), .Z(n16236) );
XOR U27062 ( .A(c5412), .B(b[5412]), .Z(n16237) );
XNOR U27063 ( .A(b[5412]), .B(n16238), .Z(c[5412]) );
XNOR U27064 ( .A(a[5412]), .B(c5412), .Z(n16238) );
XOR U27065 ( .A(c5413), .B(n16239), .Z(c5414) );
ANDN U27066 ( .B(n16240), .A(n16241), .Z(n16239) );
XOR U27067 ( .A(c5413), .B(b[5413]), .Z(n16240) );
XNOR U27068 ( .A(b[5413]), .B(n16241), .Z(c[5413]) );
XNOR U27069 ( .A(a[5413]), .B(c5413), .Z(n16241) );
XOR U27070 ( .A(c5414), .B(n16242), .Z(c5415) );
ANDN U27071 ( .B(n16243), .A(n16244), .Z(n16242) );
XOR U27072 ( .A(c5414), .B(b[5414]), .Z(n16243) );
XNOR U27073 ( .A(b[5414]), .B(n16244), .Z(c[5414]) );
XNOR U27074 ( .A(a[5414]), .B(c5414), .Z(n16244) );
XOR U27075 ( .A(c5415), .B(n16245), .Z(c5416) );
ANDN U27076 ( .B(n16246), .A(n16247), .Z(n16245) );
XOR U27077 ( .A(c5415), .B(b[5415]), .Z(n16246) );
XNOR U27078 ( .A(b[5415]), .B(n16247), .Z(c[5415]) );
XNOR U27079 ( .A(a[5415]), .B(c5415), .Z(n16247) );
XOR U27080 ( .A(c5416), .B(n16248), .Z(c5417) );
ANDN U27081 ( .B(n16249), .A(n16250), .Z(n16248) );
XOR U27082 ( .A(c5416), .B(b[5416]), .Z(n16249) );
XNOR U27083 ( .A(b[5416]), .B(n16250), .Z(c[5416]) );
XNOR U27084 ( .A(a[5416]), .B(c5416), .Z(n16250) );
XOR U27085 ( .A(c5417), .B(n16251), .Z(c5418) );
ANDN U27086 ( .B(n16252), .A(n16253), .Z(n16251) );
XOR U27087 ( .A(c5417), .B(b[5417]), .Z(n16252) );
XNOR U27088 ( .A(b[5417]), .B(n16253), .Z(c[5417]) );
XNOR U27089 ( .A(a[5417]), .B(c5417), .Z(n16253) );
XOR U27090 ( .A(c5418), .B(n16254), .Z(c5419) );
ANDN U27091 ( .B(n16255), .A(n16256), .Z(n16254) );
XOR U27092 ( .A(c5418), .B(b[5418]), .Z(n16255) );
XNOR U27093 ( .A(b[5418]), .B(n16256), .Z(c[5418]) );
XNOR U27094 ( .A(a[5418]), .B(c5418), .Z(n16256) );
XOR U27095 ( .A(c5419), .B(n16257), .Z(c5420) );
ANDN U27096 ( .B(n16258), .A(n16259), .Z(n16257) );
XOR U27097 ( .A(c5419), .B(b[5419]), .Z(n16258) );
XNOR U27098 ( .A(b[5419]), .B(n16259), .Z(c[5419]) );
XNOR U27099 ( .A(a[5419]), .B(c5419), .Z(n16259) );
XOR U27100 ( .A(c5420), .B(n16260), .Z(c5421) );
ANDN U27101 ( .B(n16261), .A(n16262), .Z(n16260) );
XOR U27102 ( .A(c5420), .B(b[5420]), .Z(n16261) );
XNOR U27103 ( .A(b[5420]), .B(n16262), .Z(c[5420]) );
XNOR U27104 ( .A(a[5420]), .B(c5420), .Z(n16262) );
XOR U27105 ( .A(c5421), .B(n16263), .Z(c5422) );
ANDN U27106 ( .B(n16264), .A(n16265), .Z(n16263) );
XOR U27107 ( .A(c5421), .B(b[5421]), .Z(n16264) );
XNOR U27108 ( .A(b[5421]), .B(n16265), .Z(c[5421]) );
XNOR U27109 ( .A(a[5421]), .B(c5421), .Z(n16265) );
XOR U27110 ( .A(c5422), .B(n16266), .Z(c5423) );
ANDN U27111 ( .B(n16267), .A(n16268), .Z(n16266) );
XOR U27112 ( .A(c5422), .B(b[5422]), .Z(n16267) );
XNOR U27113 ( .A(b[5422]), .B(n16268), .Z(c[5422]) );
XNOR U27114 ( .A(a[5422]), .B(c5422), .Z(n16268) );
XOR U27115 ( .A(c5423), .B(n16269), .Z(c5424) );
ANDN U27116 ( .B(n16270), .A(n16271), .Z(n16269) );
XOR U27117 ( .A(c5423), .B(b[5423]), .Z(n16270) );
XNOR U27118 ( .A(b[5423]), .B(n16271), .Z(c[5423]) );
XNOR U27119 ( .A(a[5423]), .B(c5423), .Z(n16271) );
XOR U27120 ( .A(c5424), .B(n16272), .Z(c5425) );
ANDN U27121 ( .B(n16273), .A(n16274), .Z(n16272) );
XOR U27122 ( .A(c5424), .B(b[5424]), .Z(n16273) );
XNOR U27123 ( .A(b[5424]), .B(n16274), .Z(c[5424]) );
XNOR U27124 ( .A(a[5424]), .B(c5424), .Z(n16274) );
XOR U27125 ( .A(c5425), .B(n16275), .Z(c5426) );
ANDN U27126 ( .B(n16276), .A(n16277), .Z(n16275) );
XOR U27127 ( .A(c5425), .B(b[5425]), .Z(n16276) );
XNOR U27128 ( .A(b[5425]), .B(n16277), .Z(c[5425]) );
XNOR U27129 ( .A(a[5425]), .B(c5425), .Z(n16277) );
XOR U27130 ( .A(c5426), .B(n16278), .Z(c5427) );
ANDN U27131 ( .B(n16279), .A(n16280), .Z(n16278) );
XOR U27132 ( .A(c5426), .B(b[5426]), .Z(n16279) );
XNOR U27133 ( .A(b[5426]), .B(n16280), .Z(c[5426]) );
XNOR U27134 ( .A(a[5426]), .B(c5426), .Z(n16280) );
XOR U27135 ( .A(c5427), .B(n16281), .Z(c5428) );
ANDN U27136 ( .B(n16282), .A(n16283), .Z(n16281) );
XOR U27137 ( .A(c5427), .B(b[5427]), .Z(n16282) );
XNOR U27138 ( .A(b[5427]), .B(n16283), .Z(c[5427]) );
XNOR U27139 ( .A(a[5427]), .B(c5427), .Z(n16283) );
XOR U27140 ( .A(c5428), .B(n16284), .Z(c5429) );
ANDN U27141 ( .B(n16285), .A(n16286), .Z(n16284) );
XOR U27142 ( .A(c5428), .B(b[5428]), .Z(n16285) );
XNOR U27143 ( .A(b[5428]), .B(n16286), .Z(c[5428]) );
XNOR U27144 ( .A(a[5428]), .B(c5428), .Z(n16286) );
XOR U27145 ( .A(c5429), .B(n16287), .Z(c5430) );
ANDN U27146 ( .B(n16288), .A(n16289), .Z(n16287) );
XOR U27147 ( .A(c5429), .B(b[5429]), .Z(n16288) );
XNOR U27148 ( .A(b[5429]), .B(n16289), .Z(c[5429]) );
XNOR U27149 ( .A(a[5429]), .B(c5429), .Z(n16289) );
XOR U27150 ( .A(c5430), .B(n16290), .Z(c5431) );
ANDN U27151 ( .B(n16291), .A(n16292), .Z(n16290) );
XOR U27152 ( .A(c5430), .B(b[5430]), .Z(n16291) );
XNOR U27153 ( .A(b[5430]), .B(n16292), .Z(c[5430]) );
XNOR U27154 ( .A(a[5430]), .B(c5430), .Z(n16292) );
XOR U27155 ( .A(c5431), .B(n16293), .Z(c5432) );
ANDN U27156 ( .B(n16294), .A(n16295), .Z(n16293) );
XOR U27157 ( .A(c5431), .B(b[5431]), .Z(n16294) );
XNOR U27158 ( .A(b[5431]), .B(n16295), .Z(c[5431]) );
XNOR U27159 ( .A(a[5431]), .B(c5431), .Z(n16295) );
XOR U27160 ( .A(c5432), .B(n16296), .Z(c5433) );
ANDN U27161 ( .B(n16297), .A(n16298), .Z(n16296) );
XOR U27162 ( .A(c5432), .B(b[5432]), .Z(n16297) );
XNOR U27163 ( .A(b[5432]), .B(n16298), .Z(c[5432]) );
XNOR U27164 ( .A(a[5432]), .B(c5432), .Z(n16298) );
XOR U27165 ( .A(c5433), .B(n16299), .Z(c5434) );
ANDN U27166 ( .B(n16300), .A(n16301), .Z(n16299) );
XOR U27167 ( .A(c5433), .B(b[5433]), .Z(n16300) );
XNOR U27168 ( .A(b[5433]), .B(n16301), .Z(c[5433]) );
XNOR U27169 ( .A(a[5433]), .B(c5433), .Z(n16301) );
XOR U27170 ( .A(c5434), .B(n16302), .Z(c5435) );
ANDN U27171 ( .B(n16303), .A(n16304), .Z(n16302) );
XOR U27172 ( .A(c5434), .B(b[5434]), .Z(n16303) );
XNOR U27173 ( .A(b[5434]), .B(n16304), .Z(c[5434]) );
XNOR U27174 ( .A(a[5434]), .B(c5434), .Z(n16304) );
XOR U27175 ( .A(c5435), .B(n16305), .Z(c5436) );
ANDN U27176 ( .B(n16306), .A(n16307), .Z(n16305) );
XOR U27177 ( .A(c5435), .B(b[5435]), .Z(n16306) );
XNOR U27178 ( .A(b[5435]), .B(n16307), .Z(c[5435]) );
XNOR U27179 ( .A(a[5435]), .B(c5435), .Z(n16307) );
XOR U27180 ( .A(c5436), .B(n16308), .Z(c5437) );
ANDN U27181 ( .B(n16309), .A(n16310), .Z(n16308) );
XOR U27182 ( .A(c5436), .B(b[5436]), .Z(n16309) );
XNOR U27183 ( .A(b[5436]), .B(n16310), .Z(c[5436]) );
XNOR U27184 ( .A(a[5436]), .B(c5436), .Z(n16310) );
XOR U27185 ( .A(c5437), .B(n16311), .Z(c5438) );
ANDN U27186 ( .B(n16312), .A(n16313), .Z(n16311) );
XOR U27187 ( .A(c5437), .B(b[5437]), .Z(n16312) );
XNOR U27188 ( .A(b[5437]), .B(n16313), .Z(c[5437]) );
XNOR U27189 ( .A(a[5437]), .B(c5437), .Z(n16313) );
XOR U27190 ( .A(c5438), .B(n16314), .Z(c5439) );
ANDN U27191 ( .B(n16315), .A(n16316), .Z(n16314) );
XOR U27192 ( .A(c5438), .B(b[5438]), .Z(n16315) );
XNOR U27193 ( .A(b[5438]), .B(n16316), .Z(c[5438]) );
XNOR U27194 ( .A(a[5438]), .B(c5438), .Z(n16316) );
XOR U27195 ( .A(c5439), .B(n16317), .Z(c5440) );
ANDN U27196 ( .B(n16318), .A(n16319), .Z(n16317) );
XOR U27197 ( .A(c5439), .B(b[5439]), .Z(n16318) );
XNOR U27198 ( .A(b[5439]), .B(n16319), .Z(c[5439]) );
XNOR U27199 ( .A(a[5439]), .B(c5439), .Z(n16319) );
XOR U27200 ( .A(c5440), .B(n16320), .Z(c5441) );
ANDN U27201 ( .B(n16321), .A(n16322), .Z(n16320) );
XOR U27202 ( .A(c5440), .B(b[5440]), .Z(n16321) );
XNOR U27203 ( .A(b[5440]), .B(n16322), .Z(c[5440]) );
XNOR U27204 ( .A(a[5440]), .B(c5440), .Z(n16322) );
XOR U27205 ( .A(c5441), .B(n16323), .Z(c5442) );
ANDN U27206 ( .B(n16324), .A(n16325), .Z(n16323) );
XOR U27207 ( .A(c5441), .B(b[5441]), .Z(n16324) );
XNOR U27208 ( .A(b[5441]), .B(n16325), .Z(c[5441]) );
XNOR U27209 ( .A(a[5441]), .B(c5441), .Z(n16325) );
XOR U27210 ( .A(c5442), .B(n16326), .Z(c5443) );
ANDN U27211 ( .B(n16327), .A(n16328), .Z(n16326) );
XOR U27212 ( .A(c5442), .B(b[5442]), .Z(n16327) );
XNOR U27213 ( .A(b[5442]), .B(n16328), .Z(c[5442]) );
XNOR U27214 ( .A(a[5442]), .B(c5442), .Z(n16328) );
XOR U27215 ( .A(c5443), .B(n16329), .Z(c5444) );
ANDN U27216 ( .B(n16330), .A(n16331), .Z(n16329) );
XOR U27217 ( .A(c5443), .B(b[5443]), .Z(n16330) );
XNOR U27218 ( .A(b[5443]), .B(n16331), .Z(c[5443]) );
XNOR U27219 ( .A(a[5443]), .B(c5443), .Z(n16331) );
XOR U27220 ( .A(c5444), .B(n16332), .Z(c5445) );
ANDN U27221 ( .B(n16333), .A(n16334), .Z(n16332) );
XOR U27222 ( .A(c5444), .B(b[5444]), .Z(n16333) );
XNOR U27223 ( .A(b[5444]), .B(n16334), .Z(c[5444]) );
XNOR U27224 ( .A(a[5444]), .B(c5444), .Z(n16334) );
XOR U27225 ( .A(c5445), .B(n16335), .Z(c5446) );
ANDN U27226 ( .B(n16336), .A(n16337), .Z(n16335) );
XOR U27227 ( .A(c5445), .B(b[5445]), .Z(n16336) );
XNOR U27228 ( .A(b[5445]), .B(n16337), .Z(c[5445]) );
XNOR U27229 ( .A(a[5445]), .B(c5445), .Z(n16337) );
XOR U27230 ( .A(c5446), .B(n16338), .Z(c5447) );
ANDN U27231 ( .B(n16339), .A(n16340), .Z(n16338) );
XOR U27232 ( .A(c5446), .B(b[5446]), .Z(n16339) );
XNOR U27233 ( .A(b[5446]), .B(n16340), .Z(c[5446]) );
XNOR U27234 ( .A(a[5446]), .B(c5446), .Z(n16340) );
XOR U27235 ( .A(c5447), .B(n16341), .Z(c5448) );
ANDN U27236 ( .B(n16342), .A(n16343), .Z(n16341) );
XOR U27237 ( .A(c5447), .B(b[5447]), .Z(n16342) );
XNOR U27238 ( .A(b[5447]), .B(n16343), .Z(c[5447]) );
XNOR U27239 ( .A(a[5447]), .B(c5447), .Z(n16343) );
XOR U27240 ( .A(c5448), .B(n16344), .Z(c5449) );
ANDN U27241 ( .B(n16345), .A(n16346), .Z(n16344) );
XOR U27242 ( .A(c5448), .B(b[5448]), .Z(n16345) );
XNOR U27243 ( .A(b[5448]), .B(n16346), .Z(c[5448]) );
XNOR U27244 ( .A(a[5448]), .B(c5448), .Z(n16346) );
XOR U27245 ( .A(c5449), .B(n16347), .Z(c5450) );
ANDN U27246 ( .B(n16348), .A(n16349), .Z(n16347) );
XOR U27247 ( .A(c5449), .B(b[5449]), .Z(n16348) );
XNOR U27248 ( .A(b[5449]), .B(n16349), .Z(c[5449]) );
XNOR U27249 ( .A(a[5449]), .B(c5449), .Z(n16349) );
XOR U27250 ( .A(c5450), .B(n16350), .Z(c5451) );
ANDN U27251 ( .B(n16351), .A(n16352), .Z(n16350) );
XOR U27252 ( .A(c5450), .B(b[5450]), .Z(n16351) );
XNOR U27253 ( .A(b[5450]), .B(n16352), .Z(c[5450]) );
XNOR U27254 ( .A(a[5450]), .B(c5450), .Z(n16352) );
XOR U27255 ( .A(c5451), .B(n16353), .Z(c5452) );
ANDN U27256 ( .B(n16354), .A(n16355), .Z(n16353) );
XOR U27257 ( .A(c5451), .B(b[5451]), .Z(n16354) );
XNOR U27258 ( .A(b[5451]), .B(n16355), .Z(c[5451]) );
XNOR U27259 ( .A(a[5451]), .B(c5451), .Z(n16355) );
XOR U27260 ( .A(c5452), .B(n16356), .Z(c5453) );
ANDN U27261 ( .B(n16357), .A(n16358), .Z(n16356) );
XOR U27262 ( .A(c5452), .B(b[5452]), .Z(n16357) );
XNOR U27263 ( .A(b[5452]), .B(n16358), .Z(c[5452]) );
XNOR U27264 ( .A(a[5452]), .B(c5452), .Z(n16358) );
XOR U27265 ( .A(c5453), .B(n16359), .Z(c5454) );
ANDN U27266 ( .B(n16360), .A(n16361), .Z(n16359) );
XOR U27267 ( .A(c5453), .B(b[5453]), .Z(n16360) );
XNOR U27268 ( .A(b[5453]), .B(n16361), .Z(c[5453]) );
XNOR U27269 ( .A(a[5453]), .B(c5453), .Z(n16361) );
XOR U27270 ( .A(c5454), .B(n16362), .Z(c5455) );
ANDN U27271 ( .B(n16363), .A(n16364), .Z(n16362) );
XOR U27272 ( .A(c5454), .B(b[5454]), .Z(n16363) );
XNOR U27273 ( .A(b[5454]), .B(n16364), .Z(c[5454]) );
XNOR U27274 ( .A(a[5454]), .B(c5454), .Z(n16364) );
XOR U27275 ( .A(c5455), .B(n16365), .Z(c5456) );
ANDN U27276 ( .B(n16366), .A(n16367), .Z(n16365) );
XOR U27277 ( .A(c5455), .B(b[5455]), .Z(n16366) );
XNOR U27278 ( .A(b[5455]), .B(n16367), .Z(c[5455]) );
XNOR U27279 ( .A(a[5455]), .B(c5455), .Z(n16367) );
XOR U27280 ( .A(c5456), .B(n16368), .Z(c5457) );
ANDN U27281 ( .B(n16369), .A(n16370), .Z(n16368) );
XOR U27282 ( .A(c5456), .B(b[5456]), .Z(n16369) );
XNOR U27283 ( .A(b[5456]), .B(n16370), .Z(c[5456]) );
XNOR U27284 ( .A(a[5456]), .B(c5456), .Z(n16370) );
XOR U27285 ( .A(c5457), .B(n16371), .Z(c5458) );
ANDN U27286 ( .B(n16372), .A(n16373), .Z(n16371) );
XOR U27287 ( .A(c5457), .B(b[5457]), .Z(n16372) );
XNOR U27288 ( .A(b[5457]), .B(n16373), .Z(c[5457]) );
XNOR U27289 ( .A(a[5457]), .B(c5457), .Z(n16373) );
XOR U27290 ( .A(c5458), .B(n16374), .Z(c5459) );
ANDN U27291 ( .B(n16375), .A(n16376), .Z(n16374) );
XOR U27292 ( .A(c5458), .B(b[5458]), .Z(n16375) );
XNOR U27293 ( .A(b[5458]), .B(n16376), .Z(c[5458]) );
XNOR U27294 ( .A(a[5458]), .B(c5458), .Z(n16376) );
XOR U27295 ( .A(c5459), .B(n16377), .Z(c5460) );
ANDN U27296 ( .B(n16378), .A(n16379), .Z(n16377) );
XOR U27297 ( .A(c5459), .B(b[5459]), .Z(n16378) );
XNOR U27298 ( .A(b[5459]), .B(n16379), .Z(c[5459]) );
XNOR U27299 ( .A(a[5459]), .B(c5459), .Z(n16379) );
XOR U27300 ( .A(c5460), .B(n16380), .Z(c5461) );
ANDN U27301 ( .B(n16381), .A(n16382), .Z(n16380) );
XOR U27302 ( .A(c5460), .B(b[5460]), .Z(n16381) );
XNOR U27303 ( .A(b[5460]), .B(n16382), .Z(c[5460]) );
XNOR U27304 ( .A(a[5460]), .B(c5460), .Z(n16382) );
XOR U27305 ( .A(c5461), .B(n16383), .Z(c5462) );
ANDN U27306 ( .B(n16384), .A(n16385), .Z(n16383) );
XOR U27307 ( .A(c5461), .B(b[5461]), .Z(n16384) );
XNOR U27308 ( .A(b[5461]), .B(n16385), .Z(c[5461]) );
XNOR U27309 ( .A(a[5461]), .B(c5461), .Z(n16385) );
XOR U27310 ( .A(c5462), .B(n16386), .Z(c5463) );
ANDN U27311 ( .B(n16387), .A(n16388), .Z(n16386) );
XOR U27312 ( .A(c5462), .B(b[5462]), .Z(n16387) );
XNOR U27313 ( .A(b[5462]), .B(n16388), .Z(c[5462]) );
XNOR U27314 ( .A(a[5462]), .B(c5462), .Z(n16388) );
XOR U27315 ( .A(c5463), .B(n16389), .Z(c5464) );
ANDN U27316 ( .B(n16390), .A(n16391), .Z(n16389) );
XOR U27317 ( .A(c5463), .B(b[5463]), .Z(n16390) );
XNOR U27318 ( .A(b[5463]), .B(n16391), .Z(c[5463]) );
XNOR U27319 ( .A(a[5463]), .B(c5463), .Z(n16391) );
XOR U27320 ( .A(c5464), .B(n16392), .Z(c5465) );
ANDN U27321 ( .B(n16393), .A(n16394), .Z(n16392) );
XOR U27322 ( .A(c5464), .B(b[5464]), .Z(n16393) );
XNOR U27323 ( .A(b[5464]), .B(n16394), .Z(c[5464]) );
XNOR U27324 ( .A(a[5464]), .B(c5464), .Z(n16394) );
XOR U27325 ( .A(c5465), .B(n16395), .Z(c5466) );
ANDN U27326 ( .B(n16396), .A(n16397), .Z(n16395) );
XOR U27327 ( .A(c5465), .B(b[5465]), .Z(n16396) );
XNOR U27328 ( .A(b[5465]), .B(n16397), .Z(c[5465]) );
XNOR U27329 ( .A(a[5465]), .B(c5465), .Z(n16397) );
XOR U27330 ( .A(c5466), .B(n16398), .Z(c5467) );
ANDN U27331 ( .B(n16399), .A(n16400), .Z(n16398) );
XOR U27332 ( .A(c5466), .B(b[5466]), .Z(n16399) );
XNOR U27333 ( .A(b[5466]), .B(n16400), .Z(c[5466]) );
XNOR U27334 ( .A(a[5466]), .B(c5466), .Z(n16400) );
XOR U27335 ( .A(c5467), .B(n16401), .Z(c5468) );
ANDN U27336 ( .B(n16402), .A(n16403), .Z(n16401) );
XOR U27337 ( .A(c5467), .B(b[5467]), .Z(n16402) );
XNOR U27338 ( .A(b[5467]), .B(n16403), .Z(c[5467]) );
XNOR U27339 ( .A(a[5467]), .B(c5467), .Z(n16403) );
XOR U27340 ( .A(c5468), .B(n16404), .Z(c5469) );
ANDN U27341 ( .B(n16405), .A(n16406), .Z(n16404) );
XOR U27342 ( .A(c5468), .B(b[5468]), .Z(n16405) );
XNOR U27343 ( .A(b[5468]), .B(n16406), .Z(c[5468]) );
XNOR U27344 ( .A(a[5468]), .B(c5468), .Z(n16406) );
XOR U27345 ( .A(c5469), .B(n16407), .Z(c5470) );
ANDN U27346 ( .B(n16408), .A(n16409), .Z(n16407) );
XOR U27347 ( .A(c5469), .B(b[5469]), .Z(n16408) );
XNOR U27348 ( .A(b[5469]), .B(n16409), .Z(c[5469]) );
XNOR U27349 ( .A(a[5469]), .B(c5469), .Z(n16409) );
XOR U27350 ( .A(c5470), .B(n16410), .Z(c5471) );
ANDN U27351 ( .B(n16411), .A(n16412), .Z(n16410) );
XOR U27352 ( .A(c5470), .B(b[5470]), .Z(n16411) );
XNOR U27353 ( .A(b[5470]), .B(n16412), .Z(c[5470]) );
XNOR U27354 ( .A(a[5470]), .B(c5470), .Z(n16412) );
XOR U27355 ( .A(c5471), .B(n16413), .Z(c5472) );
ANDN U27356 ( .B(n16414), .A(n16415), .Z(n16413) );
XOR U27357 ( .A(c5471), .B(b[5471]), .Z(n16414) );
XNOR U27358 ( .A(b[5471]), .B(n16415), .Z(c[5471]) );
XNOR U27359 ( .A(a[5471]), .B(c5471), .Z(n16415) );
XOR U27360 ( .A(c5472), .B(n16416), .Z(c5473) );
ANDN U27361 ( .B(n16417), .A(n16418), .Z(n16416) );
XOR U27362 ( .A(c5472), .B(b[5472]), .Z(n16417) );
XNOR U27363 ( .A(b[5472]), .B(n16418), .Z(c[5472]) );
XNOR U27364 ( .A(a[5472]), .B(c5472), .Z(n16418) );
XOR U27365 ( .A(c5473), .B(n16419), .Z(c5474) );
ANDN U27366 ( .B(n16420), .A(n16421), .Z(n16419) );
XOR U27367 ( .A(c5473), .B(b[5473]), .Z(n16420) );
XNOR U27368 ( .A(b[5473]), .B(n16421), .Z(c[5473]) );
XNOR U27369 ( .A(a[5473]), .B(c5473), .Z(n16421) );
XOR U27370 ( .A(c5474), .B(n16422), .Z(c5475) );
ANDN U27371 ( .B(n16423), .A(n16424), .Z(n16422) );
XOR U27372 ( .A(c5474), .B(b[5474]), .Z(n16423) );
XNOR U27373 ( .A(b[5474]), .B(n16424), .Z(c[5474]) );
XNOR U27374 ( .A(a[5474]), .B(c5474), .Z(n16424) );
XOR U27375 ( .A(c5475), .B(n16425), .Z(c5476) );
ANDN U27376 ( .B(n16426), .A(n16427), .Z(n16425) );
XOR U27377 ( .A(c5475), .B(b[5475]), .Z(n16426) );
XNOR U27378 ( .A(b[5475]), .B(n16427), .Z(c[5475]) );
XNOR U27379 ( .A(a[5475]), .B(c5475), .Z(n16427) );
XOR U27380 ( .A(c5476), .B(n16428), .Z(c5477) );
ANDN U27381 ( .B(n16429), .A(n16430), .Z(n16428) );
XOR U27382 ( .A(c5476), .B(b[5476]), .Z(n16429) );
XNOR U27383 ( .A(b[5476]), .B(n16430), .Z(c[5476]) );
XNOR U27384 ( .A(a[5476]), .B(c5476), .Z(n16430) );
XOR U27385 ( .A(c5477), .B(n16431), .Z(c5478) );
ANDN U27386 ( .B(n16432), .A(n16433), .Z(n16431) );
XOR U27387 ( .A(c5477), .B(b[5477]), .Z(n16432) );
XNOR U27388 ( .A(b[5477]), .B(n16433), .Z(c[5477]) );
XNOR U27389 ( .A(a[5477]), .B(c5477), .Z(n16433) );
XOR U27390 ( .A(c5478), .B(n16434), .Z(c5479) );
ANDN U27391 ( .B(n16435), .A(n16436), .Z(n16434) );
XOR U27392 ( .A(c5478), .B(b[5478]), .Z(n16435) );
XNOR U27393 ( .A(b[5478]), .B(n16436), .Z(c[5478]) );
XNOR U27394 ( .A(a[5478]), .B(c5478), .Z(n16436) );
XOR U27395 ( .A(c5479), .B(n16437), .Z(c5480) );
ANDN U27396 ( .B(n16438), .A(n16439), .Z(n16437) );
XOR U27397 ( .A(c5479), .B(b[5479]), .Z(n16438) );
XNOR U27398 ( .A(b[5479]), .B(n16439), .Z(c[5479]) );
XNOR U27399 ( .A(a[5479]), .B(c5479), .Z(n16439) );
XOR U27400 ( .A(c5480), .B(n16440), .Z(c5481) );
ANDN U27401 ( .B(n16441), .A(n16442), .Z(n16440) );
XOR U27402 ( .A(c5480), .B(b[5480]), .Z(n16441) );
XNOR U27403 ( .A(b[5480]), .B(n16442), .Z(c[5480]) );
XNOR U27404 ( .A(a[5480]), .B(c5480), .Z(n16442) );
XOR U27405 ( .A(c5481), .B(n16443), .Z(c5482) );
ANDN U27406 ( .B(n16444), .A(n16445), .Z(n16443) );
XOR U27407 ( .A(c5481), .B(b[5481]), .Z(n16444) );
XNOR U27408 ( .A(b[5481]), .B(n16445), .Z(c[5481]) );
XNOR U27409 ( .A(a[5481]), .B(c5481), .Z(n16445) );
XOR U27410 ( .A(c5482), .B(n16446), .Z(c5483) );
ANDN U27411 ( .B(n16447), .A(n16448), .Z(n16446) );
XOR U27412 ( .A(c5482), .B(b[5482]), .Z(n16447) );
XNOR U27413 ( .A(b[5482]), .B(n16448), .Z(c[5482]) );
XNOR U27414 ( .A(a[5482]), .B(c5482), .Z(n16448) );
XOR U27415 ( .A(c5483), .B(n16449), .Z(c5484) );
ANDN U27416 ( .B(n16450), .A(n16451), .Z(n16449) );
XOR U27417 ( .A(c5483), .B(b[5483]), .Z(n16450) );
XNOR U27418 ( .A(b[5483]), .B(n16451), .Z(c[5483]) );
XNOR U27419 ( .A(a[5483]), .B(c5483), .Z(n16451) );
XOR U27420 ( .A(c5484), .B(n16452), .Z(c5485) );
ANDN U27421 ( .B(n16453), .A(n16454), .Z(n16452) );
XOR U27422 ( .A(c5484), .B(b[5484]), .Z(n16453) );
XNOR U27423 ( .A(b[5484]), .B(n16454), .Z(c[5484]) );
XNOR U27424 ( .A(a[5484]), .B(c5484), .Z(n16454) );
XOR U27425 ( .A(c5485), .B(n16455), .Z(c5486) );
ANDN U27426 ( .B(n16456), .A(n16457), .Z(n16455) );
XOR U27427 ( .A(c5485), .B(b[5485]), .Z(n16456) );
XNOR U27428 ( .A(b[5485]), .B(n16457), .Z(c[5485]) );
XNOR U27429 ( .A(a[5485]), .B(c5485), .Z(n16457) );
XOR U27430 ( .A(c5486), .B(n16458), .Z(c5487) );
ANDN U27431 ( .B(n16459), .A(n16460), .Z(n16458) );
XOR U27432 ( .A(c5486), .B(b[5486]), .Z(n16459) );
XNOR U27433 ( .A(b[5486]), .B(n16460), .Z(c[5486]) );
XNOR U27434 ( .A(a[5486]), .B(c5486), .Z(n16460) );
XOR U27435 ( .A(c5487), .B(n16461), .Z(c5488) );
ANDN U27436 ( .B(n16462), .A(n16463), .Z(n16461) );
XOR U27437 ( .A(c5487), .B(b[5487]), .Z(n16462) );
XNOR U27438 ( .A(b[5487]), .B(n16463), .Z(c[5487]) );
XNOR U27439 ( .A(a[5487]), .B(c5487), .Z(n16463) );
XOR U27440 ( .A(c5488), .B(n16464), .Z(c5489) );
ANDN U27441 ( .B(n16465), .A(n16466), .Z(n16464) );
XOR U27442 ( .A(c5488), .B(b[5488]), .Z(n16465) );
XNOR U27443 ( .A(b[5488]), .B(n16466), .Z(c[5488]) );
XNOR U27444 ( .A(a[5488]), .B(c5488), .Z(n16466) );
XOR U27445 ( .A(c5489), .B(n16467), .Z(c5490) );
ANDN U27446 ( .B(n16468), .A(n16469), .Z(n16467) );
XOR U27447 ( .A(c5489), .B(b[5489]), .Z(n16468) );
XNOR U27448 ( .A(b[5489]), .B(n16469), .Z(c[5489]) );
XNOR U27449 ( .A(a[5489]), .B(c5489), .Z(n16469) );
XOR U27450 ( .A(c5490), .B(n16470), .Z(c5491) );
ANDN U27451 ( .B(n16471), .A(n16472), .Z(n16470) );
XOR U27452 ( .A(c5490), .B(b[5490]), .Z(n16471) );
XNOR U27453 ( .A(b[5490]), .B(n16472), .Z(c[5490]) );
XNOR U27454 ( .A(a[5490]), .B(c5490), .Z(n16472) );
XOR U27455 ( .A(c5491), .B(n16473), .Z(c5492) );
ANDN U27456 ( .B(n16474), .A(n16475), .Z(n16473) );
XOR U27457 ( .A(c5491), .B(b[5491]), .Z(n16474) );
XNOR U27458 ( .A(b[5491]), .B(n16475), .Z(c[5491]) );
XNOR U27459 ( .A(a[5491]), .B(c5491), .Z(n16475) );
XOR U27460 ( .A(c5492), .B(n16476), .Z(c5493) );
ANDN U27461 ( .B(n16477), .A(n16478), .Z(n16476) );
XOR U27462 ( .A(c5492), .B(b[5492]), .Z(n16477) );
XNOR U27463 ( .A(b[5492]), .B(n16478), .Z(c[5492]) );
XNOR U27464 ( .A(a[5492]), .B(c5492), .Z(n16478) );
XOR U27465 ( .A(c5493), .B(n16479), .Z(c5494) );
ANDN U27466 ( .B(n16480), .A(n16481), .Z(n16479) );
XOR U27467 ( .A(c5493), .B(b[5493]), .Z(n16480) );
XNOR U27468 ( .A(b[5493]), .B(n16481), .Z(c[5493]) );
XNOR U27469 ( .A(a[5493]), .B(c5493), .Z(n16481) );
XOR U27470 ( .A(c5494), .B(n16482), .Z(c5495) );
ANDN U27471 ( .B(n16483), .A(n16484), .Z(n16482) );
XOR U27472 ( .A(c5494), .B(b[5494]), .Z(n16483) );
XNOR U27473 ( .A(b[5494]), .B(n16484), .Z(c[5494]) );
XNOR U27474 ( .A(a[5494]), .B(c5494), .Z(n16484) );
XOR U27475 ( .A(c5495), .B(n16485), .Z(c5496) );
ANDN U27476 ( .B(n16486), .A(n16487), .Z(n16485) );
XOR U27477 ( .A(c5495), .B(b[5495]), .Z(n16486) );
XNOR U27478 ( .A(b[5495]), .B(n16487), .Z(c[5495]) );
XNOR U27479 ( .A(a[5495]), .B(c5495), .Z(n16487) );
XOR U27480 ( .A(c5496), .B(n16488), .Z(c5497) );
ANDN U27481 ( .B(n16489), .A(n16490), .Z(n16488) );
XOR U27482 ( .A(c5496), .B(b[5496]), .Z(n16489) );
XNOR U27483 ( .A(b[5496]), .B(n16490), .Z(c[5496]) );
XNOR U27484 ( .A(a[5496]), .B(c5496), .Z(n16490) );
XOR U27485 ( .A(c5497), .B(n16491), .Z(c5498) );
ANDN U27486 ( .B(n16492), .A(n16493), .Z(n16491) );
XOR U27487 ( .A(c5497), .B(b[5497]), .Z(n16492) );
XNOR U27488 ( .A(b[5497]), .B(n16493), .Z(c[5497]) );
XNOR U27489 ( .A(a[5497]), .B(c5497), .Z(n16493) );
XOR U27490 ( .A(c5498), .B(n16494), .Z(c5499) );
ANDN U27491 ( .B(n16495), .A(n16496), .Z(n16494) );
XOR U27492 ( .A(c5498), .B(b[5498]), .Z(n16495) );
XNOR U27493 ( .A(b[5498]), .B(n16496), .Z(c[5498]) );
XNOR U27494 ( .A(a[5498]), .B(c5498), .Z(n16496) );
XOR U27495 ( .A(c5499), .B(n16497), .Z(c5500) );
ANDN U27496 ( .B(n16498), .A(n16499), .Z(n16497) );
XOR U27497 ( .A(c5499), .B(b[5499]), .Z(n16498) );
XNOR U27498 ( .A(b[5499]), .B(n16499), .Z(c[5499]) );
XNOR U27499 ( .A(a[5499]), .B(c5499), .Z(n16499) );
XOR U27500 ( .A(c5500), .B(n16500), .Z(c5501) );
ANDN U27501 ( .B(n16501), .A(n16502), .Z(n16500) );
XOR U27502 ( .A(c5500), .B(b[5500]), .Z(n16501) );
XNOR U27503 ( .A(b[5500]), .B(n16502), .Z(c[5500]) );
XNOR U27504 ( .A(a[5500]), .B(c5500), .Z(n16502) );
XOR U27505 ( .A(c5501), .B(n16503), .Z(c5502) );
ANDN U27506 ( .B(n16504), .A(n16505), .Z(n16503) );
XOR U27507 ( .A(c5501), .B(b[5501]), .Z(n16504) );
XNOR U27508 ( .A(b[5501]), .B(n16505), .Z(c[5501]) );
XNOR U27509 ( .A(a[5501]), .B(c5501), .Z(n16505) );
XOR U27510 ( .A(c5502), .B(n16506), .Z(c5503) );
ANDN U27511 ( .B(n16507), .A(n16508), .Z(n16506) );
XOR U27512 ( .A(c5502), .B(b[5502]), .Z(n16507) );
XNOR U27513 ( .A(b[5502]), .B(n16508), .Z(c[5502]) );
XNOR U27514 ( .A(a[5502]), .B(c5502), .Z(n16508) );
XOR U27515 ( .A(c5503), .B(n16509), .Z(c5504) );
ANDN U27516 ( .B(n16510), .A(n16511), .Z(n16509) );
XOR U27517 ( .A(c5503), .B(b[5503]), .Z(n16510) );
XNOR U27518 ( .A(b[5503]), .B(n16511), .Z(c[5503]) );
XNOR U27519 ( .A(a[5503]), .B(c5503), .Z(n16511) );
XOR U27520 ( .A(c5504), .B(n16512), .Z(c5505) );
ANDN U27521 ( .B(n16513), .A(n16514), .Z(n16512) );
XOR U27522 ( .A(c5504), .B(b[5504]), .Z(n16513) );
XNOR U27523 ( .A(b[5504]), .B(n16514), .Z(c[5504]) );
XNOR U27524 ( .A(a[5504]), .B(c5504), .Z(n16514) );
XOR U27525 ( .A(c5505), .B(n16515), .Z(c5506) );
ANDN U27526 ( .B(n16516), .A(n16517), .Z(n16515) );
XOR U27527 ( .A(c5505), .B(b[5505]), .Z(n16516) );
XNOR U27528 ( .A(b[5505]), .B(n16517), .Z(c[5505]) );
XNOR U27529 ( .A(a[5505]), .B(c5505), .Z(n16517) );
XOR U27530 ( .A(c5506), .B(n16518), .Z(c5507) );
ANDN U27531 ( .B(n16519), .A(n16520), .Z(n16518) );
XOR U27532 ( .A(c5506), .B(b[5506]), .Z(n16519) );
XNOR U27533 ( .A(b[5506]), .B(n16520), .Z(c[5506]) );
XNOR U27534 ( .A(a[5506]), .B(c5506), .Z(n16520) );
XOR U27535 ( .A(c5507), .B(n16521), .Z(c5508) );
ANDN U27536 ( .B(n16522), .A(n16523), .Z(n16521) );
XOR U27537 ( .A(c5507), .B(b[5507]), .Z(n16522) );
XNOR U27538 ( .A(b[5507]), .B(n16523), .Z(c[5507]) );
XNOR U27539 ( .A(a[5507]), .B(c5507), .Z(n16523) );
XOR U27540 ( .A(c5508), .B(n16524), .Z(c5509) );
ANDN U27541 ( .B(n16525), .A(n16526), .Z(n16524) );
XOR U27542 ( .A(c5508), .B(b[5508]), .Z(n16525) );
XNOR U27543 ( .A(b[5508]), .B(n16526), .Z(c[5508]) );
XNOR U27544 ( .A(a[5508]), .B(c5508), .Z(n16526) );
XOR U27545 ( .A(c5509), .B(n16527), .Z(c5510) );
ANDN U27546 ( .B(n16528), .A(n16529), .Z(n16527) );
XOR U27547 ( .A(c5509), .B(b[5509]), .Z(n16528) );
XNOR U27548 ( .A(b[5509]), .B(n16529), .Z(c[5509]) );
XNOR U27549 ( .A(a[5509]), .B(c5509), .Z(n16529) );
XOR U27550 ( .A(c5510), .B(n16530), .Z(c5511) );
ANDN U27551 ( .B(n16531), .A(n16532), .Z(n16530) );
XOR U27552 ( .A(c5510), .B(b[5510]), .Z(n16531) );
XNOR U27553 ( .A(b[5510]), .B(n16532), .Z(c[5510]) );
XNOR U27554 ( .A(a[5510]), .B(c5510), .Z(n16532) );
XOR U27555 ( .A(c5511), .B(n16533), .Z(c5512) );
ANDN U27556 ( .B(n16534), .A(n16535), .Z(n16533) );
XOR U27557 ( .A(c5511), .B(b[5511]), .Z(n16534) );
XNOR U27558 ( .A(b[5511]), .B(n16535), .Z(c[5511]) );
XNOR U27559 ( .A(a[5511]), .B(c5511), .Z(n16535) );
XOR U27560 ( .A(c5512), .B(n16536), .Z(c5513) );
ANDN U27561 ( .B(n16537), .A(n16538), .Z(n16536) );
XOR U27562 ( .A(c5512), .B(b[5512]), .Z(n16537) );
XNOR U27563 ( .A(b[5512]), .B(n16538), .Z(c[5512]) );
XNOR U27564 ( .A(a[5512]), .B(c5512), .Z(n16538) );
XOR U27565 ( .A(c5513), .B(n16539), .Z(c5514) );
ANDN U27566 ( .B(n16540), .A(n16541), .Z(n16539) );
XOR U27567 ( .A(c5513), .B(b[5513]), .Z(n16540) );
XNOR U27568 ( .A(b[5513]), .B(n16541), .Z(c[5513]) );
XNOR U27569 ( .A(a[5513]), .B(c5513), .Z(n16541) );
XOR U27570 ( .A(c5514), .B(n16542), .Z(c5515) );
ANDN U27571 ( .B(n16543), .A(n16544), .Z(n16542) );
XOR U27572 ( .A(c5514), .B(b[5514]), .Z(n16543) );
XNOR U27573 ( .A(b[5514]), .B(n16544), .Z(c[5514]) );
XNOR U27574 ( .A(a[5514]), .B(c5514), .Z(n16544) );
XOR U27575 ( .A(c5515), .B(n16545), .Z(c5516) );
ANDN U27576 ( .B(n16546), .A(n16547), .Z(n16545) );
XOR U27577 ( .A(c5515), .B(b[5515]), .Z(n16546) );
XNOR U27578 ( .A(b[5515]), .B(n16547), .Z(c[5515]) );
XNOR U27579 ( .A(a[5515]), .B(c5515), .Z(n16547) );
XOR U27580 ( .A(c5516), .B(n16548), .Z(c5517) );
ANDN U27581 ( .B(n16549), .A(n16550), .Z(n16548) );
XOR U27582 ( .A(c5516), .B(b[5516]), .Z(n16549) );
XNOR U27583 ( .A(b[5516]), .B(n16550), .Z(c[5516]) );
XNOR U27584 ( .A(a[5516]), .B(c5516), .Z(n16550) );
XOR U27585 ( .A(c5517), .B(n16551), .Z(c5518) );
ANDN U27586 ( .B(n16552), .A(n16553), .Z(n16551) );
XOR U27587 ( .A(c5517), .B(b[5517]), .Z(n16552) );
XNOR U27588 ( .A(b[5517]), .B(n16553), .Z(c[5517]) );
XNOR U27589 ( .A(a[5517]), .B(c5517), .Z(n16553) );
XOR U27590 ( .A(c5518), .B(n16554), .Z(c5519) );
ANDN U27591 ( .B(n16555), .A(n16556), .Z(n16554) );
XOR U27592 ( .A(c5518), .B(b[5518]), .Z(n16555) );
XNOR U27593 ( .A(b[5518]), .B(n16556), .Z(c[5518]) );
XNOR U27594 ( .A(a[5518]), .B(c5518), .Z(n16556) );
XOR U27595 ( .A(c5519), .B(n16557), .Z(c5520) );
ANDN U27596 ( .B(n16558), .A(n16559), .Z(n16557) );
XOR U27597 ( .A(c5519), .B(b[5519]), .Z(n16558) );
XNOR U27598 ( .A(b[5519]), .B(n16559), .Z(c[5519]) );
XNOR U27599 ( .A(a[5519]), .B(c5519), .Z(n16559) );
XOR U27600 ( .A(c5520), .B(n16560), .Z(c5521) );
ANDN U27601 ( .B(n16561), .A(n16562), .Z(n16560) );
XOR U27602 ( .A(c5520), .B(b[5520]), .Z(n16561) );
XNOR U27603 ( .A(b[5520]), .B(n16562), .Z(c[5520]) );
XNOR U27604 ( .A(a[5520]), .B(c5520), .Z(n16562) );
XOR U27605 ( .A(c5521), .B(n16563), .Z(c5522) );
ANDN U27606 ( .B(n16564), .A(n16565), .Z(n16563) );
XOR U27607 ( .A(c5521), .B(b[5521]), .Z(n16564) );
XNOR U27608 ( .A(b[5521]), .B(n16565), .Z(c[5521]) );
XNOR U27609 ( .A(a[5521]), .B(c5521), .Z(n16565) );
XOR U27610 ( .A(c5522), .B(n16566), .Z(c5523) );
ANDN U27611 ( .B(n16567), .A(n16568), .Z(n16566) );
XOR U27612 ( .A(c5522), .B(b[5522]), .Z(n16567) );
XNOR U27613 ( .A(b[5522]), .B(n16568), .Z(c[5522]) );
XNOR U27614 ( .A(a[5522]), .B(c5522), .Z(n16568) );
XOR U27615 ( .A(c5523), .B(n16569), .Z(c5524) );
ANDN U27616 ( .B(n16570), .A(n16571), .Z(n16569) );
XOR U27617 ( .A(c5523), .B(b[5523]), .Z(n16570) );
XNOR U27618 ( .A(b[5523]), .B(n16571), .Z(c[5523]) );
XNOR U27619 ( .A(a[5523]), .B(c5523), .Z(n16571) );
XOR U27620 ( .A(c5524), .B(n16572), .Z(c5525) );
ANDN U27621 ( .B(n16573), .A(n16574), .Z(n16572) );
XOR U27622 ( .A(c5524), .B(b[5524]), .Z(n16573) );
XNOR U27623 ( .A(b[5524]), .B(n16574), .Z(c[5524]) );
XNOR U27624 ( .A(a[5524]), .B(c5524), .Z(n16574) );
XOR U27625 ( .A(c5525), .B(n16575), .Z(c5526) );
ANDN U27626 ( .B(n16576), .A(n16577), .Z(n16575) );
XOR U27627 ( .A(c5525), .B(b[5525]), .Z(n16576) );
XNOR U27628 ( .A(b[5525]), .B(n16577), .Z(c[5525]) );
XNOR U27629 ( .A(a[5525]), .B(c5525), .Z(n16577) );
XOR U27630 ( .A(c5526), .B(n16578), .Z(c5527) );
ANDN U27631 ( .B(n16579), .A(n16580), .Z(n16578) );
XOR U27632 ( .A(c5526), .B(b[5526]), .Z(n16579) );
XNOR U27633 ( .A(b[5526]), .B(n16580), .Z(c[5526]) );
XNOR U27634 ( .A(a[5526]), .B(c5526), .Z(n16580) );
XOR U27635 ( .A(c5527), .B(n16581), .Z(c5528) );
ANDN U27636 ( .B(n16582), .A(n16583), .Z(n16581) );
XOR U27637 ( .A(c5527), .B(b[5527]), .Z(n16582) );
XNOR U27638 ( .A(b[5527]), .B(n16583), .Z(c[5527]) );
XNOR U27639 ( .A(a[5527]), .B(c5527), .Z(n16583) );
XOR U27640 ( .A(c5528), .B(n16584), .Z(c5529) );
ANDN U27641 ( .B(n16585), .A(n16586), .Z(n16584) );
XOR U27642 ( .A(c5528), .B(b[5528]), .Z(n16585) );
XNOR U27643 ( .A(b[5528]), .B(n16586), .Z(c[5528]) );
XNOR U27644 ( .A(a[5528]), .B(c5528), .Z(n16586) );
XOR U27645 ( .A(c5529), .B(n16587), .Z(c5530) );
ANDN U27646 ( .B(n16588), .A(n16589), .Z(n16587) );
XOR U27647 ( .A(c5529), .B(b[5529]), .Z(n16588) );
XNOR U27648 ( .A(b[5529]), .B(n16589), .Z(c[5529]) );
XNOR U27649 ( .A(a[5529]), .B(c5529), .Z(n16589) );
XOR U27650 ( .A(c5530), .B(n16590), .Z(c5531) );
ANDN U27651 ( .B(n16591), .A(n16592), .Z(n16590) );
XOR U27652 ( .A(c5530), .B(b[5530]), .Z(n16591) );
XNOR U27653 ( .A(b[5530]), .B(n16592), .Z(c[5530]) );
XNOR U27654 ( .A(a[5530]), .B(c5530), .Z(n16592) );
XOR U27655 ( .A(c5531), .B(n16593), .Z(c5532) );
ANDN U27656 ( .B(n16594), .A(n16595), .Z(n16593) );
XOR U27657 ( .A(c5531), .B(b[5531]), .Z(n16594) );
XNOR U27658 ( .A(b[5531]), .B(n16595), .Z(c[5531]) );
XNOR U27659 ( .A(a[5531]), .B(c5531), .Z(n16595) );
XOR U27660 ( .A(c5532), .B(n16596), .Z(c5533) );
ANDN U27661 ( .B(n16597), .A(n16598), .Z(n16596) );
XOR U27662 ( .A(c5532), .B(b[5532]), .Z(n16597) );
XNOR U27663 ( .A(b[5532]), .B(n16598), .Z(c[5532]) );
XNOR U27664 ( .A(a[5532]), .B(c5532), .Z(n16598) );
XOR U27665 ( .A(c5533), .B(n16599), .Z(c5534) );
ANDN U27666 ( .B(n16600), .A(n16601), .Z(n16599) );
XOR U27667 ( .A(c5533), .B(b[5533]), .Z(n16600) );
XNOR U27668 ( .A(b[5533]), .B(n16601), .Z(c[5533]) );
XNOR U27669 ( .A(a[5533]), .B(c5533), .Z(n16601) );
XOR U27670 ( .A(c5534), .B(n16602), .Z(c5535) );
ANDN U27671 ( .B(n16603), .A(n16604), .Z(n16602) );
XOR U27672 ( .A(c5534), .B(b[5534]), .Z(n16603) );
XNOR U27673 ( .A(b[5534]), .B(n16604), .Z(c[5534]) );
XNOR U27674 ( .A(a[5534]), .B(c5534), .Z(n16604) );
XOR U27675 ( .A(c5535), .B(n16605), .Z(c5536) );
ANDN U27676 ( .B(n16606), .A(n16607), .Z(n16605) );
XOR U27677 ( .A(c5535), .B(b[5535]), .Z(n16606) );
XNOR U27678 ( .A(b[5535]), .B(n16607), .Z(c[5535]) );
XNOR U27679 ( .A(a[5535]), .B(c5535), .Z(n16607) );
XOR U27680 ( .A(c5536), .B(n16608), .Z(c5537) );
ANDN U27681 ( .B(n16609), .A(n16610), .Z(n16608) );
XOR U27682 ( .A(c5536), .B(b[5536]), .Z(n16609) );
XNOR U27683 ( .A(b[5536]), .B(n16610), .Z(c[5536]) );
XNOR U27684 ( .A(a[5536]), .B(c5536), .Z(n16610) );
XOR U27685 ( .A(c5537), .B(n16611), .Z(c5538) );
ANDN U27686 ( .B(n16612), .A(n16613), .Z(n16611) );
XOR U27687 ( .A(c5537), .B(b[5537]), .Z(n16612) );
XNOR U27688 ( .A(b[5537]), .B(n16613), .Z(c[5537]) );
XNOR U27689 ( .A(a[5537]), .B(c5537), .Z(n16613) );
XOR U27690 ( .A(c5538), .B(n16614), .Z(c5539) );
ANDN U27691 ( .B(n16615), .A(n16616), .Z(n16614) );
XOR U27692 ( .A(c5538), .B(b[5538]), .Z(n16615) );
XNOR U27693 ( .A(b[5538]), .B(n16616), .Z(c[5538]) );
XNOR U27694 ( .A(a[5538]), .B(c5538), .Z(n16616) );
XOR U27695 ( .A(c5539), .B(n16617), .Z(c5540) );
ANDN U27696 ( .B(n16618), .A(n16619), .Z(n16617) );
XOR U27697 ( .A(c5539), .B(b[5539]), .Z(n16618) );
XNOR U27698 ( .A(b[5539]), .B(n16619), .Z(c[5539]) );
XNOR U27699 ( .A(a[5539]), .B(c5539), .Z(n16619) );
XOR U27700 ( .A(c5540), .B(n16620), .Z(c5541) );
ANDN U27701 ( .B(n16621), .A(n16622), .Z(n16620) );
XOR U27702 ( .A(c5540), .B(b[5540]), .Z(n16621) );
XNOR U27703 ( .A(b[5540]), .B(n16622), .Z(c[5540]) );
XNOR U27704 ( .A(a[5540]), .B(c5540), .Z(n16622) );
XOR U27705 ( .A(c5541), .B(n16623), .Z(c5542) );
ANDN U27706 ( .B(n16624), .A(n16625), .Z(n16623) );
XOR U27707 ( .A(c5541), .B(b[5541]), .Z(n16624) );
XNOR U27708 ( .A(b[5541]), .B(n16625), .Z(c[5541]) );
XNOR U27709 ( .A(a[5541]), .B(c5541), .Z(n16625) );
XOR U27710 ( .A(c5542), .B(n16626), .Z(c5543) );
ANDN U27711 ( .B(n16627), .A(n16628), .Z(n16626) );
XOR U27712 ( .A(c5542), .B(b[5542]), .Z(n16627) );
XNOR U27713 ( .A(b[5542]), .B(n16628), .Z(c[5542]) );
XNOR U27714 ( .A(a[5542]), .B(c5542), .Z(n16628) );
XOR U27715 ( .A(c5543), .B(n16629), .Z(c5544) );
ANDN U27716 ( .B(n16630), .A(n16631), .Z(n16629) );
XOR U27717 ( .A(c5543), .B(b[5543]), .Z(n16630) );
XNOR U27718 ( .A(b[5543]), .B(n16631), .Z(c[5543]) );
XNOR U27719 ( .A(a[5543]), .B(c5543), .Z(n16631) );
XOR U27720 ( .A(c5544), .B(n16632), .Z(c5545) );
ANDN U27721 ( .B(n16633), .A(n16634), .Z(n16632) );
XOR U27722 ( .A(c5544), .B(b[5544]), .Z(n16633) );
XNOR U27723 ( .A(b[5544]), .B(n16634), .Z(c[5544]) );
XNOR U27724 ( .A(a[5544]), .B(c5544), .Z(n16634) );
XOR U27725 ( .A(c5545), .B(n16635), .Z(c5546) );
ANDN U27726 ( .B(n16636), .A(n16637), .Z(n16635) );
XOR U27727 ( .A(c5545), .B(b[5545]), .Z(n16636) );
XNOR U27728 ( .A(b[5545]), .B(n16637), .Z(c[5545]) );
XNOR U27729 ( .A(a[5545]), .B(c5545), .Z(n16637) );
XOR U27730 ( .A(c5546), .B(n16638), .Z(c5547) );
ANDN U27731 ( .B(n16639), .A(n16640), .Z(n16638) );
XOR U27732 ( .A(c5546), .B(b[5546]), .Z(n16639) );
XNOR U27733 ( .A(b[5546]), .B(n16640), .Z(c[5546]) );
XNOR U27734 ( .A(a[5546]), .B(c5546), .Z(n16640) );
XOR U27735 ( .A(c5547), .B(n16641), .Z(c5548) );
ANDN U27736 ( .B(n16642), .A(n16643), .Z(n16641) );
XOR U27737 ( .A(c5547), .B(b[5547]), .Z(n16642) );
XNOR U27738 ( .A(b[5547]), .B(n16643), .Z(c[5547]) );
XNOR U27739 ( .A(a[5547]), .B(c5547), .Z(n16643) );
XOR U27740 ( .A(c5548), .B(n16644), .Z(c5549) );
ANDN U27741 ( .B(n16645), .A(n16646), .Z(n16644) );
XOR U27742 ( .A(c5548), .B(b[5548]), .Z(n16645) );
XNOR U27743 ( .A(b[5548]), .B(n16646), .Z(c[5548]) );
XNOR U27744 ( .A(a[5548]), .B(c5548), .Z(n16646) );
XOR U27745 ( .A(c5549), .B(n16647), .Z(c5550) );
ANDN U27746 ( .B(n16648), .A(n16649), .Z(n16647) );
XOR U27747 ( .A(c5549), .B(b[5549]), .Z(n16648) );
XNOR U27748 ( .A(b[5549]), .B(n16649), .Z(c[5549]) );
XNOR U27749 ( .A(a[5549]), .B(c5549), .Z(n16649) );
XOR U27750 ( .A(c5550), .B(n16650), .Z(c5551) );
ANDN U27751 ( .B(n16651), .A(n16652), .Z(n16650) );
XOR U27752 ( .A(c5550), .B(b[5550]), .Z(n16651) );
XNOR U27753 ( .A(b[5550]), .B(n16652), .Z(c[5550]) );
XNOR U27754 ( .A(a[5550]), .B(c5550), .Z(n16652) );
XOR U27755 ( .A(c5551), .B(n16653), .Z(c5552) );
ANDN U27756 ( .B(n16654), .A(n16655), .Z(n16653) );
XOR U27757 ( .A(c5551), .B(b[5551]), .Z(n16654) );
XNOR U27758 ( .A(b[5551]), .B(n16655), .Z(c[5551]) );
XNOR U27759 ( .A(a[5551]), .B(c5551), .Z(n16655) );
XOR U27760 ( .A(c5552), .B(n16656), .Z(c5553) );
ANDN U27761 ( .B(n16657), .A(n16658), .Z(n16656) );
XOR U27762 ( .A(c5552), .B(b[5552]), .Z(n16657) );
XNOR U27763 ( .A(b[5552]), .B(n16658), .Z(c[5552]) );
XNOR U27764 ( .A(a[5552]), .B(c5552), .Z(n16658) );
XOR U27765 ( .A(c5553), .B(n16659), .Z(c5554) );
ANDN U27766 ( .B(n16660), .A(n16661), .Z(n16659) );
XOR U27767 ( .A(c5553), .B(b[5553]), .Z(n16660) );
XNOR U27768 ( .A(b[5553]), .B(n16661), .Z(c[5553]) );
XNOR U27769 ( .A(a[5553]), .B(c5553), .Z(n16661) );
XOR U27770 ( .A(c5554), .B(n16662), .Z(c5555) );
ANDN U27771 ( .B(n16663), .A(n16664), .Z(n16662) );
XOR U27772 ( .A(c5554), .B(b[5554]), .Z(n16663) );
XNOR U27773 ( .A(b[5554]), .B(n16664), .Z(c[5554]) );
XNOR U27774 ( .A(a[5554]), .B(c5554), .Z(n16664) );
XOR U27775 ( .A(c5555), .B(n16665), .Z(c5556) );
ANDN U27776 ( .B(n16666), .A(n16667), .Z(n16665) );
XOR U27777 ( .A(c5555), .B(b[5555]), .Z(n16666) );
XNOR U27778 ( .A(b[5555]), .B(n16667), .Z(c[5555]) );
XNOR U27779 ( .A(a[5555]), .B(c5555), .Z(n16667) );
XOR U27780 ( .A(c5556), .B(n16668), .Z(c5557) );
ANDN U27781 ( .B(n16669), .A(n16670), .Z(n16668) );
XOR U27782 ( .A(c5556), .B(b[5556]), .Z(n16669) );
XNOR U27783 ( .A(b[5556]), .B(n16670), .Z(c[5556]) );
XNOR U27784 ( .A(a[5556]), .B(c5556), .Z(n16670) );
XOR U27785 ( .A(c5557), .B(n16671), .Z(c5558) );
ANDN U27786 ( .B(n16672), .A(n16673), .Z(n16671) );
XOR U27787 ( .A(c5557), .B(b[5557]), .Z(n16672) );
XNOR U27788 ( .A(b[5557]), .B(n16673), .Z(c[5557]) );
XNOR U27789 ( .A(a[5557]), .B(c5557), .Z(n16673) );
XOR U27790 ( .A(c5558), .B(n16674), .Z(c5559) );
ANDN U27791 ( .B(n16675), .A(n16676), .Z(n16674) );
XOR U27792 ( .A(c5558), .B(b[5558]), .Z(n16675) );
XNOR U27793 ( .A(b[5558]), .B(n16676), .Z(c[5558]) );
XNOR U27794 ( .A(a[5558]), .B(c5558), .Z(n16676) );
XOR U27795 ( .A(c5559), .B(n16677), .Z(c5560) );
ANDN U27796 ( .B(n16678), .A(n16679), .Z(n16677) );
XOR U27797 ( .A(c5559), .B(b[5559]), .Z(n16678) );
XNOR U27798 ( .A(b[5559]), .B(n16679), .Z(c[5559]) );
XNOR U27799 ( .A(a[5559]), .B(c5559), .Z(n16679) );
XOR U27800 ( .A(c5560), .B(n16680), .Z(c5561) );
ANDN U27801 ( .B(n16681), .A(n16682), .Z(n16680) );
XOR U27802 ( .A(c5560), .B(b[5560]), .Z(n16681) );
XNOR U27803 ( .A(b[5560]), .B(n16682), .Z(c[5560]) );
XNOR U27804 ( .A(a[5560]), .B(c5560), .Z(n16682) );
XOR U27805 ( .A(c5561), .B(n16683), .Z(c5562) );
ANDN U27806 ( .B(n16684), .A(n16685), .Z(n16683) );
XOR U27807 ( .A(c5561), .B(b[5561]), .Z(n16684) );
XNOR U27808 ( .A(b[5561]), .B(n16685), .Z(c[5561]) );
XNOR U27809 ( .A(a[5561]), .B(c5561), .Z(n16685) );
XOR U27810 ( .A(c5562), .B(n16686), .Z(c5563) );
ANDN U27811 ( .B(n16687), .A(n16688), .Z(n16686) );
XOR U27812 ( .A(c5562), .B(b[5562]), .Z(n16687) );
XNOR U27813 ( .A(b[5562]), .B(n16688), .Z(c[5562]) );
XNOR U27814 ( .A(a[5562]), .B(c5562), .Z(n16688) );
XOR U27815 ( .A(c5563), .B(n16689), .Z(c5564) );
ANDN U27816 ( .B(n16690), .A(n16691), .Z(n16689) );
XOR U27817 ( .A(c5563), .B(b[5563]), .Z(n16690) );
XNOR U27818 ( .A(b[5563]), .B(n16691), .Z(c[5563]) );
XNOR U27819 ( .A(a[5563]), .B(c5563), .Z(n16691) );
XOR U27820 ( .A(c5564), .B(n16692), .Z(c5565) );
ANDN U27821 ( .B(n16693), .A(n16694), .Z(n16692) );
XOR U27822 ( .A(c5564), .B(b[5564]), .Z(n16693) );
XNOR U27823 ( .A(b[5564]), .B(n16694), .Z(c[5564]) );
XNOR U27824 ( .A(a[5564]), .B(c5564), .Z(n16694) );
XOR U27825 ( .A(c5565), .B(n16695), .Z(c5566) );
ANDN U27826 ( .B(n16696), .A(n16697), .Z(n16695) );
XOR U27827 ( .A(c5565), .B(b[5565]), .Z(n16696) );
XNOR U27828 ( .A(b[5565]), .B(n16697), .Z(c[5565]) );
XNOR U27829 ( .A(a[5565]), .B(c5565), .Z(n16697) );
XOR U27830 ( .A(c5566), .B(n16698), .Z(c5567) );
ANDN U27831 ( .B(n16699), .A(n16700), .Z(n16698) );
XOR U27832 ( .A(c5566), .B(b[5566]), .Z(n16699) );
XNOR U27833 ( .A(b[5566]), .B(n16700), .Z(c[5566]) );
XNOR U27834 ( .A(a[5566]), .B(c5566), .Z(n16700) );
XOR U27835 ( .A(c5567), .B(n16701), .Z(c5568) );
ANDN U27836 ( .B(n16702), .A(n16703), .Z(n16701) );
XOR U27837 ( .A(c5567), .B(b[5567]), .Z(n16702) );
XNOR U27838 ( .A(b[5567]), .B(n16703), .Z(c[5567]) );
XNOR U27839 ( .A(a[5567]), .B(c5567), .Z(n16703) );
XOR U27840 ( .A(c5568), .B(n16704), .Z(c5569) );
ANDN U27841 ( .B(n16705), .A(n16706), .Z(n16704) );
XOR U27842 ( .A(c5568), .B(b[5568]), .Z(n16705) );
XNOR U27843 ( .A(b[5568]), .B(n16706), .Z(c[5568]) );
XNOR U27844 ( .A(a[5568]), .B(c5568), .Z(n16706) );
XOR U27845 ( .A(c5569), .B(n16707), .Z(c5570) );
ANDN U27846 ( .B(n16708), .A(n16709), .Z(n16707) );
XOR U27847 ( .A(c5569), .B(b[5569]), .Z(n16708) );
XNOR U27848 ( .A(b[5569]), .B(n16709), .Z(c[5569]) );
XNOR U27849 ( .A(a[5569]), .B(c5569), .Z(n16709) );
XOR U27850 ( .A(c5570), .B(n16710), .Z(c5571) );
ANDN U27851 ( .B(n16711), .A(n16712), .Z(n16710) );
XOR U27852 ( .A(c5570), .B(b[5570]), .Z(n16711) );
XNOR U27853 ( .A(b[5570]), .B(n16712), .Z(c[5570]) );
XNOR U27854 ( .A(a[5570]), .B(c5570), .Z(n16712) );
XOR U27855 ( .A(c5571), .B(n16713), .Z(c5572) );
ANDN U27856 ( .B(n16714), .A(n16715), .Z(n16713) );
XOR U27857 ( .A(c5571), .B(b[5571]), .Z(n16714) );
XNOR U27858 ( .A(b[5571]), .B(n16715), .Z(c[5571]) );
XNOR U27859 ( .A(a[5571]), .B(c5571), .Z(n16715) );
XOR U27860 ( .A(c5572), .B(n16716), .Z(c5573) );
ANDN U27861 ( .B(n16717), .A(n16718), .Z(n16716) );
XOR U27862 ( .A(c5572), .B(b[5572]), .Z(n16717) );
XNOR U27863 ( .A(b[5572]), .B(n16718), .Z(c[5572]) );
XNOR U27864 ( .A(a[5572]), .B(c5572), .Z(n16718) );
XOR U27865 ( .A(c5573), .B(n16719), .Z(c5574) );
ANDN U27866 ( .B(n16720), .A(n16721), .Z(n16719) );
XOR U27867 ( .A(c5573), .B(b[5573]), .Z(n16720) );
XNOR U27868 ( .A(b[5573]), .B(n16721), .Z(c[5573]) );
XNOR U27869 ( .A(a[5573]), .B(c5573), .Z(n16721) );
XOR U27870 ( .A(c5574), .B(n16722), .Z(c5575) );
ANDN U27871 ( .B(n16723), .A(n16724), .Z(n16722) );
XOR U27872 ( .A(c5574), .B(b[5574]), .Z(n16723) );
XNOR U27873 ( .A(b[5574]), .B(n16724), .Z(c[5574]) );
XNOR U27874 ( .A(a[5574]), .B(c5574), .Z(n16724) );
XOR U27875 ( .A(c5575), .B(n16725), .Z(c5576) );
ANDN U27876 ( .B(n16726), .A(n16727), .Z(n16725) );
XOR U27877 ( .A(c5575), .B(b[5575]), .Z(n16726) );
XNOR U27878 ( .A(b[5575]), .B(n16727), .Z(c[5575]) );
XNOR U27879 ( .A(a[5575]), .B(c5575), .Z(n16727) );
XOR U27880 ( .A(c5576), .B(n16728), .Z(c5577) );
ANDN U27881 ( .B(n16729), .A(n16730), .Z(n16728) );
XOR U27882 ( .A(c5576), .B(b[5576]), .Z(n16729) );
XNOR U27883 ( .A(b[5576]), .B(n16730), .Z(c[5576]) );
XNOR U27884 ( .A(a[5576]), .B(c5576), .Z(n16730) );
XOR U27885 ( .A(c5577), .B(n16731), .Z(c5578) );
ANDN U27886 ( .B(n16732), .A(n16733), .Z(n16731) );
XOR U27887 ( .A(c5577), .B(b[5577]), .Z(n16732) );
XNOR U27888 ( .A(b[5577]), .B(n16733), .Z(c[5577]) );
XNOR U27889 ( .A(a[5577]), .B(c5577), .Z(n16733) );
XOR U27890 ( .A(c5578), .B(n16734), .Z(c5579) );
ANDN U27891 ( .B(n16735), .A(n16736), .Z(n16734) );
XOR U27892 ( .A(c5578), .B(b[5578]), .Z(n16735) );
XNOR U27893 ( .A(b[5578]), .B(n16736), .Z(c[5578]) );
XNOR U27894 ( .A(a[5578]), .B(c5578), .Z(n16736) );
XOR U27895 ( .A(c5579), .B(n16737), .Z(c5580) );
ANDN U27896 ( .B(n16738), .A(n16739), .Z(n16737) );
XOR U27897 ( .A(c5579), .B(b[5579]), .Z(n16738) );
XNOR U27898 ( .A(b[5579]), .B(n16739), .Z(c[5579]) );
XNOR U27899 ( .A(a[5579]), .B(c5579), .Z(n16739) );
XOR U27900 ( .A(c5580), .B(n16740), .Z(c5581) );
ANDN U27901 ( .B(n16741), .A(n16742), .Z(n16740) );
XOR U27902 ( .A(c5580), .B(b[5580]), .Z(n16741) );
XNOR U27903 ( .A(b[5580]), .B(n16742), .Z(c[5580]) );
XNOR U27904 ( .A(a[5580]), .B(c5580), .Z(n16742) );
XOR U27905 ( .A(c5581), .B(n16743), .Z(c5582) );
ANDN U27906 ( .B(n16744), .A(n16745), .Z(n16743) );
XOR U27907 ( .A(c5581), .B(b[5581]), .Z(n16744) );
XNOR U27908 ( .A(b[5581]), .B(n16745), .Z(c[5581]) );
XNOR U27909 ( .A(a[5581]), .B(c5581), .Z(n16745) );
XOR U27910 ( .A(c5582), .B(n16746), .Z(c5583) );
ANDN U27911 ( .B(n16747), .A(n16748), .Z(n16746) );
XOR U27912 ( .A(c5582), .B(b[5582]), .Z(n16747) );
XNOR U27913 ( .A(b[5582]), .B(n16748), .Z(c[5582]) );
XNOR U27914 ( .A(a[5582]), .B(c5582), .Z(n16748) );
XOR U27915 ( .A(c5583), .B(n16749), .Z(c5584) );
ANDN U27916 ( .B(n16750), .A(n16751), .Z(n16749) );
XOR U27917 ( .A(c5583), .B(b[5583]), .Z(n16750) );
XNOR U27918 ( .A(b[5583]), .B(n16751), .Z(c[5583]) );
XNOR U27919 ( .A(a[5583]), .B(c5583), .Z(n16751) );
XOR U27920 ( .A(c5584), .B(n16752), .Z(c5585) );
ANDN U27921 ( .B(n16753), .A(n16754), .Z(n16752) );
XOR U27922 ( .A(c5584), .B(b[5584]), .Z(n16753) );
XNOR U27923 ( .A(b[5584]), .B(n16754), .Z(c[5584]) );
XNOR U27924 ( .A(a[5584]), .B(c5584), .Z(n16754) );
XOR U27925 ( .A(c5585), .B(n16755), .Z(c5586) );
ANDN U27926 ( .B(n16756), .A(n16757), .Z(n16755) );
XOR U27927 ( .A(c5585), .B(b[5585]), .Z(n16756) );
XNOR U27928 ( .A(b[5585]), .B(n16757), .Z(c[5585]) );
XNOR U27929 ( .A(a[5585]), .B(c5585), .Z(n16757) );
XOR U27930 ( .A(c5586), .B(n16758), .Z(c5587) );
ANDN U27931 ( .B(n16759), .A(n16760), .Z(n16758) );
XOR U27932 ( .A(c5586), .B(b[5586]), .Z(n16759) );
XNOR U27933 ( .A(b[5586]), .B(n16760), .Z(c[5586]) );
XNOR U27934 ( .A(a[5586]), .B(c5586), .Z(n16760) );
XOR U27935 ( .A(c5587), .B(n16761), .Z(c5588) );
ANDN U27936 ( .B(n16762), .A(n16763), .Z(n16761) );
XOR U27937 ( .A(c5587), .B(b[5587]), .Z(n16762) );
XNOR U27938 ( .A(b[5587]), .B(n16763), .Z(c[5587]) );
XNOR U27939 ( .A(a[5587]), .B(c5587), .Z(n16763) );
XOR U27940 ( .A(c5588), .B(n16764), .Z(c5589) );
ANDN U27941 ( .B(n16765), .A(n16766), .Z(n16764) );
XOR U27942 ( .A(c5588), .B(b[5588]), .Z(n16765) );
XNOR U27943 ( .A(b[5588]), .B(n16766), .Z(c[5588]) );
XNOR U27944 ( .A(a[5588]), .B(c5588), .Z(n16766) );
XOR U27945 ( .A(c5589), .B(n16767), .Z(c5590) );
ANDN U27946 ( .B(n16768), .A(n16769), .Z(n16767) );
XOR U27947 ( .A(c5589), .B(b[5589]), .Z(n16768) );
XNOR U27948 ( .A(b[5589]), .B(n16769), .Z(c[5589]) );
XNOR U27949 ( .A(a[5589]), .B(c5589), .Z(n16769) );
XOR U27950 ( .A(c5590), .B(n16770), .Z(c5591) );
ANDN U27951 ( .B(n16771), .A(n16772), .Z(n16770) );
XOR U27952 ( .A(c5590), .B(b[5590]), .Z(n16771) );
XNOR U27953 ( .A(b[5590]), .B(n16772), .Z(c[5590]) );
XNOR U27954 ( .A(a[5590]), .B(c5590), .Z(n16772) );
XOR U27955 ( .A(c5591), .B(n16773), .Z(c5592) );
ANDN U27956 ( .B(n16774), .A(n16775), .Z(n16773) );
XOR U27957 ( .A(c5591), .B(b[5591]), .Z(n16774) );
XNOR U27958 ( .A(b[5591]), .B(n16775), .Z(c[5591]) );
XNOR U27959 ( .A(a[5591]), .B(c5591), .Z(n16775) );
XOR U27960 ( .A(c5592), .B(n16776), .Z(c5593) );
ANDN U27961 ( .B(n16777), .A(n16778), .Z(n16776) );
XOR U27962 ( .A(c5592), .B(b[5592]), .Z(n16777) );
XNOR U27963 ( .A(b[5592]), .B(n16778), .Z(c[5592]) );
XNOR U27964 ( .A(a[5592]), .B(c5592), .Z(n16778) );
XOR U27965 ( .A(c5593), .B(n16779), .Z(c5594) );
ANDN U27966 ( .B(n16780), .A(n16781), .Z(n16779) );
XOR U27967 ( .A(c5593), .B(b[5593]), .Z(n16780) );
XNOR U27968 ( .A(b[5593]), .B(n16781), .Z(c[5593]) );
XNOR U27969 ( .A(a[5593]), .B(c5593), .Z(n16781) );
XOR U27970 ( .A(c5594), .B(n16782), .Z(c5595) );
ANDN U27971 ( .B(n16783), .A(n16784), .Z(n16782) );
XOR U27972 ( .A(c5594), .B(b[5594]), .Z(n16783) );
XNOR U27973 ( .A(b[5594]), .B(n16784), .Z(c[5594]) );
XNOR U27974 ( .A(a[5594]), .B(c5594), .Z(n16784) );
XOR U27975 ( .A(c5595), .B(n16785), .Z(c5596) );
ANDN U27976 ( .B(n16786), .A(n16787), .Z(n16785) );
XOR U27977 ( .A(c5595), .B(b[5595]), .Z(n16786) );
XNOR U27978 ( .A(b[5595]), .B(n16787), .Z(c[5595]) );
XNOR U27979 ( .A(a[5595]), .B(c5595), .Z(n16787) );
XOR U27980 ( .A(c5596), .B(n16788), .Z(c5597) );
ANDN U27981 ( .B(n16789), .A(n16790), .Z(n16788) );
XOR U27982 ( .A(c5596), .B(b[5596]), .Z(n16789) );
XNOR U27983 ( .A(b[5596]), .B(n16790), .Z(c[5596]) );
XNOR U27984 ( .A(a[5596]), .B(c5596), .Z(n16790) );
XOR U27985 ( .A(c5597), .B(n16791), .Z(c5598) );
ANDN U27986 ( .B(n16792), .A(n16793), .Z(n16791) );
XOR U27987 ( .A(c5597), .B(b[5597]), .Z(n16792) );
XNOR U27988 ( .A(b[5597]), .B(n16793), .Z(c[5597]) );
XNOR U27989 ( .A(a[5597]), .B(c5597), .Z(n16793) );
XOR U27990 ( .A(c5598), .B(n16794), .Z(c5599) );
ANDN U27991 ( .B(n16795), .A(n16796), .Z(n16794) );
XOR U27992 ( .A(c5598), .B(b[5598]), .Z(n16795) );
XNOR U27993 ( .A(b[5598]), .B(n16796), .Z(c[5598]) );
XNOR U27994 ( .A(a[5598]), .B(c5598), .Z(n16796) );
XOR U27995 ( .A(c5599), .B(n16797), .Z(c5600) );
ANDN U27996 ( .B(n16798), .A(n16799), .Z(n16797) );
XOR U27997 ( .A(c5599), .B(b[5599]), .Z(n16798) );
XNOR U27998 ( .A(b[5599]), .B(n16799), .Z(c[5599]) );
XNOR U27999 ( .A(a[5599]), .B(c5599), .Z(n16799) );
XOR U28000 ( .A(c5600), .B(n16800), .Z(c5601) );
ANDN U28001 ( .B(n16801), .A(n16802), .Z(n16800) );
XOR U28002 ( .A(c5600), .B(b[5600]), .Z(n16801) );
XNOR U28003 ( .A(b[5600]), .B(n16802), .Z(c[5600]) );
XNOR U28004 ( .A(a[5600]), .B(c5600), .Z(n16802) );
XOR U28005 ( .A(c5601), .B(n16803), .Z(c5602) );
ANDN U28006 ( .B(n16804), .A(n16805), .Z(n16803) );
XOR U28007 ( .A(c5601), .B(b[5601]), .Z(n16804) );
XNOR U28008 ( .A(b[5601]), .B(n16805), .Z(c[5601]) );
XNOR U28009 ( .A(a[5601]), .B(c5601), .Z(n16805) );
XOR U28010 ( .A(c5602), .B(n16806), .Z(c5603) );
ANDN U28011 ( .B(n16807), .A(n16808), .Z(n16806) );
XOR U28012 ( .A(c5602), .B(b[5602]), .Z(n16807) );
XNOR U28013 ( .A(b[5602]), .B(n16808), .Z(c[5602]) );
XNOR U28014 ( .A(a[5602]), .B(c5602), .Z(n16808) );
XOR U28015 ( .A(c5603), .B(n16809), .Z(c5604) );
ANDN U28016 ( .B(n16810), .A(n16811), .Z(n16809) );
XOR U28017 ( .A(c5603), .B(b[5603]), .Z(n16810) );
XNOR U28018 ( .A(b[5603]), .B(n16811), .Z(c[5603]) );
XNOR U28019 ( .A(a[5603]), .B(c5603), .Z(n16811) );
XOR U28020 ( .A(c5604), .B(n16812), .Z(c5605) );
ANDN U28021 ( .B(n16813), .A(n16814), .Z(n16812) );
XOR U28022 ( .A(c5604), .B(b[5604]), .Z(n16813) );
XNOR U28023 ( .A(b[5604]), .B(n16814), .Z(c[5604]) );
XNOR U28024 ( .A(a[5604]), .B(c5604), .Z(n16814) );
XOR U28025 ( .A(c5605), .B(n16815), .Z(c5606) );
ANDN U28026 ( .B(n16816), .A(n16817), .Z(n16815) );
XOR U28027 ( .A(c5605), .B(b[5605]), .Z(n16816) );
XNOR U28028 ( .A(b[5605]), .B(n16817), .Z(c[5605]) );
XNOR U28029 ( .A(a[5605]), .B(c5605), .Z(n16817) );
XOR U28030 ( .A(c5606), .B(n16818), .Z(c5607) );
ANDN U28031 ( .B(n16819), .A(n16820), .Z(n16818) );
XOR U28032 ( .A(c5606), .B(b[5606]), .Z(n16819) );
XNOR U28033 ( .A(b[5606]), .B(n16820), .Z(c[5606]) );
XNOR U28034 ( .A(a[5606]), .B(c5606), .Z(n16820) );
XOR U28035 ( .A(c5607), .B(n16821), .Z(c5608) );
ANDN U28036 ( .B(n16822), .A(n16823), .Z(n16821) );
XOR U28037 ( .A(c5607), .B(b[5607]), .Z(n16822) );
XNOR U28038 ( .A(b[5607]), .B(n16823), .Z(c[5607]) );
XNOR U28039 ( .A(a[5607]), .B(c5607), .Z(n16823) );
XOR U28040 ( .A(c5608), .B(n16824), .Z(c5609) );
ANDN U28041 ( .B(n16825), .A(n16826), .Z(n16824) );
XOR U28042 ( .A(c5608), .B(b[5608]), .Z(n16825) );
XNOR U28043 ( .A(b[5608]), .B(n16826), .Z(c[5608]) );
XNOR U28044 ( .A(a[5608]), .B(c5608), .Z(n16826) );
XOR U28045 ( .A(c5609), .B(n16827), .Z(c5610) );
ANDN U28046 ( .B(n16828), .A(n16829), .Z(n16827) );
XOR U28047 ( .A(c5609), .B(b[5609]), .Z(n16828) );
XNOR U28048 ( .A(b[5609]), .B(n16829), .Z(c[5609]) );
XNOR U28049 ( .A(a[5609]), .B(c5609), .Z(n16829) );
XOR U28050 ( .A(c5610), .B(n16830), .Z(c5611) );
ANDN U28051 ( .B(n16831), .A(n16832), .Z(n16830) );
XOR U28052 ( .A(c5610), .B(b[5610]), .Z(n16831) );
XNOR U28053 ( .A(b[5610]), .B(n16832), .Z(c[5610]) );
XNOR U28054 ( .A(a[5610]), .B(c5610), .Z(n16832) );
XOR U28055 ( .A(c5611), .B(n16833), .Z(c5612) );
ANDN U28056 ( .B(n16834), .A(n16835), .Z(n16833) );
XOR U28057 ( .A(c5611), .B(b[5611]), .Z(n16834) );
XNOR U28058 ( .A(b[5611]), .B(n16835), .Z(c[5611]) );
XNOR U28059 ( .A(a[5611]), .B(c5611), .Z(n16835) );
XOR U28060 ( .A(c5612), .B(n16836), .Z(c5613) );
ANDN U28061 ( .B(n16837), .A(n16838), .Z(n16836) );
XOR U28062 ( .A(c5612), .B(b[5612]), .Z(n16837) );
XNOR U28063 ( .A(b[5612]), .B(n16838), .Z(c[5612]) );
XNOR U28064 ( .A(a[5612]), .B(c5612), .Z(n16838) );
XOR U28065 ( .A(c5613), .B(n16839), .Z(c5614) );
ANDN U28066 ( .B(n16840), .A(n16841), .Z(n16839) );
XOR U28067 ( .A(c5613), .B(b[5613]), .Z(n16840) );
XNOR U28068 ( .A(b[5613]), .B(n16841), .Z(c[5613]) );
XNOR U28069 ( .A(a[5613]), .B(c5613), .Z(n16841) );
XOR U28070 ( .A(c5614), .B(n16842), .Z(c5615) );
ANDN U28071 ( .B(n16843), .A(n16844), .Z(n16842) );
XOR U28072 ( .A(c5614), .B(b[5614]), .Z(n16843) );
XNOR U28073 ( .A(b[5614]), .B(n16844), .Z(c[5614]) );
XNOR U28074 ( .A(a[5614]), .B(c5614), .Z(n16844) );
XOR U28075 ( .A(c5615), .B(n16845), .Z(c5616) );
ANDN U28076 ( .B(n16846), .A(n16847), .Z(n16845) );
XOR U28077 ( .A(c5615), .B(b[5615]), .Z(n16846) );
XNOR U28078 ( .A(b[5615]), .B(n16847), .Z(c[5615]) );
XNOR U28079 ( .A(a[5615]), .B(c5615), .Z(n16847) );
XOR U28080 ( .A(c5616), .B(n16848), .Z(c5617) );
ANDN U28081 ( .B(n16849), .A(n16850), .Z(n16848) );
XOR U28082 ( .A(c5616), .B(b[5616]), .Z(n16849) );
XNOR U28083 ( .A(b[5616]), .B(n16850), .Z(c[5616]) );
XNOR U28084 ( .A(a[5616]), .B(c5616), .Z(n16850) );
XOR U28085 ( .A(c5617), .B(n16851), .Z(c5618) );
ANDN U28086 ( .B(n16852), .A(n16853), .Z(n16851) );
XOR U28087 ( .A(c5617), .B(b[5617]), .Z(n16852) );
XNOR U28088 ( .A(b[5617]), .B(n16853), .Z(c[5617]) );
XNOR U28089 ( .A(a[5617]), .B(c5617), .Z(n16853) );
XOR U28090 ( .A(c5618), .B(n16854), .Z(c5619) );
ANDN U28091 ( .B(n16855), .A(n16856), .Z(n16854) );
XOR U28092 ( .A(c5618), .B(b[5618]), .Z(n16855) );
XNOR U28093 ( .A(b[5618]), .B(n16856), .Z(c[5618]) );
XNOR U28094 ( .A(a[5618]), .B(c5618), .Z(n16856) );
XOR U28095 ( .A(c5619), .B(n16857), .Z(c5620) );
ANDN U28096 ( .B(n16858), .A(n16859), .Z(n16857) );
XOR U28097 ( .A(c5619), .B(b[5619]), .Z(n16858) );
XNOR U28098 ( .A(b[5619]), .B(n16859), .Z(c[5619]) );
XNOR U28099 ( .A(a[5619]), .B(c5619), .Z(n16859) );
XOR U28100 ( .A(c5620), .B(n16860), .Z(c5621) );
ANDN U28101 ( .B(n16861), .A(n16862), .Z(n16860) );
XOR U28102 ( .A(c5620), .B(b[5620]), .Z(n16861) );
XNOR U28103 ( .A(b[5620]), .B(n16862), .Z(c[5620]) );
XNOR U28104 ( .A(a[5620]), .B(c5620), .Z(n16862) );
XOR U28105 ( .A(c5621), .B(n16863), .Z(c5622) );
ANDN U28106 ( .B(n16864), .A(n16865), .Z(n16863) );
XOR U28107 ( .A(c5621), .B(b[5621]), .Z(n16864) );
XNOR U28108 ( .A(b[5621]), .B(n16865), .Z(c[5621]) );
XNOR U28109 ( .A(a[5621]), .B(c5621), .Z(n16865) );
XOR U28110 ( .A(c5622), .B(n16866), .Z(c5623) );
ANDN U28111 ( .B(n16867), .A(n16868), .Z(n16866) );
XOR U28112 ( .A(c5622), .B(b[5622]), .Z(n16867) );
XNOR U28113 ( .A(b[5622]), .B(n16868), .Z(c[5622]) );
XNOR U28114 ( .A(a[5622]), .B(c5622), .Z(n16868) );
XOR U28115 ( .A(c5623), .B(n16869), .Z(c5624) );
ANDN U28116 ( .B(n16870), .A(n16871), .Z(n16869) );
XOR U28117 ( .A(c5623), .B(b[5623]), .Z(n16870) );
XNOR U28118 ( .A(b[5623]), .B(n16871), .Z(c[5623]) );
XNOR U28119 ( .A(a[5623]), .B(c5623), .Z(n16871) );
XOR U28120 ( .A(c5624), .B(n16872), .Z(c5625) );
ANDN U28121 ( .B(n16873), .A(n16874), .Z(n16872) );
XOR U28122 ( .A(c5624), .B(b[5624]), .Z(n16873) );
XNOR U28123 ( .A(b[5624]), .B(n16874), .Z(c[5624]) );
XNOR U28124 ( .A(a[5624]), .B(c5624), .Z(n16874) );
XOR U28125 ( .A(c5625), .B(n16875), .Z(c5626) );
ANDN U28126 ( .B(n16876), .A(n16877), .Z(n16875) );
XOR U28127 ( .A(c5625), .B(b[5625]), .Z(n16876) );
XNOR U28128 ( .A(b[5625]), .B(n16877), .Z(c[5625]) );
XNOR U28129 ( .A(a[5625]), .B(c5625), .Z(n16877) );
XOR U28130 ( .A(c5626), .B(n16878), .Z(c5627) );
ANDN U28131 ( .B(n16879), .A(n16880), .Z(n16878) );
XOR U28132 ( .A(c5626), .B(b[5626]), .Z(n16879) );
XNOR U28133 ( .A(b[5626]), .B(n16880), .Z(c[5626]) );
XNOR U28134 ( .A(a[5626]), .B(c5626), .Z(n16880) );
XOR U28135 ( .A(c5627), .B(n16881), .Z(c5628) );
ANDN U28136 ( .B(n16882), .A(n16883), .Z(n16881) );
XOR U28137 ( .A(c5627), .B(b[5627]), .Z(n16882) );
XNOR U28138 ( .A(b[5627]), .B(n16883), .Z(c[5627]) );
XNOR U28139 ( .A(a[5627]), .B(c5627), .Z(n16883) );
XOR U28140 ( .A(c5628), .B(n16884), .Z(c5629) );
ANDN U28141 ( .B(n16885), .A(n16886), .Z(n16884) );
XOR U28142 ( .A(c5628), .B(b[5628]), .Z(n16885) );
XNOR U28143 ( .A(b[5628]), .B(n16886), .Z(c[5628]) );
XNOR U28144 ( .A(a[5628]), .B(c5628), .Z(n16886) );
XOR U28145 ( .A(c5629), .B(n16887), .Z(c5630) );
ANDN U28146 ( .B(n16888), .A(n16889), .Z(n16887) );
XOR U28147 ( .A(c5629), .B(b[5629]), .Z(n16888) );
XNOR U28148 ( .A(b[5629]), .B(n16889), .Z(c[5629]) );
XNOR U28149 ( .A(a[5629]), .B(c5629), .Z(n16889) );
XOR U28150 ( .A(c5630), .B(n16890), .Z(c5631) );
ANDN U28151 ( .B(n16891), .A(n16892), .Z(n16890) );
XOR U28152 ( .A(c5630), .B(b[5630]), .Z(n16891) );
XNOR U28153 ( .A(b[5630]), .B(n16892), .Z(c[5630]) );
XNOR U28154 ( .A(a[5630]), .B(c5630), .Z(n16892) );
XOR U28155 ( .A(c5631), .B(n16893), .Z(c5632) );
ANDN U28156 ( .B(n16894), .A(n16895), .Z(n16893) );
XOR U28157 ( .A(c5631), .B(b[5631]), .Z(n16894) );
XNOR U28158 ( .A(b[5631]), .B(n16895), .Z(c[5631]) );
XNOR U28159 ( .A(a[5631]), .B(c5631), .Z(n16895) );
XOR U28160 ( .A(c5632), .B(n16896), .Z(c5633) );
ANDN U28161 ( .B(n16897), .A(n16898), .Z(n16896) );
XOR U28162 ( .A(c5632), .B(b[5632]), .Z(n16897) );
XNOR U28163 ( .A(b[5632]), .B(n16898), .Z(c[5632]) );
XNOR U28164 ( .A(a[5632]), .B(c5632), .Z(n16898) );
XOR U28165 ( .A(c5633), .B(n16899), .Z(c5634) );
ANDN U28166 ( .B(n16900), .A(n16901), .Z(n16899) );
XOR U28167 ( .A(c5633), .B(b[5633]), .Z(n16900) );
XNOR U28168 ( .A(b[5633]), .B(n16901), .Z(c[5633]) );
XNOR U28169 ( .A(a[5633]), .B(c5633), .Z(n16901) );
XOR U28170 ( .A(c5634), .B(n16902), .Z(c5635) );
ANDN U28171 ( .B(n16903), .A(n16904), .Z(n16902) );
XOR U28172 ( .A(c5634), .B(b[5634]), .Z(n16903) );
XNOR U28173 ( .A(b[5634]), .B(n16904), .Z(c[5634]) );
XNOR U28174 ( .A(a[5634]), .B(c5634), .Z(n16904) );
XOR U28175 ( .A(c5635), .B(n16905), .Z(c5636) );
ANDN U28176 ( .B(n16906), .A(n16907), .Z(n16905) );
XOR U28177 ( .A(c5635), .B(b[5635]), .Z(n16906) );
XNOR U28178 ( .A(b[5635]), .B(n16907), .Z(c[5635]) );
XNOR U28179 ( .A(a[5635]), .B(c5635), .Z(n16907) );
XOR U28180 ( .A(c5636), .B(n16908), .Z(c5637) );
ANDN U28181 ( .B(n16909), .A(n16910), .Z(n16908) );
XOR U28182 ( .A(c5636), .B(b[5636]), .Z(n16909) );
XNOR U28183 ( .A(b[5636]), .B(n16910), .Z(c[5636]) );
XNOR U28184 ( .A(a[5636]), .B(c5636), .Z(n16910) );
XOR U28185 ( .A(c5637), .B(n16911), .Z(c5638) );
ANDN U28186 ( .B(n16912), .A(n16913), .Z(n16911) );
XOR U28187 ( .A(c5637), .B(b[5637]), .Z(n16912) );
XNOR U28188 ( .A(b[5637]), .B(n16913), .Z(c[5637]) );
XNOR U28189 ( .A(a[5637]), .B(c5637), .Z(n16913) );
XOR U28190 ( .A(c5638), .B(n16914), .Z(c5639) );
ANDN U28191 ( .B(n16915), .A(n16916), .Z(n16914) );
XOR U28192 ( .A(c5638), .B(b[5638]), .Z(n16915) );
XNOR U28193 ( .A(b[5638]), .B(n16916), .Z(c[5638]) );
XNOR U28194 ( .A(a[5638]), .B(c5638), .Z(n16916) );
XOR U28195 ( .A(c5639), .B(n16917), .Z(c5640) );
ANDN U28196 ( .B(n16918), .A(n16919), .Z(n16917) );
XOR U28197 ( .A(c5639), .B(b[5639]), .Z(n16918) );
XNOR U28198 ( .A(b[5639]), .B(n16919), .Z(c[5639]) );
XNOR U28199 ( .A(a[5639]), .B(c5639), .Z(n16919) );
XOR U28200 ( .A(c5640), .B(n16920), .Z(c5641) );
ANDN U28201 ( .B(n16921), .A(n16922), .Z(n16920) );
XOR U28202 ( .A(c5640), .B(b[5640]), .Z(n16921) );
XNOR U28203 ( .A(b[5640]), .B(n16922), .Z(c[5640]) );
XNOR U28204 ( .A(a[5640]), .B(c5640), .Z(n16922) );
XOR U28205 ( .A(c5641), .B(n16923), .Z(c5642) );
ANDN U28206 ( .B(n16924), .A(n16925), .Z(n16923) );
XOR U28207 ( .A(c5641), .B(b[5641]), .Z(n16924) );
XNOR U28208 ( .A(b[5641]), .B(n16925), .Z(c[5641]) );
XNOR U28209 ( .A(a[5641]), .B(c5641), .Z(n16925) );
XOR U28210 ( .A(c5642), .B(n16926), .Z(c5643) );
ANDN U28211 ( .B(n16927), .A(n16928), .Z(n16926) );
XOR U28212 ( .A(c5642), .B(b[5642]), .Z(n16927) );
XNOR U28213 ( .A(b[5642]), .B(n16928), .Z(c[5642]) );
XNOR U28214 ( .A(a[5642]), .B(c5642), .Z(n16928) );
XOR U28215 ( .A(c5643), .B(n16929), .Z(c5644) );
ANDN U28216 ( .B(n16930), .A(n16931), .Z(n16929) );
XOR U28217 ( .A(c5643), .B(b[5643]), .Z(n16930) );
XNOR U28218 ( .A(b[5643]), .B(n16931), .Z(c[5643]) );
XNOR U28219 ( .A(a[5643]), .B(c5643), .Z(n16931) );
XOR U28220 ( .A(c5644), .B(n16932), .Z(c5645) );
ANDN U28221 ( .B(n16933), .A(n16934), .Z(n16932) );
XOR U28222 ( .A(c5644), .B(b[5644]), .Z(n16933) );
XNOR U28223 ( .A(b[5644]), .B(n16934), .Z(c[5644]) );
XNOR U28224 ( .A(a[5644]), .B(c5644), .Z(n16934) );
XOR U28225 ( .A(c5645), .B(n16935), .Z(c5646) );
ANDN U28226 ( .B(n16936), .A(n16937), .Z(n16935) );
XOR U28227 ( .A(c5645), .B(b[5645]), .Z(n16936) );
XNOR U28228 ( .A(b[5645]), .B(n16937), .Z(c[5645]) );
XNOR U28229 ( .A(a[5645]), .B(c5645), .Z(n16937) );
XOR U28230 ( .A(c5646), .B(n16938), .Z(c5647) );
ANDN U28231 ( .B(n16939), .A(n16940), .Z(n16938) );
XOR U28232 ( .A(c5646), .B(b[5646]), .Z(n16939) );
XNOR U28233 ( .A(b[5646]), .B(n16940), .Z(c[5646]) );
XNOR U28234 ( .A(a[5646]), .B(c5646), .Z(n16940) );
XOR U28235 ( .A(c5647), .B(n16941), .Z(c5648) );
ANDN U28236 ( .B(n16942), .A(n16943), .Z(n16941) );
XOR U28237 ( .A(c5647), .B(b[5647]), .Z(n16942) );
XNOR U28238 ( .A(b[5647]), .B(n16943), .Z(c[5647]) );
XNOR U28239 ( .A(a[5647]), .B(c5647), .Z(n16943) );
XOR U28240 ( .A(c5648), .B(n16944), .Z(c5649) );
ANDN U28241 ( .B(n16945), .A(n16946), .Z(n16944) );
XOR U28242 ( .A(c5648), .B(b[5648]), .Z(n16945) );
XNOR U28243 ( .A(b[5648]), .B(n16946), .Z(c[5648]) );
XNOR U28244 ( .A(a[5648]), .B(c5648), .Z(n16946) );
XOR U28245 ( .A(c5649), .B(n16947), .Z(c5650) );
ANDN U28246 ( .B(n16948), .A(n16949), .Z(n16947) );
XOR U28247 ( .A(c5649), .B(b[5649]), .Z(n16948) );
XNOR U28248 ( .A(b[5649]), .B(n16949), .Z(c[5649]) );
XNOR U28249 ( .A(a[5649]), .B(c5649), .Z(n16949) );
XOR U28250 ( .A(c5650), .B(n16950), .Z(c5651) );
ANDN U28251 ( .B(n16951), .A(n16952), .Z(n16950) );
XOR U28252 ( .A(c5650), .B(b[5650]), .Z(n16951) );
XNOR U28253 ( .A(b[5650]), .B(n16952), .Z(c[5650]) );
XNOR U28254 ( .A(a[5650]), .B(c5650), .Z(n16952) );
XOR U28255 ( .A(c5651), .B(n16953), .Z(c5652) );
ANDN U28256 ( .B(n16954), .A(n16955), .Z(n16953) );
XOR U28257 ( .A(c5651), .B(b[5651]), .Z(n16954) );
XNOR U28258 ( .A(b[5651]), .B(n16955), .Z(c[5651]) );
XNOR U28259 ( .A(a[5651]), .B(c5651), .Z(n16955) );
XOR U28260 ( .A(c5652), .B(n16956), .Z(c5653) );
ANDN U28261 ( .B(n16957), .A(n16958), .Z(n16956) );
XOR U28262 ( .A(c5652), .B(b[5652]), .Z(n16957) );
XNOR U28263 ( .A(b[5652]), .B(n16958), .Z(c[5652]) );
XNOR U28264 ( .A(a[5652]), .B(c5652), .Z(n16958) );
XOR U28265 ( .A(c5653), .B(n16959), .Z(c5654) );
ANDN U28266 ( .B(n16960), .A(n16961), .Z(n16959) );
XOR U28267 ( .A(c5653), .B(b[5653]), .Z(n16960) );
XNOR U28268 ( .A(b[5653]), .B(n16961), .Z(c[5653]) );
XNOR U28269 ( .A(a[5653]), .B(c5653), .Z(n16961) );
XOR U28270 ( .A(c5654), .B(n16962), .Z(c5655) );
ANDN U28271 ( .B(n16963), .A(n16964), .Z(n16962) );
XOR U28272 ( .A(c5654), .B(b[5654]), .Z(n16963) );
XNOR U28273 ( .A(b[5654]), .B(n16964), .Z(c[5654]) );
XNOR U28274 ( .A(a[5654]), .B(c5654), .Z(n16964) );
XOR U28275 ( .A(c5655), .B(n16965), .Z(c5656) );
ANDN U28276 ( .B(n16966), .A(n16967), .Z(n16965) );
XOR U28277 ( .A(c5655), .B(b[5655]), .Z(n16966) );
XNOR U28278 ( .A(b[5655]), .B(n16967), .Z(c[5655]) );
XNOR U28279 ( .A(a[5655]), .B(c5655), .Z(n16967) );
XOR U28280 ( .A(c5656), .B(n16968), .Z(c5657) );
ANDN U28281 ( .B(n16969), .A(n16970), .Z(n16968) );
XOR U28282 ( .A(c5656), .B(b[5656]), .Z(n16969) );
XNOR U28283 ( .A(b[5656]), .B(n16970), .Z(c[5656]) );
XNOR U28284 ( .A(a[5656]), .B(c5656), .Z(n16970) );
XOR U28285 ( .A(c5657), .B(n16971), .Z(c5658) );
ANDN U28286 ( .B(n16972), .A(n16973), .Z(n16971) );
XOR U28287 ( .A(c5657), .B(b[5657]), .Z(n16972) );
XNOR U28288 ( .A(b[5657]), .B(n16973), .Z(c[5657]) );
XNOR U28289 ( .A(a[5657]), .B(c5657), .Z(n16973) );
XOR U28290 ( .A(c5658), .B(n16974), .Z(c5659) );
ANDN U28291 ( .B(n16975), .A(n16976), .Z(n16974) );
XOR U28292 ( .A(c5658), .B(b[5658]), .Z(n16975) );
XNOR U28293 ( .A(b[5658]), .B(n16976), .Z(c[5658]) );
XNOR U28294 ( .A(a[5658]), .B(c5658), .Z(n16976) );
XOR U28295 ( .A(c5659), .B(n16977), .Z(c5660) );
ANDN U28296 ( .B(n16978), .A(n16979), .Z(n16977) );
XOR U28297 ( .A(c5659), .B(b[5659]), .Z(n16978) );
XNOR U28298 ( .A(b[5659]), .B(n16979), .Z(c[5659]) );
XNOR U28299 ( .A(a[5659]), .B(c5659), .Z(n16979) );
XOR U28300 ( .A(c5660), .B(n16980), .Z(c5661) );
ANDN U28301 ( .B(n16981), .A(n16982), .Z(n16980) );
XOR U28302 ( .A(c5660), .B(b[5660]), .Z(n16981) );
XNOR U28303 ( .A(b[5660]), .B(n16982), .Z(c[5660]) );
XNOR U28304 ( .A(a[5660]), .B(c5660), .Z(n16982) );
XOR U28305 ( .A(c5661), .B(n16983), .Z(c5662) );
ANDN U28306 ( .B(n16984), .A(n16985), .Z(n16983) );
XOR U28307 ( .A(c5661), .B(b[5661]), .Z(n16984) );
XNOR U28308 ( .A(b[5661]), .B(n16985), .Z(c[5661]) );
XNOR U28309 ( .A(a[5661]), .B(c5661), .Z(n16985) );
XOR U28310 ( .A(c5662), .B(n16986), .Z(c5663) );
ANDN U28311 ( .B(n16987), .A(n16988), .Z(n16986) );
XOR U28312 ( .A(c5662), .B(b[5662]), .Z(n16987) );
XNOR U28313 ( .A(b[5662]), .B(n16988), .Z(c[5662]) );
XNOR U28314 ( .A(a[5662]), .B(c5662), .Z(n16988) );
XOR U28315 ( .A(c5663), .B(n16989), .Z(c5664) );
ANDN U28316 ( .B(n16990), .A(n16991), .Z(n16989) );
XOR U28317 ( .A(c5663), .B(b[5663]), .Z(n16990) );
XNOR U28318 ( .A(b[5663]), .B(n16991), .Z(c[5663]) );
XNOR U28319 ( .A(a[5663]), .B(c5663), .Z(n16991) );
XOR U28320 ( .A(c5664), .B(n16992), .Z(c5665) );
ANDN U28321 ( .B(n16993), .A(n16994), .Z(n16992) );
XOR U28322 ( .A(c5664), .B(b[5664]), .Z(n16993) );
XNOR U28323 ( .A(b[5664]), .B(n16994), .Z(c[5664]) );
XNOR U28324 ( .A(a[5664]), .B(c5664), .Z(n16994) );
XOR U28325 ( .A(c5665), .B(n16995), .Z(c5666) );
ANDN U28326 ( .B(n16996), .A(n16997), .Z(n16995) );
XOR U28327 ( .A(c5665), .B(b[5665]), .Z(n16996) );
XNOR U28328 ( .A(b[5665]), .B(n16997), .Z(c[5665]) );
XNOR U28329 ( .A(a[5665]), .B(c5665), .Z(n16997) );
XOR U28330 ( .A(c5666), .B(n16998), .Z(c5667) );
ANDN U28331 ( .B(n16999), .A(n17000), .Z(n16998) );
XOR U28332 ( .A(c5666), .B(b[5666]), .Z(n16999) );
XNOR U28333 ( .A(b[5666]), .B(n17000), .Z(c[5666]) );
XNOR U28334 ( .A(a[5666]), .B(c5666), .Z(n17000) );
XOR U28335 ( .A(c5667), .B(n17001), .Z(c5668) );
ANDN U28336 ( .B(n17002), .A(n17003), .Z(n17001) );
XOR U28337 ( .A(c5667), .B(b[5667]), .Z(n17002) );
XNOR U28338 ( .A(b[5667]), .B(n17003), .Z(c[5667]) );
XNOR U28339 ( .A(a[5667]), .B(c5667), .Z(n17003) );
XOR U28340 ( .A(c5668), .B(n17004), .Z(c5669) );
ANDN U28341 ( .B(n17005), .A(n17006), .Z(n17004) );
XOR U28342 ( .A(c5668), .B(b[5668]), .Z(n17005) );
XNOR U28343 ( .A(b[5668]), .B(n17006), .Z(c[5668]) );
XNOR U28344 ( .A(a[5668]), .B(c5668), .Z(n17006) );
XOR U28345 ( .A(c5669), .B(n17007), .Z(c5670) );
ANDN U28346 ( .B(n17008), .A(n17009), .Z(n17007) );
XOR U28347 ( .A(c5669), .B(b[5669]), .Z(n17008) );
XNOR U28348 ( .A(b[5669]), .B(n17009), .Z(c[5669]) );
XNOR U28349 ( .A(a[5669]), .B(c5669), .Z(n17009) );
XOR U28350 ( .A(c5670), .B(n17010), .Z(c5671) );
ANDN U28351 ( .B(n17011), .A(n17012), .Z(n17010) );
XOR U28352 ( .A(c5670), .B(b[5670]), .Z(n17011) );
XNOR U28353 ( .A(b[5670]), .B(n17012), .Z(c[5670]) );
XNOR U28354 ( .A(a[5670]), .B(c5670), .Z(n17012) );
XOR U28355 ( .A(c5671), .B(n17013), .Z(c5672) );
ANDN U28356 ( .B(n17014), .A(n17015), .Z(n17013) );
XOR U28357 ( .A(c5671), .B(b[5671]), .Z(n17014) );
XNOR U28358 ( .A(b[5671]), .B(n17015), .Z(c[5671]) );
XNOR U28359 ( .A(a[5671]), .B(c5671), .Z(n17015) );
XOR U28360 ( .A(c5672), .B(n17016), .Z(c5673) );
ANDN U28361 ( .B(n17017), .A(n17018), .Z(n17016) );
XOR U28362 ( .A(c5672), .B(b[5672]), .Z(n17017) );
XNOR U28363 ( .A(b[5672]), .B(n17018), .Z(c[5672]) );
XNOR U28364 ( .A(a[5672]), .B(c5672), .Z(n17018) );
XOR U28365 ( .A(c5673), .B(n17019), .Z(c5674) );
ANDN U28366 ( .B(n17020), .A(n17021), .Z(n17019) );
XOR U28367 ( .A(c5673), .B(b[5673]), .Z(n17020) );
XNOR U28368 ( .A(b[5673]), .B(n17021), .Z(c[5673]) );
XNOR U28369 ( .A(a[5673]), .B(c5673), .Z(n17021) );
XOR U28370 ( .A(c5674), .B(n17022), .Z(c5675) );
ANDN U28371 ( .B(n17023), .A(n17024), .Z(n17022) );
XOR U28372 ( .A(c5674), .B(b[5674]), .Z(n17023) );
XNOR U28373 ( .A(b[5674]), .B(n17024), .Z(c[5674]) );
XNOR U28374 ( .A(a[5674]), .B(c5674), .Z(n17024) );
XOR U28375 ( .A(c5675), .B(n17025), .Z(c5676) );
ANDN U28376 ( .B(n17026), .A(n17027), .Z(n17025) );
XOR U28377 ( .A(c5675), .B(b[5675]), .Z(n17026) );
XNOR U28378 ( .A(b[5675]), .B(n17027), .Z(c[5675]) );
XNOR U28379 ( .A(a[5675]), .B(c5675), .Z(n17027) );
XOR U28380 ( .A(c5676), .B(n17028), .Z(c5677) );
ANDN U28381 ( .B(n17029), .A(n17030), .Z(n17028) );
XOR U28382 ( .A(c5676), .B(b[5676]), .Z(n17029) );
XNOR U28383 ( .A(b[5676]), .B(n17030), .Z(c[5676]) );
XNOR U28384 ( .A(a[5676]), .B(c5676), .Z(n17030) );
XOR U28385 ( .A(c5677), .B(n17031), .Z(c5678) );
ANDN U28386 ( .B(n17032), .A(n17033), .Z(n17031) );
XOR U28387 ( .A(c5677), .B(b[5677]), .Z(n17032) );
XNOR U28388 ( .A(b[5677]), .B(n17033), .Z(c[5677]) );
XNOR U28389 ( .A(a[5677]), .B(c5677), .Z(n17033) );
XOR U28390 ( .A(c5678), .B(n17034), .Z(c5679) );
ANDN U28391 ( .B(n17035), .A(n17036), .Z(n17034) );
XOR U28392 ( .A(c5678), .B(b[5678]), .Z(n17035) );
XNOR U28393 ( .A(b[5678]), .B(n17036), .Z(c[5678]) );
XNOR U28394 ( .A(a[5678]), .B(c5678), .Z(n17036) );
XOR U28395 ( .A(c5679), .B(n17037), .Z(c5680) );
ANDN U28396 ( .B(n17038), .A(n17039), .Z(n17037) );
XOR U28397 ( .A(c5679), .B(b[5679]), .Z(n17038) );
XNOR U28398 ( .A(b[5679]), .B(n17039), .Z(c[5679]) );
XNOR U28399 ( .A(a[5679]), .B(c5679), .Z(n17039) );
XOR U28400 ( .A(c5680), .B(n17040), .Z(c5681) );
ANDN U28401 ( .B(n17041), .A(n17042), .Z(n17040) );
XOR U28402 ( .A(c5680), .B(b[5680]), .Z(n17041) );
XNOR U28403 ( .A(b[5680]), .B(n17042), .Z(c[5680]) );
XNOR U28404 ( .A(a[5680]), .B(c5680), .Z(n17042) );
XOR U28405 ( .A(c5681), .B(n17043), .Z(c5682) );
ANDN U28406 ( .B(n17044), .A(n17045), .Z(n17043) );
XOR U28407 ( .A(c5681), .B(b[5681]), .Z(n17044) );
XNOR U28408 ( .A(b[5681]), .B(n17045), .Z(c[5681]) );
XNOR U28409 ( .A(a[5681]), .B(c5681), .Z(n17045) );
XOR U28410 ( .A(c5682), .B(n17046), .Z(c5683) );
ANDN U28411 ( .B(n17047), .A(n17048), .Z(n17046) );
XOR U28412 ( .A(c5682), .B(b[5682]), .Z(n17047) );
XNOR U28413 ( .A(b[5682]), .B(n17048), .Z(c[5682]) );
XNOR U28414 ( .A(a[5682]), .B(c5682), .Z(n17048) );
XOR U28415 ( .A(c5683), .B(n17049), .Z(c5684) );
ANDN U28416 ( .B(n17050), .A(n17051), .Z(n17049) );
XOR U28417 ( .A(c5683), .B(b[5683]), .Z(n17050) );
XNOR U28418 ( .A(b[5683]), .B(n17051), .Z(c[5683]) );
XNOR U28419 ( .A(a[5683]), .B(c5683), .Z(n17051) );
XOR U28420 ( .A(c5684), .B(n17052), .Z(c5685) );
ANDN U28421 ( .B(n17053), .A(n17054), .Z(n17052) );
XOR U28422 ( .A(c5684), .B(b[5684]), .Z(n17053) );
XNOR U28423 ( .A(b[5684]), .B(n17054), .Z(c[5684]) );
XNOR U28424 ( .A(a[5684]), .B(c5684), .Z(n17054) );
XOR U28425 ( .A(c5685), .B(n17055), .Z(c5686) );
ANDN U28426 ( .B(n17056), .A(n17057), .Z(n17055) );
XOR U28427 ( .A(c5685), .B(b[5685]), .Z(n17056) );
XNOR U28428 ( .A(b[5685]), .B(n17057), .Z(c[5685]) );
XNOR U28429 ( .A(a[5685]), .B(c5685), .Z(n17057) );
XOR U28430 ( .A(c5686), .B(n17058), .Z(c5687) );
ANDN U28431 ( .B(n17059), .A(n17060), .Z(n17058) );
XOR U28432 ( .A(c5686), .B(b[5686]), .Z(n17059) );
XNOR U28433 ( .A(b[5686]), .B(n17060), .Z(c[5686]) );
XNOR U28434 ( .A(a[5686]), .B(c5686), .Z(n17060) );
XOR U28435 ( .A(c5687), .B(n17061), .Z(c5688) );
ANDN U28436 ( .B(n17062), .A(n17063), .Z(n17061) );
XOR U28437 ( .A(c5687), .B(b[5687]), .Z(n17062) );
XNOR U28438 ( .A(b[5687]), .B(n17063), .Z(c[5687]) );
XNOR U28439 ( .A(a[5687]), .B(c5687), .Z(n17063) );
XOR U28440 ( .A(c5688), .B(n17064), .Z(c5689) );
ANDN U28441 ( .B(n17065), .A(n17066), .Z(n17064) );
XOR U28442 ( .A(c5688), .B(b[5688]), .Z(n17065) );
XNOR U28443 ( .A(b[5688]), .B(n17066), .Z(c[5688]) );
XNOR U28444 ( .A(a[5688]), .B(c5688), .Z(n17066) );
XOR U28445 ( .A(c5689), .B(n17067), .Z(c5690) );
ANDN U28446 ( .B(n17068), .A(n17069), .Z(n17067) );
XOR U28447 ( .A(c5689), .B(b[5689]), .Z(n17068) );
XNOR U28448 ( .A(b[5689]), .B(n17069), .Z(c[5689]) );
XNOR U28449 ( .A(a[5689]), .B(c5689), .Z(n17069) );
XOR U28450 ( .A(c5690), .B(n17070), .Z(c5691) );
ANDN U28451 ( .B(n17071), .A(n17072), .Z(n17070) );
XOR U28452 ( .A(c5690), .B(b[5690]), .Z(n17071) );
XNOR U28453 ( .A(b[5690]), .B(n17072), .Z(c[5690]) );
XNOR U28454 ( .A(a[5690]), .B(c5690), .Z(n17072) );
XOR U28455 ( .A(c5691), .B(n17073), .Z(c5692) );
ANDN U28456 ( .B(n17074), .A(n17075), .Z(n17073) );
XOR U28457 ( .A(c5691), .B(b[5691]), .Z(n17074) );
XNOR U28458 ( .A(b[5691]), .B(n17075), .Z(c[5691]) );
XNOR U28459 ( .A(a[5691]), .B(c5691), .Z(n17075) );
XOR U28460 ( .A(c5692), .B(n17076), .Z(c5693) );
ANDN U28461 ( .B(n17077), .A(n17078), .Z(n17076) );
XOR U28462 ( .A(c5692), .B(b[5692]), .Z(n17077) );
XNOR U28463 ( .A(b[5692]), .B(n17078), .Z(c[5692]) );
XNOR U28464 ( .A(a[5692]), .B(c5692), .Z(n17078) );
XOR U28465 ( .A(c5693), .B(n17079), .Z(c5694) );
ANDN U28466 ( .B(n17080), .A(n17081), .Z(n17079) );
XOR U28467 ( .A(c5693), .B(b[5693]), .Z(n17080) );
XNOR U28468 ( .A(b[5693]), .B(n17081), .Z(c[5693]) );
XNOR U28469 ( .A(a[5693]), .B(c5693), .Z(n17081) );
XOR U28470 ( .A(c5694), .B(n17082), .Z(c5695) );
ANDN U28471 ( .B(n17083), .A(n17084), .Z(n17082) );
XOR U28472 ( .A(c5694), .B(b[5694]), .Z(n17083) );
XNOR U28473 ( .A(b[5694]), .B(n17084), .Z(c[5694]) );
XNOR U28474 ( .A(a[5694]), .B(c5694), .Z(n17084) );
XOR U28475 ( .A(c5695), .B(n17085), .Z(c5696) );
ANDN U28476 ( .B(n17086), .A(n17087), .Z(n17085) );
XOR U28477 ( .A(c5695), .B(b[5695]), .Z(n17086) );
XNOR U28478 ( .A(b[5695]), .B(n17087), .Z(c[5695]) );
XNOR U28479 ( .A(a[5695]), .B(c5695), .Z(n17087) );
XOR U28480 ( .A(c5696), .B(n17088), .Z(c5697) );
ANDN U28481 ( .B(n17089), .A(n17090), .Z(n17088) );
XOR U28482 ( .A(c5696), .B(b[5696]), .Z(n17089) );
XNOR U28483 ( .A(b[5696]), .B(n17090), .Z(c[5696]) );
XNOR U28484 ( .A(a[5696]), .B(c5696), .Z(n17090) );
XOR U28485 ( .A(c5697), .B(n17091), .Z(c5698) );
ANDN U28486 ( .B(n17092), .A(n17093), .Z(n17091) );
XOR U28487 ( .A(c5697), .B(b[5697]), .Z(n17092) );
XNOR U28488 ( .A(b[5697]), .B(n17093), .Z(c[5697]) );
XNOR U28489 ( .A(a[5697]), .B(c5697), .Z(n17093) );
XOR U28490 ( .A(c5698), .B(n17094), .Z(c5699) );
ANDN U28491 ( .B(n17095), .A(n17096), .Z(n17094) );
XOR U28492 ( .A(c5698), .B(b[5698]), .Z(n17095) );
XNOR U28493 ( .A(b[5698]), .B(n17096), .Z(c[5698]) );
XNOR U28494 ( .A(a[5698]), .B(c5698), .Z(n17096) );
XOR U28495 ( .A(c5699), .B(n17097), .Z(c5700) );
ANDN U28496 ( .B(n17098), .A(n17099), .Z(n17097) );
XOR U28497 ( .A(c5699), .B(b[5699]), .Z(n17098) );
XNOR U28498 ( .A(b[5699]), .B(n17099), .Z(c[5699]) );
XNOR U28499 ( .A(a[5699]), .B(c5699), .Z(n17099) );
XOR U28500 ( .A(c5700), .B(n17100), .Z(c5701) );
ANDN U28501 ( .B(n17101), .A(n17102), .Z(n17100) );
XOR U28502 ( .A(c5700), .B(b[5700]), .Z(n17101) );
XNOR U28503 ( .A(b[5700]), .B(n17102), .Z(c[5700]) );
XNOR U28504 ( .A(a[5700]), .B(c5700), .Z(n17102) );
XOR U28505 ( .A(c5701), .B(n17103), .Z(c5702) );
ANDN U28506 ( .B(n17104), .A(n17105), .Z(n17103) );
XOR U28507 ( .A(c5701), .B(b[5701]), .Z(n17104) );
XNOR U28508 ( .A(b[5701]), .B(n17105), .Z(c[5701]) );
XNOR U28509 ( .A(a[5701]), .B(c5701), .Z(n17105) );
XOR U28510 ( .A(c5702), .B(n17106), .Z(c5703) );
ANDN U28511 ( .B(n17107), .A(n17108), .Z(n17106) );
XOR U28512 ( .A(c5702), .B(b[5702]), .Z(n17107) );
XNOR U28513 ( .A(b[5702]), .B(n17108), .Z(c[5702]) );
XNOR U28514 ( .A(a[5702]), .B(c5702), .Z(n17108) );
XOR U28515 ( .A(c5703), .B(n17109), .Z(c5704) );
ANDN U28516 ( .B(n17110), .A(n17111), .Z(n17109) );
XOR U28517 ( .A(c5703), .B(b[5703]), .Z(n17110) );
XNOR U28518 ( .A(b[5703]), .B(n17111), .Z(c[5703]) );
XNOR U28519 ( .A(a[5703]), .B(c5703), .Z(n17111) );
XOR U28520 ( .A(c5704), .B(n17112), .Z(c5705) );
ANDN U28521 ( .B(n17113), .A(n17114), .Z(n17112) );
XOR U28522 ( .A(c5704), .B(b[5704]), .Z(n17113) );
XNOR U28523 ( .A(b[5704]), .B(n17114), .Z(c[5704]) );
XNOR U28524 ( .A(a[5704]), .B(c5704), .Z(n17114) );
XOR U28525 ( .A(c5705), .B(n17115), .Z(c5706) );
ANDN U28526 ( .B(n17116), .A(n17117), .Z(n17115) );
XOR U28527 ( .A(c5705), .B(b[5705]), .Z(n17116) );
XNOR U28528 ( .A(b[5705]), .B(n17117), .Z(c[5705]) );
XNOR U28529 ( .A(a[5705]), .B(c5705), .Z(n17117) );
XOR U28530 ( .A(c5706), .B(n17118), .Z(c5707) );
ANDN U28531 ( .B(n17119), .A(n17120), .Z(n17118) );
XOR U28532 ( .A(c5706), .B(b[5706]), .Z(n17119) );
XNOR U28533 ( .A(b[5706]), .B(n17120), .Z(c[5706]) );
XNOR U28534 ( .A(a[5706]), .B(c5706), .Z(n17120) );
XOR U28535 ( .A(c5707), .B(n17121), .Z(c5708) );
ANDN U28536 ( .B(n17122), .A(n17123), .Z(n17121) );
XOR U28537 ( .A(c5707), .B(b[5707]), .Z(n17122) );
XNOR U28538 ( .A(b[5707]), .B(n17123), .Z(c[5707]) );
XNOR U28539 ( .A(a[5707]), .B(c5707), .Z(n17123) );
XOR U28540 ( .A(c5708), .B(n17124), .Z(c5709) );
ANDN U28541 ( .B(n17125), .A(n17126), .Z(n17124) );
XOR U28542 ( .A(c5708), .B(b[5708]), .Z(n17125) );
XNOR U28543 ( .A(b[5708]), .B(n17126), .Z(c[5708]) );
XNOR U28544 ( .A(a[5708]), .B(c5708), .Z(n17126) );
XOR U28545 ( .A(c5709), .B(n17127), .Z(c5710) );
ANDN U28546 ( .B(n17128), .A(n17129), .Z(n17127) );
XOR U28547 ( .A(c5709), .B(b[5709]), .Z(n17128) );
XNOR U28548 ( .A(b[5709]), .B(n17129), .Z(c[5709]) );
XNOR U28549 ( .A(a[5709]), .B(c5709), .Z(n17129) );
XOR U28550 ( .A(c5710), .B(n17130), .Z(c5711) );
ANDN U28551 ( .B(n17131), .A(n17132), .Z(n17130) );
XOR U28552 ( .A(c5710), .B(b[5710]), .Z(n17131) );
XNOR U28553 ( .A(b[5710]), .B(n17132), .Z(c[5710]) );
XNOR U28554 ( .A(a[5710]), .B(c5710), .Z(n17132) );
XOR U28555 ( .A(c5711), .B(n17133), .Z(c5712) );
ANDN U28556 ( .B(n17134), .A(n17135), .Z(n17133) );
XOR U28557 ( .A(c5711), .B(b[5711]), .Z(n17134) );
XNOR U28558 ( .A(b[5711]), .B(n17135), .Z(c[5711]) );
XNOR U28559 ( .A(a[5711]), .B(c5711), .Z(n17135) );
XOR U28560 ( .A(c5712), .B(n17136), .Z(c5713) );
ANDN U28561 ( .B(n17137), .A(n17138), .Z(n17136) );
XOR U28562 ( .A(c5712), .B(b[5712]), .Z(n17137) );
XNOR U28563 ( .A(b[5712]), .B(n17138), .Z(c[5712]) );
XNOR U28564 ( .A(a[5712]), .B(c5712), .Z(n17138) );
XOR U28565 ( .A(c5713), .B(n17139), .Z(c5714) );
ANDN U28566 ( .B(n17140), .A(n17141), .Z(n17139) );
XOR U28567 ( .A(c5713), .B(b[5713]), .Z(n17140) );
XNOR U28568 ( .A(b[5713]), .B(n17141), .Z(c[5713]) );
XNOR U28569 ( .A(a[5713]), .B(c5713), .Z(n17141) );
XOR U28570 ( .A(c5714), .B(n17142), .Z(c5715) );
ANDN U28571 ( .B(n17143), .A(n17144), .Z(n17142) );
XOR U28572 ( .A(c5714), .B(b[5714]), .Z(n17143) );
XNOR U28573 ( .A(b[5714]), .B(n17144), .Z(c[5714]) );
XNOR U28574 ( .A(a[5714]), .B(c5714), .Z(n17144) );
XOR U28575 ( .A(c5715), .B(n17145), .Z(c5716) );
ANDN U28576 ( .B(n17146), .A(n17147), .Z(n17145) );
XOR U28577 ( .A(c5715), .B(b[5715]), .Z(n17146) );
XNOR U28578 ( .A(b[5715]), .B(n17147), .Z(c[5715]) );
XNOR U28579 ( .A(a[5715]), .B(c5715), .Z(n17147) );
XOR U28580 ( .A(c5716), .B(n17148), .Z(c5717) );
ANDN U28581 ( .B(n17149), .A(n17150), .Z(n17148) );
XOR U28582 ( .A(c5716), .B(b[5716]), .Z(n17149) );
XNOR U28583 ( .A(b[5716]), .B(n17150), .Z(c[5716]) );
XNOR U28584 ( .A(a[5716]), .B(c5716), .Z(n17150) );
XOR U28585 ( .A(c5717), .B(n17151), .Z(c5718) );
ANDN U28586 ( .B(n17152), .A(n17153), .Z(n17151) );
XOR U28587 ( .A(c5717), .B(b[5717]), .Z(n17152) );
XNOR U28588 ( .A(b[5717]), .B(n17153), .Z(c[5717]) );
XNOR U28589 ( .A(a[5717]), .B(c5717), .Z(n17153) );
XOR U28590 ( .A(c5718), .B(n17154), .Z(c5719) );
ANDN U28591 ( .B(n17155), .A(n17156), .Z(n17154) );
XOR U28592 ( .A(c5718), .B(b[5718]), .Z(n17155) );
XNOR U28593 ( .A(b[5718]), .B(n17156), .Z(c[5718]) );
XNOR U28594 ( .A(a[5718]), .B(c5718), .Z(n17156) );
XOR U28595 ( .A(c5719), .B(n17157), .Z(c5720) );
ANDN U28596 ( .B(n17158), .A(n17159), .Z(n17157) );
XOR U28597 ( .A(c5719), .B(b[5719]), .Z(n17158) );
XNOR U28598 ( .A(b[5719]), .B(n17159), .Z(c[5719]) );
XNOR U28599 ( .A(a[5719]), .B(c5719), .Z(n17159) );
XOR U28600 ( .A(c5720), .B(n17160), .Z(c5721) );
ANDN U28601 ( .B(n17161), .A(n17162), .Z(n17160) );
XOR U28602 ( .A(c5720), .B(b[5720]), .Z(n17161) );
XNOR U28603 ( .A(b[5720]), .B(n17162), .Z(c[5720]) );
XNOR U28604 ( .A(a[5720]), .B(c5720), .Z(n17162) );
XOR U28605 ( .A(c5721), .B(n17163), .Z(c5722) );
ANDN U28606 ( .B(n17164), .A(n17165), .Z(n17163) );
XOR U28607 ( .A(c5721), .B(b[5721]), .Z(n17164) );
XNOR U28608 ( .A(b[5721]), .B(n17165), .Z(c[5721]) );
XNOR U28609 ( .A(a[5721]), .B(c5721), .Z(n17165) );
XOR U28610 ( .A(c5722), .B(n17166), .Z(c5723) );
ANDN U28611 ( .B(n17167), .A(n17168), .Z(n17166) );
XOR U28612 ( .A(c5722), .B(b[5722]), .Z(n17167) );
XNOR U28613 ( .A(b[5722]), .B(n17168), .Z(c[5722]) );
XNOR U28614 ( .A(a[5722]), .B(c5722), .Z(n17168) );
XOR U28615 ( .A(c5723), .B(n17169), .Z(c5724) );
ANDN U28616 ( .B(n17170), .A(n17171), .Z(n17169) );
XOR U28617 ( .A(c5723), .B(b[5723]), .Z(n17170) );
XNOR U28618 ( .A(b[5723]), .B(n17171), .Z(c[5723]) );
XNOR U28619 ( .A(a[5723]), .B(c5723), .Z(n17171) );
XOR U28620 ( .A(c5724), .B(n17172), .Z(c5725) );
ANDN U28621 ( .B(n17173), .A(n17174), .Z(n17172) );
XOR U28622 ( .A(c5724), .B(b[5724]), .Z(n17173) );
XNOR U28623 ( .A(b[5724]), .B(n17174), .Z(c[5724]) );
XNOR U28624 ( .A(a[5724]), .B(c5724), .Z(n17174) );
XOR U28625 ( .A(c5725), .B(n17175), .Z(c5726) );
ANDN U28626 ( .B(n17176), .A(n17177), .Z(n17175) );
XOR U28627 ( .A(c5725), .B(b[5725]), .Z(n17176) );
XNOR U28628 ( .A(b[5725]), .B(n17177), .Z(c[5725]) );
XNOR U28629 ( .A(a[5725]), .B(c5725), .Z(n17177) );
XOR U28630 ( .A(c5726), .B(n17178), .Z(c5727) );
ANDN U28631 ( .B(n17179), .A(n17180), .Z(n17178) );
XOR U28632 ( .A(c5726), .B(b[5726]), .Z(n17179) );
XNOR U28633 ( .A(b[5726]), .B(n17180), .Z(c[5726]) );
XNOR U28634 ( .A(a[5726]), .B(c5726), .Z(n17180) );
XOR U28635 ( .A(c5727), .B(n17181), .Z(c5728) );
ANDN U28636 ( .B(n17182), .A(n17183), .Z(n17181) );
XOR U28637 ( .A(c5727), .B(b[5727]), .Z(n17182) );
XNOR U28638 ( .A(b[5727]), .B(n17183), .Z(c[5727]) );
XNOR U28639 ( .A(a[5727]), .B(c5727), .Z(n17183) );
XOR U28640 ( .A(c5728), .B(n17184), .Z(c5729) );
ANDN U28641 ( .B(n17185), .A(n17186), .Z(n17184) );
XOR U28642 ( .A(c5728), .B(b[5728]), .Z(n17185) );
XNOR U28643 ( .A(b[5728]), .B(n17186), .Z(c[5728]) );
XNOR U28644 ( .A(a[5728]), .B(c5728), .Z(n17186) );
XOR U28645 ( .A(c5729), .B(n17187), .Z(c5730) );
ANDN U28646 ( .B(n17188), .A(n17189), .Z(n17187) );
XOR U28647 ( .A(c5729), .B(b[5729]), .Z(n17188) );
XNOR U28648 ( .A(b[5729]), .B(n17189), .Z(c[5729]) );
XNOR U28649 ( .A(a[5729]), .B(c5729), .Z(n17189) );
XOR U28650 ( .A(c5730), .B(n17190), .Z(c5731) );
ANDN U28651 ( .B(n17191), .A(n17192), .Z(n17190) );
XOR U28652 ( .A(c5730), .B(b[5730]), .Z(n17191) );
XNOR U28653 ( .A(b[5730]), .B(n17192), .Z(c[5730]) );
XNOR U28654 ( .A(a[5730]), .B(c5730), .Z(n17192) );
XOR U28655 ( .A(c5731), .B(n17193), .Z(c5732) );
ANDN U28656 ( .B(n17194), .A(n17195), .Z(n17193) );
XOR U28657 ( .A(c5731), .B(b[5731]), .Z(n17194) );
XNOR U28658 ( .A(b[5731]), .B(n17195), .Z(c[5731]) );
XNOR U28659 ( .A(a[5731]), .B(c5731), .Z(n17195) );
XOR U28660 ( .A(c5732), .B(n17196), .Z(c5733) );
ANDN U28661 ( .B(n17197), .A(n17198), .Z(n17196) );
XOR U28662 ( .A(c5732), .B(b[5732]), .Z(n17197) );
XNOR U28663 ( .A(b[5732]), .B(n17198), .Z(c[5732]) );
XNOR U28664 ( .A(a[5732]), .B(c5732), .Z(n17198) );
XOR U28665 ( .A(c5733), .B(n17199), .Z(c5734) );
ANDN U28666 ( .B(n17200), .A(n17201), .Z(n17199) );
XOR U28667 ( .A(c5733), .B(b[5733]), .Z(n17200) );
XNOR U28668 ( .A(b[5733]), .B(n17201), .Z(c[5733]) );
XNOR U28669 ( .A(a[5733]), .B(c5733), .Z(n17201) );
XOR U28670 ( .A(c5734), .B(n17202), .Z(c5735) );
ANDN U28671 ( .B(n17203), .A(n17204), .Z(n17202) );
XOR U28672 ( .A(c5734), .B(b[5734]), .Z(n17203) );
XNOR U28673 ( .A(b[5734]), .B(n17204), .Z(c[5734]) );
XNOR U28674 ( .A(a[5734]), .B(c5734), .Z(n17204) );
XOR U28675 ( .A(c5735), .B(n17205), .Z(c5736) );
ANDN U28676 ( .B(n17206), .A(n17207), .Z(n17205) );
XOR U28677 ( .A(c5735), .B(b[5735]), .Z(n17206) );
XNOR U28678 ( .A(b[5735]), .B(n17207), .Z(c[5735]) );
XNOR U28679 ( .A(a[5735]), .B(c5735), .Z(n17207) );
XOR U28680 ( .A(c5736), .B(n17208), .Z(c5737) );
ANDN U28681 ( .B(n17209), .A(n17210), .Z(n17208) );
XOR U28682 ( .A(c5736), .B(b[5736]), .Z(n17209) );
XNOR U28683 ( .A(b[5736]), .B(n17210), .Z(c[5736]) );
XNOR U28684 ( .A(a[5736]), .B(c5736), .Z(n17210) );
XOR U28685 ( .A(c5737), .B(n17211), .Z(c5738) );
ANDN U28686 ( .B(n17212), .A(n17213), .Z(n17211) );
XOR U28687 ( .A(c5737), .B(b[5737]), .Z(n17212) );
XNOR U28688 ( .A(b[5737]), .B(n17213), .Z(c[5737]) );
XNOR U28689 ( .A(a[5737]), .B(c5737), .Z(n17213) );
XOR U28690 ( .A(c5738), .B(n17214), .Z(c5739) );
ANDN U28691 ( .B(n17215), .A(n17216), .Z(n17214) );
XOR U28692 ( .A(c5738), .B(b[5738]), .Z(n17215) );
XNOR U28693 ( .A(b[5738]), .B(n17216), .Z(c[5738]) );
XNOR U28694 ( .A(a[5738]), .B(c5738), .Z(n17216) );
XOR U28695 ( .A(c5739), .B(n17217), .Z(c5740) );
ANDN U28696 ( .B(n17218), .A(n17219), .Z(n17217) );
XOR U28697 ( .A(c5739), .B(b[5739]), .Z(n17218) );
XNOR U28698 ( .A(b[5739]), .B(n17219), .Z(c[5739]) );
XNOR U28699 ( .A(a[5739]), .B(c5739), .Z(n17219) );
XOR U28700 ( .A(c5740), .B(n17220), .Z(c5741) );
ANDN U28701 ( .B(n17221), .A(n17222), .Z(n17220) );
XOR U28702 ( .A(c5740), .B(b[5740]), .Z(n17221) );
XNOR U28703 ( .A(b[5740]), .B(n17222), .Z(c[5740]) );
XNOR U28704 ( .A(a[5740]), .B(c5740), .Z(n17222) );
XOR U28705 ( .A(c5741), .B(n17223), .Z(c5742) );
ANDN U28706 ( .B(n17224), .A(n17225), .Z(n17223) );
XOR U28707 ( .A(c5741), .B(b[5741]), .Z(n17224) );
XNOR U28708 ( .A(b[5741]), .B(n17225), .Z(c[5741]) );
XNOR U28709 ( .A(a[5741]), .B(c5741), .Z(n17225) );
XOR U28710 ( .A(c5742), .B(n17226), .Z(c5743) );
ANDN U28711 ( .B(n17227), .A(n17228), .Z(n17226) );
XOR U28712 ( .A(c5742), .B(b[5742]), .Z(n17227) );
XNOR U28713 ( .A(b[5742]), .B(n17228), .Z(c[5742]) );
XNOR U28714 ( .A(a[5742]), .B(c5742), .Z(n17228) );
XOR U28715 ( .A(c5743), .B(n17229), .Z(c5744) );
ANDN U28716 ( .B(n17230), .A(n17231), .Z(n17229) );
XOR U28717 ( .A(c5743), .B(b[5743]), .Z(n17230) );
XNOR U28718 ( .A(b[5743]), .B(n17231), .Z(c[5743]) );
XNOR U28719 ( .A(a[5743]), .B(c5743), .Z(n17231) );
XOR U28720 ( .A(c5744), .B(n17232), .Z(c5745) );
ANDN U28721 ( .B(n17233), .A(n17234), .Z(n17232) );
XOR U28722 ( .A(c5744), .B(b[5744]), .Z(n17233) );
XNOR U28723 ( .A(b[5744]), .B(n17234), .Z(c[5744]) );
XNOR U28724 ( .A(a[5744]), .B(c5744), .Z(n17234) );
XOR U28725 ( .A(c5745), .B(n17235), .Z(c5746) );
ANDN U28726 ( .B(n17236), .A(n17237), .Z(n17235) );
XOR U28727 ( .A(c5745), .B(b[5745]), .Z(n17236) );
XNOR U28728 ( .A(b[5745]), .B(n17237), .Z(c[5745]) );
XNOR U28729 ( .A(a[5745]), .B(c5745), .Z(n17237) );
XOR U28730 ( .A(c5746), .B(n17238), .Z(c5747) );
ANDN U28731 ( .B(n17239), .A(n17240), .Z(n17238) );
XOR U28732 ( .A(c5746), .B(b[5746]), .Z(n17239) );
XNOR U28733 ( .A(b[5746]), .B(n17240), .Z(c[5746]) );
XNOR U28734 ( .A(a[5746]), .B(c5746), .Z(n17240) );
XOR U28735 ( .A(c5747), .B(n17241), .Z(c5748) );
ANDN U28736 ( .B(n17242), .A(n17243), .Z(n17241) );
XOR U28737 ( .A(c5747), .B(b[5747]), .Z(n17242) );
XNOR U28738 ( .A(b[5747]), .B(n17243), .Z(c[5747]) );
XNOR U28739 ( .A(a[5747]), .B(c5747), .Z(n17243) );
XOR U28740 ( .A(c5748), .B(n17244), .Z(c5749) );
ANDN U28741 ( .B(n17245), .A(n17246), .Z(n17244) );
XOR U28742 ( .A(c5748), .B(b[5748]), .Z(n17245) );
XNOR U28743 ( .A(b[5748]), .B(n17246), .Z(c[5748]) );
XNOR U28744 ( .A(a[5748]), .B(c5748), .Z(n17246) );
XOR U28745 ( .A(c5749), .B(n17247), .Z(c5750) );
ANDN U28746 ( .B(n17248), .A(n17249), .Z(n17247) );
XOR U28747 ( .A(c5749), .B(b[5749]), .Z(n17248) );
XNOR U28748 ( .A(b[5749]), .B(n17249), .Z(c[5749]) );
XNOR U28749 ( .A(a[5749]), .B(c5749), .Z(n17249) );
XOR U28750 ( .A(c5750), .B(n17250), .Z(c5751) );
ANDN U28751 ( .B(n17251), .A(n17252), .Z(n17250) );
XOR U28752 ( .A(c5750), .B(b[5750]), .Z(n17251) );
XNOR U28753 ( .A(b[5750]), .B(n17252), .Z(c[5750]) );
XNOR U28754 ( .A(a[5750]), .B(c5750), .Z(n17252) );
XOR U28755 ( .A(c5751), .B(n17253), .Z(c5752) );
ANDN U28756 ( .B(n17254), .A(n17255), .Z(n17253) );
XOR U28757 ( .A(c5751), .B(b[5751]), .Z(n17254) );
XNOR U28758 ( .A(b[5751]), .B(n17255), .Z(c[5751]) );
XNOR U28759 ( .A(a[5751]), .B(c5751), .Z(n17255) );
XOR U28760 ( .A(c5752), .B(n17256), .Z(c5753) );
ANDN U28761 ( .B(n17257), .A(n17258), .Z(n17256) );
XOR U28762 ( .A(c5752), .B(b[5752]), .Z(n17257) );
XNOR U28763 ( .A(b[5752]), .B(n17258), .Z(c[5752]) );
XNOR U28764 ( .A(a[5752]), .B(c5752), .Z(n17258) );
XOR U28765 ( .A(c5753), .B(n17259), .Z(c5754) );
ANDN U28766 ( .B(n17260), .A(n17261), .Z(n17259) );
XOR U28767 ( .A(c5753), .B(b[5753]), .Z(n17260) );
XNOR U28768 ( .A(b[5753]), .B(n17261), .Z(c[5753]) );
XNOR U28769 ( .A(a[5753]), .B(c5753), .Z(n17261) );
XOR U28770 ( .A(c5754), .B(n17262), .Z(c5755) );
ANDN U28771 ( .B(n17263), .A(n17264), .Z(n17262) );
XOR U28772 ( .A(c5754), .B(b[5754]), .Z(n17263) );
XNOR U28773 ( .A(b[5754]), .B(n17264), .Z(c[5754]) );
XNOR U28774 ( .A(a[5754]), .B(c5754), .Z(n17264) );
XOR U28775 ( .A(c5755), .B(n17265), .Z(c5756) );
ANDN U28776 ( .B(n17266), .A(n17267), .Z(n17265) );
XOR U28777 ( .A(c5755), .B(b[5755]), .Z(n17266) );
XNOR U28778 ( .A(b[5755]), .B(n17267), .Z(c[5755]) );
XNOR U28779 ( .A(a[5755]), .B(c5755), .Z(n17267) );
XOR U28780 ( .A(c5756), .B(n17268), .Z(c5757) );
ANDN U28781 ( .B(n17269), .A(n17270), .Z(n17268) );
XOR U28782 ( .A(c5756), .B(b[5756]), .Z(n17269) );
XNOR U28783 ( .A(b[5756]), .B(n17270), .Z(c[5756]) );
XNOR U28784 ( .A(a[5756]), .B(c5756), .Z(n17270) );
XOR U28785 ( .A(c5757), .B(n17271), .Z(c5758) );
ANDN U28786 ( .B(n17272), .A(n17273), .Z(n17271) );
XOR U28787 ( .A(c5757), .B(b[5757]), .Z(n17272) );
XNOR U28788 ( .A(b[5757]), .B(n17273), .Z(c[5757]) );
XNOR U28789 ( .A(a[5757]), .B(c5757), .Z(n17273) );
XOR U28790 ( .A(c5758), .B(n17274), .Z(c5759) );
ANDN U28791 ( .B(n17275), .A(n17276), .Z(n17274) );
XOR U28792 ( .A(c5758), .B(b[5758]), .Z(n17275) );
XNOR U28793 ( .A(b[5758]), .B(n17276), .Z(c[5758]) );
XNOR U28794 ( .A(a[5758]), .B(c5758), .Z(n17276) );
XOR U28795 ( .A(c5759), .B(n17277), .Z(c5760) );
ANDN U28796 ( .B(n17278), .A(n17279), .Z(n17277) );
XOR U28797 ( .A(c5759), .B(b[5759]), .Z(n17278) );
XNOR U28798 ( .A(b[5759]), .B(n17279), .Z(c[5759]) );
XNOR U28799 ( .A(a[5759]), .B(c5759), .Z(n17279) );
XOR U28800 ( .A(c5760), .B(n17280), .Z(c5761) );
ANDN U28801 ( .B(n17281), .A(n17282), .Z(n17280) );
XOR U28802 ( .A(c5760), .B(b[5760]), .Z(n17281) );
XNOR U28803 ( .A(b[5760]), .B(n17282), .Z(c[5760]) );
XNOR U28804 ( .A(a[5760]), .B(c5760), .Z(n17282) );
XOR U28805 ( .A(c5761), .B(n17283), .Z(c5762) );
ANDN U28806 ( .B(n17284), .A(n17285), .Z(n17283) );
XOR U28807 ( .A(c5761), .B(b[5761]), .Z(n17284) );
XNOR U28808 ( .A(b[5761]), .B(n17285), .Z(c[5761]) );
XNOR U28809 ( .A(a[5761]), .B(c5761), .Z(n17285) );
XOR U28810 ( .A(c5762), .B(n17286), .Z(c5763) );
ANDN U28811 ( .B(n17287), .A(n17288), .Z(n17286) );
XOR U28812 ( .A(c5762), .B(b[5762]), .Z(n17287) );
XNOR U28813 ( .A(b[5762]), .B(n17288), .Z(c[5762]) );
XNOR U28814 ( .A(a[5762]), .B(c5762), .Z(n17288) );
XOR U28815 ( .A(c5763), .B(n17289), .Z(c5764) );
ANDN U28816 ( .B(n17290), .A(n17291), .Z(n17289) );
XOR U28817 ( .A(c5763), .B(b[5763]), .Z(n17290) );
XNOR U28818 ( .A(b[5763]), .B(n17291), .Z(c[5763]) );
XNOR U28819 ( .A(a[5763]), .B(c5763), .Z(n17291) );
XOR U28820 ( .A(c5764), .B(n17292), .Z(c5765) );
ANDN U28821 ( .B(n17293), .A(n17294), .Z(n17292) );
XOR U28822 ( .A(c5764), .B(b[5764]), .Z(n17293) );
XNOR U28823 ( .A(b[5764]), .B(n17294), .Z(c[5764]) );
XNOR U28824 ( .A(a[5764]), .B(c5764), .Z(n17294) );
XOR U28825 ( .A(c5765), .B(n17295), .Z(c5766) );
ANDN U28826 ( .B(n17296), .A(n17297), .Z(n17295) );
XOR U28827 ( .A(c5765), .B(b[5765]), .Z(n17296) );
XNOR U28828 ( .A(b[5765]), .B(n17297), .Z(c[5765]) );
XNOR U28829 ( .A(a[5765]), .B(c5765), .Z(n17297) );
XOR U28830 ( .A(c5766), .B(n17298), .Z(c5767) );
ANDN U28831 ( .B(n17299), .A(n17300), .Z(n17298) );
XOR U28832 ( .A(c5766), .B(b[5766]), .Z(n17299) );
XNOR U28833 ( .A(b[5766]), .B(n17300), .Z(c[5766]) );
XNOR U28834 ( .A(a[5766]), .B(c5766), .Z(n17300) );
XOR U28835 ( .A(c5767), .B(n17301), .Z(c5768) );
ANDN U28836 ( .B(n17302), .A(n17303), .Z(n17301) );
XOR U28837 ( .A(c5767), .B(b[5767]), .Z(n17302) );
XNOR U28838 ( .A(b[5767]), .B(n17303), .Z(c[5767]) );
XNOR U28839 ( .A(a[5767]), .B(c5767), .Z(n17303) );
XOR U28840 ( .A(c5768), .B(n17304), .Z(c5769) );
ANDN U28841 ( .B(n17305), .A(n17306), .Z(n17304) );
XOR U28842 ( .A(c5768), .B(b[5768]), .Z(n17305) );
XNOR U28843 ( .A(b[5768]), .B(n17306), .Z(c[5768]) );
XNOR U28844 ( .A(a[5768]), .B(c5768), .Z(n17306) );
XOR U28845 ( .A(c5769), .B(n17307), .Z(c5770) );
ANDN U28846 ( .B(n17308), .A(n17309), .Z(n17307) );
XOR U28847 ( .A(c5769), .B(b[5769]), .Z(n17308) );
XNOR U28848 ( .A(b[5769]), .B(n17309), .Z(c[5769]) );
XNOR U28849 ( .A(a[5769]), .B(c5769), .Z(n17309) );
XOR U28850 ( .A(c5770), .B(n17310), .Z(c5771) );
ANDN U28851 ( .B(n17311), .A(n17312), .Z(n17310) );
XOR U28852 ( .A(c5770), .B(b[5770]), .Z(n17311) );
XNOR U28853 ( .A(b[5770]), .B(n17312), .Z(c[5770]) );
XNOR U28854 ( .A(a[5770]), .B(c5770), .Z(n17312) );
XOR U28855 ( .A(c5771), .B(n17313), .Z(c5772) );
ANDN U28856 ( .B(n17314), .A(n17315), .Z(n17313) );
XOR U28857 ( .A(c5771), .B(b[5771]), .Z(n17314) );
XNOR U28858 ( .A(b[5771]), .B(n17315), .Z(c[5771]) );
XNOR U28859 ( .A(a[5771]), .B(c5771), .Z(n17315) );
XOR U28860 ( .A(c5772), .B(n17316), .Z(c5773) );
ANDN U28861 ( .B(n17317), .A(n17318), .Z(n17316) );
XOR U28862 ( .A(c5772), .B(b[5772]), .Z(n17317) );
XNOR U28863 ( .A(b[5772]), .B(n17318), .Z(c[5772]) );
XNOR U28864 ( .A(a[5772]), .B(c5772), .Z(n17318) );
XOR U28865 ( .A(c5773), .B(n17319), .Z(c5774) );
ANDN U28866 ( .B(n17320), .A(n17321), .Z(n17319) );
XOR U28867 ( .A(c5773), .B(b[5773]), .Z(n17320) );
XNOR U28868 ( .A(b[5773]), .B(n17321), .Z(c[5773]) );
XNOR U28869 ( .A(a[5773]), .B(c5773), .Z(n17321) );
XOR U28870 ( .A(c5774), .B(n17322), .Z(c5775) );
ANDN U28871 ( .B(n17323), .A(n17324), .Z(n17322) );
XOR U28872 ( .A(c5774), .B(b[5774]), .Z(n17323) );
XNOR U28873 ( .A(b[5774]), .B(n17324), .Z(c[5774]) );
XNOR U28874 ( .A(a[5774]), .B(c5774), .Z(n17324) );
XOR U28875 ( .A(c5775), .B(n17325), .Z(c5776) );
ANDN U28876 ( .B(n17326), .A(n17327), .Z(n17325) );
XOR U28877 ( .A(c5775), .B(b[5775]), .Z(n17326) );
XNOR U28878 ( .A(b[5775]), .B(n17327), .Z(c[5775]) );
XNOR U28879 ( .A(a[5775]), .B(c5775), .Z(n17327) );
XOR U28880 ( .A(c5776), .B(n17328), .Z(c5777) );
ANDN U28881 ( .B(n17329), .A(n17330), .Z(n17328) );
XOR U28882 ( .A(c5776), .B(b[5776]), .Z(n17329) );
XNOR U28883 ( .A(b[5776]), .B(n17330), .Z(c[5776]) );
XNOR U28884 ( .A(a[5776]), .B(c5776), .Z(n17330) );
XOR U28885 ( .A(c5777), .B(n17331), .Z(c5778) );
ANDN U28886 ( .B(n17332), .A(n17333), .Z(n17331) );
XOR U28887 ( .A(c5777), .B(b[5777]), .Z(n17332) );
XNOR U28888 ( .A(b[5777]), .B(n17333), .Z(c[5777]) );
XNOR U28889 ( .A(a[5777]), .B(c5777), .Z(n17333) );
XOR U28890 ( .A(c5778), .B(n17334), .Z(c5779) );
ANDN U28891 ( .B(n17335), .A(n17336), .Z(n17334) );
XOR U28892 ( .A(c5778), .B(b[5778]), .Z(n17335) );
XNOR U28893 ( .A(b[5778]), .B(n17336), .Z(c[5778]) );
XNOR U28894 ( .A(a[5778]), .B(c5778), .Z(n17336) );
XOR U28895 ( .A(c5779), .B(n17337), .Z(c5780) );
ANDN U28896 ( .B(n17338), .A(n17339), .Z(n17337) );
XOR U28897 ( .A(c5779), .B(b[5779]), .Z(n17338) );
XNOR U28898 ( .A(b[5779]), .B(n17339), .Z(c[5779]) );
XNOR U28899 ( .A(a[5779]), .B(c5779), .Z(n17339) );
XOR U28900 ( .A(c5780), .B(n17340), .Z(c5781) );
ANDN U28901 ( .B(n17341), .A(n17342), .Z(n17340) );
XOR U28902 ( .A(c5780), .B(b[5780]), .Z(n17341) );
XNOR U28903 ( .A(b[5780]), .B(n17342), .Z(c[5780]) );
XNOR U28904 ( .A(a[5780]), .B(c5780), .Z(n17342) );
XOR U28905 ( .A(c5781), .B(n17343), .Z(c5782) );
ANDN U28906 ( .B(n17344), .A(n17345), .Z(n17343) );
XOR U28907 ( .A(c5781), .B(b[5781]), .Z(n17344) );
XNOR U28908 ( .A(b[5781]), .B(n17345), .Z(c[5781]) );
XNOR U28909 ( .A(a[5781]), .B(c5781), .Z(n17345) );
XOR U28910 ( .A(c5782), .B(n17346), .Z(c5783) );
ANDN U28911 ( .B(n17347), .A(n17348), .Z(n17346) );
XOR U28912 ( .A(c5782), .B(b[5782]), .Z(n17347) );
XNOR U28913 ( .A(b[5782]), .B(n17348), .Z(c[5782]) );
XNOR U28914 ( .A(a[5782]), .B(c5782), .Z(n17348) );
XOR U28915 ( .A(c5783), .B(n17349), .Z(c5784) );
ANDN U28916 ( .B(n17350), .A(n17351), .Z(n17349) );
XOR U28917 ( .A(c5783), .B(b[5783]), .Z(n17350) );
XNOR U28918 ( .A(b[5783]), .B(n17351), .Z(c[5783]) );
XNOR U28919 ( .A(a[5783]), .B(c5783), .Z(n17351) );
XOR U28920 ( .A(c5784), .B(n17352), .Z(c5785) );
ANDN U28921 ( .B(n17353), .A(n17354), .Z(n17352) );
XOR U28922 ( .A(c5784), .B(b[5784]), .Z(n17353) );
XNOR U28923 ( .A(b[5784]), .B(n17354), .Z(c[5784]) );
XNOR U28924 ( .A(a[5784]), .B(c5784), .Z(n17354) );
XOR U28925 ( .A(c5785), .B(n17355), .Z(c5786) );
ANDN U28926 ( .B(n17356), .A(n17357), .Z(n17355) );
XOR U28927 ( .A(c5785), .B(b[5785]), .Z(n17356) );
XNOR U28928 ( .A(b[5785]), .B(n17357), .Z(c[5785]) );
XNOR U28929 ( .A(a[5785]), .B(c5785), .Z(n17357) );
XOR U28930 ( .A(c5786), .B(n17358), .Z(c5787) );
ANDN U28931 ( .B(n17359), .A(n17360), .Z(n17358) );
XOR U28932 ( .A(c5786), .B(b[5786]), .Z(n17359) );
XNOR U28933 ( .A(b[5786]), .B(n17360), .Z(c[5786]) );
XNOR U28934 ( .A(a[5786]), .B(c5786), .Z(n17360) );
XOR U28935 ( .A(c5787), .B(n17361), .Z(c5788) );
ANDN U28936 ( .B(n17362), .A(n17363), .Z(n17361) );
XOR U28937 ( .A(c5787), .B(b[5787]), .Z(n17362) );
XNOR U28938 ( .A(b[5787]), .B(n17363), .Z(c[5787]) );
XNOR U28939 ( .A(a[5787]), .B(c5787), .Z(n17363) );
XOR U28940 ( .A(c5788), .B(n17364), .Z(c5789) );
ANDN U28941 ( .B(n17365), .A(n17366), .Z(n17364) );
XOR U28942 ( .A(c5788), .B(b[5788]), .Z(n17365) );
XNOR U28943 ( .A(b[5788]), .B(n17366), .Z(c[5788]) );
XNOR U28944 ( .A(a[5788]), .B(c5788), .Z(n17366) );
XOR U28945 ( .A(c5789), .B(n17367), .Z(c5790) );
ANDN U28946 ( .B(n17368), .A(n17369), .Z(n17367) );
XOR U28947 ( .A(c5789), .B(b[5789]), .Z(n17368) );
XNOR U28948 ( .A(b[5789]), .B(n17369), .Z(c[5789]) );
XNOR U28949 ( .A(a[5789]), .B(c5789), .Z(n17369) );
XOR U28950 ( .A(c5790), .B(n17370), .Z(c5791) );
ANDN U28951 ( .B(n17371), .A(n17372), .Z(n17370) );
XOR U28952 ( .A(c5790), .B(b[5790]), .Z(n17371) );
XNOR U28953 ( .A(b[5790]), .B(n17372), .Z(c[5790]) );
XNOR U28954 ( .A(a[5790]), .B(c5790), .Z(n17372) );
XOR U28955 ( .A(c5791), .B(n17373), .Z(c5792) );
ANDN U28956 ( .B(n17374), .A(n17375), .Z(n17373) );
XOR U28957 ( .A(c5791), .B(b[5791]), .Z(n17374) );
XNOR U28958 ( .A(b[5791]), .B(n17375), .Z(c[5791]) );
XNOR U28959 ( .A(a[5791]), .B(c5791), .Z(n17375) );
XOR U28960 ( .A(c5792), .B(n17376), .Z(c5793) );
ANDN U28961 ( .B(n17377), .A(n17378), .Z(n17376) );
XOR U28962 ( .A(c5792), .B(b[5792]), .Z(n17377) );
XNOR U28963 ( .A(b[5792]), .B(n17378), .Z(c[5792]) );
XNOR U28964 ( .A(a[5792]), .B(c5792), .Z(n17378) );
XOR U28965 ( .A(c5793), .B(n17379), .Z(c5794) );
ANDN U28966 ( .B(n17380), .A(n17381), .Z(n17379) );
XOR U28967 ( .A(c5793), .B(b[5793]), .Z(n17380) );
XNOR U28968 ( .A(b[5793]), .B(n17381), .Z(c[5793]) );
XNOR U28969 ( .A(a[5793]), .B(c5793), .Z(n17381) );
XOR U28970 ( .A(c5794), .B(n17382), .Z(c5795) );
ANDN U28971 ( .B(n17383), .A(n17384), .Z(n17382) );
XOR U28972 ( .A(c5794), .B(b[5794]), .Z(n17383) );
XNOR U28973 ( .A(b[5794]), .B(n17384), .Z(c[5794]) );
XNOR U28974 ( .A(a[5794]), .B(c5794), .Z(n17384) );
XOR U28975 ( .A(c5795), .B(n17385), .Z(c5796) );
ANDN U28976 ( .B(n17386), .A(n17387), .Z(n17385) );
XOR U28977 ( .A(c5795), .B(b[5795]), .Z(n17386) );
XNOR U28978 ( .A(b[5795]), .B(n17387), .Z(c[5795]) );
XNOR U28979 ( .A(a[5795]), .B(c5795), .Z(n17387) );
XOR U28980 ( .A(c5796), .B(n17388), .Z(c5797) );
ANDN U28981 ( .B(n17389), .A(n17390), .Z(n17388) );
XOR U28982 ( .A(c5796), .B(b[5796]), .Z(n17389) );
XNOR U28983 ( .A(b[5796]), .B(n17390), .Z(c[5796]) );
XNOR U28984 ( .A(a[5796]), .B(c5796), .Z(n17390) );
XOR U28985 ( .A(c5797), .B(n17391), .Z(c5798) );
ANDN U28986 ( .B(n17392), .A(n17393), .Z(n17391) );
XOR U28987 ( .A(c5797), .B(b[5797]), .Z(n17392) );
XNOR U28988 ( .A(b[5797]), .B(n17393), .Z(c[5797]) );
XNOR U28989 ( .A(a[5797]), .B(c5797), .Z(n17393) );
XOR U28990 ( .A(c5798), .B(n17394), .Z(c5799) );
ANDN U28991 ( .B(n17395), .A(n17396), .Z(n17394) );
XOR U28992 ( .A(c5798), .B(b[5798]), .Z(n17395) );
XNOR U28993 ( .A(b[5798]), .B(n17396), .Z(c[5798]) );
XNOR U28994 ( .A(a[5798]), .B(c5798), .Z(n17396) );
XOR U28995 ( .A(c5799), .B(n17397), .Z(c5800) );
ANDN U28996 ( .B(n17398), .A(n17399), .Z(n17397) );
XOR U28997 ( .A(c5799), .B(b[5799]), .Z(n17398) );
XNOR U28998 ( .A(b[5799]), .B(n17399), .Z(c[5799]) );
XNOR U28999 ( .A(a[5799]), .B(c5799), .Z(n17399) );
XOR U29000 ( .A(c5800), .B(n17400), .Z(c5801) );
ANDN U29001 ( .B(n17401), .A(n17402), .Z(n17400) );
XOR U29002 ( .A(c5800), .B(b[5800]), .Z(n17401) );
XNOR U29003 ( .A(b[5800]), .B(n17402), .Z(c[5800]) );
XNOR U29004 ( .A(a[5800]), .B(c5800), .Z(n17402) );
XOR U29005 ( .A(c5801), .B(n17403), .Z(c5802) );
ANDN U29006 ( .B(n17404), .A(n17405), .Z(n17403) );
XOR U29007 ( .A(c5801), .B(b[5801]), .Z(n17404) );
XNOR U29008 ( .A(b[5801]), .B(n17405), .Z(c[5801]) );
XNOR U29009 ( .A(a[5801]), .B(c5801), .Z(n17405) );
XOR U29010 ( .A(c5802), .B(n17406), .Z(c5803) );
ANDN U29011 ( .B(n17407), .A(n17408), .Z(n17406) );
XOR U29012 ( .A(c5802), .B(b[5802]), .Z(n17407) );
XNOR U29013 ( .A(b[5802]), .B(n17408), .Z(c[5802]) );
XNOR U29014 ( .A(a[5802]), .B(c5802), .Z(n17408) );
XOR U29015 ( .A(c5803), .B(n17409), .Z(c5804) );
ANDN U29016 ( .B(n17410), .A(n17411), .Z(n17409) );
XOR U29017 ( .A(c5803), .B(b[5803]), .Z(n17410) );
XNOR U29018 ( .A(b[5803]), .B(n17411), .Z(c[5803]) );
XNOR U29019 ( .A(a[5803]), .B(c5803), .Z(n17411) );
XOR U29020 ( .A(c5804), .B(n17412), .Z(c5805) );
ANDN U29021 ( .B(n17413), .A(n17414), .Z(n17412) );
XOR U29022 ( .A(c5804), .B(b[5804]), .Z(n17413) );
XNOR U29023 ( .A(b[5804]), .B(n17414), .Z(c[5804]) );
XNOR U29024 ( .A(a[5804]), .B(c5804), .Z(n17414) );
XOR U29025 ( .A(c5805), .B(n17415), .Z(c5806) );
ANDN U29026 ( .B(n17416), .A(n17417), .Z(n17415) );
XOR U29027 ( .A(c5805), .B(b[5805]), .Z(n17416) );
XNOR U29028 ( .A(b[5805]), .B(n17417), .Z(c[5805]) );
XNOR U29029 ( .A(a[5805]), .B(c5805), .Z(n17417) );
XOR U29030 ( .A(c5806), .B(n17418), .Z(c5807) );
ANDN U29031 ( .B(n17419), .A(n17420), .Z(n17418) );
XOR U29032 ( .A(c5806), .B(b[5806]), .Z(n17419) );
XNOR U29033 ( .A(b[5806]), .B(n17420), .Z(c[5806]) );
XNOR U29034 ( .A(a[5806]), .B(c5806), .Z(n17420) );
XOR U29035 ( .A(c5807), .B(n17421), .Z(c5808) );
ANDN U29036 ( .B(n17422), .A(n17423), .Z(n17421) );
XOR U29037 ( .A(c5807), .B(b[5807]), .Z(n17422) );
XNOR U29038 ( .A(b[5807]), .B(n17423), .Z(c[5807]) );
XNOR U29039 ( .A(a[5807]), .B(c5807), .Z(n17423) );
XOR U29040 ( .A(c5808), .B(n17424), .Z(c5809) );
ANDN U29041 ( .B(n17425), .A(n17426), .Z(n17424) );
XOR U29042 ( .A(c5808), .B(b[5808]), .Z(n17425) );
XNOR U29043 ( .A(b[5808]), .B(n17426), .Z(c[5808]) );
XNOR U29044 ( .A(a[5808]), .B(c5808), .Z(n17426) );
XOR U29045 ( .A(c5809), .B(n17427), .Z(c5810) );
ANDN U29046 ( .B(n17428), .A(n17429), .Z(n17427) );
XOR U29047 ( .A(c5809), .B(b[5809]), .Z(n17428) );
XNOR U29048 ( .A(b[5809]), .B(n17429), .Z(c[5809]) );
XNOR U29049 ( .A(a[5809]), .B(c5809), .Z(n17429) );
XOR U29050 ( .A(c5810), .B(n17430), .Z(c5811) );
ANDN U29051 ( .B(n17431), .A(n17432), .Z(n17430) );
XOR U29052 ( .A(c5810), .B(b[5810]), .Z(n17431) );
XNOR U29053 ( .A(b[5810]), .B(n17432), .Z(c[5810]) );
XNOR U29054 ( .A(a[5810]), .B(c5810), .Z(n17432) );
XOR U29055 ( .A(c5811), .B(n17433), .Z(c5812) );
ANDN U29056 ( .B(n17434), .A(n17435), .Z(n17433) );
XOR U29057 ( .A(c5811), .B(b[5811]), .Z(n17434) );
XNOR U29058 ( .A(b[5811]), .B(n17435), .Z(c[5811]) );
XNOR U29059 ( .A(a[5811]), .B(c5811), .Z(n17435) );
XOR U29060 ( .A(c5812), .B(n17436), .Z(c5813) );
ANDN U29061 ( .B(n17437), .A(n17438), .Z(n17436) );
XOR U29062 ( .A(c5812), .B(b[5812]), .Z(n17437) );
XNOR U29063 ( .A(b[5812]), .B(n17438), .Z(c[5812]) );
XNOR U29064 ( .A(a[5812]), .B(c5812), .Z(n17438) );
XOR U29065 ( .A(c5813), .B(n17439), .Z(c5814) );
ANDN U29066 ( .B(n17440), .A(n17441), .Z(n17439) );
XOR U29067 ( .A(c5813), .B(b[5813]), .Z(n17440) );
XNOR U29068 ( .A(b[5813]), .B(n17441), .Z(c[5813]) );
XNOR U29069 ( .A(a[5813]), .B(c5813), .Z(n17441) );
XOR U29070 ( .A(c5814), .B(n17442), .Z(c5815) );
ANDN U29071 ( .B(n17443), .A(n17444), .Z(n17442) );
XOR U29072 ( .A(c5814), .B(b[5814]), .Z(n17443) );
XNOR U29073 ( .A(b[5814]), .B(n17444), .Z(c[5814]) );
XNOR U29074 ( .A(a[5814]), .B(c5814), .Z(n17444) );
XOR U29075 ( .A(c5815), .B(n17445), .Z(c5816) );
ANDN U29076 ( .B(n17446), .A(n17447), .Z(n17445) );
XOR U29077 ( .A(c5815), .B(b[5815]), .Z(n17446) );
XNOR U29078 ( .A(b[5815]), .B(n17447), .Z(c[5815]) );
XNOR U29079 ( .A(a[5815]), .B(c5815), .Z(n17447) );
XOR U29080 ( .A(c5816), .B(n17448), .Z(c5817) );
ANDN U29081 ( .B(n17449), .A(n17450), .Z(n17448) );
XOR U29082 ( .A(c5816), .B(b[5816]), .Z(n17449) );
XNOR U29083 ( .A(b[5816]), .B(n17450), .Z(c[5816]) );
XNOR U29084 ( .A(a[5816]), .B(c5816), .Z(n17450) );
XOR U29085 ( .A(c5817), .B(n17451), .Z(c5818) );
ANDN U29086 ( .B(n17452), .A(n17453), .Z(n17451) );
XOR U29087 ( .A(c5817), .B(b[5817]), .Z(n17452) );
XNOR U29088 ( .A(b[5817]), .B(n17453), .Z(c[5817]) );
XNOR U29089 ( .A(a[5817]), .B(c5817), .Z(n17453) );
XOR U29090 ( .A(c5818), .B(n17454), .Z(c5819) );
ANDN U29091 ( .B(n17455), .A(n17456), .Z(n17454) );
XOR U29092 ( .A(c5818), .B(b[5818]), .Z(n17455) );
XNOR U29093 ( .A(b[5818]), .B(n17456), .Z(c[5818]) );
XNOR U29094 ( .A(a[5818]), .B(c5818), .Z(n17456) );
XOR U29095 ( .A(c5819), .B(n17457), .Z(c5820) );
ANDN U29096 ( .B(n17458), .A(n17459), .Z(n17457) );
XOR U29097 ( .A(c5819), .B(b[5819]), .Z(n17458) );
XNOR U29098 ( .A(b[5819]), .B(n17459), .Z(c[5819]) );
XNOR U29099 ( .A(a[5819]), .B(c5819), .Z(n17459) );
XOR U29100 ( .A(c5820), .B(n17460), .Z(c5821) );
ANDN U29101 ( .B(n17461), .A(n17462), .Z(n17460) );
XOR U29102 ( .A(c5820), .B(b[5820]), .Z(n17461) );
XNOR U29103 ( .A(b[5820]), .B(n17462), .Z(c[5820]) );
XNOR U29104 ( .A(a[5820]), .B(c5820), .Z(n17462) );
XOR U29105 ( .A(c5821), .B(n17463), .Z(c5822) );
ANDN U29106 ( .B(n17464), .A(n17465), .Z(n17463) );
XOR U29107 ( .A(c5821), .B(b[5821]), .Z(n17464) );
XNOR U29108 ( .A(b[5821]), .B(n17465), .Z(c[5821]) );
XNOR U29109 ( .A(a[5821]), .B(c5821), .Z(n17465) );
XOR U29110 ( .A(c5822), .B(n17466), .Z(c5823) );
ANDN U29111 ( .B(n17467), .A(n17468), .Z(n17466) );
XOR U29112 ( .A(c5822), .B(b[5822]), .Z(n17467) );
XNOR U29113 ( .A(b[5822]), .B(n17468), .Z(c[5822]) );
XNOR U29114 ( .A(a[5822]), .B(c5822), .Z(n17468) );
XOR U29115 ( .A(c5823), .B(n17469), .Z(c5824) );
ANDN U29116 ( .B(n17470), .A(n17471), .Z(n17469) );
XOR U29117 ( .A(c5823), .B(b[5823]), .Z(n17470) );
XNOR U29118 ( .A(b[5823]), .B(n17471), .Z(c[5823]) );
XNOR U29119 ( .A(a[5823]), .B(c5823), .Z(n17471) );
XOR U29120 ( .A(c5824), .B(n17472), .Z(c5825) );
ANDN U29121 ( .B(n17473), .A(n17474), .Z(n17472) );
XOR U29122 ( .A(c5824), .B(b[5824]), .Z(n17473) );
XNOR U29123 ( .A(b[5824]), .B(n17474), .Z(c[5824]) );
XNOR U29124 ( .A(a[5824]), .B(c5824), .Z(n17474) );
XOR U29125 ( .A(c5825), .B(n17475), .Z(c5826) );
ANDN U29126 ( .B(n17476), .A(n17477), .Z(n17475) );
XOR U29127 ( .A(c5825), .B(b[5825]), .Z(n17476) );
XNOR U29128 ( .A(b[5825]), .B(n17477), .Z(c[5825]) );
XNOR U29129 ( .A(a[5825]), .B(c5825), .Z(n17477) );
XOR U29130 ( .A(c5826), .B(n17478), .Z(c5827) );
ANDN U29131 ( .B(n17479), .A(n17480), .Z(n17478) );
XOR U29132 ( .A(c5826), .B(b[5826]), .Z(n17479) );
XNOR U29133 ( .A(b[5826]), .B(n17480), .Z(c[5826]) );
XNOR U29134 ( .A(a[5826]), .B(c5826), .Z(n17480) );
XOR U29135 ( .A(c5827), .B(n17481), .Z(c5828) );
ANDN U29136 ( .B(n17482), .A(n17483), .Z(n17481) );
XOR U29137 ( .A(c5827), .B(b[5827]), .Z(n17482) );
XNOR U29138 ( .A(b[5827]), .B(n17483), .Z(c[5827]) );
XNOR U29139 ( .A(a[5827]), .B(c5827), .Z(n17483) );
XOR U29140 ( .A(c5828), .B(n17484), .Z(c5829) );
ANDN U29141 ( .B(n17485), .A(n17486), .Z(n17484) );
XOR U29142 ( .A(c5828), .B(b[5828]), .Z(n17485) );
XNOR U29143 ( .A(b[5828]), .B(n17486), .Z(c[5828]) );
XNOR U29144 ( .A(a[5828]), .B(c5828), .Z(n17486) );
XOR U29145 ( .A(c5829), .B(n17487), .Z(c5830) );
ANDN U29146 ( .B(n17488), .A(n17489), .Z(n17487) );
XOR U29147 ( .A(c5829), .B(b[5829]), .Z(n17488) );
XNOR U29148 ( .A(b[5829]), .B(n17489), .Z(c[5829]) );
XNOR U29149 ( .A(a[5829]), .B(c5829), .Z(n17489) );
XOR U29150 ( .A(c5830), .B(n17490), .Z(c5831) );
ANDN U29151 ( .B(n17491), .A(n17492), .Z(n17490) );
XOR U29152 ( .A(c5830), .B(b[5830]), .Z(n17491) );
XNOR U29153 ( .A(b[5830]), .B(n17492), .Z(c[5830]) );
XNOR U29154 ( .A(a[5830]), .B(c5830), .Z(n17492) );
XOR U29155 ( .A(c5831), .B(n17493), .Z(c5832) );
ANDN U29156 ( .B(n17494), .A(n17495), .Z(n17493) );
XOR U29157 ( .A(c5831), .B(b[5831]), .Z(n17494) );
XNOR U29158 ( .A(b[5831]), .B(n17495), .Z(c[5831]) );
XNOR U29159 ( .A(a[5831]), .B(c5831), .Z(n17495) );
XOR U29160 ( .A(c5832), .B(n17496), .Z(c5833) );
ANDN U29161 ( .B(n17497), .A(n17498), .Z(n17496) );
XOR U29162 ( .A(c5832), .B(b[5832]), .Z(n17497) );
XNOR U29163 ( .A(b[5832]), .B(n17498), .Z(c[5832]) );
XNOR U29164 ( .A(a[5832]), .B(c5832), .Z(n17498) );
XOR U29165 ( .A(c5833), .B(n17499), .Z(c5834) );
ANDN U29166 ( .B(n17500), .A(n17501), .Z(n17499) );
XOR U29167 ( .A(c5833), .B(b[5833]), .Z(n17500) );
XNOR U29168 ( .A(b[5833]), .B(n17501), .Z(c[5833]) );
XNOR U29169 ( .A(a[5833]), .B(c5833), .Z(n17501) );
XOR U29170 ( .A(c5834), .B(n17502), .Z(c5835) );
ANDN U29171 ( .B(n17503), .A(n17504), .Z(n17502) );
XOR U29172 ( .A(c5834), .B(b[5834]), .Z(n17503) );
XNOR U29173 ( .A(b[5834]), .B(n17504), .Z(c[5834]) );
XNOR U29174 ( .A(a[5834]), .B(c5834), .Z(n17504) );
XOR U29175 ( .A(c5835), .B(n17505), .Z(c5836) );
ANDN U29176 ( .B(n17506), .A(n17507), .Z(n17505) );
XOR U29177 ( .A(c5835), .B(b[5835]), .Z(n17506) );
XNOR U29178 ( .A(b[5835]), .B(n17507), .Z(c[5835]) );
XNOR U29179 ( .A(a[5835]), .B(c5835), .Z(n17507) );
XOR U29180 ( .A(c5836), .B(n17508), .Z(c5837) );
ANDN U29181 ( .B(n17509), .A(n17510), .Z(n17508) );
XOR U29182 ( .A(c5836), .B(b[5836]), .Z(n17509) );
XNOR U29183 ( .A(b[5836]), .B(n17510), .Z(c[5836]) );
XNOR U29184 ( .A(a[5836]), .B(c5836), .Z(n17510) );
XOR U29185 ( .A(c5837), .B(n17511), .Z(c5838) );
ANDN U29186 ( .B(n17512), .A(n17513), .Z(n17511) );
XOR U29187 ( .A(c5837), .B(b[5837]), .Z(n17512) );
XNOR U29188 ( .A(b[5837]), .B(n17513), .Z(c[5837]) );
XNOR U29189 ( .A(a[5837]), .B(c5837), .Z(n17513) );
XOR U29190 ( .A(c5838), .B(n17514), .Z(c5839) );
ANDN U29191 ( .B(n17515), .A(n17516), .Z(n17514) );
XOR U29192 ( .A(c5838), .B(b[5838]), .Z(n17515) );
XNOR U29193 ( .A(b[5838]), .B(n17516), .Z(c[5838]) );
XNOR U29194 ( .A(a[5838]), .B(c5838), .Z(n17516) );
XOR U29195 ( .A(c5839), .B(n17517), .Z(c5840) );
ANDN U29196 ( .B(n17518), .A(n17519), .Z(n17517) );
XOR U29197 ( .A(c5839), .B(b[5839]), .Z(n17518) );
XNOR U29198 ( .A(b[5839]), .B(n17519), .Z(c[5839]) );
XNOR U29199 ( .A(a[5839]), .B(c5839), .Z(n17519) );
XOR U29200 ( .A(c5840), .B(n17520), .Z(c5841) );
ANDN U29201 ( .B(n17521), .A(n17522), .Z(n17520) );
XOR U29202 ( .A(c5840), .B(b[5840]), .Z(n17521) );
XNOR U29203 ( .A(b[5840]), .B(n17522), .Z(c[5840]) );
XNOR U29204 ( .A(a[5840]), .B(c5840), .Z(n17522) );
XOR U29205 ( .A(c5841), .B(n17523), .Z(c5842) );
ANDN U29206 ( .B(n17524), .A(n17525), .Z(n17523) );
XOR U29207 ( .A(c5841), .B(b[5841]), .Z(n17524) );
XNOR U29208 ( .A(b[5841]), .B(n17525), .Z(c[5841]) );
XNOR U29209 ( .A(a[5841]), .B(c5841), .Z(n17525) );
XOR U29210 ( .A(c5842), .B(n17526), .Z(c5843) );
ANDN U29211 ( .B(n17527), .A(n17528), .Z(n17526) );
XOR U29212 ( .A(c5842), .B(b[5842]), .Z(n17527) );
XNOR U29213 ( .A(b[5842]), .B(n17528), .Z(c[5842]) );
XNOR U29214 ( .A(a[5842]), .B(c5842), .Z(n17528) );
XOR U29215 ( .A(c5843), .B(n17529), .Z(c5844) );
ANDN U29216 ( .B(n17530), .A(n17531), .Z(n17529) );
XOR U29217 ( .A(c5843), .B(b[5843]), .Z(n17530) );
XNOR U29218 ( .A(b[5843]), .B(n17531), .Z(c[5843]) );
XNOR U29219 ( .A(a[5843]), .B(c5843), .Z(n17531) );
XOR U29220 ( .A(c5844), .B(n17532), .Z(c5845) );
ANDN U29221 ( .B(n17533), .A(n17534), .Z(n17532) );
XOR U29222 ( .A(c5844), .B(b[5844]), .Z(n17533) );
XNOR U29223 ( .A(b[5844]), .B(n17534), .Z(c[5844]) );
XNOR U29224 ( .A(a[5844]), .B(c5844), .Z(n17534) );
XOR U29225 ( .A(c5845), .B(n17535), .Z(c5846) );
ANDN U29226 ( .B(n17536), .A(n17537), .Z(n17535) );
XOR U29227 ( .A(c5845), .B(b[5845]), .Z(n17536) );
XNOR U29228 ( .A(b[5845]), .B(n17537), .Z(c[5845]) );
XNOR U29229 ( .A(a[5845]), .B(c5845), .Z(n17537) );
XOR U29230 ( .A(c5846), .B(n17538), .Z(c5847) );
ANDN U29231 ( .B(n17539), .A(n17540), .Z(n17538) );
XOR U29232 ( .A(c5846), .B(b[5846]), .Z(n17539) );
XNOR U29233 ( .A(b[5846]), .B(n17540), .Z(c[5846]) );
XNOR U29234 ( .A(a[5846]), .B(c5846), .Z(n17540) );
XOR U29235 ( .A(c5847), .B(n17541), .Z(c5848) );
ANDN U29236 ( .B(n17542), .A(n17543), .Z(n17541) );
XOR U29237 ( .A(c5847), .B(b[5847]), .Z(n17542) );
XNOR U29238 ( .A(b[5847]), .B(n17543), .Z(c[5847]) );
XNOR U29239 ( .A(a[5847]), .B(c5847), .Z(n17543) );
XOR U29240 ( .A(c5848), .B(n17544), .Z(c5849) );
ANDN U29241 ( .B(n17545), .A(n17546), .Z(n17544) );
XOR U29242 ( .A(c5848), .B(b[5848]), .Z(n17545) );
XNOR U29243 ( .A(b[5848]), .B(n17546), .Z(c[5848]) );
XNOR U29244 ( .A(a[5848]), .B(c5848), .Z(n17546) );
XOR U29245 ( .A(c5849), .B(n17547), .Z(c5850) );
ANDN U29246 ( .B(n17548), .A(n17549), .Z(n17547) );
XOR U29247 ( .A(c5849), .B(b[5849]), .Z(n17548) );
XNOR U29248 ( .A(b[5849]), .B(n17549), .Z(c[5849]) );
XNOR U29249 ( .A(a[5849]), .B(c5849), .Z(n17549) );
XOR U29250 ( .A(c5850), .B(n17550), .Z(c5851) );
ANDN U29251 ( .B(n17551), .A(n17552), .Z(n17550) );
XOR U29252 ( .A(c5850), .B(b[5850]), .Z(n17551) );
XNOR U29253 ( .A(b[5850]), .B(n17552), .Z(c[5850]) );
XNOR U29254 ( .A(a[5850]), .B(c5850), .Z(n17552) );
XOR U29255 ( .A(c5851), .B(n17553), .Z(c5852) );
ANDN U29256 ( .B(n17554), .A(n17555), .Z(n17553) );
XOR U29257 ( .A(c5851), .B(b[5851]), .Z(n17554) );
XNOR U29258 ( .A(b[5851]), .B(n17555), .Z(c[5851]) );
XNOR U29259 ( .A(a[5851]), .B(c5851), .Z(n17555) );
XOR U29260 ( .A(c5852), .B(n17556), .Z(c5853) );
ANDN U29261 ( .B(n17557), .A(n17558), .Z(n17556) );
XOR U29262 ( .A(c5852), .B(b[5852]), .Z(n17557) );
XNOR U29263 ( .A(b[5852]), .B(n17558), .Z(c[5852]) );
XNOR U29264 ( .A(a[5852]), .B(c5852), .Z(n17558) );
XOR U29265 ( .A(c5853), .B(n17559), .Z(c5854) );
ANDN U29266 ( .B(n17560), .A(n17561), .Z(n17559) );
XOR U29267 ( .A(c5853), .B(b[5853]), .Z(n17560) );
XNOR U29268 ( .A(b[5853]), .B(n17561), .Z(c[5853]) );
XNOR U29269 ( .A(a[5853]), .B(c5853), .Z(n17561) );
XOR U29270 ( .A(c5854), .B(n17562), .Z(c5855) );
ANDN U29271 ( .B(n17563), .A(n17564), .Z(n17562) );
XOR U29272 ( .A(c5854), .B(b[5854]), .Z(n17563) );
XNOR U29273 ( .A(b[5854]), .B(n17564), .Z(c[5854]) );
XNOR U29274 ( .A(a[5854]), .B(c5854), .Z(n17564) );
XOR U29275 ( .A(c5855), .B(n17565), .Z(c5856) );
ANDN U29276 ( .B(n17566), .A(n17567), .Z(n17565) );
XOR U29277 ( .A(c5855), .B(b[5855]), .Z(n17566) );
XNOR U29278 ( .A(b[5855]), .B(n17567), .Z(c[5855]) );
XNOR U29279 ( .A(a[5855]), .B(c5855), .Z(n17567) );
XOR U29280 ( .A(c5856), .B(n17568), .Z(c5857) );
ANDN U29281 ( .B(n17569), .A(n17570), .Z(n17568) );
XOR U29282 ( .A(c5856), .B(b[5856]), .Z(n17569) );
XNOR U29283 ( .A(b[5856]), .B(n17570), .Z(c[5856]) );
XNOR U29284 ( .A(a[5856]), .B(c5856), .Z(n17570) );
XOR U29285 ( .A(c5857), .B(n17571), .Z(c5858) );
ANDN U29286 ( .B(n17572), .A(n17573), .Z(n17571) );
XOR U29287 ( .A(c5857), .B(b[5857]), .Z(n17572) );
XNOR U29288 ( .A(b[5857]), .B(n17573), .Z(c[5857]) );
XNOR U29289 ( .A(a[5857]), .B(c5857), .Z(n17573) );
XOR U29290 ( .A(c5858), .B(n17574), .Z(c5859) );
ANDN U29291 ( .B(n17575), .A(n17576), .Z(n17574) );
XOR U29292 ( .A(c5858), .B(b[5858]), .Z(n17575) );
XNOR U29293 ( .A(b[5858]), .B(n17576), .Z(c[5858]) );
XNOR U29294 ( .A(a[5858]), .B(c5858), .Z(n17576) );
XOR U29295 ( .A(c5859), .B(n17577), .Z(c5860) );
ANDN U29296 ( .B(n17578), .A(n17579), .Z(n17577) );
XOR U29297 ( .A(c5859), .B(b[5859]), .Z(n17578) );
XNOR U29298 ( .A(b[5859]), .B(n17579), .Z(c[5859]) );
XNOR U29299 ( .A(a[5859]), .B(c5859), .Z(n17579) );
XOR U29300 ( .A(c5860), .B(n17580), .Z(c5861) );
ANDN U29301 ( .B(n17581), .A(n17582), .Z(n17580) );
XOR U29302 ( .A(c5860), .B(b[5860]), .Z(n17581) );
XNOR U29303 ( .A(b[5860]), .B(n17582), .Z(c[5860]) );
XNOR U29304 ( .A(a[5860]), .B(c5860), .Z(n17582) );
XOR U29305 ( .A(c5861), .B(n17583), .Z(c5862) );
ANDN U29306 ( .B(n17584), .A(n17585), .Z(n17583) );
XOR U29307 ( .A(c5861), .B(b[5861]), .Z(n17584) );
XNOR U29308 ( .A(b[5861]), .B(n17585), .Z(c[5861]) );
XNOR U29309 ( .A(a[5861]), .B(c5861), .Z(n17585) );
XOR U29310 ( .A(c5862), .B(n17586), .Z(c5863) );
ANDN U29311 ( .B(n17587), .A(n17588), .Z(n17586) );
XOR U29312 ( .A(c5862), .B(b[5862]), .Z(n17587) );
XNOR U29313 ( .A(b[5862]), .B(n17588), .Z(c[5862]) );
XNOR U29314 ( .A(a[5862]), .B(c5862), .Z(n17588) );
XOR U29315 ( .A(c5863), .B(n17589), .Z(c5864) );
ANDN U29316 ( .B(n17590), .A(n17591), .Z(n17589) );
XOR U29317 ( .A(c5863), .B(b[5863]), .Z(n17590) );
XNOR U29318 ( .A(b[5863]), .B(n17591), .Z(c[5863]) );
XNOR U29319 ( .A(a[5863]), .B(c5863), .Z(n17591) );
XOR U29320 ( .A(c5864), .B(n17592), .Z(c5865) );
ANDN U29321 ( .B(n17593), .A(n17594), .Z(n17592) );
XOR U29322 ( .A(c5864), .B(b[5864]), .Z(n17593) );
XNOR U29323 ( .A(b[5864]), .B(n17594), .Z(c[5864]) );
XNOR U29324 ( .A(a[5864]), .B(c5864), .Z(n17594) );
XOR U29325 ( .A(c5865), .B(n17595), .Z(c5866) );
ANDN U29326 ( .B(n17596), .A(n17597), .Z(n17595) );
XOR U29327 ( .A(c5865), .B(b[5865]), .Z(n17596) );
XNOR U29328 ( .A(b[5865]), .B(n17597), .Z(c[5865]) );
XNOR U29329 ( .A(a[5865]), .B(c5865), .Z(n17597) );
XOR U29330 ( .A(c5866), .B(n17598), .Z(c5867) );
ANDN U29331 ( .B(n17599), .A(n17600), .Z(n17598) );
XOR U29332 ( .A(c5866), .B(b[5866]), .Z(n17599) );
XNOR U29333 ( .A(b[5866]), .B(n17600), .Z(c[5866]) );
XNOR U29334 ( .A(a[5866]), .B(c5866), .Z(n17600) );
XOR U29335 ( .A(c5867), .B(n17601), .Z(c5868) );
ANDN U29336 ( .B(n17602), .A(n17603), .Z(n17601) );
XOR U29337 ( .A(c5867), .B(b[5867]), .Z(n17602) );
XNOR U29338 ( .A(b[5867]), .B(n17603), .Z(c[5867]) );
XNOR U29339 ( .A(a[5867]), .B(c5867), .Z(n17603) );
XOR U29340 ( .A(c5868), .B(n17604), .Z(c5869) );
ANDN U29341 ( .B(n17605), .A(n17606), .Z(n17604) );
XOR U29342 ( .A(c5868), .B(b[5868]), .Z(n17605) );
XNOR U29343 ( .A(b[5868]), .B(n17606), .Z(c[5868]) );
XNOR U29344 ( .A(a[5868]), .B(c5868), .Z(n17606) );
XOR U29345 ( .A(c5869), .B(n17607), .Z(c5870) );
ANDN U29346 ( .B(n17608), .A(n17609), .Z(n17607) );
XOR U29347 ( .A(c5869), .B(b[5869]), .Z(n17608) );
XNOR U29348 ( .A(b[5869]), .B(n17609), .Z(c[5869]) );
XNOR U29349 ( .A(a[5869]), .B(c5869), .Z(n17609) );
XOR U29350 ( .A(c5870), .B(n17610), .Z(c5871) );
ANDN U29351 ( .B(n17611), .A(n17612), .Z(n17610) );
XOR U29352 ( .A(c5870), .B(b[5870]), .Z(n17611) );
XNOR U29353 ( .A(b[5870]), .B(n17612), .Z(c[5870]) );
XNOR U29354 ( .A(a[5870]), .B(c5870), .Z(n17612) );
XOR U29355 ( .A(c5871), .B(n17613), .Z(c5872) );
ANDN U29356 ( .B(n17614), .A(n17615), .Z(n17613) );
XOR U29357 ( .A(c5871), .B(b[5871]), .Z(n17614) );
XNOR U29358 ( .A(b[5871]), .B(n17615), .Z(c[5871]) );
XNOR U29359 ( .A(a[5871]), .B(c5871), .Z(n17615) );
XOR U29360 ( .A(c5872), .B(n17616), .Z(c5873) );
ANDN U29361 ( .B(n17617), .A(n17618), .Z(n17616) );
XOR U29362 ( .A(c5872), .B(b[5872]), .Z(n17617) );
XNOR U29363 ( .A(b[5872]), .B(n17618), .Z(c[5872]) );
XNOR U29364 ( .A(a[5872]), .B(c5872), .Z(n17618) );
XOR U29365 ( .A(c5873), .B(n17619), .Z(c5874) );
ANDN U29366 ( .B(n17620), .A(n17621), .Z(n17619) );
XOR U29367 ( .A(c5873), .B(b[5873]), .Z(n17620) );
XNOR U29368 ( .A(b[5873]), .B(n17621), .Z(c[5873]) );
XNOR U29369 ( .A(a[5873]), .B(c5873), .Z(n17621) );
XOR U29370 ( .A(c5874), .B(n17622), .Z(c5875) );
ANDN U29371 ( .B(n17623), .A(n17624), .Z(n17622) );
XOR U29372 ( .A(c5874), .B(b[5874]), .Z(n17623) );
XNOR U29373 ( .A(b[5874]), .B(n17624), .Z(c[5874]) );
XNOR U29374 ( .A(a[5874]), .B(c5874), .Z(n17624) );
XOR U29375 ( .A(c5875), .B(n17625), .Z(c5876) );
ANDN U29376 ( .B(n17626), .A(n17627), .Z(n17625) );
XOR U29377 ( .A(c5875), .B(b[5875]), .Z(n17626) );
XNOR U29378 ( .A(b[5875]), .B(n17627), .Z(c[5875]) );
XNOR U29379 ( .A(a[5875]), .B(c5875), .Z(n17627) );
XOR U29380 ( .A(c5876), .B(n17628), .Z(c5877) );
ANDN U29381 ( .B(n17629), .A(n17630), .Z(n17628) );
XOR U29382 ( .A(c5876), .B(b[5876]), .Z(n17629) );
XNOR U29383 ( .A(b[5876]), .B(n17630), .Z(c[5876]) );
XNOR U29384 ( .A(a[5876]), .B(c5876), .Z(n17630) );
XOR U29385 ( .A(c5877), .B(n17631), .Z(c5878) );
ANDN U29386 ( .B(n17632), .A(n17633), .Z(n17631) );
XOR U29387 ( .A(c5877), .B(b[5877]), .Z(n17632) );
XNOR U29388 ( .A(b[5877]), .B(n17633), .Z(c[5877]) );
XNOR U29389 ( .A(a[5877]), .B(c5877), .Z(n17633) );
XOR U29390 ( .A(c5878), .B(n17634), .Z(c5879) );
ANDN U29391 ( .B(n17635), .A(n17636), .Z(n17634) );
XOR U29392 ( .A(c5878), .B(b[5878]), .Z(n17635) );
XNOR U29393 ( .A(b[5878]), .B(n17636), .Z(c[5878]) );
XNOR U29394 ( .A(a[5878]), .B(c5878), .Z(n17636) );
XOR U29395 ( .A(c5879), .B(n17637), .Z(c5880) );
ANDN U29396 ( .B(n17638), .A(n17639), .Z(n17637) );
XOR U29397 ( .A(c5879), .B(b[5879]), .Z(n17638) );
XNOR U29398 ( .A(b[5879]), .B(n17639), .Z(c[5879]) );
XNOR U29399 ( .A(a[5879]), .B(c5879), .Z(n17639) );
XOR U29400 ( .A(c5880), .B(n17640), .Z(c5881) );
ANDN U29401 ( .B(n17641), .A(n17642), .Z(n17640) );
XOR U29402 ( .A(c5880), .B(b[5880]), .Z(n17641) );
XNOR U29403 ( .A(b[5880]), .B(n17642), .Z(c[5880]) );
XNOR U29404 ( .A(a[5880]), .B(c5880), .Z(n17642) );
XOR U29405 ( .A(c5881), .B(n17643), .Z(c5882) );
ANDN U29406 ( .B(n17644), .A(n17645), .Z(n17643) );
XOR U29407 ( .A(c5881), .B(b[5881]), .Z(n17644) );
XNOR U29408 ( .A(b[5881]), .B(n17645), .Z(c[5881]) );
XNOR U29409 ( .A(a[5881]), .B(c5881), .Z(n17645) );
XOR U29410 ( .A(c5882), .B(n17646), .Z(c5883) );
ANDN U29411 ( .B(n17647), .A(n17648), .Z(n17646) );
XOR U29412 ( .A(c5882), .B(b[5882]), .Z(n17647) );
XNOR U29413 ( .A(b[5882]), .B(n17648), .Z(c[5882]) );
XNOR U29414 ( .A(a[5882]), .B(c5882), .Z(n17648) );
XOR U29415 ( .A(c5883), .B(n17649), .Z(c5884) );
ANDN U29416 ( .B(n17650), .A(n17651), .Z(n17649) );
XOR U29417 ( .A(c5883), .B(b[5883]), .Z(n17650) );
XNOR U29418 ( .A(b[5883]), .B(n17651), .Z(c[5883]) );
XNOR U29419 ( .A(a[5883]), .B(c5883), .Z(n17651) );
XOR U29420 ( .A(c5884), .B(n17652), .Z(c5885) );
ANDN U29421 ( .B(n17653), .A(n17654), .Z(n17652) );
XOR U29422 ( .A(c5884), .B(b[5884]), .Z(n17653) );
XNOR U29423 ( .A(b[5884]), .B(n17654), .Z(c[5884]) );
XNOR U29424 ( .A(a[5884]), .B(c5884), .Z(n17654) );
XOR U29425 ( .A(c5885), .B(n17655), .Z(c5886) );
ANDN U29426 ( .B(n17656), .A(n17657), .Z(n17655) );
XOR U29427 ( .A(c5885), .B(b[5885]), .Z(n17656) );
XNOR U29428 ( .A(b[5885]), .B(n17657), .Z(c[5885]) );
XNOR U29429 ( .A(a[5885]), .B(c5885), .Z(n17657) );
XOR U29430 ( .A(c5886), .B(n17658), .Z(c5887) );
ANDN U29431 ( .B(n17659), .A(n17660), .Z(n17658) );
XOR U29432 ( .A(c5886), .B(b[5886]), .Z(n17659) );
XNOR U29433 ( .A(b[5886]), .B(n17660), .Z(c[5886]) );
XNOR U29434 ( .A(a[5886]), .B(c5886), .Z(n17660) );
XOR U29435 ( .A(c5887), .B(n17661), .Z(c5888) );
ANDN U29436 ( .B(n17662), .A(n17663), .Z(n17661) );
XOR U29437 ( .A(c5887), .B(b[5887]), .Z(n17662) );
XNOR U29438 ( .A(b[5887]), .B(n17663), .Z(c[5887]) );
XNOR U29439 ( .A(a[5887]), .B(c5887), .Z(n17663) );
XOR U29440 ( .A(c5888), .B(n17664), .Z(c5889) );
ANDN U29441 ( .B(n17665), .A(n17666), .Z(n17664) );
XOR U29442 ( .A(c5888), .B(b[5888]), .Z(n17665) );
XNOR U29443 ( .A(b[5888]), .B(n17666), .Z(c[5888]) );
XNOR U29444 ( .A(a[5888]), .B(c5888), .Z(n17666) );
XOR U29445 ( .A(c5889), .B(n17667), .Z(c5890) );
ANDN U29446 ( .B(n17668), .A(n17669), .Z(n17667) );
XOR U29447 ( .A(c5889), .B(b[5889]), .Z(n17668) );
XNOR U29448 ( .A(b[5889]), .B(n17669), .Z(c[5889]) );
XNOR U29449 ( .A(a[5889]), .B(c5889), .Z(n17669) );
XOR U29450 ( .A(c5890), .B(n17670), .Z(c5891) );
ANDN U29451 ( .B(n17671), .A(n17672), .Z(n17670) );
XOR U29452 ( .A(c5890), .B(b[5890]), .Z(n17671) );
XNOR U29453 ( .A(b[5890]), .B(n17672), .Z(c[5890]) );
XNOR U29454 ( .A(a[5890]), .B(c5890), .Z(n17672) );
XOR U29455 ( .A(c5891), .B(n17673), .Z(c5892) );
ANDN U29456 ( .B(n17674), .A(n17675), .Z(n17673) );
XOR U29457 ( .A(c5891), .B(b[5891]), .Z(n17674) );
XNOR U29458 ( .A(b[5891]), .B(n17675), .Z(c[5891]) );
XNOR U29459 ( .A(a[5891]), .B(c5891), .Z(n17675) );
XOR U29460 ( .A(c5892), .B(n17676), .Z(c5893) );
ANDN U29461 ( .B(n17677), .A(n17678), .Z(n17676) );
XOR U29462 ( .A(c5892), .B(b[5892]), .Z(n17677) );
XNOR U29463 ( .A(b[5892]), .B(n17678), .Z(c[5892]) );
XNOR U29464 ( .A(a[5892]), .B(c5892), .Z(n17678) );
XOR U29465 ( .A(c5893), .B(n17679), .Z(c5894) );
ANDN U29466 ( .B(n17680), .A(n17681), .Z(n17679) );
XOR U29467 ( .A(c5893), .B(b[5893]), .Z(n17680) );
XNOR U29468 ( .A(b[5893]), .B(n17681), .Z(c[5893]) );
XNOR U29469 ( .A(a[5893]), .B(c5893), .Z(n17681) );
XOR U29470 ( .A(c5894), .B(n17682), .Z(c5895) );
ANDN U29471 ( .B(n17683), .A(n17684), .Z(n17682) );
XOR U29472 ( .A(c5894), .B(b[5894]), .Z(n17683) );
XNOR U29473 ( .A(b[5894]), .B(n17684), .Z(c[5894]) );
XNOR U29474 ( .A(a[5894]), .B(c5894), .Z(n17684) );
XOR U29475 ( .A(c5895), .B(n17685), .Z(c5896) );
ANDN U29476 ( .B(n17686), .A(n17687), .Z(n17685) );
XOR U29477 ( .A(c5895), .B(b[5895]), .Z(n17686) );
XNOR U29478 ( .A(b[5895]), .B(n17687), .Z(c[5895]) );
XNOR U29479 ( .A(a[5895]), .B(c5895), .Z(n17687) );
XOR U29480 ( .A(c5896), .B(n17688), .Z(c5897) );
ANDN U29481 ( .B(n17689), .A(n17690), .Z(n17688) );
XOR U29482 ( .A(c5896), .B(b[5896]), .Z(n17689) );
XNOR U29483 ( .A(b[5896]), .B(n17690), .Z(c[5896]) );
XNOR U29484 ( .A(a[5896]), .B(c5896), .Z(n17690) );
XOR U29485 ( .A(c5897), .B(n17691), .Z(c5898) );
ANDN U29486 ( .B(n17692), .A(n17693), .Z(n17691) );
XOR U29487 ( .A(c5897), .B(b[5897]), .Z(n17692) );
XNOR U29488 ( .A(b[5897]), .B(n17693), .Z(c[5897]) );
XNOR U29489 ( .A(a[5897]), .B(c5897), .Z(n17693) );
XOR U29490 ( .A(c5898), .B(n17694), .Z(c5899) );
ANDN U29491 ( .B(n17695), .A(n17696), .Z(n17694) );
XOR U29492 ( .A(c5898), .B(b[5898]), .Z(n17695) );
XNOR U29493 ( .A(b[5898]), .B(n17696), .Z(c[5898]) );
XNOR U29494 ( .A(a[5898]), .B(c5898), .Z(n17696) );
XOR U29495 ( .A(c5899), .B(n17697), .Z(c5900) );
ANDN U29496 ( .B(n17698), .A(n17699), .Z(n17697) );
XOR U29497 ( .A(c5899), .B(b[5899]), .Z(n17698) );
XNOR U29498 ( .A(b[5899]), .B(n17699), .Z(c[5899]) );
XNOR U29499 ( .A(a[5899]), .B(c5899), .Z(n17699) );
XOR U29500 ( .A(c5900), .B(n17700), .Z(c5901) );
ANDN U29501 ( .B(n17701), .A(n17702), .Z(n17700) );
XOR U29502 ( .A(c5900), .B(b[5900]), .Z(n17701) );
XNOR U29503 ( .A(b[5900]), .B(n17702), .Z(c[5900]) );
XNOR U29504 ( .A(a[5900]), .B(c5900), .Z(n17702) );
XOR U29505 ( .A(c5901), .B(n17703), .Z(c5902) );
ANDN U29506 ( .B(n17704), .A(n17705), .Z(n17703) );
XOR U29507 ( .A(c5901), .B(b[5901]), .Z(n17704) );
XNOR U29508 ( .A(b[5901]), .B(n17705), .Z(c[5901]) );
XNOR U29509 ( .A(a[5901]), .B(c5901), .Z(n17705) );
XOR U29510 ( .A(c5902), .B(n17706), .Z(c5903) );
ANDN U29511 ( .B(n17707), .A(n17708), .Z(n17706) );
XOR U29512 ( .A(c5902), .B(b[5902]), .Z(n17707) );
XNOR U29513 ( .A(b[5902]), .B(n17708), .Z(c[5902]) );
XNOR U29514 ( .A(a[5902]), .B(c5902), .Z(n17708) );
XOR U29515 ( .A(c5903), .B(n17709), .Z(c5904) );
ANDN U29516 ( .B(n17710), .A(n17711), .Z(n17709) );
XOR U29517 ( .A(c5903), .B(b[5903]), .Z(n17710) );
XNOR U29518 ( .A(b[5903]), .B(n17711), .Z(c[5903]) );
XNOR U29519 ( .A(a[5903]), .B(c5903), .Z(n17711) );
XOR U29520 ( .A(c5904), .B(n17712), .Z(c5905) );
ANDN U29521 ( .B(n17713), .A(n17714), .Z(n17712) );
XOR U29522 ( .A(c5904), .B(b[5904]), .Z(n17713) );
XNOR U29523 ( .A(b[5904]), .B(n17714), .Z(c[5904]) );
XNOR U29524 ( .A(a[5904]), .B(c5904), .Z(n17714) );
XOR U29525 ( .A(c5905), .B(n17715), .Z(c5906) );
ANDN U29526 ( .B(n17716), .A(n17717), .Z(n17715) );
XOR U29527 ( .A(c5905), .B(b[5905]), .Z(n17716) );
XNOR U29528 ( .A(b[5905]), .B(n17717), .Z(c[5905]) );
XNOR U29529 ( .A(a[5905]), .B(c5905), .Z(n17717) );
XOR U29530 ( .A(c5906), .B(n17718), .Z(c5907) );
ANDN U29531 ( .B(n17719), .A(n17720), .Z(n17718) );
XOR U29532 ( .A(c5906), .B(b[5906]), .Z(n17719) );
XNOR U29533 ( .A(b[5906]), .B(n17720), .Z(c[5906]) );
XNOR U29534 ( .A(a[5906]), .B(c5906), .Z(n17720) );
XOR U29535 ( .A(c5907), .B(n17721), .Z(c5908) );
ANDN U29536 ( .B(n17722), .A(n17723), .Z(n17721) );
XOR U29537 ( .A(c5907), .B(b[5907]), .Z(n17722) );
XNOR U29538 ( .A(b[5907]), .B(n17723), .Z(c[5907]) );
XNOR U29539 ( .A(a[5907]), .B(c5907), .Z(n17723) );
XOR U29540 ( .A(c5908), .B(n17724), .Z(c5909) );
ANDN U29541 ( .B(n17725), .A(n17726), .Z(n17724) );
XOR U29542 ( .A(c5908), .B(b[5908]), .Z(n17725) );
XNOR U29543 ( .A(b[5908]), .B(n17726), .Z(c[5908]) );
XNOR U29544 ( .A(a[5908]), .B(c5908), .Z(n17726) );
XOR U29545 ( .A(c5909), .B(n17727), .Z(c5910) );
ANDN U29546 ( .B(n17728), .A(n17729), .Z(n17727) );
XOR U29547 ( .A(c5909), .B(b[5909]), .Z(n17728) );
XNOR U29548 ( .A(b[5909]), .B(n17729), .Z(c[5909]) );
XNOR U29549 ( .A(a[5909]), .B(c5909), .Z(n17729) );
XOR U29550 ( .A(c5910), .B(n17730), .Z(c5911) );
ANDN U29551 ( .B(n17731), .A(n17732), .Z(n17730) );
XOR U29552 ( .A(c5910), .B(b[5910]), .Z(n17731) );
XNOR U29553 ( .A(b[5910]), .B(n17732), .Z(c[5910]) );
XNOR U29554 ( .A(a[5910]), .B(c5910), .Z(n17732) );
XOR U29555 ( .A(c5911), .B(n17733), .Z(c5912) );
ANDN U29556 ( .B(n17734), .A(n17735), .Z(n17733) );
XOR U29557 ( .A(c5911), .B(b[5911]), .Z(n17734) );
XNOR U29558 ( .A(b[5911]), .B(n17735), .Z(c[5911]) );
XNOR U29559 ( .A(a[5911]), .B(c5911), .Z(n17735) );
XOR U29560 ( .A(c5912), .B(n17736), .Z(c5913) );
ANDN U29561 ( .B(n17737), .A(n17738), .Z(n17736) );
XOR U29562 ( .A(c5912), .B(b[5912]), .Z(n17737) );
XNOR U29563 ( .A(b[5912]), .B(n17738), .Z(c[5912]) );
XNOR U29564 ( .A(a[5912]), .B(c5912), .Z(n17738) );
XOR U29565 ( .A(c5913), .B(n17739), .Z(c5914) );
ANDN U29566 ( .B(n17740), .A(n17741), .Z(n17739) );
XOR U29567 ( .A(c5913), .B(b[5913]), .Z(n17740) );
XNOR U29568 ( .A(b[5913]), .B(n17741), .Z(c[5913]) );
XNOR U29569 ( .A(a[5913]), .B(c5913), .Z(n17741) );
XOR U29570 ( .A(c5914), .B(n17742), .Z(c5915) );
ANDN U29571 ( .B(n17743), .A(n17744), .Z(n17742) );
XOR U29572 ( .A(c5914), .B(b[5914]), .Z(n17743) );
XNOR U29573 ( .A(b[5914]), .B(n17744), .Z(c[5914]) );
XNOR U29574 ( .A(a[5914]), .B(c5914), .Z(n17744) );
XOR U29575 ( .A(c5915), .B(n17745), .Z(c5916) );
ANDN U29576 ( .B(n17746), .A(n17747), .Z(n17745) );
XOR U29577 ( .A(c5915), .B(b[5915]), .Z(n17746) );
XNOR U29578 ( .A(b[5915]), .B(n17747), .Z(c[5915]) );
XNOR U29579 ( .A(a[5915]), .B(c5915), .Z(n17747) );
XOR U29580 ( .A(c5916), .B(n17748), .Z(c5917) );
ANDN U29581 ( .B(n17749), .A(n17750), .Z(n17748) );
XOR U29582 ( .A(c5916), .B(b[5916]), .Z(n17749) );
XNOR U29583 ( .A(b[5916]), .B(n17750), .Z(c[5916]) );
XNOR U29584 ( .A(a[5916]), .B(c5916), .Z(n17750) );
XOR U29585 ( .A(c5917), .B(n17751), .Z(c5918) );
ANDN U29586 ( .B(n17752), .A(n17753), .Z(n17751) );
XOR U29587 ( .A(c5917), .B(b[5917]), .Z(n17752) );
XNOR U29588 ( .A(b[5917]), .B(n17753), .Z(c[5917]) );
XNOR U29589 ( .A(a[5917]), .B(c5917), .Z(n17753) );
XOR U29590 ( .A(c5918), .B(n17754), .Z(c5919) );
ANDN U29591 ( .B(n17755), .A(n17756), .Z(n17754) );
XOR U29592 ( .A(c5918), .B(b[5918]), .Z(n17755) );
XNOR U29593 ( .A(b[5918]), .B(n17756), .Z(c[5918]) );
XNOR U29594 ( .A(a[5918]), .B(c5918), .Z(n17756) );
XOR U29595 ( .A(c5919), .B(n17757), .Z(c5920) );
ANDN U29596 ( .B(n17758), .A(n17759), .Z(n17757) );
XOR U29597 ( .A(c5919), .B(b[5919]), .Z(n17758) );
XNOR U29598 ( .A(b[5919]), .B(n17759), .Z(c[5919]) );
XNOR U29599 ( .A(a[5919]), .B(c5919), .Z(n17759) );
XOR U29600 ( .A(c5920), .B(n17760), .Z(c5921) );
ANDN U29601 ( .B(n17761), .A(n17762), .Z(n17760) );
XOR U29602 ( .A(c5920), .B(b[5920]), .Z(n17761) );
XNOR U29603 ( .A(b[5920]), .B(n17762), .Z(c[5920]) );
XNOR U29604 ( .A(a[5920]), .B(c5920), .Z(n17762) );
XOR U29605 ( .A(c5921), .B(n17763), .Z(c5922) );
ANDN U29606 ( .B(n17764), .A(n17765), .Z(n17763) );
XOR U29607 ( .A(c5921), .B(b[5921]), .Z(n17764) );
XNOR U29608 ( .A(b[5921]), .B(n17765), .Z(c[5921]) );
XNOR U29609 ( .A(a[5921]), .B(c5921), .Z(n17765) );
XOR U29610 ( .A(c5922), .B(n17766), .Z(c5923) );
ANDN U29611 ( .B(n17767), .A(n17768), .Z(n17766) );
XOR U29612 ( .A(c5922), .B(b[5922]), .Z(n17767) );
XNOR U29613 ( .A(b[5922]), .B(n17768), .Z(c[5922]) );
XNOR U29614 ( .A(a[5922]), .B(c5922), .Z(n17768) );
XOR U29615 ( .A(c5923), .B(n17769), .Z(c5924) );
ANDN U29616 ( .B(n17770), .A(n17771), .Z(n17769) );
XOR U29617 ( .A(c5923), .B(b[5923]), .Z(n17770) );
XNOR U29618 ( .A(b[5923]), .B(n17771), .Z(c[5923]) );
XNOR U29619 ( .A(a[5923]), .B(c5923), .Z(n17771) );
XOR U29620 ( .A(c5924), .B(n17772), .Z(c5925) );
ANDN U29621 ( .B(n17773), .A(n17774), .Z(n17772) );
XOR U29622 ( .A(c5924), .B(b[5924]), .Z(n17773) );
XNOR U29623 ( .A(b[5924]), .B(n17774), .Z(c[5924]) );
XNOR U29624 ( .A(a[5924]), .B(c5924), .Z(n17774) );
XOR U29625 ( .A(c5925), .B(n17775), .Z(c5926) );
ANDN U29626 ( .B(n17776), .A(n17777), .Z(n17775) );
XOR U29627 ( .A(c5925), .B(b[5925]), .Z(n17776) );
XNOR U29628 ( .A(b[5925]), .B(n17777), .Z(c[5925]) );
XNOR U29629 ( .A(a[5925]), .B(c5925), .Z(n17777) );
XOR U29630 ( .A(c5926), .B(n17778), .Z(c5927) );
ANDN U29631 ( .B(n17779), .A(n17780), .Z(n17778) );
XOR U29632 ( .A(c5926), .B(b[5926]), .Z(n17779) );
XNOR U29633 ( .A(b[5926]), .B(n17780), .Z(c[5926]) );
XNOR U29634 ( .A(a[5926]), .B(c5926), .Z(n17780) );
XOR U29635 ( .A(c5927), .B(n17781), .Z(c5928) );
ANDN U29636 ( .B(n17782), .A(n17783), .Z(n17781) );
XOR U29637 ( .A(c5927), .B(b[5927]), .Z(n17782) );
XNOR U29638 ( .A(b[5927]), .B(n17783), .Z(c[5927]) );
XNOR U29639 ( .A(a[5927]), .B(c5927), .Z(n17783) );
XOR U29640 ( .A(c5928), .B(n17784), .Z(c5929) );
ANDN U29641 ( .B(n17785), .A(n17786), .Z(n17784) );
XOR U29642 ( .A(c5928), .B(b[5928]), .Z(n17785) );
XNOR U29643 ( .A(b[5928]), .B(n17786), .Z(c[5928]) );
XNOR U29644 ( .A(a[5928]), .B(c5928), .Z(n17786) );
XOR U29645 ( .A(c5929), .B(n17787), .Z(c5930) );
ANDN U29646 ( .B(n17788), .A(n17789), .Z(n17787) );
XOR U29647 ( .A(c5929), .B(b[5929]), .Z(n17788) );
XNOR U29648 ( .A(b[5929]), .B(n17789), .Z(c[5929]) );
XNOR U29649 ( .A(a[5929]), .B(c5929), .Z(n17789) );
XOR U29650 ( .A(c5930), .B(n17790), .Z(c5931) );
ANDN U29651 ( .B(n17791), .A(n17792), .Z(n17790) );
XOR U29652 ( .A(c5930), .B(b[5930]), .Z(n17791) );
XNOR U29653 ( .A(b[5930]), .B(n17792), .Z(c[5930]) );
XNOR U29654 ( .A(a[5930]), .B(c5930), .Z(n17792) );
XOR U29655 ( .A(c5931), .B(n17793), .Z(c5932) );
ANDN U29656 ( .B(n17794), .A(n17795), .Z(n17793) );
XOR U29657 ( .A(c5931), .B(b[5931]), .Z(n17794) );
XNOR U29658 ( .A(b[5931]), .B(n17795), .Z(c[5931]) );
XNOR U29659 ( .A(a[5931]), .B(c5931), .Z(n17795) );
XOR U29660 ( .A(c5932), .B(n17796), .Z(c5933) );
ANDN U29661 ( .B(n17797), .A(n17798), .Z(n17796) );
XOR U29662 ( .A(c5932), .B(b[5932]), .Z(n17797) );
XNOR U29663 ( .A(b[5932]), .B(n17798), .Z(c[5932]) );
XNOR U29664 ( .A(a[5932]), .B(c5932), .Z(n17798) );
XOR U29665 ( .A(c5933), .B(n17799), .Z(c5934) );
ANDN U29666 ( .B(n17800), .A(n17801), .Z(n17799) );
XOR U29667 ( .A(c5933), .B(b[5933]), .Z(n17800) );
XNOR U29668 ( .A(b[5933]), .B(n17801), .Z(c[5933]) );
XNOR U29669 ( .A(a[5933]), .B(c5933), .Z(n17801) );
XOR U29670 ( .A(c5934), .B(n17802), .Z(c5935) );
ANDN U29671 ( .B(n17803), .A(n17804), .Z(n17802) );
XOR U29672 ( .A(c5934), .B(b[5934]), .Z(n17803) );
XNOR U29673 ( .A(b[5934]), .B(n17804), .Z(c[5934]) );
XNOR U29674 ( .A(a[5934]), .B(c5934), .Z(n17804) );
XOR U29675 ( .A(c5935), .B(n17805), .Z(c5936) );
ANDN U29676 ( .B(n17806), .A(n17807), .Z(n17805) );
XOR U29677 ( .A(c5935), .B(b[5935]), .Z(n17806) );
XNOR U29678 ( .A(b[5935]), .B(n17807), .Z(c[5935]) );
XNOR U29679 ( .A(a[5935]), .B(c5935), .Z(n17807) );
XOR U29680 ( .A(c5936), .B(n17808), .Z(c5937) );
ANDN U29681 ( .B(n17809), .A(n17810), .Z(n17808) );
XOR U29682 ( .A(c5936), .B(b[5936]), .Z(n17809) );
XNOR U29683 ( .A(b[5936]), .B(n17810), .Z(c[5936]) );
XNOR U29684 ( .A(a[5936]), .B(c5936), .Z(n17810) );
XOR U29685 ( .A(c5937), .B(n17811), .Z(c5938) );
ANDN U29686 ( .B(n17812), .A(n17813), .Z(n17811) );
XOR U29687 ( .A(c5937), .B(b[5937]), .Z(n17812) );
XNOR U29688 ( .A(b[5937]), .B(n17813), .Z(c[5937]) );
XNOR U29689 ( .A(a[5937]), .B(c5937), .Z(n17813) );
XOR U29690 ( .A(c5938), .B(n17814), .Z(c5939) );
ANDN U29691 ( .B(n17815), .A(n17816), .Z(n17814) );
XOR U29692 ( .A(c5938), .B(b[5938]), .Z(n17815) );
XNOR U29693 ( .A(b[5938]), .B(n17816), .Z(c[5938]) );
XNOR U29694 ( .A(a[5938]), .B(c5938), .Z(n17816) );
XOR U29695 ( .A(c5939), .B(n17817), .Z(c5940) );
ANDN U29696 ( .B(n17818), .A(n17819), .Z(n17817) );
XOR U29697 ( .A(c5939), .B(b[5939]), .Z(n17818) );
XNOR U29698 ( .A(b[5939]), .B(n17819), .Z(c[5939]) );
XNOR U29699 ( .A(a[5939]), .B(c5939), .Z(n17819) );
XOR U29700 ( .A(c5940), .B(n17820), .Z(c5941) );
ANDN U29701 ( .B(n17821), .A(n17822), .Z(n17820) );
XOR U29702 ( .A(c5940), .B(b[5940]), .Z(n17821) );
XNOR U29703 ( .A(b[5940]), .B(n17822), .Z(c[5940]) );
XNOR U29704 ( .A(a[5940]), .B(c5940), .Z(n17822) );
XOR U29705 ( .A(c5941), .B(n17823), .Z(c5942) );
ANDN U29706 ( .B(n17824), .A(n17825), .Z(n17823) );
XOR U29707 ( .A(c5941), .B(b[5941]), .Z(n17824) );
XNOR U29708 ( .A(b[5941]), .B(n17825), .Z(c[5941]) );
XNOR U29709 ( .A(a[5941]), .B(c5941), .Z(n17825) );
XOR U29710 ( .A(c5942), .B(n17826), .Z(c5943) );
ANDN U29711 ( .B(n17827), .A(n17828), .Z(n17826) );
XOR U29712 ( .A(c5942), .B(b[5942]), .Z(n17827) );
XNOR U29713 ( .A(b[5942]), .B(n17828), .Z(c[5942]) );
XNOR U29714 ( .A(a[5942]), .B(c5942), .Z(n17828) );
XOR U29715 ( .A(c5943), .B(n17829), .Z(c5944) );
ANDN U29716 ( .B(n17830), .A(n17831), .Z(n17829) );
XOR U29717 ( .A(c5943), .B(b[5943]), .Z(n17830) );
XNOR U29718 ( .A(b[5943]), .B(n17831), .Z(c[5943]) );
XNOR U29719 ( .A(a[5943]), .B(c5943), .Z(n17831) );
XOR U29720 ( .A(c5944), .B(n17832), .Z(c5945) );
ANDN U29721 ( .B(n17833), .A(n17834), .Z(n17832) );
XOR U29722 ( .A(c5944), .B(b[5944]), .Z(n17833) );
XNOR U29723 ( .A(b[5944]), .B(n17834), .Z(c[5944]) );
XNOR U29724 ( .A(a[5944]), .B(c5944), .Z(n17834) );
XOR U29725 ( .A(c5945), .B(n17835), .Z(c5946) );
ANDN U29726 ( .B(n17836), .A(n17837), .Z(n17835) );
XOR U29727 ( .A(c5945), .B(b[5945]), .Z(n17836) );
XNOR U29728 ( .A(b[5945]), .B(n17837), .Z(c[5945]) );
XNOR U29729 ( .A(a[5945]), .B(c5945), .Z(n17837) );
XOR U29730 ( .A(c5946), .B(n17838), .Z(c5947) );
ANDN U29731 ( .B(n17839), .A(n17840), .Z(n17838) );
XOR U29732 ( .A(c5946), .B(b[5946]), .Z(n17839) );
XNOR U29733 ( .A(b[5946]), .B(n17840), .Z(c[5946]) );
XNOR U29734 ( .A(a[5946]), .B(c5946), .Z(n17840) );
XOR U29735 ( .A(c5947), .B(n17841), .Z(c5948) );
ANDN U29736 ( .B(n17842), .A(n17843), .Z(n17841) );
XOR U29737 ( .A(c5947), .B(b[5947]), .Z(n17842) );
XNOR U29738 ( .A(b[5947]), .B(n17843), .Z(c[5947]) );
XNOR U29739 ( .A(a[5947]), .B(c5947), .Z(n17843) );
XOR U29740 ( .A(c5948), .B(n17844), .Z(c5949) );
ANDN U29741 ( .B(n17845), .A(n17846), .Z(n17844) );
XOR U29742 ( .A(c5948), .B(b[5948]), .Z(n17845) );
XNOR U29743 ( .A(b[5948]), .B(n17846), .Z(c[5948]) );
XNOR U29744 ( .A(a[5948]), .B(c5948), .Z(n17846) );
XOR U29745 ( .A(c5949), .B(n17847), .Z(c5950) );
ANDN U29746 ( .B(n17848), .A(n17849), .Z(n17847) );
XOR U29747 ( .A(c5949), .B(b[5949]), .Z(n17848) );
XNOR U29748 ( .A(b[5949]), .B(n17849), .Z(c[5949]) );
XNOR U29749 ( .A(a[5949]), .B(c5949), .Z(n17849) );
XOR U29750 ( .A(c5950), .B(n17850), .Z(c5951) );
ANDN U29751 ( .B(n17851), .A(n17852), .Z(n17850) );
XOR U29752 ( .A(c5950), .B(b[5950]), .Z(n17851) );
XNOR U29753 ( .A(b[5950]), .B(n17852), .Z(c[5950]) );
XNOR U29754 ( .A(a[5950]), .B(c5950), .Z(n17852) );
XOR U29755 ( .A(c5951), .B(n17853), .Z(c5952) );
ANDN U29756 ( .B(n17854), .A(n17855), .Z(n17853) );
XOR U29757 ( .A(c5951), .B(b[5951]), .Z(n17854) );
XNOR U29758 ( .A(b[5951]), .B(n17855), .Z(c[5951]) );
XNOR U29759 ( .A(a[5951]), .B(c5951), .Z(n17855) );
XOR U29760 ( .A(c5952), .B(n17856), .Z(c5953) );
ANDN U29761 ( .B(n17857), .A(n17858), .Z(n17856) );
XOR U29762 ( .A(c5952), .B(b[5952]), .Z(n17857) );
XNOR U29763 ( .A(b[5952]), .B(n17858), .Z(c[5952]) );
XNOR U29764 ( .A(a[5952]), .B(c5952), .Z(n17858) );
XOR U29765 ( .A(c5953), .B(n17859), .Z(c5954) );
ANDN U29766 ( .B(n17860), .A(n17861), .Z(n17859) );
XOR U29767 ( .A(c5953), .B(b[5953]), .Z(n17860) );
XNOR U29768 ( .A(b[5953]), .B(n17861), .Z(c[5953]) );
XNOR U29769 ( .A(a[5953]), .B(c5953), .Z(n17861) );
XOR U29770 ( .A(c5954), .B(n17862), .Z(c5955) );
ANDN U29771 ( .B(n17863), .A(n17864), .Z(n17862) );
XOR U29772 ( .A(c5954), .B(b[5954]), .Z(n17863) );
XNOR U29773 ( .A(b[5954]), .B(n17864), .Z(c[5954]) );
XNOR U29774 ( .A(a[5954]), .B(c5954), .Z(n17864) );
XOR U29775 ( .A(c5955), .B(n17865), .Z(c5956) );
ANDN U29776 ( .B(n17866), .A(n17867), .Z(n17865) );
XOR U29777 ( .A(c5955), .B(b[5955]), .Z(n17866) );
XNOR U29778 ( .A(b[5955]), .B(n17867), .Z(c[5955]) );
XNOR U29779 ( .A(a[5955]), .B(c5955), .Z(n17867) );
XOR U29780 ( .A(c5956), .B(n17868), .Z(c5957) );
ANDN U29781 ( .B(n17869), .A(n17870), .Z(n17868) );
XOR U29782 ( .A(c5956), .B(b[5956]), .Z(n17869) );
XNOR U29783 ( .A(b[5956]), .B(n17870), .Z(c[5956]) );
XNOR U29784 ( .A(a[5956]), .B(c5956), .Z(n17870) );
XOR U29785 ( .A(c5957), .B(n17871), .Z(c5958) );
ANDN U29786 ( .B(n17872), .A(n17873), .Z(n17871) );
XOR U29787 ( .A(c5957), .B(b[5957]), .Z(n17872) );
XNOR U29788 ( .A(b[5957]), .B(n17873), .Z(c[5957]) );
XNOR U29789 ( .A(a[5957]), .B(c5957), .Z(n17873) );
XOR U29790 ( .A(c5958), .B(n17874), .Z(c5959) );
ANDN U29791 ( .B(n17875), .A(n17876), .Z(n17874) );
XOR U29792 ( .A(c5958), .B(b[5958]), .Z(n17875) );
XNOR U29793 ( .A(b[5958]), .B(n17876), .Z(c[5958]) );
XNOR U29794 ( .A(a[5958]), .B(c5958), .Z(n17876) );
XOR U29795 ( .A(c5959), .B(n17877), .Z(c5960) );
ANDN U29796 ( .B(n17878), .A(n17879), .Z(n17877) );
XOR U29797 ( .A(c5959), .B(b[5959]), .Z(n17878) );
XNOR U29798 ( .A(b[5959]), .B(n17879), .Z(c[5959]) );
XNOR U29799 ( .A(a[5959]), .B(c5959), .Z(n17879) );
XOR U29800 ( .A(c5960), .B(n17880), .Z(c5961) );
ANDN U29801 ( .B(n17881), .A(n17882), .Z(n17880) );
XOR U29802 ( .A(c5960), .B(b[5960]), .Z(n17881) );
XNOR U29803 ( .A(b[5960]), .B(n17882), .Z(c[5960]) );
XNOR U29804 ( .A(a[5960]), .B(c5960), .Z(n17882) );
XOR U29805 ( .A(c5961), .B(n17883), .Z(c5962) );
ANDN U29806 ( .B(n17884), .A(n17885), .Z(n17883) );
XOR U29807 ( .A(c5961), .B(b[5961]), .Z(n17884) );
XNOR U29808 ( .A(b[5961]), .B(n17885), .Z(c[5961]) );
XNOR U29809 ( .A(a[5961]), .B(c5961), .Z(n17885) );
XOR U29810 ( .A(c5962), .B(n17886), .Z(c5963) );
ANDN U29811 ( .B(n17887), .A(n17888), .Z(n17886) );
XOR U29812 ( .A(c5962), .B(b[5962]), .Z(n17887) );
XNOR U29813 ( .A(b[5962]), .B(n17888), .Z(c[5962]) );
XNOR U29814 ( .A(a[5962]), .B(c5962), .Z(n17888) );
XOR U29815 ( .A(c5963), .B(n17889), .Z(c5964) );
ANDN U29816 ( .B(n17890), .A(n17891), .Z(n17889) );
XOR U29817 ( .A(c5963), .B(b[5963]), .Z(n17890) );
XNOR U29818 ( .A(b[5963]), .B(n17891), .Z(c[5963]) );
XNOR U29819 ( .A(a[5963]), .B(c5963), .Z(n17891) );
XOR U29820 ( .A(c5964), .B(n17892), .Z(c5965) );
ANDN U29821 ( .B(n17893), .A(n17894), .Z(n17892) );
XOR U29822 ( .A(c5964), .B(b[5964]), .Z(n17893) );
XNOR U29823 ( .A(b[5964]), .B(n17894), .Z(c[5964]) );
XNOR U29824 ( .A(a[5964]), .B(c5964), .Z(n17894) );
XOR U29825 ( .A(c5965), .B(n17895), .Z(c5966) );
ANDN U29826 ( .B(n17896), .A(n17897), .Z(n17895) );
XOR U29827 ( .A(c5965), .B(b[5965]), .Z(n17896) );
XNOR U29828 ( .A(b[5965]), .B(n17897), .Z(c[5965]) );
XNOR U29829 ( .A(a[5965]), .B(c5965), .Z(n17897) );
XOR U29830 ( .A(c5966), .B(n17898), .Z(c5967) );
ANDN U29831 ( .B(n17899), .A(n17900), .Z(n17898) );
XOR U29832 ( .A(c5966), .B(b[5966]), .Z(n17899) );
XNOR U29833 ( .A(b[5966]), .B(n17900), .Z(c[5966]) );
XNOR U29834 ( .A(a[5966]), .B(c5966), .Z(n17900) );
XOR U29835 ( .A(c5967), .B(n17901), .Z(c5968) );
ANDN U29836 ( .B(n17902), .A(n17903), .Z(n17901) );
XOR U29837 ( .A(c5967), .B(b[5967]), .Z(n17902) );
XNOR U29838 ( .A(b[5967]), .B(n17903), .Z(c[5967]) );
XNOR U29839 ( .A(a[5967]), .B(c5967), .Z(n17903) );
XOR U29840 ( .A(c5968), .B(n17904), .Z(c5969) );
ANDN U29841 ( .B(n17905), .A(n17906), .Z(n17904) );
XOR U29842 ( .A(c5968), .B(b[5968]), .Z(n17905) );
XNOR U29843 ( .A(b[5968]), .B(n17906), .Z(c[5968]) );
XNOR U29844 ( .A(a[5968]), .B(c5968), .Z(n17906) );
XOR U29845 ( .A(c5969), .B(n17907), .Z(c5970) );
ANDN U29846 ( .B(n17908), .A(n17909), .Z(n17907) );
XOR U29847 ( .A(c5969), .B(b[5969]), .Z(n17908) );
XNOR U29848 ( .A(b[5969]), .B(n17909), .Z(c[5969]) );
XNOR U29849 ( .A(a[5969]), .B(c5969), .Z(n17909) );
XOR U29850 ( .A(c5970), .B(n17910), .Z(c5971) );
ANDN U29851 ( .B(n17911), .A(n17912), .Z(n17910) );
XOR U29852 ( .A(c5970), .B(b[5970]), .Z(n17911) );
XNOR U29853 ( .A(b[5970]), .B(n17912), .Z(c[5970]) );
XNOR U29854 ( .A(a[5970]), .B(c5970), .Z(n17912) );
XOR U29855 ( .A(c5971), .B(n17913), .Z(c5972) );
ANDN U29856 ( .B(n17914), .A(n17915), .Z(n17913) );
XOR U29857 ( .A(c5971), .B(b[5971]), .Z(n17914) );
XNOR U29858 ( .A(b[5971]), .B(n17915), .Z(c[5971]) );
XNOR U29859 ( .A(a[5971]), .B(c5971), .Z(n17915) );
XOR U29860 ( .A(c5972), .B(n17916), .Z(c5973) );
ANDN U29861 ( .B(n17917), .A(n17918), .Z(n17916) );
XOR U29862 ( .A(c5972), .B(b[5972]), .Z(n17917) );
XNOR U29863 ( .A(b[5972]), .B(n17918), .Z(c[5972]) );
XNOR U29864 ( .A(a[5972]), .B(c5972), .Z(n17918) );
XOR U29865 ( .A(c5973), .B(n17919), .Z(c5974) );
ANDN U29866 ( .B(n17920), .A(n17921), .Z(n17919) );
XOR U29867 ( .A(c5973), .B(b[5973]), .Z(n17920) );
XNOR U29868 ( .A(b[5973]), .B(n17921), .Z(c[5973]) );
XNOR U29869 ( .A(a[5973]), .B(c5973), .Z(n17921) );
XOR U29870 ( .A(c5974), .B(n17922), .Z(c5975) );
ANDN U29871 ( .B(n17923), .A(n17924), .Z(n17922) );
XOR U29872 ( .A(c5974), .B(b[5974]), .Z(n17923) );
XNOR U29873 ( .A(b[5974]), .B(n17924), .Z(c[5974]) );
XNOR U29874 ( .A(a[5974]), .B(c5974), .Z(n17924) );
XOR U29875 ( .A(c5975), .B(n17925), .Z(c5976) );
ANDN U29876 ( .B(n17926), .A(n17927), .Z(n17925) );
XOR U29877 ( .A(c5975), .B(b[5975]), .Z(n17926) );
XNOR U29878 ( .A(b[5975]), .B(n17927), .Z(c[5975]) );
XNOR U29879 ( .A(a[5975]), .B(c5975), .Z(n17927) );
XOR U29880 ( .A(c5976), .B(n17928), .Z(c5977) );
ANDN U29881 ( .B(n17929), .A(n17930), .Z(n17928) );
XOR U29882 ( .A(c5976), .B(b[5976]), .Z(n17929) );
XNOR U29883 ( .A(b[5976]), .B(n17930), .Z(c[5976]) );
XNOR U29884 ( .A(a[5976]), .B(c5976), .Z(n17930) );
XOR U29885 ( .A(c5977), .B(n17931), .Z(c5978) );
ANDN U29886 ( .B(n17932), .A(n17933), .Z(n17931) );
XOR U29887 ( .A(c5977), .B(b[5977]), .Z(n17932) );
XNOR U29888 ( .A(b[5977]), .B(n17933), .Z(c[5977]) );
XNOR U29889 ( .A(a[5977]), .B(c5977), .Z(n17933) );
XOR U29890 ( .A(c5978), .B(n17934), .Z(c5979) );
ANDN U29891 ( .B(n17935), .A(n17936), .Z(n17934) );
XOR U29892 ( .A(c5978), .B(b[5978]), .Z(n17935) );
XNOR U29893 ( .A(b[5978]), .B(n17936), .Z(c[5978]) );
XNOR U29894 ( .A(a[5978]), .B(c5978), .Z(n17936) );
XOR U29895 ( .A(c5979), .B(n17937), .Z(c5980) );
ANDN U29896 ( .B(n17938), .A(n17939), .Z(n17937) );
XOR U29897 ( .A(c5979), .B(b[5979]), .Z(n17938) );
XNOR U29898 ( .A(b[5979]), .B(n17939), .Z(c[5979]) );
XNOR U29899 ( .A(a[5979]), .B(c5979), .Z(n17939) );
XOR U29900 ( .A(c5980), .B(n17940), .Z(c5981) );
ANDN U29901 ( .B(n17941), .A(n17942), .Z(n17940) );
XOR U29902 ( .A(c5980), .B(b[5980]), .Z(n17941) );
XNOR U29903 ( .A(b[5980]), .B(n17942), .Z(c[5980]) );
XNOR U29904 ( .A(a[5980]), .B(c5980), .Z(n17942) );
XOR U29905 ( .A(c5981), .B(n17943), .Z(c5982) );
ANDN U29906 ( .B(n17944), .A(n17945), .Z(n17943) );
XOR U29907 ( .A(c5981), .B(b[5981]), .Z(n17944) );
XNOR U29908 ( .A(b[5981]), .B(n17945), .Z(c[5981]) );
XNOR U29909 ( .A(a[5981]), .B(c5981), .Z(n17945) );
XOR U29910 ( .A(c5982), .B(n17946), .Z(c5983) );
ANDN U29911 ( .B(n17947), .A(n17948), .Z(n17946) );
XOR U29912 ( .A(c5982), .B(b[5982]), .Z(n17947) );
XNOR U29913 ( .A(b[5982]), .B(n17948), .Z(c[5982]) );
XNOR U29914 ( .A(a[5982]), .B(c5982), .Z(n17948) );
XOR U29915 ( .A(c5983), .B(n17949), .Z(c5984) );
ANDN U29916 ( .B(n17950), .A(n17951), .Z(n17949) );
XOR U29917 ( .A(c5983), .B(b[5983]), .Z(n17950) );
XNOR U29918 ( .A(b[5983]), .B(n17951), .Z(c[5983]) );
XNOR U29919 ( .A(a[5983]), .B(c5983), .Z(n17951) );
XOR U29920 ( .A(c5984), .B(n17952), .Z(c5985) );
ANDN U29921 ( .B(n17953), .A(n17954), .Z(n17952) );
XOR U29922 ( .A(c5984), .B(b[5984]), .Z(n17953) );
XNOR U29923 ( .A(b[5984]), .B(n17954), .Z(c[5984]) );
XNOR U29924 ( .A(a[5984]), .B(c5984), .Z(n17954) );
XOR U29925 ( .A(c5985), .B(n17955), .Z(c5986) );
ANDN U29926 ( .B(n17956), .A(n17957), .Z(n17955) );
XOR U29927 ( .A(c5985), .B(b[5985]), .Z(n17956) );
XNOR U29928 ( .A(b[5985]), .B(n17957), .Z(c[5985]) );
XNOR U29929 ( .A(a[5985]), .B(c5985), .Z(n17957) );
XOR U29930 ( .A(c5986), .B(n17958), .Z(c5987) );
ANDN U29931 ( .B(n17959), .A(n17960), .Z(n17958) );
XOR U29932 ( .A(c5986), .B(b[5986]), .Z(n17959) );
XNOR U29933 ( .A(b[5986]), .B(n17960), .Z(c[5986]) );
XNOR U29934 ( .A(a[5986]), .B(c5986), .Z(n17960) );
XOR U29935 ( .A(c5987), .B(n17961), .Z(c5988) );
ANDN U29936 ( .B(n17962), .A(n17963), .Z(n17961) );
XOR U29937 ( .A(c5987), .B(b[5987]), .Z(n17962) );
XNOR U29938 ( .A(b[5987]), .B(n17963), .Z(c[5987]) );
XNOR U29939 ( .A(a[5987]), .B(c5987), .Z(n17963) );
XOR U29940 ( .A(c5988), .B(n17964), .Z(c5989) );
ANDN U29941 ( .B(n17965), .A(n17966), .Z(n17964) );
XOR U29942 ( .A(c5988), .B(b[5988]), .Z(n17965) );
XNOR U29943 ( .A(b[5988]), .B(n17966), .Z(c[5988]) );
XNOR U29944 ( .A(a[5988]), .B(c5988), .Z(n17966) );
XOR U29945 ( .A(c5989), .B(n17967), .Z(c5990) );
ANDN U29946 ( .B(n17968), .A(n17969), .Z(n17967) );
XOR U29947 ( .A(c5989), .B(b[5989]), .Z(n17968) );
XNOR U29948 ( .A(b[5989]), .B(n17969), .Z(c[5989]) );
XNOR U29949 ( .A(a[5989]), .B(c5989), .Z(n17969) );
XOR U29950 ( .A(c5990), .B(n17970), .Z(c5991) );
ANDN U29951 ( .B(n17971), .A(n17972), .Z(n17970) );
XOR U29952 ( .A(c5990), .B(b[5990]), .Z(n17971) );
XNOR U29953 ( .A(b[5990]), .B(n17972), .Z(c[5990]) );
XNOR U29954 ( .A(a[5990]), .B(c5990), .Z(n17972) );
XOR U29955 ( .A(c5991), .B(n17973), .Z(c5992) );
ANDN U29956 ( .B(n17974), .A(n17975), .Z(n17973) );
XOR U29957 ( .A(c5991), .B(b[5991]), .Z(n17974) );
XNOR U29958 ( .A(b[5991]), .B(n17975), .Z(c[5991]) );
XNOR U29959 ( .A(a[5991]), .B(c5991), .Z(n17975) );
XOR U29960 ( .A(c5992), .B(n17976), .Z(c5993) );
ANDN U29961 ( .B(n17977), .A(n17978), .Z(n17976) );
XOR U29962 ( .A(c5992), .B(b[5992]), .Z(n17977) );
XNOR U29963 ( .A(b[5992]), .B(n17978), .Z(c[5992]) );
XNOR U29964 ( .A(a[5992]), .B(c5992), .Z(n17978) );
XOR U29965 ( .A(c5993), .B(n17979), .Z(c5994) );
ANDN U29966 ( .B(n17980), .A(n17981), .Z(n17979) );
XOR U29967 ( .A(c5993), .B(b[5993]), .Z(n17980) );
XNOR U29968 ( .A(b[5993]), .B(n17981), .Z(c[5993]) );
XNOR U29969 ( .A(a[5993]), .B(c5993), .Z(n17981) );
XOR U29970 ( .A(c5994), .B(n17982), .Z(c5995) );
ANDN U29971 ( .B(n17983), .A(n17984), .Z(n17982) );
XOR U29972 ( .A(c5994), .B(b[5994]), .Z(n17983) );
XNOR U29973 ( .A(b[5994]), .B(n17984), .Z(c[5994]) );
XNOR U29974 ( .A(a[5994]), .B(c5994), .Z(n17984) );
XOR U29975 ( .A(c5995), .B(n17985), .Z(c5996) );
ANDN U29976 ( .B(n17986), .A(n17987), .Z(n17985) );
XOR U29977 ( .A(c5995), .B(b[5995]), .Z(n17986) );
XNOR U29978 ( .A(b[5995]), .B(n17987), .Z(c[5995]) );
XNOR U29979 ( .A(a[5995]), .B(c5995), .Z(n17987) );
XOR U29980 ( .A(c5996), .B(n17988), .Z(c5997) );
ANDN U29981 ( .B(n17989), .A(n17990), .Z(n17988) );
XOR U29982 ( .A(c5996), .B(b[5996]), .Z(n17989) );
XNOR U29983 ( .A(b[5996]), .B(n17990), .Z(c[5996]) );
XNOR U29984 ( .A(a[5996]), .B(c5996), .Z(n17990) );
XOR U29985 ( .A(c5997), .B(n17991), .Z(c5998) );
ANDN U29986 ( .B(n17992), .A(n17993), .Z(n17991) );
XOR U29987 ( .A(c5997), .B(b[5997]), .Z(n17992) );
XNOR U29988 ( .A(b[5997]), .B(n17993), .Z(c[5997]) );
XNOR U29989 ( .A(a[5997]), .B(c5997), .Z(n17993) );
XOR U29990 ( .A(c5998), .B(n17994), .Z(c5999) );
ANDN U29991 ( .B(n17995), .A(n17996), .Z(n17994) );
XOR U29992 ( .A(c5998), .B(b[5998]), .Z(n17995) );
XNOR U29993 ( .A(b[5998]), .B(n17996), .Z(c[5998]) );
XNOR U29994 ( .A(a[5998]), .B(c5998), .Z(n17996) );
XOR U29995 ( .A(c5999), .B(n17997), .Z(c6000) );
ANDN U29996 ( .B(n17998), .A(n17999), .Z(n17997) );
XOR U29997 ( .A(c5999), .B(b[5999]), .Z(n17998) );
XNOR U29998 ( .A(b[5999]), .B(n17999), .Z(c[5999]) );
XNOR U29999 ( .A(a[5999]), .B(c5999), .Z(n17999) );
XOR U30000 ( .A(c6000), .B(n18000), .Z(c6001) );
ANDN U30001 ( .B(n18001), .A(n18002), .Z(n18000) );
XOR U30002 ( .A(c6000), .B(b[6000]), .Z(n18001) );
XNOR U30003 ( .A(b[6000]), .B(n18002), .Z(c[6000]) );
XNOR U30004 ( .A(a[6000]), .B(c6000), .Z(n18002) );
XOR U30005 ( .A(c6001), .B(n18003), .Z(c6002) );
ANDN U30006 ( .B(n18004), .A(n18005), .Z(n18003) );
XOR U30007 ( .A(c6001), .B(b[6001]), .Z(n18004) );
XNOR U30008 ( .A(b[6001]), .B(n18005), .Z(c[6001]) );
XNOR U30009 ( .A(a[6001]), .B(c6001), .Z(n18005) );
XOR U30010 ( .A(c6002), .B(n18006), .Z(c6003) );
ANDN U30011 ( .B(n18007), .A(n18008), .Z(n18006) );
XOR U30012 ( .A(c6002), .B(b[6002]), .Z(n18007) );
XNOR U30013 ( .A(b[6002]), .B(n18008), .Z(c[6002]) );
XNOR U30014 ( .A(a[6002]), .B(c6002), .Z(n18008) );
XOR U30015 ( .A(c6003), .B(n18009), .Z(c6004) );
ANDN U30016 ( .B(n18010), .A(n18011), .Z(n18009) );
XOR U30017 ( .A(c6003), .B(b[6003]), .Z(n18010) );
XNOR U30018 ( .A(b[6003]), .B(n18011), .Z(c[6003]) );
XNOR U30019 ( .A(a[6003]), .B(c6003), .Z(n18011) );
XOR U30020 ( .A(c6004), .B(n18012), .Z(c6005) );
ANDN U30021 ( .B(n18013), .A(n18014), .Z(n18012) );
XOR U30022 ( .A(c6004), .B(b[6004]), .Z(n18013) );
XNOR U30023 ( .A(b[6004]), .B(n18014), .Z(c[6004]) );
XNOR U30024 ( .A(a[6004]), .B(c6004), .Z(n18014) );
XOR U30025 ( .A(c6005), .B(n18015), .Z(c6006) );
ANDN U30026 ( .B(n18016), .A(n18017), .Z(n18015) );
XOR U30027 ( .A(c6005), .B(b[6005]), .Z(n18016) );
XNOR U30028 ( .A(b[6005]), .B(n18017), .Z(c[6005]) );
XNOR U30029 ( .A(a[6005]), .B(c6005), .Z(n18017) );
XOR U30030 ( .A(c6006), .B(n18018), .Z(c6007) );
ANDN U30031 ( .B(n18019), .A(n18020), .Z(n18018) );
XOR U30032 ( .A(c6006), .B(b[6006]), .Z(n18019) );
XNOR U30033 ( .A(b[6006]), .B(n18020), .Z(c[6006]) );
XNOR U30034 ( .A(a[6006]), .B(c6006), .Z(n18020) );
XOR U30035 ( .A(c6007), .B(n18021), .Z(c6008) );
ANDN U30036 ( .B(n18022), .A(n18023), .Z(n18021) );
XOR U30037 ( .A(c6007), .B(b[6007]), .Z(n18022) );
XNOR U30038 ( .A(b[6007]), .B(n18023), .Z(c[6007]) );
XNOR U30039 ( .A(a[6007]), .B(c6007), .Z(n18023) );
XOR U30040 ( .A(c6008), .B(n18024), .Z(c6009) );
ANDN U30041 ( .B(n18025), .A(n18026), .Z(n18024) );
XOR U30042 ( .A(c6008), .B(b[6008]), .Z(n18025) );
XNOR U30043 ( .A(b[6008]), .B(n18026), .Z(c[6008]) );
XNOR U30044 ( .A(a[6008]), .B(c6008), .Z(n18026) );
XOR U30045 ( .A(c6009), .B(n18027), .Z(c6010) );
ANDN U30046 ( .B(n18028), .A(n18029), .Z(n18027) );
XOR U30047 ( .A(c6009), .B(b[6009]), .Z(n18028) );
XNOR U30048 ( .A(b[6009]), .B(n18029), .Z(c[6009]) );
XNOR U30049 ( .A(a[6009]), .B(c6009), .Z(n18029) );
XOR U30050 ( .A(c6010), .B(n18030), .Z(c6011) );
ANDN U30051 ( .B(n18031), .A(n18032), .Z(n18030) );
XOR U30052 ( .A(c6010), .B(b[6010]), .Z(n18031) );
XNOR U30053 ( .A(b[6010]), .B(n18032), .Z(c[6010]) );
XNOR U30054 ( .A(a[6010]), .B(c6010), .Z(n18032) );
XOR U30055 ( .A(c6011), .B(n18033), .Z(c6012) );
ANDN U30056 ( .B(n18034), .A(n18035), .Z(n18033) );
XOR U30057 ( .A(c6011), .B(b[6011]), .Z(n18034) );
XNOR U30058 ( .A(b[6011]), .B(n18035), .Z(c[6011]) );
XNOR U30059 ( .A(a[6011]), .B(c6011), .Z(n18035) );
XOR U30060 ( .A(c6012), .B(n18036), .Z(c6013) );
ANDN U30061 ( .B(n18037), .A(n18038), .Z(n18036) );
XOR U30062 ( .A(c6012), .B(b[6012]), .Z(n18037) );
XNOR U30063 ( .A(b[6012]), .B(n18038), .Z(c[6012]) );
XNOR U30064 ( .A(a[6012]), .B(c6012), .Z(n18038) );
XOR U30065 ( .A(c6013), .B(n18039), .Z(c6014) );
ANDN U30066 ( .B(n18040), .A(n18041), .Z(n18039) );
XOR U30067 ( .A(c6013), .B(b[6013]), .Z(n18040) );
XNOR U30068 ( .A(b[6013]), .B(n18041), .Z(c[6013]) );
XNOR U30069 ( .A(a[6013]), .B(c6013), .Z(n18041) );
XOR U30070 ( .A(c6014), .B(n18042), .Z(c6015) );
ANDN U30071 ( .B(n18043), .A(n18044), .Z(n18042) );
XOR U30072 ( .A(c6014), .B(b[6014]), .Z(n18043) );
XNOR U30073 ( .A(b[6014]), .B(n18044), .Z(c[6014]) );
XNOR U30074 ( .A(a[6014]), .B(c6014), .Z(n18044) );
XOR U30075 ( .A(c6015), .B(n18045), .Z(c6016) );
ANDN U30076 ( .B(n18046), .A(n18047), .Z(n18045) );
XOR U30077 ( .A(c6015), .B(b[6015]), .Z(n18046) );
XNOR U30078 ( .A(b[6015]), .B(n18047), .Z(c[6015]) );
XNOR U30079 ( .A(a[6015]), .B(c6015), .Z(n18047) );
XOR U30080 ( .A(c6016), .B(n18048), .Z(c6017) );
ANDN U30081 ( .B(n18049), .A(n18050), .Z(n18048) );
XOR U30082 ( .A(c6016), .B(b[6016]), .Z(n18049) );
XNOR U30083 ( .A(b[6016]), .B(n18050), .Z(c[6016]) );
XNOR U30084 ( .A(a[6016]), .B(c6016), .Z(n18050) );
XOR U30085 ( .A(c6017), .B(n18051), .Z(c6018) );
ANDN U30086 ( .B(n18052), .A(n18053), .Z(n18051) );
XOR U30087 ( .A(c6017), .B(b[6017]), .Z(n18052) );
XNOR U30088 ( .A(b[6017]), .B(n18053), .Z(c[6017]) );
XNOR U30089 ( .A(a[6017]), .B(c6017), .Z(n18053) );
XOR U30090 ( .A(c6018), .B(n18054), .Z(c6019) );
ANDN U30091 ( .B(n18055), .A(n18056), .Z(n18054) );
XOR U30092 ( .A(c6018), .B(b[6018]), .Z(n18055) );
XNOR U30093 ( .A(b[6018]), .B(n18056), .Z(c[6018]) );
XNOR U30094 ( .A(a[6018]), .B(c6018), .Z(n18056) );
XOR U30095 ( .A(c6019), .B(n18057), .Z(c6020) );
ANDN U30096 ( .B(n18058), .A(n18059), .Z(n18057) );
XOR U30097 ( .A(c6019), .B(b[6019]), .Z(n18058) );
XNOR U30098 ( .A(b[6019]), .B(n18059), .Z(c[6019]) );
XNOR U30099 ( .A(a[6019]), .B(c6019), .Z(n18059) );
XOR U30100 ( .A(c6020), .B(n18060), .Z(c6021) );
ANDN U30101 ( .B(n18061), .A(n18062), .Z(n18060) );
XOR U30102 ( .A(c6020), .B(b[6020]), .Z(n18061) );
XNOR U30103 ( .A(b[6020]), .B(n18062), .Z(c[6020]) );
XNOR U30104 ( .A(a[6020]), .B(c6020), .Z(n18062) );
XOR U30105 ( .A(c6021), .B(n18063), .Z(c6022) );
ANDN U30106 ( .B(n18064), .A(n18065), .Z(n18063) );
XOR U30107 ( .A(c6021), .B(b[6021]), .Z(n18064) );
XNOR U30108 ( .A(b[6021]), .B(n18065), .Z(c[6021]) );
XNOR U30109 ( .A(a[6021]), .B(c6021), .Z(n18065) );
XOR U30110 ( .A(c6022), .B(n18066), .Z(c6023) );
ANDN U30111 ( .B(n18067), .A(n18068), .Z(n18066) );
XOR U30112 ( .A(c6022), .B(b[6022]), .Z(n18067) );
XNOR U30113 ( .A(b[6022]), .B(n18068), .Z(c[6022]) );
XNOR U30114 ( .A(a[6022]), .B(c6022), .Z(n18068) );
XOR U30115 ( .A(c6023), .B(n18069), .Z(c6024) );
ANDN U30116 ( .B(n18070), .A(n18071), .Z(n18069) );
XOR U30117 ( .A(c6023), .B(b[6023]), .Z(n18070) );
XNOR U30118 ( .A(b[6023]), .B(n18071), .Z(c[6023]) );
XNOR U30119 ( .A(a[6023]), .B(c6023), .Z(n18071) );
XOR U30120 ( .A(c6024), .B(n18072), .Z(c6025) );
ANDN U30121 ( .B(n18073), .A(n18074), .Z(n18072) );
XOR U30122 ( .A(c6024), .B(b[6024]), .Z(n18073) );
XNOR U30123 ( .A(b[6024]), .B(n18074), .Z(c[6024]) );
XNOR U30124 ( .A(a[6024]), .B(c6024), .Z(n18074) );
XOR U30125 ( .A(c6025), .B(n18075), .Z(c6026) );
ANDN U30126 ( .B(n18076), .A(n18077), .Z(n18075) );
XOR U30127 ( .A(c6025), .B(b[6025]), .Z(n18076) );
XNOR U30128 ( .A(b[6025]), .B(n18077), .Z(c[6025]) );
XNOR U30129 ( .A(a[6025]), .B(c6025), .Z(n18077) );
XOR U30130 ( .A(c6026), .B(n18078), .Z(c6027) );
ANDN U30131 ( .B(n18079), .A(n18080), .Z(n18078) );
XOR U30132 ( .A(c6026), .B(b[6026]), .Z(n18079) );
XNOR U30133 ( .A(b[6026]), .B(n18080), .Z(c[6026]) );
XNOR U30134 ( .A(a[6026]), .B(c6026), .Z(n18080) );
XOR U30135 ( .A(c6027), .B(n18081), .Z(c6028) );
ANDN U30136 ( .B(n18082), .A(n18083), .Z(n18081) );
XOR U30137 ( .A(c6027), .B(b[6027]), .Z(n18082) );
XNOR U30138 ( .A(b[6027]), .B(n18083), .Z(c[6027]) );
XNOR U30139 ( .A(a[6027]), .B(c6027), .Z(n18083) );
XOR U30140 ( .A(c6028), .B(n18084), .Z(c6029) );
ANDN U30141 ( .B(n18085), .A(n18086), .Z(n18084) );
XOR U30142 ( .A(c6028), .B(b[6028]), .Z(n18085) );
XNOR U30143 ( .A(b[6028]), .B(n18086), .Z(c[6028]) );
XNOR U30144 ( .A(a[6028]), .B(c6028), .Z(n18086) );
XOR U30145 ( .A(c6029), .B(n18087), .Z(c6030) );
ANDN U30146 ( .B(n18088), .A(n18089), .Z(n18087) );
XOR U30147 ( .A(c6029), .B(b[6029]), .Z(n18088) );
XNOR U30148 ( .A(b[6029]), .B(n18089), .Z(c[6029]) );
XNOR U30149 ( .A(a[6029]), .B(c6029), .Z(n18089) );
XOR U30150 ( .A(c6030), .B(n18090), .Z(c6031) );
ANDN U30151 ( .B(n18091), .A(n18092), .Z(n18090) );
XOR U30152 ( .A(c6030), .B(b[6030]), .Z(n18091) );
XNOR U30153 ( .A(b[6030]), .B(n18092), .Z(c[6030]) );
XNOR U30154 ( .A(a[6030]), .B(c6030), .Z(n18092) );
XOR U30155 ( .A(c6031), .B(n18093), .Z(c6032) );
ANDN U30156 ( .B(n18094), .A(n18095), .Z(n18093) );
XOR U30157 ( .A(c6031), .B(b[6031]), .Z(n18094) );
XNOR U30158 ( .A(b[6031]), .B(n18095), .Z(c[6031]) );
XNOR U30159 ( .A(a[6031]), .B(c6031), .Z(n18095) );
XOR U30160 ( .A(c6032), .B(n18096), .Z(c6033) );
ANDN U30161 ( .B(n18097), .A(n18098), .Z(n18096) );
XOR U30162 ( .A(c6032), .B(b[6032]), .Z(n18097) );
XNOR U30163 ( .A(b[6032]), .B(n18098), .Z(c[6032]) );
XNOR U30164 ( .A(a[6032]), .B(c6032), .Z(n18098) );
XOR U30165 ( .A(c6033), .B(n18099), .Z(c6034) );
ANDN U30166 ( .B(n18100), .A(n18101), .Z(n18099) );
XOR U30167 ( .A(c6033), .B(b[6033]), .Z(n18100) );
XNOR U30168 ( .A(b[6033]), .B(n18101), .Z(c[6033]) );
XNOR U30169 ( .A(a[6033]), .B(c6033), .Z(n18101) );
XOR U30170 ( .A(c6034), .B(n18102), .Z(c6035) );
ANDN U30171 ( .B(n18103), .A(n18104), .Z(n18102) );
XOR U30172 ( .A(c6034), .B(b[6034]), .Z(n18103) );
XNOR U30173 ( .A(b[6034]), .B(n18104), .Z(c[6034]) );
XNOR U30174 ( .A(a[6034]), .B(c6034), .Z(n18104) );
XOR U30175 ( .A(c6035), .B(n18105), .Z(c6036) );
ANDN U30176 ( .B(n18106), .A(n18107), .Z(n18105) );
XOR U30177 ( .A(c6035), .B(b[6035]), .Z(n18106) );
XNOR U30178 ( .A(b[6035]), .B(n18107), .Z(c[6035]) );
XNOR U30179 ( .A(a[6035]), .B(c6035), .Z(n18107) );
XOR U30180 ( .A(c6036), .B(n18108), .Z(c6037) );
ANDN U30181 ( .B(n18109), .A(n18110), .Z(n18108) );
XOR U30182 ( .A(c6036), .B(b[6036]), .Z(n18109) );
XNOR U30183 ( .A(b[6036]), .B(n18110), .Z(c[6036]) );
XNOR U30184 ( .A(a[6036]), .B(c6036), .Z(n18110) );
XOR U30185 ( .A(c6037), .B(n18111), .Z(c6038) );
ANDN U30186 ( .B(n18112), .A(n18113), .Z(n18111) );
XOR U30187 ( .A(c6037), .B(b[6037]), .Z(n18112) );
XNOR U30188 ( .A(b[6037]), .B(n18113), .Z(c[6037]) );
XNOR U30189 ( .A(a[6037]), .B(c6037), .Z(n18113) );
XOR U30190 ( .A(c6038), .B(n18114), .Z(c6039) );
ANDN U30191 ( .B(n18115), .A(n18116), .Z(n18114) );
XOR U30192 ( .A(c6038), .B(b[6038]), .Z(n18115) );
XNOR U30193 ( .A(b[6038]), .B(n18116), .Z(c[6038]) );
XNOR U30194 ( .A(a[6038]), .B(c6038), .Z(n18116) );
XOR U30195 ( .A(c6039), .B(n18117), .Z(c6040) );
ANDN U30196 ( .B(n18118), .A(n18119), .Z(n18117) );
XOR U30197 ( .A(c6039), .B(b[6039]), .Z(n18118) );
XNOR U30198 ( .A(b[6039]), .B(n18119), .Z(c[6039]) );
XNOR U30199 ( .A(a[6039]), .B(c6039), .Z(n18119) );
XOR U30200 ( .A(c6040), .B(n18120), .Z(c6041) );
ANDN U30201 ( .B(n18121), .A(n18122), .Z(n18120) );
XOR U30202 ( .A(c6040), .B(b[6040]), .Z(n18121) );
XNOR U30203 ( .A(b[6040]), .B(n18122), .Z(c[6040]) );
XNOR U30204 ( .A(a[6040]), .B(c6040), .Z(n18122) );
XOR U30205 ( .A(c6041), .B(n18123), .Z(c6042) );
ANDN U30206 ( .B(n18124), .A(n18125), .Z(n18123) );
XOR U30207 ( .A(c6041), .B(b[6041]), .Z(n18124) );
XNOR U30208 ( .A(b[6041]), .B(n18125), .Z(c[6041]) );
XNOR U30209 ( .A(a[6041]), .B(c6041), .Z(n18125) );
XOR U30210 ( .A(c6042), .B(n18126), .Z(c6043) );
ANDN U30211 ( .B(n18127), .A(n18128), .Z(n18126) );
XOR U30212 ( .A(c6042), .B(b[6042]), .Z(n18127) );
XNOR U30213 ( .A(b[6042]), .B(n18128), .Z(c[6042]) );
XNOR U30214 ( .A(a[6042]), .B(c6042), .Z(n18128) );
XOR U30215 ( .A(c6043), .B(n18129), .Z(c6044) );
ANDN U30216 ( .B(n18130), .A(n18131), .Z(n18129) );
XOR U30217 ( .A(c6043), .B(b[6043]), .Z(n18130) );
XNOR U30218 ( .A(b[6043]), .B(n18131), .Z(c[6043]) );
XNOR U30219 ( .A(a[6043]), .B(c6043), .Z(n18131) );
XOR U30220 ( .A(c6044), .B(n18132), .Z(c6045) );
ANDN U30221 ( .B(n18133), .A(n18134), .Z(n18132) );
XOR U30222 ( .A(c6044), .B(b[6044]), .Z(n18133) );
XNOR U30223 ( .A(b[6044]), .B(n18134), .Z(c[6044]) );
XNOR U30224 ( .A(a[6044]), .B(c6044), .Z(n18134) );
XOR U30225 ( .A(c6045), .B(n18135), .Z(c6046) );
ANDN U30226 ( .B(n18136), .A(n18137), .Z(n18135) );
XOR U30227 ( .A(c6045), .B(b[6045]), .Z(n18136) );
XNOR U30228 ( .A(b[6045]), .B(n18137), .Z(c[6045]) );
XNOR U30229 ( .A(a[6045]), .B(c6045), .Z(n18137) );
XOR U30230 ( .A(c6046), .B(n18138), .Z(c6047) );
ANDN U30231 ( .B(n18139), .A(n18140), .Z(n18138) );
XOR U30232 ( .A(c6046), .B(b[6046]), .Z(n18139) );
XNOR U30233 ( .A(b[6046]), .B(n18140), .Z(c[6046]) );
XNOR U30234 ( .A(a[6046]), .B(c6046), .Z(n18140) );
XOR U30235 ( .A(c6047), .B(n18141), .Z(c6048) );
ANDN U30236 ( .B(n18142), .A(n18143), .Z(n18141) );
XOR U30237 ( .A(c6047), .B(b[6047]), .Z(n18142) );
XNOR U30238 ( .A(b[6047]), .B(n18143), .Z(c[6047]) );
XNOR U30239 ( .A(a[6047]), .B(c6047), .Z(n18143) );
XOR U30240 ( .A(c6048), .B(n18144), .Z(c6049) );
ANDN U30241 ( .B(n18145), .A(n18146), .Z(n18144) );
XOR U30242 ( .A(c6048), .B(b[6048]), .Z(n18145) );
XNOR U30243 ( .A(b[6048]), .B(n18146), .Z(c[6048]) );
XNOR U30244 ( .A(a[6048]), .B(c6048), .Z(n18146) );
XOR U30245 ( .A(c6049), .B(n18147), .Z(c6050) );
ANDN U30246 ( .B(n18148), .A(n18149), .Z(n18147) );
XOR U30247 ( .A(c6049), .B(b[6049]), .Z(n18148) );
XNOR U30248 ( .A(b[6049]), .B(n18149), .Z(c[6049]) );
XNOR U30249 ( .A(a[6049]), .B(c6049), .Z(n18149) );
XOR U30250 ( .A(c6050), .B(n18150), .Z(c6051) );
ANDN U30251 ( .B(n18151), .A(n18152), .Z(n18150) );
XOR U30252 ( .A(c6050), .B(b[6050]), .Z(n18151) );
XNOR U30253 ( .A(b[6050]), .B(n18152), .Z(c[6050]) );
XNOR U30254 ( .A(a[6050]), .B(c6050), .Z(n18152) );
XOR U30255 ( .A(c6051), .B(n18153), .Z(c6052) );
ANDN U30256 ( .B(n18154), .A(n18155), .Z(n18153) );
XOR U30257 ( .A(c6051), .B(b[6051]), .Z(n18154) );
XNOR U30258 ( .A(b[6051]), .B(n18155), .Z(c[6051]) );
XNOR U30259 ( .A(a[6051]), .B(c6051), .Z(n18155) );
XOR U30260 ( .A(c6052), .B(n18156), .Z(c6053) );
ANDN U30261 ( .B(n18157), .A(n18158), .Z(n18156) );
XOR U30262 ( .A(c6052), .B(b[6052]), .Z(n18157) );
XNOR U30263 ( .A(b[6052]), .B(n18158), .Z(c[6052]) );
XNOR U30264 ( .A(a[6052]), .B(c6052), .Z(n18158) );
XOR U30265 ( .A(c6053), .B(n18159), .Z(c6054) );
ANDN U30266 ( .B(n18160), .A(n18161), .Z(n18159) );
XOR U30267 ( .A(c6053), .B(b[6053]), .Z(n18160) );
XNOR U30268 ( .A(b[6053]), .B(n18161), .Z(c[6053]) );
XNOR U30269 ( .A(a[6053]), .B(c6053), .Z(n18161) );
XOR U30270 ( .A(c6054), .B(n18162), .Z(c6055) );
ANDN U30271 ( .B(n18163), .A(n18164), .Z(n18162) );
XOR U30272 ( .A(c6054), .B(b[6054]), .Z(n18163) );
XNOR U30273 ( .A(b[6054]), .B(n18164), .Z(c[6054]) );
XNOR U30274 ( .A(a[6054]), .B(c6054), .Z(n18164) );
XOR U30275 ( .A(c6055), .B(n18165), .Z(c6056) );
ANDN U30276 ( .B(n18166), .A(n18167), .Z(n18165) );
XOR U30277 ( .A(c6055), .B(b[6055]), .Z(n18166) );
XNOR U30278 ( .A(b[6055]), .B(n18167), .Z(c[6055]) );
XNOR U30279 ( .A(a[6055]), .B(c6055), .Z(n18167) );
XOR U30280 ( .A(c6056), .B(n18168), .Z(c6057) );
ANDN U30281 ( .B(n18169), .A(n18170), .Z(n18168) );
XOR U30282 ( .A(c6056), .B(b[6056]), .Z(n18169) );
XNOR U30283 ( .A(b[6056]), .B(n18170), .Z(c[6056]) );
XNOR U30284 ( .A(a[6056]), .B(c6056), .Z(n18170) );
XOR U30285 ( .A(c6057), .B(n18171), .Z(c6058) );
ANDN U30286 ( .B(n18172), .A(n18173), .Z(n18171) );
XOR U30287 ( .A(c6057), .B(b[6057]), .Z(n18172) );
XNOR U30288 ( .A(b[6057]), .B(n18173), .Z(c[6057]) );
XNOR U30289 ( .A(a[6057]), .B(c6057), .Z(n18173) );
XOR U30290 ( .A(c6058), .B(n18174), .Z(c6059) );
ANDN U30291 ( .B(n18175), .A(n18176), .Z(n18174) );
XOR U30292 ( .A(c6058), .B(b[6058]), .Z(n18175) );
XNOR U30293 ( .A(b[6058]), .B(n18176), .Z(c[6058]) );
XNOR U30294 ( .A(a[6058]), .B(c6058), .Z(n18176) );
XOR U30295 ( .A(c6059), .B(n18177), .Z(c6060) );
ANDN U30296 ( .B(n18178), .A(n18179), .Z(n18177) );
XOR U30297 ( .A(c6059), .B(b[6059]), .Z(n18178) );
XNOR U30298 ( .A(b[6059]), .B(n18179), .Z(c[6059]) );
XNOR U30299 ( .A(a[6059]), .B(c6059), .Z(n18179) );
XOR U30300 ( .A(c6060), .B(n18180), .Z(c6061) );
ANDN U30301 ( .B(n18181), .A(n18182), .Z(n18180) );
XOR U30302 ( .A(c6060), .B(b[6060]), .Z(n18181) );
XNOR U30303 ( .A(b[6060]), .B(n18182), .Z(c[6060]) );
XNOR U30304 ( .A(a[6060]), .B(c6060), .Z(n18182) );
XOR U30305 ( .A(c6061), .B(n18183), .Z(c6062) );
ANDN U30306 ( .B(n18184), .A(n18185), .Z(n18183) );
XOR U30307 ( .A(c6061), .B(b[6061]), .Z(n18184) );
XNOR U30308 ( .A(b[6061]), .B(n18185), .Z(c[6061]) );
XNOR U30309 ( .A(a[6061]), .B(c6061), .Z(n18185) );
XOR U30310 ( .A(c6062), .B(n18186), .Z(c6063) );
ANDN U30311 ( .B(n18187), .A(n18188), .Z(n18186) );
XOR U30312 ( .A(c6062), .B(b[6062]), .Z(n18187) );
XNOR U30313 ( .A(b[6062]), .B(n18188), .Z(c[6062]) );
XNOR U30314 ( .A(a[6062]), .B(c6062), .Z(n18188) );
XOR U30315 ( .A(c6063), .B(n18189), .Z(c6064) );
ANDN U30316 ( .B(n18190), .A(n18191), .Z(n18189) );
XOR U30317 ( .A(c6063), .B(b[6063]), .Z(n18190) );
XNOR U30318 ( .A(b[6063]), .B(n18191), .Z(c[6063]) );
XNOR U30319 ( .A(a[6063]), .B(c6063), .Z(n18191) );
XOR U30320 ( .A(c6064), .B(n18192), .Z(c6065) );
ANDN U30321 ( .B(n18193), .A(n18194), .Z(n18192) );
XOR U30322 ( .A(c6064), .B(b[6064]), .Z(n18193) );
XNOR U30323 ( .A(b[6064]), .B(n18194), .Z(c[6064]) );
XNOR U30324 ( .A(a[6064]), .B(c6064), .Z(n18194) );
XOR U30325 ( .A(c6065), .B(n18195), .Z(c6066) );
ANDN U30326 ( .B(n18196), .A(n18197), .Z(n18195) );
XOR U30327 ( .A(c6065), .B(b[6065]), .Z(n18196) );
XNOR U30328 ( .A(b[6065]), .B(n18197), .Z(c[6065]) );
XNOR U30329 ( .A(a[6065]), .B(c6065), .Z(n18197) );
XOR U30330 ( .A(c6066), .B(n18198), .Z(c6067) );
ANDN U30331 ( .B(n18199), .A(n18200), .Z(n18198) );
XOR U30332 ( .A(c6066), .B(b[6066]), .Z(n18199) );
XNOR U30333 ( .A(b[6066]), .B(n18200), .Z(c[6066]) );
XNOR U30334 ( .A(a[6066]), .B(c6066), .Z(n18200) );
XOR U30335 ( .A(c6067), .B(n18201), .Z(c6068) );
ANDN U30336 ( .B(n18202), .A(n18203), .Z(n18201) );
XOR U30337 ( .A(c6067), .B(b[6067]), .Z(n18202) );
XNOR U30338 ( .A(b[6067]), .B(n18203), .Z(c[6067]) );
XNOR U30339 ( .A(a[6067]), .B(c6067), .Z(n18203) );
XOR U30340 ( .A(c6068), .B(n18204), .Z(c6069) );
ANDN U30341 ( .B(n18205), .A(n18206), .Z(n18204) );
XOR U30342 ( .A(c6068), .B(b[6068]), .Z(n18205) );
XNOR U30343 ( .A(b[6068]), .B(n18206), .Z(c[6068]) );
XNOR U30344 ( .A(a[6068]), .B(c6068), .Z(n18206) );
XOR U30345 ( .A(c6069), .B(n18207), .Z(c6070) );
ANDN U30346 ( .B(n18208), .A(n18209), .Z(n18207) );
XOR U30347 ( .A(c6069), .B(b[6069]), .Z(n18208) );
XNOR U30348 ( .A(b[6069]), .B(n18209), .Z(c[6069]) );
XNOR U30349 ( .A(a[6069]), .B(c6069), .Z(n18209) );
XOR U30350 ( .A(c6070), .B(n18210), .Z(c6071) );
ANDN U30351 ( .B(n18211), .A(n18212), .Z(n18210) );
XOR U30352 ( .A(c6070), .B(b[6070]), .Z(n18211) );
XNOR U30353 ( .A(b[6070]), .B(n18212), .Z(c[6070]) );
XNOR U30354 ( .A(a[6070]), .B(c6070), .Z(n18212) );
XOR U30355 ( .A(c6071), .B(n18213), .Z(c6072) );
ANDN U30356 ( .B(n18214), .A(n18215), .Z(n18213) );
XOR U30357 ( .A(c6071), .B(b[6071]), .Z(n18214) );
XNOR U30358 ( .A(b[6071]), .B(n18215), .Z(c[6071]) );
XNOR U30359 ( .A(a[6071]), .B(c6071), .Z(n18215) );
XOR U30360 ( .A(c6072), .B(n18216), .Z(c6073) );
ANDN U30361 ( .B(n18217), .A(n18218), .Z(n18216) );
XOR U30362 ( .A(c6072), .B(b[6072]), .Z(n18217) );
XNOR U30363 ( .A(b[6072]), .B(n18218), .Z(c[6072]) );
XNOR U30364 ( .A(a[6072]), .B(c6072), .Z(n18218) );
XOR U30365 ( .A(c6073), .B(n18219), .Z(c6074) );
ANDN U30366 ( .B(n18220), .A(n18221), .Z(n18219) );
XOR U30367 ( .A(c6073), .B(b[6073]), .Z(n18220) );
XNOR U30368 ( .A(b[6073]), .B(n18221), .Z(c[6073]) );
XNOR U30369 ( .A(a[6073]), .B(c6073), .Z(n18221) );
XOR U30370 ( .A(c6074), .B(n18222), .Z(c6075) );
ANDN U30371 ( .B(n18223), .A(n18224), .Z(n18222) );
XOR U30372 ( .A(c6074), .B(b[6074]), .Z(n18223) );
XNOR U30373 ( .A(b[6074]), .B(n18224), .Z(c[6074]) );
XNOR U30374 ( .A(a[6074]), .B(c6074), .Z(n18224) );
XOR U30375 ( .A(c6075), .B(n18225), .Z(c6076) );
ANDN U30376 ( .B(n18226), .A(n18227), .Z(n18225) );
XOR U30377 ( .A(c6075), .B(b[6075]), .Z(n18226) );
XNOR U30378 ( .A(b[6075]), .B(n18227), .Z(c[6075]) );
XNOR U30379 ( .A(a[6075]), .B(c6075), .Z(n18227) );
XOR U30380 ( .A(c6076), .B(n18228), .Z(c6077) );
ANDN U30381 ( .B(n18229), .A(n18230), .Z(n18228) );
XOR U30382 ( .A(c6076), .B(b[6076]), .Z(n18229) );
XNOR U30383 ( .A(b[6076]), .B(n18230), .Z(c[6076]) );
XNOR U30384 ( .A(a[6076]), .B(c6076), .Z(n18230) );
XOR U30385 ( .A(c6077), .B(n18231), .Z(c6078) );
ANDN U30386 ( .B(n18232), .A(n18233), .Z(n18231) );
XOR U30387 ( .A(c6077), .B(b[6077]), .Z(n18232) );
XNOR U30388 ( .A(b[6077]), .B(n18233), .Z(c[6077]) );
XNOR U30389 ( .A(a[6077]), .B(c6077), .Z(n18233) );
XOR U30390 ( .A(c6078), .B(n18234), .Z(c6079) );
ANDN U30391 ( .B(n18235), .A(n18236), .Z(n18234) );
XOR U30392 ( .A(c6078), .B(b[6078]), .Z(n18235) );
XNOR U30393 ( .A(b[6078]), .B(n18236), .Z(c[6078]) );
XNOR U30394 ( .A(a[6078]), .B(c6078), .Z(n18236) );
XOR U30395 ( .A(c6079), .B(n18237), .Z(c6080) );
ANDN U30396 ( .B(n18238), .A(n18239), .Z(n18237) );
XOR U30397 ( .A(c6079), .B(b[6079]), .Z(n18238) );
XNOR U30398 ( .A(b[6079]), .B(n18239), .Z(c[6079]) );
XNOR U30399 ( .A(a[6079]), .B(c6079), .Z(n18239) );
XOR U30400 ( .A(c6080), .B(n18240), .Z(c6081) );
ANDN U30401 ( .B(n18241), .A(n18242), .Z(n18240) );
XOR U30402 ( .A(c6080), .B(b[6080]), .Z(n18241) );
XNOR U30403 ( .A(b[6080]), .B(n18242), .Z(c[6080]) );
XNOR U30404 ( .A(a[6080]), .B(c6080), .Z(n18242) );
XOR U30405 ( .A(c6081), .B(n18243), .Z(c6082) );
ANDN U30406 ( .B(n18244), .A(n18245), .Z(n18243) );
XOR U30407 ( .A(c6081), .B(b[6081]), .Z(n18244) );
XNOR U30408 ( .A(b[6081]), .B(n18245), .Z(c[6081]) );
XNOR U30409 ( .A(a[6081]), .B(c6081), .Z(n18245) );
XOR U30410 ( .A(c6082), .B(n18246), .Z(c6083) );
ANDN U30411 ( .B(n18247), .A(n18248), .Z(n18246) );
XOR U30412 ( .A(c6082), .B(b[6082]), .Z(n18247) );
XNOR U30413 ( .A(b[6082]), .B(n18248), .Z(c[6082]) );
XNOR U30414 ( .A(a[6082]), .B(c6082), .Z(n18248) );
XOR U30415 ( .A(c6083), .B(n18249), .Z(c6084) );
ANDN U30416 ( .B(n18250), .A(n18251), .Z(n18249) );
XOR U30417 ( .A(c6083), .B(b[6083]), .Z(n18250) );
XNOR U30418 ( .A(b[6083]), .B(n18251), .Z(c[6083]) );
XNOR U30419 ( .A(a[6083]), .B(c6083), .Z(n18251) );
XOR U30420 ( .A(c6084), .B(n18252), .Z(c6085) );
ANDN U30421 ( .B(n18253), .A(n18254), .Z(n18252) );
XOR U30422 ( .A(c6084), .B(b[6084]), .Z(n18253) );
XNOR U30423 ( .A(b[6084]), .B(n18254), .Z(c[6084]) );
XNOR U30424 ( .A(a[6084]), .B(c6084), .Z(n18254) );
XOR U30425 ( .A(c6085), .B(n18255), .Z(c6086) );
ANDN U30426 ( .B(n18256), .A(n18257), .Z(n18255) );
XOR U30427 ( .A(c6085), .B(b[6085]), .Z(n18256) );
XNOR U30428 ( .A(b[6085]), .B(n18257), .Z(c[6085]) );
XNOR U30429 ( .A(a[6085]), .B(c6085), .Z(n18257) );
XOR U30430 ( .A(c6086), .B(n18258), .Z(c6087) );
ANDN U30431 ( .B(n18259), .A(n18260), .Z(n18258) );
XOR U30432 ( .A(c6086), .B(b[6086]), .Z(n18259) );
XNOR U30433 ( .A(b[6086]), .B(n18260), .Z(c[6086]) );
XNOR U30434 ( .A(a[6086]), .B(c6086), .Z(n18260) );
XOR U30435 ( .A(c6087), .B(n18261), .Z(c6088) );
ANDN U30436 ( .B(n18262), .A(n18263), .Z(n18261) );
XOR U30437 ( .A(c6087), .B(b[6087]), .Z(n18262) );
XNOR U30438 ( .A(b[6087]), .B(n18263), .Z(c[6087]) );
XNOR U30439 ( .A(a[6087]), .B(c6087), .Z(n18263) );
XOR U30440 ( .A(c6088), .B(n18264), .Z(c6089) );
ANDN U30441 ( .B(n18265), .A(n18266), .Z(n18264) );
XOR U30442 ( .A(c6088), .B(b[6088]), .Z(n18265) );
XNOR U30443 ( .A(b[6088]), .B(n18266), .Z(c[6088]) );
XNOR U30444 ( .A(a[6088]), .B(c6088), .Z(n18266) );
XOR U30445 ( .A(c6089), .B(n18267), .Z(c6090) );
ANDN U30446 ( .B(n18268), .A(n18269), .Z(n18267) );
XOR U30447 ( .A(c6089), .B(b[6089]), .Z(n18268) );
XNOR U30448 ( .A(b[6089]), .B(n18269), .Z(c[6089]) );
XNOR U30449 ( .A(a[6089]), .B(c6089), .Z(n18269) );
XOR U30450 ( .A(c6090), .B(n18270), .Z(c6091) );
ANDN U30451 ( .B(n18271), .A(n18272), .Z(n18270) );
XOR U30452 ( .A(c6090), .B(b[6090]), .Z(n18271) );
XNOR U30453 ( .A(b[6090]), .B(n18272), .Z(c[6090]) );
XNOR U30454 ( .A(a[6090]), .B(c6090), .Z(n18272) );
XOR U30455 ( .A(c6091), .B(n18273), .Z(c6092) );
ANDN U30456 ( .B(n18274), .A(n18275), .Z(n18273) );
XOR U30457 ( .A(c6091), .B(b[6091]), .Z(n18274) );
XNOR U30458 ( .A(b[6091]), .B(n18275), .Z(c[6091]) );
XNOR U30459 ( .A(a[6091]), .B(c6091), .Z(n18275) );
XOR U30460 ( .A(c6092), .B(n18276), .Z(c6093) );
ANDN U30461 ( .B(n18277), .A(n18278), .Z(n18276) );
XOR U30462 ( .A(c6092), .B(b[6092]), .Z(n18277) );
XNOR U30463 ( .A(b[6092]), .B(n18278), .Z(c[6092]) );
XNOR U30464 ( .A(a[6092]), .B(c6092), .Z(n18278) );
XOR U30465 ( .A(c6093), .B(n18279), .Z(c6094) );
ANDN U30466 ( .B(n18280), .A(n18281), .Z(n18279) );
XOR U30467 ( .A(c6093), .B(b[6093]), .Z(n18280) );
XNOR U30468 ( .A(b[6093]), .B(n18281), .Z(c[6093]) );
XNOR U30469 ( .A(a[6093]), .B(c6093), .Z(n18281) );
XOR U30470 ( .A(c6094), .B(n18282), .Z(c6095) );
ANDN U30471 ( .B(n18283), .A(n18284), .Z(n18282) );
XOR U30472 ( .A(c6094), .B(b[6094]), .Z(n18283) );
XNOR U30473 ( .A(b[6094]), .B(n18284), .Z(c[6094]) );
XNOR U30474 ( .A(a[6094]), .B(c6094), .Z(n18284) );
XOR U30475 ( .A(c6095), .B(n18285), .Z(c6096) );
ANDN U30476 ( .B(n18286), .A(n18287), .Z(n18285) );
XOR U30477 ( .A(c6095), .B(b[6095]), .Z(n18286) );
XNOR U30478 ( .A(b[6095]), .B(n18287), .Z(c[6095]) );
XNOR U30479 ( .A(a[6095]), .B(c6095), .Z(n18287) );
XOR U30480 ( .A(c6096), .B(n18288), .Z(c6097) );
ANDN U30481 ( .B(n18289), .A(n18290), .Z(n18288) );
XOR U30482 ( .A(c6096), .B(b[6096]), .Z(n18289) );
XNOR U30483 ( .A(b[6096]), .B(n18290), .Z(c[6096]) );
XNOR U30484 ( .A(a[6096]), .B(c6096), .Z(n18290) );
XOR U30485 ( .A(c6097), .B(n18291), .Z(c6098) );
ANDN U30486 ( .B(n18292), .A(n18293), .Z(n18291) );
XOR U30487 ( .A(c6097), .B(b[6097]), .Z(n18292) );
XNOR U30488 ( .A(b[6097]), .B(n18293), .Z(c[6097]) );
XNOR U30489 ( .A(a[6097]), .B(c6097), .Z(n18293) );
XOR U30490 ( .A(c6098), .B(n18294), .Z(c6099) );
ANDN U30491 ( .B(n18295), .A(n18296), .Z(n18294) );
XOR U30492 ( .A(c6098), .B(b[6098]), .Z(n18295) );
XNOR U30493 ( .A(b[6098]), .B(n18296), .Z(c[6098]) );
XNOR U30494 ( .A(a[6098]), .B(c6098), .Z(n18296) );
XOR U30495 ( .A(c6099), .B(n18297), .Z(c6100) );
ANDN U30496 ( .B(n18298), .A(n18299), .Z(n18297) );
XOR U30497 ( .A(c6099), .B(b[6099]), .Z(n18298) );
XNOR U30498 ( .A(b[6099]), .B(n18299), .Z(c[6099]) );
XNOR U30499 ( .A(a[6099]), .B(c6099), .Z(n18299) );
XOR U30500 ( .A(c6100), .B(n18300), .Z(c6101) );
ANDN U30501 ( .B(n18301), .A(n18302), .Z(n18300) );
XOR U30502 ( .A(c6100), .B(b[6100]), .Z(n18301) );
XNOR U30503 ( .A(b[6100]), .B(n18302), .Z(c[6100]) );
XNOR U30504 ( .A(a[6100]), .B(c6100), .Z(n18302) );
XOR U30505 ( .A(c6101), .B(n18303), .Z(c6102) );
ANDN U30506 ( .B(n18304), .A(n18305), .Z(n18303) );
XOR U30507 ( .A(c6101), .B(b[6101]), .Z(n18304) );
XNOR U30508 ( .A(b[6101]), .B(n18305), .Z(c[6101]) );
XNOR U30509 ( .A(a[6101]), .B(c6101), .Z(n18305) );
XOR U30510 ( .A(c6102), .B(n18306), .Z(c6103) );
ANDN U30511 ( .B(n18307), .A(n18308), .Z(n18306) );
XOR U30512 ( .A(c6102), .B(b[6102]), .Z(n18307) );
XNOR U30513 ( .A(b[6102]), .B(n18308), .Z(c[6102]) );
XNOR U30514 ( .A(a[6102]), .B(c6102), .Z(n18308) );
XOR U30515 ( .A(c6103), .B(n18309), .Z(c6104) );
ANDN U30516 ( .B(n18310), .A(n18311), .Z(n18309) );
XOR U30517 ( .A(c6103), .B(b[6103]), .Z(n18310) );
XNOR U30518 ( .A(b[6103]), .B(n18311), .Z(c[6103]) );
XNOR U30519 ( .A(a[6103]), .B(c6103), .Z(n18311) );
XOR U30520 ( .A(c6104), .B(n18312), .Z(c6105) );
ANDN U30521 ( .B(n18313), .A(n18314), .Z(n18312) );
XOR U30522 ( .A(c6104), .B(b[6104]), .Z(n18313) );
XNOR U30523 ( .A(b[6104]), .B(n18314), .Z(c[6104]) );
XNOR U30524 ( .A(a[6104]), .B(c6104), .Z(n18314) );
XOR U30525 ( .A(c6105), .B(n18315), .Z(c6106) );
ANDN U30526 ( .B(n18316), .A(n18317), .Z(n18315) );
XOR U30527 ( .A(c6105), .B(b[6105]), .Z(n18316) );
XNOR U30528 ( .A(b[6105]), .B(n18317), .Z(c[6105]) );
XNOR U30529 ( .A(a[6105]), .B(c6105), .Z(n18317) );
XOR U30530 ( .A(c6106), .B(n18318), .Z(c6107) );
ANDN U30531 ( .B(n18319), .A(n18320), .Z(n18318) );
XOR U30532 ( .A(c6106), .B(b[6106]), .Z(n18319) );
XNOR U30533 ( .A(b[6106]), .B(n18320), .Z(c[6106]) );
XNOR U30534 ( .A(a[6106]), .B(c6106), .Z(n18320) );
XOR U30535 ( .A(c6107), .B(n18321), .Z(c6108) );
ANDN U30536 ( .B(n18322), .A(n18323), .Z(n18321) );
XOR U30537 ( .A(c6107), .B(b[6107]), .Z(n18322) );
XNOR U30538 ( .A(b[6107]), .B(n18323), .Z(c[6107]) );
XNOR U30539 ( .A(a[6107]), .B(c6107), .Z(n18323) );
XOR U30540 ( .A(c6108), .B(n18324), .Z(c6109) );
ANDN U30541 ( .B(n18325), .A(n18326), .Z(n18324) );
XOR U30542 ( .A(c6108), .B(b[6108]), .Z(n18325) );
XNOR U30543 ( .A(b[6108]), .B(n18326), .Z(c[6108]) );
XNOR U30544 ( .A(a[6108]), .B(c6108), .Z(n18326) );
XOR U30545 ( .A(c6109), .B(n18327), .Z(c6110) );
ANDN U30546 ( .B(n18328), .A(n18329), .Z(n18327) );
XOR U30547 ( .A(c6109), .B(b[6109]), .Z(n18328) );
XNOR U30548 ( .A(b[6109]), .B(n18329), .Z(c[6109]) );
XNOR U30549 ( .A(a[6109]), .B(c6109), .Z(n18329) );
XOR U30550 ( .A(c6110), .B(n18330), .Z(c6111) );
ANDN U30551 ( .B(n18331), .A(n18332), .Z(n18330) );
XOR U30552 ( .A(c6110), .B(b[6110]), .Z(n18331) );
XNOR U30553 ( .A(b[6110]), .B(n18332), .Z(c[6110]) );
XNOR U30554 ( .A(a[6110]), .B(c6110), .Z(n18332) );
XOR U30555 ( .A(c6111), .B(n18333), .Z(c6112) );
ANDN U30556 ( .B(n18334), .A(n18335), .Z(n18333) );
XOR U30557 ( .A(c6111), .B(b[6111]), .Z(n18334) );
XNOR U30558 ( .A(b[6111]), .B(n18335), .Z(c[6111]) );
XNOR U30559 ( .A(a[6111]), .B(c6111), .Z(n18335) );
XOR U30560 ( .A(c6112), .B(n18336), .Z(c6113) );
ANDN U30561 ( .B(n18337), .A(n18338), .Z(n18336) );
XOR U30562 ( .A(c6112), .B(b[6112]), .Z(n18337) );
XNOR U30563 ( .A(b[6112]), .B(n18338), .Z(c[6112]) );
XNOR U30564 ( .A(a[6112]), .B(c6112), .Z(n18338) );
XOR U30565 ( .A(c6113), .B(n18339), .Z(c6114) );
ANDN U30566 ( .B(n18340), .A(n18341), .Z(n18339) );
XOR U30567 ( .A(c6113), .B(b[6113]), .Z(n18340) );
XNOR U30568 ( .A(b[6113]), .B(n18341), .Z(c[6113]) );
XNOR U30569 ( .A(a[6113]), .B(c6113), .Z(n18341) );
XOR U30570 ( .A(c6114), .B(n18342), .Z(c6115) );
ANDN U30571 ( .B(n18343), .A(n18344), .Z(n18342) );
XOR U30572 ( .A(c6114), .B(b[6114]), .Z(n18343) );
XNOR U30573 ( .A(b[6114]), .B(n18344), .Z(c[6114]) );
XNOR U30574 ( .A(a[6114]), .B(c6114), .Z(n18344) );
XOR U30575 ( .A(c6115), .B(n18345), .Z(c6116) );
ANDN U30576 ( .B(n18346), .A(n18347), .Z(n18345) );
XOR U30577 ( .A(c6115), .B(b[6115]), .Z(n18346) );
XNOR U30578 ( .A(b[6115]), .B(n18347), .Z(c[6115]) );
XNOR U30579 ( .A(a[6115]), .B(c6115), .Z(n18347) );
XOR U30580 ( .A(c6116), .B(n18348), .Z(c6117) );
ANDN U30581 ( .B(n18349), .A(n18350), .Z(n18348) );
XOR U30582 ( .A(c6116), .B(b[6116]), .Z(n18349) );
XNOR U30583 ( .A(b[6116]), .B(n18350), .Z(c[6116]) );
XNOR U30584 ( .A(a[6116]), .B(c6116), .Z(n18350) );
XOR U30585 ( .A(c6117), .B(n18351), .Z(c6118) );
ANDN U30586 ( .B(n18352), .A(n18353), .Z(n18351) );
XOR U30587 ( .A(c6117), .B(b[6117]), .Z(n18352) );
XNOR U30588 ( .A(b[6117]), .B(n18353), .Z(c[6117]) );
XNOR U30589 ( .A(a[6117]), .B(c6117), .Z(n18353) );
XOR U30590 ( .A(c6118), .B(n18354), .Z(c6119) );
ANDN U30591 ( .B(n18355), .A(n18356), .Z(n18354) );
XOR U30592 ( .A(c6118), .B(b[6118]), .Z(n18355) );
XNOR U30593 ( .A(b[6118]), .B(n18356), .Z(c[6118]) );
XNOR U30594 ( .A(a[6118]), .B(c6118), .Z(n18356) );
XOR U30595 ( .A(c6119), .B(n18357), .Z(c6120) );
ANDN U30596 ( .B(n18358), .A(n18359), .Z(n18357) );
XOR U30597 ( .A(c6119), .B(b[6119]), .Z(n18358) );
XNOR U30598 ( .A(b[6119]), .B(n18359), .Z(c[6119]) );
XNOR U30599 ( .A(a[6119]), .B(c6119), .Z(n18359) );
XOR U30600 ( .A(c6120), .B(n18360), .Z(c6121) );
ANDN U30601 ( .B(n18361), .A(n18362), .Z(n18360) );
XOR U30602 ( .A(c6120), .B(b[6120]), .Z(n18361) );
XNOR U30603 ( .A(b[6120]), .B(n18362), .Z(c[6120]) );
XNOR U30604 ( .A(a[6120]), .B(c6120), .Z(n18362) );
XOR U30605 ( .A(c6121), .B(n18363), .Z(c6122) );
ANDN U30606 ( .B(n18364), .A(n18365), .Z(n18363) );
XOR U30607 ( .A(c6121), .B(b[6121]), .Z(n18364) );
XNOR U30608 ( .A(b[6121]), .B(n18365), .Z(c[6121]) );
XNOR U30609 ( .A(a[6121]), .B(c6121), .Z(n18365) );
XOR U30610 ( .A(c6122), .B(n18366), .Z(c6123) );
ANDN U30611 ( .B(n18367), .A(n18368), .Z(n18366) );
XOR U30612 ( .A(c6122), .B(b[6122]), .Z(n18367) );
XNOR U30613 ( .A(b[6122]), .B(n18368), .Z(c[6122]) );
XNOR U30614 ( .A(a[6122]), .B(c6122), .Z(n18368) );
XOR U30615 ( .A(c6123), .B(n18369), .Z(c6124) );
ANDN U30616 ( .B(n18370), .A(n18371), .Z(n18369) );
XOR U30617 ( .A(c6123), .B(b[6123]), .Z(n18370) );
XNOR U30618 ( .A(b[6123]), .B(n18371), .Z(c[6123]) );
XNOR U30619 ( .A(a[6123]), .B(c6123), .Z(n18371) );
XOR U30620 ( .A(c6124), .B(n18372), .Z(c6125) );
ANDN U30621 ( .B(n18373), .A(n18374), .Z(n18372) );
XOR U30622 ( .A(c6124), .B(b[6124]), .Z(n18373) );
XNOR U30623 ( .A(b[6124]), .B(n18374), .Z(c[6124]) );
XNOR U30624 ( .A(a[6124]), .B(c6124), .Z(n18374) );
XOR U30625 ( .A(c6125), .B(n18375), .Z(c6126) );
ANDN U30626 ( .B(n18376), .A(n18377), .Z(n18375) );
XOR U30627 ( .A(c6125), .B(b[6125]), .Z(n18376) );
XNOR U30628 ( .A(b[6125]), .B(n18377), .Z(c[6125]) );
XNOR U30629 ( .A(a[6125]), .B(c6125), .Z(n18377) );
XOR U30630 ( .A(c6126), .B(n18378), .Z(c6127) );
ANDN U30631 ( .B(n18379), .A(n18380), .Z(n18378) );
XOR U30632 ( .A(c6126), .B(b[6126]), .Z(n18379) );
XNOR U30633 ( .A(b[6126]), .B(n18380), .Z(c[6126]) );
XNOR U30634 ( .A(a[6126]), .B(c6126), .Z(n18380) );
XOR U30635 ( .A(c6127), .B(n18381), .Z(c6128) );
ANDN U30636 ( .B(n18382), .A(n18383), .Z(n18381) );
XOR U30637 ( .A(c6127), .B(b[6127]), .Z(n18382) );
XNOR U30638 ( .A(b[6127]), .B(n18383), .Z(c[6127]) );
XNOR U30639 ( .A(a[6127]), .B(c6127), .Z(n18383) );
XOR U30640 ( .A(c6128), .B(n18384), .Z(c6129) );
ANDN U30641 ( .B(n18385), .A(n18386), .Z(n18384) );
XOR U30642 ( .A(c6128), .B(b[6128]), .Z(n18385) );
XNOR U30643 ( .A(b[6128]), .B(n18386), .Z(c[6128]) );
XNOR U30644 ( .A(a[6128]), .B(c6128), .Z(n18386) );
XOR U30645 ( .A(c6129), .B(n18387), .Z(c6130) );
ANDN U30646 ( .B(n18388), .A(n18389), .Z(n18387) );
XOR U30647 ( .A(c6129), .B(b[6129]), .Z(n18388) );
XNOR U30648 ( .A(b[6129]), .B(n18389), .Z(c[6129]) );
XNOR U30649 ( .A(a[6129]), .B(c6129), .Z(n18389) );
XOR U30650 ( .A(c6130), .B(n18390), .Z(c6131) );
ANDN U30651 ( .B(n18391), .A(n18392), .Z(n18390) );
XOR U30652 ( .A(c6130), .B(b[6130]), .Z(n18391) );
XNOR U30653 ( .A(b[6130]), .B(n18392), .Z(c[6130]) );
XNOR U30654 ( .A(a[6130]), .B(c6130), .Z(n18392) );
XOR U30655 ( .A(c6131), .B(n18393), .Z(c6132) );
ANDN U30656 ( .B(n18394), .A(n18395), .Z(n18393) );
XOR U30657 ( .A(c6131), .B(b[6131]), .Z(n18394) );
XNOR U30658 ( .A(b[6131]), .B(n18395), .Z(c[6131]) );
XNOR U30659 ( .A(a[6131]), .B(c6131), .Z(n18395) );
XOR U30660 ( .A(c6132), .B(n18396), .Z(c6133) );
ANDN U30661 ( .B(n18397), .A(n18398), .Z(n18396) );
XOR U30662 ( .A(c6132), .B(b[6132]), .Z(n18397) );
XNOR U30663 ( .A(b[6132]), .B(n18398), .Z(c[6132]) );
XNOR U30664 ( .A(a[6132]), .B(c6132), .Z(n18398) );
XOR U30665 ( .A(c6133), .B(n18399), .Z(c6134) );
ANDN U30666 ( .B(n18400), .A(n18401), .Z(n18399) );
XOR U30667 ( .A(c6133), .B(b[6133]), .Z(n18400) );
XNOR U30668 ( .A(b[6133]), .B(n18401), .Z(c[6133]) );
XNOR U30669 ( .A(a[6133]), .B(c6133), .Z(n18401) );
XOR U30670 ( .A(c6134), .B(n18402), .Z(c6135) );
ANDN U30671 ( .B(n18403), .A(n18404), .Z(n18402) );
XOR U30672 ( .A(c6134), .B(b[6134]), .Z(n18403) );
XNOR U30673 ( .A(b[6134]), .B(n18404), .Z(c[6134]) );
XNOR U30674 ( .A(a[6134]), .B(c6134), .Z(n18404) );
XOR U30675 ( .A(c6135), .B(n18405), .Z(c6136) );
ANDN U30676 ( .B(n18406), .A(n18407), .Z(n18405) );
XOR U30677 ( .A(c6135), .B(b[6135]), .Z(n18406) );
XNOR U30678 ( .A(b[6135]), .B(n18407), .Z(c[6135]) );
XNOR U30679 ( .A(a[6135]), .B(c6135), .Z(n18407) );
XOR U30680 ( .A(c6136), .B(n18408), .Z(c6137) );
ANDN U30681 ( .B(n18409), .A(n18410), .Z(n18408) );
XOR U30682 ( .A(c6136), .B(b[6136]), .Z(n18409) );
XNOR U30683 ( .A(b[6136]), .B(n18410), .Z(c[6136]) );
XNOR U30684 ( .A(a[6136]), .B(c6136), .Z(n18410) );
XOR U30685 ( .A(c6137), .B(n18411), .Z(c6138) );
ANDN U30686 ( .B(n18412), .A(n18413), .Z(n18411) );
XOR U30687 ( .A(c6137), .B(b[6137]), .Z(n18412) );
XNOR U30688 ( .A(b[6137]), .B(n18413), .Z(c[6137]) );
XNOR U30689 ( .A(a[6137]), .B(c6137), .Z(n18413) );
XOR U30690 ( .A(c6138), .B(n18414), .Z(c6139) );
ANDN U30691 ( .B(n18415), .A(n18416), .Z(n18414) );
XOR U30692 ( .A(c6138), .B(b[6138]), .Z(n18415) );
XNOR U30693 ( .A(b[6138]), .B(n18416), .Z(c[6138]) );
XNOR U30694 ( .A(a[6138]), .B(c6138), .Z(n18416) );
XOR U30695 ( .A(c6139), .B(n18417), .Z(c6140) );
ANDN U30696 ( .B(n18418), .A(n18419), .Z(n18417) );
XOR U30697 ( .A(c6139), .B(b[6139]), .Z(n18418) );
XNOR U30698 ( .A(b[6139]), .B(n18419), .Z(c[6139]) );
XNOR U30699 ( .A(a[6139]), .B(c6139), .Z(n18419) );
XOR U30700 ( .A(c6140), .B(n18420), .Z(c6141) );
ANDN U30701 ( .B(n18421), .A(n18422), .Z(n18420) );
XOR U30702 ( .A(c6140), .B(b[6140]), .Z(n18421) );
XNOR U30703 ( .A(b[6140]), .B(n18422), .Z(c[6140]) );
XNOR U30704 ( .A(a[6140]), .B(c6140), .Z(n18422) );
XOR U30705 ( .A(c6141), .B(n18423), .Z(c6142) );
ANDN U30706 ( .B(n18424), .A(n18425), .Z(n18423) );
XOR U30707 ( .A(c6141), .B(b[6141]), .Z(n18424) );
XNOR U30708 ( .A(b[6141]), .B(n18425), .Z(c[6141]) );
XNOR U30709 ( .A(a[6141]), .B(c6141), .Z(n18425) );
XOR U30710 ( .A(c6142), .B(n18426), .Z(c6143) );
ANDN U30711 ( .B(n18427), .A(n18428), .Z(n18426) );
XOR U30712 ( .A(c6142), .B(b[6142]), .Z(n18427) );
XNOR U30713 ( .A(b[6142]), .B(n18428), .Z(c[6142]) );
XNOR U30714 ( .A(a[6142]), .B(c6142), .Z(n18428) );
XOR U30715 ( .A(c6143), .B(n18429), .Z(c6144) );
ANDN U30716 ( .B(n18430), .A(n18431), .Z(n18429) );
XOR U30717 ( .A(c6143), .B(b[6143]), .Z(n18430) );
XNOR U30718 ( .A(b[6143]), .B(n18431), .Z(c[6143]) );
XNOR U30719 ( .A(a[6143]), .B(c6143), .Z(n18431) );
XOR U30720 ( .A(c6144), .B(n18432), .Z(c6145) );
ANDN U30721 ( .B(n18433), .A(n18434), .Z(n18432) );
XOR U30722 ( .A(c6144), .B(b[6144]), .Z(n18433) );
XNOR U30723 ( .A(b[6144]), .B(n18434), .Z(c[6144]) );
XNOR U30724 ( .A(a[6144]), .B(c6144), .Z(n18434) );
XOR U30725 ( .A(c6145), .B(n18435), .Z(c6146) );
ANDN U30726 ( .B(n18436), .A(n18437), .Z(n18435) );
XOR U30727 ( .A(c6145), .B(b[6145]), .Z(n18436) );
XNOR U30728 ( .A(b[6145]), .B(n18437), .Z(c[6145]) );
XNOR U30729 ( .A(a[6145]), .B(c6145), .Z(n18437) );
XOR U30730 ( .A(c6146), .B(n18438), .Z(c6147) );
ANDN U30731 ( .B(n18439), .A(n18440), .Z(n18438) );
XOR U30732 ( .A(c6146), .B(b[6146]), .Z(n18439) );
XNOR U30733 ( .A(b[6146]), .B(n18440), .Z(c[6146]) );
XNOR U30734 ( .A(a[6146]), .B(c6146), .Z(n18440) );
XOR U30735 ( .A(c6147), .B(n18441), .Z(c6148) );
ANDN U30736 ( .B(n18442), .A(n18443), .Z(n18441) );
XOR U30737 ( .A(c6147), .B(b[6147]), .Z(n18442) );
XNOR U30738 ( .A(b[6147]), .B(n18443), .Z(c[6147]) );
XNOR U30739 ( .A(a[6147]), .B(c6147), .Z(n18443) );
XOR U30740 ( .A(c6148), .B(n18444), .Z(c6149) );
ANDN U30741 ( .B(n18445), .A(n18446), .Z(n18444) );
XOR U30742 ( .A(c6148), .B(b[6148]), .Z(n18445) );
XNOR U30743 ( .A(b[6148]), .B(n18446), .Z(c[6148]) );
XNOR U30744 ( .A(a[6148]), .B(c6148), .Z(n18446) );
XOR U30745 ( .A(c6149), .B(n18447), .Z(c6150) );
ANDN U30746 ( .B(n18448), .A(n18449), .Z(n18447) );
XOR U30747 ( .A(c6149), .B(b[6149]), .Z(n18448) );
XNOR U30748 ( .A(b[6149]), .B(n18449), .Z(c[6149]) );
XNOR U30749 ( .A(a[6149]), .B(c6149), .Z(n18449) );
XOR U30750 ( .A(c6150), .B(n18450), .Z(c6151) );
ANDN U30751 ( .B(n18451), .A(n18452), .Z(n18450) );
XOR U30752 ( .A(c6150), .B(b[6150]), .Z(n18451) );
XNOR U30753 ( .A(b[6150]), .B(n18452), .Z(c[6150]) );
XNOR U30754 ( .A(a[6150]), .B(c6150), .Z(n18452) );
XOR U30755 ( .A(c6151), .B(n18453), .Z(c6152) );
ANDN U30756 ( .B(n18454), .A(n18455), .Z(n18453) );
XOR U30757 ( .A(c6151), .B(b[6151]), .Z(n18454) );
XNOR U30758 ( .A(b[6151]), .B(n18455), .Z(c[6151]) );
XNOR U30759 ( .A(a[6151]), .B(c6151), .Z(n18455) );
XOR U30760 ( .A(c6152), .B(n18456), .Z(c6153) );
ANDN U30761 ( .B(n18457), .A(n18458), .Z(n18456) );
XOR U30762 ( .A(c6152), .B(b[6152]), .Z(n18457) );
XNOR U30763 ( .A(b[6152]), .B(n18458), .Z(c[6152]) );
XNOR U30764 ( .A(a[6152]), .B(c6152), .Z(n18458) );
XOR U30765 ( .A(c6153), .B(n18459), .Z(c6154) );
ANDN U30766 ( .B(n18460), .A(n18461), .Z(n18459) );
XOR U30767 ( .A(c6153), .B(b[6153]), .Z(n18460) );
XNOR U30768 ( .A(b[6153]), .B(n18461), .Z(c[6153]) );
XNOR U30769 ( .A(a[6153]), .B(c6153), .Z(n18461) );
XOR U30770 ( .A(c6154), .B(n18462), .Z(c6155) );
ANDN U30771 ( .B(n18463), .A(n18464), .Z(n18462) );
XOR U30772 ( .A(c6154), .B(b[6154]), .Z(n18463) );
XNOR U30773 ( .A(b[6154]), .B(n18464), .Z(c[6154]) );
XNOR U30774 ( .A(a[6154]), .B(c6154), .Z(n18464) );
XOR U30775 ( .A(c6155), .B(n18465), .Z(c6156) );
ANDN U30776 ( .B(n18466), .A(n18467), .Z(n18465) );
XOR U30777 ( .A(c6155), .B(b[6155]), .Z(n18466) );
XNOR U30778 ( .A(b[6155]), .B(n18467), .Z(c[6155]) );
XNOR U30779 ( .A(a[6155]), .B(c6155), .Z(n18467) );
XOR U30780 ( .A(c6156), .B(n18468), .Z(c6157) );
ANDN U30781 ( .B(n18469), .A(n18470), .Z(n18468) );
XOR U30782 ( .A(c6156), .B(b[6156]), .Z(n18469) );
XNOR U30783 ( .A(b[6156]), .B(n18470), .Z(c[6156]) );
XNOR U30784 ( .A(a[6156]), .B(c6156), .Z(n18470) );
XOR U30785 ( .A(c6157), .B(n18471), .Z(c6158) );
ANDN U30786 ( .B(n18472), .A(n18473), .Z(n18471) );
XOR U30787 ( .A(c6157), .B(b[6157]), .Z(n18472) );
XNOR U30788 ( .A(b[6157]), .B(n18473), .Z(c[6157]) );
XNOR U30789 ( .A(a[6157]), .B(c6157), .Z(n18473) );
XOR U30790 ( .A(c6158), .B(n18474), .Z(c6159) );
ANDN U30791 ( .B(n18475), .A(n18476), .Z(n18474) );
XOR U30792 ( .A(c6158), .B(b[6158]), .Z(n18475) );
XNOR U30793 ( .A(b[6158]), .B(n18476), .Z(c[6158]) );
XNOR U30794 ( .A(a[6158]), .B(c6158), .Z(n18476) );
XOR U30795 ( .A(c6159), .B(n18477), .Z(c6160) );
ANDN U30796 ( .B(n18478), .A(n18479), .Z(n18477) );
XOR U30797 ( .A(c6159), .B(b[6159]), .Z(n18478) );
XNOR U30798 ( .A(b[6159]), .B(n18479), .Z(c[6159]) );
XNOR U30799 ( .A(a[6159]), .B(c6159), .Z(n18479) );
XOR U30800 ( .A(c6160), .B(n18480), .Z(c6161) );
ANDN U30801 ( .B(n18481), .A(n18482), .Z(n18480) );
XOR U30802 ( .A(c6160), .B(b[6160]), .Z(n18481) );
XNOR U30803 ( .A(b[6160]), .B(n18482), .Z(c[6160]) );
XNOR U30804 ( .A(a[6160]), .B(c6160), .Z(n18482) );
XOR U30805 ( .A(c6161), .B(n18483), .Z(c6162) );
ANDN U30806 ( .B(n18484), .A(n18485), .Z(n18483) );
XOR U30807 ( .A(c6161), .B(b[6161]), .Z(n18484) );
XNOR U30808 ( .A(b[6161]), .B(n18485), .Z(c[6161]) );
XNOR U30809 ( .A(a[6161]), .B(c6161), .Z(n18485) );
XOR U30810 ( .A(c6162), .B(n18486), .Z(c6163) );
ANDN U30811 ( .B(n18487), .A(n18488), .Z(n18486) );
XOR U30812 ( .A(c6162), .B(b[6162]), .Z(n18487) );
XNOR U30813 ( .A(b[6162]), .B(n18488), .Z(c[6162]) );
XNOR U30814 ( .A(a[6162]), .B(c6162), .Z(n18488) );
XOR U30815 ( .A(c6163), .B(n18489), .Z(c6164) );
ANDN U30816 ( .B(n18490), .A(n18491), .Z(n18489) );
XOR U30817 ( .A(c6163), .B(b[6163]), .Z(n18490) );
XNOR U30818 ( .A(b[6163]), .B(n18491), .Z(c[6163]) );
XNOR U30819 ( .A(a[6163]), .B(c6163), .Z(n18491) );
XOR U30820 ( .A(c6164), .B(n18492), .Z(c6165) );
ANDN U30821 ( .B(n18493), .A(n18494), .Z(n18492) );
XOR U30822 ( .A(c6164), .B(b[6164]), .Z(n18493) );
XNOR U30823 ( .A(b[6164]), .B(n18494), .Z(c[6164]) );
XNOR U30824 ( .A(a[6164]), .B(c6164), .Z(n18494) );
XOR U30825 ( .A(c6165), .B(n18495), .Z(c6166) );
ANDN U30826 ( .B(n18496), .A(n18497), .Z(n18495) );
XOR U30827 ( .A(c6165), .B(b[6165]), .Z(n18496) );
XNOR U30828 ( .A(b[6165]), .B(n18497), .Z(c[6165]) );
XNOR U30829 ( .A(a[6165]), .B(c6165), .Z(n18497) );
XOR U30830 ( .A(c6166), .B(n18498), .Z(c6167) );
ANDN U30831 ( .B(n18499), .A(n18500), .Z(n18498) );
XOR U30832 ( .A(c6166), .B(b[6166]), .Z(n18499) );
XNOR U30833 ( .A(b[6166]), .B(n18500), .Z(c[6166]) );
XNOR U30834 ( .A(a[6166]), .B(c6166), .Z(n18500) );
XOR U30835 ( .A(c6167), .B(n18501), .Z(c6168) );
ANDN U30836 ( .B(n18502), .A(n18503), .Z(n18501) );
XOR U30837 ( .A(c6167), .B(b[6167]), .Z(n18502) );
XNOR U30838 ( .A(b[6167]), .B(n18503), .Z(c[6167]) );
XNOR U30839 ( .A(a[6167]), .B(c6167), .Z(n18503) );
XOR U30840 ( .A(c6168), .B(n18504), .Z(c6169) );
ANDN U30841 ( .B(n18505), .A(n18506), .Z(n18504) );
XOR U30842 ( .A(c6168), .B(b[6168]), .Z(n18505) );
XNOR U30843 ( .A(b[6168]), .B(n18506), .Z(c[6168]) );
XNOR U30844 ( .A(a[6168]), .B(c6168), .Z(n18506) );
XOR U30845 ( .A(c6169), .B(n18507), .Z(c6170) );
ANDN U30846 ( .B(n18508), .A(n18509), .Z(n18507) );
XOR U30847 ( .A(c6169), .B(b[6169]), .Z(n18508) );
XNOR U30848 ( .A(b[6169]), .B(n18509), .Z(c[6169]) );
XNOR U30849 ( .A(a[6169]), .B(c6169), .Z(n18509) );
XOR U30850 ( .A(c6170), .B(n18510), .Z(c6171) );
ANDN U30851 ( .B(n18511), .A(n18512), .Z(n18510) );
XOR U30852 ( .A(c6170), .B(b[6170]), .Z(n18511) );
XNOR U30853 ( .A(b[6170]), .B(n18512), .Z(c[6170]) );
XNOR U30854 ( .A(a[6170]), .B(c6170), .Z(n18512) );
XOR U30855 ( .A(c6171), .B(n18513), .Z(c6172) );
ANDN U30856 ( .B(n18514), .A(n18515), .Z(n18513) );
XOR U30857 ( .A(c6171), .B(b[6171]), .Z(n18514) );
XNOR U30858 ( .A(b[6171]), .B(n18515), .Z(c[6171]) );
XNOR U30859 ( .A(a[6171]), .B(c6171), .Z(n18515) );
XOR U30860 ( .A(c6172), .B(n18516), .Z(c6173) );
ANDN U30861 ( .B(n18517), .A(n18518), .Z(n18516) );
XOR U30862 ( .A(c6172), .B(b[6172]), .Z(n18517) );
XNOR U30863 ( .A(b[6172]), .B(n18518), .Z(c[6172]) );
XNOR U30864 ( .A(a[6172]), .B(c6172), .Z(n18518) );
XOR U30865 ( .A(c6173), .B(n18519), .Z(c6174) );
ANDN U30866 ( .B(n18520), .A(n18521), .Z(n18519) );
XOR U30867 ( .A(c6173), .B(b[6173]), .Z(n18520) );
XNOR U30868 ( .A(b[6173]), .B(n18521), .Z(c[6173]) );
XNOR U30869 ( .A(a[6173]), .B(c6173), .Z(n18521) );
XOR U30870 ( .A(c6174), .B(n18522), .Z(c6175) );
ANDN U30871 ( .B(n18523), .A(n18524), .Z(n18522) );
XOR U30872 ( .A(c6174), .B(b[6174]), .Z(n18523) );
XNOR U30873 ( .A(b[6174]), .B(n18524), .Z(c[6174]) );
XNOR U30874 ( .A(a[6174]), .B(c6174), .Z(n18524) );
XOR U30875 ( .A(c6175), .B(n18525), .Z(c6176) );
ANDN U30876 ( .B(n18526), .A(n18527), .Z(n18525) );
XOR U30877 ( .A(c6175), .B(b[6175]), .Z(n18526) );
XNOR U30878 ( .A(b[6175]), .B(n18527), .Z(c[6175]) );
XNOR U30879 ( .A(a[6175]), .B(c6175), .Z(n18527) );
XOR U30880 ( .A(c6176), .B(n18528), .Z(c6177) );
ANDN U30881 ( .B(n18529), .A(n18530), .Z(n18528) );
XOR U30882 ( .A(c6176), .B(b[6176]), .Z(n18529) );
XNOR U30883 ( .A(b[6176]), .B(n18530), .Z(c[6176]) );
XNOR U30884 ( .A(a[6176]), .B(c6176), .Z(n18530) );
XOR U30885 ( .A(c6177), .B(n18531), .Z(c6178) );
ANDN U30886 ( .B(n18532), .A(n18533), .Z(n18531) );
XOR U30887 ( .A(c6177), .B(b[6177]), .Z(n18532) );
XNOR U30888 ( .A(b[6177]), .B(n18533), .Z(c[6177]) );
XNOR U30889 ( .A(a[6177]), .B(c6177), .Z(n18533) );
XOR U30890 ( .A(c6178), .B(n18534), .Z(c6179) );
ANDN U30891 ( .B(n18535), .A(n18536), .Z(n18534) );
XOR U30892 ( .A(c6178), .B(b[6178]), .Z(n18535) );
XNOR U30893 ( .A(b[6178]), .B(n18536), .Z(c[6178]) );
XNOR U30894 ( .A(a[6178]), .B(c6178), .Z(n18536) );
XOR U30895 ( .A(c6179), .B(n18537), .Z(c6180) );
ANDN U30896 ( .B(n18538), .A(n18539), .Z(n18537) );
XOR U30897 ( .A(c6179), .B(b[6179]), .Z(n18538) );
XNOR U30898 ( .A(b[6179]), .B(n18539), .Z(c[6179]) );
XNOR U30899 ( .A(a[6179]), .B(c6179), .Z(n18539) );
XOR U30900 ( .A(c6180), .B(n18540), .Z(c6181) );
ANDN U30901 ( .B(n18541), .A(n18542), .Z(n18540) );
XOR U30902 ( .A(c6180), .B(b[6180]), .Z(n18541) );
XNOR U30903 ( .A(b[6180]), .B(n18542), .Z(c[6180]) );
XNOR U30904 ( .A(a[6180]), .B(c6180), .Z(n18542) );
XOR U30905 ( .A(c6181), .B(n18543), .Z(c6182) );
ANDN U30906 ( .B(n18544), .A(n18545), .Z(n18543) );
XOR U30907 ( .A(c6181), .B(b[6181]), .Z(n18544) );
XNOR U30908 ( .A(b[6181]), .B(n18545), .Z(c[6181]) );
XNOR U30909 ( .A(a[6181]), .B(c6181), .Z(n18545) );
XOR U30910 ( .A(c6182), .B(n18546), .Z(c6183) );
ANDN U30911 ( .B(n18547), .A(n18548), .Z(n18546) );
XOR U30912 ( .A(c6182), .B(b[6182]), .Z(n18547) );
XNOR U30913 ( .A(b[6182]), .B(n18548), .Z(c[6182]) );
XNOR U30914 ( .A(a[6182]), .B(c6182), .Z(n18548) );
XOR U30915 ( .A(c6183), .B(n18549), .Z(c6184) );
ANDN U30916 ( .B(n18550), .A(n18551), .Z(n18549) );
XOR U30917 ( .A(c6183), .B(b[6183]), .Z(n18550) );
XNOR U30918 ( .A(b[6183]), .B(n18551), .Z(c[6183]) );
XNOR U30919 ( .A(a[6183]), .B(c6183), .Z(n18551) );
XOR U30920 ( .A(c6184), .B(n18552), .Z(c6185) );
ANDN U30921 ( .B(n18553), .A(n18554), .Z(n18552) );
XOR U30922 ( .A(c6184), .B(b[6184]), .Z(n18553) );
XNOR U30923 ( .A(b[6184]), .B(n18554), .Z(c[6184]) );
XNOR U30924 ( .A(a[6184]), .B(c6184), .Z(n18554) );
XOR U30925 ( .A(c6185), .B(n18555), .Z(c6186) );
ANDN U30926 ( .B(n18556), .A(n18557), .Z(n18555) );
XOR U30927 ( .A(c6185), .B(b[6185]), .Z(n18556) );
XNOR U30928 ( .A(b[6185]), .B(n18557), .Z(c[6185]) );
XNOR U30929 ( .A(a[6185]), .B(c6185), .Z(n18557) );
XOR U30930 ( .A(c6186), .B(n18558), .Z(c6187) );
ANDN U30931 ( .B(n18559), .A(n18560), .Z(n18558) );
XOR U30932 ( .A(c6186), .B(b[6186]), .Z(n18559) );
XNOR U30933 ( .A(b[6186]), .B(n18560), .Z(c[6186]) );
XNOR U30934 ( .A(a[6186]), .B(c6186), .Z(n18560) );
XOR U30935 ( .A(c6187), .B(n18561), .Z(c6188) );
ANDN U30936 ( .B(n18562), .A(n18563), .Z(n18561) );
XOR U30937 ( .A(c6187), .B(b[6187]), .Z(n18562) );
XNOR U30938 ( .A(b[6187]), .B(n18563), .Z(c[6187]) );
XNOR U30939 ( .A(a[6187]), .B(c6187), .Z(n18563) );
XOR U30940 ( .A(c6188), .B(n18564), .Z(c6189) );
ANDN U30941 ( .B(n18565), .A(n18566), .Z(n18564) );
XOR U30942 ( .A(c6188), .B(b[6188]), .Z(n18565) );
XNOR U30943 ( .A(b[6188]), .B(n18566), .Z(c[6188]) );
XNOR U30944 ( .A(a[6188]), .B(c6188), .Z(n18566) );
XOR U30945 ( .A(c6189), .B(n18567), .Z(c6190) );
ANDN U30946 ( .B(n18568), .A(n18569), .Z(n18567) );
XOR U30947 ( .A(c6189), .B(b[6189]), .Z(n18568) );
XNOR U30948 ( .A(b[6189]), .B(n18569), .Z(c[6189]) );
XNOR U30949 ( .A(a[6189]), .B(c6189), .Z(n18569) );
XOR U30950 ( .A(c6190), .B(n18570), .Z(c6191) );
ANDN U30951 ( .B(n18571), .A(n18572), .Z(n18570) );
XOR U30952 ( .A(c6190), .B(b[6190]), .Z(n18571) );
XNOR U30953 ( .A(b[6190]), .B(n18572), .Z(c[6190]) );
XNOR U30954 ( .A(a[6190]), .B(c6190), .Z(n18572) );
XOR U30955 ( .A(c6191), .B(n18573), .Z(c6192) );
ANDN U30956 ( .B(n18574), .A(n18575), .Z(n18573) );
XOR U30957 ( .A(c6191), .B(b[6191]), .Z(n18574) );
XNOR U30958 ( .A(b[6191]), .B(n18575), .Z(c[6191]) );
XNOR U30959 ( .A(a[6191]), .B(c6191), .Z(n18575) );
XOR U30960 ( .A(c6192), .B(n18576), .Z(c6193) );
ANDN U30961 ( .B(n18577), .A(n18578), .Z(n18576) );
XOR U30962 ( .A(c6192), .B(b[6192]), .Z(n18577) );
XNOR U30963 ( .A(b[6192]), .B(n18578), .Z(c[6192]) );
XNOR U30964 ( .A(a[6192]), .B(c6192), .Z(n18578) );
XOR U30965 ( .A(c6193), .B(n18579), .Z(c6194) );
ANDN U30966 ( .B(n18580), .A(n18581), .Z(n18579) );
XOR U30967 ( .A(c6193), .B(b[6193]), .Z(n18580) );
XNOR U30968 ( .A(b[6193]), .B(n18581), .Z(c[6193]) );
XNOR U30969 ( .A(a[6193]), .B(c6193), .Z(n18581) );
XOR U30970 ( .A(c6194), .B(n18582), .Z(c6195) );
ANDN U30971 ( .B(n18583), .A(n18584), .Z(n18582) );
XOR U30972 ( .A(c6194), .B(b[6194]), .Z(n18583) );
XNOR U30973 ( .A(b[6194]), .B(n18584), .Z(c[6194]) );
XNOR U30974 ( .A(a[6194]), .B(c6194), .Z(n18584) );
XOR U30975 ( .A(c6195), .B(n18585), .Z(c6196) );
ANDN U30976 ( .B(n18586), .A(n18587), .Z(n18585) );
XOR U30977 ( .A(c6195), .B(b[6195]), .Z(n18586) );
XNOR U30978 ( .A(b[6195]), .B(n18587), .Z(c[6195]) );
XNOR U30979 ( .A(a[6195]), .B(c6195), .Z(n18587) );
XOR U30980 ( .A(c6196), .B(n18588), .Z(c6197) );
ANDN U30981 ( .B(n18589), .A(n18590), .Z(n18588) );
XOR U30982 ( .A(c6196), .B(b[6196]), .Z(n18589) );
XNOR U30983 ( .A(b[6196]), .B(n18590), .Z(c[6196]) );
XNOR U30984 ( .A(a[6196]), .B(c6196), .Z(n18590) );
XOR U30985 ( .A(c6197), .B(n18591), .Z(c6198) );
ANDN U30986 ( .B(n18592), .A(n18593), .Z(n18591) );
XOR U30987 ( .A(c6197), .B(b[6197]), .Z(n18592) );
XNOR U30988 ( .A(b[6197]), .B(n18593), .Z(c[6197]) );
XNOR U30989 ( .A(a[6197]), .B(c6197), .Z(n18593) );
XOR U30990 ( .A(c6198), .B(n18594), .Z(c6199) );
ANDN U30991 ( .B(n18595), .A(n18596), .Z(n18594) );
XOR U30992 ( .A(c6198), .B(b[6198]), .Z(n18595) );
XNOR U30993 ( .A(b[6198]), .B(n18596), .Z(c[6198]) );
XNOR U30994 ( .A(a[6198]), .B(c6198), .Z(n18596) );
XOR U30995 ( .A(c6199), .B(n18597), .Z(c6200) );
ANDN U30996 ( .B(n18598), .A(n18599), .Z(n18597) );
XOR U30997 ( .A(c6199), .B(b[6199]), .Z(n18598) );
XNOR U30998 ( .A(b[6199]), .B(n18599), .Z(c[6199]) );
XNOR U30999 ( .A(a[6199]), .B(c6199), .Z(n18599) );
XOR U31000 ( .A(c6200), .B(n18600), .Z(c6201) );
ANDN U31001 ( .B(n18601), .A(n18602), .Z(n18600) );
XOR U31002 ( .A(c6200), .B(b[6200]), .Z(n18601) );
XNOR U31003 ( .A(b[6200]), .B(n18602), .Z(c[6200]) );
XNOR U31004 ( .A(a[6200]), .B(c6200), .Z(n18602) );
XOR U31005 ( .A(c6201), .B(n18603), .Z(c6202) );
ANDN U31006 ( .B(n18604), .A(n18605), .Z(n18603) );
XOR U31007 ( .A(c6201), .B(b[6201]), .Z(n18604) );
XNOR U31008 ( .A(b[6201]), .B(n18605), .Z(c[6201]) );
XNOR U31009 ( .A(a[6201]), .B(c6201), .Z(n18605) );
XOR U31010 ( .A(c6202), .B(n18606), .Z(c6203) );
ANDN U31011 ( .B(n18607), .A(n18608), .Z(n18606) );
XOR U31012 ( .A(c6202), .B(b[6202]), .Z(n18607) );
XNOR U31013 ( .A(b[6202]), .B(n18608), .Z(c[6202]) );
XNOR U31014 ( .A(a[6202]), .B(c6202), .Z(n18608) );
XOR U31015 ( .A(c6203), .B(n18609), .Z(c6204) );
ANDN U31016 ( .B(n18610), .A(n18611), .Z(n18609) );
XOR U31017 ( .A(c6203), .B(b[6203]), .Z(n18610) );
XNOR U31018 ( .A(b[6203]), .B(n18611), .Z(c[6203]) );
XNOR U31019 ( .A(a[6203]), .B(c6203), .Z(n18611) );
XOR U31020 ( .A(c6204), .B(n18612), .Z(c6205) );
ANDN U31021 ( .B(n18613), .A(n18614), .Z(n18612) );
XOR U31022 ( .A(c6204), .B(b[6204]), .Z(n18613) );
XNOR U31023 ( .A(b[6204]), .B(n18614), .Z(c[6204]) );
XNOR U31024 ( .A(a[6204]), .B(c6204), .Z(n18614) );
XOR U31025 ( .A(c6205), .B(n18615), .Z(c6206) );
ANDN U31026 ( .B(n18616), .A(n18617), .Z(n18615) );
XOR U31027 ( .A(c6205), .B(b[6205]), .Z(n18616) );
XNOR U31028 ( .A(b[6205]), .B(n18617), .Z(c[6205]) );
XNOR U31029 ( .A(a[6205]), .B(c6205), .Z(n18617) );
XOR U31030 ( .A(c6206), .B(n18618), .Z(c6207) );
ANDN U31031 ( .B(n18619), .A(n18620), .Z(n18618) );
XOR U31032 ( .A(c6206), .B(b[6206]), .Z(n18619) );
XNOR U31033 ( .A(b[6206]), .B(n18620), .Z(c[6206]) );
XNOR U31034 ( .A(a[6206]), .B(c6206), .Z(n18620) );
XOR U31035 ( .A(c6207), .B(n18621), .Z(c6208) );
ANDN U31036 ( .B(n18622), .A(n18623), .Z(n18621) );
XOR U31037 ( .A(c6207), .B(b[6207]), .Z(n18622) );
XNOR U31038 ( .A(b[6207]), .B(n18623), .Z(c[6207]) );
XNOR U31039 ( .A(a[6207]), .B(c6207), .Z(n18623) );
XOR U31040 ( .A(c6208), .B(n18624), .Z(c6209) );
ANDN U31041 ( .B(n18625), .A(n18626), .Z(n18624) );
XOR U31042 ( .A(c6208), .B(b[6208]), .Z(n18625) );
XNOR U31043 ( .A(b[6208]), .B(n18626), .Z(c[6208]) );
XNOR U31044 ( .A(a[6208]), .B(c6208), .Z(n18626) );
XOR U31045 ( .A(c6209), .B(n18627), .Z(c6210) );
ANDN U31046 ( .B(n18628), .A(n18629), .Z(n18627) );
XOR U31047 ( .A(c6209), .B(b[6209]), .Z(n18628) );
XNOR U31048 ( .A(b[6209]), .B(n18629), .Z(c[6209]) );
XNOR U31049 ( .A(a[6209]), .B(c6209), .Z(n18629) );
XOR U31050 ( .A(c6210), .B(n18630), .Z(c6211) );
ANDN U31051 ( .B(n18631), .A(n18632), .Z(n18630) );
XOR U31052 ( .A(c6210), .B(b[6210]), .Z(n18631) );
XNOR U31053 ( .A(b[6210]), .B(n18632), .Z(c[6210]) );
XNOR U31054 ( .A(a[6210]), .B(c6210), .Z(n18632) );
XOR U31055 ( .A(c6211), .B(n18633), .Z(c6212) );
ANDN U31056 ( .B(n18634), .A(n18635), .Z(n18633) );
XOR U31057 ( .A(c6211), .B(b[6211]), .Z(n18634) );
XNOR U31058 ( .A(b[6211]), .B(n18635), .Z(c[6211]) );
XNOR U31059 ( .A(a[6211]), .B(c6211), .Z(n18635) );
XOR U31060 ( .A(c6212), .B(n18636), .Z(c6213) );
ANDN U31061 ( .B(n18637), .A(n18638), .Z(n18636) );
XOR U31062 ( .A(c6212), .B(b[6212]), .Z(n18637) );
XNOR U31063 ( .A(b[6212]), .B(n18638), .Z(c[6212]) );
XNOR U31064 ( .A(a[6212]), .B(c6212), .Z(n18638) );
XOR U31065 ( .A(c6213), .B(n18639), .Z(c6214) );
ANDN U31066 ( .B(n18640), .A(n18641), .Z(n18639) );
XOR U31067 ( .A(c6213), .B(b[6213]), .Z(n18640) );
XNOR U31068 ( .A(b[6213]), .B(n18641), .Z(c[6213]) );
XNOR U31069 ( .A(a[6213]), .B(c6213), .Z(n18641) );
XOR U31070 ( .A(c6214), .B(n18642), .Z(c6215) );
ANDN U31071 ( .B(n18643), .A(n18644), .Z(n18642) );
XOR U31072 ( .A(c6214), .B(b[6214]), .Z(n18643) );
XNOR U31073 ( .A(b[6214]), .B(n18644), .Z(c[6214]) );
XNOR U31074 ( .A(a[6214]), .B(c6214), .Z(n18644) );
XOR U31075 ( .A(c6215), .B(n18645), .Z(c6216) );
ANDN U31076 ( .B(n18646), .A(n18647), .Z(n18645) );
XOR U31077 ( .A(c6215), .B(b[6215]), .Z(n18646) );
XNOR U31078 ( .A(b[6215]), .B(n18647), .Z(c[6215]) );
XNOR U31079 ( .A(a[6215]), .B(c6215), .Z(n18647) );
XOR U31080 ( .A(c6216), .B(n18648), .Z(c6217) );
ANDN U31081 ( .B(n18649), .A(n18650), .Z(n18648) );
XOR U31082 ( .A(c6216), .B(b[6216]), .Z(n18649) );
XNOR U31083 ( .A(b[6216]), .B(n18650), .Z(c[6216]) );
XNOR U31084 ( .A(a[6216]), .B(c6216), .Z(n18650) );
XOR U31085 ( .A(c6217), .B(n18651), .Z(c6218) );
ANDN U31086 ( .B(n18652), .A(n18653), .Z(n18651) );
XOR U31087 ( .A(c6217), .B(b[6217]), .Z(n18652) );
XNOR U31088 ( .A(b[6217]), .B(n18653), .Z(c[6217]) );
XNOR U31089 ( .A(a[6217]), .B(c6217), .Z(n18653) );
XOR U31090 ( .A(c6218), .B(n18654), .Z(c6219) );
ANDN U31091 ( .B(n18655), .A(n18656), .Z(n18654) );
XOR U31092 ( .A(c6218), .B(b[6218]), .Z(n18655) );
XNOR U31093 ( .A(b[6218]), .B(n18656), .Z(c[6218]) );
XNOR U31094 ( .A(a[6218]), .B(c6218), .Z(n18656) );
XOR U31095 ( .A(c6219), .B(n18657), .Z(c6220) );
ANDN U31096 ( .B(n18658), .A(n18659), .Z(n18657) );
XOR U31097 ( .A(c6219), .B(b[6219]), .Z(n18658) );
XNOR U31098 ( .A(b[6219]), .B(n18659), .Z(c[6219]) );
XNOR U31099 ( .A(a[6219]), .B(c6219), .Z(n18659) );
XOR U31100 ( .A(c6220), .B(n18660), .Z(c6221) );
ANDN U31101 ( .B(n18661), .A(n18662), .Z(n18660) );
XOR U31102 ( .A(c6220), .B(b[6220]), .Z(n18661) );
XNOR U31103 ( .A(b[6220]), .B(n18662), .Z(c[6220]) );
XNOR U31104 ( .A(a[6220]), .B(c6220), .Z(n18662) );
XOR U31105 ( .A(c6221), .B(n18663), .Z(c6222) );
ANDN U31106 ( .B(n18664), .A(n18665), .Z(n18663) );
XOR U31107 ( .A(c6221), .B(b[6221]), .Z(n18664) );
XNOR U31108 ( .A(b[6221]), .B(n18665), .Z(c[6221]) );
XNOR U31109 ( .A(a[6221]), .B(c6221), .Z(n18665) );
XOR U31110 ( .A(c6222), .B(n18666), .Z(c6223) );
ANDN U31111 ( .B(n18667), .A(n18668), .Z(n18666) );
XOR U31112 ( .A(c6222), .B(b[6222]), .Z(n18667) );
XNOR U31113 ( .A(b[6222]), .B(n18668), .Z(c[6222]) );
XNOR U31114 ( .A(a[6222]), .B(c6222), .Z(n18668) );
XOR U31115 ( .A(c6223), .B(n18669), .Z(c6224) );
ANDN U31116 ( .B(n18670), .A(n18671), .Z(n18669) );
XOR U31117 ( .A(c6223), .B(b[6223]), .Z(n18670) );
XNOR U31118 ( .A(b[6223]), .B(n18671), .Z(c[6223]) );
XNOR U31119 ( .A(a[6223]), .B(c6223), .Z(n18671) );
XOR U31120 ( .A(c6224), .B(n18672), .Z(c6225) );
ANDN U31121 ( .B(n18673), .A(n18674), .Z(n18672) );
XOR U31122 ( .A(c6224), .B(b[6224]), .Z(n18673) );
XNOR U31123 ( .A(b[6224]), .B(n18674), .Z(c[6224]) );
XNOR U31124 ( .A(a[6224]), .B(c6224), .Z(n18674) );
XOR U31125 ( .A(c6225), .B(n18675), .Z(c6226) );
ANDN U31126 ( .B(n18676), .A(n18677), .Z(n18675) );
XOR U31127 ( .A(c6225), .B(b[6225]), .Z(n18676) );
XNOR U31128 ( .A(b[6225]), .B(n18677), .Z(c[6225]) );
XNOR U31129 ( .A(a[6225]), .B(c6225), .Z(n18677) );
XOR U31130 ( .A(c6226), .B(n18678), .Z(c6227) );
ANDN U31131 ( .B(n18679), .A(n18680), .Z(n18678) );
XOR U31132 ( .A(c6226), .B(b[6226]), .Z(n18679) );
XNOR U31133 ( .A(b[6226]), .B(n18680), .Z(c[6226]) );
XNOR U31134 ( .A(a[6226]), .B(c6226), .Z(n18680) );
XOR U31135 ( .A(c6227), .B(n18681), .Z(c6228) );
ANDN U31136 ( .B(n18682), .A(n18683), .Z(n18681) );
XOR U31137 ( .A(c6227), .B(b[6227]), .Z(n18682) );
XNOR U31138 ( .A(b[6227]), .B(n18683), .Z(c[6227]) );
XNOR U31139 ( .A(a[6227]), .B(c6227), .Z(n18683) );
XOR U31140 ( .A(c6228), .B(n18684), .Z(c6229) );
ANDN U31141 ( .B(n18685), .A(n18686), .Z(n18684) );
XOR U31142 ( .A(c6228), .B(b[6228]), .Z(n18685) );
XNOR U31143 ( .A(b[6228]), .B(n18686), .Z(c[6228]) );
XNOR U31144 ( .A(a[6228]), .B(c6228), .Z(n18686) );
XOR U31145 ( .A(c6229), .B(n18687), .Z(c6230) );
ANDN U31146 ( .B(n18688), .A(n18689), .Z(n18687) );
XOR U31147 ( .A(c6229), .B(b[6229]), .Z(n18688) );
XNOR U31148 ( .A(b[6229]), .B(n18689), .Z(c[6229]) );
XNOR U31149 ( .A(a[6229]), .B(c6229), .Z(n18689) );
XOR U31150 ( .A(c6230), .B(n18690), .Z(c6231) );
ANDN U31151 ( .B(n18691), .A(n18692), .Z(n18690) );
XOR U31152 ( .A(c6230), .B(b[6230]), .Z(n18691) );
XNOR U31153 ( .A(b[6230]), .B(n18692), .Z(c[6230]) );
XNOR U31154 ( .A(a[6230]), .B(c6230), .Z(n18692) );
XOR U31155 ( .A(c6231), .B(n18693), .Z(c6232) );
ANDN U31156 ( .B(n18694), .A(n18695), .Z(n18693) );
XOR U31157 ( .A(c6231), .B(b[6231]), .Z(n18694) );
XNOR U31158 ( .A(b[6231]), .B(n18695), .Z(c[6231]) );
XNOR U31159 ( .A(a[6231]), .B(c6231), .Z(n18695) );
XOR U31160 ( .A(c6232), .B(n18696), .Z(c6233) );
ANDN U31161 ( .B(n18697), .A(n18698), .Z(n18696) );
XOR U31162 ( .A(c6232), .B(b[6232]), .Z(n18697) );
XNOR U31163 ( .A(b[6232]), .B(n18698), .Z(c[6232]) );
XNOR U31164 ( .A(a[6232]), .B(c6232), .Z(n18698) );
XOR U31165 ( .A(c6233), .B(n18699), .Z(c6234) );
ANDN U31166 ( .B(n18700), .A(n18701), .Z(n18699) );
XOR U31167 ( .A(c6233), .B(b[6233]), .Z(n18700) );
XNOR U31168 ( .A(b[6233]), .B(n18701), .Z(c[6233]) );
XNOR U31169 ( .A(a[6233]), .B(c6233), .Z(n18701) );
XOR U31170 ( .A(c6234), .B(n18702), .Z(c6235) );
ANDN U31171 ( .B(n18703), .A(n18704), .Z(n18702) );
XOR U31172 ( .A(c6234), .B(b[6234]), .Z(n18703) );
XNOR U31173 ( .A(b[6234]), .B(n18704), .Z(c[6234]) );
XNOR U31174 ( .A(a[6234]), .B(c6234), .Z(n18704) );
XOR U31175 ( .A(c6235), .B(n18705), .Z(c6236) );
ANDN U31176 ( .B(n18706), .A(n18707), .Z(n18705) );
XOR U31177 ( .A(c6235), .B(b[6235]), .Z(n18706) );
XNOR U31178 ( .A(b[6235]), .B(n18707), .Z(c[6235]) );
XNOR U31179 ( .A(a[6235]), .B(c6235), .Z(n18707) );
XOR U31180 ( .A(c6236), .B(n18708), .Z(c6237) );
ANDN U31181 ( .B(n18709), .A(n18710), .Z(n18708) );
XOR U31182 ( .A(c6236), .B(b[6236]), .Z(n18709) );
XNOR U31183 ( .A(b[6236]), .B(n18710), .Z(c[6236]) );
XNOR U31184 ( .A(a[6236]), .B(c6236), .Z(n18710) );
XOR U31185 ( .A(c6237), .B(n18711), .Z(c6238) );
ANDN U31186 ( .B(n18712), .A(n18713), .Z(n18711) );
XOR U31187 ( .A(c6237), .B(b[6237]), .Z(n18712) );
XNOR U31188 ( .A(b[6237]), .B(n18713), .Z(c[6237]) );
XNOR U31189 ( .A(a[6237]), .B(c6237), .Z(n18713) );
XOR U31190 ( .A(c6238), .B(n18714), .Z(c6239) );
ANDN U31191 ( .B(n18715), .A(n18716), .Z(n18714) );
XOR U31192 ( .A(c6238), .B(b[6238]), .Z(n18715) );
XNOR U31193 ( .A(b[6238]), .B(n18716), .Z(c[6238]) );
XNOR U31194 ( .A(a[6238]), .B(c6238), .Z(n18716) );
XOR U31195 ( .A(c6239), .B(n18717), .Z(c6240) );
ANDN U31196 ( .B(n18718), .A(n18719), .Z(n18717) );
XOR U31197 ( .A(c6239), .B(b[6239]), .Z(n18718) );
XNOR U31198 ( .A(b[6239]), .B(n18719), .Z(c[6239]) );
XNOR U31199 ( .A(a[6239]), .B(c6239), .Z(n18719) );
XOR U31200 ( .A(c6240), .B(n18720), .Z(c6241) );
ANDN U31201 ( .B(n18721), .A(n18722), .Z(n18720) );
XOR U31202 ( .A(c6240), .B(b[6240]), .Z(n18721) );
XNOR U31203 ( .A(b[6240]), .B(n18722), .Z(c[6240]) );
XNOR U31204 ( .A(a[6240]), .B(c6240), .Z(n18722) );
XOR U31205 ( .A(c6241), .B(n18723), .Z(c6242) );
ANDN U31206 ( .B(n18724), .A(n18725), .Z(n18723) );
XOR U31207 ( .A(c6241), .B(b[6241]), .Z(n18724) );
XNOR U31208 ( .A(b[6241]), .B(n18725), .Z(c[6241]) );
XNOR U31209 ( .A(a[6241]), .B(c6241), .Z(n18725) );
XOR U31210 ( .A(c6242), .B(n18726), .Z(c6243) );
ANDN U31211 ( .B(n18727), .A(n18728), .Z(n18726) );
XOR U31212 ( .A(c6242), .B(b[6242]), .Z(n18727) );
XNOR U31213 ( .A(b[6242]), .B(n18728), .Z(c[6242]) );
XNOR U31214 ( .A(a[6242]), .B(c6242), .Z(n18728) );
XOR U31215 ( .A(c6243), .B(n18729), .Z(c6244) );
ANDN U31216 ( .B(n18730), .A(n18731), .Z(n18729) );
XOR U31217 ( .A(c6243), .B(b[6243]), .Z(n18730) );
XNOR U31218 ( .A(b[6243]), .B(n18731), .Z(c[6243]) );
XNOR U31219 ( .A(a[6243]), .B(c6243), .Z(n18731) );
XOR U31220 ( .A(c6244), .B(n18732), .Z(c6245) );
ANDN U31221 ( .B(n18733), .A(n18734), .Z(n18732) );
XOR U31222 ( .A(c6244), .B(b[6244]), .Z(n18733) );
XNOR U31223 ( .A(b[6244]), .B(n18734), .Z(c[6244]) );
XNOR U31224 ( .A(a[6244]), .B(c6244), .Z(n18734) );
XOR U31225 ( .A(c6245), .B(n18735), .Z(c6246) );
ANDN U31226 ( .B(n18736), .A(n18737), .Z(n18735) );
XOR U31227 ( .A(c6245), .B(b[6245]), .Z(n18736) );
XNOR U31228 ( .A(b[6245]), .B(n18737), .Z(c[6245]) );
XNOR U31229 ( .A(a[6245]), .B(c6245), .Z(n18737) );
XOR U31230 ( .A(c6246), .B(n18738), .Z(c6247) );
ANDN U31231 ( .B(n18739), .A(n18740), .Z(n18738) );
XOR U31232 ( .A(c6246), .B(b[6246]), .Z(n18739) );
XNOR U31233 ( .A(b[6246]), .B(n18740), .Z(c[6246]) );
XNOR U31234 ( .A(a[6246]), .B(c6246), .Z(n18740) );
XOR U31235 ( .A(c6247), .B(n18741), .Z(c6248) );
ANDN U31236 ( .B(n18742), .A(n18743), .Z(n18741) );
XOR U31237 ( .A(c6247), .B(b[6247]), .Z(n18742) );
XNOR U31238 ( .A(b[6247]), .B(n18743), .Z(c[6247]) );
XNOR U31239 ( .A(a[6247]), .B(c6247), .Z(n18743) );
XOR U31240 ( .A(c6248), .B(n18744), .Z(c6249) );
ANDN U31241 ( .B(n18745), .A(n18746), .Z(n18744) );
XOR U31242 ( .A(c6248), .B(b[6248]), .Z(n18745) );
XNOR U31243 ( .A(b[6248]), .B(n18746), .Z(c[6248]) );
XNOR U31244 ( .A(a[6248]), .B(c6248), .Z(n18746) );
XOR U31245 ( .A(c6249), .B(n18747), .Z(c6250) );
ANDN U31246 ( .B(n18748), .A(n18749), .Z(n18747) );
XOR U31247 ( .A(c6249), .B(b[6249]), .Z(n18748) );
XNOR U31248 ( .A(b[6249]), .B(n18749), .Z(c[6249]) );
XNOR U31249 ( .A(a[6249]), .B(c6249), .Z(n18749) );
XOR U31250 ( .A(c6250), .B(n18750), .Z(c6251) );
ANDN U31251 ( .B(n18751), .A(n18752), .Z(n18750) );
XOR U31252 ( .A(c6250), .B(b[6250]), .Z(n18751) );
XNOR U31253 ( .A(b[6250]), .B(n18752), .Z(c[6250]) );
XNOR U31254 ( .A(a[6250]), .B(c6250), .Z(n18752) );
XOR U31255 ( .A(c6251), .B(n18753), .Z(c6252) );
ANDN U31256 ( .B(n18754), .A(n18755), .Z(n18753) );
XOR U31257 ( .A(c6251), .B(b[6251]), .Z(n18754) );
XNOR U31258 ( .A(b[6251]), .B(n18755), .Z(c[6251]) );
XNOR U31259 ( .A(a[6251]), .B(c6251), .Z(n18755) );
XOR U31260 ( .A(c6252), .B(n18756), .Z(c6253) );
ANDN U31261 ( .B(n18757), .A(n18758), .Z(n18756) );
XOR U31262 ( .A(c6252), .B(b[6252]), .Z(n18757) );
XNOR U31263 ( .A(b[6252]), .B(n18758), .Z(c[6252]) );
XNOR U31264 ( .A(a[6252]), .B(c6252), .Z(n18758) );
XOR U31265 ( .A(c6253), .B(n18759), .Z(c6254) );
ANDN U31266 ( .B(n18760), .A(n18761), .Z(n18759) );
XOR U31267 ( .A(c6253), .B(b[6253]), .Z(n18760) );
XNOR U31268 ( .A(b[6253]), .B(n18761), .Z(c[6253]) );
XNOR U31269 ( .A(a[6253]), .B(c6253), .Z(n18761) );
XOR U31270 ( .A(c6254), .B(n18762), .Z(c6255) );
ANDN U31271 ( .B(n18763), .A(n18764), .Z(n18762) );
XOR U31272 ( .A(c6254), .B(b[6254]), .Z(n18763) );
XNOR U31273 ( .A(b[6254]), .B(n18764), .Z(c[6254]) );
XNOR U31274 ( .A(a[6254]), .B(c6254), .Z(n18764) );
XOR U31275 ( .A(c6255), .B(n18765), .Z(c6256) );
ANDN U31276 ( .B(n18766), .A(n18767), .Z(n18765) );
XOR U31277 ( .A(c6255), .B(b[6255]), .Z(n18766) );
XNOR U31278 ( .A(b[6255]), .B(n18767), .Z(c[6255]) );
XNOR U31279 ( .A(a[6255]), .B(c6255), .Z(n18767) );
XOR U31280 ( .A(c6256), .B(n18768), .Z(c6257) );
ANDN U31281 ( .B(n18769), .A(n18770), .Z(n18768) );
XOR U31282 ( .A(c6256), .B(b[6256]), .Z(n18769) );
XNOR U31283 ( .A(b[6256]), .B(n18770), .Z(c[6256]) );
XNOR U31284 ( .A(a[6256]), .B(c6256), .Z(n18770) );
XOR U31285 ( .A(c6257), .B(n18771), .Z(c6258) );
ANDN U31286 ( .B(n18772), .A(n18773), .Z(n18771) );
XOR U31287 ( .A(c6257), .B(b[6257]), .Z(n18772) );
XNOR U31288 ( .A(b[6257]), .B(n18773), .Z(c[6257]) );
XNOR U31289 ( .A(a[6257]), .B(c6257), .Z(n18773) );
XOR U31290 ( .A(c6258), .B(n18774), .Z(c6259) );
ANDN U31291 ( .B(n18775), .A(n18776), .Z(n18774) );
XOR U31292 ( .A(c6258), .B(b[6258]), .Z(n18775) );
XNOR U31293 ( .A(b[6258]), .B(n18776), .Z(c[6258]) );
XNOR U31294 ( .A(a[6258]), .B(c6258), .Z(n18776) );
XOR U31295 ( .A(c6259), .B(n18777), .Z(c6260) );
ANDN U31296 ( .B(n18778), .A(n18779), .Z(n18777) );
XOR U31297 ( .A(c6259), .B(b[6259]), .Z(n18778) );
XNOR U31298 ( .A(b[6259]), .B(n18779), .Z(c[6259]) );
XNOR U31299 ( .A(a[6259]), .B(c6259), .Z(n18779) );
XOR U31300 ( .A(c6260), .B(n18780), .Z(c6261) );
ANDN U31301 ( .B(n18781), .A(n18782), .Z(n18780) );
XOR U31302 ( .A(c6260), .B(b[6260]), .Z(n18781) );
XNOR U31303 ( .A(b[6260]), .B(n18782), .Z(c[6260]) );
XNOR U31304 ( .A(a[6260]), .B(c6260), .Z(n18782) );
XOR U31305 ( .A(c6261), .B(n18783), .Z(c6262) );
ANDN U31306 ( .B(n18784), .A(n18785), .Z(n18783) );
XOR U31307 ( .A(c6261), .B(b[6261]), .Z(n18784) );
XNOR U31308 ( .A(b[6261]), .B(n18785), .Z(c[6261]) );
XNOR U31309 ( .A(a[6261]), .B(c6261), .Z(n18785) );
XOR U31310 ( .A(c6262), .B(n18786), .Z(c6263) );
ANDN U31311 ( .B(n18787), .A(n18788), .Z(n18786) );
XOR U31312 ( .A(c6262), .B(b[6262]), .Z(n18787) );
XNOR U31313 ( .A(b[6262]), .B(n18788), .Z(c[6262]) );
XNOR U31314 ( .A(a[6262]), .B(c6262), .Z(n18788) );
XOR U31315 ( .A(c6263), .B(n18789), .Z(c6264) );
ANDN U31316 ( .B(n18790), .A(n18791), .Z(n18789) );
XOR U31317 ( .A(c6263), .B(b[6263]), .Z(n18790) );
XNOR U31318 ( .A(b[6263]), .B(n18791), .Z(c[6263]) );
XNOR U31319 ( .A(a[6263]), .B(c6263), .Z(n18791) );
XOR U31320 ( .A(c6264), .B(n18792), .Z(c6265) );
ANDN U31321 ( .B(n18793), .A(n18794), .Z(n18792) );
XOR U31322 ( .A(c6264), .B(b[6264]), .Z(n18793) );
XNOR U31323 ( .A(b[6264]), .B(n18794), .Z(c[6264]) );
XNOR U31324 ( .A(a[6264]), .B(c6264), .Z(n18794) );
XOR U31325 ( .A(c6265), .B(n18795), .Z(c6266) );
ANDN U31326 ( .B(n18796), .A(n18797), .Z(n18795) );
XOR U31327 ( .A(c6265), .B(b[6265]), .Z(n18796) );
XNOR U31328 ( .A(b[6265]), .B(n18797), .Z(c[6265]) );
XNOR U31329 ( .A(a[6265]), .B(c6265), .Z(n18797) );
XOR U31330 ( .A(c6266), .B(n18798), .Z(c6267) );
ANDN U31331 ( .B(n18799), .A(n18800), .Z(n18798) );
XOR U31332 ( .A(c6266), .B(b[6266]), .Z(n18799) );
XNOR U31333 ( .A(b[6266]), .B(n18800), .Z(c[6266]) );
XNOR U31334 ( .A(a[6266]), .B(c6266), .Z(n18800) );
XOR U31335 ( .A(c6267), .B(n18801), .Z(c6268) );
ANDN U31336 ( .B(n18802), .A(n18803), .Z(n18801) );
XOR U31337 ( .A(c6267), .B(b[6267]), .Z(n18802) );
XNOR U31338 ( .A(b[6267]), .B(n18803), .Z(c[6267]) );
XNOR U31339 ( .A(a[6267]), .B(c6267), .Z(n18803) );
XOR U31340 ( .A(c6268), .B(n18804), .Z(c6269) );
ANDN U31341 ( .B(n18805), .A(n18806), .Z(n18804) );
XOR U31342 ( .A(c6268), .B(b[6268]), .Z(n18805) );
XNOR U31343 ( .A(b[6268]), .B(n18806), .Z(c[6268]) );
XNOR U31344 ( .A(a[6268]), .B(c6268), .Z(n18806) );
XOR U31345 ( .A(c6269), .B(n18807), .Z(c6270) );
ANDN U31346 ( .B(n18808), .A(n18809), .Z(n18807) );
XOR U31347 ( .A(c6269), .B(b[6269]), .Z(n18808) );
XNOR U31348 ( .A(b[6269]), .B(n18809), .Z(c[6269]) );
XNOR U31349 ( .A(a[6269]), .B(c6269), .Z(n18809) );
XOR U31350 ( .A(c6270), .B(n18810), .Z(c6271) );
ANDN U31351 ( .B(n18811), .A(n18812), .Z(n18810) );
XOR U31352 ( .A(c6270), .B(b[6270]), .Z(n18811) );
XNOR U31353 ( .A(b[6270]), .B(n18812), .Z(c[6270]) );
XNOR U31354 ( .A(a[6270]), .B(c6270), .Z(n18812) );
XOR U31355 ( .A(c6271), .B(n18813), .Z(c6272) );
ANDN U31356 ( .B(n18814), .A(n18815), .Z(n18813) );
XOR U31357 ( .A(c6271), .B(b[6271]), .Z(n18814) );
XNOR U31358 ( .A(b[6271]), .B(n18815), .Z(c[6271]) );
XNOR U31359 ( .A(a[6271]), .B(c6271), .Z(n18815) );
XOR U31360 ( .A(c6272), .B(n18816), .Z(c6273) );
ANDN U31361 ( .B(n18817), .A(n18818), .Z(n18816) );
XOR U31362 ( .A(c6272), .B(b[6272]), .Z(n18817) );
XNOR U31363 ( .A(b[6272]), .B(n18818), .Z(c[6272]) );
XNOR U31364 ( .A(a[6272]), .B(c6272), .Z(n18818) );
XOR U31365 ( .A(c6273), .B(n18819), .Z(c6274) );
ANDN U31366 ( .B(n18820), .A(n18821), .Z(n18819) );
XOR U31367 ( .A(c6273), .B(b[6273]), .Z(n18820) );
XNOR U31368 ( .A(b[6273]), .B(n18821), .Z(c[6273]) );
XNOR U31369 ( .A(a[6273]), .B(c6273), .Z(n18821) );
XOR U31370 ( .A(c6274), .B(n18822), .Z(c6275) );
ANDN U31371 ( .B(n18823), .A(n18824), .Z(n18822) );
XOR U31372 ( .A(c6274), .B(b[6274]), .Z(n18823) );
XNOR U31373 ( .A(b[6274]), .B(n18824), .Z(c[6274]) );
XNOR U31374 ( .A(a[6274]), .B(c6274), .Z(n18824) );
XOR U31375 ( .A(c6275), .B(n18825), .Z(c6276) );
ANDN U31376 ( .B(n18826), .A(n18827), .Z(n18825) );
XOR U31377 ( .A(c6275), .B(b[6275]), .Z(n18826) );
XNOR U31378 ( .A(b[6275]), .B(n18827), .Z(c[6275]) );
XNOR U31379 ( .A(a[6275]), .B(c6275), .Z(n18827) );
XOR U31380 ( .A(c6276), .B(n18828), .Z(c6277) );
ANDN U31381 ( .B(n18829), .A(n18830), .Z(n18828) );
XOR U31382 ( .A(c6276), .B(b[6276]), .Z(n18829) );
XNOR U31383 ( .A(b[6276]), .B(n18830), .Z(c[6276]) );
XNOR U31384 ( .A(a[6276]), .B(c6276), .Z(n18830) );
XOR U31385 ( .A(c6277), .B(n18831), .Z(c6278) );
ANDN U31386 ( .B(n18832), .A(n18833), .Z(n18831) );
XOR U31387 ( .A(c6277), .B(b[6277]), .Z(n18832) );
XNOR U31388 ( .A(b[6277]), .B(n18833), .Z(c[6277]) );
XNOR U31389 ( .A(a[6277]), .B(c6277), .Z(n18833) );
XOR U31390 ( .A(c6278), .B(n18834), .Z(c6279) );
ANDN U31391 ( .B(n18835), .A(n18836), .Z(n18834) );
XOR U31392 ( .A(c6278), .B(b[6278]), .Z(n18835) );
XNOR U31393 ( .A(b[6278]), .B(n18836), .Z(c[6278]) );
XNOR U31394 ( .A(a[6278]), .B(c6278), .Z(n18836) );
XOR U31395 ( .A(c6279), .B(n18837), .Z(c6280) );
ANDN U31396 ( .B(n18838), .A(n18839), .Z(n18837) );
XOR U31397 ( .A(c6279), .B(b[6279]), .Z(n18838) );
XNOR U31398 ( .A(b[6279]), .B(n18839), .Z(c[6279]) );
XNOR U31399 ( .A(a[6279]), .B(c6279), .Z(n18839) );
XOR U31400 ( .A(c6280), .B(n18840), .Z(c6281) );
ANDN U31401 ( .B(n18841), .A(n18842), .Z(n18840) );
XOR U31402 ( .A(c6280), .B(b[6280]), .Z(n18841) );
XNOR U31403 ( .A(b[6280]), .B(n18842), .Z(c[6280]) );
XNOR U31404 ( .A(a[6280]), .B(c6280), .Z(n18842) );
XOR U31405 ( .A(c6281), .B(n18843), .Z(c6282) );
ANDN U31406 ( .B(n18844), .A(n18845), .Z(n18843) );
XOR U31407 ( .A(c6281), .B(b[6281]), .Z(n18844) );
XNOR U31408 ( .A(b[6281]), .B(n18845), .Z(c[6281]) );
XNOR U31409 ( .A(a[6281]), .B(c6281), .Z(n18845) );
XOR U31410 ( .A(c6282), .B(n18846), .Z(c6283) );
ANDN U31411 ( .B(n18847), .A(n18848), .Z(n18846) );
XOR U31412 ( .A(c6282), .B(b[6282]), .Z(n18847) );
XNOR U31413 ( .A(b[6282]), .B(n18848), .Z(c[6282]) );
XNOR U31414 ( .A(a[6282]), .B(c6282), .Z(n18848) );
XOR U31415 ( .A(c6283), .B(n18849), .Z(c6284) );
ANDN U31416 ( .B(n18850), .A(n18851), .Z(n18849) );
XOR U31417 ( .A(c6283), .B(b[6283]), .Z(n18850) );
XNOR U31418 ( .A(b[6283]), .B(n18851), .Z(c[6283]) );
XNOR U31419 ( .A(a[6283]), .B(c6283), .Z(n18851) );
XOR U31420 ( .A(c6284), .B(n18852), .Z(c6285) );
ANDN U31421 ( .B(n18853), .A(n18854), .Z(n18852) );
XOR U31422 ( .A(c6284), .B(b[6284]), .Z(n18853) );
XNOR U31423 ( .A(b[6284]), .B(n18854), .Z(c[6284]) );
XNOR U31424 ( .A(a[6284]), .B(c6284), .Z(n18854) );
XOR U31425 ( .A(c6285), .B(n18855), .Z(c6286) );
ANDN U31426 ( .B(n18856), .A(n18857), .Z(n18855) );
XOR U31427 ( .A(c6285), .B(b[6285]), .Z(n18856) );
XNOR U31428 ( .A(b[6285]), .B(n18857), .Z(c[6285]) );
XNOR U31429 ( .A(a[6285]), .B(c6285), .Z(n18857) );
XOR U31430 ( .A(c6286), .B(n18858), .Z(c6287) );
ANDN U31431 ( .B(n18859), .A(n18860), .Z(n18858) );
XOR U31432 ( .A(c6286), .B(b[6286]), .Z(n18859) );
XNOR U31433 ( .A(b[6286]), .B(n18860), .Z(c[6286]) );
XNOR U31434 ( .A(a[6286]), .B(c6286), .Z(n18860) );
XOR U31435 ( .A(c6287), .B(n18861), .Z(c6288) );
ANDN U31436 ( .B(n18862), .A(n18863), .Z(n18861) );
XOR U31437 ( .A(c6287), .B(b[6287]), .Z(n18862) );
XNOR U31438 ( .A(b[6287]), .B(n18863), .Z(c[6287]) );
XNOR U31439 ( .A(a[6287]), .B(c6287), .Z(n18863) );
XOR U31440 ( .A(c6288), .B(n18864), .Z(c6289) );
ANDN U31441 ( .B(n18865), .A(n18866), .Z(n18864) );
XOR U31442 ( .A(c6288), .B(b[6288]), .Z(n18865) );
XNOR U31443 ( .A(b[6288]), .B(n18866), .Z(c[6288]) );
XNOR U31444 ( .A(a[6288]), .B(c6288), .Z(n18866) );
XOR U31445 ( .A(c6289), .B(n18867), .Z(c6290) );
ANDN U31446 ( .B(n18868), .A(n18869), .Z(n18867) );
XOR U31447 ( .A(c6289), .B(b[6289]), .Z(n18868) );
XNOR U31448 ( .A(b[6289]), .B(n18869), .Z(c[6289]) );
XNOR U31449 ( .A(a[6289]), .B(c6289), .Z(n18869) );
XOR U31450 ( .A(c6290), .B(n18870), .Z(c6291) );
ANDN U31451 ( .B(n18871), .A(n18872), .Z(n18870) );
XOR U31452 ( .A(c6290), .B(b[6290]), .Z(n18871) );
XNOR U31453 ( .A(b[6290]), .B(n18872), .Z(c[6290]) );
XNOR U31454 ( .A(a[6290]), .B(c6290), .Z(n18872) );
XOR U31455 ( .A(c6291), .B(n18873), .Z(c6292) );
ANDN U31456 ( .B(n18874), .A(n18875), .Z(n18873) );
XOR U31457 ( .A(c6291), .B(b[6291]), .Z(n18874) );
XNOR U31458 ( .A(b[6291]), .B(n18875), .Z(c[6291]) );
XNOR U31459 ( .A(a[6291]), .B(c6291), .Z(n18875) );
XOR U31460 ( .A(c6292), .B(n18876), .Z(c6293) );
ANDN U31461 ( .B(n18877), .A(n18878), .Z(n18876) );
XOR U31462 ( .A(c6292), .B(b[6292]), .Z(n18877) );
XNOR U31463 ( .A(b[6292]), .B(n18878), .Z(c[6292]) );
XNOR U31464 ( .A(a[6292]), .B(c6292), .Z(n18878) );
XOR U31465 ( .A(c6293), .B(n18879), .Z(c6294) );
ANDN U31466 ( .B(n18880), .A(n18881), .Z(n18879) );
XOR U31467 ( .A(c6293), .B(b[6293]), .Z(n18880) );
XNOR U31468 ( .A(b[6293]), .B(n18881), .Z(c[6293]) );
XNOR U31469 ( .A(a[6293]), .B(c6293), .Z(n18881) );
XOR U31470 ( .A(c6294), .B(n18882), .Z(c6295) );
ANDN U31471 ( .B(n18883), .A(n18884), .Z(n18882) );
XOR U31472 ( .A(c6294), .B(b[6294]), .Z(n18883) );
XNOR U31473 ( .A(b[6294]), .B(n18884), .Z(c[6294]) );
XNOR U31474 ( .A(a[6294]), .B(c6294), .Z(n18884) );
XOR U31475 ( .A(c6295), .B(n18885), .Z(c6296) );
ANDN U31476 ( .B(n18886), .A(n18887), .Z(n18885) );
XOR U31477 ( .A(c6295), .B(b[6295]), .Z(n18886) );
XNOR U31478 ( .A(b[6295]), .B(n18887), .Z(c[6295]) );
XNOR U31479 ( .A(a[6295]), .B(c6295), .Z(n18887) );
XOR U31480 ( .A(c6296), .B(n18888), .Z(c6297) );
ANDN U31481 ( .B(n18889), .A(n18890), .Z(n18888) );
XOR U31482 ( .A(c6296), .B(b[6296]), .Z(n18889) );
XNOR U31483 ( .A(b[6296]), .B(n18890), .Z(c[6296]) );
XNOR U31484 ( .A(a[6296]), .B(c6296), .Z(n18890) );
XOR U31485 ( .A(c6297), .B(n18891), .Z(c6298) );
ANDN U31486 ( .B(n18892), .A(n18893), .Z(n18891) );
XOR U31487 ( .A(c6297), .B(b[6297]), .Z(n18892) );
XNOR U31488 ( .A(b[6297]), .B(n18893), .Z(c[6297]) );
XNOR U31489 ( .A(a[6297]), .B(c6297), .Z(n18893) );
XOR U31490 ( .A(c6298), .B(n18894), .Z(c6299) );
ANDN U31491 ( .B(n18895), .A(n18896), .Z(n18894) );
XOR U31492 ( .A(c6298), .B(b[6298]), .Z(n18895) );
XNOR U31493 ( .A(b[6298]), .B(n18896), .Z(c[6298]) );
XNOR U31494 ( .A(a[6298]), .B(c6298), .Z(n18896) );
XOR U31495 ( .A(c6299), .B(n18897), .Z(c6300) );
ANDN U31496 ( .B(n18898), .A(n18899), .Z(n18897) );
XOR U31497 ( .A(c6299), .B(b[6299]), .Z(n18898) );
XNOR U31498 ( .A(b[6299]), .B(n18899), .Z(c[6299]) );
XNOR U31499 ( .A(a[6299]), .B(c6299), .Z(n18899) );
XOR U31500 ( .A(c6300), .B(n18900), .Z(c6301) );
ANDN U31501 ( .B(n18901), .A(n18902), .Z(n18900) );
XOR U31502 ( .A(c6300), .B(b[6300]), .Z(n18901) );
XNOR U31503 ( .A(b[6300]), .B(n18902), .Z(c[6300]) );
XNOR U31504 ( .A(a[6300]), .B(c6300), .Z(n18902) );
XOR U31505 ( .A(c6301), .B(n18903), .Z(c6302) );
ANDN U31506 ( .B(n18904), .A(n18905), .Z(n18903) );
XOR U31507 ( .A(c6301), .B(b[6301]), .Z(n18904) );
XNOR U31508 ( .A(b[6301]), .B(n18905), .Z(c[6301]) );
XNOR U31509 ( .A(a[6301]), .B(c6301), .Z(n18905) );
XOR U31510 ( .A(c6302), .B(n18906), .Z(c6303) );
ANDN U31511 ( .B(n18907), .A(n18908), .Z(n18906) );
XOR U31512 ( .A(c6302), .B(b[6302]), .Z(n18907) );
XNOR U31513 ( .A(b[6302]), .B(n18908), .Z(c[6302]) );
XNOR U31514 ( .A(a[6302]), .B(c6302), .Z(n18908) );
XOR U31515 ( .A(c6303), .B(n18909), .Z(c6304) );
ANDN U31516 ( .B(n18910), .A(n18911), .Z(n18909) );
XOR U31517 ( .A(c6303), .B(b[6303]), .Z(n18910) );
XNOR U31518 ( .A(b[6303]), .B(n18911), .Z(c[6303]) );
XNOR U31519 ( .A(a[6303]), .B(c6303), .Z(n18911) );
XOR U31520 ( .A(c6304), .B(n18912), .Z(c6305) );
ANDN U31521 ( .B(n18913), .A(n18914), .Z(n18912) );
XOR U31522 ( .A(c6304), .B(b[6304]), .Z(n18913) );
XNOR U31523 ( .A(b[6304]), .B(n18914), .Z(c[6304]) );
XNOR U31524 ( .A(a[6304]), .B(c6304), .Z(n18914) );
XOR U31525 ( .A(c6305), .B(n18915), .Z(c6306) );
ANDN U31526 ( .B(n18916), .A(n18917), .Z(n18915) );
XOR U31527 ( .A(c6305), .B(b[6305]), .Z(n18916) );
XNOR U31528 ( .A(b[6305]), .B(n18917), .Z(c[6305]) );
XNOR U31529 ( .A(a[6305]), .B(c6305), .Z(n18917) );
XOR U31530 ( .A(c6306), .B(n18918), .Z(c6307) );
ANDN U31531 ( .B(n18919), .A(n18920), .Z(n18918) );
XOR U31532 ( .A(c6306), .B(b[6306]), .Z(n18919) );
XNOR U31533 ( .A(b[6306]), .B(n18920), .Z(c[6306]) );
XNOR U31534 ( .A(a[6306]), .B(c6306), .Z(n18920) );
XOR U31535 ( .A(c6307), .B(n18921), .Z(c6308) );
ANDN U31536 ( .B(n18922), .A(n18923), .Z(n18921) );
XOR U31537 ( .A(c6307), .B(b[6307]), .Z(n18922) );
XNOR U31538 ( .A(b[6307]), .B(n18923), .Z(c[6307]) );
XNOR U31539 ( .A(a[6307]), .B(c6307), .Z(n18923) );
XOR U31540 ( .A(c6308), .B(n18924), .Z(c6309) );
ANDN U31541 ( .B(n18925), .A(n18926), .Z(n18924) );
XOR U31542 ( .A(c6308), .B(b[6308]), .Z(n18925) );
XNOR U31543 ( .A(b[6308]), .B(n18926), .Z(c[6308]) );
XNOR U31544 ( .A(a[6308]), .B(c6308), .Z(n18926) );
XOR U31545 ( .A(c6309), .B(n18927), .Z(c6310) );
ANDN U31546 ( .B(n18928), .A(n18929), .Z(n18927) );
XOR U31547 ( .A(c6309), .B(b[6309]), .Z(n18928) );
XNOR U31548 ( .A(b[6309]), .B(n18929), .Z(c[6309]) );
XNOR U31549 ( .A(a[6309]), .B(c6309), .Z(n18929) );
XOR U31550 ( .A(c6310), .B(n18930), .Z(c6311) );
ANDN U31551 ( .B(n18931), .A(n18932), .Z(n18930) );
XOR U31552 ( .A(c6310), .B(b[6310]), .Z(n18931) );
XNOR U31553 ( .A(b[6310]), .B(n18932), .Z(c[6310]) );
XNOR U31554 ( .A(a[6310]), .B(c6310), .Z(n18932) );
XOR U31555 ( .A(c6311), .B(n18933), .Z(c6312) );
ANDN U31556 ( .B(n18934), .A(n18935), .Z(n18933) );
XOR U31557 ( .A(c6311), .B(b[6311]), .Z(n18934) );
XNOR U31558 ( .A(b[6311]), .B(n18935), .Z(c[6311]) );
XNOR U31559 ( .A(a[6311]), .B(c6311), .Z(n18935) );
XOR U31560 ( .A(c6312), .B(n18936), .Z(c6313) );
ANDN U31561 ( .B(n18937), .A(n18938), .Z(n18936) );
XOR U31562 ( .A(c6312), .B(b[6312]), .Z(n18937) );
XNOR U31563 ( .A(b[6312]), .B(n18938), .Z(c[6312]) );
XNOR U31564 ( .A(a[6312]), .B(c6312), .Z(n18938) );
XOR U31565 ( .A(c6313), .B(n18939), .Z(c6314) );
ANDN U31566 ( .B(n18940), .A(n18941), .Z(n18939) );
XOR U31567 ( .A(c6313), .B(b[6313]), .Z(n18940) );
XNOR U31568 ( .A(b[6313]), .B(n18941), .Z(c[6313]) );
XNOR U31569 ( .A(a[6313]), .B(c6313), .Z(n18941) );
XOR U31570 ( .A(c6314), .B(n18942), .Z(c6315) );
ANDN U31571 ( .B(n18943), .A(n18944), .Z(n18942) );
XOR U31572 ( .A(c6314), .B(b[6314]), .Z(n18943) );
XNOR U31573 ( .A(b[6314]), .B(n18944), .Z(c[6314]) );
XNOR U31574 ( .A(a[6314]), .B(c6314), .Z(n18944) );
XOR U31575 ( .A(c6315), .B(n18945), .Z(c6316) );
ANDN U31576 ( .B(n18946), .A(n18947), .Z(n18945) );
XOR U31577 ( .A(c6315), .B(b[6315]), .Z(n18946) );
XNOR U31578 ( .A(b[6315]), .B(n18947), .Z(c[6315]) );
XNOR U31579 ( .A(a[6315]), .B(c6315), .Z(n18947) );
XOR U31580 ( .A(c6316), .B(n18948), .Z(c6317) );
ANDN U31581 ( .B(n18949), .A(n18950), .Z(n18948) );
XOR U31582 ( .A(c6316), .B(b[6316]), .Z(n18949) );
XNOR U31583 ( .A(b[6316]), .B(n18950), .Z(c[6316]) );
XNOR U31584 ( .A(a[6316]), .B(c6316), .Z(n18950) );
XOR U31585 ( .A(c6317), .B(n18951), .Z(c6318) );
ANDN U31586 ( .B(n18952), .A(n18953), .Z(n18951) );
XOR U31587 ( .A(c6317), .B(b[6317]), .Z(n18952) );
XNOR U31588 ( .A(b[6317]), .B(n18953), .Z(c[6317]) );
XNOR U31589 ( .A(a[6317]), .B(c6317), .Z(n18953) );
XOR U31590 ( .A(c6318), .B(n18954), .Z(c6319) );
ANDN U31591 ( .B(n18955), .A(n18956), .Z(n18954) );
XOR U31592 ( .A(c6318), .B(b[6318]), .Z(n18955) );
XNOR U31593 ( .A(b[6318]), .B(n18956), .Z(c[6318]) );
XNOR U31594 ( .A(a[6318]), .B(c6318), .Z(n18956) );
XOR U31595 ( .A(c6319), .B(n18957), .Z(c6320) );
ANDN U31596 ( .B(n18958), .A(n18959), .Z(n18957) );
XOR U31597 ( .A(c6319), .B(b[6319]), .Z(n18958) );
XNOR U31598 ( .A(b[6319]), .B(n18959), .Z(c[6319]) );
XNOR U31599 ( .A(a[6319]), .B(c6319), .Z(n18959) );
XOR U31600 ( .A(c6320), .B(n18960), .Z(c6321) );
ANDN U31601 ( .B(n18961), .A(n18962), .Z(n18960) );
XOR U31602 ( .A(c6320), .B(b[6320]), .Z(n18961) );
XNOR U31603 ( .A(b[6320]), .B(n18962), .Z(c[6320]) );
XNOR U31604 ( .A(a[6320]), .B(c6320), .Z(n18962) );
XOR U31605 ( .A(c6321), .B(n18963), .Z(c6322) );
ANDN U31606 ( .B(n18964), .A(n18965), .Z(n18963) );
XOR U31607 ( .A(c6321), .B(b[6321]), .Z(n18964) );
XNOR U31608 ( .A(b[6321]), .B(n18965), .Z(c[6321]) );
XNOR U31609 ( .A(a[6321]), .B(c6321), .Z(n18965) );
XOR U31610 ( .A(c6322), .B(n18966), .Z(c6323) );
ANDN U31611 ( .B(n18967), .A(n18968), .Z(n18966) );
XOR U31612 ( .A(c6322), .B(b[6322]), .Z(n18967) );
XNOR U31613 ( .A(b[6322]), .B(n18968), .Z(c[6322]) );
XNOR U31614 ( .A(a[6322]), .B(c6322), .Z(n18968) );
XOR U31615 ( .A(c6323), .B(n18969), .Z(c6324) );
ANDN U31616 ( .B(n18970), .A(n18971), .Z(n18969) );
XOR U31617 ( .A(c6323), .B(b[6323]), .Z(n18970) );
XNOR U31618 ( .A(b[6323]), .B(n18971), .Z(c[6323]) );
XNOR U31619 ( .A(a[6323]), .B(c6323), .Z(n18971) );
XOR U31620 ( .A(c6324), .B(n18972), .Z(c6325) );
ANDN U31621 ( .B(n18973), .A(n18974), .Z(n18972) );
XOR U31622 ( .A(c6324), .B(b[6324]), .Z(n18973) );
XNOR U31623 ( .A(b[6324]), .B(n18974), .Z(c[6324]) );
XNOR U31624 ( .A(a[6324]), .B(c6324), .Z(n18974) );
XOR U31625 ( .A(c6325), .B(n18975), .Z(c6326) );
ANDN U31626 ( .B(n18976), .A(n18977), .Z(n18975) );
XOR U31627 ( .A(c6325), .B(b[6325]), .Z(n18976) );
XNOR U31628 ( .A(b[6325]), .B(n18977), .Z(c[6325]) );
XNOR U31629 ( .A(a[6325]), .B(c6325), .Z(n18977) );
XOR U31630 ( .A(c6326), .B(n18978), .Z(c6327) );
ANDN U31631 ( .B(n18979), .A(n18980), .Z(n18978) );
XOR U31632 ( .A(c6326), .B(b[6326]), .Z(n18979) );
XNOR U31633 ( .A(b[6326]), .B(n18980), .Z(c[6326]) );
XNOR U31634 ( .A(a[6326]), .B(c6326), .Z(n18980) );
XOR U31635 ( .A(c6327), .B(n18981), .Z(c6328) );
ANDN U31636 ( .B(n18982), .A(n18983), .Z(n18981) );
XOR U31637 ( .A(c6327), .B(b[6327]), .Z(n18982) );
XNOR U31638 ( .A(b[6327]), .B(n18983), .Z(c[6327]) );
XNOR U31639 ( .A(a[6327]), .B(c6327), .Z(n18983) );
XOR U31640 ( .A(c6328), .B(n18984), .Z(c6329) );
ANDN U31641 ( .B(n18985), .A(n18986), .Z(n18984) );
XOR U31642 ( .A(c6328), .B(b[6328]), .Z(n18985) );
XNOR U31643 ( .A(b[6328]), .B(n18986), .Z(c[6328]) );
XNOR U31644 ( .A(a[6328]), .B(c6328), .Z(n18986) );
XOR U31645 ( .A(c6329), .B(n18987), .Z(c6330) );
ANDN U31646 ( .B(n18988), .A(n18989), .Z(n18987) );
XOR U31647 ( .A(c6329), .B(b[6329]), .Z(n18988) );
XNOR U31648 ( .A(b[6329]), .B(n18989), .Z(c[6329]) );
XNOR U31649 ( .A(a[6329]), .B(c6329), .Z(n18989) );
XOR U31650 ( .A(c6330), .B(n18990), .Z(c6331) );
ANDN U31651 ( .B(n18991), .A(n18992), .Z(n18990) );
XOR U31652 ( .A(c6330), .B(b[6330]), .Z(n18991) );
XNOR U31653 ( .A(b[6330]), .B(n18992), .Z(c[6330]) );
XNOR U31654 ( .A(a[6330]), .B(c6330), .Z(n18992) );
XOR U31655 ( .A(c6331), .B(n18993), .Z(c6332) );
ANDN U31656 ( .B(n18994), .A(n18995), .Z(n18993) );
XOR U31657 ( .A(c6331), .B(b[6331]), .Z(n18994) );
XNOR U31658 ( .A(b[6331]), .B(n18995), .Z(c[6331]) );
XNOR U31659 ( .A(a[6331]), .B(c6331), .Z(n18995) );
XOR U31660 ( .A(c6332), .B(n18996), .Z(c6333) );
ANDN U31661 ( .B(n18997), .A(n18998), .Z(n18996) );
XOR U31662 ( .A(c6332), .B(b[6332]), .Z(n18997) );
XNOR U31663 ( .A(b[6332]), .B(n18998), .Z(c[6332]) );
XNOR U31664 ( .A(a[6332]), .B(c6332), .Z(n18998) );
XOR U31665 ( .A(c6333), .B(n18999), .Z(c6334) );
ANDN U31666 ( .B(n19000), .A(n19001), .Z(n18999) );
XOR U31667 ( .A(c6333), .B(b[6333]), .Z(n19000) );
XNOR U31668 ( .A(b[6333]), .B(n19001), .Z(c[6333]) );
XNOR U31669 ( .A(a[6333]), .B(c6333), .Z(n19001) );
XOR U31670 ( .A(c6334), .B(n19002), .Z(c6335) );
ANDN U31671 ( .B(n19003), .A(n19004), .Z(n19002) );
XOR U31672 ( .A(c6334), .B(b[6334]), .Z(n19003) );
XNOR U31673 ( .A(b[6334]), .B(n19004), .Z(c[6334]) );
XNOR U31674 ( .A(a[6334]), .B(c6334), .Z(n19004) );
XOR U31675 ( .A(c6335), .B(n19005), .Z(c6336) );
ANDN U31676 ( .B(n19006), .A(n19007), .Z(n19005) );
XOR U31677 ( .A(c6335), .B(b[6335]), .Z(n19006) );
XNOR U31678 ( .A(b[6335]), .B(n19007), .Z(c[6335]) );
XNOR U31679 ( .A(a[6335]), .B(c6335), .Z(n19007) );
XOR U31680 ( .A(c6336), .B(n19008), .Z(c6337) );
ANDN U31681 ( .B(n19009), .A(n19010), .Z(n19008) );
XOR U31682 ( .A(c6336), .B(b[6336]), .Z(n19009) );
XNOR U31683 ( .A(b[6336]), .B(n19010), .Z(c[6336]) );
XNOR U31684 ( .A(a[6336]), .B(c6336), .Z(n19010) );
XOR U31685 ( .A(c6337), .B(n19011), .Z(c6338) );
ANDN U31686 ( .B(n19012), .A(n19013), .Z(n19011) );
XOR U31687 ( .A(c6337), .B(b[6337]), .Z(n19012) );
XNOR U31688 ( .A(b[6337]), .B(n19013), .Z(c[6337]) );
XNOR U31689 ( .A(a[6337]), .B(c6337), .Z(n19013) );
XOR U31690 ( .A(c6338), .B(n19014), .Z(c6339) );
ANDN U31691 ( .B(n19015), .A(n19016), .Z(n19014) );
XOR U31692 ( .A(c6338), .B(b[6338]), .Z(n19015) );
XNOR U31693 ( .A(b[6338]), .B(n19016), .Z(c[6338]) );
XNOR U31694 ( .A(a[6338]), .B(c6338), .Z(n19016) );
XOR U31695 ( .A(c6339), .B(n19017), .Z(c6340) );
ANDN U31696 ( .B(n19018), .A(n19019), .Z(n19017) );
XOR U31697 ( .A(c6339), .B(b[6339]), .Z(n19018) );
XNOR U31698 ( .A(b[6339]), .B(n19019), .Z(c[6339]) );
XNOR U31699 ( .A(a[6339]), .B(c6339), .Z(n19019) );
XOR U31700 ( .A(c6340), .B(n19020), .Z(c6341) );
ANDN U31701 ( .B(n19021), .A(n19022), .Z(n19020) );
XOR U31702 ( .A(c6340), .B(b[6340]), .Z(n19021) );
XNOR U31703 ( .A(b[6340]), .B(n19022), .Z(c[6340]) );
XNOR U31704 ( .A(a[6340]), .B(c6340), .Z(n19022) );
XOR U31705 ( .A(c6341), .B(n19023), .Z(c6342) );
ANDN U31706 ( .B(n19024), .A(n19025), .Z(n19023) );
XOR U31707 ( .A(c6341), .B(b[6341]), .Z(n19024) );
XNOR U31708 ( .A(b[6341]), .B(n19025), .Z(c[6341]) );
XNOR U31709 ( .A(a[6341]), .B(c6341), .Z(n19025) );
XOR U31710 ( .A(c6342), .B(n19026), .Z(c6343) );
ANDN U31711 ( .B(n19027), .A(n19028), .Z(n19026) );
XOR U31712 ( .A(c6342), .B(b[6342]), .Z(n19027) );
XNOR U31713 ( .A(b[6342]), .B(n19028), .Z(c[6342]) );
XNOR U31714 ( .A(a[6342]), .B(c6342), .Z(n19028) );
XOR U31715 ( .A(c6343), .B(n19029), .Z(c6344) );
ANDN U31716 ( .B(n19030), .A(n19031), .Z(n19029) );
XOR U31717 ( .A(c6343), .B(b[6343]), .Z(n19030) );
XNOR U31718 ( .A(b[6343]), .B(n19031), .Z(c[6343]) );
XNOR U31719 ( .A(a[6343]), .B(c6343), .Z(n19031) );
XOR U31720 ( .A(c6344), .B(n19032), .Z(c6345) );
ANDN U31721 ( .B(n19033), .A(n19034), .Z(n19032) );
XOR U31722 ( .A(c6344), .B(b[6344]), .Z(n19033) );
XNOR U31723 ( .A(b[6344]), .B(n19034), .Z(c[6344]) );
XNOR U31724 ( .A(a[6344]), .B(c6344), .Z(n19034) );
XOR U31725 ( .A(c6345), .B(n19035), .Z(c6346) );
ANDN U31726 ( .B(n19036), .A(n19037), .Z(n19035) );
XOR U31727 ( .A(c6345), .B(b[6345]), .Z(n19036) );
XNOR U31728 ( .A(b[6345]), .B(n19037), .Z(c[6345]) );
XNOR U31729 ( .A(a[6345]), .B(c6345), .Z(n19037) );
XOR U31730 ( .A(c6346), .B(n19038), .Z(c6347) );
ANDN U31731 ( .B(n19039), .A(n19040), .Z(n19038) );
XOR U31732 ( .A(c6346), .B(b[6346]), .Z(n19039) );
XNOR U31733 ( .A(b[6346]), .B(n19040), .Z(c[6346]) );
XNOR U31734 ( .A(a[6346]), .B(c6346), .Z(n19040) );
XOR U31735 ( .A(c6347), .B(n19041), .Z(c6348) );
ANDN U31736 ( .B(n19042), .A(n19043), .Z(n19041) );
XOR U31737 ( .A(c6347), .B(b[6347]), .Z(n19042) );
XNOR U31738 ( .A(b[6347]), .B(n19043), .Z(c[6347]) );
XNOR U31739 ( .A(a[6347]), .B(c6347), .Z(n19043) );
XOR U31740 ( .A(c6348), .B(n19044), .Z(c6349) );
ANDN U31741 ( .B(n19045), .A(n19046), .Z(n19044) );
XOR U31742 ( .A(c6348), .B(b[6348]), .Z(n19045) );
XNOR U31743 ( .A(b[6348]), .B(n19046), .Z(c[6348]) );
XNOR U31744 ( .A(a[6348]), .B(c6348), .Z(n19046) );
XOR U31745 ( .A(c6349), .B(n19047), .Z(c6350) );
ANDN U31746 ( .B(n19048), .A(n19049), .Z(n19047) );
XOR U31747 ( .A(c6349), .B(b[6349]), .Z(n19048) );
XNOR U31748 ( .A(b[6349]), .B(n19049), .Z(c[6349]) );
XNOR U31749 ( .A(a[6349]), .B(c6349), .Z(n19049) );
XOR U31750 ( .A(c6350), .B(n19050), .Z(c6351) );
ANDN U31751 ( .B(n19051), .A(n19052), .Z(n19050) );
XOR U31752 ( .A(c6350), .B(b[6350]), .Z(n19051) );
XNOR U31753 ( .A(b[6350]), .B(n19052), .Z(c[6350]) );
XNOR U31754 ( .A(a[6350]), .B(c6350), .Z(n19052) );
XOR U31755 ( .A(c6351), .B(n19053), .Z(c6352) );
ANDN U31756 ( .B(n19054), .A(n19055), .Z(n19053) );
XOR U31757 ( .A(c6351), .B(b[6351]), .Z(n19054) );
XNOR U31758 ( .A(b[6351]), .B(n19055), .Z(c[6351]) );
XNOR U31759 ( .A(a[6351]), .B(c6351), .Z(n19055) );
XOR U31760 ( .A(c6352), .B(n19056), .Z(c6353) );
ANDN U31761 ( .B(n19057), .A(n19058), .Z(n19056) );
XOR U31762 ( .A(c6352), .B(b[6352]), .Z(n19057) );
XNOR U31763 ( .A(b[6352]), .B(n19058), .Z(c[6352]) );
XNOR U31764 ( .A(a[6352]), .B(c6352), .Z(n19058) );
XOR U31765 ( .A(c6353), .B(n19059), .Z(c6354) );
ANDN U31766 ( .B(n19060), .A(n19061), .Z(n19059) );
XOR U31767 ( .A(c6353), .B(b[6353]), .Z(n19060) );
XNOR U31768 ( .A(b[6353]), .B(n19061), .Z(c[6353]) );
XNOR U31769 ( .A(a[6353]), .B(c6353), .Z(n19061) );
XOR U31770 ( .A(c6354), .B(n19062), .Z(c6355) );
ANDN U31771 ( .B(n19063), .A(n19064), .Z(n19062) );
XOR U31772 ( .A(c6354), .B(b[6354]), .Z(n19063) );
XNOR U31773 ( .A(b[6354]), .B(n19064), .Z(c[6354]) );
XNOR U31774 ( .A(a[6354]), .B(c6354), .Z(n19064) );
XOR U31775 ( .A(c6355), .B(n19065), .Z(c6356) );
ANDN U31776 ( .B(n19066), .A(n19067), .Z(n19065) );
XOR U31777 ( .A(c6355), .B(b[6355]), .Z(n19066) );
XNOR U31778 ( .A(b[6355]), .B(n19067), .Z(c[6355]) );
XNOR U31779 ( .A(a[6355]), .B(c6355), .Z(n19067) );
XOR U31780 ( .A(c6356), .B(n19068), .Z(c6357) );
ANDN U31781 ( .B(n19069), .A(n19070), .Z(n19068) );
XOR U31782 ( .A(c6356), .B(b[6356]), .Z(n19069) );
XNOR U31783 ( .A(b[6356]), .B(n19070), .Z(c[6356]) );
XNOR U31784 ( .A(a[6356]), .B(c6356), .Z(n19070) );
XOR U31785 ( .A(c6357), .B(n19071), .Z(c6358) );
ANDN U31786 ( .B(n19072), .A(n19073), .Z(n19071) );
XOR U31787 ( .A(c6357), .B(b[6357]), .Z(n19072) );
XNOR U31788 ( .A(b[6357]), .B(n19073), .Z(c[6357]) );
XNOR U31789 ( .A(a[6357]), .B(c6357), .Z(n19073) );
XOR U31790 ( .A(c6358), .B(n19074), .Z(c6359) );
ANDN U31791 ( .B(n19075), .A(n19076), .Z(n19074) );
XOR U31792 ( .A(c6358), .B(b[6358]), .Z(n19075) );
XNOR U31793 ( .A(b[6358]), .B(n19076), .Z(c[6358]) );
XNOR U31794 ( .A(a[6358]), .B(c6358), .Z(n19076) );
XOR U31795 ( .A(c6359), .B(n19077), .Z(c6360) );
ANDN U31796 ( .B(n19078), .A(n19079), .Z(n19077) );
XOR U31797 ( .A(c6359), .B(b[6359]), .Z(n19078) );
XNOR U31798 ( .A(b[6359]), .B(n19079), .Z(c[6359]) );
XNOR U31799 ( .A(a[6359]), .B(c6359), .Z(n19079) );
XOR U31800 ( .A(c6360), .B(n19080), .Z(c6361) );
ANDN U31801 ( .B(n19081), .A(n19082), .Z(n19080) );
XOR U31802 ( .A(c6360), .B(b[6360]), .Z(n19081) );
XNOR U31803 ( .A(b[6360]), .B(n19082), .Z(c[6360]) );
XNOR U31804 ( .A(a[6360]), .B(c6360), .Z(n19082) );
XOR U31805 ( .A(c6361), .B(n19083), .Z(c6362) );
ANDN U31806 ( .B(n19084), .A(n19085), .Z(n19083) );
XOR U31807 ( .A(c6361), .B(b[6361]), .Z(n19084) );
XNOR U31808 ( .A(b[6361]), .B(n19085), .Z(c[6361]) );
XNOR U31809 ( .A(a[6361]), .B(c6361), .Z(n19085) );
XOR U31810 ( .A(c6362), .B(n19086), .Z(c6363) );
ANDN U31811 ( .B(n19087), .A(n19088), .Z(n19086) );
XOR U31812 ( .A(c6362), .B(b[6362]), .Z(n19087) );
XNOR U31813 ( .A(b[6362]), .B(n19088), .Z(c[6362]) );
XNOR U31814 ( .A(a[6362]), .B(c6362), .Z(n19088) );
XOR U31815 ( .A(c6363), .B(n19089), .Z(c6364) );
ANDN U31816 ( .B(n19090), .A(n19091), .Z(n19089) );
XOR U31817 ( .A(c6363), .B(b[6363]), .Z(n19090) );
XNOR U31818 ( .A(b[6363]), .B(n19091), .Z(c[6363]) );
XNOR U31819 ( .A(a[6363]), .B(c6363), .Z(n19091) );
XOR U31820 ( .A(c6364), .B(n19092), .Z(c6365) );
ANDN U31821 ( .B(n19093), .A(n19094), .Z(n19092) );
XOR U31822 ( .A(c6364), .B(b[6364]), .Z(n19093) );
XNOR U31823 ( .A(b[6364]), .B(n19094), .Z(c[6364]) );
XNOR U31824 ( .A(a[6364]), .B(c6364), .Z(n19094) );
XOR U31825 ( .A(c6365), .B(n19095), .Z(c6366) );
ANDN U31826 ( .B(n19096), .A(n19097), .Z(n19095) );
XOR U31827 ( .A(c6365), .B(b[6365]), .Z(n19096) );
XNOR U31828 ( .A(b[6365]), .B(n19097), .Z(c[6365]) );
XNOR U31829 ( .A(a[6365]), .B(c6365), .Z(n19097) );
XOR U31830 ( .A(c6366), .B(n19098), .Z(c6367) );
ANDN U31831 ( .B(n19099), .A(n19100), .Z(n19098) );
XOR U31832 ( .A(c6366), .B(b[6366]), .Z(n19099) );
XNOR U31833 ( .A(b[6366]), .B(n19100), .Z(c[6366]) );
XNOR U31834 ( .A(a[6366]), .B(c6366), .Z(n19100) );
XOR U31835 ( .A(c6367), .B(n19101), .Z(c6368) );
ANDN U31836 ( .B(n19102), .A(n19103), .Z(n19101) );
XOR U31837 ( .A(c6367), .B(b[6367]), .Z(n19102) );
XNOR U31838 ( .A(b[6367]), .B(n19103), .Z(c[6367]) );
XNOR U31839 ( .A(a[6367]), .B(c6367), .Z(n19103) );
XOR U31840 ( .A(c6368), .B(n19104), .Z(c6369) );
ANDN U31841 ( .B(n19105), .A(n19106), .Z(n19104) );
XOR U31842 ( .A(c6368), .B(b[6368]), .Z(n19105) );
XNOR U31843 ( .A(b[6368]), .B(n19106), .Z(c[6368]) );
XNOR U31844 ( .A(a[6368]), .B(c6368), .Z(n19106) );
XOR U31845 ( .A(c6369), .B(n19107), .Z(c6370) );
ANDN U31846 ( .B(n19108), .A(n19109), .Z(n19107) );
XOR U31847 ( .A(c6369), .B(b[6369]), .Z(n19108) );
XNOR U31848 ( .A(b[6369]), .B(n19109), .Z(c[6369]) );
XNOR U31849 ( .A(a[6369]), .B(c6369), .Z(n19109) );
XOR U31850 ( .A(c6370), .B(n19110), .Z(c6371) );
ANDN U31851 ( .B(n19111), .A(n19112), .Z(n19110) );
XOR U31852 ( .A(c6370), .B(b[6370]), .Z(n19111) );
XNOR U31853 ( .A(b[6370]), .B(n19112), .Z(c[6370]) );
XNOR U31854 ( .A(a[6370]), .B(c6370), .Z(n19112) );
XOR U31855 ( .A(c6371), .B(n19113), .Z(c6372) );
ANDN U31856 ( .B(n19114), .A(n19115), .Z(n19113) );
XOR U31857 ( .A(c6371), .B(b[6371]), .Z(n19114) );
XNOR U31858 ( .A(b[6371]), .B(n19115), .Z(c[6371]) );
XNOR U31859 ( .A(a[6371]), .B(c6371), .Z(n19115) );
XOR U31860 ( .A(c6372), .B(n19116), .Z(c6373) );
ANDN U31861 ( .B(n19117), .A(n19118), .Z(n19116) );
XOR U31862 ( .A(c6372), .B(b[6372]), .Z(n19117) );
XNOR U31863 ( .A(b[6372]), .B(n19118), .Z(c[6372]) );
XNOR U31864 ( .A(a[6372]), .B(c6372), .Z(n19118) );
XOR U31865 ( .A(c6373), .B(n19119), .Z(c6374) );
ANDN U31866 ( .B(n19120), .A(n19121), .Z(n19119) );
XOR U31867 ( .A(c6373), .B(b[6373]), .Z(n19120) );
XNOR U31868 ( .A(b[6373]), .B(n19121), .Z(c[6373]) );
XNOR U31869 ( .A(a[6373]), .B(c6373), .Z(n19121) );
XOR U31870 ( .A(c6374), .B(n19122), .Z(c6375) );
ANDN U31871 ( .B(n19123), .A(n19124), .Z(n19122) );
XOR U31872 ( .A(c6374), .B(b[6374]), .Z(n19123) );
XNOR U31873 ( .A(b[6374]), .B(n19124), .Z(c[6374]) );
XNOR U31874 ( .A(a[6374]), .B(c6374), .Z(n19124) );
XOR U31875 ( .A(c6375), .B(n19125), .Z(c6376) );
ANDN U31876 ( .B(n19126), .A(n19127), .Z(n19125) );
XOR U31877 ( .A(c6375), .B(b[6375]), .Z(n19126) );
XNOR U31878 ( .A(b[6375]), .B(n19127), .Z(c[6375]) );
XNOR U31879 ( .A(a[6375]), .B(c6375), .Z(n19127) );
XOR U31880 ( .A(c6376), .B(n19128), .Z(c6377) );
ANDN U31881 ( .B(n19129), .A(n19130), .Z(n19128) );
XOR U31882 ( .A(c6376), .B(b[6376]), .Z(n19129) );
XNOR U31883 ( .A(b[6376]), .B(n19130), .Z(c[6376]) );
XNOR U31884 ( .A(a[6376]), .B(c6376), .Z(n19130) );
XOR U31885 ( .A(c6377), .B(n19131), .Z(c6378) );
ANDN U31886 ( .B(n19132), .A(n19133), .Z(n19131) );
XOR U31887 ( .A(c6377), .B(b[6377]), .Z(n19132) );
XNOR U31888 ( .A(b[6377]), .B(n19133), .Z(c[6377]) );
XNOR U31889 ( .A(a[6377]), .B(c6377), .Z(n19133) );
XOR U31890 ( .A(c6378), .B(n19134), .Z(c6379) );
ANDN U31891 ( .B(n19135), .A(n19136), .Z(n19134) );
XOR U31892 ( .A(c6378), .B(b[6378]), .Z(n19135) );
XNOR U31893 ( .A(b[6378]), .B(n19136), .Z(c[6378]) );
XNOR U31894 ( .A(a[6378]), .B(c6378), .Z(n19136) );
XOR U31895 ( .A(c6379), .B(n19137), .Z(c6380) );
ANDN U31896 ( .B(n19138), .A(n19139), .Z(n19137) );
XOR U31897 ( .A(c6379), .B(b[6379]), .Z(n19138) );
XNOR U31898 ( .A(b[6379]), .B(n19139), .Z(c[6379]) );
XNOR U31899 ( .A(a[6379]), .B(c6379), .Z(n19139) );
XOR U31900 ( .A(c6380), .B(n19140), .Z(c6381) );
ANDN U31901 ( .B(n19141), .A(n19142), .Z(n19140) );
XOR U31902 ( .A(c6380), .B(b[6380]), .Z(n19141) );
XNOR U31903 ( .A(b[6380]), .B(n19142), .Z(c[6380]) );
XNOR U31904 ( .A(a[6380]), .B(c6380), .Z(n19142) );
XOR U31905 ( .A(c6381), .B(n19143), .Z(c6382) );
ANDN U31906 ( .B(n19144), .A(n19145), .Z(n19143) );
XOR U31907 ( .A(c6381), .B(b[6381]), .Z(n19144) );
XNOR U31908 ( .A(b[6381]), .B(n19145), .Z(c[6381]) );
XNOR U31909 ( .A(a[6381]), .B(c6381), .Z(n19145) );
XOR U31910 ( .A(c6382), .B(n19146), .Z(c6383) );
ANDN U31911 ( .B(n19147), .A(n19148), .Z(n19146) );
XOR U31912 ( .A(c6382), .B(b[6382]), .Z(n19147) );
XNOR U31913 ( .A(b[6382]), .B(n19148), .Z(c[6382]) );
XNOR U31914 ( .A(a[6382]), .B(c6382), .Z(n19148) );
XOR U31915 ( .A(c6383), .B(n19149), .Z(c6384) );
ANDN U31916 ( .B(n19150), .A(n19151), .Z(n19149) );
XOR U31917 ( .A(c6383), .B(b[6383]), .Z(n19150) );
XNOR U31918 ( .A(b[6383]), .B(n19151), .Z(c[6383]) );
XNOR U31919 ( .A(a[6383]), .B(c6383), .Z(n19151) );
XOR U31920 ( .A(c6384), .B(n19152), .Z(c6385) );
ANDN U31921 ( .B(n19153), .A(n19154), .Z(n19152) );
XOR U31922 ( .A(c6384), .B(b[6384]), .Z(n19153) );
XNOR U31923 ( .A(b[6384]), .B(n19154), .Z(c[6384]) );
XNOR U31924 ( .A(a[6384]), .B(c6384), .Z(n19154) );
XOR U31925 ( .A(c6385), .B(n19155), .Z(c6386) );
ANDN U31926 ( .B(n19156), .A(n19157), .Z(n19155) );
XOR U31927 ( .A(c6385), .B(b[6385]), .Z(n19156) );
XNOR U31928 ( .A(b[6385]), .B(n19157), .Z(c[6385]) );
XNOR U31929 ( .A(a[6385]), .B(c6385), .Z(n19157) );
XOR U31930 ( .A(c6386), .B(n19158), .Z(c6387) );
ANDN U31931 ( .B(n19159), .A(n19160), .Z(n19158) );
XOR U31932 ( .A(c6386), .B(b[6386]), .Z(n19159) );
XNOR U31933 ( .A(b[6386]), .B(n19160), .Z(c[6386]) );
XNOR U31934 ( .A(a[6386]), .B(c6386), .Z(n19160) );
XOR U31935 ( .A(c6387), .B(n19161), .Z(c6388) );
ANDN U31936 ( .B(n19162), .A(n19163), .Z(n19161) );
XOR U31937 ( .A(c6387), .B(b[6387]), .Z(n19162) );
XNOR U31938 ( .A(b[6387]), .B(n19163), .Z(c[6387]) );
XNOR U31939 ( .A(a[6387]), .B(c6387), .Z(n19163) );
XOR U31940 ( .A(c6388), .B(n19164), .Z(c6389) );
ANDN U31941 ( .B(n19165), .A(n19166), .Z(n19164) );
XOR U31942 ( .A(c6388), .B(b[6388]), .Z(n19165) );
XNOR U31943 ( .A(b[6388]), .B(n19166), .Z(c[6388]) );
XNOR U31944 ( .A(a[6388]), .B(c6388), .Z(n19166) );
XOR U31945 ( .A(c6389), .B(n19167), .Z(c6390) );
ANDN U31946 ( .B(n19168), .A(n19169), .Z(n19167) );
XOR U31947 ( .A(c6389), .B(b[6389]), .Z(n19168) );
XNOR U31948 ( .A(b[6389]), .B(n19169), .Z(c[6389]) );
XNOR U31949 ( .A(a[6389]), .B(c6389), .Z(n19169) );
XOR U31950 ( .A(c6390), .B(n19170), .Z(c6391) );
ANDN U31951 ( .B(n19171), .A(n19172), .Z(n19170) );
XOR U31952 ( .A(c6390), .B(b[6390]), .Z(n19171) );
XNOR U31953 ( .A(b[6390]), .B(n19172), .Z(c[6390]) );
XNOR U31954 ( .A(a[6390]), .B(c6390), .Z(n19172) );
XOR U31955 ( .A(c6391), .B(n19173), .Z(c6392) );
ANDN U31956 ( .B(n19174), .A(n19175), .Z(n19173) );
XOR U31957 ( .A(c6391), .B(b[6391]), .Z(n19174) );
XNOR U31958 ( .A(b[6391]), .B(n19175), .Z(c[6391]) );
XNOR U31959 ( .A(a[6391]), .B(c6391), .Z(n19175) );
XOR U31960 ( .A(c6392), .B(n19176), .Z(c6393) );
ANDN U31961 ( .B(n19177), .A(n19178), .Z(n19176) );
XOR U31962 ( .A(c6392), .B(b[6392]), .Z(n19177) );
XNOR U31963 ( .A(b[6392]), .B(n19178), .Z(c[6392]) );
XNOR U31964 ( .A(a[6392]), .B(c6392), .Z(n19178) );
XOR U31965 ( .A(c6393), .B(n19179), .Z(c6394) );
ANDN U31966 ( .B(n19180), .A(n19181), .Z(n19179) );
XOR U31967 ( .A(c6393), .B(b[6393]), .Z(n19180) );
XNOR U31968 ( .A(b[6393]), .B(n19181), .Z(c[6393]) );
XNOR U31969 ( .A(a[6393]), .B(c6393), .Z(n19181) );
XOR U31970 ( .A(c6394), .B(n19182), .Z(c6395) );
ANDN U31971 ( .B(n19183), .A(n19184), .Z(n19182) );
XOR U31972 ( .A(c6394), .B(b[6394]), .Z(n19183) );
XNOR U31973 ( .A(b[6394]), .B(n19184), .Z(c[6394]) );
XNOR U31974 ( .A(a[6394]), .B(c6394), .Z(n19184) );
XOR U31975 ( .A(c6395), .B(n19185), .Z(c6396) );
ANDN U31976 ( .B(n19186), .A(n19187), .Z(n19185) );
XOR U31977 ( .A(c6395), .B(b[6395]), .Z(n19186) );
XNOR U31978 ( .A(b[6395]), .B(n19187), .Z(c[6395]) );
XNOR U31979 ( .A(a[6395]), .B(c6395), .Z(n19187) );
XOR U31980 ( .A(c6396), .B(n19188), .Z(c6397) );
ANDN U31981 ( .B(n19189), .A(n19190), .Z(n19188) );
XOR U31982 ( .A(c6396), .B(b[6396]), .Z(n19189) );
XNOR U31983 ( .A(b[6396]), .B(n19190), .Z(c[6396]) );
XNOR U31984 ( .A(a[6396]), .B(c6396), .Z(n19190) );
XOR U31985 ( .A(c6397), .B(n19191), .Z(c6398) );
ANDN U31986 ( .B(n19192), .A(n19193), .Z(n19191) );
XOR U31987 ( .A(c6397), .B(b[6397]), .Z(n19192) );
XNOR U31988 ( .A(b[6397]), .B(n19193), .Z(c[6397]) );
XNOR U31989 ( .A(a[6397]), .B(c6397), .Z(n19193) );
XOR U31990 ( .A(c6398), .B(n19194), .Z(c6399) );
ANDN U31991 ( .B(n19195), .A(n19196), .Z(n19194) );
XOR U31992 ( .A(c6398), .B(b[6398]), .Z(n19195) );
XNOR U31993 ( .A(b[6398]), .B(n19196), .Z(c[6398]) );
XNOR U31994 ( .A(a[6398]), .B(c6398), .Z(n19196) );
XOR U31995 ( .A(c6399), .B(n19197), .Z(c6400) );
ANDN U31996 ( .B(n19198), .A(n19199), .Z(n19197) );
XOR U31997 ( .A(c6399), .B(b[6399]), .Z(n19198) );
XNOR U31998 ( .A(b[6399]), .B(n19199), .Z(c[6399]) );
XNOR U31999 ( .A(a[6399]), .B(c6399), .Z(n19199) );
XOR U32000 ( .A(c6400), .B(n19200), .Z(c6401) );
ANDN U32001 ( .B(n19201), .A(n19202), .Z(n19200) );
XOR U32002 ( .A(c6400), .B(b[6400]), .Z(n19201) );
XNOR U32003 ( .A(b[6400]), .B(n19202), .Z(c[6400]) );
XNOR U32004 ( .A(a[6400]), .B(c6400), .Z(n19202) );
XOR U32005 ( .A(c6401), .B(n19203), .Z(c6402) );
ANDN U32006 ( .B(n19204), .A(n19205), .Z(n19203) );
XOR U32007 ( .A(c6401), .B(b[6401]), .Z(n19204) );
XNOR U32008 ( .A(b[6401]), .B(n19205), .Z(c[6401]) );
XNOR U32009 ( .A(a[6401]), .B(c6401), .Z(n19205) );
XOR U32010 ( .A(c6402), .B(n19206), .Z(c6403) );
ANDN U32011 ( .B(n19207), .A(n19208), .Z(n19206) );
XOR U32012 ( .A(c6402), .B(b[6402]), .Z(n19207) );
XNOR U32013 ( .A(b[6402]), .B(n19208), .Z(c[6402]) );
XNOR U32014 ( .A(a[6402]), .B(c6402), .Z(n19208) );
XOR U32015 ( .A(c6403), .B(n19209), .Z(c6404) );
ANDN U32016 ( .B(n19210), .A(n19211), .Z(n19209) );
XOR U32017 ( .A(c6403), .B(b[6403]), .Z(n19210) );
XNOR U32018 ( .A(b[6403]), .B(n19211), .Z(c[6403]) );
XNOR U32019 ( .A(a[6403]), .B(c6403), .Z(n19211) );
XOR U32020 ( .A(c6404), .B(n19212), .Z(c6405) );
ANDN U32021 ( .B(n19213), .A(n19214), .Z(n19212) );
XOR U32022 ( .A(c6404), .B(b[6404]), .Z(n19213) );
XNOR U32023 ( .A(b[6404]), .B(n19214), .Z(c[6404]) );
XNOR U32024 ( .A(a[6404]), .B(c6404), .Z(n19214) );
XOR U32025 ( .A(c6405), .B(n19215), .Z(c6406) );
ANDN U32026 ( .B(n19216), .A(n19217), .Z(n19215) );
XOR U32027 ( .A(c6405), .B(b[6405]), .Z(n19216) );
XNOR U32028 ( .A(b[6405]), .B(n19217), .Z(c[6405]) );
XNOR U32029 ( .A(a[6405]), .B(c6405), .Z(n19217) );
XOR U32030 ( .A(c6406), .B(n19218), .Z(c6407) );
ANDN U32031 ( .B(n19219), .A(n19220), .Z(n19218) );
XOR U32032 ( .A(c6406), .B(b[6406]), .Z(n19219) );
XNOR U32033 ( .A(b[6406]), .B(n19220), .Z(c[6406]) );
XNOR U32034 ( .A(a[6406]), .B(c6406), .Z(n19220) );
XOR U32035 ( .A(c6407), .B(n19221), .Z(c6408) );
ANDN U32036 ( .B(n19222), .A(n19223), .Z(n19221) );
XOR U32037 ( .A(c6407), .B(b[6407]), .Z(n19222) );
XNOR U32038 ( .A(b[6407]), .B(n19223), .Z(c[6407]) );
XNOR U32039 ( .A(a[6407]), .B(c6407), .Z(n19223) );
XOR U32040 ( .A(c6408), .B(n19224), .Z(c6409) );
ANDN U32041 ( .B(n19225), .A(n19226), .Z(n19224) );
XOR U32042 ( .A(c6408), .B(b[6408]), .Z(n19225) );
XNOR U32043 ( .A(b[6408]), .B(n19226), .Z(c[6408]) );
XNOR U32044 ( .A(a[6408]), .B(c6408), .Z(n19226) );
XOR U32045 ( .A(c6409), .B(n19227), .Z(c6410) );
ANDN U32046 ( .B(n19228), .A(n19229), .Z(n19227) );
XOR U32047 ( .A(c6409), .B(b[6409]), .Z(n19228) );
XNOR U32048 ( .A(b[6409]), .B(n19229), .Z(c[6409]) );
XNOR U32049 ( .A(a[6409]), .B(c6409), .Z(n19229) );
XOR U32050 ( .A(c6410), .B(n19230), .Z(c6411) );
ANDN U32051 ( .B(n19231), .A(n19232), .Z(n19230) );
XOR U32052 ( .A(c6410), .B(b[6410]), .Z(n19231) );
XNOR U32053 ( .A(b[6410]), .B(n19232), .Z(c[6410]) );
XNOR U32054 ( .A(a[6410]), .B(c6410), .Z(n19232) );
XOR U32055 ( .A(c6411), .B(n19233), .Z(c6412) );
ANDN U32056 ( .B(n19234), .A(n19235), .Z(n19233) );
XOR U32057 ( .A(c6411), .B(b[6411]), .Z(n19234) );
XNOR U32058 ( .A(b[6411]), .B(n19235), .Z(c[6411]) );
XNOR U32059 ( .A(a[6411]), .B(c6411), .Z(n19235) );
XOR U32060 ( .A(c6412), .B(n19236), .Z(c6413) );
ANDN U32061 ( .B(n19237), .A(n19238), .Z(n19236) );
XOR U32062 ( .A(c6412), .B(b[6412]), .Z(n19237) );
XNOR U32063 ( .A(b[6412]), .B(n19238), .Z(c[6412]) );
XNOR U32064 ( .A(a[6412]), .B(c6412), .Z(n19238) );
XOR U32065 ( .A(c6413), .B(n19239), .Z(c6414) );
ANDN U32066 ( .B(n19240), .A(n19241), .Z(n19239) );
XOR U32067 ( .A(c6413), .B(b[6413]), .Z(n19240) );
XNOR U32068 ( .A(b[6413]), .B(n19241), .Z(c[6413]) );
XNOR U32069 ( .A(a[6413]), .B(c6413), .Z(n19241) );
XOR U32070 ( .A(c6414), .B(n19242), .Z(c6415) );
ANDN U32071 ( .B(n19243), .A(n19244), .Z(n19242) );
XOR U32072 ( .A(c6414), .B(b[6414]), .Z(n19243) );
XNOR U32073 ( .A(b[6414]), .B(n19244), .Z(c[6414]) );
XNOR U32074 ( .A(a[6414]), .B(c6414), .Z(n19244) );
XOR U32075 ( .A(c6415), .B(n19245), .Z(c6416) );
ANDN U32076 ( .B(n19246), .A(n19247), .Z(n19245) );
XOR U32077 ( .A(c6415), .B(b[6415]), .Z(n19246) );
XNOR U32078 ( .A(b[6415]), .B(n19247), .Z(c[6415]) );
XNOR U32079 ( .A(a[6415]), .B(c6415), .Z(n19247) );
XOR U32080 ( .A(c6416), .B(n19248), .Z(c6417) );
ANDN U32081 ( .B(n19249), .A(n19250), .Z(n19248) );
XOR U32082 ( .A(c6416), .B(b[6416]), .Z(n19249) );
XNOR U32083 ( .A(b[6416]), .B(n19250), .Z(c[6416]) );
XNOR U32084 ( .A(a[6416]), .B(c6416), .Z(n19250) );
XOR U32085 ( .A(c6417), .B(n19251), .Z(c6418) );
ANDN U32086 ( .B(n19252), .A(n19253), .Z(n19251) );
XOR U32087 ( .A(c6417), .B(b[6417]), .Z(n19252) );
XNOR U32088 ( .A(b[6417]), .B(n19253), .Z(c[6417]) );
XNOR U32089 ( .A(a[6417]), .B(c6417), .Z(n19253) );
XOR U32090 ( .A(c6418), .B(n19254), .Z(c6419) );
ANDN U32091 ( .B(n19255), .A(n19256), .Z(n19254) );
XOR U32092 ( .A(c6418), .B(b[6418]), .Z(n19255) );
XNOR U32093 ( .A(b[6418]), .B(n19256), .Z(c[6418]) );
XNOR U32094 ( .A(a[6418]), .B(c6418), .Z(n19256) );
XOR U32095 ( .A(c6419), .B(n19257), .Z(c6420) );
ANDN U32096 ( .B(n19258), .A(n19259), .Z(n19257) );
XOR U32097 ( .A(c6419), .B(b[6419]), .Z(n19258) );
XNOR U32098 ( .A(b[6419]), .B(n19259), .Z(c[6419]) );
XNOR U32099 ( .A(a[6419]), .B(c6419), .Z(n19259) );
XOR U32100 ( .A(c6420), .B(n19260), .Z(c6421) );
ANDN U32101 ( .B(n19261), .A(n19262), .Z(n19260) );
XOR U32102 ( .A(c6420), .B(b[6420]), .Z(n19261) );
XNOR U32103 ( .A(b[6420]), .B(n19262), .Z(c[6420]) );
XNOR U32104 ( .A(a[6420]), .B(c6420), .Z(n19262) );
XOR U32105 ( .A(c6421), .B(n19263), .Z(c6422) );
ANDN U32106 ( .B(n19264), .A(n19265), .Z(n19263) );
XOR U32107 ( .A(c6421), .B(b[6421]), .Z(n19264) );
XNOR U32108 ( .A(b[6421]), .B(n19265), .Z(c[6421]) );
XNOR U32109 ( .A(a[6421]), .B(c6421), .Z(n19265) );
XOR U32110 ( .A(c6422), .B(n19266), .Z(c6423) );
ANDN U32111 ( .B(n19267), .A(n19268), .Z(n19266) );
XOR U32112 ( .A(c6422), .B(b[6422]), .Z(n19267) );
XNOR U32113 ( .A(b[6422]), .B(n19268), .Z(c[6422]) );
XNOR U32114 ( .A(a[6422]), .B(c6422), .Z(n19268) );
XOR U32115 ( .A(c6423), .B(n19269), .Z(c6424) );
ANDN U32116 ( .B(n19270), .A(n19271), .Z(n19269) );
XOR U32117 ( .A(c6423), .B(b[6423]), .Z(n19270) );
XNOR U32118 ( .A(b[6423]), .B(n19271), .Z(c[6423]) );
XNOR U32119 ( .A(a[6423]), .B(c6423), .Z(n19271) );
XOR U32120 ( .A(c6424), .B(n19272), .Z(c6425) );
ANDN U32121 ( .B(n19273), .A(n19274), .Z(n19272) );
XOR U32122 ( .A(c6424), .B(b[6424]), .Z(n19273) );
XNOR U32123 ( .A(b[6424]), .B(n19274), .Z(c[6424]) );
XNOR U32124 ( .A(a[6424]), .B(c6424), .Z(n19274) );
XOR U32125 ( .A(c6425), .B(n19275), .Z(c6426) );
ANDN U32126 ( .B(n19276), .A(n19277), .Z(n19275) );
XOR U32127 ( .A(c6425), .B(b[6425]), .Z(n19276) );
XNOR U32128 ( .A(b[6425]), .B(n19277), .Z(c[6425]) );
XNOR U32129 ( .A(a[6425]), .B(c6425), .Z(n19277) );
XOR U32130 ( .A(c6426), .B(n19278), .Z(c6427) );
ANDN U32131 ( .B(n19279), .A(n19280), .Z(n19278) );
XOR U32132 ( .A(c6426), .B(b[6426]), .Z(n19279) );
XNOR U32133 ( .A(b[6426]), .B(n19280), .Z(c[6426]) );
XNOR U32134 ( .A(a[6426]), .B(c6426), .Z(n19280) );
XOR U32135 ( .A(c6427), .B(n19281), .Z(c6428) );
ANDN U32136 ( .B(n19282), .A(n19283), .Z(n19281) );
XOR U32137 ( .A(c6427), .B(b[6427]), .Z(n19282) );
XNOR U32138 ( .A(b[6427]), .B(n19283), .Z(c[6427]) );
XNOR U32139 ( .A(a[6427]), .B(c6427), .Z(n19283) );
XOR U32140 ( .A(c6428), .B(n19284), .Z(c6429) );
ANDN U32141 ( .B(n19285), .A(n19286), .Z(n19284) );
XOR U32142 ( .A(c6428), .B(b[6428]), .Z(n19285) );
XNOR U32143 ( .A(b[6428]), .B(n19286), .Z(c[6428]) );
XNOR U32144 ( .A(a[6428]), .B(c6428), .Z(n19286) );
XOR U32145 ( .A(c6429), .B(n19287), .Z(c6430) );
ANDN U32146 ( .B(n19288), .A(n19289), .Z(n19287) );
XOR U32147 ( .A(c6429), .B(b[6429]), .Z(n19288) );
XNOR U32148 ( .A(b[6429]), .B(n19289), .Z(c[6429]) );
XNOR U32149 ( .A(a[6429]), .B(c6429), .Z(n19289) );
XOR U32150 ( .A(c6430), .B(n19290), .Z(c6431) );
ANDN U32151 ( .B(n19291), .A(n19292), .Z(n19290) );
XOR U32152 ( .A(c6430), .B(b[6430]), .Z(n19291) );
XNOR U32153 ( .A(b[6430]), .B(n19292), .Z(c[6430]) );
XNOR U32154 ( .A(a[6430]), .B(c6430), .Z(n19292) );
XOR U32155 ( .A(c6431), .B(n19293), .Z(c6432) );
ANDN U32156 ( .B(n19294), .A(n19295), .Z(n19293) );
XOR U32157 ( .A(c6431), .B(b[6431]), .Z(n19294) );
XNOR U32158 ( .A(b[6431]), .B(n19295), .Z(c[6431]) );
XNOR U32159 ( .A(a[6431]), .B(c6431), .Z(n19295) );
XOR U32160 ( .A(c6432), .B(n19296), .Z(c6433) );
ANDN U32161 ( .B(n19297), .A(n19298), .Z(n19296) );
XOR U32162 ( .A(c6432), .B(b[6432]), .Z(n19297) );
XNOR U32163 ( .A(b[6432]), .B(n19298), .Z(c[6432]) );
XNOR U32164 ( .A(a[6432]), .B(c6432), .Z(n19298) );
XOR U32165 ( .A(c6433), .B(n19299), .Z(c6434) );
ANDN U32166 ( .B(n19300), .A(n19301), .Z(n19299) );
XOR U32167 ( .A(c6433), .B(b[6433]), .Z(n19300) );
XNOR U32168 ( .A(b[6433]), .B(n19301), .Z(c[6433]) );
XNOR U32169 ( .A(a[6433]), .B(c6433), .Z(n19301) );
XOR U32170 ( .A(c6434), .B(n19302), .Z(c6435) );
ANDN U32171 ( .B(n19303), .A(n19304), .Z(n19302) );
XOR U32172 ( .A(c6434), .B(b[6434]), .Z(n19303) );
XNOR U32173 ( .A(b[6434]), .B(n19304), .Z(c[6434]) );
XNOR U32174 ( .A(a[6434]), .B(c6434), .Z(n19304) );
XOR U32175 ( .A(c6435), .B(n19305), .Z(c6436) );
ANDN U32176 ( .B(n19306), .A(n19307), .Z(n19305) );
XOR U32177 ( .A(c6435), .B(b[6435]), .Z(n19306) );
XNOR U32178 ( .A(b[6435]), .B(n19307), .Z(c[6435]) );
XNOR U32179 ( .A(a[6435]), .B(c6435), .Z(n19307) );
XOR U32180 ( .A(c6436), .B(n19308), .Z(c6437) );
ANDN U32181 ( .B(n19309), .A(n19310), .Z(n19308) );
XOR U32182 ( .A(c6436), .B(b[6436]), .Z(n19309) );
XNOR U32183 ( .A(b[6436]), .B(n19310), .Z(c[6436]) );
XNOR U32184 ( .A(a[6436]), .B(c6436), .Z(n19310) );
XOR U32185 ( .A(c6437), .B(n19311), .Z(c6438) );
ANDN U32186 ( .B(n19312), .A(n19313), .Z(n19311) );
XOR U32187 ( .A(c6437), .B(b[6437]), .Z(n19312) );
XNOR U32188 ( .A(b[6437]), .B(n19313), .Z(c[6437]) );
XNOR U32189 ( .A(a[6437]), .B(c6437), .Z(n19313) );
XOR U32190 ( .A(c6438), .B(n19314), .Z(c6439) );
ANDN U32191 ( .B(n19315), .A(n19316), .Z(n19314) );
XOR U32192 ( .A(c6438), .B(b[6438]), .Z(n19315) );
XNOR U32193 ( .A(b[6438]), .B(n19316), .Z(c[6438]) );
XNOR U32194 ( .A(a[6438]), .B(c6438), .Z(n19316) );
XOR U32195 ( .A(c6439), .B(n19317), .Z(c6440) );
ANDN U32196 ( .B(n19318), .A(n19319), .Z(n19317) );
XOR U32197 ( .A(c6439), .B(b[6439]), .Z(n19318) );
XNOR U32198 ( .A(b[6439]), .B(n19319), .Z(c[6439]) );
XNOR U32199 ( .A(a[6439]), .B(c6439), .Z(n19319) );
XOR U32200 ( .A(c6440), .B(n19320), .Z(c6441) );
ANDN U32201 ( .B(n19321), .A(n19322), .Z(n19320) );
XOR U32202 ( .A(c6440), .B(b[6440]), .Z(n19321) );
XNOR U32203 ( .A(b[6440]), .B(n19322), .Z(c[6440]) );
XNOR U32204 ( .A(a[6440]), .B(c6440), .Z(n19322) );
XOR U32205 ( .A(c6441), .B(n19323), .Z(c6442) );
ANDN U32206 ( .B(n19324), .A(n19325), .Z(n19323) );
XOR U32207 ( .A(c6441), .B(b[6441]), .Z(n19324) );
XNOR U32208 ( .A(b[6441]), .B(n19325), .Z(c[6441]) );
XNOR U32209 ( .A(a[6441]), .B(c6441), .Z(n19325) );
XOR U32210 ( .A(c6442), .B(n19326), .Z(c6443) );
ANDN U32211 ( .B(n19327), .A(n19328), .Z(n19326) );
XOR U32212 ( .A(c6442), .B(b[6442]), .Z(n19327) );
XNOR U32213 ( .A(b[6442]), .B(n19328), .Z(c[6442]) );
XNOR U32214 ( .A(a[6442]), .B(c6442), .Z(n19328) );
XOR U32215 ( .A(c6443), .B(n19329), .Z(c6444) );
ANDN U32216 ( .B(n19330), .A(n19331), .Z(n19329) );
XOR U32217 ( .A(c6443), .B(b[6443]), .Z(n19330) );
XNOR U32218 ( .A(b[6443]), .B(n19331), .Z(c[6443]) );
XNOR U32219 ( .A(a[6443]), .B(c6443), .Z(n19331) );
XOR U32220 ( .A(c6444), .B(n19332), .Z(c6445) );
ANDN U32221 ( .B(n19333), .A(n19334), .Z(n19332) );
XOR U32222 ( .A(c6444), .B(b[6444]), .Z(n19333) );
XNOR U32223 ( .A(b[6444]), .B(n19334), .Z(c[6444]) );
XNOR U32224 ( .A(a[6444]), .B(c6444), .Z(n19334) );
XOR U32225 ( .A(c6445), .B(n19335), .Z(c6446) );
ANDN U32226 ( .B(n19336), .A(n19337), .Z(n19335) );
XOR U32227 ( .A(c6445), .B(b[6445]), .Z(n19336) );
XNOR U32228 ( .A(b[6445]), .B(n19337), .Z(c[6445]) );
XNOR U32229 ( .A(a[6445]), .B(c6445), .Z(n19337) );
XOR U32230 ( .A(c6446), .B(n19338), .Z(c6447) );
ANDN U32231 ( .B(n19339), .A(n19340), .Z(n19338) );
XOR U32232 ( .A(c6446), .B(b[6446]), .Z(n19339) );
XNOR U32233 ( .A(b[6446]), .B(n19340), .Z(c[6446]) );
XNOR U32234 ( .A(a[6446]), .B(c6446), .Z(n19340) );
XOR U32235 ( .A(c6447), .B(n19341), .Z(c6448) );
ANDN U32236 ( .B(n19342), .A(n19343), .Z(n19341) );
XOR U32237 ( .A(c6447), .B(b[6447]), .Z(n19342) );
XNOR U32238 ( .A(b[6447]), .B(n19343), .Z(c[6447]) );
XNOR U32239 ( .A(a[6447]), .B(c6447), .Z(n19343) );
XOR U32240 ( .A(c6448), .B(n19344), .Z(c6449) );
ANDN U32241 ( .B(n19345), .A(n19346), .Z(n19344) );
XOR U32242 ( .A(c6448), .B(b[6448]), .Z(n19345) );
XNOR U32243 ( .A(b[6448]), .B(n19346), .Z(c[6448]) );
XNOR U32244 ( .A(a[6448]), .B(c6448), .Z(n19346) );
XOR U32245 ( .A(c6449), .B(n19347), .Z(c6450) );
ANDN U32246 ( .B(n19348), .A(n19349), .Z(n19347) );
XOR U32247 ( .A(c6449), .B(b[6449]), .Z(n19348) );
XNOR U32248 ( .A(b[6449]), .B(n19349), .Z(c[6449]) );
XNOR U32249 ( .A(a[6449]), .B(c6449), .Z(n19349) );
XOR U32250 ( .A(c6450), .B(n19350), .Z(c6451) );
ANDN U32251 ( .B(n19351), .A(n19352), .Z(n19350) );
XOR U32252 ( .A(c6450), .B(b[6450]), .Z(n19351) );
XNOR U32253 ( .A(b[6450]), .B(n19352), .Z(c[6450]) );
XNOR U32254 ( .A(a[6450]), .B(c6450), .Z(n19352) );
XOR U32255 ( .A(c6451), .B(n19353), .Z(c6452) );
ANDN U32256 ( .B(n19354), .A(n19355), .Z(n19353) );
XOR U32257 ( .A(c6451), .B(b[6451]), .Z(n19354) );
XNOR U32258 ( .A(b[6451]), .B(n19355), .Z(c[6451]) );
XNOR U32259 ( .A(a[6451]), .B(c6451), .Z(n19355) );
XOR U32260 ( .A(c6452), .B(n19356), .Z(c6453) );
ANDN U32261 ( .B(n19357), .A(n19358), .Z(n19356) );
XOR U32262 ( .A(c6452), .B(b[6452]), .Z(n19357) );
XNOR U32263 ( .A(b[6452]), .B(n19358), .Z(c[6452]) );
XNOR U32264 ( .A(a[6452]), .B(c6452), .Z(n19358) );
XOR U32265 ( .A(c6453), .B(n19359), .Z(c6454) );
ANDN U32266 ( .B(n19360), .A(n19361), .Z(n19359) );
XOR U32267 ( .A(c6453), .B(b[6453]), .Z(n19360) );
XNOR U32268 ( .A(b[6453]), .B(n19361), .Z(c[6453]) );
XNOR U32269 ( .A(a[6453]), .B(c6453), .Z(n19361) );
XOR U32270 ( .A(c6454), .B(n19362), .Z(c6455) );
ANDN U32271 ( .B(n19363), .A(n19364), .Z(n19362) );
XOR U32272 ( .A(c6454), .B(b[6454]), .Z(n19363) );
XNOR U32273 ( .A(b[6454]), .B(n19364), .Z(c[6454]) );
XNOR U32274 ( .A(a[6454]), .B(c6454), .Z(n19364) );
XOR U32275 ( .A(c6455), .B(n19365), .Z(c6456) );
ANDN U32276 ( .B(n19366), .A(n19367), .Z(n19365) );
XOR U32277 ( .A(c6455), .B(b[6455]), .Z(n19366) );
XNOR U32278 ( .A(b[6455]), .B(n19367), .Z(c[6455]) );
XNOR U32279 ( .A(a[6455]), .B(c6455), .Z(n19367) );
XOR U32280 ( .A(c6456), .B(n19368), .Z(c6457) );
ANDN U32281 ( .B(n19369), .A(n19370), .Z(n19368) );
XOR U32282 ( .A(c6456), .B(b[6456]), .Z(n19369) );
XNOR U32283 ( .A(b[6456]), .B(n19370), .Z(c[6456]) );
XNOR U32284 ( .A(a[6456]), .B(c6456), .Z(n19370) );
XOR U32285 ( .A(c6457), .B(n19371), .Z(c6458) );
ANDN U32286 ( .B(n19372), .A(n19373), .Z(n19371) );
XOR U32287 ( .A(c6457), .B(b[6457]), .Z(n19372) );
XNOR U32288 ( .A(b[6457]), .B(n19373), .Z(c[6457]) );
XNOR U32289 ( .A(a[6457]), .B(c6457), .Z(n19373) );
XOR U32290 ( .A(c6458), .B(n19374), .Z(c6459) );
ANDN U32291 ( .B(n19375), .A(n19376), .Z(n19374) );
XOR U32292 ( .A(c6458), .B(b[6458]), .Z(n19375) );
XNOR U32293 ( .A(b[6458]), .B(n19376), .Z(c[6458]) );
XNOR U32294 ( .A(a[6458]), .B(c6458), .Z(n19376) );
XOR U32295 ( .A(c6459), .B(n19377), .Z(c6460) );
ANDN U32296 ( .B(n19378), .A(n19379), .Z(n19377) );
XOR U32297 ( .A(c6459), .B(b[6459]), .Z(n19378) );
XNOR U32298 ( .A(b[6459]), .B(n19379), .Z(c[6459]) );
XNOR U32299 ( .A(a[6459]), .B(c6459), .Z(n19379) );
XOR U32300 ( .A(c6460), .B(n19380), .Z(c6461) );
ANDN U32301 ( .B(n19381), .A(n19382), .Z(n19380) );
XOR U32302 ( .A(c6460), .B(b[6460]), .Z(n19381) );
XNOR U32303 ( .A(b[6460]), .B(n19382), .Z(c[6460]) );
XNOR U32304 ( .A(a[6460]), .B(c6460), .Z(n19382) );
XOR U32305 ( .A(c6461), .B(n19383), .Z(c6462) );
ANDN U32306 ( .B(n19384), .A(n19385), .Z(n19383) );
XOR U32307 ( .A(c6461), .B(b[6461]), .Z(n19384) );
XNOR U32308 ( .A(b[6461]), .B(n19385), .Z(c[6461]) );
XNOR U32309 ( .A(a[6461]), .B(c6461), .Z(n19385) );
XOR U32310 ( .A(c6462), .B(n19386), .Z(c6463) );
ANDN U32311 ( .B(n19387), .A(n19388), .Z(n19386) );
XOR U32312 ( .A(c6462), .B(b[6462]), .Z(n19387) );
XNOR U32313 ( .A(b[6462]), .B(n19388), .Z(c[6462]) );
XNOR U32314 ( .A(a[6462]), .B(c6462), .Z(n19388) );
XOR U32315 ( .A(c6463), .B(n19389), .Z(c6464) );
ANDN U32316 ( .B(n19390), .A(n19391), .Z(n19389) );
XOR U32317 ( .A(c6463), .B(b[6463]), .Z(n19390) );
XNOR U32318 ( .A(b[6463]), .B(n19391), .Z(c[6463]) );
XNOR U32319 ( .A(a[6463]), .B(c6463), .Z(n19391) );
XOR U32320 ( .A(c6464), .B(n19392), .Z(c6465) );
ANDN U32321 ( .B(n19393), .A(n19394), .Z(n19392) );
XOR U32322 ( .A(c6464), .B(b[6464]), .Z(n19393) );
XNOR U32323 ( .A(b[6464]), .B(n19394), .Z(c[6464]) );
XNOR U32324 ( .A(a[6464]), .B(c6464), .Z(n19394) );
XOR U32325 ( .A(c6465), .B(n19395), .Z(c6466) );
ANDN U32326 ( .B(n19396), .A(n19397), .Z(n19395) );
XOR U32327 ( .A(c6465), .B(b[6465]), .Z(n19396) );
XNOR U32328 ( .A(b[6465]), .B(n19397), .Z(c[6465]) );
XNOR U32329 ( .A(a[6465]), .B(c6465), .Z(n19397) );
XOR U32330 ( .A(c6466), .B(n19398), .Z(c6467) );
ANDN U32331 ( .B(n19399), .A(n19400), .Z(n19398) );
XOR U32332 ( .A(c6466), .B(b[6466]), .Z(n19399) );
XNOR U32333 ( .A(b[6466]), .B(n19400), .Z(c[6466]) );
XNOR U32334 ( .A(a[6466]), .B(c6466), .Z(n19400) );
XOR U32335 ( .A(c6467), .B(n19401), .Z(c6468) );
ANDN U32336 ( .B(n19402), .A(n19403), .Z(n19401) );
XOR U32337 ( .A(c6467), .B(b[6467]), .Z(n19402) );
XNOR U32338 ( .A(b[6467]), .B(n19403), .Z(c[6467]) );
XNOR U32339 ( .A(a[6467]), .B(c6467), .Z(n19403) );
XOR U32340 ( .A(c6468), .B(n19404), .Z(c6469) );
ANDN U32341 ( .B(n19405), .A(n19406), .Z(n19404) );
XOR U32342 ( .A(c6468), .B(b[6468]), .Z(n19405) );
XNOR U32343 ( .A(b[6468]), .B(n19406), .Z(c[6468]) );
XNOR U32344 ( .A(a[6468]), .B(c6468), .Z(n19406) );
XOR U32345 ( .A(c6469), .B(n19407), .Z(c6470) );
ANDN U32346 ( .B(n19408), .A(n19409), .Z(n19407) );
XOR U32347 ( .A(c6469), .B(b[6469]), .Z(n19408) );
XNOR U32348 ( .A(b[6469]), .B(n19409), .Z(c[6469]) );
XNOR U32349 ( .A(a[6469]), .B(c6469), .Z(n19409) );
XOR U32350 ( .A(c6470), .B(n19410), .Z(c6471) );
ANDN U32351 ( .B(n19411), .A(n19412), .Z(n19410) );
XOR U32352 ( .A(c6470), .B(b[6470]), .Z(n19411) );
XNOR U32353 ( .A(b[6470]), .B(n19412), .Z(c[6470]) );
XNOR U32354 ( .A(a[6470]), .B(c6470), .Z(n19412) );
XOR U32355 ( .A(c6471), .B(n19413), .Z(c6472) );
ANDN U32356 ( .B(n19414), .A(n19415), .Z(n19413) );
XOR U32357 ( .A(c6471), .B(b[6471]), .Z(n19414) );
XNOR U32358 ( .A(b[6471]), .B(n19415), .Z(c[6471]) );
XNOR U32359 ( .A(a[6471]), .B(c6471), .Z(n19415) );
XOR U32360 ( .A(c6472), .B(n19416), .Z(c6473) );
ANDN U32361 ( .B(n19417), .A(n19418), .Z(n19416) );
XOR U32362 ( .A(c6472), .B(b[6472]), .Z(n19417) );
XNOR U32363 ( .A(b[6472]), .B(n19418), .Z(c[6472]) );
XNOR U32364 ( .A(a[6472]), .B(c6472), .Z(n19418) );
XOR U32365 ( .A(c6473), .B(n19419), .Z(c6474) );
ANDN U32366 ( .B(n19420), .A(n19421), .Z(n19419) );
XOR U32367 ( .A(c6473), .B(b[6473]), .Z(n19420) );
XNOR U32368 ( .A(b[6473]), .B(n19421), .Z(c[6473]) );
XNOR U32369 ( .A(a[6473]), .B(c6473), .Z(n19421) );
XOR U32370 ( .A(c6474), .B(n19422), .Z(c6475) );
ANDN U32371 ( .B(n19423), .A(n19424), .Z(n19422) );
XOR U32372 ( .A(c6474), .B(b[6474]), .Z(n19423) );
XNOR U32373 ( .A(b[6474]), .B(n19424), .Z(c[6474]) );
XNOR U32374 ( .A(a[6474]), .B(c6474), .Z(n19424) );
XOR U32375 ( .A(c6475), .B(n19425), .Z(c6476) );
ANDN U32376 ( .B(n19426), .A(n19427), .Z(n19425) );
XOR U32377 ( .A(c6475), .B(b[6475]), .Z(n19426) );
XNOR U32378 ( .A(b[6475]), .B(n19427), .Z(c[6475]) );
XNOR U32379 ( .A(a[6475]), .B(c6475), .Z(n19427) );
XOR U32380 ( .A(c6476), .B(n19428), .Z(c6477) );
ANDN U32381 ( .B(n19429), .A(n19430), .Z(n19428) );
XOR U32382 ( .A(c6476), .B(b[6476]), .Z(n19429) );
XNOR U32383 ( .A(b[6476]), .B(n19430), .Z(c[6476]) );
XNOR U32384 ( .A(a[6476]), .B(c6476), .Z(n19430) );
XOR U32385 ( .A(c6477), .B(n19431), .Z(c6478) );
ANDN U32386 ( .B(n19432), .A(n19433), .Z(n19431) );
XOR U32387 ( .A(c6477), .B(b[6477]), .Z(n19432) );
XNOR U32388 ( .A(b[6477]), .B(n19433), .Z(c[6477]) );
XNOR U32389 ( .A(a[6477]), .B(c6477), .Z(n19433) );
XOR U32390 ( .A(c6478), .B(n19434), .Z(c6479) );
ANDN U32391 ( .B(n19435), .A(n19436), .Z(n19434) );
XOR U32392 ( .A(c6478), .B(b[6478]), .Z(n19435) );
XNOR U32393 ( .A(b[6478]), .B(n19436), .Z(c[6478]) );
XNOR U32394 ( .A(a[6478]), .B(c6478), .Z(n19436) );
XOR U32395 ( .A(c6479), .B(n19437), .Z(c6480) );
ANDN U32396 ( .B(n19438), .A(n19439), .Z(n19437) );
XOR U32397 ( .A(c6479), .B(b[6479]), .Z(n19438) );
XNOR U32398 ( .A(b[6479]), .B(n19439), .Z(c[6479]) );
XNOR U32399 ( .A(a[6479]), .B(c6479), .Z(n19439) );
XOR U32400 ( .A(c6480), .B(n19440), .Z(c6481) );
ANDN U32401 ( .B(n19441), .A(n19442), .Z(n19440) );
XOR U32402 ( .A(c6480), .B(b[6480]), .Z(n19441) );
XNOR U32403 ( .A(b[6480]), .B(n19442), .Z(c[6480]) );
XNOR U32404 ( .A(a[6480]), .B(c6480), .Z(n19442) );
XOR U32405 ( .A(c6481), .B(n19443), .Z(c6482) );
ANDN U32406 ( .B(n19444), .A(n19445), .Z(n19443) );
XOR U32407 ( .A(c6481), .B(b[6481]), .Z(n19444) );
XNOR U32408 ( .A(b[6481]), .B(n19445), .Z(c[6481]) );
XNOR U32409 ( .A(a[6481]), .B(c6481), .Z(n19445) );
XOR U32410 ( .A(c6482), .B(n19446), .Z(c6483) );
ANDN U32411 ( .B(n19447), .A(n19448), .Z(n19446) );
XOR U32412 ( .A(c6482), .B(b[6482]), .Z(n19447) );
XNOR U32413 ( .A(b[6482]), .B(n19448), .Z(c[6482]) );
XNOR U32414 ( .A(a[6482]), .B(c6482), .Z(n19448) );
XOR U32415 ( .A(c6483), .B(n19449), .Z(c6484) );
ANDN U32416 ( .B(n19450), .A(n19451), .Z(n19449) );
XOR U32417 ( .A(c6483), .B(b[6483]), .Z(n19450) );
XNOR U32418 ( .A(b[6483]), .B(n19451), .Z(c[6483]) );
XNOR U32419 ( .A(a[6483]), .B(c6483), .Z(n19451) );
XOR U32420 ( .A(c6484), .B(n19452), .Z(c6485) );
ANDN U32421 ( .B(n19453), .A(n19454), .Z(n19452) );
XOR U32422 ( .A(c6484), .B(b[6484]), .Z(n19453) );
XNOR U32423 ( .A(b[6484]), .B(n19454), .Z(c[6484]) );
XNOR U32424 ( .A(a[6484]), .B(c6484), .Z(n19454) );
XOR U32425 ( .A(c6485), .B(n19455), .Z(c6486) );
ANDN U32426 ( .B(n19456), .A(n19457), .Z(n19455) );
XOR U32427 ( .A(c6485), .B(b[6485]), .Z(n19456) );
XNOR U32428 ( .A(b[6485]), .B(n19457), .Z(c[6485]) );
XNOR U32429 ( .A(a[6485]), .B(c6485), .Z(n19457) );
XOR U32430 ( .A(c6486), .B(n19458), .Z(c6487) );
ANDN U32431 ( .B(n19459), .A(n19460), .Z(n19458) );
XOR U32432 ( .A(c6486), .B(b[6486]), .Z(n19459) );
XNOR U32433 ( .A(b[6486]), .B(n19460), .Z(c[6486]) );
XNOR U32434 ( .A(a[6486]), .B(c6486), .Z(n19460) );
XOR U32435 ( .A(c6487), .B(n19461), .Z(c6488) );
ANDN U32436 ( .B(n19462), .A(n19463), .Z(n19461) );
XOR U32437 ( .A(c6487), .B(b[6487]), .Z(n19462) );
XNOR U32438 ( .A(b[6487]), .B(n19463), .Z(c[6487]) );
XNOR U32439 ( .A(a[6487]), .B(c6487), .Z(n19463) );
XOR U32440 ( .A(c6488), .B(n19464), .Z(c6489) );
ANDN U32441 ( .B(n19465), .A(n19466), .Z(n19464) );
XOR U32442 ( .A(c6488), .B(b[6488]), .Z(n19465) );
XNOR U32443 ( .A(b[6488]), .B(n19466), .Z(c[6488]) );
XNOR U32444 ( .A(a[6488]), .B(c6488), .Z(n19466) );
XOR U32445 ( .A(c6489), .B(n19467), .Z(c6490) );
ANDN U32446 ( .B(n19468), .A(n19469), .Z(n19467) );
XOR U32447 ( .A(c6489), .B(b[6489]), .Z(n19468) );
XNOR U32448 ( .A(b[6489]), .B(n19469), .Z(c[6489]) );
XNOR U32449 ( .A(a[6489]), .B(c6489), .Z(n19469) );
XOR U32450 ( .A(c6490), .B(n19470), .Z(c6491) );
ANDN U32451 ( .B(n19471), .A(n19472), .Z(n19470) );
XOR U32452 ( .A(c6490), .B(b[6490]), .Z(n19471) );
XNOR U32453 ( .A(b[6490]), .B(n19472), .Z(c[6490]) );
XNOR U32454 ( .A(a[6490]), .B(c6490), .Z(n19472) );
XOR U32455 ( .A(c6491), .B(n19473), .Z(c6492) );
ANDN U32456 ( .B(n19474), .A(n19475), .Z(n19473) );
XOR U32457 ( .A(c6491), .B(b[6491]), .Z(n19474) );
XNOR U32458 ( .A(b[6491]), .B(n19475), .Z(c[6491]) );
XNOR U32459 ( .A(a[6491]), .B(c6491), .Z(n19475) );
XOR U32460 ( .A(c6492), .B(n19476), .Z(c6493) );
ANDN U32461 ( .B(n19477), .A(n19478), .Z(n19476) );
XOR U32462 ( .A(c6492), .B(b[6492]), .Z(n19477) );
XNOR U32463 ( .A(b[6492]), .B(n19478), .Z(c[6492]) );
XNOR U32464 ( .A(a[6492]), .B(c6492), .Z(n19478) );
XOR U32465 ( .A(c6493), .B(n19479), .Z(c6494) );
ANDN U32466 ( .B(n19480), .A(n19481), .Z(n19479) );
XOR U32467 ( .A(c6493), .B(b[6493]), .Z(n19480) );
XNOR U32468 ( .A(b[6493]), .B(n19481), .Z(c[6493]) );
XNOR U32469 ( .A(a[6493]), .B(c6493), .Z(n19481) );
XOR U32470 ( .A(c6494), .B(n19482), .Z(c6495) );
ANDN U32471 ( .B(n19483), .A(n19484), .Z(n19482) );
XOR U32472 ( .A(c6494), .B(b[6494]), .Z(n19483) );
XNOR U32473 ( .A(b[6494]), .B(n19484), .Z(c[6494]) );
XNOR U32474 ( .A(a[6494]), .B(c6494), .Z(n19484) );
XOR U32475 ( .A(c6495), .B(n19485), .Z(c6496) );
ANDN U32476 ( .B(n19486), .A(n19487), .Z(n19485) );
XOR U32477 ( .A(c6495), .B(b[6495]), .Z(n19486) );
XNOR U32478 ( .A(b[6495]), .B(n19487), .Z(c[6495]) );
XNOR U32479 ( .A(a[6495]), .B(c6495), .Z(n19487) );
XOR U32480 ( .A(c6496), .B(n19488), .Z(c6497) );
ANDN U32481 ( .B(n19489), .A(n19490), .Z(n19488) );
XOR U32482 ( .A(c6496), .B(b[6496]), .Z(n19489) );
XNOR U32483 ( .A(b[6496]), .B(n19490), .Z(c[6496]) );
XNOR U32484 ( .A(a[6496]), .B(c6496), .Z(n19490) );
XOR U32485 ( .A(c6497), .B(n19491), .Z(c6498) );
ANDN U32486 ( .B(n19492), .A(n19493), .Z(n19491) );
XOR U32487 ( .A(c6497), .B(b[6497]), .Z(n19492) );
XNOR U32488 ( .A(b[6497]), .B(n19493), .Z(c[6497]) );
XNOR U32489 ( .A(a[6497]), .B(c6497), .Z(n19493) );
XOR U32490 ( .A(c6498), .B(n19494), .Z(c6499) );
ANDN U32491 ( .B(n19495), .A(n19496), .Z(n19494) );
XOR U32492 ( .A(c6498), .B(b[6498]), .Z(n19495) );
XNOR U32493 ( .A(b[6498]), .B(n19496), .Z(c[6498]) );
XNOR U32494 ( .A(a[6498]), .B(c6498), .Z(n19496) );
XOR U32495 ( .A(c6499), .B(n19497), .Z(c6500) );
ANDN U32496 ( .B(n19498), .A(n19499), .Z(n19497) );
XOR U32497 ( .A(c6499), .B(b[6499]), .Z(n19498) );
XNOR U32498 ( .A(b[6499]), .B(n19499), .Z(c[6499]) );
XNOR U32499 ( .A(a[6499]), .B(c6499), .Z(n19499) );
XOR U32500 ( .A(c6500), .B(n19500), .Z(c6501) );
ANDN U32501 ( .B(n19501), .A(n19502), .Z(n19500) );
XOR U32502 ( .A(c6500), .B(b[6500]), .Z(n19501) );
XNOR U32503 ( .A(b[6500]), .B(n19502), .Z(c[6500]) );
XNOR U32504 ( .A(a[6500]), .B(c6500), .Z(n19502) );
XOR U32505 ( .A(c6501), .B(n19503), .Z(c6502) );
ANDN U32506 ( .B(n19504), .A(n19505), .Z(n19503) );
XOR U32507 ( .A(c6501), .B(b[6501]), .Z(n19504) );
XNOR U32508 ( .A(b[6501]), .B(n19505), .Z(c[6501]) );
XNOR U32509 ( .A(a[6501]), .B(c6501), .Z(n19505) );
XOR U32510 ( .A(c6502), .B(n19506), .Z(c6503) );
ANDN U32511 ( .B(n19507), .A(n19508), .Z(n19506) );
XOR U32512 ( .A(c6502), .B(b[6502]), .Z(n19507) );
XNOR U32513 ( .A(b[6502]), .B(n19508), .Z(c[6502]) );
XNOR U32514 ( .A(a[6502]), .B(c6502), .Z(n19508) );
XOR U32515 ( .A(c6503), .B(n19509), .Z(c6504) );
ANDN U32516 ( .B(n19510), .A(n19511), .Z(n19509) );
XOR U32517 ( .A(c6503), .B(b[6503]), .Z(n19510) );
XNOR U32518 ( .A(b[6503]), .B(n19511), .Z(c[6503]) );
XNOR U32519 ( .A(a[6503]), .B(c6503), .Z(n19511) );
XOR U32520 ( .A(c6504), .B(n19512), .Z(c6505) );
ANDN U32521 ( .B(n19513), .A(n19514), .Z(n19512) );
XOR U32522 ( .A(c6504), .B(b[6504]), .Z(n19513) );
XNOR U32523 ( .A(b[6504]), .B(n19514), .Z(c[6504]) );
XNOR U32524 ( .A(a[6504]), .B(c6504), .Z(n19514) );
XOR U32525 ( .A(c6505), .B(n19515), .Z(c6506) );
ANDN U32526 ( .B(n19516), .A(n19517), .Z(n19515) );
XOR U32527 ( .A(c6505), .B(b[6505]), .Z(n19516) );
XNOR U32528 ( .A(b[6505]), .B(n19517), .Z(c[6505]) );
XNOR U32529 ( .A(a[6505]), .B(c6505), .Z(n19517) );
XOR U32530 ( .A(c6506), .B(n19518), .Z(c6507) );
ANDN U32531 ( .B(n19519), .A(n19520), .Z(n19518) );
XOR U32532 ( .A(c6506), .B(b[6506]), .Z(n19519) );
XNOR U32533 ( .A(b[6506]), .B(n19520), .Z(c[6506]) );
XNOR U32534 ( .A(a[6506]), .B(c6506), .Z(n19520) );
XOR U32535 ( .A(c6507), .B(n19521), .Z(c6508) );
ANDN U32536 ( .B(n19522), .A(n19523), .Z(n19521) );
XOR U32537 ( .A(c6507), .B(b[6507]), .Z(n19522) );
XNOR U32538 ( .A(b[6507]), .B(n19523), .Z(c[6507]) );
XNOR U32539 ( .A(a[6507]), .B(c6507), .Z(n19523) );
XOR U32540 ( .A(c6508), .B(n19524), .Z(c6509) );
ANDN U32541 ( .B(n19525), .A(n19526), .Z(n19524) );
XOR U32542 ( .A(c6508), .B(b[6508]), .Z(n19525) );
XNOR U32543 ( .A(b[6508]), .B(n19526), .Z(c[6508]) );
XNOR U32544 ( .A(a[6508]), .B(c6508), .Z(n19526) );
XOR U32545 ( .A(c6509), .B(n19527), .Z(c6510) );
ANDN U32546 ( .B(n19528), .A(n19529), .Z(n19527) );
XOR U32547 ( .A(c6509), .B(b[6509]), .Z(n19528) );
XNOR U32548 ( .A(b[6509]), .B(n19529), .Z(c[6509]) );
XNOR U32549 ( .A(a[6509]), .B(c6509), .Z(n19529) );
XOR U32550 ( .A(c6510), .B(n19530), .Z(c6511) );
ANDN U32551 ( .B(n19531), .A(n19532), .Z(n19530) );
XOR U32552 ( .A(c6510), .B(b[6510]), .Z(n19531) );
XNOR U32553 ( .A(b[6510]), .B(n19532), .Z(c[6510]) );
XNOR U32554 ( .A(a[6510]), .B(c6510), .Z(n19532) );
XOR U32555 ( .A(c6511), .B(n19533), .Z(c6512) );
ANDN U32556 ( .B(n19534), .A(n19535), .Z(n19533) );
XOR U32557 ( .A(c6511), .B(b[6511]), .Z(n19534) );
XNOR U32558 ( .A(b[6511]), .B(n19535), .Z(c[6511]) );
XNOR U32559 ( .A(a[6511]), .B(c6511), .Z(n19535) );
XOR U32560 ( .A(c6512), .B(n19536), .Z(c6513) );
ANDN U32561 ( .B(n19537), .A(n19538), .Z(n19536) );
XOR U32562 ( .A(c6512), .B(b[6512]), .Z(n19537) );
XNOR U32563 ( .A(b[6512]), .B(n19538), .Z(c[6512]) );
XNOR U32564 ( .A(a[6512]), .B(c6512), .Z(n19538) );
XOR U32565 ( .A(c6513), .B(n19539), .Z(c6514) );
ANDN U32566 ( .B(n19540), .A(n19541), .Z(n19539) );
XOR U32567 ( .A(c6513), .B(b[6513]), .Z(n19540) );
XNOR U32568 ( .A(b[6513]), .B(n19541), .Z(c[6513]) );
XNOR U32569 ( .A(a[6513]), .B(c6513), .Z(n19541) );
XOR U32570 ( .A(c6514), .B(n19542), .Z(c6515) );
ANDN U32571 ( .B(n19543), .A(n19544), .Z(n19542) );
XOR U32572 ( .A(c6514), .B(b[6514]), .Z(n19543) );
XNOR U32573 ( .A(b[6514]), .B(n19544), .Z(c[6514]) );
XNOR U32574 ( .A(a[6514]), .B(c6514), .Z(n19544) );
XOR U32575 ( .A(c6515), .B(n19545), .Z(c6516) );
ANDN U32576 ( .B(n19546), .A(n19547), .Z(n19545) );
XOR U32577 ( .A(c6515), .B(b[6515]), .Z(n19546) );
XNOR U32578 ( .A(b[6515]), .B(n19547), .Z(c[6515]) );
XNOR U32579 ( .A(a[6515]), .B(c6515), .Z(n19547) );
XOR U32580 ( .A(c6516), .B(n19548), .Z(c6517) );
ANDN U32581 ( .B(n19549), .A(n19550), .Z(n19548) );
XOR U32582 ( .A(c6516), .B(b[6516]), .Z(n19549) );
XNOR U32583 ( .A(b[6516]), .B(n19550), .Z(c[6516]) );
XNOR U32584 ( .A(a[6516]), .B(c6516), .Z(n19550) );
XOR U32585 ( .A(c6517), .B(n19551), .Z(c6518) );
ANDN U32586 ( .B(n19552), .A(n19553), .Z(n19551) );
XOR U32587 ( .A(c6517), .B(b[6517]), .Z(n19552) );
XNOR U32588 ( .A(b[6517]), .B(n19553), .Z(c[6517]) );
XNOR U32589 ( .A(a[6517]), .B(c6517), .Z(n19553) );
XOR U32590 ( .A(c6518), .B(n19554), .Z(c6519) );
ANDN U32591 ( .B(n19555), .A(n19556), .Z(n19554) );
XOR U32592 ( .A(c6518), .B(b[6518]), .Z(n19555) );
XNOR U32593 ( .A(b[6518]), .B(n19556), .Z(c[6518]) );
XNOR U32594 ( .A(a[6518]), .B(c6518), .Z(n19556) );
XOR U32595 ( .A(c6519), .B(n19557), .Z(c6520) );
ANDN U32596 ( .B(n19558), .A(n19559), .Z(n19557) );
XOR U32597 ( .A(c6519), .B(b[6519]), .Z(n19558) );
XNOR U32598 ( .A(b[6519]), .B(n19559), .Z(c[6519]) );
XNOR U32599 ( .A(a[6519]), .B(c6519), .Z(n19559) );
XOR U32600 ( .A(c6520), .B(n19560), .Z(c6521) );
ANDN U32601 ( .B(n19561), .A(n19562), .Z(n19560) );
XOR U32602 ( .A(c6520), .B(b[6520]), .Z(n19561) );
XNOR U32603 ( .A(b[6520]), .B(n19562), .Z(c[6520]) );
XNOR U32604 ( .A(a[6520]), .B(c6520), .Z(n19562) );
XOR U32605 ( .A(c6521), .B(n19563), .Z(c6522) );
ANDN U32606 ( .B(n19564), .A(n19565), .Z(n19563) );
XOR U32607 ( .A(c6521), .B(b[6521]), .Z(n19564) );
XNOR U32608 ( .A(b[6521]), .B(n19565), .Z(c[6521]) );
XNOR U32609 ( .A(a[6521]), .B(c6521), .Z(n19565) );
XOR U32610 ( .A(c6522), .B(n19566), .Z(c6523) );
ANDN U32611 ( .B(n19567), .A(n19568), .Z(n19566) );
XOR U32612 ( .A(c6522), .B(b[6522]), .Z(n19567) );
XNOR U32613 ( .A(b[6522]), .B(n19568), .Z(c[6522]) );
XNOR U32614 ( .A(a[6522]), .B(c6522), .Z(n19568) );
XOR U32615 ( .A(c6523), .B(n19569), .Z(c6524) );
ANDN U32616 ( .B(n19570), .A(n19571), .Z(n19569) );
XOR U32617 ( .A(c6523), .B(b[6523]), .Z(n19570) );
XNOR U32618 ( .A(b[6523]), .B(n19571), .Z(c[6523]) );
XNOR U32619 ( .A(a[6523]), .B(c6523), .Z(n19571) );
XOR U32620 ( .A(c6524), .B(n19572), .Z(c6525) );
ANDN U32621 ( .B(n19573), .A(n19574), .Z(n19572) );
XOR U32622 ( .A(c6524), .B(b[6524]), .Z(n19573) );
XNOR U32623 ( .A(b[6524]), .B(n19574), .Z(c[6524]) );
XNOR U32624 ( .A(a[6524]), .B(c6524), .Z(n19574) );
XOR U32625 ( .A(c6525), .B(n19575), .Z(c6526) );
ANDN U32626 ( .B(n19576), .A(n19577), .Z(n19575) );
XOR U32627 ( .A(c6525), .B(b[6525]), .Z(n19576) );
XNOR U32628 ( .A(b[6525]), .B(n19577), .Z(c[6525]) );
XNOR U32629 ( .A(a[6525]), .B(c6525), .Z(n19577) );
XOR U32630 ( .A(c6526), .B(n19578), .Z(c6527) );
ANDN U32631 ( .B(n19579), .A(n19580), .Z(n19578) );
XOR U32632 ( .A(c6526), .B(b[6526]), .Z(n19579) );
XNOR U32633 ( .A(b[6526]), .B(n19580), .Z(c[6526]) );
XNOR U32634 ( .A(a[6526]), .B(c6526), .Z(n19580) );
XOR U32635 ( .A(c6527), .B(n19581), .Z(c6528) );
ANDN U32636 ( .B(n19582), .A(n19583), .Z(n19581) );
XOR U32637 ( .A(c6527), .B(b[6527]), .Z(n19582) );
XNOR U32638 ( .A(b[6527]), .B(n19583), .Z(c[6527]) );
XNOR U32639 ( .A(a[6527]), .B(c6527), .Z(n19583) );
XOR U32640 ( .A(c6528), .B(n19584), .Z(c6529) );
ANDN U32641 ( .B(n19585), .A(n19586), .Z(n19584) );
XOR U32642 ( .A(c6528), .B(b[6528]), .Z(n19585) );
XNOR U32643 ( .A(b[6528]), .B(n19586), .Z(c[6528]) );
XNOR U32644 ( .A(a[6528]), .B(c6528), .Z(n19586) );
XOR U32645 ( .A(c6529), .B(n19587), .Z(c6530) );
ANDN U32646 ( .B(n19588), .A(n19589), .Z(n19587) );
XOR U32647 ( .A(c6529), .B(b[6529]), .Z(n19588) );
XNOR U32648 ( .A(b[6529]), .B(n19589), .Z(c[6529]) );
XNOR U32649 ( .A(a[6529]), .B(c6529), .Z(n19589) );
XOR U32650 ( .A(c6530), .B(n19590), .Z(c6531) );
ANDN U32651 ( .B(n19591), .A(n19592), .Z(n19590) );
XOR U32652 ( .A(c6530), .B(b[6530]), .Z(n19591) );
XNOR U32653 ( .A(b[6530]), .B(n19592), .Z(c[6530]) );
XNOR U32654 ( .A(a[6530]), .B(c6530), .Z(n19592) );
XOR U32655 ( .A(c6531), .B(n19593), .Z(c6532) );
ANDN U32656 ( .B(n19594), .A(n19595), .Z(n19593) );
XOR U32657 ( .A(c6531), .B(b[6531]), .Z(n19594) );
XNOR U32658 ( .A(b[6531]), .B(n19595), .Z(c[6531]) );
XNOR U32659 ( .A(a[6531]), .B(c6531), .Z(n19595) );
XOR U32660 ( .A(c6532), .B(n19596), .Z(c6533) );
ANDN U32661 ( .B(n19597), .A(n19598), .Z(n19596) );
XOR U32662 ( .A(c6532), .B(b[6532]), .Z(n19597) );
XNOR U32663 ( .A(b[6532]), .B(n19598), .Z(c[6532]) );
XNOR U32664 ( .A(a[6532]), .B(c6532), .Z(n19598) );
XOR U32665 ( .A(c6533), .B(n19599), .Z(c6534) );
ANDN U32666 ( .B(n19600), .A(n19601), .Z(n19599) );
XOR U32667 ( .A(c6533), .B(b[6533]), .Z(n19600) );
XNOR U32668 ( .A(b[6533]), .B(n19601), .Z(c[6533]) );
XNOR U32669 ( .A(a[6533]), .B(c6533), .Z(n19601) );
XOR U32670 ( .A(c6534), .B(n19602), .Z(c6535) );
ANDN U32671 ( .B(n19603), .A(n19604), .Z(n19602) );
XOR U32672 ( .A(c6534), .B(b[6534]), .Z(n19603) );
XNOR U32673 ( .A(b[6534]), .B(n19604), .Z(c[6534]) );
XNOR U32674 ( .A(a[6534]), .B(c6534), .Z(n19604) );
XOR U32675 ( .A(c6535), .B(n19605), .Z(c6536) );
ANDN U32676 ( .B(n19606), .A(n19607), .Z(n19605) );
XOR U32677 ( .A(c6535), .B(b[6535]), .Z(n19606) );
XNOR U32678 ( .A(b[6535]), .B(n19607), .Z(c[6535]) );
XNOR U32679 ( .A(a[6535]), .B(c6535), .Z(n19607) );
XOR U32680 ( .A(c6536), .B(n19608), .Z(c6537) );
ANDN U32681 ( .B(n19609), .A(n19610), .Z(n19608) );
XOR U32682 ( .A(c6536), .B(b[6536]), .Z(n19609) );
XNOR U32683 ( .A(b[6536]), .B(n19610), .Z(c[6536]) );
XNOR U32684 ( .A(a[6536]), .B(c6536), .Z(n19610) );
XOR U32685 ( .A(c6537), .B(n19611), .Z(c6538) );
ANDN U32686 ( .B(n19612), .A(n19613), .Z(n19611) );
XOR U32687 ( .A(c6537), .B(b[6537]), .Z(n19612) );
XNOR U32688 ( .A(b[6537]), .B(n19613), .Z(c[6537]) );
XNOR U32689 ( .A(a[6537]), .B(c6537), .Z(n19613) );
XOR U32690 ( .A(c6538), .B(n19614), .Z(c6539) );
ANDN U32691 ( .B(n19615), .A(n19616), .Z(n19614) );
XOR U32692 ( .A(c6538), .B(b[6538]), .Z(n19615) );
XNOR U32693 ( .A(b[6538]), .B(n19616), .Z(c[6538]) );
XNOR U32694 ( .A(a[6538]), .B(c6538), .Z(n19616) );
XOR U32695 ( .A(c6539), .B(n19617), .Z(c6540) );
ANDN U32696 ( .B(n19618), .A(n19619), .Z(n19617) );
XOR U32697 ( .A(c6539), .B(b[6539]), .Z(n19618) );
XNOR U32698 ( .A(b[6539]), .B(n19619), .Z(c[6539]) );
XNOR U32699 ( .A(a[6539]), .B(c6539), .Z(n19619) );
XOR U32700 ( .A(c6540), .B(n19620), .Z(c6541) );
ANDN U32701 ( .B(n19621), .A(n19622), .Z(n19620) );
XOR U32702 ( .A(c6540), .B(b[6540]), .Z(n19621) );
XNOR U32703 ( .A(b[6540]), .B(n19622), .Z(c[6540]) );
XNOR U32704 ( .A(a[6540]), .B(c6540), .Z(n19622) );
XOR U32705 ( .A(c6541), .B(n19623), .Z(c6542) );
ANDN U32706 ( .B(n19624), .A(n19625), .Z(n19623) );
XOR U32707 ( .A(c6541), .B(b[6541]), .Z(n19624) );
XNOR U32708 ( .A(b[6541]), .B(n19625), .Z(c[6541]) );
XNOR U32709 ( .A(a[6541]), .B(c6541), .Z(n19625) );
XOR U32710 ( .A(c6542), .B(n19626), .Z(c6543) );
ANDN U32711 ( .B(n19627), .A(n19628), .Z(n19626) );
XOR U32712 ( .A(c6542), .B(b[6542]), .Z(n19627) );
XNOR U32713 ( .A(b[6542]), .B(n19628), .Z(c[6542]) );
XNOR U32714 ( .A(a[6542]), .B(c6542), .Z(n19628) );
XOR U32715 ( .A(c6543), .B(n19629), .Z(c6544) );
ANDN U32716 ( .B(n19630), .A(n19631), .Z(n19629) );
XOR U32717 ( .A(c6543), .B(b[6543]), .Z(n19630) );
XNOR U32718 ( .A(b[6543]), .B(n19631), .Z(c[6543]) );
XNOR U32719 ( .A(a[6543]), .B(c6543), .Z(n19631) );
XOR U32720 ( .A(c6544), .B(n19632), .Z(c6545) );
ANDN U32721 ( .B(n19633), .A(n19634), .Z(n19632) );
XOR U32722 ( .A(c6544), .B(b[6544]), .Z(n19633) );
XNOR U32723 ( .A(b[6544]), .B(n19634), .Z(c[6544]) );
XNOR U32724 ( .A(a[6544]), .B(c6544), .Z(n19634) );
XOR U32725 ( .A(c6545), .B(n19635), .Z(c6546) );
ANDN U32726 ( .B(n19636), .A(n19637), .Z(n19635) );
XOR U32727 ( .A(c6545), .B(b[6545]), .Z(n19636) );
XNOR U32728 ( .A(b[6545]), .B(n19637), .Z(c[6545]) );
XNOR U32729 ( .A(a[6545]), .B(c6545), .Z(n19637) );
XOR U32730 ( .A(c6546), .B(n19638), .Z(c6547) );
ANDN U32731 ( .B(n19639), .A(n19640), .Z(n19638) );
XOR U32732 ( .A(c6546), .B(b[6546]), .Z(n19639) );
XNOR U32733 ( .A(b[6546]), .B(n19640), .Z(c[6546]) );
XNOR U32734 ( .A(a[6546]), .B(c6546), .Z(n19640) );
XOR U32735 ( .A(c6547), .B(n19641), .Z(c6548) );
ANDN U32736 ( .B(n19642), .A(n19643), .Z(n19641) );
XOR U32737 ( .A(c6547), .B(b[6547]), .Z(n19642) );
XNOR U32738 ( .A(b[6547]), .B(n19643), .Z(c[6547]) );
XNOR U32739 ( .A(a[6547]), .B(c6547), .Z(n19643) );
XOR U32740 ( .A(c6548), .B(n19644), .Z(c6549) );
ANDN U32741 ( .B(n19645), .A(n19646), .Z(n19644) );
XOR U32742 ( .A(c6548), .B(b[6548]), .Z(n19645) );
XNOR U32743 ( .A(b[6548]), .B(n19646), .Z(c[6548]) );
XNOR U32744 ( .A(a[6548]), .B(c6548), .Z(n19646) );
XOR U32745 ( .A(c6549), .B(n19647), .Z(c6550) );
ANDN U32746 ( .B(n19648), .A(n19649), .Z(n19647) );
XOR U32747 ( .A(c6549), .B(b[6549]), .Z(n19648) );
XNOR U32748 ( .A(b[6549]), .B(n19649), .Z(c[6549]) );
XNOR U32749 ( .A(a[6549]), .B(c6549), .Z(n19649) );
XOR U32750 ( .A(c6550), .B(n19650), .Z(c6551) );
ANDN U32751 ( .B(n19651), .A(n19652), .Z(n19650) );
XOR U32752 ( .A(c6550), .B(b[6550]), .Z(n19651) );
XNOR U32753 ( .A(b[6550]), .B(n19652), .Z(c[6550]) );
XNOR U32754 ( .A(a[6550]), .B(c6550), .Z(n19652) );
XOR U32755 ( .A(c6551), .B(n19653), .Z(c6552) );
ANDN U32756 ( .B(n19654), .A(n19655), .Z(n19653) );
XOR U32757 ( .A(c6551), .B(b[6551]), .Z(n19654) );
XNOR U32758 ( .A(b[6551]), .B(n19655), .Z(c[6551]) );
XNOR U32759 ( .A(a[6551]), .B(c6551), .Z(n19655) );
XOR U32760 ( .A(c6552), .B(n19656), .Z(c6553) );
ANDN U32761 ( .B(n19657), .A(n19658), .Z(n19656) );
XOR U32762 ( .A(c6552), .B(b[6552]), .Z(n19657) );
XNOR U32763 ( .A(b[6552]), .B(n19658), .Z(c[6552]) );
XNOR U32764 ( .A(a[6552]), .B(c6552), .Z(n19658) );
XOR U32765 ( .A(c6553), .B(n19659), .Z(c6554) );
ANDN U32766 ( .B(n19660), .A(n19661), .Z(n19659) );
XOR U32767 ( .A(c6553), .B(b[6553]), .Z(n19660) );
XNOR U32768 ( .A(b[6553]), .B(n19661), .Z(c[6553]) );
XNOR U32769 ( .A(a[6553]), .B(c6553), .Z(n19661) );
XOR U32770 ( .A(c6554), .B(n19662), .Z(c6555) );
ANDN U32771 ( .B(n19663), .A(n19664), .Z(n19662) );
XOR U32772 ( .A(c6554), .B(b[6554]), .Z(n19663) );
XNOR U32773 ( .A(b[6554]), .B(n19664), .Z(c[6554]) );
XNOR U32774 ( .A(a[6554]), .B(c6554), .Z(n19664) );
XOR U32775 ( .A(c6555), .B(n19665), .Z(c6556) );
ANDN U32776 ( .B(n19666), .A(n19667), .Z(n19665) );
XOR U32777 ( .A(c6555), .B(b[6555]), .Z(n19666) );
XNOR U32778 ( .A(b[6555]), .B(n19667), .Z(c[6555]) );
XNOR U32779 ( .A(a[6555]), .B(c6555), .Z(n19667) );
XOR U32780 ( .A(c6556), .B(n19668), .Z(c6557) );
ANDN U32781 ( .B(n19669), .A(n19670), .Z(n19668) );
XOR U32782 ( .A(c6556), .B(b[6556]), .Z(n19669) );
XNOR U32783 ( .A(b[6556]), .B(n19670), .Z(c[6556]) );
XNOR U32784 ( .A(a[6556]), .B(c6556), .Z(n19670) );
XOR U32785 ( .A(c6557), .B(n19671), .Z(c6558) );
ANDN U32786 ( .B(n19672), .A(n19673), .Z(n19671) );
XOR U32787 ( .A(c6557), .B(b[6557]), .Z(n19672) );
XNOR U32788 ( .A(b[6557]), .B(n19673), .Z(c[6557]) );
XNOR U32789 ( .A(a[6557]), .B(c6557), .Z(n19673) );
XOR U32790 ( .A(c6558), .B(n19674), .Z(c6559) );
ANDN U32791 ( .B(n19675), .A(n19676), .Z(n19674) );
XOR U32792 ( .A(c6558), .B(b[6558]), .Z(n19675) );
XNOR U32793 ( .A(b[6558]), .B(n19676), .Z(c[6558]) );
XNOR U32794 ( .A(a[6558]), .B(c6558), .Z(n19676) );
XOR U32795 ( .A(c6559), .B(n19677), .Z(c6560) );
ANDN U32796 ( .B(n19678), .A(n19679), .Z(n19677) );
XOR U32797 ( .A(c6559), .B(b[6559]), .Z(n19678) );
XNOR U32798 ( .A(b[6559]), .B(n19679), .Z(c[6559]) );
XNOR U32799 ( .A(a[6559]), .B(c6559), .Z(n19679) );
XOR U32800 ( .A(c6560), .B(n19680), .Z(c6561) );
ANDN U32801 ( .B(n19681), .A(n19682), .Z(n19680) );
XOR U32802 ( .A(c6560), .B(b[6560]), .Z(n19681) );
XNOR U32803 ( .A(b[6560]), .B(n19682), .Z(c[6560]) );
XNOR U32804 ( .A(a[6560]), .B(c6560), .Z(n19682) );
XOR U32805 ( .A(c6561), .B(n19683), .Z(c6562) );
ANDN U32806 ( .B(n19684), .A(n19685), .Z(n19683) );
XOR U32807 ( .A(c6561), .B(b[6561]), .Z(n19684) );
XNOR U32808 ( .A(b[6561]), .B(n19685), .Z(c[6561]) );
XNOR U32809 ( .A(a[6561]), .B(c6561), .Z(n19685) );
XOR U32810 ( .A(c6562), .B(n19686), .Z(c6563) );
ANDN U32811 ( .B(n19687), .A(n19688), .Z(n19686) );
XOR U32812 ( .A(c6562), .B(b[6562]), .Z(n19687) );
XNOR U32813 ( .A(b[6562]), .B(n19688), .Z(c[6562]) );
XNOR U32814 ( .A(a[6562]), .B(c6562), .Z(n19688) );
XOR U32815 ( .A(c6563), .B(n19689), .Z(c6564) );
ANDN U32816 ( .B(n19690), .A(n19691), .Z(n19689) );
XOR U32817 ( .A(c6563), .B(b[6563]), .Z(n19690) );
XNOR U32818 ( .A(b[6563]), .B(n19691), .Z(c[6563]) );
XNOR U32819 ( .A(a[6563]), .B(c6563), .Z(n19691) );
XOR U32820 ( .A(c6564), .B(n19692), .Z(c6565) );
ANDN U32821 ( .B(n19693), .A(n19694), .Z(n19692) );
XOR U32822 ( .A(c6564), .B(b[6564]), .Z(n19693) );
XNOR U32823 ( .A(b[6564]), .B(n19694), .Z(c[6564]) );
XNOR U32824 ( .A(a[6564]), .B(c6564), .Z(n19694) );
XOR U32825 ( .A(c6565), .B(n19695), .Z(c6566) );
ANDN U32826 ( .B(n19696), .A(n19697), .Z(n19695) );
XOR U32827 ( .A(c6565), .B(b[6565]), .Z(n19696) );
XNOR U32828 ( .A(b[6565]), .B(n19697), .Z(c[6565]) );
XNOR U32829 ( .A(a[6565]), .B(c6565), .Z(n19697) );
XOR U32830 ( .A(c6566), .B(n19698), .Z(c6567) );
ANDN U32831 ( .B(n19699), .A(n19700), .Z(n19698) );
XOR U32832 ( .A(c6566), .B(b[6566]), .Z(n19699) );
XNOR U32833 ( .A(b[6566]), .B(n19700), .Z(c[6566]) );
XNOR U32834 ( .A(a[6566]), .B(c6566), .Z(n19700) );
XOR U32835 ( .A(c6567), .B(n19701), .Z(c6568) );
ANDN U32836 ( .B(n19702), .A(n19703), .Z(n19701) );
XOR U32837 ( .A(c6567), .B(b[6567]), .Z(n19702) );
XNOR U32838 ( .A(b[6567]), .B(n19703), .Z(c[6567]) );
XNOR U32839 ( .A(a[6567]), .B(c6567), .Z(n19703) );
XOR U32840 ( .A(c6568), .B(n19704), .Z(c6569) );
ANDN U32841 ( .B(n19705), .A(n19706), .Z(n19704) );
XOR U32842 ( .A(c6568), .B(b[6568]), .Z(n19705) );
XNOR U32843 ( .A(b[6568]), .B(n19706), .Z(c[6568]) );
XNOR U32844 ( .A(a[6568]), .B(c6568), .Z(n19706) );
XOR U32845 ( .A(c6569), .B(n19707), .Z(c6570) );
ANDN U32846 ( .B(n19708), .A(n19709), .Z(n19707) );
XOR U32847 ( .A(c6569), .B(b[6569]), .Z(n19708) );
XNOR U32848 ( .A(b[6569]), .B(n19709), .Z(c[6569]) );
XNOR U32849 ( .A(a[6569]), .B(c6569), .Z(n19709) );
XOR U32850 ( .A(c6570), .B(n19710), .Z(c6571) );
ANDN U32851 ( .B(n19711), .A(n19712), .Z(n19710) );
XOR U32852 ( .A(c6570), .B(b[6570]), .Z(n19711) );
XNOR U32853 ( .A(b[6570]), .B(n19712), .Z(c[6570]) );
XNOR U32854 ( .A(a[6570]), .B(c6570), .Z(n19712) );
XOR U32855 ( .A(c6571), .B(n19713), .Z(c6572) );
ANDN U32856 ( .B(n19714), .A(n19715), .Z(n19713) );
XOR U32857 ( .A(c6571), .B(b[6571]), .Z(n19714) );
XNOR U32858 ( .A(b[6571]), .B(n19715), .Z(c[6571]) );
XNOR U32859 ( .A(a[6571]), .B(c6571), .Z(n19715) );
XOR U32860 ( .A(c6572), .B(n19716), .Z(c6573) );
ANDN U32861 ( .B(n19717), .A(n19718), .Z(n19716) );
XOR U32862 ( .A(c6572), .B(b[6572]), .Z(n19717) );
XNOR U32863 ( .A(b[6572]), .B(n19718), .Z(c[6572]) );
XNOR U32864 ( .A(a[6572]), .B(c6572), .Z(n19718) );
XOR U32865 ( .A(c6573), .B(n19719), .Z(c6574) );
ANDN U32866 ( .B(n19720), .A(n19721), .Z(n19719) );
XOR U32867 ( .A(c6573), .B(b[6573]), .Z(n19720) );
XNOR U32868 ( .A(b[6573]), .B(n19721), .Z(c[6573]) );
XNOR U32869 ( .A(a[6573]), .B(c6573), .Z(n19721) );
XOR U32870 ( .A(c6574), .B(n19722), .Z(c6575) );
ANDN U32871 ( .B(n19723), .A(n19724), .Z(n19722) );
XOR U32872 ( .A(c6574), .B(b[6574]), .Z(n19723) );
XNOR U32873 ( .A(b[6574]), .B(n19724), .Z(c[6574]) );
XNOR U32874 ( .A(a[6574]), .B(c6574), .Z(n19724) );
XOR U32875 ( .A(c6575), .B(n19725), .Z(c6576) );
ANDN U32876 ( .B(n19726), .A(n19727), .Z(n19725) );
XOR U32877 ( .A(c6575), .B(b[6575]), .Z(n19726) );
XNOR U32878 ( .A(b[6575]), .B(n19727), .Z(c[6575]) );
XNOR U32879 ( .A(a[6575]), .B(c6575), .Z(n19727) );
XOR U32880 ( .A(c6576), .B(n19728), .Z(c6577) );
ANDN U32881 ( .B(n19729), .A(n19730), .Z(n19728) );
XOR U32882 ( .A(c6576), .B(b[6576]), .Z(n19729) );
XNOR U32883 ( .A(b[6576]), .B(n19730), .Z(c[6576]) );
XNOR U32884 ( .A(a[6576]), .B(c6576), .Z(n19730) );
XOR U32885 ( .A(c6577), .B(n19731), .Z(c6578) );
ANDN U32886 ( .B(n19732), .A(n19733), .Z(n19731) );
XOR U32887 ( .A(c6577), .B(b[6577]), .Z(n19732) );
XNOR U32888 ( .A(b[6577]), .B(n19733), .Z(c[6577]) );
XNOR U32889 ( .A(a[6577]), .B(c6577), .Z(n19733) );
XOR U32890 ( .A(c6578), .B(n19734), .Z(c6579) );
ANDN U32891 ( .B(n19735), .A(n19736), .Z(n19734) );
XOR U32892 ( .A(c6578), .B(b[6578]), .Z(n19735) );
XNOR U32893 ( .A(b[6578]), .B(n19736), .Z(c[6578]) );
XNOR U32894 ( .A(a[6578]), .B(c6578), .Z(n19736) );
XOR U32895 ( .A(c6579), .B(n19737), .Z(c6580) );
ANDN U32896 ( .B(n19738), .A(n19739), .Z(n19737) );
XOR U32897 ( .A(c6579), .B(b[6579]), .Z(n19738) );
XNOR U32898 ( .A(b[6579]), .B(n19739), .Z(c[6579]) );
XNOR U32899 ( .A(a[6579]), .B(c6579), .Z(n19739) );
XOR U32900 ( .A(c6580), .B(n19740), .Z(c6581) );
ANDN U32901 ( .B(n19741), .A(n19742), .Z(n19740) );
XOR U32902 ( .A(c6580), .B(b[6580]), .Z(n19741) );
XNOR U32903 ( .A(b[6580]), .B(n19742), .Z(c[6580]) );
XNOR U32904 ( .A(a[6580]), .B(c6580), .Z(n19742) );
XOR U32905 ( .A(c6581), .B(n19743), .Z(c6582) );
ANDN U32906 ( .B(n19744), .A(n19745), .Z(n19743) );
XOR U32907 ( .A(c6581), .B(b[6581]), .Z(n19744) );
XNOR U32908 ( .A(b[6581]), .B(n19745), .Z(c[6581]) );
XNOR U32909 ( .A(a[6581]), .B(c6581), .Z(n19745) );
XOR U32910 ( .A(c6582), .B(n19746), .Z(c6583) );
ANDN U32911 ( .B(n19747), .A(n19748), .Z(n19746) );
XOR U32912 ( .A(c6582), .B(b[6582]), .Z(n19747) );
XNOR U32913 ( .A(b[6582]), .B(n19748), .Z(c[6582]) );
XNOR U32914 ( .A(a[6582]), .B(c6582), .Z(n19748) );
XOR U32915 ( .A(c6583), .B(n19749), .Z(c6584) );
ANDN U32916 ( .B(n19750), .A(n19751), .Z(n19749) );
XOR U32917 ( .A(c6583), .B(b[6583]), .Z(n19750) );
XNOR U32918 ( .A(b[6583]), .B(n19751), .Z(c[6583]) );
XNOR U32919 ( .A(a[6583]), .B(c6583), .Z(n19751) );
XOR U32920 ( .A(c6584), .B(n19752), .Z(c6585) );
ANDN U32921 ( .B(n19753), .A(n19754), .Z(n19752) );
XOR U32922 ( .A(c6584), .B(b[6584]), .Z(n19753) );
XNOR U32923 ( .A(b[6584]), .B(n19754), .Z(c[6584]) );
XNOR U32924 ( .A(a[6584]), .B(c6584), .Z(n19754) );
XOR U32925 ( .A(c6585), .B(n19755), .Z(c6586) );
ANDN U32926 ( .B(n19756), .A(n19757), .Z(n19755) );
XOR U32927 ( .A(c6585), .B(b[6585]), .Z(n19756) );
XNOR U32928 ( .A(b[6585]), .B(n19757), .Z(c[6585]) );
XNOR U32929 ( .A(a[6585]), .B(c6585), .Z(n19757) );
XOR U32930 ( .A(c6586), .B(n19758), .Z(c6587) );
ANDN U32931 ( .B(n19759), .A(n19760), .Z(n19758) );
XOR U32932 ( .A(c6586), .B(b[6586]), .Z(n19759) );
XNOR U32933 ( .A(b[6586]), .B(n19760), .Z(c[6586]) );
XNOR U32934 ( .A(a[6586]), .B(c6586), .Z(n19760) );
XOR U32935 ( .A(c6587), .B(n19761), .Z(c6588) );
ANDN U32936 ( .B(n19762), .A(n19763), .Z(n19761) );
XOR U32937 ( .A(c6587), .B(b[6587]), .Z(n19762) );
XNOR U32938 ( .A(b[6587]), .B(n19763), .Z(c[6587]) );
XNOR U32939 ( .A(a[6587]), .B(c6587), .Z(n19763) );
XOR U32940 ( .A(c6588), .B(n19764), .Z(c6589) );
ANDN U32941 ( .B(n19765), .A(n19766), .Z(n19764) );
XOR U32942 ( .A(c6588), .B(b[6588]), .Z(n19765) );
XNOR U32943 ( .A(b[6588]), .B(n19766), .Z(c[6588]) );
XNOR U32944 ( .A(a[6588]), .B(c6588), .Z(n19766) );
XOR U32945 ( .A(c6589), .B(n19767), .Z(c6590) );
ANDN U32946 ( .B(n19768), .A(n19769), .Z(n19767) );
XOR U32947 ( .A(c6589), .B(b[6589]), .Z(n19768) );
XNOR U32948 ( .A(b[6589]), .B(n19769), .Z(c[6589]) );
XNOR U32949 ( .A(a[6589]), .B(c6589), .Z(n19769) );
XOR U32950 ( .A(c6590), .B(n19770), .Z(c6591) );
ANDN U32951 ( .B(n19771), .A(n19772), .Z(n19770) );
XOR U32952 ( .A(c6590), .B(b[6590]), .Z(n19771) );
XNOR U32953 ( .A(b[6590]), .B(n19772), .Z(c[6590]) );
XNOR U32954 ( .A(a[6590]), .B(c6590), .Z(n19772) );
XOR U32955 ( .A(c6591), .B(n19773), .Z(c6592) );
ANDN U32956 ( .B(n19774), .A(n19775), .Z(n19773) );
XOR U32957 ( .A(c6591), .B(b[6591]), .Z(n19774) );
XNOR U32958 ( .A(b[6591]), .B(n19775), .Z(c[6591]) );
XNOR U32959 ( .A(a[6591]), .B(c6591), .Z(n19775) );
XOR U32960 ( .A(c6592), .B(n19776), .Z(c6593) );
ANDN U32961 ( .B(n19777), .A(n19778), .Z(n19776) );
XOR U32962 ( .A(c6592), .B(b[6592]), .Z(n19777) );
XNOR U32963 ( .A(b[6592]), .B(n19778), .Z(c[6592]) );
XNOR U32964 ( .A(a[6592]), .B(c6592), .Z(n19778) );
XOR U32965 ( .A(c6593), .B(n19779), .Z(c6594) );
ANDN U32966 ( .B(n19780), .A(n19781), .Z(n19779) );
XOR U32967 ( .A(c6593), .B(b[6593]), .Z(n19780) );
XNOR U32968 ( .A(b[6593]), .B(n19781), .Z(c[6593]) );
XNOR U32969 ( .A(a[6593]), .B(c6593), .Z(n19781) );
XOR U32970 ( .A(c6594), .B(n19782), .Z(c6595) );
ANDN U32971 ( .B(n19783), .A(n19784), .Z(n19782) );
XOR U32972 ( .A(c6594), .B(b[6594]), .Z(n19783) );
XNOR U32973 ( .A(b[6594]), .B(n19784), .Z(c[6594]) );
XNOR U32974 ( .A(a[6594]), .B(c6594), .Z(n19784) );
XOR U32975 ( .A(c6595), .B(n19785), .Z(c6596) );
ANDN U32976 ( .B(n19786), .A(n19787), .Z(n19785) );
XOR U32977 ( .A(c6595), .B(b[6595]), .Z(n19786) );
XNOR U32978 ( .A(b[6595]), .B(n19787), .Z(c[6595]) );
XNOR U32979 ( .A(a[6595]), .B(c6595), .Z(n19787) );
XOR U32980 ( .A(c6596), .B(n19788), .Z(c6597) );
ANDN U32981 ( .B(n19789), .A(n19790), .Z(n19788) );
XOR U32982 ( .A(c6596), .B(b[6596]), .Z(n19789) );
XNOR U32983 ( .A(b[6596]), .B(n19790), .Z(c[6596]) );
XNOR U32984 ( .A(a[6596]), .B(c6596), .Z(n19790) );
XOR U32985 ( .A(c6597), .B(n19791), .Z(c6598) );
ANDN U32986 ( .B(n19792), .A(n19793), .Z(n19791) );
XOR U32987 ( .A(c6597), .B(b[6597]), .Z(n19792) );
XNOR U32988 ( .A(b[6597]), .B(n19793), .Z(c[6597]) );
XNOR U32989 ( .A(a[6597]), .B(c6597), .Z(n19793) );
XOR U32990 ( .A(c6598), .B(n19794), .Z(c6599) );
ANDN U32991 ( .B(n19795), .A(n19796), .Z(n19794) );
XOR U32992 ( .A(c6598), .B(b[6598]), .Z(n19795) );
XNOR U32993 ( .A(b[6598]), .B(n19796), .Z(c[6598]) );
XNOR U32994 ( .A(a[6598]), .B(c6598), .Z(n19796) );
XOR U32995 ( .A(c6599), .B(n19797), .Z(c6600) );
ANDN U32996 ( .B(n19798), .A(n19799), .Z(n19797) );
XOR U32997 ( .A(c6599), .B(b[6599]), .Z(n19798) );
XNOR U32998 ( .A(b[6599]), .B(n19799), .Z(c[6599]) );
XNOR U32999 ( .A(a[6599]), .B(c6599), .Z(n19799) );
XOR U33000 ( .A(c6600), .B(n19800), .Z(c6601) );
ANDN U33001 ( .B(n19801), .A(n19802), .Z(n19800) );
XOR U33002 ( .A(c6600), .B(b[6600]), .Z(n19801) );
XNOR U33003 ( .A(b[6600]), .B(n19802), .Z(c[6600]) );
XNOR U33004 ( .A(a[6600]), .B(c6600), .Z(n19802) );
XOR U33005 ( .A(c6601), .B(n19803), .Z(c6602) );
ANDN U33006 ( .B(n19804), .A(n19805), .Z(n19803) );
XOR U33007 ( .A(c6601), .B(b[6601]), .Z(n19804) );
XNOR U33008 ( .A(b[6601]), .B(n19805), .Z(c[6601]) );
XNOR U33009 ( .A(a[6601]), .B(c6601), .Z(n19805) );
XOR U33010 ( .A(c6602), .B(n19806), .Z(c6603) );
ANDN U33011 ( .B(n19807), .A(n19808), .Z(n19806) );
XOR U33012 ( .A(c6602), .B(b[6602]), .Z(n19807) );
XNOR U33013 ( .A(b[6602]), .B(n19808), .Z(c[6602]) );
XNOR U33014 ( .A(a[6602]), .B(c6602), .Z(n19808) );
XOR U33015 ( .A(c6603), .B(n19809), .Z(c6604) );
ANDN U33016 ( .B(n19810), .A(n19811), .Z(n19809) );
XOR U33017 ( .A(c6603), .B(b[6603]), .Z(n19810) );
XNOR U33018 ( .A(b[6603]), .B(n19811), .Z(c[6603]) );
XNOR U33019 ( .A(a[6603]), .B(c6603), .Z(n19811) );
XOR U33020 ( .A(c6604), .B(n19812), .Z(c6605) );
ANDN U33021 ( .B(n19813), .A(n19814), .Z(n19812) );
XOR U33022 ( .A(c6604), .B(b[6604]), .Z(n19813) );
XNOR U33023 ( .A(b[6604]), .B(n19814), .Z(c[6604]) );
XNOR U33024 ( .A(a[6604]), .B(c6604), .Z(n19814) );
XOR U33025 ( .A(c6605), .B(n19815), .Z(c6606) );
ANDN U33026 ( .B(n19816), .A(n19817), .Z(n19815) );
XOR U33027 ( .A(c6605), .B(b[6605]), .Z(n19816) );
XNOR U33028 ( .A(b[6605]), .B(n19817), .Z(c[6605]) );
XNOR U33029 ( .A(a[6605]), .B(c6605), .Z(n19817) );
XOR U33030 ( .A(c6606), .B(n19818), .Z(c6607) );
ANDN U33031 ( .B(n19819), .A(n19820), .Z(n19818) );
XOR U33032 ( .A(c6606), .B(b[6606]), .Z(n19819) );
XNOR U33033 ( .A(b[6606]), .B(n19820), .Z(c[6606]) );
XNOR U33034 ( .A(a[6606]), .B(c6606), .Z(n19820) );
XOR U33035 ( .A(c6607), .B(n19821), .Z(c6608) );
ANDN U33036 ( .B(n19822), .A(n19823), .Z(n19821) );
XOR U33037 ( .A(c6607), .B(b[6607]), .Z(n19822) );
XNOR U33038 ( .A(b[6607]), .B(n19823), .Z(c[6607]) );
XNOR U33039 ( .A(a[6607]), .B(c6607), .Z(n19823) );
XOR U33040 ( .A(c6608), .B(n19824), .Z(c6609) );
ANDN U33041 ( .B(n19825), .A(n19826), .Z(n19824) );
XOR U33042 ( .A(c6608), .B(b[6608]), .Z(n19825) );
XNOR U33043 ( .A(b[6608]), .B(n19826), .Z(c[6608]) );
XNOR U33044 ( .A(a[6608]), .B(c6608), .Z(n19826) );
XOR U33045 ( .A(c6609), .B(n19827), .Z(c6610) );
ANDN U33046 ( .B(n19828), .A(n19829), .Z(n19827) );
XOR U33047 ( .A(c6609), .B(b[6609]), .Z(n19828) );
XNOR U33048 ( .A(b[6609]), .B(n19829), .Z(c[6609]) );
XNOR U33049 ( .A(a[6609]), .B(c6609), .Z(n19829) );
XOR U33050 ( .A(c6610), .B(n19830), .Z(c6611) );
ANDN U33051 ( .B(n19831), .A(n19832), .Z(n19830) );
XOR U33052 ( .A(c6610), .B(b[6610]), .Z(n19831) );
XNOR U33053 ( .A(b[6610]), .B(n19832), .Z(c[6610]) );
XNOR U33054 ( .A(a[6610]), .B(c6610), .Z(n19832) );
XOR U33055 ( .A(c6611), .B(n19833), .Z(c6612) );
ANDN U33056 ( .B(n19834), .A(n19835), .Z(n19833) );
XOR U33057 ( .A(c6611), .B(b[6611]), .Z(n19834) );
XNOR U33058 ( .A(b[6611]), .B(n19835), .Z(c[6611]) );
XNOR U33059 ( .A(a[6611]), .B(c6611), .Z(n19835) );
XOR U33060 ( .A(c6612), .B(n19836), .Z(c6613) );
ANDN U33061 ( .B(n19837), .A(n19838), .Z(n19836) );
XOR U33062 ( .A(c6612), .B(b[6612]), .Z(n19837) );
XNOR U33063 ( .A(b[6612]), .B(n19838), .Z(c[6612]) );
XNOR U33064 ( .A(a[6612]), .B(c6612), .Z(n19838) );
XOR U33065 ( .A(c6613), .B(n19839), .Z(c6614) );
ANDN U33066 ( .B(n19840), .A(n19841), .Z(n19839) );
XOR U33067 ( .A(c6613), .B(b[6613]), .Z(n19840) );
XNOR U33068 ( .A(b[6613]), .B(n19841), .Z(c[6613]) );
XNOR U33069 ( .A(a[6613]), .B(c6613), .Z(n19841) );
XOR U33070 ( .A(c6614), .B(n19842), .Z(c6615) );
ANDN U33071 ( .B(n19843), .A(n19844), .Z(n19842) );
XOR U33072 ( .A(c6614), .B(b[6614]), .Z(n19843) );
XNOR U33073 ( .A(b[6614]), .B(n19844), .Z(c[6614]) );
XNOR U33074 ( .A(a[6614]), .B(c6614), .Z(n19844) );
XOR U33075 ( .A(c6615), .B(n19845), .Z(c6616) );
ANDN U33076 ( .B(n19846), .A(n19847), .Z(n19845) );
XOR U33077 ( .A(c6615), .B(b[6615]), .Z(n19846) );
XNOR U33078 ( .A(b[6615]), .B(n19847), .Z(c[6615]) );
XNOR U33079 ( .A(a[6615]), .B(c6615), .Z(n19847) );
XOR U33080 ( .A(c6616), .B(n19848), .Z(c6617) );
ANDN U33081 ( .B(n19849), .A(n19850), .Z(n19848) );
XOR U33082 ( .A(c6616), .B(b[6616]), .Z(n19849) );
XNOR U33083 ( .A(b[6616]), .B(n19850), .Z(c[6616]) );
XNOR U33084 ( .A(a[6616]), .B(c6616), .Z(n19850) );
XOR U33085 ( .A(c6617), .B(n19851), .Z(c6618) );
ANDN U33086 ( .B(n19852), .A(n19853), .Z(n19851) );
XOR U33087 ( .A(c6617), .B(b[6617]), .Z(n19852) );
XNOR U33088 ( .A(b[6617]), .B(n19853), .Z(c[6617]) );
XNOR U33089 ( .A(a[6617]), .B(c6617), .Z(n19853) );
XOR U33090 ( .A(c6618), .B(n19854), .Z(c6619) );
ANDN U33091 ( .B(n19855), .A(n19856), .Z(n19854) );
XOR U33092 ( .A(c6618), .B(b[6618]), .Z(n19855) );
XNOR U33093 ( .A(b[6618]), .B(n19856), .Z(c[6618]) );
XNOR U33094 ( .A(a[6618]), .B(c6618), .Z(n19856) );
XOR U33095 ( .A(c6619), .B(n19857), .Z(c6620) );
ANDN U33096 ( .B(n19858), .A(n19859), .Z(n19857) );
XOR U33097 ( .A(c6619), .B(b[6619]), .Z(n19858) );
XNOR U33098 ( .A(b[6619]), .B(n19859), .Z(c[6619]) );
XNOR U33099 ( .A(a[6619]), .B(c6619), .Z(n19859) );
XOR U33100 ( .A(c6620), .B(n19860), .Z(c6621) );
ANDN U33101 ( .B(n19861), .A(n19862), .Z(n19860) );
XOR U33102 ( .A(c6620), .B(b[6620]), .Z(n19861) );
XNOR U33103 ( .A(b[6620]), .B(n19862), .Z(c[6620]) );
XNOR U33104 ( .A(a[6620]), .B(c6620), .Z(n19862) );
XOR U33105 ( .A(c6621), .B(n19863), .Z(c6622) );
ANDN U33106 ( .B(n19864), .A(n19865), .Z(n19863) );
XOR U33107 ( .A(c6621), .B(b[6621]), .Z(n19864) );
XNOR U33108 ( .A(b[6621]), .B(n19865), .Z(c[6621]) );
XNOR U33109 ( .A(a[6621]), .B(c6621), .Z(n19865) );
XOR U33110 ( .A(c6622), .B(n19866), .Z(c6623) );
ANDN U33111 ( .B(n19867), .A(n19868), .Z(n19866) );
XOR U33112 ( .A(c6622), .B(b[6622]), .Z(n19867) );
XNOR U33113 ( .A(b[6622]), .B(n19868), .Z(c[6622]) );
XNOR U33114 ( .A(a[6622]), .B(c6622), .Z(n19868) );
XOR U33115 ( .A(c6623), .B(n19869), .Z(c6624) );
ANDN U33116 ( .B(n19870), .A(n19871), .Z(n19869) );
XOR U33117 ( .A(c6623), .B(b[6623]), .Z(n19870) );
XNOR U33118 ( .A(b[6623]), .B(n19871), .Z(c[6623]) );
XNOR U33119 ( .A(a[6623]), .B(c6623), .Z(n19871) );
XOR U33120 ( .A(c6624), .B(n19872), .Z(c6625) );
ANDN U33121 ( .B(n19873), .A(n19874), .Z(n19872) );
XOR U33122 ( .A(c6624), .B(b[6624]), .Z(n19873) );
XNOR U33123 ( .A(b[6624]), .B(n19874), .Z(c[6624]) );
XNOR U33124 ( .A(a[6624]), .B(c6624), .Z(n19874) );
XOR U33125 ( .A(c6625), .B(n19875), .Z(c6626) );
ANDN U33126 ( .B(n19876), .A(n19877), .Z(n19875) );
XOR U33127 ( .A(c6625), .B(b[6625]), .Z(n19876) );
XNOR U33128 ( .A(b[6625]), .B(n19877), .Z(c[6625]) );
XNOR U33129 ( .A(a[6625]), .B(c6625), .Z(n19877) );
XOR U33130 ( .A(c6626), .B(n19878), .Z(c6627) );
ANDN U33131 ( .B(n19879), .A(n19880), .Z(n19878) );
XOR U33132 ( .A(c6626), .B(b[6626]), .Z(n19879) );
XNOR U33133 ( .A(b[6626]), .B(n19880), .Z(c[6626]) );
XNOR U33134 ( .A(a[6626]), .B(c6626), .Z(n19880) );
XOR U33135 ( .A(c6627), .B(n19881), .Z(c6628) );
ANDN U33136 ( .B(n19882), .A(n19883), .Z(n19881) );
XOR U33137 ( .A(c6627), .B(b[6627]), .Z(n19882) );
XNOR U33138 ( .A(b[6627]), .B(n19883), .Z(c[6627]) );
XNOR U33139 ( .A(a[6627]), .B(c6627), .Z(n19883) );
XOR U33140 ( .A(c6628), .B(n19884), .Z(c6629) );
ANDN U33141 ( .B(n19885), .A(n19886), .Z(n19884) );
XOR U33142 ( .A(c6628), .B(b[6628]), .Z(n19885) );
XNOR U33143 ( .A(b[6628]), .B(n19886), .Z(c[6628]) );
XNOR U33144 ( .A(a[6628]), .B(c6628), .Z(n19886) );
XOR U33145 ( .A(c6629), .B(n19887), .Z(c6630) );
ANDN U33146 ( .B(n19888), .A(n19889), .Z(n19887) );
XOR U33147 ( .A(c6629), .B(b[6629]), .Z(n19888) );
XNOR U33148 ( .A(b[6629]), .B(n19889), .Z(c[6629]) );
XNOR U33149 ( .A(a[6629]), .B(c6629), .Z(n19889) );
XOR U33150 ( .A(c6630), .B(n19890), .Z(c6631) );
ANDN U33151 ( .B(n19891), .A(n19892), .Z(n19890) );
XOR U33152 ( .A(c6630), .B(b[6630]), .Z(n19891) );
XNOR U33153 ( .A(b[6630]), .B(n19892), .Z(c[6630]) );
XNOR U33154 ( .A(a[6630]), .B(c6630), .Z(n19892) );
XOR U33155 ( .A(c6631), .B(n19893), .Z(c6632) );
ANDN U33156 ( .B(n19894), .A(n19895), .Z(n19893) );
XOR U33157 ( .A(c6631), .B(b[6631]), .Z(n19894) );
XNOR U33158 ( .A(b[6631]), .B(n19895), .Z(c[6631]) );
XNOR U33159 ( .A(a[6631]), .B(c6631), .Z(n19895) );
XOR U33160 ( .A(c6632), .B(n19896), .Z(c6633) );
ANDN U33161 ( .B(n19897), .A(n19898), .Z(n19896) );
XOR U33162 ( .A(c6632), .B(b[6632]), .Z(n19897) );
XNOR U33163 ( .A(b[6632]), .B(n19898), .Z(c[6632]) );
XNOR U33164 ( .A(a[6632]), .B(c6632), .Z(n19898) );
XOR U33165 ( .A(c6633), .B(n19899), .Z(c6634) );
ANDN U33166 ( .B(n19900), .A(n19901), .Z(n19899) );
XOR U33167 ( .A(c6633), .B(b[6633]), .Z(n19900) );
XNOR U33168 ( .A(b[6633]), .B(n19901), .Z(c[6633]) );
XNOR U33169 ( .A(a[6633]), .B(c6633), .Z(n19901) );
XOR U33170 ( .A(c6634), .B(n19902), .Z(c6635) );
ANDN U33171 ( .B(n19903), .A(n19904), .Z(n19902) );
XOR U33172 ( .A(c6634), .B(b[6634]), .Z(n19903) );
XNOR U33173 ( .A(b[6634]), .B(n19904), .Z(c[6634]) );
XNOR U33174 ( .A(a[6634]), .B(c6634), .Z(n19904) );
XOR U33175 ( .A(c6635), .B(n19905), .Z(c6636) );
ANDN U33176 ( .B(n19906), .A(n19907), .Z(n19905) );
XOR U33177 ( .A(c6635), .B(b[6635]), .Z(n19906) );
XNOR U33178 ( .A(b[6635]), .B(n19907), .Z(c[6635]) );
XNOR U33179 ( .A(a[6635]), .B(c6635), .Z(n19907) );
XOR U33180 ( .A(c6636), .B(n19908), .Z(c6637) );
ANDN U33181 ( .B(n19909), .A(n19910), .Z(n19908) );
XOR U33182 ( .A(c6636), .B(b[6636]), .Z(n19909) );
XNOR U33183 ( .A(b[6636]), .B(n19910), .Z(c[6636]) );
XNOR U33184 ( .A(a[6636]), .B(c6636), .Z(n19910) );
XOR U33185 ( .A(c6637), .B(n19911), .Z(c6638) );
ANDN U33186 ( .B(n19912), .A(n19913), .Z(n19911) );
XOR U33187 ( .A(c6637), .B(b[6637]), .Z(n19912) );
XNOR U33188 ( .A(b[6637]), .B(n19913), .Z(c[6637]) );
XNOR U33189 ( .A(a[6637]), .B(c6637), .Z(n19913) );
XOR U33190 ( .A(c6638), .B(n19914), .Z(c6639) );
ANDN U33191 ( .B(n19915), .A(n19916), .Z(n19914) );
XOR U33192 ( .A(c6638), .B(b[6638]), .Z(n19915) );
XNOR U33193 ( .A(b[6638]), .B(n19916), .Z(c[6638]) );
XNOR U33194 ( .A(a[6638]), .B(c6638), .Z(n19916) );
XOR U33195 ( .A(c6639), .B(n19917), .Z(c6640) );
ANDN U33196 ( .B(n19918), .A(n19919), .Z(n19917) );
XOR U33197 ( .A(c6639), .B(b[6639]), .Z(n19918) );
XNOR U33198 ( .A(b[6639]), .B(n19919), .Z(c[6639]) );
XNOR U33199 ( .A(a[6639]), .B(c6639), .Z(n19919) );
XOR U33200 ( .A(c6640), .B(n19920), .Z(c6641) );
ANDN U33201 ( .B(n19921), .A(n19922), .Z(n19920) );
XOR U33202 ( .A(c6640), .B(b[6640]), .Z(n19921) );
XNOR U33203 ( .A(b[6640]), .B(n19922), .Z(c[6640]) );
XNOR U33204 ( .A(a[6640]), .B(c6640), .Z(n19922) );
XOR U33205 ( .A(c6641), .B(n19923), .Z(c6642) );
ANDN U33206 ( .B(n19924), .A(n19925), .Z(n19923) );
XOR U33207 ( .A(c6641), .B(b[6641]), .Z(n19924) );
XNOR U33208 ( .A(b[6641]), .B(n19925), .Z(c[6641]) );
XNOR U33209 ( .A(a[6641]), .B(c6641), .Z(n19925) );
XOR U33210 ( .A(c6642), .B(n19926), .Z(c6643) );
ANDN U33211 ( .B(n19927), .A(n19928), .Z(n19926) );
XOR U33212 ( .A(c6642), .B(b[6642]), .Z(n19927) );
XNOR U33213 ( .A(b[6642]), .B(n19928), .Z(c[6642]) );
XNOR U33214 ( .A(a[6642]), .B(c6642), .Z(n19928) );
XOR U33215 ( .A(c6643), .B(n19929), .Z(c6644) );
ANDN U33216 ( .B(n19930), .A(n19931), .Z(n19929) );
XOR U33217 ( .A(c6643), .B(b[6643]), .Z(n19930) );
XNOR U33218 ( .A(b[6643]), .B(n19931), .Z(c[6643]) );
XNOR U33219 ( .A(a[6643]), .B(c6643), .Z(n19931) );
XOR U33220 ( .A(c6644), .B(n19932), .Z(c6645) );
ANDN U33221 ( .B(n19933), .A(n19934), .Z(n19932) );
XOR U33222 ( .A(c6644), .B(b[6644]), .Z(n19933) );
XNOR U33223 ( .A(b[6644]), .B(n19934), .Z(c[6644]) );
XNOR U33224 ( .A(a[6644]), .B(c6644), .Z(n19934) );
XOR U33225 ( .A(c6645), .B(n19935), .Z(c6646) );
ANDN U33226 ( .B(n19936), .A(n19937), .Z(n19935) );
XOR U33227 ( .A(c6645), .B(b[6645]), .Z(n19936) );
XNOR U33228 ( .A(b[6645]), .B(n19937), .Z(c[6645]) );
XNOR U33229 ( .A(a[6645]), .B(c6645), .Z(n19937) );
XOR U33230 ( .A(c6646), .B(n19938), .Z(c6647) );
ANDN U33231 ( .B(n19939), .A(n19940), .Z(n19938) );
XOR U33232 ( .A(c6646), .B(b[6646]), .Z(n19939) );
XNOR U33233 ( .A(b[6646]), .B(n19940), .Z(c[6646]) );
XNOR U33234 ( .A(a[6646]), .B(c6646), .Z(n19940) );
XOR U33235 ( .A(c6647), .B(n19941), .Z(c6648) );
ANDN U33236 ( .B(n19942), .A(n19943), .Z(n19941) );
XOR U33237 ( .A(c6647), .B(b[6647]), .Z(n19942) );
XNOR U33238 ( .A(b[6647]), .B(n19943), .Z(c[6647]) );
XNOR U33239 ( .A(a[6647]), .B(c6647), .Z(n19943) );
XOR U33240 ( .A(c6648), .B(n19944), .Z(c6649) );
ANDN U33241 ( .B(n19945), .A(n19946), .Z(n19944) );
XOR U33242 ( .A(c6648), .B(b[6648]), .Z(n19945) );
XNOR U33243 ( .A(b[6648]), .B(n19946), .Z(c[6648]) );
XNOR U33244 ( .A(a[6648]), .B(c6648), .Z(n19946) );
XOR U33245 ( .A(c6649), .B(n19947), .Z(c6650) );
ANDN U33246 ( .B(n19948), .A(n19949), .Z(n19947) );
XOR U33247 ( .A(c6649), .B(b[6649]), .Z(n19948) );
XNOR U33248 ( .A(b[6649]), .B(n19949), .Z(c[6649]) );
XNOR U33249 ( .A(a[6649]), .B(c6649), .Z(n19949) );
XOR U33250 ( .A(c6650), .B(n19950), .Z(c6651) );
ANDN U33251 ( .B(n19951), .A(n19952), .Z(n19950) );
XOR U33252 ( .A(c6650), .B(b[6650]), .Z(n19951) );
XNOR U33253 ( .A(b[6650]), .B(n19952), .Z(c[6650]) );
XNOR U33254 ( .A(a[6650]), .B(c6650), .Z(n19952) );
XOR U33255 ( .A(c6651), .B(n19953), .Z(c6652) );
ANDN U33256 ( .B(n19954), .A(n19955), .Z(n19953) );
XOR U33257 ( .A(c6651), .B(b[6651]), .Z(n19954) );
XNOR U33258 ( .A(b[6651]), .B(n19955), .Z(c[6651]) );
XNOR U33259 ( .A(a[6651]), .B(c6651), .Z(n19955) );
XOR U33260 ( .A(c6652), .B(n19956), .Z(c6653) );
ANDN U33261 ( .B(n19957), .A(n19958), .Z(n19956) );
XOR U33262 ( .A(c6652), .B(b[6652]), .Z(n19957) );
XNOR U33263 ( .A(b[6652]), .B(n19958), .Z(c[6652]) );
XNOR U33264 ( .A(a[6652]), .B(c6652), .Z(n19958) );
XOR U33265 ( .A(c6653), .B(n19959), .Z(c6654) );
ANDN U33266 ( .B(n19960), .A(n19961), .Z(n19959) );
XOR U33267 ( .A(c6653), .B(b[6653]), .Z(n19960) );
XNOR U33268 ( .A(b[6653]), .B(n19961), .Z(c[6653]) );
XNOR U33269 ( .A(a[6653]), .B(c6653), .Z(n19961) );
XOR U33270 ( .A(c6654), .B(n19962), .Z(c6655) );
ANDN U33271 ( .B(n19963), .A(n19964), .Z(n19962) );
XOR U33272 ( .A(c6654), .B(b[6654]), .Z(n19963) );
XNOR U33273 ( .A(b[6654]), .B(n19964), .Z(c[6654]) );
XNOR U33274 ( .A(a[6654]), .B(c6654), .Z(n19964) );
XOR U33275 ( .A(c6655), .B(n19965), .Z(c6656) );
ANDN U33276 ( .B(n19966), .A(n19967), .Z(n19965) );
XOR U33277 ( .A(c6655), .B(b[6655]), .Z(n19966) );
XNOR U33278 ( .A(b[6655]), .B(n19967), .Z(c[6655]) );
XNOR U33279 ( .A(a[6655]), .B(c6655), .Z(n19967) );
XOR U33280 ( .A(c6656), .B(n19968), .Z(c6657) );
ANDN U33281 ( .B(n19969), .A(n19970), .Z(n19968) );
XOR U33282 ( .A(c6656), .B(b[6656]), .Z(n19969) );
XNOR U33283 ( .A(b[6656]), .B(n19970), .Z(c[6656]) );
XNOR U33284 ( .A(a[6656]), .B(c6656), .Z(n19970) );
XOR U33285 ( .A(c6657), .B(n19971), .Z(c6658) );
ANDN U33286 ( .B(n19972), .A(n19973), .Z(n19971) );
XOR U33287 ( .A(c6657), .B(b[6657]), .Z(n19972) );
XNOR U33288 ( .A(b[6657]), .B(n19973), .Z(c[6657]) );
XNOR U33289 ( .A(a[6657]), .B(c6657), .Z(n19973) );
XOR U33290 ( .A(c6658), .B(n19974), .Z(c6659) );
ANDN U33291 ( .B(n19975), .A(n19976), .Z(n19974) );
XOR U33292 ( .A(c6658), .B(b[6658]), .Z(n19975) );
XNOR U33293 ( .A(b[6658]), .B(n19976), .Z(c[6658]) );
XNOR U33294 ( .A(a[6658]), .B(c6658), .Z(n19976) );
XOR U33295 ( .A(c6659), .B(n19977), .Z(c6660) );
ANDN U33296 ( .B(n19978), .A(n19979), .Z(n19977) );
XOR U33297 ( .A(c6659), .B(b[6659]), .Z(n19978) );
XNOR U33298 ( .A(b[6659]), .B(n19979), .Z(c[6659]) );
XNOR U33299 ( .A(a[6659]), .B(c6659), .Z(n19979) );
XOR U33300 ( .A(c6660), .B(n19980), .Z(c6661) );
ANDN U33301 ( .B(n19981), .A(n19982), .Z(n19980) );
XOR U33302 ( .A(c6660), .B(b[6660]), .Z(n19981) );
XNOR U33303 ( .A(b[6660]), .B(n19982), .Z(c[6660]) );
XNOR U33304 ( .A(a[6660]), .B(c6660), .Z(n19982) );
XOR U33305 ( .A(c6661), .B(n19983), .Z(c6662) );
ANDN U33306 ( .B(n19984), .A(n19985), .Z(n19983) );
XOR U33307 ( .A(c6661), .B(b[6661]), .Z(n19984) );
XNOR U33308 ( .A(b[6661]), .B(n19985), .Z(c[6661]) );
XNOR U33309 ( .A(a[6661]), .B(c6661), .Z(n19985) );
XOR U33310 ( .A(c6662), .B(n19986), .Z(c6663) );
ANDN U33311 ( .B(n19987), .A(n19988), .Z(n19986) );
XOR U33312 ( .A(c6662), .B(b[6662]), .Z(n19987) );
XNOR U33313 ( .A(b[6662]), .B(n19988), .Z(c[6662]) );
XNOR U33314 ( .A(a[6662]), .B(c6662), .Z(n19988) );
XOR U33315 ( .A(c6663), .B(n19989), .Z(c6664) );
ANDN U33316 ( .B(n19990), .A(n19991), .Z(n19989) );
XOR U33317 ( .A(c6663), .B(b[6663]), .Z(n19990) );
XNOR U33318 ( .A(b[6663]), .B(n19991), .Z(c[6663]) );
XNOR U33319 ( .A(a[6663]), .B(c6663), .Z(n19991) );
XOR U33320 ( .A(c6664), .B(n19992), .Z(c6665) );
ANDN U33321 ( .B(n19993), .A(n19994), .Z(n19992) );
XOR U33322 ( .A(c6664), .B(b[6664]), .Z(n19993) );
XNOR U33323 ( .A(b[6664]), .B(n19994), .Z(c[6664]) );
XNOR U33324 ( .A(a[6664]), .B(c6664), .Z(n19994) );
XOR U33325 ( .A(c6665), .B(n19995), .Z(c6666) );
ANDN U33326 ( .B(n19996), .A(n19997), .Z(n19995) );
XOR U33327 ( .A(c6665), .B(b[6665]), .Z(n19996) );
XNOR U33328 ( .A(b[6665]), .B(n19997), .Z(c[6665]) );
XNOR U33329 ( .A(a[6665]), .B(c6665), .Z(n19997) );
XOR U33330 ( .A(c6666), .B(n19998), .Z(c6667) );
ANDN U33331 ( .B(n19999), .A(n20000), .Z(n19998) );
XOR U33332 ( .A(c6666), .B(b[6666]), .Z(n19999) );
XNOR U33333 ( .A(b[6666]), .B(n20000), .Z(c[6666]) );
XNOR U33334 ( .A(a[6666]), .B(c6666), .Z(n20000) );
XOR U33335 ( .A(c6667), .B(n20001), .Z(c6668) );
ANDN U33336 ( .B(n20002), .A(n20003), .Z(n20001) );
XOR U33337 ( .A(c6667), .B(b[6667]), .Z(n20002) );
XNOR U33338 ( .A(b[6667]), .B(n20003), .Z(c[6667]) );
XNOR U33339 ( .A(a[6667]), .B(c6667), .Z(n20003) );
XOR U33340 ( .A(c6668), .B(n20004), .Z(c6669) );
ANDN U33341 ( .B(n20005), .A(n20006), .Z(n20004) );
XOR U33342 ( .A(c6668), .B(b[6668]), .Z(n20005) );
XNOR U33343 ( .A(b[6668]), .B(n20006), .Z(c[6668]) );
XNOR U33344 ( .A(a[6668]), .B(c6668), .Z(n20006) );
XOR U33345 ( .A(c6669), .B(n20007), .Z(c6670) );
ANDN U33346 ( .B(n20008), .A(n20009), .Z(n20007) );
XOR U33347 ( .A(c6669), .B(b[6669]), .Z(n20008) );
XNOR U33348 ( .A(b[6669]), .B(n20009), .Z(c[6669]) );
XNOR U33349 ( .A(a[6669]), .B(c6669), .Z(n20009) );
XOR U33350 ( .A(c6670), .B(n20010), .Z(c6671) );
ANDN U33351 ( .B(n20011), .A(n20012), .Z(n20010) );
XOR U33352 ( .A(c6670), .B(b[6670]), .Z(n20011) );
XNOR U33353 ( .A(b[6670]), .B(n20012), .Z(c[6670]) );
XNOR U33354 ( .A(a[6670]), .B(c6670), .Z(n20012) );
XOR U33355 ( .A(c6671), .B(n20013), .Z(c6672) );
ANDN U33356 ( .B(n20014), .A(n20015), .Z(n20013) );
XOR U33357 ( .A(c6671), .B(b[6671]), .Z(n20014) );
XNOR U33358 ( .A(b[6671]), .B(n20015), .Z(c[6671]) );
XNOR U33359 ( .A(a[6671]), .B(c6671), .Z(n20015) );
XOR U33360 ( .A(c6672), .B(n20016), .Z(c6673) );
ANDN U33361 ( .B(n20017), .A(n20018), .Z(n20016) );
XOR U33362 ( .A(c6672), .B(b[6672]), .Z(n20017) );
XNOR U33363 ( .A(b[6672]), .B(n20018), .Z(c[6672]) );
XNOR U33364 ( .A(a[6672]), .B(c6672), .Z(n20018) );
XOR U33365 ( .A(c6673), .B(n20019), .Z(c6674) );
ANDN U33366 ( .B(n20020), .A(n20021), .Z(n20019) );
XOR U33367 ( .A(c6673), .B(b[6673]), .Z(n20020) );
XNOR U33368 ( .A(b[6673]), .B(n20021), .Z(c[6673]) );
XNOR U33369 ( .A(a[6673]), .B(c6673), .Z(n20021) );
XOR U33370 ( .A(c6674), .B(n20022), .Z(c6675) );
ANDN U33371 ( .B(n20023), .A(n20024), .Z(n20022) );
XOR U33372 ( .A(c6674), .B(b[6674]), .Z(n20023) );
XNOR U33373 ( .A(b[6674]), .B(n20024), .Z(c[6674]) );
XNOR U33374 ( .A(a[6674]), .B(c6674), .Z(n20024) );
XOR U33375 ( .A(c6675), .B(n20025), .Z(c6676) );
ANDN U33376 ( .B(n20026), .A(n20027), .Z(n20025) );
XOR U33377 ( .A(c6675), .B(b[6675]), .Z(n20026) );
XNOR U33378 ( .A(b[6675]), .B(n20027), .Z(c[6675]) );
XNOR U33379 ( .A(a[6675]), .B(c6675), .Z(n20027) );
XOR U33380 ( .A(c6676), .B(n20028), .Z(c6677) );
ANDN U33381 ( .B(n20029), .A(n20030), .Z(n20028) );
XOR U33382 ( .A(c6676), .B(b[6676]), .Z(n20029) );
XNOR U33383 ( .A(b[6676]), .B(n20030), .Z(c[6676]) );
XNOR U33384 ( .A(a[6676]), .B(c6676), .Z(n20030) );
XOR U33385 ( .A(c6677), .B(n20031), .Z(c6678) );
ANDN U33386 ( .B(n20032), .A(n20033), .Z(n20031) );
XOR U33387 ( .A(c6677), .B(b[6677]), .Z(n20032) );
XNOR U33388 ( .A(b[6677]), .B(n20033), .Z(c[6677]) );
XNOR U33389 ( .A(a[6677]), .B(c6677), .Z(n20033) );
XOR U33390 ( .A(c6678), .B(n20034), .Z(c6679) );
ANDN U33391 ( .B(n20035), .A(n20036), .Z(n20034) );
XOR U33392 ( .A(c6678), .B(b[6678]), .Z(n20035) );
XNOR U33393 ( .A(b[6678]), .B(n20036), .Z(c[6678]) );
XNOR U33394 ( .A(a[6678]), .B(c6678), .Z(n20036) );
XOR U33395 ( .A(c6679), .B(n20037), .Z(c6680) );
ANDN U33396 ( .B(n20038), .A(n20039), .Z(n20037) );
XOR U33397 ( .A(c6679), .B(b[6679]), .Z(n20038) );
XNOR U33398 ( .A(b[6679]), .B(n20039), .Z(c[6679]) );
XNOR U33399 ( .A(a[6679]), .B(c6679), .Z(n20039) );
XOR U33400 ( .A(c6680), .B(n20040), .Z(c6681) );
ANDN U33401 ( .B(n20041), .A(n20042), .Z(n20040) );
XOR U33402 ( .A(c6680), .B(b[6680]), .Z(n20041) );
XNOR U33403 ( .A(b[6680]), .B(n20042), .Z(c[6680]) );
XNOR U33404 ( .A(a[6680]), .B(c6680), .Z(n20042) );
XOR U33405 ( .A(c6681), .B(n20043), .Z(c6682) );
ANDN U33406 ( .B(n20044), .A(n20045), .Z(n20043) );
XOR U33407 ( .A(c6681), .B(b[6681]), .Z(n20044) );
XNOR U33408 ( .A(b[6681]), .B(n20045), .Z(c[6681]) );
XNOR U33409 ( .A(a[6681]), .B(c6681), .Z(n20045) );
XOR U33410 ( .A(c6682), .B(n20046), .Z(c6683) );
ANDN U33411 ( .B(n20047), .A(n20048), .Z(n20046) );
XOR U33412 ( .A(c6682), .B(b[6682]), .Z(n20047) );
XNOR U33413 ( .A(b[6682]), .B(n20048), .Z(c[6682]) );
XNOR U33414 ( .A(a[6682]), .B(c6682), .Z(n20048) );
XOR U33415 ( .A(c6683), .B(n20049), .Z(c6684) );
ANDN U33416 ( .B(n20050), .A(n20051), .Z(n20049) );
XOR U33417 ( .A(c6683), .B(b[6683]), .Z(n20050) );
XNOR U33418 ( .A(b[6683]), .B(n20051), .Z(c[6683]) );
XNOR U33419 ( .A(a[6683]), .B(c6683), .Z(n20051) );
XOR U33420 ( .A(c6684), .B(n20052), .Z(c6685) );
ANDN U33421 ( .B(n20053), .A(n20054), .Z(n20052) );
XOR U33422 ( .A(c6684), .B(b[6684]), .Z(n20053) );
XNOR U33423 ( .A(b[6684]), .B(n20054), .Z(c[6684]) );
XNOR U33424 ( .A(a[6684]), .B(c6684), .Z(n20054) );
XOR U33425 ( .A(c6685), .B(n20055), .Z(c6686) );
ANDN U33426 ( .B(n20056), .A(n20057), .Z(n20055) );
XOR U33427 ( .A(c6685), .B(b[6685]), .Z(n20056) );
XNOR U33428 ( .A(b[6685]), .B(n20057), .Z(c[6685]) );
XNOR U33429 ( .A(a[6685]), .B(c6685), .Z(n20057) );
XOR U33430 ( .A(c6686), .B(n20058), .Z(c6687) );
ANDN U33431 ( .B(n20059), .A(n20060), .Z(n20058) );
XOR U33432 ( .A(c6686), .B(b[6686]), .Z(n20059) );
XNOR U33433 ( .A(b[6686]), .B(n20060), .Z(c[6686]) );
XNOR U33434 ( .A(a[6686]), .B(c6686), .Z(n20060) );
XOR U33435 ( .A(c6687), .B(n20061), .Z(c6688) );
ANDN U33436 ( .B(n20062), .A(n20063), .Z(n20061) );
XOR U33437 ( .A(c6687), .B(b[6687]), .Z(n20062) );
XNOR U33438 ( .A(b[6687]), .B(n20063), .Z(c[6687]) );
XNOR U33439 ( .A(a[6687]), .B(c6687), .Z(n20063) );
XOR U33440 ( .A(c6688), .B(n20064), .Z(c6689) );
ANDN U33441 ( .B(n20065), .A(n20066), .Z(n20064) );
XOR U33442 ( .A(c6688), .B(b[6688]), .Z(n20065) );
XNOR U33443 ( .A(b[6688]), .B(n20066), .Z(c[6688]) );
XNOR U33444 ( .A(a[6688]), .B(c6688), .Z(n20066) );
XOR U33445 ( .A(c6689), .B(n20067), .Z(c6690) );
ANDN U33446 ( .B(n20068), .A(n20069), .Z(n20067) );
XOR U33447 ( .A(c6689), .B(b[6689]), .Z(n20068) );
XNOR U33448 ( .A(b[6689]), .B(n20069), .Z(c[6689]) );
XNOR U33449 ( .A(a[6689]), .B(c6689), .Z(n20069) );
XOR U33450 ( .A(c6690), .B(n20070), .Z(c6691) );
ANDN U33451 ( .B(n20071), .A(n20072), .Z(n20070) );
XOR U33452 ( .A(c6690), .B(b[6690]), .Z(n20071) );
XNOR U33453 ( .A(b[6690]), .B(n20072), .Z(c[6690]) );
XNOR U33454 ( .A(a[6690]), .B(c6690), .Z(n20072) );
XOR U33455 ( .A(c6691), .B(n20073), .Z(c6692) );
ANDN U33456 ( .B(n20074), .A(n20075), .Z(n20073) );
XOR U33457 ( .A(c6691), .B(b[6691]), .Z(n20074) );
XNOR U33458 ( .A(b[6691]), .B(n20075), .Z(c[6691]) );
XNOR U33459 ( .A(a[6691]), .B(c6691), .Z(n20075) );
XOR U33460 ( .A(c6692), .B(n20076), .Z(c6693) );
ANDN U33461 ( .B(n20077), .A(n20078), .Z(n20076) );
XOR U33462 ( .A(c6692), .B(b[6692]), .Z(n20077) );
XNOR U33463 ( .A(b[6692]), .B(n20078), .Z(c[6692]) );
XNOR U33464 ( .A(a[6692]), .B(c6692), .Z(n20078) );
XOR U33465 ( .A(c6693), .B(n20079), .Z(c6694) );
ANDN U33466 ( .B(n20080), .A(n20081), .Z(n20079) );
XOR U33467 ( .A(c6693), .B(b[6693]), .Z(n20080) );
XNOR U33468 ( .A(b[6693]), .B(n20081), .Z(c[6693]) );
XNOR U33469 ( .A(a[6693]), .B(c6693), .Z(n20081) );
XOR U33470 ( .A(c6694), .B(n20082), .Z(c6695) );
ANDN U33471 ( .B(n20083), .A(n20084), .Z(n20082) );
XOR U33472 ( .A(c6694), .B(b[6694]), .Z(n20083) );
XNOR U33473 ( .A(b[6694]), .B(n20084), .Z(c[6694]) );
XNOR U33474 ( .A(a[6694]), .B(c6694), .Z(n20084) );
XOR U33475 ( .A(c6695), .B(n20085), .Z(c6696) );
ANDN U33476 ( .B(n20086), .A(n20087), .Z(n20085) );
XOR U33477 ( .A(c6695), .B(b[6695]), .Z(n20086) );
XNOR U33478 ( .A(b[6695]), .B(n20087), .Z(c[6695]) );
XNOR U33479 ( .A(a[6695]), .B(c6695), .Z(n20087) );
XOR U33480 ( .A(c6696), .B(n20088), .Z(c6697) );
ANDN U33481 ( .B(n20089), .A(n20090), .Z(n20088) );
XOR U33482 ( .A(c6696), .B(b[6696]), .Z(n20089) );
XNOR U33483 ( .A(b[6696]), .B(n20090), .Z(c[6696]) );
XNOR U33484 ( .A(a[6696]), .B(c6696), .Z(n20090) );
XOR U33485 ( .A(c6697), .B(n20091), .Z(c6698) );
ANDN U33486 ( .B(n20092), .A(n20093), .Z(n20091) );
XOR U33487 ( .A(c6697), .B(b[6697]), .Z(n20092) );
XNOR U33488 ( .A(b[6697]), .B(n20093), .Z(c[6697]) );
XNOR U33489 ( .A(a[6697]), .B(c6697), .Z(n20093) );
XOR U33490 ( .A(c6698), .B(n20094), .Z(c6699) );
ANDN U33491 ( .B(n20095), .A(n20096), .Z(n20094) );
XOR U33492 ( .A(c6698), .B(b[6698]), .Z(n20095) );
XNOR U33493 ( .A(b[6698]), .B(n20096), .Z(c[6698]) );
XNOR U33494 ( .A(a[6698]), .B(c6698), .Z(n20096) );
XOR U33495 ( .A(c6699), .B(n20097), .Z(c6700) );
ANDN U33496 ( .B(n20098), .A(n20099), .Z(n20097) );
XOR U33497 ( .A(c6699), .B(b[6699]), .Z(n20098) );
XNOR U33498 ( .A(b[6699]), .B(n20099), .Z(c[6699]) );
XNOR U33499 ( .A(a[6699]), .B(c6699), .Z(n20099) );
XOR U33500 ( .A(c6700), .B(n20100), .Z(c6701) );
ANDN U33501 ( .B(n20101), .A(n20102), .Z(n20100) );
XOR U33502 ( .A(c6700), .B(b[6700]), .Z(n20101) );
XNOR U33503 ( .A(b[6700]), .B(n20102), .Z(c[6700]) );
XNOR U33504 ( .A(a[6700]), .B(c6700), .Z(n20102) );
XOR U33505 ( .A(c6701), .B(n20103), .Z(c6702) );
ANDN U33506 ( .B(n20104), .A(n20105), .Z(n20103) );
XOR U33507 ( .A(c6701), .B(b[6701]), .Z(n20104) );
XNOR U33508 ( .A(b[6701]), .B(n20105), .Z(c[6701]) );
XNOR U33509 ( .A(a[6701]), .B(c6701), .Z(n20105) );
XOR U33510 ( .A(c6702), .B(n20106), .Z(c6703) );
ANDN U33511 ( .B(n20107), .A(n20108), .Z(n20106) );
XOR U33512 ( .A(c6702), .B(b[6702]), .Z(n20107) );
XNOR U33513 ( .A(b[6702]), .B(n20108), .Z(c[6702]) );
XNOR U33514 ( .A(a[6702]), .B(c6702), .Z(n20108) );
XOR U33515 ( .A(c6703), .B(n20109), .Z(c6704) );
ANDN U33516 ( .B(n20110), .A(n20111), .Z(n20109) );
XOR U33517 ( .A(c6703), .B(b[6703]), .Z(n20110) );
XNOR U33518 ( .A(b[6703]), .B(n20111), .Z(c[6703]) );
XNOR U33519 ( .A(a[6703]), .B(c6703), .Z(n20111) );
XOR U33520 ( .A(c6704), .B(n20112), .Z(c6705) );
ANDN U33521 ( .B(n20113), .A(n20114), .Z(n20112) );
XOR U33522 ( .A(c6704), .B(b[6704]), .Z(n20113) );
XNOR U33523 ( .A(b[6704]), .B(n20114), .Z(c[6704]) );
XNOR U33524 ( .A(a[6704]), .B(c6704), .Z(n20114) );
XOR U33525 ( .A(c6705), .B(n20115), .Z(c6706) );
ANDN U33526 ( .B(n20116), .A(n20117), .Z(n20115) );
XOR U33527 ( .A(c6705), .B(b[6705]), .Z(n20116) );
XNOR U33528 ( .A(b[6705]), .B(n20117), .Z(c[6705]) );
XNOR U33529 ( .A(a[6705]), .B(c6705), .Z(n20117) );
XOR U33530 ( .A(c6706), .B(n20118), .Z(c6707) );
ANDN U33531 ( .B(n20119), .A(n20120), .Z(n20118) );
XOR U33532 ( .A(c6706), .B(b[6706]), .Z(n20119) );
XNOR U33533 ( .A(b[6706]), .B(n20120), .Z(c[6706]) );
XNOR U33534 ( .A(a[6706]), .B(c6706), .Z(n20120) );
XOR U33535 ( .A(c6707), .B(n20121), .Z(c6708) );
ANDN U33536 ( .B(n20122), .A(n20123), .Z(n20121) );
XOR U33537 ( .A(c6707), .B(b[6707]), .Z(n20122) );
XNOR U33538 ( .A(b[6707]), .B(n20123), .Z(c[6707]) );
XNOR U33539 ( .A(a[6707]), .B(c6707), .Z(n20123) );
XOR U33540 ( .A(c6708), .B(n20124), .Z(c6709) );
ANDN U33541 ( .B(n20125), .A(n20126), .Z(n20124) );
XOR U33542 ( .A(c6708), .B(b[6708]), .Z(n20125) );
XNOR U33543 ( .A(b[6708]), .B(n20126), .Z(c[6708]) );
XNOR U33544 ( .A(a[6708]), .B(c6708), .Z(n20126) );
XOR U33545 ( .A(c6709), .B(n20127), .Z(c6710) );
ANDN U33546 ( .B(n20128), .A(n20129), .Z(n20127) );
XOR U33547 ( .A(c6709), .B(b[6709]), .Z(n20128) );
XNOR U33548 ( .A(b[6709]), .B(n20129), .Z(c[6709]) );
XNOR U33549 ( .A(a[6709]), .B(c6709), .Z(n20129) );
XOR U33550 ( .A(c6710), .B(n20130), .Z(c6711) );
ANDN U33551 ( .B(n20131), .A(n20132), .Z(n20130) );
XOR U33552 ( .A(c6710), .B(b[6710]), .Z(n20131) );
XNOR U33553 ( .A(b[6710]), .B(n20132), .Z(c[6710]) );
XNOR U33554 ( .A(a[6710]), .B(c6710), .Z(n20132) );
XOR U33555 ( .A(c6711), .B(n20133), .Z(c6712) );
ANDN U33556 ( .B(n20134), .A(n20135), .Z(n20133) );
XOR U33557 ( .A(c6711), .B(b[6711]), .Z(n20134) );
XNOR U33558 ( .A(b[6711]), .B(n20135), .Z(c[6711]) );
XNOR U33559 ( .A(a[6711]), .B(c6711), .Z(n20135) );
XOR U33560 ( .A(c6712), .B(n20136), .Z(c6713) );
ANDN U33561 ( .B(n20137), .A(n20138), .Z(n20136) );
XOR U33562 ( .A(c6712), .B(b[6712]), .Z(n20137) );
XNOR U33563 ( .A(b[6712]), .B(n20138), .Z(c[6712]) );
XNOR U33564 ( .A(a[6712]), .B(c6712), .Z(n20138) );
XOR U33565 ( .A(c6713), .B(n20139), .Z(c6714) );
ANDN U33566 ( .B(n20140), .A(n20141), .Z(n20139) );
XOR U33567 ( .A(c6713), .B(b[6713]), .Z(n20140) );
XNOR U33568 ( .A(b[6713]), .B(n20141), .Z(c[6713]) );
XNOR U33569 ( .A(a[6713]), .B(c6713), .Z(n20141) );
XOR U33570 ( .A(c6714), .B(n20142), .Z(c6715) );
ANDN U33571 ( .B(n20143), .A(n20144), .Z(n20142) );
XOR U33572 ( .A(c6714), .B(b[6714]), .Z(n20143) );
XNOR U33573 ( .A(b[6714]), .B(n20144), .Z(c[6714]) );
XNOR U33574 ( .A(a[6714]), .B(c6714), .Z(n20144) );
XOR U33575 ( .A(c6715), .B(n20145), .Z(c6716) );
ANDN U33576 ( .B(n20146), .A(n20147), .Z(n20145) );
XOR U33577 ( .A(c6715), .B(b[6715]), .Z(n20146) );
XNOR U33578 ( .A(b[6715]), .B(n20147), .Z(c[6715]) );
XNOR U33579 ( .A(a[6715]), .B(c6715), .Z(n20147) );
XOR U33580 ( .A(c6716), .B(n20148), .Z(c6717) );
ANDN U33581 ( .B(n20149), .A(n20150), .Z(n20148) );
XOR U33582 ( .A(c6716), .B(b[6716]), .Z(n20149) );
XNOR U33583 ( .A(b[6716]), .B(n20150), .Z(c[6716]) );
XNOR U33584 ( .A(a[6716]), .B(c6716), .Z(n20150) );
XOR U33585 ( .A(c6717), .B(n20151), .Z(c6718) );
ANDN U33586 ( .B(n20152), .A(n20153), .Z(n20151) );
XOR U33587 ( .A(c6717), .B(b[6717]), .Z(n20152) );
XNOR U33588 ( .A(b[6717]), .B(n20153), .Z(c[6717]) );
XNOR U33589 ( .A(a[6717]), .B(c6717), .Z(n20153) );
XOR U33590 ( .A(c6718), .B(n20154), .Z(c6719) );
ANDN U33591 ( .B(n20155), .A(n20156), .Z(n20154) );
XOR U33592 ( .A(c6718), .B(b[6718]), .Z(n20155) );
XNOR U33593 ( .A(b[6718]), .B(n20156), .Z(c[6718]) );
XNOR U33594 ( .A(a[6718]), .B(c6718), .Z(n20156) );
XOR U33595 ( .A(c6719), .B(n20157), .Z(c6720) );
ANDN U33596 ( .B(n20158), .A(n20159), .Z(n20157) );
XOR U33597 ( .A(c6719), .B(b[6719]), .Z(n20158) );
XNOR U33598 ( .A(b[6719]), .B(n20159), .Z(c[6719]) );
XNOR U33599 ( .A(a[6719]), .B(c6719), .Z(n20159) );
XOR U33600 ( .A(c6720), .B(n20160), .Z(c6721) );
ANDN U33601 ( .B(n20161), .A(n20162), .Z(n20160) );
XOR U33602 ( .A(c6720), .B(b[6720]), .Z(n20161) );
XNOR U33603 ( .A(b[6720]), .B(n20162), .Z(c[6720]) );
XNOR U33604 ( .A(a[6720]), .B(c6720), .Z(n20162) );
XOR U33605 ( .A(c6721), .B(n20163), .Z(c6722) );
ANDN U33606 ( .B(n20164), .A(n20165), .Z(n20163) );
XOR U33607 ( .A(c6721), .B(b[6721]), .Z(n20164) );
XNOR U33608 ( .A(b[6721]), .B(n20165), .Z(c[6721]) );
XNOR U33609 ( .A(a[6721]), .B(c6721), .Z(n20165) );
XOR U33610 ( .A(c6722), .B(n20166), .Z(c6723) );
ANDN U33611 ( .B(n20167), .A(n20168), .Z(n20166) );
XOR U33612 ( .A(c6722), .B(b[6722]), .Z(n20167) );
XNOR U33613 ( .A(b[6722]), .B(n20168), .Z(c[6722]) );
XNOR U33614 ( .A(a[6722]), .B(c6722), .Z(n20168) );
XOR U33615 ( .A(c6723), .B(n20169), .Z(c6724) );
ANDN U33616 ( .B(n20170), .A(n20171), .Z(n20169) );
XOR U33617 ( .A(c6723), .B(b[6723]), .Z(n20170) );
XNOR U33618 ( .A(b[6723]), .B(n20171), .Z(c[6723]) );
XNOR U33619 ( .A(a[6723]), .B(c6723), .Z(n20171) );
XOR U33620 ( .A(c6724), .B(n20172), .Z(c6725) );
ANDN U33621 ( .B(n20173), .A(n20174), .Z(n20172) );
XOR U33622 ( .A(c6724), .B(b[6724]), .Z(n20173) );
XNOR U33623 ( .A(b[6724]), .B(n20174), .Z(c[6724]) );
XNOR U33624 ( .A(a[6724]), .B(c6724), .Z(n20174) );
XOR U33625 ( .A(c6725), .B(n20175), .Z(c6726) );
ANDN U33626 ( .B(n20176), .A(n20177), .Z(n20175) );
XOR U33627 ( .A(c6725), .B(b[6725]), .Z(n20176) );
XNOR U33628 ( .A(b[6725]), .B(n20177), .Z(c[6725]) );
XNOR U33629 ( .A(a[6725]), .B(c6725), .Z(n20177) );
XOR U33630 ( .A(c6726), .B(n20178), .Z(c6727) );
ANDN U33631 ( .B(n20179), .A(n20180), .Z(n20178) );
XOR U33632 ( .A(c6726), .B(b[6726]), .Z(n20179) );
XNOR U33633 ( .A(b[6726]), .B(n20180), .Z(c[6726]) );
XNOR U33634 ( .A(a[6726]), .B(c6726), .Z(n20180) );
XOR U33635 ( .A(c6727), .B(n20181), .Z(c6728) );
ANDN U33636 ( .B(n20182), .A(n20183), .Z(n20181) );
XOR U33637 ( .A(c6727), .B(b[6727]), .Z(n20182) );
XNOR U33638 ( .A(b[6727]), .B(n20183), .Z(c[6727]) );
XNOR U33639 ( .A(a[6727]), .B(c6727), .Z(n20183) );
XOR U33640 ( .A(c6728), .B(n20184), .Z(c6729) );
ANDN U33641 ( .B(n20185), .A(n20186), .Z(n20184) );
XOR U33642 ( .A(c6728), .B(b[6728]), .Z(n20185) );
XNOR U33643 ( .A(b[6728]), .B(n20186), .Z(c[6728]) );
XNOR U33644 ( .A(a[6728]), .B(c6728), .Z(n20186) );
XOR U33645 ( .A(c6729), .B(n20187), .Z(c6730) );
ANDN U33646 ( .B(n20188), .A(n20189), .Z(n20187) );
XOR U33647 ( .A(c6729), .B(b[6729]), .Z(n20188) );
XNOR U33648 ( .A(b[6729]), .B(n20189), .Z(c[6729]) );
XNOR U33649 ( .A(a[6729]), .B(c6729), .Z(n20189) );
XOR U33650 ( .A(c6730), .B(n20190), .Z(c6731) );
ANDN U33651 ( .B(n20191), .A(n20192), .Z(n20190) );
XOR U33652 ( .A(c6730), .B(b[6730]), .Z(n20191) );
XNOR U33653 ( .A(b[6730]), .B(n20192), .Z(c[6730]) );
XNOR U33654 ( .A(a[6730]), .B(c6730), .Z(n20192) );
XOR U33655 ( .A(c6731), .B(n20193), .Z(c6732) );
ANDN U33656 ( .B(n20194), .A(n20195), .Z(n20193) );
XOR U33657 ( .A(c6731), .B(b[6731]), .Z(n20194) );
XNOR U33658 ( .A(b[6731]), .B(n20195), .Z(c[6731]) );
XNOR U33659 ( .A(a[6731]), .B(c6731), .Z(n20195) );
XOR U33660 ( .A(c6732), .B(n20196), .Z(c6733) );
ANDN U33661 ( .B(n20197), .A(n20198), .Z(n20196) );
XOR U33662 ( .A(c6732), .B(b[6732]), .Z(n20197) );
XNOR U33663 ( .A(b[6732]), .B(n20198), .Z(c[6732]) );
XNOR U33664 ( .A(a[6732]), .B(c6732), .Z(n20198) );
XOR U33665 ( .A(c6733), .B(n20199), .Z(c6734) );
ANDN U33666 ( .B(n20200), .A(n20201), .Z(n20199) );
XOR U33667 ( .A(c6733), .B(b[6733]), .Z(n20200) );
XNOR U33668 ( .A(b[6733]), .B(n20201), .Z(c[6733]) );
XNOR U33669 ( .A(a[6733]), .B(c6733), .Z(n20201) );
XOR U33670 ( .A(c6734), .B(n20202), .Z(c6735) );
ANDN U33671 ( .B(n20203), .A(n20204), .Z(n20202) );
XOR U33672 ( .A(c6734), .B(b[6734]), .Z(n20203) );
XNOR U33673 ( .A(b[6734]), .B(n20204), .Z(c[6734]) );
XNOR U33674 ( .A(a[6734]), .B(c6734), .Z(n20204) );
XOR U33675 ( .A(c6735), .B(n20205), .Z(c6736) );
ANDN U33676 ( .B(n20206), .A(n20207), .Z(n20205) );
XOR U33677 ( .A(c6735), .B(b[6735]), .Z(n20206) );
XNOR U33678 ( .A(b[6735]), .B(n20207), .Z(c[6735]) );
XNOR U33679 ( .A(a[6735]), .B(c6735), .Z(n20207) );
XOR U33680 ( .A(c6736), .B(n20208), .Z(c6737) );
ANDN U33681 ( .B(n20209), .A(n20210), .Z(n20208) );
XOR U33682 ( .A(c6736), .B(b[6736]), .Z(n20209) );
XNOR U33683 ( .A(b[6736]), .B(n20210), .Z(c[6736]) );
XNOR U33684 ( .A(a[6736]), .B(c6736), .Z(n20210) );
XOR U33685 ( .A(c6737), .B(n20211), .Z(c6738) );
ANDN U33686 ( .B(n20212), .A(n20213), .Z(n20211) );
XOR U33687 ( .A(c6737), .B(b[6737]), .Z(n20212) );
XNOR U33688 ( .A(b[6737]), .B(n20213), .Z(c[6737]) );
XNOR U33689 ( .A(a[6737]), .B(c6737), .Z(n20213) );
XOR U33690 ( .A(c6738), .B(n20214), .Z(c6739) );
ANDN U33691 ( .B(n20215), .A(n20216), .Z(n20214) );
XOR U33692 ( .A(c6738), .B(b[6738]), .Z(n20215) );
XNOR U33693 ( .A(b[6738]), .B(n20216), .Z(c[6738]) );
XNOR U33694 ( .A(a[6738]), .B(c6738), .Z(n20216) );
XOR U33695 ( .A(c6739), .B(n20217), .Z(c6740) );
ANDN U33696 ( .B(n20218), .A(n20219), .Z(n20217) );
XOR U33697 ( .A(c6739), .B(b[6739]), .Z(n20218) );
XNOR U33698 ( .A(b[6739]), .B(n20219), .Z(c[6739]) );
XNOR U33699 ( .A(a[6739]), .B(c6739), .Z(n20219) );
XOR U33700 ( .A(c6740), .B(n20220), .Z(c6741) );
ANDN U33701 ( .B(n20221), .A(n20222), .Z(n20220) );
XOR U33702 ( .A(c6740), .B(b[6740]), .Z(n20221) );
XNOR U33703 ( .A(b[6740]), .B(n20222), .Z(c[6740]) );
XNOR U33704 ( .A(a[6740]), .B(c6740), .Z(n20222) );
XOR U33705 ( .A(c6741), .B(n20223), .Z(c6742) );
ANDN U33706 ( .B(n20224), .A(n20225), .Z(n20223) );
XOR U33707 ( .A(c6741), .B(b[6741]), .Z(n20224) );
XNOR U33708 ( .A(b[6741]), .B(n20225), .Z(c[6741]) );
XNOR U33709 ( .A(a[6741]), .B(c6741), .Z(n20225) );
XOR U33710 ( .A(c6742), .B(n20226), .Z(c6743) );
ANDN U33711 ( .B(n20227), .A(n20228), .Z(n20226) );
XOR U33712 ( .A(c6742), .B(b[6742]), .Z(n20227) );
XNOR U33713 ( .A(b[6742]), .B(n20228), .Z(c[6742]) );
XNOR U33714 ( .A(a[6742]), .B(c6742), .Z(n20228) );
XOR U33715 ( .A(c6743), .B(n20229), .Z(c6744) );
ANDN U33716 ( .B(n20230), .A(n20231), .Z(n20229) );
XOR U33717 ( .A(c6743), .B(b[6743]), .Z(n20230) );
XNOR U33718 ( .A(b[6743]), .B(n20231), .Z(c[6743]) );
XNOR U33719 ( .A(a[6743]), .B(c6743), .Z(n20231) );
XOR U33720 ( .A(c6744), .B(n20232), .Z(c6745) );
ANDN U33721 ( .B(n20233), .A(n20234), .Z(n20232) );
XOR U33722 ( .A(c6744), .B(b[6744]), .Z(n20233) );
XNOR U33723 ( .A(b[6744]), .B(n20234), .Z(c[6744]) );
XNOR U33724 ( .A(a[6744]), .B(c6744), .Z(n20234) );
XOR U33725 ( .A(c6745), .B(n20235), .Z(c6746) );
ANDN U33726 ( .B(n20236), .A(n20237), .Z(n20235) );
XOR U33727 ( .A(c6745), .B(b[6745]), .Z(n20236) );
XNOR U33728 ( .A(b[6745]), .B(n20237), .Z(c[6745]) );
XNOR U33729 ( .A(a[6745]), .B(c6745), .Z(n20237) );
XOR U33730 ( .A(c6746), .B(n20238), .Z(c6747) );
ANDN U33731 ( .B(n20239), .A(n20240), .Z(n20238) );
XOR U33732 ( .A(c6746), .B(b[6746]), .Z(n20239) );
XNOR U33733 ( .A(b[6746]), .B(n20240), .Z(c[6746]) );
XNOR U33734 ( .A(a[6746]), .B(c6746), .Z(n20240) );
XOR U33735 ( .A(c6747), .B(n20241), .Z(c6748) );
ANDN U33736 ( .B(n20242), .A(n20243), .Z(n20241) );
XOR U33737 ( .A(c6747), .B(b[6747]), .Z(n20242) );
XNOR U33738 ( .A(b[6747]), .B(n20243), .Z(c[6747]) );
XNOR U33739 ( .A(a[6747]), .B(c6747), .Z(n20243) );
XOR U33740 ( .A(c6748), .B(n20244), .Z(c6749) );
ANDN U33741 ( .B(n20245), .A(n20246), .Z(n20244) );
XOR U33742 ( .A(c6748), .B(b[6748]), .Z(n20245) );
XNOR U33743 ( .A(b[6748]), .B(n20246), .Z(c[6748]) );
XNOR U33744 ( .A(a[6748]), .B(c6748), .Z(n20246) );
XOR U33745 ( .A(c6749), .B(n20247), .Z(c6750) );
ANDN U33746 ( .B(n20248), .A(n20249), .Z(n20247) );
XOR U33747 ( .A(c6749), .B(b[6749]), .Z(n20248) );
XNOR U33748 ( .A(b[6749]), .B(n20249), .Z(c[6749]) );
XNOR U33749 ( .A(a[6749]), .B(c6749), .Z(n20249) );
XOR U33750 ( .A(c6750), .B(n20250), .Z(c6751) );
ANDN U33751 ( .B(n20251), .A(n20252), .Z(n20250) );
XOR U33752 ( .A(c6750), .B(b[6750]), .Z(n20251) );
XNOR U33753 ( .A(b[6750]), .B(n20252), .Z(c[6750]) );
XNOR U33754 ( .A(a[6750]), .B(c6750), .Z(n20252) );
XOR U33755 ( .A(c6751), .B(n20253), .Z(c6752) );
ANDN U33756 ( .B(n20254), .A(n20255), .Z(n20253) );
XOR U33757 ( .A(c6751), .B(b[6751]), .Z(n20254) );
XNOR U33758 ( .A(b[6751]), .B(n20255), .Z(c[6751]) );
XNOR U33759 ( .A(a[6751]), .B(c6751), .Z(n20255) );
XOR U33760 ( .A(c6752), .B(n20256), .Z(c6753) );
ANDN U33761 ( .B(n20257), .A(n20258), .Z(n20256) );
XOR U33762 ( .A(c6752), .B(b[6752]), .Z(n20257) );
XNOR U33763 ( .A(b[6752]), .B(n20258), .Z(c[6752]) );
XNOR U33764 ( .A(a[6752]), .B(c6752), .Z(n20258) );
XOR U33765 ( .A(c6753), .B(n20259), .Z(c6754) );
ANDN U33766 ( .B(n20260), .A(n20261), .Z(n20259) );
XOR U33767 ( .A(c6753), .B(b[6753]), .Z(n20260) );
XNOR U33768 ( .A(b[6753]), .B(n20261), .Z(c[6753]) );
XNOR U33769 ( .A(a[6753]), .B(c6753), .Z(n20261) );
XOR U33770 ( .A(c6754), .B(n20262), .Z(c6755) );
ANDN U33771 ( .B(n20263), .A(n20264), .Z(n20262) );
XOR U33772 ( .A(c6754), .B(b[6754]), .Z(n20263) );
XNOR U33773 ( .A(b[6754]), .B(n20264), .Z(c[6754]) );
XNOR U33774 ( .A(a[6754]), .B(c6754), .Z(n20264) );
XOR U33775 ( .A(c6755), .B(n20265), .Z(c6756) );
ANDN U33776 ( .B(n20266), .A(n20267), .Z(n20265) );
XOR U33777 ( .A(c6755), .B(b[6755]), .Z(n20266) );
XNOR U33778 ( .A(b[6755]), .B(n20267), .Z(c[6755]) );
XNOR U33779 ( .A(a[6755]), .B(c6755), .Z(n20267) );
XOR U33780 ( .A(c6756), .B(n20268), .Z(c6757) );
ANDN U33781 ( .B(n20269), .A(n20270), .Z(n20268) );
XOR U33782 ( .A(c6756), .B(b[6756]), .Z(n20269) );
XNOR U33783 ( .A(b[6756]), .B(n20270), .Z(c[6756]) );
XNOR U33784 ( .A(a[6756]), .B(c6756), .Z(n20270) );
XOR U33785 ( .A(c6757), .B(n20271), .Z(c6758) );
ANDN U33786 ( .B(n20272), .A(n20273), .Z(n20271) );
XOR U33787 ( .A(c6757), .B(b[6757]), .Z(n20272) );
XNOR U33788 ( .A(b[6757]), .B(n20273), .Z(c[6757]) );
XNOR U33789 ( .A(a[6757]), .B(c6757), .Z(n20273) );
XOR U33790 ( .A(c6758), .B(n20274), .Z(c6759) );
ANDN U33791 ( .B(n20275), .A(n20276), .Z(n20274) );
XOR U33792 ( .A(c6758), .B(b[6758]), .Z(n20275) );
XNOR U33793 ( .A(b[6758]), .B(n20276), .Z(c[6758]) );
XNOR U33794 ( .A(a[6758]), .B(c6758), .Z(n20276) );
XOR U33795 ( .A(c6759), .B(n20277), .Z(c6760) );
ANDN U33796 ( .B(n20278), .A(n20279), .Z(n20277) );
XOR U33797 ( .A(c6759), .B(b[6759]), .Z(n20278) );
XNOR U33798 ( .A(b[6759]), .B(n20279), .Z(c[6759]) );
XNOR U33799 ( .A(a[6759]), .B(c6759), .Z(n20279) );
XOR U33800 ( .A(c6760), .B(n20280), .Z(c6761) );
ANDN U33801 ( .B(n20281), .A(n20282), .Z(n20280) );
XOR U33802 ( .A(c6760), .B(b[6760]), .Z(n20281) );
XNOR U33803 ( .A(b[6760]), .B(n20282), .Z(c[6760]) );
XNOR U33804 ( .A(a[6760]), .B(c6760), .Z(n20282) );
XOR U33805 ( .A(c6761), .B(n20283), .Z(c6762) );
ANDN U33806 ( .B(n20284), .A(n20285), .Z(n20283) );
XOR U33807 ( .A(c6761), .B(b[6761]), .Z(n20284) );
XNOR U33808 ( .A(b[6761]), .B(n20285), .Z(c[6761]) );
XNOR U33809 ( .A(a[6761]), .B(c6761), .Z(n20285) );
XOR U33810 ( .A(c6762), .B(n20286), .Z(c6763) );
ANDN U33811 ( .B(n20287), .A(n20288), .Z(n20286) );
XOR U33812 ( .A(c6762), .B(b[6762]), .Z(n20287) );
XNOR U33813 ( .A(b[6762]), .B(n20288), .Z(c[6762]) );
XNOR U33814 ( .A(a[6762]), .B(c6762), .Z(n20288) );
XOR U33815 ( .A(c6763), .B(n20289), .Z(c6764) );
ANDN U33816 ( .B(n20290), .A(n20291), .Z(n20289) );
XOR U33817 ( .A(c6763), .B(b[6763]), .Z(n20290) );
XNOR U33818 ( .A(b[6763]), .B(n20291), .Z(c[6763]) );
XNOR U33819 ( .A(a[6763]), .B(c6763), .Z(n20291) );
XOR U33820 ( .A(c6764), .B(n20292), .Z(c6765) );
ANDN U33821 ( .B(n20293), .A(n20294), .Z(n20292) );
XOR U33822 ( .A(c6764), .B(b[6764]), .Z(n20293) );
XNOR U33823 ( .A(b[6764]), .B(n20294), .Z(c[6764]) );
XNOR U33824 ( .A(a[6764]), .B(c6764), .Z(n20294) );
XOR U33825 ( .A(c6765), .B(n20295), .Z(c6766) );
ANDN U33826 ( .B(n20296), .A(n20297), .Z(n20295) );
XOR U33827 ( .A(c6765), .B(b[6765]), .Z(n20296) );
XNOR U33828 ( .A(b[6765]), .B(n20297), .Z(c[6765]) );
XNOR U33829 ( .A(a[6765]), .B(c6765), .Z(n20297) );
XOR U33830 ( .A(c6766), .B(n20298), .Z(c6767) );
ANDN U33831 ( .B(n20299), .A(n20300), .Z(n20298) );
XOR U33832 ( .A(c6766), .B(b[6766]), .Z(n20299) );
XNOR U33833 ( .A(b[6766]), .B(n20300), .Z(c[6766]) );
XNOR U33834 ( .A(a[6766]), .B(c6766), .Z(n20300) );
XOR U33835 ( .A(c6767), .B(n20301), .Z(c6768) );
ANDN U33836 ( .B(n20302), .A(n20303), .Z(n20301) );
XOR U33837 ( .A(c6767), .B(b[6767]), .Z(n20302) );
XNOR U33838 ( .A(b[6767]), .B(n20303), .Z(c[6767]) );
XNOR U33839 ( .A(a[6767]), .B(c6767), .Z(n20303) );
XOR U33840 ( .A(c6768), .B(n20304), .Z(c6769) );
ANDN U33841 ( .B(n20305), .A(n20306), .Z(n20304) );
XOR U33842 ( .A(c6768), .B(b[6768]), .Z(n20305) );
XNOR U33843 ( .A(b[6768]), .B(n20306), .Z(c[6768]) );
XNOR U33844 ( .A(a[6768]), .B(c6768), .Z(n20306) );
XOR U33845 ( .A(c6769), .B(n20307), .Z(c6770) );
ANDN U33846 ( .B(n20308), .A(n20309), .Z(n20307) );
XOR U33847 ( .A(c6769), .B(b[6769]), .Z(n20308) );
XNOR U33848 ( .A(b[6769]), .B(n20309), .Z(c[6769]) );
XNOR U33849 ( .A(a[6769]), .B(c6769), .Z(n20309) );
XOR U33850 ( .A(c6770), .B(n20310), .Z(c6771) );
ANDN U33851 ( .B(n20311), .A(n20312), .Z(n20310) );
XOR U33852 ( .A(c6770), .B(b[6770]), .Z(n20311) );
XNOR U33853 ( .A(b[6770]), .B(n20312), .Z(c[6770]) );
XNOR U33854 ( .A(a[6770]), .B(c6770), .Z(n20312) );
XOR U33855 ( .A(c6771), .B(n20313), .Z(c6772) );
ANDN U33856 ( .B(n20314), .A(n20315), .Z(n20313) );
XOR U33857 ( .A(c6771), .B(b[6771]), .Z(n20314) );
XNOR U33858 ( .A(b[6771]), .B(n20315), .Z(c[6771]) );
XNOR U33859 ( .A(a[6771]), .B(c6771), .Z(n20315) );
XOR U33860 ( .A(c6772), .B(n20316), .Z(c6773) );
ANDN U33861 ( .B(n20317), .A(n20318), .Z(n20316) );
XOR U33862 ( .A(c6772), .B(b[6772]), .Z(n20317) );
XNOR U33863 ( .A(b[6772]), .B(n20318), .Z(c[6772]) );
XNOR U33864 ( .A(a[6772]), .B(c6772), .Z(n20318) );
XOR U33865 ( .A(c6773), .B(n20319), .Z(c6774) );
ANDN U33866 ( .B(n20320), .A(n20321), .Z(n20319) );
XOR U33867 ( .A(c6773), .B(b[6773]), .Z(n20320) );
XNOR U33868 ( .A(b[6773]), .B(n20321), .Z(c[6773]) );
XNOR U33869 ( .A(a[6773]), .B(c6773), .Z(n20321) );
XOR U33870 ( .A(c6774), .B(n20322), .Z(c6775) );
ANDN U33871 ( .B(n20323), .A(n20324), .Z(n20322) );
XOR U33872 ( .A(c6774), .B(b[6774]), .Z(n20323) );
XNOR U33873 ( .A(b[6774]), .B(n20324), .Z(c[6774]) );
XNOR U33874 ( .A(a[6774]), .B(c6774), .Z(n20324) );
XOR U33875 ( .A(c6775), .B(n20325), .Z(c6776) );
ANDN U33876 ( .B(n20326), .A(n20327), .Z(n20325) );
XOR U33877 ( .A(c6775), .B(b[6775]), .Z(n20326) );
XNOR U33878 ( .A(b[6775]), .B(n20327), .Z(c[6775]) );
XNOR U33879 ( .A(a[6775]), .B(c6775), .Z(n20327) );
XOR U33880 ( .A(c6776), .B(n20328), .Z(c6777) );
ANDN U33881 ( .B(n20329), .A(n20330), .Z(n20328) );
XOR U33882 ( .A(c6776), .B(b[6776]), .Z(n20329) );
XNOR U33883 ( .A(b[6776]), .B(n20330), .Z(c[6776]) );
XNOR U33884 ( .A(a[6776]), .B(c6776), .Z(n20330) );
XOR U33885 ( .A(c6777), .B(n20331), .Z(c6778) );
ANDN U33886 ( .B(n20332), .A(n20333), .Z(n20331) );
XOR U33887 ( .A(c6777), .B(b[6777]), .Z(n20332) );
XNOR U33888 ( .A(b[6777]), .B(n20333), .Z(c[6777]) );
XNOR U33889 ( .A(a[6777]), .B(c6777), .Z(n20333) );
XOR U33890 ( .A(c6778), .B(n20334), .Z(c6779) );
ANDN U33891 ( .B(n20335), .A(n20336), .Z(n20334) );
XOR U33892 ( .A(c6778), .B(b[6778]), .Z(n20335) );
XNOR U33893 ( .A(b[6778]), .B(n20336), .Z(c[6778]) );
XNOR U33894 ( .A(a[6778]), .B(c6778), .Z(n20336) );
XOR U33895 ( .A(c6779), .B(n20337), .Z(c6780) );
ANDN U33896 ( .B(n20338), .A(n20339), .Z(n20337) );
XOR U33897 ( .A(c6779), .B(b[6779]), .Z(n20338) );
XNOR U33898 ( .A(b[6779]), .B(n20339), .Z(c[6779]) );
XNOR U33899 ( .A(a[6779]), .B(c6779), .Z(n20339) );
XOR U33900 ( .A(c6780), .B(n20340), .Z(c6781) );
ANDN U33901 ( .B(n20341), .A(n20342), .Z(n20340) );
XOR U33902 ( .A(c6780), .B(b[6780]), .Z(n20341) );
XNOR U33903 ( .A(b[6780]), .B(n20342), .Z(c[6780]) );
XNOR U33904 ( .A(a[6780]), .B(c6780), .Z(n20342) );
XOR U33905 ( .A(c6781), .B(n20343), .Z(c6782) );
ANDN U33906 ( .B(n20344), .A(n20345), .Z(n20343) );
XOR U33907 ( .A(c6781), .B(b[6781]), .Z(n20344) );
XNOR U33908 ( .A(b[6781]), .B(n20345), .Z(c[6781]) );
XNOR U33909 ( .A(a[6781]), .B(c6781), .Z(n20345) );
XOR U33910 ( .A(c6782), .B(n20346), .Z(c6783) );
ANDN U33911 ( .B(n20347), .A(n20348), .Z(n20346) );
XOR U33912 ( .A(c6782), .B(b[6782]), .Z(n20347) );
XNOR U33913 ( .A(b[6782]), .B(n20348), .Z(c[6782]) );
XNOR U33914 ( .A(a[6782]), .B(c6782), .Z(n20348) );
XOR U33915 ( .A(c6783), .B(n20349), .Z(c6784) );
ANDN U33916 ( .B(n20350), .A(n20351), .Z(n20349) );
XOR U33917 ( .A(c6783), .B(b[6783]), .Z(n20350) );
XNOR U33918 ( .A(b[6783]), .B(n20351), .Z(c[6783]) );
XNOR U33919 ( .A(a[6783]), .B(c6783), .Z(n20351) );
XOR U33920 ( .A(c6784), .B(n20352), .Z(c6785) );
ANDN U33921 ( .B(n20353), .A(n20354), .Z(n20352) );
XOR U33922 ( .A(c6784), .B(b[6784]), .Z(n20353) );
XNOR U33923 ( .A(b[6784]), .B(n20354), .Z(c[6784]) );
XNOR U33924 ( .A(a[6784]), .B(c6784), .Z(n20354) );
XOR U33925 ( .A(c6785), .B(n20355), .Z(c6786) );
ANDN U33926 ( .B(n20356), .A(n20357), .Z(n20355) );
XOR U33927 ( .A(c6785), .B(b[6785]), .Z(n20356) );
XNOR U33928 ( .A(b[6785]), .B(n20357), .Z(c[6785]) );
XNOR U33929 ( .A(a[6785]), .B(c6785), .Z(n20357) );
XOR U33930 ( .A(c6786), .B(n20358), .Z(c6787) );
ANDN U33931 ( .B(n20359), .A(n20360), .Z(n20358) );
XOR U33932 ( .A(c6786), .B(b[6786]), .Z(n20359) );
XNOR U33933 ( .A(b[6786]), .B(n20360), .Z(c[6786]) );
XNOR U33934 ( .A(a[6786]), .B(c6786), .Z(n20360) );
XOR U33935 ( .A(c6787), .B(n20361), .Z(c6788) );
ANDN U33936 ( .B(n20362), .A(n20363), .Z(n20361) );
XOR U33937 ( .A(c6787), .B(b[6787]), .Z(n20362) );
XNOR U33938 ( .A(b[6787]), .B(n20363), .Z(c[6787]) );
XNOR U33939 ( .A(a[6787]), .B(c6787), .Z(n20363) );
XOR U33940 ( .A(c6788), .B(n20364), .Z(c6789) );
ANDN U33941 ( .B(n20365), .A(n20366), .Z(n20364) );
XOR U33942 ( .A(c6788), .B(b[6788]), .Z(n20365) );
XNOR U33943 ( .A(b[6788]), .B(n20366), .Z(c[6788]) );
XNOR U33944 ( .A(a[6788]), .B(c6788), .Z(n20366) );
XOR U33945 ( .A(c6789), .B(n20367), .Z(c6790) );
ANDN U33946 ( .B(n20368), .A(n20369), .Z(n20367) );
XOR U33947 ( .A(c6789), .B(b[6789]), .Z(n20368) );
XNOR U33948 ( .A(b[6789]), .B(n20369), .Z(c[6789]) );
XNOR U33949 ( .A(a[6789]), .B(c6789), .Z(n20369) );
XOR U33950 ( .A(c6790), .B(n20370), .Z(c6791) );
ANDN U33951 ( .B(n20371), .A(n20372), .Z(n20370) );
XOR U33952 ( .A(c6790), .B(b[6790]), .Z(n20371) );
XNOR U33953 ( .A(b[6790]), .B(n20372), .Z(c[6790]) );
XNOR U33954 ( .A(a[6790]), .B(c6790), .Z(n20372) );
XOR U33955 ( .A(c6791), .B(n20373), .Z(c6792) );
ANDN U33956 ( .B(n20374), .A(n20375), .Z(n20373) );
XOR U33957 ( .A(c6791), .B(b[6791]), .Z(n20374) );
XNOR U33958 ( .A(b[6791]), .B(n20375), .Z(c[6791]) );
XNOR U33959 ( .A(a[6791]), .B(c6791), .Z(n20375) );
XOR U33960 ( .A(c6792), .B(n20376), .Z(c6793) );
ANDN U33961 ( .B(n20377), .A(n20378), .Z(n20376) );
XOR U33962 ( .A(c6792), .B(b[6792]), .Z(n20377) );
XNOR U33963 ( .A(b[6792]), .B(n20378), .Z(c[6792]) );
XNOR U33964 ( .A(a[6792]), .B(c6792), .Z(n20378) );
XOR U33965 ( .A(c6793), .B(n20379), .Z(c6794) );
ANDN U33966 ( .B(n20380), .A(n20381), .Z(n20379) );
XOR U33967 ( .A(c6793), .B(b[6793]), .Z(n20380) );
XNOR U33968 ( .A(b[6793]), .B(n20381), .Z(c[6793]) );
XNOR U33969 ( .A(a[6793]), .B(c6793), .Z(n20381) );
XOR U33970 ( .A(c6794), .B(n20382), .Z(c6795) );
ANDN U33971 ( .B(n20383), .A(n20384), .Z(n20382) );
XOR U33972 ( .A(c6794), .B(b[6794]), .Z(n20383) );
XNOR U33973 ( .A(b[6794]), .B(n20384), .Z(c[6794]) );
XNOR U33974 ( .A(a[6794]), .B(c6794), .Z(n20384) );
XOR U33975 ( .A(c6795), .B(n20385), .Z(c6796) );
ANDN U33976 ( .B(n20386), .A(n20387), .Z(n20385) );
XOR U33977 ( .A(c6795), .B(b[6795]), .Z(n20386) );
XNOR U33978 ( .A(b[6795]), .B(n20387), .Z(c[6795]) );
XNOR U33979 ( .A(a[6795]), .B(c6795), .Z(n20387) );
XOR U33980 ( .A(c6796), .B(n20388), .Z(c6797) );
ANDN U33981 ( .B(n20389), .A(n20390), .Z(n20388) );
XOR U33982 ( .A(c6796), .B(b[6796]), .Z(n20389) );
XNOR U33983 ( .A(b[6796]), .B(n20390), .Z(c[6796]) );
XNOR U33984 ( .A(a[6796]), .B(c6796), .Z(n20390) );
XOR U33985 ( .A(c6797), .B(n20391), .Z(c6798) );
ANDN U33986 ( .B(n20392), .A(n20393), .Z(n20391) );
XOR U33987 ( .A(c6797), .B(b[6797]), .Z(n20392) );
XNOR U33988 ( .A(b[6797]), .B(n20393), .Z(c[6797]) );
XNOR U33989 ( .A(a[6797]), .B(c6797), .Z(n20393) );
XOR U33990 ( .A(c6798), .B(n20394), .Z(c6799) );
ANDN U33991 ( .B(n20395), .A(n20396), .Z(n20394) );
XOR U33992 ( .A(c6798), .B(b[6798]), .Z(n20395) );
XNOR U33993 ( .A(b[6798]), .B(n20396), .Z(c[6798]) );
XNOR U33994 ( .A(a[6798]), .B(c6798), .Z(n20396) );
XOR U33995 ( .A(c6799), .B(n20397), .Z(c6800) );
ANDN U33996 ( .B(n20398), .A(n20399), .Z(n20397) );
XOR U33997 ( .A(c6799), .B(b[6799]), .Z(n20398) );
XNOR U33998 ( .A(b[6799]), .B(n20399), .Z(c[6799]) );
XNOR U33999 ( .A(a[6799]), .B(c6799), .Z(n20399) );
XOR U34000 ( .A(c6800), .B(n20400), .Z(c6801) );
ANDN U34001 ( .B(n20401), .A(n20402), .Z(n20400) );
XOR U34002 ( .A(c6800), .B(b[6800]), .Z(n20401) );
XNOR U34003 ( .A(b[6800]), .B(n20402), .Z(c[6800]) );
XNOR U34004 ( .A(a[6800]), .B(c6800), .Z(n20402) );
XOR U34005 ( .A(c6801), .B(n20403), .Z(c6802) );
ANDN U34006 ( .B(n20404), .A(n20405), .Z(n20403) );
XOR U34007 ( .A(c6801), .B(b[6801]), .Z(n20404) );
XNOR U34008 ( .A(b[6801]), .B(n20405), .Z(c[6801]) );
XNOR U34009 ( .A(a[6801]), .B(c6801), .Z(n20405) );
XOR U34010 ( .A(c6802), .B(n20406), .Z(c6803) );
ANDN U34011 ( .B(n20407), .A(n20408), .Z(n20406) );
XOR U34012 ( .A(c6802), .B(b[6802]), .Z(n20407) );
XNOR U34013 ( .A(b[6802]), .B(n20408), .Z(c[6802]) );
XNOR U34014 ( .A(a[6802]), .B(c6802), .Z(n20408) );
XOR U34015 ( .A(c6803), .B(n20409), .Z(c6804) );
ANDN U34016 ( .B(n20410), .A(n20411), .Z(n20409) );
XOR U34017 ( .A(c6803), .B(b[6803]), .Z(n20410) );
XNOR U34018 ( .A(b[6803]), .B(n20411), .Z(c[6803]) );
XNOR U34019 ( .A(a[6803]), .B(c6803), .Z(n20411) );
XOR U34020 ( .A(c6804), .B(n20412), .Z(c6805) );
ANDN U34021 ( .B(n20413), .A(n20414), .Z(n20412) );
XOR U34022 ( .A(c6804), .B(b[6804]), .Z(n20413) );
XNOR U34023 ( .A(b[6804]), .B(n20414), .Z(c[6804]) );
XNOR U34024 ( .A(a[6804]), .B(c6804), .Z(n20414) );
XOR U34025 ( .A(c6805), .B(n20415), .Z(c6806) );
ANDN U34026 ( .B(n20416), .A(n20417), .Z(n20415) );
XOR U34027 ( .A(c6805), .B(b[6805]), .Z(n20416) );
XNOR U34028 ( .A(b[6805]), .B(n20417), .Z(c[6805]) );
XNOR U34029 ( .A(a[6805]), .B(c6805), .Z(n20417) );
XOR U34030 ( .A(c6806), .B(n20418), .Z(c6807) );
ANDN U34031 ( .B(n20419), .A(n20420), .Z(n20418) );
XOR U34032 ( .A(c6806), .B(b[6806]), .Z(n20419) );
XNOR U34033 ( .A(b[6806]), .B(n20420), .Z(c[6806]) );
XNOR U34034 ( .A(a[6806]), .B(c6806), .Z(n20420) );
XOR U34035 ( .A(c6807), .B(n20421), .Z(c6808) );
ANDN U34036 ( .B(n20422), .A(n20423), .Z(n20421) );
XOR U34037 ( .A(c6807), .B(b[6807]), .Z(n20422) );
XNOR U34038 ( .A(b[6807]), .B(n20423), .Z(c[6807]) );
XNOR U34039 ( .A(a[6807]), .B(c6807), .Z(n20423) );
XOR U34040 ( .A(c6808), .B(n20424), .Z(c6809) );
ANDN U34041 ( .B(n20425), .A(n20426), .Z(n20424) );
XOR U34042 ( .A(c6808), .B(b[6808]), .Z(n20425) );
XNOR U34043 ( .A(b[6808]), .B(n20426), .Z(c[6808]) );
XNOR U34044 ( .A(a[6808]), .B(c6808), .Z(n20426) );
XOR U34045 ( .A(c6809), .B(n20427), .Z(c6810) );
ANDN U34046 ( .B(n20428), .A(n20429), .Z(n20427) );
XOR U34047 ( .A(c6809), .B(b[6809]), .Z(n20428) );
XNOR U34048 ( .A(b[6809]), .B(n20429), .Z(c[6809]) );
XNOR U34049 ( .A(a[6809]), .B(c6809), .Z(n20429) );
XOR U34050 ( .A(c6810), .B(n20430), .Z(c6811) );
ANDN U34051 ( .B(n20431), .A(n20432), .Z(n20430) );
XOR U34052 ( .A(c6810), .B(b[6810]), .Z(n20431) );
XNOR U34053 ( .A(b[6810]), .B(n20432), .Z(c[6810]) );
XNOR U34054 ( .A(a[6810]), .B(c6810), .Z(n20432) );
XOR U34055 ( .A(c6811), .B(n20433), .Z(c6812) );
ANDN U34056 ( .B(n20434), .A(n20435), .Z(n20433) );
XOR U34057 ( .A(c6811), .B(b[6811]), .Z(n20434) );
XNOR U34058 ( .A(b[6811]), .B(n20435), .Z(c[6811]) );
XNOR U34059 ( .A(a[6811]), .B(c6811), .Z(n20435) );
XOR U34060 ( .A(c6812), .B(n20436), .Z(c6813) );
ANDN U34061 ( .B(n20437), .A(n20438), .Z(n20436) );
XOR U34062 ( .A(c6812), .B(b[6812]), .Z(n20437) );
XNOR U34063 ( .A(b[6812]), .B(n20438), .Z(c[6812]) );
XNOR U34064 ( .A(a[6812]), .B(c6812), .Z(n20438) );
XOR U34065 ( .A(c6813), .B(n20439), .Z(c6814) );
ANDN U34066 ( .B(n20440), .A(n20441), .Z(n20439) );
XOR U34067 ( .A(c6813), .B(b[6813]), .Z(n20440) );
XNOR U34068 ( .A(b[6813]), .B(n20441), .Z(c[6813]) );
XNOR U34069 ( .A(a[6813]), .B(c6813), .Z(n20441) );
XOR U34070 ( .A(c6814), .B(n20442), .Z(c6815) );
ANDN U34071 ( .B(n20443), .A(n20444), .Z(n20442) );
XOR U34072 ( .A(c6814), .B(b[6814]), .Z(n20443) );
XNOR U34073 ( .A(b[6814]), .B(n20444), .Z(c[6814]) );
XNOR U34074 ( .A(a[6814]), .B(c6814), .Z(n20444) );
XOR U34075 ( .A(c6815), .B(n20445), .Z(c6816) );
ANDN U34076 ( .B(n20446), .A(n20447), .Z(n20445) );
XOR U34077 ( .A(c6815), .B(b[6815]), .Z(n20446) );
XNOR U34078 ( .A(b[6815]), .B(n20447), .Z(c[6815]) );
XNOR U34079 ( .A(a[6815]), .B(c6815), .Z(n20447) );
XOR U34080 ( .A(c6816), .B(n20448), .Z(c6817) );
ANDN U34081 ( .B(n20449), .A(n20450), .Z(n20448) );
XOR U34082 ( .A(c6816), .B(b[6816]), .Z(n20449) );
XNOR U34083 ( .A(b[6816]), .B(n20450), .Z(c[6816]) );
XNOR U34084 ( .A(a[6816]), .B(c6816), .Z(n20450) );
XOR U34085 ( .A(c6817), .B(n20451), .Z(c6818) );
ANDN U34086 ( .B(n20452), .A(n20453), .Z(n20451) );
XOR U34087 ( .A(c6817), .B(b[6817]), .Z(n20452) );
XNOR U34088 ( .A(b[6817]), .B(n20453), .Z(c[6817]) );
XNOR U34089 ( .A(a[6817]), .B(c6817), .Z(n20453) );
XOR U34090 ( .A(c6818), .B(n20454), .Z(c6819) );
ANDN U34091 ( .B(n20455), .A(n20456), .Z(n20454) );
XOR U34092 ( .A(c6818), .B(b[6818]), .Z(n20455) );
XNOR U34093 ( .A(b[6818]), .B(n20456), .Z(c[6818]) );
XNOR U34094 ( .A(a[6818]), .B(c6818), .Z(n20456) );
XOR U34095 ( .A(c6819), .B(n20457), .Z(c6820) );
ANDN U34096 ( .B(n20458), .A(n20459), .Z(n20457) );
XOR U34097 ( .A(c6819), .B(b[6819]), .Z(n20458) );
XNOR U34098 ( .A(b[6819]), .B(n20459), .Z(c[6819]) );
XNOR U34099 ( .A(a[6819]), .B(c6819), .Z(n20459) );
XOR U34100 ( .A(c6820), .B(n20460), .Z(c6821) );
ANDN U34101 ( .B(n20461), .A(n20462), .Z(n20460) );
XOR U34102 ( .A(c6820), .B(b[6820]), .Z(n20461) );
XNOR U34103 ( .A(b[6820]), .B(n20462), .Z(c[6820]) );
XNOR U34104 ( .A(a[6820]), .B(c6820), .Z(n20462) );
XOR U34105 ( .A(c6821), .B(n20463), .Z(c6822) );
ANDN U34106 ( .B(n20464), .A(n20465), .Z(n20463) );
XOR U34107 ( .A(c6821), .B(b[6821]), .Z(n20464) );
XNOR U34108 ( .A(b[6821]), .B(n20465), .Z(c[6821]) );
XNOR U34109 ( .A(a[6821]), .B(c6821), .Z(n20465) );
XOR U34110 ( .A(c6822), .B(n20466), .Z(c6823) );
ANDN U34111 ( .B(n20467), .A(n20468), .Z(n20466) );
XOR U34112 ( .A(c6822), .B(b[6822]), .Z(n20467) );
XNOR U34113 ( .A(b[6822]), .B(n20468), .Z(c[6822]) );
XNOR U34114 ( .A(a[6822]), .B(c6822), .Z(n20468) );
XOR U34115 ( .A(c6823), .B(n20469), .Z(c6824) );
ANDN U34116 ( .B(n20470), .A(n20471), .Z(n20469) );
XOR U34117 ( .A(c6823), .B(b[6823]), .Z(n20470) );
XNOR U34118 ( .A(b[6823]), .B(n20471), .Z(c[6823]) );
XNOR U34119 ( .A(a[6823]), .B(c6823), .Z(n20471) );
XOR U34120 ( .A(c6824), .B(n20472), .Z(c6825) );
ANDN U34121 ( .B(n20473), .A(n20474), .Z(n20472) );
XOR U34122 ( .A(c6824), .B(b[6824]), .Z(n20473) );
XNOR U34123 ( .A(b[6824]), .B(n20474), .Z(c[6824]) );
XNOR U34124 ( .A(a[6824]), .B(c6824), .Z(n20474) );
XOR U34125 ( .A(c6825), .B(n20475), .Z(c6826) );
ANDN U34126 ( .B(n20476), .A(n20477), .Z(n20475) );
XOR U34127 ( .A(c6825), .B(b[6825]), .Z(n20476) );
XNOR U34128 ( .A(b[6825]), .B(n20477), .Z(c[6825]) );
XNOR U34129 ( .A(a[6825]), .B(c6825), .Z(n20477) );
XOR U34130 ( .A(c6826), .B(n20478), .Z(c6827) );
ANDN U34131 ( .B(n20479), .A(n20480), .Z(n20478) );
XOR U34132 ( .A(c6826), .B(b[6826]), .Z(n20479) );
XNOR U34133 ( .A(b[6826]), .B(n20480), .Z(c[6826]) );
XNOR U34134 ( .A(a[6826]), .B(c6826), .Z(n20480) );
XOR U34135 ( .A(c6827), .B(n20481), .Z(c6828) );
ANDN U34136 ( .B(n20482), .A(n20483), .Z(n20481) );
XOR U34137 ( .A(c6827), .B(b[6827]), .Z(n20482) );
XNOR U34138 ( .A(b[6827]), .B(n20483), .Z(c[6827]) );
XNOR U34139 ( .A(a[6827]), .B(c6827), .Z(n20483) );
XOR U34140 ( .A(c6828), .B(n20484), .Z(c6829) );
ANDN U34141 ( .B(n20485), .A(n20486), .Z(n20484) );
XOR U34142 ( .A(c6828), .B(b[6828]), .Z(n20485) );
XNOR U34143 ( .A(b[6828]), .B(n20486), .Z(c[6828]) );
XNOR U34144 ( .A(a[6828]), .B(c6828), .Z(n20486) );
XOR U34145 ( .A(c6829), .B(n20487), .Z(c6830) );
ANDN U34146 ( .B(n20488), .A(n20489), .Z(n20487) );
XOR U34147 ( .A(c6829), .B(b[6829]), .Z(n20488) );
XNOR U34148 ( .A(b[6829]), .B(n20489), .Z(c[6829]) );
XNOR U34149 ( .A(a[6829]), .B(c6829), .Z(n20489) );
XOR U34150 ( .A(c6830), .B(n20490), .Z(c6831) );
ANDN U34151 ( .B(n20491), .A(n20492), .Z(n20490) );
XOR U34152 ( .A(c6830), .B(b[6830]), .Z(n20491) );
XNOR U34153 ( .A(b[6830]), .B(n20492), .Z(c[6830]) );
XNOR U34154 ( .A(a[6830]), .B(c6830), .Z(n20492) );
XOR U34155 ( .A(c6831), .B(n20493), .Z(c6832) );
ANDN U34156 ( .B(n20494), .A(n20495), .Z(n20493) );
XOR U34157 ( .A(c6831), .B(b[6831]), .Z(n20494) );
XNOR U34158 ( .A(b[6831]), .B(n20495), .Z(c[6831]) );
XNOR U34159 ( .A(a[6831]), .B(c6831), .Z(n20495) );
XOR U34160 ( .A(c6832), .B(n20496), .Z(c6833) );
ANDN U34161 ( .B(n20497), .A(n20498), .Z(n20496) );
XOR U34162 ( .A(c6832), .B(b[6832]), .Z(n20497) );
XNOR U34163 ( .A(b[6832]), .B(n20498), .Z(c[6832]) );
XNOR U34164 ( .A(a[6832]), .B(c6832), .Z(n20498) );
XOR U34165 ( .A(c6833), .B(n20499), .Z(c6834) );
ANDN U34166 ( .B(n20500), .A(n20501), .Z(n20499) );
XOR U34167 ( .A(c6833), .B(b[6833]), .Z(n20500) );
XNOR U34168 ( .A(b[6833]), .B(n20501), .Z(c[6833]) );
XNOR U34169 ( .A(a[6833]), .B(c6833), .Z(n20501) );
XOR U34170 ( .A(c6834), .B(n20502), .Z(c6835) );
ANDN U34171 ( .B(n20503), .A(n20504), .Z(n20502) );
XOR U34172 ( .A(c6834), .B(b[6834]), .Z(n20503) );
XNOR U34173 ( .A(b[6834]), .B(n20504), .Z(c[6834]) );
XNOR U34174 ( .A(a[6834]), .B(c6834), .Z(n20504) );
XOR U34175 ( .A(c6835), .B(n20505), .Z(c6836) );
ANDN U34176 ( .B(n20506), .A(n20507), .Z(n20505) );
XOR U34177 ( .A(c6835), .B(b[6835]), .Z(n20506) );
XNOR U34178 ( .A(b[6835]), .B(n20507), .Z(c[6835]) );
XNOR U34179 ( .A(a[6835]), .B(c6835), .Z(n20507) );
XOR U34180 ( .A(c6836), .B(n20508), .Z(c6837) );
ANDN U34181 ( .B(n20509), .A(n20510), .Z(n20508) );
XOR U34182 ( .A(c6836), .B(b[6836]), .Z(n20509) );
XNOR U34183 ( .A(b[6836]), .B(n20510), .Z(c[6836]) );
XNOR U34184 ( .A(a[6836]), .B(c6836), .Z(n20510) );
XOR U34185 ( .A(c6837), .B(n20511), .Z(c6838) );
ANDN U34186 ( .B(n20512), .A(n20513), .Z(n20511) );
XOR U34187 ( .A(c6837), .B(b[6837]), .Z(n20512) );
XNOR U34188 ( .A(b[6837]), .B(n20513), .Z(c[6837]) );
XNOR U34189 ( .A(a[6837]), .B(c6837), .Z(n20513) );
XOR U34190 ( .A(c6838), .B(n20514), .Z(c6839) );
ANDN U34191 ( .B(n20515), .A(n20516), .Z(n20514) );
XOR U34192 ( .A(c6838), .B(b[6838]), .Z(n20515) );
XNOR U34193 ( .A(b[6838]), .B(n20516), .Z(c[6838]) );
XNOR U34194 ( .A(a[6838]), .B(c6838), .Z(n20516) );
XOR U34195 ( .A(c6839), .B(n20517), .Z(c6840) );
ANDN U34196 ( .B(n20518), .A(n20519), .Z(n20517) );
XOR U34197 ( .A(c6839), .B(b[6839]), .Z(n20518) );
XNOR U34198 ( .A(b[6839]), .B(n20519), .Z(c[6839]) );
XNOR U34199 ( .A(a[6839]), .B(c6839), .Z(n20519) );
XOR U34200 ( .A(c6840), .B(n20520), .Z(c6841) );
ANDN U34201 ( .B(n20521), .A(n20522), .Z(n20520) );
XOR U34202 ( .A(c6840), .B(b[6840]), .Z(n20521) );
XNOR U34203 ( .A(b[6840]), .B(n20522), .Z(c[6840]) );
XNOR U34204 ( .A(a[6840]), .B(c6840), .Z(n20522) );
XOR U34205 ( .A(c6841), .B(n20523), .Z(c6842) );
ANDN U34206 ( .B(n20524), .A(n20525), .Z(n20523) );
XOR U34207 ( .A(c6841), .B(b[6841]), .Z(n20524) );
XNOR U34208 ( .A(b[6841]), .B(n20525), .Z(c[6841]) );
XNOR U34209 ( .A(a[6841]), .B(c6841), .Z(n20525) );
XOR U34210 ( .A(c6842), .B(n20526), .Z(c6843) );
ANDN U34211 ( .B(n20527), .A(n20528), .Z(n20526) );
XOR U34212 ( .A(c6842), .B(b[6842]), .Z(n20527) );
XNOR U34213 ( .A(b[6842]), .B(n20528), .Z(c[6842]) );
XNOR U34214 ( .A(a[6842]), .B(c6842), .Z(n20528) );
XOR U34215 ( .A(c6843), .B(n20529), .Z(c6844) );
ANDN U34216 ( .B(n20530), .A(n20531), .Z(n20529) );
XOR U34217 ( .A(c6843), .B(b[6843]), .Z(n20530) );
XNOR U34218 ( .A(b[6843]), .B(n20531), .Z(c[6843]) );
XNOR U34219 ( .A(a[6843]), .B(c6843), .Z(n20531) );
XOR U34220 ( .A(c6844), .B(n20532), .Z(c6845) );
ANDN U34221 ( .B(n20533), .A(n20534), .Z(n20532) );
XOR U34222 ( .A(c6844), .B(b[6844]), .Z(n20533) );
XNOR U34223 ( .A(b[6844]), .B(n20534), .Z(c[6844]) );
XNOR U34224 ( .A(a[6844]), .B(c6844), .Z(n20534) );
XOR U34225 ( .A(c6845), .B(n20535), .Z(c6846) );
ANDN U34226 ( .B(n20536), .A(n20537), .Z(n20535) );
XOR U34227 ( .A(c6845), .B(b[6845]), .Z(n20536) );
XNOR U34228 ( .A(b[6845]), .B(n20537), .Z(c[6845]) );
XNOR U34229 ( .A(a[6845]), .B(c6845), .Z(n20537) );
XOR U34230 ( .A(c6846), .B(n20538), .Z(c6847) );
ANDN U34231 ( .B(n20539), .A(n20540), .Z(n20538) );
XOR U34232 ( .A(c6846), .B(b[6846]), .Z(n20539) );
XNOR U34233 ( .A(b[6846]), .B(n20540), .Z(c[6846]) );
XNOR U34234 ( .A(a[6846]), .B(c6846), .Z(n20540) );
XOR U34235 ( .A(c6847), .B(n20541), .Z(c6848) );
ANDN U34236 ( .B(n20542), .A(n20543), .Z(n20541) );
XOR U34237 ( .A(c6847), .B(b[6847]), .Z(n20542) );
XNOR U34238 ( .A(b[6847]), .B(n20543), .Z(c[6847]) );
XNOR U34239 ( .A(a[6847]), .B(c6847), .Z(n20543) );
XOR U34240 ( .A(c6848), .B(n20544), .Z(c6849) );
ANDN U34241 ( .B(n20545), .A(n20546), .Z(n20544) );
XOR U34242 ( .A(c6848), .B(b[6848]), .Z(n20545) );
XNOR U34243 ( .A(b[6848]), .B(n20546), .Z(c[6848]) );
XNOR U34244 ( .A(a[6848]), .B(c6848), .Z(n20546) );
XOR U34245 ( .A(c6849), .B(n20547), .Z(c6850) );
ANDN U34246 ( .B(n20548), .A(n20549), .Z(n20547) );
XOR U34247 ( .A(c6849), .B(b[6849]), .Z(n20548) );
XNOR U34248 ( .A(b[6849]), .B(n20549), .Z(c[6849]) );
XNOR U34249 ( .A(a[6849]), .B(c6849), .Z(n20549) );
XOR U34250 ( .A(c6850), .B(n20550), .Z(c6851) );
ANDN U34251 ( .B(n20551), .A(n20552), .Z(n20550) );
XOR U34252 ( .A(c6850), .B(b[6850]), .Z(n20551) );
XNOR U34253 ( .A(b[6850]), .B(n20552), .Z(c[6850]) );
XNOR U34254 ( .A(a[6850]), .B(c6850), .Z(n20552) );
XOR U34255 ( .A(c6851), .B(n20553), .Z(c6852) );
ANDN U34256 ( .B(n20554), .A(n20555), .Z(n20553) );
XOR U34257 ( .A(c6851), .B(b[6851]), .Z(n20554) );
XNOR U34258 ( .A(b[6851]), .B(n20555), .Z(c[6851]) );
XNOR U34259 ( .A(a[6851]), .B(c6851), .Z(n20555) );
XOR U34260 ( .A(c6852), .B(n20556), .Z(c6853) );
ANDN U34261 ( .B(n20557), .A(n20558), .Z(n20556) );
XOR U34262 ( .A(c6852), .B(b[6852]), .Z(n20557) );
XNOR U34263 ( .A(b[6852]), .B(n20558), .Z(c[6852]) );
XNOR U34264 ( .A(a[6852]), .B(c6852), .Z(n20558) );
XOR U34265 ( .A(c6853), .B(n20559), .Z(c6854) );
ANDN U34266 ( .B(n20560), .A(n20561), .Z(n20559) );
XOR U34267 ( .A(c6853), .B(b[6853]), .Z(n20560) );
XNOR U34268 ( .A(b[6853]), .B(n20561), .Z(c[6853]) );
XNOR U34269 ( .A(a[6853]), .B(c6853), .Z(n20561) );
XOR U34270 ( .A(c6854), .B(n20562), .Z(c6855) );
ANDN U34271 ( .B(n20563), .A(n20564), .Z(n20562) );
XOR U34272 ( .A(c6854), .B(b[6854]), .Z(n20563) );
XNOR U34273 ( .A(b[6854]), .B(n20564), .Z(c[6854]) );
XNOR U34274 ( .A(a[6854]), .B(c6854), .Z(n20564) );
XOR U34275 ( .A(c6855), .B(n20565), .Z(c6856) );
ANDN U34276 ( .B(n20566), .A(n20567), .Z(n20565) );
XOR U34277 ( .A(c6855), .B(b[6855]), .Z(n20566) );
XNOR U34278 ( .A(b[6855]), .B(n20567), .Z(c[6855]) );
XNOR U34279 ( .A(a[6855]), .B(c6855), .Z(n20567) );
XOR U34280 ( .A(c6856), .B(n20568), .Z(c6857) );
ANDN U34281 ( .B(n20569), .A(n20570), .Z(n20568) );
XOR U34282 ( .A(c6856), .B(b[6856]), .Z(n20569) );
XNOR U34283 ( .A(b[6856]), .B(n20570), .Z(c[6856]) );
XNOR U34284 ( .A(a[6856]), .B(c6856), .Z(n20570) );
XOR U34285 ( .A(c6857), .B(n20571), .Z(c6858) );
ANDN U34286 ( .B(n20572), .A(n20573), .Z(n20571) );
XOR U34287 ( .A(c6857), .B(b[6857]), .Z(n20572) );
XNOR U34288 ( .A(b[6857]), .B(n20573), .Z(c[6857]) );
XNOR U34289 ( .A(a[6857]), .B(c6857), .Z(n20573) );
XOR U34290 ( .A(c6858), .B(n20574), .Z(c6859) );
ANDN U34291 ( .B(n20575), .A(n20576), .Z(n20574) );
XOR U34292 ( .A(c6858), .B(b[6858]), .Z(n20575) );
XNOR U34293 ( .A(b[6858]), .B(n20576), .Z(c[6858]) );
XNOR U34294 ( .A(a[6858]), .B(c6858), .Z(n20576) );
XOR U34295 ( .A(c6859), .B(n20577), .Z(c6860) );
ANDN U34296 ( .B(n20578), .A(n20579), .Z(n20577) );
XOR U34297 ( .A(c6859), .B(b[6859]), .Z(n20578) );
XNOR U34298 ( .A(b[6859]), .B(n20579), .Z(c[6859]) );
XNOR U34299 ( .A(a[6859]), .B(c6859), .Z(n20579) );
XOR U34300 ( .A(c6860), .B(n20580), .Z(c6861) );
ANDN U34301 ( .B(n20581), .A(n20582), .Z(n20580) );
XOR U34302 ( .A(c6860), .B(b[6860]), .Z(n20581) );
XNOR U34303 ( .A(b[6860]), .B(n20582), .Z(c[6860]) );
XNOR U34304 ( .A(a[6860]), .B(c6860), .Z(n20582) );
XOR U34305 ( .A(c6861), .B(n20583), .Z(c6862) );
ANDN U34306 ( .B(n20584), .A(n20585), .Z(n20583) );
XOR U34307 ( .A(c6861), .B(b[6861]), .Z(n20584) );
XNOR U34308 ( .A(b[6861]), .B(n20585), .Z(c[6861]) );
XNOR U34309 ( .A(a[6861]), .B(c6861), .Z(n20585) );
XOR U34310 ( .A(c6862), .B(n20586), .Z(c6863) );
ANDN U34311 ( .B(n20587), .A(n20588), .Z(n20586) );
XOR U34312 ( .A(c6862), .B(b[6862]), .Z(n20587) );
XNOR U34313 ( .A(b[6862]), .B(n20588), .Z(c[6862]) );
XNOR U34314 ( .A(a[6862]), .B(c6862), .Z(n20588) );
XOR U34315 ( .A(c6863), .B(n20589), .Z(c6864) );
ANDN U34316 ( .B(n20590), .A(n20591), .Z(n20589) );
XOR U34317 ( .A(c6863), .B(b[6863]), .Z(n20590) );
XNOR U34318 ( .A(b[6863]), .B(n20591), .Z(c[6863]) );
XNOR U34319 ( .A(a[6863]), .B(c6863), .Z(n20591) );
XOR U34320 ( .A(c6864), .B(n20592), .Z(c6865) );
ANDN U34321 ( .B(n20593), .A(n20594), .Z(n20592) );
XOR U34322 ( .A(c6864), .B(b[6864]), .Z(n20593) );
XNOR U34323 ( .A(b[6864]), .B(n20594), .Z(c[6864]) );
XNOR U34324 ( .A(a[6864]), .B(c6864), .Z(n20594) );
XOR U34325 ( .A(c6865), .B(n20595), .Z(c6866) );
ANDN U34326 ( .B(n20596), .A(n20597), .Z(n20595) );
XOR U34327 ( .A(c6865), .B(b[6865]), .Z(n20596) );
XNOR U34328 ( .A(b[6865]), .B(n20597), .Z(c[6865]) );
XNOR U34329 ( .A(a[6865]), .B(c6865), .Z(n20597) );
XOR U34330 ( .A(c6866), .B(n20598), .Z(c6867) );
ANDN U34331 ( .B(n20599), .A(n20600), .Z(n20598) );
XOR U34332 ( .A(c6866), .B(b[6866]), .Z(n20599) );
XNOR U34333 ( .A(b[6866]), .B(n20600), .Z(c[6866]) );
XNOR U34334 ( .A(a[6866]), .B(c6866), .Z(n20600) );
XOR U34335 ( .A(c6867), .B(n20601), .Z(c6868) );
ANDN U34336 ( .B(n20602), .A(n20603), .Z(n20601) );
XOR U34337 ( .A(c6867), .B(b[6867]), .Z(n20602) );
XNOR U34338 ( .A(b[6867]), .B(n20603), .Z(c[6867]) );
XNOR U34339 ( .A(a[6867]), .B(c6867), .Z(n20603) );
XOR U34340 ( .A(c6868), .B(n20604), .Z(c6869) );
ANDN U34341 ( .B(n20605), .A(n20606), .Z(n20604) );
XOR U34342 ( .A(c6868), .B(b[6868]), .Z(n20605) );
XNOR U34343 ( .A(b[6868]), .B(n20606), .Z(c[6868]) );
XNOR U34344 ( .A(a[6868]), .B(c6868), .Z(n20606) );
XOR U34345 ( .A(c6869), .B(n20607), .Z(c6870) );
ANDN U34346 ( .B(n20608), .A(n20609), .Z(n20607) );
XOR U34347 ( .A(c6869), .B(b[6869]), .Z(n20608) );
XNOR U34348 ( .A(b[6869]), .B(n20609), .Z(c[6869]) );
XNOR U34349 ( .A(a[6869]), .B(c6869), .Z(n20609) );
XOR U34350 ( .A(c6870), .B(n20610), .Z(c6871) );
ANDN U34351 ( .B(n20611), .A(n20612), .Z(n20610) );
XOR U34352 ( .A(c6870), .B(b[6870]), .Z(n20611) );
XNOR U34353 ( .A(b[6870]), .B(n20612), .Z(c[6870]) );
XNOR U34354 ( .A(a[6870]), .B(c6870), .Z(n20612) );
XOR U34355 ( .A(c6871), .B(n20613), .Z(c6872) );
ANDN U34356 ( .B(n20614), .A(n20615), .Z(n20613) );
XOR U34357 ( .A(c6871), .B(b[6871]), .Z(n20614) );
XNOR U34358 ( .A(b[6871]), .B(n20615), .Z(c[6871]) );
XNOR U34359 ( .A(a[6871]), .B(c6871), .Z(n20615) );
XOR U34360 ( .A(c6872), .B(n20616), .Z(c6873) );
ANDN U34361 ( .B(n20617), .A(n20618), .Z(n20616) );
XOR U34362 ( .A(c6872), .B(b[6872]), .Z(n20617) );
XNOR U34363 ( .A(b[6872]), .B(n20618), .Z(c[6872]) );
XNOR U34364 ( .A(a[6872]), .B(c6872), .Z(n20618) );
XOR U34365 ( .A(c6873), .B(n20619), .Z(c6874) );
ANDN U34366 ( .B(n20620), .A(n20621), .Z(n20619) );
XOR U34367 ( .A(c6873), .B(b[6873]), .Z(n20620) );
XNOR U34368 ( .A(b[6873]), .B(n20621), .Z(c[6873]) );
XNOR U34369 ( .A(a[6873]), .B(c6873), .Z(n20621) );
XOR U34370 ( .A(c6874), .B(n20622), .Z(c6875) );
ANDN U34371 ( .B(n20623), .A(n20624), .Z(n20622) );
XOR U34372 ( .A(c6874), .B(b[6874]), .Z(n20623) );
XNOR U34373 ( .A(b[6874]), .B(n20624), .Z(c[6874]) );
XNOR U34374 ( .A(a[6874]), .B(c6874), .Z(n20624) );
XOR U34375 ( .A(c6875), .B(n20625), .Z(c6876) );
ANDN U34376 ( .B(n20626), .A(n20627), .Z(n20625) );
XOR U34377 ( .A(c6875), .B(b[6875]), .Z(n20626) );
XNOR U34378 ( .A(b[6875]), .B(n20627), .Z(c[6875]) );
XNOR U34379 ( .A(a[6875]), .B(c6875), .Z(n20627) );
XOR U34380 ( .A(c6876), .B(n20628), .Z(c6877) );
ANDN U34381 ( .B(n20629), .A(n20630), .Z(n20628) );
XOR U34382 ( .A(c6876), .B(b[6876]), .Z(n20629) );
XNOR U34383 ( .A(b[6876]), .B(n20630), .Z(c[6876]) );
XNOR U34384 ( .A(a[6876]), .B(c6876), .Z(n20630) );
XOR U34385 ( .A(c6877), .B(n20631), .Z(c6878) );
ANDN U34386 ( .B(n20632), .A(n20633), .Z(n20631) );
XOR U34387 ( .A(c6877), .B(b[6877]), .Z(n20632) );
XNOR U34388 ( .A(b[6877]), .B(n20633), .Z(c[6877]) );
XNOR U34389 ( .A(a[6877]), .B(c6877), .Z(n20633) );
XOR U34390 ( .A(c6878), .B(n20634), .Z(c6879) );
ANDN U34391 ( .B(n20635), .A(n20636), .Z(n20634) );
XOR U34392 ( .A(c6878), .B(b[6878]), .Z(n20635) );
XNOR U34393 ( .A(b[6878]), .B(n20636), .Z(c[6878]) );
XNOR U34394 ( .A(a[6878]), .B(c6878), .Z(n20636) );
XOR U34395 ( .A(c6879), .B(n20637), .Z(c6880) );
ANDN U34396 ( .B(n20638), .A(n20639), .Z(n20637) );
XOR U34397 ( .A(c6879), .B(b[6879]), .Z(n20638) );
XNOR U34398 ( .A(b[6879]), .B(n20639), .Z(c[6879]) );
XNOR U34399 ( .A(a[6879]), .B(c6879), .Z(n20639) );
XOR U34400 ( .A(c6880), .B(n20640), .Z(c6881) );
ANDN U34401 ( .B(n20641), .A(n20642), .Z(n20640) );
XOR U34402 ( .A(c6880), .B(b[6880]), .Z(n20641) );
XNOR U34403 ( .A(b[6880]), .B(n20642), .Z(c[6880]) );
XNOR U34404 ( .A(a[6880]), .B(c6880), .Z(n20642) );
XOR U34405 ( .A(c6881), .B(n20643), .Z(c6882) );
ANDN U34406 ( .B(n20644), .A(n20645), .Z(n20643) );
XOR U34407 ( .A(c6881), .B(b[6881]), .Z(n20644) );
XNOR U34408 ( .A(b[6881]), .B(n20645), .Z(c[6881]) );
XNOR U34409 ( .A(a[6881]), .B(c6881), .Z(n20645) );
XOR U34410 ( .A(c6882), .B(n20646), .Z(c6883) );
ANDN U34411 ( .B(n20647), .A(n20648), .Z(n20646) );
XOR U34412 ( .A(c6882), .B(b[6882]), .Z(n20647) );
XNOR U34413 ( .A(b[6882]), .B(n20648), .Z(c[6882]) );
XNOR U34414 ( .A(a[6882]), .B(c6882), .Z(n20648) );
XOR U34415 ( .A(c6883), .B(n20649), .Z(c6884) );
ANDN U34416 ( .B(n20650), .A(n20651), .Z(n20649) );
XOR U34417 ( .A(c6883), .B(b[6883]), .Z(n20650) );
XNOR U34418 ( .A(b[6883]), .B(n20651), .Z(c[6883]) );
XNOR U34419 ( .A(a[6883]), .B(c6883), .Z(n20651) );
XOR U34420 ( .A(c6884), .B(n20652), .Z(c6885) );
ANDN U34421 ( .B(n20653), .A(n20654), .Z(n20652) );
XOR U34422 ( .A(c6884), .B(b[6884]), .Z(n20653) );
XNOR U34423 ( .A(b[6884]), .B(n20654), .Z(c[6884]) );
XNOR U34424 ( .A(a[6884]), .B(c6884), .Z(n20654) );
XOR U34425 ( .A(c6885), .B(n20655), .Z(c6886) );
ANDN U34426 ( .B(n20656), .A(n20657), .Z(n20655) );
XOR U34427 ( .A(c6885), .B(b[6885]), .Z(n20656) );
XNOR U34428 ( .A(b[6885]), .B(n20657), .Z(c[6885]) );
XNOR U34429 ( .A(a[6885]), .B(c6885), .Z(n20657) );
XOR U34430 ( .A(c6886), .B(n20658), .Z(c6887) );
ANDN U34431 ( .B(n20659), .A(n20660), .Z(n20658) );
XOR U34432 ( .A(c6886), .B(b[6886]), .Z(n20659) );
XNOR U34433 ( .A(b[6886]), .B(n20660), .Z(c[6886]) );
XNOR U34434 ( .A(a[6886]), .B(c6886), .Z(n20660) );
XOR U34435 ( .A(c6887), .B(n20661), .Z(c6888) );
ANDN U34436 ( .B(n20662), .A(n20663), .Z(n20661) );
XOR U34437 ( .A(c6887), .B(b[6887]), .Z(n20662) );
XNOR U34438 ( .A(b[6887]), .B(n20663), .Z(c[6887]) );
XNOR U34439 ( .A(a[6887]), .B(c6887), .Z(n20663) );
XOR U34440 ( .A(c6888), .B(n20664), .Z(c6889) );
ANDN U34441 ( .B(n20665), .A(n20666), .Z(n20664) );
XOR U34442 ( .A(c6888), .B(b[6888]), .Z(n20665) );
XNOR U34443 ( .A(b[6888]), .B(n20666), .Z(c[6888]) );
XNOR U34444 ( .A(a[6888]), .B(c6888), .Z(n20666) );
XOR U34445 ( .A(c6889), .B(n20667), .Z(c6890) );
ANDN U34446 ( .B(n20668), .A(n20669), .Z(n20667) );
XOR U34447 ( .A(c6889), .B(b[6889]), .Z(n20668) );
XNOR U34448 ( .A(b[6889]), .B(n20669), .Z(c[6889]) );
XNOR U34449 ( .A(a[6889]), .B(c6889), .Z(n20669) );
XOR U34450 ( .A(c6890), .B(n20670), .Z(c6891) );
ANDN U34451 ( .B(n20671), .A(n20672), .Z(n20670) );
XOR U34452 ( .A(c6890), .B(b[6890]), .Z(n20671) );
XNOR U34453 ( .A(b[6890]), .B(n20672), .Z(c[6890]) );
XNOR U34454 ( .A(a[6890]), .B(c6890), .Z(n20672) );
XOR U34455 ( .A(c6891), .B(n20673), .Z(c6892) );
ANDN U34456 ( .B(n20674), .A(n20675), .Z(n20673) );
XOR U34457 ( .A(c6891), .B(b[6891]), .Z(n20674) );
XNOR U34458 ( .A(b[6891]), .B(n20675), .Z(c[6891]) );
XNOR U34459 ( .A(a[6891]), .B(c6891), .Z(n20675) );
XOR U34460 ( .A(c6892), .B(n20676), .Z(c6893) );
ANDN U34461 ( .B(n20677), .A(n20678), .Z(n20676) );
XOR U34462 ( .A(c6892), .B(b[6892]), .Z(n20677) );
XNOR U34463 ( .A(b[6892]), .B(n20678), .Z(c[6892]) );
XNOR U34464 ( .A(a[6892]), .B(c6892), .Z(n20678) );
XOR U34465 ( .A(c6893), .B(n20679), .Z(c6894) );
ANDN U34466 ( .B(n20680), .A(n20681), .Z(n20679) );
XOR U34467 ( .A(c6893), .B(b[6893]), .Z(n20680) );
XNOR U34468 ( .A(b[6893]), .B(n20681), .Z(c[6893]) );
XNOR U34469 ( .A(a[6893]), .B(c6893), .Z(n20681) );
XOR U34470 ( .A(c6894), .B(n20682), .Z(c6895) );
ANDN U34471 ( .B(n20683), .A(n20684), .Z(n20682) );
XOR U34472 ( .A(c6894), .B(b[6894]), .Z(n20683) );
XNOR U34473 ( .A(b[6894]), .B(n20684), .Z(c[6894]) );
XNOR U34474 ( .A(a[6894]), .B(c6894), .Z(n20684) );
XOR U34475 ( .A(c6895), .B(n20685), .Z(c6896) );
ANDN U34476 ( .B(n20686), .A(n20687), .Z(n20685) );
XOR U34477 ( .A(c6895), .B(b[6895]), .Z(n20686) );
XNOR U34478 ( .A(b[6895]), .B(n20687), .Z(c[6895]) );
XNOR U34479 ( .A(a[6895]), .B(c6895), .Z(n20687) );
XOR U34480 ( .A(c6896), .B(n20688), .Z(c6897) );
ANDN U34481 ( .B(n20689), .A(n20690), .Z(n20688) );
XOR U34482 ( .A(c6896), .B(b[6896]), .Z(n20689) );
XNOR U34483 ( .A(b[6896]), .B(n20690), .Z(c[6896]) );
XNOR U34484 ( .A(a[6896]), .B(c6896), .Z(n20690) );
XOR U34485 ( .A(c6897), .B(n20691), .Z(c6898) );
ANDN U34486 ( .B(n20692), .A(n20693), .Z(n20691) );
XOR U34487 ( .A(c6897), .B(b[6897]), .Z(n20692) );
XNOR U34488 ( .A(b[6897]), .B(n20693), .Z(c[6897]) );
XNOR U34489 ( .A(a[6897]), .B(c6897), .Z(n20693) );
XOR U34490 ( .A(c6898), .B(n20694), .Z(c6899) );
ANDN U34491 ( .B(n20695), .A(n20696), .Z(n20694) );
XOR U34492 ( .A(c6898), .B(b[6898]), .Z(n20695) );
XNOR U34493 ( .A(b[6898]), .B(n20696), .Z(c[6898]) );
XNOR U34494 ( .A(a[6898]), .B(c6898), .Z(n20696) );
XOR U34495 ( .A(c6899), .B(n20697), .Z(c6900) );
ANDN U34496 ( .B(n20698), .A(n20699), .Z(n20697) );
XOR U34497 ( .A(c6899), .B(b[6899]), .Z(n20698) );
XNOR U34498 ( .A(b[6899]), .B(n20699), .Z(c[6899]) );
XNOR U34499 ( .A(a[6899]), .B(c6899), .Z(n20699) );
XOR U34500 ( .A(c6900), .B(n20700), .Z(c6901) );
ANDN U34501 ( .B(n20701), .A(n20702), .Z(n20700) );
XOR U34502 ( .A(c6900), .B(b[6900]), .Z(n20701) );
XNOR U34503 ( .A(b[6900]), .B(n20702), .Z(c[6900]) );
XNOR U34504 ( .A(a[6900]), .B(c6900), .Z(n20702) );
XOR U34505 ( .A(c6901), .B(n20703), .Z(c6902) );
ANDN U34506 ( .B(n20704), .A(n20705), .Z(n20703) );
XOR U34507 ( .A(c6901), .B(b[6901]), .Z(n20704) );
XNOR U34508 ( .A(b[6901]), .B(n20705), .Z(c[6901]) );
XNOR U34509 ( .A(a[6901]), .B(c6901), .Z(n20705) );
XOR U34510 ( .A(c6902), .B(n20706), .Z(c6903) );
ANDN U34511 ( .B(n20707), .A(n20708), .Z(n20706) );
XOR U34512 ( .A(c6902), .B(b[6902]), .Z(n20707) );
XNOR U34513 ( .A(b[6902]), .B(n20708), .Z(c[6902]) );
XNOR U34514 ( .A(a[6902]), .B(c6902), .Z(n20708) );
XOR U34515 ( .A(c6903), .B(n20709), .Z(c6904) );
ANDN U34516 ( .B(n20710), .A(n20711), .Z(n20709) );
XOR U34517 ( .A(c6903), .B(b[6903]), .Z(n20710) );
XNOR U34518 ( .A(b[6903]), .B(n20711), .Z(c[6903]) );
XNOR U34519 ( .A(a[6903]), .B(c6903), .Z(n20711) );
XOR U34520 ( .A(c6904), .B(n20712), .Z(c6905) );
ANDN U34521 ( .B(n20713), .A(n20714), .Z(n20712) );
XOR U34522 ( .A(c6904), .B(b[6904]), .Z(n20713) );
XNOR U34523 ( .A(b[6904]), .B(n20714), .Z(c[6904]) );
XNOR U34524 ( .A(a[6904]), .B(c6904), .Z(n20714) );
XOR U34525 ( .A(c6905), .B(n20715), .Z(c6906) );
ANDN U34526 ( .B(n20716), .A(n20717), .Z(n20715) );
XOR U34527 ( .A(c6905), .B(b[6905]), .Z(n20716) );
XNOR U34528 ( .A(b[6905]), .B(n20717), .Z(c[6905]) );
XNOR U34529 ( .A(a[6905]), .B(c6905), .Z(n20717) );
XOR U34530 ( .A(c6906), .B(n20718), .Z(c6907) );
ANDN U34531 ( .B(n20719), .A(n20720), .Z(n20718) );
XOR U34532 ( .A(c6906), .B(b[6906]), .Z(n20719) );
XNOR U34533 ( .A(b[6906]), .B(n20720), .Z(c[6906]) );
XNOR U34534 ( .A(a[6906]), .B(c6906), .Z(n20720) );
XOR U34535 ( .A(c6907), .B(n20721), .Z(c6908) );
ANDN U34536 ( .B(n20722), .A(n20723), .Z(n20721) );
XOR U34537 ( .A(c6907), .B(b[6907]), .Z(n20722) );
XNOR U34538 ( .A(b[6907]), .B(n20723), .Z(c[6907]) );
XNOR U34539 ( .A(a[6907]), .B(c6907), .Z(n20723) );
XOR U34540 ( .A(c6908), .B(n20724), .Z(c6909) );
ANDN U34541 ( .B(n20725), .A(n20726), .Z(n20724) );
XOR U34542 ( .A(c6908), .B(b[6908]), .Z(n20725) );
XNOR U34543 ( .A(b[6908]), .B(n20726), .Z(c[6908]) );
XNOR U34544 ( .A(a[6908]), .B(c6908), .Z(n20726) );
XOR U34545 ( .A(c6909), .B(n20727), .Z(c6910) );
ANDN U34546 ( .B(n20728), .A(n20729), .Z(n20727) );
XOR U34547 ( .A(c6909), .B(b[6909]), .Z(n20728) );
XNOR U34548 ( .A(b[6909]), .B(n20729), .Z(c[6909]) );
XNOR U34549 ( .A(a[6909]), .B(c6909), .Z(n20729) );
XOR U34550 ( .A(c6910), .B(n20730), .Z(c6911) );
ANDN U34551 ( .B(n20731), .A(n20732), .Z(n20730) );
XOR U34552 ( .A(c6910), .B(b[6910]), .Z(n20731) );
XNOR U34553 ( .A(b[6910]), .B(n20732), .Z(c[6910]) );
XNOR U34554 ( .A(a[6910]), .B(c6910), .Z(n20732) );
XOR U34555 ( .A(c6911), .B(n20733), .Z(c6912) );
ANDN U34556 ( .B(n20734), .A(n20735), .Z(n20733) );
XOR U34557 ( .A(c6911), .B(b[6911]), .Z(n20734) );
XNOR U34558 ( .A(b[6911]), .B(n20735), .Z(c[6911]) );
XNOR U34559 ( .A(a[6911]), .B(c6911), .Z(n20735) );
XOR U34560 ( .A(c6912), .B(n20736), .Z(c6913) );
ANDN U34561 ( .B(n20737), .A(n20738), .Z(n20736) );
XOR U34562 ( .A(c6912), .B(b[6912]), .Z(n20737) );
XNOR U34563 ( .A(b[6912]), .B(n20738), .Z(c[6912]) );
XNOR U34564 ( .A(a[6912]), .B(c6912), .Z(n20738) );
XOR U34565 ( .A(c6913), .B(n20739), .Z(c6914) );
ANDN U34566 ( .B(n20740), .A(n20741), .Z(n20739) );
XOR U34567 ( .A(c6913), .B(b[6913]), .Z(n20740) );
XNOR U34568 ( .A(b[6913]), .B(n20741), .Z(c[6913]) );
XNOR U34569 ( .A(a[6913]), .B(c6913), .Z(n20741) );
XOR U34570 ( .A(c6914), .B(n20742), .Z(c6915) );
ANDN U34571 ( .B(n20743), .A(n20744), .Z(n20742) );
XOR U34572 ( .A(c6914), .B(b[6914]), .Z(n20743) );
XNOR U34573 ( .A(b[6914]), .B(n20744), .Z(c[6914]) );
XNOR U34574 ( .A(a[6914]), .B(c6914), .Z(n20744) );
XOR U34575 ( .A(c6915), .B(n20745), .Z(c6916) );
ANDN U34576 ( .B(n20746), .A(n20747), .Z(n20745) );
XOR U34577 ( .A(c6915), .B(b[6915]), .Z(n20746) );
XNOR U34578 ( .A(b[6915]), .B(n20747), .Z(c[6915]) );
XNOR U34579 ( .A(a[6915]), .B(c6915), .Z(n20747) );
XOR U34580 ( .A(c6916), .B(n20748), .Z(c6917) );
ANDN U34581 ( .B(n20749), .A(n20750), .Z(n20748) );
XOR U34582 ( .A(c6916), .B(b[6916]), .Z(n20749) );
XNOR U34583 ( .A(b[6916]), .B(n20750), .Z(c[6916]) );
XNOR U34584 ( .A(a[6916]), .B(c6916), .Z(n20750) );
XOR U34585 ( .A(c6917), .B(n20751), .Z(c6918) );
ANDN U34586 ( .B(n20752), .A(n20753), .Z(n20751) );
XOR U34587 ( .A(c6917), .B(b[6917]), .Z(n20752) );
XNOR U34588 ( .A(b[6917]), .B(n20753), .Z(c[6917]) );
XNOR U34589 ( .A(a[6917]), .B(c6917), .Z(n20753) );
XOR U34590 ( .A(c6918), .B(n20754), .Z(c6919) );
ANDN U34591 ( .B(n20755), .A(n20756), .Z(n20754) );
XOR U34592 ( .A(c6918), .B(b[6918]), .Z(n20755) );
XNOR U34593 ( .A(b[6918]), .B(n20756), .Z(c[6918]) );
XNOR U34594 ( .A(a[6918]), .B(c6918), .Z(n20756) );
XOR U34595 ( .A(c6919), .B(n20757), .Z(c6920) );
ANDN U34596 ( .B(n20758), .A(n20759), .Z(n20757) );
XOR U34597 ( .A(c6919), .B(b[6919]), .Z(n20758) );
XNOR U34598 ( .A(b[6919]), .B(n20759), .Z(c[6919]) );
XNOR U34599 ( .A(a[6919]), .B(c6919), .Z(n20759) );
XOR U34600 ( .A(c6920), .B(n20760), .Z(c6921) );
ANDN U34601 ( .B(n20761), .A(n20762), .Z(n20760) );
XOR U34602 ( .A(c6920), .B(b[6920]), .Z(n20761) );
XNOR U34603 ( .A(b[6920]), .B(n20762), .Z(c[6920]) );
XNOR U34604 ( .A(a[6920]), .B(c6920), .Z(n20762) );
XOR U34605 ( .A(c6921), .B(n20763), .Z(c6922) );
ANDN U34606 ( .B(n20764), .A(n20765), .Z(n20763) );
XOR U34607 ( .A(c6921), .B(b[6921]), .Z(n20764) );
XNOR U34608 ( .A(b[6921]), .B(n20765), .Z(c[6921]) );
XNOR U34609 ( .A(a[6921]), .B(c6921), .Z(n20765) );
XOR U34610 ( .A(c6922), .B(n20766), .Z(c6923) );
ANDN U34611 ( .B(n20767), .A(n20768), .Z(n20766) );
XOR U34612 ( .A(c6922), .B(b[6922]), .Z(n20767) );
XNOR U34613 ( .A(b[6922]), .B(n20768), .Z(c[6922]) );
XNOR U34614 ( .A(a[6922]), .B(c6922), .Z(n20768) );
XOR U34615 ( .A(c6923), .B(n20769), .Z(c6924) );
ANDN U34616 ( .B(n20770), .A(n20771), .Z(n20769) );
XOR U34617 ( .A(c6923), .B(b[6923]), .Z(n20770) );
XNOR U34618 ( .A(b[6923]), .B(n20771), .Z(c[6923]) );
XNOR U34619 ( .A(a[6923]), .B(c6923), .Z(n20771) );
XOR U34620 ( .A(c6924), .B(n20772), .Z(c6925) );
ANDN U34621 ( .B(n20773), .A(n20774), .Z(n20772) );
XOR U34622 ( .A(c6924), .B(b[6924]), .Z(n20773) );
XNOR U34623 ( .A(b[6924]), .B(n20774), .Z(c[6924]) );
XNOR U34624 ( .A(a[6924]), .B(c6924), .Z(n20774) );
XOR U34625 ( .A(c6925), .B(n20775), .Z(c6926) );
ANDN U34626 ( .B(n20776), .A(n20777), .Z(n20775) );
XOR U34627 ( .A(c6925), .B(b[6925]), .Z(n20776) );
XNOR U34628 ( .A(b[6925]), .B(n20777), .Z(c[6925]) );
XNOR U34629 ( .A(a[6925]), .B(c6925), .Z(n20777) );
XOR U34630 ( .A(c6926), .B(n20778), .Z(c6927) );
ANDN U34631 ( .B(n20779), .A(n20780), .Z(n20778) );
XOR U34632 ( .A(c6926), .B(b[6926]), .Z(n20779) );
XNOR U34633 ( .A(b[6926]), .B(n20780), .Z(c[6926]) );
XNOR U34634 ( .A(a[6926]), .B(c6926), .Z(n20780) );
XOR U34635 ( .A(c6927), .B(n20781), .Z(c6928) );
ANDN U34636 ( .B(n20782), .A(n20783), .Z(n20781) );
XOR U34637 ( .A(c6927), .B(b[6927]), .Z(n20782) );
XNOR U34638 ( .A(b[6927]), .B(n20783), .Z(c[6927]) );
XNOR U34639 ( .A(a[6927]), .B(c6927), .Z(n20783) );
XOR U34640 ( .A(c6928), .B(n20784), .Z(c6929) );
ANDN U34641 ( .B(n20785), .A(n20786), .Z(n20784) );
XOR U34642 ( .A(c6928), .B(b[6928]), .Z(n20785) );
XNOR U34643 ( .A(b[6928]), .B(n20786), .Z(c[6928]) );
XNOR U34644 ( .A(a[6928]), .B(c6928), .Z(n20786) );
XOR U34645 ( .A(c6929), .B(n20787), .Z(c6930) );
ANDN U34646 ( .B(n20788), .A(n20789), .Z(n20787) );
XOR U34647 ( .A(c6929), .B(b[6929]), .Z(n20788) );
XNOR U34648 ( .A(b[6929]), .B(n20789), .Z(c[6929]) );
XNOR U34649 ( .A(a[6929]), .B(c6929), .Z(n20789) );
XOR U34650 ( .A(c6930), .B(n20790), .Z(c6931) );
ANDN U34651 ( .B(n20791), .A(n20792), .Z(n20790) );
XOR U34652 ( .A(c6930), .B(b[6930]), .Z(n20791) );
XNOR U34653 ( .A(b[6930]), .B(n20792), .Z(c[6930]) );
XNOR U34654 ( .A(a[6930]), .B(c6930), .Z(n20792) );
XOR U34655 ( .A(c6931), .B(n20793), .Z(c6932) );
ANDN U34656 ( .B(n20794), .A(n20795), .Z(n20793) );
XOR U34657 ( .A(c6931), .B(b[6931]), .Z(n20794) );
XNOR U34658 ( .A(b[6931]), .B(n20795), .Z(c[6931]) );
XNOR U34659 ( .A(a[6931]), .B(c6931), .Z(n20795) );
XOR U34660 ( .A(c6932), .B(n20796), .Z(c6933) );
ANDN U34661 ( .B(n20797), .A(n20798), .Z(n20796) );
XOR U34662 ( .A(c6932), .B(b[6932]), .Z(n20797) );
XNOR U34663 ( .A(b[6932]), .B(n20798), .Z(c[6932]) );
XNOR U34664 ( .A(a[6932]), .B(c6932), .Z(n20798) );
XOR U34665 ( .A(c6933), .B(n20799), .Z(c6934) );
ANDN U34666 ( .B(n20800), .A(n20801), .Z(n20799) );
XOR U34667 ( .A(c6933), .B(b[6933]), .Z(n20800) );
XNOR U34668 ( .A(b[6933]), .B(n20801), .Z(c[6933]) );
XNOR U34669 ( .A(a[6933]), .B(c6933), .Z(n20801) );
XOR U34670 ( .A(c6934), .B(n20802), .Z(c6935) );
ANDN U34671 ( .B(n20803), .A(n20804), .Z(n20802) );
XOR U34672 ( .A(c6934), .B(b[6934]), .Z(n20803) );
XNOR U34673 ( .A(b[6934]), .B(n20804), .Z(c[6934]) );
XNOR U34674 ( .A(a[6934]), .B(c6934), .Z(n20804) );
XOR U34675 ( .A(c6935), .B(n20805), .Z(c6936) );
ANDN U34676 ( .B(n20806), .A(n20807), .Z(n20805) );
XOR U34677 ( .A(c6935), .B(b[6935]), .Z(n20806) );
XNOR U34678 ( .A(b[6935]), .B(n20807), .Z(c[6935]) );
XNOR U34679 ( .A(a[6935]), .B(c6935), .Z(n20807) );
XOR U34680 ( .A(c6936), .B(n20808), .Z(c6937) );
ANDN U34681 ( .B(n20809), .A(n20810), .Z(n20808) );
XOR U34682 ( .A(c6936), .B(b[6936]), .Z(n20809) );
XNOR U34683 ( .A(b[6936]), .B(n20810), .Z(c[6936]) );
XNOR U34684 ( .A(a[6936]), .B(c6936), .Z(n20810) );
XOR U34685 ( .A(c6937), .B(n20811), .Z(c6938) );
ANDN U34686 ( .B(n20812), .A(n20813), .Z(n20811) );
XOR U34687 ( .A(c6937), .B(b[6937]), .Z(n20812) );
XNOR U34688 ( .A(b[6937]), .B(n20813), .Z(c[6937]) );
XNOR U34689 ( .A(a[6937]), .B(c6937), .Z(n20813) );
XOR U34690 ( .A(c6938), .B(n20814), .Z(c6939) );
ANDN U34691 ( .B(n20815), .A(n20816), .Z(n20814) );
XOR U34692 ( .A(c6938), .B(b[6938]), .Z(n20815) );
XNOR U34693 ( .A(b[6938]), .B(n20816), .Z(c[6938]) );
XNOR U34694 ( .A(a[6938]), .B(c6938), .Z(n20816) );
XOR U34695 ( .A(c6939), .B(n20817), .Z(c6940) );
ANDN U34696 ( .B(n20818), .A(n20819), .Z(n20817) );
XOR U34697 ( .A(c6939), .B(b[6939]), .Z(n20818) );
XNOR U34698 ( .A(b[6939]), .B(n20819), .Z(c[6939]) );
XNOR U34699 ( .A(a[6939]), .B(c6939), .Z(n20819) );
XOR U34700 ( .A(c6940), .B(n20820), .Z(c6941) );
ANDN U34701 ( .B(n20821), .A(n20822), .Z(n20820) );
XOR U34702 ( .A(c6940), .B(b[6940]), .Z(n20821) );
XNOR U34703 ( .A(b[6940]), .B(n20822), .Z(c[6940]) );
XNOR U34704 ( .A(a[6940]), .B(c6940), .Z(n20822) );
XOR U34705 ( .A(c6941), .B(n20823), .Z(c6942) );
ANDN U34706 ( .B(n20824), .A(n20825), .Z(n20823) );
XOR U34707 ( .A(c6941), .B(b[6941]), .Z(n20824) );
XNOR U34708 ( .A(b[6941]), .B(n20825), .Z(c[6941]) );
XNOR U34709 ( .A(a[6941]), .B(c6941), .Z(n20825) );
XOR U34710 ( .A(c6942), .B(n20826), .Z(c6943) );
ANDN U34711 ( .B(n20827), .A(n20828), .Z(n20826) );
XOR U34712 ( .A(c6942), .B(b[6942]), .Z(n20827) );
XNOR U34713 ( .A(b[6942]), .B(n20828), .Z(c[6942]) );
XNOR U34714 ( .A(a[6942]), .B(c6942), .Z(n20828) );
XOR U34715 ( .A(c6943), .B(n20829), .Z(c6944) );
ANDN U34716 ( .B(n20830), .A(n20831), .Z(n20829) );
XOR U34717 ( .A(c6943), .B(b[6943]), .Z(n20830) );
XNOR U34718 ( .A(b[6943]), .B(n20831), .Z(c[6943]) );
XNOR U34719 ( .A(a[6943]), .B(c6943), .Z(n20831) );
XOR U34720 ( .A(c6944), .B(n20832), .Z(c6945) );
ANDN U34721 ( .B(n20833), .A(n20834), .Z(n20832) );
XOR U34722 ( .A(c6944), .B(b[6944]), .Z(n20833) );
XNOR U34723 ( .A(b[6944]), .B(n20834), .Z(c[6944]) );
XNOR U34724 ( .A(a[6944]), .B(c6944), .Z(n20834) );
XOR U34725 ( .A(c6945), .B(n20835), .Z(c6946) );
ANDN U34726 ( .B(n20836), .A(n20837), .Z(n20835) );
XOR U34727 ( .A(c6945), .B(b[6945]), .Z(n20836) );
XNOR U34728 ( .A(b[6945]), .B(n20837), .Z(c[6945]) );
XNOR U34729 ( .A(a[6945]), .B(c6945), .Z(n20837) );
XOR U34730 ( .A(c6946), .B(n20838), .Z(c6947) );
ANDN U34731 ( .B(n20839), .A(n20840), .Z(n20838) );
XOR U34732 ( .A(c6946), .B(b[6946]), .Z(n20839) );
XNOR U34733 ( .A(b[6946]), .B(n20840), .Z(c[6946]) );
XNOR U34734 ( .A(a[6946]), .B(c6946), .Z(n20840) );
XOR U34735 ( .A(c6947), .B(n20841), .Z(c6948) );
ANDN U34736 ( .B(n20842), .A(n20843), .Z(n20841) );
XOR U34737 ( .A(c6947), .B(b[6947]), .Z(n20842) );
XNOR U34738 ( .A(b[6947]), .B(n20843), .Z(c[6947]) );
XNOR U34739 ( .A(a[6947]), .B(c6947), .Z(n20843) );
XOR U34740 ( .A(c6948), .B(n20844), .Z(c6949) );
ANDN U34741 ( .B(n20845), .A(n20846), .Z(n20844) );
XOR U34742 ( .A(c6948), .B(b[6948]), .Z(n20845) );
XNOR U34743 ( .A(b[6948]), .B(n20846), .Z(c[6948]) );
XNOR U34744 ( .A(a[6948]), .B(c6948), .Z(n20846) );
XOR U34745 ( .A(c6949), .B(n20847), .Z(c6950) );
ANDN U34746 ( .B(n20848), .A(n20849), .Z(n20847) );
XOR U34747 ( .A(c6949), .B(b[6949]), .Z(n20848) );
XNOR U34748 ( .A(b[6949]), .B(n20849), .Z(c[6949]) );
XNOR U34749 ( .A(a[6949]), .B(c6949), .Z(n20849) );
XOR U34750 ( .A(c6950), .B(n20850), .Z(c6951) );
ANDN U34751 ( .B(n20851), .A(n20852), .Z(n20850) );
XOR U34752 ( .A(c6950), .B(b[6950]), .Z(n20851) );
XNOR U34753 ( .A(b[6950]), .B(n20852), .Z(c[6950]) );
XNOR U34754 ( .A(a[6950]), .B(c6950), .Z(n20852) );
XOR U34755 ( .A(c6951), .B(n20853), .Z(c6952) );
ANDN U34756 ( .B(n20854), .A(n20855), .Z(n20853) );
XOR U34757 ( .A(c6951), .B(b[6951]), .Z(n20854) );
XNOR U34758 ( .A(b[6951]), .B(n20855), .Z(c[6951]) );
XNOR U34759 ( .A(a[6951]), .B(c6951), .Z(n20855) );
XOR U34760 ( .A(c6952), .B(n20856), .Z(c6953) );
ANDN U34761 ( .B(n20857), .A(n20858), .Z(n20856) );
XOR U34762 ( .A(c6952), .B(b[6952]), .Z(n20857) );
XNOR U34763 ( .A(b[6952]), .B(n20858), .Z(c[6952]) );
XNOR U34764 ( .A(a[6952]), .B(c6952), .Z(n20858) );
XOR U34765 ( .A(c6953), .B(n20859), .Z(c6954) );
ANDN U34766 ( .B(n20860), .A(n20861), .Z(n20859) );
XOR U34767 ( .A(c6953), .B(b[6953]), .Z(n20860) );
XNOR U34768 ( .A(b[6953]), .B(n20861), .Z(c[6953]) );
XNOR U34769 ( .A(a[6953]), .B(c6953), .Z(n20861) );
XOR U34770 ( .A(c6954), .B(n20862), .Z(c6955) );
ANDN U34771 ( .B(n20863), .A(n20864), .Z(n20862) );
XOR U34772 ( .A(c6954), .B(b[6954]), .Z(n20863) );
XNOR U34773 ( .A(b[6954]), .B(n20864), .Z(c[6954]) );
XNOR U34774 ( .A(a[6954]), .B(c6954), .Z(n20864) );
XOR U34775 ( .A(c6955), .B(n20865), .Z(c6956) );
ANDN U34776 ( .B(n20866), .A(n20867), .Z(n20865) );
XOR U34777 ( .A(c6955), .B(b[6955]), .Z(n20866) );
XNOR U34778 ( .A(b[6955]), .B(n20867), .Z(c[6955]) );
XNOR U34779 ( .A(a[6955]), .B(c6955), .Z(n20867) );
XOR U34780 ( .A(c6956), .B(n20868), .Z(c6957) );
ANDN U34781 ( .B(n20869), .A(n20870), .Z(n20868) );
XOR U34782 ( .A(c6956), .B(b[6956]), .Z(n20869) );
XNOR U34783 ( .A(b[6956]), .B(n20870), .Z(c[6956]) );
XNOR U34784 ( .A(a[6956]), .B(c6956), .Z(n20870) );
XOR U34785 ( .A(c6957), .B(n20871), .Z(c6958) );
ANDN U34786 ( .B(n20872), .A(n20873), .Z(n20871) );
XOR U34787 ( .A(c6957), .B(b[6957]), .Z(n20872) );
XNOR U34788 ( .A(b[6957]), .B(n20873), .Z(c[6957]) );
XNOR U34789 ( .A(a[6957]), .B(c6957), .Z(n20873) );
XOR U34790 ( .A(c6958), .B(n20874), .Z(c6959) );
ANDN U34791 ( .B(n20875), .A(n20876), .Z(n20874) );
XOR U34792 ( .A(c6958), .B(b[6958]), .Z(n20875) );
XNOR U34793 ( .A(b[6958]), .B(n20876), .Z(c[6958]) );
XNOR U34794 ( .A(a[6958]), .B(c6958), .Z(n20876) );
XOR U34795 ( .A(c6959), .B(n20877), .Z(c6960) );
ANDN U34796 ( .B(n20878), .A(n20879), .Z(n20877) );
XOR U34797 ( .A(c6959), .B(b[6959]), .Z(n20878) );
XNOR U34798 ( .A(b[6959]), .B(n20879), .Z(c[6959]) );
XNOR U34799 ( .A(a[6959]), .B(c6959), .Z(n20879) );
XOR U34800 ( .A(c6960), .B(n20880), .Z(c6961) );
ANDN U34801 ( .B(n20881), .A(n20882), .Z(n20880) );
XOR U34802 ( .A(c6960), .B(b[6960]), .Z(n20881) );
XNOR U34803 ( .A(b[6960]), .B(n20882), .Z(c[6960]) );
XNOR U34804 ( .A(a[6960]), .B(c6960), .Z(n20882) );
XOR U34805 ( .A(c6961), .B(n20883), .Z(c6962) );
ANDN U34806 ( .B(n20884), .A(n20885), .Z(n20883) );
XOR U34807 ( .A(c6961), .B(b[6961]), .Z(n20884) );
XNOR U34808 ( .A(b[6961]), .B(n20885), .Z(c[6961]) );
XNOR U34809 ( .A(a[6961]), .B(c6961), .Z(n20885) );
XOR U34810 ( .A(c6962), .B(n20886), .Z(c6963) );
ANDN U34811 ( .B(n20887), .A(n20888), .Z(n20886) );
XOR U34812 ( .A(c6962), .B(b[6962]), .Z(n20887) );
XNOR U34813 ( .A(b[6962]), .B(n20888), .Z(c[6962]) );
XNOR U34814 ( .A(a[6962]), .B(c6962), .Z(n20888) );
XOR U34815 ( .A(c6963), .B(n20889), .Z(c6964) );
ANDN U34816 ( .B(n20890), .A(n20891), .Z(n20889) );
XOR U34817 ( .A(c6963), .B(b[6963]), .Z(n20890) );
XNOR U34818 ( .A(b[6963]), .B(n20891), .Z(c[6963]) );
XNOR U34819 ( .A(a[6963]), .B(c6963), .Z(n20891) );
XOR U34820 ( .A(c6964), .B(n20892), .Z(c6965) );
ANDN U34821 ( .B(n20893), .A(n20894), .Z(n20892) );
XOR U34822 ( .A(c6964), .B(b[6964]), .Z(n20893) );
XNOR U34823 ( .A(b[6964]), .B(n20894), .Z(c[6964]) );
XNOR U34824 ( .A(a[6964]), .B(c6964), .Z(n20894) );
XOR U34825 ( .A(c6965), .B(n20895), .Z(c6966) );
ANDN U34826 ( .B(n20896), .A(n20897), .Z(n20895) );
XOR U34827 ( .A(c6965), .B(b[6965]), .Z(n20896) );
XNOR U34828 ( .A(b[6965]), .B(n20897), .Z(c[6965]) );
XNOR U34829 ( .A(a[6965]), .B(c6965), .Z(n20897) );
XOR U34830 ( .A(c6966), .B(n20898), .Z(c6967) );
ANDN U34831 ( .B(n20899), .A(n20900), .Z(n20898) );
XOR U34832 ( .A(c6966), .B(b[6966]), .Z(n20899) );
XNOR U34833 ( .A(b[6966]), .B(n20900), .Z(c[6966]) );
XNOR U34834 ( .A(a[6966]), .B(c6966), .Z(n20900) );
XOR U34835 ( .A(c6967), .B(n20901), .Z(c6968) );
ANDN U34836 ( .B(n20902), .A(n20903), .Z(n20901) );
XOR U34837 ( .A(c6967), .B(b[6967]), .Z(n20902) );
XNOR U34838 ( .A(b[6967]), .B(n20903), .Z(c[6967]) );
XNOR U34839 ( .A(a[6967]), .B(c6967), .Z(n20903) );
XOR U34840 ( .A(c6968), .B(n20904), .Z(c6969) );
ANDN U34841 ( .B(n20905), .A(n20906), .Z(n20904) );
XOR U34842 ( .A(c6968), .B(b[6968]), .Z(n20905) );
XNOR U34843 ( .A(b[6968]), .B(n20906), .Z(c[6968]) );
XNOR U34844 ( .A(a[6968]), .B(c6968), .Z(n20906) );
XOR U34845 ( .A(c6969), .B(n20907), .Z(c6970) );
ANDN U34846 ( .B(n20908), .A(n20909), .Z(n20907) );
XOR U34847 ( .A(c6969), .B(b[6969]), .Z(n20908) );
XNOR U34848 ( .A(b[6969]), .B(n20909), .Z(c[6969]) );
XNOR U34849 ( .A(a[6969]), .B(c6969), .Z(n20909) );
XOR U34850 ( .A(c6970), .B(n20910), .Z(c6971) );
ANDN U34851 ( .B(n20911), .A(n20912), .Z(n20910) );
XOR U34852 ( .A(c6970), .B(b[6970]), .Z(n20911) );
XNOR U34853 ( .A(b[6970]), .B(n20912), .Z(c[6970]) );
XNOR U34854 ( .A(a[6970]), .B(c6970), .Z(n20912) );
XOR U34855 ( .A(c6971), .B(n20913), .Z(c6972) );
ANDN U34856 ( .B(n20914), .A(n20915), .Z(n20913) );
XOR U34857 ( .A(c6971), .B(b[6971]), .Z(n20914) );
XNOR U34858 ( .A(b[6971]), .B(n20915), .Z(c[6971]) );
XNOR U34859 ( .A(a[6971]), .B(c6971), .Z(n20915) );
XOR U34860 ( .A(c6972), .B(n20916), .Z(c6973) );
ANDN U34861 ( .B(n20917), .A(n20918), .Z(n20916) );
XOR U34862 ( .A(c6972), .B(b[6972]), .Z(n20917) );
XNOR U34863 ( .A(b[6972]), .B(n20918), .Z(c[6972]) );
XNOR U34864 ( .A(a[6972]), .B(c6972), .Z(n20918) );
XOR U34865 ( .A(c6973), .B(n20919), .Z(c6974) );
ANDN U34866 ( .B(n20920), .A(n20921), .Z(n20919) );
XOR U34867 ( .A(c6973), .B(b[6973]), .Z(n20920) );
XNOR U34868 ( .A(b[6973]), .B(n20921), .Z(c[6973]) );
XNOR U34869 ( .A(a[6973]), .B(c6973), .Z(n20921) );
XOR U34870 ( .A(c6974), .B(n20922), .Z(c6975) );
ANDN U34871 ( .B(n20923), .A(n20924), .Z(n20922) );
XOR U34872 ( .A(c6974), .B(b[6974]), .Z(n20923) );
XNOR U34873 ( .A(b[6974]), .B(n20924), .Z(c[6974]) );
XNOR U34874 ( .A(a[6974]), .B(c6974), .Z(n20924) );
XOR U34875 ( .A(c6975), .B(n20925), .Z(c6976) );
ANDN U34876 ( .B(n20926), .A(n20927), .Z(n20925) );
XOR U34877 ( .A(c6975), .B(b[6975]), .Z(n20926) );
XNOR U34878 ( .A(b[6975]), .B(n20927), .Z(c[6975]) );
XNOR U34879 ( .A(a[6975]), .B(c6975), .Z(n20927) );
XOR U34880 ( .A(c6976), .B(n20928), .Z(c6977) );
ANDN U34881 ( .B(n20929), .A(n20930), .Z(n20928) );
XOR U34882 ( .A(c6976), .B(b[6976]), .Z(n20929) );
XNOR U34883 ( .A(b[6976]), .B(n20930), .Z(c[6976]) );
XNOR U34884 ( .A(a[6976]), .B(c6976), .Z(n20930) );
XOR U34885 ( .A(c6977), .B(n20931), .Z(c6978) );
ANDN U34886 ( .B(n20932), .A(n20933), .Z(n20931) );
XOR U34887 ( .A(c6977), .B(b[6977]), .Z(n20932) );
XNOR U34888 ( .A(b[6977]), .B(n20933), .Z(c[6977]) );
XNOR U34889 ( .A(a[6977]), .B(c6977), .Z(n20933) );
XOR U34890 ( .A(c6978), .B(n20934), .Z(c6979) );
ANDN U34891 ( .B(n20935), .A(n20936), .Z(n20934) );
XOR U34892 ( .A(c6978), .B(b[6978]), .Z(n20935) );
XNOR U34893 ( .A(b[6978]), .B(n20936), .Z(c[6978]) );
XNOR U34894 ( .A(a[6978]), .B(c6978), .Z(n20936) );
XOR U34895 ( .A(c6979), .B(n20937), .Z(c6980) );
ANDN U34896 ( .B(n20938), .A(n20939), .Z(n20937) );
XOR U34897 ( .A(c6979), .B(b[6979]), .Z(n20938) );
XNOR U34898 ( .A(b[6979]), .B(n20939), .Z(c[6979]) );
XNOR U34899 ( .A(a[6979]), .B(c6979), .Z(n20939) );
XOR U34900 ( .A(c6980), .B(n20940), .Z(c6981) );
ANDN U34901 ( .B(n20941), .A(n20942), .Z(n20940) );
XOR U34902 ( .A(c6980), .B(b[6980]), .Z(n20941) );
XNOR U34903 ( .A(b[6980]), .B(n20942), .Z(c[6980]) );
XNOR U34904 ( .A(a[6980]), .B(c6980), .Z(n20942) );
XOR U34905 ( .A(c6981), .B(n20943), .Z(c6982) );
ANDN U34906 ( .B(n20944), .A(n20945), .Z(n20943) );
XOR U34907 ( .A(c6981), .B(b[6981]), .Z(n20944) );
XNOR U34908 ( .A(b[6981]), .B(n20945), .Z(c[6981]) );
XNOR U34909 ( .A(a[6981]), .B(c6981), .Z(n20945) );
XOR U34910 ( .A(c6982), .B(n20946), .Z(c6983) );
ANDN U34911 ( .B(n20947), .A(n20948), .Z(n20946) );
XOR U34912 ( .A(c6982), .B(b[6982]), .Z(n20947) );
XNOR U34913 ( .A(b[6982]), .B(n20948), .Z(c[6982]) );
XNOR U34914 ( .A(a[6982]), .B(c6982), .Z(n20948) );
XOR U34915 ( .A(c6983), .B(n20949), .Z(c6984) );
ANDN U34916 ( .B(n20950), .A(n20951), .Z(n20949) );
XOR U34917 ( .A(c6983), .B(b[6983]), .Z(n20950) );
XNOR U34918 ( .A(b[6983]), .B(n20951), .Z(c[6983]) );
XNOR U34919 ( .A(a[6983]), .B(c6983), .Z(n20951) );
XOR U34920 ( .A(c6984), .B(n20952), .Z(c6985) );
ANDN U34921 ( .B(n20953), .A(n20954), .Z(n20952) );
XOR U34922 ( .A(c6984), .B(b[6984]), .Z(n20953) );
XNOR U34923 ( .A(b[6984]), .B(n20954), .Z(c[6984]) );
XNOR U34924 ( .A(a[6984]), .B(c6984), .Z(n20954) );
XOR U34925 ( .A(c6985), .B(n20955), .Z(c6986) );
ANDN U34926 ( .B(n20956), .A(n20957), .Z(n20955) );
XOR U34927 ( .A(c6985), .B(b[6985]), .Z(n20956) );
XNOR U34928 ( .A(b[6985]), .B(n20957), .Z(c[6985]) );
XNOR U34929 ( .A(a[6985]), .B(c6985), .Z(n20957) );
XOR U34930 ( .A(c6986), .B(n20958), .Z(c6987) );
ANDN U34931 ( .B(n20959), .A(n20960), .Z(n20958) );
XOR U34932 ( .A(c6986), .B(b[6986]), .Z(n20959) );
XNOR U34933 ( .A(b[6986]), .B(n20960), .Z(c[6986]) );
XNOR U34934 ( .A(a[6986]), .B(c6986), .Z(n20960) );
XOR U34935 ( .A(c6987), .B(n20961), .Z(c6988) );
ANDN U34936 ( .B(n20962), .A(n20963), .Z(n20961) );
XOR U34937 ( .A(c6987), .B(b[6987]), .Z(n20962) );
XNOR U34938 ( .A(b[6987]), .B(n20963), .Z(c[6987]) );
XNOR U34939 ( .A(a[6987]), .B(c6987), .Z(n20963) );
XOR U34940 ( .A(c6988), .B(n20964), .Z(c6989) );
ANDN U34941 ( .B(n20965), .A(n20966), .Z(n20964) );
XOR U34942 ( .A(c6988), .B(b[6988]), .Z(n20965) );
XNOR U34943 ( .A(b[6988]), .B(n20966), .Z(c[6988]) );
XNOR U34944 ( .A(a[6988]), .B(c6988), .Z(n20966) );
XOR U34945 ( .A(c6989), .B(n20967), .Z(c6990) );
ANDN U34946 ( .B(n20968), .A(n20969), .Z(n20967) );
XOR U34947 ( .A(c6989), .B(b[6989]), .Z(n20968) );
XNOR U34948 ( .A(b[6989]), .B(n20969), .Z(c[6989]) );
XNOR U34949 ( .A(a[6989]), .B(c6989), .Z(n20969) );
XOR U34950 ( .A(c6990), .B(n20970), .Z(c6991) );
ANDN U34951 ( .B(n20971), .A(n20972), .Z(n20970) );
XOR U34952 ( .A(c6990), .B(b[6990]), .Z(n20971) );
XNOR U34953 ( .A(b[6990]), .B(n20972), .Z(c[6990]) );
XNOR U34954 ( .A(a[6990]), .B(c6990), .Z(n20972) );
XOR U34955 ( .A(c6991), .B(n20973), .Z(c6992) );
ANDN U34956 ( .B(n20974), .A(n20975), .Z(n20973) );
XOR U34957 ( .A(c6991), .B(b[6991]), .Z(n20974) );
XNOR U34958 ( .A(b[6991]), .B(n20975), .Z(c[6991]) );
XNOR U34959 ( .A(a[6991]), .B(c6991), .Z(n20975) );
XOR U34960 ( .A(c6992), .B(n20976), .Z(c6993) );
ANDN U34961 ( .B(n20977), .A(n20978), .Z(n20976) );
XOR U34962 ( .A(c6992), .B(b[6992]), .Z(n20977) );
XNOR U34963 ( .A(b[6992]), .B(n20978), .Z(c[6992]) );
XNOR U34964 ( .A(a[6992]), .B(c6992), .Z(n20978) );
XOR U34965 ( .A(c6993), .B(n20979), .Z(c6994) );
ANDN U34966 ( .B(n20980), .A(n20981), .Z(n20979) );
XOR U34967 ( .A(c6993), .B(b[6993]), .Z(n20980) );
XNOR U34968 ( .A(b[6993]), .B(n20981), .Z(c[6993]) );
XNOR U34969 ( .A(a[6993]), .B(c6993), .Z(n20981) );
XOR U34970 ( .A(c6994), .B(n20982), .Z(c6995) );
ANDN U34971 ( .B(n20983), .A(n20984), .Z(n20982) );
XOR U34972 ( .A(c6994), .B(b[6994]), .Z(n20983) );
XNOR U34973 ( .A(b[6994]), .B(n20984), .Z(c[6994]) );
XNOR U34974 ( .A(a[6994]), .B(c6994), .Z(n20984) );
XOR U34975 ( .A(c6995), .B(n20985), .Z(c6996) );
ANDN U34976 ( .B(n20986), .A(n20987), .Z(n20985) );
XOR U34977 ( .A(c6995), .B(b[6995]), .Z(n20986) );
XNOR U34978 ( .A(b[6995]), .B(n20987), .Z(c[6995]) );
XNOR U34979 ( .A(a[6995]), .B(c6995), .Z(n20987) );
XOR U34980 ( .A(c6996), .B(n20988), .Z(c6997) );
ANDN U34981 ( .B(n20989), .A(n20990), .Z(n20988) );
XOR U34982 ( .A(c6996), .B(b[6996]), .Z(n20989) );
XNOR U34983 ( .A(b[6996]), .B(n20990), .Z(c[6996]) );
XNOR U34984 ( .A(a[6996]), .B(c6996), .Z(n20990) );
XOR U34985 ( .A(c6997), .B(n20991), .Z(c6998) );
ANDN U34986 ( .B(n20992), .A(n20993), .Z(n20991) );
XOR U34987 ( .A(c6997), .B(b[6997]), .Z(n20992) );
XNOR U34988 ( .A(b[6997]), .B(n20993), .Z(c[6997]) );
XNOR U34989 ( .A(a[6997]), .B(c6997), .Z(n20993) );
XOR U34990 ( .A(c6998), .B(n20994), .Z(c6999) );
ANDN U34991 ( .B(n20995), .A(n20996), .Z(n20994) );
XOR U34992 ( .A(c6998), .B(b[6998]), .Z(n20995) );
XNOR U34993 ( .A(b[6998]), .B(n20996), .Z(c[6998]) );
XNOR U34994 ( .A(a[6998]), .B(c6998), .Z(n20996) );
XOR U34995 ( .A(c6999), .B(n20997), .Z(c7000) );
ANDN U34996 ( .B(n20998), .A(n20999), .Z(n20997) );
XOR U34997 ( .A(c6999), .B(b[6999]), .Z(n20998) );
XNOR U34998 ( .A(b[6999]), .B(n20999), .Z(c[6999]) );
XNOR U34999 ( .A(a[6999]), .B(c6999), .Z(n20999) );
XOR U35000 ( .A(c7000), .B(n21000), .Z(c7001) );
ANDN U35001 ( .B(n21001), .A(n21002), .Z(n21000) );
XOR U35002 ( .A(c7000), .B(b[7000]), .Z(n21001) );
XNOR U35003 ( .A(b[7000]), .B(n21002), .Z(c[7000]) );
XNOR U35004 ( .A(a[7000]), .B(c7000), .Z(n21002) );
XOR U35005 ( .A(c7001), .B(n21003), .Z(c7002) );
ANDN U35006 ( .B(n21004), .A(n21005), .Z(n21003) );
XOR U35007 ( .A(c7001), .B(b[7001]), .Z(n21004) );
XNOR U35008 ( .A(b[7001]), .B(n21005), .Z(c[7001]) );
XNOR U35009 ( .A(a[7001]), .B(c7001), .Z(n21005) );
XOR U35010 ( .A(c7002), .B(n21006), .Z(c7003) );
ANDN U35011 ( .B(n21007), .A(n21008), .Z(n21006) );
XOR U35012 ( .A(c7002), .B(b[7002]), .Z(n21007) );
XNOR U35013 ( .A(b[7002]), .B(n21008), .Z(c[7002]) );
XNOR U35014 ( .A(a[7002]), .B(c7002), .Z(n21008) );
XOR U35015 ( .A(c7003), .B(n21009), .Z(c7004) );
ANDN U35016 ( .B(n21010), .A(n21011), .Z(n21009) );
XOR U35017 ( .A(c7003), .B(b[7003]), .Z(n21010) );
XNOR U35018 ( .A(b[7003]), .B(n21011), .Z(c[7003]) );
XNOR U35019 ( .A(a[7003]), .B(c7003), .Z(n21011) );
XOR U35020 ( .A(c7004), .B(n21012), .Z(c7005) );
ANDN U35021 ( .B(n21013), .A(n21014), .Z(n21012) );
XOR U35022 ( .A(c7004), .B(b[7004]), .Z(n21013) );
XNOR U35023 ( .A(b[7004]), .B(n21014), .Z(c[7004]) );
XNOR U35024 ( .A(a[7004]), .B(c7004), .Z(n21014) );
XOR U35025 ( .A(c7005), .B(n21015), .Z(c7006) );
ANDN U35026 ( .B(n21016), .A(n21017), .Z(n21015) );
XOR U35027 ( .A(c7005), .B(b[7005]), .Z(n21016) );
XNOR U35028 ( .A(b[7005]), .B(n21017), .Z(c[7005]) );
XNOR U35029 ( .A(a[7005]), .B(c7005), .Z(n21017) );
XOR U35030 ( .A(c7006), .B(n21018), .Z(c7007) );
ANDN U35031 ( .B(n21019), .A(n21020), .Z(n21018) );
XOR U35032 ( .A(c7006), .B(b[7006]), .Z(n21019) );
XNOR U35033 ( .A(b[7006]), .B(n21020), .Z(c[7006]) );
XNOR U35034 ( .A(a[7006]), .B(c7006), .Z(n21020) );
XOR U35035 ( .A(c7007), .B(n21021), .Z(c7008) );
ANDN U35036 ( .B(n21022), .A(n21023), .Z(n21021) );
XOR U35037 ( .A(c7007), .B(b[7007]), .Z(n21022) );
XNOR U35038 ( .A(b[7007]), .B(n21023), .Z(c[7007]) );
XNOR U35039 ( .A(a[7007]), .B(c7007), .Z(n21023) );
XOR U35040 ( .A(c7008), .B(n21024), .Z(c7009) );
ANDN U35041 ( .B(n21025), .A(n21026), .Z(n21024) );
XOR U35042 ( .A(c7008), .B(b[7008]), .Z(n21025) );
XNOR U35043 ( .A(b[7008]), .B(n21026), .Z(c[7008]) );
XNOR U35044 ( .A(a[7008]), .B(c7008), .Z(n21026) );
XOR U35045 ( .A(c7009), .B(n21027), .Z(c7010) );
ANDN U35046 ( .B(n21028), .A(n21029), .Z(n21027) );
XOR U35047 ( .A(c7009), .B(b[7009]), .Z(n21028) );
XNOR U35048 ( .A(b[7009]), .B(n21029), .Z(c[7009]) );
XNOR U35049 ( .A(a[7009]), .B(c7009), .Z(n21029) );
XOR U35050 ( .A(c7010), .B(n21030), .Z(c7011) );
ANDN U35051 ( .B(n21031), .A(n21032), .Z(n21030) );
XOR U35052 ( .A(c7010), .B(b[7010]), .Z(n21031) );
XNOR U35053 ( .A(b[7010]), .B(n21032), .Z(c[7010]) );
XNOR U35054 ( .A(a[7010]), .B(c7010), .Z(n21032) );
XOR U35055 ( .A(c7011), .B(n21033), .Z(c7012) );
ANDN U35056 ( .B(n21034), .A(n21035), .Z(n21033) );
XOR U35057 ( .A(c7011), .B(b[7011]), .Z(n21034) );
XNOR U35058 ( .A(b[7011]), .B(n21035), .Z(c[7011]) );
XNOR U35059 ( .A(a[7011]), .B(c7011), .Z(n21035) );
XOR U35060 ( .A(c7012), .B(n21036), .Z(c7013) );
ANDN U35061 ( .B(n21037), .A(n21038), .Z(n21036) );
XOR U35062 ( .A(c7012), .B(b[7012]), .Z(n21037) );
XNOR U35063 ( .A(b[7012]), .B(n21038), .Z(c[7012]) );
XNOR U35064 ( .A(a[7012]), .B(c7012), .Z(n21038) );
XOR U35065 ( .A(c7013), .B(n21039), .Z(c7014) );
ANDN U35066 ( .B(n21040), .A(n21041), .Z(n21039) );
XOR U35067 ( .A(c7013), .B(b[7013]), .Z(n21040) );
XNOR U35068 ( .A(b[7013]), .B(n21041), .Z(c[7013]) );
XNOR U35069 ( .A(a[7013]), .B(c7013), .Z(n21041) );
XOR U35070 ( .A(c7014), .B(n21042), .Z(c7015) );
ANDN U35071 ( .B(n21043), .A(n21044), .Z(n21042) );
XOR U35072 ( .A(c7014), .B(b[7014]), .Z(n21043) );
XNOR U35073 ( .A(b[7014]), .B(n21044), .Z(c[7014]) );
XNOR U35074 ( .A(a[7014]), .B(c7014), .Z(n21044) );
XOR U35075 ( .A(c7015), .B(n21045), .Z(c7016) );
ANDN U35076 ( .B(n21046), .A(n21047), .Z(n21045) );
XOR U35077 ( .A(c7015), .B(b[7015]), .Z(n21046) );
XNOR U35078 ( .A(b[7015]), .B(n21047), .Z(c[7015]) );
XNOR U35079 ( .A(a[7015]), .B(c7015), .Z(n21047) );
XOR U35080 ( .A(c7016), .B(n21048), .Z(c7017) );
ANDN U35081 ( .B(n21049), .A(n21050), .Z(n21048) );
XOR U35082 ( .A(c7016), .B(b[7016]), .Z(n21049) );
XNOR U35083 ( .A(b[7016]), .B(n21050), .Z(c[7016]) );
XNOR U35084 ( .A(a[7016]), .B(c7016), .Z(n21050) );
XOR U35085 ( .A(c7017), .B(n21051), .Z(c7018) );
ANDN U35086 ( .B(n21052), .A(n21053), .Z(n21051) );
XOR U35087 ( .A(c7017), .B(b[7017]), .Z(n21052) );
XNOR U35088 ( .A(b[7017]), .B(n21053), .Z(c[7017]) );
XNOR U35089 ( .A(a[7017]), .B(c7017), .Z(n21053) );
XOR U35090 ( .A(c7018), .B(n21054), .Z(c7019) );
ANDN U35091 ( .B(n21055), .A(n21056), .Z(n21054) );
XOR U35092 ( .A(c7018), .B(b[7018]), .Z(n21055) );
XNOR U35093 ( .A(b[7018]), .B(n21056), .Z(c[7018]) );
XNOR U35094 ( .A(a[7018]), .B(c7018), .Z(n21056) );
XOR U35095 ( .A(c7019), .B(n21057), .Z(c7020) );
ANDN U35096 ( .B(n21058), .A(n21059), .Z(n21057) );
XOR U35097 ( .A(c7019), .B(b[7019]), .Z(n21058) );
XNOR U35098 ( .A(b[7019]), .B(n21059), .Z(c[7019]) );
XNOR U35099 ( .A(a[7019]), .B(c7019), .Z(n21059) );
XOR U35100 ( .A(c7020), .B(n21060), .Z(c7021) );
ANDN U35101 ( .B(n21061), .A(n21062), .Z(n21060) );
XOR U35102 ( .A(c7020), .B(b[7020]), .Z(n21061) );
XNOR U35103 ( .A(b[7020]), .B(n21062), .Z(c[7020]) );
XNOR U35104 ( .A(a[7020]), .B(c7020), .Z(n21062) );
XOR U35105 ( .A(c7021), .B(n21063), .Z(c7022) );
ANDN U35106 ( .B(n21064), .A(n21065), .Z(n21063) );
XOR U35107 ( .A(c7021), .B(b[7021]), .Z(n21064) );
XNOR U35108 ( .A(b[7021]), .B(n21065), .Z(c[7021]) );
XNOR U35109 ( .A(a[7021]), .B(c7021), .Z(n21065) );
XOR U35110 ( .A(c7022), .B(n21066), .Z(c7023) );
ANDN U35111 ( .B(n21067), .A(n21068), .Z(n21066) );
XOR U35112 ( .A(c7022), .B(b[7022]), .Z(n21067) );
XNOR U35113 ( .A(b[7022]), .B(n21068), .Z(c[7022]) );
XNOR U35114 ( .A(a[7022]), .B(c7022), .Z(n21068) );
XOR U35115 ( .A(c7023), .B(n21069), .Z(c7024) );
ANDN U35116 ( .B(n21070), .A(n21071), .Z(n21069) );
XOR U35117 ( .A(c7023), .B(b[7023]), .Z(n21070) );
XNOR U35118 ( .A(b[7023]), .B(n21071), .Z(c[7023]) );
XNOR U35119 ( .A(a[7023]), .B(c7023), .Z(n21071) );
XOR U35120 ( .A(c7024), .B(n21072), .Z(c7025) );
ANDN U35121 ( .B(n21073), .A(n21074), .Z(n21072) );
XOR U35122 ( .A(c7024), .B(b[7024]), .Z(n21073) );
XNOR U35123 ( .A(b[7024]), .B(n21074), .Z(c[7024]) );
XNOR U35124 ( .A(a[7024]), .B(c7024), .Z(n21074) );
XOR U35125 ( .A(c7025), .B(n21075), .Z(c7026) );
ANDN U35126 ( .B(n21076), .A(n21077), .Z(n21075) );
XOR U35127 ( .A(c7025), .B(b[7025]), .Z(n21076) );
XNOR U35128 ( .A(b[7025]), .B(n21077), .Z(c[7025]) );
XNOR U35129 ( .A(a[7025]), .B(c7025), .Z(n21077) );
XOR U35130 ( .A(c7026), .B(n21078), .Z(c7027) );
ANDN U35131 ( .B(n21079), .A(n21080), .Z(n21078) );
XOR U35132 ( .A(c7026), .B(b[7026]), .Z(n21079) );
XNOR U35133 ( .A(b[7026]), .B(n21080), .Z(c[7026]) );
XNOR U35134 ( .A(a[7026]), .B(c7026), .Z(n21080) );
XOR U35135 ( .A(c7027), .B(n21081), .Z(c7028) );
ANDN U35136 ( .B(n21082), .A(n21083), .Z(n21081) );
XOR U35137 ( .A(c7027), .B(b[7027]), .Z(n21082) );
XNOR U35138 ( .A(b[7027]), .B(n21083), .Z(c[7027]) );
XNOR U35139 ( .A(a[7027]), .B(c7027), .Z(n21083) );
XOR U35140 ( .A(c7028), .B(n21084), .Z(c7029) );
ANDN U35141 ( .B(n21085), .A(n21086), .Z(n21084) );
XOR U35142 ( .A(c7028), .B(b[7028]), .Z(n21085) );
XNOR U35143 ( .A(b[7028]), .B(n21086), .Z(c[7028]) );
XNOR U35144 ( .A(a[7028]), .B(c7028), .Z(n21086) );
XOR U35145 ( .A(c7029), .B(n21087), .Z(c7030) );
ANDN U35146 ( .B(n21088), .A(n21089), .Z(n21087) );
XOR U35147 ( .A(c7029), .B(b[7029]), .Z(n21088) );
XNOR U35148 ( .A(b[7029]), .B(n21089), .Z(c[7029]) );
XNOR U35149 ( .A(a[7029]), .B(c7029), .Z(n21089) );
XOR U35150 ( .A(c7030), .B(n21090), .Z(c7031) );
ANDN U35151 ( .B(n21091), .A(n21092), .Z(n21090) );
XOR U35152 ( .A(c7030), .B(b[7030]), .Z(n21091) );
XNOR U35153 ( .A(b[7030]), .B(n21092), .Z(c[7030]) );
XNOR U35154 ( .A(a[7030]), .B(c7030), .Z(n21092) );
XOR U35155 ( .A(c7031), .B(n21093), .Z(c7032) );
ANDN U35156 ( .B(n21094), .A(n21095), .Z(n21093) );
XOR U35157 ( .A(c7031), .B(b[7031]), .Z(n21094) );
XNOR U35158 ( .A(b[7031]), .B(n21095), .Z(c[7031]) );
XNOR U35159 ( .A(a[7031]), .B(c7031), .Z(n21095) );
XOR U35160 ( .A(c7032), .B(n21096), .Z(c7033) );
ANDN U35161 ( .B(n21097), .A(n21098), .Z(n21096) );
XOR U35162 ( .A(c7032), .B(b[7032]), .Z(n21097) );
XNOR U35163 ( .A(b[7032]), .B(n21098), .Z(c[7032]) );
XNOR U35164 ( .A(a[7032]), .B(c7032), .Z(n21098) );
XOR U35165 ( .A(c7033), .B(n21099), .Z(c7034) );
ANDN U35166 ( .B(n21100), .A(n21101), .Z(n21099) );
XOR U35167 ( .A(c7033), .B(b[7033]), .Z(n21100) );
XNOR U35168 ( .A(b[7033]), .B(n21101), .Z(c[7033]) );
XNOR U35169 ( .A(a[7033]), .B(c7033), .Z(n21101) );
XOR U35170 ( .A(c7034), .B(n21102), .Z(c7035) );
ANDN U35171 ( .B(n21103), .A(n21104), .Z(n21102) );
XOR U35172 ( .A(c7034), .B(b[7034]), .Z(n21103) );
XNOR U35173 ( .A(b[7034]), .B(n21104), .Z(c[7034]) );
XNOR U35174 ( .A(a[7034]), .B(c7034), .Z(n21104) );
XOR U35175 ( .A(c7035), .B(n21105), .Z(c7036) );
ANDN U35176 ( .B(n21106), .A(n21107), .Z(n21105) );
XOR U35177 ( .A(c7035), .B(b[7035]), .Z(n21106) );
XNOR U35178 ( .A(b[7035]), .B(n21107), .Z(c[7035]) );
XNOR U35179 ( .A(a[7035]), .B(c7035), .Z(n21107) );
XOR U35180 ( .A(c7036), .B(n21108), .Z(c7037) );
ANDN U35181 ( .B(n21109), .A(n21110), .Z(n21108) );
XOR U35182 ( .A(c7036), .B(b[7036]), .Z(n21109) );
XNOR U35183 ( .A(b[7036]), .B(n21110), .Z(c[7036]) );
XNOR U35184 ( .A(a[7036]), .B(c7036), .Z(n21110) );
XOR U35185 ( .A(c7037), .B(n21111), .Z(c7038) );
ANDN U35186 ( .B(n21112), .A(n21113), .Z(n21111) );
XOR U35187 ( .A(c7037), .B(b[7037]), .Z(n21112) );
XNOR U35188 ( .A(b[7037]), .B(n21113), .Z(c[7037]) );
XNOR U35189 ( .A(a[7037]), .B(c7037), .Z(n21113) );
XOR U35190 ( .A(c7038), .B(n21114), .Z(c7039) );
ANDN U35191 ( .B(n21115), .A(n21116), .Z(n21114) );
XOR U35192 ( .A(c7038), .B(b[7038]), .Z(n21115) );
XNOR U35193 ( .A(b[7038]), .B(n21116), .Z(c[7038]) );
XNOR U35194 ( .A(a[7038]), .B(c7038), .Z(n21116) );
XOR U35195 ( .A(c7039), .B(n21117), .Z(c7040) );
ANDN U35196 ( .B(n21118), .A(n21119), .Z(n21117) );
XOR U35197 ( .A(c7039), .B(b[7039]), .Z(n21118) );
XNOR U35198 ( .A(b[7039]), .B(n21119), .Z(c[7039]) );
XNOR U35199 ( .A(a[7039]), .B(c7039), .Z(n21119) );
XOR U35200 ( .A(c7040), .B(n21120), .Z(c7041) );
ANDN U35201 ( .B(n21121), .A(n21122), .Z(n21120) );
XOR U35202 ( .A(c7040), .B(b[7040]), .Z(n21121) );
XNOR U35203 ( .A(b[7040]), .B(n21122), .Z(c[7040]) );
XNOR U35204 ( .A(a[7040]), .B(c7040), .Z(n21122) );
XOR U35205 ( .A(c7041), .B(n21123), .Z(c7042) );
ANDN U35206 ( .B(n21124), .A(n21125), .Z(n21123) );
XOR U35207 ( .A(c7041), .B(b[7041]), .Z(n21124) );
XNOR U35208 ( .A(b[7041]), .B(n21125), .Z(c[7041]) );
XNOR U35209 ( .A(a[7041]), .B(c7041), .Z(n21125) );
XOR U35210 ( .A(c7042), .B(n21126), .Z(c7043) );
ANDN U35211 ( .B(n21127), .A(n21128), .Z(n21126) );
XOR U35212 ( .A(c7042), .B(b[7042]), .Z(n21127) );
XNOR U35213 ( .A(b[7042]), .B(n21128), .Z(c[7042]) );
XNOR U35214 ( .A(a[7042]), .B(c7042), .Z(n21128) );
XOR U35215 ( .A(c7043), .B(n21129), .Z(c7044) );
ANDN U35216 ( .B(n21130), .A(n21131), .Z(n21129) );
XOR U35217 ( .A(c7043), .B(b[7043]), .Z(n21130) );
XNOR U35218 ( .A(b[7043]), .B(n21131), .Z(c[7043]) );
XNOR U35219 ( .A(a[7043]), .B(c7043), .Z(n21131) );
XOR U35220 ( .A(c7044), .B(n21132), .Z(c7045) );
ANDN U35221 ( .B(n21133), .A(n21134), .Z(n21132) );
XOR U35222 ( .A(c7044), .B(b[7044]), .Z(n21133) );
XNOR U35223 ( .A(b[7044]), .B(n21134), .Z(c[7044]) );
XNOR U35224 ( .A(a[7044]), .B(c7044), .Z(n21134) );
XOR U35225 ( .A(c7045), .B(n21135), .Z(c7046) );
ANDN U35226 ( .B(n21136), .A(n21137), .Z(n21135) );
XOR U35227 ( .A(c7045), .B(b[7045]), .Z(n21136) );
XNOR U35228 ( .A(b[7045]), .B(n21137), .Z(c[7045]) );
XNOR U35229 ( .A(a[7045]), .B(c7045), .Z(n21137) );
XOR U35230 ( .A(c7046), .B(n21138), .Z(c7047) );
ANDN U35231 ( .B(n21139), .A(n21140), .Z(n21138) );
XOR U35232 ( .A(c7046), .B(b[7046]), .Z(n21139) );
XNOR U35233 ( .A(b[7046]), .B(n21140), .Z(c[7046]) );
XNOR U35234 ( .A(a[7046]), .B(c7046), .Z(n21140) );
XOR U35235 ( .A(c7047), .B(n21141), .Z(c7048) );
ANDN U35236 ( .B(n21142), .A(n21143), .Z(n21141) );
XOR U35237 ( .A(c7047), .B(b[7047]), .Z(n21142) );
XNOR U35238 ( .A(b[7047]), .B(n21143), .Z(c[7047]) );
XNOR U35239 ( .A(a[7047]), .B(c7047), .Z(n21143) );
XOR U35240 ( .A(c7048), .B(n21144), .Z(c7049) );
ANDN U35241 ( .B(n21145), .A(n21146), .Z(n21144) );
XOR U35242 ( .A(c7048), .B(b[7048]), .Z(n21145) );
XNOR U35243 ( .A(b[7048]), .B(n21146), .Z(c[7048]) );
XNOR U35244 ( .A(a[7048]), .B(c7048), .Z(n21146) );
XOR U35245 ( .A(c7049), .B(n21147), .Z(c7050) );
ANDN U35246 ( .B(n21148), .A(n21149), .Z(n21147) );
XOR U35247 ( .A(c7049), .B(b[7049]), .Z(n21148) );
XNOR U35248 ( .A(b[7049]), .B(n21149), .Z(c[7049]) );
XNOR U35249 ( .A(a[7049]), .B(c7049), .Z(n21149) );
XOR U35250 ( .A(c7050), .B(n21150), .Z(c7051) );
ANDN U35251 ( .B(n21151), .A(n21152), .Z(n21150) );
XOR U35252 ( .A(c7050), .B(b[7050]), .Z(n21151) );
XNOR U35253 ( .A(b[7050]), .B(n21152), .Z(c[7050]) );
XNOR U35254 ( .A(a[7050]), .B(c7050), .Z(n21152) );
XOR U35255 ( .A(c7051), .B(n21153), .Z(c7052) );
ANDN U35256 ( .B(n21154), .A(n21155), .Z(n21153) );
XOR U35257 ( .A(c7051), .B(b[7051]), .Z(n21154) );
XNOR U35258 ( .A(b[7051]), .B(n21155), .Z(c[7051]) );
XNOR U35259 ( .A(a[7051]), .B(c7051), .Z(n21155) );
XOR U35260 ( .A(c7052), .B(n21156), .Z(c7053) );
ANDN U35261 ( .B(n21157), .A(n21158), .Z(n21156) );
XOR U35262 ( .A(c7052), .B(b[7052]), .Z(n21157) );
XNOR U35263 ( .A(b[7052]), .B(n21158), .Z(c[7052]) );
XNOR U35264 ( .A(a[7052]), .B(c7052), .Z(n21158) );
XOR U35265 ( .A(c7053), .B(n21159), .Z(c7054) );
ANDN U35266 ( .B(n21160), .A(n21161), .Z(n21159) );
XOR U35267 ( .A(c7053), .B(b[7053]), .Z(n21160) );
XNOR U35268 ( .A(b[7053]), .B(n21161), .Z(c[7053]) );
XNOR U35269 ( .A(a[7053]), .B(c7053), .Z(n21161) );
XOR U35270 ( .A(c7054), .B(n21162), .Z(c7055) );
ANDN U35271 ( .B(n21163), .A(n21164), .Z(n21162) );
XOR U35272 ( .A(c7054), .B(b[7054]), .Z(n21163) );
XNOR U35273 ( .A(b[7054]), .B(n21164), .Z(c[7054]) );
XNOR U35274 ( .A(a[7054]), .B(c7054), .Z(n21164) );
XOR U35275 ( .A(c7055), .B(n21165), .Z(c7056) );
ANDN U35276 ( .B(n21166), .A(n21167), .Z(n21165) );
XOR U35277 ( .A(c7055), .B(b[7055]), .Z(n21166) );
XNOR U35278 ( .A(b[7055]), .B(n21167), .Z(c[7055]) );
XNOR U35279 ( .A(a[7055]), .B(c7055), .Z(n21167) );
XOR U35280 ( .A(c7056), .B(n21168), .Z(c7057) );
ANDN U35281 ( .B(n21169), .A(n21170), .Z(n21168) );
XOR U35282 ( .A(c7056), .B(b[7056]), .Z(n21169) );
XNOR U35283 ( .A(b[7056]), .B(n21170), .Z(c[7056]) );
XNOR U35284 ( .A(a[7056]), .B(c7056), .Z(n21170) );
XOR U35285 ( .A(c7057), .B(n21171), .Z(c7058) );
ANDN U35286 ( .B(n21172), .A(n21173), .Z(n21171) );
XOR U35287 ( .A(c7057), .B(b[7057]), .Z(n21172) );
XNOR U35288 ( .A(b[7057]), .B(n21173), .Z(c[7057]) );
XNOR U35289 ( .A(a[7057]), .B(c7057), .Z(n21173) );
XOR U35290 ( .A(c7058), .B(n21174), .Z(c7059) );
ANDN U35291 ( .B(n21175), .A(n21176), .Z(n21174) );
XOR U35292 ( .A(c7058), .B(b[7058]), .Z(n21175) );
XNOR U35293 ( .A(b[7058]), .B(n21176), .Z(c[7058]) );
XNOR U35294 ( .A(a[7058]), .B(c7058), .Z(n21176) );
XOR U35295 ( .A(c7059), .B(n21177), .Z(c7060) );
ANDN U35296 ( .B(n21178), .A(n21179), .Z(n21177) );
XOR U35297 ( .A(c7059), .B(b[7059]), .Z(n21178) );
XNOR U35298 ( .A(b[7059]), .B(n21179), .Z(c[7059]) );
XNOR U35299 ( .A(a[7059]), .B(c7059), .Z(n21179) );
XOR U35300 ( .A(c7060), .B(n21180), .Z(c7061) );
ANDN U35301 ( .B(n21181), .A(n21182), .Z(n21180) );
XOR U35302 ( .A(c7060), .B(b[7060]), .Z(n21181) );
XNOR U35303 ( .A(b[7060]), .B(n21182), .Z(c[7060]) );
XNOR U35304 ( .A(a[7060]), .B(c7060), .Z(n21182) );
XOR U35305 ( .A(c7061), .B(n21183), .Z(c7062) );
ANDN U35306 ( .B(n21184), .A(n21185), .Z(n21183) );
XOR U35307 ( .A(c7061), .B(b[7061]), .Z(n21184) );
XNOR U35308 ( .A(b[7061]), .B(n21185), .Z(c[7061]) );
XNOR U35309 ( .A(a[7061]), .B(c7061), .Z(n21185) );
XOR U35310 ( .A(c7062), .B(n21186), .Z(c7063) );
ANDN U35311 ( .B(n21187), .A(n21188), .Z(n21186) );
XOR U35312 ( .A(c7062), .B(b[7062]), .Z(n21187) );
XNOR U35313 ( .A(b[7062]), .B(n21188), .Z(c[7062]) );
XNOR U35314 ( .A(a[7062]), .B(c7062), .Z(n21188) );
XOR U35315 ( .A(c7063), .B(n21189), .Z(c7064) );
ANDN U35316 ( .B(n21190), .A(n21191), .Z(n21189) );
XOR U35317 ( .A(c7063), .B(b[7063]), .Z(n21190) );
XNOR U35318 ( .A(b[7063]), .B(n21191), .Z(c[7063]) );
XNOR U35319 ( .A(a[7063]), .B(c7063), .Z(n21191) );
XOR U35320 ( .A(c7064), .B(n21192), .Z(c7065) );
ANDN U35321 ( .B(n21193), .A(n21194), .Z(n21192) );
XOR U35322 ( .A(c7064), .B(b[7064]), .Z(n21193) );
XNOR U35323 ( .A(b[7064]), .B(n21194), .Z(c[7064]) );
XNOR U35324 ( .A(a[7064]), .B(c7064), .Z(n21194) );
XOR U35325 ( .A(c7065), .B(n21195), .Z(c7066) );
ANDN U35326 ( .B(n21196), .A(n21197), .Z(n21195) );
XOR U35327 ( .A(c7065), .B(b[7065]), .Z(n21196) );
XNOR U35328 ( .A(b[7065]), .B(n21197), .Z(c[7065]) );
XNOR U35329 ( .A(a[7065]), .B(c7065), .Z(n21197) );
XOR U35330 ( .A(c7066), .B(n21198), .Z(c7067) );
ANDN U35331 ( .B(n21199), .A(n21200), .Z(n21198) );
XOR U35332 ( .A(c7066), .B(b[7066]), .Z(n21199) );
XNOR U35333 ( .A(b[7066]), .B(n21200), .Z(c[7066]) );
XNOR U35334 ( .A(a[7066]), .B(c7066), .Z(n21200) );
XOR U35335 ( .A(c7067), .B(n21201), .Z(c7068) );
ANDN U35336 ( .B(n21202), .A(n21203), .Z(n21201) );
XOR U35337 ( .A(c7067), .B(b[7067]), .Z(n21202) );
XNOR U35338 ( .A(b[7067]), .B(n21203), .Z(c[7067]) );
XNOR U35339 ( .A(a[7067]), .B(c7067), .Z(n21203) );
XOR U35340 ( .A(c7068), .B(n21204), .Z(c7069) );
ANDN U35341 ( .B(n21205), .A(n21206), .Z(n21204) );
XOR U35342 ( .A(c7068), .B(b[7068]), .Z(n21205) );
XNOR U35343 ( .A(b[7068]), .B(n21206), .Z(c[7068]) );
XNOR U35344 ( .A(a[7068]), .B(c7068), .Z(n21206) );
XOR U35345 ( .A(c7069), .B(n21207), .Z(c7070) );
ANDN U35346 ( .B(n21208), .A(n21209), .Z(n21207) );
XOR U35347 ( .A(c7069), .B(b[7069]), .Z(n21208) );
XNOR U35348 ( .A(b[7069]), .B(n21209), .Z(c[7069]) );
XNOR U35349 ( .A(a[7069]), .B(c7069), .Z(n21209) );
XOR U35350 ( .A(c7070), .B(n21210), .Z(c7071) );
ANDN U35351 ( .B(n21211), .A(n21212), .Z(n21210) );
XOR U35352 ( .A(c7070), .B(b[7070]), .Z(n21211) );
XNOR U35353 ( .A(b[7070]), .B(n21212), .Z(c[7070]) );
XNOR U35354 ( .A(a[7070]), .B(c7070), .Z(n21212) );
XOR U35355 ( .A(c7071), .B(n21213), .Z(c7072) );
ANDN U35356 ( .B(n21214), .A(n21215), .Z(n21213) );
XOR U35357 ( .A(c7071), .B(b[7071]), .Z(n21214) );
XNOR U35358 ( .A(b[7071]), .B(n21215), .Z(c[7071]) );
XNOR U35359 ( .A(a[7071]), .B(c7071), .Z(n21215) );
XOR U35360 ( .A(c7072), .B(n21216), .Z(c7073) );
ANDN U35361 ( .B(n21217), .A(n21218), .Z(n21216) );
XOR U35362 ( .A(c7072), .B(b[7072]), .Z(n21217) );
XNOR U35363 ( .A(b[7072]), .B(n21218), .Z(c[7072]) );
XNOR U35364 ( .A(a[7072]), .B(c7072), .Z(n21218) );
XOR U35365 ( .A(c7073), .B(n21219), .Z(c7074) );
ANDN U35366 ( .B(n21220), .A(n21221), .Z(n21219) );
XOR U35367 ( .A(c7073), .B(b[7073]), .Z(n21220) );
XNOR U35368 ( .A(b[7073]), .B(n21221), .Z(c[7073]) );
XNOR U35369 ( .A(a[7073]), .B(c7073), .Z(n21221) );
XOR U35370 ( .A(c7074), .B(n21222), .Z(c7075) );
ANDN U35371 ( .B(n21223), .A(n21224), .Z(n21222) );
XOR U35372 ( .A(c7074), .B(b[7074]), .Z(n21223) );
XNOR U35373 ( .A(b[7074]), .B(n21224), .Z(c[7074]) );
XNOR U35374 ( .A(a[7074]), .B(c7074), .Z(n21224) );
XOR U35375 ( .A(c7075), .B(n21225), .Z(c7076) );
ANDN U35376 ( .B(n21226), .A(n21227), .Z(n21225) );
XOR U35377 ( .A(c7075), .B(b[7075]), .Z(n21226) );
XNOR U35378 ( .A(b[7075]), .B(n21227), .Z(c[7075]) );
XNOR U35379 ( .A(a[7075]), .B(c7075), .Z(n21227) );
XOR U35380 ( .A(c7076), .B(n21228), .Z(c7077) );
ANDN U35381 ( .B(n21229), .A(n21230), .Z(n21228) );
XOR U35382 ( .A(c7076), .B(b[7076]), .Z(n21229) );
XNOR U35383 ( .A(b[7076]), .B(n21230), .Z(c[7076]) );
XNOR U35384 ( .A(a[7076]), .B(c7076), .Z(n21230) );
XOR U35385 ( .A(c7077), .B(n21231), .Z(c7078) );
ANDN U35386 ( .B(n21232), .A(n21233), .Z(n21231) );
XOR U35387 ( .A(c7077), .B(b[7077]), .Z(n21232) );
XNOR U35388 ( .A(b[7077]), .B(n21233), .Z(c[7077]) );
XNOR U35389 ( .A(a[7077]), .B(c7077), .Z(n21233) );
XOR U35390 ( .A(c7078), .B(n21234), .Z(c7079) );
ANDN U35391 ( .B(n21235), .A(n21236), .Z(n21234) );
XOR U35392 ( .A(c7078), .B(b[7078]), .Z(n21235) );
XNOR U35393 ( .A(b[7078]), .B(n21236), .Z(c[7078]) );
XNOR U35394 ( .A(a[7078]), .B(c7078), .Z(n21236) );
XOR U35395 ( .A(c7079), .B(n21237), .Z(c7080) );
ANDN U35396 ( .B(n21238), .A(n21239), .Z(n21237) );
XOR U35397 ( .A(c7079), .B(b[7079]), .Z(n21238) );
XNOR U35398 ( .A(b[7079]), .B(n21239), .Z(c[7079]) );
XNOR U35399 ( .A(a[7079]), .B(c7079), .Z(n21239) );
XOR U35400 ( .A(c7080), .B(n21240), .Z(c7081) );
ANDN U35401 ( .B(n21241), .A(n21242), .Z(n21240) );
XOR U35402 ( .A(c7080), .B(b[7080]), .Z(n21241) );
XNOR U35403 ( .A(b[7080]), .B(n21242), .Z(c[7080]) );
XNOR U35404 ( .A(a[7080]), .B(c7080), .Z(n21242) );
XOR U35405 ( .A(c7081), .B(n21243), .Z(c7082) );
ANDN U35406 ( .B(n21244), .A(n21245), .Z(n21243) );
XOR U35407 ( .A(c7081), .B(b[7081]), .Z(n21244) );
XNOR U35408 ( .A(b[7081]), .B(n21245), .Z(c[7081]) );
XNOR U35409 ( .A(a[7081]), .B(c7081), .Z(n21245) );
XOR U35410 ( .A(c7082), .B(n21246), .Z(c7083) );
ANDN U35411 ( .B(n21247), .A(n21248), .Z(n21246) );
XOR U35412 ( .A(c7082), .B(b[7082]), .Z(n21247) );
XNOR U35413 ( .A(b[7082]), .B(n21248), .Z(c[7082]) );
XNOR U35414 ( .A(a[7082]), .B(c7082), .Z(n21248) );
XOR U35415 ( .A(c7083), .B(n21249), .Z(c7084) );
ANDN U35416 ( .B(n21250), .A(n21251), .Z(n21249) );
XOR U35417 ( .A(c7083), .B(b[7083]), .Z(n21250) );
XNOR U35418 ( .A(b[7083]), .B(n21251), .Z(c[7083]) );
XNOR U35419 ( .A(a[7083]), .B(c7083), .Z(n21251) );
XOR U35420 ( .A(c7084), .B(n21252), .Z(c7085) );
ANDN U35421 ( .B(n21253), .A(n21254), .Z(n21252) );
XOR U35422 ( .A(c7084), .B(b[7084]), .Z(n21253) );
XNOR U35423 ( .A(b[7084]), .B(n21254), .Z(c[7084]) );
XNOR U35424 ( .A(a[7084]), .B(c7084), .Z(n21254) );
XOR U35425 ( .A(c7085), .B(n21255), .Z(c7086) );
ANDN U35426 ( .B(n21256), .A(n21257), .Z(n21255) );
XOR U35427 ( .A(c7085), .B(b[7085]), .Z(n21256) );
XNOR U35428 ( .A(b[7085]), .B(n21257), .Z(c[7085]) );
XNOR U35429 ( .A(a[7085]), .B(c7085), .Z(n21257) );
XOR U35430 ( .A(c7086), .B(n21258), .Z(c7087) );
ANDN U35431 ( .B(n21259), .A(n21260), .Z(n21258) );
XOR U35432 ( .A(c7086), .B(b[7086]), .Z(n21259) );
XNOR U35433 ( .A(b[7086]), .B(n21260), .Z(c[7086]) );
XNOR U35434 ( .A(a[7086]), .B(c7086), .Z(n21260) );
XOR U35435 ( .A(c7087), .B(n21261), .Z(c7088) );
ANDN U35436 ( .B(n21262), .A(n21263), .Z(n21261) );
XOR U35437 ( .A(c7087), .B(b[7087]), .Z(n21262) );
XNOR U35438 ( .A(b[7087]), .B(n21263), .Z(c[7087]) );
XNOR U35439 ( .A(a[7087]), .B(c7087), .Z(n21263) );
XOR U35440 ( .A(c7088), .B(n21264), .Z(c7089) );
ANDN U35441 ( .B(n21265), .A(n21266), .Z(n21264) );
XOR U35442 ( .A(c7088), .B(b[7088]), .Z(n21265) );
XNOR U35443 ( .A(b[7088]), .B(n21266), .Z(c[7088]) );
XNOR U35444 ( .A(a[7088]), .B(c7088), .Z(n21266) );
XOR U35445 ( .A(c7089), .B(n21267), .Z(c7090) );
ANDN U35446 ( .B(n21268), .A(n21269), .Z(n21267) );
XOR U35447 ( .A(c7089), .B(b[7089]), .Z(n21268) );
XNOR U35448 ( .A(b[7089]), .B(n21269), .Z(c[7089]) );
XNOR U35449 ( .A(a[7089]), .B(c7089), .Z(n21269) );
XOR U35450 ( .A(c7090), .B(n21270), .Z(c7091) );
ANDN U35451 ( .B(n21271), .A(n21272), .Z(n21270) );
XOR U35452 ( .A(c7090), .B(b[7090]), .Z(n21271) );
XNOR U35453 ( .A(b[7090]), .B(n21272), .Z(c[7090]) );
XNOR U35454 ( .A(a[7090]), .B(c7090), .Z(n21272) );
XOR U35455 ( .A(c7091), .B(n21273), .Z(c7092) );
ANDN U35456 ( .B(n21274), .A(n21275), .Z(n21273) );
XOR U35457 ( .A(c7091), .B(b[7091]), .Z(n21274) );
XNOR U35458 ( .A(b[7091]), .B(n21275), .Z(c[7091]) );
XNOR U35459 ( .A(a[7091]), .B(c7091), .Z(n21275) );
XOR U35460 ( .A(c7092), .B(n21276), .Z(c7093) );
ANDN U35461 ( .B(n21277), .A(n21278), .Z(n21276) );
XOR U35462 ( .A(c7092), .B(b[7092]), .Z(n21277) );
XNOR U35463 ( .A(b[7092]), .B(n21278), .Z(c[7092]) );
XNOR U35464 ( .A(a[7092]), .B(c7092), .Z(n21278) );
XOR U35465 ( .A(c7093), .B(n21279), .Z(c7094) );
ANDN U35466 ( .B(n21280), .A(n21281), .Z(n21279) );
XOR U35467 ( .A(c7093), .B(b[7093]), .Z(n21280) );
XNOR U35468 ( .A(b[7093]), .B(n21281), .Z(c[7093]) );
XNOR U35469 ( .A(a[7093]), .B(c7093), .Z(n21281) );
XOR U35470 ( .A(c7094), .B(n21282), .Z(c7095) );
ANDN U35471 ( .B(n21283), .A(n21284), .Z(n21282) );
XOR U35472 ( .A(c7094), .B(b[7094]), .Z(n21283) );
XNOR U35473 ( .A(b[7094]), .B(n21284), .Z(c[7094]) );
XNOR U35474 ( .A(a[7094]), .B(c7094), .Z(n21284) );
XOR U35475 ( .A(c7095), .B(n21285), .Z(c7096) );
ANDN U35476 ( .B(n21286), .A(n21287), .Z(n21285) );
XOR U35477 ( .A(c7095), .B(b[7095]), .Z(n21286) );
XNOR U35478 ( .A(b[7095]), .B(n21287), .Z(c[7095]) );
XNOR U35479 ( .A(a[7095]), .B(c7095), .Z(n21287) );
XOR U35480 ( .A(c7096), .B(n21288), .Z(c7097) );
ANDN U35481 ( .B(n21289), .A(n21290), .Z(n21288) );
XOR U35482 ( .A(c7096), .B(b[7096]), .Z(n21289) );
XNOR U35483 ( .A(b[7096]), .B(n21290), .Z(c[7096]) );
XNOR U35484 ( .A(a[7096]), .B(c7096), .Z(n21290) );
XOR U35485 ( .A(c7097), .B(n21291), .Z(c7098) );
ANDN U35486 ( .B(n21292), .A(n21293), .Z(n21291) );
XOR U35487 ( .A(c7097), .B(b[7097]), .Z(n21292) );
XNOR U35488 ( .A(b[7097]), .B(n21293), .Z(c[7097]) );
XNOR U35489 ( .A(a[7097]), .B(c7097), .Z(n21293) );
XOR U35490 ( .A(c7098), .B(n21294), .Z(c7099) );
ANDN U35491 ( .B(n21295), .A(n21296), .Z(n21294) );
XOR U35492 ( .A(c7098), .B(b[7098]), .Z(n21295) );
XNOR U35493 ( .A(b[7098]), .B(n21296), .Z(c[7098]) );
XNOR U35494 ( .A(a[7098]), .B(c7098), .Z(n21296) );
XOR U35495 ( .A(c7099), .B(n21297), .Z(c7100) );
ANDN U35496 ( .B(n21298), .A(n21299), .Z(n21297) );
XOR U35497 ( .A(c7099), .B(b[7099]), .Z(n21298) );
XNOR U35498 ( .A(b[7099]), .B(n21299), .Z(c[7099]) );
XNOR U35499 ( .A(a[7099]), .B(c7099), .Z(n21299) );
XOR U35500 ( .A(c7100), .B(n21300), .Z(c7101) );
ANDN U35501 ( .B(n21301), .A(n21302), .Z(n21300) );
XOR U35502 ( .A(c7100), .B(b[7100]), .Z(n21301) );
XNOR U35503 ( .A(b[7100]), .B(n21302), .Z(c[7100]) );
XNOR U35504 ( .A(a[7100]), .B(c7100), .Z(n21302) );
XOR U35505 ( .A(c7101), .B(n21303), .Z(c7102) );
ANDN U35506 ( .B(n21304), .A(n21305), .Z(n21303) );
XOR U35507 ( .A(c7101), .B(b[7101]), .Z(n21304) );
XNOR U35508 ( .A(b[7101]), .B(n21305), .Z(c[7101]) );
XNOR U35509 ( .A(a[7101]), .B(c7101), .Z(n21305) );
XOR U35510 ( .A(c7102), .B(n21306), .Z(c7103) );
ANDN U35511 ( .B(n21307), .A(n21308), .Z(n21306) );
XOR U35512 ( .A(c7102), .B(b[7102]), .Z(n21307) );
XNOR U35513 ( .A(b[7102]), .B(n21308), .Z(c[7102]) );
XNOR U35514 ( .A(a[7102]), .B(c7102), .Z(n21308) );
XOR U35515 ( .A(c7103), .B(n21309), .Z(c7104) );
ANDN U35516 ( .B(n21310), .A(n21311), .Z(n21309) );
XOR U35517 ( .A(c7103), .B(b[7103]), .Z(n21310) );
XNOR U35518 ( .A(b[7103]), .B(n21311), .Z(c[7103]) );
XNOR U35519 ( .A(a[7103]), .B(c7103), .Z(n21311) );
XOR U35520 ( .A(c7104), .B(n21312), .Z(c7105) );
ANDN U35521 ( .B(n21313), .A(n21314), .Z(n21312) );
XOR U35522 ( .A(c7104), .B(b[7104]), .Z(n21313) );
XNOR U35523 ( .A(b[7104]), .B(n21314), .Z(c[7104]) );
XNOR U35524 ( .A(a[7104]), .B(c7104), .Z(n21314) );
XOR U35525 ( .A(c7105), .B(n21315), .Z(c7106) );
ANDN U35526 ( .B(n21316), .A(n21317), .Z(n21315) );
XOR U35527 ( .A(c7105), .B(b[7105]), .Z(n21316) );
XNOR U35528 ( .A(b[7105]), .B(n21317), .Z(c[7105]) );
XNOR U35529 ( .A(a[7105]), .B(c7105), .Z(n21317) );
XOR U35530 ( .A(c7106), .B(n21318), .Z(c7107) );
ANDN U35531 ( .B(n21319), .A(n21320), .Z(n21318) );
XOR U35532 ( .A(c7106), .B(b[7106]), .Z(n21319) );
XNOR U35533 ( .A(b[7106]), .B(n21320), .Z(c[7106]) );
XNOR U35534 ( .A(a[7106]), .B(c7106), .Z(n21320) );
XOR U35535 ( .A(c7107), .B(n21321), .Z(c7108) );
ANDN U35536 ( .B(n21322), .A(n21323), .Z(n21321) );
XOR U35537 ( .A(c7107), .B(b[7107]), .Z(n21322) );
XNOR U35538 ( .A(b[7107]), .B(n21323), .Z(c[7107]) );
XNOR U35539 ( .A(a[7107]), .B(c7107), .Z(n21323) );
XOR U35540 ( .A(c7108), .B(n21324), .Z(c7109) );
ANDN U35541 ( .B(n21325), .A(n21326), .Z(n21324) );
XOR U35542 ( .A(c7108), .B(b[7108]), .Z(n21325) );
XNOR U35543 ( .A(b[7108]), .B(n21326), .Z(c[7108]) );
XNOR U35544 ( .A(a[7108]), .B(c7108), .Z(n21326) );
XOR U35545 ( .A(c7109), .B(n21327), .Z(c7110) );
ANDN U35546 ( .B(n21328), .A(n21329), .Z(n21327) );
XOR U35547 ( .A(c7109), .B(b[7109]), .Z(n21328) );
XNOR U35548 ( .A(b[7109]), .B(n21329), .Z(c[7109]) );
XNOR U35549 ( .A(a[7109]), .B(c7109), .Z(n21329) );
XOR U35550 ( .A(c7110), .B(n21330), .Z(c7111) );
ANDN U35551 ( .B(n21331), .A(n21332), .Z(n21330) );
XOR U35552 ( .A(c7110), .B(b[7110]), .Z(n21331) );
XNOR U35553 ( .A(b[7110]), .B(n21332), .Z(c[7110]) );
XNOR U35554 ( .A(a[7110]), .B(c7110), .Z(n21332) );
XOR U35555 ( .A(c7111), .B(n21333), .Z(c7112) );
ANDN U35556 ( .B(n21334), .A(n21335), .Z(n21333) );
XOR U35557 ( .A(c7111), .B(b[7111]), .Z(n21334) );
XNOR U35558 ( .A(b[7111]), .B(n21335), .Z(c[7111]) );
XNOR U35559 ( .A(a[7111]), .B(c7111), .Z(n21335) );
XOR U35560 ( .A(c7112), .B(n21336), .Z(c7113) );
ANDN U35561 ( .B(n21337), .A(n21338), .Z(n21336) );
XOR U35562 ( .A(c7112), .B(b[7112]), .Z(n21337) );
XNOR U35563 ( .A(b[7112]), .B(n21338), .Z(c[7112]) );
XNOR U35564 ( .A(a[7112]), .B(c7112), .Z(n21338) );
XOR U35565 ( .A(c7113), .B(n21339), .Z(c7114) );
ANDN U35566 ( .B(n21340), .A(n21341), .Z(n21339) );
XOR U35567 ( .A(c7113), .B(b[7113]), .Z(n21340) );
XNOR U35568 ( .A(b[7113]), .B(n21341), .Z(c[7113]) );
XNOR U35569 ( .A(a[7113]), .B(c7113), .Z(n21341) );
XOR U35570 ( .A(c7114), .B(n21342), .Z(c7115) );
ANDN U35571 ( .B(n21343), .A(n21344), .Z(n21342) );
XOR U35572 ( .A(c7114), .B(b[7114]), .Z(n21343) );
XNOR U35573 ( .A(b[7114]), .B(n21344), .Z(c[7114]) );
XNOR U35574 ( .A(a[7114]), .B(c7114), .Z(n21344) );
XOR U35575 ( .A(c7115), .B(n21345), .Z(c7116) );
ANDN U35576 ( .B(n21346), .A(n21347), .Z(n21345) );
XOR U35577 ( .A(c7115), .B(b[7115]), .Z(n21346) );
XNOR U35578 ( .A(b[7115]), .B(n21347), .Z(c[7115]) );
XNOR U35579 ( .A(a[7115]), .B(c7115), .Z(n21347) );
XOR U35580 ( .A(c7116), .B(n21348), .Z(c7117) );
ANDN U35581 ( .B(n21349), .A(n21350), .Z(n21348) );
XOR U35582 ( .A(c7116), .B(b[7116]), .Z(n21349) );
XNOR U35583 ( .A(b[7116]), .B(n21350), .Z(c[7116]) );
XNOR U35584 ( .A(a[7116]), .B(c7116), .Z(n21350) );
XOR U35585 ( .A(c7117), .B(n21351), .Z(c7118) );
ANDN U35586 ( .B(n21352), .A(n21353), .Z(n21351) );
XOR U35587 ( .A(c7117), .B(b[7117]), .Z(n21352) );
XNOR U35588 ( .A(b[7117]), .B(n21353), .Z(c[7117]) );
XNOR U35589 ( .A(a[7117]), .B(c7117), .Z(n21353) );
XOR U35590 ( .A(c7118), .B(n21354), .Z(c7119) );
ANDN U35591 ( .B(n21355), .A(n21356), .Z(n21354) );
XOR U35592 ( .A(c7118), .B(b[7118]), .Z(n21355) );
XNOR U35593 ( .A(b[7118]), .B(n21356), .Z(c[7118]) );
XNOR U35594 ( .A(a[7118]), .B(c7118), .Z(n21356) );
XOR U35595 ( .A(c7119), .B(n21357), .Z(c7120) );
ANDN U35596 ( .B(n21358), .A(n21359), .Z(n21357) );
XOR U35597 ( .A(c7119), .B(b[7119]), .Z(n21358) );
XNOR U35598 ( .A(b[7119]), .B(n21359), .Z(c[7119]) );
XNOR U35599 ( .A(a[7119]), .B(c7119), .Z(n21359) );
XOR U35600 ( .A(c7120), .B(n21360), .Z(c7121) );
ANDN U35601 ( .B(n21361), .A(n21362), .Z(n21360) );
XOR U35602 ( .A(c7120), .B(b[7120]), .Z(n21361) );
XNOR U35603 ( .A(b[7120]), .B(n21362), .Z(c[7120]) );
XNOR U35604 ( .A(a[7120]), .B(c7120), .Z(n21362) );
XOR U35605 ( .A(c7121), .B(n21363), .Z(c7122) );
ANDN U35606 ( .B(n21364), .A(n21365), .Z(n21363) );
XOR U35607 ( .A(c7121), .B(b[7121]), .Z(n21364) );
XNOR U35608 ( .A(b[7121]), .B(n21365), .Z(c[7121]) );
XNOR U35609 ( .A(a[7121]), .B(c7121), .Z(n21365) );
XOR U35610 ( .A(c7122), .B(n21366), .Z(c7123) );
ANDN U35611 ( .B(n21367), .A(n21368), .Z(n21366) );
XOR U35612 ( .A(c7122), .B(b[7122]), .Z(n21367) );
XNOR U35613 ( .A(b[7122]), .B(n21368), .Z(c[7122]) );
XNOR U35614 ( .A(a[7122]), .B(c7122), .Z(n21368) );
XOR U35615 ( .A(c7123), .B(n21369), .Z(c7124) );
ANDN U35616 ( .B(n21370), .A(n21371), .Z(n21369) );
XOR U35617 ( .A(c7123), .B(b[7123]), .Z(n21370) );
XNOR U35618 ( .A(b[7123]), .B(n21371), .Z(c[7123]) );
XNOR U35619 ( .A(a[7123]), .B(c7123), .Z(n21371) );
XOR U35620 ( .A(c7124), .B(n21372), .Z(c7125) );
ANDN U35621 ( .B(n21373), .A(n21374), .Z(n21372) );
XOR U35622 ( .A(c7124), .B(b[7124]), .Z(n21373) );
XNOR U35623 ( .A(b[7124]), .B(n21374), .Z(c[7124]) );
XNOR U35624 ( .A(a[7124]), .B(c7124), .Z(n21374) );
XOR U35625 ( .A(c7125), .B(n21375), .Z(c7126) );
ANDN U35626 ( .B(n21376), .A(n21377), .Z(n21375) );
XOR U35627 ( .A(c7125), .B(b[7125]), .Z(n21376) );
XNOR U35628 ( .A(b[7125]), .B(n21377), .Z(c[7125]) );
XNOR U35629 ( .A(a[7125]), .B(c7125), .Z(n21377) );
XOR U35630 ( .A(c7126), .B(n21378), .Z(c7127) );
ANDN U35631 ( .B(n21379), .A(n21380), .Z(n21378) );
XOR U35632 ( .A(c7126), .B(b[7126]), .Z(n21379) );
XNOR U35633 ( .A(b[7126]), .B(n21380), .Z(c[7126]) );
XNOR U35634 ( .A(a[7126]), .B(c7126), .Z(n21380) );
XOR U35635 ( .A(c7127), .B(n21381), .Z(c7128) );
ANDN U35636 ( .B(n21382), .A(n21383), .Z(n21381) );
XOR U35637 ( .A(c7127), .B(b[7127]), .Z(n21382) );
XNOR U35638 ( .A(b[7127]), .B(n21383), .Z(c[7127]) );
XNOR U35639 ( .A(a[7127]), .B(c7127), .Z(n21383) );
XOR U35640 ( .A(c7128), .B(n21384), .Z(c7129) );
ANDN U35641 ( .B(n21385), .A(n21386), .Z(n21384) );
XOR U35642 ( .A(c7128), .B(b[7128]), .Z(n21385) );
XNOR U35643 ( .A(b[7128]), .B(n21386), .Z(c[7128]) );
XNOR U35644 ( .A(a[7128]), .B(c7128), .Z(n21386) );
XOR U35645 ( .A(c7129), .B(n21387), .Z(c7130) );
ANDN U35646 ( .B(n21388), .A(n21389), .Z(n21387) );
XOR U35647 ( .A(c7129), .B(b[7129]), .Z(n21388) );
XNOR U35648 ( .A(b[7129]), .B(n21389), .Z(c[7129]) );
XNOR U35649 ( .A(a[7129]), .B(c7129), .Z(n21389) );
XOR U35650 ( .A(c7130), .B(n21390), .Z(c7131) );
ANDN U35651 ( .B(n21391), .A(n21392), .Z(n21390) );
XOR U35652 ( .A(c7130), .B(b[7130]), .Z(n21391) );
XNOR U35653 ( .A(b[7130]), .B(n21392), .Z(c[7130]) );
XNOR U35654 ( .A(a[7130]), .B(c7130), .Z(n21392) );
XOR U35655 ( .A(c7131), .B(n21393), .Z(c7132) );
ANDN U35656 ( .B(n21394), .A(n21395), .Z(n21393) );
XOR U35657 ( .A(c7131), .B(b[7131]), .Z(n21394) );
XNOR U35658 ( .A(b[7131]), .B(n21395), .Z(c[7131]) );
XNOR U35659 ( .A(a[7131]), .B(c7131), .Z(n21395) );
XOR U35660 ( .A(c7132), .B(n21396), .Z(c7133) );
ANDN U35661 ( .B(n21397), .A(n21398), .Z(n21396) );
XOR U35662 ( .A(c7132), .B(b[7132]), .Z(n21397) );
XNOR U35663 ( .A(b[7132]), .B(n21398), .Z(c[7132]) );
XNOR U35664 ( .A(a[7132]), .B(c7132), .Z(n21398) );
XOR U35665 ( .A(c7133), .B(n21399), .Z(c7134) );
ANDN U35666 ( .B(n21400), .A(n21401), .Z(n21399) );
XOR U35667 ( .A(c7133), .B(b[7133]), .Z(n21400) );
XNOR U35668 ( .A(b[7133]), .B(n21401), .Z(c[7133]) );
XNOR U35669 ( .A(a[7133]), .B(c7133), .Z(n21401) );
XOR U35670 ( .A(c7134), .B(n21402), .Z(c7135) );
ANDN U35671 ( .B(n21403), .A(n21404), .Z(n21402) );
XOR U35672 ( .A(c7134), .B(b[7134]), .Z(n21403) );
XNOR U35673 ( .A(b[7134]), .B(n21404), .Z(c[7134]) );
XNOR U35674 ( .A(a[7134]), .B(c7134), .Z(n21404) );
XOR U35675 ( .A(c7135), .B(n21405), .Z(c7136) );
ANDN U35676 ( .B(n21406), .A(n21407), .Z(n21405) );
XOR U35677 ( .A(c7135), .B(b[7135]), .Z(n21406) );
XNOR U35678 ( .A(b[7135]), .B(n21407), .Z(c[7135]) );
XNOR U35679 ( .A(a[7135]), .B(c7135), .Z(n21407) );
XOR U35680 ( .A(c7136), .B(n21408), .Z(c7137) );
ANDN U35681 ( .B(n21409), .A(n21410), .Z(n21408) );
XOR U35682 ( .A(c7136), .B(b[7136]), .Z(n21409) );
XNOR U35683 ( .A(b[7136]), .B(n21410), .Z(c[7136]) );
XNOR U35684 ( .A(a[7136]), .B(c7136), .Z(n21410) );
XOR U35685 ( .A(c7137), .B(n21411), .Z(c7138) );
ANDN U35686 ( .B(n21412), .A(n21413), .Z(n21411) );
XOR U35687 ( .A(c7137), .B(b[7137]), .Z(n21412) );
XNOR U35688 ( .A(b[7137]), .B(n21413), .Z(c[7137]) );
XNOR U35689 ( .A(a[7137]), .B(c7137), .Z(n21413) );
XOR U35690 ( .A(c7138), .B(n21414), .Z(c7139) );
ANDN U35691 ( .B(n21415), .A(n21416), .Z(n21414) );
XOR U35692 ( .A(c7138), .B(b[7138]), .Z(n21415) );
XNOR U35693 ( .A(b[7138]), .B(n21416), .Z(c[7138]) );
XNOR U35694 ( .A(a[7138]), .B(c7138), .Z(n21416) );
XOR U35695 ( .A(c7139), .B(n21417), .Z(c7140) );
ANDN U35696 ( .B(n21418), .A(n21419), .Z(n21417) );
XOR U35697 ( .A(c7139), .B(b[7139]), .Z(n21418) );
XNOR U35698 ( .A(b[7139]), .B(n21419), .Z(c[7139]) );
XNOR U35699 ( .A(a[7139]), .B(c7139), .Z(n21419) );
XOR U35700 ( .A(c7140), .B(n21420), .Z(c7141) );
ANDN U35701 ( .B(n21421), .A(n21422), .Z(n21420) );
XOR U35702 ( .A(c7140), .B(b[7140]), .Z(n21421) );
XNOR U35703 ( .A(b[7140]), .B(n21422), .Z(c[7140]) );
XNOR U35704 ( .A(a[7140]), .B(c7140), .Z(n21422) );
XOR U35705 ( .A(c7141), .B(n21423), .Z(c7142) );
ANDN U35706 ( .B(n21424), .A(n21425), .Z(n21423) );
XOR U35707 ( .A(c7141), .B(b[7141]), .Z(n21424) );
XNOR U35708 ( .A(b[7141]), .B(n21425), .Z(c[7141]) );
XNOR U35709 ( .A(a[7141]), .B(c7141), .Z(n21425) );
XOR U35710 ( .A(c7142), .B(n21426), .Z(c7143) );
ANDN U35711 ( .B(n21427), .A(n21428), .Z(n21426) );
XOR U35712 ( .A(c7142), .B(b[7142]), .Z(n21427) );
XNOR U35713 ( .A(b[7142]), .B(n21428), .Z(c[7142]) );
XNOR U35714 ( .A(a[7142]), .B(c7142), .Z(n21428) );
XOR U35715 ( .A(c7143), .B(n21429), .Z(c7144) );
ANDN U35716 ( .B(n21430), .A(n21431), .Z(n21429) );
XOR U35717 ( .A(c7143), .B(b[7143]), .Z(n21430) );
XNOR U35718 ( .A(b[7143]), .B(n21431), .Z(c[7143]) );
XNOR U35719 ( .A(a[7143]), .B(c7143), .Z(n21431) );
XOR U35720 ( .A(c7144), .B(n21432), .Z(c7145) );
ANDN U35721 ( .B(n21433), .A(n21434), .Z(n21432) );
XOR U35722 ( .A(c7144), .B(b[7144]), .Z(n21433) );
XNOR U35723 ( .A(b[7144]), .B(n21434), .Z(c[7144]) );
XNOR U35724 ( .A(a[7144]), .B(c7144), .Z(n21434) );
XOR U35725 ( .A(c7145), .B(n21435), .Z(c7146) );
ANDN U35726 ( .B(n21436), .A(n21437), .Z(n21435) );
XOR U35727 ( .A(c7145), .B(b[7145]), .Z(n21436) );
XNOR U35728 ( .A(b[7145]), .B(n21437), .Z(c[7145]) );
XNOR U35729 ( .A(a[7145]), .B(c7145), .Z(n21437) );
XOR U35730 ( .A(c7146), .B(n21438), .Z(c7147) );
ANDN U35731 ( .B(n21439), .A(n21440), .Z(n21438) );
XOR U35732 ( .A(c7146), .B(b[7146]), .Z(n21439) );
XNOR U35733 ( .A(b[7146]), .B(n21440), .Z(c[7146]) );
XNOR U35734 ( .A(a[7146]), .B(c7146), .Z(n21440) );
XOR U35735 ( .A(c7147), .B(n21441), .Z(c7148) );
ANDN U35736 ( .B(n21442), .A(n21443), .Z(n21441) );
XOR U35737 ( .A(c7147), .B(b[7147]), .Z(n21442) );
XNOR U35738 ( .A(b[7147]), .B(n21443), .Z(c[7147]) );
XNOR U35739 ( .A(a[7147]), .B(c7147), .Z(n21443) );
XOR U35740 ( .A(c7148), .B(n21444), .Z(c7149) );
ANDN U35741 ( .B(n21445), .A(n21446), .Z(n21444) );
XOR U35742 ( .A(c7148), .B(b[7148]), .Z(n21445) );
XNOR U35743 ( .A(b[7148]), .B(n21446), .Z(c[7148]) );
XNOR U35744 ( .A(a[7148]), .B(c7148), .Z(n21446) );
XOR U35745 ( .A(c7149), .B(n21447), .Z(c7150) );
ANDN U35746 ( .B(n21448), .A(n21449), .Z(n21447) );
XOR U35747 ( .A(c7149), .B(b[7149]), .Z(n21448) );
XNOR U35748 ( .A(b[7149]), .B(n21449), .Z(c[7149]) );
XNOR U35749 ( .A(a[7149]), .B(c7149), .Z(n21449) );
XOR U35750 ( .A(c7150), .B(n21450), .Z(c7151) );
ANDN U35751 ( .B(n21451), .A(n21452), .Z(n21450) );
XOR U35752 ( .A(c7150), .B(b[7150]), .Z(n21451) );
XNOR U35753 ( .A(b[7150]), .B(n21452), .Z(c[7150]) );
XNOR U35754 ( .A(a[7150]), .B(c7150), .Z(n21452) );
XOR U35755 ( .A(c7151), .B(n21453), .Z(c7152) );
ANDN U35756 ( .B(n21454), .A(n21455), .Z(n21453) );
XOR U35757 ( .A(c7151), .B(b[7151]), .Z(n21454) );
XNOR U35758 ( .A(b[7151]), .B(n21455), .Z(c[7151]) );
XNOR U35759 ( .A(a[7151]), .B(c7151), .Z(n21455) );
XOR U35760 ( .A(c7152), .B(n21456), .Z(c7153) );
ANDN U35761 ( .B(n21457), .A(n21458), .Z(n21456) );
XOR U35762 ( .A(c7152), .B(b[7152]), .Z(n21457) );
XNOR U35763 ( .A(b[7152]), .B(n21458), .Z(c[7152]) );
XNOR U35764 ( .A(a[7152]), .B(c7152), .Z(n21458) );
XOR U35765 ( .A(c7153), .B(n21459), .Z(c7154) );
ANDN U35766 ( .B(n21460), .A(n21461), .Z(n21459) );
XOR U35767 ( .A(c7153), .B(b[7153]), .Z(n21460) );
XNOR U35768 ( .A(b[7153]), .B(n21461), .Z(c[7153]) );
XNOR U35769 ( .A(a[7153]), .B(c7153), .Z(n21461) );
XOR U35770 ( .A(c7154), .B(n21462), .Z(c7155) );
ANDN U35771 ( .B(n21463), .A(n21464), .Z(n21462) );
XOR U35772 ( .A(c7154), .B(b[7154]), .Z(n21463) );
XNOR U35773 ( .A(b[7154]), .B(n21464), .Z(c[7154]) );
XNOR U35774 ( .A(a[7154]), .B(c7154), .Z(n21464) );
XOR U35775 ( .A(c7155), .B(n21465), .Z(c7156) );
ANDN U35776 ( .B(n21466), .A(n21467), .Z(n21465) );
XOR U35777 ( .A(c7155), .B(b[7155]), .Z(n21466) );
XNOR U35778 ( .A(b[7155]), .B(n21467), .Z(c[7155]) );
XNOR U35779 ( .A(a[7155]), .B(c7155), .Z(n21467) );
XOR U35780 ( .A(c7156), .B(n21468), .Z(c7157) );
ANDN U35781 ( .B(n21469), .A(n21470), .Z(n21468) );
XOR U35782 ( .A(c7156), .B(b[7156]), .Z(n21469) );
XNOR U35783 ( .A(b[7156]), .B(n21470), .Z(c[7156]) );
XNOR U35784 ( .A(a[7156]), .B(c7156), .Z(n21470) );
XOR U35785 ( .A(c7157), .B(n21471), .Z(c7158) );
ANDN U35786 ( .B(n21472), .A(n21473), .Z(n21471) );
XOR U35787 ( .A(c7157), .B(b[7157]), .Z(n21472) );
XNOR U35788 ( .A(b[7157]), .B(n21473), .Z(c[7157]) );
XNOR U35789 ( .A(a[7157]), .B(c7157), .Z(n21473) );
XOR U35790 ( .A(c7158), .B(n21474), .Z(c7159) );
ANDN U35791 ( .B(n21475), .A(n21476), .Z(n21474) );
XOR U35792 ( .A(c7158), .B(b[7158]), .Z(n21475) );
XNOR U35793 ( .A(b[7158]), .B(n21476), .Z(c[7158]) );
XNOR U35794 ( .A(a[7158]), .B(c7158), .Z(n21476) );
XOR U35795 ( .A(c7159), .B(n21477), .Z(c7160) );
ANDN U35796 ( .B(n21478), .A(n21479), .Z(n21477) );
XOR U35797 ( .A(c7159), .B(b[7159]), .Z(n21478) );
XNOR U35798 ( .A(b[7159]), .B(n21479), .Z(c[7159]) );
XNOR U35799 ( .A(a[7159]), .B(c7159), .Z(n21479) );
XOR U35800 ( .A(c7160), .B(n21480), .Z(c7161) );
ANDN U35801 ( .B(n21481), .A(n21482), .Z(n21480) );
XOR U35802 ( .A(c7160), .B(b[7160]), .Z(n21481) );
XNOR U35803 ( .A(b[7160]), .B(n21482), .Z(c[7160]) );
XNOR U35804 ( .A(a[7160]), .B(c7160), .Z(n21482) );
XOR U35805 ( .A(c7161), .B(n21483), .Z(c7162) );
ANDN U35806 ( .B(n21484), .A(n21485), .Z(n21483) );
XOR U35807 ( .A(c7161), .B(b[7161]), .Z(n21484) );
XNOR U35808 ( .A(b[7161]), .B(n21485), .Z(c[7161]) );
XNOR U35809 ( .A(a[7161]), .B(c7161), .Z(n21485) );
XOR U35810 ( .A(c7162), .B(n21486), .Z(c7163) );
ANDN U35811 ( .B(n21487), .A(n21488), .Z(n21486) );
XOR U35812 ( .A(c7162), .B(b[7162]), .Z(n21487) );
XNOR U35813 ( .A(b[7162]), .B(n21488), .Z(c[7162]) );
XNOR U35814 ( .A(a[7162]), .B(c7162), .Z(n21488) );
XOR U35815 ( .A(c7163), .B(n21489), .Z(c7164) );
ANDN U35816 ( .B(n21490), .A(n21491), .Z(n21489) );
XOR U35817 ( .A(c7163), .B(b[7163]), .Z(n21490) );
XNOR U35818 ( .A(b[7163]), .B(n21491), .Z(c[7163]) );
XNOR U35819 ( .A(a[7163]), .B(c7163), .Z(n21491) );
XOR U35820 ( .A(c7164), .B(n21492), .Z(c7165) );
ANDN U35821 ( .B(n21493), .A(n21494), .Z(n21492) );
XOR U35822 ( .A(c7164), .B(b[7164]), .Z(n21493) );
XNOR U35823 ( .A(b[7164]), .B(n21494), .Z(c[7164]) );
XNOR U35824 ( .A(a[7164]), .B(c7164), .Z(n21494) );
XOR U35825 ( .A(c7165), .B(n21495), .Z(c7166) );
ANDN U35826 ( .B(n21496), .A(n21497), .Z(n21495) );
XOR U35827 ( .A(c7165), .B(b[7165]), .Z(n21496) );
XNOR U35828 ( .A(b[7165]), .B(n21497), .Z(c[7165]) );
XNOR U35829 ( .A(a[7165]), .B(c7165), .Z(n21497) );
XOR U35830 ( .A(c7166), .B(n21498), .Z(c7167) );
ANDN U35831 ( .B(n21499), .A(n21500), .Z(n21498) );
XOR U35832 ( .A(c7166), .B(b[7166]), .Z(n21499) );
XNOR U35833 ( .A(b[7166]), .B(n21500), .Z(c[7166]) );
XNOR U35834 ( .A(a[7166]), .B(c7166), .Z(n21500) );
XOR U35835 ( .A(c7167), .B(n21501), .Z(c7168) );
ANDN U35836 ( .B(n21502), .A(n21503), .Z(n21501) );
XOR U35837 ( .A(c7167), .B(b[7167]), .Z(n21502) );
XNOR U35838 ( .A(b[7167]), .B(n21503), .Z(c[7167]) );
XNOR U35839 ( .A(a[7167]), .B(c7167), .Z(n21503) );
XOR U35840 ( .A(c7168), .B(n21504), .Z(c7169) );
ANDN U35841 ( .B(n21505), .A(n21506), .Z(n21504) );
XOR U35842 ( .A(c7168), .B(b[7168]), .Z(n21505) );
XNOR U35843 ( .A(b[7168]), .B(n21506), .Z(c[7168]) );
XNOR U35844 ( .A(a[7168]), .B(c7168), .Z(n21506) );
XOR U35845 ( .A(c7169), .B(n21507), .Z(c7170) );
ANDN U35846 ( .B(n21508), .A(n21509), .Z(n21507) );
XOR U35847 ( .A(c7169), .B(b[7169]), .Z(n21508) );
XNOR U35848 ( .A(b[7169]), .B(n21509), .Z(c[7169]) );
XNOR U35849 ( .A(a[7169]), .B(c7169), .Z(n21509) );
XOR U35850 ( .A(c7170), .B(n21510), .Z(c7171) );
ANDN U35851 ( .B(n21511), .A(n21512), .Z(n21510) );
XOR U35852 ( .A(c7170), .B(b[7170]), .Z(n21511) );
XNOR U35853 ( .A(b[7170]), .B(n21512), .Z(c[7170]) );
XNOR U35854 ( .A(a[7170]), .B(c7170), .Z(n21512) );
XOR U35855 ( .A(c7171), .B(n21513), .Z(c7172) );
ANDN U35856 ( .B(n21514), .A(n21515), .Z(n21513) );
XOR U35857 ( .A(c7171), .B(b[7171]), .Z(n21514) );
XNOR U35858 ( .A(b[7171]), .B(n21515), .Z(c[7171]) );
XNOR U35859 ( .A(a[7171]), .B(c7171), .Z(n21515) );
XOR U35860 ( .A(c7172), .B(n21516), .Z(c7173) );
ANDN U35861 ( .B(n21517), .A(n21518), .Z(n21516) );
XOR U35862 ( .A(c7172), .B(b[7172]), .Z(n21517) );
XNOR U35863 ( .A(b[7172]), .B(n21518), .Z(c[7172]) );
XNOR U35864 ( .A(a[7172]), .B(c7172), .Z(n21518) );
XOR U35865 ( .A(c7173), .B(n21519), .Z(c7174) );
ANDN U35866 ( .B(n21520), .A(n21521), .Z(n21519) );
XOR U35867 ( .A(c7173), .B(b[7173]), .Z(n21520) );
XNOR U35868 ( .A(b[7173]), .B(n21521), .Z(c[7173]) );
XNOR U35869 ( .A(a[7173]), .B(c7173), .Z(n21521) );
XOR U35870 ( .A(c7174), .B(n21522), .Z(c7175) );
ANDN U35871 ( .B(n21523), .A(n21524), .Z(n21522) );
XOR U35872 ( .A(c7174), .B(b[7174]), .Z(n21523) );
XNOR U35873 ( .A(b[7174]), .B(n21524), .Z(c[7174]) );
XNOR U35874 ( .A(a[7174]), .B(c7174), .Z(n21524) );
XOR U35875 ( .A(c7175), .B(n21525), .Z(c7176) );
ANDN U35876 ( .B(n21526), .A(n21527), .Z(n21525) );
XOR U35877 ( .A(c7175), .B(b[7175]), .Z(n21526) );
XNOR U35878 ( .A(b[7175]), .B(n21527), .Z(c[7175]) );
XNOR U35879 ( .A(a[7175]), .B(c7175), .Z(n21527) );
XOR U35880 ( .A(c7176), .B(n21528), .Z(c7177) );
ANDN U35881 ( .B(n21529), .A(n21530), .Z(n21528) );
XOR U35882 ( .A(c7176), .B(b[7176]), .Z(n21529) );
XNOR U35883 ( .A(b[7176]), .B(n21530), .Z(c[7176]) );
XNOR U35884 ( .A(a[7176]), .B(c7176), .Z(n21530) );
XOR U35885 ( .A(c7177), .B(n21531), .Z(c7178) );
ANDN U35886 ( .B(n21532), .A(n21533), .Z(n21531) );
XOR U35887 ( .A(c7177), .B(b[7177]), .Z(n21532) );
XNOR U35888 ( .A(b[7177]), .B(n21533), .Z(c[7177]) );
XNOR U35889 ( .A(a[7177]), .B(c7177), .Z(n21533) );
XOR U35890 ( .A(c7178), .B(n21534), .Z(c7179) );
ANDN U35891 ( .B(n21535), .A(n21536), .Z(n21534) );
XOR U35892 ( .A(c7178), .B(b[7178]), .Z(n21535) );
XNOR U35893 ( .A(b[7178]), .B(n21536), .Z(c[7178]) );
XNOR U35894 ( .A(a[7178]), .B(c7178), .Z(n21536) );
XOR U35895 ( .A(c7179), .B(n21537), .Z(c7180) );
ANDN U35896 ( .B(n21538), .A(n21539), .Z(n21537) );
XOR U35897 ( .A(c7179), .B(b[7179]), .Z(n21538) );
XNOR U35898 ( .A(b[7179]), .B(n21539), .Z(c[7179]) );
XNOR U35899 ( .A(a[7179]), .B(c7179), .Z(n21539) );
XOR U35900 ( .A(c7180), .B(n21540), .Z(c7181) );
ANDN U35901 ( .B(n21541), .A(n21542), .Z(n21540) );
XOR U35902 ( .A(c7180), .B(b[7180]), .Z(n21541) );
XNOR U35903 ( .A(b[7180]), .B(n21542), .Z(c[7180]) );
XNOR U35904 ( .A(a[7180]), .B(c7180), .Z(n21542) );
XOR U35905 ( .A(c7181), .B(n21543), .Z(c7182) );
ANDN U35906 ( .B(n21544), .A(n21545), .Z(n21543) );
XOR U35907 ( .A(c7181), .B(b[7181]), .Z(n21544) );
XNOR U35908 ( .A(b[7181]), .B(n21545), .Z(c[7181]) );
XNOR U35909 ( .A(a[7181]), .B(c7181), .Z(n21545) );
XOR U35910 ( .A(c7182), .B(n21546), .Z(c7183) );
ANDN U35911 ( .B(n21547), .A(n21548), .Z(n21546) );
XOR U35912 ( .A(c7182), .B(b[7182]), .Z(n21547) );
XNOR U35913 ( .A(b[7182]), .B(n21548), .Z(c[7182]) );
XNOR U35914 ( .A(a[7182]), .B(c7182), .Z(n21548) );
XOR U35915 ( .A(c7183), .B(n21549), .Z(c7184) );
ANDN U35916 ( .B(n21550), .A(n21551), .Z(n21549) );
XOR U35917 ( .A(c7183), .B(b[7183]), .Z(n21550) );
XNOR U35918 ( .A(b[7183]), .B(n21551), .Z(c[7183]) );
XNOR U35919 ( .A(a[7183]), .B(c7183), .Z(n21551) );
XOR U35920 ( .A(c7184), .B(n21552), .Z(c7185) );
ANDN U35921 ( .B(n21553), .A(n21554), .Z(n21552) );
XOR U35922 ( .A(c7184), .B(b[7184]), .Z(n21553) );
XNOR U35923 ( .A(b[7184]), .B(n21554), .Z(c[7184]) );
XNOR U35924 ( .A(a[7184]), .B(c7184), .Z(n21554) );
XOR U35925 ( .A(c7185), .B(n21555), .Z(c7186) );
ANDN U35926 ( .B(n21556), .A(n21557), .Z(n21555) );
XOR U35927 ( .A(c7185), .B(b[7185]), .Z(n21556) );
XNOR U35928 ( .A(b[7185]), .B(n21557), .Z(c[7185]) );
XNOR U35929 ( .A(a[7185]), .B(c7185), .Z(n21557) );
XOR U35930 ( .A(c7186), .B(n21558), .Z(c7187) );
ANDN U35931 ( .B(n21559), .A(n21560), .Z(n21558) );
XOR U35932 ( .A(c7186), .B(b[7186]), .Z(n21559) );
XNOR U35933 ( .A(b[7186]), .B(n21560), .Z(c[7186]) );
XNOR U35934 ( .A(a[7186]), .B(c7186), .Z(n21560) );
XOR U35935 ( .A(c7187), .B(n21561), .Z(c7188) );
ANDN U35936 ( .B(n21562), .A(n21563), .Z(n21561) );
XOR U35937 ( .A(c7187), .B(b[7187]), .Z(n21562) );
XNOR U35938 ( .A(b[7187]), .B(n21563), .Z(c[7187]) );
XNOR U35939 ( .A(a[7187]), .B(c7187), .Z(n21563) );
XOR U35940 ( .A(c7188), .B(n21564), .Z(c7189) );
ANDN U35941 ( .B(n21565), .A(n21566), .Z(n21564) );
XOR U35942 ( .A(c7188), .B(b[7188]), .Z(n21565) );
XNOR U35943 ( .A(b[7188]), .B(n21566), .Z(c[7188]) );
XNOR U35944 ( .A(a[7188]), .B(c7188), .Z(n21566) );
XOR U35945 ( .A(c7189), .B(n21567), .Z(c7190) );
ANDN U35946 ( .B(n21568), .A(n21569), .Z(n21567) );
XOR U35947 ( .A(c7189), .B(b[7189]), .Z(n21568) );
XNOR U35948 ( .A(b[7189]), .B(n21569), .Z(c[7189]) );
XNOR U35949 ( .A(a[7189]), .B(c7189), .Z(n21569) );
XOR U35950 ( .A(c7190), .B(n21570), .Z(c7191) );
ANDN U35951 ( .B(n21571), .A(n21572), .Z(n21570) );
XOR U35952 ( .A(c7190), .B(b[7190]), .Z(n21571) );
XNOR U35953 ( .A(b[7190]), .B(n21572), .Z(c[7190]) );
XNOR U35954 ( .A(a[7190]), .B(c7190), .Z(n21572) );
XOR U35955 ( .A(c7191), .B(n21573), .Z(c7192) );
ANDN U35956 ( .B(n21574), .A(n21575), .Z(n21573) );
XOR U35957 ( .A(c7191), .B(b[7191]), .Z(n21574) );
XNOR U35958 ( .A(b[7191]), .B(n21575), .Z(c[7191]) );
XNOR U35959 ( .A(a[7191]), .B(c7191), .Z(n21575) );
XOR U35960 ( .A(c7192), .B(n21576), .Z(c7193) );
ANDN U35961 ( .B(n21577), .A(n21578), .Z(n21576) );
XOR U35962 ( .A(c7192), .B(b[7192]), .Z(n21577) );
XNOR U35963 ( .A(b[7192]), .B(n21578), .Z(c[7192]) );
XNOR U35964 ( .A(a[7192]), .B(c7192), .Z(n21578) );
XOR U35965 ( .A(c7193), .B(n21579), .Z(c7194) );
ANDN U35966 ( .B(n21580), .A(n21581), .Z(n21579) );
XOR U35967 ( .A(c7193), .B(b[7193]), .Z(n21580) );
XNOR U35968 ( .A(b[7193]), .B(n21581), .Z(c[7193]) );
XNOR U35969 ( .A(a[7193]), .B(c7193), .Z(n21581) );
XOR U35970 ( .A(c7194), .B(n21582), .Z(c7195) );
ANDN U35971 ( .B(n21583), .A(n21584), .Z(n21582) );
XOR U35972 ( .A(c7194), .B(b[7194]), .Z(n21583) );
XNOR U35973 ( .A(b[7194]), .B(n21584), .Z(c[7194]) );
XNOR U35974 ( .A(a[7194]), .B(c7194), .Z(n21584) );
XOR U35975 ( .A(c7195), .B(n21585), .Z(c7196) );
ANDN U35976 ( .B(n21586), .A(n21587), .Z(n21585) );
XOR U35977 ( .A(c7195), .B(b[7195]), .Z(n21586) );
XNOR U35978 ( .A(b[7195]), .B(n21587), .Z(c[7195]) );
XNOR U35979 ( .A(a[7195]), .B(c7195), .Z(n21587) );
XOR U35980 ( .A(c7196), .B(n21588), .Z(c7197) );
ANDN U35981 ( .B(n21589), .A(n21590), .Z(n21588) );
XOR U35982 ( .A(c7196), .B(b[7196]), .Z(n21589) );
XNOR U35983 ( .A(b[7196]), .B(n21590), .Z(c[7196]) );
XNOR U35984 ( .A(a[7196]), .B(c7196), .Z(n21590) );
XOR U35985 ( .A(c7197), .B(n21591), .Z(c7198) );
ANDN U35986 ( .B(n21592), .A(n21593), .Z(n21591) );
XOR U35987 ( .A(c7197), .B(b[7197]), .Z(n21592) );
XNOR U35988 ( .A(b[7197]), .B(n21593), .Z(c[7197]) );
XNOR U35989 ( .A(a[7197]), .B(c7197), .Z(n21593) );
XOR U35990 ( .A(c7198), .B(n21594), .Z(c7199) );
ANDN U35991 ( .B(n21595), .A(n21596), .Z(n21594) );
XOR U35992 ( .A(c7198), .B(b[7198]), .Z(n21595) );
XNOR U35993 ( .A(b[7198]), .B(n21596), .Z(c[7198]) );
XNOR U35994 ( .A(a[7198]), .B(c7198), .Z(n21596) );
XOR U35995 ( .A(c7199), .B(n21597), .Z(c7200) );
ANDN U35996 ( .B(n21598), .A(n21599), .Z(n21597) );
XOR U35997 ( .A(c7199), .B(b[7199]), .Z(n21598) );
XNOR U35998 ( .A(b[7199]), .B(n21599), .Z(c[7199]) );
XNOR U35999 ( .A(a[7199]), .B(c7199), .Z(n21599) );
XOR U36000 ( .A(c7200), .B(n21600), .Z(c7201) );
ANDN U36001 ( .B(n21601), .A(n21602), .Z(n21600) );
XOR U36002 ( .A(c7200), .B(b[7200]), .Z(n21601) );
XNOR U36003 ( .A(b[7200]), .B(n21602), .Z(c[7200]) );
XNOR U36004 ( .A(a[7200]), .B(c7200), .Z(n21602) );
XOR U36005 ( .A(c7201), .B(n21603), .Z(c7202) );
ANDN U36006 ( .B(n21604), .A(n21605), .Z(n21603) );
XOR U36007 ( .A(c7201), .B(b[7201]), .Z(n21604) );
XNOR U36008 ( .A(b[7201]), .B(n21605), .Z(c[7201]) );
XNOR U36009 ( .A(a[7201]), .B(c7201), .Z(n21605) );
XOR U36010 ( .A(c7202), .B(n21606), .Z(c7203) );
ANDN U36011 ( .B(n21607), .A(n21608), .Z(n21606) );
XOR U36012 ( .A(c7202), .B(b[7202]), .Z(n21607) );
XNOR U36013 ( .A(b[7202]), .B(n21608), .Z(c[7202]) );
XNOR U36014 ( .A(a[7202]), .B(c7202), .Z(n21608) );
XOR U36015 ( .A(c7203), .B(n21609), .Z(c7204) );
ANDN U36016 ( .B(n21610), .A(n21611), .Z(n21609) );
XOR U36017 ( .A(c7203), .B(b[7203]), .Z(n21610) );
XNOR U36018 ( .A(b[7203]), .B(n21611), .Z(c[7203]) );
XNOR U36019 ( .A(a[7203]), .B(c7203), .Z(n21611) );
XOR U36020 ( .A(c7204), .B(n21612), .Z(c7205) );
ANDN U36021 ( .B(n21613), .A(n21614), .Z(n21612) );
XOR U36022 ( .A(c7204), .B(b[7204]), .Z(n21613) );
XNOR U36023 ( .A(b[7204]), .B(n21614), .Z(c[7204]) );
XNOR U36024 ( .A(a[7204]), .B(c7204), .Z(n21614) );
XOR U36025 ( .A(c7205), .B(n21615), .Z(c7206) );
ANDN U36026 ( .B(n21616), .A(n21617), .Z(n21615) );
XOR U36027 ( .A(c7205), .B(b[7205]), .Z(n21616) );
XNOR U36028 ( .A(b[7205]), .B(n21617), .Z(c[7205]) );
XNOR U36029 ( .A(a[7205]), .B(c7205), .Z(n21617) );
XOR U36030 ( .A(c7206), .B(n21618), .Z(c7207) );
ANDN U36031 ( .B(n21619), .A(n21620), .Z(n21618) );
XOR U36032 ( .A(c7206), .B(b[7206]), .Z(n21619) );
XNOR U36033 ( .A(b[7206]), .B(n21620), .Z(c[7206]) );
XNOR U36034 ( .A(a[7206]), .B(c7206), .Z(n21620) );
XOR U36035 ( .A(c7207), .B(n21621), .Z(c7208) );
ANDN U36036 ( .B(n21622), .A(n21623), .Z(n21621) );
XOR U36037 ( .A(c7207), .B(b[7207]), .Z(n21622) );
XNOR U36038 ( .A(b[7207]), .B(n21623), .Z(c[7207]) );
XNOR U36039 ( .A(a[7207]), .B(c7207), .Z(n21623) );
XOR U36040 ( .A(c7208), .B(n21624), .Z(c7209) );
ANDN U36041 ( .B(n21625), .A(n21626), .Z(n21624) );
XOR U36042 ( .A(c7208), .B(b[7208]), .Z(n21625) );
XNOR U36043 ( .A(b[7208]), .B(n21626), .Z(c[7208]) );
XNOR U36044 ( .A(a[7208]), .B(c7208), .Z(n21626) );
XOR U36045 ( .A(c7209), .B(n21627), .Z(c7210) );
ANDN U36046 ( .B(n21628), .A(n21629), .Z(n21627) );
XOR U36047 ( .A(c7209), .B(b[7209]), .Z(n21628) );
XNOR U36048 ( .A(b[7209]), .B(n21629), .Z(c[7209]) );
XNOR U36049 ( .A(a[7209]), .B(c7209), .Z(n21629) );
XOR U36050 ( .A(c7210), .B(n21630), .Z(c7211) );
ANDN U36051 ( .B(n21631), .A(n21632), .Z(n21630) );
XOR U36052 ( .A(c7210), .B(b[7210]), .Z(n21631) );
XNOR U36053 ( .A(b[7210]), .B(n21632), .Z(c[7210]) );
XNOR U36054 ( .A(a[7210]), .B(c7210), .Z(n21632) );
XOR U36055 ( .A(c7211), .B(n21633), .Z(c7212) );
ANDN U36056 ( .B(n21634), .A(n21635), .Z(n21633) );
XOR U36057 ( .A(c7211), .B(b[7211]), .Z(n21634) );
XNOR U36058 ( .A(b[7211]), .B(n21635), .Z(c[7211]) );
XNOR U36059 ( .A(a[7211]), .B(c7211), .Z(n21635) );
XOR U36060 ( .A(c7212), .B(n21636), .Z(c7213) );
ANDN U36061 ( .B(n21637), .A(n21638), .Z(n21636) );
XOR U36062 ( .A(c7212), .B(b[7212]), .Z(n21637) );
XNOR U36063 ( .A(b[7212]), .B(n21638), .Z(c[7212]) );
XNOR U36064 ( .A(a[7212]), .B(c7212), .Z(n21638) );
XOR U36065 ( .A(c7213), .B(n21639), .Z(c7214) );
ANDN U36066 ( .B(n21640), .A(n21641), .Z(n21639) );
XOR U36067 ( .A(c7213), .B(b[7213]), .Z(n21640) );
XNOR U36068 ( .A(b[7213]), .B(n21641), .Z(c[7213]) );
XNOR U36069 ( .A(a[7213]), .B(c7213), .Z(n21641) );
XOR U36070 ( .A(c7214), .B(n21642), .Z(c7215) );
ANDN U36071 ( .B(n21643), .A(n21644), .Z(n21642) );
XOR U36072 ( .A(c7214), .B(b[7214]), .Z(n21643) );
XNOR U36073 ( .A(b[7214]), .B(n21644), .Z(c[7214]) );
XNOR U36074 ( .A(a[7214]), .B(c7214), .Z(n21644) );
XOR U36075 ( .A(c7215), .B(n21645), .Z(c7216) );
ANDN U36076 ( .B(n21646), .A(n21647), .Z(n21645) );
XOR U36077 ( .A(c7215), .B(b[7215]), .Z(n21646) );
XNOR U36078 ( .A(b[7215]), .B(n21647), .Z(c[7215]) );
XNOR U36079 ( .A(a[7215]), .B(c7215), .Z(n21647) );
XOR U36080 ( .A(c7216), .B(n21648), .Z(c7217) );
ANDN U36081 ( .B(n21649), .A(n21650), .Z(n21648) );
XOR U36082 ( .A(c7216), .B(b[7216]), .Z(n21649) );
XNOR U36083 ( .A(b[7216]), .B(n21650), .Z(c[7216]) );
XNOR U36084 ( .A(a[7216]), .B(c7216), .Z(n21650) );
XOR U36085 ( .A(c7217), .B(n21651), .Z(c7218) );
ANDN U36086 ( .B(n21652), .A(n21653), .Z(n21651) );
XOR U36087 ( .A(c7217), .B(b[7217]), .Z(n21652) );
XNOR U36088 ( .A(b[7217]), .B(n21653), .Z(c[7217]) );
XNOR U36089 ( .A(a[7217]), .B(c7217), .Z(n21653) );
XOR U36090 ( .A(c7218), .B(n21654), .Z(c7219) );
ANDN U36091 ( .B(n21655), .A(n21656), .Z(n21654) );
XOR U36092 ( .A(c7218), .B(b[7218]), .Z(n21655) );
XNOR U36093 ( .A(b[7218]), .B(n21656), .Z(c[7218]) );
XNOR U36094 ( .A(a[7218]), .B(c7218), .Z(n21656) );
XOR U36095 ( .A(c7219), .B(n21657), .Z(c7220) );
ANDN U36096 ( .B(n21658), .A(n21659), .Z(n21657) );
XOR U36097 ( .A(c7219), .B(b[7219]), .Z(n21658) );
XNOR U36098 ( .A(b[7219]), .B(n21659), .Z(c[7219]) );
XNOR U36099 ( .A(a[7219]), .B(c7219), .Z(n21659) );
XOR U36100 ( .A(c7220), .B(n21660), .Z(c7221) );
ANDN U36101 ( .B(n21661), .A(n21662), .Z(n21660) );
XOR U36102 ( .A(c7220), .B(b[7220]), .Z(n21661) );
XNOR U36103 ( .A(b[7220]), .B(n21662), .Z(c[7220]) );
XNOR U36104 ( .A(a[7220]), .B(c7220), .Z(n21662) );
XOR U36105 ( .A(c7221), .B(n21663), .Z(c7222) );
ANDN U36106 ( .B(n21664), .A(n21665), .Z(n21663) );
XOR U36107 ( .A(c7221), .B(b[7221]), .Z(n21664) );
XNOR U36108 ( .A(b[7221]), .B(n21665), .Z(c[7221]) );
XNOR U36109 ( .A(a[7221]), .B(c7221), .Z(n21665) );
XOR U36110 ( .A(c7222), .B(n21666), .Z(c7223) );
ANDN U36111 ( .B(n21667), .A(n21668), .Z(n21666) );
XOR U36112 ( .A(c7222), .B(b[7222]), .Z(n21667) );
XNOR U36113 ( .A(b[7222]), .B(n21668), .Z(c[7222]) );
XNOR U36114 ( .A(a[7222]), .B(c7222), .Z(n21668) );
XOR U36115 ( .A(c7223), .B(n21669), .Z(c7224) );
ANDN U36116 ( .B(n21670), .A(n21671), .Z(n21669) );
XOR U36117 ( .A(c7223), .B(b[7223]), .Z(n21670) );
XNOR U36118 ( .A(b[7223]), .B(n21671), .Z(c[7223]) );
XNOR U36119 ( .A(a[7223]), .B(c7223), .Z(n21671) );
XOR U36120 ( .A(c7224), .B(n21672), .Z(c7225) );
ANDN U36121 ( .B(n21673), .A(n21674), .Z(n21672) );
XOR U36122 ( .A(c7224), .B(b[7224]), .Z(n21673) );
XNOR U36123 ( .A(b[7224]), .B(n21674), .Z(c[7224]) );
XNOR U36124 ( .A(a[7224]), .B(c7224), .Z(n21674) );
XOR U36125 ( .A(c7225), .B(n21675), .Z(c7226) );
ANDN U36126 ( .B(n21676), .A(n21677), .Z(n21675) );
XOR U36127 ( .A(c7225), .B(b[7225]), .Z(n21676) );
XNOR U36128 ( .A(b[7225]), .B(n21677), .Z(c[7225]) );
XNOR U36129 ( .A(a[7225]), .B(c7225), .Z(n21677) );
XOR U36130 ( .A(c7226), .B(n21678), .Z(c7227) );
ANDN U36131 ( .B(n21679), .A(n21680), .Z(n21678) );
XOR U36132 ( .A(c7226), .B(b[7226]), .Z(n21679) );
XNOR U36133 ( .A(b[7226]), .B(n21680), .Z(c[7226]) );
XNOR U36134 ( .A(a[7226]), .B(c7226), .Z(n21680) );
XOR U36135 ( .A(c7227), .B(n21681), .Z(c7228) );
ANDN U36136 ( .B(n21682), .A(n21683), .Z(n21681) );
XOR U36137 ( .A(c7227), .B(b[7227]), .Z(n21682) );
XNOR U36138 ( .A(b[7227]), .B(n21683), .Z(c[7227]) );
XNOR U36139 ( .A(a[7227]), .B(c7227), .Z(n21683) );
XOR U36140 ( .A(c7228), .B(n21684), .Z(c7229) );
ANDN U36141 ( .B(n21685), .A(n21686), .Z(n21684) );
XOR U36142 ( .A(c7228), .B(b[7228]), .Z(n21685) );
XNOR U36143 ( .A(b[7228]), .B(n21686), .Z(c[7228]) );
XNOR U36144 ( .A(a[7228]), .B(c7228), .Z(n21686) );
XOR U36145 ( .A(c7229), .B(n21687), .Z(c7230) );
ANDN U36146 ( .B(n21688), .A(n21689), .Z(n21687) );
XOR U36147 ( .A(c7229), .B(b[7229]), .Z(n21688) );
XNOR U36148 ( .A(b[7229]), .B(n21689), .Z(c[7229]) );
XNOR U36149 ( .A(a[7229]), .B(c7229), .Z(n21689) );
XOR U36150 ( .A(c7230), .B(n21690), .Z(c7231) );
ANDN U36151 ( .B(n21691), .A(n21692), .Z(n21690) );
XOR U36152 ( .A(c7230), .B(b[7230]), .Z(n21691) );
XNOR U36153 ( .A(b[7230]), .B(n21692), .Z(c[7230]) );
XNOR U36154 ( .A(a[7230]), .B(c7230), .Z(n21692) );
XOR U36155 ( .A(c7231), .B(n21693), .Z(c7232) );
ANDN U36156 ( .B(n21694), .A(n21695), .Z(n21693) );
XOR U36157 ( .A(c7231), .B(b[7231]), .Z(n21694) );
XNOR U36158 ( .A(b[7231]), .B(n21695), .Z(c[7231]) );
XNOR U36159 ( .A(a[7231]), .B(c7231), .Z(n21695) );
XOR U36160 ( .A(c7232), .B(n21696), .Z(c7233) );
ANDN U36161 ( .B(n21697), .A(n21698), .Z(n21696) );
XOR U36162 ( .A(c7232), .B(b[7232]), .Z(n21697) );
XNOR U36163 ( .A(b[7232]), .B(n21698), .Z(c[7232]) );
XNOR U36164 ( .A(a[7232]), .B(c7232), .Z(n21698) );
XOR U36165 ( .A(c7233), .B(n21699), .Z(c7234) );
ANDN U36166 ( .B(n21700), .A(n21701), .Z(n21699) );
XOR U36167 ( .A(c7233), .B(b[7233]), .Z(n21700) );
XNOR U36168 ( .A(b[7233]), .B(n21701), .Z(c[7233]) );
XNOR U36169 ( .A(a[7233]), .B(c7233), .Z(n21701) );
XOR U36170 ( .A(c7234), .B(n21702), .Z(c7235) );
ANDN U36171 ( .B(n21703), .A(n21704), .Z(n21702) );
XOR U36172 ( .A(c7234), .B(b[7234]), .Z(n21703) );
XNOR U36173 ( .A(b[7234]), .B(n21704), .Z(c[7234]) );
XNOR U36174 ( .A(a[7234]), .B(c7234), .Z(n21704) );
XOR U36175 ( .A(c7235), .B(n21705), .Z(c7236) );
ANDN U36176 ( .B(n21706), .A(n21707), .Z(n21705) );
XOR U36177 ( .A(c7235), .B(b[7235]), .Z(n21706) );
XNOR U36178 ( .A(b[7235]), .B(n21707), .Z(c[7235]) );
XNOR U36179 ( .A(a[7235]), .B(c7235), .Z(n21707) );
XOR U36180 ( .A(c7236), .B(n21708), .Z(c7237) );
ANDN U36181 ( .B(n21709), .A(n21710), .Z(n21708) );
XOR U36182 ( .A(c7236), .B(b[7236]), .Z(n21709) );
XNOR U36183 ( .A(b[7236]), .B(n21710), .Z(c[7236]) );
XNOR U36184 ( .A(a[7236]), .B(c7236), .Z(n21710) );
XOR U36185 ( .A(c7237), .B(n21711), .Z(c7238) );
ANDN U36186 ( .B(n21712), .A(n21713), .Z(n21711) );
XOR U36187 ( .A(c7237), .B(b[7237]), .Z(n21712) );
XNOR U36188 ( .A(b[7237]), .B(n21713), .Z(c[7237]) );
XNOR U36189 ( .A(a[7237]), .B(c7237), .Z(n21713) );
XOR U36190 ( .A(c7238), .B(n21714), .Z(c7239) );
ANDN U36191 ( .B(n21715), .A(n21716), .Z(n21714) );
XOR U36192 ( .A(c7238), .B(b[7238]), .Z(n21715) );
XNOR U36193 ( .A(b[7238]), .B(n21716), .Z(c[7238]) );
XNOR U36194 ( .A(a[7238]), .B(c7238), .Z(n21716) );
XOR U36195 ( .A(c7239), .B(n21717), .Z(c7240) );
ANDN U36196 ( .B(n21718), .A(n21719), .Z(n21717) );
XOR U36197 ( .A(c7239), .B(b[7239]), .Z(n21718) );
XNOR U36198 ( .A(b[7239]), .B(n21719), .Z(c[7239]) );
XNOR U36199 ( .A(a[7239]), .B(c7239), .Z(n21719) );
XOR U36200 ( .A(c7240), .B(n21720), .Z(c7241) );
ANDN U36201 ( .B(n21721), .A(n21722), .Z(n21720) );
XOR U36202 ( .A(c7240), .B(b[7240]), .Z(n21721) );
XNOR U36203 ( .A(b[7240]), .B(n21722), .Z(c[7240]) );
XNOR U36204 ( .A(a[7240]), .B(c7240), .Z(n21722) );
XOR U36205 ( .A(c7241), .B(n21723), .Z(c7242) );
ANDN U36206 ( .B(n21724), .A(n21725), .Z(n21723) );
XOR U36207 ( .A(c7241), .B(b[7241]), .Z(n21724) );
XNOR U36208 ( .A(b[7241]), .B(n21725), .Z(c[7241]) );
XNOR U36209 ( .A(a[7241]), .B(c7241), .Z(n21725) );
XOR U36210 ( .A(c7242), .B(n21726), .Z(c7243) );
ANDN U36211 ( .B(n21727), .A(n21728), .Z(n21726) );
XOR U36212 ( .A(c7242), .B(b[7242]), .Z(n21727) );
XNOR U36213 ( .A(b[7242]), .B(n21728), .Z(c[7242]) );
XNOR U36214 ( .A(a[7242]), .B(c7242), .Z(n21728) );
XOR U36215 ( .A(c7243), .B(n21729), .Z(c7244) );
ANDN U36216 ( .B(n21730), .A(n21731), .Z(n21729) );
XOR U36217 ( .A(c7243), .B(b[7243]), .Z(n21730) );
XNOR U36218 ( .A(b[7243]), .B(n21731), .Z(c[7243]) );
XNOR U36219 ( .A(a[7243]), .B(c7243), .Z(n21731) );
XOR U36220 ( .A(c7244), .B(n21732), .Z(c7245) );
ANDN U36221 ( .B(n21733), .A(n21734), .Z(n21732) );
XOR U36222 ( .A(c7244), .B(b[7244]), .Z(n21733) );
XNOR U36223 ( .A(b[7244]), .B(n21734), .Z(c[7244]) );
XNOR U36224 ( .A(a[7244]), .B(c7244), .Z(n21734) );
XOR U36225 ( .A(c7245), .B(n21735), .Z(c7246) );
ANDN U36226 ( .B(n21736), .A(n21737), .Z(n21735) );
XOR U36227 ( .A(c7245), .B(b[7245]), .Z(n21736) );
XNOR U36228 ( .A(b[7245]), .B(n21737), .Z(c[7245]) );
XNOR U36229 ( .A(a[7245]), .B(c7245), .Z(n21737) );
XOR U36230 ( .A(c7246), .B(n21738), .Z(c7247) );
ANDN U36231 ( .B(n21739), .A(n21740), .Z(n21738) );
XOR U36232 ( .A(c7246), .B(b[7246]), .Z(n21739) );
XNOR U36233 ( .A(b[7246]), .B(n21740), .Z(c[7246]) );
XNOR U36234 ( .A(a[7246]), .B(c7246), .Z(n21740) );
XOR U36235 ( .A(c7247), .B(n21741), .Z(c7248) );
ANDN U36236 ( .B(n21742), .A(n21743), .Z(n21741) );
XOR U36237 ( .A(c7247), .B(b[7247]), .Z(n21742) );
XNOR U36238 ( .A(b[7247]), .B(n21743), .Z(c[7247]) );
XNOR U36239 ( .A(a[7247]), .B(c7247), .Z(n21743) );
XOR U36240 ( .A(c7248), .B(n21744), .Z(c7249) );
ANDN U36241 ( .B(n21745), .A(n21746), .Z(n21744) );
XOR U36242 ( .A(c7248), .B(b[7248]), .Z(n21745) );
XNOR U36243 ( .A(b[7248]), .B(n21746), .Z(c[7248]) );
XNOR U36244 ( .A(a[7248]), .B(c7248), .Z(n21746) );
XOR U36245 ( .A(c7249), .B(n21747), .Z(c7250) );
ANDN U36246 ( .B(n21748), .A(n21749), .Z(n21747) );
XOR U36247 ( .A(c7249), .B(b[7249]), .Z(n21748) );
XNOR U36248 ( .A(b[7249]), .B(n21749), .Z(c[7249]) );
XNOR U36249 ( .A(a[7249]), .B(c7249), .Z(n21749) );
XOR U36250 ( .A(c7250), .B(n21750), .Z(c7251) );
ANDN U36251 ( .B(n21751), .A(n21752), .Z(n21750) );
XOR U36252 ( .A(c7250), .B(b[7250]), .Z(n21751) );
XNOR U36253 ( .A(b[7250]), .B(n21752), .Z(c[7250]) );
XNOR U36254 ( .A(a[7250]), .B(c7250), .Z(n21752) );
XOR U36255 ( .A(c7251), .B(n21753), .Z(c7252) );
ANDN U36256 ( .B(n21754), .A(n21755), .Z(n21753) );
XOR U36257 ( .A(c7251), .B(b[7251]), .Z(n21754) );
XNOR U36258 ( .A(b[7251]), .B(n21755), .Z(c[7251]) );
XNOR U36259 ( .A(a[7251]), .B(c7251), .Z(n21755) );
XOR U36260 ( .A(c7252), .B(n21756), .Z(c7253) );
ANDN U36261 ( .B(n21757), .A(n21758), .Z(n21756) );
XOR U36262 ( .A(c7252), .B(b[7252]), .Z(n21757) );
XNOR U36263 ( .A(b[7252]), .B(n21758), .Z(c[7252]) );
XNOR U36264 ( .A(a[7252]), .B(c7252), .Z(n21758) );
XOR U36265 ( .A(c7253), .B(n21759), .Z(c7254) );
ANDN U36266 ( .B(n21760), .A(n21761), .Z(n21759) );
XOR U36267 ( .A(c7253), .B(b[7253]), .Z(n21760) );
XNOR U36268 ( .A(b[7253]), .B(n21761), .Z(c[7253]) );
XNOR U36269 ( .A(a[7253]), .B(c7253), .Z(n21761) );
XOR U36270 ( .A(c7254), .B(n21762), .Z(c7255) );
ANDN U36271 ( .B(n21763), .A(n21764), .Z(n21762) );
XOR U36272 ( .A(c7254), .B(b[7254]), .Z(n21763) );
XNOR U36273 ( .A(b[7254]), .B(n21764), .Z(c[7254]) );
XNOR U36274 ( .A(a[7254]), .B(c7254), .Z(n21764) );
XOR U36275 ( .A(c7255), .B(n21765), .Z(c7256) );
ANDN U36276 ( .B(n21766), .A(n21767), .Z(n21765) );
XOR U36277 ( .A(c7255), .B(b[7255]), .Z(n21766) );
XNOR U36278 ( .A(b[7255]), .B(n21767), .Z(c[7255]) );
XNOR U36279 ( .A(a[7255]), .B(c7255), .Z(n21767) );
XOR U36280 ( .A(c7256), .B(n21768), .Z(c7257) );
ANDN U36281 ( .B(n21769), .A(n21770), .Z(n21768) );
XOR U36282 ( .A(c7256), .B(b[7256]), .Z(n21769) );
XNOR U36283 ( .A(b[7256]), .B(n21770), .Z(c[7256]) );
XNOR U36284 ( .A(a[7256]), .B(c7256), .Z(n21770) );
XOR U36285 ( .A(c7257), .B(n21771), .Z(c7258) );
ANDN U36286 ( .B(n21772), .A(n21773), .Z(n21771) );
XOR U36287 ( .A(c7257), .B(b[7257]), .Z(n21772) );
XNOR U36288 ( .A(b[7257]), .B(n21773), .Z(c[7257]) );
XNOR U36289 ( .A(a[7257]), .B(c7257), .Z(n21773) );
XOR U36290 ( .A(c7258), .B(n21774), .Z(c7259) );
ANDN U36291 ( .B(n21775), .A(n21776), .Z(n21774) );
XOR U36292 ( .A(c7258), .B(b[7258]), .Z(n21775) );
XNOR U36293 ( .A(b[7258]), .B(n21776), .Z(c[7258]) );
XNOR U36294 ( .A(a[7258]), .B(c7258), .Z(n21776) );
XOR U36295 ( .A(c7259), .B(n21777), .Z(c7260) );
ANDN U36296 ( .B(n21778), .A(n21779), .Z(n21777) );
XOR U36297 ( .A(c7259), .B(b[7259]), .Z(n21778) );
XNOR U36298 ( .A(b[7259]), .B(n21779), .Z(c[7259]) );
XNOR U36299 ( .A(a[7259]), .B(c7259), .Z(n21779) );
XOR U36300 ( .A(c7260), .B(n21780), .Z(c7261) );
ANDN U36301 ( .B(n21781), .A(n21782), .Z(n21780) );
XOR U36302 ( .A(c7260), .B(b[7260]), .Z(n21781) );
XNOR U36303 ( .A(b[7260]), .B(n21782), .Z(c[7260]) );
XNOR U36304 ( .A(a[7260]), .B(c7260), .Z(n21782) );
XOR U36305 ( .A(c7261), .B(n21783), .Z(c7262) );
ANDN U36306 ( .B(n21784), .A(n21785), .Z(n21783) );
XOR U36307 ( .A(c7261), .B(b[7261]), .Z(n21784) );
XNOR U36308 ( .A(b[7261]), .B(n21785), .Z(c[7261]) );
XNOR U36309 ( .A(a[7261]), .B(c7261), .Z(n21785) );
XOR U36310 ( .A(c7262), .B(n21786), .Z(c7263) );
ANDN U36311 ( .B(n21787), .A(n21788), .Z(n21786) );
XOR U36312 ( .A(c7262), .B(b[7262]), .Z(n21787) );
XNOR U36313 ( .A(b[7262]), .B(n21788), .Z(c[7262]) );
XNOR U36314 ( .A(a[7262]), .B(c7262), .Z(n21788) );
XOR U36315 ( .A(c7263), .B(n21789), .Z(c7264) );
ANDN U36316 ( .B(n21790), .A(n21791), .Z(n21789) );
XOR U36317 ( .A(c7263), .B(b[7263]), .Z(n21790) );
XNOR U36318 ( .A(b[7263]), .B(n21791), .Z(c[7263]) );
XNOR U36319 ( .A(a[7263]), .B(c7263), .Z(n21791) );
XOR U36320 ( .A(c7264), .B(n21792), .Z(c7265) );
ANDN U36321 ( .B(n21793), .A(n21794), .Z(n21792) );
XOR U36322 ( .A(c7264), .B(b[7264]), .Z(n21793) );
XNOR U36323 ( .A(b[7264]), .B(n21794), .Z(c[7264]) );
XNOR U36324 ( .A(a[7264]), .B(c7264), .Z(n21794) );
XOR U36325 ( .A(c7265), .B(n21795), .Z(c7266) );
ANDN U36326 ( .B(n21796), .A(n21797), .Z(n21795) );
XOR U36327 ( .A(c7265), .B(b[7265]), .Z(n21796) );
XNOR U36328 ( .A(b[7265]), .B(n21797), .Z(c[7265]) );
XNOR U36329 ( .A(a[7265]), .B(c7265), .Z(n21797) );
XOR U36330 ( .A(c7266), .B(n21798), .Z(c7267) );
ANDN U36331 ( .B(n21799), .A(n21800), .Z(n21798) );
XOR U36332 ( .A(c7266), .B(b[7266]), .Z(n21799) );
XNOR U36333 ( .A(b[7266]), .B(n21800), .Z(c[7266]) );
XNOR U36334 ( .A(a[7266]), .B(c7266), .Z(n21800) );
XOR U36335 ( .A(c7267), .B(n21801), .Z(c7268) );
ANDN U36336 ( .B(n21802), .A(n21803), .Z(n21801) );
XOR U36337 ( .A(c7267), .B(b[7267]), .Z(n21802) );
XNOR U36338 ( .A(b[7267]), .B(n21803), .Z(c[7267]) );
XNOR U36339 ( .A(a[7267]), .B(c7267), .Z(n21803) );
XOR U36340 ( .A(c7268), .B(n21804), .Z(c7269) );
ANDN U36341 ( .B(n21805), .A(n21806), .Z(n21804) );
XOR U36342 ( .A(c7268), .B(b[7268]), .Z(n21805) );
XNOR U36343 ( .A(b[7268]), .B(n21806), .Z(c[7268]) );
XNOR U36344 ( .A(a[7268]), .B(c7268), .Z(n21806) );
XOR U36345 ( .A(c7269), .B(n21807), .Z(c7270) );
ANDN U36346 ( .B(n21808), .A(n21809), .Z(n21807) );
XOR U36347 ( .A(c7269), .B(b[7269]), .Z(n21808) );
XNOR U36348 ( .A(b[7269]), .B(n21809), .Z(c[7269]) );
XNOR U36349 ( .A(a[7269]), .B(c7269), .Z(n21809) );
XOR U36350 ( .A(c7270), .B(n21810), .Z(c7271) );
ANDN U36351 ( .B(n21811), .A(n21812), .Z(n21810) );
XOR U36352 ( .A(c7270), .B(b[7270]), .Z(n21811) );
XNOR U36353 ( .A(b[7270]), .B(n21812), .Z(c[7270]) );
XNOR U36354 ( .A(a[7270]), .B(c7270), .Z(n21812) );
XOR U36355 ( .A(c7271), .B(n21813), .Z(c7272) );
ANDN U36356 ( .B(n21814), .A(n21815), .Z(n21813) );
XOR U36357 ( .A(c7271), .B(b[7271]), .Z(n21814) );
XNOR U36358 ( .A(b[7271]), .B(n21815), .Z(c[7271]) );
XNOR U36359 ( .A(a[7271]), .B(c7271), .Z(n21815) );
XOR U36360 ( .A(c7272), .B(n21816), .Z(c7273) );
ANDN U36361 ( .B(n21817), .A(n21818), .Z(n21816) );
XOR U36362 ( .A(c7272), .B(b[7272]), .Z(n21817) );
XNOR U36363 ( .A(b[7272]), .B(n21818), .Z(c[7272]) );
XNOR U36364 ( .A(a[7272]), .B(c7272), .Z(n21818) );
XOR U36365 ( .A(c7273), .B(n21819), .Z(c7274) );
ANDN U36366 ( .B(n21820), .A(n21821), .Z(n21819) );
XOR U36367 ( .A(c7273), .B(b[7273]), .Z(n21820) );
XNOR U36368 ( .A(b[7273]), .B(n21821), .Z(c[7273]) );
XNOR U36369 ( .A(a[7273]), .B(c7273), .Z(n21821) );
XOR U36370 ( .A(c7274), .B(n21822), .Z(c7275) );
ANDN U36371 ( .B(n21823), .A(n21824), .Z(n21822) );
XOR U36372 ( .A(c7274), .B(b[7274]), .Z(n21823) );
XNOR U36373 ( .A(b[7274]), .B(n21824), .Z(c[7274]) );
XNOR U36374 ( .A(a[7274]), .B(c7274), .Z(n21824) );
XOR U36375 ( .A(c7275), .B(n21825), .Z(c7276) );
ANDN U36376 ( .B(n21826), .A(n21827), .Z(n21825) );
XOR U36377 ( .A(c7275), .B(b[7275]), .Z(n21826) );
XNOR U36378 ( .A(b[7275]), .B(n21827), .Z(c[7275]) );
XNOR U36379 ( .A(a[7275]), .B(c7275), .Z(n21827) );
XOR U36380 ( .A(c7276), .B(n21828), .Z(c7277) );
ANDN U36381 ( .B(n21829), .A(n21830), .Z(n21828) );
XOR U36382 ( .A(c7276), .B(b[7276]), .Z(n21829) );
XNOR U36383 ( .A(b[7276]), .B(n21830), .Z(c[7276]) );
XNOR U36384 ( .A(a[7276]), .B(c7276), .Z(n21830) );
XOR U36385 ( .A(c7277), .B(n21831), .Z(c7278) );
ANDN U36386 ( .B(n21832), .A(n21833), .Z(n21831) );
XOR U36387 ( .A(c7277), .B(b[7277]), .Z(n21832) );
XNOR U36388 ( .A(b[7277]), .B(n21833), .Z(c[7277]) );
XNOR U36389 ( .A(a[7277]), .B(c7277), .Z(n21833) );
XOR U36390 ( .A(c7278), .B(n21834), .Z(c7279) );
ANDN U36391 ( .B(n21835), .A(n21836), .Z(n21834) );
XOR U36392 ( .A(c7278), .B(b[7278]), .Z(n21835) );
XNOR U36393 ( .A(b[7278]), .B(n21836), .Z(c[7278]) );
XNOR U36394 ( .A(a[7278]), .B(c7278), .Z(n21836) );
XOR U36395 ( .A(c7279), .B(n21837), .Z(c7280) );
ANDN U36396 ( .B(n21838), .A(n21839), .Z(n21837) );
XOR U36397 ( .A(c7279), .B(b[7279]), .Z(n21838) );
XNOR U36398 ( .A(b[7279]), .B(n21839), .Z(c[7279]) );
XNOR U36399 ( .A(a[7279]), .B(c7279), .Z(n21839) );
XOR U36400 ( .A(c7280), .B(n21840), .Z(c7281) );
ANDN U36401 ( .B(n21841), .A(n21842), .Z(n21840) );
XOR U36402 ( .A(c7280), .B(b[7280]), .Z(n21841) );
XNOR U36403 ( .A(b[7280]), .B(n21842), .Z(c[7280]) );
XNOR U36404 ( .A(a[7280]), .B(c7280), .Z(n21842) );
XOR U36405 ( .A(c7281), .B(n21843), .Z(c7282) );
ANDN U36406 ( .B(n21844), .A(n21845), .Z(n21843) );
XOR U36407 ( .A(c7281), .B(b[7281]), .Z(n21844) );
XNOR U36408 ( .A(b[7281]), .B(n21845), .Z(c[7281]) );
XNOR U36409 ( .A(a[7281]), .B(c7281), .Z(n21845) );
XOR U36410 ( .A(c7282), .B(n21846), .Z(c7283) );
ANDN U36411 ( .B(n21847), .A(n21848), .Z(n21846) );
XOR U36412 ( .A(c7282), .B(b[7282]), .Z(n21847) );
XNOR U36413 ( .A(b[7282]), .B(n21848), .Z(c[7282]) );
XNOR U36414 ( .A(a[7282]), .B(c7282), .Z(n21848) );
XOR U36415 ( .A(c7283), .B(n21849), .Z(c7284) );
ANDN U36416 ( .B(n21850), .A(n21851), .Z(n21849) );
XOR U36417 ( .A(c7283), .B(b[7283]), .Z(n21850) );
XNOR U36418 ( .A(b[7283]), .B(n21851), .Z(c[7283]) );
XNOR U36419 ( .A(a[7283]), .B(c7283), .Z(n21851) );
XOR U36420 ( .A(c7284), .B(n21852), .Z(c7285) );
ANDN U36421 ( .B(n21853), .A(n21854), .Z(n21852) );
XOR U36422 ( .A(c7284), .B(b[7284]), .Z(n21853) );
XNOR U36423 ( .A(b[7284]), .B(n21854), .Z(c[7284]) );
XNOR U36424 ( .A(a[7284]), .B(c7284), .Z(n21854) );
XOR U36425 ( .A(c7285), .B(n21855), .Z(c7286) );
ANDN U36426 ( .B(n21856), .A(n21857), .Z(n21855) );
XOR U36427 ( .A(c7285), .B(b[7285]), .Z(n21856) );
XNOR U36428 ( .A(b[7285]), .B(n21857), .Z(c[7285]) );
XNOR U36429 ( .A(a[7285]), .B(c7285), .Z(n21857) );
XOR U36430 ( .A(c7286), .B(n21858), .Z(c7287) );
ANDN U36431 ( .B(n21859), .A(n21860), .Z(n21858) );
XOR U36432 ( .A(c7286), .B(b[7286]), .Z(n21859) );
XNOR U36433 ( .A(b[7286]), .B(n21860), .Z(c[7286]) );
XNOR U36434 ( .A(a[7286]), .B(c7286), .Z(n21860) );
XOR U36435 ( .A(c7287), .B(n21861), .Z(c7288) );
ANDN U36436 ( .B(n21862), .A(n21863), .Z(n21861) );
XOR U36437 ( .A(c7287), .B(b[7287]), .Z(n21862) );
XNOR U36438 ( .A(b[7287]), .B(n21863), .Z(c[7287]) );
XNOR U36439 ( .A(a[7287]), .B(c7287), .Z(n21863) );
XOR U36440 ( .A(c7288), .B(n21864), .Z(c7289) );
ANDN U36441 ( .B(n21865), .A(n21866), .Z(n21864) );
XOR U36442 ( .A(c7288), .B(b[7288]), .Z(n21865) );
XNOR U36443 ( .A(b[7288]), .B(n21866), .Z(c[7288]) );
XNOR U36444 ( .A(a[7288]), .B(c7288), .Z(n21866) );
XOR U36445 ( .A(c7289), .B(n21867), .Z(c7290) );
ANDN U36446 ( .B(n21868), .A(n21869), .Z(n21867) );
XOR U36447 ( .A(c7289), .B(b[7289]), .Z(n21868) );
XNOR U36448 ( .A(b[7289]), .B(n21869), .Z(c[7289]) );
XNOR U36449 ( .A(a[7289]), .B(c7289), .Z(n21869) );
XOR U36450 ( .A(c7290), .B(n21870), .Z(c7291) );
ANDN U36451 ( .B(n21871), .A(n21872), .Z(n21870) );
XOR U36452 ( .A(c7290), .B(b[7290]), .Z(n21871) );
XNOR U36453 ( .A(b[7290]), .B(n21872), .Z(c[7290]) );
XNOR U36454 ( .A(a[7290]), .B(c7290), .Z(n21872) );
XOR U36455 ( .A(c7291), .B(n21873), .Z(c7292) );
ANDN U36456 ( .B(n21874), .A(n21875), .Z(n21873) );
XOR U36457 ( .A(c7291), .B(b[7291]), .Z(n21874) );
XNOR U36458 ( .A(b[7291]), .B(n21875), .Z(c[7291]) );
XNOR U36459 ( .A(a[7291]), .B(c7291), .Z(n21875) );
XOR U36460 ( .A(c7292), .B(n21876), .Z(c7293) );
ANDN U36461 ( .B(n21877), .A(n21878), .Z(n21876) );
XOR U36462 ( .A(c7292), .B(b[7292]), .Z(n21877) );
XNOR U36463 ( .A(b[7292]), .B(n21878), .Z(c[7292]) );
XNOR U36464 ( .A(a[7292]), .B(c7292), .Z(n21878) );
XOR U36465 ( .A(c7293), .B(n21879), .Z(c7294) );
ANDN U36466 ( .B(n21880), .A(n21881), .Z(n21879) );
XOR U36467 ( .A(c7293), .B(b[7293]), .Z(n21880) );
XNOR U36468 ( .A(b[7293]), .B(n21881), .Z(c[7293]) );
XNOR U36469 ( .A(a[7293]), .B(c7293), .Z(n21881) );
XOR U36470 ( .A(c7294), .B(n21882), .Z(c7295) );
ANDN U36471 ( .B(n21883), .A(n21884), .Z(n21882) );
XOR U36472 ( .A(c7294), .B(b[7294]), .Z(n21883) );
XNOR U36473 ( .A(b[7294]), .B(n21884), .Z(c[7294]) );
XNOR U36474 ( .A(a[7294]), .B(c7294), .Z(n21884) );
XOR U36475 ( .A(c7295), .B(n21885), .Z(c7296) );
ANDN U36476 ( .B(n21886), .A(n21887), .Z(n21885) );
XOR U36477 ( .A(c7295), .B(b[7295]), .Z(n21886) );
XNOR U36478 ( .A(b[7295]), .B(n21887), .Z(c[7295]) );
XNOR U36479 ( .A(a[7295]), .B(c7295), .Z(n21887) );
XOR U36480 ( .A(c7296), .B(n21888), .Z(c7297) );
ANDN U36481 ( .B(n21889), .A(n21890), .Z(n21888) );
XOR U36482 ( .A(c7296), .B(b[7296]), .Z(n21889) );
XNOR U36483 ( .A(b[7296]), .B(n21890), .Z(c[7296]) );
XNOR U36484 ( .A(a[7296]), .B(c7296), .Z(n21890) );
XOR U36485 ( .A(c7297), .B(n21891), .Z(c7298) );
ANDN U36486 ( .B(n21892), .A(n21893), .Z(n21891) );
XOR U36487 ( .A(c7297), .B(b[7297]), .Z(n21892) );
XNOR U36488 ( .A(b[7297]), .B(n21893), .Z(c[7297]) );
XNOR U36489 ( .A(a[7297]), .B(c7297), .Z(n21893) );
XOR U36490 ( .A(c7298), .B(n21894), .Z(c7299) );
ANDN U36491 ( .B(n21895), .A(n21896), .Z(n21894) );
XOR U36492 ( .A(c7298), .B(b[7298]), .Z(n21895) );
XNOR U36493 ( .A(b[7298]), .B(n21896), .Z(c[7298]) );
XNOR U36494 ( .A(a[7298]), .B(c7298), .Z(n21896) );
XOR U36495 ( .A(c7299), .B(n21897), .Z(c7300) );
ANDN U36496 ( .B(n21898), .A(n21899), .Z(n21897) );
XOR U36497 ( .A(c7299), .B(b[7299]), .Z(n21898) );
XNOR U36498 ( .A(b[7299]), .B(n21899), .Z(c[7299]) );
XNOR U36499 ( .A(a[7299]), .B(c7299), .Z(n21899) );
XOR U36500 ( .A(c7300), .B(n21900), .Z(c7301) );
ANDN U36501 ( .B(n21901), .A(n21902), .Z(n21900) );
XOR U36502 ( .A(c7300), .B(b[7300]), .Z(n21901) );
XNOR U36503 ( .A(b[7300]), .B(n21902), .Z(c[7300]) );
XNOR U36504 ( .A(a[7300]), .B(c7300), .Z(n21902) );
XOR U36505 ( .A(c7301), .B(n21903), .Z(c7302) );
ANDN U36506 ( .B(n21904), .A(n21905), .Z(n21903) );
XOR U36507 ( .A(c7301), .B(b[7301]), .Z(n21904) );
XNOR U36508 ( .A(b[7301]), .B(n21905), .Z(c[7301]) );
XNOR U36509 ( .A(a[7301]), .B(c7301), .Z(n21905) );
XOR U36510 ( .A(c7302), .B(n21906), .Z(c7303) );
ANDN U36511 ( .B(n21907), .A(n21908), .Z(n21906) );
XOR U36512 ( .A(c7302), .B(b[7302]), .Z(n21907) );
XNOR U36513 ( .A(b[7302]), .B(n21908), .Z(c[7302]) );
XNOR U36514 ( .A(a[7302]), .B(c7302), .Z(n21908) );
XOR U36515 ( .A(c7303), .B(n21909), .Z(c7304) );
ANDN U36516 ( .B(n21910), .A(n21911), .Z(n21909) );
XOR U36517 ( .A(c7303), .B(b[7303]), .Z(n21910) );
XNOR U36518 ( .A(b[7303]), .B(n21911), .Z(c[7303]) );
XNOR U36519 ( .A(a[7303]), .B(c7303), .Z(n21911) );
XOR U36520 ( .A(c7304), .B(n21912), .Z(c7305) );
ANDN U36521 ( .B(n21913), .A(n21914), .Z(n21912) );
XOR U36522 ( .A(c7304), .B(b[7304]), .Z(n21913) );
XNOR U36523 ( .A(b[7304]), .B(n21914), .Z(c[7304]) );
XNOR U36524 ( .A(a[7304]), .B(c7304), .Z(n21914) );
XOR U36525 ( .A(c7305), .B(n21915), .Z(c7306) );
ANDN U36526 ( .B(n21916), .A(n21917), .Z(n21915) );
XOR U36527 ( .A(c7305), .B(b[7305]), .Z(n21916) );
XNOR U36528 ( .A(b[7305]), .B(n21917), .Z(c[7305]) );
XNOR U36529 ( .A(a[7305]), .B(c7305), .Z(n21917) );
XOR U36530 ( .A(c7306), .B(n21918), .Z(c7307) );
ANDN U36531 ( .B(n21919), .A(n21920), .Z(n21918) );
XOR U36532 ( .A(c7306), .B(b[7306]), .Z(n21919) );
XNOR U36533 ( .A(b[7306]), .B(n21920), .Z(c[7306]) );
XNOR U36534 ( .A(a[7306]), .B(c7306), .Z(n21920) );
XOR U36535 ( .A(c7307), .B(n21921), .Z(c7308) );
ANDN U36536 ( .B(n21922), .A(n21923), .Z(n21921) );
XOR U36537 ( .A(c7307), .B(b[7307]), .Z(n21922) );
XNOR U36538 ( .A(b[7307]), .B(n21923), .Z(c[7307]) );
XNOR U36539 ( .A(a[7307]), .B(c7307), .Z(n21923) );
XOR U36540 ( .A(c7308), .B(n21924), .Z(c7309) );
ANDN U36541 ( .B(n21925), .A(n21926), .Z(n21924) );
XOR U36542 ( .A(c7308), .B(b[7308]), .Z(n21925) );
XNOR U36543 ( .A(b[7308]), .B(n21926), .Z(c[7308]) );
XNOR U36544 ( .A(a[7308]), .B(c7308), .Z(n21926) );
XOR U36545 ( .A(c7309), .B(n21927), .Z(c7310) );
ANDN U36546 ( .B(n21928), .A(n21929), .Z(n21927) );
XOR U36547 ( .A(c7309), .B(b[7309]), .Z(n21928) );
XNOR U36548 ( .A(b[7309]), .B(n21929), .Z(c[7309]) );
XNOR U36549 ( .A(a[7309]), .B(c7309), .Z(n21929) );
XOR U36550 ( .A(c7310), .B(n21930), .Z(c7311) );
ANDN U36551 ( .B(n21931), .A(n21932), .Z(n21930) );
XOR U36552 ( .A(c7310), .B(b[7310]), .Z(n21931) );
XNOR U36553 ( .A(b[7310]), .B(n21932), .Z(c[7310]) );
XNOR U36554 ( .A(a[7310]), .B(c7310), .Z(n21932) );
XOR U36555 ( .A(c7311), .B(n21933), .Z(c7312) );
ANDN U36556 ( .B(n21934), .A(n21935), .Z(n21933) );
XOR U36557 ( .A(c7311), .B(b[7311]), .Z(n21934) );
XNOR U36558 ( .A(b[7311]), .B(n21935), .Z(c[7311]) );
XNOR U36559 ( .A(a[7311]), .B(c7311), .Z(n21935) );
XOR U36560 ( .A(c7312), .B(n21936), .Z(c7313) );
ANDN U36561 ( .B(n21937), .A(n21938), .Z(n21936) );
XOR U36562 ( .A(c7312), .B(b[7312]), .Z(n21937) );
XNOR U36563 ( .A(b[7312]), .B(n21938), .Z(c[7312]) );
XNOR U36564 ( .A(a[7312]), .B(c7312), .Z(n21938) );
XOR U36565 ( .A(c7313), .B(n21939), .Z(c7314) );
ANDN U36566 ( .B(n21940), .A(n21941), .Z(n21939) );
XOR U36567 ( .A(c7313), .B(b[7313]), .Z(n21940) );
XNOR U36568 ( .A(b[7313]), .B(n21941), .Z(c[7313]) );
XNOR U36569 ( .A(a[7313]), .B(c7313), .Z(n21941) );
XOR U36570 ( .A(c7314), .B(n21942), .Z(c7315) );
ANDN U36571 ( .B(n21943), .A(n21944), .Z(n21942) );
XOR U36572 ( .A(c7314), .B(b[7314]), .Z(n21943) );
XNOR U36573 ( .A(b[7314]), .B(n21944), .Z(c[7314]) );
XNOR U36574 ( .A(a[7314]), .B(c7314), .Z(n21944) );
XOR U36575 ( .A(c7315), .B(n21945), .Z(c7316) );
ANDN U36576 ( .B(n21946), .A(n21947), .Z(n21945) );
XOR U36577 ( .A(c7315), .B(b[7315]), .Z(n21946) );
XNOR U36578 ( .A(b[7315]), .B(n21947), .Z(c[7315]) );
XNOR U36579 ( .A(a[7315]), .B(c7315), .Z(n21947) );
XOR U36580 ( .A(c7316), .B(n21948), .Z(c7317) );
ANDN U36581 ( .B(n21949), .A(n21950), .Z(n21948) );
XOR U36582 ( .A(c7316), .B(b[7316]), .Z(n21949) );
XNOR U36583 ( .A(b[7316]), .B(n21950), .Z(c[7316]) );
XNOR U36584 ( .A(a[7316]), .B(c7316), .Z(n21950) );
XOR U36585 ( .A(c7317), .B(n21951), .Z(c7318) );
ANDN U36586 ( .B(n21952), .A(n21953), .Z(n21951) );
XOR U36587 ( .A(c7317), .B(b[7317]), .Z(n21952) );
XNOR U36588 ( .A(b[7317]), .B(n21953), .Z(c[7317]) );
XNOR U36589 ( .A(a[7317]), .B(c7317), .Z(n21953) );
XOR U36590 ( .A(c7318), .B(n21954), .Z(c7319) );
ANDN U36591 ( .B(n21955), .A(n21956), .Z(n21954) );
XOR U36592 ( .A(c7318), .B(b[7318]), .Z(n21955) );
XNOR U36593 ( .A(b[7318]), .B(n21956), .Z(c[7318]) );
XNOR U36594 ( .A(a[7318]), .B(c7318), .Z(n21956) );
XOR U36595 ( .A(c7319), .B(n21957), .Z(c7320) );
ANDN U36596 ( .B(n21958), .A(n21959), .Z(n21957) );
XOR U36597 ( .A(c7319), .B(b[7319]), .Z(n21958) );
XNOR U36598 ( .A(b[7319]), .B(n21959), .Z(c[7319]) );
XNOR U36599 ( .A(a[7319]), .B(c7319), .Z(n21959) );
XOR U36600 ( .A(c7320), .B(n21960), .Z(c7321) );
ANDN U36601 ( .B(n21961), .A(n21962), .Z(n21960) );
XOR U36602 ( .A(c7320), .B(b[7320]), .Z(n21961) );
XNOR U36603 ( .A(b[7320]), .B(n21962), .Z(c[7320]) );
XNOR U36604 ( .A(a[7320]), .B(c7320), .Z(n21962) );
XOR U36605 ( .A(c7321), .B(n21963), .Z(c7322) );
ANDN U36606 ( .B(n21964), .A(n21965), .Z(n21963) );
XOR U36607 ( .A(c7321), .B(b[7321]), .Z(n21964) );
XNOR U36608 ( .A(b[7321]), .B(n21965), .Z(c[7321]) );
XNOR U36609 ( .A(a[7321]), .B(c7321), .Z(n21965) );
XOR U36610 ( .A(c7322), .B(n21966), .Z(c7323) );
ANDN U36611 ( .B(n21967), .A(n21968), .Z(n21966) );
XOR U36612 ( .A(c7322), .B(b[7322]), .Z(n21967) );
XNOR U36613 ( .A(b[7322]), .B(n21968), .Z(c[7322]) );
XNOR U36614 ( .A(a[7322]), .B(c7322), .Z(n21968) );
XOR U36615 ( .A(c7323), .B(n21969), .Z(c7324) );
ANDN U36616 ( .B(n21970), .A(n21971), .Z(n21969) );
XOR U36617 ( .A(c7323), .B(b[7323]), .Z(n21970) );
XNOR U36618 ( .A(b[7323]), .B(n21971), .Z(c[7323]) );
XNOR U36619 ( .A(a[7323]), .B(c7323), .Z(n21971) );
XOR U36620 ( .A(c7324), .B(n21972), .Z(c7325) );
ANDN U36621 ( .B(n21973), .A(n21974), .Z(n21972) );
XOR U36622 ( .A(c7324), .B(b[7324]), .Z(n21973) );
XNOR U36623 ( .A(b[7324]), .B(n21974), .Z(c[7324]) );
XNOR U36624 ( .A(a[7324]), .B(c7324), .Z(n21974) );
XOR U36625 ( .A(c7325), .B(n21975), .Z(c7326) );
ANDN U36626 ( .B(n21976), .A(n21977), .Z(n21975) );
XOR U36627 ( .A(c7325), .B(b[7325]), .Z(n21976) );
XNOR U36628 ( .A(b[7325]), .B(n21977), .Z(c[7325]) );
XNOR U36629 ( .A(a[7325]), .B(c7325), .Z(n21977) );
XOR U36630 ( .A(c7326), .B(n21978), .Z(c7327) );
ANDN U36631 ( .B(n21979), .A(n21980), .Z(n21978) );
XOR U36632 ( .A(c7326), .B(b[7326]), .Z(n21979) );
XNOR U36633 ( .A(b[7326]), .B(n21980), .Z(c[7326]) );
XNOR U36634 ( .A(a[7326]), .B(c7326), .Z(n21980) );
XOR U36635 ( .A(c7327), .B(n21981), .Z(c7328) );
ANDN U36636 ( .B(n21982), .A(n21983), .Z(n21981) );
XOR U36637 ( .A(c7327), .B(b[7327]), .Z(n21982) );
XNOR U36638 ( .A(b[7327]), .B(n21983), .Z(c[7327]) );
XNOR U36639 ( .A(a[7327]), .B(c7327), .Z(n21983) );
XOR U36640 ( .A(c7328), .B(n21984), .Z(c7329) );
ANDN U36641 ( .B(n21985), .A(n21986), .Z(n21984) );
XOR U36642 ( .A(c7328), .B(b[7328]), .Z(n21985) );
XNOR U36643 ( .A(b[7328]), .B(n21986), .Z(c[7328]) );
XNOR U36644 ( .A(a[7328]), .B(c7328), .Z(n21986) );
XOR U36645 ( .A(c7329), .B(n21987), .Z(c7330) );
ANDN U36646 ( .B(n21988), .A(n21989), .Z(n21987) );
XOR U36647 ( .A(c7329), .B(b[7329]), .Z(n21988) );
XNOR U36648 ( .A(b[7329]), .B(n21989), .Z(c[7329]) );
XNOR U36649 ( .A(a[7329]), .B(c7329), .Z(n21989) );
XOR U36650 ( .A(c7330), .B(n21990), .Z(c7331) );
ANDN U36651 ( .B(n21991), .A(n21992), .Z(n21990) );
XOR U36652 ( .A(c7330), .B(b[7330]), .Z(n21991) );
XNOR U36653 ( .A(b[7330]), .B(n21992), .Z(c[7330]) );
XNOR U36654 ( .A(a[7330]), .B(c7330), .Z(n21992) );
XOR U36655 ( .A(c7331), .B(n21993), .Z(c7332) );
ANDN U36656 ( .B(n21994), .A(n21995), .Z(n21993) );
XOR U36657 ( .A(c7331), .B(b[7331]), .Z(n21994) );
XNOR U36658 ( .A(b[7331]), .B(n21995), .Z(c[7331]) );
XNOR U36659 ( .A(a[7331]), .B(c7331), .Z(n21995) );
XOR U36660 ( .A(c7332), .B(n21996), .Z(c7333) );
ANDN U36661 ( .B(n21997), .A(n21998), .Z(n21996) );
XOR U36662 ( .A(c7332), .B(b[7332]), .Z(n21997) );
XNOR U36663 ( .A(b[7332]), .B(n21998), .Z(c[7332]) );
XNOR U36664 ( .A(a[7332]), .B(c7332), .Z(n21998) );
XOR U36665 ( .A(c7333), .B(n21999), .Z(c7334) );
ANDN U36666 ( .B(n22000), .A(n22001), .Z(n21999) );
XOR U36667 ( .A(c7333), .B(b[7333]), .Z(n22000) );
XNOR U36668 ( .A(b[7333]), .B(n22001), .Z(c[7333]) );
XNOR U36669 ( .A(a[7333]), .B(c7333), .Z(n22001) );
XOR U36670 ( .A(c7334), .B(n22002), .Z(c7335) );
ANDN U36671 ( .B(n22003), .A(n22004), .Z(n22002) );
XOR U36672 ( .A(c7334), .B(b[7334]), .Z(n22003) );
XNOR U36673 ( .A(b[7334]), .B(n22004), .Z(c[7334]) );
XNOR U36674 ( .A(a[7334]), .B(c7334), .Z(n22004) );
XOR U36675 ( .A(c7335), .B(n22005), .Z(c7336) );
ANDN U36676 ( .B(n22006), .A(n22007), .Z(n22005) );
XOR U36677 ( .A(c7335), .B(b[7335]), .Z(n22006) );
XNOR U36678 ( .A(b[7335]), .B(n22007), .Z(c[7335]) );
XNOR U36679 ( .A(a[7335]), .B(c7335), .Z(n22007) );
XOR U36680 ( .A(c7336), .B(n22008), .Z(c7337) );
ANDN U36681 ( .B(n22009), .A(n22010), .Z(n22008) );
XOR U36682 ( .A(c7336), .B(b[7336]), .Z(n22009) );
XNOR U36683 ( .A(b[7336]), .B(n22010), .Z(c[7336]) );
XNOR U36684 ( .A(a[7336]), .B(c7336), .Z(n22010) );
XOR U36685 ( .A(c7337), .B(n22011), .Z(c7338) );
ANDN U36686 ( .B(n22012), .A(n22013), .Z(n22011) );
XOR U36687 ( .A(c7337), .B(b[7337]), .Z(n22012) );
XNOR U36688 ( .A(b[7337]), .B(n22013), .Z(c[7337]) );
XNOR U36689 ( .A(a[7337]), .B(c7337), .Z(n22013) );
XOR U36690 ( .A(c7338), .B(n22014), .Z(c7339) );
ANDN U36691 ( .B(n22015), .A(n22016), .Z(n22014) );
XOR U36692 ( .A(c7338), .B(b[7338]), .Z(n22015) );
XNOR U36693 ( .A(b[7338]), .B(n22016), .Z(c[7338]) );
XNOR U36694 ( .A(a[7338]), .B(c7338), .Z(n22016) );
XOR U36695 ( .A(c7339), .B(n22017), .Z(c7340) );
ANDN U36696 ( .B(n22018), .A(n22019), .Z(n22017) );
XOR U36697 ( .A(c7339), .B(b[7339]), .Z(n22018) );
XNOR U36698 ( .A(b[7339]), .B(n22019), .Z(c[7339]) );
XNOR U36699 ( .A(a[7339]), .B(c7339), .Z(n22019) );
XOR U36700 ( .A(c7340), .B(n22020), .Z(c7341) );
ANDN U36701 ( .B(n22021), .A(n22022), .Z(n22020) );
XOR U36702 ( .A(c7340), .B(b[7340]), .Z(n22021) );
XNOR U36703 ( .A(b[7340]), .B(n22022), .Z(c[7340]) );
XNOR U36704 ( .A(a[7340]), .B(c7340), .Z(n22022) );
XOR U36705 ( .A(c7341), .B(n22023), .Z(c7342) );
ANDN U36706 ( .B(n22024), .A(n22025), .Z(n22023) );
XOR U36707 ( .A(c7341), .B(b[7341]), .Z(n22024) );
XNOR U36708 ( .A(b[7341]), .B(n22025), .Z(c[7341]) );
XNOR U36709 ( .A(a[7341]), .B(c7341), .Z(n22025) );
XOR U36710 ( .A(c7342), .B(n22026), .Z(c7343) );
ANDN U36711 ( .B(n22027), .A(n22028), .Z(n22026) );
XOR U36712 ( .A(c7342), .B(b[7342]), .Z(n22027) );
XNOR U36713 ( .A(b[7342]), .B(n22028), .Z(c[7342]) );
XNOR U36714 ( .A(a[7342]), .B(c7342), .Z(n22028) );
XOR U36715 ( .A(c7343), .B(n22029), .Z(c7344) );
ANDN U36716 ( .B(n22030), .A(n22031), .Z(n22029) );
XOR U36717 ( .A(c7343), .B(b[7343]), .Z(n22030) );
XNOR U36718 ( .A(b[7343]), .B(n22031), .Z(c[7343]) );
XNOR U36719 ( .A(a[7343]), .B(c7343), .Z(n22031) );
XOR U36720 ( .A(c7344), .B(n22032), .Z(c7345) );
ANDN U36721 ( .B(n22033), .A(n22034), .Z(n22032) );
XOR U36722 ( .A(c7344), .B(b[7344]), .Z(n22033) );
XNOR U36723 ( .A(b[7344]), .B(n22034), .Z(c[7344]) );
XNOR U36724 ( .A(a[7344]), .B(c7344), .Z(n22034) );
XOR U36725 ( .A(c7345), .B(n22035), .Z(c7346) );
ANDN U36726 ( .B(n22036), .A(n22037), .Z(n22035) );
XOR U36727 ( .A(c7345), .B(b[7345]), .Z(n22036) );
XNOR U36728 ( .A(b[7345]), .B(n22037), .Z(c[7345]) );
XNOR U36729 ( .A(a[7345]), .B(c7345), .Z(n22037) );
XOR U36730 ( .A(c7346), .B(n22038), .Z(c7347) );
ANDN U36731 ( .B(n22039), .A(n22040), .Z(n22038) );
XOR U36732 ( .A(c7346), .B(b[7346]), .Z(n22039) );
XNOR U36733 ( .A(b[7346]), .B(n22040), .Z(c[7346]) );
XNOR U36734 ( .A(a[7346]), .B(c7346), .Z(n22040) );
XOR U36735 ( .A(c7347), .B(n22041), .Z(c7348) );
ANDN U36736 ( .B(n22042), .A(n22043), .Z(n22041) );
XOR U36737 ( .A(c7347), .B(b[7347]), .Z(n22042) );
XNOR U36738 ( .A(b[7347]), .B(n22043), .Z(c[7347]) );
XNOR U36739 ( .A(a[7347]), .B(c7347), .Z(n22043) );
XOR U36740 ( .A(c7348), .B(n22044), .Z(c7349) );
ANDN U36741 ( .B(n22045), .A(n22046), .Z(n22044) );
XOR U36742 ( .A(c7348), .B(b[7348]), .Z(n22045) );
XNOR U36743 ( .A(b[7348]), .B(n22046), .Z(c[7348]) );
XNOR U36744 ( .A(a[7348]), .B(c7348), .Z(n22046) );
XOR U36745 ( .A(c7349), .B(n22047), .Z(c7350) );
ANDN U36746 ( .B(n22048), .A(n22049), .Z(n22047) );
XOR U36747 ( .A(c7349), .B(b[7349]), .Z(n22048) );
XNOR U36748 ( .A(b[7349]), .B(n22049), .Z(c[7349]) );
XNOR U36749 ( .A(a[7349]), .B(c7349), .Z(n22049) );
XOR U36750 ( .A(c7350), .B(n22050), .Z(c7351) );
ANDN U36751 ( .B(n22051), .A(n22052), .Z(n22050) );
XOR U36752 ( .A(c7350), .B(b[7350]), .Z(n22051) );
XNOR U36753 ( .A(b[7350]), .B(n22052), .Z(c[7350]) );
XNOR U36754 ( .A(a[7350]), .B(c7350), .Z(n22052) );
XOR U36755 ( .A(c7351), .B(n22053), .Z(c7352) );
ANDN U36756 ( .B(n22054), .A(n22055), .Z(n22053) );
XOR U36757 ( .A(c7351), .B(b[7351]), .Z(n22054) );
XNOR U36758 ( .A(b[7351]), .B(n22055), .Z(c[7351]) );
XNOR U36759 ( .A(a[7351]), .B(c7351), .Z(n22055) );
XOR U36760 ( .A(c7352), .B(n22056), .Z(c7353) );
ANDN U36761 ( .B(n22057), .A(n22058), .Z(n22056) );
XOR U36762 ( .A(c7352), .B(b[7352]), .Z(n22057) );
XNOR U36763 ( .A(b[7352]), .B(n22058), .Z(c[7352]) );
XNOR U36764 ( .A(a[7352]), .B(c7352), .Z(n22058) );
XOR U36765 ( .A(c7353), .B(n22059), .Z(c7354) );
ANDN U36766 ( .B(n22060), .A(n22061), .Z(n22059) );
XOR U36767 ( .A(c7353), .B(b[7353]), .Z(n22060) );
XNOR U36768 ( .A(b[7353]), .B(n22061), .Z(c[7353]) );
XNOR U36769 ( .A(a[7353]), .B(c7353), .Z(n22061) );
XOR U36770 ( .A(c7354), .B(n22062), .Z(c7355) );
ANDN U36771 ( .B(n22063), .A(n22064), .Z(n22062) );
XOR U36772 ( .A(c7354), .B(b[7354]), .Z(n22063) );
XNOR U36773 ( .A(b[7354]), .B(n22064), .Z(c[7354]) );
XNOR U36774 ( .A(a[7354]), .B(c7354), .Z(n22064) );
XOR U36775 ( .A(c7355), .B(n22065), .Z(c7356) );
ANDN U36776 ( .B(n22066), .A(n22067), .Z(n22065) );
XOR U36777 ( .A(c7355), .B(b[7355]), .Z(n22066) );
XNOR U36778 ( .A(b[7355]), .B(n22067), .Z(c[7355]) );
XNOR U36779 ( .A(a[7355]), .B(c7355), .Z(n22067) );
XOR U36780 ( .A(c7356), .B(n22068), .Z(c7357) );
ANDN U36781 ( .B(n22069), .A(n22070), .Z(n22068) );
XOR U36782 ( .A(c7356), .B(b[7356]), .Z(n22069) );
XNOR U36783 ( .A(b[7356]), .B(n22070), .Z(c[7356]) );
XNOR U36784 ( .A(a[7356]), .B(c7356), .Z(n22070) );
XOR U36785 ( .A(c7357), .B(n22071), .Z(c7358) );
ANDN U36786 ( .B(n22072), .A(n22073), .Z(n22071) );
XOR U36787 ( .A(c7357), .B(b[7357]), .Z(n22072) );
XNOR U36788 ( .A(b[7357]), .B(n22073), .Z(c[7357]) );
XNOR U36789 ( .A(a[7357]), .B(c7357), .Z(n22073) );
XOR U36790 ( .A(c7358), .B(n22074), .Z(c7359) );
ANDN U36791 ( .B(n22075), .A(n22076), .Z(n22074) );
XOR U36792 ( .A(c7358), .B(b[7358]), .Z(n22075) );
XNOR U36793 ( .A(b[7358]), .B(n22076), .Z(c[7358]) );
XNOR U36794 ( .A(a[7358]), .B(c7358), .Z(n22076) );
XOR U36795 ( .A(c7359), .B(n22077), .Z(c7360) );
ANDN U36796 ( .B(n22078), .A(n22079), .Z(n22077) );
XOR U36797 ( .A(c7359), .B(b[7359]), .Z(n22078) );
XNOR U36798 ( .A(b[7359]), .B(n22079), .Z(c[7359]) );
XNOR U36799 ( .A(a[7359]), .B(c7359), .Z(n22079) );
XOR U36800 ( .A(c7360), .B(n22080), .Z(c7361) );
ANDN U36801 ( .B(n22081), .A(n22082), .Z(n22080) );
XOR U36802 ( .A(c7360), .B(b[7360]), .Z(n22081) );
XNOR U36803 ( .A(b[7360]), .B(n22082), .Z(c[7360]) );
XNOR U36804 ( .A(a[7360]), .B(c7360), .Z(n22082) );
XOR U36805 ( .A(c7361), .B(n22083), .Z(c7362) );
ANDN U36806 ( .B(n22084), .A(n22085), .Z(n22083) );
XOR U36807 ( .A(c7361), .B(b[7361]), .Z(n22084) );
XNOR U36808 ( .A(b[7361]), .B(n22085), .Z(c[7361]) );
XNOR U36809 ( .A(a[7361]), .B(c7361), .Z(n22085) );
XOR U36810 ( .A(c7362), .B(n22086), .Z(c7363) );
ANDN U36811 ( .B(n22087), .A(n22088), .Z(n22086) );
XOR U36812 ( .A(c7362), .B(b[7362]), .Z(n22087) );
XNOR U36813 ( .A(b[7362]), .B(n22088), .Z(c[7362]) );
XNOR U36814 ( .A(a[7362]), .B(c7362), .Z(n22088) );
XOR U36815 ( .A(c7363), .B(n22089), .Z(c7364) );
ANDN U36816 ( .B(n22090), .A(n22091), .Z(n22089) );
XOR U36817 ( .A(c7363), .B(b[7363]), .Z(n22090) );
XNOR U36818 ( .A(b[7363]), .B(n22091), .Z(c[7363]) );
XNOR U36819 ( .A(a[7363]), .B(c7363), .Z(n22091) );
XOR U36820 ( .A(c7364), .B(n22092), .Z(c7365) );
ANDN U36821 ( .B(n22093), .A(n22094), .Z(n22092) );
XOR U36822 ( .A(c7364), .B(b[7364]), .Z(n22093) );
XNOR U36823 ( .A(b[7364]), .B(n22094), .Z(c[7364]) );
XNOR U36824 ( .A(a[7364]), .B(c7364), .Z(n22094) );
XOR U36825 ( .A(c7365), .B(n22095), .Z(c7366) );
ANDN U36826 ( .B(n22096), .A(n22097), .Z(n22095) );
XOR U36827 ( .A(c7365), .B(b[7365]), .Z(n22096) );
XNOR U36828 ( .A(b[7365]), .B(n22097), .Z(c[7365]) );
XNOR U36829 ( .A(a[7365]), .B(c7365), .Z(n22097) );
XOR U36830 ( .A(c7366), .B(n22098), .Z(c7367) );
ANDN U36831 ( .B(n22099), .A(n22100), .Z(n22098) );
XOR U36832 ( .A(c7366), .B(b[7366]), .Z(n22099) );
XNOR U36833 ( .A(b[7366]), .B(n22100), .Z(c[7366]) );
XNOR U36834 ( .A(a[7366]), .B(c7366), .Z(n22100) );
XOR U36835 ( .A(c7367), .B(n22101), .Z(c7368) );
ANDN U36836 ( .B(n22102), .A(n22103), .Z(n22101) );
XOR U36837 ( .A(c7367), .B(b[7367]), .Z(n22102) );
XNOR U36838 ( .A(b[7367]), .B(n22103), .Z(c[7367]) );
XNOR U36839 ( .A(a[7367]), .B(c7367), .Z(n22103) );
XOR U36840 ( .A(c7368), .B(n22104), .Z(c7369) );
ANDN U36841 ( .B(n22105), .A(n22106), .Z(n22104) );
XOR U36842 ( .A(c7368), .B(b[7368]), .Z(n22105) );
XNOR U36843 ( .A(b[7368]), .B(n22106), .Z(c[7368]) );
XNOR U36844 ( .A(a[7368]), .B(c7368), .Z(n22106) );
XOR U36845 ( .A(c7369), .B(n22107), .Z(c7370) );
ANDN U36846 ( .B(n22108), .A(n22109), .Z(n22107) );
XOR U36847 ( .A(c7369), .B(b[7369]), .Z(n22108) );
XNOR U36848 ( .A(b[7369]), .B(n22109), .Z(c[7369]) );
XNOR U36849 ( .A(a[7369]), .B(c7369), .Z(n22109) );
XOR U36850 ( .A(c7370), .B(n22110), .Z(c7371) );
ANDN U36851 ( .B(n22111), .A(n22112), .Z(n22110) );
XOR U36852 ( .A(c7370), .B(b[7370]), .Z(n22111) );
XNOR U36853 ( .A(b[7370]), .B(n22112), .Z(c[7370]) );
XNOR U36854 ( .A(a[7370]), .B(c7370), .Z(n22112) );
XOR U36855 ( .A(c7371), .B(n22113), .Z(c7372) );
ANDN U36856 ( .B(n22114), .A(n22115), .Z(n22113) );
XOR U36857 ( .A(c7371), .B(b[7371]), .Z(n22114) );
XNOR U36858 ( .A(b[7371]), .B(n22115), .Z(c[7371]) );
XNOR U36859 ( .A(a[7371]), .B(c7371), .Z(n22115) );
XOR U36860 ( .A(c7372), .B(n22116), .Z(c7373) );
ANDN U36861 ( .B(n22117), .A(n22118), .Z(n22116) );
XOR U36862 ( .A(c7372), .B(b[7372]), .Z(n22117) );
XNOR U36863 ( .A(b[7372]), .B(n22118), .Z(c[7372]) );
XNOR U36864 ( .A(a[7372]), .B(c7372), .Z(n22118) );
XOR U36865 ( .A(c7373), .B(n22119), .Z(c7374) );
ANDN U36866 ( .B(n22120), .A(n22121), .Z(n22119) );
XOR U36867 ( .A(c7373), .B(b[7373]), .Z(n22120) );
XNOR U36868 ( .A(b[7373]), .B(n22121), .Z(c[7373]) );
XNOR U36869 ( .A(a[7373]), .B(c7373), .Z(n22121) );
XOR U36870 ( .A(c7374), .B(n22122), .Z(c7375) );
ANDN U36871 ( .B(n22123), .A(n22124), .Z(n22122) );
XOR U36872 ( .A(c7374), .B(b[7374]), .Z(n22123) );
XNOR U36873 ( .A(b[7374]), .B(n22124), .Z(c[7374]) );
XNOR U36874 ( .A(a[7374]), .B(c7374), .Z(n22124) );
XOR U36875 ( .A(c7375), .B(n22125), .Z(c7376) );
ANDN U36876 ( .B(n22126), .A(n22127), .Z(n22125) );
XOR U36877 ( .A(c7375), .B(b[7375]), .Z(n22126) );
XNOR U36878 ( .A(b[7375]), .B(n22127), .Z(c[7375]) );
XNOR U36879 ( .A(a[7375]), .B(c7375), .Z(n22127) );
XOR U36880 ( .A(c7376), .B(n22128), .Z(c7377) );
ANDN U36881 ( .B(n22129), .A(n22130), .Z(n22128) );
XOR U36882 ( .A(c7376), .B(b[7376]), .Z(n22129) );
XNOR U36883 ( .A(b[7376]), .B(n22130), .Z(c[7376]) );
XNOR U36884 ( .A(a[7376]), .B(c7376), .Z(n22130) );
XOR U36885 ( .A(c7377), .B(n22131), .Z(c7378) );
ANDN U36886 ( .B(n22132), .A(n22133), .Z(n22131) );
XOR U36887 ( .A(c7377), .B(b[7377]), .Z(n22132) );
XNOR U36888 ( .A(b[7377]), .B(n22133), .Z(c[7377]) );
XNOR U36889 ( .A(a[7377]), .B(c7377), .Z(n22133) );
XOR U36890 ( .A(c7378), .B(n22134), .Z(c7379) );
ANDN U36891 ( .B(n22135), .A(n22136), .Z(n22134) );
XOR U36892 ( .A(c7378), .B(b[7378]), .Z(n22135) );
XNOR U36893 ( .A(b[7378]), .B(n22136), .Z(c[7378]) );
XNOR U36894 ( .A(a[7378]), .B(c7378), .Z(n22136) );
XOR U36895 ( .A(c7379), .B(n22137), .Z(c7380) );
ANDN U36896 ( .B(n22138), .A(n22139), .Z(n22137) );
XOR U36897 ( .A(c7379), .B(b[7379]), .Z(n22138) );
XNOR U36898 ( .A(b[7379]), .B(n22139), .Z(c[7379]) );
XNOR U36899 ( .A(a[7379]), .B(c7379), .Z(n22139) );
XOR U36900 ( .A(c7380), .B(n22140), .Z(c7381) );
ANDN U36901 ( .B(n22141), .A(n22142), .Z(n22140) );
XOR U36902 ( .A(c7380), .B(b[7380]), .Z(n22141) );
XNOR U36903 ( .A(b[7380]), .B(n22142), .Z(c[7380]) );
XNOR U36904 ( .A(a[7380]), .B(c7380), .Z(n22142) );
XOR U36905 ( .A(c7381), .B(n22143), .Z(c7382) );
ANDN U36906 ( .B(n22144), .A(n22145), .Z(n22143) );
XOR U36907 ( .A(c7381), .B(b[7381]), .Z(n22144) );
XNOR U36908 ( .A(b[7381]), .B(n22145), .Z(c[7381]) );
XNOR U36909 ( .A(a[7381]), .B(c7381), .Z(n22145) );
XOR U36910 ( .A(c7382), .B(n22146), .Z(c7383) );
ANDN U36911 ( .B(n22147), .A(n22148), .Z(n22146) );
XOR U36912 ( .A(c7382), .B(b[7382]), .Z(n22147) );
XNOR U36913 ( .A(b[7382]), .B(n22148), .Z(c[7382]) );
XNOR U36914 ( .A(a[7382]), .B(c7382), .Z(n22148) );
XOR U36915 ( .A(c7383), .B(n22149), .Z(c7384) );
ANDN U36916 ( .B(n22150), .A(n22151), .Z(n22149) );
XOR U36917 ( .A(c7383), .B(b[7383]), .Z(n22150) );
XNOR U36918 ( .A(b[7383]), .B(n22151), .Z(c[7383]) );
XNOR U36919 ( .A(a[7383]), .B(c7383), .Z(n22151) );
XOR U36920 ( .A(c7384), .B(n22152), .Z(c7385) );
ANDN U36921 ( .B(n22153), .A(n22154), .Z(n22152) );
XOR U36922 ( .A(c7384), .B(b[7384]), .Z(n22153) );
XNOR U36923 ( .A(b[7384]), .B(n22154), .Z(c[7384]) );
XNOR U36924 ( .A(a[7384]), .B(c7384), .Z(n22154) );
XOR U36925 ( .A(c7385), .B(n22155), .Z(c7386) );
ANDN U36926 ( .B(n22156), .A(n22157), .Z(n22155) );
XOR U36927 ( .A(c7385), .B(b[7385]), .Z(n22156) );
XNOR U36928 ( .A(b[7385]), .B(n22157), .Z(c[7385]) );
XNOR U36929 ( .A(a[7385]), .B(c7385), .Z(n22157) );
XOR U36930 ( .A(c7386), .B(n22158), .Z(c7387) );
ANDN U36931 ( .B(n22159), .A(n22160), .Z(n22158) );
XOR U36932 ( .A(c7386), .B(b[7386]), .Z(n22159) );
XNOR U36933 ( .A(b[7386]), .B(n22160), .Z(c[7386]) );
XNOR U36934 ( .A(a[7386]), .B(c7386), .Z(n22160) );
XOR U36935 ( .A(c7387), .B(n22161), .Z(c7388) );
ANDN U36936 ( .B(n22162), .A(n22163), .Z(n22161) );
XOR U36937 ( .A(c7387), .B(b[7387]), .Z(n22162) );
XNOR U36938 ( .A(b[7387]), .B(n22163), .Z(c[7387]) );
XNOR U36939 ( .A(a[7387]), .B(c7387), .Z(n22163) );
XOR U36940 ( .A(c7388), .B(n22164), .Z(c7389) );
ANDN U36941 ( .B(n22165), .A(n22166), .Z(n22164) );
XOR U36942 ( .A(c7388), .B(b[7388]), .Z(n22165) );
XNOR U36943 ( .A(b[7388]), .B(n22166), .Z(c[7388]) );
XNOR U36944 ( .A(a[7388]), .B(c7388), .Z(n22166) );
XOR U36945 ( .A(c7389), .B(n22167), .Z(c7390) );
ANDN U36946 ( .B(n22168), .A(n22169), .Z(n22167) );
XOR U36947 ( .A(c7389), .B(b[7389]), .Z(n22168) );
XNOR U36948 ( .A(b[7389]), .B(n22169), .Z(c[7389]) );
XNOR U36949 ( .A(a[7389]), .B(c7389), .Z(n22169) );
XOR U36950 ( .A(c7390), .B(n22170), .Z(c7391) );
ANDN U36951 ( .B(n22171), .A(n22172), .Z(n22170) );
XOR U36952 ( .A(c7390), .B(b[7390]), .Z(n22171) );
XNOR U36953 ( .A(b[7390]), .B(n22172), .Z(c[7390]) );
XNOR U36954 ( .A(a[7390]), .B(c7390), .Z(n22172) );
XOR U36955 ( .A(c7391), .B(n22173), .Z(c7392) );
ANDN U36956 ( .B(n22174), .A(n22175), .Z(n22173) );
XOR U36957 ( .A(c7391), .B(b[7391]), .Z(n22174) );
XNOR U36958 ( .A(b[7391]), .B(n22175), .Z(c[7391]) );
XNOR U36959 ( .A(a[7391]), .B(c7391), .Z(n22175) );
XOR U36960 ( .A(c7392), .B(n22176), .Z(c7393) );
ANDN U36961 ( .B(n22177), .A(n22178), .Z(n22176) );
XOR U36962 ( .A(c7392), .B(b[7392]), .Z(n22177) );
XNOR U36963 ( .A(b[7392]), .B(n22178), .Z(c[7392]) );
XNOR U36964 ( .A(a[7392]), .B(c7392), .Z(n22178) );
XOR U36965 ( .A(c7393), .B(n22179), .Z(c7394) );
ANDN U36966 ( .B(n22180), .A(n22181), .Z(n22179) );
XOR U36967 ( .A(c7393), .B(b[7393]), .Z(n22180) );
XNOR U36968 ( .A(b[7393]), .B(n22181), .Z(c[7393]) );
XNOR U36969 ( .A(a[7393]), .B(c7393), .Z(n22181) );
XOR U36970 ( .A(c7394), .B(n22182), .Z(c7395) );
ANDN U36971 ( .B(n22183), .A(n22184), .Z(n22182) );
XOR U36972 ( .A(c7394), .B(b[7394]), .Z(n22183) );
XNOR U36973 ( .A(b[7394]), .B(n22184), .Z(c[7394]) );
XNOR U36974 ( .A(a[7394]), .B(c7394), .Z(n22184) );
XOR U36975 ( .A(c7395), .B(n22185), .Z(c7396) );
ANDN U36976 ( .B(n22186), .A(n22187), .Z(n22185) );
XOR U36977 ( .A(c7395), .B(b[7395]), .Z(n22186) );
XNOR U36978 ( .A(b[7395]), .B(n22187), .Z(c[7395]) );
XNOR U36979 ( .A(a[7395]), .B(c7395), .Z(n22187) );
XOR U36980 ( .A(c7396), .B(n22188), .Z(c7397) );
ANDN U36981 ( .B(n22189), .A(n22190), .Z(n22188) );
XOR U36982 ( .A(c7396), .B(b[7396]), .Z(n22189) );
XNOR U36983 ( .A(b[7396]), .B(n22190), .Z(c[7396]) );
XNOR U36984 ( .A(a[7396]), .B(c7396), .Z(n22190) );
XOR U36985 ( .A(c7397), .B(n22191), .Z(c7398) );
ANDN U36986 ( .B(n22192), .A(n22193), .Z(n22191) );
XOR U36987 ( .A(c7397), .B(b[7397]), .Z(n22192) );
XNOR U36988 ( .A(b[7397]), .B(n22193), .Z(c[7397]) );
XNOR U36989 ( .A(a[7397]), .B(c7397), .Z(n22193) );
XOR U36990 ( .A(c7398), .B(n22194), .Z(c7399) );
ANDN U36991 ( .B(n22195), .A(n22196), .Z(n22194) );
XOR U36992 ( .A(c7398), .B(b[7398]), .Z(n22195) );
XNOR U36993 ( .A(b[7398]), .B(n22196), .Z(c[7398]) );
XNOR U36994 ( .A(a[7398]), .B(c7398), .Z(n22196) );
XOR U36995 ( .A(c7399), .B(n22197), .Z(c7400) );
ANDN U36996 ( .B(n22198), .A(n22199), .Z(n22197) );
XOR U36997 ( .A(c7399), .B(b[7399]), .Z(n22198) );
XNOR U36998 ( .A(b[7399]), .B(n22199), .Z(c[7399]) );
XNOR U36999 ( .A(a[7399]), .B(c7399), .Z(n22199) );
XOR U37000 ( .A(c7400), .B(n22200), .Z(c7401) );
ANDN U37001 ( .B(n22201), .A(n22202), .Z(n22200) );
XOR U37002 ( .A(c7400), .B(b[7400]), .Z(n22201) );
XNOR U37003 ( .A(b[7400]), .B(n22202), .Z(c[7400]) );
XNOR U37004 ( .A(a[7400]), .B(c7400), .Z(n22202) );
XOR U37005 ( .A(c7401), .B(n22203), .Z(c7402) );
ANDN U37006 ( .B(n22204), .A(n22205), .Z(n22203) );
XOR U37007 ( .A(c7401), .B(b[7401]), .Z(n22204) );
XNOR U37008 ( .A(b[7401]), .B(n22205), .Z(c[7401]) );
XNOR U37009 ( .A(a[7401]), .B(c7401), .Z(n22205) );
XOR U37010 ( .A(c7402), .B(n22206), .Z(c7403) );
ANDN U37011 ( .B(n22207), .A(n22208), .Z(n22206) );
XOR U37012 ( .A(c7402), .B(b[7402]), .Z(n22207) );
XNOR U37013 ( .A(b[7402]), .B(n22208), .Z(c[7402]) );
XNOR U37014 ( .A(a[7402]), .B(c7402), .Z(n22208) );
XOR U37015 ( .A(c7403), .B(n22209), .Z(c7404) );
ANDN U37016 ( .B(n22210), .A(n22211), .Z(n22209) );
XOR U37017 ( .A(c7403), .B(b[7403]), .Z(n22210) );
XNOR U37018 ( .A(b[7403]), .B(n22211), .Z(c[7403]) );
XNOR U37019 ( .A(a[7403]), .B(c7403), .Z(n22211) );
XOR U37020 ( .A(c7404), .B(n22212), .Z(c7405) );
ANDN U37021 ( .B(n22213), .A(n22214), .Z(n22212) );
XOR U37022 ( .A(c7404), .B(b[7404]), .Z(n22213) );
XNOR U37023 ( .A(b[7404]), .B(n22214), .Z(c[7404]) );
XNOR U37024 ( .A(a[7404]), .B(c7404), .Z(n22214) );
XOR U37025 ( .A(c7405), .B(n22215), .Z(c7406) );
ANDN U37026 ( .B(n22216), .A(n22217), .Z(n22215) );
XOR U37027 ( .A(c7405), .B(b[7405]), .Z(n22216) );
XNOR U37028 ( .A(b[7405]), .B(n22217), .Z(c[7405]) );
XNOR U37029 ( .A(a[7405]), .B(c7405), .Z(n22217) );
XOR U37030 ( .A(c7406), .B(n22218), .Z(c7407) );
ANDN U37031 ( .B(n22219), .A(n22220), .Z(n22218) );
XOR U37032 ( .A(c7406), .B(b[7406]), .Z(n22219) );
XNOR U37033 ( .A(b[7406]), .B(n22220), .Z(c[7406]) );
XNOR U37034 ( .A(a[7406]), .B(c7406), .Z(n22220) );
XOR U37035 ( .A(c7407), .B(n22221), .Z(c7408) );
ANDN U37036 ( .B(n22222), .A(n22223), .Z(n22221) );
XOR U37037 ( .A(c7407), .B(b[7407]), .Z(n22222) );
XNOR U37038 ( .A(b[7407]), .B(n22223), .Z(c[7407]) );
XNOR U37039 ( .A(a[7407]), .B(c7407), .Z(n22223) );
XOR U37040 ( .A(c7408), .B(n22224), .Z(c7409) );
ANDN U37041 ( .B(n22225), .A(n22226), .Z(n22224) );
XOR U37042 ( .A(c7408), .B(b[7408]), .Z(n22225) );
XNOR U37043 ( .A(b[7408]), .B(n22226), .Z(c[7408]) );
XNOR U37044 ( .A(a[7408]), .B(c7408), .Z(n22226) );
XOR U37045 ( .A(c7409), .B(n22227), .Z(c7410) );
ANDN U37046 ( .B(n22228), .A(n22229), .Z(n22227) );
XOR U37047 ( .A(c7409), .B(b[7409]), .Z(n22228) );
XNOR U37048 ( .A(b[7409]), .B(n22229), .Z(c[7409]) );
XNOR U37049 ( .A(a[7409]), .B(c7409), .Z(n22229) );
XOR U37050 ( .A(c7410), .B(n22230), .Z(c7411) );
ANDN U37051 ( .B(n22231), .A(n22232), .Z(n22230) );
XOR U37052 ( .A(c7410), .B(b[7410]), .Z(n22231) );
XNOR U37053 ( .A(b[7410]), .B(n22232), .Z(c[7410]) );
XNOR U37054 ( .A(a[7410]), .B(c7410), .Z(n22232) );
XOR U37055 ( .A(c7411), .B(n22233), .Z(c7412) );
ANDN U37056 ( .B(n22234), .A(n22235), .Z(n22233) );
XOR U37057 ( .A(c7411), .B(b[7411]), .Z(n22234) );
XNOR U37058 ( .A(b[7411]), .B(n22235), .Z(c[7411]) );
XNOR U37059 ( .A(a[7411]), .B(c7411), .Z(n22235) );
XOR U37060 ( .A(c7412), .B(n22236), .Z(c7413) );
ANDN U37061 ( .B(n22237), .A(n22238), .Z(n22236) );
XOR U37062 ( .A(c7412), .B(b[7412]), .Z(n22237) );
XNOR U37063 ( .A(b[7412]), .B(n22238), .Z(c[7412]) );
XNOR U37064 ( .A(a[7412]), .B(c7412), .Z(n22238) );
XOR U37065 ( .A(c7413), .B(n22239), .Z(c7414) );
ANDN U37066 ( .B(n22240), .A(n22241), .Z(n22239) );
XOR U37067 ( .A(c7413), .B(b[7413]), .Z(n22240) );
XNOR U37068 ( .A(b[7413]), .B(n22241), .Z(c[7413]) );
XNOR U37069 ( .A(a[7413]), .B(c7413), .Z(n22241) );
XOR U37070 ( .A(c7414), .B(n22242), .Z(c7415) );
ANDN U37071 ( .B(n22243), .A(n22244), .Z(n22242) );
XOR U37072 ( .A(c7414), .B(b[7414]), .Z(n22243) );
XNOR U37073 ( .A(b[7414]), .B(n22244), .Z(c[7414]) );
XNOR U37074 ( .A(a[7414]), .B(c7414), .Z(n22244) );
XOR U37075 ( .A(c7415), .B(n22245), .Z(c7416) );
ANDN U37076 ( .B(n22246), .A(n22247), .Z(n22245) );
XOR U37077 ( .A(c7415), .B(b[7415]), .Z(n22246) );
XNOR U37078 ( .A(b[7415]), .B(n22247), .Z(c[7415]) );
XNOR U37079 ( .A(a[7415]), .B(c7415), .Z(n22247) );
XOR U37080 ( .A(c7416), .B(n22248), .Z(c7417) );
ANDN U37081 ( .B(n22249), .A(n22250), .Z(n22248) );
XOR U37082 ( .A(c7416), .B(b[7416]), .Z(n22249) );
XNOR U37083 ( .A(b[7416]), .B(n22250), .Z(c[7416]) );
XNOR U37084 ( .A(a[7416]), .B(c7416), .Z(n22250) );
XOR U37085 ( .A(c7417), .B(n22251), .Z(c7418) );
ANDN U37086 ( .B(n22252), .A(n22253), .Z(n22251) );
XOR U37087 ( .A(c7417), .B(b[7417]), .Z(n22252) );
XNOR U37088 ( .A(b[7417]), .B(n22253), .Z(c[7417]) );
XNOR U37089 ( .A(a[7417]), .B(c7417), .Z(n22253) );
XOR U37090 ( .A(c7418), .B(n22254), .Z(c7419) );
ANDN U37091 ( .B(n22255), .A(n22256), .Z(n22254) );
XOR U37092 ( .A(c7418), .B(b[7418]), .Z(n22255) );
XNOR U37093 ( .A(b[7418]), .B(n22256), .Z(c[7418]) );
XNOR U37094 ( .A(a[7418]), .B(c7418), .Z(n22256) );
XOR U37095 ( .A(c7419), .B(n22257), .Z(c7420) );
ANDN U37096 ( .B(n22258), .A(n22259), .Z(n22257) );
XOR U37097 ( .A(c7419), .B(b[7419]), .Z(n22258) );
XNOR U37098 ( .A(b[7419]), .B(n22259), .Z(c[7419]) );
XNOR U37099 ( .A(a[7419]), .B(c7419), .Z(n22259) );
XOR U37100 ( .A(c7420), .B(n22260), .Z(c7421) );
ANDN U37101 ( .B(n22261), .A(n22262), .Z(n22260) );
XOR U37102 ( .A(c7420), .B(b[7420]), .Z(n22261) );
XNOR U37103 ( .A(b[7420]), .B(n22262), .Z(c[7420]) );
XNOR U37104 ( .A(a[7420]), .B(c7420), .Z(n22262) );
XOR U37105 ( .A(c7421), .B(n22263), .Z(c7422) );
ANDN U37106 ( .B(n22264), .A(n22265), .Z(n22263) );
XOR U37107 ( .A(c7421), .B(b[7421]), .Z(n22264) );
XNOR U37108 ( .A(b[7421]), .B(n22265), .Z(c[7421]) );
XNOR U37109 ( .A(a[7421]), .B(c7421), .Z(n22265) );
XOR U37110 ( .A(c7422), .B(n22266), .Z(c7423) );
ANDN U37111 ( .B(n22267), .A(n22268), .Z(n22266) );
XOR U37112 ( .A(c7422), .B(b[7422]), .Z(n22267) );
XNOR U37113 ( .A(b[7422]), .B(n22268), .Z(c[7422]) );
XNOR U37114 ( .A(a[7422]), .B(c7422), .Z(n22268) );
XOR U37115 ( .A(c7423), .B(n22269), .Z(c7424) );
ANDN U37116 ( .B(n22270), .A(n22271), .Z(n22269) );
XOR U37117 ( .A(c7423), .B(b[7423]), .Z(n22270) );
XNOR U37118 ( .A(b[7423]), .B(n22271), .Z(c[7423]) );
XNOR U37119 ( .A(a[7423]), .B(c7423), .Z(n22271) );
XOR U37120 ( .A(c7424), .B(n22272), .Z(c7425) );
ANDN U37121 ( .B(n22273), .A(n22274), .Z(n22272) );
XOR U37122 ( .A(c7424), .B(b[7424]), .Z(n22273) );
XNOR U37123 ( .A(b[7424]), .B(n22274), .Z(c[7424]) );
XNOR U37124 ( .A(a[7424]), .B(c7424), .Z(n22274) );
XOR U37125 ( .A(c7425), .B(n22275), .Z(c7426) );
ANDN U37126 ( .B(n22276), .A(n22277), .Z(n22275) );
XOR U37127 ( .A(c7425), .B(b[7425]), .Z(n22276) );
XNOR U37128 ( .A(b[7425]), .B(n22277), .Z(c[7425]) );
XNOR U37129 ( .A(a[7425]), .B(c7425), .Z(n22277) );
XOR U37130 ( .A(c7426), .B(n22278), .Z(c7427) );
ANDN U37131 ( .B(n22279), .A(n22280), .Z(n22278) );
XOR U37132 ( .A(c7426), .B(b[7426]), .Z(n22279) );
XNOR U37133 ( .A(b[7426]), .B(n22280), .Z(c[7426]) );
XNOR U37134 ( .A(a[7426]), .B(c7426), .Z(n22280) );
XOR U37135 ( .A(c7427), .B(n22281), .Z(c7428) );
ANDN U37136 ( .B(n22282), .A(n22283), .Z(n22281) );
XOR U37137 ( .A(c7427), .B(b[7427]), .Z(n22282) );
XNOR U37138 ( .A(b[7427]), .B(n22283), .Z(c[7427]) );
XNOR U37139 ( .A(a[7427]), .B(c7427), .Z(n22283) );
XOR U37140 ( .A(c7428), .B(n22284), .Z(c7429) );
ANDN U37141 ( .B(n22285), .A(n22286), .Z(n22284) );
XOR U37142 ( .A(c7428), .B(b[7428]), .Z(n22285) );
XNOR U37143 ( .A(b[7428]), .B(n22286), .Z(c[7428]) );
XNOR U37144 ( .A(a[7428]), .B(c7428), .Z(n22286) );
XOR U37145 ( .A(c7429), .B(n22287), .Z(c7430) );
ANDN U37146 ( .B(n22288), .A(n22289), .Z(n22287) );
XOR U37147 ( .A(c7429), .B(b[7429]), .Z(n22288) );
XNOR U37148 ( .A(b[7429]), .B(n22289), .Z(c[7429]) );
XNOR U37149 ( .A(a[7429]), .B(c7429), .Z(n22289) );
XOR U37150 ( .A(c7430), .B(n22290), .Z(c7431) );
ANDN U37151 ( .B(n22291), .A(n22292), .Z(n22290) );
XOR U37152 ( .A(c7430), .B(b[7430]), .Z(n22291) );
XNOR U37153 ( .A(b[7430]), .B(n22292), .Z(c[7430]) );
XNOR U37154 ( .A(a[7430]), .B(c7430), .Z(n22292) );
XOR U37155 ( .A(c7431), .B(n22293), .Z(c7432) );
ANDN U37156 ( .B(n22294), .A(n22295), .Z(n22293) );
XOR U37157 ( .A(c7431), .B(b[7431]), .Z(n22294) );
XNOR U37158 ( .A(b[7431]), .B(n22295), .Z(c[7431]) );
XNOR U37159 ( .A(a[7431]), .B(c7431), .Z(n22295) );
XOR U37160 ( .A(c7432), .B(n22296), .Z(c7433) );
ANDN U37161 ( .B(n22297), .A(n22298), .Z(n22296) );
XOR U37162 ( .A(c7432), .B(b[7432]), .Z(n22297) );
XNOR U37163 ( .A(b[7432]), .B(n22298), .Z(c[7432]) );
XNOR U37164 ( .A(a[7432]), .B(c7432), .Z(n22298) );
XOR U37165 ( .A(c7433), .B(n22299), .Z(c7434) );
ANDN U37166 ( .B(n22300), .A(n22301), .Z(n22299) );
XOR U37167 ( .A(c7433), .B(b[7433]), .Z(n22300) );
XNOR U37168 ( .A(b[7433]), .B(n22301), .Z(c[7433]) );
XNOR U37169 ( .A(a[7433]), .B(c7433), .Z(n22301) );
XOR U37170 ( .A(c7434), .B(n22302), .Z(c7435) );
ANDN U37171 ( .B(n22303), .A(n22304), .Z(n22302) );
XOR U37172 ( .A(c7434), .B(b[7434]), .Z(n22303) );
XNOR U37173 ( .A(b[7434]), .B(n22304), .Z(c[7434]) );
XNOR U37174 ( .A(a[7434]), .B(c7434), .Z(n22304) );
XOR U37175 ( .A(c7435), .B(n22305), .Z(c7436) );
ANDN U37176 ( .B(n22306), .A(n22307), .Z(n22305) );
XOR U37177 ( .A(c7435), .B(b[7435]), .Z(n22306) );
XNOR U37178 ( .A(b[7435]), .B(n22307), .Z(c[7435]) );
XNOR U37179 ( .A(a[7435]), .B(c7435), .Z(n22307) );
XOR U37180 ( .A(c7436), .B(n22308), .Z(c7437) );
ANDN U37181 ( .B(n22309), .A(n22310), .Z(n22308) );
XOR U37182 ( .A(c7436), .B(b[7436]), .Z(n22309) );
XNOR U37183 ( .A(b[7436]), .B(n22310), .Z(c[7436]) );
XNOR U37184 ( .A(a[7436]), .B(c7436), .Z(n22310) );
XOR U37185 ( .A(c7437), .B(n22311), .Z(c7438) );
ANDN U37186 ( .B(n22312), .A(n22313), .Z(n22311) );
XOR U37187 ( .A(c7437), .B(b[7437]), .Z(n22312) );
XNOR U37188 ( .A(b[7437]), .B(n22313), .Z(c[7437]) );
XNOR U37189 ( .A(a[7437]), .B(c7437), .Z(n22313) );
XOR U37190 ( .A(c7438), .B(n22314), .Z(c7439) );
ANDN U37191 ( .B(n22315), .A(n22316), .Z(n22314) );
XOR U37192 ( .A(c7438), .B(b[7438]), .Z(n22315) );
XNOR U37193 ( .A(b[7438]), .B(n22316), .Z(c[7438]) );
XNOR U37194 ( .A(a[7438]), .B(c7438), .Z(n22316) );
XOR U37195 ( .A(c7439), .B(n22317), .Z(c7440) );
ANDN U37196 ( .B(n22318), .A(n22319), .Z(n22317) );
XOR U37197 ( .A(c7439), .B(b[7439]), .Z(n22318) );
XNOR U37198 ( .A(b[7439]), .B(n22319), .Z(c[7439]) );
XNOR U37199 ( .A(a[7439]), .B(c7439), .Z(n22319) );
XOR U37200 ( .A(c7440), .B(n22320), .Z(c7441) );
ANDN U37201 ( .B(n22321), .A(n22322), .Z(n22320) );
XOR U37202 ( .A(c7440), .B(b[7440]), .Z(n22321) );
XNOR U37203 ( .A(b[7440]), .B(n22322), .Z(c[7440]) );
XNOR U37204 ( .A(a[7440]), .B(c7440), .Z(n22322) );
XOR U37205 ( .A(c7441), .B(n22323), .Z(c7442) );
ANDN U37206 ( .B(n22324), .A(n22325), .Z(n22323) );
XOR U37207 ( .A(c7441), .B(b[7441]), .Z(n22324) );
XNOR U37208 ( .A(b[7441]), .B(n22325), .Z(c[7441]) );
XNOR U37209 ( .A(a[7441]), .B(c7441), .Z(n22325) );
XOR U37210 ( .A(c7442), .B(n22326), .Z(c7443) );
ANDN U37211 ( .B(n22327), .A(n22328), .Z(n22326) );
XOR U37212 ( .A(c7442), .B(b[7442]), .Z(n22327) );
XNOR U37213 ( .A(b[7442]), .B(n22328), .Z(c[7442]) );
XNOR U37214 ( .A(a[7442]), .B(c7442), .Z(n22328) );
XOR U37215 ( .A(c7443), .B(n22329), .Z(c7444) );
ANDN U37216 ( .B(n22330), .A(n22331), .Z(n22329) );
XOR U37217 ( .A(c7443), .B(b[7443]), .Z(n22330) );
XNOR U37218 ( .A(b[7443]), .B(n22331), .Z(c[7443]) );
XNOR U37219 ( .A(a[7443]), .B(c7443), .Z(n22331) );
XOR U37220 ( .A(c7444), .B(n22332), .Z(c7445) );
ANDN U37221 ( .B(n22333), .A(n22334), .Z(n22332) );
XOR U37222 ( .A(c7444), .B(b[7444]), .Z(n22333) );
XNOR U37223 ( .A(b[7444]), .B(n22334), .Z(c[7444]) );
XNOR U37224 ( .A(a[7444]), .B(c7444), .Z(n22334) );
XOR U37225 ( .A(c7445), .B(n22335), .Z(c7446) );
ANDN U37226 ( .B(n22336), .A(n22337), .Z(n22335) );
XOR U37227 ( .A(c7445), .B(b[7445]), .Z(n22336) );
XNOR U37228 ( .A(b[7445]), .B(n22337), .Z(c[7445]) );
XNOR U37229 ( .A(a[7445]), .B(c7445), .Z(n22337) );
XOR U37230 ( .A(c7446), .B(n22338), .Z(c7447) );
ANDN U37231 ( .B(n22339), .A(n22340), .Z(n22338) );
XOR U37232 ( .A(c7446), .B(b[7446]), .Z(n22339) );
XNOR U37233 ( .A(b[7446]), .B(n22340), .Z(c[7446]) );
XNOR U37234 ( .A(a[7446]), .B(c7446), .Z(n22340) );
XOR U37235 ( .A(c7447), .B(n22341), .Z(c7448) );
ANDN U37236 ( .B(n22342), .A(n22343), .Z(n22341) );
XOR U37237 ( .A(c7447), .B(b[7447]), .Z(n22342) );
XNOR U37238 ( .A(b[7447]), .B(n22343), .Z(c[7447]) );
XNOR U37239 ( .A(a[7447]), .B(c7447), .Z(n22343) );
XOR U37240 ( .A(c7448), .B(n22344), .Z(c7449) );
ANDN U37241 ( .B(n22345), .A(n22346), .Z(n22344) );
XOR U37242 ( .A(c7448), .B(b[7448]), .Z(n22345) );
XNOR U37243 ( .A(b[7448]), .B(n22346), .Z(c[7448]) );
XNOR U37244 ( .A(a[7448]), .B(c7448), .Z(n22346) );
XOR U37245 ( .A(c7449), .B(n22347), .Z(c7450) );
ANDN U37246 ( .B(n22348), .A(n22349), .Z(n22347) );
XOR U37247 ( .A(c7449), .B(b[7449]), .Z(n22348) );
XNOR U37248 ( .A(b[7449]), .B(n22349), .Z(c[7449]) );
XNOR U37249 ( .A(a[7449]), .B(c7449), .Z(n22349) );
XOR U37250 ( .A(c7450), .B(n22350), .Z(c7451) );
ANDN U37251 ( .B(n22351), .A(n22352), .Z(n22350) );
XOR U37252 ( .A(c7450), .B(b[7450]), .Z(n22351) );
XNOR U37253 ( .A(b[7450]), .B(n22352), .Z(c[7450]) );
XNOR U37254 ( .A(a[7450]), .B(c7450), .Z(n22352) );
XOR U37255 ( .A(c7451), .B(n22353), .Z(c7452) );
ANDN U37256 ( .B(n22354), .A(n22355), .Z(n22353) );
XOR U37257 ( .A(c7451), .B(b[7451]), .Z(n22354) );
XNOR U37258 ( .A(b[7451]), .B(n22355), .Z(c[7451]) );
XNOR U37259 ( .A(a[7451]), .B(c7451), .Z(n22355) );
XOR U37260 ( .A(c7452), .B(n22356), .Z(c7453) );
ANDN U37261 ( .B(n22357), .A(n22358), .Z(n22356) );
XOR U37262 ( .A(c7452), .B(b[7452]), .Z(n22357) );
XNOR U37263 ( .A(b[7452]), .B(n22358), .Z(c[7452]) );
XNOR U37264 ( .A(a[7452]), .B(c7452), .Z(n22358) );
XOR U37265 ( .A(c7453), .B(n22359), .Z(c7454) );
ANDN U37266 ( .B(n22360), .A(n22361), .Z(n22359) );
XOR U37267 ( .A(c7453), .B(b[7453]), .Z(n22360) );
XNOR U37268 ( .A(b[7453]), .B(n22361), .Z(c[7453]) );
XNOR U37269 ( .A(a[7453]), .B(c7453), .Z(n22361) );
XOR U37270 ( .A(c7454), .B(n22362), .Z(c7455) );
ANDN U37271 ( .B(n22363), .A(n22364), .Z(n22362) );
XOR U37272 ( .A(c7454), .B(b[7454]), .Z(n22363) );
XNOR U37273 ( .A(b[7454]), .B(n22364), .Z(c[7454]) );
XNOR U37274 ( .A(a[7454]), .B(c7454), .Z(n22364) );
XOR U37275 ( .A(c7455), .B(n22365), .Z(c7456) );
ANDN U37276 ( .B(n22366), .A(n22367), .Z(n22365) );
XOR U37277 ( .A(c7455), .B(b[7455]), .Z(n22366) );
XNOR U37278 ( .A(b[7455]), .B(n22367), .Z(c[7455]) );
XNOR U37279 ( .A(a[7455]), .B(c7455), .Z(n22367) );
XOR U37280 ( .A(c7456), .B(n22368), .Z(c7457) );
ANDN U37281 ( .B(n22369), .A(n22370), .Z(n22368) );
XOR U37282 ( .A(c7456), .B(b[7456]), .Z(n22369) );
XNOR U37283 ( .A(b[7456]), .B(n22370), .Z(c[7456]) );
XNOR U37284 ( .A(a[7456]), .B(c7456), .Z(n22370) );
XOR U37285 ( .A(c7457), .B(n22371), .Z(c7458) );
ANDN U37286 ( .B(n22372), .A(n22373), .Z(n22371) );
XOR U37287 ( .A(c7457), .B(b[7457]), .Z(n22372) );
XNOR U37288 ( .A(b[7457]), .B(n22373), .Z(c[7457]) );
XNOR U37289 ( .A(a[7457]), .B(c7457), .Z(n22373) );
XOR U37290 ( .A(c7458), .B(n22374), .Z(c7459) );
ANDN U37291 ( .B(n22375), .A(n22376), .Z(n22374) );
XOR U37292 ( .A(c7458), .B(b[7458]), .Z(n22375) );
XNOR U37293 ( .A(b[7458]), .B(n22376), .Z(c[7458]) );
XNOR U37294 ( .A(a[7458]), .B(c7458), .Z(n22376) );
XOR U37295 ( .A(c7459), .B(n22377), .Z(c7460) );
ANDN U37296 ( .B(n22378), .A(n22379), .Z(n22377) );
XOR U37297 ( .A(c7459), .B(b[7459]), .Z(n22378) );
XNOR U37298 ( .A(b[7459]), .B(n22379), .Z(c[7459]) );
XNOR U37299 ( .A(a[7459]), .B(c7459), .Z(n22379) );
XOR U37300 ( .A(c7460), .B(n22380), .Z(c7461) );
ANDN U37301 ( .B(n22381), .A(n22382), .Z(n22380) );
XOR U37302 ( .A(c7460), .B(b[7460]), .Z(n22381) );
XNOR U37303 ( .A(b[7460]), .B(n22382), .Z(c[7460]) );
XNOR U37304 ( .A(a[7460]), .B(c7460), .Z(n22382) );
XOR U37305 ( .A(c7461), .B(n22383), .Z(c7462) );
ANDN U37306 ( .B(n22384), .A(n22385), .Z(n22383) );
XOR U37307 ( .A(c7461), .B(b[7461]), .Z(n22384) );
XNOR U37308 ( .A(b[7461]), .B(n22385), .Z(c[7461]) );
XNOR U37309 ( .A(a[7461]), .B(c7461), .Z(n22385) );
XOR U37310 ( .A(c7462), .B(n22386), .Z(c7463) );
ANDN U37311 ( .B(n22387), .A(n22388), .Z(n22386) );
XOR U37312 ( .A(c7462), .B(b[7462]), .Z(n22387) );
XNOR U37313 ( .A(b[7462]), .B(n22388), .Z(c[7462]) );
XNOR U37314 ( .A(a[7462]), .B(c7462), .Z(n22388) );
XOR U37315 ( .A(c7463), .B(n22389), .Z(c7464) );
ANDN U37316 ( .B(n22390), .A(n22391), .Z(n22389) );
XOR U37317 ( .A(c7463), .B(b[7463]), .Z(n22390) );
XNOR U37318 ( .A(b[7463]), .B(n22391), .Z(c[7463]) );
XNOR U37319 ( .A(a[7463]), .B(c7463), .Z(n22391) );
XOR U37320 ( .A(c7464), .B(n22392), .Z(c7465) );
ANDN U37321 ( .B(n22393), .A(n22394), .Z(n22392) );
XOR U37322 ( .A(c7464), .B(b[7464]), .Z(n22393) );
XNOR U37323 ( .A(b[7464]), .B(n22394), .Z(c[7464]) );
XNOR U37324 ( .A(a[7464]), .B(c7464), .Z(n22394) );
XOR U37325 ( .A(c7465), .B(n22395), .Z(c7466) );
ANDN U37326 ( .B(n22396), .A(n22397), .Z(n22395) );
XOR U37327 ( .A(c7465), .B(b[7465]), .Z(n22396) );
XNOR U37328 ( .A(b[7465]), .B(n22397), .Z(c[7465]) );
XNOR U37329 ( .A(a[7465]), .B(c7465), .Z(n22397) );
XOR U37330 ( .A(c7466), .B(n22398), .Z(c7467) );
ANDN U37331 ( .B(n22399), .A(n22400), .Z(n22398) );
XOR U37332 ( .A(c7466), .B(b[7466]), .Z(n22399) );
XNOR U37333 ( .A(b[7466]), .B(n22400), .Z(c[7466]) );
XNOR U37334 ( .A(a[7466]), .B(c7466), .Z(n22400) );
XOR U37335 ( .A(c7467), .B(n22401), .Z(c7468) );
ANDN U37336 ( .B(n22402), .A(n22403), .Z(n22401) );
XOR U37337 ( .A(c7467), .B(b[7467]), .Z(n22402) );
XNOR U37338 ( .A(b[7467]), .B(n22403), .Z(c[7467]) );
XNOR U37339 ( .A(a[7467]), .B(c7467), .Z(n22403) );
XOR U37340 ( .A(c7468), .B(n22404), .Z(c7469) );
ANDN U37341 ( .B(n22405), .A(n22406), .Z(n22404) );
XOR U37342 ( .A(c7468), .B(b[7468]), .Z(n22405) );
XNOR U37343 ( .A(b[7468]), .B(n22406), .Z(c[7468]) );
XNOR U37344 ( .A(a[7468]), .B(c7468), .Z(n22406) );
XOR U37345 ( .A(c7469), .B(n22407), .Z(c7470) );
ANDN U37346 ( .B(n22408), .A(n22409), .Z(n22407) );
XOR U37347 ( .A(c7469), .B(b[7469]), .Z(n22408) );
XNOR U37348 ( .A(b[7469]), .B(n22409), .Z(c[7469]) );
XNOR U37349 ( .A(a[7469]), .B(c7469), .Z(n22409) );
XOR U37350 ( .A(c7470), .B(n22410), .Z(c7471) );
ANDN U37351 ( .B(n22411), .A(n22412), .Z(n22410) );
XOR U37352 ( .A(c7470), .B(b[7470]), .Z(n22411) );
XNOR U37353 ( .A(b[7470]), .B(n22412), .Z(c[7470]) );
XNOR U37354 ( .A(a[7470]), .B(c7470), .Z(n22412) );
XOR U37355 ( .A(c7471), .B(n22413), .Z(c7472) );
ANDN U37356 ( .B(n22414), .A(n22415), .Z(n22413) );
XOR U37357 ( .A(c7471), .B(b[7471]), .Z(n22414) );
XNOR U37358 ( .A(b[7471]), .B(n22415), .Z(c[7471]) );
XNOR U37359 ( .A(a[7471]), .B(c7471), .Z(n22415) );
XOR U37360 ( .A(c7472), .B(n22416), .Z(c7473) );
ANDN U37361 ( .B(n22417), .A(n22418), .Z(n22416) );
XOR U37362 ( .A(c7472), .B(b[7472]), .Z(n22417) );
XNOR U37363 ( .A(b[7472]), .B(n22418), .Z(c[7472]) );
XNOR U37364 ( .A(a[7472]), .B(c7472), .Z(n22418) );
XOR U37365 ( .A(c7473), .B(n22419), .Z(c7474) );
ANDN U37366 ( .B(n22420), .A(n22421), .Z(n22419) );
XOR U37367 ( .A(c7473), .B(b[7473]), .Z(n22420) );
XNOR U37368 ( .A(b[7473]), .B(n22421), .Z(c[7473]) );
XNOR U37369 ( .A(a[7473]), .B(c7473), .Z(n22421) );
XOR U37370 ( .A(c7474), .B(n22422), .Z(c7475) );
ANDN U37371 ( .B(n22423), .A(n22424), .Z(n22422) );
XOR U37372 ( .A(c7474), .B(b[7474]), .Z(n22423) );
XNOR U37373 ( .A(b[7474]), .B(n22424), .Z(c[7474]) );
XNOR U37374 ( .A(a[7474]), .B(c7474), .Z(n22424) );
XOR U37375 ( .A(c7475), .B(n22425), .Z(c7476) );
ANDN U37376 ( .B(n22426), .A(n22427), .Z(n22425) );
XOR U37377 ( .A(c7475), .B(b[7475]), .Z(n22426) );
XNOR U37378 ( .A(b[7475]), .B(n22427), .Z(c[7475]) );
XNOR U37379 ( .A(a[7475]), .B(c7475), .Z(n22427) );
XOR U37380 ( .A(c7476), .B(n22428), .Z(c7477) );
ANDN U37381 ( .B(n22429), .A(n22430), .Z(n22428) );
XOR U37382 ( .A(c7476), .B(b[7476]), .Z(n22429) );
XNOR U37383 ( .A(b[7476]), .B(n22430), .Z(c[7476]) );
XNOR U37384 ( .A(a[7476]), .B(c7476), .Z(n22430) );
XOR U37385 ( .A(c7477), .B(n22431), .Z(c7478) );
ANDN U37386 ( .B(n22432), .A(n22433), .Z(n22431) );
XOR U37387 ( .A(c7477), .B(b[7477]), .Z(n22432) );
XNOR U37388 ( .A(b[7477]), .B(n22433), .Z(c[7477]) );
XNOR U37389 ( .A(a[7477]), .B(c7477), .Z(n22433) );
XOR U37390 ( .A(c7478), .B(n22434), .Z(c7479) );
ANDN U37391 ( .B(n22435), .A(n22436), .Z(n22434) );
XOR U37392 ( .A(c7478), .B(b[7478]), .Z(n22435) );
XNOR U37393 ( .A(b[7478]), .B(n22436), .Z(c[7478]) );
XNOR U37394 ( .A(a[7478]), .B(c7478), .Z(n22436) );
XOR U37395 ( .A(c7479), .B(n22437), .Z(c7480) );
ANDN U37396 ( .B(n22438), .A(n22439), .Z(n22437) );
XOR U37397 ( .A(c7479), .B(b[7479]), .Z(n22438) );
XNOR U37398 ( .A(b[7479]), .B(n22439), .Z(c[7479]) );
XNOR U37399 ( .A(a[7479]), .B(c7479), .Z(n22439) );
XOR U37400 ( .A(c7480), .B(n22440), .Z(c7481) );
ANDN U37401 ( .B(n22441), .A(n22442), .Z(n22440) );
XOR U37402 ( .A(c7480), .B(b[7480]), .Z(n22441) );
XNOR U37403 ( .A(b[7480]), .B(n22442), .Z(c[7480]) );
XNOR U37404 ( .A(a[7480]), .B(c7480), .Z(n22442) );
XOR U37405 ( .A(c7481), .B(n22443), .Z(c7482) );
ANDN U37406 ( .B(n22444), .A(n22445), .Z(n22443) );
XOR U37407 ( .A(c7481), .B(b[7481]), .Z(n22444) );
XNOR U37408 ( .A(b[7481]), .B(n22445), .Z(c[7481]) );
XNOR U37409 ( .A(a[7481]), .B(c7481), .Z(n22445) );
XOR U37410 ( .A(c7482), .B(n22446), .Z(c7483) );
ANDN U37411 ( .B(n22447), .A(n22448), .Z(n22446) );
XOR U37412 ( .A(c7482), .B(b[7482]), .Z(n22447) );
XNOR U37413 ( .A(b[7482]), .B(n22448), .Z(c[7482]) );
XNOR U37414 ( .A(a[7482]), .B(c7482), .Z(n22448) );
XOR U37415 ( .A(c7483), .B(n22449), .Z(c7484) );
ANDN U37416 ( .B(n22450), .A(n22451), .Z(n22449) );
XOR U37417 ( .A(c7483), .B(b[7483]), .Z(n22450) );
XNOR U37418 ( .A(b[7483]), .B(n22451), .Z(c[7483]) );
XNOR U37419 ( .A(a[7483]), .B(c7483), .Z(n22451) );
XOR U37420 ( .A(c7484), .B(n22452), .Z(c7485) );
ANDN U37421 ( .B(n22453), .A(n22454), .Z(n22452) );
XOR U37422 ( .A(c7484), .B(b[7484]), .Z(n22453) );
XNOR U37423 ( .A(b[7484]), .B(n22454), .Z(c[7484]) );
XNOR U37424 ( .A(a[7484]), .B(c7484), .Z(n22454) );
XOR U37425 ( .A(c7485), .B(n22455), .Z(c7486) );
ANDN U37426 ( .B(n22456), .A(n22457), .Z(n22455) );
XOR U37427 ( .A(c7485), .B(b[7485]), .Z(n22456) );
XNOR U37428 ( .A(b[7485]), .B(n22457), .Z(c[7485]) );
XNOR U37429 ( .A(a[7485]), .B(c7485), .Z(n22457) );
XOR U37430 ( .A(c7486), .B(n22458), .Z(c7487) );
ANDN U37431 ( .B(n22459), .A(n22460), .Z(n22458) );
XOR U37432 ( .A(c7486), .B(b[7486]), .Z(n22459) );
XNOR U37433 ( .A(b[7486]), .B(n22460), .Z(c[7486]) );
XNOR U37434 ( .A(a[7486]), .B(c7486), .Z(n22460) );
XOR U37435 ( .A(c7487), .B(n22461), .Z(c7488) );
ANDN U37436 ( .B(n22462), .A(n22463), .Z(n22461) );
XOR U37437 ( .A(c7487), .B(b[7487]), .Z(n22462) );
XNOR U37438 ( .A(b[7487]), .B(n22463), .Z(c[7487]) );
XNOR U37439 ( .A(a[7487]), .B(c7487), .Z(n22463) );
XOR U37440 ( .A(c7488), .B(n22464), .Z(c7489) );
ANDN U37441 ( .B(n22465), .A(n22466), .Z(n22464) );
XOR U37442 ( .A(c7488), .B(b[7488]), .Z(n22465) );
XNOR U37443 ( .A(b[7488]), .B(n22466), .Z(c[7488]) );
XNOR U37444 ( .A(a[7488]), .B(c7488), .Z(n22466) );
XOR U37445 ( .A(c7489), .B(n22467), .Z(c7490) );
ANDN U37446 ( .B(n22468), .A(n22469), .Z(n22467) );
XOR U37447 ( .A(c7489), .B(b[7489]), .Z(n22468) );
XNOR U37448 ( .A(b[7489]), .B(n22469), .Z(c[7489]) );
XNOR U37449 ( .A(a[7489]), .B(c7489), .Z(n22469) );
XOR U37450 ( .A(c7490), .B(n22470), .Z(c7491) );
ANDN U37451 ( .B(n22471), .A(n22472), .Z(n22470) );
XOR U37452 ( .A(c7490), .B(b[7490]), .Z(n22471) );
XNOR U37453 ( .A(b[7490]), .B(n22472), .Z(c[7490]) );
XNOR U37454 ( .A(a[7490]), .B(c7490), .Z(n22472) );
XOR U37455 ( .A(c7491), .B(n22473), .Z(c7492) );
ANDN U37456 ( .B(n22474), .A(n22475), .Z(n22473) );
XOR U37457 ( .A(c7491), .B(b[7491]), .Z(n22474) );
XNOR U37458 ( .A(b[7491]), .B(n22475), .Z(c[7491]) );
XNOR U37459 ( .A(a[7491]), .B(c7491), .Z(n22475) );
XOR U37460 ( .A(c7492), .B(n22476), .Z(c7493) );
ANDN U37461 ( .B(n22477), .A(n22478), .Z(n22476) );
XOR U37462 ( .A(c7492), .B(b[7492]), .Z(n22477) );
XNOR U37463 ( .A(b[7492]), .B(n22478), .Z(c[7492]) );
XNOR U37464 ( .A(a[7492]), .B(c7492), .Z(n22478) );
XOR U37465 ( .A(c7493), .B(n22479), .Z(c7494) );
ANDN U37466 ( .B(n22480), .A(n22481), .Z(n22479) );
XOR U37467 ( .A(c7493), .B(b[7493]), .Z(n22480) );
XNOR U37468 ( .A(b[7493]), .B(n22481), .Z(c[7493]) );
XNOR U37469 ( .A(a[7493]), .B(c7493), .Z(n22481) );
XOR U37470 ( .A(c7494), .B(n22482), .Z(c7495) );
ANDN U37471 ( .B(n22483), .A(n22484), .Z(n22482) );
XOR U37472 ( .A(c7494), .B(b[7494]), .Z(n22483) );
XNOR U37473 ( .A(b[7494]), .B(n22484), .Z(c[7494]) );
XNOR U37474 ( .A(a[7494]), .B(c7494), .Z(n22484) );
XOR U37475 ( .A(c7495), .B(n22485), .Z(c7496) );
ANDN U37476 ( .B(n22486), .A(n22487), .Z(n22485) );
XOR U37477 ( .A(c7495), .B(b[7495]), .Z(n22486) );
XNOR U37478 ( .A(b[7495]), .B(n22487), .Z(c[7495]) );
XNOR U37479 ( .A(a[7495]), .B(c7495), .Z(n22487) );
XOR U37480 ( .A(c7496), .B(n22488), .Z(c7497) );
ANDN U37481 ( .B(n22489), .A(n22490), .Z(n22488) );
XOR U37482 ( .A(c7496), .B(b[7496]), .Z(n22489) );
XNOR U37483 ( .A(b[7496]), .B(n22490), .Z(c[7496]) );
XNOR U37484 ( .A(a[7496]), .B(c7496), .Z(n22490) );
XOR U37485 ( .A(c7497), .B(n22491), .Z(c7498) );
ANDN U37486 ( .B(n22492), .A(n22493), .Z(n22491) );
XOR U37487 ( .A(c7497), .B(b[7497]), .Z(n22492) );
XNOR U37488 ( .A(b[7497]), .B(n22493), .Z(c[7497]) );
XNOR U37489 ( .A(a[7497]), .B(c7497), .Z(n22493) );
XOR U37490 ( .A(c7498), .B(n22494), .Z(c7499) );
ANDN U37491 ( .B(n22495), .A(n22496), .Z(n22494) );
XOR U37492 ( .A(c7498), .B(b[7498]), .Z(n22495) );
XNOR U37493 ( .A(b[7498]), .B(n22496), .Z(c[7498]) );
XNOR U37494 ( .A(a[7498]), .B(c7498), .Z(n22496) );
XOR U37495 ( .A(c7499), .B(n22497), .Z(c7500) );
ANDN U37496 ( .B(n22498), .A(n22499), .Z(n22497) );
XOR U37497 ( .A(c7499), .B(b[7499]), .Z(n22498) );
XNOR U37498 ( .A(b[7499]), .B(n22499), .Z(c[7499]) );
XNOR U37499 ( .A(a[7499]), .B(c7499), .Z(n22499) );
XOR U37500 ( .A(c7500), .B(n22500), .Z(c7501) );
ANDN U37501 ( .B(n22501), .A(n22502), .Z(n22500) );
XOR U37502 ( .A(c7500), .B(b[7500]), .Z(n22501) );
XNOR U37503 ( .A(b[7500]), .B(n22502), .Z(c[7500]) );
XNOR U37504 ( .A(a[7500]), .B(c7500), .Z(n22502) );
XOR U37505 ( .A(c7501), .B(n22503), .Z(c7502) );
ANDN U37506 ( .B(n22504), .A(n22505), .Z(n22503) );
XOR U37507 ( .A(c7501), .B(b[7501]), .Z(n22504) );
XNOR U37508 ( .A(b[7501]), .B(n22505), .Z(c[7501]) );
XNOR U37509 ( .A(a[7501]), .B(c7501), .Z(n22505) );
XOR U37510 ( .A(c7502), .B(n22506), .Z(c7503) );
ANDN U37511 ( .B(n22507), .A(n22508), .Z(n22506) );
XOR U37512 ( .A(c7502), .B(b[7502]), .Z(n22507) );
XNOR U37513 ( .A(b[7502]), .B(n22508), .Z(c[7502]) );
XNOR U37514 ( .A(a[7502]), .B(c7502), .Z(n22508) );
XOR U37515 ( .A(c7503), .B(n22509), .Z(c7504) );
ANDN U37516 ( .B(n22510), .A(n22511), .Z(n22509) );
XOR U37517 ( .A(c7503), .B(b[7503]), .Z(n22510) );
XNOR U37518 ( .A(b[7503]), .B(n22511), .Z(c[7503]) );
XNOR U37519 ( .A(a[7503]), .B(c7503), .Z(n22511) );
XOR U37520 ( .A(c7504), .B(n22512), .Z(c7505) );
ANDN U37521 ( .B(n22513), .A(n22514), .Z(n22512) );
XOR U37522 ( .A(c7504), .B(b[7504]), .Z(n22513) );
XNOR U37523 ( .A(b[7504]), .B(n22514), .Z(c[7504]) );
XNOR U37524 ( .A(a[7504]), .B(c7504), .Z(n22514) );
XOR U37525 ( .A(c7505), .B(n22515), .Z(c7506) );
ANDN U37526 ( .B(n22516), .A(n22517), .Z(n22515) );
XOR U37527 ( .A(c7505), .B(b[7505]), .Z(n22516) );
XNOR U37528 ( .A(b[7505]), .B(n22517), .Z(c[7505]) );
XNOR U37529 ( .A(a[7505]), .B(c7505), .Z(n22517) );
XOR U37530 ( .A(c7506), .B(n22518), .Z(c7507) );
ANDN U37531 ( .B(n22519), .A(n22520), .Z(n22518) );
XOR U37532 ( .A(c7506), .B(b[7506]), .Z(n22519) );
XNOR U37533 ( .A(b[7506]), .B(n22520), .Z(c[7506]) );
XNOR U37534 ( .A(a[7506]), .B(c7506), .Z(n22520) );
XOR U37535 ( .A(c7507), .B(n22521), .Z(c7508) );
ANDN U37536 ( .B(n22522), .A(n22523), .Z(n22521) );
XOR U37537 ( .A(c7507), .B(b[7507]), .Z(n22522) );
XNOR U37538 ( .A(b[7507]), .B(n22523), .Z(c[7507]) );
XNOR U37539 ( .A(a[7507]), .B(c7507), .Z(n22523) );
XOR U37540 ( .A(c7508), .B(n22524), .Z(c7509) );
ANDN U37541 ( .B(n22525), .A(n22526), .Z(n22524) );
XOR U37542 ( .A(c7508), .B(b[7508]), .Z(n22525) );
XNOR U37543 ( .A(b[7508]), .B(n22526), .Z(c[7508]) );
XNOR U37544 ( .A(a[7508]), .B(c7508), .Z(n22526) );
XOR U37545 ( .A(c7509), .B(n22527), .Z(c7510) );
ANDN U37546 ( .B(n22528), .A(n22529), .Z(n22527) );
XOR U37547 ( .A(c7509), .B(b[7509]), .Z(n22528) );
XNOR U37548 ( .A(b[7509]), .B(n22529), .Z(c[7509]) );
XNOR U37549 ( .A(a[7509]), .B(c7509), .Z(n22529) );
XOR U37550 ( .A(c7510), .B(n22530), .Z(c7511) );
ANDN U37551 ( .B(n22531), .A(n22532), .Z(n22530) );
XOR U37552 ( .A(c7510), .B(b[7510]), .Z(n22531) );
XNOR U37553 ( .A(b[7510]), .B(n22532), .Z(c[7510]) );
XNOR U37554 ( .A(a[7510]), .B(c7510), .Z(n22532) );
XOR U37555 ( .A(c7511), .B(n22533), .Z(c7512) );
ANDN U37556 ( .B(n22534), .A(n22535), .Z(n22533) );
XOR U37557 ( .A(c7511), .B(b[7511]), .Z(n22534) );
XNOR U37558 ( .A(b[7511]), .B(n22535), .Z(c[7511]) );
XNOR U37559 ( .A(a[7511]), .B(c7511), .Z(n22535) );
XOR U37560 ( .A(c7512), .B(n22536), .Z(c7513) );
ANDN U37561 ( .B(n22537), .A(n22538), .Z(n22536) );
XOR U37562 ( .A(c7512), .B(b[7512]), .Z(n22537) );
XNOR U37563 ( .A(b[7512]), .B(n22538), .Z(c[7512]) );
XNOR U37564 ( .A(a[7512]), .B(c7512), .Z(n22538) );
XOR U37565 ( .A(c7513), .B(n22539), .Z(c7514) );
ANDN U37566 ( .B(n22540), .A(n22541), .Z(n22539) );
XOR U37567 ( .A(c7513), .B(b[7513]), .Z(n22540) );
XNOR U37568 ( .A(b[7513]), .B(n22541), .Z(c[7513]) );
XNOR U37569 ( .A(a[7513]), .B(c7513), .Z(n22541) );
XOR U37570 ( .A(c7514), .B(n22542), .Z(c7515) );
ANDN U37571 ( .B(n22543), .A(n22544), .Z(n22542) );
XOR U37572 ( .A(c7514), .B(b[7514]), .Z(n22543) );
XNOR U37573 ( .A(b[7514]), .B(n22544), .Z(c[7514]) );
XNOR U37574 ( .A(a[7514]), .B(c7514), .Z(n22544) );
XOR U37575 ( .A(c7515), .B(n22545), .Z(c7516) );
ANDN U37576 ( .B(n22546), .A(n22547), .Z(n22545) );
XOR U37577 ( .A(c7515), .B(b[7515]), .Z(n22546) );
XNOR U37578 ( .A(b[7515]), .B(n22547), .Z(c[7515]) );
XNOR U37579 ( .A(a[7515]), .B(c7515), .Z(n22547) );
XOR U37580 ( .A(c7516), .B(n22548), .Z(c7517) );
ANDN U37581 ( .B(n22549), .A(n22550), .Z(n22548) );
XOR U37582 ( .A(c7516), .B(b[7516]), .Z(n22549) );
XNOR U37583 ( .A(b[7516]), .B(n22550), .Z(c[7516]) );
XNOR U37584 ( .A(a[7516]), .B(c7516), .Z(n22550) );
XOR U37585 ( .A(c7517), .B(n22551), .Z(c7518) );
ANDN U37586 ( .B(n22552), .A(n22553), .Z(n22551) );
XOR U37587 ( .A(c7517), .B(b[7517]), .Z(n22552) );
XNOR U37588 ( .A(b[7517]), .B(n22553), .Z(c[7517]) );
XNOR U37589 ( .A(a[7517]), .B(c7517), .Z(n22553) );
XOR U37590 ( .A(c7518), .B(n22554), .Z(c7519) );
ANDN U37591 ( .B(n22555), .A(n22556), .Z(n22554) );
XOR U37592 ( .A(c7518), .B(b[7518]), .Z(n22555) );
XNOR U37593 ( .A(b[7518]), .B(n22556), .Z(c[7518]) );
XNOR U37594 ( .A(a[7518]), .B(c7518), .Z(n22556) );
XOR U37595 ( .A(c7519), .B(n22557), .Z(c7520) );
ANDN U37596 ( .B(n22558), .A(n22559), .Z(n22557) );
XOR U37597 ( .A(c7519), .B(b[7519]), .Z(n22558) );
XNOR U37598 ( .A(b[7519]), .B(n22559), .Z(c[7519]) );
XNOR U37599 ( .A(a[7519]), .B(c7519), .Z(n22559) );
XOR U37600 ( .A(c7520), .B(n22560), .Z(c7521) );
ANDN U37601 ( .B(n22561), .A(n22562), .Z(n22560) );
XOR U37602 ( .A(c7520), .B(b[7520]), .Z(n22561) );
XNOR U37603 ( .A(b[7520]), .B(n22562), .Z(c[7520]) );
XNOR U37604 ( .A(a[7520]), .B(c7520), .Z(n22562) );
XOR U37605 ( .A(c7521), .B(n22563), .Z(c7522) );
ANDN U37606 ( .B(n22564), .A(n22565), .Z(n22563) );
XOR U37607 ( .A(c7521), .B(b[7521]), .Z(n22564) );
XNOR U37608 ( .A(b[7521]), .B(n22565), .Z(c[7521]) );
XNOR U37609 ( .A(a[7521]), .B(c7521), .Z(n22565) );
XOR U37610 ( .A(c7522), .B(n22566), .Z(c7523) );
ANDN U37611 ( .B(n22567), .A(n22568), .Z(n22566) );
XOR U37612 ( .A(c7522), .B(b[7522]), .Z(n22567) );
XNOR U37613 ( .A(b[7522]), .B(n22568), .Z(c[7522]) );
XNOR U37614 ( .A(a[7522]), .B(c7522), .Z(n22568) );
XOR U37615 ( .A(c7523), .B(n22569), .Z(c7524) );
ANDN U37616 ( .B(n22570), .A(n22571), .Z(n22569) );
XOR U37617 ( .A(c7523), .B(b[7523]), .Z(n22570) );
XNOR U37618 ( .A(b[7523]), .B(n22571), .Z(c[7523]) );
XNOR U37619 ( .A(a[7523]), .B(c7523), .Z(n22571) );
XOR U37620 ( .A(c7524), .B(n22572), .Z(c7525) );
ANDN U37621 ( .B(n22573), .A(n22574), .Z(n22572) );
XOR U37622 ( .A(c7524), .B(b[7524]), .Z(n22573) );
XNOR U37623 ( .A(b[7524]), .B(n22574), .Z(c[7524]) );
XNOR U37624 ( .A(a[7524]), .B(c7524), .Z(n22574) );
XOR U37625 ( .A(c7525), .B(n22575), .Z(c7526) );
ANDN U37626 ( .B(n22576), .A(n22577), .Z(n22575) );
XOR U37627 ( .A(c7525), .B(b[7525]), .Z(n22576) );
XNOR U37628 ( .A(b[7525]), .B(n22577), .Z(c[7525]) );
XNOR U37629 ( .A(a[7525]), .B(c7525), .Z(n22577) );
XOR U37630 ( .A(c7526), .B(n22578), .Z(c7527) );
ANDN U37631 ( .B(n22579), .A(n22580), .Z(n22578) );
XOR U37632 ( .A(c7526), .B(b[7526]), .Z(n22579) );
XNOR U37633 ( .A(b[7526]), .B(n22580), .Z(c[7526]) );
XNOR U37634 ( .A(a[7526]), .B(c7526), .Z(n22580) );
XOR U37635 ( .A(c7527), .B(n22581), .Z(c7528) );
ANDN U37636 ( .B(n22582), .A(n22583), .Z(n22581) );
XOR U37637 ( .A(c7527), .B(b[7527]), .Z(n22582) );
XNOR U37638 ( .A(b[7527]), .B(n22583), .Z(c[7527]) );
XNOR U37639 ( .A(a[7527]), .B(c7527), .Z(n22583) );
XOR U37640 ( .A(c7528), .B(n22584), .Z(c7529) );
ANDN U37641 ( .B(n22585), .A(n22586), .Z(n22584) );
XOR U37642 ( .A(c7528), .B(b[7528]), .Z(n22585) );
XNOR U37643 ( .A(b[7528]), .B(n22586), .Z(c[7528]) );
XNOR U37644 ( .A(a[7528]), .B(c7528), .Z(n22586) );
XOR U37645 ( .A(c7529), .B(n22587), .Z(c7530) );
ANDN U37646 ( .B(n22588), .A(n22589), .Z(n22587) );
XOR U37647 ( .A(c7529), .B(b[7529]), .Z(n22588) );
XNOR U37648 ( .A(b[7529]), .B(n22589), .Z(c[7529]) );
XNOR U37649 ( .A(a[7529]), .B(c7529), .Z(n22589) );
XOR U37650 ( .A(c7530), .B(n22590), .Z(c7531) );
ANDN U37651 ( .B(n22591), .A(n22592), .Z(n22590) );
XOR U37652 ( .A(c7530), .B(b[7530]), .Z(n22591) );
XNOR U37653 ( .A(b[7530]), .B(n22592), .Z(c[7530]) );
XNOR U37654 ( .A(a[7530]), .B(c7530), .Z(n22592) );
XOR U37655 ( .A(c7531), .B(n22593), .Z(c7532) );
ANDN U37656 ( .B(n22594), .A(n22595), .Z(n22593) );
XOR U37657 ( .A(c7531), .B(b[7531]), .Z(n22594) );
XNOR U37658 ( .A(b[7531]), .B(n22595), .Z(c[7531]) );
XNOR U37659 ( .A(a[7531]), .B(c7531), .Z(n22595) );
XOR U37660 ( .A(c7532), .B(n22596), .Z(c7533) );
ANDN U37661 ( .B(n22597), .A(n22598), .Z(n22596) );
XOR U37662 ( .A(c7532), .B(b[7532]), .Z(n22597) );
XNOR U37663 ( .A(b[7532]), .B(n22598), .Z(c[7532]) );
XNOR U37664 ( .A(a[7532]), .B(c7532), .Z(n22598) );
XOR U37665 ( .A(c7533), .B(n22599), .Z(c7534) );
ANDN U37666 ( .B(n22600), .A(n22601), .Z(n22599) );
XOR U37667 ( .A(c7533), .B(b[7533]), .Z(n22600) );
XNOR U37668 ( .A(b[7533]), .B(n22601), .Z(c[7533]) );
XNOR U37669 ( .A(a[7533]), .B(c7533), .Z(n22601) );
XOR U37670 ( .A(c7534), .B(n22602), .Z(c7535) );
ANDN U37671 ( .B(n22603), .A(n22604), .Z(n22602) );
XOR U37672 ( .A(c7534), .B(b[7534]), .Z(n22603) );
XNOR U37673 ( .A(b[7534]), .B(n22604), .Z(c[7534]) );
XNOR U37674 ( .A(a[7534]), .B(c7534), .Z(n22604) );
XOR U37675 ( .A(c7535), .B(n22605), .Z(c7536) );
ANDN U37676 ( .B(n22606), .A(n22607), .Z(n22605) );
XOR U37677 ( .A(c7535), .B(b[7535]), .Z(n22606) );
XNOR U37678 ( .A(b[7535]), .B(n22607), .Z(c[7535]) );
XNOR U37679 ( .A(a[7535]), .B(c7535), .Z(n22607) );
XOR U37680 ( .A(c7536), .B(n22608), .Z(c7537) );
ANDN U37681 ( .B(n22609), .A(n22610), .Z(n22608) );
XOR U37682 ( .A(c7536), .B(b[7536]), .Z(n22609) );
XNOR U37683 ( .A(b[7536]), .B(n22610), .Z(c[7536]) );
XNOR U37684 ( .A(a[7536]), .B(c7536), .Z(n22610) );
XOR U37685 ( .A(c7537), .B(n22611), .Z(c7538) );
ANDN U37686 ( .B(n22612), .A(n22613), .Z(n22611) );
XOR U37687 ( .A(c7537), .B(b[7537]), .Z(n22612) );
XNOR U37688 ( .A(b[7537]), .B(n22613), .Z(c[7537]) );
XNOR U37689 ( .A(a[7537]), .B(c7537), .Z(n22613) );
XOR U37690 ( .A(c7538), .B(n22614), .Z(c7539) );
ANDN U37691 ( .B(n22615), .A(n22616), .Z(n22614) );
XOR U37692 ( .A(c7538), .B(b[7538]), .Z(n22615) );
XNOR U37693 ( .A(b[7538]), .B(n22616), .Z(c[7538]) );
XNOR U37694 ( .A(a[7538]), .B(c7538), .Z(n22616) );
XOR U37695 ( .A(c7539), .B(n22617), .Z(c7540) );
ANDN U37696 ( .B(n22618), .A(n22619), .Z(n22617) );
XOR U37697 ( .A(c7539), .B(b[7539]), .Z(n22618) );
XNOR U37698 ( .A(b[7539]), .B(n22619), .Z(c[7539]) );
XNOR U37699 ( .A(a[7539]), .B(c7539), .Z(n22619) );
XOR U37700 ( .A(c7540), .B(n22620), .Z(c7541) );
ANDN U37701 ( .B(n22621), .A(n22622), .Z(n22620) );
XOR U37702 ( .A(c7540), .B(b[7540]), .Z(n22621) );
XNOR U37703 ( .A(b[7540]), .B(n22622), .Z(c[7540]) );
XNOR U37704 ( .A(a[7540]), .B(c7540), .Z(n22622) );
XOR U37705 ( .A(c7541), .B(n22623), .Z(c7542) );
ANDN U37706 ( .B(n22624), .A(n22625), .Z(n22623) );
XOR U37707 ( .A(c7541), .B(b[7541]), .Z(n22624) );
XNOR U37708 ( .A(b[7541]), .B(n22625), .Z(c[7541]) );
XNOR U37709 ( .A(a[7541]), .B(c7541), .Z(n22625) );
XOR U37710 ( .A(c7542), .B(n22626), .Z(c7543) );
ANDN U37711 ( .B(n22627), .A(n22628), .Z(n22626) );
XOR U37712 ( .A(c7542), .B(b[7542]), .Z(n22627) );
XNOR U37713 ( .A(b[7542]), .B(n22628), .Z(c[7542]) );
XNOR U37714 ( .A(a[7542]), .B(c7542), .Z(n22628) );
XOR U37715 ( .A(c7543), .B(n22629), .Z(c7544) );
ANDN U37716 ( .B(n22630), .A(n22631), .Z(n22629) );
XOR U37717 ( .A(c7543), .B(b[7543]), .Z(n22630) );
XNOR U37718 ( .A(b[7543]), .B(n22631), .Z(c[7543]) );
XNOR U37719 ( .A(a[7543]), .B(c7543), .Z(n22631) );
XOR U37720 ( .A(c7544), .B(n22632), .Z(c7545) );
ANDN U37721 ( .B(n22633), .A(n22634), .Z(n22632) );
XOR U37722 ( .A(c7544), .B(b[7544]), .Z(n22633) );
XNOR U37723 ( .A(b[7544]), .B(n22634), .Z(c[7544]) );
XNOR U37724 ( .A(a[7544]), .B(c7544), .Z(n22634) );
XOR U37725 ( .A(c7545), .B(n22635), .Z(c7546) );
ANDN U37726 ( .B(n22636), .A(n22637), .Z(n22635) );
XOR U37727 ( .A(c7545), .B(b[7545]), .Z(n22636) );
XNOR U37728 ( .A(b[7545]), .B(n22637), .Z(c[7545]) );
XNOR U37729 ( .A(a[7545]), .B(c7545), .Z(n22637) );
XOR U37730 ( .A(c7546), .B(n22638), .Z(c7547) );
ANDN U37731 ( .B(n22639), .A(n22640), .Z(n22638) );
XOR U37732 ( .A(c7546), .B(b[7546]), .Z(n22639) );
XNOR U37733 ( .A(b[7546]), .B(n22640), .Z(c[7546]) );
XNOR U37734 ( .A(a[7546]), .B(c7546), .Z(n22640) );
XOR U37735 ( .A(c7547), .B(n22641), .Z(c7548) );
ANDN U37736 ( .B(n22642), .A(n22643), .Z(n22641) );
XOR U37737 ( .A(c7547), .B(b[7547]), .Z(n22642) );
XNOR U37738 ( .A(b[7547]), .B(n22643), .Z(c[7547]) );
XNOR U37739 ( .A(a[7547]), .B(c7547), .Z(n22643) );
XOR U37740 ( .A(c7548), .B(n22644), .Z(c7549) );
ANDN U37741 ( .B(n22645), .A(n22646), .Z(n22644) );
XOR U37742 ( .A(c7548), .B(b[7548]), .Z(n22645) );
XNOR U37743 ( .A(b[7548]), .B(n22646), .Z(c[7548]) );
XNOR U37744 ( .A(a[7548]), .B(c7548), .Z(n22646) );
XOR U37745 ( .A(c7549), .B(n22647), .Z(c7550) );
ANDN U37746 ( .B(n22648), .A(n22649), .Z(n22647) );
XOR U37747 ( .A(c7549), .B(b[7549]), .Z(n22648) );
XNOR U37748 ( .A(b[7549]), .B(n22649), .Z(c[7549]) );
XNOR U37749 ( .A(a[7549]), .B(c7549), .Z(n22649) );
XOR U37750 ( .A(c7550), .B(n22650), .Z(c7551) );
ANDN U37751 ( .B(n22651), .A(n22652), .Z(n22650) );
XOR U37752 ( .A(c7550), .B(b[7550]), .Z(n22651) );
XNOR U37753 ( .A(b[7550]), .B(n22652), .Z(c[7550]) );
XNOR U37754 ( .A(a[7550]), .B(c7550), .Z(n22652) );
XOR U37755 ( .A(c7551), .B(n22653), .Z(c7552) );
ANDN U37756 ( .B(n22654), .A(n22655), .Z(n22653) );
XOR U37757 ( .A(c7551), .B(b[7551]), .Z(n22654) );
XNOR U37758 ( .A(b[7551]), .B(n22655), .Z(c[7551]) );
XNOR U37759 ( .A(a[7551]), .B(c7551), .Z(n22655) );
XOR U37760 ( .A(c7552), .B(n22656), .Z(c7553) );
ANDN U37761 ( .B(n22657), .A(n22658), .Z(n22656) );
XOR U37762 ( .A(c7552), .B(b[7552]), .Z(n22657) );
XNOR U37763 ( .A(b[7552]), .B(n22658), .Z(c[7552]) );
XNOR U37764 ( .A(a[7552]), .B(c7552), .Z(n22658) );
XOR U37765 ( .A(c7553), .B(n22659), .Z(c7554) );
ANDN U37766 ( .B(n22660), .A(n22661), .Z(n22659) );
XOR U37767 ( .A(c7553), .B(b[7553]), .Z(n22660) );
XNOR U37768 ( .A(b[7553]), .B(n22661), .Z(c[7553]) );
XNOR U37769 ( .A(a[7553]), .B(c7553), .Z(n22661) );
XOR U37770 ( .A(c7554), .B(n22662), .Z(c7555) );
ANDN U37771 ( .B(n22663), .A(n22664), .Z(n22662) );
XOR U37772 ( .A(c7554), .B(b[7554]), .Z(n22663) );
XNOR U37773 ( .A(b[7554]), .B(n22664), .Z(c[7554]) );
XNOR U37774 ( .A(a[7554]), .B(c7554), .Z(n22664) );
XOR U37775 ( .A(c7555), .B(n22665), .Z(c7556) );
ANDN U37776 ( .B(n22666), .A(n22667), .Z(n22665) );
XOR U37777 ( .A(c7555), .B(b[7555]), .Z(n22666) );
XNOR U37778 ( .A(b[7555]), .B(n22667), .Z(c[7555]) );
XNOR U37779 ( .A(a[7555]), .B(c7555), .Z(n22667) );
XOR U37780 ( .A(c7556), .B(n22668), .Z(c7557) );
ANDN U37781 ( .B(n22669), .A(n22670), .Z(n22668) );
XOR U37782 ( .A(c7556), .B(b[7556]), .Z(n22669) );
XNOR U37783 ( .A(b[7556]), .B(n22670), .Z(c[7556]) );
XNOR U37784 ( .A(a[7556]), .B(c7556), .Z(n22670) );
XOR U37785 ( .A(c7557), .B(n22671), .Z(c7558) );
ANDN U37786 ( .B(n22672), .A(n22673), .Z(n22671) );
XOR U37787 ( .A(c7557), .B(b[7557]), .Z(n22672) );
XNOR U37788 ( .A(b[7557]), .B(n22673), .Z(c[7557]) );
XNOR U37789 ( .A(a[7557]), .B(c7557), .Z(n22673) );
XOR U37790 ( .A(c7558), .B(n22674), .Z(c7559) );
ANDN U37791 ( .B(n22675), .A(n22676), .Z(n22674) );
XOR U37792 ( .A(c7558), .B(b[7558]), .Z(n22675) );
XNOR U37793 ( .A(b[7558]), .B(n22676), .Z(c[7558]) );
XNOR U37794 ( .A(a[7558]), .B(c7558), .Z(n22676) );
XOR U37795 ( .A(c7559), .B(n22677), .Z(c7560) );
ANDN U37796 ( .B(n22678), .A(n22679), .Z(n22677) );
XOR U37797 ( .A(c7559), .B(b[7559]), .Z(n22678) );
XNOR U37798 ( .A(b[7559]), .B(n22679), .Z(c[7559]) );
XNOR U37799 ( .A(a[7559]), .B(c7559), .Z(n22679) );
XOR U37800 ( .A(c7560), .B(n22680), .Z(c7561) );
ANDN U37801 ( .B(n22681), .A(n22682), .Z(n22680) );
XOR U37802 ( .A(c7560), .B(b[7560]), .Z(n22681) );
XNOR U37803 ( .A(b[7560]), .B(n22682), .Z(c[7560]) );
XNOR U37804 ( .A(a[7560]), .B(c7560), .Z(n22682) );
XOR U37805 ( .A(c7561), .B(n22683), .Z(c7562) );
ANDN U37806 ( .B(n22684), .A(n22685), .Z(n22683) );
XOR U37807 ( .A(c7561), .B(b[7561]), .Z(n22684) );
XNOR U37808 ( .A(b[7561]), .B(n22685), .Z(c[7561]) );
XNOR U37809 ( .A(a[7561]), .B(c7561), .Z(n22685) );
XOR U37810 ( .A(c7562), .B(n22686), .Z(c7563) );
ANDN U37811 ( .B(n22687), .A(n22688), .Z(n22686) );
XOR U37812 ( .A(c7562), .B(b[7562]), .Z(n22687) );
XNOR U37813 ( .A(b[7562]), .B(n22688), .Z(c[7562]) );
XNOR U37814 ( .A(a[7562]), .B(c7562), .Z(n22688) );
XOR U37815 ( .A(c7563), .B(n22689), .Z(c7564) );
ANDN U37816 ( .B(n22690), .A(n22691), .Z(n22689) );
XOR U37817 ( .A(c7563), .B(b[7563]), .Z(n22690) );
XNOR U37818 ( .A(b[7563]), .B(n22691), .Z(c[7563]) );
XNOR U37819 ( .A(a[7563]), .B(c7563), .Z(n22691) );
XOR U37820 ( .A(c7564), .B(n22692), .Z(c7565) );
ANDN U37821 ( .B(n22693), .A(n22694), .Z(n22692) );
XOR U37822 ( .A(c7564), .B(b[7564]), .Z(n22693) );
XNOR U37823 ( .A(b[7564]), .B(n22694), .Z(c[7564]) );
XNOR U37824 ( .A(a[7564]), .B(c7564), .Z(n22694) );
XOR U37825 ( .A(c7565), .B(n22695), .Z(c7566) );
ANDN U37826 ( .B(n22696), .A(n22697), .Z(n22695) );
XOR U37827 ( .A(c7565), .B(b[7565]), .Z(n22696) );
XNOR U37828 ( .A(b[7565]), .B(n22697), .Z(c[7565]) );
XNOR U37829 ( .A(a[7565]), .B(c7565), .Z(n22697) );
XOR U37830 ( .A(c7566), .B(n22698), .Z(c7567) );
ANDN U37831 ( .B(n22699), .A(n22700), .Z(n22698) );
XOR U37832 ( .A(c7566), .B(b[7566]), .Z(n22699) );
XNOR U37833 ( .A(b[7566]), .B(n22700), .Z(c[7566]) );
XNOR U37834 ( .A(a[7566]), .B(c7566), .Z(n22700) );
XOR U37835 ( .A(c7567), .B(n22701), .Z(c7568) );
ANDN U37836 ( .B(n22702), .A(n22703), .Z(n22701) );
XOR U37837 ( .A(c7567), .B(b[7567]), .Z(n22702) );
XNOR U37838 ( .A(b[7567]), .B(n22703), .Z(c[7567]) );
XNOR U37839 ( .A(a[7567]), .B(c7567), .Z(n22703) );
XOR U37840 ( .A(c7568), .B(n22704), .Z(c7569) );
ANDN U37841 ( .B(n22705), .A(n22706), .Z(n22704) );
XOR U37842 ( .A(c7568), .B(b[7568]), .Z(n22705) );
XNOR U37843 ( .A(b[7568]), .B(n22706), .Z(c[7568]) );
XNOR U37844 ( .A(a[7568]), .B(c7568), .Z(n22706) );
XOR U37845 ( .A(c7569), .B(n22707), .Z(c7570) );
ANDN U37846 ( .B(n22708), .A(n22709), .Z(n22707) );
XOR U37847 ( .A(c7569), .B(b[7569]), .Z(n22708) );
XNOR U37848 ( .A(b[7569]), .B(n22709), .Z(c[7569]) );
XNOR U37849 ( .A(a[7569]), .B(c7569), .Z(n22709) );
XOR U37850 ( .A(c7570), .B(n22710), .Z(c7571) );
ANDN U37851 ( .B(n22711), .A(n22712), .Z(n22710) );
XOR U37852 ( .A(c7570), .B(b[7570]), .Z(n22711) );
XNOR U37853 ( .A(b[7570]), .B(n22712), .Z(c[7570]) );
XNOR U37854 ( .A(a[7570]), .B(c7570), .Z(n22712) );
XOR U37855 ( .A(c7571), .B(n22713), .Z(c7572) );
ANDN U37856 ( .B(n22714), .A(n22715), .Z(n22713) );
XOR U37857 ( .A(c7571), .B(b[7571]), .Z(n22714) );
XNOR U37858 ( .A(b[7571]), .B(n22715), .Z(c[7571]) );
XNOR U37859 ( .A(a[7571]), .B(c7571), .Z(n22715) );
XOR U37860 ( .A(c7572), .B(n22716), .Z(c7573) );
ANDN U37861 ( .B(n22717), .A(n22718), .Z(n22716) );
XOR U37862 ( .A(c7572), .B(b[7572]), .Z(n22717) );
XNOR U37863 ( .A(b[7572]), .B(n22718), .Z(c[7572]) );
XNOR U37864 ( .A(a[7572]), .B(c7572), .Z(n22718) );
XOR U37865 ( .A(c7573), .B(n22719), .Z(c7574) );
ANDN U37866 ( .B(n22720), .A(n22721), .Z(n22719) );
XOR U37867 ( .A(c7573), .B(b[7573]), .Z(n22720) );
XNOR U37868 ( .A(b[7573]), .B(n22721), .Z(c[7573]) );
XNOR U37869 ( .A(a[7573]), .B(c7573), .Z(n22721) );
XOR U37870 ( .A(c7574), .B(n22722), .Z(c7575) );
ANDN U37871 ( .B(n22723), .A(n22724), .Z(n22722) );
XOR U37872 ( .A(c7574), .B(b[7574]), .Z(n22723) );
XNOR U37873 ( .A(b[7574]), .B(n22724), .Z(c[7574]) );
XNOR U37874 ( .A(a[7574]), .B(c7574), .Z(n22724) );
XOR U37875 ( .A(c7575), .B(n22725), .Z(c7576) );
ANDN U37876 ( .B(n22726), .A(n22727), .Z(n22725) );
XOR U37877 ( .A(c7575), .B(b[7575]), .Z(n22726) );
XNOR U37878 ( .A(b[7575]), .B(n22727), .Z(c[7575]) );
XNOR U37879 ( .A(a[7575]), .B(c7575), .Z(n22727) );
XOR U37880 ( .A(c7576), .B(n22728), .Z(c7577) );
ANDN U37881 ( .B(n22729), .A(n22730), .Z(n22728) );
XOR U37882 ( .A(c7576), .B(b[7576]), .Z(n22729) );
XNOR U37883 ( .A(b[7576]), .B(n22730), .Z(c[7576]) );
XNOR U37884 ( .A(a[7576]), .B(c7576), .Z(n22730) );
XOR U37885 ( .A(c7577), .B(n22731), .Z(c7578) );
ANDN U37886 ( .B(n22732), .A(n22733), .Z(n22731) );
XOR U37887 ( .A(c7577), .B(b[7577]), .Z(n22732) );
XNOR U37888 ( .A(b[7577]), .B(n22733), .Z(c[7577]) );
XNOR U37889 ( .A(a[7577]), .B(c7577), .Z(n22733) );
XOR U37890 ( .A(c7578), .B(n22734), .Z(c7579) );
ANDN U37891 ( .B(n22735), .A(n22736), .Z(n22734) );
XOR U37892 ( .A(c7578), .B(b[7578]), .Z(n22735) );
XNOR U37893 ( .A(b[7578]), .B(n22736), .Z(c[7578]) );
XNOR U37894 ( .A(a[7578]), .B(c7578), .Z(n22736) );
XOR U37895 ( .A(c7579), .B(n22737), .Z(c7580) );
ANDN U37896 ( .B(n22738), .A(n22739), .Z(n22737) );
XOR U37897 ( .A(c7579), .B(b[7579]), .Z(n22738) );
XNOR U37898 ( .A(b[7579]), .B(n22739), .Z(c[7579]) );
XNOR U37899 ( .A(a[7579]), .B(c7579), .Z(n22739) );
XOR U37900 ( .A(c7580), .B(n22740), .Z(c7581) );
ANDN U37901 ( .B(n22741), .A(n22742), .Z(n22740) );
XOR U37902 ( .A(c7580), .B(b[7580]), .Z(n22741) );
XNOR U37903 ( .A(b[7580]), .B(n22742), .Z(c[7580]) );
XNOR U37904 ( .A(a[7580]), .B(c7580), .Z(n22742) );
XOR U37905 ( .A(c7581), .B(n22743), .Z(c7582) );
ANDN U37906 ( .B(n22744), .A(n22745), .Z(n22743) );
XOR U37907 ( .A(c7581), .B(b[7581]), .Z(n22744) );
XNOR U37908 ( .A(b[7581]), .B(n22745), .Z(c[7581]) );
XNOR U37909 ( .A(a[7581]), .B(c7581), .Z(n22745) );
XOR U37910 ( .A(c7582), .B(n22746), .Z(c7583) );
ANDN U37911 ( .B(n22747), .A(n22748), .Z(n22746) );
XOR U37912 ( .A(c7582), .B(b[7582]), .Z(n22747) );
XNOR U37913 ( .A(b[7582]), .B(n22748), .Z(c[7582]) );
XNOR U37914 ( .A(a[7582]), .B(c7582), .Z(n22748) );
XOR U37915 ( .A(c7583), .B(n22749), .Z(c7584) );
ANDN U37916 ( .B(n22750), .A(n22751), .Z(n22749) );
XOR U37917 ( .A(c7583), .B(b[7583]), .Z(n22750) );
XNOR U37918 ( .A(b[7583]), .B(n22751), .Z(c[7583]) );
XNOR U37919 ( .A(a[7583]), .B(c7583), .Z(n22751) );
XOR U37920 ( .A(c7584), .B(n22752), .Z(c7585) );
ANDN U37921 ( .B(n22753), .A(n22754), .Z(n22752) );
XOR U37922 ( .A(c7584), .B(b[7584]), .Z(n22753) );
XNOR U37923 ( .A(b[7584]), .B(n22754), .Z(c[7584]) );
XNOR U37924 ( .A(a[7584]), .B(c7584), .Z(n22754) );
XOR U37925 ( .A(c7585), .B(n22755), .Z(c7586) );
ANDN U37926 ( .B(n22756), .A(n22757), .Z(n22755) );
XOR U37927 ( .A(c7585), .B(b[7585]), .Z(n22756) );
XNOR U37928 ( .A(b[7585]), .B(n22757), .Z(c[7585]) );
XNOR U37929 ( .A(a[7585]), .B(c7585), .Z(n22757) );
XOR U37930 ( .A(c7586), .B(n22758), .Z(c7587) );
ANDN U37931 ( .B(n22759), .A(n22760), .Z(n22758) );
XOR U37932 ( .A(c7586), .B(b[7586]), .Z(n22759) );
XNOR U37933 ( .A(b[7586]), .B(n22760), .Z(c[7586]) );
XNOR U37934 ( .A(a[7586]), .B(c7586), .Z(n22760) );
XOR U37935 ( .A(c7587), .B(n22761), .Z(c7588) );
ANDN U37936 ( .B(n22762), .A(n22763), .Z(n22761) );
XOR U37937 ( .A(c7587), .B(b[7587]), .Z(n22762) );
XNOR U37938 ( .A(b[7587]), .B(n22763), .Z(c[7587]) );
XNOR U37939 ( .A(a[7587]), .B(c7587), .Z(n22763) );
XOR U37940 ( .A(c7588), .B(n22764), .Z(c7589) );
ANDN U37941 ( .B(n22765), .A(n22766), .Z(n22764) );
XOR U37942 ( .A(c7588), .B(b[7588]), .Z(n22765) );
XNOR U37943 ( .A(b[7588]), .B(n22766), .Z(c[7588]) );
XNOR U37944 ( .A(a[7588]), .B(c7588), .Z(n22766) );
XOR U37945 ( .A(c7589), .B(n22767), .Z(c7590) );
ANDN U37946 ( .B(n22768), .A(n22769), .Z(n22767) );
XOR U37947 ( .A(c7589), .B(b[7589]), .Z(n22768) );
XNOR U37948 ( .A(b[7589]), .B(n22769), .Z(c[7589]) );
XNOR U37949 ( .A(a[7589]), .B(c7589), .Z(n22769) );
XOR U37950 ( .A(c7590), .B(n22770), .Z(c7591) );
ANDN U37951 ( .B(n22771), .A(n22772), .Z(n22770) );
XOR U37952 ( .A(c7590), .B(b[7590]), .Z(n22771) );
XNOR U37953 ( .A(b[7590]), .B(n22772), .Z(c[7590]) );
XNOR U37954 ( .A(a[7590]), .B(c7590), .Z(n22772) );
XOR U37955 ( .A(c7591), .B(n22773), .Z(c7592) );
ANDN U37956 ( .B(n22774), .A(n22775), .Z(n22773) );
XOR U37957 ( .A(c7591), .B(b[7591]), .Z(n22774) );
XNOR U37958 ( .A(b[7591]), .B(n22775), .Z(c[7591]) );
XNOR U37959 ( .A(a[7591]), .B(c7591), .Z(n22775) );
XOR U37960 ( .A(c7592), .B(n22776), .Z(c7593) );
ANDN U37961 ( .B(n22777), .A(n22778), .Z(n22776) );
XOR U37962 ( .A(c7592), .B(b[7592]), .Z(n22777) );
XNOR U37963 ( .A(b[7592]), .B(n22778), .Z(c[7592]) );
XNOR U37964 ( .A(a[7592]), .B(c7592), .Z(n22778) );
XOR U37965 ( .A(c7593), .B(n22779), .Z(c7594) );
ANDN U37966 ( .B(n22780), .A(n22781), .Z(n22779) );
XOR U37967 ( .A(c7593), .B(b[7593]), .Z(n22780) );
XNOR U37968 ( .A(b[7593]), .B(n22781), .Z(c[7593]) );
XNOR U37969 ( .A(a[7593]), .B(c7593), .Z(n22781) );
XOR U37970 ( .A(c7594), .B(n22782), .Z(c7595) );
ANDN U37971 ( .B(n22783), .A(n22784), .Z(n22782) );
XOR U37972 ( .A(c7594), .B(b[7594]), .Z(n22783) );
XNOR U37973 ( .A(b[7594]), .B(n22784), .Z(c[7594]) );
XNOR U37974 ( .A(a[7594]), .B(c7594), .Z(n22784) );
XOR U37975 ( .A(c7595), .B(n22785), .Z(c7596) );
ANDN U37976 ( .B(n22786), .A(n22787), .Z(n22785) );
XOR U37977 ( .A(c7595), .B(b[7595]), .Z(n22786) );
XNOR U37978 ( .A(b[7595]), .B(n22787), .Z(c[7595]) );
XNOR U37979 ( .A(a[7595]), .B(c7595), .Z(n22787) );
XOR U37980 ( .A(c7596), .B(n22788), .Z(c7597) );
ANDN U37981 ( .B(n22789), .A(n22790), .Z(n22788) );
XOR U37982 ( .A(c7596), .B(b[7596]), .Z(n22789) );
XNOR U37983 ( .A(b[7596]), .B(n22790), .Z(c[7596]) );
XNOR U37984 ( .A(a[7596]), .B(c7596), .Z(n22790) );
XOR U37985 ( .A(c7597), .B(n22791), .Z(c7598) );
ANDN U37986 ( .B(n22792), .A(n22793), .Z(n22791) );
XOR U37987 ( .A(c7597), .B(b[7597]), .Z(n22792) );
XNOR U37988 ( .A(b[7597]), .B(n22793), .Z(c[7597]) );
XNOR U37989 ( .A(a[7597]), .B(c7597), .Z(n22793) );
XOR U37990 ( .A(c7598), .B(n22794), .Z(c7599) );
ANDN U37991 ( .B(n22795), .A(n22796), .Z(n22794) );
XOR U37992 ( .A(c7598), .B(b[7598]), .Z(n22795) );
XNOR U37993 ( .A(b[7598]), .B(n22796), .Z(c[7598]) );
XNOR U37994 ( .A(a[7598]), .B(c7598), .Z(n22796) );
XOR U37995 ( .A(c7599), .B(n22797), .Z(c7600) );
ANDN U37996 ( .B(n22798), .A(n22799), .Z(n22797) );
XOR U37997 ( .A(c7599), .B(b[7599]), .Z(n22798) );
XNOR U37998 ( .A(b[7599]), .B(n22799), .Z(c[7599]) );
XNOR U37999 ( .A(a[7599]), .B(c7599), .Z(n22799) );
XOR U38000 ( .A(c7600), .B(n22800), .Z(c7601) );
ANDN U38001 ( .B(n22801), .A(n22802), .Z(n22800) );
XOR U38002 ( .A(c7600), .B(b[7600]), .Z(n22801) );
XNOR U38003 ( .A(b[7600]), .B(n22802), .Z(c[7600]) );
XNOR U38004 ( .A(a[7600]), .B(c7600), .Z(n22802) );
XOR U38005 ( .A(c7601), .B(n22803), .Z(c7602) );
ANDN U38006 ( .B(n22804), .A(n22805), .Z(n22803) );
XOR U38007 ( .A(c7601), .B(b[7601]), .Z(n22804) );
XNOR U38008 ( .A(b[7601]), .B(n22805), .Z(c[7601]) );
XNOR U38009 ( .A(a[7601]), .B(c7601), .Z(n22805) );
XOR U38010 ( .A(c7602), .B(n22806), .Z(c7603) );
ANDN U38011 ( .B(n22807), .A(n22808), .Z(n22806) );
XOR U38012 ( .A(c7602), .B(b[7602]), .Z(n22807) );
XNOR U38013 ( .A(b[7602]), .B(n22808), .Z(c[7602]) );
XNOR U38014 ( .A(a[7602]), .B(c7602), .Z(n22808) );
XOR U38015 ( .A(c7603), .B(n22809), .Z(c7604) );
ANDN U38016 ( .B(n22810), .A(n22811), .Z(n22809) );
XOR U38017 ( .A(c7603), .B(b[7603]), .Z(n22810) );
XNOR U38018 ( .A(b[7603]), .B(n22811), .Z(c[7603]) );
XNOR U38019 ( .A(a[7603]), .B(c7603), .Z(n22811) );
XOR U38020 ( .A(c7604), .B(n22812), .Z(c7605) );
ANDN U38021 ( .B(n22813), .A(n22814), .Z(n22812) );
XOR U38022 ( .A(c7604), .B(b[7604]), .Z(n22813) );
XNOR U38023 ( .A(b[7604]), .B(n22814), .Z(c[7604]) );
XNOR U38024 ( .A(a[7604]), .B(c7604), .Z(n22814) );
XOR U38025 ( .A(c7605), .B(n22815), .Z(c7606) );
ANDN U38026 ( .B(n22816), .A(n22817), .Z(n22815) );
XOR U38027 ( .A(c7605), .B(b[7605]), .Z(n22816) );
XNOR U38028 ( .A(b[7605]), .B(n22817), .Z(c[7605]) );
XNOR U38029 ( .A(a[7605]), .B(c7605), .Z(n22817) );
XOR U38030 ( .A(c7606), .B(n22818), .Z(c7607) );
ANDN U38031 ( .B(n22819), .A(n22820), .Z(n22818) );
XOR U38032 ( .A(c7606), .B(b[7606]), .Z(n22819) );
XNOR U38033 ( .A(b[7606]), .B(n22820), .Z(c[7606]) );
XNOR U38034 ( .A(a[7606]), .B(c7606), .Z(n22820) );
XOR U38035 ( .A(c7607), .B(n22821), .Z(c7608) );
ANDN U38036 ( .B(n22822), .A(n22823), .Z(n22821) );
XOR U38037 ( .A(c7607), .B(b[7607]), .Z(n22822) );
XNOR U38038 ( .A(b[7607]), .B(n22823), .Z(c[7607]) );
XNOR U38039 ( .A(a[7607]), .B(c7607), .Z(n22823) );
XOR U38040 ( .A(c7608), .B(n22824), .Z(c7609) );
ANDN U38041 ( .B(n22825), .A(n22826), .Z(n22824) );
XOR U38042 ( .A(c7608), .B(b[7608]), .Z(n22825) );
XNOR U38043 ( .A(b[7608]), .B(n22826), .Z(c[7608]) );
XNOR U38044 ( .A(a[7608]), .B(c7608), .Z(n22826) );
XOR U38045 ( .A(c7609), .B(n22827), .Z(c7610) );
ANDN U38046 ( .B(n22828), .A(n22829), .Z(n22827) );
XOR U38047 ( .A(c7609), .B(b[7609]), .Z(n22828) );
XNOR U38048 ( .A(b[7609]), .B(n22829), .Z(c[7609]) );
XNOR U38049 ( .A(a[7609]), .B(c7609), .Z(n22829) );
XOR U38050 ( .A(c7610), .B(n22830), .Z(c7611) );
ANDN U38051 ( .B(n22831), .A(n22832), .Z(n22830) );
XOR U38052 ( .A(c7610), .B(b[7610]), .Z(n22831) );
XNOR U38053 ( .A(b[7610]), .B(n22832), .Z(c[7610]) );
XNOR U38054 ( .A(a[7610]), .B(c7610), .Z(n22832) );
XOR U38055 ( .A(c7611), .B(n22833), .Z(c7612) );
ANDN U38056 ( .B(n22834), .A(n22835), .Z(n22833) );
XOR U38057 ( .A(c7611), .B(b[7611]), .Z(n22834) );
XNOR U38058 ( .A(b[7611]), .B(n22835), .Z(c[7611]) );
XNOR U38059 ( .A(a[7611]), .B(c7611), .Z(n22835) );
XOR U38060 ( .A(c7612), .B(n22836), .Z(c7613) );
ANDN U38061 ( .B(n22837), .A(n22838), .Z(n22836) );
XOR U38062 ( .A(c7612), .B(b[7612]), .Z(n22837) );
XNOR U38063 ( .A(b[7612]), .B(n22838), .Z(c[7612]) );
XNOR U38064 ( .A(a[7612]), .B(c7612), .Z(n22838) );
XOR U38065 ( .A(c7613), .B(n22839), .Z(c7614) );
ANDN U38066 ( .B(n22840), .A(n22841), .Z(n22839) );
XOR U38067 ( .A(c7613), .B(b[7613]), .Z(n22840) );
XNOR U38068 ( .A(b[7613]), .B(n22841), .Z(c[7613]) );
XNOR U38069 ( .A(a[7613]), .B(c7613), .Z(n22841) );
XOR U38070 ( .A(c7614), .B(n22842), .Z(c7615) );
ANDN U38071 ( .B(n22843), .A(n22844), .Z(n22842) );
XOR U38072 ( .A(c7614), .B(b[7614]), .Z(n22843) );
XNOR U38073 ( .A(b[7614]), .B(n22844), .Z(c[7614]) );
XNOR U38074 ( .A(a[7614]), .B(c7614), .Z(n22844) );
XOR U38075 ( .A(c7615), .B(n22845), .Z(c7616) );
ANDN U38076 ( .B(n22846), .A(n22847), .Z(n22845) );
XOR U38077 ( .A(c7615), .B(b[7615]), .Z(n22846) );
XNOR U38078 ( .A(b[7615]), .B(n22847), .Z(c[7615]) );
XNOR U38079 ( .A(a[7615]), .B(c7615), .Z(n22847) );
XOR U38080 ( .A(c7616), .B(n22848), .Z(c7617) );
ANDN U38081 ( .B(n22849), .A(n22850), .Z(n22848) );
XOR U38082 ( .A(c7616), .B(b[7616]), .Z(n22849) );
XNOR U38083 ( .A(b[7616]), .B(n22850), .Z(c[7616]) );
XNOR U38084 ( .A(a[7616]), .B(c7616), .Z(n22850) );
XOR U38085 ( .A(c7617), .B(n22851), .Z(c7618) );
ANDN U38086 ( .B(n22852), .A(n22853), .Z(n22851) );
XOR U38087 ( .A(c7617), .B(b[7617]), .Z(n22852) );
XNOR U38088 ( .A(b[7617]), .B(n22853), .Z(c[7617]) );
XNOR U38089 ( .A(a[7617]), .B(c7617), .Z(n22853) );
XOR U38090 ( .A(c7618), .B(n22854), .Z(c7619) );
ANDN U38091 ( .B(n22855), .A(n22856), .Z(n22854) );
XOR U38092 ( .A(c7618), .B(b[7618]), .Z(n22855) );
XNOR U38093 ( .A(b[7618]), .B(n22856), .Z(c[7618]) );
XNOR U38094 ( .A(a[7618]), .B(c7618), .Z(n22856) );
XOR U38095 ( .A(c7619), .B(n22857), .Z(c7620) );
ANDN U38096 ( .B(n22858), .A(n22859), .Z(n22857) );
XOR U38097 ( .A(c7619), .B(b[7619]), .Z(n22858) );
XNOR U38098 ( .A(b[7619]), .B(n22859), .Z(c[7619]) );
XNOR U38099 ( .A(a[7619]), .B(c7619), .Z(n22859) );
XOR U38100 ( .A(c7620), .B(n22860), .Z(c7621) );
ANDN U38101 ( .B(n22861), .A(n22862), .Z(n22860) );
XOR U38102 ( .A(c7620), .B(b[7620]), .Z(n22861) );
XNOR U38103 ( .A(b[7620]), .B(n22862), .Z(c[7620]) );
XNOR U38104 ( .A(a[7620]), .B(c7620), .Z(n22862) );
XOR U38105 ( .A(c7621), .B(n22863), .Z(c7622) );
ANDN U38106 ( .B(n22864), .A(n22865), .Z(n22863) );
XOR U38107 ( .A(c7621), .B(b[7621]), .Z(n22864) );
XNOR U38108 ( .A(b[7621]), .B(n22865), .Z(c[7621]) );
XNOR U38109 ( .A(a[7621]), .B(c7621), .Z(n22865) );
XOR U38110 ( .A(c7622), .B(n22866), .Z(c7623) );
ANDN U38111 ( .B(n22867), .A(n22868), .Z(n22866) );
XOR U38112 ( .A(c7622), .B(b[7622]), .Z(n22867) );
XNOR U38113 ( .A(b[7622]), .B(n22868), .Z(c[7622]) );
XNOR U38114 ( .A(a[7622]), .B(c7622), .Z(n22868) );
XOR U38115 ( .A(c7623), .B(n22869), .Z(c7624) );
ANDN U38116 ( .B(n22870), .A(n22871), .Z(n22869) );
XOR U38117 ( .A(c7623), .B(b[7623]), .Z(n22870) );
XNOR U38118 ( .A(b[7623]), .B(n22871), .Z(c[7623]) );
XNOR U38119 ( .A(a[7623]), .B(c7623), .Z(n22871) );
XOR U38120 ( .A(c7624), .B(n22872), .Z(c7625) );
ANDN U38121 ( .B(n22873), .A(n22874), .Z(n22872) );
XOR U38122 ( .A(c7624), .B(b[7624]), .Z(n22873) );
XNOR U38123 ( .A(b[7624]), .B(n22874), .Z(c[7624]) );
XNOR U38124 ( .A(a[7624]), .B(c7624), .Z(n22874) );
XOR U38125 ( .A(c7625), .B(n22875), .Z(c7626) );
ANDN U38126 ( .B(n22876), .A(n22877), .Z(n22875) );
XOR U38127 ( .A(c7625), .B(b[7625]), .Z(n22876) );
XNOR U38128 ( .A(b[7625]), .B(n22877), .Z(c[7625]) );
XNOR U38129 ( .A(a[7625]), .B(c7625), .Z(n22877) );
XOR U38130 ( .A(c7626), .B(n22878), .Z(c7627) );
ANDN U38131 ( .B(n22879), .A(n22880), .Z(n22878) );
XOR U38132 ( .A(c7626), .B(b[7626]), .Z(n22879) );
XNOR U38133 ( .A(b[7626]), .B(n22880), .Z(c[7626]) );
XNOR U38134 ( .A(a[7626]), .B(c7626), .Z(n22880) );
XOR U38135 ( .A(c7627), .B(n22881), .Z(c7628) );
ANDN U38136 ( .B(n22882), .A(n22883), .Z(n22881) );
XOR U38137 ( .A(c7627), .B(b[7627]), .Z(n22882) );
XNOR U38138 ( .A(b[7627]), .B(n22883), .Z(c[7627]) );
XNOR U38139 ( .A(a[7627]), .B(c7627), .Z(n22883) );
XOR U38140 ( .A(c7628), .B(n22884), .Z(c7629) );
ANDN U38141 ( .B(n22885), .A(n22886), .Z(n22884) );
XOR U38142 ( .A(c7628), .B(b[7628]), .Z(n22885) );
XNOR U38143 ( .A(b[7628]), .B(n22886), .Z(c[7628]) );
XNOR U38144 ( .A(a[7628]), .B(c7628), .Z(n22886) );
XOR U38145 ( .A(c7629), .B(n22887), .Z(c7630) );
ANDN U38146 ( .B(n22888), .A(n22889), .Z(n22887) );
XOR U38147 ( .A(c7629), .B(b[7629]), .Z(n22888) );
XNOR U38148 ( .A(b[7629]), .B(n22889), .Z(c[7629]) );
XNOR U38149 ( .A(a[7629]), .B(c7629), .Z(n22889) );
XOR U38150 ( .A(c7630), .B(n22890), .Z(c7631) );
ANDN U38151 ( .B(n22891), .A(n22892), .Z(n22890) );
XOR U38152 ( .A(c7630), .B(b[7630]), .Z(n22891) );
XNOR U38153 ( .A(b[7630]), .B(n22892), .Z(c[7630]) );
XNOR U38154 ( .A(a[7630]), .B(c7630), .Z(n22892) );
XOR U38155 ( .A(c7631), .B(n22893), .Z(c7632) );
ANDN U38156 ( .B(n22894), .A(n22895), .Z(n22893) );
XOR U38157 ( .A(c7631), .B(b[7631]), .Z(n22894) );
XNOR U38158 ( .A(b[7631]), .B(n22895), .Z(c[7631]) );
XNOR U38159 ( .A(a[7631]), .B(c7631), .Z(n22895) );
XOR U38160 ( .A(c7632), .B(n22896), .Z(c7633) );
ANDN U38161 ( .B(n22897), .A(n22898), .Z(n22896) );
XOR U38162 ( .A(c7632), .B(b[7632]), .Z(n22897) );
XNOR U38163 ( .A(b[7632]), .B(n22898), .Z(c[7632]) );
XNOR U38164 ( .A(a[7632]), .B(c7632), .Z(n22898) );
XOR U38165 ( .A(c7633), .B(n22899), .Z(c7634) );
ANDN U38166 ( .B(n22900), .A(n22901), .Z(n22899) );
XOR U38167 ( .A(c7633), .B(b[7633]), .Z(n22900) );
XNOR U38168 ( .A(b[7633]), .B(n22901), .Z(c[7633]) );
XNOR U38169 ( .A(a[7633]), .B(c7633), .Z(n22901) );
XOR U38170 ( .A(c7634), .B(n22902), .Z(c7635) );
ANDN U38171 ( .B(n22903), .A(n22904), .Z(n22902) );
XOR U38172 ( .A(c7634), .B(b[7634]), .Z(n22903) );
XNOR U38173 ( .A(b[7634]), .B(n22904), .Z(c[7634]) );
XNOR U38174 ( .A(a[7634]), .B(c7634), .Z(n22904) );
XOR U38175 ( .A(c7635), .B(n22905), .Z(c7636) );
ANDN U38176 ( .B(n22906), .A(n22907), .Z(n22905) );
XOR U38177 ( .A(c7635), .B(b[7635]), .Z(n22906) );
XNOR U38178 ( .A(b[7635]), .B(n22907), .Z(c[7635]) );
XNOR U38179 ( .A(a[7635]), .B(c7635), .Z(n22907) );
XOR U38180 ( .A(c7636), .B(n22908), .Z(c7637) );
ANDN U38181 ( .B(n22909), .A(n22910), .Z(n22908) );
XOR U38182 ( .A(c7636), .B(b[7636]), .Z(n22909) );
XNOR U38183 ( .A(b[7636]), .B(n22910), .Z(c[7636]) );
XNOR U38184 ( .A(a[7636]), .B(c7636), .Z(n22910) );
XOR U38185 ( .A(c7637), .B(n22911), .Z(c7638) );
ANDN U38186 ( .B(n22912), .A(n22913), .Z(n22911) );
XOR U38187 ( .A(c7637), .B(b[7637]), .Z(n22912) );
XNOR U38188 ( .A(b[7637]), .B(n22913), .Z(c[7637]) );
XNOR U38189 ( .A(a[7637]), .B(c7637), .Z(n22913) );
XOR U38190 ( .A(c7638), .B(n22914), .Z(c7639) );
ANDN U38191 ( .B(n22915), .A(n22916), .Z(n22914) );
XOR U38192 ( .A(c7638), .B(b[7638]), .Z(n22915) );
XNOR U38193 ( .A(b[7638]), .B(n22916), .Z(c[7638]) );
XNOR U38194 ( .A(a[7638]), .B(c7638), .Z(n22916) );
XOR U38195 ( .A(c7639), .B(n22917), .Z(c7640) );
ANDN U38196 ( .B(n22918), .A(n22919), .Z(n22917) );
XOR U38197 ( .A(c7639), .B(b[7639]), .Z(n22918) );
XNOR U38198 ( .A(b[7639]), .B(n22919), .Z(c[7639]) );
XNOR U38199 ( .A(a[7639]), .B(c7639), .Z(n22919) );
XOR U38200 ( .A(c7640), .B(n22920), .Z(c7641) );
ANDN U38201 ( .B(n22921), .A(n22922), .Z(n22920) );
XOR U38202 ( .A(c7640), .B(b[7640]), .Z(n22921) );
XNOR U38203 ( .A(b[7640]), .B(n22922), .Z(c[7640]) );
XNOR U38204 ( .A(a[7640]), .B(c7640), .Z(n22922) );
XOR U38205 ( .A(c7641), .B(n22923), .Z(c7642) );
ANDN U38206 ( .B(n22924), .A(n22925), .Z(n22923) );
XOR U38207 ( .A(c7641), .B(b[7641]), .Z(n22924) );
XNOR U38208 ( .A(b[7641]), .B(n22925), .Z(c[7641]) );
XNOR U38209 ( .A(a[7641]), .B(c7641), .Z(n22925) );
XOR U38210 ( .A(c7642), .B(n22926), .Z(c7643) );
ANDN U38211 ( .B(n22927), .A(n22928), .Z(n22926) );
XOR U38212 ( .A(c7642), .B(b[7642]), .Z(n22927) );
XNOR U38213 ( .A(b[7642]), .B(n22928), .Z(c[7642]) );
XNOR U38214 ( .A(a[7642]), .B(c7642), .Z(n22928) );
XOR U38215 ( .A(c7643), .B(n22929), .Z(c7644) );
ANDN U38216 ( .B(n22930), .A(n22931), .Z(n22929) );
XOR U38217 ( .A(c7643), .B(b[7643]), .Z(n22930) );
XNOR U38218 ( .A(b[7643]), .B(n22931), .Z(c[7643]) );
XNOR U38219 ( .A(a[7643]), .B(c7643), .Z(n22931) );
XOR U38220 ( .A(c7644), .B(n22932), .Z(c7645) );
ANDN U38221 ( .B(n22933), .A(n22934), .Z(n22932) );
XOR U38222 ( .A(c7644), .B(b[7644]), .Z(n22933) );
XNOR U38223 ( .A(b[7644]), .B(n22934), .Z(c[7644]) );
XNOR U38224 ( .A(a[7644]), .B(c7644), .Z(n22934) );
XOR U38225 ( .A(c7645), .B(n22935), .Z(c7646) );
ANDN U38226 ( .B(n22936), .A(n22937), .Z(n22935) );
XOR U38227 ( .A(c7645), .B(b[7645]), .Z(n22936) );
XNOR U38228 ( .A(b[7645]), .B(n22937), .Z(c[7645]) );
XNOR U38229 ( .A(a[7645]), .B(c7645), .Z(n22937) );
XOR U38230 ( .A(c7646), .B(n22938), .Z(c7647) );
ANDN U38231 ( .B(n22939), .A(n22940), .Z(n22938) );
XOR U38232 ( .A(c7646), .B(b[7646]), .Z(n22939) );
XNOR U38233 ( .A(b[7646]), .B(n22940), .Z(c[7646]) );
XNOR U38234 ( .A(a[7646]), .B(c7646), .Z(n22940) );
XOR U38235 ( .A(c7647), .B(n22941), .Z(c7648) );
ANDN U38236 ( .B(n22942), .A(n22943), .Z(n22941) );
XOR U38237 ( .A(c7647), .B(b[7647]), .Z(n22942) );
XNOR U38238 ( .A(b[7647]), .B(n22943), .Z(c[7647]) );
XNOR U38239 ( .A(a[7647]), .B(c7647), .Z(n22943) );
XOR U38240 ( .A(c7648), .B(n22944), .Z(c7649) );
ANDN U38241 ( .B(n22945), .A(n22946), .Z(n22944) );
XOR U38242 ( .A(c7648), .B(b[7648]), .Z(n22945) );
XNOR U38243 ( .A(b[7648]), .B(n22946), .Z(c[7648]) );
XNOR U38244 ( .A(a[7648]), .B(c7648), .Z(n22946) );
XOR U38245 ( .A(c7649), .B(n22947), .Z(c7650) );
ANDN U38246 ( .B(n22948), .A(n22949), .Z(n22947) );
XOR U38247 ( .A(c7649), .B(b[7649]), .Z(n22948) );
XNOR U38248 ( .A(b[7649]), .B(n22949), .Z(c[7649]) );
XNOR U38249 ( .A(a[7649]), .B(c7649), .Z(n22949) );
XOR U38250 ( .A(c7650), .B(n22950), .Z(c7651) );
ANDN U38251 ( .B(n22951), .A(n22952), .Z(n22950) );
XOR U38252 ( .A(c7650), .B(b[7650]), .Z(n22951) );
XNOR U38253 ( .A(b[7650]), .B(n22952), .Z(c[7650]) );
XNOR U38254 ( .A(a[7650]), .B(c7650), .Z(n22952) );
XOR U38255 ( .A(c7651), .B(n22953), .Z(c7652) );
ANDN U38256 ( .B(n22954), .A(n22955), .Z(n22953) );
XOR U38257 ( .A(c7651), .B(b[7651]), .Z(n22954) );
XNOR U38258 ( .A(b[7651]), .B(n22955), .Z(c[7651]) );
XNOR U38259 ( .A(a[7651]), .B(c7651), .Z(n22955) );
XOR U38260 ( .A(c7652), .B(n22956), .Z(c7653) );
ANDN U38261 ( .B(n22957), .A(n22958), .Z(n22956) );
XOR U38262 ( .A(c7652), .B(b[7652]), .Z(n22957) );
XNOR U38263 ( .A(b[7652]), .B(n22958), .Z(c[7652]) );
XNOR U38264 ( .A(a[7652]), .B(c7652), .Z(n22958) );
XOR U38265 ( .A(c7653), .B(n22959), .Z(c7654) );
ANDN U38266 ( .B(n22960), .A(n22961), .Z(n22959) );
XOR U38267 ( .A(c7653), .B(b[7653]), .Z(n22960) );
XNOR U38268 ( .A(b[7653]), .B(n22961), .Z(c[7653]) );
XNOR U38269 ( .A(a[7653]), .B(c7653), .Z(n22961) );
XOR U38270 ( .A(c7654), .B(n22962), .Z(c7655) );
ANDN U38271 ( .B(n22963), .A(n22964), .Z(n22962) );
XOR U38272 ( .A(c7654), .B(b[7654]), .Z(n22963) );
XNOR U38273 ( .A(b[7654]), .B(n22964), .Z(c[7654]) );
XNOR U38274 ( .A(a[7654]), .B(c7654), .Z(n22964) );
XOR U38275 ( .A(c7655), .B(n22965), .Z(c7656) );
ANDN U38276 ( .B(n22966), .A(n22967), .Z(n22965) );
XOR U38277 ( .A(c7655), .B(b[7655]), .Z(n22966) );
XNOR U38278 ( .A(b[7655]), .B(n22967), .Z(c[7655]) );
XNOR U38279 ( .A(a[7655]), .B(c7655), .Z(n22967) );
XOR U38280 ( .A(c7656), .B(n22968), .Z(c7657) );
ANDN U38281 ( .B(n22969), .A(n22970), .Z(n22968) );
XOR U38282 ( .A(c7656), .B(b[7656]), .Z(n22969) );
XNOR U38283 ( .A(b[7656]), .B(n22970), .Z(c[7656]) );
XNOR U38284 ( .A(a[7656]), .B(c7656), .Z(n22970) );
XOR U38285 ( .A(c7657), .B(n22971), .Z(c7658) );
ANDN U38286 ( .B(n22972), .A(n22973), .Z(n22971) );
XOR U38287 ( .A(c7657), .B(b[7657]), .Z(n22972) );
XNOR U38288 ( .A(b[7657]), .B(n22973), .Z(c[7657]) );
XNOR U38289 ( .A(a[7657]), .B(c7657), .Z(n22973) );
XOR U38290 ( .A(c7658), .B(n22974), .Z(c7659) );
ANDN U38291 ( .B(n22975), .A(n22976), .Z(n22974) );
XOR U38292 ( .A(c7658), .B(b[7658]), .Z(n22975) );
XNOR U38293 ( .A(b[7658]), .B(n22976), .Z(c[7658]) );
XNOR U38294 ( .A(a[7658]), .B(c7658), .Z(n22976) );
XOR U38295 ( .A(c7659), .B(n22977), .Z(c7660) );
ANDN U38296 ( .B(n22978), .A(n22979), .Z(n22977) );
XOR U38297 ( .A(c7659), .B(b[7659]), .Z(n22978) );
XNOR U38298 ( .A(b[7659]), .B(n22979), .Z(c[7659]) );
XNOR U38299 ( .A(a[7659]), .B(c7659), .Z(n22979) );
XOR U38300 ( .A(c7660), .B(n22980), .Z(c7661) );
ANDN U38301 ( .B(n22981), .A(n22982), .Z(n22980) );
XOR U38302 ( .A(c7660), .B(b[7660]), .Z(n22981) );
XNOR U38303 ( .A(b[7660]), .B(n22982), .Z(c[7660]) );
XNOR U38304 ( .A(a[7660]), .B(c7660), .Z(n22982) );
XOR U38305 ( .A(c7661), .B(n22983), .Z(c7662) );
ANDN U38306 ( .B(n22984), .A(n22985), .Z(n22983) );
XOR U38307 ( .A(c7661), .B(b[7661]), .Z(n22984) );
XNOR U38308 ( .A(b[7661]), .B(n22985), .Z(c[7661]) );
XNOR U38309 ( .A(a[7661]), .B(c7661), .Z(n22985) );
XOR U38310 ( .A(c7662), .B(n22986), .Z(c7663) );
ANDN U38311 ( .B(n22987), .A(n22988), .Z(n22986) );
XOR U38312 ( .A(c7662), .B(b[7662]), .Z(n22987) );
XNOR U38313 ( .A(b[7662]), .B(n22988), .Z(c[7662]) );
XNOR U38314 ( .A(a[7662]), .B(c7662), .Z(n22988) );
XOR U38315 ( .A(c7663), .B(n22989), .Z(c7664) );
ANDN U38316 ( .B(n22990), .A(n22991), .Z(n22989) );
XOR U38317 ( .A(c7663), .B(b[7663]), .Z(n22990) );
XNOR U38318 ( .A(b[7663]), .B(n22991), .Z(c[7663]) );
XNOR U38319 ( .A(a[7663]), .B(c7663), .Z(n22991) );
XOR U38320 ( .A(c7664), .B(n22992), .Z(c7665) );
ANDN U38321 ( .B(n22993), .A(n22994), .Z(n22992) );
XOR U38322 ( .A(c7664), .B(b[7664]), .Z(n22993) );
XNOR U38323 ( .A(b[7664]), .B(n22994), .Z(c[7664]) );
XNOR U38324 ( .A(a[7664]), .B(c7664), .Z(n22994) );
XOR U38325 ( .A(c7665), .B(n22995), .Z(c7666) );
ANDN U38326 ( .B(n22996), .A(n22997), .Z(n22995) );
XOR U38327 ( .A(c7665), .B(b[7665]), .Z(n22996) );
XNOR U38328 ( .A(b[7665]), .B(n22997), .Z(c[7665]) );
XNOR U38329 ( .A(a[7665]), .B(c7665), .Z(n22997) );
XOR U38330 ( .A(c7666), .B(n22998), .Z(c7667) );
ANDN U38331 ( .B(n22999), .A(n23000), .Z(n22998) );
XOR U38332 ( .A(c7666), .B(b[7666]), .Z(n22999) );
XNOR U38333 ( .A(b[7666]), .B(n23000), .Z(c[7666]) );
XNOR U38334 ( .A(a[7666]), .B(c7666), .Z(n23000) );
XOR U38335 ( .A(c7667), .B(n23001), .Z(c7668) );
ANDN U38336 ( .B(n23002), .A(n23003), .Z(n23001) );
XOR U38337 ( .A(c7667), .B(b[7667]), .Z(n23002) );
XNOR U38338 ( .A(b[7667]), .B(n23003), .Z(c[7667]) );
XNOR U38339 ( .A(a[7667]), .B(c7667), .Z(n23003) );
XOR U38340 ( .A(c7668), .B(n23004), .Z(c7669) );
ANDN U38341 ( .B(n23005), .A(n23006), .Z(n23004) );
XOR U38342 ( .A(c7668), .B(b[7668]), .Z(n23005) );
XNOR U38343 ( .A(b[7668]), .B(n23006), .Z(c[7668]) );
XNOR U38344 ( .A(a[7668]), .B(c7668), .Z(n23006) );
XOR U38345 ( .A(c7669), .B(n23007), .Z(c7670) );
ANDN U38346 ( .B(n23008), .A(n23009), .Z(n23007) );
XOR U38347 ( .A(c7669), .B(b[7669]), .Z(n23008) );
XNOR U38348 ( .A(b[7669]), .B(n23009), .Z(c[7669]) );
XNOR U38349 ( .A(a[7669]), .B(c7669), .Z(n23009) );
XOR U38350 ( .A(c7670), .B(n23010), .Z(c7671) );
ANDN U38351 ( .B(n23011), .A(n23012), .Z(n23010) );
XOR U38352 ( .A(c7670), .B(b[7670]), .Z(n23011) );
XNOR U38353 ( .A(b[7670]), .B(n23012), .Z(c[7670]) );
XNOR U38354 ( .A(a[7670]), .B(c7670), .Z(n23012) );
XOR U38355 ( .A(c7671), .B(n23013), .Z(c7672) );
ANDN U38356 ( .B(n23014), .A(n23015), .Z(n23013) );
XOR U38357 ( .A(c7671), .B(b[7671]), .Z(n23014) );
XNOR U38358 ( .A(b[7671]), .B(n23015), .Z(c[7671]) );
XNOR U38359 ( .A(a[7671]), .B(c7671), .Z(n23015) );
XOR U38360 ( .A(c7672), .B(n23016), .Z(c7673) );
ANDN U38361 ( .B(n23017), .A(n23018), .Z(n23016) );
XOR U38362 ( .A(c7672), .B(b[7672]), .Z(n23017) );
XNOR U38363 ( .A(b[7672]), .B(n23018), .Z(c[7672]) );
XNOR U38364 ( .A(a[7672]), .B(c7672), .Z(n23018) );
XOR U38365 ( .A(c7673), .B(n23019), .Z(c7674) );
ANDN U38366 ( .B(n23020), .A(n23021), .Z(n23019) );
XOR U38367 ( .A(c7673), .B(b[7673]), .Z(n23020) );
XNOR U38368 ( .A(b[7673]), .B(n23021), .Z(c[7673]) );
XNOR U38369 ( .A(a[7673]), .B(c7673), .Z(n23021) );
XOR U38370 ( .A(c7674), .B(n23022), .Z(c7675) );
ANDN U38371 ( .B(n23023), .A(n23024), .Z(n23022) );
XOR U38372 ( .A(c7674), .B(b[7674]), .Z(n23023) );
XNOR U38373 ( .A(b[7674]), .B(n23024), .Z(c[7674]) );
XNOR U38374 ( .A(a[7674]), .B(c7674), .Z(n23024) );
XOR U38375 ( .A(c7675), .B(n23025), .Z(c7676) );
ANDN U38376 ( .B(n23026), .A(n23027), .Z(n23025) );
XOR U38377 ( .A(c7675), .B(b[7675]), .Z(n23026) );
XNOR U38378 ( .A(b[7675]), .B(n23027), .Z(c[7675]) );
XNOR U38379 ( .A(a[7675]), .B(c7675), .Z(n23027) );
XOR U38380 ( .A(c7676), .B(n23028), .Z(c7677) );
ANDN U38381 ( .B(n23029), .A(n23030), .Z(n23028) );
XOR U38382 ( .A(c7676), .B(b[7676]), .Z(n23029) );
XNOR U38383 ( .A(b[7676]), .B(n23030), .Z(c[7676]) );
XNOR U38384 ( .A(a[7676]), .B(c7676), .Z(n23030) );
XOR U38385 ( .A(c7677), .B(n23031), .Z(c7678) );
ANDN U38386 ( .B(n23032), .A(n23033), .Z(n23031) );
XOR U38387 ( .A(c7677), .B(b[7677]), .Z(n23032) );
XNOR U38388 ( .A(b[7677]), .B(n23033), .Z(c[7677]) );
XNOR U38389 ( .A(a[7677]), .B(c7677), .Z(n23033) );
XOR U38390 ( .A(c7678), .B(n23034), .Z(c7679) );
ANDN U38391 ( .B(n23035), .A(n23036), .Z(n23034) );
XOR U38392 ( .A(c7678), .B(b[7678]), .Z(n23035) );
XNOR U38393 ( .A(b[7678]), .B(n23036), .Z(c[7678]) );
XNOR U38394 ( .A(a[7678]), .B(c7678), .Z(n23036) );
XOR U38395 ( .A(c7679), .B(n23037), .Z(c7680) );
ANDN U38396 ( .B(n23038), .A(n23039), .Z(n23037) );
XOR U38397 ( .A(c7679), .B(b[7679]), .Z(n23038) );
XNOR U38398 ( .A(b[7679]), .B(n23039), .Z(c[7679]) );
XNOR U38399 ( .A(a[7679]), .B(c7679), .Z(n23039) );
XOR U38400 ( .A(c7680), .B(n23040), .Z(c7681) );
ANDN U38401 ( .B(n23041), .A(n23042), .Z(n23040) );
XOR U38402 ( .A(c7680), .B(b[7680]), .Z(n23041) );
XNOR U38403 ( .A(b[7680]), .B(n23042), .Z(c[7680]) );
XNOR U38404 ( .A(a[7680]), .B(c7680), .Z(n23042) );
XOR U38405 ( .A(c7681), .B(n23043), .Z(c7682) );
ANDN U38406 ( .B(n23044), .A(n23045), .Z(n23043) );
XOR U38407 ( .A(c7681), .B(b[7681]), .Z(n23044) );
XNOR U38408 ( .A(b[7681]), .B(n23045), .Z(c[7681]) );
XNOR U38409 ( .A(a[7681]), .B(c7681), .Z(n23045) );
XOR U38410 ( .A(c7682), .B(n23046), .Z(c7683) );
ANDN U38411 ( .B(n23047), .A(n23048), .Z(n23046) );
XOR U38412 ( .A(c7682), .B(b[7682]), .Z(n23047) );
XNOR U38413 ( .A(b[7682]), .B(n23048), .Z(c[7682]) );
XNOR U38414 ( .A(a[7682]), .B(c7682), .Z(n23048) );
XOR U38415 ( .A(c7683), .B(n23049), .Z(c7684) );
ANDN U38416 ( .B(n23050), .A(n23051), .Z(n23049) );
XOR U38417 ( .A(c7683), .B(b[7683]), .Z(n23050) );
XNOR U38418 ( .A(b[7683]), .B(n23051), .Z(c[7683]) );
XNOR U38419 ( .A(a[7683]), .B(c7683), .Z(n23051) );
XOR U38420 ( .A(c7684), .B(n23052), .Z(c7685) );
ANDN U38421 ( .B(n23053), .A(n23054), .Z(n23052) );
XOR U38422 ( .A(c7684), .B(b[7684]), .Z(n23053) );
XNOR U38423 ( .A(b[7684]), .B(n23054), .Z(c[7684]) );
XNOR U38424 ( .A(a[7684]), .B(c7684), .Z(n23054) );
XOR U38425 ( .A(c7685), .B(n23055), .Z(c7686) );
ANDN U38426 ( .B(n23056), .A(n23057), .Z(n23055) );
XOR U38427 ( .A(c7685), .B(b[7685]), .Z(n23056) );
XNOR U38428 ( .A(b[7685]), .B(n23057), .Z(c[7685]) );
XNOR U38429 ( .A(a[7685]), .B(c7685), .Z(n23057) );
XOR U38430 ( .A(c7686), .B(n23058), .Z(c7687) );
ANDN U38431 ( .B(n23059), .A(n23060), .Z(n23058) );
XOR U38432 ( .A(c7686), .B(b[7686]), .Z(n23059) );
XNOR U38433 ( .A(b[7686]), .B(n23060), .Z(c[7686]) );
XNOR U38434 ( .A(a[7686]), .B(c7686), .Z(n23060) );
XOR U38435 ( .A(c7687), .B(n23061), .Z(c7688) );
ANDN U38436 ( .B(n23062), .A(n23063), .Z(n23061) );
XOR U38437 ( .A(c7687), .B(b[7687]), .Z(n23062) );
XNOR U38438 ( .A(b[7687]), .B(n23063), .Z(c[7687]) );
XNOR U38439 ( .A(a[7687]), .B(c7687), .Z(n23063) );
XOR U38440 ( .A(c7688), .B(n23064), .Z(c7689) );
ANDN U38441 ( .B(n23065), .A(n23066), .Z(n23064) );
XOR U38442 ( .A(c7688), .B(b[7688]), .Z(n23065) );
XNOR U38443 ( .A(b[7688]), .B(n23066), .Z(c[7688]) );
XNOR U38444 ( .A(a[7688]), .B(c7688), .Z(n23066) );
XOR U38445 ( .A(c7689), .B(n23067), .Z(c7690) );
ANDN U38446 ( .B(n23068), .A(n23069), .Z(n23067) );
XOR U38447 ( .A(c7689), .B(b[7689]), .Z(n23068) );
XNOR U38448 ( .A(b[7689]), .B(n23069), .Z(c[7689]) );
XNOR U38449 ( .A(a[7689]), .B(c7689), .Z(n23069) );
XOR U38450 ( .A(c7690), .B(n23070), .Z(c7691) );
ANDN U38451 ( .B(n23071), .A(n23072), .Z(n23070) );
XOR U38452 ( .A(c7690), .B(b[7690]), .Z(n23071) );
XNOR U38453 ( .A(b[7690]), .B(n23072), .Z(c[7690]) );
XNOR U38454 ( .A(a[7690]), .B(c7690), .Z(n23072) );
XOR U38455 ( .A(c7691), .B(n23073), .Z(c7692) );
ANDN U38456 ( .B(n23074), .A(n23075), .Z(n23073) );
XOR U38457 ( .A(c7691), .B(b[7691]), .Z(n23074) );
XNOR U38458 ( .A(b[7691]), .B(n23075), .Z(c[7691]) );
XNOR U38459 ( .A(a[7691]), .B(c7691), .Z(n23075) );
XOR U38460 ( .A(c7692), .B(n23076), .Z(c7693) );
ANDN U38461 ( .B(n23077), .A(n23078), .Z(n23076) );
XOR U38462 ( .A(c7692), .B(b[7692]), .Z(n23077) );
XNOR U38463 ( .A(b[7692]), .B(n23078), .Z(c[7692]) );
XNOR U38464 ( .A(a[7692]), .B(c7692), .Z(n23078) );
XOR U38465 ( .A(c7693), .B(n23079), .Z(c7694) );
ANDN U38466 ( .B(n23080), .A(n23081), .Z(n23079) );
XOR U38467 ( .A(c7693), .B(b[7693]), .Z(n23080) );
XNOR U38468 ( .A(b[7693]), .B(n23081), .Z(c[7693]) );
XNOR U38469 ( .A(a[7693]), .B(c7693), .Z(n23081) );
XOR U38470 ( .A(c7694), .B(n23082), .Z(c7695) );
ANDN U38471 ( .B(n23083), .A(n23084), .Z(n23082) );
XOR U38472 ( .A(c7694), .B(b[7694]), .Z(n23083) );
XNOR U38473 ( .A(b[7694]), .B(n23084), .Z(c[7694]) );
XNOR U38474 ( .A(a[7694]), .B(c7694), .Z(n23084) );
XOR U38475 ( .A(c7695), .B(n23085), .Z(c7696) );
ANDN U38476 ( .B(n23086), .A(n23087), .Z(n23085) );
XOR U38477 ( .A(c7695), .B(b[7695]), .Z(n23086) );
XNOR U38478 ( .A(b[7695]), .B(n23087), .Z(c[7695]) );
XNOR U38479 ( .A(a[7695]), .B(c7695), .Z(n23087) );
XOR U38480 ( .A(c7696), .B(n23088), .Z(c7697) );
ANDN U38481 ( .B(n23089), .A(n23090), .Z(n23088) );
XOR U38482 ( .A(c7696), .B(b[7696]), .Z(n23089) );
XNOR U38483 ( .A(b[7696]), .B(n23090), .Z(c[7696]) );
XNOR U38484 ( .A(a[7696]), .B(c7696), .Z(n23090) );
XOR U38485 ( .A(c7697), .B(n23091), .Z(c7698) );
ANDN U38486 ( .B(n23092), .A(n23093), .Z(n23091) );
XOR U38487 ( .A(c7697), .B(b[7697]), .Z(n23092) );
XNOR U38488 ( .A(b[7697]), .B(n23093), .Z(c[7697]) );
XNOR U38489 ( .A(a[7697]), .B(c7697), .Z(n23093) );
XOR U38490 ( .A(c7698), .B(n23094), .Z(c7699) );
ANDN U38491 ( .B(n23095), .A(n23096), .Z(n23094) );
XOR U38492 ( .A(c7698), .B(b[7698]), .Z(n23095) );
XNOR U38493 ( .A(b[7698]), .B(n23096), .Z(c[7698]) );
XNOR U38494 ( .A(a[7698]), .B(c7698), .Z(n23096) );
XOR U38495 ( .A(c7699), .B(n23097), .Z(c7700) );
ANDN U38496 ( .B(n23098), .A(n23099), .Z(n23097) );
XOR U38497 ( .A(c7699), .B(b[7699]), .Z(n23098) );
XNOR U38498 ( .A(b[7699]), .B(n23099), .Z(c[7699]) );
XNOR U38499 ( .A(a[7699]), .B(c7699), .Z(n23099) );
XOR U38500 ( .A(c7700), .B(n23100), .Z(c7701) );
ANDN U38501 ( .B(n23101), .A(n23102), .Z(n23100) );
XOR U38502 ( .A(c7700), .B(b[7700]), .Z(n23101) );
XNOR U38503 ( .A(b[7700]), .B(n23102), .Z(c[7700]) );
XNOR U38504 ( .A(a[7700]), .B(c7700), .Z(n23102) );
XOR U38505 ( .A(c7701), .B(n23103), .Z(c7702) );
ANDN U38506 ( .B(n23104), .A(n23105), .Z(n23103) );
XOR U38507 ( .A(c7701), .B(b[7701]), .Z(n23104) );
XNOR U38508 ( .A(b[7701]), .B(n23105), .Z(c[7701]) );
XNOR U38509 ( .A(a[7701]), .B(c7701), .Z(n23105) );
XOR U38510 ( .A(c7702), .B(n23106), .Z(c7703) );
ANDN U38511 ( .B(n23107), .A(n23108), .Z(n23106) );
XOR U38512 ( .A(c7702), .B(b[7702]), .Z(n23107) );
XNOR U38513 ( .A(b[7702]), .B(n23108), .Z(c[7702]) );
XNOR U38514 ( .A(a[7702]), .B(c7702), .Z(n23108) );
XOR U38515 ( .A(c7703), .B(n23109), .Z(c7704) );
ANDN U38516 ( .B(n23110), .A(n23111), .Z(n23109) );
XOR U38517 ( .A(c7703), .B(b[7703]), .Z(n23110) );
XNOR U38518 ( .A(b[7703]), .B(n23111), .Z(c[7703]) );
XNOR U38519 ( .A(a[7703]), .B(c7703), .Z(n23111) );
XOR U38520 ( .A(c7704), .B(n23112), .Z(c7705) );
ANDN U38521 ( .B(n23113), .A(n23114), .Z(n23112) );
XOR U38522 ( .A(c7704), .B(b[7704]), .Z(n23113) );
XNOR U38523 ( .A(b[7704]), .B(n23114), .Z(c[7704]) );
XNOR U38524 ( .A(a[7704]), .B(c7704), .Z(n23114) );
XOR U38525 ( .A(c7705), .B(n23115), .Z(c7706) );
ANDN U38526 ( .B(n23116), .A(n23117), .Z(n23115) );
XOR U38527 ( .A(c7705), .B(b[7705]), .Z(n23116) );
XNOR U38528 ( .A(b[7705]), .B(n23117), .Z(c[7705]) );
XNOR U38529 ( .A(a[7705]), .B(c7705), .Z(n23117) );
XOR U38530 ( .A(c7706), .B(n23118), .Z(c7707) );
ANDN U38531 ( .B(n23119), .A(n23120), .Z(n23118) );
XOR U38532 ( .A(c7706), .B(b[7706]), .Z(n23119) );
XNOR U38533 ( .A(b[7706]), .B(n23120), .Z(c[7706]) );
XNOR U38534 ( .A(a[7706]), .B(c7706), .Z(n23120) );
XOR U38535 ( .A(c7707), .B(n23121), .Z(c7708) );
ANDN U38536 ( .B(n23122), .A(n23123), .Z(n23121) );
XOR U38537 ( .A(c7707), .B(b[7707]), .Z(n23122) );
XNOR U38538 ( .A(b[7707]), .B(n23123), .Z(c[7707]) );
XNOR U38539 ( .A(a[7707]), .B(c7707), .Z(n23123) );
XOR U38540 ( .A(c7708), .B(n23124), .Z(c7709) );
ANDN U38541 ( .B(n23125), .A(n23126), .Z(n23124) );
XOR U38542 ( .A(c7708), .B(b[7708]), .Z(n23125) );
XNOR U38543 ( .A(b[7708]), .B(n23126), .Z(c[7708]) );
XNOR U38544 ( .A(a[7708]), .B(c7708), .Z(n23126) );
XOR U38545 ( .A(c7709), .B(n23127), .Z(c7710) );
ANDN U38546 ( .B(n23128), .A(n23129), .Z(n23127) );
XOR U38547 ( .A(c7709), .B(b[7709]), .Z(n23128) );
XNOR U38548 ( .A(b[7709]), .B(n23129), .Z(c[7709]) );
XNOR U38549 ( .A(a[7709]), .B(c7709), .Z(n23129) );
XOR U38550 ( .A(c7710), .B(n23130), .Z(c7711) );
ANDN U38551 ( .B(n23131), .A(n23132), .Z(n23130) );
XOR U38552 ( .A(c7710), .B(b[7710]), .Z(n23131) );
XNOR U38553 ( .A(b[7710]), .B(n23132), .Z(c[7710]) );
XNOR U38554 ( .A(a[7710]), .B(c7710), .Z(n23132) );
XOR U38555 ( .A(c7711), .B(n23133), .Z(c7712) );
ANDN U38556 ( .B(n23134), .A(n23135), .Z(n23133) );
XOR U38557 ( .A(c7711), .B(b[7711]), .Z(n23134) );
XNOR U38558 ( .A(b[7711]), .B(n23135), .Z(c[7711]) );
XNOR U38559 ( .A(a[7711]), .B(c7711), .Z(n23135) );
XOR U38560 ( .A(c7712), .B(n23136), .Z(c7713) );
ANDN U38561 ( .B(n23137), .A(n23138), .Z(n23136) );
XOR U38562 ( .A(c7712), .B(b[7712]), .Z(n23137) );
XNOR U38563 ( .A(b[7712]), .B(n23138), .Z(c[7712]) );
XNOR U38564 ( .A(a[7712]), .B(c7712), .Z(n23138) );
XOR U38565 ( .A(c7713), .B(n23139), .Z(c7714) );
ANDN U38566 ( .B(n23140), .A(n23141), .Z(n23139) );
XOR U38567 ( .A(c7713), .B(b[7713]), .Z(n23140) );
XNOR U38568 ( .A(b[7713]), .B(n23141), .Z(c[7713]) );
XNOR U38569 ( .A(a[7713]), .B(c7713), .Z(n23141) );
XOR U38570 ( .A(c7714), .B(n23142), .Z(c7715) );
ANDN U38571 ( .B(n23143), .A(n23144), .Z(n23142) );
XOR U38572 ( .A(c7714), .B(b[7714]), .Z(n23143) );
XNOR U38573 ( .A(b[7714]), .B(n23144), .Z(c[7714]) );
XNOR U38574 ( .A(a[7714]), .B(c7714), .Z(n23144) );
XOR U38575 ( .A(c7715), .B(n23145), .Z(c7716) );
ANDN U38576 ( .B(n23146), .A(n23147), .Z(n23145) );
XOR U38577 ( .A(c7715), .B(b[7715]), .Z(n23146) );
XNOR U38578 ( .A(b[7715]), .B(n23147), .Z(c[7715]) );
XNOR U38579 ( .A(a[7715]), .B(c7715), .Z(n23147) );
XOR U38580 ( .A(c7716), .B(n23148), .Z(c7717) );
ANDN U38581 ( .B(n23149), .A(n23150), .Z(n23148) );
XOR U38582 ( .A(c7716), .B(b[7716]), .Z(n23149) );
XNOR U38583 ( .A(b[7716]), .B(n23150), .Z(c[7716]) );
XNOR U38584 ( .A(a[7716]), .B(c7716), .Z(n23150) );
XOR U38585 ( .A(c7717), .B(n23151), .Z(c7718) );
ANDN U38586 ( .B(n23152), .A(n23153), .Z(n23151) );
XOR U38587 ( .A(c7717), .B(b[7717]), .Z(n23152) );
XNOR U38588 ( .A(b[7717]), .B(n23153), .Z(c[7717]) );
XNOR U38589 ( .A(a[7717]), .B(c7717), .Z(n23153) );
XOR U38590 ( .A(c7718), .B(n23154), .Z(c7719) );
ANDN U38591 ( .B(n23155), .A(n23156), .Z(n23154) );
XOR U38592 ( .A(c7718), .B(b[7718]), .Z(n23155) );
XNOR U38593 ( .A(b[7718]), .B(n23156), .Z(c[7718]) );
XNOR U38594 ( .A(a[7718]), .B(c7718), .Z(n23156) );
XOR U38595 ( .A(c7719), .B(n23157), .Z(c7720) );
ANDN U38596 ( .B(n23158), .A(n23159), .Z(n23157) );
XOR U38597 ( .A(c7719), .B(b[7719]), .Z(n23158) );
XNOR U38598 ( .A(b[7719]), .B(n23159), .Z(c[7719]) );
XNOR U38599 ( .A(a[7719]), .B(c7719), .Z(n23159) );
XOR U38600 ( .A(c7720), .B(n23160), .Z(c7721) );
ANDN U38601 ( .B(n23161), .A(n23162), .Z(n23160) );
XOR U38602 ( .A(c7720), .B(b[7720]), .Z(n23161) );
XNOR U38603 ( .A(b[7720]), .B(n23162), .Z(c[7720]) );
XNOR U38604 ( .A(a[7720]), .B(c7720), .Z(n23162) );
XOR U38605 ( .A(c7721), .B(n23163), .Z(c7722) );
ANDN U38606 ( .B(n23164), .A(n23165), .Z(n23163) );
XOR U38607 ( .A(c7721), .B(b[7721]), .Z(n23164) );
XNOR U38608 ( .A(b[7721]), .B(n23165), .Z(c[7721]) );
XNOR U38609 ( .A(a[7721]), .B(c7721), .Z(n23165) );
XOR U38610 ( .A(c7722), .B(n23166), .Z(c7723) );
ANDN U38611 ( .B(n23167), .A(n23168), .Z(n23166) );
XOR U38612 ( .A(c7722), .B(b[7722]), .Z(n23167) );
XNOR U38613 ( .A(b[7722]), .B(n23168), .Z(c[7722]) );
XNOR U38614 ( .A(a[7722]), .B(c7722), .Z(n23168) );
XOR U38615 ( .A(c7723), .B(n23169), .Z(c7724) );
ANDN U38616 ( .B(n23170), .A(n23171), .Z(n23169) );
XOR U38617 ( .A(c7723), .B(b[7723]), .Z(n23170) );
XNOR U38618 ( .A(b[7723]), .B(n23171), .Z(c[7723]) );
XNOR U38619 ( .A(a[7723]), .B(c7723), .Z(n23171) );
XOR U38620 ( .A(c7724), .B(n23172), .Z(c7725) );
ANDN U38621 ( .B(n23173), .A(n23174), .Z(n23172) );
XOR U38622 ( .A(c7724), .B(b[7724]), .Z(n23173) );
XNOR U38623 ( .A(b[7724]), .B(n23174), .Z(c[7724]) );
XNOR U38624 ( .A(a[7724]), .B(c7724), .Z(n23174) );
XOR U38625 ( .A(c7725), .B(n23175), .Z(c7726) );
ANDN U38626 ( .B(n23176), .A(n23177), .Z(n23175) );
XOR U38627 ( .A(c7725), .B(b[7725]), .Z(n23176) );
XNOR U38628 ( .A(b[7725]), .B(n23177), .Z(c[7725]) );
XNOR U38629 ( .A(a[7725]), .B(c7725), .Z(n23177) );
XOR U38630 ( .A(c7726), .B(n23178), .Z(c7727) );
ANDN U38631 ( .B(n23179), .A(n23180), .Z(n23178) );
XOR U38632 ( .A(c7726), .B(b[7726]), .Z(n23179) );
XNOR U38633 ( .A(b[7726]), .B(n23180), .Z(c[7726]) );
XNOR U38634 ( .A(a[7726]), .B(c7726), .Z(n23180) );
XOR U38635 ( .A(c7727), .B(n23181), .Z(c7728) );
ANDN U38636 ( .B(n23182), .A(n23183), .Z(n23181) );
XOR U38637 ( .A(c7727), .B(b[7727]), .Z(n23182) );
XNOR U38638 ( .A(b[7727]), .B(n23183), .Z(c[7727]) );
XNOR U38639 ( .A(a[7727]), .B(c7727), .Z(n23183) );
XOR U38640 ( .A(c7728), .B(n23184), .Z(c7729) );
ANDN U38641 ( .B(n23185), .A(n23186), .Z(n23184) );
XOR U38642 ( .A(c7728), .B(b[7728]), .Z(n23185) );
XNOR U38643 ( .A(b[7728]), .B(n23186), .Z(c[7728]) );
XNOR U38644 ( .A(a[7728]), .B(c7728), .Z(n23186) );
XOR U38645 ( .A(c7729), .B(n23187), .Z(c7730) );
ANDN U38646 ( .B(n23188), .A(n23189), .Z(n23187) );
XOR U38647 ( .A(c7729), .B(b[7729]), .Z(n23188) );
XNOR U38648 ( .A(b[7729]), .B(n23189), .Z(c[7729]) );
XNOR U38649 ( .A(a[7729]), .B(c7729), .Z(n23189) );
XOR U38650 ( .A(c7730), .B(n23190), .Z(c7731) );
ANDN U38651 ( .B(n23191), .A(n23192), .Z(n23190) );
XOR U38652 ( .A(c7730), .B(b[7730]), .Z(n23191) );
XNOR U38653 ( .A(b[7730]), .B(n23192), .Z(c[7730]) );
XNOR U38654 ( .A(a[7730]), .B(c7730), .Z(n23192) );
XOR U38655 ( .A(c7731), .B(n23193), .Z(c7732) );
ANDN U38656 ( .B(n23194), .A(n23195), .Z(n23193) );
XOR U38657 ( .A(c7731), .B(b[7731]), .Z(n23194) );
XNOR U38658 ( .A(b[7731]), .B(n23195), .Z(c[7731]) );
XNOR U38659 ( .A(a[7731]), .B(c7731), .Z(n23195) );
XOR U38660 ( .A(c7732), .B(n23196), .Z(c7733) );
ANDN U38661 ( .B(n23197), .A(n23198), .Z(n23196) );
XOR U38662 ( .A(c7732), .B(b[7732]), .Z(n23197) );
XNOR U38663 ( .A(b[7732]), .B(n23198), .Z(c[7732]) );
XNOR U38664 ( .A(a[7732]), .B(c7732), .Z(n23198) );
XOR U38665 ( .A(c7733), .B(n23199), .Z(c7734) );
ANDN U38666 ( .B(n23200), .A(n23201), .Z(n23199) );
XOR U38667 ( .A(c7733), .B(b[7733]), .Z(n23200) );
XNOR U38668 ( .A(b[7733]), .B(n23201), .Z(c[7733]) );
XNOR U38669 ( .A(a[7733]), .B(c7733), .Z(n23201) );
XOR U38670 ( .A(c7734), .B(n23202), .Z(c7735) );
ANDN U38671 ( .B(n23203), .A(n23204), .Z(n23202) );
XOR U38672 ( .A(c7734), .B(b[7734]), .Z(n23203) );
XNOR U38673 ( .A(b[7734]), .B(n23204), .Z(c[7734]) );
XNOR U38674 ( .A(a[7734]), .B(c7734), .Z(n23204) );
XOR U38675 ( .A(c7735), .B(n23205), .Z(c7736) );
ANDN U38676 ( .B(n23206), .A(n23207), .Z(n23205) );
XOR U38677 ( .A(c7735), .B(b[7735]), .Z(n23206) );
XNOR U38678 ( .A(b[7735]), .B(n23207), .Z(c[7735]) );
XNOR U38679 ( .A(a[7735]), .B(c7735), .Z(n23207) );
XOR U38680 ( .A(c7736), .B(n23208), .Z(c7737) );
ANDN U38681 ( .B(n23209), .A(n23210), .Z(n23208) );
XOR U38682 ( .A(c7736), .B(b[7736]), .Z(n23209) );
XNOR U38683 ( .A(b[7736]), .B(n23210), .Z(c[7736]) );
XNOR U38684 ( .A(a[7736]), .B(c7736), .Z(n23210) );
XOR U38685 ( .A(c7737), .B(n23211), .Z(c7738) );
ANDN U38686 ( .B(n23212), .A(n23213), .Z(n23211) );
XOR U38687 ( .A(c7737), .B(b[7737]), .Z(n23212) );
XNOR U38688 ( .A(b[7737]), .B(n23213), .Z(c[7737]) );
XNOR U38689 ( .A(a[7737]), .B(c7737), .Z(n23213) );
XOR U38690 ( .A(c7738), .B(n23214), .Z(c7739) );
ANDN U38691 ( .B(n23215), .A(n23216), .Z(n23214) );
XOR U38692 ( .A(c7738), .B(b[7738]), .Z(n23215) );
XNOR U38693 ( .A(b[7738]), .B(n23216), .Z(c[7738]) );
XNOR U38694 ( .A(a[7738]), .B(c7738), .Z(n23216) );
XOR U38695 ( .A(c7739), .B(n23217), .Z(c7740) );
ANDN U38696 ( .B(n23218), .A(n23219), .Z(n23217) );
XOR U38697 ( .A(c7739), .B(b[7739]), .Z(n23218) );
XNOR U38698 ( .A(b[7739]), .B(n23219), .Z(c[7739]) );
XNOR U38699 ( .A(a[7739]), .B(c7739), .Z(n23219) );
XOR U38700 ( .A(c7740), .B(n23220), .Z(c7741) );
ANDN U38701 ( .B(n23221), .A(n23222), .Z(n23220) );
XOR U38702 ( .A(c7740), .B(b[7740]), .Z(n23221) );
XNOR U38703 ( .A(b[7740]), .B(n23222), .Z(c[7740]) );
XNOR U38704 ( .A(a[7740]), .B(c7740), .Z(n23222) );
XOR U38705 ( .A(c7741), .B(n23223), .Z(c7742) );
ANDN U38706 ( .B(n23224), .A(n23225), .Z(n23223) );
XOR U38707 ( .A(c7741), .B(b[7741]), .Z(n23224) );
XNOR U38708 ( .A(b[7741]), .B(n23225), .Z(c[7741]) );
XNOR U38709 ( .A(a[7741]), .B(c7741), .Z(n23225) );
XOR U38710 ( .A(c7742), .B(n23226), .Z(c7743) );
ANDN U38711 ( .B(n23227), .A(n23228), .Z(n23226) );
XOR U38712 ( .A(c7742), .B(b[7742]), .Z(n23227) );
XNOR U38713 ( .A(b[7742]), .B(n23228), .Z(c[7742]) );
XNOR U38714 ( .A(a[7742]), .B(c7742), .Z(n23228) );
XOR U38715 ( .A(c7743), .B(n23229), .Z(c7744) );
ANDN U38716 ( .B(n23230), .A(n23231), .Z(n23229) );
XOR U38717 ( .A(c7743), .B(b[7743]), .Z(n23230) );
XNOR U38718 ( .A(b[7743]), .B(n23231), .Z(c[7743]) );
XNOR U38719 ( .A(a[7743]), .B(c7743), .Z(n23231) );
XOR U38720 ( .A(c7744), .B(n23232), .Z(c7745) );
ANDN U38721 ( .B(n23233), .A(n23234), .Z(n23232) );
XOR U38722 ( .A(c7744), .B(b[7744]), .Z(n23233) );
XNOR U38723 ( .A(b[7744]), .B(n23234), .Z(c[7744]) );
XNOR U38724 ( .A(a[7744]), .B(c7744), .Z(n23234) );
XOR U38725 ( .A(c7745), .B(n23235), .Z(c7746) );
ANDN U38726 ( .B(n23236), .A(n23237), .Z(n23235) );
XOR U38727 ( .A(c7745), .B(b[7745]), .Z(n23236) );
XNOR U38728 ( .A(b[7745]), .B(n23237), .Z(c[7745]) );
XNOR U38729 ( .A(a[7745]), .B(c7745), .Z(n23237) );
XOR U38730 ( .A(c7746), .B(n23238), .Z(c7747) );
ANDN U38731 ( .B(n23239), .A(n23240), .Z(n23238) );
XOR U38732 ( .A(c7746), .B(b[7746]), .Z(n23239) );
XNOR U38733 ( .A(b[7746]), .B(n23240), .Z(c[7746]) );
XNOR U38734 ( .A(a[7746]), .B(c7746), .Z(n23240) );
XOR U38735 ( .A(c7747), .B(n23241), .Z(c7748) );
ANDN U38736 ( .B(n23242), .A(n23243), .Z(n23241) );
XOR U38737 ( .A(c7747), .B(b[7747]), .Z(n23242) );
XNOR U38738 ( .A(b[7747]), .B(n23243), .Z(c[7747]) );
XNOR U38739 ( .A(a[7747]), .B(c7747), .Z(n23243) );
XOR U38740 ( .A(c7748), .B(n23244), .Z(c7749) );
ANDN U38741 ( .B(n23245), .A(n23246), .Z(n23244) );
XOR U38742 ( .A(c7748), .B(b[7748]), .Z(n23245) );
XNOR U38743 ( .A(b[7748]), .B(n23246), .Z(c[7748]) );
XNOR U38744 ( .A(a[7748]), .B(c7748), .Z(n23246) );
XOR U38745 ( .A(c7749), .B(n23247), .Z(c7750) );
ANDN U38746 ( .B(n23248), .A(n23249), .Z(n23247) );
XOR U38747 ( .A(c7749), .B(b[7749]), .Z(n23248) );
XNOR U38748 ( .A(b[7749]), .B(n23249), .Z(c[7749]) );
XNOR U38749 ( .A(a[7749]), .B(c7749), .Z(n23249) );
XOR U38750 ( .A(c7750), .B(n23250), .Z(c7751) );
ANDN U38751 ( .B(n23251), .A(n23252), .Z(n23250) );
XOR U38752 ( .A(c7750), .B(b[7750]), .Z(n23251) );
XNOR U38753 ( .A(b[7750]), .B(n23252), .Z(c[7750]) );
XNOR U38754 ( .A(a[7750]), .B(c7750), .Z(n23252) );
XOR U38755 ( .A(c7751), .B(n23253), .Z(c7752) );
ANDN U38756 ( .B(n23254), .A(n23255), .Z(n23253) );
XOR U38757 ( .A(c7751), .B(b[7751]), .Z(n23254) );
XNOR U38758 ( .A(b[7751]), .B(n23255), .Z(c[7751]) );
XNOR U38759 ( .A(a[7751]), .B(c7751), .Z(n23255) );
XOR U38760 ( .A(c7752), .B(n23256), .Z(c7753) );
ANDN U38761 ( .B(n23257), .A(n23258), .Z(n23256) );
XOR U38762 ( .A(c7752), .B(b[7752]), .Z(n23257) );
XNOR U38763 ( .A(b[7752]), .B(n23258), .Z(c[7752]) );
XNOR U38764 ( .A(a[7752]), .B(c7752), .Z(n23258) );
XOR U38765 ( .A(c7753), .B(n23259), .Z(c7754) );
ANDN U38766 ( .B(n23260), .A(n23261), .Z(n23259) );
XOR U38767 ( .A(c7753), .B(b[7753]), .Z(n23260) );
XNOR U38768 ( .A(b[7753]), .B(n23261), .Z(c[7753]) );
XNOR U38769 ( .A(a[7753]), .B(c7753), .Z(n23261) );
XOR U38770 ( .A(c7754), .B(n23262), .Z(c7755) );
ANDN U38771 ( .B(n23263), .A(n23264), .Z(n23262) );
XOR U38772 ( .A(c7754), .B(b[7754]), .Z(n23263) );
XNOR U38773 ( .A(b[7754]), .B(n23264), .Z(c[7754]) );
XNOR U38774 ( .A(a[7754]), .B(c7754), .Z(n23264) );
XOR U38775 ( .A(c7755), .B(n23265), .Z(c7756) );
ANDN U38776 ( .B(n23266), .A(n23267), .Z(n23265) );
XOR U38777 ( .A(c7755), .B(b[7755]), .Z(n23266) );
XNOR U38778 ( .A(b[7755]), .B(n23267), .Z(c[7755]) );
XNOR U38779 ( .A(a[7755]), .B(c7755), .Z(n23267) );
XOR U38780 ( .A(c7756), .B(n23268), .Z(c7757) );
ANDN U38781 ( .B(n23269), .A(n23270), .Z(n23268) );
XOR U38782 ( .A(c7756), .B(b[7756]), .Z(n23269) );
XNOR U38783 ( .A(b[7756]), .B(n23270), .Z(c[7756]) );
XNOR U38784 ( .A(a[7756]), .B(c7756), .Z(n23270) );
XOR U38785 ( .A(c7757), .B(n23271), .Z(c7758) );
ANDN U38786 ( .B(n23272), .A(n23273), .Z(n23271) );
XOR U38787 ( .A(c7757), .B(b[7757]), .Z(n23272) );
XNOR U38788 ( .A(b[7757]), .B(n23273), .Z(c[7757]) );
XNOR U38789 ( .A(a[7757]), .B(c7757), .Z(n23273) );
XOR U38790 ( .A(c7758), .B(n23274), .Z(c7759) );
ANDN U38791 ( .B(n23275), .A(n23276), .Z(n23274) );
XOR U38792 ( .A(c7758), .B(b[7758]), .Z(n23275) );
XNOR U38793 ( .A(b[7758]), .B(n23276), .Z(c[7758]) );
XNOR U38794 ( .A(a[7758]), .B(c7758), .Z(n23276) );
XOR U38795 ( .A(c7759), .B(n23277), .Z(c7760) );
ANDN U38796 ( .B(n23278), .A(n23279), .Z(n23277) );
XOR U38797 ( .A(c7759), .B(b[7759]), .Z(n23278) );
XNOR U38798 ( .A(b[7759]), .B(n23279), .Z(c[7759]) );
XNOR U38799 ( .A(a[7759]), .B(c7759), .Z(n23279) );
XOR U38800 ( .A(c7760), .B(n23280), .Z(c7761) );
ANDN U38801 ( .B(n23281), .A(n23282), .Z(n23280) );
XOR U38802 ( .A(c7760), .B(b[7760]), .Z(n23281) );
XNOR U38803 ( .A(b[7760]), .B(n23282), .Z(c[7760]) );
XNOR U38804 ( .A(a[7760]), .B(c7760), .Z(n23282) );
XOR U38805 ( .A(c7761), .B(n23283), .Z(c7762) );
ANDN U38806 ( .B(n23284), .A(n23285), .Z(n23283) );
XOR U38807 ( .A(c7761), .B(b[7761]), .Z(n23284) );
XNOR U38808 ( .A(b[7761]), .B(n23285), .Z(c[7761]) );
XNOR U38809 ( .A(a[7761]), .B(c7761), .Z(n23285) );
XOR U38810 ( .A(c7762), .B(n23286), .Z(c7763) );
ANDN U38811 ( .B(n23287), .A(n23288), .Z(n23286) );
XOR U38812 ( .A(c7762), .B(b[7762]), .Z(n23287) );
XNOR U38813 ( .A(b[7762]), .B(n23288), .Z(c[7762]) );
XNOR U38814 ( .A(a[7762]), .B(c7762), .Z(n23288) );
XOR U38815 ( .A(c7763), .B(n23289), .Z(c7764) );
ANDN U38816 ( .B(n23290), .A(n23291), .Z(n23289) );
XOR U38817 ( .A(c7763), .B(b[7763]), .Z(n23290) );
XNOR U38818 ( .A(b[7763]), .B(n23291), .Z(c[7763]) );
XNOR U38819 ( .A(a[7763]), .B(c7763), .Z(n23291) );
XOR U38820 ( .A(c7764), .B(n23292), .Z(c7765) );
ANDN U38821 ( .B(n23293), .A(n23294), .Z(n23292) );
XOR U38822 ( .A(c7764), .B(b[7764]), .Z(n23293) );
XNOR U38823 ( .A(b[7764]), .B(n23294), .Z(c[7764]) );
XNOR U38824 ( .A(a[7764]), .B(c7764), .Z(n23294) );
XOR U38825 ( .A(c7765), .B(n23295), .Z(c7766) );
ANDN U38826 ( .B(n23296), .A(n23297), .Z(n23295) );
XOR U38827 ( .A(c7765), .B(b[7765]), .Z(n23296) );
XNOR U38828 ( .A(b[7765]), .B(n23297), .Z(c[7765]) );
XNOR U38829 ( .A(a[7765]), .B(c7765), .Z(n23297) );
XOR U38830 ( .A(c7766), .B(n23298), .Z(c7767) );
ANDN U38831 ( .B(n23299), .A(n23300), .Z(n23298) );
XOR U38832 ( .A(c7766), .B(b[7766]), .Z(n23299) );
XNOR U38833 ( .A(b[7766]), .B(n23300), .Z(c[7766]) );
XNOR U38834 ( .A(a[7766]), .B(c7766), .Z(n23300) );
XOR U38835 ( .A(c7767), .B(n23301), .Z(c7768) );
ANDN U38836 ( .B(n23302), .A(n23303), .Z(n23301) );
XOR U38837 ( .A(c7767), .B(b[7767]), .Z(n23302) );
XNOR U38838 ( .A(b[7767]), .B(n23303), .Z(c[7767]) );
XNOR U38839 ( .A(a[7767]), .B(c7767), .Z(n23303) );
XOR U38840 ( .A(c7768), .B(n23304), .Z(c7769) );
ANDN U38841 ( .B(n23305), .A(n23306), .Z(n23304) );
XOR U38842 ( .A(c7768), .B(b[7768]), .Z(n23305) );
XNOR U38843 ( .A(b[7768]), .B(n23306), .Z(c[7768]) );
XNOR U38844 ( .A(a[7768]), .B(c7768), .Z(n23306) );
XOR U38845 ( .A(c7769), .B(n23307), .Z(c7770) );
ANDN U38846 ( .B(n23308), .A(n23309), .Z(n23307) );
XOR U38847 ( .A(c7769), .B(b[7769]), .Z(n23308) );
XNOR U38848 ( .A(b[7769]), .B(n23309), .Z(c[7769]) );
XNOR U38849 ( .A(a[7769]), .B(c7769), .Z(n23309) );
XOR U38850 ( .A(c7770), .B(n23310), .Z(c7771) );
ANDN U38851 ( .B(n23311), .A(n23312), .Z(n23310) );
XOR U38852 ( .A(c7770), .B(b[7770]), .Z(n23311) );
XNOR U38853 ( .A(b[7770]), .B(n23312), .Z(c[7770]) );
XNOR U38854 ( .A(a[7770]), .B(c7770), .Z(n23312) );
XOR U38855 ( .A(c7771), .B(n23313), .Z(c7772) );
ANDN U38856 ( .B(n23314), .A(n23315), .Z(n23313) );
XOR U38857 ( .A(c7771), .B(b[7771]), .Z(n23314) );
XNOR U38858 ( .A(b[7771]), .B(n23315), .Z(c[7771]) );
XNOR U38859 ( .A(a[7771]), .B(c7771), .Z(n23315) );
XOR U38860 ( .A(c7772), .B(n23316), .Z(c7773) );
ANDN U38861 ( .B(n23317), .A(n23318), .Z(n23316) );
XOR U38862 ( .A(c7772), .B(b[7772]), .Z(n23317) );
XNOR U38863 ( .A(b[7772]), .B(n23318), .Z(c[7772]) );
XNOR U38864 ( .A(a[7772]), .B(c7772), .Z(n23318) );
XOR U38865 ( .A(c7773), .B(n23319), .Z(c7774) );
ANDN U38866 ( .B(n23320), .A(n23321), .Z(n23319) );
XOR U38867 ( .A(c7773), .B(b[7773]), .Z(n23320) );
XNOR U38868 ( .A(b[7773]), .B(n23321), .Z(c[7773]) );
XNOR U38869 ( .A(a[7773]), .B(c7773), .Z(n23321) );
XOR U38870 ( .A(c7774), .B(n23322), .Z(c7775) );
ANDN U38871 ( .B(n23323), .A(n23324), .Z(n23322) );
XOR U38872 ( .A(c7774), .B(b[7774]), .Z(n23323) );
XNOR U38873 ( .A(b[7774]), .B(n23324), .Z(c[7774]) );
XNOR U38874 ( .A(a[7774]), .B(c7774), .Z(n23324) );
XOR U38875 ( .A(c7775), .B(n23325), .Z(c7776) );
ANDN U38876 ( .B(n23326), .A(n23327), .Z(n23325) );
XOR U38877 ( .A(c7775), .B(b[7775]), .Z(n23326) );
XNOR U38878 ( .A(b[7775]), .B(n23327), .Z(c[7775]) );
XNOR U38879 ( .A(a[7775]), .B(c7775), .Z(n23327) );
XOR U38880 ( .A(c7776), .B(n23328), .Z(c7777) );
ANDN U38881 ( .B(n23329), .A(n23330), .Z(n23328) );
XOR U38882 ( .A(c7776), .B(b[7776]), .Z(n23329) );
XNOR U38883 ( .A(b[7776]), .B(n23330), .Z(c[7776]) );
XNOR U38884 ( .A(a[7776]), .B(c7776), .Z(n23330) );
XOR U38885 ( .A(c7777), .B(n23331), .Z(c7778) );
ANDN U38886 ( .B(n23332), .A(n23333), .Z(n23331) );
XOR U38887 ( .A(c7777), .B(b[7777]), .Z(n23332) );
XNOR U38888 ( .A(b[7777]), .B(n23333), .Z(c[7777]) );
XNOR U38889 ( .A(a[7777]), .B(c7777), .Z(n23333) );
XOR U38890 ( .A(c7778), .B(n23334), .Z(c7779) );
ANDN U38891 ( .B(n23335), .A(n23336), .Z(n23334) );
XOR U38892 ( .A(c7778), .B(b[7778]), .Z(n23335) );
XNOR U38893 ( .A(b[7778]), .B(n23336), .Z(c[7778]) );
XNOR U38894 ( .A(a[7778]), .B(c7778), .Z(n23336) );
XOR U38895 ( .A(c7779), .B(n23337), .Z(c7780) );
ANDN U38896 ( .B(n23338), .A(n23339), .Z(n23337) );
XOR U38897 ( .A(c7779), .B(b[7779]), .Z(n23338) );
XNOR U38898 ( .A(b[7779]), .B(n23339), .Z(c[7779]) );
XNOR U38899 ( .A(a[7779]), .B(c7779), .Z(n23339) );
XOR U38900 ( .A(c7780), .B(n23340), .Z(c7781) );
ANDN U38901 ( .B(n23341), .A(n23342), .Z(n23340) );
XOR U38902 ( .A(c7780), .B(b[7780]), .Z(n23341) );
XNOR U38903 ( .A(b[7780]), .B(n23342), .Z(c[7780]) );
XNOR U38904 ( .A(a[7780]), .B(c7780), .Z(n23342) );
XOR U38905 ( .A(c7781), .B(n23343), .Z(c7782) );
ANDN U38906 ( .B(n23344), .A(n23345), .Z(n23343) );
XOR U38907 ( .A(c7781), .B(b[7781]), .Z(n23344) );
XNOR U38908 ( .A(b[7781]), .B(n23345), .Z(c[7781]) );
XNOR U38909 ( .A(a[7781]), .B(c7781), .Z(n23345) );
XOR U38910 ( .A(c7782), .B(n23346), .Z(c7783) );
ANDN U38911 ( .B(n23347), .A(n23348), .Z(n23346) );
XOR U38912 ( .A(c7782), .B(b[7782]), .Z(n23347) );
XNOR U38913 ( .A(b[7782]), .B(n23348), .Z(c[7782]) );
XNOR U38914 ( .A(a[7782]), .B(c7782), .Z(n23348) );
XOR U38915 ( .A(c7783), .B(n23349), .Z(c7784) );
ANDN U38916 ( .B(n23350), .A(n23351), .Z(n23349) );
XOR U38917 ( .A(c7783), .B(b[7783]), .Z(n23350) );
XNOR U38918 ( .A(b[7783]), .B(n23351), .Z(c[7783]) );
XNOR U38919 ( .A(a[7783]), .B(c7783), .Z(n23351) );
XOR U38920 ( .A(c7784), .B(n23352), .Z(c7785) );
ANDN U38921 ( .B(n23353), .A(n23354), .Z(n23352) );
XOR U38922 ( .A(c7784), .B(b[7784]), .Z(n23353) );
XNOR U38923 ( .A(b[7784]), .B(n23354), .Z(c[7784]) );
XNOR U38924 ( .A(a[7784]), .B(c7784), .Z(n23354) );
XOR U38925 ( .A(c7785), .B(n23355), .Z(c7786) );
ANDN U38926 ( .B(n23356), .A(n23357), .Z(n23355) );
XOR U38927 ( .A(c7785), .B(b[7785]), .Z(n23356) );
XNOR U38928 ( .A(b[7785]), .B(n23357), .Z(c[7785]) );
XNOR U38929 ( .A(a[7785]), .B(c7785), .Z(n23357) );
XOR U38930 ( .A(c7786), .B(n23358), .Z(c7787) );
ANDN U38931 ( .B(n23359), .A(n23360), .Z(n23358) );
XOR U38932 ( .A(c7786), .B(b[7786]), .Z(n23359) );
XNOR U38933 ( .A(b[7786]), .B(n23360), .Z(c[7786]) );
XNOR U38934 ( .A(a[7786]), .B(c7786), .Z(n23360) );
XOR U38935 ( .A(c7787), .B(n23361), .Z(c7788) );
ANDN U38936 ( .B(n23362), .A(n23363), .Z(n23361) );
XOR U38937 ( .A(c7787), .B(b[7787]), .Z(n23362) );
XNOR U38938 ( .A(b[7787]), .B(n23363), .Z(c[7787]) );
XNOR U38939 ( .A(a[7787]), .B(c7787), .Z(n23363) );
XOR U38940 ( .A(c7788), .B(n23364), .Z(c7789) );
ANDN U38941 ( .B(n23365), .A(n23366), .Z(n23364) );
XOR U38942 ( .A(c7788), .B(b[7788]), .Z(n23365) );
XNOR U38943 ( .A(b[7788]), .B(n23366), .Z(c[7788]) );
XNOR U38944 ( .A(a[7788]), .B(c7788), .Z(n23366) );
XOR U38945 ( .A(c7789), .B(n23367), .Z(c7790) );
ANDN U38946 ( .B(n23368), .A(n23369), .Z(n23367) );
XOR U38947 ( .A(c7789), .B(b[7789]), .Z(n23368) );
XNOR U38948 ( .A(b[7789]), .B(n23369), .Z(c[7789]) );
XNOR U38949 ( .A(a[7789]), .B(c7789), .Z(n23369) );
XOR U38950 ( .A(c7790), .B(n23370), .Z(c7791) );
ANDN U38951 ( .B(n23371), .A(n23372), .Z(n23370) );
XOR U38952 ( .A(c7790), .B(b[7790]), .Z(n23371) );
XNOR U38953 ( .A(b[7790]), .B(n23372), .Z(c[7790]) );
XNOR U38954 ( .A(a[7790]), .B(c7790), .Z(n23372) );
XOR U38955 ( .A(c7791), .B(n23373), .Z(c7792) );
ANDN U38956 ( .B(n23374), .A(n23375), .Z(n23373) );
XOR U38957 ( .A(c7791), .B(b[7791]), .Z(n23374) );
XNOR U38958 ( .A(b[7791]), .B(n23375), .Z(c[7791]) );
XNOR U38959 ( .A(a[7791]), .B(c7791), .Z(n23375) );
XOR U38960 ( .A(c7792), .B(n23376), .Z(c7793) );
ANDN U38961 ( .B(n23377), .A(n23378), .Z(n23376) );
XOR U38962 ( .A(c7792), .B(b[7792]), .Z(n23377) );
XNOR U38963 ( .A(b[7792]), .B(n23378), .Z(c[7792]) );
XNOR U38964 ( .A(a[7792]), .B(c7792), .Z(n23378) );
XOR U38965 ( .A(c7793), .B(n23379), .Z(c7794) );
ANDN U38966 ( .B(n23380), .A(n23381), .Z(n23379) );
XOR U38967 ( .A(c7793), .B(b[7793]), .Z(n23380) );
XNOR U38968 ( .A(b[7793]), .B(n23381), .Z(c[7793]) );
XNOR U38969 ( .A(a[7793]), .B(c7793), .Z(n23381) );
XOR U38970 ( .A(c7794), .B(n23382), .Z(c7795) );
ANDN U38971 ( .B(n23383), .A(n23384), .Z(n23382) );
XOR U38972 ( .A(c7794), .B(b[7794]), .Z(n23383) );
XNOR U38973 ( .A(b[7794]), .B(n23384), .Z(c[7794]) );
XNOR U38974 ( .A(a[7794]), .B(c7794), .Z(n23384) );
XOR U38975 ( .A(c7795), .B(n23385), .Z(c7796) );
ANDN U38976 ( .B(n23386), .A(n23387), .Z(n23385) );
XOR U38977 ( .A(c7795), .B(b[7795]), .Z(n23386) );
XNOR U38978 ( .A(b[7795]), .B(n23387), .Z(c[7795]) );
XNOR U38979 ( .A(a[7795]), .B(c7795), .Z(n23387) );
XOR U38980 ( .A(c7796), .B(n23388), .Z(c7797) );
ANDN U38981 ( .B(n23389), .A(n23390), .Z(n23388) );
XOR U38982 ( .A(c7796), .B(b[7796]), .Z(n23389) );
XNOR U38983 ( .A(b[7796]), .B(n23390), .Z(c[7796]) );
XNOR U38984 ( .A(a[7796]), .B(c7796), .Z(n23390) );
XOR U38985 ( .A(c7797), .B(n23391), .Z(c7798) );
ANDN U38986 ( .B(n23392), .A(n23393), .Z(n23391) );
XOR U38987 ( .A(c7797), .B(b[7797]), .Z(n23392) );
XNOR U38988 ( .A(b[7797]), .B(n23393), .Z(c[7797]) );
XNOR U38989 ( .A(a[7797]), .B(c7797), .Z(n23393) );
XOR U38990 ( .A(c7798), .B(n23394), .Z(c7799) );
ANDN U38991 ( .B(n23395), .A(n23396), .Z(n23394) );
XOR U38992 ( .A(c7798), .B(b[7798]), .Z(n23395) );
XNOR U38993 ( .A(b[7798]), .B(n23396), .Z(c[7798]) );
XNOR U38994 ( .A(a[7798]), .B(c7798), .Z(n23396) );
XOR U38995 ( .A(c7799), .B(n23397), .Z(c7800) );
ANDN U38996 ( .B(n23398), .A(n23399), .Z(n23397) );
XOR U38997 ( .A(c7799), .B(b[7799]), .Z(n23398) );
XNOR U38998 ( .A(b[7799]), .B(n23399), .Z(c[7799]) );
XNOR U38999 ( .A(a[7799]), .B(c7799), .Z(n23399) );
XOR U39000 ( .A(c7800), .B(n23400), .Z(c7801) );
ANDN U39001 ( .B(n23401), .A(n23402), .Z(n23400) );
XOR U39002 ( .A(c7800), .B(b[7800]), .Z(n23401) );
XNOR U39003 ( .A(b[7800]), .B(n23402), .Z(c[7800]) );
XNOR U39004 ( .A(a[7800]), .B(c7800), .Z(n23402) );
XOR U39005 ( .A(c7801), .B(n23403), .Z(c7802) );
ANDN U39006 ( .B(n23404), .A(n23405), .Z(n23403) );
XOR U39007 ( .A(c7801), .B(b[7801]), .Z(n23404) );
XNOR U39008 ( .A(b[7801]), .B(n23405), .Z(c[7801]) );
XNOR U39009 ( .A(a[7801]), .B(c7801), .Z(n23405) );
XOR U39010 ( .A(c7802), .B(n23406), .Z(c7803) );
ANDN U39011 ( .B(n23407), .A(n23408), .Z(n23406) );
XOR U39012 ( .A(c7802), .B(b[7802]), .Z(n23407) );
XNOR U39013 ( .A(b[7802]), .B(n23408), .Z(c[7802]) );
XNOR U39014 ( .A(a[7802]), .B(c7802), .Z(n23408) );
XOR U39015 ( .A(c7803), .B(n23409), .Z(c7804) );
ANDN U39016 ( .B(n23410), .A(n23411), .Z(n23409) );
XOR U39017 ( .A(c7803), .B(b[7803]), .Z(n23410) );
XNOR U39018 ( .A(b[7803]), .B(n23411), .Z(c[7803]) );
XNOR U39019 ( .A(a[7803]), .B(c7803), .Z(n23411) );
XOR U39020 ( .A(c7804), .B(n23412), .Z(c7805) );
ANDN U39021 ( .B(n23413), .A(n23414), .Z(n23412) );
XOR U39022 ( .A(c7804), .B(b[7804]), .Z(n23413) );
XNOR U39023 ( .A(b[7804]), .B(n23414), .Z(c[7804]) );
XNOR U39024 ( .A(a[7804]), .B(c7804), .Z(n23414) );
XOR U39025 ( .A(c7805), .B(n23415), .Z(c7806) );
ANDN U39026 ( .B(n23416), .A(n23417), .Z(n23415) );
XOR U39027 ( .A(c7805), .B(b[7805]), .Z(n23416) );
XNOR U39028 ( .A(b[7805]), .B(n23417), .Z(c[7805]) );
XNOR U39029 ( .A(a[7805]), .B(c7805), .Z(n23417) );
XOR U39030 ( .A(c7806), .B(n23418), .Z(c7807) );
ANDN U39031 ( .B(n23419), .A(n23420), .Z(n23418) );
XOR U39032 ( .A(c7806), .B(b[7806]), .Z(n23419) );
XNOR U39033 ( .A(b[7806]), .B(n23420), .Z(c[7806]) );
XNOR U39034 ( .A(a[7806]), .B(c7806), .Z(n23420) );
XOR U39035 ( .A(c7807), .B(n23421), .Z(c7808) );
ANDN U39036 ( .B(n23422), .A(n23423), .Z(n23421) );
XOR U39037 ( .A(c7807), .B(b[7807]), .Z(n23422) );
XNOR U39038 ( .A(b[7807]), .B(n23423), .Z(c[7807]) );
XNOR U39039 ( .A(a[7807]), .B(c7807), .Z(n23423) );
XOR U39040 ( .A(c7808), .B(n23424), .Z(c7809) );
ANDN U39041 ( .B(n23425), .A(n23426), .Z(n23424) );
XOR U39042 ( .A(c7808), .B(b[7808]), .Z(n23425) );
XNOR U39043 ( .A(b[7808]), .B(n23426), .Z(c[7808]) );
XNOR U39044 ( .A(a[7808]), .B(c7808), .Z(n23426) );
XOR U39045 ( .A(c7809), .B(n23427), .Z(c7810) );
ANDN U39046 ( .B(n23428), .A(n23429), .Z(n23427) );
XOR U39047 ( .A(c7809), .B(b[7809]), .Z(n23428) );
XNOR U39048 ( .A(b[7809]), .B(n23429), .Z(c[7809]) );
XNOR U39049 ( .A(a[7809]), .B(c7809), .Z(n23429) );
XOR U39050 ( .A(c7810), .B(n23430), .Z(c7811) );
ANDN U39051 ( .B(n23431), .A(n23432), .Z(n23430) );
XOR U39052 ( .A(c7810), .B(b[7810]), .Z(n23431) );
XNOR U39053 ( .A(b[7810]), .B(n23432), .Z(c[7810]) );
XNOR U39054 ( .A(a[7810]), .B(c7810), .Z(n23432) );
XOR U39055 ( .A(c7811), .B(n23433), .Z(c7812) );
ANDN U39056 ( .B(n23434), .A(n23435), .Z(n23433) );
XOR U39057 ( .A(c7811), .B(b[7811]), .Z(n23434) );
XNOR U39058 ( .A(b[7811]), .B(n23435), .Z(c[7811]) );
XNOR U39059 ( .A(a[7811]), .B(c7811), .Z(n23435) );
XOR U39060 ( .A(c7812), .B(n23436), .Z(c7813) );
ANDN U39061 ( .B(n23437), .A(n23438), .Z(n23436) );
XOR U39062 ( .A(c7812), .B(b[7812]), .Z(n23437) );
XNOR U39063 ( .A(b[7812]), .B(n23438), .Z(c[7812]) );
XNOR U39064 ( .A(a[7812]), .B(c7812), .Z(n23438) );
XOR U39065 ( .A(c7813), .B(n23439), .Z(c7814) );
ANDN U39066 ( .B(n23440), .A(n23441), .Z(n23439) );
XOR U39067 ( .A(c7813), .B(b[7813]), .Z(n23440) );
XNOR U39068 ( .A(b[7813]), .B(n23441), .Z(c[7813]) );
XNOR U39069 ( .A(a[7813]), .B(c7813), .Z(n23441) );
XOR U39070 ( .A(c7814), .B(n23442), .Z(c7815) );
ANDN U39071 ( .B(n23443), .A(n23444), .Z(n23442) );
XOR U39072 ( .A(c7814), .B(b[7814]), .Z(n23443) );
XNOR U39073 ( .A(b[7814]), .B(n23444), .Z(c[7814]) );
XNOR U39074 ( .A(a[7814]), .B(c7814), .Z(n23444) );
XOR U39075 ( .A(c7815), .B(n23445), .Z(c7816) );
ANDN U39076 ( .B(n23446), .A(n23447), .Z(n23445) );
XOR U39077 ( .A(c7815), .B(b[7815]), .Z(n23446) );
XNOR U39078 ( .A(b[7815]), .B(n23447), .Z(c[7815]) );
XNOR U39079 ( .A(a[7815]), .B(c7815), .Z(n23447) );
XOR U39080 ( .A(c7816), .B(n23448), .Z(c7817) );
ANDN U39081 ( .B(n23449), .A(n23450), .Z(n23448) );
XOR U39082 ( .A(c7816), .B(b[7816]), .Z(n23449) );
XNOR U39083 ( .A(b[7816]), .B(n23450), .Z(c[7816]) );
XNOR U39084 ( .A(a[7816]), .B(c7816), .Z(n23450) );
XOR U39085 ( .A(c7817), .B(n23451), .Z(c7818) );
ANDN U39086 ( .B(n23452), .A(n23453), .Z(n23451) );
XOR U39087 ( .A(c7817), .B(b[7817]), .Z(n23452) );
XNOR U39088 ( .A(b[7817]), .B(n23453), .Z(c[7817]) );
XNOR U39089 ( .A(a[7817]), .B(c7817), .Z(n23453) );
XOR U39090 ( .A(c7818), .B(n23454), .Z(c7819) );
ANDN U39091 ( .B(n23455), .A(n23456), .Z(n23454) );
XOR U39092 ( .A(c7818), .B(b[7818]), .Z(n23455) );
XNOR U39093 ( .A(b[7818]), .B(n23456), .Z(c[7818]) );
XNOR U39094 ( .A(a[7818]), .B(c7818), .Z(n23456) );
XOR U39095 ( .A(c7819), .B(n23457), .Z(c7820) );
ANDN U39096 ( .B(n23458), .A(n23459), .Z(n23457) );
XOR U39097 ( .A(c7819), .B(b[7819]), .Z(n23458) );
XNOR U39098 ( .A(b[7819]), .B(n23459), .Z(c[7819]) );
XNOR U39099 ( .A(a[7819]), .B(c7819), .Z(n23459) );
XOR U39100 ( .A(c7820), .B(n23460), .Z(c7821) );
ANDN U39101 ( .B(n23461), .A(n23462), .Z(n23460) );
XOR U39102 ( .A(c7820), .B(b[7820]), .Z(n23461) );
XNOR U39103 ( .A(b[7820]), .B(n23462), .Z(c[7820]) );
XNOR U39104 ( .A(a[7820]), .B(c7820), .Z(n23462) );
XOR U39105 ( .A(c7821), .B(n23463), .Z(c7822) );
ANDN U39106 ( .B(n23464), .A(n23465), .Z(n23463) );
XOR U39107 ( .A(c7821), .B(b[7821]), .Z(n23464) );
XNOR U39108 ( .A(b[7821]), .B(n23465), .Z(c[7821]) );
XNOR U39109 ( .A(a[7821]), .B(c7821), .Z(n23465) );
XOR U39110 ( .A(c7822), .B(n23466), .Z(c7823) );
ANDN U39111 ( .B(n23467), .A(n23468), .Z(n23466) );
XOR U39112 ( .A(c7822), .B(b[7822]), .Z(n23467) );
XNOR U39113 ( .A(b[7822]), .B(n23468), .Z(c[7822]) );
XNOR U39114 ( .A(a[7822]), .B(c7822), .Z(n23468) );
XOR U39115 ( .A(c7823), .B(n23469), .Z(c7824) );
ANDN U39116 ( .B(n23470), .A(n23471), .Z(n23469) );
XOR U39117 ( .A(c7823), .B(b[7823]), .Z(n23470) );
XNOR U39118 ( .A(b[7823]), .B(n23471), .Z(c[7823]) );
XNOR U39119 ( .A(a[7823]), .B(c7823), .Z(n23471) );
XOR U39120 ( .A(c7824), .B(n23472), .Z(c7825) );
ANDN U39121 ( .B(n23473), .A(n23474), .Z(n23472) );
XOR U39122 ( .A(c7824), .B(b[7824]), .Z(n23473) );
XNOR U39123 ( .A(b[7824]), .B(n23474), .Z(c[7824]) );
XNOR U39124 ( .A(a[7824]), .B(c7824), .Z(n23474) );
XOR U39125 ( .A(c7825), .B(n23475), .Z(c7826) );
ANDN U39126 ( .B(n23476), .A(n23477), .Z(n23475) );
XOR U39127 ( .A(c7825), .B(b[7825]), .Z(n23476) );
XNOR U39128 ( .A(b[7825]), .B(n23477), .Z(c[7825]) );
XNOR U39129 ( .A(a[7825]), .B(c7825), .Z(n23477) );
XOR U39130 ( .A(c7826), .B(n23478), .Z(c7827) );
ANDN U39131 ( .B(n23479), .A(n23480), .Z(n23478) );
XOR U39132 ( .A(c7826), .B(b[7826]), .Z(n23479) );
XNOR U39133 ( .A(b[7826]), .B(n23480), .Z(c[7826]) );
XNOR U39134 ( .A(a[7826]), .B(c7826), .Z(n23480) );
XOR U39135 ( .A(c7827), .B(n23481), .Z(c7828) );
ANDN U39136 ( .B(n23482), .A(n23483), .Z(n23481) );
XOR U39137 ( .A(c7827), .B(b[7827]), .Z(n23482) );
XNOR U39138 ( .A(b[7827]), .B(n23483), .Z(c[7827]) );
XNOR U39139 ( .A(a[7827]), .B(c7827), .Z(n23483) );
XOR U39140 ( .A(c7828), .B(n23484), .Z(c7829) );
ANDN U39141 ( .B(n23485), .A(n23486), .Z(n23484) );
XOR U39142 ( .A(c7828), .B(b[7828]), .Z(n23485) );
XNOR U39143 ( .A(b[7828]), .B(n23486), .Z(c[7828]) );
XNOR U39144 ( .A(a[7828]), .B(c7828), .Z(n23486) );
XOR U39145 ( .A(c7829), .B(n23487), .Z(c7830) );
ANDN U39146 ( .B(n23488), .A(n23489), .Z(n23487) );
XOR U39147 ( .A(c7829), .B(b[7829]), .Z(n23488) );
XNOR U39148 ( .A(b[7829]), .B(n23489), .Z(c[7829]) );
XNOR U39149 ( .A(a[7829]), .B(c7829), .Z(n23489) );
XOR U39150 ( .A(c7830), .B(n23490), .Z(c7831) );
ANDN U39151 ( .B(n23491), .A(n23492), .Z(n23490) );
XOR U39152 ( .A(c7830), .B(b[7830]), .Z(n23491) );
XNOR U39153 ( .A(b[7830]), .B(n23492), .Z(c[7830]) );
XNOR U39154 ( .A(a[7830]), .B(c7830), .Z(n23492) );
XOR U39155 ( .A(c7831), .B(n23493), .Z(c7832) );
ANDN U39156 ( .B(n23494), .A(n23495), .Z(n23493) );
XOR U39157 ( .A(c7831), .B(b[7831]), .Z(n23494) );
XNOR U39158 ( .A(b[7831]), .B(n23495), .Z(c[7831]) );
XNOR U39159 ( .A(a[7831]), .B(c7831), .Z(n23495) );
XOR U39160 ( .A(c7832), .B(n23496), .Z(c7833) );
ANDN U39161 ( .B(n23497), .A(n23498), .Z(n23496) );
XOR U39162 ( .A(c7832), .B(b[7832]), .Z(n23497) );
XNOR U39163 ( .A(b[7832]), .B(n23498), .Z(c[7832]) );
XNOR U39164 ( .A(a[7832]), .B(c7832), .Z(n23498) );
XOR U39165 ( .A(c7833), .B(n23499), .Z(c7834) );
ANDN U39166 ( .B(n23500), .A(n23501), .Z(n23499) );
XOR U39167 ( .A(c7833), .B(b[7833]), .Z(n23500) );
XNOR U39168 ( .A(b[7833]), .B(n23501), .Z(c[7833]) );
XNOR U39169 ( .A(a[7833]), .B(c7833), .Z(n23501) );
XOR U39170 ( .A(c7834), .B(n23502), .Z(c7835) );
ANDN U39171 ( .B(n23503), .A(n23504), .Z(n23502) );
XOR U39172 ( .A(c7834), .B(b[7834]), .Z(n23503) );
XNOR U39173 ( .A(b[7834]), .B(n23504), .Z(c[7834]) );
XNOR U39174 ( .A(a[7834]), .B(c7834), .Z(n23504) );
XOR U39175 ( .A(c7835), .B(n23505), .Z(c7836) );
ANDN U39176 ( .B(n23506), .A(n23507), .Z(n23505) );
XOR U39177 ( .A(c7835), .B(b[7835]), .Z(n23506) );
XNOR U39178 ( .A(b[7835]), .B(n23507), .Z(c[7835]) );
XNOR U39179 ( .A(a[7835]), .B(c7835), .Z(n23507) );
XOR U39180 ( .A(c7836), .B(n23508), .Z(c7837) );
ANDN U39181 ( .B(n23509), .A(n23510), .Z(n23508) );
XOR U39182 ( .A(c7836), .B(b[7836]), .Z(n23509) );
XNOR U39183 ( .A(b[7836]), .B(n23510), .Z(c[7836]) );
XNOR U39184 ( .A(a[7836]), .B(c7836), .Z(n23510) );
XOR U39185 ( .A(c7837), .B(n23511), .Z(c7838) );
ANDN U39186 ( .B(n23512), .A(n23513), .Z(n23511) );
XOR U39187 ( .A(c7837), .B(b[7837]), .Z(n23512) );
XNOR U39188 ( .A(b[7837]), .B(n23513), .Z(c[7837]) );
XNOR U39189 ( .A(a[7837]), .B(c7837), .Z(n23513) );
XOR U39190 ( .A(c7838), .B(n23514), .Z(c7839) );
ANDN U39191 ( .B(n23515), .A(n23516), .Z(n23514) );
XOR U39192 ( .A(c7838), .B(b[7838]), .Z(n23515) );
XNOR U39193 ( .A(b[7838]), .B(n23516), .Z(c[7838]) );
XNOR U39194 ( .A(a[7838]), .B(c7838), .Z(n23516) );
XOR U39195 ( .A(c7839), .B(n23517), .Z(c7840) );
ANDN U39196 ( .B(n23518), .A(n23519), .Z(n23517) );
XOR U39197 ( .A(c7839), .B(b[7839]), .Z(n23518) );
XNOR U39198 ( .A(b[7839]), .B(n23519), .Z(c[7839]) );
XNOR U39199 ( .A(a[7839]), .B(c7839), .Z(n23519) );
XOR U39200 ( .A(c7840), .B(n23520), .Z(c7841) );
ANDN U39201 ( .B(n23521), .A(n23522), .Z(n23520) );
XOR U39202 ( .A(c7840), .B(b[7840]), .Z(n23521) );
XNOR U39203 ( .A(b[7840]), .B(n23522), .Z(c[7840]) );
XNOR U39204 ( .A(a[7840]), .B(c7840), .Z(n23522) );
XOR U39205 ( .A(c7841), .B(n23523), .Z(c7842) );
ANDN U39206 ( .B(n23524), .A(n23525), .Z(n23523) );
XOR U39207 ( .A(c7841), .B(b[7841]), .Z(n23524) );
XNOR U39208 ( .A(b[7841]), .B(n23525), .Z(c[7841]) );
XNOR U39209 ( .A(a[7841]), .B(c7841), .Z(n23525) );
XOR U39210 ( .A(c7842), .B(n23526), .Z(c7843) );
ANDN U39211 ( .B(n23527), .A(n23528), .Z(n23526) );
XOR U39212 ( .A(c7842), .B(b[7842]), .Z(n23527) );
XNOR U39213 ( .A(b[7842]), .B(n23528), .Z(c[7842]) );
XNOR U39214 ( .A(a[7842]), .B(c7842), .Z(n23528) );
XOR U39215 ( .A(c7843), .B(n23529), .Z(c7844) );
ANDN U39216 ( .B(n23530), .A(n23531), .Z(n23529) );
XOR U39217 ( .A(c7843), .B(b[7843]), .Z(n23530) );
XNOR U39218 ( .A(b[7843]), .B(n23531), .Z(c[7843]) );
XNOR U39219 ( .A(a[7843]), .B(c7843), .Z(n23531) );
XOR U39220 ( .A(c7844), .B(n23532), .Z(c7845) );
ANDN U39221 ( .B(n23533), .A(n23534), .Z(n23532) );
XOR U39222 ( .A(c7844), .B(b[7844]), .Z(n23533) );
XNOR U39223 ( .A(b[7844]), .B(n23534), .Z(c[7844]) );
XNOR U39224 ( .A(a[7844]), .B(c7844), .Z(n23534) );
XOR U39225 ( .A(c7845), .B(n23535), .Z(c7846) );
ANDN U39226 ( .B(n23536), .A(n23537), .Z(n23535) );
XOR U39227 ( .A(c7845), .B(b[7845]), .Z(n23536) );
XNOR U39228 ( .A(b[7845]), .B(n23537), .Z(c[7845]) );
XNOR U39229 ( .A(a[7845]), .B(c7845), .Z(n23537) );
XOR U39230 ( .A(c7846), .B(n23538), .Z(c7847) );
ANDN U39231 ( .B(n23539), .A(n23540), .Z(n23538) );
XOR U39232 ( .A(c7846), .B(b[7846]), .Z(n23539) );
XNOR U39233 ( .A(b[7846]), .B(n23540), .Z(c[7846]) );
XNOR U39234 ( .A(a[7846]), .B(c7846), .Z(n23540) );
XOR U39235 ( .A(c7847), .B(n23541), .Z(c7848) );
ANDN U39236 ( .B(n23542), .A(n23543), .Z(n23541) );
XOR U39237 ( .A(c7847), .B(b[7847]), .Z(n23542) );
XNOR U39238 ( .A(b[7847]), .B(n23543), .Z(c[7847]) );
XNOR U39239 ( .A(a[7847]), .B(c7847), .Z(n23543) );
XOR U39240 ( .A(c7848), .B(n23544), .Z(c7849) );
ANDN U39241 ( .B(n23545), .A(n23546), .Z(n23544) );
XOR U39242 ( .A(c7848), .B(b[7848]), .Z(n23545) );
XNOR U39243 ( .A(b[7848]), .B(n23546), .Z(c[7848]) );
XNOR U39244 ( .A(a[7848]), .B(c7848), .Z(n23546) );
XOR U39245 ( .A(c7849), .B(n23547), .Z(c7850) );
ANDN U39246 ( .B(n23548), .A(n23549), .Z(n23547) );
XOR U39247 ( .A(c7849), .B(b[7849]), .Z(n23548) );
XNOR U39248 ( .A(b[7849]), .B(n23549), .Z(c[7849]) );
XNOR U39249 ( .A(a[7849]), .B(c7849), .Z(n23549) );
XOR U39250 ( .A(c7850), .B(n23550), .Z(c7851) );
ANDN U39251 ( .B(n23551), .A(n23552), .Z(n23550) );
XOR U39252 ( .A(c7850), .B(b[7850]), .Z(n23551) );
XNOR U39253 ( .A(b[7850]), .B(n23552), .Z(c[7850]) );
XNOR U39254 ( .A(a[7850]), .B(c7850), .Z(n23552) );
XOR U39255 ( .A(c7851), .B(n23553), .Z(c7852) );
ANDN U39256 ( .B(n23554), .A(n23555), .Z(n23553) );
XOR U39257 ( .A(c7851), .B(b[7851]), .Z(n23554) );
XNOR U39258 ( .A(b[7851]), .B(n23555), .Z(c[7851]) );
XNOR U39259 ( .A(a[7851]), .B(c7851), .Z(n23555) );
XOR U39260 ( .A(c7852), .B(n23556), .Z(c7853) );
ANDN U39261 ( .B(n23557), .A(n23558), .Z(n23556) );
XOR U39262 ( .A(c7852), .B(b[7852]), .Z(n23557) );
XNOR U39263 ( .A(b[7852]), .B(n23558), .Z(c[7852]) );
XNOR U39264 ( .A(a[7852]), .B(c7852), .Z(n23558) );
XOR U39265 ( .A(c7853), .B(n23559), .Z(c7854) );
ANDN U39266 ( .B(n23560), .A(n23561), .Z(n23559) );
XOR U39267 ( .A(c7853), .B(b[7853]), .Z(n23560) );
XNOR U39268 ( .A(b[7853]), .B(n23561), .Z(c[7853]) );
XNOR U39269 ( .A(a[7853]), .B(c7853), .Z(n23561) );
XOR U39270 ( .A(c7854), .B(n23562), .Z(c7855) );
ANDN U39271 ( .B(n23563), .A(n23564), .Z(n23562) );
XOR U39272 ( .A(c7854), .B(b[7854]), .Z(n23563) );
XNOR U39273 ( .A(b[7854]), .B(n23564), .Z(c[7854]) );
XNOR U39274 ( .A(a[7854]), .B(c7854), .Z(n23564) );
XOR U39275 ( .A(c7855), .B(n23565), .Z(c7856) );
ANDN U39276 ( .B(n23566), .A(n23567), .Z(n23565) );
XOR U39277 ( .A(c7855), .B(b[7855]), .Z(n23566) );
XNOR U39278 ( .A(b[7855]), .B(n23567), .Z(c[7855]) );
XNOR U39279 ( .A(a[7855]), .B(c7855), .Z(n23567) );
XOR U39280 ( .A(c7856), .B(n23568), .Z(c7857) );
ANDN U39281 ( .B(n23569), .A(n23570), .Z(n23568) );
XOR U39282 ( .A(c7856), .B(b[7856]), .Z(n23569) );
XNOR U39283 ( .A(b[7856]), .B(n23570), .Z(c[7856]) );
XNOR U39284 ( .A(a[7856]), .B(c7856), .Z(n23570) );
XOR U39285 ( .A(c7857), .B(n23571), .Z(c7858) );
ANDN U39286 ( .B(n23572), .A(n23573), .Z(n23571) );
XOR U39287 ( .A(c7857), .B(b[7857]), .Z(n23572) );
XNOR U39288 ( .A(b[7857]), .B(n23573), .Z(c[7857]) );
XNOR U39289 ( .A(a[7857]), .B(c7857), .Z(n23573) );
XOR U39290 ( .A(c7858), .B(n23574), .Z(c7859) );
ANDN U39291 ( .B(n23575), .A(n23576), .Z(n23574) );
XOR U39292 ( .A(c7858), .B(b[7858]), .Z(n23575) );
XNOR U39293 ( .A(b[7858]), .B(n23576), .Z(c[7858]) );
XNOR U39294 ( .A(a[7858]), .B(c7858), .Z(n23576) );
XOR U39295 ( .A(c7859), .B(n23577), .Z(c7860) );
ANDN U39296 ( .B(n23578), .A(n23579), .Z(n23577) );
XOR U39297 ( .A(c7859), .B(b[7859]), .Z(n23578) );
XNOR U39298 ( .A(b[7859]), .B(n23579), .Z(c[7859]) );
XNOR U39299 ( .A(a[7859]), .B(c7859), .Z(n23579) );
XOR U39300 ( .A(c7860), .B(n23580), .Z(c7861) );
ANDN U39301 ( .B(n23581), .A(n23582), .Z(n23580) );
XOR U39302 ( .A(c7860), .B(b[7860]), .Z(n23581) );
XNOR U39303 ( .A(b[7860]), .B(n23582), .Z(c[7860]) );
XNOR U39304 ( .A(a[7860]), .B(c7860), .Z(n23582) );
XOR U39305 ( .A(c7861), .B(n23583), .Z(c7862) );
ANDN U39306 ( .B(n23584), .A(n23585), .Z(n23583) );
XOR U39307 ( .A(c7861), .B(b[7861]), .Z(n23584) );
XNOR U39308 ( .A(b[7861]), .B(n23585), .Z(c[7861]) );
XNOR U39309 ( .A(a[7861]), .B(c7861), .Z(n23585) );
XOR U39310 ( .A(c7862), .B(n23586), .Z(c7863) );
ANDN U39311 ( .B(n23587), .A(n23588), .Z(n23586) );
XOR U39312 ( .A(c7862), .B(b[7862]), .Z(n23587) );
XNOR U39313 ( .A(b[7862]), .B(n23588), .Z(c[7862]) );
XNOR U39314 ( .A(a[7862]), .B(c7862), .Z(n23588) );
XOR U39315 ( .A(c7863), .B(n23589), .Z(c7864) );
ANDN U39316 ( .B(n23590), .A(n23591), .Z(n23589) );
XOR U39317 ( .A(c7863), .B(b[7863]), .Z(n23590) );
XNOR U39318 ( .A(b[7863]), .B(n23591), .Z(c[7863]) );
XNOR U39319 ( .A(a[7863]), .B(c7863), .Z(n23591) );
XOR U39320 ( .A(c7864), .B(n23592), .Z(c7865) );
ANDN U39321 ( .B(n23593), .A(n23594), .Z(n23592) );
XOR U39322 ( .A(c7864), .B(b[7864]), .Z(n23593) );
XNOR U39323 ( .A(b[7864]), .B(n23594), .Z(c[7864]) );
XNOR U39324 ( .A(a[7864]), .B(c7864), .Z(n23594) );
XOR U39325 ( .A(c7865), .B(n23595), .Z(c7866) );
ANDN U39326 ( .B(n23596), .A(n23597), .Z(n23595) );
XOR U39327 ( .A(c7865), .B(b[7865]), .Z(n23596) );
XNOR U39328 ( .A(b[7865]), .B(n23597), .Z(c[7865]) );
XNOR U39329 ( .A(a[7865]), .B(c7865), .Z(n23597) );
XOR U39330 ( .A(c7866), .B(n23598), .Z(c7867) );
ANDN U39331 ( .B(n23599), .A(n23600), .Z(n23598) );
XOR U39332 ( .A(c7866), .B(b[7866]), .Z(n23599) );
XNOR U39333 ( .A(b[7866]), .B(n23600), .Z(c[7866]) );
XNOR U39334 ( .A(a[7866]), .B(c7866), .Z(n23600) );
XOR U39335 ( .A(c7867), .B(n23601), .Z(c7868) );
ANDN U39336 ( .B(n23602), .A(n23603), .Z(n23601) );
XOR U39337 ( .A(c7867), .B(b[7867]), .Z(n23602) );
XNOR U39338 ( .A(b[7867]), .B(n23603), .Z(c[7867]) );
XNOR U39339 ( .A(a[7867]), .B(c7867), .Z(n23603) );
XOR U39340 ( .A(c7868), .B(n23604), .Z(c7869) );
ANDN U39341 ( .B(n23605), .A(n23606), .Z(n23604) );
XOR U39342 ( .A(c7868), .B(b[7868]), .Z(n23605) );
XNOR U39343 ( .A(b[7868]), .B(n23606), .Z(c[7868]) );
XNOR U39344 ( .A(a[7868]), .B(c7868), .Z(n23606) );
XOR U39345 ( .A(c7869), .B(n23607), .Z(c7870) );
ANDN U39346 ( .B(n23608), .A(n23609), .Z(n23607) );
XOR U39347 ( .A(c7869), .B(b[7869]), .Z(n23608) );
XNOR U39348 ( .A(b[7869]), .B(n23609), .Z(c[7869]) );
XNOR U39349 ( .A(a[7869]), .B(c7869), .Z(n23609) );
XOR U39350 ( .A(c7870), .B(n23610), .Z(c7871) );
ANDN U39351 ( .B(n23611), .A(n23612), .Z(n23610) );
XOR U39352 ( .A(c7870), .B(b[7870]), .Z(n23611) );
XNOR U39353 ( .A(b[7870]), .B(n23612), .Z(c[7870]) );
XNOR U39354 ( .A(a[7870]), .B(c7870), .Z(n23612) );
XOR U39355 ( .A(c7871), .B(n23613), .Z(c7872) );
ANDN U39356 ( .B(n23614), .A(n23615), .Z(n23613) );
XOR U39357 ( .A(c7871), .B(b[7871]), .Z(n23614) );
XNOR U39358 ( .A(b[7871]), .B(n23615), .Z(c[7871]) );
XNOR U39359 ( .A(a[7871]), .B(c7871), .Z(n23615) );
XOR U39360 ( .A(c7872), .B(n23616), .Z(c7873) );
ANDN U39361 ( .B(n23617), .A(n23618), .Z(n23616) );
XOR U39362 ( .A(c7872), .B(b[7872]), .Z(n23617) );
XNOR U39363 ( .A(b[7872]), .B(n23618), .Z(c[7872]) );
XNOR U39364 ( .A(a[7872]), .B(c7872), .Z(n23618) );
XOR U39365 ( .A(c7873), .B(n23619), .Z(c7874) );
ANDN U39366 ( .B(n23620), .A(n23621), .Z(n23619) );
XOR U39367 ( .A(c7873), .B(b[7873]), .Z(n23620) );
XNOR U39368 ( .A(b[7873]), .B(n23621), .Z(c[7873]) );
XNOR U39369 ( .A(a[7873]), .B(c7873), .Z(n23621) );
XOR U39370 ( .A(c7874), .B(n23622), .Z(c7875) );
ANDN U39371 ( .B(n23623), .A(n23624), .Z(n23622) );
XOR U39372 ( .A(c7874), .B(b[7874]), .Z(n23623) );
XNOR U39373 ( .A(b[7874]), .B(n23624), .Z(c[7874]) );
XNOR U39374 ( .A(a[7874]), .B(c7874), .Z(n23624) );
XOR U39375 ( .A(c7875), .B(n23625), .Z(c7876) );
ANDN U39376 ( .B(n23626), .A(n23627), .Z(n23625) );
XOR U39377 ( .A(c7875), .B(b[7875]), .Z(n23626) );
XNOR U39378 ( .A(b[7875]), .B(n23627), .Z(c[7875]) );
XNOR U39379 ( .A(a[7875]), .B(c7875), .Z(n23627) );
XOR U39380 ( .A(c7876), .B(n23628), .Z(c7877) );
ANDN U39381 ( .B(n23629), .A(n23630), .Z(n23628) );
XOR U39382 ( .A(c7876), .B(b[7876]), .Z(n23629) );
XNOR U39383 ( .A(b[7876]), .B(n23630), .Z(c[7876]) );
XNOR U39384 ( .A(a[7876]), .B(c7876), .Z(n23630) );
XOR U39385 ( .A(c7877), .B(n23631), .Z(c7878) );
ANDN U39386 ( .B(n23632), .A(n23633), .Z(n23631) );
XOR U39387 ( .A(c7877), .B(b[7877]), .Z(n23632) );
XNOR U39388 ( .A(b[7877]), .B(n23633), .Z(c[7877]) );
XNOR U39389 ( .A(a[7877]), .B(c7877), .Z(n23633) );
XOR U39390 ( .A(c7878), .B(n23634), .Z(c7879) );
ANDN U39391 ( .B(n23635), .A(n23636), .Z(n23634) );
XOR U39392 ( .A(c7878), .B(b[7878]), .Z(n23635) );
XNOR U39393 ( .A(b[7878]), .B(n23636), .Z(c[7878]) );
XNOR U39394 ( .A(a[7878]), .B(c7878), .Z(n23636) );
XOR U39395 ( .A(c7879), .B(n23637), .Z(c7880) );
ANDN U39396 ( .B(n23638), .A(n23639), .Z(n23637) );
XOR U39397 ( .A(c7879), .B(b[7879]), .Z(n23638) );
XNOR U39398 ( .A(b[7879]), .B(n23639), .Z(c[7879]) );
XNOR U39399 ( .A(a[7879]), .B(c7879), .Z(n23639) );
XOR U39400 ( .A(c7880), .B(n23640), .Z(c7881) );
ANDN U39401 ( .B(n23641), .A(n23642), .Z(n23640) );
XOR U39402 ( .A(c7880), .B(b[7880]), .Z(n23641) );
XNOR U39403 ( .A(b[7880]), .B(n23642), .Z(c[7880]) );
XNOR U39404 ( .A(a[7880]), .B(c7880), .Z(n23642) );
XOR U39405 ( .A(c7881), .B(n23643), .Z(c7882) );
ANDN U39406 ( .B(n23644), .A(n23645), .Z(n23643) );
XOR U39407 ( .A(c7881), .B(b[7881]), .Z(n23644) );
XNOR U39408 ( .A(b[7881]), .B(n23645), .Z(c[7881]) );
XNOR U39409 ( .A(a[7881]), .B(c7881), .Z(n23645) );
XOR U39410 ( .A(c7882), .B(n23646), .Z(c7883) );
ANDN U39411 ( .B(n23647), .A(n23648), .Z(n23646) );
XOR U39412 ( .A(c7882), .B(b[7882]), .Z(n23647) );
XNOR U39413 ( .A(b[7882]), .B(n23648), .Z(c[7882]) );
XNOR U39414 ( .A(a[7882]), .B(c7882), .Z(n23648) );
XOR U39415 ( .A(c7883), .B(n23649), .Z(c7884) );
ANDN U39416 ( .B(n23650), .A(n23651), .Z(n23649) );
XOR U39417 ( .A(c7883), .B(b[7883]), .Z(n23650) );
XNOR U39418 ( .A(b[7883]), .B(n23651), .Z(c[7883]) );
XNOR U39419 ( .A(a[7883]), .B(c7883), .Z(n23651) );
XOR U39420 ( .A(c7884), .B(n23652), .Z(c7885) );
ANDN U39421 ( .B(n23653), .A(n23654), .Z(n23652) );
XOR U39422 ( .A(c7884), .B(b[7884]), .Z(n23653) );
XNOR U39423 ( .A(b[7884]), .B(n23654), .Z(c[7884]) );
XNOR U39424 ( .A(a[7884]), .B(c7884), .Z(n23654) );
XOR U39425 ( .A(c7885), .B(n23655), .Z(c7886) );
ANDN U39426 ( .B(n23656), .A(n23657), .Z(n23655) );
XOR U39427 ( .A(c7885), .B(b[7885]), .Z(n23656) );
XNOR U39428 ( .A(b[7885]), .B(n23657), .Z(c[7885]) );
XNOR U39429 ( .A(a[7885]), .B(c7885), .Z(n23657) );
XOR U39430 ( .A(c7886), .B(n23658), .Z(c7887) );
ANDN U39431 ( .B(n23659), .A(n23660), .Z(n23658) );
XOR U39432 ( .A(c7886), .B(b[7886]), .Z(n23659) );
XNOR U39433 ( .A(b[7886]), .B(n23660), .Z(c[7886]) );
XNOR U39434 ( .A(a[7886]), .B(c7886), .Z(n23660) );
XOR U39435 ( .A(c7887), .B(n23661), .Z(c7888) );
ANDN U39436 ( .B(n23662), .A(n23663), .Z(n23661) );
XOR U39437 ( .A(c7887), .B(b[7887]), .Z(n23662) );
XNOR U39438 ( .A(b[7887]), .B(n23663), .Z(c[7887]) );
XNOR U39439 ( .A(a[7887]), .B(c7887), .Z(n23663) );
XOR U39440 ( .A(c7888), .B(n23664), .Z(c7889) );
ANDN U39441 ( .B(n23665), .A(n23666), .Z(n23664) );
XOR U39442 ( .A(c7888), .B(b[7888]), .Z(n23665) );
XNOR U39443 ( .A(b[7888]), .B(n23666), .Z(c[7888]) );
XNOR U39444 ( .A(a[7888]), .B(c7888), .Z(n23666) );
XOR U39445 ( .A(c7889), .B(n23667), .Z(c7890) );
ANDN U39446 ( .B(n23668), .A(n23669), .Z(n23667) );
XOR U39447 ( .A(c7889), .B(b[7889]), .Z(n23668) );
XNOR U39448 ( .A(b[7889]), .B(n23669), .Z(c[7889]) );
XNOR U39449 ( .A(a[7889]), .B(c7889), .Z(n23669) );
XOR U39450 ( .A(c7890), .B(n23670), .Z(c7891) );
ANDN U39451 ( .B(n23671), .A(n23672), .Z(n23670) );
XOR U39452 ( .A(c7890), .B(b[7890]), .Z(n23671) );
XNOR U39453 ( .A(b[7890]), .B(n23672), .Z(c[7890]) );
XNOR U39454 ( .A(a[7890]), .B(c7890), .Z(n23672) );
XOR U39455 ( .A(c7891), .B(n23673), .Z(c7892) );
ANDN U39456 ( .B(n23674), .A(n23675), .Z(n23673) );
XOR U39457 ( .A(c7891), .B(b[7891]), .Z(n23674) );
XNOR U39458 ( .A(b[7891]), .B(n23675), .Z(c[7891]) );
XNOR U39459 ( .A(a[7891]), .B(c7891), .Z(n23675) );
XOR U39460 ( .A(c7892), .B(n23676), .Z(c7893) );
ANDN U39461 ( .B(n23677), .A(n23678), .Z(n23676) );
XOR U39462 ( .A(c7892), .B(b[7892]), .Z(n23677) );
XNOR U39463 ( .A(b[7892]), .B(n23678), .Z(c[7892]) );
XNOR U39464 ( .A(a[7892]), .B(c7892), .Z(n23678) );
XOR U39465 ( .A(c7893), .B(n23679), .Z(c7894) );
ANDN U39466 ( .B(n23680), .A(n23681), .Z(n23679) );
XOR U39467 ( .A(c7893), .B(b[7893]), .Z(n23680) );
XNOR U39468 ( .A(b[7893]), .B(n23681), .Z(c[7893]) );
XNOR U39469 ( .A(a[7893]), .B(c7893), .Z(n23681) );
XOR U39470 ( .A(c7894), .B(n23682), .Z(c7895) );
ANDN U39471 ( .B(n23683), .A(n23684), .Z(n23682) );
XOR U39472 ( .A(c7894), .B(b[7894]), .Z(n23683) );
XNOR U39473 ( .A(b[7894]), .B(n23684), .Z(c[7894]) );
XNOR U39474 ( .A(a[7894]), .B(c7894), .Z(n23684) );
XOR U39475 ( .A(c7895), .B(n23685), .Z(c7896) );
ANDN U39476 ( .B(n23686), .A(n23687), .Z(n23685) );
XOR U39477 ( .A(c7895), .B(b[7895]), .Z(n23686) );
XNOR U39478 ( .A(b[7895]), .B(n23687), .Z(c[7895]) );
XNOR U39479 ( .A(a[7895]), .B(c7895), .Z(n23687) );
XOR U39480 ( .A(c7896), .B(n23688), .Z(c7897) );
ANDN U39481 ( .B(n23689), .A(n23690), .Z(n23688) );
XOR U39482 ( .A(c7896), .B(b[7896]), .Z(n23689) );
XNOR U39483 ( .A(b[7896]), .B(n23690), .Z(c[7896]) );
XNOR U39484 ( .A(a[7896]), .B(c7896), .Z(n23690) );
XOR U39485 ( .A(c7897), .B(n23691), .Z(c7898) );
ANDN U39486 ( .B(n23692), .A(n23693), .Z(n23691) );
XOR U39487 ( .A(c7897), .B(b[7897]), .Z(n23692) );
XNOR U39488 ( .A(b[7897]), .B(n23693), .Z(c[7897]) );
XNOR U39489 ( .A(a[7897]), .B(c7897), .Z(n23693) );
XOR U39490 ( .A(c7898), .B(n23694), .Z(c7899) );
ANDN U39491 ( .B(n23695), .A(n23696), .Z(n23694) );
XOR U39492 ( .A(c7898), .B(b[7898]), .Z(n23695) );
XNOR U39493 ( .A(b[7898]), .B(n23696), .Z(c[7898]) );
XNOR U39494 ( .A(a[7898]), .B(c7898), .Z(n23696) );
XOR U39495 ( .A(c7899), .B(n23697), .Z(c7900) );
ANDN U39496 ( .B(n23698), .A(n23699), .Z(n23697) );
XOR U39497 ( .A(c7899), .B(b[7899]), .Z(n23698) );
XNOR U39498 ( .A(b[7899]), .B(n23699), .Z(c[7899]) );
XNOR U39499 ( .A(a[7899]), .B(c7899), .Z(n23699) );
XOR U39500 ( .A(c7900), .B(n23700), .Z(c7901) );
ANDN U39501 ( .B(n23701), .A(n23702), .Z(n23700) );
XOR U39502 ( .A(c7900), .B(b[7900]), .Z(n23701) );
XNOR U39503 ( .A(b[7900]), .B(n23702), .Z(c[7900]) );
XNOR U39504 ( .A(a[7900]), .B(c7900), .Z(n23702) );
XOR U39505 ( .A(c7901), .B(n23703), .Z(c7902) );
ANDN U39506 ( .B(n23704), .A(n23705), .Z(n23703) );
XOR U39507 ( .A(c7901), .B(b[7901]), .Z(n23704) );
XNOR U39508 ( .A(b[7901]), .B(n23705), .Z(c[7901]) );
XNOR U39509 ( .A(a[7901]), .B(c7901), .Z(n23705) );
XOR U39510 ( .A(c7902), .B(n23706), .Z(c7903) );
ANDN U39511 ( .B(n23707), .A(n23708), .Z(n23706) );
XOR U39512 ( .A(c7902), .B(b[7902]), .Z(n23707) );
XNOR U39513 ( .A(b[7902]), .B(n23708), .Z(c[7902]) );
XNOR U39514 ( .A(a[7902]), .B(c7902), .Z(n23708) );
XOR U39515 ( .A(c7903), .B(n23709), .Z(c7904) );
ANDN U39516 ( .B(n23710), .A(n23711), .Z(n23709) );
XOR U39517 ( .A(c7903), .B(b[7903]), .Z(n23710) );
XNOR U39518 ( .A(b[7903]), .B(n23711), .Z(c[7903]) );
XNOR U39519 ( .A(a[7903]), .B(c7903), .Z(n23711) );
XOR U39520 ( .A(c7904), .B(n23712), .Z(c7905) );
ANDN U39521 ( .B(n23713), .A(n23714), .Z(n23712) );
XOR U39522 ( .A(c7904), .B(b[7904]), .Z(n23713) );
XNOR U39523 ( .A(b[7904]), .B(n23714), .Z(c[7904]) );
XNOR U39524 ( .A(a[7904]), .B(c7904), .Z(n23714) );
XOR U39525 ( .A(c7905), .B(n23715), .Z(c7906) );
ANDN U39526 ( .B(n23716), .A(n23717), .Z(n23715) );
XOR U39527 ( .A(c7905), .B(b[7905]), .Z(n23716) );
XNOR U39528 ( .A(b[7905]), .B(n23717), .Z(c[7905]) );
XNOR U39529 ( .A(a[7905]), .B(c7905), .Z(n23717) );
XOR U39530 ( .A(c7906), .B(n23718), .Z(c7907) );
ANDN U39531 ( .B(n23719), .A(n23720), .Z(n23718) );
XOR U39532 ( .A(c7906), .B(b[7906]), .Z(n23719) );
XNOR U39533 ( .A(b[7906]), .B(n23720), .Z(c[7906]) );
XNOR U39534 ( .A(a[7906]), .B(c7906), .Z(n23720) );
XOR U39535 ( .A(c7907), .B(n23721), .Z(c7908) );
ANDN U39536 ( .B(n23722), .A(n23723), .Z(n23721) );
XOR U39537 ( .A(c7907), .B(b[7907]), .Z(n23722) );
XNOR U39538 ( .A(b[7907]), .B(n23723), .Z(c[7907]) );
XNOR U39539 ( .A(a[7907]), .B(c7907), .Z(n23723) );
XOR U39540 ( .A(c7908), .B(n23724), .Z(c7909) );
ANDN U39541 ( .B(n23725), .A(n23726), .Z(n23724) );
XOR U39542 ( .A(c7908), .B(b[7908]), .Z(n23725) );
XNOR U39543 ( .A(b[7908]), .B(n23726), .Z(c[7908]) );
XNOR U39544 ( .A(a[7908]), .B(c7908), .Z(n23726) );
XOR U39545 ( .A(c7909), .B(n23727), .Z(c7910) );
ANDN U39546 ( .B(n23728), .A(n23729), .Z(n23727) );
XOR U39547 ( .A(c7909), .B(b[7909]), .Z(n23728) );
XNOR U39548 ( .A(b[7909]), .B(n23729), .Z(c[7909]) );
XNOR U39549 ( .A(a[7909]), .B(c7909), .Z(n23729) );
XOR U39550 ( .A(c7910), .B(n23730), .Z(c7911) );
ANDN U39551 ( .B(n23731), .A(n23732), .Z(n23730) );
XOR U39552 ( .A(c7910), .B(b[7910]), .Z(n23731) );
XNOR U39553 ( .A(b[7910]), .B(n23732), .Z(c[7910]) );
XNOR U39554 ( .A(a[7910]), .B(c7910), .Z(n23732) );
XOR U39555 ( .A(c7911), .B(n23733), .Z(c7912) );
ANDN U39556 ( .B(n23734), .A(n23735), .Z(n23733) );
XOR U39557 ( .A(c7911), .B(b[7911]), .Z(n23734) );
XNOR U39558 ( .A(b[7911]), .B(n23735), .Z(c[7911]) );
XNOR U39559 ( .A(a[7911]), .B(c7911), .Z(n23735) );
XOR U39560 ( .A(c7912), .B(n23736), .Z(c7913) );
ANDN U39561 ( .B(n23737), .A(n23738), .Z(n23736) );
XOR U39562 ( .A(c7912), .B(b[7912]), .Z(n23737) );
XNOR U39563 ( .A(b[7912]), .B(n23738), .Z(c[7912]) );
XNOR U39564 ( .A(a[7912]), .B(c7912), .Z(n23738) );
XOR U39565 ( .A(c7913), .B(n23739), .Z(c7914) );
ANDN U39566 ( .B(n23740), .A(n23741), .Z(n23739) );
XOR U39567 ( .A(c7913), .B(b[7913]), .Z(n23740) );
XNOR U39568 ( .A(b[7913]), .B(n23741), .Z(c[7913]) );
XNOR U39569 ( .A(a[7913]), .B(c7913), .Z(n23741) );
XOR U39570 ( .A(c7914), .B(n23742), .Z(c7915) );
ANDN U39571 ( .B(n23743), .A(n23744), .Z(n23742) );
XOR U39572 ( .A(c7914), .B(b[7914]), .Z(n23743) );
XNOR U39573 ( .A(b[7914]), .B(n23744), .Z(c[7914]) );
XNOR U39574 ( .A(a[7914]), .B(c7914), .Z(n23744) );
XOR U39575 ( .A(c7915), .B(n23745), .Z(c7916) );
ANDN U39576 ( .B(n23746), .A(n23747), .Z(n23745) );
XOR U39577 ( .A(c7915), .B(b[7915]), .Z(n23746) );
XNOR U39578 ( .A(b[7915]), .B(n23747), .Z(c[7915]) );
XNOR U39579 ( .A(a[7915]), .B(c7915), .Z(n23747) );
XOR U39580 ( .A(c7916), .B(n23748), .Z(c7917) );
ANDN U39581 ( .B(n23749), .A(n23750), .Z(n23748) );
XOR U39582 ( .A(c7916), .B(b[7916]), .Z(n23749) );
XNOR U39583 ( .A(b[7916]), .B(n23750), .Z(c[7916]) );
XNOR U39584 ( .A(a[7916]), .B(c7916), .Z(n23750) );
XOR U39585 ( .A(c7917), .B(n23751), .Z(c7918) );
ANDN U39586 ( .B(n23752), .A(n23753), .Z(n23751) );
XOR U39587 ( .A(c7917), .B(b[7917]), .Z(n23752) );
XNOR U39588 ( .A(b[7917]), .B(n23753), .Z(c[7917]) );
XNOR U39589 ( .A(a[7917]), .B(c7917), .Z(n23753) );
XOR U39590 ( .A(c7918), .B(n23754), .Z(c7919) );
ANDN U39591 ( .B(n23755), .A(n23756), .Z(n23754) );
XOR U39592 ( .A(c7918), .B(b[7918]), .Z(n23755) );
XNOR U39593 ( .A(b[7918]), .B(n23756), .Z(c[7918]) );
XNOR U39594 ( .A(a[7918]), .B(c7918), .Z(n23756) );
XOR U39595 ( .A(c7919), .B(n23757), .Z(c7920) );
ANDN U39596 ( .B(n23758), .A(n23759), .Z(n23757) );
XOR U39597 ( .A(c7919), .B(b[7919]), .Z(n23758) );
XNOR U39598 ( .A(b[7919]), .B(n23759), .Z(c[7919]) );
XNOR U39599 ( .A(a[7919]), .B(c7919), .Z(n23759) );
XOR U39600 ( .A(c7920), .B(n23760), .Z(c7921) );
ANDN U39601 ( .B(n23761), .A(n23762), .Z(n23760) );
XOR U39602 ( .A(c7920), .B(b[7920]), .Z(n23761) );
XNOR U39603 ( .A(b[7920]), .B(n23762), .Z(c[7920]) );
XNOR U39604 ( .A(a[7920]), .B(c7920), .Z(n23762) );
XOR U39605 ( .A(c7921), .B(n23763), .Z(c7922) );
ANDN U39606 ( .B(n23764), .A(n23765), .Z(n23763) );
XOR U39607 ( .A(c7921), .B(b[7921]), .Z(n23764) );
XNOR U39608 ( .A(b[7921]), .B(n23765), .Z(c[7921]) );
XNOR U39609 ( .A(a[7921]), .B(c7921), .Z(n23765) );
XOR U39610 ( .A(c7922), .B(n23766), .Z(c7923) );
ANDN U39611 ( .B(n23767), .A(n23768), .Z(n23766) );
XOR U39612 ( .A(c7922), .B(b[7922]), .Z(n23767) );
XNOR U39613 ( .A(b[7922]), .B(n23768), .Z(c[7922]) );
XNOR U39614 ( .A(a[7922]), .B(c7922), .Z(n23768) );
XOR U39615 ( .A(c7923), .B(n23769), .Z(c7924) );
ANDN U39616 ( .B(n23770), .A(n23771), .Z(n23769) );
XOR U39617 ( .A(c7923), .B(b[7923]), .Z(n23770) );
XNOR U39618 ( .A(b[7923]), .B(n23771), .Z(c[7923]) );
XNOR U39619 ( .A(a[7923]), .B(c7923), .Z(n23771) );
XOR U39620 ( .A(c7924), .B(n23772), .Z(c7925) );
ANDN U39621 ( .B(n23773), .A(n23774), .Z(n23772) );
XOR U39622 ( .A(c7924), .B(b[7924]), .Z(n23773) );
XNOR U39623 ( .A(b[7924]), .B(n23774), .Z(c[7924]) );
XNOR U39624 ( .A(a[7924]), .B(c7924), .Z(n23774) );
XOR U39625 ( .A(c7925), .B(n23775), .Z(c7926) );
ANDN U39626 ( .B(n23776), .A(n23777), .Z(n23775) );
XOR U39627 ( .A(c7925), .B(b[7925]), .Z(n23776) );
XNOR U39628 ( .A(b[7925]), .B(n23777), .Z(c[7925]) );
XNOR U39629 ( .A(a[7925]), .B(c7925), .Z(n23777) );
XOR U39630 ( .A(c7926), .B(n23778), .Z(c7927) );
ANDN U39631 ( .B(n23779), .A(n23780), .Z(n23778) );
XOR U39632 ( .A(c7926), .B(b[7926]), .Z(n23779) );
XNOR U39633 ( .A(b[7926]), .B(n23780), .Z(c[7926]) );
XNOR U39634 ( .A(a[7926]), .B(c7926), .Z(n23780) );
XOR U39635 ( .A(c7927), .B(n23781), .Z(c7928) );
ANDN U39636 ( .B(n23782), .A(n23783), .Z(n23781) );
XOR U39637 ( .A(c7927), .B(b[7927]), .Z(n23782) );
XNOR U39638 ( .A(b[7927]), .B(n23783), .Z(c[7927]) );
XNOR U39639 ( .A(a[7927]), .B(c7927), .Z(n23783) );
XOR U39640 ( .A(c7928), .B(n23784), .Z(c7929) );
ANDN U39641 ( .B(n23785), .A(n23786), .Z(n23784) );
XOR U39642 ( .A(c7928), .B(b[7928]), .Z(n23785) );
XNOR U39643 ( .A(b[7928]), .B(n23786), .Z(c[7928]) );
XNOR U39644 ( .A(a[7928]), .B(c7928), .Z(n23786) );
XOR U39645 ( .A(c7929), .B(n23787), .Z(c7930) );
ANDN U39646 ( .B(n23788), .A(n23789), .Z(n23787) );
XOR U39647 ( .A(c7929), .B(b[7929]), .Z(n23788) );
XNOR U39648 ( .A(b[7929]), .B(n23789), .Z(c[7929]) );
XNOR U39649 ( .A(a[7929]), .B(c7929), .Z(n23789) );
XOR U39650 ( .A(c7930), .B(n23790), .Z(c7931) );
ANDN U39651 ( .B(n23791), .A(n23792), .Z(n23790) );
XOR U39652 ( .A(c7930), .B(b[7930]), .Z(n23791) );
XNOR U39653 ( .A(b[7930]), .B(n23792), .Z(c[7930]) );
XNOR U39654 ( .A(a[7930]), .B(c7930), .Z(n23792) );
XOR U39655 ( .A(c7931), .B(n23793), .Z(c7932) );
ANDN U39656 ( .B(n23794), .A(n23795), .Z(n23793) );
XOR U39657 ( .A(c7931), .B(b[7931]), .Z(n23794) );
XNOR U39658 ( .A(b[7931]), .B(n23795), .Z(c[7931]) );
XNOR U39659 ( .A(a[7931]), .B(c7931), .Z(n23795) );
XOR U39660 ( .A(c7932), .B(n23796), .Z(c7933) );
ANDN U39661 ( .B(n23797), .A(n23798), .Z(n23796) );
XOR U39662 ( .A(c7932), .B(b[7932]), .Z(n23797) );
XNOR U39663 ( .A(b[7932]), .B(n23798), .Z(c[7932]) );
XNOR U39664 ( .A(a[7932]), .B(c7932), .Z(n23798) );
XOR U39665 ( .A(c7933), .B(n23799), .Z(c7934) );
ANDN U39666 ( .B(n23800), .A(n23801), .Z(n23799) );
XOR U39667 ( .A(c7933), .B(b[7933]), .Z(n23800) );
XNOR U39668 ( .A(b[7933]), .B(n23801), .Z(c[7933]) );
XNOR U39669 ( .A(a[7933]), .B(c7933), .Z(n23801) );
XOR U39670 ( .A(c7934), .B(n23802), .Z(c7935) );
ANDN U39671 ( .B(n23803), .A(n23804), .Z(n23802) );
XOR U39672 ( .A(c7934), .B(b[7934]), .Z(n23803) );
XNOR U39673 ( .A(b[7934]), .B(n23804), .Z(c[7934]) );
XNOR U39674 ( .A(a[7934]), .B(c7934), .Z(n23804) );
XOR U39675 ( .A(c7935), .B(n23805), .Z(c7936) );
ANDN U39676 ( .B(n23806), .A(n23807), .Z(n23805) );
XOR U39677 ( .A(c7935), .B(b[7935]), .Z(n23806) );
XNOR U39678 ( .A(b[7935]), .B(n23807), .Z(c[7935]) );
XNOR U39679 ( .A(a[7935]), .B(c7935), .Z(n23807) );
XOR U39680 ( .A(c7936), .B(n23808), .Z(c7937) );
ANDN U39681 ( .B(n23809), .A(n23810), .Z(n23808) );
XOR U39682 ( .A(c7936), .B(b[7936]), .Z(n23809) );
XNOR U39683 ( .A(b[7936]), .B(n23810), .Z(c[7936]) );
XNOR U39684 ( .A(a[7936]), .B(c7936), .Z(n23810) );
XOR U39685 ( .A(c7937), .B(n23811), .Z(c7938) );
ANDN U39686 ( .B(n23812), .A(n23813), .Z(n23811) );
XOR U39687 ( .A(c7937), .B(b[7937]), .Z(n23812) );
XNOR U39688 ( .A(b[7937]), .B(n23813), .Z(c[7937]) );
XNOR U39689 ( .A(a[7937]), .B(c7937), .Z(n23813) );
XOR U39690 ( .A(c7938), .B(n23814), .Z(c7939) );
ANDN U39691 ( .B(n23815), .A(n23816), .Z(n23814) );
XOR U39692 ( .A(c7938), .B(b[7938]), .Z(n23815) );
XNOR U39693 ( .A(b[7938]), .B(n23816), .Z(c[7938]) );
XNOR U39694 ( .A(a[7938]), .B(c7938), .Z(n23816) );
XOR U39695 ( .A(c7939), .B(n23817), .Z(c7940) );
ANDN U39696 ( .B(n23818), .A(n23819), .Z(n23817) );
XOR U39697 ( .A(c7939), .B(b[7939]), .Z(n23818) );
XNOR U39698 ( .A(b[7939]), .B(n23819), .Z(c[7939]) );
XNOR U39699 ( .A(a[7939]), .B(c7939), .Z(n23819) );
XOR U39700 ( .A(c7940), .B(n23820), .Z(c7941) );
ANDN U39701 ( .B(n23821), .A(n23822), .Z(n23820) );
XOR U39702 ( .A(c7940), .B(b[7940]), .Z(n23821) );
XNOR U39703 ( .A(b[7940]), .B(n23822), .Z(c[7940]) );
XNOR U39704 ( .A(a[7940]), .B(c7940), .Z(n23822) );
XOR U39705 ( .A(c7941), .B(n23823), .Z(c7942) );
ANDN U39706 ( .B(n23824), .A(n23825), .Z(n23823) );
XOR U39707 ( .A(c7941), .B(b[7941]), .Z(n23824) );
XNOR U39708 ( .A(b[7941]), .B(n23825), .Z(c[7941]) );
XNOR U39709 ( .A(a[7941]), .B(c7941), .Z(n23825) );
XOR U39710 ( .A(c7942), .B(n23826), .Z(c7943) );
ANDN U39711 ( .B(n23827), .A(n23828), .Z(n23826) );
XOR U39712 ( .A(c7942), .B(b[7942]), .Z(n23827) );
XNOR U39713 ( .A(b[7942]), .B(n23828), .Z(c[7942]) );
XNOR U39714 ( .A(a[7942]), .B(c7942), .Z(n23828) );
XOR U39715 ( .A(c7943), .B(n23829), .Z(c7944) );
ANDN U39716 ( .B(n23830), .A(n23831), .Z(n23829) );
XOR U39717 ( .A(c7943), .B(b[7943]), .Z(n23830) );
XNOR U39718 ( .A(b[7943]), .B(n23831), .Z(c[7943]) );
XNOR U39719 ( .A(a[7943]), .B(c7943), .Z(n23831) );
XOR U39720 ( .A(c7944), .B(n23832), .Z(c7945) );
ANDN U39721 ( .B(n23833), .A(n23834), .Z(n23832) );
XOR U39722 ( .A(c7944), .B(b[7944]), .Z(n23833) );
XNOR U39723 ( .A(b[7944]), .B(n23834), .Z(c[7944]) );
XNOR U39724 ( .A(a[7944]), .B(c7944), .Z(n23834) );
XOR U39725 ( .A(c7945), .B(n23835), .Z(c7946) );
ANDN U39726 ( .B(n23836), .A(n23837), .Z(n23835) );
XOR U39727 ( .A(c7945), .B(b[7945]), .Z(n23836) );
XNOR U39728 ( .A(b[7945]), .B(n23837), .Z(c[7945]) );
XNOR U39729 ( .A(a[7945]), .B(c7945), .Z(n23837) );
XOR U39730 ( .A(c7946), .B(n23838), .Z(c7947) );
ANDN U39731 ( .B(n23839), .A(n23840), .Z(n23838) );
XOR U39732 ( .A(c7946), .B(b[7946]), .Z(n23839) );
XNOR U39733 ( .A(b[7946]), .B(n23840), .Z(c[7946]) );
XNOR U39734 ( .A(a[7946]), .B(c7946), .Z(n23840) );
XOR U39735 ( .A(c7947), .B(n23841), .Z(c7948) );
ANDN U39736 ( .B(n23842), .A(n23843), .Z(n23841) );
XOR U39737 ( .A(c7947), .B(b[7947]), .Z(n23842) );
XNOR U39738 ( .A(b[7947]), .B(n23843), .Z(c[7947]) );
XNOR U39739 ( .A(a[7947]), .B(c7947), .Z(n23843) );
XOR U39740 ( .A(c7948), .B(n23844), .Z(c7949) );
ANDN U39741 ( .B(n23845), .A(n23846), .Z(n23844) );
XOR U39742 ( .A(c7948), .B(b[7948]), .Z(n23845) );
XNOR U39743 ( .A(b[7948]), .B(n23846), .Z(c[7948]) );
XNOR U39744 ( .A(a[7948]), .B(c7948), .Z(n23846) );
XOR U39745 ( .A(c7949), .B(n23847), .Z(c7950) );
ANDN U39746 ( .B(n23848), .A(n23849), .Z(n23847) );
XOR U39747 ( .A(c7949), .B(b[7949]), .Z(n23848) );
XNOR U39748 ( .A(b[7949]), .B(n23849), .Z(c[7949]) );
XNOR U39749 ( .A(a[7949]), .B(c7949), .Z(n23849) );
XOR U39750 ( .A(c7950), .B(n23850), .Z(c7951) );
ANDN U39751 ( .B(n23851), .A(n23852), .Z(n23850) );
XOR U39752 ( .A(c7950), .B(b[7950]), .Z(n23851) );
XNOR U39753 ( .A(b[7950]), .B(n23852), .Z(c[7950]) );
XNOR U39754 ( .A(a[7950]), .B(c7950), .Z(n23852) );
XOR U39755 ( .A(c7951), .B(n23853), .Z(c7952) );
ANDN U39756 ( .B(n23854), .A(n23855), .Z(n23853) );
XOR U39757 ( .A(c7951), .B(b[7951]), .Z(n23854) );
XNOR U39758 ( .A(b[7951]), .B(n23855), .Z(c[7951]) );
XNOR U39759 ( .A(a[7951]), .B(c7951), .Z(n23855) );
XOR U39760 ( .A(c7952), .B(n23856), .Z(c7953) );
ANDN U39761 ( .B(n23857), .A(n23858), .Z(n23856) );
XOR U39762 ( .A(c7952), .B(b[7952]), .Z(n23857) );
XNOR U39763 ( .A(b[7952]), .B(n23858), .Z(c[7952]) );
XNOR U39764 ( .A(a[7952]), .B(c7952), .Z(n23858) );
XOR U39765 ( .A(c7953), .B(n23859), .Z(c7954) );
ANDN U39766 ( .B(n23860), .A(n23861), .Z(n23859) );
XOR U39767 ( .A(c7953), .B(b[7953]), .Z(n23860) );
XNOR U39768 ( .A(b[7953]), .B(n23861), .Z(c[7953]) );
XNOR U39769 ( .A(a[7953]), .B(c7953), .Z(n23861) );
XOR U39770 ( .A(c7954), .B(n23862), .Z(c7955) );
ANDN U39771 ( .B(n23863), .A(n23864), .Z(n23862) );
XOR U39772 ( .A(c7954), .B(b[7954]), .Z(n23863) );
XNOR U39773 ( .A(b[7954]), .B(n23864), .Z(c[7954]) );
XNOR U39774 ( .A(a[7954]), .B(c7954), .Z(n23864) );
XOR U39775 ( .A(c7955), .B(n23865), .Z(c7956) );
ANDN U39776 ( .B(n23866), .A(n23867), .Z(n23865) );
XOR U39777 ( .A(c7955), .B(b[7955]), .Z(n23866) );
XNOR U39778 ( .A(b[7955]), .B(n23867), .Z(c[7955]) );
XNOR U39779 ( .A(a[7955]), .B(c7955), .Z(n23867) );
XOR U39780 ( .A(c7956), .B(n23868), .Z(c7957) );
ANDN U39781 ( .B(n23869), .A(n23870), .Z(n23868) );
XOR U39782 ( .A(c7956), .B(b[7956]), .Z(n23869) );
XNOR U39783 ( .A(b[7956]), .B(n23870), .Z(c[7956]) );
XNOR U39784 ( .A(a[7956]), .B(c7956), .Z(n23870) );
XOR U39785 ( .A(c7957), .B(n23871), .Z(c7958) );
ANDN U39786 ( .B(n23872), .A(n23873), .Z(n23871) );
XOR U39787 ( .A(c7957), .B(b[7957]), .Z(n23872) );
XNOR U39788 ( .A(b[7957]), .B(n23873), .Z(c[7957]) );
XNOR U39789 ( .A(a[7957]), .B(c7957), .Z(n23873) );
XOR U39790 ( .A(c7958), .B(n23874), .Z(c7959) );
ANDN U39791 ( .B(n23875), .A(n23876), .Z(n23874) );
XOR U39792 ( .A(c7958), .B(b[7958]), .Z(n23875) );
XNOR U39793 ( .A(b[7958]), .B(n23876), .Z(c[7958]) );
XNOR U39794 ( .A(a[7958]), .B(c7958), .Z(n23876) );
XOR U39795 ( .A(c7959), .B(n23877), .Z(c7960) );
ANDN U39796 ( .B(n23878), .A(n23879), .Z(n23877) );
XOR U39797 ( .A(c7959), .B(b[7959]), .Z(n23878) );
XNOR U39798 ( .A(b[7959]), .B(n23879), .Z(c[7959]) );
XNOR U39799 ( .A(a[7959]), .B(c7959), .Z(n23879) );
XOR U39800 ( .A(c7960), .B(n23880), .Z(c7961) );
ANDN U39801 ( .B(n23881), .A(n23882), .Z(n23880) );
XOR U39802 ( .A(c7960), .B(b[7960]), .Z(n23881) );
XNOR U39803 ( .A(b[7960]), .B(n23882), .Z(c[7960]) );
XNOR U39804 ( .A(a[7960]), .B(c7960), .Z(n23882) );
XOR U39805 ( .A(c7961), .B(n23883), .Z(c7962) );
ANDN U39806 ( .B(n23884), .A(n23885), .Z(n23883) );
XOR U39807 ( .A(c7961), .B(b[7961]), .Z(n23884) );
XNOR U39808 ( .A(b[7961]), .B(n23885), .Z(c[7961]) );
XNOR U39809 ( .A(a[7961]), .B(c7961), .Z(n23885) );
XOR U39810 ( .A(c7962), .B(n23886), .Z(c7963) );
ANDN U39811 ( .B(n23887), .A(n23888), .Z(n23886) );
XOR U39812 ( .A(c7962), .B(b[7962]), .Z(n23887) );
XNOR U39813 ( .A(b[7962]), .B(n23888), .Z(c[7962]) );
XNOR U39814 ( .A(a[7962]), .B(c7962), .Z(n23888) );
XOR U39815 ( .A(c7963), .B(n23889), .Z(c7964) );
ANDN U39816 ( .B(n23890), .A(n23891), .Z(n23889) );
XOR U39817 ( .A(c7963), .B(b[7963]), .Z(n23890) );
XNOR U39818 ( .A(b[7963]), .B(n23891), .Z(c[7963]) );
XNOR U39819 ( .A(a[7963]), .B(c7963), .Z(n23891) );
XOR U39820 ( .A(c7964), .B(n23892), .Z(c7965) );
ANDN U39821 ( .B(n23893), .A(n23894), .Z(n23892) );
XOR U39822 ( .A(c7964), .B(b[7964]), .Z(n23893) );
XNOR U39823 ( .A(b[7964]), .B(n23894), .Z(c[7964]) );
XNOR U39824 ( .A(a[7964]), .B(c7964), .Z(n23894) );
XOR U39825 ( .A(c7965), .B(n23895), .Z(c7966) );
ANDN U39826 ( .B(n23896), .A(n23897), .Z(n23895) );
XOR U39827 ( .A(c7965), .B(b[7965]), .Z(n23896) );
XNOR U39828 ( .A(b[7965]), .B(n23897), .Z(c[7965]) );
XNOR U39829 ( .A(a[7965]), .B(c7965), .Z(n23897) );
XOR U39830 ( .A(c7966), .B(n23898), .Z(c7967) );
ANDN U39831 ( .B(n23899), .A(n23900), .Z(n23898) );
XOR U39832 ( .A(c7966), .B(b[7966]), .Z(n23899) );
XNOR U39833 ( .A(b[7966]), .B(n23900), .Z(c[7966]) );
XNOR U39834 ( .A(a[7966]), .B(c7966), .Z(n23900) );
XOR U39835 ( .A(c7967), .B(n23901), .Z(c7968) );
ANDN U39836 ( .B(n23902), .A(n23903), .Z(n23901) );
XOR U39837 ( .A(c7967), .B(b[7967]), .Z(n23902) );
XNOR U39838 ( .A(b[7967]), .B(n23903), .Z(c[7967]) );
XNOR U39839 ( .A(a[7967]), .B(c7967), .Z(n23903) );
XOR U39840 ( .A(c7968), .B(n23904), .Z(c7969) );
ANDN U39841 ( .B(n23905), .A(n23906), .Z(n23904) );
XOR U39842 ( .A(c7968), .B(b[7968]), .Z(n23905) );
XNOR U39843 ( .A(b[7968]), .B(n23906), .Z(c[7968]) );
XNOR U39844 ( .A(a[7968]), .B(c7968), .Z(n23906) );
XOR U39845 ( .A(c7969), .B(n23907), .Z(c7970) );
ANDN U39846 ( .B(n23908), .A(n23909), .Z(n23907) );
XOR U39847 ( .A(c7969), .B(b[7969]), .Z(n23908) );
XNOR U39848 ( .A(b[7969]), .B(n23909), .Z(c[7969]) );
XNOR U39849 ( .A(a[7969]), .B(c7969), .Z(n23909) );
XOR U39850 ( .A(c7970), .B(n23910), .Z(c7971) );
ANDN U39851 ( .B(n23911), .A(n23912), .Z(n23910) );
XOR U39852 ( .A(c7970), .B(b[7970]), .Z(n23911) );
XNOR U39853 ( .A(b[7970]), .B(n23912), .Z(c[7970]) );
XNOR U39854 ( .A(a[7970]), .B(c7970), .Z(n23912) );
XOR U39855 ( .A(c7971), .B(n23913), .Z(c7972) );
ANDN U39856 ( .B(n23914), .A(n23915), .Z(n23913) );
XOR U39857 ( .A(c7971), .B(b[7971]), .Z(n23914) );
XNOR U39858 ( .A(b[7971]), .B(n23915), .Z(c[7971]) );
XNOR U39859 ( .A(a[7971]), .B(c7971), .Z(n23915) );
XOR U39860 ( .A(c7972), .B(n23916), .Z(c7973) );
ANDN U39861 ( .B(n23917), .A(n23918), .Z(n23916) );
XOR U39862 ( .A(c7972), .B(b[7972]), .Z(n23917) );
XNOR U39863 ( .A(b[7972]), .B(n23918), .Z(c[7972]) );
XNOR U39864 ( .A(a[7972]), .B(c7972), .Z(n23918) );
XOR U39865 ( .A(c7973), .B(n23919), .Z(c7974) );
ANDN U39866 ( .B(n23920), .A(n23921), .Z(n23919) );
XOR U39867 ( .A(c7973), .B(b[7973]), .Z(n23920) );
XNOR U39868 ( .A(b[7973]), .B(n23921), .Z(c[7973]) );
XNOR U39869 ( .A(a[7973]), .B(c7973), .Z(n23921) );
XOR U39870 ( .A(c7974), .B(n23922), .Z(c7975) );
ANDN U39871 ( .B(n23923), .A(n23924), .Z(n23922) );
XOR U39872 ( .A(c7974), .B(b[7974]), .Z(n23923) );
XNOR U39873 ( .A(b[7974]), .B(n23924), .Z(c[7974]) );
XNOR U39874 ( .A(a[7974]), .B(c7974), .Z(n23924) );
XOR U39875 ( .A(c7975), .B(n23925), .Z(c7976) );
ANDN U39876 ( .B(n23926), .A(n23927), .Z(n23925) );
XOR U39877 ( .A(c7975), .B(b[7975]), .Z(n23926) );
XNOR U39878 ( .A(b[7975]), .B(n23927), .Z(c[7975]) );
XNOR U39879 ( .A(a[7975]), .B(c7975), .Z(n23927) );
XOR U39880 ( .A(c7976), .B(n23928), .Z(c7977) );
ANDN U39881 ( .B(n23929), .A(n23930), .Z(n23928) );
XOR U39882 ( .A(c7976), .B(b[7976]), .Z(n23929) );
XNOR U39883 ( .A(b[7976]), .B(n23930), .Z(c[7976]) );
XNOR U39884 ( .A(a[7976]), .B(c7976), .Z(n23930) );
XOR U39885 ( .A(c7977), .B(n23931), .Z(c7978) );
ANDN U39886 ( .B(n23932), .A(n23933), .Z(n23931) );
XOR U39887 ( .A(c7977), .B(b[7977]), .Z(n23932) );
XNOR U39888 ( .A(b[7977]), .B(n23933), .Z(c[7977]) );
XNOR U39889 ( .A(a[7977]), .B(c7977), .Z(n23933) );
XOR U39890 ( .A(c7978), .B(n23934), .Z(c7979) );
ANDN U39891 ( .B(n23935), .A(n23936), .Z(n23934) );
XOR U39892 ( .A(c7978), .B(b[7978]), .Z(n23935) );
XNOR U39893 ( .A(b[7978]), .B(n23936), .Z(c[7978]) );
XNOR U39894 ( .A(a[7978]), .B(c7978), .Z(n23936) );
XOR U39895 ( .A(c7979), .B(n23937), .Z(c7980) );
ANDN U39896 ( .B(n23938), .A(n23939), .Z(n23937) );
XOR U39897 ( .A(c7979), .B(b[7979]), .Z(n23938) );
XNOR U39898 ( .A(b[7979]), .B(n23939), .Z(c[7979]) );
XNOR U39899 ( .A(a[7979]), .B(c7979), .Z(n23939) );
XOR U39900 ( .A(c7980), .B(n23940), .Z(c7981) );
ANDN U39901 ( .B(n23941), .A(n23942), .Z(n23940) );
XOR U39902 ( .A(c7980), .B(b[7980]), .Z(n23941) );
XNOR U39903 ( .A(b[7980]), .B(n23942), .Z(c[7980]) );
XNOR U39904 ( .A(a[7980]), .B(c7980), .Z(n23942) );
XOR U39905 ( .A(c7981), .B(n23943), .Z(c7982) );
ANDN U39906 ( .B(n23944), .A(n23945), .Z(n23943) );
XOR U39907 ( .A(c7981), .B(b[7981]), .Z(n23944) );
XNOR U39908 ( .A(b[7981]), .B(n23945), .Z(c[7981]) );
XNOR U39909 ( .A(a[7981]), .B(c7981), .Z(n23945) );
XOR U39910 ( .A(c7982), .B(n23946), .Z(c7983) );
ANDN U39911 ( .B(n23947), .A(n23948), .Z(n23946) );
XOR U39912 ( .A(c7982), .B(b[7982]), .Z(n23947) );
XNOR U39913 ( .A(b[7982]), .B(n23948), .Z(c[7982]) );
XNOR U39914 ( .A(a[7982]), .B(c7982), .Z(n23948) );
XOR U39915 ( .A(c7983), .B(n23949), .Z(c7984) );
ANDN U39916 ( .B(n23950), .A(n23951), .Z(n23949) );
XOR U39917 ( .A(c7983), .B(b[7983]), .Z(n23950) );
XNOR U39918 ( .A(b[7983]), .B(n23951), .Z(c[7983]) );
XNOR U39919 ( .A(a[7983]), .B(c7983), .Z(n23951) );
XOR U39920 ( .A(c7984), .B(n23952), .Z(c7985) );
ANDN U39921 ( .B(n23953), .A(n23954), .Z(n23952) );
XOR U39922 ( .A(c7984), .B(b[7984]), .Z(n23953) );
XNOR U39923 ( .A(b[7984]), .B(n23954), .Z(c[7984]) );
XNOR U39924 ( .A(a[7984]), .B(c7984), .Z(n23954) );
XOR U39925 ( .A(c7985), .B(n23955), .Z(c7986) );
ANDN U39926 ( .B(n23956), .A(n23957), .Z(n23955) );
XOR U39927 ( .A(c7985), .B(b[7985]), .Z(n23956) );
XNOR U39928 ( .A(b[7985]), .B(n23957), .Z(c[7985]) );
XNOR U39929 ( .A(a[7985]), .B(c7985), .Z(n23957) );
XOR U39930 ( .A(c7986), .B(n23958), .Z(c7987) );
ANDN U39931 ( .B(n23959), .A(n23960), .Z(n23958) );
XOR U39932 ( .A(c7986), .B(b[7986]), .Z(n23959) );
XNOR U39933 ( .A(b[7986]), .B(n23960), .Z(c[7986]) );
XNOR U39934 ( .A(a[7986]), .B(c7986), .Z(n23960) );
XOR U39935 ( .A(c7987), .B(n23961), .Z(c7988) );
ANDN U39936 ( .B(n23962), .A(n23963), .Z(n23961) );
XOR U39937 ( .A(c7987), .B(b[7987]), .Z(n23962) );
XNOR U39938 ( .A(b[7987]), .B(n23963), .Z(c[7987]) );
XNOR U39939 ( .A(a[7987]), .B(c7987), .Z(n23963) );
XOR U39940 ( .A(c7988), .B(n23964), .Z(c7989) );
ANDN U39941 ( .B(n23965), .A(n23966), .Z(n23964) );
XOR U39942 ( .A(c7988), .B(b[7988]), .Z(n23965) );
XNOR U39943 ( .A(b[7988]), .B(n23966), .Z(c[7988]) );
XNOR U39944 ( .A(a[7988]), .B(c7988), .Z(n23966) );
XOR U39945 ( .A(c7989), .B(n23967), .Z(c7990) );
ANDN U39946 ( .B(n23968), .A(n23969), .Z(n23967) );
XOR U39947 ( .A(c7989), .B(b[7989]), .Z(n23968) );
XNOR U39948 ( .A(b[7989]), .B(n23969), .Z(c[7989]) );
XNOR U39949 ( .A(a[7989]), .B(c7989), .Z(n23969) );
XOR U39950 ( .A(c7990), .B(n23970), .Z(c7991) );
ANDN U39951 ( .B(n23971), .A(n23972), .Z(n23970) );
XOR U39952 ( .A(c7990), .B(b[7990]), .Z(n23971) );
XNOR U39953 ( .A(b[7990]), .B(n23972), .Z(c[7990]) );
XNOR U39954 ( .A(a[7990]), .B(c7990), .Z(n23972) );
XOR U39955 ( .A(c7991), .B(n23973), .Z(c7992) );
ANDN U39956 ( .B(n23974), .A(n23975), .Z(n23973) );
XOR U39957 ( .A(c7991), .B(b[7991]), .Z(n23974) );
XNOR U39958 ( .A(b[7991]), .B(n23975), .Z(c[7991]) );
XNOR U39959 ( .A(a[7991]), .B(c7991), .Z(n23975) );
XOR U39960 ( .A(c7992), .B(n23976), .Z(c7993) );
ANDN U39961 ( .B(n23977), .A(n23978), .Z(n23976) );
XOR U39962 ( .A(c7992), .B(b[7992]), .Z(n23977) );
XNOR U39963 ( .A(b[7992]), .B(n23978), .Z(c[7992]) );
XNOR U39964 ( .A(a[7992]), .B(c7992), .Z(n23978) );
XOR U39965 ( .A(c7993), .B(n23979), .Z(c7994) );
ANDN U39966 ( .B(n23980), .A(n23981), .Z(n23979) );
XOR U39967 ( .A(c7993), .B(b[7993]), .Z(n23980) );
XNOR U39968 ( .A(b[7993]), .B(n23981), .Z(c[7993]) );
XNOR U39969 ( .A(a[7993]), .B(c7993), .Z(n23981) );
XOR U39970 ( .A(c7994), .B(n23982), .Z(c7995) );
ANDN U39971 ( .B(n23983), .A(n23984), .Z(n23982) );
XOR U39972 ( .A(c7994), .B(b[7994]), .Z(n23983) );
XNOR U39973 ( .A(b[7994]), .B(n23984), .Z(c[7994]) );
XNOR U39974 ( .A(a[7994]), .B(c7994), .Z(n23984) );
XOR U39975 ( .A(c7995), .B(n23985), .Z(c7996) );
ANDN U39976 ( .B(n23986), .A(n23987), .Z(n23985) );
XOR U39977 ( .A(c7995), .B(b[7995]), .Z(n23986) );
XNOR U39978 ( .A(b[7995]), .B(n23987), .Z(c[7995]) );
XNOR U39979 ( .A(a[7995]), .B(c7995), .Z(n23987) );
XOR U39980 ( .A(c7996), .B(n23988), .Z(c7997) );
ANDN U39981 ( .B(n23989), .A(n23990), .Z(n23988) );
XOR U39982 ( .A(c7996), .B(b[7996]), .Z(n23989) );
XNOR U39983 ( .A(b[7996]), .B(n23990), .Z(c[7996]) );
XNOR U39984 ( .A(a[7996]), .B(c7996), .Z(n23990) );
XOR U39985 ( .A(c7997), .B(n23991), .Z(c7998) );
ANDN U39986 ( .B(n23992), .A(n23993), .Z(n23991) );
XOR U39987 ( .A(c7997), .B(b[7997]), .Z(n23992) );
XNOR U39988 ( .A(b[7997]), .B(n23993), .Z(c[7997]) );
XNOR U39989 ( .A(a[7997]), .B(c7997), .Z(n23993) );
XOR U39990 ( .A(c7998), .B(n23994), .Z(c7999) );
ANDN U39991 ( .B(n23995), .A(n23996), .Z(n23994) );
XOR U39992 ( .A(c7998), .B(b[7998]), .Z(n23995) );
XNOR U39993 ( .A(b[7998]), .B(n23996), .Z(c[7998]) );
XNOR U39994 ( .A(a[7998]), .B(c7998), .Z(n23996) );
XOR U39995 ( .A(c7999), .B(n23997), .Z(c8000) );
ANDN U39996 ( .B(n23998), .A(n23999), .Z(n23997) );
XOR U39997 ( .A(c7999), .B(b[7999]), .Z(n23998) );
XNOR U39998 ( .A(b[7999]), .B(n23999), .Z(c[7999]) );
XNOR U39999 ( .A(a[7999]), .B(c7999), .Z(n23999) );
XOR U40000 ( .A(c8000), .B(n24000), .Z(c8001) );
ANDN U40001 ( .B(n24001), .A(n24002), .Z(n24000) );
XOR U40002 ( .A(c8000), .B(b[8000]), .Z(n24001) );
XNOR U40003 ( .A(b[8000]), .B(n24002), .Z(c[8000]) );
XNOR U40004 ( .A(a[8000]), .B(c8000), .Z(n24002) );
XOR U40005 ( .A(c8001), .B(n24003), .Z(c8002) );
ANDN U40006 ( .B(n24004), .A(n24005), .Z(n24003) );
XOR U40007 ( .A(c8001), .B(b[8001]), .Z(n24004) );
XNOR U40008 ( .A(b[8001]), .B(n24005), .Z(c[8001]) );
XNOR U40009 ( .A(a[8001]), .B(c8001), .Z(n24005) );
XOR U40010 ( .A(c8002), .B(n24006), .Z(c8003) );
ANDN U40011 ( .B(n24007), .A(n24008), .Z(n24006) );
XOR U40012 ( .A(c8002), .B(b[8002]), .Z(n24007) );
XNOR U40013 ( .A(b[8002]), .B(n24008), .Z(c[8002]) );
XNOR U40014 ( .A(a[8002]), .B(c8002), .Z(n24008) );
XOR U40015 ( .A(c8003), .B(n24009), .Z(c8004) );
ANDN U40016 ( .B(n24010), .A(n24011), .Z(n24009) );
XOR U40017 ( .A(c8003), .B(b[8003]), .Z(n24010) );
XNOR U40018 ( .A(b[8003]), .B(n24011), .Z(c[8003]) );
XNOR U40019 ( .A(a[8003]), .B(c8003), .Z(n24011) );
XOR U40020 ( .A(c8004), .B(n24012), .Z(c8005) );
ANDN U40021 ( .B(n24013), .A(n24014), .Z(n24012) );
XOR U40022 ( .A(c8004), .B(b[8004]), .Z(n24013) );
XNOR U40023 ( .A(b[8004]), .B(n24014), .Z(c[8004]) );
XNOR U40024 ( .A(a[8004]), .B(c8004), .Z(n24014) );
XOR U40025 ( .A(c8005), .B(n24015), .Z(c8006) );
ANDN U40026 ( .B(n24016), .A(n24017), .Z(n24015) );
XOR U40027 ( .A(c8005), .B(b[8005]), .Z(n24016) );
XNOR U40028 ( .A(b[8005]), .B(n24017), .Z(c[8005]) );
XNOR U40029 ( .A(a[8005]), .B(c8005), .Z(n24017) );
XOR U40030 ( .A(c8006), .B(n24018), .Z(c8007) );
ANDN U40031 ( .B(n24019), .A(n24020), .Z(n24018) );
XOR U40032 ( .A(c8006), .B(b[8006]), .Z(n24019) );
XNOR U40033 ( .A(b[8006]), .B(n24020), .Z(c[8006]) );
XNOR U40034 ( .A(a[8006]), .B(c8006), .Z(n24020) );
XOR U40035 ( .A(c8007), .B(n24021), .Z(c8008) );
ANDN U40036 ( .B(n24022), .A(n24023), .Z(n24021) );
XOR U40037 ( .A(c8007), .B(b[8007]), .Z(n24022) );
XNOR U40038 ( .A(b[8007]), .B(n24023), .Z(c[8007]) );
XNOR U40039 ( .A(a[8007]), .B(c8007), .Z(n24023) );
XOR U40040 ( .A(c8008), .B(n24024), .Z(c8009) );
ANDN U40041 ( .B(n24025), .A(n24026), .Z(n24024) );
XOR U40042 ( .A(c8008), .B(b[8008]), .Z(n24025) );
XNOR U40043 ( .A(b[8008]), .B(n24026), .Z(c[8008]) );
XNOR U40044 ( .A(a[8008]), .B(c8008), .Z(n24026) );
XOR U40045 ( .A(c8009), .B(n24027), .Z(c8010) );
ANDN U40046 ( .B(n24028), .A(n24029), .Z(n24027) );
XOR U40047 ( .A(c8009), .B(b[8009]), .Z(n24028) );
XNOR U40048 ( .A(b[8009]), .B(n24029), .Z(c[8009]) );
XNOR U40049 ( .A(a[8009]), .B(c8009), .Z(n24029) );
XOR U40050 ( .A(c8010), .B(n24030), .Z(c8011) );
ANDN U40051 ( .B(n24031), .A(n24032), .Z(n24030) );
XOR U40052 ( .A(c8010), .B(b[8010]), .Z(n24031) );
XNOR U40053 ( .A(b[8010]), .B(n24032), .Z(c[8010]) );
XNOR U40054 ( .A(a[8010]), .B(c8010), .Z(n24032) );
XOR U40055 ( .A(c8011), .B(n24033), .Z(c8012) );
ANDN U40056 ( .B(n24034), .A(n24035), .Z(n24033) );
XOR U40057 ( .A(c8011), .B(b[8011]), .Z(n24034) );
XNOR U40058 ( .A(b[8011]), .B(n24035), .Z(c[8011]) );
XNOR U40059 ( .A(a[8011]), .B(c8011), .Z(n24035) );
XOR U40060 ( .A(c8012), .B(n24036), .Z(c8013) );
ANDN U40061 ( .B(n24037), .A(n24038), .Z(n24036) );
XOR U40062 ( .A(c8012), .B(b[8012]), .Z(n24037) );
XNOR U40063 ( .A(b[8012]), .B(n24038), .Z(c[8012]) );
XNOR U40064 ( .A(a[8012]), .B(c8012), .Z(n24038) );
XOR U40065 ( .A(c8013), .B(n24039), .Z(c8014) );
ANDN U40066 ( .B(n24040), .A(n24041), .Z(n24039) );
XOR U40067 ( .A(c8013), .B(b[8013]), .Z(n24040) );
XNOR U40068 ( .A(b[8013]), .B(n24041), .Z(c[8013]) );
XNOR U40069 ( .A(a[8013]), .B(c8013), .Z(n24041) );
XOR U40070 ( .A(c8014), .B(n24042), .Z(c8015) );
ANDN U40071 ( .B(n24043), .A(n24044), .Z(n24042) );
XOR U40072 ( .A(c8014), .B(b[8014]), .Z(n24043) );
XNOR U40073 ( .A(b[8014]), .B(n24044), .Z(c[8014]) );
XNOR U40074 ( .A(a[8014]), .B(c8014), .Z(n24044) );
XOR U40075 ( .A(c8015), .B(n24045), .Z(c8016) );
ANDN U40076 ( .B(n24046), .A(n24047), .Z(n24045) );
XOR U40077 ( .A(c8015), .B(b[8015]), .Z(n24046) );
XNOR U40078 ( .A(b[8015]), .B(n24047), .Z(c[8015]) );
XNOR U40079 ( .A(a[8015]), .B(c8015), .Z(n24047) );
XOR U40080 ( .A(c8016), .B(n24048), .Z(c8017) );
ANDN U40081 ( .B(n24049), .A(n24050), .Z(n24048) );
XOR U40082 ( .A(c8016), .B(b[8016]), .Z(n24049) );
XNOR U40083 ( .A(b[8016]), .B(n24050), .Z(c[8016]) );
XNOR U40084 ( .A(a[8016]), .B(c8016), .Z(n24050) );
XOR U40085 ( .A(c8017), .B(n24051), .Z(c8018) );
ANDN U40086 ( .B(n24052), .A(n24053), .Z(n24051) );
XOR U40087 ( .A(c8017), .B(b[8017]), .Z(n24052) );
XNOR U40088 ( .A(b[8017]), .B(n24053), .Z(c[8017]) );
XNOR U40089 ( .A(a[8017]), .B(c8017), .Z(n24053) );
XOR U40090 ( .A(c8018), .B(n24054), .Z(c8019) );
ANDN U40091 ( .B(n24055), .A(n24056), .Z(n24054) );
XOR U40092 ( .A(c8018), .B(b[8018]), .Z(n24055) );
XNOR U40093 ( .A(b[8018]), .B(n24056), .Z(c[8018]) );
XNOR U40094 ( .A(a[8018]), .B(c8018), .Z(n24056) );
XOR U40095 ( .A(c8019), .B(n24057), .Z(c8020) );
ANDN U40096 ( .B(n24058), .A(n24059), .Z(n24057) );
XOR U40097 ( .A(c8019), .B(b[8019]), .Z(n24058) );
XNOR U40098 ( .A(b[8019]), .B(n24059), .Z(c[8019]) );
XNOR U40099 ( .A(a[8019]), .B(c8019), .Z(n24059) );
XOR U40100 ( .A(c8020), .B(n24060), .Z(c8021) );
ANDN U40101 ( .B(n24061), .A(n24062), .Z(n24060) );
XOR U40102 ( .A(c8020), .B(b[8020]), .Z(n24061) );
XNOR U40103 ( .A(b[8020]), .B(n24062), .Z(c[8020]) );
XNOR U40104 ( .A(a[8020]), .B(c8020), .Z(n24062) );
XOR U40105 ( .A(c8021), .B(n24063), .Z(c8022) );
ANDN U40106 ( .B(n24064), .A(n24065), .Z(n24063) );
XOR U40107 ( .A(c8021), .B(b[8021]), .Z(n24064) );
XNOR U40108 ( .A(b[8021]), .B(n24065), .Z(c[8021]) );
XNOR U40109 ( .A(a[8021]), .B(c8021), .Z(n24065) );
XOR U40110 ( .A(c8022), .B(n24066), .Z(c8023) );
ANDN U40111 ( .B(n24067), .A(n24068), .Z(n24066) );
XOR U40112 ( .A(c8022), .B(b[8022]), .Z(n24067) );
XNOR U40113 ( .A(b[8022]), .B(n24068), .Z(c[8022]) );
XNOR U40114 ( .A(a[8022]), .B(c8022), .Z(n24068) );
XOR U40115 ( .A(c8023), .B(n24069), .Z(c8024) );
ANDN U40116 ( .B(n24070), .A(n24071), .Z(n24069) );
XOR U40117 ( .A(c8023), .B(b[8023]), .Z(n24070) );
XNOR U40118 ( .A(b[8023]), .B(n24071), .Z(c[8023]) );
XNOR U40119 ( .A(a[8023]), .B(c8023), .Z(n24071) );
XOR U40120 ( .A(c8024), .B(n24072), .Z(c8025) );
ANDN U40121 ( .B(n24073), .A(n24074), .Z(n24072) );
XOR U40122 ( .A(c8024), .B(b[8024]), .Z(n24073) );
XNOR U40123 ( .A(b[8024]), .B(n24074), .Z(c[8024]) );
XNOR U40124 ( .A(a[8024]), .B(c8024), .Z(n24074) );
XOR U40125 ( .A(c8025), .B(n24075), .Z(c8026) );
ANDN U40126 ( .B(n24076), .A(n24077), .Z(n24075) );
XOR U40127 ( .A(c8025), .B(b[8025]), .Z(n24076) );
XNOR U40128 ( .A(b[8025]), .B(n24077), .Z(c[8025]) );
XNOR U40129 ( .A(a[8025]), .B(c8025), .Z(n24077) );
XOR U40130 ( .A(c8026), .B(n24078), .Z(c8027) );
ANDN U40131 ( .B(n24079), .A(n24080), .Z(n24078) );
XOR U40132 ( .A(c8026), .B(b[8026]), .Z(n24079) );
XNOR U40133 ( .A(b[8026]), .B(n24080), .Z(c[8026]) );
XNOR U40134 ( .A(a[8026]), .B(c8026), .Z(n24080) );
XOR U40135 ( .A(c8027), .B(n24081), .Z(c8028) );
ANDN U40136 ( .B(n24082), .A(n24083), .Z(n24081) );
XOR U40137 ( .A(c8027), .B(b[8027]), .Z(n24082) );
XNOR U40138 ( .A(b[8027]), .B(n24083), .Z(c[8027]) );
XNOR U40139 ( .A(a[8027]), .B(c8027), .Z(n24083) );
XOR U40140 ( .A(c8028), .B(n24084), .Z(c8029) );
ANDN U40141 ( .B(n24085), .A(n24086), .Z(n24084) );
XOR U40142 ( .A(c8028), .B(b[8028]), .Z(n24085) );
XNOR U40143 ( .A(b[8028]), .B(n24086), .Z(c[8028]) );
XNOR U40144 ( .A(a[8028]), .B(c8028), .Z(n24086) );
XOR U40145 ( .A(c8029), .B(n24087), .Z(c8030) );
ANDN U40146 ( .B(n24088), .A(n24089), .Z(n24087) );
XOR U40147 ( .A(c8029), .B(b[8029]), .Z(n24088) );
XNOR U40148 ( .A(b[8029]), .B(n24089), .Z(c[8029]) );
XNOR U40149 ( .A(a[8029]), .B(c8029), .Z(n24089) );
XOR U40150 ( .A(c8030), .B(n24090), .Z(c8031) );
ANDN U40151 ( .B(n24091), .A(n24092), .Z(n24090) );
XOR U40152 ( .A(c8030), .B(b[8030]), .Z(n24091) );
XNOR U40153 ( .A(b[8030]), .B(n24092), .Z(c[8030]) );
XNOR U40154 ( .A(a[8030]), .B(c8030), .Z(n24092) );
XOR U40155 ( .A(c8031), .B(n24093), .Z(c8032) );
ANDN U40156 ( .B(n24094), .A(n24095), .Z(n24093) );
XOR U40157 ( .A(c8031), .B(b[8031]), .Z(n24094) );
XNOR U40158 ( .A(b[8031]), .B(n24095), .Z(c[8031]) );
XNOR U40159 ( .A(a[8031]), .B(c8031), .Z(n24095) );
XOR U40160 ( .A(c8032), .B(n24096), .Z(c8033) );
ANDN U40161 ( .B(n24097), .A(n24098), .Z(n24096) );
XOR U40162 ( .A(c8032), .B(b[8032]), .Z(n24097) );
XNOR U40163 ( .A(b[8032]), .B(n24098), .Z(c[8032]) );
XNOR U40164 ( .A(a[8032]), .B(c8032), .Z(n24098) );
XOR U40165 ( .A(c8033), .B(n24099), .Z(c8034) );
ANDN U40166 ( .B(n24100), .A(n24101), .Z(n24099) );
XOR U40167 ( .A(c8033), .B(b[8033]), .Z(n24100) );
XNOR U40168 ( .A(b[8033]), .B(n24101), .Z(c[8033]) );
XNOR U40169 ( .A(a[8033]), .B(c8033), .Z(n24101) );
XOR U40170 ( .A(c8034), .B(n24102), .Z(c8035) );
ANDN U40171 ( .B(n24103), .A(n24104), .Z(n24102) );
XOR U40172 ( .A(c8034), .B(b[8034]), .Z(n24103) );
XNOR U40173 ( .A(b[8034]), .B(n24104), .Z(c[8034]) );
XNOR U40174 ( .A(a[8034]), .B(c8034), .Z(n24104) );
XOR U40175 ( .A(c8035), .B(n24105), .Z(c8036) );
ANDN U40176 ( .B(n24106), .A(n24107), .Z(n24105) );
XOR U40177 ( .A(c8035), .B(b[8035]), .Z(n24106) );
XNOR U40178 ( .A(b[8035]), .B(n24107), .Z(c[8035]) );
XNOR U40179 ( .A(a[8035]), .B(c8035), .Z(n24107) );
XOR U40180 ( .A(c8036), .B(n24108), .Z(c8037) );
ANDN U40181 ( .B(n24109), .A(n24110), .Z(n24108) );
XOR U40182 ( .A(c8036), .B(b[8036]), .Z(n24109) );
XNOR U40183 ( .A(b[8036]), .B(n24110), .Z(c[8036]) );
XNOR U40184 ( .A(a[8036]), .B(c8036), .Z(n24110) );
XOR U40185 ( .A(c8037), .B(n24111), .Z(c8038) );
ANDN U40186 ( .B(n24112), .A(n24113), .Z(n24111) );
XOR U40187 ( .A(c8037), .B(b[8037]), .Z(n24112) );
XNOR U40188 ( .A(b[8037]), .B(n24113), .Z(c[8037]) );
XNOR U40189 ( .A(a[8037]), .B(c8037), .Z(n24113) );
XOR U40190 ( .A(c8038), .B(n24114), .Z(c8039) );
ANDN U40191 ( .B(n24115), .A(n24116), .Z(n24114) );
XOR U40192 ( .A(c8038), .B(b[8038]), .Z(n24115) );
XNOR U40193 ( .A(b[8038]), .B(n24116), .Z(c[8038]) );
XNOR U40194 ( .A(a[8038]), .B(c8038), .Z(n24116) );
XOR U40195 ( .A(c8039), .B(n24117), .Z(c8040) );
ANDN U40196 ( .B(n24118), .A(n24119), .Z(n24117) );
XOR U40197 ( .A(c8039), .B(b[8039]), .Z(n24118) );
XNOR U40198 ( .A(b[8039]), .B(n24119), .Z(c[8039]) );
XNOR U40199 ( .A(a[8039]), .B(c8039), .Z(n24119) );
XOR U40200 ( .A(c8040), .B(n24120), .Z(c8041) );
ANDN U40201 ( .B(n24121), .A(n24122), .Z(n24120) );
XOR U40202 ( .A(c8040), .B(b[8040]), .Z(n24121) );
XNOR U40203 ( .A(b[8040]), .B(n24122), .Z(c[8040]) );
XNOR U40204 ( .A(a[8040]), .B(c8040), .Z(n24122) );
XOR U40205 ( .A(c8041), .B(n24123), .Z(c8042) );
ANDN U40206 ( .B(n24124), .A(n24125), .Z(n24123) );
XOR U40207 ( .A(c8041), .B(b[8041]), .Z(n24124) );
XNOR U40208 ( .A(b[8041]), .B(n24125), .Z(c[8041]) );
XNOR U40209 ( .A(a[8041]), .B(c8041), .Z(n24125) );
XOR U40210 ( .A(c8042), .B(n24126), .Z(c8043) );
ANDN U40211 ( .B(n24127), .A(n24128), .Z(n24126) );
XOR U40212 ( .A(c8042), .B(b[8042]), .Z(n24127) );
XNOR U40213 ( .A(b[8042]), .B(n24128), .Z(c[8042]) );
XNOR U40214 ( .A(a[8042]), .B(c8042), .Z(n24128) );
XOR U40215 ( .A(c8043), .B(n24129), .Z(c8044) );
ANDN U40216 ( .B(n24130), .A(n24131), .Z(n24129) );
XOR U40217 ( .A(c8043), .B(b[8043]), .Z(n24130) );
XNOR U40218 ( .A(b[8043]), .B(n24131), .Z(c[8043]) );
XNOR U40219 ( .A(a[8043]), .B(c8043), .Z(n24131) );
XOR U40220 ( .A(c8044), .B(n24132), .Z(c8045) );
ANDN U40221 ( .B(n24133), .A(n24134), .Z(n24132) );
XOR U40222 ( .A(c8044), .B(b[8044]), .Z(n24133) );
XNOR U40223 ( .A(b[8044]), .B(n24134), .Z(c[8044]) );
XNOR U40224 ( .A(a[8044]), .B(c8044), .Z(n24134) );
XOR U40225 ( .A(c8045), .B(n24135), .Z(c8046) );
ANDN U40226 ( .B(n24136), .A(n24137), .Z(n24135) );
XOR U40227 ( .A(c8045), .B(b[8045]), .Z(n24136) );
XNOR U40228 ( .A(b[8045]), .B(n24137), .Z(c[8045]) );
XNOR U40229 ( .A(a[8045]), .B(c8045), .Z(n24137) );
XOR U40230 ( .A(c8046), .B(n24138), .Z(c8047) );
ANDN U40231 ( .B(n24139), .A(n24140), .Z(n24138) );
XOR U40232 ( .A(c8046), .B(b[8046]), .Z(n24139) );
XNOR U40233 ( .A(b[8046]), .B(n24140), .Z(c[8046]) );
XNOR U40234 ( .A(a[8046]), .B(c8046), .Z(n24140) );
XOR U40235 ( .A(c8047), .B(n24141), .Z(c8048) );
ANDN U40236 ( .B(n24142), .A(n24143), .Z(n24141) );
XOR U40237 ( .A(c8047), .B(b[8047]), .Z(n24142) );
XNOR U40238 ( .A(b[8047]), .B(n24143), .Z(c[8047]) );
XNOR U40239 ( .A(a[8047]), .B(c8047), .Z(n24143) );
XOR U40240 ( .A(c8048), .B(n24144), .Z(c8049) );
ANDN U40241 ( .B(n24145), .A(n24146), .Z(n24144) );
XOR U40242 ( .A(c8048), .B(b[8048]), .Z(n24145) );
XNOR U40243 ( .A(b[8048]), .B(n24146), .Z(c[8048]) );
XNOR U40244 ( .A(a[8048]), .B(c8048), .Z(n24146) );
XOR U40245 ( .A(c8049), .B(n24147), .Z(c8050) );
ANDN U40246 ( .B(n24148), .A(n24149), .Z(n24147) );
XOR U40247 ( .A(c8049), .B(b[8049]), .Z(n24148) );
XNOR U40248 ( .A(b[8049]), .B(n24149), .Z(c[8049]) );
XNOR U40249 ( .A(a[8049]), .B(c8049), .Z(n24149) );
XOR U40250 ( .A(c8050), .B(n24150), .Z(c8051) );
ANDN U40251 ( .B(n24151), .A(n24152), .Z(n24150) );
XOR U40252 ( .A(c8050), .B(b[8050]), .Z(n24151) );
XNOR U40253 ( .A(b[8050]), .B(n24152), .Z(c[8050]) );
XNOR U40254 ( .A(a[8050]), .B(c8050), .Z(n24152) );
XOR U40255 ( .A(c8051), .B(n24153), .Z(c8052) );
ANDN U40256 ( .B(n24154), .A(n24155), .Z(n24153) );
XOR U40257 ( .A(c8051), .B(b[8051]), .Z(n24154) );
XNOR U40258 ( .A(b[8051]), .B(n24155), .Z(c[8051]) );
XNOR U40259 ( .A(a[8051]), .B(c8051), .Z(n24155) );
XOR U40260 ( .A(c8052), .B(n24156), .Z(c8053) );
ANDN U40261 ( .B(n24157), .A(n24158), .Z(n24156) );
XOR U40262 ( .A(c8052), .B(b[8052]), .Z(n24157) );
XNOR U40263 ( .A(b[8052]), .B(n24158), .Z(c[8052]) );
XNOR U40264 ( .A(a[8052]), .B(c8052), .Z(n24158) );
XOR U40265 ( .A(c8053), .B(n24159), .Z(c8054) );
ANDN U40266 ( .B(n24160), .A(n24161), .Z(n24159) );
XOR U40267 ( .A(c8053), .B(b[8053]), .Z(n24160) );
XNOR U40268 ( .A(b[8053]), .B(n24161), .Z(c[8053]) );
XNOR U40269 ( .A(a[8053]), .B(c8053), .Z(n24161) );
XOR U40270 ( .A(c8054), .B(n24162), .Z(c8055) );
ANDN U40271 ( .B(n24163), .A(n24164), .Z(n24162) );
XOR U40272 ( .A(c8054), .B(b[8054]), .Z(n24163) );
XNOR U40273 ( .A(b[8054]), .B(n24164), .Z(c[8054]) );
XNOR U40274 ( .A(a[8054]), .B(c8054), .Z(n24164) );
XOR U40275 ( .A(c8055), .B(n24165), .Z(c8056) );
ANDN U40276 ( .B(n24166), .A(n24167), .Z(n24165) );
XOR U40277 ( .A(c8055), .B(b[8055]), .Z(n24166) );
XNOR U40278 ( .A(b[8055]), .B(n24167), .Z(c[8055]) );
XNOR U40279 ( .A(a[8055]), .B(c8055), .Z(n24167) );
XOR U40280 ( .A(c8056), .B(n24168), .Z(c8057) );
ANDN U40281 ( .B(n24169), .A(n24170), .Z(n24168) );
XOR U40282 ( .A(c8056), .B(b[8056]), .Z(n24169) );
XNOR U40283 ( .A(b[8056]), .B(n24170), .Z(c[8056]) );
XNOR U40284 ( .A(a[8056]), .B(c8056), .Z(n24170) );
XOR U40285 ( .A(c8057), .B(n24171), .Z(c8058) );
ANDN U40286 ( .B(n24172), .A(n24173), .Z(n24171) );
XOR U40287 ( .A(c8057), .B(b[8057]), .Z(n24172) );
XNOR U40288 ( .A(b[8057]), .B(n24173), .Z(c[8057]) );
XNOR U40289 ( .A(a[8057]), .B(c8057), .Z(n24173) );
XOR U40290 ( .A(c8058), .B(n24174), .Z(c8059) );
ANDN U40291 ( .B(n24175), .A(n24176), .Z(n24174) );
XOR U40292 ( .A(c8058), .B(b[8058]), .Z(n24175) );
XNOR U40293 ( .A(b[8058]), .B(n24176), .Z(c[8058]) );
XNOR U40294 ( .A(a[8058]), .B(c8058), .Z(n24176) );
XOR U40295 ( .A(c8059), .B(n24177), .Z(c8060) );
ANDN U40296 ( .B(n24178), .A(n24179), .Z(n24177) );
XOR U40297 ( .A(c8059), .B(b[8059]), .Z(n24178) );
XNOR U40298 ( .A(b[8059]), .B(n24179), .Z(c[8059]) );
XNOR U40299 ( .A(a[8059]), .B(c8059), .Z(n24179) );
XOR U40300 ( .A(c8060), .B(n24180), .Z(c8061) );
ANDN U40301 ( .B(n24181), .A(n24182), .Z(n24180) );
XOR U40302 ( .A(c8060), .B(b[8060]), .Z(n24181) );
XNOR U40303 ( .A(b[8060]), .B(n24182), .Z(c[8060]) );
XNOR U40304 ( .A(a[8060]), .B(c8060), .Z(n24182) );
XOR U40305 ( .A(c8061), .B(n24183), .Z(c8062) );
ANDN U40306 ( .B(n24184), .A(n24185), .Z(n24183) );
XOR U40307 ( .A(c8061), .B(b[8061]), .Z(n24184) );
XNOR U40308 ( .A(b[8061]), .B(n24185), .Z(c[8061]) );
XNOR U40309 ( .A(a[8061]), .B(c8061), .Z(n24185) );
XOR U40310 ( .A(c8062), .B(n24186), .Z(c8063) );
ANDN U40311 ( .B(n24187), .A(n24188), .Z(n24186) );
XOR U40312 ( .A(c8062), .B(b[8062]), .Z(n24187) );
XNOR U40313 ( .A(b[8062]), .B(n24188), .Z(c[8062]) );
XNOR U40314 ( .A(a[8062]), .B(c8062), .Z(n24188) );
XOR U40315 ( .A(c8063), .B(n24189), .Z(c8064) );
ANDN U40316 ( .B(n24190), .A(n24191), .Z(n24189) );
XOR U40317 ( .A(c8063), .B(b[8063]), .Z(n24190) );
XNOR U40318 ( .A(b[8063]), .B(n24191), .Z(c[8063]) );
XNOR U40319 ( .A(a[8063]), .B(c8063), .Z(n24191) );
XOR U40320 ( .A(c8064), .B(n24192), .Z(c8065) );
ANDN U40321 ( .B(n24193), .A(n24194), .Z(n24192) );
XOR U40322 ( .A(c8064), .B(b[8064]), .Z(n24193) );
XNOR U40323 ( .A(b[8064]), .B(n24194), .Z(c[8064]) );
XNOR U40324 ( .A(a[8064]), .B(c8064), .Z(n24194) );
XOR U40325 ( .A(c8065), .B(n24195), .Z(c8066) );
ANDN U40326 ( .B(n24196), .A(n24197), .Z(n24195) );
XOR U40327 ( .A(c8065), .B(b[8065]), .Z(n24196) );
XNOR U40328 ( .A(b[8065]), .B(n24197), .Z(c[8065]) );
XNOR U40329 ( .A(a[8065]), .B(c8065), .Z(n24197) );
XOR U40330 ( .A(c8066), .B(n24198), .Z(c8067) );
ANDN U40331 ( .B(n24199), .A(n24200), .Z(n24198) );
XOR U40332 ( .A(c8066), .B(b[8066]), .Z(n24199) );
XNOR U40333 ( .A(b[8066]), .B(n24200), .Z(c[8066]) );
XNOR U40334 ( .A(a[8066]), .B(c8066), .Z(n24200) );
XOR U40335 ( .A(c8067), .B(n24201), .Z(c8068) );
ANDN U40336 ( .B(n24202), .A(n24203), .Z(n24201) );
XOR U40337 ( .A(c8067), .B(b[8067]), .Z(n24202) );
XNOR U40338 ( .A(b[8067]), .B(n24203), .Z(c[8067]) );
XNOR U40339 ( .A(a[8067]), .B(c8067), .Z(n24203) );
XOR U40340 ( .A(c8068), .B(n24204), .Z(c8069) );
ANDN U40341 ( .B(n24205), .A(n24206), .Z(n24204) );
XOR U40342 ( .A(c8068), .B(b[8068]), .Z(n24205) );
XNOR U40343 ( .A(b[8068]), .B(n24206), .Z(c[8068]) );
XNOR U40344 ( .A(a[8068]), .B(c8068), .Z(n24206) );
XOR U40345 ( .A(c8069), .B(n24207), .Z(c8070) );
ANDN U40346 ( .B(n24208), .A(n24209), .Z(n24207) );
XOR U40347 ( .A(c8069), .B(b[8069]), .Z(n24208) );
XNOR U40348 ( .A(b[8069]), .B(n24209), .Z(c[8069]) );
XNOR U40349 ( .A(a[8069]), .B(c8069), .Z(n24209) );
XOR U40350 ( .A(c8070), .B(n24210), .Z(c8071) );
ANDN U40351 ( .B(n24211), .A(n24212), .Z(n24210) );
XOR U40352 ( .A(c8070), .B(b[8070]), .Z(n24211) );
XNOR U40353 ( .A(b[8070]), .B(n24212), .Z(c[8070]) );
XNOR U40354 ( .A(a[8070]), .B(c8070), .Z(n24212) );
XOR U40355 ( .A(c8071), .B(n24213), .Z(c8072) );
ANDN U40356 ( .B(n24214), .A(n24215), .Z(n24213) );
XOR U40357 ( .A(c8071), .B(b[8071]), .Z(n24214) );
XNOR U40358 ( .A(b[8071]), .B(n24215), .Z(c[8071]) );
XNOR U40359 ( .A(a[8071]), .B(c8071), .Z(n24215) );
XOR U40360 ( .A(c8072), .B(n24216), .Z(c8073) );
ANDN U40361 ( .B(n24217), .A(n24218), .Z(n24216) );
XOR U40362 ( .A(c8072), .B(b[8072]), .Z(n24217) );
XNOR U40363 ( .A(b[8072]), .B(n24218), .Z(c[8072]) );
XNOR U40364 ( .A(a[8072]), .B(c8072), .Z(n24218) );
XOR U40365 ( .A(c8073), .B(n24219), .Z(c8074) );
ANDN U40366 ( .B(n24220), .A(n24221), .Z(n24219) );
XOR U40367 ( .A(c8073), .B(b[8073]), .Z(n24220) );
XNOR U40368 ( .A(b[8073]), .B(n24221), .Z(c[8073]) );
XNOR U40369 ( .A(a[8073]), .B(c8073), .Z(n24221) );
XOR U40370 ( .A(c8074), .B(n24222), .Z(c8075) );
ANDN U40371 ( .B(n24223), .A(n24224), .Z(n24222) );
XOR U40372 ( .A(c8074), .B(b[8074]), .Z(n24223) );
XNOR U40373 ( .A(b[8074]), .B(n24224), .Z(c[8074]) );
XNOR U40374 ( .A(a[8074]), .B(c8074), .Z(n24224) );
XOR U40375 ( .A(c8075), .B(n24225), .Z(c8076) );
ANDN U40376 ( .B(n24226), .A(n24227), .Z(n24225) );
XOR U40377 ( .A(c8075), .B(b[8075]), .Z(n24226) );
XNOR U40378 ( .A(b[8075]), .B(n24227), .Z(c[8075]) );
XNOR U40379 ( .A(a[8075]), .B(c8075), .Z(n24227) );
XOR U40380 ( .A(c8076), .B(n24228), .Z(c8077) );
ANDN U40381 ( .B(n24229), .A(n24230), .Z(n24228) );
XOR U40382 ( .A(c8076), .B(b[8076]), .Z(n24229) );
XNOR U40383 ( .A(b[8076]), .B(n24230), .Z(c[8076]) );
XNOR U40384 ( .A(a[8076]), .B(c8076), .Z(n24230) );
XOR U40385 ( .A(c8077), .B(n24231), .Z(c8078) );
ANDN U40386 ( .B(n24232), .A(n24233), .Z(n24231) );
XOR U40387 ( .A(c8077), .B(b[8077]), .Z(n24232) );
XNOR U40388 ( .A(b[8077]), .B(n24233), .Z(c[8077]) );
XNOR U40389 ( .A(a[8077]), .B(c8077), .Z(n24233) );
XOR U40390 ( .A(c8078), .B(n24234), .Z(c8079) );
ANDN U40391 ( .B(n24235), .A(n24236), .Z(n24234) );
XOR U40392 ( .A(c8078), .B(b[8078]), .Z(n24235) );
XNOR U40393 ( .A(b[8078]), .B(n24236), .Z(c[8078]) );
XNOR U40394 ( .A(a[8078]), .B(c8078), .Z(n24236) );
XOR U40395 ( .A(c8079), .B(n24237), .Z(c8080) );
ANDN U40396 ( .B(n24238), .A(n24239), .Z(n24237) );
XOR U40397 ( .A(c8079), .B(b[8079]), .Z(n24238) );
XNOR U40398 ( .A(b[8079]), .B(n24239), .Z(c[8079]) );
XNOR U40399 ( .A(a[8079]), .B(c8079), .Z(n24239) );
XOR U40400 ( .A(c8080), .B(n24240), .Z(c8081) );
ANDN U40401 ( .B(n24241), .A(n24242), .Z(n24240) );
XOR U40402 ( .A(c8080), .B(b[8080]), .Z(n24241) );
XNOR U40403 ( .A(b[8080]), .B(n24242), .Z(c[8080]) );
XNOR U40404 ( .A(a[8080]), .B(c8080), .Z(n24242) );
XOR U40405 ( .A(c8081), .B(n24243), .Z(c8082) );
ANDN U40406 ( .B(n24244), .A(n24245), .Z(n24243) );
XOR U40407 ( .A(c8081), .B(b[8081]), .Z(n24244) );
XNOR U40408 ( .A(b[8081]), .B(n24245), .Z(c[8081]) );
XNOR U40409 ( .A(a[8081]), .B(c8081), .Z(n24245) );
XOR U40410 ( .A(c8082), .B(n24246), .Z(c8083) );
ANDN U40411 ( .B(n24247), .A(n24248), .Z(n24246) );
XOR U40412 ( .A(c8082), .B(b[8082]), .Z(n24247) );
XNOR U40413 ( .A(b[8082]), .B(n24248), .Z(c[8082]) );
XNOR U40414 ( .A(a[8082]), .B(c8082), .Z(n24248) );
XOR U40415 ( .A(c8083), .B(n24249), .Z(c8084) );
ANDN U40416 ( .B(n24250), .A(n24251), .Z(n24249) );
XOR U40417 ( .A(c8083), .B(b[8083]), .Z(n24250) );
XNOR U40418 ( .A(b[8083]), .B(n24251), .Z(c[8083]) );
XNOR U40419 ( .A(a[8083]), .B(c8083), .Z(n24251) );
XOR U40420 ( .A(c8084), .B(n24252), .Z(c8085) );
ANDN U40421 ( .B(n24253), .A(n24254), .Z(n24252) );
XOR U40422 ( .A(c8084), .B(b[8084]), .Z(n24253) );
XNOR U40423 ( .A(b[8084]), .B(n24254), .Z(c[8084]) );
XNOR U40424 ( .A(a[8084]), .B(c8084), .Z(n24254) );
XOR U40425 ( .A(c8085), .B(n24255), .Z(c8086) );
ANDN U40426 ( .B(n24256), .A(n24257), .Z(n24255) );
XOR U40427 ( .A(c8085), .B(b[8085]), .Z(n24256) );
XNOR U40428 ( .A(b[8085]), .B(n24257), .Z(c[8085]) );
XNOR U40429 ( .A(a[8085]), .B(c8085), .Z(n24257) );
XOR U40430 ( .A(c8086), .B(n24258), .Z(c8087) );
ANDN U40431 ( .B(n24259), .A(n24260), .Z(n24258) );
XOR U40432 ( .A(c8086), .B(b[8086]), .Z(n24259) );
XNOR U40433 ( .A(b[8086]), .B(n24260), .Z(c[8086]) );
XNOR U40434 ( .A(a[8086]), .B(c8086), .Z(n24260) );
XOR U40435 ( .A(c8087), .B(n24261), .Z(c8088) );
ANDN U40436 ( .B(n24262), .A(n24263), .Z(n24261) );
XOR U40437 ( .A(c8087), .B(b[8087]), .Z(n24262) );
XNOR U40438 ( .A(b[8087]), .B(n24263), .Z(c[8087]) );
XNOR U40439 ( .A(a[8087]), .B(c8087), .Z(n24263) );
XOR U40440 ( .A(c8088), .B(n24264), .Z(c8089) );
ANDN U40441 ( .B(n24265), .A(n24266), .Z(n24264) );
XOR U40442 ( .A(c8088), .B(b[8088]), .Z(n24265) );
XNOR U40443 ( .A(b[8088]), .B(n24266), .Z(c[8088]) );
XNOR U40444 ( .A(a[8088]), .B(c8088), .Z(n24266) );
XOR U40445 ( .A(c8089), .B(n24267), .Z(c8090) );
ANDN U40446 ( .B(n24268), .A(n24269), .Z(n24267) );
XOR U40447 ( .A(c8089), .B(b[8089]), .Z(n24268) );
XNOR U40448 ( .A(b[8089]), .B(n24269), .Z(c[8089]) );
XNOR U40449 ( .A(a[8089]), .B(c8089), .Z(n24269) );
XOR U40450 ( .A(c8090), .B(n24270), .Z(c8091) );
ANDN U40451 ( .B(n24271), .A(n24272), .Z(n24270) );
XOR U40452 ( .A(c8090), .B(b[8090]), .Z(n24271) );
XNOR U40453 ( .A(b[8090]), .B(n24272), .Z(c[8090]) );
XNOR U40454 ( .A(a[8090]), .B(c8090), .Z(n24272) );
XOR U40455 ( .A(c8091), .B(n24273), .Z(c8092) );
ANDN U40456 ( .B(n24274), .A(n24275), .Z(n24273) );
XOR U40457 ( .A(c8091), .B(b[8091]), .Z(n24274) );
XNOR U40458 ( .A(b[8091]), .B(n24275), .Z(c[8091]) );
XNOR U40459 ( .A(a[8091]), .B(c8091), .Z(n24275) );
XOR U40460 ( .A(c8092), .B(n24276), .Z(c8093) );
ANDN U40461 ( .B(n24277), .A(n24278), .Z(n24276) );
XOR U40462 ( .A(c8092), .B(b[8092]), .Z(n24277) );
XNOR U40463 ( .A(b[8092]), .B(n24278), .Z(c[8092]) );
XNOR U40464 ( .A(a[8092]), .B(c8092), .Z(n24278) );
XOR U40465 ( .A(c8093), .B(n24279), .Z(c8094) );
ANDN U40466 ( .B(n24280), .A(n24281), .Z(n24279) );
XOR U40467 ( .A(c8093), .B(b[8093]), .Z(n24280) );
XNOR U40468 ( .A(b[8093]), .B(n24281), .Z(c[8093]) );
XNOR U40469 ( .A(a[8093]), .B(c8093), .Z(n24281) );
XOR U40470 ( .A(c8094), .B(n24282), .Z(c8095) );
ANDN U40471 ( .B(n24283), .A(n24284), .Z(n24282) );
XOR U40472 ( .A(c8094), .B(b[8094]), .Z(n24283) );
XNOR U40473 ( .A(b[8094]), .B(n24284), .Z(c[8094]) );
XNOR U40474 ( .A(a[8094]), .B(c8094), .Z(n24284) );
XOR U40475 ( .A(c8095), .B(n24285), .Z(c8096) );
ANDN U40476 ( .B(n24286), .A(n24287), .Z(n24285) );
XOR U40477 ( .A(c8095), .B(b[8095]), .Z(n24286) );
XNOR U40478 ( .A(b[8095]), .B(n24287), .Z(c[8095]) );
XNOR U40479 ( .A(a[8095]), .B(c8095), .Z(n24287) );
XOR U40480 ( .A(c8096), .B(n24288), .Z(c8097) );
ANDN U40481 ( .B(n24289), .A(n24290), .Z(n24288) );
XOR U40482 ( .A(c8096), .B(b[8096]), .Z(n24289) );
XNOR U40483 ( .A(b[8096]), .B(n24290), .Z(c[8096]) );
XNOR U40484 ( .A(a[8096]), .B(c8096), .Z(n24290) );
XOR U40485 ( .A(c8097), .B(n24291), .Z(c8098) );
ANDN U40486 ( .B(n24292), .A(n24293), .Z(n24291) );
XOR U40487 ( .A(c8097), .B(b[8097]), .Z(n24292) );
XNOR U40488 ( .A(b[8097]), .B(n24293), .Z(c[8097]) );
XNOR U40489 ( .A(a[8097]), .B(c8097), .Z(n24293) );
XOR U40490 ( .A(c8098), .B(n24294), .Z(c8099) );
ANDN U40491 ( .B(n24295), .A(n24296), .Z(n24294) );
XOR U40492 ( .A(c8098), .B(b[8098]), .Z(n24295) );
XNOR U40493 ( .A(b[8098]), .B(n24296), .Z(c[8098]) );
XNOR U40494 ( .A(a[8098]), .B(c8098), .Z(n24296) );
XOR U40495 ( .A(c8099), .B(n24297), .Z(c8100) );
ANDN U40496 ( .B(n24298), .A(n24299), .Z(n24297) );
XOR U40497 ( .A(c8099), .B(b[8099]), .Z(n24298) );
XNOR U40498 ( .A(b[8099]), .B(n24299), .Z(c[8099]) );
XNOR U40499 ( .A(a[8099]), .B(c8099), .Z(n24299) );
XOR U40500 ( .A(c8100), .B(n24300), .Z(c8101) );
ANDN U40501 ( .B(n24301), .A(n24302), .Z(n24300) );
XOR U40502 ( .A(c8100), .B(b[8100]), .Z(n24301) );
XNOR U40503 ( .A(b[8100]), .B(n24302), .Z(c[8100]) );
XNOR U40504 ( .A(a[8100]), .B(c8100), .Z(n24302) );
XOR U40505 ( .A(c8101), .B(n24303), .Z(c8102) );
ANDN U40506 ( .B(n24304), .A(n24305), .Z(n24303) );
XOR U40507 ( .A(c8101), .B(b[8101]), .Z(n24304) );
XNOR U40508 ( .A(b[8101]), .B(n24305), .Z(c[8101]) );
XNOR U40509 ( .A(a[8101]), .B(c8101), .Z(n24305) );
XOR U40510 ( .A(c8102), .B(n24306), .Z(c8103) );
ANDN U40511 ( .B(n24307), .A(n24308), .Z(n24306) );
XOR U40512 ( .A(c8102), .B(b[8102]), .Z(n24307) );
XNOR U40513 ( .A(b[8102]), .B(n24308), .Z(c[8102]) );
XNOR U40514 ( .A(a[8102]), .B(c8102), .Z(n24308) );
XOR U40515 ( .A(c8103), .B(n24309), .Z(c8104) );
ANDN U40516 ( .B(n24310), .A(n24311), .Z(n24309) );
XOR U40517 ( .A(c8103), .B(b[8103]), .Z(n24310) );
XNOR U40518 ( .A(b[8103]), .B(n24311), .Z(c[8103]) );
XNOR U40519 ( .A(a[8103]), .B(c8103), .Z(n24311) );
XOR U40520 ( .A(c8104), .B(n24312), .Z(c8105) );
ANDN U40521 ( .B(n24313), .A(n24314), .Z(n24312) );
XOR U40522 ( .A(c8104), .B(b[8104]), .Z(n24313) );
XNOR U40523 ( .A(b[8104]), .B(n24314), .Z(c[8104]) );
XNOR U40524 ( .A(a[8104]), .B(c8104), .Z(n24314) );
XOR U40525 ( .A(c8105), .B(n24315), .Z(c8106) );
ANDN U40526 ( .B(n24316), .A(n24317), .Z(n24315) );
XOR U40527 ( .A(c8105), .B(b[8105]), .Z(n24316) );
XNOR U40528 ( .A(b[8105]), .B(n24317), .Z(c[8105]) );
XNOR U40529 ( .A(a[8105]), .B(c8105), .Z(n24317) );
XOR U40530 ( .A(c8106), .B(n24318), .Z(c8107) );
ANDN U40531 ( .B(n24319), .A(n24320), .Z(n24318) );
XOR U40532 ( .A(c8106), .B(b[8106]), .Z(n24319) );
XNOR U40533 ( .A(b[8106]), .B(n24320), .Z(c[8106]) );
XNOR U40534 ( .A(a[8106]), .B(c8106), .Z(n24320) );
XOR U40535 ( .A(c8107), .B(n24321), .Z(c8108) );
ANDN U40536 ( .B(n24322), .A(n24323), .Z(n24321) );
XOR U40537 ( .A(c8107), .B(b[8107]), .Z(n24322) );
XNOR U40538 ( .A(b[8107]), .B(n24323), .Z(c[8107]) );
XNOR U40539 ( .A(a[8107]), .B(c8107), .Z(n24323) );
XOR U40540 ( .A(c8108), .B(n24324), .Z(c8109) );
ANDN U40541 ( .B(n24325), .A(n24326), .Z(n24324) );
XOR U40542 ( .A(c8108), .B(b[8108]), .Z(n24325) );
XNOR U40543 ( .A(b[8108]), .B(n24326), .Z(c[8108]) );
XNOR U40544 ( .A(a[8108]), .B(c8108), .Z(n24326) );
XOR U40545 ( .A(c8109), .B(n24327), .Z(c8110) );
ANDN U40546 ( .B(n24328), .A(n24329), .Z(n24327) );
XOR U40547 ( .A(c8109), .B(b[8109]), .Z(n24328) );
XNOR U40548 ( .A(b[8109]), .B(n24329), .Z(c[8109]) );
XNOR U40549 ( .A(a[8109]), .B(c8109), .Z(n24329) );
XOR U40550 ( .A(c8110), .B(n24330), .Z(c8111) );
ANDN U40551 ( .B(n24331), .A(n24332), .Z(n24330) );
XOR U40552 ( .A(c8110), .B(b[8110]), .Z(n24331) );
XNOR U40553 ( .A(b[8110]), .B(n24332), .Z(c[8110]) );
XNOR U40554 ( .A(a[8110]), .B(c8110), .Z(n24332) );
XOR U40555 ( .A(c8111), .B(n24333), .Z(c8112) );
ANDN U40556 ( .B(n24334), .A(n24335), .Z(n24333) );
XOR U40557 ( .A(c8111), .B(b[8111]), .Z(n24334) );
XNOR U40558 ( .A(b[8111]), .B(n24335), .Z(c[8111]) );
XNOR U40559 ( .A(a[8111]), .B(c8111), .Z(n24335) );
XOR U40560 ( .A(c8112), .B(n24336), .Z(c8113) );
ANDN U40561 ( .B(n24337), .A(n24338), .Z(n24336) );
XOR U40562 ( .A(c8112), .B(b[8112]), .Z(n24337) );
XNOR U40563 ( .A(b[8112]), .B(n24338), .Z(c[8112]) );
XNOR U40564 ( .A(a[8112]), .B(c8112), .Z(n24338) );
XOR U40565 ( .A(c8113), .B(n24339), .Z(c8114) );
ANDN U40566 ( .B(n24340), .A(n24341), .Z(n24339) );
XOR U40567 ( .A(c8113), .B(b[8113]), .Z(n24340) );
XNOR U40568 ( .A(b[8113]), .B(n24341), .Z(c[8113]) );
XNOR U40569 ( .A(a[8113]), .B(c8113), .Z(n24341) );
XOR U40570 ( .A(c8114), .B(n24342), .Z(c8115) );
ANDN U40571 ( .B(n24343), .A(n24344), .Z(n24342) );
XOR U40572 ( .A(c8114), .B(b[8114]), .Z(n24343) );
XNOR U40573 ( .A(b[8114]), .B(n24344), .Z(c[8114]) );
XNOR U40574 ( .A(a[8114]), .B(c8114), .Z(n24344) );
XOR U40575 ( .A(c8115), .B(n24345), .Z(c8116) );
ANDN U40576 ( .B(n24346), .A(n24347), .Z(n24345) );
XOR U40577 ( .A(c8115), .B(b[8115]), .Z(n24346) );
XNOR U40578 ( .A(b[8115]), .B(n24347), .Z(c[8115]) );
XNOR U40579 ( .A(a[8115]), .B(c8115), .Z(n24347) );
XOR U40580 ( .A(c8116), .B(n24348), .Z(c8117) );
ANDN U40581 ( .B(n24349), .A(n24350), .Z(n24348) );
XOR U40582 ( .A(c8116), .B(b[8116]), .Z(n24349) );
XNOR U40583 ( .A(b[8116]), .B(n24350), .Z(c[8116]) );
XNOR U40584 ( .A(a[8116]), .B(c8116), .Z(n24350) );
XOR U40585 ( .A(c8117), .B(n24351), .Z(c8118) );
ANDN U40586 ( .B(n24352), .A(n24353), .Z(n24351) );
XOR U40587 ( .A(c8117), .B(b[8117]), .Z(n24352) );
XNOR U40588 ( .A(b[8117]), .B(n24353), .Z(c[8117]) );
XNOR U40589 ( .A(a[8117]), .B(c8117), .Z(n24353) );
XOR U40590 ( .A(c8118), .B(n24354), .Z(c8119) );
ANDN U40591 ( .B(n24355), .A(n24356), .Z(n24354) );
XOR U40592 ( .A(c8118), .B(b[8118]), .Z(n24355) );
XNOR U40593 ( .A(b[8118]), .B(n24356), .Z(c[8118]) );
XNOR U40594 ( .A(a[8118]), .B(c8118), .Z(n24356) );
XOR U40595 ( .A(c8119), .B(n24357), .Z(c8120) );
ANDN U40596 ( .B(n24358), .A(n24359), .Z(n24357) );
XOR U40597 ( .A(c8119), .B(b[8119]), .Z(n24358) );
XNOR U40598 ( .A(b[8119]), .B(n24359), .Z(c[8119]) );
XNOR U40599 ( .A(a[8119]), .B(c8119), .Z(n24359) );
XOR U40600 ( .A(c8120), .B(n24360), .Z(c8121) );
ANDN U40601 ( .B(n24361), .A(n24362), .Z(n24360) );
XOR U40602 ( .A(c8120), .B(b[8120]), .Z(n24361) );
XNOR U40603 ( .A(b[8120]), .B(n24362), .Z(c[8120]) );
XNOR U40604 ( .A(a[8120]), .B(c8120), .Z(n24362) );
XOR U40605 ( .A(c8121), .B(n24363), .Z(c8122) );
ANDN U40606 ( .B(n24364), .A(n24365), .Z(n24363) );
XOR U40607 ( .A(c8121), .B(b[8121]), .Z(n24364) );
XNOR U40608 ( .A(b[8121]), .B(n24365), .Z(c[8121]) );
XNOR U40609 ( .A(a[8121]), .B(c8121), .Z(n24365) );
XOR U40610 ( .A(c8122), .B(n24366), .Z(c8123) );
ANDN U40611 ( .B(n24367), .A(n24368), .Z(n24366) );
XOR U40612 ( .A(c8122), .B(b[8122]), .Z(n24367) );
XNOR U40613 ( .A(b[8122]), .B(n24368), .Z(c[8122]) );
XNOR U40614 ( .A(a[8122]), .B(c8122), .Z(n24368) );
XOR U40615 ( .A(c8123), .B(n24369), .Z(c8124) );
ANDN U40616 ( .B(n24370), .A(n24371), .Z(n24369) );
XOR U40617 ( .A(c8123), .B(b[8123]), .Z(n24370) );
XNOR U40618 ( .A(b[8123]), .B(n24371), .Z(c[8123]) );
XNOR U40619 ( .A(a[8123]), .B(c8123), .Z(n24371) );
XOR U40620 ( .A(c8124), .B(n24372), .Z(c8125) );
ANDN U40621 ( .B(n24373), .A(n24374), .Z(n24372) );
XOR U40622 ( .A(c8124), .B(b[8124]), .Z(n24373) );
XNOR U40623 ( .A(b[8124]), .B(n24374), .Z(c[8124]) );
XNOR U40624 ( .A(a[8124]), .B(c8124), .Z(n24374) );
XOR U40625 ( .A(c8125), .B(n24375), .Z(c8126) );
ANDN U40626 ( .B(n24376), .A(n24377), .Z(n24375) );
XOR U40627 ( .A(c8125), .B(b[8125]), .Z(n24376) );
XNOR U40628 ( .A(b[8125]), .B(n24377), .Z(c[8125]) );
XNOR U40629 ( .A(a[8125]), .B(c8125), .Z(n24377) );
XOR U40630 ( .A(c8126), .B(n24378), .Z(c8127) );
ANDN U40631 ( .B(n24379), .A(n24380), .Z(n24378) );
XOR U40632 ( .A(c8126), .B(b[8126]), .Z(n24379) );
XNOR U40633 ( .A(b[8126]), .B(n24380), .Z(c[8126]) );
XNOR U40634 ( .A(a[8126]), .B(c8126), .Z(n24380) );
XOR U40635 ( .A(c8127), .B(n24381), .Z(c8128) );
ANDN U40636 ( .B(n24382), .A(n24383), .Z(n24381) );
XOR U40637 ( .A(c8127), .B(b[8127]), .Z(n24382) );
XNOR U40638 ( .A(b[8127]), .B(n24383), .Z(c[8127]) );
XNOR U40639 ( .A(a[8127]), .B(c8127), .Z(n24383) );
XOR U40640 ( .A(c8128), .B(n24384), .Z(c8129) );
ANDN U40641 ( .B(n24385), .A(n24386), .Z(n24384) );
XOR U40642 ( .A(c8128), .B(b[8128]), .Z(n24385) );
XNOR U40643 ( .A(b[8128]), .B(n24386), .Z(c[8128]) );
XNOR U40644 ( .A(a[8128]), .B(c8128), .Z(n24386) );
XOR U40645 ( .A(c8129), .B(n24387), .Z(c8130) );
ANDN U40646 ( .B(n24388), .A(n24389), .Z(n24387) );
XOR U40647 ( .A(c8129), .B(b[8129]), .Z(n24388) );
XNOR U40648 ( .A(b[8129]), .B(n24389), .Z(c[8129]) );
XNOR U40649 ( .A(a[8129]), .B(c8129), .Z(n24389) );
XOR U40650 ( .A(c8130), .B(n24390), .Z(c8131) );
ANDN U40651 ( .B(n24391), .A(n24392), .Z(n24390) );
XOR U40652 ( .A(c8130), .B(b[8130]), .Z(n24391) );
XNOR U40653 ( .A(b[8130]), .B(n24392), .Z(c[8130]) );
XNOR U40654 ( .A(a[8130]), .B(c8130), .Z(n24392) );
XOR U40655 ( .A(c8131), .B(n24393), .Z(c8132) );
ANDN U40656 ( .B(n24394), .A(n24395), .Z(n24393) );
XOR U40657 ( .A(c8131), .B(b[8131]), .Z(n24394) );
XNOR U40658 ( .A(b[8131]), .B(n24395), .Z(c[8131]) );
XNOR U40659 ( .A(a[8131]), .B(c8131), .Z(n24395) );
XOR U40660 ( .A(c8132), .B(n24396), .Z(c8133) );
ANDN U40661 ( .B(n24397), .A(n24398), .Z(n24396) );
XOR U40662 ( .A(c8132), .B(b[8132]), .Z(n24397) );
XNOR U40663 ( .A(b[8132]), .B(n24398), .Z(c[8132]) );
XNOR U40664 ( .A(a[8132]), .B(c8132), .Z(n24398) );
XOR U40665 ( .A(c8133), .B(n24399), .Z(c8134) );
ANDN U40666 ( .B(n24400), .A(n24401), .Z(n24399) );
XOR U40667 ( .A(c8133), .B(b[8133]), .Z(n24400) );
XNOR U40668 ( .A(b[8133]), .B(n24401), .Z(c[8133]) );
XNOR U40669 ( .A(a[8133]), .B(c8133), .Z(n24401) );
XOR U40670 ( .A(c8134), .B(n24402), .Z(c8135) );
ANDN U40671 ( .B(n24403), .A(n24404), .Z(n24402) );
XOR U40672 ( .A(c8134), .B(b[8134]), .Z(n24403) );
XNOR U40673 ( .A(b[8134]), .B(n24404), .Z(c[8134]) );
XNOR U40674 ( .A(a[8134]), .B(c8134), .Z(n24404) );
XOR U40675 ( .A(c8135), .B(n24405), .Z(c8136) );
ANDN U40676 ( .B(n24406), .A(n24407), .Z(n24405) );
XOR U40677 ( .A(c8135), .B(b[8135]), .Z(n24406) );
XNOR U40678 ( .A(b[8135]), .B(n24407), .Z(c[8135]) );
XNOR U40679 ( .A(a[8135]), .B(c8135), .Z(n24407) );
XOR U40680 ( .A(c8136), .B(n24408), .Z(c8137) );
ANDN U40681 ( .B(n24409), .A(n24410), .Z(n24408) );
XOR U40682 ( .A(c8136), .B(b[8136]), .Z(n24409) );
XNOR U40683 ( .A(b[8136]), .B(n24410), .Z(c[8136]) );
XNOR U40684 ( .A(a[8136]), .B(c8136), .Z(n24410) );
XOR U40685 ( .A(c8137), .B(n24411), .Z(c8138) );
ANDN U40686 ( .B(n24412), .A(n24413), .Z(n24411) );
XOR U40687 ( .A(c8137), .B(b[8137]), .Z(n24412) );
XNOR U40688 ( .A(b[8137]), .B(n24413), .Z(c[8137]) );
XNOR U40689 ( .A(a[8137]), .B(c8137), .Z(n24413) );
XOR U40690 ( .A(c8138), .B(n24414), .Z(c8139) );
ANDN U40691 ( .B(n24415), .A(n24416), .Z(n24414) );
XOR U40692 ( .A(c8138), .B(b[8138]), .Z(n24415) );
XNOR U40693 ( .A(b[8138]), .B(n24416), .Z(c[8138]) );
XNOR U40694 ( .A(a[8138]), .B(c8138), .Z(n24416) );
XOR U40695 ( .A(c8139), .B(n24417), .Z(c8140) );
ANDN U40696 ( .B(n24418), .A(n24419), .Z(n24417) );
XOR U40697 ( .A(c8139), .B(b[8139]), .Z(n24418) );
XNOR U40698 ( .A(b[8139]), .B(n24419), .Z(c[8139]) );
XNOR U40699 ( .A(a[8139]), .B(c8139), .Z(n24419) );
XOR U40700 ( .A(c8140), .B(n24420), .Z(c8141) );
ANDN U40701 ( .B(n24421), .A(n24422), .Z(n24420) );
XOR U40702 ( .A(c8140), .B(b[8140]), .Z(n24421) );
XNOR U40703 ( .A(b[8140]), .B(n24422), .Z(c[8140]) );
XNOR U40704 ( .A(a[8140]), .B(c8140), .Z(n24422) );
XOR U40705 ( .A(c8141), .B(n24423), .Z(c8142) );
ANDN U40706 ( .B(n24424), .A(n24425), .Z(n24423) );
XOR U40707 ( .A(c8141), .B(b[8141]), .Z(n24424) );
XNOR U40708 ( .A(b[8141]), .B(n24425), .Z(c[8141]) );
XNOR U40709 ( .A(a[8141]), .B(c8141), .Z(n24425) );
XOR U40710 ( .A(c8142), .B(n24426), .Z(c8143) );
ANDN U40711 ( .B(n24427), .A(n24428), .Z(n24426) );
XOR U40712 ( .A(c8142), .B(b[8142]), .Z(n24427) );
XNOR U40713 ( .A(b[8142]), .B(n24428), .Z(c[8142]) );
XNOR U40714 ( .A(a[8142]), .B(c8142), .Z(n24428) );
XOR U40715 ( .A(c8143), .B(n24429), .Z(c8144) );
ANDN U40716 ( .B(n24430), .A(n24431), .Z(n24429) );
XOR U40717 ( .A(c8143), .B(b[8143]), .Z(n24430) );
XNOR U40718 ( .A(b[8143]), .B(n24431), .Z(c[8143]) );
XNOR U40719 ( .A(a[8143]), .B(c8143), .Z(n24431) );
XOR U40720 ( .A(c8144), .B(n24432), .Z(c8145) );
ANDN U40721 ( .B(n24433), .A(n24434), .Z(n24432) );
XOR U40722 ( .A(c8144), .B(b[8144]), .Z(n24433) );
XNOR U40723 ( .A(b[8144]), .B(n24434), .Z(c[8144]) );
XNOR U40724 ( .A(a[8144]), .B(c8144), .Z(n24434) );
XOR U40725 ( .A(c8145), .B(n24435), .Z(c8146) );
ANDN U40726 ( .B(n24436), .A(n24437), .Z(n24435) );
XOR U40727 ( .A(c8145), .B(b[8145]), .Z(n24436) );
XNOR U40728 ( .A(b[8145]), .B(n24437), .Z(c[8145]) );
XNOR U40729 ( .A(a[8145]), .B(c8145), .Z(n24437) );
XOR U40730 ( .A(c8146), .B(n24438), .Z(c8147) );
ANDN U40731 ( .B(n24439), .A(n24440), .Z(n24438) );
XOR U40732 ( .A(c8146), .B(b[8146]), .Z(n24439) );
XNOR U40733 ( .A(b[8146]), .B(n24440), .Z(c[8146]) );
XNOR U40734 ( .A(a[8146]), .B(c8146), .Z(n24440) );
XOR U40735 ( .A(c8147), .B(n24441), .Z(c8148) );
ANDN U40736 ( .B(n24442), .A(n24443), .Z(n24441) );
XOR U40737 ( .A(c8147), .B(b[8147]), .Z(n24442) );
XNOR U40738 ( .A(b[8147]), .B(n24443), .Z(c[8147]) );
XNOR U40739 ( .A(a[8147]), .B(c8147), .Z(n24443) );
XOR U40740 ( .A(c8148), .B(n24444), .Z(c8149) );
ANDN U40741 ( .B(n24445), .A(n24446), .Z(n24444) );
XOR U40742 ( .A(c8148), .B(b[8148]), .Z(n24445) );
XNOR U40743 ( .A(b[8148]), .B(n24446), .Z(c[8148]) );
XNOR U40744 ( .A(a[8148]), .B(c8148), .Z(n24446) );
XOR U40745 ( .A(c8149), .B(n24447), .Z(c8150) );
ANDN U40746 ( .B(n24448), .A(n24449), .Z(n24447) );
XOR U40747 ( .A(c8149), .B(b[8149]), .Z(n24448) );
XNOR U40748 ( .A(b[8149]), .B(n24449), .Z(c[8149]) );
XNOR U40749 ( .A(a[8149]), .B(c8149), .Z(n24449) );
XOR U40750 ( .A(c8150), .B(n24450), .Z(c8151) );
ANDN U40751 ( .B(n24451), .A(n24452), .Z(n24450) );
XOR U40752 ( .A(c8150), .B(b[8150]), .Z(n24451) );
XNOR U40753 ( .A(b[8150]), .B(n24452), .Z(c[8150]) );
XNOR U40754 ( .A(a[8150]), .B(c8150), .Z(n24452) );
XOR U40755 ( .A(c8151), .B(n24453), .Z(c8152) );
ANDN U40756 ( .B(n24454), .A(n24455), .Z(n24453) );
XOR U40757 ( .A(c8151), .B(b[8151]), .Z(n24454) );
XNOR U40758 ( .A(b[8151]), .B(n24455), .Z(c[8151]) );
XNOR U40759 ( .A(a[8151]), .B(c8151), .Z(n24455) );
XOR U40760 ( .A(c8152), .B(n24456), .Z(c8153) );
ANDN U40761 ( .B(n24457), .A(n24458), .Z(n24456) );
XOR U40762 ( .A(c8152), .B(b[8152]), .Z(n24457) );
XNOR U40763 ( .A(b[8152]), .B(n24458), .Z(c[8152]) );
XNOR U40764 ( .A(a[8152]), .B(c8152), .Z(n24458) );
XOR U40765 ( .A(c8153), .B(n24459), .Z(c8154) );
ANDN U40766 ( .B(n24460), .A(n24461), .Z(n24459) );
XOR U40767 ( .A(c8153), .B(b[8153]), .Z(n24460) );
XNOR U40768 ( .A(b[8153]), .B(n24461), .Z(c[8153]) );
XNOR U40769 ( .A(a[8153]), .B(c8153), .Z(n24461) );
XOR U40770 ( .A(c8154), .B(n24462), .Z(c8155) );
ANDN U40771 ( .B(n24463), .A(n24464), .Z(n24462) );
XOR U40772 ( .A(c8154), .B(b[8154]), .Z(n24463) );
XNOR U40773 ( .A(b[8154]), .B(n24464), .Z(c[8154]) );
XNOR U40774 ( .A(a[8154]), .B(c8154), .Z(n24464) );
XOR U40775 ( .A(c8155), .B(n24465), .Z(c8156) );
ANDN U40776 ( .B(n24466), .A(n24467), .Z(n24465) );
XOR U40777 ( .A(c8155), .B(b[8155]), .Z(n24466) );
XNOR U40778 ( .A(b[8155]), .B(n24467), .Z(c[8155]) );
XNOR U40779 ( .A(a[8155]), .B(c8155), .Z(n24467) );
XOR U40780 ( .A(c8156), .B(n24468), .Z(c8157) );
ANDN U40781 ( .B(n24469), .A(n24470), .Z(n24468) );
XOR U40782 ( .A(c8156), .B(b[8156]), .Z(n24469) );
XNOR U40783 ( .A(b[8156]), .B(n24470), .Z(c[8156]) );
XNOR U40784 ( .A(a[8156]), .B(c8156), .Z(n24470) );
XOR U40785 ( .A(c8157), .B(n24471), .Z(c8158) );
ANDN U40786 ( .B(n24472), .A(n24473), .Z(n24471) );
XOR U40787 ( .A(c8157), .B(b[8157]), .Z(n24472) );
XNOR U40788 ( .A(b[8157]), .B(n24473), .Z(c[8157]) );
XNOR U40789 ( .A(a[8157]), .B(c8157), .Z(n24473) );
XOR U40790 ( .A(c8158), .B(n24474), .Z(c8159) );
ANDN U40791 ( .B(n24475), .A(n24476), .Z(n24474) );
XOR U40792 ( .A(c8158), .B(b[8158]), .Z(n24475) );
XNOR U40793 ( .A(b[8158]), .B(n24476), .Z(c[8158]) );
XNOR U40794 ( .A(a[8158]), .B(c8158), .Z(n24476) );
XOR U40795 ( .A(c8159), .B(n24477), .Z(c8160) );
ANDN U40796 ( .B(n24478), .A(n24479), .Z(n24477) );
XOR U40797 ( .A(c8159), .B(b[8159]), .Z(n24478) );
XNOR U40798 ( .A(b[8159]), .B(n24479), .Z(c[8159]) );
XNOR U40799 ( .A(a[8159]), .B(c8159), .Z(n24479) );
XOR U40800 ( .A(c8160), .B(n24480), .Z(c8161) );
ANDN U40801 ( .B(n24481), .A(n24482), .Z(n24480) );
XOR U40802 ( .A(c8160), .B(b[8160]), .Z(n24481) );
XNOR U40803 ( .A(b[8160]), .B(n24482), .Z(c[8160]) );
XNOR U40804 ( .A(a[8160]), .B(c8160), .Z(n24482) );
XOR U40805 ( .A(c8161), .B(n24483), .Z(c8162) );
ANDN U40806 ( .B(n24484), .A(n24485), .Z(n24483) );
XOR U40807 ( .A(c8161), .B(b[8161]), .Z(n24484) );
XNOR U40808 ( .A(b[8161]), .B(n24485), .Z(c[8161]) );
XNOR U40809 ( .A(a[8161]), .B(c8161), .Z(n24485) );
XOR U40810 ( .A(c8162), .B(n24486), .Z(c8163) );
ANDN U40811 ( .B(n24487), .A(n24488), .Z(n24486) );
XOR U40812 ( .A(c8162), .B(b[8162]), .Z(n24487) );
XNOR U40813 ( .A(b[8162]), .B(n24488), .Z(c[8162]) );
XNOR U40814 ( .A(a[8162]), .B(c8162), .Z(n24488) );
XOR U40815 ( .A(c8163), .B(n24489), .Z(c8164) );
ANDN U40816 ( .B(n24490), .A(n24491), .Z(n24489) );
XOR U40817 ( .A(c8163), .B(b[8163]), .Z(n24490) );
XNOR U40818 ( .A(b[8163]), .B(n24491), .Z(c[8163]) );
XNOR U40819 ( .A(a[8163]), .B(c8163), .Z(n24491) );
XOR U40820 ( .A(c8164), .B(n24492), .Z(c8165) );
ANDN U40821 ( .B(n24493), .A(n24494), .Z(n24492) );
XOR U40822 ( .A(c8164), .B(b[8164]), .Z(n24493) );
XNOR U40823 ( .A(b[8164]), .B(n24494), .Z(c[8164]) );
XNOR U40824 ( .A(a[8164]), .B(c8164), .Z(n24494) );
XOR U40825 ( .A(c8165), .B(n24495), .Z(c8166) );
ANDN U40826 ( .B(n24496), .A(n24497), .Z(n24495) );
XOR U40827 ( .A(c8165), .B(b[8165]), .Z(n24496) );
XNOR U40828 ( .A(b[8165]), .B(n24497), .Z(c[8165]) );
XNOR U40829 ( .A(a[8165]), .B(c8165), .Z(n24497) );
XOR U40830 ( .A(c8166), .B(n24498), .Z(c8167) );
ANDN U40831 ( .B(n24499), .A(n24500), .Z(n24498) );
XOR U40832 ( .A(c8166), .B(b[8166]), .Z(n24499) );
XNOR U40833 ( .A(b[8166]), .B(n24500), .Z(c[8166]) );
XNOR U40834 ( .A(a[8166]), .B(c8166), .Z(n24500) );
XOR U40835 ( .A(c8167), .B(n24501), .Z(c8168) );
ANDN U40836 ( .B(n24502), .A(n24503), .Z(n24501) );
XOR U40837 ( .A(c8167), .B(b[8167]), .Z(n24502) );
XNOR U40838 ( .A(b[8167]), .B(n24503), .Z(c[8167]) );
XNOR U40839 ( .A(a[8167]), .B(c8167), .Z(n24503) );
XOR U40840 ( .A(c8168), .B(n24504), .Z(c8169) );
ANDN U40841 ( .B(n24505), .A(n24506), .Z(n24504) );
XOR U40842 ( .A(c8168), .B(b[8168]), .Z(n24505) );
XNOR U40843 ( .A(b[8168]), .B(n24506), .Z(c[8168]) );
XNOR U40844 ( .A(a[8168]), .B(c8168), .Z(n24506) );
XOR U40845 ( .A(c8169), .B(n24507), .Z(c8170) );
ANDN U40846 ( .B(n24508), .A(n24509), .Z(n24507) );
XOR U40847 ( .A(c8169), .B(b[8169]), .Z(n24508) );
XNOR U40848 ( .A(b[8169]), .B(n24509), .Z(c[8169]) );
XNOR U40849 ( .A(a[8169]), .B(c8169), .Z(n24509) );
XOR U40850 ( .A(c8170), .B(n24510), .Z(c8171) );
ANDN U40851 ( .B(n24511), .A(n24512), .Z(n24510) );
XOR U40852 ( .A(c8170), .B(b[8170]), .Z(n24511) );
XNOR U40853 ( .A(b[8170]), .B(n24512), .Z(c[8170]) );
XNOR U40854 ( .A(a[8170]), .B(c8170), .Z(n24512) );
XOR U40855 ( .A(c8171), .B(n24513), .Z(c8172) );
ANDN U40856 ( .B(n24514), .A(n24515), .Z(n24513) );
XOR U40857 ( .A(c8171), .B(b[8171]), .Z(n24514) );
XNOR U40858 ( .A(b[8171]), .B(n24515), .Z(c[8171]) );
XNOR U40859 ( .A(a[8171]), .B(c8171), .Z(n24515) );
XOR U40860 ( .A(c8172), .B(n24516), .Z(c8173) );
ANDN U40861 ( .B(n24517), .A(n24518), .Z(n24516) );
XOR U40862 ( .A(c8172), .B(b[8172]), .Z(n24517) );
XNOR U40863 ( .A(b[8172]), .B(n24518), .Z(c[8172]) );
XNOR U40864 ( .A(a[8172]), .B(c8172), .Z(n24518) );
XOR U40865 ( .A(c8173), .B(n24519), .Z(c8174) );
ANDN U40866 ( .B(n24520), .A(n24521), .Z(n24519) );
XOR U40867 ( .A(c8173), .B(b[8173]), .Z(n24520) );
XNOR U40868 ( .A(b[8173]), .B(n24521), .Z(c[8173]) );
XNOR U40869 ( .A(a[8173]), .B(c8173), .Z(n24521) );
XOR U40870 ( .A(c8174), .B(n24522), .Z(c8175) );
ANDN U40871 ( .B(n24523), .A(n24524), .Z(n24522) );
XOR U40872 ( .A(c8174), .B(b[8174]), .Z(n24523) );
XNOR U40873 ( .A(b[8174]), .B(n24524), .Z(c[8174]) );
XNOR U40874 ( .A(a[8174]), .B(c8174), .Z(n24524) );
XOR U40875 ( .A(c8175), .B(n24525), .Z(c8176) );
ANDN U40876 ( .B(n24526), .A(n24527), .Z(n24525) );
XOR U40877 ( .A(c8175), .B(b[8175]), .Z(n24526) );
XNOR U40878 ( .A(b[8175]), .B(n24527), .Z(c[8175]) );
XNOR U40879 ( .A(a[8175]), .B(c8175), .Z(n24527) );
XOR U40880 ( .A(c8176), .B(n24528), .Z(c8177) );
ANDN U40881 ( .B(n24529), .A(n24530), .Z(n24528) );
XOR U40882 ( .A(c8176), .B(b[8176]), .Z(n24529) );
XNOR U40883 ( .A(b[8176]), .B(n24530), .Z(c[8176]) );
XNOR U40884 ( .A(a[8176]), .B(c8176), .Z(n24530) );
XOR U40885 ( .A(c8177), .B(n24531), .Z(c8178) );
ANDN U40886 ( .B(n24532), .A(n24533), .Z(n24531) );
XOR U40887 ( .A(c8177), .B(b[8177]), .Z(n24532) );
XNOR U40888 ( .A(b[8177]), .B(n24533), .Z(c[8177]) );
XNOR U40889 ( .A(a[8177]), .B(c8177), .Z(n24533) );
XOR U40890 ( .A(c8178), .B(n24534), .Z(c8179) );
ANDN U40891 ( .B(n24535), .A(n24536), .Z(n24534) );
XOR U40892 ( .A(c8178), .B(b[8178]), .Z(n24535) );
XNOR U40893 ( .A(b[8178]), .B(n24536), .Z(c[8178]) );
XNOR U40894 ( .A(a[8178]), .B(c8178), .Z(n24536) );
XOR U40895 ( .A(c8179), .B(n24537), .Z(c8180) );
ANDN U40896 ( .B(n24538), .A(n24539), .Z(n24537) );
XOR U40897 ( .A(c8179), .B(b[8179]), .Z(n24538) );
XNOR U40898 ( .A(b[8179]), .B(n24539), .Z(c[8179]) );
XNOR U40899 ( .A(a[8179]), .B(c8179), .Z(n24539) );
XOR U40900 ( .A(c8180), .B(n24540), .Z(c8181) );
ANDN U40901 ( .B(n24541), .A(n24542), .Z(n24540) );
XOR U40902 ( .A(c8180), .B(b[8180]), .Z(n24541) );
XNOR U40903 ( .A(b[8180]), .B(n24542), .Z(c[8180]) );
XNOR U40904 ( .A(a[8180]), .B(c8180), .Z(n24542) );
XOR U40905 ( .A(c8181), .B(n24543), .Z(c8182) );
ANDN U40906 ( .B(n24544), .A(n24545), .Z(n24543) );
XOR U40907 ( .A(c8181), .B(b[8181]), .Z(n24544) );
XNOR U40908 ( .A(b[8181]), .B(n24545), .Z(c[8181]) );
XNOR U40909 ( .A(a[8181]), .B(c8181), .Z(n24545) );
XOR U40910 ( .A(c8182), .B(n24546), .Z(c8183) );
ANDN U40911 ( .B(n24547), .A(n24548), .Z(n24546) );
XOR U40912 ( .A(c8182), .B(b[8182]), .Z(n24547) );
XNOR U40913 ( .A(b[8182]), .B(n24548), .Z(c[8182]) );
XNOR U40914 ( .A(a[8182]), .B(c8182), .Z(n24548) );
XOR U40915 ( .A(c8183), .B(n24549), .Z(c8184) );
ANDN U40916 ( .B(n24550), .A(n24551), .Z(n24549) );
XOR U40917 ( .A(c8183), .B(b[8183]), .Z(n24550) );
XNOR U40918 ( .A(b[8183]), .B(n24551), .Z(c[8183]) );
XNOR U40919 ( .A(a[8183]), .B(c8183), .Z(n24551) );
XOR U40920 ( .A(c8184), .B(n24552), .Z(c8185) );
ANDN U40921 ( .B(n24553), .A(n24554), .Z(n24552) );
XOR U40922 ( .A(c8184), .B(b[8184]), .Z(n24553) );
XNOR U40923 ( .A(b[8184]), .B(n24554), .Z(c[8184]) );
XNOR U40924 ( .A(a[8184]), .B(c8184), .Z(n24554) );
XOR U40925 ( .A(c8185), .B(n24555), .Z(c8186) );
ANDN U40926 ( .B(n24556), .A(n24557), .Z(n24555) );
XOR U40927 ( .A(c8185), .B(b[8185]), .Z(n24556) );
XNOR U40928 ( .A(b[8185]), .B(n24557), .Z(c[8185]) );
XNOR U40929 ( .A(a[8185]), .B(c8185), .Z(n24557) );
XOR U40930 ( .A(c8186), .B(n24558), .Z(c8187) );
ANDN U40931 ( .B(n24559), .A(n24560), .Z(n24558) );
XOR U40932 ( .A(c8186), .B(b[8186]), .Z(n24559) );
XNOR U40933 ( .A(b[8186]), .B(n24560), .Z(c[8186]) );
XNOR U40934 ( .A(a[8186]), .B(c8186), .Z(n24560) );
XOR U40935 ( .A(c8187), .B(n24561), .Z(c8188) );
ANDN U40936 ( .B(n24562), .A(n24563), .Z(n24561) );
XOR U40937 ( .A(c8187), .B(b[8187]), .Z(n24562) );
XNOR U40938 ( .A(b[8187]), .B(n24563), .Z(c[8187]) );
XNOR U40939 ( .A(a[8187]), .B(c8187), .Z(n24563) );
XOR U40940 ( .A(c8188), .B(n24564), .Z(c8189) );
ANDN U40941 ( .B(n24565), .A(n24566), .Z(n24564) );
XOR U40942 ( .A(c8188), .B(b[8188]), .Z(n24565) );
XNOR U40943 ( .A(b[8188]), .B(n24566), .Z(c[8188]) );
XNOR U40944 ( .A(a[8188]), .B(c8188), .Z(n24566) );
XOR U40945 ( .A(c8189), .B(n24567), .Z(c8190) );
ANDN U40946 ( .B(n24568), .A(n24569), .Z(n24567) );
XOR U40947 ( .A(c8189), .B(b[8189]), .Z(n24568) );
XNOR U40948 ( .A(b[8189]), .B(n24569), .Z(c[8189]) );
XNOR U40949 ( .A(a[8189]), .B(c8189), .Z(n24569) );
XOR U40950 ( .A(c8190), .B(n24570), .Z(c8191) );
ANDN U40951 ( .B(n24571), .A(n24572), .Z(n24570) );
XOR U40952 ( .A(c8190), .B(b[8190]), .Z(n24571) );
XNOR U40953 ( .A(b[8190]), .B(n24572), .Z(c[8190]) );
XNOR U40954 ( .A(a[8190]), .B(c8190), .Z(n24572) );
XOR U40955 ( .A(c8191), .B(n24573), .Z(c8192) );
ANDN U40956 ( .B(n24574), .A(n24575), .Z(n24573) );
XOR U40957 ( .A(c8191), .B(b[8191]), .Z(n24574) );
XNOR U40958 ( .A(b[8191]), .B(n24575), .Z(c[8191]) );
XNOR U40959 ( .A(a[8191]), .B(c8191), .Z(n24575) );


endmodule
