
module hamming_N1600_CC1 ( clk, rst, x, y, o );
  input [1599:0] x;
  input [1599:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567;

  NAND U1601 ( .A(n1290), .B(n1289), .Z(n1) );
  NAND U1602 ( .A(n1287), .B(n1288), .Z(n2) );
  NAND U1603 ( .A(n1), .B(n2), .Z(n5955) );
  NAND U1604 ( .A(n1053), .B(n1052), .Z(n3) );
  NAND U1605 ( .A(n1050), .B(n1051), .Z(n4) );
  AND U1606 ( .A(n3), .B(n4), .Z(n5948) );
  NAND U1607 ( .A(n3421), .B(n3420), .Z(n5) );
  NAND U1608 ( .A(n3418), .B(n3419), .Z(n6) );
  AND U1609 ( .A(n5), .B(n6), .Z(n6853) );
  NAND U1610 ( .A(n3489), .B(n3488), .Z(n7) );
  NAND U1611 ( .A(n3486), .B(n3487), .Z(n8) );
  NAND U1612 ( .A(n7), .B(n8), .Z(n6442) );
  NAND U1613 ( .A(n4303), .B(n4302), .Z(n9) );
  NAND U1614 ( .A(n4300), .B(n4301), .Z(n10) );
  AND U1615 ( .A(n9), .B(n10), .Z(n5561) );
  NAND U1616 ( .A(n3477), .B(n3476), .Z(n11) );
  NAND U1617 ( .A(n3474), .B(n3475), .Z(n12) );
  NAND U1618 ( .A(n11), .B(n12), .Z(n6112) );
  NAND U1619 ( .A(n3507), .B(n3506), .Z(n13) );
  NAND U1620 ( .A(n3504), .B(n3505), .Z(n14) );
  NAND U1621 ( .A(n13), .B(n14), .Z(n6106) );
  NAND U1622 ( .A(n5235), .B(n5234), .Z(n15) );
  NAND U1623 ( .A(n5232), .B(n5233), .Z(n16) );
  NAND U1624 ( .A(n15), .B(n16), .Z(n5869) );
  NAND U1625 ( .A(n4295), .B(n4294), .Z(n17) );
  NAND U1626 ( .A(n4292), .B(n4293), .Z(n18) );
  AND U1627 ( .A(n17), .B(n18), .Z(n5800) );
  NAND U1628 ( .A(n5624), .B(n5623), .Z(n19) );
  NAND U1629 ( .A(n5622), .B(n5621), .Z(n20) );
  NAND U1630 ( .A(n19), .B(n20), .Z(n7514) );
  NAND U1631 ( .A(n5757), .B(n5756), .Z(n21) );
  NAND U1632 ( .A(n5755), .B(n5754), .Z(n22) );
  NAND U1633 ( .A(n21), .B(n22), .Z(n8452) );
  NAND U1634 ( .A(n6750), .B(n6749), .Z(n23) );
  NAND U1635 ( .A(n6748), .B(n6747), .Z(n24) );
  NAND U1636 ( .A(n23), .B(n24), .Z(n8031) );
  NAND U1637 ( .A(n5349), .B(n5348), .Z(n25) );
  NAND U1638 ( .A(n5347), .B(n5346), .Z(n26) );
  NAND U1639 ( .A(n25), .B(n26), .Z(n8050) );
  NAND U1640 ( .A(n7094), .B(n7093), .Z(n27) );
  NAND U1641 ( .A(n7092), .B(n7091), .Z(n28) );
  NAND U1642 ( .A(n27), .B(n28), .Z(n8038) );
  NAND U1643 ( .A(n6412), .B(n6411), .Z(n29) );
  NAND U1644 ( .A(n6410), .B(n6409), .Z(n30) );
  AND U1645 ( .A(n29), .B(n30), .Z(n8260) );
  NAND U1646 ( .A(n5307), .B(n5306), .Z(n31) );
  NAND U1647 ( .A(n5305), .B(n5304), .Z(n32) );
  AND U1648 ( .A(n31), .B(n32), .Z(n8302) );
  NAND U1649 ( .A(n7566), .B(n7565), .Z(n33) );
  NAND U1650 ( .A(n7564), .B(n7563), .Z(n34) );
  AND U1651 ( .A(n33), .B(n34), .Z(n9029) );
  NAND U1652 ( .A(n8066), .B(n8065), .Z(n35) );
  NAND U1653 ( .A(n8064), .B(n8063), .Z(n36) );
  NAND U1654 ( .A(n35), .B(n36), .Z(n8788) );
  NAND U1655 ( .A(n7836), .B(n7835), .Z(n37) );
  NAND U1656 ( .A(n7834), .B(n7833), .Z(n38) );
  NAND U1657 ( .A(n37), .B(n38), .Z(n8657) );
  OR U1658 ( .A(n7679), .B(n7680), .Z(n39) );
  NAND U1659 ( .A(n7678), .B(n7677), .Z(n40) );
  NAND U1660 ( .A(n39), .B(n40), .Z(n8813) );
  NAND U1661 ( .A(n8462), .B(n8461), .Z(n41) );
  NAND U1662 ( .A(n8460), .B(n8459), .Z(n42) );
  NAND U1663 ( .A(n41), .B(n42), .Z(n9168) );
  NAND U1664 ( .A(n8651), .B(n8650), .Z(n43) );
  NAND U1665 ( .A(n8648), .B(n8649), .Z(n44) );
  AND U1666 ( .A(n43), .B(n44), .Z(n9179) );
  NAND U1667 ( .A(n9186), .B(n9187), .Z(n45) );
  NANDN U1668 ( .A(n9189), .B(n9188), .Z(n46) );
  NAND U1669 ( .A(n45), .B(n46), .Z(n9393) );
  NAND U1670 ( .A(n9475), .B(n9474), .Z(n47) );
  NAND U1671 ( .A(n9472), .B(n9473), .Z(n48) );
  AND U1672 ( .A(n47), .B(n48), .Z(n9530) );
  NAND U1673 ( .A(n9534), .B(n9533), .Z(n49) );
  NAND U1674 ( .A(n9532), .B(n9531), .Z(n50) );
  NAND U1675 ( .A(n49), .B(n50), .Z(n9560) );
  NAND U1676 ( .A(n3703), .B(n3702), .Z(n51) );
  NAND U1677 ( .A(n3700), .B(n3701), .Z(n52) );
  NAND U1678 ( .A(n51), .B(n52), .Z(n6770) );
  NAND U1679 ( .A(n1286), .B(n1285), .Z(n53) );
  NAND U1680 ( .A(n1283), .B(n1284), .Z(n54) );
  AND U1681 ( .A(n53), .B(n54), .Z(n5954) );
  NAND U1682 ( .A(n1064), .B(n1063), .Z(n55) );
  NAND U1683 ( .A(n1061), .B(n1062), .Z(n56) );
  NAND U1684 ( .A(n55), .B(n56), .Z(n5951) );
  NAND U1685 ( .A(n4771), .B(n4770), .Z(n57) );
  NAND U1686 ( .A(n4768), .B(n4769), .Z(n58) );
  AND U1687 ( .A(n57), .B(n58), .Z(n6669) );
  NAND U1688 ( .A(n1037), .B(n1036), .Z(n59) );
  NAND U1689 ( .A(n1034), .B(n1035), .Z(n60) );
  AND U1690 ( .A(n59), .B(n60), .Z(n6847) );
  NAND U1691 ( .A(n2993), .B(n2992), .Z(n61) );
  NAND U1692 ( .A(n2990), .B(n2991), .Z(n62) );
  AND U1693 ( .A(n61), .B(n62), .Z(n5907) );
  NAND U1694 ( .A(n2505), .B(n2504), .Z(n63) );
  NAND U1695 ( .A(n2502), .B(n2503), .Z(n64) );
  AND U1696 ( .A(n63), .B(n64), .Z(n6452) );
  NAND U1697 ( .A(n3485), .B(n3484), .Z(n65) );
  NAND U1698 ( .A(n3482), .B(n3483), .Z(n66) );
  AND U1699 ( .A(n65), .B(n66), .Z(n6441) );
  NAND U1700 ( .A(n4307), .B(n4306), .Z(n67) );
  NAND U1701 ( .A(n4304), .B(n4305), .Z(n68) );
  AND U1702 ( .A(n67), .B(n68), .Z(n5560) );
  NAND U1703 ( .A(n3473), .B(n3472), .Z(n69) );
  NAND U1704 ( .A(n3470), .B(n3471), .Z(n70) );
  AND U1705 ( .A(n69), .B(n70), .Z(n6111) );
  NAND U1706 ( .A(n3503), .B(n3502), .Z(n71) );
  NAND U1707 ( .A(n3500), .B(n3501), .Z(n72) );
  AND U1708 ( .A(n71), .B(n72), .Z(n6105) );
  NAND U1709 ( .A(n3589), .B(n3588), .Z(n73) );
  NAND U1710 ( .A(n3586), .B(n3587), .Z(n74) );
  AND U1711 ( .A(n73), .B(n74), .Z(n6707) );
  NAND U1712 ( .A(n4775), .B(n4774), .Z(n75) );
  NAND U1713 ( .A(n4772), .B(n4773), .Z(n76) );
  AND U1714 ( .A(n75), .B(n76), .Z(n6654) );
  NAND U1715 ( .A(n3581), .B(n3580), .Z(n77) );
  NAND U1716 ( .A(n3578), .B(n3579), .Z(n78) );
  NAND U1717 ( .A(n77), .B(n78), .Z(n6642) );
  NAND U1718 ( .A(n3915), .B(n3914), .Z(n79) );
  NAND U1719 ( .A(n3912), .B(n3913), .Z(n80) );
  NAND U1720 ( .A(n79), .B(n80), .Z(n5893) );
  NAND U1721 ( .A(n5231), .B(n5230), .Z(n81) );
  NAND U1722 ( .A(n5228), .B(n5229), .Z(n82) );
  AND U1723 ( .A(n81), .B(n82), .Z(n5868) );
  NAND U1724 ( .A(n1981), .B(n1980), .Z(n83) );
  NAND U1725 ( .A(n1978), .B(n1979), .Z(n84) );
  NAND U1726 ( .A(n83), .B(n84), .Z(n5989) );
  NAND U1727 ( .A(n991), .B(n990), .Z(n85) );
  NAND U1728 ( .A(n988), .B(n989), .Z(n86) );
  AND U1729 ( .A(n85), .B(n86), .Z(n6329) );
  NAND U1730 ( .A(n2419), .B(n2418), .Z(n87) );
  NAND U1731 ( .A(n2416), .B(n2417), .Z(n88) );
  AND U1732 ( .A(n87), .B(n88), .Z(n6913) );
  NAND U1733 ( .A(n1862), .B(n1861), .Z(n89) );
  NAND U1734 ( .A(n1859), .B(n1860), .Z(n90) );
  NAND U1735 ( .A(n89), .B(n90), .Z(n6046) );
  NAND U1736 ( .A(n3033), .B(n3032), .Z(n91) );
  NAND U1737 ( .A(n3031), .B(n3030), .Z(n92) );
  NAND U1738 ( .A(n91), .B(n92), .Z(n5782) );
  NAND U1739 ( .A(n1638), .B(n1637), .Z(n93) );
  NANDN U1740 ( .A(n1636), .B(n1635), .Z(n94) );
  NAND U1741 ( .A(n93), .B(n94), .Z(n5695) );
  NAND U1742 ( .A(n1537), .B(n1538), .Z(n95) );
  NANDN U1743 ( .A(n1540), .B(n1539), .Z(n96) );
  NAND U1744 ( .A(n95), .B(n96), .Z(n7205) );
  NAND U1745 ( .A(n4955), .B(n4954), .Z(n97) );
  NANDN U1746 ( .A(n4953), .B(n4952), .Z(n98) );
  NAND U1747 ( .A(n97), .B(n98), .Z(n5536) );
  NAND U1748 ( .A(n5031), .B(n5030), .Z(n99) );
  NAND U1749 ( .A(n5028), .B(n5029), .Z(n100) );
  AND U1750 ( .A(n99), .B(n100), .Z(n6044) );
  NAND U1751 ( .A(n1905), .B(n1904), .Z(n101) );
  NAND U1752 ( .A(n1902), .B(n1903), .Z(n102) );
  NAND U1753 ( .A(n101), .B(n102), .Z(n6084) );
  NAND U1754 ( .A(n5173), .B(n5172), .Z(n103) );
  NANDN U1755 ( .A(n5171), .B(n5170), .Z(n104) );
  NAND U1756 ( .A(n103), .B(n104), .Z(n6905) );
  NAND U1757 ( .A(n5285), .B(n5284), .Z(n105) );
  NAND U1758 ( .A(n5283), .B(n5282), .Z(n106) );
  NAND U1759 ( .A(n105), .B(n106), .Z(n6360) );
  NAND U1760 ( .A(n4901), .B(n4900), .Z(n107) );
  NAND U1761 ( .A(n4899), .B(n4898), .Z(n108) );
  NAND U1762 ( .A(n107), .B(n108), .Z(n5944) );
  NAND U1763 ( .A(n6856), .B(n6855), .Z(n109) );
  NAND U1764 ( .A(n6854), .B(n6853), .Z(n110) );
  NAND U1765 ( .A(n109), .B(n110), .Z(n8251) );
  NAND U1766 ( .A(n7146), .B(n7145), .Z(n111) );
  NAND U1767 ( .A(n7144), .B(n7143), .Z(n112) );
  NAND U1768 ( .A(n111), .B(n112), .Z(n8179) );
  NAND U1769 ( .A(n7262), .B(n7261), .Z(n113) );
  NAND U1770 ( .A(n7260), .B(n7259), .Z(n114) );
  NAND U1771 ( .A(n113), .B(n114), .Z(n7586) );
  NAND U1772 ( .A(n6001), .B(n6000), .Z(n115) );
  NAND U1773 ( .A(n5999), .B(n5998), .Z(n116) );
  NAND U1774 ( .A(n115), .B(n116), .Z(n7630) );
  NAND U1775 ( .A(n6746), .B(n6745), .Z(n117) );
  NAND U1776 ( .A(n6743), .B(n6744), .Z(n118) );
  AND U1777 ( .A(n117), .B(n118), .Z(n8032) );
  NAND U1778 ( .A(n6055), .B(n6054), .Z(n119) );
  NAND U1779 ( .A(n6053), .B(n6052), .Z(n120) );
  NAND U1780 ( .A(n119), .B(n120), .Z(n8456) );
  XNOR U1781 ( .A(n7674), .B(n7673), .Z(n8055) );
  NAND U1782 ( .A(n5345), .B(n5344), .Z(n121) );
  NAND U1783 ( .A(n5343), .B(n5342), .Z(n122) );
  AND U1784 ( .A(n121), .B(n122), .Z(n8049) );
  NAND U1785 ( .A(n7090), .B(n7089), .Z(n123) );
  NAND U1786 ( .A(n7088), .B(n7087), .Z(n124) );
  AND U1787 ( .A(n123), .B(n124), .Z(n8037) );
  NAND U1788 ( .A(n7370), .B(n7369), .Z(n125) );
  NAND U1789 ( .A(n7368), .B(n7367), .Z(n126) );
  AND U1790 ( .A(n125), .B(n126), .Z(n8278) );
  XNOR U1791 ( .A(n8440), .B(n8439), .Z(n8259) );
  NAND U1792 ( .A(n6392), .B(n6391), .Z(n127) );
  NANDN U1793 ( .A(n6390), .B(n6389), .Z(n128) );
  AND U1794 ( .A(n127), .B(n128), .Z(n7499) );
  NAND U1795 ( .A(n5583), .B(n5582), .Z(n129) );
  NAND U1796 ( .A(n5580), .B(n5581), .Z(n130) );
  AND U1797 ( .A(n129), .B(n130), .Z(n7996) );
  NAND U1798 ( .A(n6082), .B(n6081), .Z(n131) );
  NAND U1799 ( .A(n6080), .B(n6079), .Z(n132) );
  NAND U1800 ( .A(n131), .B(n132), .Z(n7683) );
  NAND U1801 ( .A(n5317), .B(n5316), .Z(n133) );
  NAND U1802 ( .A(n5315), .B(n5314), .Z(n134) );
  AND U1803 ( .A(n133), .B(n134), .Z(n8303) );
  NAND U1804 ( .A(n5327), .B(n5326), .Z(n135) );
  NAND U1805 ( .A(n5325), .B(n5324), .Z(n136) );
  AND U1806 ( .A(n135), .B(n136), .Z(n8292) );
  NAND U1807 ( .A(n7470), .B(n7469), .Z(n137) );
  NAND U1808 ( .A(n7468), .B(n7467), .Z(n138) );
  AND U1809 ( .A(n137), .B(n138), .Z(n9020) );
  NAND U1810 ( .A(n7637), .B(n7638), .Z(n139) );
  NANDN U1811 ( .A(n7640), .B(n7639), .Z(n140) );
  NAND U1812 ( .A(n139), .B(n140), .Z(n8577) );
  NAND U1813 ( .A(n7546), .B(n7545), .Z(n141) );
  NAND U1814 ( .A(n7544), .B(n7543), .Z(n142) );
  AND U1815 ( .A(n141), .B(n142), .Z(n8570) );
  NAND U1816 ( .A(n5775), .B(n5774), .Z(n143) );
  NAND U1817 ( .A(n5773), .B(n5772), .Z(n144) );
  NAND U1818 ( .A(n143), .B(n144), .Z(n8460) );
  NAND U1819 ( .A(n8110), .B(n8109), .Z(n145) );
  NAND U1820 ( .A(n8108), .B(n8107), .Z(n146) );
  NAND U1821 ( .A(n145), .B(n146), .Z(n8616) );
  XNOR U1822 ( .A(n8825), .B(n8824), .Z(n8826) );
  NAND U1823 ( .A(n8258), .B(n8257), .Z(n147) );
  NAND U1824 ( .A(n8256), .B(n8255), .Z(n148) );
  AND U1825 ( .A(n147), .B(n148), .Z(n8964) );
  NAND U1826 ( .A(n7616), .B(n7615), .Z(n149) );
  NAND U1827 ( .A(n7613), .B(n7614), .Z(n150) );
  AND U1828 ( .A(n149), .B(n150), .Z(n8729) );
  NAND U1829 ( .A(n8963), .B(n8962), .Z(n151) );
  NAND U1830 ( .A(n8961), .B(n8960), .Z(n152) );
  NAND U1831 ( .A(n151), .B(n152), .Z(n9172) );
  AND U1832 ( .A(n8640), .B(n8641), .Z(n9171) );
  NAND U1833 ( .A(n8655), .B(n8654), .Z(n153) );
  NAND U1834 ( .A(n8652), .B(n8653), .Z(n154) );
  AND U1835 ( .A(n153), .B(n154), .Z(n9178) );
  NAND U1836 ( .A(n8656), .B(n8657), .Z(n155) );
  NANDN U1837 ( .A(n8659), .B(n8658), .Z(n156) );
  AND U1838 ( .A(n155), .B(n156), .Z(n9221) );
  NAND U1839 ( .A(n9185), .B(n9184), .Z(n157) );
  NAND U1840 ( .A(n9183), .B(n9182), .Z(n158) );
  AND U1841 ( .A(n157), .B(n158), .Z(n9385) );
  NAND U1842 ( .A(n9227), .B(n9226), .Z(n159) );
  NAND U1843 ( .A(n9225), .B(n9224), .Z(n160) );
  AND U1844 ( .A(n159), .B(n160), .Z(n9396) );
  NAND U1845 ( .A(n7694), .B(n7693), .Z(n161) );
  NAND U1846 ( .A(n7691), .B(n7692), .Z(n162) );
  NAND U1847 ( .A(n161), .B(n162), .Z(n8670) );
  NAND U1848 ( .A(n9394), .B(n9393), .Z(n163) );
  NAND U1849 ( .A(n9392), .B(n9391), .Z(n164) );
  NAND U1850 ( .A(n163), .B(n164), .Z(n9492) );
  NAND U1851 ( .A(n9530), .B(n9529), .Z(n165) );
  NAND U1852 ( .A(n9527), .B(n9528), .Z(n166) );
  NAND U1853 ( .A(n165), .B(n166), .Z(n9562) );
  XOR U1854 ( .A(n9469), .B(n9468), .Z(n9523) );
  XNOR U1855 ( .A(n1478), .B(n1477), .Z(n1479) );
  XNOR U1856 ( .A(n5153), .B(n5152), .Z(n5154) );
  NAND U1857 ( .A(n2175), .B(n2174), .Z(n167) );
  NAND U1858 ( .A(n2172), .B(n2173), .Z(n168) );
  NAND U1859 ( .A(n167), .B(n168), .Z(n5720) );
  NAND U1860 ( .A(n1710), .B(n1709), .Z(n169) );
  NAND U1861 ( .A(n1707), .B(n1708), .Z(n170) );
  AND U1862 ( .A(n169), .B(n170), .Z(n6777) );
  NAND U1863 ( .A(n3699), .B(n3698), .Z(n171) );
  NAND U1864 ( .A(n3696), .B(n3697), .Z(n172) );
  AND U1865 ( .A(n171), .B(n172), .Z(n6769) );
  NAND U1866 ( .A(n3759), .B(n3758), .Z(n173) );
  NAND U1867 ( .A(n3756), .B(n3757), .Z(n174) );
  NAND U1868 ( .A(n173), .B(n174), .Z(n6764) );
  NAND U1869 ( .A(n2715), .B(n2714), .Z(n175) );
  NAND U1870 ( .A(n2712), .B(n2713), .Z(n176) );
  AND U1871 ( .A(n175), .B(n176), .Z(n7303) );
  NAND U1872 ( .A(n3551), .B(n3550), .Z(n177) );
  NAND U1873 ( .A(n3548), .B(n3549), .Z(n178) );
  NAND U1874 ( .A(n177), .B(n178), .Z(n6662) );
  NAND U1875 ( .A(n1298), .B(n1297), .Z(n179) );
  NAND U1876 ( .A(n1295), .B(n1296), .Z(n180) );
  AND U1877 ( .A(n179), .B(n180), .Z(n6801) );
  NAND U1878 ( .A(n2545), .B(n2544), .Z(n181) );
  NAND U1879 ( .A(n2542), .B(n2543), .Z(n182) );
  NAND U1880 ( .A(n181), .B(n182), .Z(n6404) );
  NAND U1881 ( .A(n2861), .B(n2860), .Z(n183) );
  NAND U1882 ( .A(n2858), .B(n2859), .Z(n184) );
  AND U1883 ( .A(n183), .B(n184), .Z(n5904) );
  NAND U1884 ( .A(n4367), .B(n4366), .Z(n185) );
  NAND U1885 ( .A(n4364), .B(n4365), .Z(n186) );
  AND U1886 ( .A(n185), .B(n186), .Z(n5898) );
  NAND U1887 ( .A(n3493), .B(n3492), .Z(n187) );
  NAND U1888 ( .A(n3490), .B(n3491), .Z(n188) );
  NAND U1889 ( .A(n187), .B(n188), .Z(n6444) );
  NAND U1890 ( .A(n4311), .B(n4310), .Z(n189) );
  NAND U1891 ( .A(n4308), .B(n4309), .Z(n190) );
  AND U1892 ( .A(n189), .B(n190), .Z(n5562) );
  NAND U1893 ( .A(n4795), .B(n4794), .Z(n191) );
  NAND U1894 ( .A(n4792), .B(n4793), .Z(n192) );
  NAND U1895 ( .A(n191), .B(n192), .Z(n6118) );
  NAND U1896 ( .A(n3481), .B(n3480), .Z(n193) );
  NAND U1897 ( .A(n3478), .B(n3479), .Z(n194) );
  NAND U1898 ( .A(n193), .B(n194), .Z(n6114) );
  NAND U1899 ( .A(n3511), .B(n3510), .Z(n195) );
  NAND U1900 ( .A(n3508), .B(n3509), .Z(n196) );
  NAND U1901 ( .A(n195), .B(n196), .Z(n6108) );
  NAND U1902 ( .A(n5063), .B(n5062), .Z(n197) );
  NAND U1903 ( .A(n5060), .B(n5061), .Z(n198) );
  AND U1904 ( .A(n197), .B(n198), .Z(n6717) );
  NAND U1905 ( .A(n4509), .B(n4508), .Z(n199) );
  NAND U1906 ( .A(n4506), .B(n4507), .Z(n200) );
  AND U1907 ( .A(n199), .B(n200), .Z(n6713) );
  NAND U1908 ( .A(n4783), .B(n4782), .Z(n201) );
  NAND U1909 ( .A(n4780), .B(n4781), .Z(n202) );
  AND U1910 ( .A(n201), .B(n202), .Z(n6655) );
  NAND U1911 ( .A(n3919), .B(n3918), .Z(n203) );
  NAND U1912 ( .A(n3916), .B(n3917), .Z(n204) );
  NAND U1913 ( .A(n203), .B(n204), .Z(n5895) );
  NAND U1914 ( .A(n4219), .B(n4218), .Z(n205) );
  NAND U1915 ( .A(n4216), .B(n4217), .Z(n206) );
  AND U1916 ( .A(n205), .B(n206), .Z(n5751) );
  NAND U1917 ( .A(n1886), .B(n1885), .Z(n207) );
  NAND U1918 ( .A(n1883), .B(n1884), .Z(n208) );
  AND U1919 ( .A(n207), .B(n208), .Z(n6063) );
  AND U1920 ( .A(n1881), .B(n1882), .Z(n6062) );
  NAND U1921 ( .A(n3875), .B(n3874), .Z(n209) );
  NAND U1922 ( .A(n3872), .B(n3873), .Z(n210) );
  AND U1923 ( .A(n209), .B(n210), .Z(n6145) );
  NAND U1924 ( .A(n4139), .B(n4138), .Z(n211) );
  NAND U1925 ( .A(n4136), .B(n4137), .Z(n212) );
  NAND U1926 ( .A(n211), .B(n212), .Z(n5879) );
  NAND U1927 ( .A(n4019), .B(n4018), .Z(n213) );
  NAND U1928 ( .A(n4016), .B(n4017), .Z(n214) );
  AND U1929 ( .A(n213), .B(n214), .Z(n7333) );
  NAND U1930 ( .A(n4727), .B(n4726), .Z(n215) );
  NAND U1931 ( .A(n4724), .B(n4725), .Z(n216) );
  AND U1932 ( .A(n215), .B(n216), .Z(n5444) );
  NAND U1933 ( .A(n4731), .B(n4730), .Z(n217) );
  NAND U1934 ( .A(n4728), .B(n4729), .Z(n218) );
  AND U1935 ( .A(n217), .B(n218), .Z(n5439) );
  NAND U1936 ( .A(n987), .B(n986), .Z(n219) );
  NAND U1937 ( .A(n984), .B(n985), .Z(n220) );
  AND U1938 ( .A(n219), .B(n220), .Z(n6327) );
  NAND U1939 ( .A(n4929), .B(n4928), .Z(n221) );
  NAND U1940 ( .A(n4926), .B(n4927), .Z(n222) );
  AND U1941 ( .A(n221), .B(n222), .Z(n6053) );
  NAND U1942 ( .A(n3011), .B(n3010), .Z(n223) );
  NAND U1943 ( .A(n3008), .B(n3009), .Z(n224) );
  AND U1944 ( .A(n223), .B(n224), .Z(n5785) );
  NAND U1945 ( .A(n1634), .B(n1633), .Z(n225) );
  NAND U1946 ( .A(n1631), .B(n1632), .Z(n226) );
  AND U1947 ( .A(n225), .B(n226), .Z(n5696) );
  NAND U1948 ( .A(n1536), .B(n1535), .Z(n227) );
  NAND U1949 ( .A(n1533), .B(n1534), .Z(n228) );
  AND U1950 ( .A(n227), .B(n228), .Z(n7206) );
  NAND U1951 ( .A(n2079), .B(n2078), .Z(n229) );
  NAND U1952 ( .A(n2077), .B(n2076), .Z(n230) );
  NAND U1953 ( .A(n229), .B(n230), .Z(n6841) );
  NAND U1954 ( .A(n1172), .B(n1171), .Z(n231) );
  NAND U1955 ( .A(n1170), .B(n1169), .Z(n232) );
  NAND U1956 ( .A(n231), .B(n232), .Z(n6723) );
  NAND U1957 ( .A(n4569), .B(n4568), .Z(n233) );
  NAND U1958 ( .A(n4567), .B(n4566), .Z(n234) );
  NAND U1959 ( .A(n233), .B(n234), .Z(n7165) );
  NAND U1960 ( .A(n4339), .B(n4338), .Z(n235) );
  NAND U1961 ( .A(n4336), .B(n4337), .Z(n236) );
  AND U1962 ( .A(n235), .B(n236), .Z(n5580) );
  NAND U1963 ( .A(n1901), .B(n1900), .Z(n237) );
  NAND U1964 ( .A(n1898), .B(n1899), .Z(n238) );
  AND U1965 ( .A(n237), .B(n238), .Z(n6083) );
  NAND U1966 ( .A(n4823), .B(n4822), .Z(n239) );
  NAND U1967 ( .A(n4821), .B(n4820), .Z(n240) );
  NAND U1968 ( .A(n239), .B(n240), .Z(n6899) );
  NAND U1969 ( .A(n2355), .B(n2354), .Z(n241) );
  NAND U1970 ( .A(n2353), .B(n2352), .Z(n242) );
  NAND U1971 ( .A(n241), .B(n242), .Z(n6337) );
  NAND U1972 ( .A(n1810), .B(n1809), .Z(n243) );
  NAND U1973 ( .A(n1808), .B(n1807), .Z(n244) );
  NAND U1974 ( .A(n243), .B(n244), .Z(n5941) );
  NAND U1975 ( .A(n5103), .B(n5102), .Z(n245) );
  NAND U1976 ( .A(n5101), .B(n5100), .Z(n246) );
  NAND U1977 ( .A(n245), .B(n246), .Z(n6791) );
  NAND U1978 ( .A(n6670), .B(n6669), .Z(n247) );
  NAND U1979 ( .A(n6668), .B(n6667), .Z(n248) );
  NAND U1980 ( .A(n247), .B(n248), .Z(n7461) );
  NAND U1981 ( .A(n6800), .B(n6799), .Z(n249) );
  NAND U1982 ( .A(n6798), .B(n6797), .Z(n250) );
  NAND U1983 ( .A(n249), .B(n250), .Z(n8249) );
  NAND U1984 ( .A(n6640), .B(n6639), .Z(n251) );
  NAND U1985 ( .A(n6638), .B(n6637), .Z(n252) );
  NAND U1986 ( .A(n251), .B(n252), .Z(n7641) );
  NAND U1987 ( .A(n5909), .B(n5908), .Z(n253) );
  NAND U1988 ( .A(n5907), .B(n5906), .Z(n254) );
  NAND U1989 ( .A(n253), .B(n254), .Z(n7547) );
  NAND U1990 ( .A(n6454), .B(n6453), .Z(n255) );
  NAND U1991 ( .A(n6452), .B(n6451), .Z(n256) );
  NAND U1992 ( .A(n255), .B(n256), .Z(n7510) );
  NAND U1993 ( .A(n5891), .B(n5890), .Z(n257) );
  NAND U1994 ( .A(n5888), .B(n5889), .Z(n258) );
  AND U1995 ( .A(n257), .B(n258), .Z(n7596) );
  NAND U1996 ( .A(n6916), .B(n6915), .Z(n259) );
  NAND U1997 ( .A(n6914), .B(n6913), .Z(n260) );
  AND U1998 ( .A(n259), .B(n260), .Z(n8432) );
  NAND U1999 ( .A(n6434), .B(n6433), .Z(n261) );
  NANDN U2000 ( .A(n6432), .B(n6431), .Z(n262) );
  NAND U2001 ( .A(n261), .B(n262), .Z(n8262) );
  NAND U2002 ( .A(n6388), .B(n6387), .Z(n263) );
  NAND U2003 ( .A(n6386), .B(n6385), .Z(n264) );
  AND U2004 ( .A(n263), .B(n264), .Z(n7501) );
  XNOR U2005 ( .A(n6370), .B(n6369), .Z(n6372) );
  NAND U2006 ( .A(n5579), .B(n5578), .Z(n265) );
  NAND U2007 ( .A(n5576), .B(n5577), .Z(n266) );
  AND U2008 ( .A(n265), .B(n266), .Z(n7998) );
  NAND U2009 ( .A(n5803), .B(n5802), .Z(n267) );
  NAND U2010 ( .A(n5800), .B(n5801), .Z(n268) );
  AND U2011 ( .A(n267), .B(n268), .Z(n7672) );
  NAND U2012 ( .A(n6908), .B(n6907), .Z(n269) );
  NAND U2013 ( .A(n6906), .B(n6905), .Z(n270) );
  AND U2014 ( .A(n269), .B(n270), .Z(n8295) );
  NAND U2015 ( .A(n5337), .B(n5336), .Z(n271) );
  NAND U2016 ( .A(n5335), .B(n5334), .Z(n272) );
  AND U2017 ( .A(n271), .B(n272), .Z(n8293) );
  NAND U2018 ( .A(n6362), .B(n6361), .Z(n273) );
  NAND U2019 ( .A(n6360), .B(n6359), .Z(n274) );
  AND U2020 ( .A(n273), .B(n274), .Z(n8085) );
  NAND U2021 ( .A(n7102), .B(n7101), .Z(n275) );
  NAND U2022 ( .A(n7100), .B(n7099), .Z(n276) );
  AND U2023 ( .A(n275), .B(n276), .Z(n8077) );
  NAND U2024 ( .A(n5367), .B(n5366), .Z(n277) );
  NAND U2025 ( .A(n5365), .B(n5364), .Z(n278) );
  AND U2026 ( .A(n277), .B(n278), .Z(n8075) );
  NAND U2027 ( .A(n5947), .B(n5946), .Z(n279) );
  NAND U2028 ( .A(n5945), .B(n5944), .Z(n280) );
  AND U2029 ( .A(n279), .B(n280), .Z(n7576) );
  NAND U2030 ( .A(n7183), .B(n7184), .Z(n281) );
  NANDN U2031 ( .A(n7186), .B(n7185), .Z(n282) );
  AND U2032 ( .A(n281), .B(n282), .Z(n8336) );
  NAND U2033 ( .A(n7060), .B(n7059), .Z(n283) );
  NAND U2034 ( .A(n7058), .B(n7057), .Z(n284) );
  NAND U2035 ( .A(n283), .B(n284), .Z(n8412) );
  NAND U2036 ( .A(n5825), .B(n5824), .Z(n285) );
  NAND U2037 ( .A(n5822), .B(n5823), .Z(n286) );
  AND U2038 ( .A(n285), .B(n286), .Z(n7456) );
  NAND U2039 ( .A(n7076), .B(n7075), .Z(n287) );
  NAND U2040 ( .A(n7074), .B(n7073), .Z(n288) );
  AND U2041 ( .A(n287), .B(n288), .Z(n7811) );
  NAND U2042 ( .A(n6866), .B(n6865), .Z(n289) );
  NAND U2043 ( .A(n6864), .B(n6863), .Z(n290) );
  NAND U2044 ( .A(n289), .B(n290), .Z(n7705) );
  NAND U2045 ( .A(n7574), .B(n7573), .Z(n291) );
  NAND U2046 ( .A(n7572), .B(n7571), .Z(n292) );
  AND U2047 ( .A(n291), .B(n292), .Z(n9031) );
  NAND U2048 ( .A(n7474), .B(n7473), .Z(n293) );
  NAND U2049 ( .A(n7472), .B(n7471), .Z(n294) );
  AND U2050 ( .A(n293), .B(n294), .Z(n9022) );
  NAND U2051 ( .A(n8254), .B(n8253), .Z(n295) );
  NAND U2052 ( .A(n8252), .B(n8251), .Z(n296) );
  NAND U2053 ( .A(n295), .B(n296), .Z(n8585) );
  NAND U2054 ( .A(n7636), .B(n7635), .Z(n297) );
  NAND U2055 ( .A(n7634), .B(n7633), .Z(n298) );
  AND U2056 ( .A(n297), .B(n298), .Z(n8576) );
  NAND U2057 ( .A(n7553), .B(n7554), .Z(n299) );
  NANDN U2058 ( .A(n7556), .B(n7555), .Z(n300) );
  AND U2059 ( .A(n299), .B(n300), .Z(n8572) );
  NAND U2060 ( .A(n7516), .B(n7515), .Z(n301) );
  NAND U2061 ( .A(n7514), .B(n7513), .Z(n302) );
  AND U2062 ( .A(n301), .B(n302), .Z(n8960) );
  NAND U2063 ( .A(n7588), .B(n7587), .Z(n303) );
  NAND U2064 ( .A(n7586), .B(n7585), .Z(n304) );
  AND U2065 ( .A(n303), .B(n304), .Z(n8953) );
  NAND U2066 ( .A(n7632), .B(n7631), .Z(n305) );
  NAND U2067 ( .A(n7630), .B(n7629), .Z(n306) );
  NAND U2068 ( .A(n305), .B(n306), .Z(n8803) );
  NAND U2069 ( .A(n8430), .B(n8429), .Z(n307) );
  NAND U2070 ( .A(n8428), .B(n8427), .Z(n308) );
  AND U2071 ( .A(n307), .B(n308), .Z(n8652) );
  NAND U2072 ( .A(n8062), .B(n8061), .Z(n309) );
  NAND U2073 ( .A(n8059), .B(n8060), .Z(n310) );
  AND U2074 ( .A(n309), .B(n310), .Z(n8789) );
  NAND U2075 ( .A(n7936), .B(n7935), .Z(n311) );
  NAND U2076 ( .A(n7934), .B(n7933), .Z(n312) );
  NAND U2077 ( .A(n311), .B(n312), .Z(n8782) );
  NAND U2078 ( .A(n8106), .B(n8105), .Z(n313) );
  NAND U2079 ( .A(n8103), .B(n8104), .Z(n314) );
  AND U2080 ( .A(n313), .B(n314), .Z(n8617) );
  NAND U2081 ( .A(n8280), .B(n8279), .Z(n315) );
  NAND U2082 ( .A(n8278), .B(n8277), .Z(n316) );
  NAND U2083 ( .A(n315), .B(n316), .Z(n8986) );
  NAND U2084 ( .A(n7508), .B(n7507), .Z(n317) );
  NAND U2085 ( .A(n7506), .B(n7505), .Z(n318) );
  NAND U2086 ( .A(n317), .B(n318), .Z(n8996) );
  NAND U2087 ( .A(n6998), .B(n6997), .Z(n319) );
  NANDN U2088 ( .A(n6996), .B(n6995), .Z(n320) );
  AND U2089 ( .A(n319), .B(n320), .Z(n7527) );
  NAND U2090 ( .A(n8304), .B(n8303), .Z(n321) );
  NAND U2091 ( .A(n8302), .B(n8301), .Z(n322) );
  NAND U2092 ( .A(n321), .B(n322), .Z(n9013) );
  NAND U2093 ( .A(n7968), .B(n7967), .Z(n323) );
  NAND U2094 ( .A(n7966), .B(n7965), .Z(n324) );
  NAND U2095 ( .A(n323), .B(n324), .Z(n8830) );
  NAND U2096 ( .A(n8240), .B(n8239), .Z(n325) );
  NAND U2097 ( .A(n8238), .B(n8237), .Z(n326) );
  NAND U2098 ( .A(n325), .B(n326), .Z(n8966) );
  NAND U2099 ( .A(n7524), .B(n7523), .Z(n327) );
  NAND U2100 ( .A(n7522), .B(n7521), .Z(n328) );
  NAND U2101 ( .A(n327), .B(n328), .Z(n8751) );
  NAND U2102 ( .A(n9027), .B(n9026), .Z(n329) );
  NAND U2103 ( .A(n9025), .B(n9024), .Z(n330) );
  NAND U2104 ( .A(n329), .B(n330), .Z(n9194) );
  NAND U2105 ( .A(n8959), .B(n8958), .Z(n331) );
  NAND U2106 ( .A(n8956), .B(n8957), .Z(n332) );
  AND U2107 ( .A(n331), .B(n332), .Z(n9173) );
  NAND U2108 ( .A(n8992), .B(n8993), .Z(n333) );
  NANDN U2109 ( .A(n8995), .B(n8994), .Z(n334) );
  AND U2110 ( .A(n333), .B(n334), .Z(n9232) );
  XNOR U2111 ( .A(n8761), .B(n8760), .Z(n8763) );
  OR U2112 ( .A(n9018), .B(n9019), .Z(n335) );
  NAND U2113 ( .A(n9016), .B(n9017), .Z(n336) );
  AND U2114 ( .A(n335), .B(n336), .Z(n9214) );
  OR U2115 ( .A(n9010), .B(n9011), .Z(n337) );
  NAND U2116 ( .A(n9009), .B(n9008), .Z(n338) );
  NAND U2117 ( .A(n337), .B(n338), .Z(n9204) );
  NAND U2118 ( .A(n8947), .B(n8946), .Z(n339) );
  NAND U2119 ( .A(n8945), .B(n8944), .Z(n340) );
  NAND U2120 ( .A(n339), .B(n340), .Z(n9140) );
  NAND U2121 ( .A(n9223), .B(n9222), .Z(n341) );
  NAND U2122 ( .A(n9221), .B(n9220), .Z(n342) );
  NAND U2123 ( .A(n341), .B(n342), .Z(n9395) );
  XNOR U2124 ( .A(n9253), .B(n9252), .Z(n9255) );
  NAND U2125 ( .A(n7026), .B(n7025), .Z(n343) );
  NAND U2126 ( .A(n7023), .B(n7024), .Z(n344) );
  NAND U2127 ( .A(n343), .B(n344), .Z(n7691) );
  XNOR U2128 ( .A(n9454), .B(n9453), .Z(n9455) );
  NAND U2129 ( .A(n9416), .B(n9415), .Z(n345) );
  NAND U2130 ( .A(n9413), .B(n9414), .Z(n346) );
  AND U2131 ( .A(n345), .B(n346), .Z(n9481) );
  XOR U2132 ( .A(n9329), .B(n9328), .Z(n9331) );
  NAND U2133 ( .A(n9307), .B(n9308), .Z(n347) );
  XOR U2134 ( .A(n9307), .B(n9308), .Z(n348) );
  NANDN U2135 ( .A(n9306), .B(n348), .Z(n349) );
  NAND U2136 ( .A(n347), .B(n349), .Z(n9359) );
  NAND U2137 ( .A(n9546), .B(n9547), .Z(n350) );
  XOR U2138 ( .A(n9546), .B(n9547), .Z(n351) );
  NAND U2139 ( .A(n351), .B(n9545), .Z(n352) );
  NAND U2140 ( .A(n350), .B(n352), .Z(n9556) );
  NANDN U2141 ( .A(n9563), .B(n9562), .Z(n353) );
  NANDN U2142 ( .A(n9561), .B(n9560), .Z(n354) );
  AND U2143 ( .A(n353), .B(n354), .Z(n9564) );
  XNOR U2144 ( .A(n1644), .B(n1643), .Z(n1645) );
  XNOR U2145 ( .A(n1506), .B(n1505), .Z(n1507) );
  XNOR U2146 ( .A(n1490), .B(n1489), .Z(n1491) );
  XNOR U2147 ( .A(n5147), .B(n5146), .Z(n5148) );
  XNOR U2148 ( .A(n2527), .B(n2526), .Z(n2528) );
  XNOR U2149 ( .A(n3435), .B(n3434), .Z(n3436) );
  NAND U2150 ( .A(n1294), .B(n1293), .Z(n355) );
  NAND U2151 ( .A(n1291), .B(n1292), .Z(n356) );
  AND U2152 ( .A(n355), .B(n356), .Z(n5956) );
  NAND U2153 ( .A(n2797), .B(n2796), .Z(n357) );
  NAND U2154 ( .A(n2794), .B(n2795), .Z(n358) );
  AND U2155 ( .A(n357), .B(n358), .Z(n7319) );
  NAND U2156 ( .A(n4759), .B(n4758), .Z(n359) );
  NAND U2157 ( .A(n4756), .B(n4757), .Z(n360) );
  AND U2158 ( .A(n359), .B(n360), .Z(n7293) );
  NAND U2159 ( .A(n4763), .B(n4762), .Z(n361) );
  NAND U2160 ( .A(n4760), .B(n4761), .Z(n362) );
  AND U2161 ( .A(n361), .B(n362), .Z(n6668) );
  NAND U2162 ( .A(n3547), .B(n3546), .Z(n363) );
  NAND U2163 ( .A(n3544), .B(n3545), .Z(n364) );
  AND U2164 ( .A(n363), .B(n364), .Z(n6661) );
  NAND U2165 ( .A(n3515), .B(n3514), .Z(n365) );
  NAND U2166 ( .A(n3512), .B(n3513), .Z(n366) );
  AND U2167 ( .A(n365), .B(n366), .Z(n6397) );
  NAND U2168 ( .A(n3425), .B(n3424), .Z(n367) );
  NAND U2169 ( .A(n3422), .B(n3423), .Z(n368) );
  AND U2170 ( .A(n367), .B(n368), .Z(n6855) );
  NAND U2171 ( .A(n2997), .B(n2996), .Z(n369) );
  NAND U2172 ( .A(n2994), .B(n2995), .Z(n370) );
  AND U2173 ( .A(n369), .B(n370), .Z(n5906) );
  NAND U2174 ( .A(n1398), .B(n1397), .Z(n371) );
  NAND U2175 ( .A(n1395), .B(n1396), .Z(n372) );
  AND U2176 ( .A(n371), .B(n372), .Z(n6034) );
  NAND U2177 ( .A(n4353), .B(n4352), .Z(n373) );
  NAND U2178 ( .A(n4350), .B(n4351), .Z(n374) );
  AND U2179 ( .A(n373), .B(n374), .Z(n5621) );
  NAND U2180 ( .A(n4005), .B(n4004), .Z(n375) );
  NAND U2181 ( .A(n4002), .B(n4003), .Z(n376) );
  AND U2182 ( .A(n375), .B(n376), .Z(n7144) );
  NAND U2183 ( .A(n1580), .B(n1579), .Z(n377) );
  NAND U2184 ( .A(n1577), .B(n1578), .Z(n378) );
  AND U2185 ( .A(n377), .B(n378), .Z(n7136) );
  NAND U2186 ( .A(n4791), .B(n4790), .Z(n379) );
  NAND U2187 ( .A(n4788), .B(n4789), .Z(n380) );
  AND U2188 ( .A(n379), .B(n380), .Z(n6117) );
  NAND U2189 ( .A(n5071), .B(n5070), .Z(n381) );
  NAND U2190 ( .A(n5068), .B(n5069), .Z(n382) );
  AND U2191 ( .A(n381), .B(n382), .Z(n6719) );
  NAND U2192 ( .A(n4779), .B(n4778), .Z(n383) );
  NAND U2193 ( .A(n4776), .B(n4777), .Z(n384) );
  AND U2194 ( .A(n383), .B(n384), .Z(n6653) );
  NAND U2195 ( .A(n3577), .B(n3576), .Z(n385) );
  NAND U2196 ( .A(n3574), .B(n3575), .Z(n386) );
  AND U2197 ( .A(n385), .B(n386), .Z(n6641) );
  NAND U2198 ( .A(n3911), .B(n3910), .Z(n387) );
  NAND U2199 ( .A(n3908), .B(n3909), .Z(n388) );
  AND U2200 ( .A(n387), .B(n388), .Z(n5892) );
  NAND U2201 ( .A(n4419), .B(n4418), .Z(n389) );
  NAND U2202 ( .A(n4416), .B(n4417), .Z(n390) );
  AND U2203 ( .A(n389), .B(n390), .Z(n5888) );
  NAND U2204 ( .A(n1897), .B(n1896), .Z(n391) );
  NAND U2205 ( .A(n1895), .B(n1894), .Z(n392) );
  NAND U2206 ( .A(n391), .B(n392), .Z(n6066) );
  NAND U2207 ( .A(n1158), .B(n1157), .Z(n393) );
  NAND U2208 ( .A(n1155), .B(n1156), .Z(n394) );
  AND U2209 ( .A(n393), .B(n394), .Z(n5605) );
  NAND U2210 ( .A(n4135), .B(n4134), .Z(n395) );
  NAND U2211 ( .A(n4132), .B(n4133), .Z(n396) );
  AND U2212 ( .A(n395), .B(n396), .Z(n5878) );
  NAND U2213 ( .A(n1985), .B(n1984), .Z(n397) );
  NAND U2214 ( .A(n1982), .B(n1983), .Z(n398) );
  AND U2215 ( .A(n397), .B(n398), .Z(n5990) );
  NAND U2216 ( .A(n4023), .B(n4022), .Z(n399) );
  NAND U2217 ( .A(n4020), .B(n4021), .Z(n400) );
  NAND U2218 ( .A(n399), .B(n400), .Z(n7334) );
  NAND U2219 ( .A(n1098), .B(n1097), .Z(n401) );
  NAND U2220 ( .A(n1095), .B(n1096), .Z(n402) );
  NAND U2221 ( .A(n401), .B(n402), .Z(n6332) );
  NAND U2222 ( .A(n3953), .B(n3952), .Z(n403) );
  NAND U2223 ( .A(n3950), .B(n3951), .Z(n404) );
  AND U2224 ( .A(n403), .B(n404), .Z(n6324) );
  NAND U2225 ( .A(n4933), .B(n4932), .Z(n405) );
  NAND U2226 ( .A(n4930), .B(n4931), .Z(n406) );
  AND U2227 ( .A(n405), .B(n406), .Z(n6052) );
  NAND U2228 ( .A(n4057), .B(n4056), .Z(n407) );
  NAND U2229 ( .A(n4055), .B(n4054), .Z(n408) );
  NAND U2230 ( .A(n407), .B(n408), .Z(n5570) );
  NAND U2231 ( .A(n1560), .B(n1559), .Z(n409) );
  NAND U2232 ( .A(n1558), .B(n1557), .Z(n410) );
  AND U2233 ( .A(n409), .B(n410), .Z(n5726) );
  NAND U2234 ( .A(n1458), .B(n1457), .Z(n411) );
  NAND U2235 ( .A(n1456), .B(n1455), .Z(n412) );
  AND U2236 ( .A(n411), .B(n412), .Z(n5738) );
  NAND U2237 ( .A(n1627), .B(n1628), .Z(n413) );
  NANDN U2238 ( .A(n1630), .B(n1629), .Z(n414) );
  AND U2239 ( .A(n413), .B(n414), .Z(n5698) );
  NAND U2240 ( .A(n1529), .B(n1530), .Z(n415) );
  NANDN U2241 ( .A(n1532), .B(n1531), .Z(n416) );
  AND U2242 ( .A(n415), .B(n416), .Z(n7208) );
  NAND U2243 ( .A(n2075), .B(n2074), .Z(n417) );
  NAND U2244 ( .A(n2072), .B(n2073), .Z(n418) );
  AND U2245 ( .A(n417), .B(n418), .Z(n6842) );
  NAND U2246 ( .A(n1989), .B(n1988), .Z(n419) );
  NAND U2247 ( .A(n1987), .B(n1986), .Z(n420) );
  NAND U2248 ( .A(n419), .B(n420), .Z(n6835) );
  NAND U2249 ( .A(n4805), .B(n4804), .Z(n421) );
  NAND U2250 ( .A(n4802), .B(n4803), .Z(n422) );
  AND U2251 ( .A(n421), .B(n422), .Z(n6702) );
  NAND U2252 ( .A(n4787), .B(n4786), .Z(n423) );
  NAND U2253 ( .A(n4785), .B(n4784), .Z(n424) );
  NAND U2254 ( .A(n423), .B(n424), .Z(n6099) );
  NAND U2255 ( .A(n4557), .B(n4556), .Z(n425) );
  NAND U2256 ( .A(n4555), .B(n4554), .Z(n426) );
  NAND U2257 ( .A(n425), .B(n426), .Z(n7177) );
  NAND U2258 ( .A(n4699), .B(n4698), .Z(n427) );
  NAND U2259 ( .A(n4697), .B(n4696), .Z(n428) );
  NAND U2260 ( .A(n427), .B(n428), .Z(n7171) );
  NAND U2261 ( .A(n4565), .B(n4564), .Z(n429) );
  NAND U2262 ( .A(n4562), .B(n4563), .Z(n430) );
  AND U2263 ( .A(n429), .B(n430), .Z(n7166) );
  NAND U2264 ( .A(n4235), .B(n4234), .Z(n431) );
  NAND U2265 ( .A(n4233), .B(n4232), .Z(n432) );
  NAND U2266 ( .A(n431), .B(n432), .Z(n6193) );
  NAND U2267 ( .A(n2203), .B(n2202), .Z(n433) );
  NAND U2268 ( .A(n2201), .B(n2200), .Z(n434) );
  NAND U2269 ( .A(n433), .B(n434), .Z(n6677) );
  NAND U2270 ( .A(n2241), .B(n2240), .Z(n435) );
  NAND U2271 ( .A(n2239), .B(n2238), .Z(n436) );
  NAND U2272 ( .A(n435), .B(n436), .Z(n6671) );
  NAND U2273 ( .A(n4951), .B(n4950), .Z(n437) );
  NANDN U2274 ( .A(n4949), .B(n4948), .Z(n438) );
  AND U2275 ( .A(n437), .B(n438), .Z(n5537) );
  NAND U2276 ( .A(n2747), .B(n2746), .Z(n439) );
  NAND U2277 ( .A(n2745), .B(n2744), .Z(n440) );
  NAND U2278 ( .A(n439), .B(n440), .Z(n5380) );
  NAND U2279 ( .A(n2817), .B(n2816), .Z(n441) );
  NAND U2280 ( .A(n2815), .B(n2814), .Z(n442) );
  NAND U2281 ( .A(n441), .B(n442), .Z(n7423) );
  NAND U2282 ( .A(n5227), .B(n5226), .Z(n443) );
  NAND U2283 ( .A(n5225), .B(n5224), .Z(n444) );
  NAND U2284 ( .A(n443), .B(n444), .Z(n6387) );
  NAND U2285 ( .A(n4849), .B(n4848), .Z(n445) );
  NAND U2286 ( .A(n4847), .B(n4846), .Z(n446) );
  NAND U2287 ( .A(n445), .B(n446), .Z(n6295) );
  NAND U2288 ( .A(n1642), .B(n1641), .Z(n447) );
  NAND U2289 ( .A(n1639), .B(n1640), .Z(n448) );
  AND U2290 ( .A(n447), .B(n448), .Z(n5838) );
  NAND U2291 ( .A(n1504), .B(n1503), .Z(n449) );
  NAND U2292 ( .A(n1501), .B(n1502), .Z(n450) );
  AND U2293 ( .A(n449), .B(n450), .Z(n5832) );
  NAND U2294 ( .A(n4343), .B(n4342), .Z(n451) );
  NAND U2295 ( .A(n4340), .B(n4341), .Z(n452) );
  AND U2296 ( .A(n451), .B(n452), .Z(n5582) );
  NAND U2297 ( .A(n4445), .B(n4444), .Z(n453) );
  NAND U2298 ( .A(n4442), .B(n4443), .Z(n454) );
  NAND U2299 ( .A(n453), .B(n454), .Z(n5863) );
  NAND U2300 ( .A(n4147), .B(n4146), .Z(n455) );
  NAND U2301 ( .A(n4144), .B(n4145), .Z(n456) );
  AND U2302 ( .A(n455), .B(n456), .Z(n5856) );
  XNOR U2303 ( .A(n6420), .B(n6419), .Z(n6422) );
  NAND U2304 ( .A(n4819), .B(n4818), .Z(n457) );
  NAND U2305 ( .A(n4817), .B(n4816), .Z(n458) );
  AND U2306 ( .A(n457), .B(n458), .Z(n6900) );
  NAND U2307 ( .A(n2913), .B(n2912), .Z(n459) );
  NAND U2308 ( .A(n2911), .B(n2910), .Z(n460) );
  NAND U2309 ( .A(n459), .B(n460), .Z(n6205) );
  NAND U2310 ( .A(n1910), .B(n1911), .Z(n461) );
  NANDN U2311 ( .A(n1913), .B(n1912), .Z(n462) );
  AND U2312 ( .A(n461), .B(n462), .Z(n7269) );
  NAND U2313 ( .A(n2267), .B(n2266), .Z(n463) );
  NAND U2314 ( .A(n2265), .B(n2264), .Z(n464) );
  NAND U2315 ( .A(n463), .B(n464), .Z(n7241) );
  NAND U2316 ( .A(n5075), .B(n5074), .Z(n465) );
  NAND U2317 ( .A(n5073), .B(n5072), .Z(n466) );
  NAND U2318 ( .A(n465), .B(n466), .Z(n7129) );
  NAND U2319 ( .A(n4943), .B(n4942), .Z(n467) );
  NAND U2320 ( .A(n4941), .B(n4940), .Z(n468) );
  NAND U2321 ( .A(n467), .B(n468), .Z(n6751) );
  NAND U2322 ( .A(n1990), .B(n1991), .Z(n469) );
  NANDN U2323 ( .A(n1993), .B(n1992), .Z(n470) );
  AND U2324 ( .A(n469), .B(n470), .Z(n5985) );
  NAND U2325 ( .A(n5053), .B(n5052), .Z(n471) );
  NAND U2326 ( .A(n5051), .B(n5050), .Z(n472) );
  NAND U2327 ( .A(n471), .B(n472), .Z(n6020) );
  NAND U2328 ( .A(n3092), .B(n3093), .Z(n473) );
  NANDN U2329 ( .A(n3095), .B(n3094), .Z(n474) );
  AND U2330 ( .A(n473), .B(n474), .Z(n6989) );
  NAND U2331 ( .A(n4675), .B(n4674), .Z(n475) );
  NAND U2332 ( .A(n4673), .B(n4672), .Z(n476) );
  AND U2333 ( .A(n475), .B(n476), .Z(n6924) );
  NAND U2334 ( .A(n2917), .B(n2916), .Z(n477) );
  NAND U2335 ( .A(n2915), .B(n2914), .Z(n478) );
  NAND U2336 ( .A(n477), .B(n478), .Z(n6571) );
  NAND U2337 ( .A(n7318), .B(n7317), .Z(n479) );
  NAND U2338 ( .A(n7315), .B(n7316), .Z(n480) );
  AND U2339 ( .A(n479), .B(n480), .Z(n7488) );
  NAND U2340 ( .A(n7304), .B(n7303), .Z(n481) );
  NAND U2341 ( .A(n7302), .B(n7301), .Z(n482) );
  NAND U2342 ( .A(n481), .B(n482), .Z(n7481) );
  NAND U2343 ( .A(n6015), .B(n6014), .Z(n483) );
  NAND U2344 ( .A(n6013), .B(n6012), .Z(n484) );
  NAND U2345 ( .A(n483), .B(n484), .Z(n7638) );
  NAND U2346 ( .A(n6636), .B(n6635), .Z(n485) );
  NAND U2347 ( .A(n6633), .B(n6634), .Z(n486) );
  AND U2348 ( .A(n485), .B(n486), .Z(n7642) );
  NAND U2349 ( .A(n5905), .B(n5904), .Z(n487) );
  NAND U2350 ( .A(n5902), .B(n5903), .Z(n488) );
  AND U2351 ( .A(n487), .B(n488), .Z(n7548) );
  NAND U2352 ( .A(n6045), .B(n6044), .Z(n489) );
  NAND U2353 ( .A(n6043), .B(n6042), .Z(n490) );
  NAND U2354 ( .A(n489), .B(n490), .Z(n7554) );
  NAND U2355 ( .A(n5620), .B(n5619), .Z(n491) );
  NAND U2356 ( .A(n5618), .B(n5617), .Z(n492) );
  NAND U2357 ( .A(n491), .B(n492), .Z(n7513) );
  NAND U2358 ( .A(n5563), .B(n5562), .Z(n493) );
  NAND U2359 ( .A(n5561), .B(n5560), .Z(n494) );
  NAND U2360 ( .A(n493), .B(n494), .Z(n7518) );
  NAND U2361 ( .A(n7142), .B(n7141), .Z(n495) );
  NAND U2362 ( .A(n7139), .B(n7140), .Z(n496) );
  AND U2363 ( .A(n495), .B(n496), .Z(n8180) );
  NAND U2364 ( .A(n6716), .B(n6715), .Z(n497) );
  NAND U2365 ( .A(n6713), .B(n6714), .Z(n498) );
  AND U2366 ( .A(n497), .B(n498), .Z(n8174) );
  NAND U2367 ( .A(n4263), .B(n4262), .Z(n499) );
  NAND U2368 ( .A(n4260), .B(n4261), .Z(n500) );
  AND U2369 ( .A(n499), .B(n500), .Z(n5772) );
  NAND U2370 ( .A(n2257), .B(n2256), .Z(n501) );
  NAND U2371 ( .A(n2254), .B(n2255), .Z(n502) );
  AND U2372 ( .A(n501), .B(n502), .Z(n5766) );
  NAND U2373 ( .A(n5598), .B(n5597), .Z(n503) );
  NAND U2374 ( .A(n5595), .B(n5596), .Z(n504) );
  AND U2375 ( .A(n503), .B(n504), .Z(n8266) );
  NAND U2376 ( .A(n5640), .B(n5639), .Z(n505) );
  NAND U2377 ( .A(n5638), .B(n5637), .Z(n506) );
  NAND U2378 ( .A(n505), .B(n506), .Z(n7617) );
  NAND U2379 ( .A(n5997), .B(n5996), .Z(n507) );
  NAND U2380 ( .A(n5995), .B(n5994), .Z(n508) );
  NAND U2381 ( .A(n507), .B(n508), .Z(n7629) );
  NAND U2382 ( .A(n7332), .B(n7331), .Z(n509) );
  NAND U2383 ( .A(n7329), .B(n7330), .Z(n510) );
  AND U2384 ( .A(n509), .B(n510), .Z(n8026) );
  NAND U2385 ( .A(n5445), .B(n5444), .Z(n511) );
  NAND U2386 ( .A(n5442), .B(n5443), .Z(n512) );
  AND U2387 ( .A(n511), .B(n512), .Z(n8020) );
  NAND U2388 ( .A(n6742), .B(n6741), .Z(n513) );
  NAND U2389 ( .A(n6739), .B(n6740), .Z(n514) );
  AND U2390 ( .A(n513), .B(n514), .Z(n8034) );
  NAND U2391 ( .A(n6480), .B(n6479), .Z(n515) );
  NAND U2392 ( .A(n6477), .B(n6478), .Z(n516) );
  AND U2393 ( .A(n515), .B(n516), .Z(n8220) );
  NAND U2394 ( .A(n6330), .B(n6329), .Z(n517) );
  NAND U2395 ( .A(n6327), .B(n6328), .Z(n518) );
  AND U2396 ( .A(n517), .B(n518), .Z(n8422) );
  NAND U2397 ( .A(n6912), .B(n6911), .Z(n519) );
  NAND U2398 ( .A(n6909), .B(n6910), .Z(n520) );
  AND U2399 ( .A(n519), .B(n520), .Z(n8434) );
  NAND U2400 ( .A(n6056), .B(n6057), .Z(n521) );
  NANDN U2401 ( .A(n6059), .B(n6058), .Z(n522) );
  AND U2402 ( .A(n521), .B(n522), .Z(n8455) );
  NAND U2403 ( .A(n7371), .B(n7372), .Z(n523) );
  NANDN U2404 ( .A(n7374), .B(n7373), .Z(n524) );
  AND U2405 ( .A(n523), .B(n524), .Z(n8277) );
  NAND U2406 ( .A(n1758), .B(n1757), .Z(n525) );
  NAND U2407 ( .A(n1756), .B(n1755), .Z(n526) );
  NAND U2408 ( .A(n525), .B(n526), .Z(n7061) );
  NAND U2409 ( .A(n5587), .B(n5586), .Z(n527) );
  NAND U2410 ( .A(n5585), .B(n5584), .Z(n528) );
  NAND U2411 ( .A(n527), .B(n528), .Z(n7995) );
  XNOR U2412 ( .A(n7672), .B(n7671), .Z(n7673) );
  NAND U2413 ( .A(n5407), .B(n5406), .Z(n529) );
  NAND U2414 ( .A(n5405), .B(n5404), .Z(n530) );
  NAND U2415 ( .A(n529), .B(n530), .Z(n8014) );
  NAND U2416 ( .A(n7106), .B(n7105), .Z(n531) );
  NAND U2417 ( .A(n7104), .B(n7103), .Z(n532) );
  NAND U2418 ( .A(n531), .B(n532), .Z(n8078) );
  NAND U2419 ( .A(n5363), .B(n5362), .Z(n533) );
  NAND U2420 ( .A(n5361), .B(n5360), .Z(n534) );
  AND U2421 ( .A(n533), .B(n534), .Z(n8073) );
  NAND U2422 ( .A(n5943), .B(n5942), .Z(n535) );
  NAND U2423 ( .A(n5941), .B(n5940), .Z(n536) );
  AND U2424 ( .A(n535), .B(n536), .Z(n7581) );
  NAND U2425 ( .A(n7266), .B(n7265), .Z(n537) );
  NANDN U2426 ( .A(n7264), .B(n7263), .Z(n538) );
  AND U2427 ( .A(n537), .B(n538), .Z(n7971) );
  NAND U2428 ( .A(n6870), .B(n6869), .Z(n539) );
  NAND U2429 ( .A(n6868), .B(n6867), .Z(n540) );
  NAND U2430 ( .A(n539), .B(n540), .Z(n7538) );
  NAND U2431 ( .A(n6564), .B(n6563), .Z(n541) );
  NAND U2432 ( .A(n6562), .B(n6561), .Z(n542) );
  AND U2433 ( .A(n541), .B(n542), .Z(n7718) );
  NAND U2434 ( .A(n6626), .B(n6625), .Z(n543) );
  NAND U2435 ( .A(n6623), .B(n6624), .Z(n544) );
  AND U2436 ( .A(n543), .B(n544), .Z(n7711) );
  NAND U2437 ( .A(n6834), .B(n6833), .Z(n545) );
  NAND U2438 ( .A(n6832), .B(n6831), .Z(n546) );
  AND U2439 ( .A(n545), .B(n546), .Z(n7708) );
  NAND U2440 ( .A(n6548), .B(n6547), .Z(n547) );
  NAND U2441 ( .A(n6546), .B(n6545), .Z(n548) );
  NAND U2442 ( .A(n547), .B(n548), .Z(n7777) );
  NAND U2443 ( .A(n6598), .B(n6597), .Z(n549) );
  NAND U2444 ( .A(n6596), .B(n6595), .Z(n550) );
  AND U2445 ( .A(n549), .B(n550), .Z(n7601) );
  NAND U2446 ( .A(n7570), .B(n7569), .Z(n551) );
  NAND U2447 ( .A(n7568), .B(n7567), .Z(n552) );
  AND U2448 ( .A(n551), .B(n552), .Z(n9028) );
  NAND U2449 ( .A(n7512), .B(n7511), .Z(n553) );
  NAND U2450 ( .A(n7510), .B(n7509), .Z(n554) );
  AND U2451 ( .A(n553), .B(n554), .Z(n8961) );
  NAND U2452 ( .A(n5771), .B(n5770), .Z(n555) );
  NAND U2453 ( .A(n5769), .B(n5768), .Z(n556) );
  NAND U2454 ( .A(n555), .B(n556), .Z(n8459) );
  NAND U2455 ( .A(n8454), .B(n8453), .Z(n557) );
  NAND U2456 ( .A(n8452), .B(n8451), .Z(n558) );
  AND U2457 ( .A(n557), .B(n558), .Z(n8640) );
  NAND U2458 ( .A(n8269), .B(n8270), .Z(n559) );
  NANDN U2459 ( .A(n8272), .B(n8271), .Z(n560) );
  NAND U2460 ( .A(n559), .B(n560), .Z(n8807) );
  NAND U2461 ( .A(n7932), .B(n7931), .Z(n561) );
  NAND U2462 ( .A(n7929), .B(n7930), .Z(n562) );
  AND U2463 ( .A(n561), .B(n562), .Z(n8783) );
  NAND U2464 ( .A(n8259), .B(n8260), .Z(n563) );
  NANDN U2465 ( .A(n8262), .B(n8261), .Z(n564) );
  AND U2466 ( .A(n563), .B(n564), .Z(n8988) );
  NAND U2467 ( .A(n5217), .B(n5216), .Z(n565) );
  NANDN U2468 ( .A(n5215), .B(n5214), .Z(n566) );
  AND U2469 ( .A(n565), .B(n566), .Z(n6966) );
  XNOR U2470 ( .A(n7404), .B(n7403), .Z(n7405) );
  NAND U2471 ( .A(n4061), .B(n4060), .Z(n567) );
  NANDN U2472 ( .A(n4059), .B(n4058), .Z(n568) );
  AND U2473 ( .A(n567), .B(n568), .Z(n6607) );
  NAND U2474 ( .A(n7684), .B(n7683), .Z(n569) );
  NAND U2475 ( .A(n7682), .B(n7681), .Z(n570) );
  AND U2476 ( .A(n569), .B(n570), .Z(n8814) );
  NAND U2477 ( .A(n8086), .B(n8085), .Z(n571) );
  NAND U2478 ( .A(n8084), .B(n8083), .Z(n572) );
  NAND U2479 ( .A(n571), .B(n572), .Z(n9002) );
  NAND U2480 ( .A(n7578), .B(n7577), .Z(n573) );
  NAND U2481 ( .A(n7575), .B(n7576), .Z(n574) );
  AND U2482 ( .A(n573), .B(n574), .Z(n8590) );
  NAND U2483 ( .A(n7982), .B(n7981), .Z(n575) );
  NAND U2484 ( .A(n7980), .B(n7979), .Z(n576) );
  NAND U2485 ( .A(n575), .B(n576), .Z(n8945) );
  NAND U2486 ( .A(n8290), .B(n8289), .Z(n577) );
  NANDN U2487 ( .A(n8288), .B(n8287), .Z(n578) );
  AND U2488 ( .A(n577), .B(n578), .Z(n8705) );
  NAND U2489 ( .A(n8411), .B(n8412), .Z(n579) );
  NANDN U2490 ( .A(n8414), .B(n8413), .Z(n580) );
  NAND U2491 ( .A(n579), .B(n580), .Z(n8739) );
  NAND U2492 ( .A(n9038), .B(n9037), .Z(n581) );
  NAND U2493 ( .A(n9035), .B(n9036), .Z(n582) );
  AND U2494 ( .A(n581), .B(n582), .Z(n9187) );
  NAND U2495 ( .A(n9023), .B(n9022), .Z(n583) );
  NAND U2496 ( .A(n9021), .B(n9020), .Z(n584) );
  NAND U2497 ( .A(n583), .B(n584), .Z(n9196) );
  NAND U2498 ( .A(n8955), .B(n8954), .Z(n585) );
  NAND U2499 ( .A(n8952), .B(n8953), .Z(n586) );
  AND U2500 ( .A(n585), .B(n586), .Z(n9174) );
  NAND U2501 ( .A(n8781), .B(n8780), .Z(n587) );
  NAND U2502 ( .A(n8779), .B(n8778), .Z(n588) );
  NAND U2503 ( .A(n587), .B(n588), .Z(n9226) );
  NAND U2504 ( .A(n8663), .B(n8662), .Z(n589) );
  NAND U2505 ( .A(n8661), .B(n8660), .Z(n590) );
  AND U2506 ( .A(n589), .B(n590), .Z(n9222) );
  XNOR U2507 ( .A(n7862), .B(n7861), .Z(n7863) );
  XOR U2508 ( .A(n8983), .B(n8982), .Z(n8873) );
  XNOR U2509 ( .A(n8394), .B(n8393), .Z(n8395) );
  XNOR U2510 ( .A(n9050), .B(n9049), .Z(n9051) );
  NAND U2511 ( .A(n9012), .B(n9013), .Z(n591) );
  NANDN U2512 ( .A(n9015), .B(n9014), .Z(n592) );
  AND U2513 ( .A(n591), .B(n592), .Z(n9215) );
  NAND U2514 ( .A(n8964), .B(n8965), .Z(n593) );
  NANDN U2515 ( .A(n8967), .B(n8966), .Z(n594) );
  NAND U2516 ( .A(n593), .B(n594), .Z(n9146) );
  NAND U2517 ( .A(n8943), .B(n8942), .Z(n595) );
  NAND U2518 ( .A(n8941), .B(n8940), .Z(n596) );
  AND U2519 ( .A(n595), .B(n596), .Z(n9141) );
  NAND U2520 ( .A(n8600), .B(n8601), .Z(n597) );
  NANDN U2521 ( .A(n8603), .B(n8602), .Z(n598) );
  AND U2522 ( .A(n597), .B(n598), .Z(n9282) );
  NAND U2523 ( .A(n8935), .B(n8934), .Z(n599) );
  NAND U2524 ( .A(n8932), .B(n8933), .Z(n600) );
  AND U2525 ( .A(n599), .B(n600), .Z(n9096) );
  NAND U2526 ( .A(n8703), .B(n8702), .Z(n601) );
  NAND U2527 ( .A(n8701), .B(n8700), .Z(n602) );
  AND U2528 ( .A(n601), .B(n602), .Z(n9095) );
  NAND U2529 ( .A(n8734), .B(n8735), .Z(n603) );
  NANDN U2530 ( .A(n8737), .B(n8736), .Z(n604) );
  AND U2531 ( .A(n603), .B(n604), .Z(n9087) );
  NAND U2532 ( .A(n8750), .B(n8751), .Z(n605) );
  NANDN U2533 ( .A(n8753), .B(n8752), .Z(n606) );
  NAND U2534 ( .A(n605), .B(n606), .Z(n9136) );
  NAND U2535 ( .A(n9193), .B(n9192), .Z(n607) );
  NAND U2536 ( .A(n9191), .B(n9190), .Z(n608) );
  AND U2537 ( .A(n607), .B(n608), .Z(n9392) );
  NAND U2538 ( .A(n9178), .B(n9179), .Z(n609) );
  NANDN U2539 ( .A(n9181), .B(n9180), .Z(n610) );
  NAND U2540 ( .A(n609), .B(n610), .Z(n9386) );
  NAND U2541 ( .A(n9231), .B(n9230), .Z(n611) );
  NAND U2542 ( .A(n9229), .B(n9228), .Z(n612) );
  AND U2543 ( .A(n611), .B(n612), .Z(n9397) );
  NAND U2544 ( .A(n9239), .B(n9238), .Z(n613) );
  NAND U2545 ( .A(n9237), .B(n9236), .Z(n614) );
  NAND U2546 ( .A(n613), .B(n614), .Z(n9380) );
  XNOR U2547 ( .A(n7028), .B(n7027), .Z(n7029) );
  NAND U2548 ( .A(n7116), .B(n7115), .Z(n615) );
  NANDN U2549 ( .A(n7114), .B(n7113), .Z(n616) );
  AND U2550 ( .A(n615), .B(n616), .Z(n8401) );
  XNOR U2551 ( .A(n9131), .B(n9130), .Z(n9132) );
  XNOR U2552 ( .A(n9125), .B(n9124), .Z(n9126) );
  NAND U2553 ( .A(n9213), .B(n9212), .Z(n617) );
  NAND U2554 ( .A(n9211), .B(n9210), .Z(n618) );
  NAND U2555 ( .A(n617), .B(n618), .Z(n9410) );
  XNOR U2556 ( .A(n8511), .B(n8510), .Z(n8512) );
  XOR U2557 ( .A(n8390), .B(n8389), .Z(n7692) );
  XNOR U2558 ( .A(n9075), .B(n9074), .Z(n9077) );
  XNOR U2559 ( .A(n8529), .B(n8528), .Z(n8531) );
  XOR U2560 ( .A(n9343), .B(n9342), .Z(n9362) );
  XNOR U2561 ( .A(n9518), .B(n9517), .Z(n9519) );
  NAND U2562 ( .A(n9479), .B(n9478), .Z(n619) );
  NANDN U2563 ( .A(n9477), .B(n9476), .Z(n620) );
  AND U2564 ( .A(n619), .B(n620), .Z(n9538) );
  ANDN U2565 ( .B(n9535), .A(n9536), .Z(n9542) );
  XNOR U2566 ( .A(n9467), .B(n9466), .Z(n9468) );
  NAND U2567 ( .A(n9358), .B(n9360), .Z(n621) );
  XOR U2568 ( .A(n9358), .B(n9360), .Z(n622) );
  NANDN U2569 ( .A(n9359), .B(n622), .Z(n623) );
  NAND U2570 ( .A(n621), .B(n623), .Z(n9524) );
  NAND U2571 ( .A(n9556), .B(n9557), .Z(n624) );
  XOR U2572 ( .A(n9556), .B(n9557), .Z(n625) );
  NANDN U2573 ( .A(n9555), .B(n625), .Z(n626) );
  NAND U2574 ( .A(n624), .B(n626), .Z(n9566) );
  XNOR U2575 ( .A(n1818), .B(n1817), .Z(n1819) );
  XNOR U2576 ( .A(n5141), .B(n5140), .Z(n5142) );
  XNOR U2577 ( .A(n3557), .B(n3556), .Z(n3558) );
  NAND U2578 ( .A(n2171), .B(n2170), .Z(n627) );
  NAND U2579 ( .A(n2168), .B(n2169), .Z(n628) );
  AND U2580 ( .A(n627), .B(n628), .Z(n5719) );
  NAND U2581 ( .A(n1194), .B(n1193), .Z(n629) );
  NAND U2582 ( .A(n1191), .B(n1192), .Z(n630) );
  AND U2583 ( .A(n629), .B(n630), .Z(n6467) );
  NAND U2584 ( .A(n4087), .B(n4086), .Z(n631) );
  NAND U2585 ( .A(n4084), .B(n4085), .Z(n632) );
  AND U2586 ( .A(n631), .B(n632), .Z(n5683) );
  NAND U2587 ( .A(n1700), .B(n1699), .Z(n633) );
  NAND U2588 ( .A(n1697), .B(n1698), .Z(n634) );
  AND U2589 ( .A(n633), .B(n634), .Z(n6775) );
  NAND U2590 ( .A(n3707), .B(n3706), .Z(n635) );
  NAND U2591 ( .A(n3704), .B(n3705), .Z(n636) );
  NAND U2592 ( .A(n635), .B(n636), .Z(n6772) );
  NAND U2593 ( .A(n3763), .B(n3762), .Z(n637) );
  NAND U2594 ( .A(n3760), .B(n3761), .Z(n638) );
  NAND U2595 ( .A(n637), .B(n638), .Z(n6766) );
  NAND U2596 ( .A(n2801), .B(n2800), .Z(n639) );
  NAND U2597 ( .A(n2798), .B(n2799), .Z(n640) );
  NAND U2598 ( .A(n639), .B(n640), .Z(n7320) );
  NAND U2599 ( .A(n4767), .B(n4766), .Z(n641) );
  NAND U2600 ( .A(n4764), .B(n4765), .Z(n642) );
  AND U2601 ( .A(n641), .B(n642), .Z(n6667) );
  NAND U2602 ( .A(n3555), .B(n3554), .Z(n643) );
  NAND U2603 ( .A(n3552), .B(n3553), .Z(n644) );
  NAND U2604 ( .A(n643), .B(n644), .Z(n6664) );
  NAND U2605 ( .A(n2541), .B(n2540), .Z(n645) );
  NAND U2606 ( .A(n2538), .B(n2539), .Z(n646) );
  AND U2607 ( .A(n645), .B(n646), .Z(n6403) );
  NAND U2608 ( .A(n3525), .B(n3524), .Z(n647) );
  NAND U2609 ( .A(n3522), .B(n3523), .Z(n648) );
  NAND U2610 ( .A(n647), .B(n648), .Z(n6400) );
  NAND U2611 ( .A(n3605), .B(n3604), .Z(n649) );
  NAND U2612 ( .A(n3602), .B(n3603), .Z(n650) );
  AND U2613 ( .A(n649), .B(n650), .Z(n6002) );
  NAND U2614 ( .A(n4683), .B(n4682), .Z(n651) );
  NAND U2615 ( .A(n4680), .B(n4681), .Z(n652) );
  AND U2616 ( .A(n651), .B(n652), .Z(n6627) );
  NAND U2617 ( .A(n3001), .B(n3000), .Z(n653) );
  NAND U2618 ( .A(n2998), .B(n2999), .Z(n654) );
  AND U2619 ( .A(n653), .B(n654), .Z(n5908) );
  NAND U2620 ( .A(n2851), .B(n2850), .Z(n655) );
  NAND U2621 ( .A(n2848), .B(n2849), .Z(n656) );
  AND U2622 ( .A(n655), .B(n656), .Z(n5903) );
  NAND U2623 ( .A(n4357), .B(n4356), .Z(n657) );
  NAND U2624 ( .A(n4354), .B(n4355), .Z(n658) );
  AND U2625 ( .A(n657), .B(n658), .Z(n5623) );
  NAND U2626 ( .A(n2515), .B(n2514), .Z(n659) );
  NAND U2627 ( .A(n2512), .B(n2513), .Z(n660) );
  AND U2628 ( .A(n659), .B(n660), .Z(n6453) );
  NAND U2629 ( .A(n4009), .B(n4008), .Z(n661) );
  NAND U2630 ( .A(n4006), .B(n4007), .Z(n662) );
  AND U2631 ( .A(n661), .B(n662), .Z(n7143) );
  NAND U2632 ( .A(n5067), .B(n5066), .Z(n663) );
  NAND U2633 ( .A(n5064), .B(n5065), .Z(n664) );
  NAND U2634 ( .A(n663), .B(n664), .Z(n6718) );
  NAND U2635 ( .A(n4513), .B(n4512), .Z(n665) );
  NAND U2636 ( .A(n4510), .B(n4511), .Z(n666) );
  AND U2637 ( .A(n665), .B(n666), .Z(n6715) );
  NAND U2638 ( .A(n3585), .B(n3584), .Z(n667) );
  NAND U2639 ( .A(n3582), .B(n3583), .Z(n668) );
  AND U2640 ( .A(n667), .B(n668), .Z(n6643) );
  NAND U2641 ( .A(n4423), .B(n4422), .Z(n669) );
  NAND U2642 ( .A(n4420), .B(n4421), .Z(n670) );
  AND U2643 ( .A(n669), .B(n670), .Z(n5890) );
  NAND U2644 ( .A(n2237), .B(n2236), .Z(n671) );
  NAND U2645 ( .A(n2234), .B(n2235), .Z(n672) );
  AND U2646 ( .A(n671), .B(n672), .Z(n5756) );
  NAND U2647 ( .A(n3895), .B(n3894), .Z(n673) );
  NAND U2648 ( .A(n3892), .B(n3893), .Z(n674) );
  NAND U2649 ( .A(n673), .B(n674), .Z(n6152) );
  NAND U2650 ( .A(n3885), .B(n3884), .Z(n675) );
  NAND U2651 ( .A(n3882), .B(n3883), .Z(n676) );
  NAND U2652 ( .A(n675), .B(n676), .Z(n6148) );
  NAND U2653 ( .A(n1162), .B(n1161), .Z(n677) );
  NAND U2654 ( .A(n1159), .B(n1160), .Z(n678) );
  NAND U2655 ( .A(n677), .B(n678), .Z(n5606) );
  NAND U2656 ( .A(n4143), .B(n4142), .Z(n679) );
  NAND U2657 ( .A(n4140), .B(n4141), .Z(n680) );
  AND U2658 ( .A(n679), .B(n680), .Z(n5880) );
  NAND U2659 ( .A(n5239), .B(n5238), .Z(n681) );
  NAND U2660 ( .A(n5236), .B(n5237), .Z(n682) );
  NAND U2661 ( .A(n681), .B(n682), .Z(n5871) );
  NAND U2662 ( .A(n2003), .B(n2002), .Z(n683) );
  NAND U2663 ( .A(n2000), .B(n2001), .Z(n684) );
  AND U2664 ( .A(n683), .B(n684), .Z(n5998) );
  NAND U2665 ( .A(n4027), .B(n4026), .Z(n685) );
  NAND U2666 ( .A(n4024), .B(n4025), .Z(n686) );
  AND U2667 ( .A(n685), .B(n686), .Z(n7335) );
  NAND U2668 ( .A(n1744), .B(n1743), .Z(n687) );
  NAND U2669 ( .A(n1741), .B(n1742), .Z(n688) );
  AND U2670 ( .A(n687), .B(n688), .Z(n6747) );
  NAND U2671 ( .A(n1102), .B(n1101), .Z(n689) );
  NAND U2672 ( .A(n1099), .B(n1100), .Z(n690) );
  AND U2673 ( .A(n689), .B(n690), .Z(n6333) );
  NAND U2674 ( .A(n1614), .B(n1613), .Z(n691) );
  NAND U2675 ( .A(n1612), .B(n1611), .Z(n692) );
  NAND U2676 ( .A(n691), .B(n692), .Z(n5701) );
  NAND U2677 ( .A(n1412), .B(n1411), .Z(n693) );
  NAND U2678 ( .A(n1409), .B(n1410), .Z(n694) );
  AND U2679 ( .A(n693), .B(n694), .Z(n5733) );
  NAND U2680 ( .A(n4173), .B(n4172), .Z(n695) );
  NAND U2681 ( .A(n4170), .B(n4171), .Z(n696) );
  AND U2682 ( .A(n695), .B(n696), .Z(n5644) );
  NAND U2683 ( .A(n4131), .B(n4130), .Z(n697) );
  NAND U2684 ( .A(n4129), .B(n4128), .Z(n698) );
  NAND U2685 ( .A(n697), .B(n698), .Z(n7199) );
  NAND U2686 ( .A(n1216), .B(n1215), .Z(n699) );
  NAND U2687 ( .A(n1213), .B(n1214), .Z(n700) );
  AND U2688 ( .A(n699), .B(n700), .Z(n7388) );
  NAND U2689 ( .A(n4163), .B(n4162), .Z(n701) );
  NAND U2690 ( .A(n4161), .B(n4160), .Z(n702) );
  NAND U2691 ( .A(n701), .B(n702), .Z(n5452) );
  NAND U2692 ( .A(n2519), .B(n2518), .Z(n703) );
  NAND U2693 ( .A(n2517), .B(n2516), .Z(n704) );
  NAND U2694 ( .A(n703), .B(n704), .Z(n6123) );
  NAND U2695 ( .A(n4553), .B(n4552), .Z(n705) );
  NAND U2696 ( .A(n4550), .B(n4551), .Z(n706) );
  AND U2697 ( .A(n705), .B(n706), .Z(n7178) );
  NAND U2698 ( .A(n4679), .B(n4678), .Z(n707) );
  NAND U2699 ( .A(n4676), .B(n4677), .Z(n708) );
  AND U2700 ( .A(n707), .B(n708), .Z(n7173) );
  NAND U2701 ( .A(n4561), .B(n4560), .Z(n709) );
  NAND U2702 ( .A(n4558), .B(n4559), .Z(n710) );
  AND U2703 ( .A(n709), .B(n710), .Z(n7168) );
  NAND U2704 ( .A(n4031), .B(n4030), .Z(n711) );
  NAND U2705 ( .A(n4029), .B(n4028), .Z(n712) );
  NAND U2706 ( .A(n711), .B(n712), .Z(n5542) );
  NAND U2707 ( .A(n2597), .B(n2596), .Z(n713) );
  NAND U2708 ( .A(n2595), .B(n2594), .Z(n714) );
  NAND U2709 ( .A(n713), .B(n714), .Z(n5512) );
  NAND U2710 ( .A(n4947), .B(n4946), .Z(n715) );
  NAND U2711 ( .A(n4945), .B(n4944), .Z(n716) );
  AND U2712 ( .A(n715), .B(n716), .Z(n5539) );
  NAND U2713 ( .A(n2483), .B(n2482), .Z(n717) );
  NAND U2714 ( .A(n2481), .B(n2480), .Z(n718) );
  NAND U2715 ( .A(n717), .B(n718), .Z(n5386) );
  NAND U2716 ( .A(n2725), .B(n2724), .Z(n719) );
  NAND U2717 ( .A(n2722), .B(n2723), .Z(n720) );
  AND U2718 ( .A(n719), .B(n720), .Z(n5383) );
  NAND U2719 ( .A(n2053), .B(n2052), .Z(n721) );
  NAND U2720 ( .A(n2051), .B(n2050), .Z(n722) );
  NAND U2721 ( .A(n721), .B(n722), .Z(n6410) );
  NAND U2722 ( .A(n3429), .B(n3428), .Z(n723) );
  NAND U2723 ( .A(n3427), .B(n3426), .Z(n724) );
  NAND U2724 ( .A(n723), .B(n724), .Z(n7357) );
  NAND U2725 ( .A(n3433), .B(n3432), .Z(n725) );
  NAND U2726 ( .A(n3430), .B(n3431), .Z(n726) );
  AND U2727 ( .A(n725), .B(n726), .Z(n7348) );
  NAND U2728 ( .A(n4035), .B(n4034), .Z(n727) );
  NAND U2729 ( .A(n4032), .B(n4033), .Z(n728) );
  AND U2730 ( .A(n727), .B(n728), .Z(n5573) );
  NAND U2731 ( .A(n4827), .B(n4826), .Z(n729) );
  NAND U2732 ( .A(n4824), .B(n4825), .Z(n730) );
  AND U2733 ( .A(n729), .B(n730), .Z(n6298) );
  XNOR U2734 ( .A(n5839), .B(n5838), .Z(n5841) );
  XNOR U2735 ( .A(n5833), .B(n5832), .Z(n5835) );
  XNOR U2736 ( .A(n5863), .B(n5862), .Z(n5865) );
  XNOR U2737 ( .A(n5857), .B(n5856), .Z(n5859) );
  NAND U2738 ( .A(n4299), .B(n4298), .Z(n731) );
  NAND U2739 ( .A(n4296), .B(n4297), .Z(n732) );
  AND U2740 ( .A(n731), .B(n732), .Z(n5802) );
  XNOR U2741 ( .A(n6070), .B(n6069), .Z(n6072) );
  XNOR U2742 ( .A(n6090), .B(n6089), .Z(n6092) );
  NAND U2743 ( .A(n1909), .B(n1908), .Z(n733) );
  NAND U2744 ( .A(n1906), .B(n1907), .Z(n734) );
  NAND U2745 ( .A(n733), .B(n734), .Z(n6086) );
  XNOR U2746 ( .A(n6354), .B(n6353), .Z(n6356) );
  NAND U2747 ( .A(n3099), .B(n3098), .Z(n735) );
  NAND U2748 ( .A(n3097), .B(n3096), .Z(n736) );
  AND U2749 ( .A(n735), .B(n736), .Z(n5311) );
  NAND U2750 ( .A(n4815), .B(n4814), .Z(n737) );
  NAND U2751 ( .A(n4812), .B(n4813), .Z(n738) );
  AND U2752 ( .A(n737), .B(n738), .Z(n6902) );
  NAND U2753 ( .A(n1402), .B(n1401), .Z(n739) );
  NAND U2754 ( .A(n1400), .B(n1399), .Z(n740) );
  NAND U2755 ( .A(n739), .B(n740), .Z(n6235) );
  NAND U2756 ( .A(n2107), .B(n2106), .Z(n741) );
  NAND U2757 ( .A(n2105), .B(n2104), .Z(n742) );
  NAND U2758 ( .A(n741), .B(n742), .Z(n6311) );
  NAND U2759 ( .A(n4109), .B(n4108), .Z(n743) );
  NAND U2760 ( .A(n4106), .B(n4107), .Z(n744) );
  AND U2761 ( .A(n743), .B(n744), .Z(n5910) );
  NAND U2762 ( .A(n1917), .B(n1916), .Z(n745) );
  NAND U2763 ( .A(n1914), .B(n1915), .Z(n746) );
  AND U2764 ( .A(n745), .B(n746), .Z(n7268) );
  NAND U2765 ( .A(n2013), .B(n2012), .Z(n747) );
  NAND U2766 ( .A(n2011), .B(n2010), .Z(n748) );
  NAND U2767 ( .A(n747), .B(n748), .Z(n5982) );
  NAND U2768 ( .A(n1754), .B(n1753), .Z(n749) );
  NAND U2769 ( .A(n1752), .B(n1751), .Z(n750) );
  NAND U2770 ( .A(n749), .B(n750), .Z(n6026) );
  NAND U2771 ( .A(n1136), .B(n1135), .Z(n751) );
  NAND U2772 ( .A(n1133), .B(n1134), .Z(n752) );
  AND U2773 ( .A(n751), .B(n752), .Z(n7380) );
  NAND U2774 ( .A(n1576), .B(n1575), .Z(n753) );
  NAND U2775 ( .A(n1574), .B(n1573), .Z(n754) );
  AND U2776 ( .A(n753), .B(n754), .Z(n7005) );
  NAND U2777 ( .A(n3091), .B(n3090), .Z(n755) );
  NAND U2778 ( .A(n3089), .B(n3088), .Z(n756) );
  AND U2779 ( .A(n755), .B(n756), .Z(n6991) );
  NAND U2780 ( .A(n2748), .B(n2749), .Z(n757) );
  NANDN U2781 ( .A(n2751), .B(n2750), .Z(n758) );
  AND U2782 ( .A(n757), .B(n758), .Z(n6962) );
  NAND U2783 ( .A(n5963), .B(n5962), .Z(n759) );
  NAND U2784 ( .A(n5961), .B(n5960), .Z(n760) );
  NAND U2785 ( .A(n759), .B(n760), .Z(n7572) );
  NAND U2786 ( .A(n7314), .B(n7313), .Z(n761) );
  NAND U2787 ( .A(n7311), .B(n7312), .Z(n762) );
  AND U2788 ( .A(n761), .B(n762), .Z(n7490) );
  NAND U2789 ( .A(n7294), .B(n7293), .Z(n763) );
  NAND U2790 ( .A(n7291), .B(n7292), .Z(n764) );
  AND U2791 ( .A(n763), .B(n764), .Z(n7484) );
  NAND U2792 ( .A(n6660), .B(n6659), .Z(n765) );
  NAND U2793 ( .A(n6657), .B(n6658), .Z(n766) );
  AND U2794 ( .A(n765), .B(n766), .Z(n7464) );
  NAND U2795 ( .A(n6396), .B(n6395), .Z(n767) );
  NAND U2796 ( .A(n6393), .B(n6394), .Z(n768) );
  AND U2797 ( .A(n767), .B(n768), .Z(n8244) );
  NAND U2798 ( .A(n6011), .B(n6010), .Z(n769) );
  NAND U2799 ( .A(n6009), .B(n6008), .Z(n770) );
  NAND U2800 ( .A(n769), .B(n770), .Z(n7637) );
  NAND U2801 ( .A(n5901), .B(n5900), .Z(n771) );
  NAND U2802 ( .A(n5898), .B(n5899), .Z(n772) );
  AND U2803 ( .A(n771), .B(n772), .Z(n7550) );
  NAND U2804 ( .A(n6035), .B(n6034), .Z(n773) );
  NAND U2805 ( .A(n6033), .B(n6032), .Z(n774) );
  NAND U2806 ( .A(n773), .B(n774), .Z(n7555) );
  NAND U2807 ( .A(n6450), .B(n6449), .Z(n775) );
  NAND U2808 ( .A(n6448), .B(n6447), .Z(n776) );
  NAND U2809 ( .A(n775), .B(n776), .Z(n7509) );
  NAND U2810 ( .A(n7138), .B(n7137), .Z(n777) );
  NAND U2811 ( .A(n7135), .B(n7136), .Z(n778) );
  AND U2812 ( .A(n777), .B(n778), .Z(n8182) );
  NAND U2813 ( .A(n6656), .B(n6655), .Z(n779) );
  NAND U2814 ( .A(n6654), .B(n6653), .Z(n780) );
  NAND U2815 ( .A(n779), .B(n780), .Z(n7589) );
  NAND U2816 ( .A(n5887), .B(n5886), .Z(n781) );
  NAND U2817 ( .A(n5884), .B(n5885), .Z(n782) );
  AND U2818 ( .A(n781), .B(n782), .Z(n7598) );
  NAND U2819 ( .A(n4267), .B(n4266), .Z(n783) );
  NAND U2820 ( .A(n4264), .B(n4265), .Z(n784) );
  AND U2821 ( .A(n783), .B(n784), .Z(n5774) );
  NAND U2822 ( .A(n5753), .B(n5752), .Z(n785) );
  NAND U2823 ( .A(n5751), .B(n5750), .Z(n786) );
  NAND U2824 ( .A(n785), .B(n786), .Z(n8451) );
  NAND U2825 ( .A(n5877), .B(n5876), .Z(n787) );
  NAND U2826 ( .A(n5875), .B(n5874), .Z(n788) );
  AND U2827 ( .A(n787), .B(n788), .Z(n7624) );
  NAND U2828 ( .A(n7328), .B(n7327), .Z(n789) );
  NAND U2829 ( .A(n7325), .B(n7326), .Z(n790) );
  AND U2830 ( .A(n789), .B(n790), .Z(n8028) );
  NAND U2831 ( .A(n5441), .B(n5440), .Z(n791) );
  NAND U2832 ( .A(n5438), .B(n5439), .Z(n792) );
  AND U2833 ( .A(n791), .B(n792), .Z(n8022) );
  NAND U2834 ( .A(n6476), .B(n6475), .Z(n793) );
  NAND U2835 ( .A(n6473), .B(n6474), .Z(n794) );
  AND U2836 ( .A(n793), .B(n794), .Z(n8222) );
  NAND U2837 ( .A(n6326), .B(n6325), .Z(n795) );
  NAND U2838 ( .A(n6323), .B(n6324), .Z(n796) );
  AND U2839 ( .A(n795), .B(n796), .Z(n8424) );
  NAND U2840 ( .A(n5353), .B(n5352), .Z(n797) );
  NAND U2841 ( .A(n5351), .B(n5350), .Z(n798) );
  AND U2842 ( .A(n797), .B(n798), .Z(n8051) );
  NAND U2843 ( .A(n7424), .B(n7423), .Z(n799) );
  NAND U2844 ( .A(n7422), .B(n7421), .Z(n800) );
  AND U2845 ( .A(n799), .B(n800), .Z(n8043) );
  NAND U2846 ( .A(n7086), .B(n7085), .Z(n801) );
  NAND U2847 ( .A(n7084), .B(n7083), .Z(n802) );
  AND U2848 ( .A(n801), .B(n802), .Z(n8039) );
  NAND U2849 ( .A(n7378), .B(n7377), .Z(n803) );
  NANDN U2850 ( .A(n7376), .B(n7375), .Z(n804) );
  AND U2851 ( .A(n803), .B(n804), .Z(n8279) );
  NAND U2852 ( .A(n1550), .B(n1549), .Z(n805) );
  NAND U2853 ( .A(n1548), .B(n1547), .Z(n806) );
  AND U2854 ( .A(n805), .B(n806), .Z(n6953) );
  NAND U2855 ( .A(n4062), .B(n4063), .Z(n807) );
  NANDN U2856 ( .A(n4065), .B(n4064), .Z(n808) );
  AND U2857 ( .A(n807), .B(n808), .Z(n6605) );
  NAND U2858 ( .A(n5189), .B(n5188), .Z(n809) );
  NAND U2859 ( .A(n5186), .B(n5187), .Z(n810) );
  AND U2860 ( .A(n809), .B(n810), .Z(n6971) );
  XNOR U2861 ( .A(n7996), .B(n7995), .Z(n7997) );
  NAND U2862 ( .A(n6078), .B(n6077), .Z(n811) );
  NAND U2863 ( .A(n6076), .B(n6075), .Z(n812) );
  NAND U2864 ( .A(n811), .B(n812), .Z(n7678) );
  XNOR U2865 ( .A(n8438), .B(n8437), .Z(n8439) );
  NAND U2866 ( .A(n6340), .B(n6339), .Z(n813) );
  NAND U2867 ( .A(n6338), .B(n6337), .Z(n814) );
  AND U2868 ( .A(n813), .B(n814), .Z(n8084) );
  NAND U2869 ( .A(n7098), .B(n7097), .Z(n815) );
  NAND U2870 ( .A(n7096), .B(n7095), .Z(n816) );
  AND U2871 ( .A(n815), .B(n816), .Z(n8079) );
  NAND U2872 ( .A(n6095), .B(n6096), .Z(n817) );
  NANDN U2873 ( .A(n6098), .B(n6097), .Z(n818) );
  AND U2874 ( .A(n817), .B(n818), .Z(n7892) );
  NAND U2875 ( .A(n7366), .B(n7365), .Z(n819) );
  NAND U2876 ( .A(n7364), .B(n7363), .Z(n820) );
  NAND U2877 ( .A(n819), .B(n820), .Z(n8093) );
  NAND U2878 ( .A(n6019), .B(n6018), .Z(n821) );
  NAND U2879 ( .A(n6016), .B(n6017), .Z(n822) );
  AND U2880 ( .A(n821), .B(n822), .Z(n7990) );
  NAND U2881 ( .A(n6790), .B(n6789), .Z(n823) );
  NAND U2882 ( .A(n6787), .B(n6788), .Z(n824) );
  AND U2883 ( .A(n823), .B(n824), .Z(n7736) );
  NAND U2884 ( .A(n6732), .B(n6731), .Z(n825) );
  NAND U2885 ( .A(n6729), .B(n6730), .Z(n826) );
  AND U2886 ( .A(n825), .B(n826), .Z(n7730) );
  NAND U2887 ( .A(n6304), .B(n6303), .Z(n827) );
  NAND U2888 ( .A(n6301), .B(n6302), .Z(n828) );
  AND U2889 ( .A(n827), .B(n828), .Z(n7724) );
  NAND U2890 ( .A(n5341), .B(n5340), .Z(n829) );
  NAND U2891 ( .A(n5339), .B(n5338), .Z(n830) );
  AND U2892 ( .A(n829), .B(n830), .Z(n8472) );
  NAND U2893 ( .A(n6520), .B(n6519), .Z(n831) );
  NAND U2894 ( .A(n6518), .B(n6517), .Z(n832) );
  NAND U2895 ( .A(n831), .B(n832), .Z(n8087) );
  NAND U2896 ( .A(n6381), .B(n6382), .Z(n833) );
  NANDN U2897 ( .A(n6384), .B(n6383), .Z(n834) );
  AND U2898 ( .A(n833), .B(n834), .Z(n8067) );
  NAND U2899 ( .A(n6895), .B(n6896), .Z(n835) );
  NANDN U2900 ( .A(n6898), .B(n6897), .Z(n836) );
  AND U2901 ( .A(n835), .B(n836), .Z(n7773) );
  XNOR U2902 ( .A(n7602), .B(n7601), .Z(n7603) );
  NAND U2903 ( .A(n8250), .B(n8249), .Z(n837) );
  NAND U2904 ( .A(n8248), .B(n8247), .Z(n838) );
  NAND U2905 ( .A(n837), .B(n838), .Z(n8583) );
  NAND U2906 ( .A(n7517), .B(n7518), .Z(n839) );
  NANDN U2907 ( .A(n7520), .B(n7519), .Z(n840) );
  AND U2908 ( .A(n839), .B(n840), .Z(n8962) );
  NAND U2909 ( .A(n8185), .B(n8186), .Z(n841) );
  NANDN U2910 ( .A(n8188), .B(n8187), .Z(n842) );
  AND U2911 ( .A(n841), .B(n842), .Z(n8956) );
  NAND U2912 ( .A(n5767), .B(n5766), .Z(n843) );
  NAND U2913 ( .A(n5765), .B(n5764), .Z(n844) );
  NAND U2914 ( .A(n843), .B(n844), .Z(n8461) );
  AND U2915 ( .A(n8449), .B(n8450), .Z(n8641) );
  NAND U2916 ( .A(n8273), .B(n8274), .Z(n845) );
  NANDN U2917 ( .A(n8276), .B(n8275), .Z(n846) );
  AND U2918 ( .A(n845), .B(n846), .Z(n8808) );
  NAND U2919 ( .A(n8455), .B(n8456), .Z(n847) );
  NANDN U2920 ( .A(n8458), .B(n8457), .Z(n848) );
  NAND U2921 ( .A(n847), .B(n848), .Z(n8643) );
  NAND U2922 ( .A(n8058), .B(n8057), .Z(n849) );
  NAND U2923 ( .A(n8055), .B(n8056), .Z(n850) );
  AND U2924 ( .A(n849), .B(n850), .Z(n8790) );
  NAND U2925 ( .A(n7928), .B(n7927), .Z(n851) );
  NAND U2926 ( .A(n7925), .B(n7926), .Z(n852) );
  AND U2927 ( .A(n851), .B(n852), .Z(n8784) );
  NAND U2928 ( .A(n7912), .B(n7911), .Z(n853) );
  NAND U2929 ( .A(n7910), .B(n7909), .Z(n854) );
  NAND U2930 ( .A(n853), .B(n854), .Z(n8778) );
  NAND U2931 ( .A(n7826), .B(n7825), .Z(n855) );
  NAND U2932 ( .A(n7824), .B(n7823), .Z(n856) );
  NAND U2933 ( .A(n855), .B(n856), .Z(n8658) );
  NAND U2934 ( .A(n8132), .B(n8131), .Z(n857) );
  NAND U2935 ( .A(n8130), .B(n8129), .Z(n858) );
  NAND U2936 ( .A(n857), .B(n858), .Z(n8662) );
  NAND U2937 ( .A(n8320), .B(n8319), .Z(n859) );
  NAND U2938 ( .A(n8317), .B(n8318), .Z(n860) );
  AND U2939 ( .A(n859), .B(n860), .Z(n8567) );
  NAND U2940 ( .A(n8479), .B(n8478), .Z(n861) );
  NAND U2941 ( .A(n8477), .B(n8476), .Z(n862) );
  AND U2942 ( .A(n861), .B(n862), .Z(n8625) );
  NAND U2943 ( .A(n8102), .B(n8101), .Z(n863) );
  NAND U2944 ( .A(n8099), .B(n8100), .Z(n864) );
  AND U2945 ( .A(n863), .B(n864), .Z(n8619) );
  XNOR U2946 ( .A(n6600), .B(n6599), .Z(n6601) );
  NAND U2947 ( .A(n6132), .B(n6131), .Z(n865) );
  NAND U2948 ( .A(n6130), .B(n6129), .Z(n866) );
  AND U2949 ( .A(n865), .B(n866), .Z(n8118) );
  XNOR U2950 ( .A(n8827), .B(n8826), .Z(n9018) );
  NAND U2951 ( .A(n8294), .B(n8293), .Z(n867) );
  NAND U2952 ( .A(n8292), .B(n8291), .Z(n868) );
  NAND U2953 ( .A(n867), .B(n868), .Z(n9014) );
  NAND U2954 ( .A(n7964), .B(n7963), .Z(n869) );
  NAND U2955 ( .A(n7961), .B(n7962), .Z(n870) );
  AND U2956 ( .A(n869), .B(n870), .Z(n8831) );
  NAND U2957 ( .A(n8076), .B(n8075), .Z(n871) );
  NAND U2958 ( .A(n8073), .B(n8074), .Z(n872) );
  AND U2959 ( .A(n871), .B(n872), .Z(n9005) );
  NAND U2960 ( .A(n7972), .B(n7971), .Z(n873) );
  NAND U2961 ( .A(n7970), .B(n7969), .Z(n874) );
  NAND U2962 ( .A(n873), .B(n874), .Z(n8946) );
  NAND U2963 ( .A(n8154), .B(n8153), .Z(n875) );
  NAND U2964 ( .A(n8152), .B(n8151), .Z(n876) );
  NAND U2965 ( .A(n875), .B(n876), .Z(n8940) );
  NAND U2966 ( .A(n7701), .B(n7702), .Z(n877) );
  NANDN U2967 ( .A(n7704), .B(n7703), .Z(n878) );
  AND U2968 ( .A(n877), .B(n878), .Z(n8724) );
  NAND U2969 ( .A(n7780), .B(n7779), .Z(n879) );
  NAND U2970 ( .A(n7778), .B(n7777), .Z(n880) );
  AND U2971 ( .A(n879), .B(n880), .Z(n8884) );
  NAND U2972 ( .A(n9042), .B(n9041), .Z(n881) );
  NAND U2973 ( .A(n9039), .B(n9040), .Z(n882) );
  AND U2974 ( .A(n881), .B(n882), .Z(n9186) );
  XNOR U2975 ( .A(n7406), .B(n7405), .Z(n6819) );
  XNOR U2976 ( .A(n8917), .B(n8916), .Z(n8918) );
  XNOR U2977 ( .A(n8683), .B(n8682), .Z(n8685) );
  NAND U2978 ( .A(n8951), .B(n8950), .Z(n883) );
  NAND U2979 ( .A(n8949), .B(n8948), .Z(n884) );
  AND U2980 ( .A(n883), .B(n884), .Z(n9148) );
  NAND U2981 ( .A(n8939), .B(n8938), .Z(n885) );
  NAND U2982 ( .A(n8937), .B(n8936), .Z(n886) );
  AND U2983 ( .A(n885), .B(n886), .Z(n9142) );
  NAND U2984 ( .A(n8928), .B(n8929), .Z(n887) );
  NANDN U2985 ( .A(n8931), .B(n8930), .Z(n888) );
  AND U2986 ( .A(n887), .B(n888), .Z(n9097) );
  NAND U2987 ( .A(n8845), .B(n8844), .Z(n889) );
  NAND U2988 ( .A(n8842), .B(n8843), .Z(n890) );
  AND U2989 ( .A(n889), .B(n890), .Z(n9112) );
  NAND U2990 ( .A(n8891), .B(n8890), .Z(n891) );
  NAND U2991 ( .A(n8888), .B(n8889), .Z(n892) );
  AND U2992 ( .A(n891), .B(n892), .Z(n9247) );
  NAND U2993 ( .A(n9197), .B(n9196), .Z(n893) );
  NAND U2994 ( .A(n9195), .B(n9194), .Z(n894) );
  AND U2995 ( .A(n893), .B(n894), .Z(n9391) );
  NAND U2996 ( .A(n9235), .B(n9234), .Z(n895) );
  NAND U2997 ( .A(n9232), .B(n9233), .Z(n896) );
  AND U2998 ( .A(n895), .B(n896), .Z(n9379) );
  XNOR U2999 ( .A(n6268), .B(n6267), .Z(n7437) );
  XNOR U3000 ( .A(n8388), .B(n8387), .Z(n8389) );
  XOR U3001 ( .A(n7864), .B(n7863), .Z(n7686) );
  XNOR U3002 ( .A(n8400), .B(n8399), .Z(n8402) );
  XOR U3003 ( .A(n8396), .B(n8395), .Z(n7800) );
  XNOR U3004 ( .A(n9295), .B(n9294), .Z(n9296) );
  NAND U3005 ( .A(n9155), .B(n9154), .Z(n897) );
  NAND U3006 ( .A(n9152), .B(n9153), .Z(n898) );
  AND U3007 ( .A(n897), .B(n898), .Z(n9417) );
  NAND U3008 ( .A(n9095), .B(n9094), .Z(n899) );
  NAND U3009 ( .A(n9092), .B(n9093), .Z(n900) );
  AND U3010 ( .A(n899), .B(n900), .Z(n9400) );
  NAND U3011 ( .A(n9108), .B(n9109), .Z(n901) );
  NANDN U3012 ( .A(n9111), .B(n9110), .Z(n902) );
  AND U3013 ( .A(n901), .B(n902), .Z(n9449) );
  NAND U3014 ( .A(n9136), .B(n9137), .Z(n903) );
  NANDN U3015 ( .A(n9139), .B(n9138), .Z(n904) );
  AND U3016 ( .A(n903), .B(n904), .Z(n9431) );
  OR U3017 ( .A(n9387), .B(n9388), .Z(n905) );
  NAND U3018 ( .A(n9386), .B(n9385), .Z(n906) );
  NAND U3019 ( .A(n905), .B(n906), .Z(n9495) );
  NAND U3020 ( .A(n9398), .B(n9397), .Z(n907) );
  NAND U3021 ( .A(n9396), .B(n9395), .Z(n908) );
  NAND U3022 ( .A(n907), .B(n908), .Z(n9486) );
  XOR U3023 ( .A(n7030), .B(n7029), .Z(n7024) );
  XOR U3024 ( .A(n9133), .B(n9132), .Z(n9315) );
  NAND U3025 ( .A(n9409), .B(n9410), .Z(n909) );
  NANDN U3026 ( .A(n9412), .B(n9411), .Z(n910) );
  NAND U3027 ( .A(n909), .B(n910), .Z(n9480) );
  NAND U3028 ( .A(n9408), .B(n9407), .Z(n911) );
  NAND U3029 ( .A(n9405), .B(n9406), .Z(n912) );
  NAND U3030 ( .A(n911), .B(n912), .Z(n9504) );
  XNOR U3031 ( .A(n9303), .B(n9302), .Z(n9321) );
  XOR U3032 ( .A(n9349), .B(n9348), .Z(n9363) );
  XOR U3033 ( .A(n9549), .B(n9548), .Z(n9551) );
  XNOR U3034 ( .A(n8378), .B(n8377), .Z(n7451) );
  XNOR U3035 ( .A(n9065), .B(n9064), .Z(n9308) );
  NAND U3036 ( .A(n9523), .B(n9525), .Z(n913) );
  XOR U3037 ( .A(n9523), .B(n9525), .Z(n914) );
  NAND U3038 ( .A(n914), .B(n9524), .Z(n915) );
  NAND U3039 ( .A(n913), .B(n915), .Z(n9545) );
  NAND U3040 ( .A(n9564), .B(n9565), .Z(n916) );
  NANDN U3041 ( .A(n9567), .B(n9566), .Z(n917) );
  NAND U3042 ( .A(n916), .B(n917), .Z(o[10]) );
  XOR U3043 ( .A(x[1139]), .B(y[1139]), .Z(n3734) );
  XOR U3044 ( .A(x[79]), .B(y[79]), .Z(n3732) );
  XNOR U3045 ( .A(x[1141]), .B(y[1141]), .Z(n3733) );
  XOR U3046 ( .A(n3732), .B(n3733), .Z(n3735) );
  XNOR U3047 ( .A(n3734), .B(n3735), .Z(n1628) );
  XOR U3048 ( .A(x[1143]), .B(y[1143]), .Z(n3703) );
  XOR U3049 ( .A(x[1145]), .B(y[1145]), .Z(n3701) );
  XOR U3050 ( .A(x[1546]), .B(y[1546]), .Z(n3700) );
  XOR U3051 ( .A(n3701), .B(n3700), .Z(n3702) );
  XOR U3052 ( .A(n3703), .B(n3702), .Z(n1627) );
  XOR U3053 ( .A(n1628), .B(n1627), .Z(n1629) );
  XOR U3054 ( .A(x[1147]), .B(y[1147]), .Z(n3638) );
  XOR U3055 ( .A(x[286]), .B(y[286]), .Z(n3636) );
  XNOR U3056 ( .A(x[1149]), .B(y[1149]), .Z(n3637) );
  XOR U3057 ( .A(n3636), .B(n3637), .Z(n3639) );
  XOR U3058 ( .A(n3638), .B(n3639), .Z(n1630) );
  XOR U3059 ( .A(n1629), .B(n1630), .Z(n3090) );
  XOR U3060 ( .A(x[1159]), .B(y[1159]), .Z(n956) );
  XOR U3061 ( .A(x[91]), .B(y[91]), .Z(n954) );
  XNOR U3062 ( .A(x[1161]), .B(y[1161]), .Z(n955) );
  XOR U3063 ( .A(n954), .B(n955), .Z(n957) );
  XNOR U3064 ( .A(n956), .B(n957), .Z(n2082) );
  XOR U3065 ( .A(x[1151]), .B(y[1151]), .Z(n3614) );
  XOR U3066 ( .A(x[85]), .B(y[85]), .Z(n3612) );
  XNOR U3067 ( .A(x[1153]), .B(y[1153]), .Z(n3613) );
  XOR U3068 ( .A(n3612), .B(n3613), .Z(n3615) );
  XNOR U3069 ( .A(n3614), .B(n3615), .Z(n2080) );
  XOR U3070 ( .A(x[1155]), .B(y[1155]), .Z(n3608) );
  XOR U3071 ( .A(x[280]), .B(y[280]), .Z(n3606) );
  XNOR U3072 ( .A(x[1157]), .B(y[1157]), .Z(n3607) );
  XOR U3073 ( .A(n3606), .B(n3607), .Z(n3609) );
  XOR U3074 ( .A(n3608), .B(n3609), .Z(n2081) );
  XOR U3075 ( .A(n2080), .B(n2081), .Z(n2083) );
  XOR U3076 ( .A(n2082), .B(n2083), .Z(n3088) );
  XOR U3077 ( .A(x[1163]), .B(y[1163]), .Z(n1307) );
  XOR U3078 ( .A(x[95]), .B(y[95]), .Z(n1305) );
  XNOR U3079 ( .A(x[1165]), .B(y[1165]), .Z(n1306) );
  XOR U3080 ( .A(n1305), .B(n1306), .Z(n1308) );
  XNOR U3081 ( .A(n1307), .B(n1308), .Z(n2353) );
  XOR U3082 ( .A(x[1167]), .B(y[1167]), .Z(n1047) );
  XOR U3083 ( .A(x[1169]), .B(y[1169]), .Z(n1044) );
  XNOR U3084 ( .A(x[1548]), .B(y[1548]), .Z(n1045) );
  XNOR U3085 ( .A(n1044), .B(n1045), .Z(n1046) );
  XOR U3086 ( .A(n1047), .B(n1046), .Z(n2352) );
  XOR U3087 ( .A(n2353), .B(n2352), .Z(n2355) );
  XOR U3088 ( .A(x[1171]), .B(y[1171]), .Z(n1040) );
  XOR U3089 ( .A(x[101]), .B(y[101]), .Z(n1038) );
  XNOR U3090 ( .A(x[1173]), .B(y[1173]), .Z(n1039) );
  XOR U3091 ( .A(n1038), .B(n1039), .Z(n1041) );
  XNOR U3092 ( .A(n1040), .B(n1041), .Z(n2354) );
  XNOR U3093 ( .A(n2355), .B(n2354), .Z(n3089) );
  XOR U3094 ( .A(n3088), .B(n3089), .Z(n3091) );
  XOR U3095 ( .A(n3090), .B(n3091), .Z(n1124) );
  XOR U3096 ( .A(x[1319]), .B(y[1319]), .Z(n1642) );
  XOR U3097 ( .A(x[201]), .B(y[201]), .Z(n1640) );
  XOR U3098 ( .A(x[1321]), .B(y[1321]), .Z(n1639) );
  XOR U3099 ( .A(n1640), .B(n1639), .Z(n1641) );
  XOR U3100 ( .A(n1642), .B(n1641), .Z(n1172) );
  XOR U3101 ( .A(x[1315]), .B(y[1315]), .Z(n4933) );
  XOR U3102 ( .A(x[180]), .B(y[180]), .Z(n4931) );
  XOR U3103 ( .A(x[1317]), .B(y[1317]), .Z(n4930) );
  XOR U3104 ( .A(n4931), .B(n4930), .Z(n4932) );
  XOR U3105 ( .A(n4933), .B(n4932), .Z(n1170) );
  XOR U3106 ( .A(x[1427]), .B(y[1427]), .Z(n4767) );
  XOR U3107 ( .A(x[277]), .B(y[277]), .Z(n4765) );
  XOR U3108 ( .A(x[1429]), .B(y[1429]), .Z(n4764) );
  XOR U3109 ( .A(n4765), .B(n4764), .Z(n4766) );
  XOR U3110 ( .A(n4767), .B(n4766), .Z(n1169) );
  XOR U3111 ( .A(n1170), .B(n1169), .Z(n1171) );
  XOR U3112 ( .A(n1172), .B(n1171), .Z(n5131) );
  XOR U3113 ( .A(x[1323]), .B(y[1323]), .Z(n4911) );
  XOR U3114 ( .A(x[205]), .B(y[205]), .Z(n4909) );
  XOR U3115 ( .A(x[1325]), .B(y[1325]), .Z(n4908) );
  XOR U3116 ( .A(n4909), .B(n4908), .Z(n4910) );
  XOR U3117 ( .A(n4911), .B(n4910), .Z(n4803) );
  XOR U3118 ( .A(x[1423]), .B(y[1423]), .Z(n4783) );
  XOR U3119 ( .A(x[1425]), .B(y[1425]), .Z(n4781) );
  XOR U3120 ( .A(x[1580]), .B(y[1580]), .Z(n4780) );
  XOR U3121 ( .A(n4781), .B(n4780), .Z(n4782) );
  XOR U3122 ( .A(n4783), .B(n4782), .Z(n4802) );
  XOR U3123 ( .A(n4803), .B(n4802), .Z(n4805) );
  XOR U3124 ( .A(x[1419]), .B(y[1419]), .Z(n5031) );
  XOR U3125 ( .A(x[271]), .B(y[271]), .Z(n5029) );
  XOR U3126 ( .A(x[1421]), .B(y[1421]), .Z(n5028) );
  XOR U3127 ( .A(n5029), .B(n5028), .Z(n5030) );
  XOR U3128 ( .A(n5031), .B(n5030), .Z(n4804) );
  XOR U3129 ( .A(n4805), .B(n4804), .Z(n5129) );
  XOR U3130 ( .A(x[1327]), .B(y[1327]), .Z(n4135) );
  XOR U3131 ( .A(x[1329]), .B(y[1329]), .Z(n4133) );
  XOR U3132 ( .A(x[1568]), .B(y[1568]), .Z(n4132) );
  XOR U3133 ( .A(n4133), .B(n4132), .Z(n4134) );
  XOR U3134 ( .A(n4135), .B(n4134), .Z(n2517) );
  XOR U3135 ( .A(x[1363]), .B(y[1363]), .Z(n1897) );
  XOR U3136 ( .A(x[233]), .B(y[233]), .Z(n1895) );
  XOR U3137 ( .A(x[1365]), .B(y[1365]), .Z(n1894) );
  XOR U3138 ( .A(n1895), .B(n1894), .Z(n1896) );
  XOR U3139 ( .A(n1897), .B(n1896), .Z(n2516) );
  XOR U3140 ( .A(n2517), .B(n2516), .Z(n2519) );
  XOR U3141 ( .A(x[1331]), .B(y[1331]), .Z(n4147) );
  XOR U3142 ( .A(x[211]), .B(y[211]), .Z(n4145) );
  XOR U3143 ( .A(x[1333]), .B(y[1333]), .Z(n4144) );
  XOR U3144 ( .A(n4145), .B(n4144), .Z(n4146) );
  XOR U3145 ( .A(n4147), .B(n4146), .Z(n2518) );
  XNOR U3146 ( .A(n2519), .B(n2518), .Z(n5128) );
  XNOR U3147 ( .A(n5129), .B(n5128), .Z(n5130) );
  XNOR U3148 ( .A(n5131), .B(n5130), .Z(n1121) );
  XOR U3149 ( .A(x[1103]), .B(y[1103]), .Z(n2882) );
  XOR U3150 ( .A(x[1105]), .B(y[1105]), .Z(n2880) );
  XNOR U3151 ( .A(x[1540]), .B(y[1540]), .Z(n2881) );
  XOR U3152 ( .A(n2880), .B(n2881), .Z(n2883) );
  XNOR U3153 ( .A(n2882), .B(n2883), .Z(n1558) );
  XOR U3154 ( .A(x[1107]), .B(y[1107]), .Z(n2515) );
  XOR U3155 ( .A(x[57]), .B(y[57]), .Z(n2513) );
  XOR U3156 ( .A(x[1109]), .B(y[1109]), .Z(n2512) );
  XOR U3157 ( .A(n2513), .B(n2512), .Z(n2514) );
  XOR U3158 ( .A(n2515), .B(n2514), .Z(n1557) );
  XOR U3159 ( .A(n1558), .B(n1557), .Z(n1560) );
  XOR U3160 ( .A(x[1111]), .B(y[1111]), .Z(n4771) );
  XOR U3161 ( .A(x[1113]), .B(y[1113]), .Z(n4769) );
  XOR U3162 ( .A(x[1542]), .B(y[1542]), .Z(n4768) );
  XOR U3163 ( .A(n4769), .B(n4768), .Z(n4770) );
  XOR U3164 ( .A(n4771), .B(n4770), .Z(n1559) );
  XOR U3165 ( .A(n1560), .B(n1559), .Z(n2751) );
  XOR U3166 ( .A(x[1115]), .B(y[1115]), .Z(n4050) );
  XOR U3167 ( .A(x[306]), .B(y[306]), .Z(n4048) );
  XNOR U3168 ( .A(x[1117]), .B(y[1117]), .Z(n4049) );
  XOR U3169 ( .A(n4048), .B(n4049), .Z(n4051) );
  XNOR U3170 ( .A(n4050), .B(n4051), .Z(n5174) );
  XOR U3171 ( .A(x[1119]), .B(y[1119]), .Z(n4044) );
  XOR U3172 ( .A(x[63]), .B(y[63]), .Z(n4042) );
  XNOR U3173 ( .A(x[1121]), .B(y[1121]), .Z(n4043) );
  XOR U3174 ( .A(n4042), .B(n4043), .Z(n4045) );
  XOR U3175 ( .A(n4044), .B(n4045), .Z(n5175) );
  XNOR U3176 ( .A(n5174), .B(n5175), .Z(n5176) );
  XOR U3177 ( .A(x[1123]), .B(y[1123]), .Z(n3814) );
  XOR U3178 ( .A(x[300]), .B(y[300]), .Z(n3812) );
  XNOR U3179 ( .A(x[1125]), .B(y[1125]), .Z(n3813) );
  XOR U3180 ( .A(n3812), .B(n3813), .Z(n3815) );
  XOR U3181 ( .A(n3814), .B(n3815), .Z(n5177) );
  XOR U3182 ( .A(n5176), .B(n5177), .Z(n2748) );
  XOR U3183 ( .A(x[1127]), .B(y[1127]), .Z(n3885) );
  XOR U3184 ( .A(x[69]), .B(y[69]), .Z(n3883) );
  XOR U3185 ( .A(x[1129]), .B(y[1129]), .Z(n3882) );
  XOR U3186 ( .A(n3883), .B(n3882), .Z(n3884) );
  XOR U3187 ( .A(n3885), .B(n3884), .Z(n2258) );
  XOR U3188 ( .A(x[1131]), .B(y[1131]), .Z(n3790) );
  XOR U3189 ( .A(x[73]), .B(y[73]), .Z(n3788) );
  XNOR U3190 ( .A(x[1133]), .B(y[1133]), .Z(n3789) );
  XOR U3191 ( .A(n3788), .B(n3789), .Z(n3791) );
  XOR U3192 ( .A(n3790), .B(n3791), .Z(n2259) );
  XNOR U3193 ( .A(n2258), .B(n2259), .Z(n2261) );
  XOR U3194 ( .A(x[1135]), .B(y[1135]), .Z(n3759) );
  XOR U3195 ( .A(x[1137]), .B(y[1137]), .Z(n3757) );
  XOR U3196 ( .A(x[1544]), .B(y[1544]), .Z(n3756) );
  XOR U3197 ( .A(n3757), .B(n3756), .Z(n3758) );
  XOR U3198 ( .A(n3759), .B(n3758), .Z(n2260) );
  XNOR U3199 ( .A(n2261), .B(n2260), .Z(n2749) );
  XOR U3200 ( .A(n2748), .B(n2749), .Z(n2750) );
  XOR U3201 ( .A(n2751), .B(n2750), .Z(n1122) );
  XNOR U3202 ( .A(n1121), .B(n1122), .Z(n1123) );
  XOR U3203 ( .A(n1124), .B(n1123), .Z(n5210) );
  XOR U3204 ( .A(x[1267]), .B(y[1267]), .Z(n5063) );
  XOR U3205 ( .A(x[167]), .B(y[167]), .Z(n5061) );
  XOR U3206 ( .A(x[1269]), .B(y[1269]), .Z(n5060) );
  XOR U3207 ( .A(n5061), .B(n5060), .Z(n5062) );
  XOR U3208 ( .A(n5063), .B(n5062), .Z(n4945) );
  XOR U3209 ( .A(x[1451]), .B(y[1451]), .Z(n3911) );
  XOR U3210 ( .A(x[293]), .B(y[293]), .Z(n3909) );
  XOR U3211 ( .A(x[1453]), .B(y[1453]), .Z(n3908) );
  XOR U3212 ( .A(n3909), .B(n3908), .Z(n3910) );
  XOR U3213 ( .A(n3911), .B(n3910), .Z(n4944) );
  XOR U3214 ( .A(n4945), .B(n4944), .Z(n4947) );
  XOR U3215 ( .A(x[1271]), .B(y[1271]), .Z(n4791) );
  XOR U3216 ( .A(x[1273]), .B(y[1273]), .Z(n4789) );
  XOR U3217 ( .A(x[1562]), .B(y[1562]), .Z(n4788) );
  XOR U3218 ( .A(n4789), .B(n4788), .Z(n4790) );
  XOR U3219 ( .A(n4791), .B(n4790), .Z(n4946) );
  XOR U3220 ( .A(n4947), .B(n4946), .Z(n4166) );
  XOR U3221 ( .A(x[1275]), .B(y[1275]), .Z(n5018) );
  XOR U3222 ( .A(x[206]), .B(y[206]), .Z(n5016) );
  XNOR U3223 ( .A(x[1277]), .B(y[1277]), .Z(n5017) );
  XOR U3224 ( .A(n5016), .B(n5017), .Z(n5019) );
  XNOR U3225 ( .A(n5018), .B(n5019), .Z(n1960) );
  XOR U3226 ( .A(x[1447]), .B(y[1447]), .Z(n1165) );
  XOR U3227 ( .A(x[289]), .B(y[289]), .Z(n1163) );
  XNOR U3228 ( .A(x[1449]), .B(y[1449]), .Z(n1164) );
  XOR U3229 ( .A(n1163), .B(n1164), .Z(n1166) );
  XOR U3230 ( .A(n1165), .B(n1166), .Z(n1961) );
  XNOR U3231 ( .A(n1960), .B(n1961), .Z(n1962) );
  XOR U3232 ( .A(x[1279]), .B(y[1279]), .Z(n1731) );
  XOR U3233 ( .A(x[173]), .B(y[173]), .Z(n1729) );
  XNOR U3234 ( .A(x[1281]), .B(y[1281]), .Z(n1730) );
  XOR U3235 ( .A(n1729), .B(n1730), .Z(n1732) );
  XOR U3236 ( .A(n1731), .B(n1732), .Z(n1963) );
  XOR U3237 ( .A(n1962), .B(n1963), .Z(n4164) );
  XOR U3238 ( .A(x[1283]), .B(y[1283]), .Z(n1744) );
  XOR U3239 ( .A(x[200]), .B(y[200]), .Z(n1742) );
  XOR U3240 ( .A(x[1285]), .B(y[1285]), .Z(n1741) );
  XOR U3241 ( .A(n1742), .B(n1741), .Z(n1743) );
  XOR U3242 ( .A(n1744), .B(n1743), .Z(n4952) );
  XOR U3243 ( .A(x[1443]), .B(y[1443]), .Z(n1181) );
  XOR U3244 ( .A(x[100]), .B(y[100]), .Z(n1179) );
  XNOR U3245 ( .A(x[1445]), .B(y[1445]), .Z(n1180) );
  XOR U3246 ( .A(n1179), .B(n1180), .Z(n1182) );
  XOR U3247 ( .A(n1181), .B(n1182), .Z(n4953) );
  XNOR U3248 ( .A(n4952), .B(n4953), .Z(n4955) );
  XOR U3249 ( .A(x[1287]), .B(y[1287]), .Z(n2003) );
  XOR U3250 ( .A(x[179]), .B(y[179]), .Z(n2001) );
  XOR U3251 ( .A(x[1289]), .B(y[1289]), .Z(n2000) );
  XOR U3252 ( .A(n2001), .B(n2000), .Z(n2002) );
  XOR U3253 ( .A(n2003), .B(n2002), .Z(n4954) );
  XOR U3254 ( .A(n4955), .B(n4954), .Z(n4165) );
  XOR U3255 ( .A(n4164), .B(n4165), .Z(n4167) );
  XOR U3256 ( .A(n4166), .B(n4167), .Z(n5209) );
  XOR U3257 ( .A(x[1243]), .B(y[1243]), .Z(n4798) );
  XOR U3258 ( .A(x[226]), .B(y[226]), .Z(n4796) );
  XNOR U3259 ( .A(x[1245]), .B(y[1245]), .Z(n4797) );
  XOR U3260 ( .A(n4796), .B(n4797), .Z(n4799) );
  XNOR U3261 ( .A(n4798), .B(n4799), .Z(n4986) );
  XOR U3262 ( .A(x[1463]), .B(y[1463]), .Z(n4102) );
  XOR U3263 ( .A(x[1465]), .B(y[1465]), .Z(n4100) );
  XNOR U3264 ( .A(x[1586]), .B(y[1586]), .Z(n4101) );
  XOR U3265 ( .A(n4100), .B(n4101), .Z(n4103) );
  XOR U3266 ( .A(n4102), .B(n4103), .Z(n4987) );
  XNOR U3267 ( .A(n4986), .B(n4987), .Z(n4988) );
  XOR U3268 ( .A(x[1247]), .B(y[1247]), .Z(n5024) );
  XOR U3269 ( .A(x[151]), .B(y[151]), .Z(n5022) );
  XNOR U3270 ( .A(x[1249]), .B(y[1249]), .Z(n5023) );
  XOR U3271 ( .A(n5022), .B(n5023), .Z(n5025) );
  XOR U3272 ( .A(n5024), .B(n5025), .Z(n4989) );
  XOR U3273 ( .A(n4988), .B(n4989), .Z(n3992) );
  XOR U3274 ( .A(x[1251]), .B(y[1251]), .Z(n4775) );
  XOR U3275 ( .A(x[220]), .B(y[220]), .Z(n4773) );
  XOR U3276 ( .A(x[1253]), .B(y[1253]), .Z(n4772) );
  XOR U3277 ( .A(n4773), .B(n4772), .Z(n4774) );
  XOR U3278 ( .A(n4775), .B(n4774), .Z(n1808) );
  XOR U3279 ( .A(x[1459]), .B(y[1459]), .Z(n4005) );
  XOR U3280 ( .A(x[299]), .B(y[299]), .Z(n4003) );
  XOR U3281 ( .A(x[1461]), .B(y[1461]), .Z(n4002) );
  XOR U3282 ( .A(n4003), .B(n4002), .Z(n4004) );
  XOR U3283 ( .A(n4005), .B(n4004), .Z(n1807) );
  XOR U3284 ( .A(n1808), .B(n1807), .Z(n1810) );
  XOR U3285 ( .A(x[1255]), .B(y[1255]), .Z(n4763) );
  XOR U3286 ( .A(x[157]), .B(y[157]), .Z(n4761) );
  XOR U3287 ( .A(x[1257]), .B(y[1257]), .Z(n4760) );
  XOR U3288 ( .A(n4761), .B(n4760), .Z(n4762) );
  XOR U3289 ( .A(n4763), .B(n4762), .Z(n1809) );
  XOR U3290 ( .A(n1810), .B(n1809), .Z(n3991) );
  XOR U3291 ( .A(x[1259]), .B(y[1259]), .Z(n2505) );
  XOR U3292 ( .A(x[161]), .B(y[161]), .Z(n2503) );
  XOR U3293 ( .A(x[1261]), .B(y[1261]), .Z(n2502) );
  XOR U3294 ( .A(n2503), .B(n2502), .Z(n2504) );
  XOR U3295 ( .A(n2505), .B(n2504), .Z(n4948) );
  XOR U3296 ( .A(x[1455]), .B(y[1455]), .Z(n2820) );
  XOR U3297 ( .A(x[1457]), .B(y[1457]), .Z(n2818) );
  XNOR U3298 ( .A(x[1584]), .B(y[1584]), .Z(n2819) );
  XOR U3299 ( .A(n2818), .B(n2819), .Z(n2821) );
  XOR U3300 ( .A(n2820), .B(n2821), .Z(n4949) );
  XNOR U3301 ( .A(n4948), .B(n4949), .Z(n4951) );
  XOR U3302 ( .A(x[1263]), .B(y[1263]), .Z(n1194) );
  XOR U3303 ( .A(x[1265]), .B(y[1265]), .Z(n1192) );
  XOR U3304 ( .A(x[1560]), .B(y[1560]), .Z(n1191) );
  XOR U3305 ( .A(n1192), .B(n1191), .Z(n1193) );
  XOR U3306 ( .A(n1194), .B(n1193), .Z(n4950) );
  XOR U3307 ( .A(n4951), .B(n4950), .Z(n3990) );
  XNOR U3308 ( .A(n3991), .B(n3990), .Z(n3993) );
  XOR U3309 ( .A(n3992), .B(n3993), .Z(n5208) );
  XOR U3310 ( .A(n5209), .B(n5208), .Z(n5211) );
  XOR U3311 ( .A(n5210), .B(n5211), .Z(n1337) );
  XOR U3312 ( .A(x[919]), .B(y[919]), .Z(n2797) );
  XOR U3313 ( .A(x[921]), .B(y[921]), .Z(n2795) );
  XOR U3314 ( .A(x[1518]), .B(y[1518]), .Z(n2794) );
  XOR U3315 ( .A(n2795), .B(n2794), .Z(n2796) );
  XOR U3316 ( .A(n2797), .B(n2796), .Z(n1410) );
  XOR U3317 ( .A(x[927]), .B(y[927]), .Z(n1710) );
  XOR U3318 ( .A(x[82]), .B(y[82]), .Z(n1708) );
  XOR U3319 ( .A(x[929]), .B(y[929]), .Z(n1707) );
  XOR U3320 ( .A(n1708), .B(n1707), .Z(n1709) );
  XOR U3321 ( .A(n1710), .B(n1709), .Z(n1409) );
  XOR U3322 ( .A(n1410), .B(n1409), .Z(n1412) );
  XOR U3323 ( .A(x[935]), .B(y[935]), .Z(n1791) );
  XOR U3324 ( .A(x[74]), .B(y[74]), .Z(n1789) );
  XNOR U3325 ( .A(x[937]), .B(y[937]), .Z(n1790) );
  XOR U3326 ( .A(n1789), .B(n1790), .Z(n1792) );
  XNOR U3327 ( .A(n1791), .B(n1792), .Z(n1411) );
  XOR U3328 ( .A(n1412), .B(n1411), .Z(n3998) );
  XOR U3329 ( .A(x[943]), .B(y[943]), .Z(n4888) );
  XOR U3330 ( .A(x[945]), .B(y[945]), .Z(n4886) );
  XNOR U3331 ( .A(x[1520]), .B(y[1520]), .Z(n4887) );
  XOR U3332 ( .A(n4886), .B(n4887), .Z(n4889) );
  XNOR U3333 ( .A(n4888), .B(n4889), .Z(n1413) );
  XOR U3334 ( .A(x[951]), .B(y[951]), .Z(n4894) );
  XOR U3335 ( .A(x[953]), .B(y[953]), .Z(n4892) );
  XNOR U3336 ( .A(x[1522]), .B(y[1522]), .Z(n4893) );
  XOR U3337 ( .A(n4892), .B(n4893), .Z(n4895) );
  XOR U3338 ( .A(n4894), .B(n4895), .Z(n1414) );
  XNOR U3339 ( .A(n1413), .B(n1414), .Z(n1416) );
  XOR U3340 ( .A(x[959]), .B(y[959]), .Z(n1926) );
  XOR U3341 ( .A(x[54]), .B(y[54]), .Z(n1924) );
  XNOR U3342 ( .A(x[961]), .B(y[961]), .Z(n1925) );
  XOR U3343 ( .A(n1924), .B(n1925), .Z(n1927) );
  XNOR U3344 ( .A(n1926), .B(n1927), .Z(n1415) );
  XOR U3345 ( .A(n1416), .B(n1415), .Z(n3997) );
  XOR U3346 ( .A(x[967]), .B(y[967]), .Z(n1950) );
  XOR U3347 ( .A(x[48]), .B(y[48]), .Z(n1948) );
  XNOR U3348 ( .A(x[969]), .B(y[969]), .Z(n1949) );
  XOR U3349 ( .A(n1948), .B(n1949), .Z(n1951) );
  XNOR U3350 ( .A(n1950), .B(n1951), .Z(n1449) );
  XOR U3351 ( .A(x[975]), .B(y[975]), .Z(n1944) );
  XOR U3352 ( .A(x[977]), .B(y[977]), .Z(n1942) );
  XNOR U3353 ( .A(x[1524]), .B(y[1524]), .Z(n1943) );
  XOR U3354 ( .A(n1942), .B(n1943), .Z(n1945) );
  XOR U3355 ( .A(n1944), .B(n1945), .Z(n1450) );
  XNOR U3356 ( .A(n1449), .B(n1450), .Z(n1452) );
  XOR U3357 ( .A(x[983]), .B(y[983]), .Z(n2529) );
  XOR U3358 ( .A(x[985]), .B(y[985]), .Z(n2526) );
  XNOR U3359 ( .A(x[1526]), .B(y[1526]), .Z(n2527) );
  XOR U3360 ( .A(n2529), .B(n2528), .Z(n1451) );
  XNOR U3361 ( .A(n1452), .B(n1451), .Z(n3996) );
  XOR U3362 ( .A(n3997), .B(n3996), .Z(n3999) );
  XOR U3363 ( .A(n3998), .B(n3999), .Z(n2486) );
  XOR U3364 ( .A(x[847]), .B(y[847]), .Z(n2950) );
  XOR U3365 ( .A(x[849]), .B(y[849]), .Z(n2948) );
  XNOR U3366 ( .A(x[1508]), .B(y[1508]), .Z(n2949) );
  XOR U3367 ( .A(n2948), .B(n2949), .Z(n2951) );
  XNOR U3368 ( .A(n2950), .B(n2951), .Z(n4192) );
  XOR U3369 ( .A(x[855]), .B(y[855]), .Z(n4746) );
  XOR U3370 ( .A(x[857]), .B(y[857]), .Z(n4744) );
  XNOR U3371 ( .A(x[1510]), .B(y[1510]), .Z(n4745) );
  XOR U3372 ( .A(n4744), .B(n4745), .Z(n4747) );
  XOR U3373 ( .A(n4746), .B(n4747), .Z(n4193) );
  XNOR U3374 ( .A(n4192), .B(n4193), .Z(n4195) );
  XOR U3375 ( .A(x[863]), .B(y[863]), .Z(n4360) );
  XOR U3376 ( .A(x[136]), .B(y[136]), .Z(n4358) );
  XNOR U3377 ( .A(x[865]), .B(y[865]), .Z(n4359) );
  XOR U3378 ( .A(n4358), .B(n4359), .Z(n4361) );
  XNOR U3379 ( .A(n4360), .B(n4361), .Z(n4194) );
  XOR U3380 ( .A(n4195), .B(n4194), .Z(n2754) );
  XOR U3381 ( .A(x[871]), .B(y[871]), .Z(n4270) );
  XOR U3382 ( .A(x[130]), .B(y[130]), .Z(n4268) );
  XNOR U3383 ( .A(x[873]), .B(y[873]), .Z(n4269) );
  XOR U3384 ( .A(n4268), .B(n4269), .Z(n4271) );
  XNOR U3385 ( .A(n4270), .B(n4271), .Z(n4171) );
  XOR U3386 ( .A(x[879]), .B(y[879]), .Z(n2993) );
  XOR U3387 ( .A(x[881]), .B(y[881]), .Z(n2991) );
  XOR U3388 ( .A(x[1512]), .B(y[1512]), .Z(n2990) );
  XOR U3389 ( .A(n2991), .B(n2990), .Z(n2992) );
  XOR U3390 ( .A(n2993), .B(n2992), .Z(n4170) );
  XOR U3391 ( .A(n4171), .B(n4170), .Z(n4173) );
  XOR U3392 ( .A(x[887]), .B(y[887]), .Z(n3072) );
  XOR U3393 ( .A(x[889]), .B(y[889]), .Z(n3070) );
  XNOR U3394 ( .A(x[1514]), .B(y[1514]), .Z(n3071) );
  XOR U3395 ( .A(n3070), .B(n3071), .Z(n3073) );
  XNOR U3396 ( .A(n3072), .B(n3073), .Z(n4172) );
  XOR U3397 ( .A(n4173), .B(n4172), .Z(n2753) );
  XOR U3398 ( .A(x[911]), .B(y[911]), .Z(n2766) );
  XOR U3399 ( .A(x[913]), .B(y[913]), .Z(n2764) );
  XNOR U3400 ( .A(x[1516]), .B(y[1516]), .Z(n2765) );
  XOR U3401 ( .A(n2764), .B(n2765), .Z(n2767) );
  XNOR U3402 ( .A(n2766), .B(n2767), .Z(n4235) );
  XOR U3403 ( .A(x[895]), .B(y[895]), .Z(n4019) );
  XOR U3404 ( .A(x[110]), .B(y[110]), .Z(n4017) );
  XOR U3405 ( .A(x[897]), .B(y[897]), .Z(n4016) );
  XOR U3406 ( .A(n4017), .B(n4016), .Z(n4018) );
  XOR U3407 ( .A(n4019), .B(n4018), .Z(n4233) );
  XOR U3408 ( .A(x[903]), .B(y[903]), .Z(n2851) );
  XOR U3409 ( .A(x[102]), .B(y[102]), .Z(n2849) );
  XOR U3410 ( .A(x[905]), .B(y[905]), .Z(n2848) );
  XOR U3411 ( .A(n2849), .B(n2848), .Z(n2850) );
  XOR U3412 ( .A(n2851), .B(n2850), .Z(n4232) );
  XOR U3413 ( .A(n4233), .B(n4232), .Z(n4234) );
  XNOR U3414 ( .A(n4235), .B(n4234), .Z(n2752) );
  XOR U3415 ( .A(n2753), .B(n2752), .Z(n2755) );
  XOR U3416 ( .A(n2754), .B(n2755), .Z(n2485) );
  XOR U3417 ( .A(x[1411]), .B(y[1411]), .Z(n5046) );
  XOR U3418 ( .A(x[120]), .B(y[120]), .Z(n5044) );
  XNOR U3419 ( .A(x[1413]), .B(y[1413]), .Z(n5045) );
  XOR U3420 ( .A(n5044), .B(n5045), .Z(n5047) );
  XNOR U3421 ( .A(n5046), .B(n5047), .Z(n5073) );
  XOR U3422 ( .A(x[1359]), .B(y[1359]), .Z(n1856) );
  XOR U3423 ( .A(x[1361]), .B(y[1361]), .Z(n1853) );
  XNOR U3424 ( .A(x[1572]), .B(y[1572]), .Z(n1854) );
  XNOR U3425 ( .A(n1853), .B(n1854), .Z(n1855) );
  XOR U3426 ( .A(n1856), .B(n1855), .Z(n5072) );
  XOR U3427 ( .A(n5073), .B(n5072), .Z(n5075) );
  XOR U3428 ( .A(x[1339]), .B(y[1339]), .Z(n4936) );
  XOR U3429 ( .A(x[166]), .B(y[166]), .Z(n4934) );
  XNOR U3430 ( .A(x[1341]), .B(y[1341]), .Z(n4935) );
  XOR U3431 ( .A(n4934), .B(n4935), .Z(n4937) );
  XNOR U3432 ( .A(n4936), .B(n4937), .Z(n5074) );
  XOR U3433 ( .A(n5075), .B(n5074), .Z(n1111) );
  XOR U3434 ( .A(x[1379]), .B(y[1379]), .Z(n1646) );
  XOR U3435 ( .A(x[140]), .B(y[140]), .Z(n1643) );
  XNOR U3436 ( .A(x[1381]), .B(y[1381]), .Z(n1644) );
  XOR U3437 ( .A(n1646), .B(n1645), .Z(n1673) );
  XOR U3438 ( .A(x[1399]), .B(y[1399]), .Z(n1737) );
  XOR U3439 ( .A(x[1401]), .B(y[1401]), .Z(n1735) );
  XNOR U3440 ( .A(x[1578]), .B(y[1578]), .Z(n1736) );
  XOR U3441 ( .A(n1735), .B(n1736), .Z(n1738) );
  XOR U3442 ( .A(n1737), .B(n1738), .Z(n1674) );
  XNOR U3443 ( .A(n1673), .B(n1674), .Z(n1676) );
  XOR U3444 ( .A(x[1395]), .B(y[1395]), .Z(n1747) );
  XOR U3445 ( .A(x[255]), .B(y[255]), .Z(n1745) );
  XNOR U3446 ( .A(x[1397]), .B(y[1397]), .Z(n1746) );
  XOR U3447 ( .A(n1745), .B(n1746), .Z(n1748) );
  XNOR U3448 ( .A(n1747), .B(n1748), .Z(n1675) );
  XOR U3449 ( .A(n1676), .B(n1675), .Z(n1110) );
  XOR U3450 ( .A(x[1355]), .B(y[1355]), .Z(n5034) );
  XOR U3451 ( .A(x[227]), .B(y[227]), .Z(n5032) );
  XNOR U3452 ( .A(x[1357]), .B(y[1357]), .Z(n5033) );
  XOR U3453 ( .A(n5032), .B(n5033), .Z(n5035) );
  XNOR U3454 ( .A(n5034), .B(n5035), .Z(n2011) );
  XOR U3455 ( .A(x[1371]), .B(y[1371]), .Z(n4923) );
  XOR U3456 ( .A(x[146]), .B(y[146]), .Z(n4921) );
  XOR U3457 ( .A(x[1373]), .B(y[1373]), .Z(n4920) );
  XOR U3458 ( .A(n4921), .B(n4920), .Z(n4922) );
  XOR U3459 ( .A(n4923), .B(n4922), .Z(n2010) );
  XOR U3460 ( .A(n2011), .B(n2010), .Z(n2013) );
  XOR U3461 ( .A(x[1407]), .B(y[1407]), .Z(n1719) );
  XOR U3462 ( .A(x[261]), .B(y[261]), .Z(n1717) );
  XNOR U3463 ( .A(x[1409]), .B(y[1409]), .Z(n1718) );
  XOR U3464 ( .A(n1717), .B(n1718), .Z(n1720) );
  XNOR U3465 ( .A(n1719), .B(n1720), .Z(n2012) );
  XNOR U3466 ( .A(n2013), .B(n2012), .Z(n1109) );
  XOR U3467 ( .A(n1110), .B(n1109), .Z(n1112) );
  XNOR U3468 ( .A(n1111), .B(n1112), .Z(n2484) );
  XOR U3469 ( .A(n2485), .B(n2484), .Z(n2487) );
  XOR U3470 ( .A(n2486), .B(n2487), .Z(n1336) );
  XOR U3471 ( .A(x[609]), .B(y[609]), .Z(n2237) );
  XOR U3472 ( .A(x[611]), .B(y[611]), .Z(n2235) );
  XOR U3473 ( .A(x[620]), .B(y[620]), .Z(n2234) );
  XOR U3474 ( .A(n2235), .B(n2234), .Z(n2236) );
  XOR U3475 ( .A(n2237), .B(n2236), .Z(n2745) );
  XOR U3476 ( .A(x[613]), .B(y[613]), .Z(n2175) );
  XOR U3477 ( .A(x[350]), .B(y[350]), .Z(n2173) );
  XOR U3478 ( .A(x[615]), .B(y[615]), .Z(n2172) );
  XOR U3479 ( .A(n2173), .B(n2172), .Z(n2174) );
  XOR U3480 ( .A(n2175), .B(n2174), .Z(n2744) );
  XOR U3481 ( .A(n2745), .B(n2744), .Z(n2747) );
  XOR U3482 ( .A(x[617]), .B(y[617]), .Z(n2171) );
  XOR U3483 ( .A(x[344]), .B(y[344]), .Z(n2169) );
  XOR U3484 ( .A(x[619]), .B(y[619]), .Z(n2168) );
  XOR U3485 ( .A(n2169), .B(n2168), .Z(n2170) );
  XOR U3486 ( .A(n2171), .B(n2170), .Z(n2746) );
  XOR U3487 ( .A(n2747), .B(n2746), .Z(n5221) );
  XOR U3488 ( .A(x[621]), .B(y[621]), .Z(n2178) );
  XOR U3489 ( .A(x[623]), .B(y[623]), .Z(n2176) );
  XNOR U3490 ( .A(x[1480]), .B(y[1480]), .Z(n2177) );
  XOR U3491 ( .A(n2176), .B(n2177), .Z(n2179) );
  XNOR U3492 ( .A(n2178), .B(n2179), .Z(n2788) );
  XOR U3493 ( .A(x[625]), .B(y[625]), .Z(n2190) );
  XOR U3494 ( .A(x[336]), .B(y[336]), .Z(n2188) );
  XNOR U3495 ( .A(x[627]), .B(y[627]), .Z(n2189) );
  XOR U3496 ( .A(n2188), .B(n2189), .Z(n2191) );
  XOR U3497 ( .A(n2190), .B(n2191), .Z(n2789) );
  XNOR U3498 ( .A(n2788), .B(n2789), .Z(n2791) );
  XOR U3499 ( .A(x[629]), .B(y[629]), .Z(n2184) );
  XOR U3500 ( .A(x[631]), .B(y[631]), .Z(n2182) );
  XNOR U3501 ( .A(x[1482]), .B(y[1482]), .Z(n2183) );
  XOR U3502 ( .A(n2182), .B(n2183), .Z(n2185) );
  XNOR U3503 ( .A(n2184), .B(n2185), .Z(n2790) );
  XOR U3504 ( .A(n2791), .B(n2790), .Z(n5219) );
  XOR U3505 ( .A(x[633]), .B(y[633]), .Z(n2196) );
  XOR U3506 ( .A(x[606]), .B(y[606]), .Z(n2194) );
  XNOR U3507 ( .A(x[635]), .B(y[635]), .Z(n2195) );
  XOR U3508 ( .A(n2194), .B(n2195), .Z(n2197) );
  XNOR U3509 ( .A(n2196), .B(n2197), .Z(n2808) );
  XOR U3510 ( .A(x[637]), .B(y[637]), .Z(n2094) );
  XOR U3511 ( .A(x[330]), .B(y[330]), .Z(n2092) );
  XNOR U3512 ( .A(x[639]), .B(y[639]), .Z(n2093) );
  XOR U3513 ( .A(n2092), .B(n2093), .Z(n2095) );
  XOR U3514 ( .A(n2094), .B(n2095), .Z(n2809) );
  XNOR U3515 ( .A(n2808), .B(n2809), .Z(n2811) );
  XOR U3516 ( .A(x[641]), .B(y[641]), .Z(n4584) );
  XOR U3517 ( .A(x[600]), .B(y[600]), .Z(n4582) );
  XNOR U3518 ( .A(x[643]), .B(y[643]), .Z(n4583) );
  XOR U3519 ( .A(n4582), .B(n4583), .Z(n4585) );
  XNOR U3520 ( .A(n4584), .B(n4585), .Z(n2810) );
  XNOR U3521 ( .A(n2811), .B(n2810), .Z(n5218) );
  XNOR U3522 ( .A(n5219), .B(n5218), .Z(n5220) );
  XNOR U3523 ( .A(n5221), .B(n5220), .Z(n1329) );
  XOR U3524 ( .A(x[645]), .B(y[645]), .Z(n4068) );
  XOR U3525 ( .A(x[322]), .B(y[322]), .Z(n4066) );
  XNOR U3526 ( .A(x[647]), .B(y[647]), .Z(n4067) );
  XOR U3527 ( .A(n4066), .B(n4067), .Z(n4069) );
  XNOR U3528 ( .A(n4068), .B(n4069), .Z(n2782) );
  XOR U3529 ( .A(x[649]), .B(y[649]), .Z(n2088) );
  XOR U3530 ( .A(x[316]), .B(y[316]), .Z(n2086) );
  XNOR U3531 ( .A(x[651]), .B(y[651]), .Z(n2087) );
  XOR U3532 ( .A(n2086), .B(n2087), .Z(n2089) );
  XOR U3533 ( .A(n2088), .B(n2089), .Z(n2783) );
  XNOR U3534 ( .A(n2782), .B(n2783), .Z(n2785) );
  XOR U3535 ( .A(x[653]), .B(y[653]), .Z(n3020) );
  XOR U3536 ( .A(x[655]), .B(y[655]), .Z(n3018) );
  XNOR U3537 ( .A(x[1484]), .B(y[1484]), .Z(n3019) );
  XOR U3538 ( .A(n3018), .B(n3019), .Z(n3021) );
  XNOR U3539 ( .A(n3020), .B(n3021), .Z(n2784) );
  XOR U3540 ( .A(n2785), .B(n2784), .Z(n1780) );
  XOR U3541 ( .A(x[657]), .B(y[657]), .Z(n4038) );
  XOR U3542 ( .A(x[310]), .B(y[310]), .Z(n4036) );
  XNOR U3543 ( .A(x[659]), .B(y[659]), .Z(n4037) );
  XOR U3544 ( .A(n4036), .B(n4037), .Z(n4039) );
  XNOR U3545 ( .A(n4038), .B(n4039), .Z(n4029) );
  XOR U3546 ( .A(x[661]), .B(y[661]), .Z(n3027) );
  XOR U3547 ( .A(x[663]), .B(y[663]), .Z(n3024) );
  XNOR U3548 ( .A(x[1486]), .B(y[1486]), .Z(n3025) );
  XNOR U3549 ( .A(n3024), .B(n3025), .Z(n3026) );
  XOR U3550 ( .A(n3027), .B(n3026), .Z(n4028) );
  XOR U3551 ( .A(n4029), .B(n4028), .Z(n4031) );
  XOR U3552 ( .A(x[665]), .B(y[665]), .Z(n3928) );
  XOR U3553 ( .A(x[586]), .B(y[586]), .Z(n3926) );
  XNOR U3554 ( .A(x[667]), .B(y[667]), .Z(n3927) );
  XOR U3555 ( .A(n3926), .B(n3927), .Z(n3929) );
  XNOR U3556 ( .A(n3928), .B(n3929), .Z(n4030) );
  XOR U3557 ( .A(n4031), .B(n4030), .Z(n1778) );
  XOR U3558 ( .A(x[669]), .B(y[669]), .Z(n3875) );
  XOR U3559 ( .A(x[302]), .B(y[302]), .Z(n3873) );
  XOR U3560 ( .A(x[671]), .B(y[671]), .Z(n3872) );
  XOR U3561 ( .A(n3873), .B(n3872), .Z(n3874) );
  XOR U3562 ( .A(n3875), .B(n3874), .Z(n2758) );
  XOR U3563 ( .A(x[673]), .B(y[673]), .Z(n3934) );
  XOR U3564 ( .A(x[580]), .B(y[580]), .Z(n3932) );
  XNOR U3565 ( .A(x[675]), .B(y[675]), .Z(n3933) );
  XOR U3566 ( .A(n3932), .B(n3933), .Z(n3935) );
  XOR U3567 ( .A(n3934), .B(n3935), .Z(n2759) );
  XNOR U3568 ( .A(n2758), .B(n2759), .Z(n2761) );
  XOR U3569 ( .A(x[677]), .B(y[677]), .Z(n3895) );
  XOR U3570 ( .A(x[294]), .B(y[294]), .Z(n3893) );
  XOR U3571 ( .A(x[679]), .B(y[679]), .Z(n3892) );
  XOR U3572 ( .A(n3893), .B(n3892), .Z(n3894) );
  XOR U3573 ( .A(n3895), .B(n3894), .Z(n2760) );
  XNOR U3574 ( .A(n2761), .B(n2760), .Z(n1777) );
  XNOR U3575 ( .A(n1778), .B(n1777), .Z(n1779) );
  XOR U3576 ( .A(n1780), .B(n1779), .Z(n1330) );
  XNOR U3577 ( .A(n1329), .B(n1330), .Z(n1331) );
  XOR U3578 ( .A(x[681]), .B(y[681]), .Z(n1249) );
  XOR U3579 ( .A(x[290]), .B(y[290]), .Z(n1247) );
  XNOR U3580 ( .A(x[683]), .B(y[683]), .Z(n1248) );
  XOR U3581 ( .A(n1247), .B(n1248), .Z(n1250) );
  XNOR U3582 ( .A(n1249), .B(n1250), .Z(n2836) );
  XOR U3583 ( .A(x[685]), .B(y[685]), .Z(n1261) );
  XOR U3584 ( .A(x[687]), .B(y[687]), .Z(n1259) );
  XNOR U3585 ( .A(x[1488]), .B(y[1488]), .Z(n1260) );
  XOR U3586 ( .A(n1259), .B(n1260), .Z(n1262) );
  XOR U3587 ( .A(n1261), .B(n1262), .Z(n2837) );
  XNOR U3588 ( .A(n2836), .B(n2837), .Z(n2839) );
  XOR U3589 ( .A(x[689]), .B(y[689]), .Z(n3820) );
  XOR U3590 ( .A(x[282]), .B(y[282]), .Z(n3818) );
  XNOR U3591 ( .A(x[691]), .B(y[691]), .Z(n3819) );
  XOR U3592 ( .A(n3818), .B(n3819), .Z(n3821) );
  XNOR U3593 ( .A(n3820), .B(n3821), .Z(n2838) );
  XOR U3594 ( .A(n2839), .B(n2838), .Z(n2331) );
  XOR U3595 ( .A(x[693]), .B(y[693]), .Z(n3778) );
  XOR U3596 ( .A(x[695]), .B(y[695]), .Z(n3776) );
  XNOR U3597 ( .A(x[1490]), .B(y[1490]), .Z(n3777) );
  XOR U3598 ( .A(n3776), .B(n3777), .Z(n3779) );
  XNOR U3599 ( .A(n3778), .B(n3779), .Z(n2842) );
  XOR U3600 ( .A(x[697]), .B(y[697]), .Z(n1255) );
  XOR U3601 ( .A(x[566]), .B(y[566]), .Z(n1253) );
  XNOR U3602 ( .A(x[699]), .B(y[699]), .Z(n1254) );
  XOR U3603 ( .A(n1253), .B(n1254), .Z(n1256) );
  XOR U3604 ( .A(n1255), .B(n1256), .Z(n2843) );
  XNOR U3605 ( .A(n2842), .B(n2843), .Z(n2845) );
  XOR U3606 ( .A(x[701]), .B(y[701]), .Z(n3763) );
  XOR U3607 ( .A(x[274]), .B(y[274]), .Z(n3761) );
  XOR U3608 ( .A(x[703]), .B(y[703]), .Z(n3760) );
  XOR U3609 ( .A(n3761), .B(n3760), .Z(n3762) );
  XOR U3610 ( .A(n3763), .B(n3762), .Z(n2844) );
  XOR U3611 ( .A(n2845), .B(n2844), .Z(n2329) );
  XOR U3612 ( .A(x[705]), .B(y[705]), .Z(n3722) );
  XOR U3613 ( .A(x[560]), .B(y[560]), .Z(n3720) );
  XNOR U3614 ( .A(x[707]), .B(y[707]), .Z(n3721) );
  XOR U3615 ( .A(n3720), .B(n3721), .Z(n3723) );
  XNOR U3616 ( .A(n3722), .B(n3723), .Z(n2862) );
  XOR U3617 ( .A(x[709]), .B(y[709]), .Z(n3898) );
  XOR U3618 ( .A(x[268]), .B(y[268]), .Z(n3896) );
  XNOR U3619 ( .A(x[711]), .B(y[711]), .Z(n3897) );
  XOR U3620 ( .A(n3896), .B(n3897), .Z(n3899) );
  XOR U3621 ( .A(n3898), .B(n3899), .Z(n2863) );
  XNOR U3622 ( .A(n2862), .B(n2863), .Z(n2865) );
  XOR U3623 ( .A(x[713]), .B(y[713]), .Z(n3707) );
  XOR U3624 ( .A(x[262]), .B(y[262]), .Z(n3705) );
  XOR U3625 ( .A(x[715]), .B(y[715]), .Z(n3704) );
  XOR U3626 ( .A(n3705), .B(n3704), .Z(n3706) );
  XOR U3627 ( .A(n3707), .B(n3706), .Z(n2864) );
  XNOR U3628 ( .A(n2865), .B(n2864), .Z(n2328) );
  XNOR U3629 ( .A(n2329), .B(n2328), .Z(n2330) );
  XOR U3630 ( .A(n2331), .B(n2330), .Z(n1332) );
  XNOR U3631 ( .A(n1331), .B(n1332), .Z(n1335) );
  XOR U3632 ( .A(n1336), .B(n1335), .Z(n1338) );
  XOR U3633 ( .A(n1337), .B(n1338), .Z(n1349) );
  XOR U3634 ( .A(x[1232]), .B(y[1232]), .Z(n4650) );
  XOR U3635 ( .A(x[1228]), .B(y[1228]), .Z(n4648) );
  XNOR U3636 ( .A(x[1230]), .B(y[1230]), .Z(n4649) );
  XOR U3637 ( .A(n4648), .B(n4649), .Z(n4651) );
  XNOR U3638 ( .A(n4650), .B(n4651), .Z(n2298) );
  XOR U3639 ( .A(x[1226]), .B(y[1226]), .Z(n4644) );
  XOR U3640 ( .A(x[1222]), .B(y[1222]), .Z(n4642) );
  XNOR U3641 ( .A(x[1224]), .B(y[1224]), .Z(n4643) );
  XOR U3642 ( .A(n4642), .B(n4643), .Z(n4645) );
  XOR U3643 ( .A(n4644), .B(n4645), .Z(n2299) );
  XNOR U3644 ( .A(n2298), .B(n2299), .Z(n2301) );
  XOR U3645 ( .A(x[1220]), .B(y[1220]), .Z(n4656) );
  XOR U3646 ( .A(x[1216]), .B(y[1216]), .Z(n4654) );
  XNOR U3647 ( .A(x[1218]), .B(y[1218]), .Z(n4655) );
  XOR U3648 ( .A(n4654), .B(n4655), .Z(n4657) );
  XNOR U3649 ( .A(n4656), .B(n4657), .Z(n2300) );
  XOR U3650 ( .A(n2301), .B(n2300), .Z(n1474) );
  XOR U3651 ( .A(x[1244]), .B(y[1244]), .Z(n4686) );
  XOR U3652 ( .A(x[1240]), .B(y[1240]), .Z(n4684) );
  XNOR U3653 ( .A(x[1242]), .B(y[1242]), .Z(n4685) );
  XOR U3654 ( .A(n4684), .B(n4685), .Z(n4687) );
  XNOR U3655 ( .A(n4686), .B(n4687), .Z(n1711) );
  XOR U3656 ( .A(x[362]), .B(y[362]), .Z(n2900) );
  XOR U3657 ( .A(x[354]), .B(y[354]), .Z(n2898) );
  XNOR U3658 ( .A(x[750]), .B(y[750]), .Z(n2899) );
  XOR U3659 ( .A(n2898), .B(n2899), .Z(n2901) );
  XOR U3660 ( .A(n2900), .B(n2901), .Z(n1712) );
  XNOR U3661 ( .A(n1711), .B(n1712), .Z(n1714) );
  XOR U3662 ( .A(x[1238]), .B(y[1238]), .Z(n4692) );
  XOR U3663 ( .A(x[1234]), .B(y[1234]), .Z(n4690) );
  XNOR U3664 ( .A(x[1236]), .B(y[1236]), .Z(n4691) );
  XOR U3665 ( .A(n4690), .B(n4691), .Z(n4693) );
  XNOR U3666 ( .A(n4692), .B(n4693), .Z(n1713) );
  XOR U3667 ( .A(n1714), .B(n1713), .Z(n1472) );
  XOR U3668 ( .A(x[1058]), .B(y[1058]), .Z(n3460) );
  XOR U3669 ( .A(x[1054]), .B(y[1054]), .Z(n3458) );
  XNOR U3670 ( .A(x[1056]), .B(y[1056]), .Z(n3459) );
  XOR U3671 ( .A(n3458), .B(n3459), .Z(n3461) );
  XNOR U3672 ( .A(n3460), .B(n3461), .Z(n1632) );
  XOR U3673 ( .A(x[138]), .B(y[138]), .Z(n2997) );
  XOR U3674 ( .A(x[132]), .B(y[132]), .Z(n2995) );
  XOR U3675 ( .A(x[134]), .B(y[134]), .Z(n2994) );
  XOR U3676 ( .A(n2995), .B(n2994), .Z(n2996) );
  XOR U3677 ( .A(n2997), .B(n2996), .Z(n1631) );
  XOR U3678 ( .A(n1632), .B(n1631), .Z(n1634) );
  XOR U3679 ( .A(x[1052]), .B(y[1052]), .Z(n3466) );
  XOR U3680 ( .A(x[1048]), .B(y[1048]), .Z(n3464) );
  XNOR U3681 ( .A(x[1050]), .B(y[1050]), .Z(n3465) );
  XOR U3682 ( .A(n3464), .B(n3465), .Z(n3467) );
  XNOR U3683 ( .A(n3466), .B(n3467), .Z(n1633) );
  XNOR U3684 ( .A(n1634), .B(n1633), .Z(n1471) );
  XNOR U3685 ( .A(n1472), .B(n1471), .Z(n1473) );
  XNOR U3686 ( .A(n1474), .B(n1473), .Z(n2652) );
  XOR U3687 ( .A(x[1072]), .B(y[1072]), .Z(n3551) );
  XOR U3688 ( .A(x[1066]), .B(y[1066]), .Z(n3549) );
  XOR U3689 ( .A(x[1068]), .B(y[1068]), .Z(n3548) );
  XOR U3690 ( .A(n3549), .B(n3548), .Z(n3550) );
  XOR U3691 ( .A(n3551), .B(n3550), .Z(n4618) );
  XOR U3692 ( .A(x[162]), .B(y[162]), .Z(n4212) );
  XOR U3693 ( .A(x[158]), .B(y[158]), .Z(n4210) );
  XNOR U3694 ( .A(x[678]), .B(y[678]), .Z(n4211) );
  XOR U3695 ( .A(n4210), .B(n4211), .Z(n4213) );
  XOR U3696 ( .A(n4212), .B(n4213), .Z(n4619) );
  XNOR U3697 ( .A(n4618), .B(n4619), .Z(n4621) );
  XOR U3698 ( .A(x[1064]), .B(y[1064]), .Z(n3555) );
  XOR U3699 ( .A(x[1060]), .B(y[1060]), .Z(n3553) );
  XOR U3700 ( .A(x[1062]), .B(y[1062]), .Z(n3552) );
  XOR U3701 ( .A(n3553), .B(n3552), .Z(n3554) );
  XOR U3702 ( .A(n3555), .B(n3554), .Z(n4620) );
  XOR U3703 ( .A(n4621), .B(n4620), .Z(n1468) );
  XOR U3704 ( .A(x[1168]), .B(y[1168]), .Z(n3592) );
  XOR U3705 ( .A(x[1160]), .B(y[1160]), .Z(n3590) );
  XNOR U3706 ( .A(x[1164]), .B(y[1164]), .Z(n3591) );
  XOR U3707 ( .A(n3590), .B(n3591), .Z(n3593) );
  XNOR U3708 ( .A(n3592), .B(n3593), .Z(n5283) );
  XOR U3709 ( .A(x[250]), .B(y[250]), .Z(n4371) );
  XOR U3710 ( .A(x[244]), .B(y[244]), .Z(n4368) );
  XNOR U3711 ( .A(x[710]), .B(y[710]), .Z(n4369) );
  XNOR U3712 ( .A(n4368), .B(n4369), .Z(n4370) );
  XOR U3713 ( .A(n4371), .B(n4370), .Z(n5282) );
  XOR U3714 ( .A(n5283), .B(n5282), .Z(n5285) );
  XOR U3715 ( .A(x[1156]), .B(y[1156]), .Z(n3598) );
  XOR U3716 ( .A(x[1148]), .B(y[1148]), .Z(n3596) );
  XNOR U3717 ( .A(x[1152]), .B(y[1152]), .Z(n3597) );
  XOR U3718 ( .A(n3596), .B(n3597), .Z(n3599) );
  XNOR U3719 ( .A(n3598), .B(n3599), .Z(n5284) );
  XOR U3720 ( .A(n5285), .B(n5284), .Z(n1466) );
  XOR U3721 ( .A(x[1214]), .B(y[1214]), .Z(n3477) );
  XOR U3722 ( .A(x[1210]), .B(y[1210]), .Z(n3475) );
  XOR U3723 ( .A(x[1212]), .B(y[1212]), .Z(n3474) );
  XOR U3724 ( .A(n3475), .B(n3474), .Z(n3476) );
  XOR U3725 ( .A(n3477), .B(n3476), .Z(n2201) );
  XOR U3726 ( .A(x[1208]), .B(y[1208]), .Z(n3473) );
  XOR U3727 ( .A(x[1204]), .B(y[1204]), .Z(n3471) );
  XOR U3728 ( .A(x[1206]), .B(y[1206]), .Z(n3470) );
  XOR U3729 ( .A(n3471), .B(n3470), .Z(n3472) );
  XOR U3730 ( .A(n3473), .B(n3472), .Z(n2200) );
  XOR U3731 ( .A(n2201), .B(n2200), .Z(n2203) );
  XOR U3732 ( .A(x[1202]), .B(y[1202]), .Z(n3481) );
  XOR U3733 ( .A(x[1196]), .B(y[1196]), .Z(n3479) );
  XOR U3734 ( .A(x[1200]), .B(y[1200]), .Z(n3478) );
  XOR U3735 ( .A(n3479), .B(n3478), .Z(n3480) );
  XOR U3736 ( .A(n3481), .B(n3480), .Z(n2202) );
  XNOR U3737 ( .A(n2203), .B(n2202), .Z(n1465) );
  XNOR U3738 ( .A(n1466), .B(n1465), .Z(n1467) );
  XOR U3739 ( .A(n1468), .B(n1467), .Z(n2653) );
  XNOR U3740 ( .A(n2652), .B(n2653), .Z(n2655) );
  XOR U3741 ( .A(x[1046]), .B(y[1046]), .Z(n3489) );
  XOR U3742 ( .A(x[1042]), .B(y[1042]), .Z(n3487) );
  XOR U3743 ( .A(x[1044]), .B(y[1044]), .Z(n3486) );
  XOR U3744 ( .A(n3487), .B(n3486), .Z(n3488) );
  XOR U3745 ( .A(n3489), .B(n3488), .Z(n1612) );
  XOR U3746 ( .A(x[1040]), .B(y[1040]), .Z(n3485) );
  XOR U3747 ( .A(x[1036]), .B(y[1036]), .Z(n3483) );
  XOR U3748 ( .A(x[1038]), .B(y[1038]), .Z(n3482) );
  XOR U3749 ( .A(n3483), .B(n3482), .Z(n3484) );
  XOR U3750 ( .A(n3485), .B(n3484), .Z(n1611) );
  XOR U3751 ( .A(n1612), .B(n1611), .Z(n1614) );
  XOR U3752 ( .A(x[1034]), .B(y[1034]), .Z(n3493) );
  XOR U3753 ( .A(x[1030]), .B(y[1030]), .Z(n3491) );
  XOR U3754 ( .A(x[1032]), .B(y[1032]), .Z(n3490) );
  XOR U3755 ( .A(n3491), .B(n3490), .Z(n3492) );
  XOR U3756 ( .A(n3493), .B(n3492), .Z(n1613) );
  XOR U3757 ( .A(n1614), .B(n1613), .Z(n1520) );
  XOR U3758 ( .A(x[1256]), .B(y[1256]), .Z(n4836) );
  XOR U3759 ( .A(x[1252]), .B(y[1252]), .Z(n4834) );
  XNOR U3760 ( .A(x[1254]), .B(y[1254]), .Z(n4835) );
  XOR U3761 ( .A(n4834), .B(n4835), .Z(n4837) );
  XNOR U3762 ( .A(n4836), .B(n4837), .Z(n4902) );
  XOR U3763 ( .A(x[390]), .B(y[390]), .Z(n2962) );
  XOR U3764 ( .A(x[382]), .B(y[382]), .Z(n2960) );
  XNOR U3765 ( .A(x[388]), .B(y[388]), .Z(n2961) );
  XOR U3766 ( .A(n2960), .B(n2961), .Z(n2963) );
  XOR U3767 ( .A(n2962), .B(n2963), .Z(n4903) );
  XNOR U3768 ( .A(n4902), .B(n4903), .Z(n4905) );
  XOR U3769 ( .A(x[1250]), .B(y[1250]), .Z(n4842) );
  XOR U3770 ( .A(x[1246]), .B(y[1246]), .Z(n4840) );
  XNOR U3771 ( .A(x[1248]), .B(y[1248]), .Z(n4841) );
  XOR U3772 ( .A(n4840), .B(n4841), .Z(n4843) );
  XNOR U3773 ( .A(n4842), .B(n4843), .Z(n4904) );
  XOR U3774 ( .A(n4905), .B(n4904), .Z(n1518) );
  XOR U3775 ( .A(x[1028]), .B(y[1028]), .Z(n3402) );
  XOR U3776 ( .A(x[1024]), .B(y[1024]), .Z(n3400) );
  XNOR U3777 ( .A(x[1026]), .B(y[1026]), .Z(n3401) );
  XOR U3778 ( .A(n3400), .B(n3401), .Z(n3403) );
  XNOR U3779 ( .A(n3402), .B(n3403), .Z(n1561) );
  XOR U3780 ( .A(x[1022]), .B(y[1022]), .Z(n3396) );
  XOR U3781 ( .A(x[1018]), .B(y[1018]), .Z(n3394) );
  XNOR U3782 ( .A(x[1020]), .B(y[1020]), .Z(n3395) );
  XOR U3783 ( .A(n3394), .B(n3395), .Z(n3397) );
  XOR U3784 ( .A(n3396), .B(n3397), .Z(n1562) );
  XNOR U3785 ( .A(n1561), .B(n1562), .Z(n1564) );
  XOR U3786 ( .A(x[1016]), .B(y[1016]), .Z(n3408) );
  XOR U3787 ( .A(x[1012]), .B(y[1012]), .Z(n3406) );
  XNOR U3788 ( .A(x[1014]), .B(y[1014]), .Z(n3407) );
  XOR U3789 ( .A(n3406), .B(n3407), .Z(n3409) );
  XNOR U3790 ( .A(n3408), .B(n3409), .Z(n1563) );
  XNOR U3791 ( .A(n1564), .B(n1563), .Z(n1517) );
  XNOR U3792 ( .A(n1518), .B(n1517), .Z(n1519) );
  XNOR U3793 ( .A(n1520), .B(n1519), .Z(n2654) );
  XOR U3794 ( .A(n2655), .B(n2654), .Z(n5111) );
  XOR U3795 ( .A(x[844]), .B(y[844]), .Z(n1237) );
  XOR U3796 ( .A(x[842]), .B(y[842]), .Z(n1235) );
  XNOR U3797 ( .A(x[1424]), .B(y[1424]), .Z(n1236) );
  XOR U3798 ( .A(n1235), .B(n1236), .Z(n1238) );
  XNOR U3799 ( .A(n1237), .B(n1238), .Z(n4122) );
  XOR U3800 ( .A(x[838]), .B(y[838]), .Z(n1231) );
  XOR U3801 ( .A(x[834]), .B(y[834]), .Z(n1229) );
  XNOR U3802 ( .A(x[1154]), .B(y[1154]), .Z(n1230) );
  XOR U3803 ( .A(n1229), .B(n1230), .Z(n1232) );
  XOR U3804 ( .A(n1231), .B(n1232), .Z(n4123) );
  XNOR U3805 ( .A(n4122), .B(n4123), .Z(n4125) );
  XOR U3806 ( .A(x[832]), .B(y[832]), .Z(n1243) );
  XOR U3807 ( .A(x[830]), .B(y[830]), .Z(n1241) );
  XNOR U3808 ( .A(x[1426]), .B(y[1426]), .Z(n1242) );
  XOR U3809 ( .A(n1241), .B(n1242), .Z(n1244) );
  XNOR U3810 ( .A(n1243), .B(n1244), .Z(n4124) );
  XOR U3811 ( .A(n4125), .B(n4124), .Z(n4522) );
  XOR U3812 ( .A(x[1354]), .B(y[1354]), .Z(n5149) );
  XOR U3813 ( .A(x[1342]), .B(y[1342]), .Z(n5146) );
  XNOR U3814 ( .A(x[1356]), .B(y[1356]), .Z(n5147) );
  XOR U3815 ( .A(n5149), .B(n5148), .Z(n4161) );
  XOR U3816 ( .A(x[548]), .B(y[548]), .Z(n1492) );
  XOR U3817 ( .A(x[542]), .B(y[542]), .Z(n1489) );
  XNOR U3818 ( .A(x[840]), .B(y[840]), .Z(n1490) );
  XOR U3819 ( .A(n1492), .B(n1491), .Z(n4160) );
  XOR U3820 ( .A(n4161), .B(n4160), .Z(n4163) );
  XOR U3821 ( .A(x[1314]), .B(y[1314]), .Z(n5155) );
  XOR U3822 ( .A(x[1322]), .B(y[1322]), .Z(n5152) );
  XNOR U3823 ( .A(x[1358]), .B(y[1358]), .Z(n5153) );
  XOR U3824 ( .A(n5155), .B(n5154), .Z(n4162) );
  XOR U3825 ( .A(n4163), .B(n4162), .Z(n4521) );
  XOR U3826 ( .A(x[828]), .B(y[828]), .Z(n3974) );
  XOR U3827 ( .A(x[826]), .B(y[826]), .Z(n3972) );
  XNOR U3828 ( .A(x[1150]), .B(y[1150]), .Z(n3973) );
  XOR U3829 ( .A(n3972), .B(n3973), .Z(n3975) );
  XNOR U3830 ( .A(n3974), .B(n3975), .Z(n1217) );
  XOR U3831 ( .A(x[824]), .B(y[824]), .Z(n3968) );
  XOR U3832 ( .A(x[820]), .B(y[820]), .Z(n3966) );
  XNOR U3833 ( .A(x[1428]), .B(y[1428]), .Z(n3967) );
  XOR U3834 ( .A(n3966), .B(n3967), .Z(n3969) );
  XOR U3835 ( .A(n3968), .B(n3969), .Z(n1218) );
  XNOR U3836 ( .A(n1217), .B(n1218), .Z(n1220) );
  XOR U3837 ( .A(x[816]), .B(y[816]), .Z(n3980) );
  XOR U3838 ( .A(x[814]), .B(y[814]), .Z(n3978) );
  XNOR U3839 ( .A(x[1146]), .B(y[1146]), .Z(n3979) );
  XOR U3840 ( .A(n3978), .B(n3979), .Z(n3981) );
  XNOR U3841 ( .A(n3980), .B(n3981), .Z(n1219) );
  XNOR U3842 ( .A(n1220), .B(n1219), .Z(n4520) );
  XOR U3843 ( .A(n4521), .B(n4520), .Z(n4523) );
  XOR U3844 ( .A(n4522), .B(n4523), .Z(n4703) );
  XOR U3845 ( .A(x[860]), .B(y[860]), .Z(n991) );
  XOR U3846 ( .A(x[856]), .B(y[856]), .Z(n989) );
  XOR U3847 ( .A(x[1162]), .B(y[1162]), .Z(n988) );
  XOR U3848 ( .A(n989), .B(n988), .Z(n990) );
  XOR U3849 ( .A(n991), .B(n990), .Z(n2483) );
  XOR U3850 ( .A(x[864]), .B(y[864]), .Z(n987) );
  XOR U3851 ( .A(x[862]), .B(y[862]), .Z(n985) );
  XOR U3852 ( .A(x[1420]), .B(y[1420]), .Z(n984) );
  XOR U3853 ( .A(n985), .B(n984), .Z(n986) );
  XOR U3854 ( .A(n987), .B(n986), .Z(n2481) );
  XOR U3855 ( .A(x[171]), .B(y[171]), .Z(n2715) );
  XOR U3856 ( .A(x[175]), .B(y[175]), .Z(n2713) );
  XOR U3857 ( .A(x[476]), .B(y[476]), .Z(n2712) );
  XOR U3858 ( .A(n2713), .B(n2712), .Z(n2714) );
  XOR U3859 ( .A(n2715), .B(n2714), .Z(n2480) );
  XOR U3860 ( .A(n2481), .B(n2480), .Z(n2482) );
  XOR U3861 ( .A(n2483), .B(n2482), .Z(n1355) );
  XOR U3862 ( .A(x[1294]), .B(y[1294]), .Z(n1831) );
  XOR U3863 ( .A(x[1318]), .B(y[1318]), .Z(n1829) );
  XNOR U3864 ( .A(x[1360]), .B(y[1360]), .Z(n1830) );
  XOR U3865 ( .A(n1829), .B(n1830), .Z(n1832) );
  XNOR U3866 ( .A(n1831), .B(n1832), .Z(n1754) );
  XOR U3867 ( .A(x[1312]), .B(y[1312]), .Z(n1825) );
  XOR U3868 ( .A(x[1298]), .B(y[1298]), .Z(n1823) );
  XNOR U3869 ( .A(x[1316]), .B(y[1316]), .Z(n1824) );
  XOR U3870 ( .A(n1823), .B(n1824), .Z(n1826) );
  XNOR U3871 ( .A(n1825), .B(n1826), .Z(n1752) );
  XOR U3872 ( .A(x[532]), .B(y[532]), .Z(n1504) );
  XOR U3873 ( .A(x[528]), .B(y[528]), .Z(n1502) );
  XOR U3874 ( .A(x[530]), .B(y[530]), .Z(n1501) );
  XOR U3875 ( .A(n1502), .B(n1501), .Z(n1503) );
  XOR U3876 ( .A(n1504), .B(n1503), .Z(n1751) );
  XOR U3877 ( .A(n1752), .B(n1751), .Z(n1753) );
  XOR U3878 ( .A(n1754), .B(n1753), .Z(n1354) );
  XOR U3879 ( .A(x[848]), .B(y[848]), .Z(n3962) );
  XOR U3880 ( .A(x[846]), .B(y[846]), .Z(n3960) );
  XNOR U3881 ( .A(x[1158]), .B(y[1158]), .Z(n3961) );
  XOR U3882 ( .A(n3960), .B(n3961), .Z(n3963) );
  XNOR U3883 ( .A(n3962), .B(n3963), .Z(n1031) );
  XOR U3884 ( .A(x[852]), .B(y[852]), .Z(n3956) );
  XOR U3885 ( .A(x[850]), .B(y[850]), .Z(n3954) );
  XNOR U3886 ( .A(x[1422]), .B(y[1422]), .Z(n3955) );
  XOR U3887 ( .A(n3954), .B(n3955), .Z(n3957) );
  XNOR U3888 ( .A(n3956), .B(n3957), .Z(n1028) );
  XOR U3889 ( .A(x[185]), .B(y[185]), .Z(n3108) );
  XOR U3890 ( .A(x[187]), .B(y[187]), .Z(n3106) );
  XNOR U3891 ( .A(x[191]), .B(y[191]), .Z(n3107) );
  XOR U3892 ( .A(n3106), .B(n3107), .Z(n3109) );
  XOR U3893 ( .A(n3108), .B(n3109), .Z(n1029) );
  XNOR U3894 ( .A(n1028), .B(n1029), .Z(n1030) );
  XNOR U3895 ( .A(n1031), .B(n1030), .Z(n1353) );
  XOR U3896 ( .A(n1354), .B(n1353), .Z(n1356) );
  XOR U3897 ( .A(n1355), .B(n1356), .Z(n4701) );
  XOR U3898 ( .A(x[890]), .B(y[890]), .Z(n1290) );
  XOR U3899 ( .A(x[888]), .B(y[888]), .Z(n1288) );
  XOR U3900 ( .A(x[1414]), .B(y[1414]), .Z(n1287) );
  XOR U3901 ( .A(n1288), .B(n1287), .Z(n1289) );
  XOR U3902 ( .A(n1290), .B(n1289), .Z(n3431) );
  XOR U3903 ( .A(x[886]), .B(y[886]), .Z(n1286) );
  XOR U3904 ( .A(x[884]), .B(y[884]), .Z(n1284) );
  XOR U3905 ( .A(x[1174]), .B(y[1174]), .Z(n1283) );
  XOR U3906 ( .A(n1284), .B(n1283), .Z(n1285) );
  XOR U3907 ( .A(n1286), .B(n1285), .Z(n3430) );
  XOR U3908 ( .A(n3431), .B(n3430), .Z(n3433) );
  XOR U3909 ( .A(x[882]), .B(y[882]), .Z(n1294) );
  XOR U3910 ( .A(x[880]), .B(y[880]), .Z(n1292) );
  XOR U3911 ( .A(x[1416]), .B(y[1416]), .Z(n1291) );
  XOR U3912 ( .A(n1292), .B(n1291), .Z(n1293) );
  XOR U3913 ( .A(n1294), .B(n1293), .Z(n3432) );
  XOR U3914 ( .A(n3433), .B(n3432), .Z(n1427) );
  XOR U3915 ( .A(x[1286]), .B(y[1286]), .Z(n4864) );
  XOR U3916 ( .A(x[1284]), .B(y[1284]), .Z(n4862) );
  XNOR U3917 ( .A(x[1320]), .B(y[1320]), .Z(n4863) );
  XOR U3918 ( .A(n4862), .B(n4863), .Z(n4865) );
  XNOR U3919 ( .A(n4864), .B(n4865), .Z(n4806) );
  XOR U3920 ( .A(x[1362]), .B(y[1362]), .Z(n4858) );
  XOR U3921 ( .A(x[1324]), .B(y[1324]), .Z(n4856) );
  XNOR U3922 ( .A(x[1364]), .B(y[1364]), .Z(n4857) );
  XOR U3923 ( .A(n4856), .B(n4857), .Z(n4859) );
  XOR U3924 ( .A(n4858), .B(n4859), .Z(n4807) );
  XNOR U3925 ( .A(n4806), .B(n4807), .Z(n4809) );
  XOR U3926 ( .A(x[1366]), .B(y[1366]), .Z(n4870) );
  XOR U3927 ( .A(x[1282]), .B(y[1282]), .Z(n4868) );
  XNOR U3928 ( .A(x[1326]), .B(y[1326]), .Z(n4869) );
  XOR U3929 ( .A(n4868), .B(n4869), .Z(n4871) );
  XNOR U3930 ( .A(n4870), .B(n4871), .Z(n4808) );
  XOR U3931 ( .A(n4809), .B(n4808), .Z(n1426) );
  XOR U3932 ( .A(x[878]), .B(y[878]), .Z(n1057) );
  XOR U3933 ( .A(x[876]), .B(y[876]), .Z(n1055) );
  XOR U3934 ( .A(x[1170]), .B(y[1170]), .Z(n1054) );
  XOR U3935 ( .A(n1055), .B(n1054), .Z(n1056) );
  XOR U3936 ( .A(n1057), .B(n1056), .Z(n3427) );
  XOR U3937 ( .A(x[874]), .B(y[874]), .Z(n1053) );
  XOR U3938 ( .A(x[870]), .B(y[870]), .Z(n1051) );
  XOR U3939 ( .A(x[1418]), .B(y[1418]), .Z(n1050) );
  XOR U3940 ( .A(n1051), .B(n1050), .Z(n1052) );
  XOR U3941 ( .A(n1053), .B(n1052), .Z(n3426) );
  XOR U3942 ( .A(n3427), .B(n3426), .Z(n3429) );
  XOR U3943 ( .A(x[868]), .B(y[868]), .Z(n1064) );
  XOR U3944 ( .A(x[866]), .B(y[866]), .Z(n1062) );
  XOR U3945 ( .A(x[1166]), .B(y[1166]), .Z(n1061) );
  XOR U3946 ( .A(n1062), .B(n1061), .Z(n1063) );
  XOR U3947 ( .A(n1064), .B(n1063), .Z(n3428) );
  XNOR U3948 ( .A(n3429), .B(n3428), .Z(n1425) );
  XOR U3949 ( .A(n1426), .B(n1425), .Z(n1428) );
  XNOR U3950 ( .A(n1427), .B(n1428), .Z(n4700) );
  XNOR U3951 ( .A(n4701), .B(n4700), .Z(n4702) );
  XNOR U3952 ( .A(n4703), .B(n4702), .Z(n5110) );
  XNOR U3953 ( .A(n5111), .B(n5110), .Z(n5112) );
  XOR U3954 ( .A(x[906]), .B(y[906]), .Z(n968) );
  XOR U3955 ( .A(x[904]), .B(y[904]), .Z(n966) );
  XNOR U3956 ( .A(x[1410]), .B(y[1410]), .Z(n967) );
  XOR U3957 ( .A(n966), .B(n967), .Z(n969) );
  XNOR U3958 ( .A(n968), .B(n969), .Z(n2911) );
  XOR U3959 ( .A(x[99]), .B(y[99]), .Z(n2801) );
  XOR U3960 ( .A(x[103]), .B(y[103]), .Z(n2799) );
  XOR U3961 ( .A(x[105]), .B(y[105]), .Z(n2798) );
  XOR U3962 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3963 ( .A(n2801), .B(n2800), .Z(n2910) );
  XOR U3964 ( .A(n2911), .B(n2910), .Z(n2913) );
  XOR U3965 ( .A(x[902]), .B(y[902]), .Z(n974) );
  XOR U3966 ( .A(x[900]), .B(y[900]), .Z(n972) );
  XNOR U3967 ( .A(x[1182]), .B(y[1182]), .Z(n973) );
  XOR U3968 ( .A(n972), .B(n973), .Z(n975) );
  XNOR U3969 ( .A(n974), .B(n975), .Z(n2912) );
  XOR U3970 ( .A(n2913), .B(n2912), .Z(n1405) );
  XOR U3971 ( .A(x[1280]), .B(y[1280]), .Z(n5235) );
  XOR U3972 ( .A(x[1278]), .B(y[1278]), .Z(n5233) );
  XOR U3973 ( .A(x[1290]), .B(y[1290]), .Z(n5232) );
  XOR U3974 ( .A(n5233), .B(n5232), .Z(n5234) );
  XOR U3975 ( .A(n5235), .B(n5234), .Z(n4785) );
  XOR U3976 ( .A(x[1276]), .B(y[1276]), .Z(n5231) );
  XOR U3977 ( .A(x[1288]), .B(y[1288]), .Z(n5229) );
  XOR U3978 ( .A(x[1368]), .B(y[1368]), .Z(n5228) );
  XOR U3979 ( .A(n5229), .B(n5228), .Z(n5230) );
  XOR U3980 ( .A(n5231), .B(n5230), .Z(n4784) );
  XOR U3981 ( .A(n4785), .B(n4784), .Z(n4787) );
  XOR U3982 ( .A(x[1370]), .B(y[1370]), .Z(n5239) );
  XOR U3983 ( .A(x[1292]), .B(y[1292]), .Z(n5237) );
  XOR U3984 ( .A(x[1372]), .B(y[1372]), .Z(n5236) );
  XOR U3985 ( .A(n5237), .B(n5236), .Z(n5238) );
  XOR U3986 ( .A(n5239), .B(n5238), .Z(n4786) );
  XOR U3987 ( .A(n4787), .B(n4786), .Z(n1404) );
  XOR U3988 ( .A(x[898]), .B(y[898]), .Z(n1018) );
  XOR U3989 ( .A(x[896]), .B(y[896]), .Z(n1016) );
  XNOR U3990 ( .A(x[1412]), .B(y[1412]), .Z(n1017) );
  XOR U3991 ( .A(n1016), .B(n1017), .Z(n1019) );
  XNOR U3992 ( .A(n1018), .B(n1019), .Z(n3494) );
  XOR U3993 ( .A(x[115]), .B(y[115]), .Z(n2804) );
  XOR U3994 ( .A(x[119]), .B(y[119]), .Z(n2802) );
  XNOR U3995 ( .A(x[516]), .B(y[516]), .Z(n2803) );
  XOR U3996 ( .A(n2802), .B(n2803), .Z(n2805) );
  XOR U3997 ( .A(n2804), .B(n2805), .Z(n3495) );
  XNOR U3998 ( .A(n3494), .B(n3495), .Z(n3497) );
  XOR U3999 ( .A(x[894]), .B(y[894]), .Z(n1024) );
  XOR U4000 ( .A(x[892]), .B(y[892]), .Z(n1022) );
  XNOR U4001 ( .A(x[1178]), .B(y[1178]), .Z(n1023) );
  XOR U4002 ( .A(n1022), .B(n1023), .Z(n1025) );
  XNOR U4003 ( .A(n1024), .B(n1025), .Z(n3496) );
  XNOR U4004 ( .A(n3497), .B(n3496), .Z(n1403) );
  XOR U4005 ( .A(n1404), .B(n1403), .Z(n1406) );
  XOR U4006 ( .A(n1405), .B(n1406), .Z(n2063) );
  XOR U4007 ( .A(x[930]), .B(y[930]), .Z(n1273) );
  XOR U4008 ( .A(x[928]), .B(y[928]), .Z(n1271) );
  XNOR U4009 ( .A(x[1404]), .B(y[1404]), .Z(n1272) );
  XOR U4010 ( .A(n1271), .B(n1272), .Z(n1274) );
  XNOR U4011 ( .A(n1273), .B(n1274), .Z(n4470) );
  XOR U4012 ( .A(x[926]), .B(y[926]), .Z(n1267) );
  XOR U4013 ( .A(x[924]), .B(y[924]), .Z(n1265) );
  XNOR U4014 ( .A(x[1194]), .B(y[1194]), .Z(n1266) );
  XOR U4015 ( .A(n1265), .B(n1266), .Z(n1268) );
  XOR U4016 ( .A(n1267), .B(n1268), .Z(n4471) );
  XNOR U4017 ( .A(n4470), .B(n4471), .Z(n4473) );
  XOR U4018 ( .A(x[922]), .B(y[922]), .Z(n1279) );
  XOR U4019 ( .A(x[920]), .B(y[920]), .Z(n1277) );
  XNOR U4020 ( .A(x[1406]), .B(y[1406]), .Z(n1278) );
  XOR U4021 ( .A(n1277), .B(n1278), .Z(n1280) );
  XNOR U4022 ( .A(n1279), .B(n1280), .Z(n4472) );
  XOR U4023 ( .A(n4473), .B(n4472), .Z(n1623) );
  XOR U4024 ( .A(x[1378]), .B(y[1378]), .Z(n2140) );
  XOR U4025 ( .A(x[1308]), .B(y[1308]), .Z(n2138) );
  XNOR U4026 ( .A(x[1380]), .B(y[1380]), .Z(n2139) );
  XOR U4027 ( .A(n2138), .B(n2139), .Z(n2141) );
  XNOR U4028 ( .A(n2140), .B(n2141), .Z(n1210) );
  XOR U4029 ( .A(x[1374]), .B(y[1374]), .Z(n2134) );
  XOR U4030 ( .A(x[1296]), .B(y[1296]), .Z(n2132) );
  XNOR U4031 ( .A(x[1376]), .B(y[1376]), .Z(n2133) );
  XOR U4032 ( .A(n2132), .B(n2133), .Z(n2135) );
  XNOR U4033 ( .A(n2134), .B(n2135), .Z(n1207) );
  XOR U4034 ( .A(x[474]), .B(y[474]), .Z(n1391) );
  XOR U4035 ( .A(x[470]), .B(y[470]), .Z(n1389) );
  XNOR U4036 ( .A(x[800]), .B(y[800]), .Z(n1390) );
  XOR U4037 ( .A(n1389), .B(n1390), .Z(n1392) );
  XOR U4038 ( .A(n1391), .B(n1392), .Z(n1208) );
  XNOR U4039 ( .A(n1207), .B(n1208), .Z(n1209) );
  XOR U4040 ( .A(n1210), .B(n1209), .Z(n1622) );
  XOR U4041 ( .A(x[918]), .B(y[918]), .Z(n932) );
  XOR U4042 ( .A(x[916]), .B(y[916]), .Z(n930) );
  XNOR U4043 ( .A(x[1190]), .B(y[1190]), .Z(n931) );
  XOR U4044 ( .A(n930), .B(n931), .Z(n933) );
  XNOR U4045 ( .A(n932), .B(n933), .Z(n2966) );
  XOR U4046 ( .A(x[914]), .B(y[914]), .Z(n926) );
  XOR U4047 ( .A(x[912]), .B(y[912]), .Z(n924) );
  XNOR U4048 ( .A(x[1408]), .B(y[1408]), .Z(n925) );
  XOR U4049 ( .A(n924), .B(n925), .Z(n927) );
  XOR U4050 ( .A(n926), .B(n927), .Z(n2967) );
  XNOR U4051 ( .A(n2966), .B(n2967), .Z(n2969) );
  XOR U4052 ( .A(x[910]), .B(y[910]), .Z(n938) );
  XOR U4053 ( .A(x[908]), .B(y[908]), .Z(n936) );
  XNOR U4054 ( .A(x[1186]), .B(y[1186]), .Z(n937) );
  XOR U4055 ( .A(n936), .B(n937), .Z(n939) );
  XNOR U4056 ( .A(n938), .B(n939), .Z(n2968) );
  XNOR U4057 ( .A(n2969), .B(n2968), .Z(n1621) );
  XOR U4058 ( .A(n1622), .B(n1621), .Z(n1624) );
  XOR U4059 ( .A(n1623), .B(n1624), .Z(n2061) );
  XOR U4060 ( .A(x[944]), .B(y[944]), .Z(n3390) );
  XOR U4061 ( .A(x[940]), .B(y[940]), .Z(n3388) );
  XNOR U4062 ( .A(x[942]), .B(y[942]), .Z(n3389) );
  XOR U4063 ( .A(n3388), .B(n3389), .Z(n3391) );
  XNOR U4064 ( .A(n3390), .B(n3391), .Z(n1402) );
  XOR U4065 ( .A(x[950]), .B(y[950]), .Z(n3384) );
  XOR U4066 ( .A(x[946]), .B(y[946]), .Z(n3382) );
  XNOR U4067 ( .A(x[948]), .B(y[948]), .Z(n3383) );
  XOR U4068 ( .A(n3382), .B(n3383), .Z(n3385) );
  XNOR U4069 ( .A(n3384), .B(n3385), .Z(n1400) );
  XOR U4070 ( .A(x[27]), .B(y[27]), .Z(n2861) );
  XOR U4071 ( .A(x[31]), .B(y[31]), .Z(n2859) );
  XOR U4072 ( .A(x[33]), .B(y[33]), .Z(n2858) );
  XOR U4073 ( .A(n2859), .B(n2858), .Z(n2860) );
  XOR U4074 ( .A(n2861), .B(n2860), .Z(n1399) );
  XOR U4075 ( .A(n1400), .B(n1399), .Z(n1401) );
  XOR U4076 ( .A(n1402), .B(n1401), .Z(n1543) );
  XOR U4077 ( .A(x[1274]), .B(y[1274]), .Z(n1981) );
  XOR U4078 ( .A(x[1300]), .B(y[1300]), .Z(n1979) );
  XOR U4079 ( .A(x[1382]), .B(y[1382]), .Z(n1978) );
  XOR U4080 ( .A(n1979), .B(n1978), .Z(n1980) );
  XOR U4081 ( .A(n1981), .B(n1980), .Z(n2595) );
  XOR U4082 ( .A(x[458]), .B(y[458]), .Z(n1398) );
  XOR U4083 ( .A(x[452]), .B(y[452]), .Z(n1396) );
  XOR U4084 ( .A(x[456]), .B(y[456]), .Z(n1395) );
  XOR U4085 ( .A(n1396), .B(n1395), .Z(n1397) );
  XOR U4086 ( .A(n1398), .B(n1397), .Z(n2594) );
  XOR U4087 ( .A(n2595), .B(n2594), .Z(n2597) );
  XOR U4088 ( .A(x[1384]), .B(y[1384]), .Z(n1985) );
  XOR U4089 ( .A(x[1310]), .B(y[1310]), .Z(n1983) );
  XOR U4090 ( .A(x[1386]), .B(y[1386]), .Z(n1982) );
  XOR U4091 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U4092 ( .A(n1985), .B(n1984), .Z(n2596) );
  XOR U4093 ( .A(n2597), .B(n2596), .Z(n1542) );
  XOR U4094 ( .A(x[938]), .B(y[938]), .Z(n3348) );
  XOR U4095 ( .A(x[936]), .B(y[936]), .Z(n3346) );
  XNOR U4096 ( .A(x[1402]), .B(y[1402]), .Z(n3347) );
  XOR U4097 ( .A(n3346), .B(n3347), .Z(n3349) );
  XNOR U4098 ( .A(n3348), .B(n3349), .Z(n4514) );
  XOR U4099 ( .A(x[45]), .B(y[45]), .Z(n2826) );
  XOR U4100 ( .A(x[49]), .B(y[49]), .Z(n2824) );
  XNOR U4101 ( .A(x[568]), .B(y[568]), .Z(n2825) );
  XOR U4102 ( .A(n2824), .B(n2825), .Z(n2827) );
  XOR U4103 ( .A(n2826), .B(n2827), .Z(n4515) );
  XNOR U4104 ( .A(n4514), .B(n4515), .Z(n4517) );
  XOR U4105 ( .A(x[934]), .B(y[934]), .Z(n3354) );
  XOR U4106 ( .A(x[932]), .B(y[932]), .Z(n3352) );
  XNOR U4107 ( .A(x[1198]), .B(y[1198]), .Z(n3353) );
  XOR U4108 ( .A(n3352), .B(n3353), .Z(n3355) );
  XNOR U4109 ( .A(n3354), .B(n3355), .Z(n4516) );
  XNOR U4110 ( .A(n4517), .B(n4516), .Z(n1541) );
  XOR U4111 ( .A(n1542), .B(n1541), .Z(n1544) );
  XNOR U4112 ( .A(n1543), .B(n1544), .Z(n2060) );
  XNOR U4113 ( .A(n2061), .B(n2060), .Z(n2062) );
  XOR U4114 ( .A(n2063), .B(n2062), .Z(n5113) );
  XNOR U4115 ( .A(n5112), .B(n5113), .Z(n1347) );
  XOR U4116 ( .A(x[273]), .B(y[273]), .Z(n3132) );
  XOR U4117 ( .A(x[275]), .B(y[275]), .Z(n3130) );
  XNOR U4118 ( .A(x[394]), .B(y[394]), .Z(n3131) );
  XOR U4119 ( .A(n3130), .B(n3131), .Z(n3133) );
  XNOR U4120 ( .A(n3132), .B(n3133), .Z(n3690) );
  XOR U4121 ( .A(x[1511]), .B(y[1511]), .Z(n2932) );
  XOR U4122 ( .A(x[333]), .B(y[333]), .Z(n2930) );
  XNOR U4123 ( .A(x[1513]), .B(y[1513]), .Z(n2931) );
  XOR U4124 ( .A(n2930), .B(n2931), .Z(n2933) );
  XOR U4125 ( .A(n2932), .B(n2933), .Z(n3691) );
  XNOR U4126 ( .A(n3690), .B(n3691), .Z(n3692) );
  XOR U4127 ( .A(x[279]), .B(y[279]), .Z(n3144) );
  XOR U4128 ( .A(x[281]), .B(y[281]), .Z(n3142) );
  XNOR U4129 ( .A(x[285]), .B(y[285]), .Z(n3143) );
  XOR U4130 ( .A(n3142), .B(n3143), .Z(n3145) );
  XOR U4131 ( .A(n3144), .B(n3145), .Z(n3693) );
  XOR U4132 ( .A(n3692), .B(n3693), .Z(n2916) );
  XOR U4133 ( .A(x[287]), .B(y[287]), .Z(n3198) );
  XOR U4134 ( .A(x[291]), .B(y[291]), .Z(n3196) );
  XNOR U4135 ( .A(x[295]), .B(y[295]), .Z(n3197) );
  XOR U4136 ( .A(n3196), .B(n3197), .Z(n3199) );
  XNOR U4137 ( .A(n3198), .B(n3199), .Z(n3678) );
  XOR U4138 ( .A(x[987]), .B(y[987]), .Z(n2522) );
  XOR U4139 ( .A(x[386]), .B(y[386]), .Z(n2520) );
  XNOR U4140 ( .A(x[989]), .B(y[989]), .Z(n2521) );
  XOR U4141 ( .A(n2520), .B(n2521), .Z(n2523) );
  XOR U4142 ( .A(n2522), .B(n2523), .Z(n3679) );
  XNOR U4143 ( .A(n3678), .B(n3679), .Z(n3680) );
  XOR U4144 ( .A(x[297]), .B(y[297]), .Z(n3192) );
  XOR U4145 ( .A(x[301]), .B(y[301]), .Z(n3190) );
  XNOR U4146 ( .A(x[368]), .B(y[368]), .Z(n3191) );
  XOR U4147 ( .A(n3190), .B(n3191), .Z(n3193) );
  XOR U4148 ( .A(n3192), .B(n3193), .Z(n3681) );
  XOR U4149 ( .A(n3680), .B(n3681), .Z(n2914) );
  XOR U4150 ( .A(x[303]), .B(y[303]), .Z(n3204) );
  XOR U4151 ( .A(x[307]), .B(y[307]), .Z(n3202) );
  XNOR U4152 ( .A(x[358]), .B(y[358]), .Z(n3203) );
  XOR U4153 ( .A(n3202), .B(n3203), .Z(n3205) );
  XNOR U4154 ( .A(n3204), .B(n3205), .Z(n3714) );
  XOR U4155 ( .A(x[1507]), .B(y[1507]), .Z(n4602) );
  XOR U4156 ( .A(x[60]), .B(y[60]), .Z(n4600) );
  XNOR U4157 ( .A(x[1509]), .B(y[1509]), .Z(n4601) );
  XOR U4158 ( .A(n4600), .B(n4601), .Z(n4603) );
  XOR U4159 ( .A(n4602), .B(n4603), .Z(n3715) );
  XNOR U4160 ( .A(n3714), .B(n3715), .Z(n3717) );
  XOR U4161 ( .A(x[319]), .B(y[319]), .Z(n3162) );
  XOR U4162 ( .A(x[323]), .B(y[323]), .Z(n3160) );
  XNOR U4163 ( .A(x[325]), .B(y[325]), .Z(n3161) );
  XOR U4164 ( .A(n3160), .B(n3161), .Z(n3163) );
  XNOR U4165 ( .A(n3162), .B(n3163), .Z(n3716) );
  XNOR U4166 ( .A(n3717), .B(n3716), .Z(n2915) );
  XOR U4167 ( .A(n2914), .B(n2915), .Z(n2917) );
  XOR U4168 ( .A(n2916), .B(n2917), .Z(n5187) );
  XOR U4169 ( .A(x[335]), .B(y[335]), .Z(n3856) );
  XOR U4170 ( .A(x[324]), .B(y[324]), .Z(n3854) );
  XNOR U4171 ( .A(x[339]), .B(y[339]), .Z(n3855) );
  XOR U4172 ( .A(n3854), .B(n3855), .Z(n3857) );
  XNOR U4173 ( .A(n3856), .B(n3857), .Z(n3744) );
  XOR U4174 ( .A(x[995]), .B(y[995]), .Z(n2534) );
  XOR U4175 ( .A(x[380]), .B(y[380]), .Z(n2532) );
  XNOR U4176 ( .A(x[997]), .B(y[997]), .Z(n2533) );
  XOR U4177 ( .A(n2532), .B(n2533), .Z(n2535) );
  XOR U4178 ( .A(n2534), .B(n2535), .Z(n3745) );
  XNOR U4179 ( .A(n3744), .B(n3745), .Z(n3746) );
  XOR U4180 ( .A(x[341]), .B(y[341]), .Z(n3850) );
  XOR U4181 ( .A(x[345]), .B(y[345]), .Z(n3848) );
  XNOR U4182 ( .A(x[347]), .B(y[347]), .Z(n3849) );
  XOR U4183 ( .A(n3848), .B(n3849), .Z(n3851) );
  XOR U4184 ( .A(n3850), .B(n3851), .Z(n3747) );
  XOR U4185 ( .A(n3746), .B(n3747), .Z(n4674) );
  XOR U4186 ( .A(x[351]), .B(y[351]), .Z(n3862) );
  XOR U4187 ( .A(x[353]), .B(y[353]), .Z(n3860) );
  XNOR U4188 ( .A(x[357]), .B(y[357]), .Z(n3861) );
  XOR U4189 ( .A(n3860), .B(n3861), .Z(n3863) );
  XNOR U4190 ( .A(n3862), .B(n3863), .Z(n3764) );
  XOR U4191 ( .A(x[1503]), .B(y[1503]), .Z(n1595) );
  XOR U4192 ( .A(x[327]), .B(y[327]), .Z(n1593) );
  XNOR U4193 ( .A(x[1505]), .B(y[1505]), .Z(n1594) );
  XOR U4194 ( .A(n1593), .B(n1594), .Z(n1596) );
  XOR U4195 ( .A(n1595), .B(n1596), .Z(n3765) );
  XNOR U4196 ( .A(n3764), .B(n3765), .Z(n3766) );
  XOR U4197 ( .A(x[361]), .B(y[361]), .Z(n3838) );
  XOR U4198 ( .A(x[296]), .B(y[296]), .Z(n3836) );
  XNOR U4199 ( .A(x[363]), .B(y[363]), .Z(n3837) );
  XOR U4200 ( .A(n3836), .B(n3837), .Z(n3839) );
  XOR U4201 ( .A(n3838), .B(n3839), .Z(n3767) );
  XOR U4202 ( .A(n3766), .B(n3767), .Z(n4672) );
  XOR U4203 ( .A(x[367]), .B(y[367]), .Z(n3832) );
  XOR U4204 ( .A(x[288]), .B(y[288]), .Z(n3830) );
  XNOR U4205 ( .A(x[369]), .B(y[369]), .Z(n3831) );
  XOR U4206 ( .A(n3830), .B(n3831), .Z(n3833) );
  XNOR U4207 ( .A(n3832), .B(n3833), .Z(n3738) );
  XOR U4208 ( .A(x[1003]), .B(y[1003]), .Z(n4376) );
  XOR U4209 ( .A(x[14]), .B(y[14]), .Z(n4374) );
  XNOR U4210 ( .A(x[1005]), .B(y[1005]), .Z(n4375) );
  XOR U4211 ( .A(n4374), .B(n4375), .Z(n4377) );
  XOR U4212 ( .A(n4376), .B(n4377), .Z(n3739) );
  XNOR U4213 ( .A(n3738), .B(n3739), .Z(n3741) );
  XOR U4214 ( .A(x[373]), .B(y[373]), .Z(n3844) );
  XOR U4215 ( .A(x[375]), .B(y[375]), .Z(n3842) );
  XNOR U4216 ( .A(x[379]), .B(y[379]), .Z(n3843) );
  XOR U4217 ( .A(n3842), .B(n3843), .Z(n3845) );
  XNOR U4218 ( .A(n3844), .B(n3845), .Z(n3740) );
  XNOR U4219 ( .A(n3741), .B(n3740), .Z(n4673) );
  XOR U4220 ( .A(n4672), .B(n4673), .Z(n4675) );
  XOR U4221 ( .A(n4674), .B(n4675), .Z(n5186) );
  XOR U4222 ( .A(n5187), .B(n5186), .Z(n5189) );
  XOR U4223 ( .A(x[383]), .B(y[383]), .Z(n3330) );
  XOR U4224 ( .A(x[385]), .B(y[385]), .Z(n3328) );
  XNOR U4225 ( .A(x[387]), .B(y[387]), .Z(n3329) );
  XOR U4226 ( .A(n3328), .B(n3329), .Z(n3331) );
  XNOR U4227 ( .A(n3330), .B(n3331), .Z(n3794) );
  XOR U4228 ( .A(x[1499]), .B(y[1499]), .Z(n1485) );
  XOR U4229 ( .A(x[66]), .B(y[66]), .Z(n1483) );
  XNOR U4230 ( .A(x[1501]), .B(y[1501]), .Z(n1484) );
  XOR U4231 ( .A(n1483), .B(n1484), .Z(n1486) );
  XOR U4232 ( .A(n1485), .B(n1486), .Z(n3795) );
  XNOR U4233 ( .A(n3794), .B(n3795), .Z(n3797) );
  XOR U4234 ( .A(x[389]), .B(y[389]), .Z(n3324) );
  XOR U4235 ( .A(x[258]), .B(y[258]), .Z(n3322) );
  XNOR U4236 ( .A(x[391]), .B(y[391]), .Z(n3323) );
  XOR U4237 ( .A(n3322), .B(n3323), .Z(n3325) );
  XNOR U4238 ( .A(n3324), .B(n3325), .Z(n3796) );
  XOR U4239 ( .A(n3797), .B(n3796), .Z(n4627) );
  XOR U4240 ( .A(x[393]), .B(y[393]), .Z(n3336) );
  XOR U4241 ( .A(x[252]), .B(y[252]), .Z(n3334) );
  XNOR U4242 ( .A(x[395]), .B(y[395]), .Z(n3335) );
  XOR U4243 ( .A(n3334), .B(n3335), .Z(n3337) );
  XNOR U4244 ( .A(n3336), .B(n3337), .Z(n3800) );
  XOR U4245 ( .A(x[1011]), .B(y[1011]), .Z(n2548) );
  XOR U4246 ( .A(x[8]), .B(y[8]), .Z(n2546) );
  XNOR U4247 ( .A(x[1013]), .B(y[1013]), .Z(n2547) );
  XOR U4248 ( .A(n2546), .B(n2547), .Z(n2549) );
  XOR U4249 ( .A(n2548), .B(n2549), .Z(n3801) );
  XNOR U4250 ( .A(n3800), .B(n3801), .Z(n3803) );
  XOR U4251 ( .A(x[397]), .B(y[397]), .Z(n3306) );
  XOR U4252 ( .A(x[399]), .B(y[399]), .Z(n3304) );
  XNOR U4253 ( .A(x[401]), .B(y[401]), .Z(n3305) );
  XOR U4254 ( .A(n3304), .B(n3305), .Z(n3307) );
  XNOR U4255 ( .A(n3306), .B(n3307), .Z(n3802) );
  XOR U4256 ( .A(n3803), .B(n3802), .Z(n4625) );
  XOR U4257 ( .A(x[403]), .B(y[403]), .Z(n3300) );
  XOR U4258 ( .A(x[405]), .B(y[405]), .Z(n3298) );
  XNOR U4259 ( .A(x[407]), .B(y[407]), .Z(n3299) );
  XOR U4260 ( .A(n3298), .B(n3299), .Z(n3301) );
  XNOR U4261 ( .A(n3300), .B(n3301), .Z(n3824) );
  XOR U4262 ( .A(x[1495]), .B(y[1495]), .Z(n4484) );
  XOR U4263 ( .A(x[1497]), .B(y[1497]), .Z(n4482) );
  XNOR U4264 ( .A(x[1590]), .B(y[1590]), .Z(n4483) );
  XOR U4265 ( .A(n4482), .B(n4483), .Z(n4485) );
  XOR U4266 ( .A(n4484), .B(n4485), .Z(n3825) );
  XNOR U4267 ( .A(n3824), .B(n3825), .Z(n3827) );
  XOR U4268 ( .A(x[409]), .B(y[409]), .Z(n3312) );
  XOR U4269 ( .A(x[224]), .B(y[224]), .Z(n3310) );
  XNOR U4270 ( .A(x[411]), .B(y[411]), .Z(n3311) );
  XOR U4271 ( .A(n3310), .B(n3311), .Z(n3313) );
  XNOR U4272 ( .A(n3312), .B(n3313), .Z(n3826) );
  XNOR U4273 ( .A(n3827), .B(n3826), .Z(n4624) );
  XNOR U4274 ( .A(n4625), .B(n4624), .Z(n4626) );
  XNOR U4275 ( .A(n4627), .B(n4626), .Z(n5188) );
  XOR U4276 ( .A(n5189), .B(n5188), .Z(n2661) );
  XOR U4277 ( .A(x[413]), .B(y[413]), .Z(n3282) );
  XOR U4278 ( .A(x[216]), .B(y[216]), .Z(n3280) );
  XNOR U4279 ( .A(x[415]), .B(y[415]), .Z(n3281) );
  XOR U4280 ( .A(n3280), .B(n3281), .Z(n3283) );
  XNOR U4281 ( .A(n3282), .B(n3283), .Z(n3902) );
  XOR U4282 ( .A(x[1019]), .B(y[1019]), .Z(n4994) );
  XOR U4283 ( .A(x[366]), .B(y[366]), .Z(n4992) );
  XNOR U4284 ( .A(x[1021]), .B(y[1021]), .Z(n4993) );
  XOR U4285 ( .A(n4992), .B(n4993), .Z(n4995) );
  XOR U4286 ( .A(n4994), .B(n4995), .Z(n3903) );
  XNOR U4287 ( .A(n3902), .B(n3903), .Z(n3905) );
  XOR U4288 ( .A(x[417]), .B(y[417]), .Z(n3276) );
  XOR U4289 ( .A(x[419]), .B(y[419]), .Z(n3274) );
  XNOR U4290 ( .A(x[421]), .B(y[421]), .Z(n3275) );
  XOR U4291 ( .A(n3274), .B(n3275), .Z(n3277) );
  XNOR U4292 ( .A(n3276), .B(n3277), .Z(n3904) );
  XOR U4293 ( .A(n3905), .B(n3904), .Z(n1618) );
  XOR U4294 ( .A(x[423]), .B(y[423]), .Z(n3288) );
  XOR U4295 ( .A(x[425]), .B(y[425]), .Z(n3286) );
  XNOR U4296 ( .A(x[427]), .B(y[427]), .Z(n3287) );
  XOR U4297 ( .A(n3286), .B(n3287), .Z(n3289) );
  XNOR U4298 ( .A(n3288), .B(n3289), .Z(n3770) );
  XOR U4299 ( .A(x[1491]), .B(y[1491]), .Z(n1385) );
  XOR U4300 ( .A(x[321]), .B(y[321]), .Z(n1383) );
  XNOR U4301 ( .A(x[1493]), .B(y[1493]), .Z(n1384) );
  XOR U4302 ( .A(n1383), .B(n1384), .Z(n1386) );
  XOR U4303 ( .A(n1385), .B(n1386), .Z(n3771) );
  XNOR U4304 ( .A(n3770), .B(n3771), .Z(n3773) );
  XOR U4305 ( .A(x[429]), .B(y[429]), .Z(n3264) );
  XOR U4306 ( .A(x[190]), .B(y[190]), .Z(n3262) );
  XNOR U4307 ( .A(x[431]), .B(y[431]), .Z(n3263) );
  XOR U4308 ( .A(n3262), .B(n3263), .Z(n3265) );
  XNOR U4309 ( .A(n3264), .B(n3265), .Z(n3772) );
  XOR U4310 ( .A(n3773), .B(n3772), .Z(n1616) );
  XOR U4311 ( .A(x[433]), .B(y[433]), .Z(n3258) );
  XOR U4312 ( .A(x[182]), .B(y[182]), .Z(n3256) );
  XNOR U4313 ( .A(x[435]), .B(y[435]), .Z(n3257) );
  XOR U4314 ( .A(n3256), .B(n3257), .Z(n3259) );
  XNOR U4315 ( .A(n3258), .B(n3259), .Z(n3938) );
  XOR U4316 ( .A(x[1027]), .B(y[1027]), .Z(n1079) );
  XOR U4317 ( .A(x[360]), .B(y[360]), .Z(n1077) );
  XNOR U4318 ( .A(x[1029]), .B(y[1029]), .Z(n1078) );
  XOR U4319 ( .A(n1077), .B(n1078), .Z(n1080) );
  XOR U4320 ( .A(n1079), .B(n1080), .Z(n3939) );
  XNOR U4321 ( .A(n3938), .B(n3939), .Z(n3941) );
  XOR U4322 ( .A(x[437]), .B(y[437]), .Z(n3270) );
  XOR U4323 ( .A(x[439]), .B(y[439]), .Z(n3268) );
  XNOR U4324 ( .A(x[441]), .B(y[441]), .Z(n3269) );
  XOR U4325 ( .A(n3268), .B(n3269), .Z(n3271) );
  XNOR U4326 ( .A(n3270), .B(n3271), .Z(n3940) );
  XNOR U4327 ( .A(n3941), .B(n3940), .Z(n1615) );
  XNOR U4328 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U4329 ( .A(n1618), .B(n1617), .Z(n2054) );
  XOR U4330 ( .A(x[443]), .B(y[443]), .Z(n3240) );
  XOR U4331 ( .A(x[445]), .B(y[445]), .Z(n3238) );
  XNOR U4332 ( .A(x[447]), .B(y[447]), .Z(n3239) );
  XOR U4333 ( .A(n3238), .B(n3239), .Z(n3241) );
  XNOR U4334 ( .A(n3240), .B(n3241), .Z(n3866) );
  XOR U4335 ( .A(x[1487]), .B(y[1487]), .Z(n4454) );
  XOR U4336 ( .A(x[1489]), .B(y[1489]), .Z(n4452) );
  XNOR U4337 ( .A(x[1588]), .B(y[1588]), .Z(n4453) );
  XOR U4338 ( .A(n4452), .B(n4453), .Z(n4455) );
  XOR U4339 ( .A(n4454), .B(n4455), .Z(n3867) );
  XNOR U4340 ( .A(n3866), .B(n3867), .Z(n3869) );
  XOR U4341 ( .A(x[449]), .B(y[449]), .Z(n3234) );
  XOR U4342 ( .A(x[154]), .B(y[154]), .Z(n3232) );
  XNOR U4343 ( .A(x[451]), .B(y[451]), .Z(n3233) );
  XOR U4344 ( .A(n3232), .B(n3233), .Z(n3235) );
  XNOR U4345 ( .A(n3234), .B(n3235), .Z(n3868) );
  XOR U4346 ( .A(n3869), .B(n3868), .Z(n4579) );
  XOR U4347 ( .A(x[453]), .B(y[453]), .Z(n3246) );
  XOR U4348 ( .A(x[148]), .B(y[148]), .Z(n3244) );
  XNOR U4349 ( .A(x[455]), .B(y[455]), .Z(n3245) );
  XOR U4350 ( .A(n3244), .B(n3245), .Z(n3247) );
  XNOR U4351 ( .A(n3246), .B(n3247), .Z(n3316) );
  XOR U4352 ( .A(x[1035]), .B(y[1035]), .Z(n1085) );
  XOR U4353 ( .A(x[7]), .B(y[7]), .Z(n1083) );
  XNOR U4354 ( .A(x[1037]), .B(y[1037]), .Z(n1084) );
  XOR U4355 ( .A(n1083), .B(n1084), .Z(n1086) );
  XOR U4356 ( .A(n1085), .B(n1086), .Z(n3317) );
  XNOR U4357 ( .A(n3316), .B(n3317), .Z(n3319) );
  XOR U4358 ( .A(x[457]), .B(y[457]), .Z(n3222) );
  XOR U4359 ( .A(x[459]), .B(y[459]), .Z(n3220) );
  XNOR U4360 ( .A(x[461]), .B(y[461]), .Z(n3221) );
  XOR U4361 ( .A(n3220), .B(n3221), .Z(n3223) );
  XNOR U4362 ( .A(n3222), .B(n3223), .Z(n3318) );
  XOR U4363 ( .A(n3319), .B(n3318), .Z(n4577) );
  XOR U4364 ( .A(x[463]), .B(y[463]), .Z(n3216) );
  XOR U4365 ( .A(x[465]), .B(y[465]), .Z(n3214) );
  XNOR U4366 ( .A(x[467]), .B(y[467]), .Z(n3215) );
  XOR U4367 ( .A(n3214), .B(n3215), .Z(n3217) );
  XNOR U4368 ( .A(n3216), .B(n3217), .Z(n3292) );
  XOR U4369 ( .A(x[1483]), .B(y[1483]), .Z(n2894) );
  XOR U4370 ( .A(x[315]), .B(y[315]), .Z(n2892) );
  XNOR U4371 ( .A(x[1485]), .B(y[1485]), .Z(n2893) );
  XOR U4372 ( .A(n2892), .B(n2893), .Z(n2895) );
  XOR U4373 ( .A(n2894), .B(n2895), .Z(n3293) );
  XNOR U4374 ( .A(n3292), .B(n3293), .Z(n3295) );
  XOR U4375 ( .A(x[469]), .B(y[469]), .Z(n3228) );
  XOR U4376 ( .A(x[118]), .B(y[118]), .Z(n3226) );
  XNOR U4377 ( .A(x[471]), .B(y[471]), .Z(n3227) );
  XOR U4378 ( .A(n3226), .B(n3227), .Z(n3229) );
  XNOR U4379 ( .A(n3228), .B(n3229), .Z(n3294) );
  XNOR U4380 ( .A(n3295), .B(n3294), .Z(n4576) );
  XNOR U4381 ( .A(n4577), .B(n4576), .Z(n4578) );
  XOR U4382 ( .A(n4579), .B(n4578), .Z(n2055) );
  XNOR U4383 ( .A(n2054), .B(n2055), .Z(n2057) );
  XOR U4384 ( .A(x[473]), .B(y[473]), .Z(n2116) );
  XOR U4385 ( .A(x[112]), .B(y[112]), .Z(n2114) );
  XNOR U4386 ( .A(x[475]), .B(y[475]), .Z(n2115) );
  XOR U4387 ( .A(n2114), .B(n2115), .Z(n2117) );
  XNOR U4388 ( .A(n2116), .B(n2117), .Z(n3250) );
  XOR U4389 ( .A(x[1043]), .B(y[1043]), .Z(n1091) );
  XOR U4390 ( .A(x[13]), .B(y[13]), .Z(n1089) );
  XNOR U4391 ( .A(x[1045]), .B(y[1045]), .Z(n1090) );
  XOR U4392 ( .A(n1089), .B(n1090), .Z(n1092) );
  XOR U4393 ( .A(n1091), .B(n1092), .Z(n3251) );
  XNOR U4394 ( .A(n3250), .B(n3251), .Z(n3253) );
  XOR U4395 ( .A(x[477]), .B(y[477]), .Z(n2110) );
  XOR U4396 ( .A(x[479]), .B(y[479]), .Z(n2108) );
  XNOR U4397 ( .A(x[481]), .B(y[481]), .Z(n2109) );
  XOR U4398 ( .A(n2108), .B(n2109), .Z(n2111) );
  XNOR U4399 ( .A(n2110), .B(n2111), .Z(n3252) );
  XOR U4400 ( .A(n3253), .B(n3252), .Z(n4573) );
  XOR U4401 ( .A(x[483]), .B(y[483]), .Z(n2122) );
  XOR U4402 ( .A(x[485]), .B(y[485]), .Z(n2120) );
  XNOR U4403 ( .A(x[487]), .B(y[487]), .Z(n2121) );
  XOR U4404 ( .A(n2120), .B(n2121), .Z(n2123) );
  XNOR U4405 ( .A(n2122), .B(n2123), .Z(n3154) );
  XOR U4406 ( .A(x[1479]), .B(y[1479]), .Z(n4412) );
  XOR U4407 ( .A(x[311]), .B(y[311]), .Z(n4410) );
  XNOR U4408 ( .A(x[1481]), .B(y[1481]), .Z(n4411) );
  XOR U4409 ( .A(n4410), .B(n4411), .Z(n4413) );
  XOR U4410 ( .A(n4412), .B(n4413), .Z(n3155) );
  XNOR U4411 ( .A(n3154), .B(n3155), .Z(n3157) );
  XOR U4412 ( .A(x[489]), .B(y[489]), .Z(n2152) );
  XOR U4413 ( .A(x[84]), .B(y[84]), .Z(n2150) );
  XNOR U4414 ( .A(x[491]), .B(y[491]), .Z(n2151) );
  XOR U4415 ( .A(n2150), .B(n2151), .Z(n2153) );
  XNOR U4416 ( .A(n2152), .B(n2153), .Z(n3156) );
  XOR U4417 ( .A(n3157), .B(n3156), .Z(n4571) );
  XOR U4418 ( .A(x[493]), .B(y[493]), .Z(n2146) );
  XOR U4419 ( .A(x[76]), .B(y[76]), .Z(n2144) );
  XNOR U4420 ( .A(x[495]), .B(y[495]), .Z(n2145) );
  XOR U4421 ( .A(n2144), .B(n2145), .Z(n2147) );
  XNOR U4422 ( .A(n2146), .B(n2147), .Z(n3178) );
  XOR U4423 ( .A(x[1051]), .B(y[1051]), .Z(n2566) );
  XOR U4424 ( .A(x[346]), .B(y[346]), .Z(n2564) );
  XNOR U4425 ( .A(x[1053]), .B(y[1053]), .Z(n2565) );
  XOR U4426 ( .A(n2564), .B(n2565), .Z(n2567) );
  XOR U4427 ( .A(n2566), .B(n2567), .Z(n3179) );
  XNOR U4428 ( .A(n3178), .B(n3179), .Z(n3181) );
  XOR U4429 ( .A(x[497]), .B(y[497]), .Z(n2158) );
  XOR U4430 ( .A(x[499]), .B(y[499]), .Z(n2156) );
  XNOR U4431 ( .A(x[501]), .B(y[501]), .Z(n2157) );
  XOR U4432 ( .A(n2156), .B(n2157), .Z(n2159) );
  XNOR U4433 ( .A(n2158), .B(n2159), .Z(n3180) );
  XNOR U4434 ( .A(n3181), .B(n3180), .Z(n4570) );
  XNOR U4435 ( .A(n4571), .B(n4570), .Z(n4572) );
  XNOR U4436 ( .A(n4573), .B(n4572), .Z(n2056) );
  XOR U4437 ( .A(n2057), .B(n2056), .Z(n2659) );
  XOR U4438 ( .A(x[561]), .B(y[561]), .Z(n2364) );
  XOR U4439 ( .A(x[384]), .B(y[384]), .Z(n2362) );
  XNOR U4440 ( .A(x[563]), .B(y[563]), .Z(n2363) );
  XOR U4441 ( .A(n2362), .B(n2363), .Z(n2365) );
  XNOR U4442 ( .A(n2364), .B(n2365), .Z(n3119) );
  XOR U4443 ( .A(x[565]), .B(y[565]), .Z(n2251) );
  XOR U4444 ( .A(x[567]), .B(y[567]), .Z(n2248) );
  XNOR U4445 ( .A(x[640]), .B(y[640]), .Z(n2249) );
  XNOR U4446 ( .A(n2248), .B(n2249), .Z(n2250) );
  XOR U4447 ( .A(n2251), .B(n2250), .Z(n3118) );
  XOR U4448 ( .A(n3119), .B(n3118), .Z(n3121) );
  XOR U4449 ( .A(x[569]), .B(y[569]), .Z(n2244) );
  XOR U4450 ( .A(x[376]), .B(y[376]), .Z(n2242) );
  XNOR U4451 ( .A(x[571]), .B(y[571]), .Z(n2243) );
  XOR U4452 ( .A(n2242), .B(n2243), .Z(n2245) );
  XNOR U4453 ( .A(n2244), .B(n2245), .Z(n3120) );
  XOR U4454 ( .A(n3121), .B(n3120), .Z(n2271) );
  XOR U4455 ( .A(x[585]), .B(y[585]), .Z(n2218) );
  XOR U4456 ( .A(x[593]), .B(y[593]), .Z(n2216) );
  XNOR U4457 ( .A(x[1478]), .B(y[1478]), .Z(n2217) );
  XOR U4458 ( .A(n2216), .B(n2217), .Z(n2219) );
  XNOR U4459 ( .A(n2218), .B(n2219), .Z(n2716) );
  XOR U4460 ( .A(x[601]), .B(y[601]), .Z(n2230) );
  XOR U4461 ( .A(x[603]), .B(y[603]), .Z(n2228) );
  XNOR U4462 ( .A(x[626]), .B(y[626]), .Z(n2229) );
  XOR U4463 ( .A(n2228), .B(n2229), .Z(n2231) );
  XOR U4464 ( .A(n2230), .B(n2231), .Z(n2717) );
  XNOR U4465 ( .A(n2716), .B(n2717), .Z(n2719) );
  XOR U4466 ( .A(x[605]), .B(y[605]), .Z(n2224) );
  XOR U4467 ( .A(x[356]), .B(y[356]), .Z(n2222) );
  XNOR U4468 ( .A(x[607]), .B(y[607]), .Z(n2223) );
  XOR U4469 ( .A(n2222), .B(n2223), .Z(n2225) );
  XNOR U4470 ( .A(n2224), .B(n2225), .Z(n2718) );
  XOR U4471 ( .A(n2719), .B(n2718), .Z(n2269) );
  XOR U4472 ( .A(x[573]), .B(y[573]), .Z(n2257) );
  XOR U4473 ( .A(x[372]), .B(y[372]), .Z(n2255) );
  XOR U4474 ( .A(x[575]), .B(y[575]), .Z(n2254) );
  XOR U4475 ( .A(n2255), .B(n2254), .Z(n2256) );
  XOR U4476 ( .A(n2257), .B(n2256), .Z(n2694) );
  XOR U4477 ( .A(x[577]), .B(y[577]), .Z(n2212) );
  XOR U4478 ( .A(x[579]), .B(y[579]), .Z(n2210) );
  XNOR U4479 ( .A(x[1476]), .B(y[1476]), .Z(n2211) );
  XOR U4480 ( .A(n2210), .B(n2211), .Z(n2213) );
  XOR U4481 ( .A(n2212), .B(n2213), .Z(n2695) );
  XNOR U4482 ( .A(n2694), .B(n2695), .Z(n2697) );
  XOR U4483 ( .A(x[581]), .B(y[581]), .Z(n2206) );
  XOR U4484 ( .A(x[364]), .B(y[364]), .Z(n2204) );
  XNOR U4485 ( .A(x[583]), .B(y[583]), .Z(n2205) );
  XOR U4486 ( .A(n2204), .B(n2205), .Z(n2207) );
  XNOR U4487 ( .A(n2206), .B(n2207), .Z(n2696) );
  XNOR U4488 ( .A(n2697), .B(n2696), .Z(n2268) );
  XNOR U4489 ( .A(n2269), .B(n2268), .Z(n2270) );
  XOR U4490 ( .A(n2271), .B(n2270), .Z(n1434) );
  XOR U4491 ( .A(x[503]), .B(y[503]), .Z(n1843) );
  XOR U4492 ( .A(x[505]), .B(y[505]), .Z(n1841) );
  XNOR U4493 ( .A(x[507]), .B(y[507]), .Z(n1842) );
  XOR U4494 ( .A(n1841), .B(n1842), .Z(n1844) );
  XNOR U4495 ( .A(n1843), .B(n1844), .Z(n3184) );
  XOR U4496 ( .A(x[1475]), .B(y[1475]), .Z(n4320) );
  XOR U4497 ( .A(x[80]), .B(y[80]), .Z(n4318) );
  XNOR U4498 ( .A(x[1477]), .B(y[1477]), .Z(n4319) );
  XOR U4499 ( .A(n4318), .B(n4319), .Z(n4321) );
  XOR U4500 ( .A(n4320), .B(n4321), .Z(n3185) );
  XNOR U4501 ( .A(n3184), .B(n3185), .Z(n3187) );
  XOR U4502 ( .A(x[509]), .B(y[509]), .Z(n1837) );
  XOR U4503 ( .A(x[50]), .B(y[50]), .Z(n1835) );
  XNOR U4504 ( .A(x[511]), .B(y[511]), .Z(n1836) );
  XOR U4505 ( .A(n1835), .B(n1836), .Z(n1838) );
  XNOR U4506 ( .A(n1837), .B(n1838), .Z(n3186) );
  XOR U4507 ( .A(n3187), .B(n3186), .Z(n4633) );
  XOR U4508 ( .A(x[513]), .B(y[513]), .Z(n1849) );
  XOR U4509 ( .A(x[515]), .B(y[515]), .Z(n1847) );
  XNOR U4510 ( .A(x[1468]), .B(y[1468]), .Z(n1848) );
  XOR U4511 ( .A(n1847), .B(n1848), .Z(n1850) );
  XNOR U4512 ( .A(n1849), .B(n1850), .Z(n3208) );
  XOR U4513 ( .A(x[1059]), .B(y[1059]), .Z(n2572) );
  XOR U4514 ( .A(x[340]), .B(y[340]), .Z(n2570) );
  XNOR U4515 ( .A(x[1061]), .B(y[1061]), .Z(n2571) );
  XOR U4516 ( .A(n2570), .B(n2571), .Z(n2573) );
  XOR U4517 ( .A(n2572), .B(n2573), .Z(n3209) );
  XNOR U4518 ( .A(n3208), .B(n3209), .Z(n3211) );
  XOR U4519 ( .A(x[517]), .B(y[517]), .Z(n5254) );
  XOR U4520 ( .A(x[418]), .B(y[418]), .Z(n5252) );
  XNOR U4521 ( .A(x[519]), .B(y[519]), .Z(n5253) );
  XOR U4522 ( .A(n5252), .B(n5253), .Z(n5255) );
  XNOR U4523 ( .A(n5254), .B(n5255), .Z(n3210) );
  XOR U4524 ( .A(n3211), .B(n3210), .Z(n4631) );
  XOR U4525 ( .A(x[521]), .B(y[521]), .Z(n5248) );
  XOR U4526 ( .A(x[523]), .B(y[523]), .Z(n5246) );
  XNOR U4527 ( .A(x[1470]), .B(y[1470]), .Z(n5247) );
  XOR U4528 ( .A(n5246), .B(n5247), .Z(n5249) );
  XNOR U4529 ( .A(n5248), .B(n5249), .Z(n3124) );
  XOR U4530 ( .A(x[1471]), .B(y[1471]), .Z(n4200) );
  XOR U4531 ( .A(x[305]), .B(y[305]), .Z(n4198) );
  XNOR U4532 ( .A(x[1473]), .B(y[1473]), .Z(n4199) );
  XOR U4533 ( .A(n4198), .B(n4199), .Z(n4201) );
  XOR U4534 ( .A(n4200), .B(n4201), .Z(n3125) );
  XNOR U4535 ( .A(n3124), .B(n3125), .Z(n3127) );
  XOR U4536 ( .A(x[525]), .B(y[525]), .Z(n5260) );
  XOR U4537 ( .A(x[527]), .B(y[527]), .Z(n5258) );
  XNOR U4538 ( .A(x[666]), .B(y[666]), .Z(n5259) );
  XOR U4539 ( .A(n5258), .B(n5259), .Z(n5261) );
  XNOR U4540 ( .A(n5260), .B(n5261), .Z(n3126) );
  XNOR U4541 ( .A(n3127), .B(n3126), .Z(n4630) );
  XNOR U4542 ( .A(n4631), .B(n4630), .Z(n4632) );
  XOR U4543 ( .A(n4633), .B(n4632), .Z(n1432) );
  XOR U4544 ( .A(x[529]), .B(y[529]), .Z(n5272) );
  XOR U4545 ( .A(x[412]), .B(y[412]), .Z(n5270) );
  XNOR U4546 ( .A(x[531]), .B(y[531]), .Z(n5271) );
  XOR U4547 ( .A(n5270), .B(n5271), .Z(n5273) );
  XNOR U4548 ( .A(n5272), .B(n5273), .Z(n3148) );
  XOR U4549 ( .A(x[1067]), .B(y[1067]), .Z(n2578) );
  XOR U4550 ( .A(x[29]), .B(y[29]), .Z(n2576) );
  XNOR U4551 ( .A(x[1069]), .B(y[1069]), .Z(n2577) );
  XOR U4552 ( .A(n2576), .B(n2577), .Z(n2579) );
  XOR U4553 ( .A(n2578), .B(n2579), .Z(n3149) );
  XNOR U4554 ( .A(n3148), .B(n3149), .Z(n3151) );
  XOR U4555 ( .A(x[533]), .B(y[533]), .Z(n5266) );
  XOR U4556 ( .A(x[535]), .B(y[535]), .Z(n5264) );
  XNOR U4557 ( .A(x[660]), .B(y[660]), .Z(n5265) );
  XOR U4558 ( .A(n5264), .B(n5265), .Z(n5267) );
  XNOR U4559 ( .A(n5266), .B(n5267), .Z(n3150) );
  XOR U4560 ( .A(n3151), .B(n3150), .Z(n4668) );
  XOR U4561 ( .A(x[537]), .B(y[537]), .Z(n5278) );
  XOR U4562 ( .A(x[404]), .B(y[404]), .Z(n5276) );
  XNOR U4563 ( .A(x[539]), .B(y[539]), .Z(n5277) );
  XOR U4564 ( .A(n5276), .B(n5277), .Z(n5279) );
  XNOR U4565 ( .A(n5278), .B(n5279), .Z(n2664) );
  XOR U4566 ( .A(x[541]), .B(y[541]), .Z(n2336) );
  XOR U4567 ( .A(x[398]), .B(y[398]), .Z(n2334) );
  XNOR U4568 ( .A(x[543]), .B(y[543]), .Z(n2335) );
  XOR U4569 ( .A(n2334), .B(n2335), .Z(n2337) );
  XOR U4570 ( .A(n2336), .B(n2337), .Z(n2665) );
  XNOR U4571 ( .A(n2664), .B(n2665), .Z(n2667) );
  XOR U4572 ( .A(x[545]), .B(y[545]), .Z(n2348) );
  XOR U4573 ( .A(x[547]), .B(y[547]), .Z(n2346) );
  XNOR U4574 ( .A(x[1472]), .B(y[1472]), .Z(n2347) );
  XOR U4575 ( .A(n2346), .B(n2347), .Z(n2349) );
  XNOR U4576 ( .A(n2348), .B(n2349), .Z(n2666) );
  XOR U4577 ( .A(n2667), .B(n2666), .Z(n4667) );
  XOR U4578 ( .A(x[549]), .B(y[549]), .Z(n2342) );
  XOR U4579 ( .A(x[392]), .B(y[392]), .Z(n2340) );
  XNOR U4580 ( .A(x[551]), .B(y[551]), .Z(n2341) );
  XOR U4581 ( .A(n2340), .B(n2341), .Z(n2343) );
  XNOR U4582 ( .A(n2342), .B(n2343), .Z(n2688) );
  XOR U4583 ( .A(x[553]), .B(y[553]), .Z(n2358) );
  XOR U4584 ( .A(x[555]), .B(y[555]), .Z(n2356) );
  XNOR U4585 ( .A(x[1474]), .B(y[1474]), .Z(n2357) );
  XOR U4586 ( .A(n2356), .B(n2357), .Z(n2359) );
  XOR U4587 ( .A(n2358), .B(n2359), .Z(n2689) );
  XNOR U4588 ( .A(n2688), .B(n2689), .Z(n2691) );
  XOR U4589 ( .A(x[557]), .B(y[557]), .Z(n2370) );
  XOR U4590 ( .A(x[559]), .B(y[559]), .Z(n2368) );
  XNOR U4591 ( .A(x[646]), .B(y[646]), .Z(n2369) );
  XOR U4592 ( .A(n2368), .B(n2369), .Z(n2371) );
  XNOR U4593 ( .A(n2370), .B(n2371), .Z(n2690) );
  XNOR U4594 ( .A(n2691), .B(n2690), .Z(n4666) );
  XOR U4595 ( .A(n4667), .B(n4666), .Z(n4669) );
  XNOR U4596 ( .A(n4668), .B(n4669), .Z(n1431) );
  XOR U4597 ( .A(n1432), .B(n1431), .Z(n1433) );
  XOR U4598 ( .A(n1434), .B(n1433), .Z(n2658) );
  XNOR U4599 ( .A(n2659), .B(n2658), .Z(n2660) );
  XOR U4600 ( .A(n2661), .B(n2660), .Z(n1348) );
  XOR U4601 ( .A(n1347), .B(n1348), .Z(n1350) );
  XOR U4602 ( .A(n1349), .B(n1350), .Z(n919) );
  XOR U4603 ( .A(x[717]), .B(y[717]), .Z(n3662) );
  XOR U4604 ( .A(x[719]), .B(y[719]), .Z(n3660) );
  XNOR U4605 ( .A(x[1492]), .B(y[1492]), .Z(n3661) );
  XOR U4606 ( .A(n3660), .B(n3661), .Z(n3663) );
  XNOR U4607 ( .A(n3662), .B(n3663), .Z(n3031) );
  XOR U4608 ( .A(x[721]), .B(y[721]), .Z(n3675) );
  XOR U4609 ( .A(x[254]), .B(y[254]), .Z(n3672) );
  XNOR U4610 ( .A(x[723]), .B(y[723]), .Z(n3673) );
  XNOR U4611 ( .A(n3672), .B(n3673), .Z(n3674) );
  XOR U4612 ( .A(n3675), .B(n3674), .Z(n3030) );
  XOR U4613 ( .A(n3031), .B(n3030), .Z(n3033) );
  XOR U4614 ( .A(x[725]), .B(y[725]), .Z(n3644) );
  XOR U4615 ( .A(x[727]), .B(y[727]), .Z(n3642) );
  XNOR U4616 ( .A(x[1494]), .B(y[1494]), .Z(n3643) );
  XOR U4617 ( .A(n3642), .B(n3643), .Z(n3645) );
  XNOR U4618 ( .A(n3644), .B(n3645), .Z(n3032) );
  XOR U4619 ( .A(n3033), .B(n3032), .Z(n5193) );
  XOR U4620 ( .A(x[729]), .B(y[729]), .Z(n3605) );
  XOR U4621 ( .A(x[546]), .B(y[546]), .Z(n3603) );
  XOR U4622 ( .A(x[731]), .B(y[731]), .Z(n3602) );
  XOR U4623 ( .A(n3603), .B(n3602), .Z(n3604) );
  XOR U4624 ( .A(n3605), .B(n3604), .Z(n3009) );
  XOR U4625 ( .A(x[733]), .B(y[733]), .Z(n3669) );
  XOR U4626 ( .A(x[248]), .B(y[248]), .Z(n3666) );
  XNOR U4627 ( .A(x[735]), .B(y[735]), .Z(n3667) );
  XNOR U4628 ( .A(n3666), .B(n3667), .Z(n3668) );
  XOR U4629 ( .A(n3669), .B(n3668), .Z(n3008) );
  XOR U4630 ( .A(n3009), .B(n3008), .Z(n3011) );
  XOR U4631 ( .A(x[737]), .B(y[737]), .Z(n950) );
  XOR U4632 ( .A(x[540]), .B(y[540]), .Z(n948) );
  XNOR U4633 ( .A(x[739]), .B(y[739]), .Z(n949) );
  XOR U4634 ( .A(n948), .B(n949), .Z(n951) );
  XNOR U4635 ( .A(n950), .B(n951), .Z(n3010) );
  XOR U4636 ( .A(n3011), .B(n3010), .Z(n5191) );
  XOR U4637 ( .A(x[741]), .B(y[741]), .Z(n1298) );
  XOR U4638 ( .A(x[238]), .B(y[238]), .Z(n1296) );
  XOR U4639 ( .A(x[743]), .B(y[743]), .Z(n1295) );
  XOR U4640 ( .A(n1296), .B(n1295), .Z(n1297) );
  XOR U4641 ( .A(n1298), .B(n1297), .Z(n4055) );
  XOR U4642 ( .A(x[745]), .B(y[745]), .Z(n3037) );
  XOR U4643 ( .A(x[234]), .B(y[234]), .Z(n3034) );
  XNOR U4644 ( .A(x[747]), .B(y[747]), .Z(n3035) );
  XNOR U4645 ( .A(n3034), .B(n3035), .Z(n3036) );
  XOR U4646 ( .A(n3037), .B(n3036), .Z(n4054) );
  XOR U4647 ( .A(n4055), .B(n4054), .Z(n4057) );
  XOR U4648 ( .A(x[749]), .B(y[749]), .Z(n4731) );
  XOR U4649 ( .A(x[751]), .B(y[751]), .Z(n4729) );
  XOR U4650 ( .A(x[1496]), .B(y[1496]), .Z(n4728) );
  XOR U4651 ( .A(n4729), .B(n4728), .Z(n4730) );
  XOR U4652 ( .A(n4731), .B(n4730), .Z(n4056) );
  XNOR U4653 ( .A(n4057), .B(n4056), .Z(n5190) );
  XNOR U4654 ( .A(n5191), .B(n5190), .Z(n5192) );
  XNOR U4655 ( .A(n5193), .B(n5192), .Z(n1065) );
  XOR U4656 ( .A(x[753]), .B(y[753]), .Z(n4176) );
  XOR U4657 ( .A(x[228]), .B(y[228]), .Z(n4174) );
  XNOR U4658 ( .A(x[755]), .B(y[755]), .Z(n4175) );
  XOR U4659 ( .A(n4174), .B(n4175), .Z(n4177) );
  XNOR U4660 ( .A(n4176), .B(n4177), .Z(n4033) );
  XOR U4661 ( .A(x[757]), .B(y[757]), .Z(n1580) );
  XOR U4662 ( .A(x[759]), .B(y[759]), .Z(n1578) );
  XOR U4663 ( .A(x[1498]), .B(y[1498]), .Z(n1577) );
  XOR U4664 ( .A(n1578), .B(n1577), .Z(n1579) );
  XOR U4665 ( .A(n1580), .B(n1579), .Z(n4032) );
  XOR U4666 ( .A(n4033), .B(n4032), .Z(n4035) );
  XOR U4667 ( .A(x[761]), .B(y[761]), .Z(n3571) );
  XOR U4668 ( .A(x[526]), .B(y[526]), .Z(n3569) );
  XOR U4669 ( .A(x[763]), .B(y[763]), .Z(n3568) );
  XOR U4670 ( .A(n3569), .B(n3568), .Z(n3570) );
  XOR U4671 ( .A(n3571), .B(n3570), .Z(n4034) );
  XOR U4672 ( .A(n4035), .B(n4034), .Z(n5205) );
  XOR U4673 ( .A(x[765]), .B(y[765]), .Z(n3372) );
  XOR U4674 ( .A(x[218]), .B(y[218]), .Z(n3370) );
  XNOR U4675 ( .A(x[767]), .B(y[767]), .Z(n3371) );
  XOR U4676 ( .A(n3370), .B(n3371), .Z(n3373) );
  XNOR U4677 ( .A(n3372), .B(n3373), .Z(n2815) );
  XOR U4678 ( .A(x[769]), .B(y[769]), .Z(n3367) );
  XOR U4679 ( .A(x[520]), .B(y[520]), .Z(n3364) );
  XNOR U4680 ( .A(x[771]), .B(y[771]), .Z(n3365) );
  XNOR U4681 ( .A(n3364), .B(n3365), .Z(n3366) );
  XOR U4682 ( .A(n3367), .B(n3366), .Z(n2814) );
  XOR U4683 ( .A(n2815), .B(n2814), .Z(n2817) );
  XOR U4684 ( .A(x[773]), .B(y[773]), .Z(n3525) );
  XOR U4685 ( .A(x[212]), .B(y[212]), .Z(n3523) );
  XOR U4686 ( .A(x[775]), .B(y[775]), .Z(n3522) );
  XOR U4687 ( .A(n3523), .B(n3522), .Z(n3524) );
  XOR U4688 ( .A(n3525), .B(n3524), .Z(n2816) );
  XOR U4689 ( .A(n2817), .B(n2816), .Z(n5203) );
  XOR U4690 ( .A(x[777]), .B(y[777]), .Z(n3565) );
  XOR U4691 ( .A(x[208]), .B(y[208]), .Z(n3563) );
  XOR U4692 ( .A(x[779]), .B(y[779]), .Z(n3562) );
  XOR U4693 ( .A(n3563), .B(n3562), .Z(n3564) );
  XOR U4694 ( .A(n3565), .B(n3564), .Z(n2723) );
  XOR U4695 ( .A(x[781]), .B(y[781]), .Z(n3421) );
  XOR U4696 ( .A(x[783]), .B(y[783]), .Z(n3419) );
  XOR U4697 ( .A(x[1500]), .B(y[1500]), .Z(n3418) );
  XOR U4698 ( .A(n3419), .B(n3418), .Z(n3420) );
  XOR U4699 ( .A(n3421), .B(n3420), .Z(n2722) );
  XOR U4700 ( .A(n2723), .B(n2722), .Z(n2725) );
  XOR U4701 ( .A(x[785]), .B(y[785]), .Z(n3425) );
  XOR U4702 ( .A(x[198]), .B(y[198]), .Z(n3423) );
  XOR U4703 ( .A(x[787]), .B(y[787]), .Z(n3422) );
  XOR U4704 ( .A(n3423), .B(n3422), .Z(n3424) );
  XOR U4705 ( .A(n3425), .B(n3424), .Z(n2724) );
  XNOR U4706 ( .A(n2725), .B(n2724), .Z(n5202) );
  XNOR U4707 ( .A(n5203), .B(n5202), .Z(n5204) );
  XOR U4708 ( .A(n5205), .B(n5204), .Z(n1066) );
  XNOR U4709 ( .A(n1065), .B(n1066), .Z(n1068) );
  XOR U4710 ( .A(x[791]), .B(y[791]), .Z(n4238) );
  XOR U4711 ( .A(x[793]), .B(y[793]), .Z(n4236) );
  XNOR U4712 ( .A(x[1502]), .B(y[1502]), .Z(n4237) );
  XOR U4713 ( .A(n4236), .B(n4237), .Z(n4239) );
  XNOR U4714 ( .A(n4238), .B(n4239), .Z(n3097) );
  XOR U4715 ( .A(x[795]), .B(y[795]), .Z(n2101) );
  XOR U4716 ( .A(x[506]), .B(y[506]), .Z(n2098) );
  XNOR U4717 ( .A(x[797]), .B(y[797]), .Z(n2099) );
  XNOR U4718 ( .A(n2098), .B(n2099), .Z(n2100) );
  XOR U4719 ( .A(n2101), .B(n2100), .Z(n3096) );
  XOR U4720 ( .A(n3097), .B(n3096), .Z(n3099) );
  XOR U4721 ( .A(x[799]), .B(y[799]), .Z(n4289) );
  XOR U4722 ( .A(x[192]), .B(y[192]), .Z(n4286) );
  XNOR U4723 ( .A(x[801]), .B(y[801]), .Z(n4287) );
  XNOR U4724 ( .A(n4286), .B(n4287), .Z(n4288) );
  XOR U4725 ( .A(n4289), .B(n4288), .Z(n3098) );
  XOR U4726 ( .A(n3099), .B(n3098), .Z(n3095) );
  XOR U4727 ( .A(x[803]), .B(y[803]), .Z(n4394) );
  XOR U4728 ( .A(x[500]), .B(y[500]), .Z(n4392) );
  XNOR U4729 ( .A(x[805]), .B(y[805]), .Z(n4393) );
  XOR U4730 ( .A(n4392), .B(n4393), .Z(n4395) );
  XNOR U4731 ( .A(n4394), .B(n4395), .Z(n3002) );
  XOR U4732 ( .A(x[807]), .B(y[807]), .Z(n4332) );
  XOR U4733 ( .A(x[184]), .B(y[184]), .Z(n4330) );
  XNOR U4734 ( .A(x[809]), .B(y[809]), .Z(n4331) );
  XOR U4735 ( .A(n4330), .B(n4331), .Z(n4333) );
  XOR U4736 ( .A(n4332), .B(n4333), .Z(n3003) );
  XNOR U4737 ( .A(n3002), .B(n3003), .Z(n3004) );
  XOR U4738 ( .A(x[815]), .B(y[815]), .Z(n1865) );
  XOR U4739 ( .A(x[817]), .B(y[817]), .Z(n1863) );
  XNOR U4740 ( .A(x[1504]), .B(y[1504]), .Z(n1864) );
  XOR U4741 ( .A(n1863), .B(n1864), .Z(n1866) );
  XOR U4742 ( .A(n1865), .B(n1866), .Z(n3005) );
  XOR U4743 ( .A(n3004), .B(n3005), .Z(n3092) );
  XOR U4744 ( .A(x[823]), .B(y[823]), .Z(n1513) );
  XOR U4745 ( .A(x[825]), .B(y[825]), .Z(n1511) );
  XNOR U4746 ( .A(x[1506]), .B(y[1506]), .Z(n1512) );
  XOR U4747 ( .A(n1511), .B(n1512), .Z(n1514) );
  XNOR U4748 ( .A(n1513), .B(n1514), .Z(n1915) );
  XOR U4749 ( .A(x[831]), .B(y[831]), .Z(n1368) );
  XOR U4750 ( .A(x[164]), .B(y[164]), .Z(n1365) );
  XNOR U4751 ( .A(x[833]), .B(y[833]), .Z(n1366) );
  XNOR U4752 ( .A(n1365), .B(n1366), .Z(n1367) );
  XOR U4753 ( .A(n1368), .B(n1367), .Z(n1914) );
  XOR U4754 ( .A(n1915), .B(n1914), .Z(n1917) );
  XOR U4755 ( .A(x[839]), .B(y[839]), .Z(n4502) );
  XOR U4756 ( .A(x[156]), .B(y[156]), .Z(n4500) );
  XNOR U4757 ( .A(x[841]), .B(y[841]), .Z(n4501) );
  XOR U4758 ( .A(n4500), .B(n4501), .Z(n4503) );
  XNOR U4759 ( .A(n4502), .B(n4503), .Z(n1916) );
  XNOR U4760 ( .A(n1917), .B(n1916), .Z(n3093) );
  XOR U4761 ( .A(n3092), .B(n3093), .Z(n3094) );
  XNOR U4762 ( .A(n3095), .B(n3094), .Z(n1067) );
  XOR U4763 ( .A(n1068), .B(n1067), .Z(n2312) );
  XOR U4764 ( .A(x[1403]), .B(y[1403]), .Z(n1725) );
  XOR U4765 ( .A(x[126]), .B(y[126]), .Z(n1723) );
  XNOR U4766 ( .A(x[1405]), .B(y[1405]), .Z(n1724) );
  XOR U4767 ( .A(n1723), .B(n1724), .Z(n1726) );
  XNOR U4768 ( .A(n1725), .B(n1726), .Z(n1635) );
  XOR U4769 ( .A(x[1391]), .B(y[1391]), .Z(n2006) );
  XOR U4770 ( .A(x[1393]), .B(y[1393]), .Z(n2004) );
  XNOR U4771 ( .A(x[1576]), .B(y[1576]), .Z(n2005) );
  XOR U4772 ( .A(n2004), .B(n2005), .Z(n2007) );
  XOR U4773 ( .A(n2006), .B(n2007), .Z(n1636) );
  XNOR U4774 ( .A(n1635), .B(n1636), .Z(n1638) );
  XOR U4775 ( .A(x[1375]), .B(y[1375]), .Z(n4917) );
  XOR U4776 ( .A(x[239]), .B(y[239]), .Z(n4915) );
  XOR U4777 ( .A(x[1377]), .B(y[1377]), .Z(n4914) );
  XOR U4778 ( .A(n4915), .B(n4914), .Z(n4916) );
  XOR U4779 ( .A(n4917), .B(n4916), .Z(n1637) );
  XOR U4780 ( .A(n1638), .B(n1637), .Z(n1913) );
  XOR U4781 ( .A(x[1383]), .B(y[1383]), .Z(n4156) );
  XOR U4782 ( .A(x[245]), .B(y[245]), .Z(n4154) );
  XNOR U4783 ( .A(x[1385]), .B(y[1385]), .Z(n4155) );
  XOR U4784 ( .A(n4154), .B(n4155), .Z(n4157) );
  XOR U4785 ( .A(n4156), .B(n4157), .Z(n1910) );
  XOR U4786 ( .A(x[1387]), .B(y[1387]), .Z(n4151) );
  XOR U4787 ( .A(x[249]), .B(y[249]), .Z(n4148) );
  XNOR U4788 ( .A(x[1389]), .B(y[1389]), .Z(n4149) );
  XNOR U4789 ( .A(n4148), .B(n4149), .Z(n4150) );
  XNOR U4790 ( .A(n4151), .B(n4150), .Z(n1911) );
  XOR U4791 ( .A(n1910), .B(n1911), .Z(n1912) );
  XOR U4792 ( .A(n1913), .B(n1912), .Z(n1136) );
  XOR U4793 ( .A(x[1343]), .B(y[1343]), .Z(n1862) );
  XOR U4794 ( .A(x[217]), .B(y[217]), .Z(n1860) );
  XOR U4795 ( .A(x[1345]), .B(y[1345]), .Z(n1859) );
  XOR U4796 ( .A(n1860), .B(n1859), .Z(n1861) );
  XOR U4797 ( .A(n1862), .B(n1861), .Z(n5051) );
  XOR U4798 ( .A(x[1351]), .B(y[1351]), .Z(n4929) );
  XOR U4799 ( .A(x[223]), .B(y[223]), .Z(n4927) );
  XOR U4800 ( .A(x[1353]), .B(y[1353]), .Z(n4926) );
  XOR U4801 ( .A(n4927), .B(n4926), .Z(n4928) );
  XOR U4802 ( .A(n4929), .B(n4928), .Z(n5050) );
  XOR U4803 ( .A(n5051), .B(n5050), .Z(n5053) );
  XOR U4804 ( .A(x[1347]), .B(y[1347]), .Z(n1886) );
  XOR U4805 ( .A(x[160]), .B(y[160]), .Z(n1884) );
  XOR U4806 ( .A(x[1349]), .B(y[1349]), .Z(n1883) );
  XOR U4807 ( .A(n1884), .B(n1883), .Z(n1885) );
  XOR U4808 ( .A(n1886), .B(n1885), .Z(n5052) );
  XOR U4809 ( .A(n5053), .B(n5052), .Z(n1134) );
  XOR U4810 ( .A(x[1335]), .B(y[1335]), .Z(n1996) );
  XOR U4811 ( .A(x[1337]), .B(y[1337]), .Z(n1994) );
  XNOR U4812 ( .A(x[1570]), .B(y[1570]), .Z(n1995) );
  XOR U4813 ( .A(n1994), .B(n1995), .Z(n1997) );
  XNOR U4814 ( .A(n1996), .B(n1997), .Z(n1991) );
  XOR U4815 ( .A(x[1367]), .B(y[1367]), .Z(n1890) );
  XOR U4816 ( .A(x[1369]), .B(y[1369]), .Z(n1888) );
  XOR U4817 ( .A(x[1574]), .B(y[1574]), .Z(n1887) );
  XOR U4818 ( .A(n1888), .B(n1887), .Z(n1889) );
  XOR U4819 ( .A(n1890), .B(n1889), .Z(n1990) );
  XOR U4820 ( .A(n1991), .B(n1990), .Z(n1992) );
  XOR U4821 ( .A(x[1415]), .B(y[1415]), .Z(n5040) );
  XOR U4822 ( .A(x[267]), .B(y[267]), .Z(n5038) );
  XNOR U4823 ( .A(x[1417]), .B(y[1417]), .Z(n5039) );
  XOR U4824 ( .A(n5038), .B(n5039), .Z(n5041) );
  XOR U4825 ( .A(n5040), .B(n5041), .Z(n1993) );
  XNOR U4826 ( .A(n1992), .B(n1993), .Z(n1133) );
  XOR U4827 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U4828 ( .A(n1136), .B(n1135), .Z(n1128) );
  XOR U4829 ( .A(x[991]), .B(y[991]), .Z(n4714) );
  XOR U4830 ( .A(x[28]), .B(y[28]), .Z(n4712) );
  XNOR U4831 ( .A(x[993]), .B(y[993]), .Z(n4713) );
  XOR U4832 ( .A(n4712), .B(n4713), .Z(n4715) );
  XNOR U4833 ( .A(n4714), .B(n4715), .Z(n1456) );
  XOR U4834 ( .A(x[999]), .B(y[999]), .Z(n2545) );
  XOR U4835 ( .A(x[18]), .B(y[18]), .Z(n2543) );
  XOR U4836 ( .A(x[1001]), .B(y[1001]), .Z(n2542) );
  XOR U4837 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U4838 ( .A(n2545), .B(n2544), .Z(n1455) );
  XOR U4839 ( .A(n1456), .B(n1455), .Z(n1458) );
  XOR U4840 ( .A(x[1007]), .B(y[1007]), .Z(n2541) );
  XOR U4841 ( .A(x[1009]), .B(y[1009]), .Z(n2539) );
  XOR U4842 ( .A(x[1528]), .B(y[1528]), .Z(n2538) );
  XOR U4843 ( .A(n2539), .B(n2538), .Z(n2540) );
  XOR U4844 ( .A(n2541), .B(n2540), .Z(n1457) );
  XOR U4845 ( .A(n1458), .B(n1457), .Z(n4065) );
  XOR U4846 ( .A(x[1015]), .B(y[1015]), .Z(n5001) );
  XOR U4847 ( .A(x[1017]), .B(y[1017]), .Z(n4999) );
  XOR U4848 ( .A(x[1530]), .B(y[1530]), .Z(n4998) );
  XOR U4849 ( .A(n4999), .B(n4998), .Z(n5000) );
  XOR U4850 ( .A(n5001), .B(n5000), .Z(n1530) );
  XOR U4851 ( .A(x[1023]), .B(y[1023]), .Z(n5007) );
  XOR U4852 ( .A(x[2]), .B(y[2]), .Z(n5005) );
  XOR U4853 ( .A(x[1025]), .B(y[1025]), .Z(n5004) );
  XOR U4854 ( .A(n5005), .B(n5004), .Z(n5006) );
  XOR U4855 ( .A(n5007), .B(n5006), .Z(n1529) );
  XOR U4856 ( .A(n1530), .B(n1529), .Z(n1531) );
  XOR U4857 ( .A(x[1031]), .B(y[1031]), .Z(n1073) );
  XOR U4858 ( .A(x[3]), .B(y[3]), .Z(n1071) );
  XNOR U4859 ( .A(x[1033]), .B(y[1033]), .Z(n1072) );
  XOR U4860 ( .A(n1071), .B(n1072), .Z(n1074) );
  XOR U4861 ( .A(n1073), .B(n1074), .Z(n1532) );
  XOR U4862 ( .A(n1531), .B(n1532), .Z(n4062) );
  XOR U4863 ( .A(x[1039]), .B(y[1039]), .Z(n1098) );
  XOR U4864 ( .A(x[1041]), .B(y[1041]), .Z(n1096) );
  XOR U4865 ( .A(x[1532]), .B(y[1532]), .Z(n1095) );
  XOR U4866 ( .A(n1096), .B(n1095), .Z(n1097) );
  XOR U4867 ( .A(n1098), .B(n1097), .Z(n1534) );
  XOR U4868 ( .A(x[1047]), .B(y[1047]), .Z(n1102) );
  XOR U4869 ( .A(x[1049]), .B(y[1049]), .Z(n1100) );
  XOR U4870 ( .A(x[1534]), .B(y[1534]), .Z(n1099) );
  XOR U4871 ( .A(n1100), .B(n1099), .Z(n1101) );
  XOR U4872 ( .A(n1102), .B(n1101), .Z(n1533) );
  XOR U4873 ( .A(n1534), .B(n1533), .Z(n1536) );
  XOR U4874 ( .A(x[1055]), .B(y[1055]), .Z(n2560) );
  XOR U4875 ( .A(x[19]), .B(y[19]), .Z(n2558) );
  XNOR U4876 ( .A(x[1057]), .B(y[1057]), .Z(n2559) );
  XOR U4877 ( .A(n2558), .B(n2559), .Z(n2561) );
  XNOR U4878 ( .A(n2560), .B(n2561), .Z(n1535) );
  XNOR U4879 ( .A(n1536), .B(n1535), .Z(n4063) );
  XOR U4880 ( .A(n4062), .B(n4063), .Z(n4064) );
  XNOR U4881 ( .A(n4065), .B(n4064), .Z(n1127) );
  XOR U4882 ( .A(n1128), .B(n1127), .Z(n1130) );
  XOR U4883 ( .A(x[1063]), .B(y[1063]), .Z(n2584) );
  XOR U4884 ( .A(x[25]), .B(y[25]), .Z(n2582) );
  XNOR U4885 ( .A(x[1065]), .B(y[1065]), .Z(n2583) );
  XOR U4886 ( .A(n2582), .B(n2583), .Z(n2585) );
  XNOR U4887 ( .A(n2584), .B(n2585), .Z(n1551) );
  XOR U4888 ( .A(x[1071]), .B(y[1071]), .Z(n2590) );
  XOR U4889 ( .A(x[1073]), .B(y[1073]), .Z(n2588) );
  XNOR U4890 ( .A(x[1536]), .B(y[1536]), .Z(n2589) );
  XOR U4891 ( .A(n2588), .B(n2589), .Z(n2591) );
  XOR U4892 ( .A(n2590), .B(n2591), .Z(n1552) );
  XNOR U4893 ( .A(n1551), .B(n1552), .Z(n1553) );
  XOR U4894 ( .A(x[1075]), .B(y[1075]), .Z(n1145) );
  XOR U4895 ( .A(x[35]), .B(y[35]), .Z(n1143) );
  XNOR U4896 ( .A(x[1077]), .B(y[1077]), .Z(n1144) );
  XOR U4897 ( .A(n1143), .B(n1144), .Z(n1146) );
  XOR U4898 ( .A(n1145), .B(n1146), .Z(n1554) );
  XOR U4899 ( .A(n1553), .B(n1554), .Z(n4060) );
  XOR U4900 ( .A(x[1079]), .B(y[1079]), .Z(n1139) );
  XOR U4901 ( .A(x[1081]), .B(y[1081]), .Z(n1137) );
  XNOR U4902 ( .A(x[1538]), .B(y[1538]), .Z(n1138) );
  XOR U4903 ( .A(n1137), .B(n1138), .Z(n1140) );
  XNOR U4904 ( .A(n1139), .B(n1140), .Z(n5170) );
  XOR U4905 ( .A(x[1083]), .B(y[1083]), .Z(n1151) );
  XOR U4906 ( .A(x[326]), .B(y[326]), .Z(n1149) );
  XNOR U4907 ( .A(x[1085]), .B(y[1085]), .Z(n1150) );
  XOR U4908 ( .A(n1149), .B(n1150), .Z(n1152) );
  XOR U4909 ( .A(n1151), .B(n1152), .Z(n5171) );
  XNOR U4910 ( .A(n5170), .B(n5171), .Z(n5173) );
  XOR U4911 ( .A(x[1087]), .B(y[1087]), .Z(n1162) );
  XOR U4912 ( .A(x[41]), .B(y[41]), .Z(n1160) );
  XOR U4913 ( .A(x[1089]), .B(y[1089]), .Z(n1159) );
  XOR U4914 ( .A(n1160), .B(n1159), .Z(n1161) );
  XOR U4915 ( .A(n1162), .B(n1161), .Z(n5172) );
  XOR U4916 ( .A(n5173), .B(n5172), .Z(n4059) );
  XOR U4917 ( .A(x[1091]), .B(y[1091]), .Z(n1158) );
  XOR U4918 ( .A(x[320]), .B(y[320]), .Z(n1156) );
  XOR U4919 ( .A(x[1093]), .B(y[1093]), .Z(n1155) );
  XOR U4920 ( .A(n1156), .B(n1155), .Z(n1157) );
  XOR U4921 ( .A(n1158), .B(n1157), .Z(n5164) );
  XOR U4922 ( .A(x[1095]), .B(y[1095]), .Z(n1175) );
  XOR U4923 ( .A(x[47]), .B(y[47]), .Z(n1173) );
  XNOR U4924 ( .A(x[1097]), .B(y[1097]), .Z(n1174) );
  XOR U4925 ( .A(n1173), .B(n1174), .Z(n1176) );
  XOR U4926 ( .A(n1175), .B(n1176), .Z(n5165) );
  XNOR U4927 ( .A(n5164), .B(n5165), .Z(n5167) );
  XOR U4928 ( .A(x[1099]), .B(y[1099]), .Z(n1187) );
  XOR U4929 ( .A(x[51]), .B(y[51]), .Z(n1185) );
  XNOR U4930 ( .A(x[1101]), .B(y[1101]), .Z(n1186) );
  XOR U4931 ( .A(n1185), .B(n1186), .Z(n1188) );
  XNOR U4932 ( .A(n1187), .B(n1188), .Z(n5166) );
  XNOR U4933 ( .A(n5167), .B(n5166), .Z(n4058) );
  XNOR U4934 ( .A(n4059), .B(n4058), .Z(n4061) );
  XOR U4935 ( .A(n4060), .B(n4061), .Z(n1129) );
  XOR U4936 ( .A(n1130), .B(n1129), .Z(n2311) );
  XOR U4937 ( .A(x[1291]), .B(y[1291]), .Z(n4139) );
  XOR U4938 ( .A(x[183]), .B(y[183]), .Z(n4137) );
  XOR U4939 ( .A(x[1293]), .B(y[1293]), .Z(n4136) );
  XOR U4940 ( .A(n4137), .B(n4136), .Z(n4138) );
  XOR U4941 ( .A(n4139), .B(n4138), .Z(n2496) );
  XOR U4942 ( .A(x[1439]), .B(y[1439]), .Z(n1197) );
  XOR U4943 ( .A(x[283]), .B(y[283]), .Z(n1195) );
  XNOR U4944 ( .A(x[1441]), .B(y[1441]), .Z(n1196) );
  XOR U4945 ( .A(n1195), .B(n1196), .Z(n1198) );
  XOR U4946 ( .A(n1197), .B(n1198), .Z(n2497) );
  XNOR U4947 ( .A(n2496), .B(n2497), .Z(n2499) );
  XOR U4948 ( .A(x[1295]), .B(y[1295]), .Z(n4143) );
  XOR U4949 ( .A(x[1297]), .B(y[1297]), .Z(n4141) );
  XOR U4950 ( .A(x[1564]), .B(y[1564]), .Z(n4140) );
  XOR U4951 ( .A(n4141), .B(n4140), .Z(n4142) );
  XOR U4952 ( .A(n4143), .B(n4142), .Z(n2498) );
  XOR U4953 ( .A(n2499), .B(n2498), .Z(n3947) );
  XOR U4954 ( .A(x[1299]), .B(y[1299]), .Z(n1651) );
  XOR U4955 ( .A(x[189]), .B(y[189]), .Z(n1649) );
  XNOR U4956 ( .A(x[1301]), .B(y[1301]), .Z(n1650) );
  XOR U4957 ( .A(n1649), .B(n1650), .Z(n1652) );
  XNOR U4958 ( .A(n1651), .B(n1652), .Z(n5010) );
  XOR U4959 ( .A(x[1435]), .B(y[1435]), .Z(n1203) );
  XOR U4960 ( .A(x[106]), .B(y[106]), .Z(n1201) );
  XNOR U4961 ( .A(x[1437]), .B(y[1437]), .Z(n1202) );
  XOR U4962 ( .A(n1201), .B(n1202), .Z(n1204) );
  XOR U4963 ( .A(n1203), .B(n1204), .Z(n5011) );
  XNOR U4964 ( .A(n5010), .B(n5011), .Z(n5013) );
  XOR U4965 ( .A(x[1303]), .B(y[1303]), .Z(n1657) );
  XOR U4966 ( .A(x[1305]), .B(y[1305]), .Z(n1655) );
  XNOR U4967 ( .A(x[1566]), .B(y[1566]), .Z(n1656) );
  XOR U4968 ( .A(n1655), .B(n1656), .Z(n1658) );
  XNOR U4969 ( .A(n1657), .B(n1658), .Z(n5012) );
  XOR U4970 ( .A(n5013), .B(n5012), .Z(n3945) );
  XOR U4971 ( .A(x[1307]), .B(y[1307]), .Z(n1669) );
  XOR U4972 ( .A(x[186]), .B(y[186]), .Z(n1667) );
  XNOR U4973 ( .A(x[1309]), .B(y[1309]), .Z(n1668) );
  XOR U4974 ( .A(n1667), .B(n1668), .Z(n1670) );
  XNOR U4975 ( .A(n1669), .B(n1670), .Z(n5054) );
  XOR U4976 ( .A(x[1431]), .B(y[1431]), .Z(n2508) );
  XOR U4977 ( .A(x[1433]), .B(y[1433]), .Z(n2506) );
  XNOR U4978 ( .A(x[1582]), .B(y[1582]), .Z(n2507) );
  XOR U4979 ( .A(n2506), .B(n2507), .Z(n2509) );
  XOR U4980 ( .A(n2508), .B(n2509), .Z(n5055) );
  XNOR U4981 ( .A(n5054), .B(n5055), .Z(n5057) );
  XOR U4982 ( .A(x[1311]), .B(y[1311]), .Z(n1663) );
  XOR U4983 ( .A(x[195]), .B(y[195]), .Z(n1661) );
  XNOR U4984 ( .A(x[1313]), .B(y[1313]), .Z(n1662) );
  XOR U4985 ( .A(n1661), .B(n1662), .Z(n1664) );
  XNOR U4986 ( .A(n1663), .B(n1664), .Z(n5056) );
  XNOR U4987 ( .A(n5057), .B(n5056), .Z(n3944) );
  XNOR U4988 ( .A(n3945), .B(n3944), .Z(n3946) );
  XNOR U4989 ( .A(n3947), .B(n3946), .Z(n2380) );
  XOR U4990 ( .A(x[1183]), .B(y[1183]), .Z(n3518) );
  XOR U4991 ( .A(x[107]), .B(y[107]), .Z(n3516) );
  XNOR U4992 ( .A(x[1185]), .B(y[1185]), .Z(n3517) );
  XOR U4993 ( .A(n3516), .B(n3517), .Z(n3519) );
  XNOR U4994 ( .A(n3518), .B(n3519), .Z(n2295) );
  XOR U4995 ( .A(x[1175]), .B(y[1175]), .Z(n2476) );
  XOR U4996 ( .A(x[1177]), .B(y[1177]), .Z(n2474) );
  XNOR U4997 ( .A(x[1550]), .B(y[1550]), .Z(n2475) );
  XOR U4998 ( .A(n2474), .B(n2475), .Z(n2477) );
  XNOR U4999 ( .A(n2476), .B(n2477), .Z(n2292) );
  XOR U5000 ( .A(x[1179]), .B(y[1179]), .Z(n2470) );
  XOR U5001 ( .A(x[266]), .B(y[266]), .Z(n2468) );
  XNOR U5002 ( .A(x[1181]), .B(y[1181]), .Z(n2469) );
  XOR U5003 ( .A(n2468), .B(n2469), .Z(n2471) );
  XOR U5004 ( .A(n2470), .B(n2471), .Z(n2293) );
  XNOR U5005 ( .A(n2292), .B(n2293), .Z(n2294) );
  XOR U5006 ( .A(n2295), .B(n2294), .Z(n3687) );
  XOR U5007 ( .A(x[1195]), .B(y[1195]), .Z(n3442) );
  XOR U5008 ( .A(x[117]), .B(y[117]), .Z(n3441) );
  XOR U5009 ( .A(x[1197]), .B(y[1197]), .Z(n3440) );
  XOR U5010 ( .A(n3441), .B(n3440), .Z(n3443) );
  XOR U5011 ( .A(n3442), .B(n3443), .Z(n2241) );
  XOR U5012 ( .A(x[1187]), .B(y[1187]), .Z(n2419) );
  XOR U5013 ( .A(x[260]), .B(y[260]), .Z(n2417) );
  XOR U5014 ( .A(x[1189]), .B(y[1189]), .Z(n2416) );
  XOR U5015 ( .A(n2417), .B(n2416), .Z(n2418) );
  XOR U5016 ( .A(n2419), .B(n2418), .Z(n2239) );
  XOR U5017 ( .A(x[1191]), .B(y[1191]), .Z(n3448) );
  XOR U5018 ( .A(x[113]), .B(y[113]), .Z(n3447) );
  XOR U5019 ( .A(x[1193]), .B(y[1193]), .Z(n3446) );
  XOR U5020 ( .A(n3447), .B(n3446), .Z(n3449) );
  XOR U5021 ( .A(n3448), .B(n3449), .Z(n2238) );
  XOR U5022 ( .A(n2239), .B(n2238), .Z(n2240) );
  XOR U5023 ( .A(n2241), .B(n2240), .Z(n3685) );
  XOR U5024 ( .A(x[1207]), .B(y[1207]), .Z(n3728) );
  XOR U5025 ( .A(x[1209]), .B(y[1209]), .Z(n3726) );
  XNOR U5026 ( .A(x[1554]), .B(y[1554]), .Z(n3727) );
  XOR U5027 ( .A(n3726), .B(n3727), .Z(n3729) );
  XNOR U5028 ( .A(n3728), .B(n3729), .Z(n1786) );
  XOR U5029 ( .A(x[1199]), .B(y[1199]), .Z(n2422) );
  XOR U5030 ( .A(x[1201]), .B(y[1201]), .Z(n2420) );
  XNOR U5031 ( .A(x[1552]), .B(y[1552]), .Z(n2421) );
  XOR U5032 ( .A(n2420), .B(n2421), .Z(n2423) );
  XNOR U5033 ( .A(n2422), .B(n2423), .Z(n1783) );
  XOR U5034 ( .A(x[1203]), .B(y[1203]), .Z(n1301) );
  XOR U5035 ( .A(x[123]), .B(y[123]), .Z(n1299) );
  XNOR U5036 ( .A(x[1205]), .B(y[1205]), .Z(n1300) );
  XOR U5037 ( .A(n1299), .B(n1300), .Z(n1302) );
  XOR U5038 ( .A(n1301), .B(n1302), .Z(n1784) );
  XNOR U5039 ( .A(n1783), .B(n1784), .Z(n1785) );
  XNOR U5040 ( .A(n1786), .B(n1785), .Z(n3684) );
  XNOR U5041 ( .A(n3685), .B(n3684), .Z(n3686) );
  XOR U5042 ( .A(n3687), .B(n3686), .Z(n2381) );
  XNOR U5043 ( .A(n2380), .B(n2381), .Z(n2383) );
  XOR U5044 ( .A(x[1211]), .B(y[1211]), .Z(n3784) );
  XOR U5045 ( .A(x[246]), .B(y[246]), .Z(n3782) );
  XNOR U5046 ( .A(x[1213]), .B(y[1213]), .Z(n3783) );
  XOR U5047 ( .A(n3782), .B(n3783), .Z(n3785) );
  XNOR U5048 ( .A(n3784), .B(n3785), .Z(n2105) );
  XOR U5049 ( .A(x[1215]), .B(y[1215]), .Z(n3879) );
  XOR U5050 ( .A(x[129]), .B(y[129]), .Z(n3876) );
  XNOR U5051 ( .A(x[1217]), .B(y[1217]), .Z(n3877) );
  XNOR U5052 ( .A(n3876), .B(n3877), .Z(n3878) );
  XOR U5053 ( .A(n3879), .B(n3878), .Z(n2104) );
  XOR U5054 ( .A(n2105), .B(n2104), .Z(n2107) );
  XOR U5055 ( .A(x[1219]), .B(y[1219]), .Z(n4406) );
  XOR U5056 ( .A(x[240]), .B(y[240]), .Z(n4404) );
  XNOR U5057 ( .A(x[1221]), .B(y[1221]), .Z(n4405) );
  XOR U5058 ( .A(n4404), .B(n4405), .Z(n4407) );
  XNOR U5059 ( .A(n4406), .B(n4407), .Z(n2106) );
  XOR U5060 ( .A(n2107), .B(n2106), .Z(n2389) );
  XOR U5061 ( .A(x[1223]), .B(y[1223]), .Z(n4400) );
  XOR U5062 ( .A(x[135]), .B(y[135]), .Z(n4398) );
  XNOR U5063 ( .A(x[1225]), .B(y[1225]), .Z(n4399) );
  XOR U5064 ( .A(n4398), .B(n4399), .Z(n4401) );
  XNOR U5065 ( .A(n4400), .B(n4401), .Z(n4899) );
  XOR U5066 ( .A(x[1227]), .B(y[1227]), .Z(n4779) );
  XOR U5067 ( .A(x[139]), .B(y[139]), .Z(n4777) );
  XOR U5068 ( .A(x[1229]), .B(y[1229]), .Z(n4776) );
  XOR U5069 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U5070 ( .A(n4779), .B(n4778), .Z(n4898) );
  XOR U5071 ( .A(n4899), .B(n4898), .Z(n4901) );
  XOR U5072 ( .A(x[1231]), .B(y[1231]), .Z(n5067) );
  XOR U5073 ( .A(x[1233]), .B(y[1233]), .Z(n5065) );
  XOR U5074 ( .A(x[1556]), .B(y[1556]), .Z(n5064) );
  XOR U5075 ( .A(n5065), .B(n5064), .Z(n5066) );
  XOR U5076 ( .A(n5067), .B(n5066), .Z(n4900) );
  XOR U5077 ( .A(n4901), .B(n4900), .Z(n2387) );
  XOR U5078 ( .A(x[1235]), .B(y[1235]), .Z(n5071) );
  XOR U5079 ( .A(x[145]), .B(y[145]), .Z(n5069) );
  XOR U5080 ( .A(x[1237]), .B(y[1237]), .Z(n5068) );
  XOR U5081 ( .A(n5069), .B(n5068), .Z(n5070) );
  XOR U5082 ( .A(n5071), .B(n5070), .Z(n2051) );
  XOR U5083 ( .A(x[1467]), .B(y[1467]), .Z(n2975) );
  XOR U5084 ( .A(x[86]), .B(y[86]), .Z(n2972) );
  XNOR U5085 ( .A(x[1469]), .B(y[1469]), .Z(n2973) );
  XNOR U5086 ( .A(n2972), .B(n2973), .Z(n2974) );
  XOR U5087 ( .A(n2975), .B(n2974), .Z(n2050) );
  XOR U5088 ( .A(n2051), .B(n2050), .Z(n2053) );
  XOR U5089 ( .A(x[1239]), .B(y[1239]), .Z(n4795) );
  XOR U5090 ( .A(x[1241]), .B(y[1241]), .Z(n4793) );
  XOR U5091 ( .A(x[1558]), .B(y[1558]), .Z(n4792) );
  XOR U5092 ( .A(n4793), .B(n4792), .Z(n4794) );
  XOR U5093 ( .A(n4795), .B(n4794), .Z(n2052) );
  XNOR U5094 ( .A(n2053), .B(n2052), .Z(n2386) );
  XNOR U5095 ( .A(n2387), .B(n2386), .Z(n2388) );
  XNOR U5096 ( .A(n2389), .B(n2388), .Z(n2382) );
  XNOR U5097 ( .A(n2383), .B(n2382), .Z(n2310) );
  XOR U5098 ( .A(n2311), .B(n2310), .Z(n2313) );
  XNOR U5099 ( .A(n2312), .B(n2313), .Z(n918) );
  XNOR U5100 ( .A(n919), .B(n918), .Z(n921) );
  XOR U5101 ( .A(x[424]), .B(y[424]), .Z(n4466) );
  XOR U5102 ( .A(x[416]), .B(y[416]), .Z(n4464) );
  XNOR U5103 ( .A(x[422]), .B(y[422]), .Z(n4465) );
  XOR U5104 ( .A(n4464), .B(n4465), .Z(n4467) );
  XNOR U5105 ( .A(n4466), .B(n4467), .Z(n4697) );
  XOR U5106 ( .A(x[875]), .B(y[875]), .Z(n2035) );
  XOR U5107 ( .A(x[124]), .B(y[124]), .Z(n2032) );
  XNOR U5108 ( .A(x[877]), .B(y[877]), .Z(n2033) );
  XNOR U5109 ( .A(n2032), .B(n2033), .Z(n2034) );
  XOR U5110 ( .A(n2035), .B(n2034), .Z(n4696) );
  XOR U5111 ( .A(n4697), .B(n4696), .Z(n4699) );
  XOR U5112 ( .A(x[414]), .B(y[414]), .Z(n2956) );
  XOR U5113 ( .A(x[410]), .B(y[410]), .Z(n2954) );
  XNOR U5114 ( .A(x[768]), .B(y[768]), .Z(n2955) );
  XOR U5115 ( .A(n2954), .B(n2955), .Z(n2957) );
  XNOR U5116 ( .A(n2956), .B(n2957), .Z(n4698) );
  XOR U5117 ( .A(n4699), .B(n4698), .Z(n1570) );
  XOR U5118 ( .A(x[408]), .B(y[408]), .Z(n4830) );
  XOR U5119 ( .A(x[396]), .B(y[396]), .Z(n4828) );
  XNOR U5120 ( .A(x[764]), .B(y[764]), .Z(n4829) );
  XOR U5121 ( .A(n4828), .B(n4829), .Z(n4831) );
  XNOR U5122 ( .A(n4830), .B(n4831), .Z(n4847) );
  XOR U5123 ( .A(x[1563]), .B(y[1563]), .Z(n4087) );
  XOR U5124 ( .A(x[26]), .B(y[26]), .Z(n4085) );
  XOR U5125 ( .A(x[1565]), .B(y[1565]), .Z(n4084) );
  XOR U5126 ( .A(n4085), .B(n4084), .Z(n4086) );
  XOR U5127 ( .A(n4087), .B(n4086), .Z(n4846) );
  XOR U5128 ( .A(n4847), .B(n4846), .Z(n4849) );
  XOR U5129 ( .A(x[378]), .B(y[378]), .Z(n4683) );
  XOR U5130 ( .A(x[370]), .B(y[370]), .Z(n4681) );
  XOR U5131 ( .A(x[374]), .B(y[374]), .Z(n4680) );
  XOR U5132 ( .A(n4681), .B(n4680), .Z(n4682) );
  XOR U5133 ( .A(n4683), .B(n4682), .Z(n4848) );
  XOR U5134 ( .A(n4849), .B(n4848), .Z(n1568) );
  XOR U5135 ( .A(x[352]), .B(y[352]), .Z(n2906) );
  XOR U5136 ( .A(x[348]), .B(y[348]), .Z(n2904) );
  XNOR U5137 ( .A(x[746]), .B(y[746]), .Z(n2905) );
  XOR U5138 ( .A(n2904), .B(n2905), .Z(n2907) );
  XNOR U5139 ( .A(n2906), .B(n2907), .Z(n4980) );
  XOR U5140 ( .A(x[883]), .B(y[883]), .Z(n2046) );
  XOR U5141 ( .A(x[116]), .B(y[116]), .Z(n2044) );
  XNOR U5142 ( .A(x[885]), .B(y[885]), .Z(n2045) );
  XOR U5143 ( .A(n2044), .B(n2045), .Z(n2047) );
  XOR U5144 ( .A(n2046), .B(n2047), .Z(n4981) );
  XNOR U5145 ( .A(n4980), .B(n4981), .Z(n4983) );
  XOR U5146 ( .A(x[342]), .B(y[342]), .Z(n4752) );
  XOR U5147 ( .A(x[334]), .B(y[334]), .Z(n4750) );
  XNOR U5148 ( .A(x[338]), .B(y[338]), .Z(n4751) );
  XOR U5149 ( .A(n4750), .B(n4751), .Z(n4753) );
  XNOR U5150 ( .A(n4752), .B(n4753), .Z(n4982) );
  XNOR U5151 ( .A(n4983), .B(n4982), .Z(n1567) );
  XNOR U5152 ( .A(n1568), .B(n1567), .Z(n1569) );
  XNOR U5153 ( .A(n1570), .B(n1569), .Z(n2316) );
  XOR U5154 ( .A(x[328]), .B(y[328]), .Z(n4759) );
  XOR U5155 ( .A(x[314]), .B(y[314]), .Z(n4757) );
  XOR U5156 ( .A(x[318]), .B(y[318]), .Z(n4756) );
  XOR U5157 ( .A(n4757), .B(n4756), .Z(n4758) );
  XOR U5158 ( .A(n4759), .B(n4758), .Z(n5101) );
  XOR U5159 ( .A(x[1559]), .B(y[1559]), .Z(n3055) );
  XOR U5160 ( .A(x[1561]), .B(y[1561]), .Z(n3052) );
  XNOR U5161 ( .A(x[1598]), .B(y[1598]), .Z(n3053) );
  XNOR U5162 ( .A(n3052), .B(n3053), .Z(n3054) );
  XOR U5163 ( .A(n3055), .B(n3054), .Z(n5100) );
  XOR U5164 ( .A(n5101), .B(n5100), .Z(n5103) );
  XOR U5165 ( .A(x[312]), .B(y[312]), .Z(n4419) );
  XOR U5166 ( .A(x[308]), .B(y[308]), .Z(n4417) );
  XOR U5167 ( .A(x[732]), .B(y[732]), .Z(n4416) );
  XOR U5168 ( .A(n4417), .B(n4416), .Z(n4418) );
  XOR U5169 ( .A(n4419), .B(n4418), .Z(n5102) );
  XOR U5170 ( .A(n5103), .B(n5102), .Z(n5199) );
  XOR U5171 ( .A(x[304]), .B(y[304]), .Z(n4423) );
  XOR U5172 ( .A(x[298]), .B(y[298]), .Z(n4421) );
  XOR U5173 ( .A(x[728]), .B(y[728]), .Z(n4420) );
  XOR U5174 ( .A(n4421), .B(n4420), .Z(n4422) );
  XOR U5175 ( .A(n4423), .B(n4422), .Z(n1987) );
  XOR U5176 ( .A(x[891]), .B(y[891]), .Z(n1688) );
  XOR U5177 ( .A(x[446]), .B(y[446]), .Z(n1685) );
  XNOR U5178 ( .A(x[893]), .B(y[893]), .Z(n1686) );
  XNOR U5179 ( .A(n1685), .B(n1686), .Z(n1687) );
  XOR U5180 ( .A(n1688), .B(n1687), .Z(n1986) );
  XOR U5181 ( .A(n1987), .B(n1986), .Z(n1989) );
  XOR U5182 ( .A(x[292]), .B(y[292]), .Z(n3503) );
  XOR U5183 ( .A(x[278]), .B(y[278]), .Z(n3501) );
  XOR U5184 ( .A(x[284]), .B(y[284]), .Z(n3500) );
  XOR U5185 ( .A(n3501), .B(n3500), .Z(n3502) );
  XOR U5186 ( .A(n3503), .B(n3502), .Z(n1988) );
  XOR U5187 ( .A(n1989), .B(n1988), .Z(n5197) );
  XOR U5188 ( .A(x[264]), .B(y[264]), .Z(n3589) );
  XOR U5189 ( .A(x[256]), .B(y[256]), .Z(n3587) );
  XOR U5190 ( .A(x[714]), .B(y[714]), .Z(n3586) );
  XOR U5191 ( .A(n3587), .B(n3586), .Z(n3588) );
  XOR U5192 ( .A(n3589), .B(n3588), .Z(n2073) );
  XOR U5193 ( .A(x[1555]), .B(y[1555]), .Z(n4219) );
  XOR U5194 ( .A(x[365]), .B(y[365]), .Z(n4217) );
  XOR U5195 ( .A(x[1557]), .B(y[1557]), .Z(n4216) );
  XOR U5196 ( .A(n4217), .B(n4216), .Z(n4218) );
  XOR U5197 ( .A(n4219), .B(n4218), .Z(n2072) );
  XOR U5198 ( .A(n2073), .B(n2072), .Z(n2075) );
  XOR U5199 ( .A(x[242]), .B(y[242]), .Z(n4315) );
  XOR U5200 ( .A(x[232]), .B(y[232]), .Z(n4313) );
  XOR U5201 ( .A(x[236]), .B(y[236]), .Z(n4312) );
  XOR U5202 ( .A(n4313), .B(n4312), .Z(n4314) );
  XOR U5203 ( .A(n4315), .B(n4314), .Z(n2074) );
  XNOR U5204 ( .A(n2075), .B(n2074), .Z(n5196) );
  XNOR U5205 ( .A(n5197), .B(n5196), .Z(n5198) );
  XOR U5206 ( .A(n5199), .B(n5198), .Z(n2317) );
  XNOR U5207 ( .A(n2316), .B(n2317), .Z(n2319) );
  XOR U5208 ( .A(x[230]), .B(y[230]), .Z(n4326) );
  XOR U5209 ( .A(x[214]), .B(y[214]), .Z(n4324) );
  XNOR U5210 ( .A(x[222]), .B(y[222]), .Z(n4325) );
  XOR U5211 ( .A(n4324), .B(n4325), .Z(n4327) );
  XNOR U5212 ( .A(n4326), .B(n4327), .Z(n5240) );
  XOR U5213 ( .A(x[899]), .B(y[899]), .Z(n1681) );
  XOR U5214 ( .A(x[440]), .B(y[440]), .Z(n1679) );
  XNOR U5215 ( .A(x[901]), .B(y[901]), .Z(n1680) );
  XOR U5216 ( .A(n1679), .B(n1680), .Z(n1682) );
  XOR U5217 ( .A(n1681), .B(n1682), .Z(n5241) );
  XNOR U5218 ( .A(n5240), .B(n5241), .Z(n5243) );
  XOR U5219 ( .A(x[210]), .B(y[210]), .Z(n4276) );
  XOR U5220 ( .A(x[204]), .B(y[204]), .Z(n4274) );
  XNOR U5221 ( .A(x[696]), .B(y[696]), .Z(n4275) );
  XOR U5222 ( .A(n4274), .B(n4275), .Z(n4277) );
  XNOR U5223 ( .A(n4276), .B(n4277), .Z(n5242) );
  XOR U5224 ( .A(n5243), .B(n5242), .Z(n2307) );
  XOR U5225 ( .A(x[202]), .B(y[202]), .Z(n4282) );
  XOR U5226 ( .A(x[196]), .B(y[196]), .Z(n4280) );
  XNOR U5227 ( .A(x[692]), .B(y[692]), .Z(n4281) );
  XOR U5228 ( .A(n4280), .B(n4281), .Z(n4283) );
  XNOR U5229 ( .A(n4282), .B(n4283), .Z(n4874) );
  XOR U5230 ( .A(x[1551]), .B(y[1551]), .Z(n4256) );
  XOR U5231 ( .A(x[1553]), .B(y[1553]), .Z(n4254) );
  XNOR U5232 ( .A(x[1596]), .B(y[1596]), .Z(n4255) );
  XOR U5233 ( .A(n4254), .B(n4255), .Z(n4257) );
  XOR U5234 ( .A(n4256), .B(n4257), .Z(n4875) );
  XNOR U5235 ( .A(n4874), .B(n4875), .Z(n4877) );
  XOR U5236 ( .A(x[194]), .B(y[194]), .Z(n4206) );
  XOR U5237 ( .A(x[176]), .B(y[176]), .Z(n4204) );
  XNOR U5238 ( .A(x[188]), .B(y[188]), .Z(n4205) );
  XOR U5239 ( .A(n4204), .B(n4205), .Z(n4207) );
  XNOR U5240 ( .A(n4206), .B(n4207), .Z(n4876) );
  XOR U5241 ( .A(n4877), .B(n4876), .Z(n2305) );
  XOR U5242 ( .A(x[174]), .B(y[174]), .Z(n3547) );
  XOR U5243 ( .A(x[168]), .B(y[168]), .Z(n3545) );
  XOR U5244 ( .A(x[170]), .B(y[170]), .Z(n3544) );
  XOR U5245 ( .A(n3545), .B(n3544), .Z(n3546) );
  XOR U5246 ( .A(n3547), .B(n3546), .Z(n1811) );
  XOR U5247 ( .A(x[907]), .B(y[907]), .Z(n1693) );
  XOR U5248 ( .A(x[96]), .B(y[96]), .Z(n1691) );
  XNOR U5249 ( .A(x[909]), .B(y[909]), .Z(n1692) );
  XOR U5250 ( .A(n1691), .B(n1692), .Z(n1694) );
  XOR U5251 ( .A(n1693), .B(n1694), .Z(n1812) );
  XNOR U5252 ( .A(n1811), .B(n1812), .Z(n1814) );
  XOR U5253 ( .A(x[150]), .B(y[150]), .Z(n3454) );
  XOR U5254 ( .A(x[142]), .B(y[142]), .Z(n3452) );
  XNOR U5255 ( .A(x[674]), .B(y[674]), .Z(n3453) );
  XOR U5256 ( .A(n3452), .B(n3453), .Z(n3455) );
  XNOR U5257 ( .A(n3454), .B(n3455), .Z(n1813) );
  XNOR U5258 ( .A(n1814), .B(n1813), .Z(n2304) );
  XNOR U5259 ( .A(n2305), .B(n2304), .Z(n2306) );
  XNOR U5260 ( .A(n2307), .B(n2306), .Z(n2318) );
  XOR U5261 ( .A(n2319), .B(n2318), .Z(n2493) );
  XOR U5262 ( .A(x[128]), .B(y[128]), .Z(n3001) );
  XOR U5263 ( .A(x[114]), .B(y[114]), .Z(n2999) );
  XOR U5264 ( .A(x[122]), .B(y[122]), .Z(n2998) );
  XOR U5265 ( .A(n2999), .B(n2998), .Z(n3000) );
  XOR U5266 ( .A(n3001), .B(n3000), .Z(n5159) );
  XOR U5267 ( .A(x[1547]), .B(y[1547]), .Z(n4303) );
  XOR U5268 ( .A(x[359]), .B(y[359]), .Z(n4301) );
  XOR U5269 ( .A(x[1549]), .B(y[1549]), .Z(n4300) );
  XOR U5270 ( .A(n4301), .B(n4300), .Z(n4302) );
  XOR U5271 ( .A(n4303), .B(n4302), .Z(n5158) );
  XOR U5272 ( .A(n5159), .B(n5158), .Z(n5161) );
  XOR U5273 ( .A(x[108]), .B(y[108]), .Z(n2980) );
  XOR U5274 ( .A(x[104]), .B(y[104]), .Z(n2978) );
  XNOR U5275 ( .A(x[656]), .B(y[656]), .Z(n2979) );
  XOR U5276 ( .A(n2978), .B(n2979), .Z(n2981) );
  XNOR U5277 ( .A(n2980), .B(n2981), .Z(n5160) );
  XOR U5278 ( .A(n5161), .B(n5160), .Z(n2165) );
  XOR U5279 ( .A(x[98]), .B(y[98]), .Z(n2986) );
  XOR U5280 ( .A(x[94]), .B(y[94]), .Z(n2984) );
  XNOR U5281 ( .A(x[652]), .B(y[652]), .Z(n2985) );
  XOR U5282 ( .A(n2984), .B(n2985), .Z(n2987) );
  XNOR U5283 ( .A(n2986), .B(n2987), .Z(n4821) );
  XOR U5284 ( .A(x[915]), .B(y[915]), .Z(n1704) );
  XOR U5285 ( .A(x[90]), .B(y[90]), .Z(n1701) );
  XNOR U5286 ( .A(x[917]), .B(y[917]), .Z(n1702) );
  XNOR U5287 ( .A(n1701), .B(n1702), .Z(n1703) );
  XOR U5288 ( .A(n1704), .B(n1703), .Z(n4820) );
  XOR U5289 ( .A(n4821), .B(n4820), .Z(n4823) );
  XOR U5290 ( .A(x[92]), .B(y[92]), .Z(n3078) );
  XOR U5291 ( .A(x[78]), .B(y[78]), .Z(n3076) );
  XNOR U5292 ( .A(x[88]), .B(y[88]), .Z(n3077) );
  XOR U5293 ( .A(n3076), .B(n3077), .Z(n3079) );
  XNOR U5294 ( .A(n3078), .B(n3079), .Z(n4822) );
  XOR U5295 ( .A(n4823), .B(n4822), .Z(n2163) );
  XOR U5296 ( .A(x[72]), .B(y[72]), .Z(n3084) );
  XOR U5297 ( .A(x[64]), .B(y[64]), .Z(n3082) );
  XNOR U5298 ( .A(x[68]), .B(y[68]), .Z(n3083) );
  XOR U5299 ( .A(n3082), .B(n3083), .Z(n3085) );
  XNOR U5300 ( .A(n3084), .B(n3085), .Z(n4813) );
  XOR U5301 ( .A(x[1543]), .B(y[1543]), .Z(n4347) );
  XOR U5302 ( .A(x[355]), .B(y[355]), .Z(n4344) );
  XNOR U5303 ( .A(x[1545]), .B(y[1545]), .Z(n4345) );
  XNOR U5304 ( .A(n4344), .B(n4345), .Z(n4346) );
  XOR U5305 ( .A(n4347), .B(n4346), .Z(n4812) );
  XOR U5306 ( .A(n4813), .B(n4812), .Z(n4815) );
  XOR U5307 ( .A(x[58]), .B(y[58]), .Z(n2394) );
  XOR U5308 ( .A(x[56]), .B(y[56]), .Z(n2392) );
  XNOR U5309 ( .A(x[634]), .B(y[634]), .Z(n2393) );
  XOR U5310 ( .A(n2392), .B(n2393), .Z(n2395) );
  XNOR U5311 ( .A(n2394), .B(n2395), .Z(n4814) );
  XNOR U5312 ( .A(n4815), .B(n4814), .Z(n2162) );
  XNOR U5313 ( .A(n2163), .B(n2162), .Z(n2164) );
  XNOR U5314 ( .A(n2165), .B(n2164), .Z(n2374) );
  XOR U5315 ( .A(x[38]), .B(y[38]), .Z(n2428) );
  XOR U5316 ( .A(x[32]), .B(y[32]), .Z(n2426) );
  XNOR U5317 ( .A(x[36]), .B(y[36]), .Z(n2427) );
  XOR U5318 ( .A(n2426), .B(n2427), .Z(n2429) );
  XNOR U5319 ( .A(n2428), .B(n2429), .Z(n5135) );
  XOR U5320 ( .A(x[923]), .B(y[923]), .Z(n1700) );
  XOR U5321 ( .A(x[426]), .B(y[426]), .Z(n1698) );
  XOR U5322 ( .A(x[925]), .B(y[925]), .Z(n1697) );
  XOR U5323 ( .A(n1698), .B(n1697), .Z(n1699) );
  XOR U5324 ( .A(n1700), .B(n1699), .Z(n5134) );
  XOR U5325 ( .A(n5135), .B(n5134), .Z(n5137) );
  XOR U5326 ( .A(x[16]), .B(y[16]), .Z(n4023) );
  XOR U5327 ( .A(x[12]), .B(y[12]), .Z(n4021) );
  XOR U5328 ( .A(x[612]), .B(y[612]), .Z(n4020) );
  XOR U5329 ( .A(n4021), .B(n4020), .Z(n4022) );
  XOR U5330 ( .A(n4023), .B(n4022), .Z(n5136) );
  XOR U5331 ( .A(n5137), .B(n5136), .Z(n1762) );
  XOR U5332 ( .A(x[10]), .B(y[10]), .Z(n4027) );
  XOR U5333 ( .A(x[6]), .B(y[6]), .Z(n4025) );
  XOR U5334 ( .A(x[608]), .B(y[608]), .Z(n4024) );
  XOR U5335 ( .A(n4025), .B(n4024), .Z(n4026) );
  XOR U5336 ( .A(n4027), .B(n4026), .Z(n4850) );
  XOR U5337 ( .A(x[1539]), .B(y[1539]), .Z(n4382) );
  XOR U5338 ( .A(x[40]), .B(y[40]), .Z(n4380) );
  XNOR U5339 ( .A(x[1541]), .B(y[1541]), .Z(n4381) );
  XOR U5340 ( .A(n4380), .B(n4381), .Z(n4383) );
  XOR U5341 ( .A(n4382), .B(n4383), .Z(n4851) );
  XNOR U5342 ( .A(n4850), .B(n4851), .Z(n4853) );
  XOR U5343 ( .A(x[4]), .B(y[4]), .Z(n4009) );
  XOR U5344 ( .A(x[0]), .B(y[0]), .Z(n4007) );
  XOR U5345 ( .A(x[1]), .B(y[1]), .Z(n4006) );
  XOR U5346 ( .A(n4007), .B(n4006), .Z(n4008) );
  XOR U5347 ( .A(n4009), .B(n4008), .Z(n4852) );
  XOR U5348 ( .A(n4853), .B(n4852), .Z(n1760) );
  XOR U5349 ( .A(x[5]), .B(y[5]), .Z(n4012) );
  XOR U5350 ( .A(x[9]), .B(y[9]), .Z(n4010) );
  XNOR U5351 ( .A(x[11]), .B(y[11]), .Z(n4011) );
  XOR U5352 ( .A(n4010), .B(n4011), .Z(n4013) );
  XNOR U5353 ( .A(n4012), .B(n4013), .Z(n5225) );
  XOR U5354 ( .A(x[931]), .B(y[931]), .Z(n1798) );
  XOR U5355 ( .A(x[420]), .B(y[420]), .Z(n1795) );
  XNOR U5356 ( .A(x[933]), .B(y[933]), .Z(n1796) );
  XNOR U5357 ( .A(n1795), .B(n1796), .Z(n1797) );
  XOR U5358 ( .A(n1798), .B(n1797), .Z(n5224) );
  XOR U5359 ( .A(n5225), .B(n5224), .Z(n5227) );
  XOR U5360 ( .A(x[15]), .B(y[15]), .Z(n2854) );
  XOR U5361 ( .A(x[17]), .B(y[17]), .Z(n2852) );
  XNOR U5362 ( .A(x[590]), .B(y[590]), .Z(n2853) );
  XOR U5363 ( .A(n2852), .B(n2853), .Z(n2855) );
  XNOR U5364 ( .A(n2854), .B(n2855), .Z(n5226) );
  XNOR U5365 ( .A(n5227), .B(n5226), .Z(n1759) );
  XNOR U5366 ( .A(n1760), .B(n1759), .Z(n1761) );
  XOR U5367 ( .A(n1762), .B(n1761), .Z(n2375) );
  XNOR U5368 ( .A(n2374), .B(n2375), .Z(n2377) );
  XOR U5369 ( .A(x[21]), .B(y[21]), .Z(n3378) );
  XOR U5370 ( .A(x[23]), .B(y[23]), .Z(n3376) );
  XNOR U5371 ( .A(x[584]), .B(y[584]), .Z(n3377) );
  XOR U5372 ( .A(n3376), .B(n3377), .Z(n3379) );
  XNOR U5373 ( .A(n3378), .B(n3379), .Z(n2066) );
  XOR U5374 ( .A(x[1535]), .B(y[1535]), .Z(n4388) );
  XOR U5375 ( .A(x[349]), .B(y[349]), .Z(n4386) );
  XNOR U5376 ( .A(x[1537]), .B(y[1537]), .Z(n4387) );
  XOR U5377 ( .A(n4386), .B(n4387), .Z(n4389) );
  XOR U5378 ( .A(n4388), .B(n4389), .Z(n2067) );
  XNOR U5379 ( .A(n2066), .B(n2067), .Z(n2069) );
  XOR U5380 ( .A(x[37]), .B(y[37]), .Z(n3342) );
  XOR U5381 ( .A(x[39]), .B(y[39]), .Z(n3340) );
  XNOR U5382 ( .A(x[43]), .B(y[43]), .Z(n3341) );
  XOR U5383 ( .A(n3340), .B(n3341), .Z(n3343) );
  XNOR U5384 ( .A(n3342), .B(n3343), .Z(n2068) );
  XOR U5385 ( .A(n2069), .B(n2068), .Z(n2325) );
  XOR U5386 ( .A(x[53]), .B(y[53]), .Z(n2832) );
  XOR U5387 ( .A(x[55]), .B(y[55]), .Z(n2830) );
  XNOR U5388 ( .A(x[562]), .B(y[562]), .Z(n2831) );
  XOR U5389 ( .A(n2830), .B(n2831), .Z(n2833) );
  XNOR U5390 ( .A(n2832), .B(n2833), .Z(n1966) );
  XOR U5391 ( .A(x[939]), .B(y[939]), .Z(n1803) );
  XOR U5392 ( .A(x[70]), .B(y[70]), .Z(n1801) );
  XNOR U5393 ( .A(x[941]), .B(y[941]), .Z(n1802) );
  XOR U5394 ( .A(n1801), .B(n1802), .Z(n1804) );
  XOR U5395 ( .A(n1803), .B(n1804), .Z(n1967) );
  XNOR U5396 ( .A(n1966), .B(n1967), .Z(n1969) );
  XOR U5397 ( .A(x[59]), .B(y[59]), .Z(n2772) );
  XOR U5398 ( .A(x[61]), .B(y[61]), .Z(n2770) );
  XNOR U5399 ( .A(x[65]), .B(y[65]), .Z(n2771) );
  XOR U5400 ( .A(n2770), .B(n2771), .Z(n2773) );
  XNOR U5401 ( .A(n2772), .B(n2773), .Z(n1968) );
  XOR U5402 ( .A(n1969), .B(n1968), .Z(n2323) );
  XOR U5403 ( .A(x[67]), .B(y[67]), .Z(n2778) );
  XOR U5404 ( .A(x[71]), .B(y[71]), .Z(n2776) );
  XNOR U5405 ( .A(x[75]), .B(y[75]), .Z(n2777) );
  XOR U5406 ( .A(n2776), .B(n2777), .Z(n2779) );
  XNOR U5407 ( .A(n2778), .B(n2779), .Z(n5076) );
  XOR U5408 ( .A(x[1531]), .B(y[1531]), .Z(n4720) );
  XOR U5409 ( .A(x[46]), .B(y[46]), .Z(n4718) );
  XNOR U5410 ( .A(x[1533]), .B(y[1533]), .Z(n4719) );
  XOR U5411 ( .A(n4718), .B(n4719), .Z(n4721) );
  XOR U5412 ( .A(n4720), .B(n4721), .Z(n5077) );
  XNOR U5413 ( .A(n5076), .B(n5077), .Z(n5079) );
  XOR U5414 ( .A(x[77]), .B(y[77]), .Z(n3915) );
  XOR U5415 ( .A(x[81]), .B(y[81]), .Z(n3913) );
  XOR U5416 ( .A(x[544]), .B(y[544]), .Z(n3912) );
  XOR U5417 ( .A(n3913), .B(n3912), .Z(n3914) );
  XOR U5418 ( .A(n3915), .B(n3914), .Z(n5078) );
  XNOR U5419 ( .A(n5079), .B(n5078), .Z(n2322) );
  XNOR U5420 ( .A(n2323), .B(n2322), .Z(n2324) );
  XNOR U5421 ( .A(n2325), .B(n2324), .Z(n2376) );
  XOR U5422 ( .A(n2377), .B(n2376), .Z(n2491) );
  XOR U5423 ( .A(x[209]), .B(y[209]), .Z(n2678) );
  XOR U5424 ( .A(x[213]), .B(y[213]), .Z(n2676) );
  XNOR U5425 ( .A(x[450]), .B(y[450]), .Z(n2677) );
  XOR U5426 ( .A(n2676), .B(n2677), .Z(n2679) );
  XNOR U5427 ( .A(n2678), .B(n2679), .Z(n3648) );
  XOR U5428 ( .A(x[971]), .B(y[971]), .Z(n2876) );
  XOR U5429 ( .A(x[42]), .B(y[42]), .Z(n2874) );
  XNOR U5430 ( .A(x[973]), .B(y[973]), .Z(n2875) );
  XOR U5431 ( .A(n2874), .B(n2875), .Z(n2877) );
  XOR U5432 ( .A(n2876), .B(n2877), .Z(n3649) );
  XNOR U5433 ( .A(n3648), .B(n3649), .Z(n3650) );
  XOR U5434 ( .A(x[215]), .B(y[215]), .Z(n2672) );
  XOR U5435 ( .A(x[219]), .B(y[219]), .Z(n2670) );
  XNOR U5436 ( .A(x[221]), .B(y[221]), .Z(n2671) );
  XOR U5437 ( .A(n2670), .B(n2671), .Z(n2673) );
  XOR U5438 ( .A(n2672), .B(n2673), .Z(n3651) );
  XNOR U5439 ( .A(n3650), .B(n3651), .Z(n4709) );
  XOR U5440 ( .A(x[225]), .B(y[225]), .Z(n2684) );
  XOR U5441 ( .A(x[229]), .B(y[229]), .Z(n2682) );
  XNOR U5442 ( .A(x[231]), .B(y[231]), .Z(n2683) );
  XOR U5443 ( .A(n2682), .B(n2683), .Z(n2685) );
  XNOR U5444 ( .A(n2684), .B(n2685), .Z(n3654) );
  XOR U5445 ( .A(x[1515]), .B(y[1515]), .Z(n2888) );
  XOR U5446 ( .A(x[337]), .B(y[337]), .Z(n2886) );
  XNOR U5447 ( .A(x[1517]), .B(y[1517]), .Z(n2887) );
  XOR U5448 ( .A(n2886), .B(n2887), .Z(n2889) );
  XOR U5449 ( .A(n2888), .B(n2889), .Z(n3655) );
  XNOR U5450 ( .A(n3654), .B(n3655), .Z(n3656) );
  XOR U5451 ( .A(x[235]), .B(y[235]), .Z(n994) );
  XOR U5452 ( .A(x[237]), .B(y[237]), .Z(n992) );
  XNOR U5453 ( .A(x[432]), .B(y[432]), .Z(n993) );
  XOR U5454 ( .A(n992), .B(n993), .Z(n995) );
  XOR U5455 ( .A(n994), .B(n995), .Z(n3657) );
  XNOR U5456 ( .A(n3656), .B(n3657), .Z(n4707) );
  XOR U5457 ( .A(x[247]), .B(y[247]), .Z(n3360) );
  XOR U5458 ( .A(x[251]), .B(y[251]), .Z(n3358) );
  XNOR U5459 ( .A(x[253]), .B(y[253]), .Z(n3359) );
  XOR U5460 ( .A(n3358), .B(n3359), .Z(n3361) );
  XNOR U5461 ( .A(n3360), .B(n3361), .Z(n3708) );
  XOR U5462 ( .A(x[979]), .B(y[979]), .Z(n1956) );
  XOR U5463 ( .A(x[34]), .B(y[34]), .Z(n1954) );
  XNOR U5464 ( .A(x[981]), .B(y[981]), .Z(n1955) );
  XOR U5465 ( .A(n1954), .B(n1955), .Z(n1957) );
  XOR U5466 ( .A(n1956), .B(n1957), .Z(n3709) );
  XNOR U5467 ( .A(n3708), .B(n3709), .Z(n3710) );
  XOR U5468 ( .A(x[265]), .B(y[265]), .Z(n3138) );
  XOR U5469 ( .A(x[269]), .B(y[269]), .Z(n3136) );
  XNOR U5470 ( .A(x[402]), .B(y[402]), .Z(n3137) );
  XOR U5471 ( .A(n3136), .B(n3137), .Z(n3139) );
  XOR U5472 ( .A(n3138), .B(n3139), .Z(n3711) );
  XNOR U5473 ( .A(n3710), .B(n3711), .Z(n4706) );
  XOR U5474 ( .A(n4707), .B(n4706), .Z(n4708) );
  XOR U5475 ( .A(n4709), .B(n4708), .Z(n5216) );
  XOR U5476 ( .A(x[147]), .B(y[147]), .Z(n2708) );
  XOR U5477 ( .A(x[149]), .B(y[149]), .Z(n2706) );
  XNOR U5478 ( .A(x[494]), .B(y[494]), .Z(n2707) );
  XOR U5479 ( .A(n2706), .B(n2707), .Z(n2709) );
  XNOR U5480 ( .A(n2708), .B(n2709), .Z(n4636) );
  XOR U5481 ( .A(x[1523]), .B(y[1523]), .Z(n4734) );
  XOR U5482 ( .A(x[343]), .B(y[343]), .Z(n4732) );
  XNOR U5483 ( .A(x[1525]), .B(y[1525]), .Z(n4733) );
  XOR U5484 ( .A(n4732), .B(n4733), .Z(n4735) );
  XOR U5485 ( .A(n4734), .B(n4735), .Z(n4637) );
  XNOR U5486 ( .A(n4636), .B(n4637), .Z(n4639) );
  XOR U5487 ( .A(x[153]), .B(y[153]), .Z(n2702) );
  XOR U5488 ( .A(x[155]), .B(y[155]), .Z(n2700) );
  XNOR U5489 ( .A(x[159]), .B(y[159]), .Z(n2701) );
  XOR U5490 ( .A(n2700), .B(n2701), .Z(n2703) );
  XNOR U5491 ( .A(n2702), .B(n2703), .Z(n4638) );
  XOR U5492 ( .A(n4639), .B(n4638), .Z(n1773) );
  XOR U5493 ( .A(x[163]), .B(y[163]), .Z(n980) );
  XOR U5494 ( .A(x[165]), .B(y[165]), .Z(n978) );
  XNOR U5495 ( .A(x[169]), .B(y[169]), .Z(n979) );
  XOR U5496 ( .A(n978), .B(n979), .Z(n981) );
  XNOR U5497 ( .A(n980), .B(n981), .Z(n4116) );
  XOR U5498 ( .A(x[963]), .B(y[963]), .Z(n1938) );
  XOR U5499 ( .A(x[400]), .B(y[400]), .Z(n1936) );
  XNOR U5500 ( .A(x[965]), .B(y[965]), .Z(n1937) );
  XOR U5501 ( .A(n1936), .B(n1937), .Z(n1939) );
  XOR U5502 ( .A(n1938), .B(n1939), .Z(n4117) );
  XNOR U5503 ( .A(n4116), .B(n4117), .Z(n4119) );
  XOR U5504 ( .A(x[177]), .B(y[177]), .Z(n3953) );
  XOR U5505 ( .A(x[181]), .B(y[181]), .Z(n3951) );
  XOR U5506 ( .A(x[472]), .B(y[472]), .Z(n3950) );
  XOR U5507 ( .A(n3951), .B(n3950), .Z(n3952) );
  XOR U5508 ( .A(n3953), .B(n3952), .Z(n4118) );
  XOR U5509 ( .A(n4119), .B(n4118), .Z(n1772) );
  XOR U5510 ( .A(x[193]), .B(y[193]), .Z(n3102) );
  XOR U5511 ( .A(x[197]), .B(y[197]), .Z(n3100) );
  XNOR U5512 ( .A(x[199]), .B(y[199]), .Z(n3101) );
  XOR U5513 ( .A(n3100), .B(n3101), .Z(n3103) );
  XNOR U5514 ( .A(n3102), .B(n3103), .Z(n3624) );
  XOR U5515 ( .A(x[1519]), .B(y[1519]), .Z(n4740) );
  XOR U5516 ( .A(x[1521]), .B(y[1521]), .Z(n4738) );
  XNOR U5517 ( .A(x[1592]), .B(y[1592]), .Z(n4739) );
  XOR U5518 ( .A(n4738), .B(n4739), .Z(n4741) );
  XOR U5519 ( .A(n4740), .B(n4741), .Z(n3625) );
  XNOR U5520 ( .A(n3624), .B(n3625), .Z(n3627) );
  XOR U5521 ( .A(x[203]), .B(y[203]), .Z(n3114) );
  XOR U5522 ( .A(x[207]), .B(y[207]), .Z(n3112) );
  XNOR U5523 ( .A(x[454]), .B(y[454]), .Z(n3113) );
  XOR U5524 ( .A(n3112), .B(n3113), .Z(n3115) );
  XNOR U5525 ( .A(n3114), .B(n3115), .Z(n3626) );
  XNOR U5526 ( .A(n3627), .B(n3626), .Z(n1771) );
  XOR U5527 ( .A(n1772), .B(n1771), .Z(n1774) );
  XOR U5528 ( .A(n1773), .B(n1774), .Z(n5215) );
  XOR U5529 ( .A(x[83]), .B(y[83]), .Z(n3919) );
  XOR U5530 ( .A(x[87]), .B(y[87]), .Z(n3917) );
  XOR U5531 ( .A(x[538]), .B(y[538]), .Z(n3916) );
  XOR U5532 ( .A(n3917), .B(n3916), .Z(n3918) );
  XOR U5533 ( .A(n3919), .B(n3918), .Z(n4956) );
  XOR U5534 ( .A(x[947]), .B(y[947]), .Z(n4882) );
  XOR U5535 ( .A(x[62]), .B(y[62]), .Z(n4880) );
  XNOR U5536 ( .A(x[949]), .B(y[949]), .Z(n4881) );
  XOR U5537 ( .A(n4880), .B(n4881), .Z(n4883) );
  XOR U5538 ( .A(n4882), .B(n4883), .Z(n4957) );
  XNOR U5539 ( .A(n4956), .B(n4957), .Z(n4959) );
  XOR U5540 ( .A(x[89]), .B(y[89]), .Z(n962) );
  XOR U5541 ( .A(x[93]), .B(y[93]), .Z(n960) );
  XNOR U5542 ( .A(x[97]), .B(y[97]), .Z(n961) );
  XOR U5543 ( .A(n960), .B(n961), .Z(n963) );
  XNOR U5544 ( .A(n962), .B(n963), .Z(n4958) );
  XOR U5545 ( .A(n4959), .B(n4958), .Z(n1767) );
  XOR U5546 ( .A(x[131]), .B(y[131]), .Z(n2728) );
  XOR U5547 ( .A(x[133]), .B(y[133]), .Z(n2726) );
  XNOR U5548 ( .A(x[137]), .B(y[137]), .Z(n2727) );
  XOR U5549 ( .A(n2726), .B(n2727), .Z(n2729) );
  XNOR U5550 ( .A(n2728), .B(n2729), .Z(n4677) );
  XOR U5551 ( .A(x[955]), .B(y[955]), .Z(n1933) );
  XOR U5552 ( .A(x[406]), .B(y[406]), .Z(n1930) );
  XNOR U5553 ( .A(x[957]), .B(y[957]), .Z(n1931) );
  XNOR U5554 ( .A(n1930), .B(n1931), .Z(n1932) );
  XOR U5555 ( .A(n1933), .B(n1932), .Z(n4676) );
  XOR U5556 ( .A(n4677), .B(n4676), .Z(n4679) );
  XOR U5557 ( .A(x[141]), .B(y[141]), .Z(n2740) );
  XOR U5558 ( .A(x[143]), .B(y[143]), .Z(n2738) );
  XNOR U5559 ( .A(x[498]), .B(y[498]), .Z(n2739) );
  XOR U5560 ( .A(n2738), .B(n2739), .Z(n2741) );
  XNOR U5561 ( .A(n2740), .B(n2741), .Z(n4678) );
  XOR U5562 ( .A(n4679), .B(n4678), .Z(n1766) );
  XOR U5563 ( .A(x[109]), .B(y[109]), .Z(n1012) );
  XOR U5564 ( .A(x[111]), .B(y[111]), .Z(n1010) );
  XNOR U5565 ( .A(x[522]), .B(y[522]), .Z(n1011) );
  XOR U5566 ( .A(n1010), .B(n1011), .Z(n1013) );
  XNOR U5567 ( .A(n1012), .B(n1013), .Z(n4825) );
  XOR U5568 ( .A(x[1527]), .B(y[1527]), .Z(n4727) );
  XOR U5569 ( .A(x[1529]), .B(y[1529]), .Z(n4725) );
  XOR U5570 ( .A(x[1594]), .B(y[1594]), .Z(n4724) );
  XOR U5571 ( .A(n4725), .B(n4724), .Z(n4726) );
  XOR U5572 ( .A(n4727), .B(n4726), .Z(n4824) );
  XOR U5573 ( .A(n4825), .B(n4824), .Z(n4827) );
  XOR U5574 ( .A(x[121]), .B(y[121]), .Z(n2734) );
  XOR U5575 ( .A(x[125]), .B(y[125]), .Z(n2732) );
  XNOR U5576 ( .A(x[127]), .B(y[127]), .Z(n2733) );
  XOR U5577 ( .A(n2732), .B(n2733), .Z(n2735) );
  XNOR U5578 ( .A(n2734), .B(n2735), .Z(n4826) );
  XNOR U5579 ( .A(n4827), .B(n4826), .Z(n1765) );
  XOR U5580 ( .A(n1766), .B(n1765), .Z(n1768) );
  XNOR U5581 ( .A(n1767), .B(n1768), .Z(n5214) );
  XNOR U5582 ( .A(n5215), .B(n5214), .Z(n5217) );
  XOR U5583 ( .A(n5216), .B(n5217), .Z(n2490) );
  XNOR U5584 ( .A(n2491), .B(n2490), .Z(n2492) );
  XOR U5585 ( .A(n2493), .B(n2492), .Z(n1344) );
  XOR U5586 ( .A(x[616]), .B(y[616]), .Z(n1583) );
  XOR U5587 ( .A(x[614]), .B(y[614]), .Z(n1581) );
  XNOR U5588 ( .A(x[1466]), .B(y[1466]), .Z(n1582) );
  XOR U5589 ( .A(n1581), .B(n1582), .Z(n1584) );
  XNOR U5590 ( .A(n1583), .B(n1584), .Z(n4551) );
  XOR U5591 ( .A(x[1583]), .B(y[1583]), .Z(n3753) );
  XOR U5592 ( .A(x[789]), .B(y[789]), .Z(n3750) );
  XNOR U5593 ( .A(x[1585]), .B(y[1585]), .Z(n3751) );
  XNOR U5594 ( .A(n3750), .B(n3751), .Z(n3752) );
  XOR U5595 ( .A(n3753), .B(n3752), .Z(n4550) );
  XOR U5596 ( .A(n4551), .B(n4550), .Z(n4553) );
  XOR U5597 ( .A(x[610]), .B(y[610]), .Z(n1589) );
  XOR U5598 ( .A(x[604]), .B(y[604]), .Z(n1587) );
  XNOR U5599 ( .A(x[1070]), .B(y[1070]), .Z(n1588) );
  XOR U5600 ( .A(n1587), .B(n1588), .Z(n1590) );
  XNOR U5601 ( .A(n1589), .B(n1590), .Z(n4552) );
  XOR U5602 ( .A(n4553), .B(n4552), .Z(n1362) );
  XOR U5603 ( .A(x[602]), .B(y[602]), .Z(n1601) );
  XOR U5604 ( .A(x[598]), .B(y[598]), .Z(n1599) );
  XNOR U5605 ( .A(x[872]), .B(y[872]), .Z(n1600) );
  XOR U5606 ( .A(n1599), .B(n1600), .Z(n1602) );
  XNOR U5607 ( .A(n1601), .B(n1602), .Z(n4532) );
  XOR U5608 ( .A(x[843]), .B(y[843]), .Z(n2022) );
  XOR U5609 ( .A(x[152]), .B(y[152]), .Z(n2020) );
  XNOR U5610 ( .A(x[845]), .B(y[845]), .Z(n2021) );
  XOR U5611 ( .A(n2020), .B(n2021), .Z(n2023) );
  XOR U5612 ( .A(n2022), .B(n2023), .Z(n4533) );
  XNOR U5613 ( .A(n4532), .B(n4533), .Z(n4535) );
  XOR U5614 ( .A(x[596]), .B(y[596]), .Z(n1607) );
  XOR U5615 ( .A(x[592]), .B(y[592]), .Z(n1605) );
  XNOR U5616 ( .A(x[594]), .B(y[594]), .Z(n1606) );
  XOR U5617 ( .A(n1605), .B(n1606), .Z(n1608) );
  XNOR U5618 ( .A(n1607), .B(n1608), .Z(n4534) );
  XOR U5619 ( .A(n4535), .B(n4534), .Z(n1360) );
  XOR U5620 ( .A(x[588]), .B(y[588]), .Z(n4438) );
  XOR U5621 ( .A(x[578]), .B(y[578]), .Z(n4436) );
  XNOR U5622 ( .A(x[582]), .B(y[582]), .Z(n4437) );
  XOR U5623 ( .A(n4436), .B(n4437), .Z(n4439) );
  XNOR U5624 ( .A(n4438), .B(n4439), .Z(n4555) );
  XOR U5625 ( .A(x[1579]), .B(y[1579]), .Z(n3809) );
  XOR U5626 ( .A(x[381]), .B(y[381]), .Z(n3806) );
  XNOR U5627 ( .A(x[1581]), .B(y[1581]), .Z(n3807) );
  XNOR U5628 ( .A(n3806), .B(n3807), .Z(n3808) );
  XOR U5629 ( .A(n3809), .B(n3808), .Z(n4554) );
  XOR U5630 ( .A(n4555), .B(n4554), .Z(n4557) );
  XOR U5631 ( .A(x[564]), .B(y[564]), .Z(n1480) );
  XOR U5632 ( .A(x[556]), .B(y[556]), .Z(n1477) );
  XNOR U5633 ( .A(x[558]), .B(y[558]), .Z(n1478) );
  XOR U5634 ( .A(n1480), .B(n1479), .Z(n4556) );
  XNOR U5635 ( .A(n4557), .B(n4556), .Z(n1359) );
  XNOR U5636 ( .A(n1360), .B(n1359), .Z(n1361) );
  XNOR U5637 ( .A(n1362), .B(n1361), .Z(n5116) );
  XOR U5638 ( .A(x[554]), .B(y[554]), .Z(n5143) );
  XOR U5639 ( .A(x[550]), .B(y[550]), .Z(n5140) );
  XNOR U5640 ( .A(x[552]), .B(y[552]), .Z(n5141) );
  XOR U5641 ( .A(n5143), .B(n5142), .Z(n4567) );
  XOR U5642 ( .A(x[851]), .B(y[851]), .Z(n2017) );
  XOR U5643 ( .A(x[144]), .B(y[144]), .Z(n2014) );
  XNOR U5644 ( .A(x[853]), .B(y[853]), .Z(n2015) );
  XNOR U5645 ( .A(n2014), .B(n2015), .Z(n2016) );
  XOR U5646 ( .A(n2017), .B(n2016), .Z(n4566) );
  XOR U5647 ( .A(n4567), .B(n4566), .Z(n4569) );
  XOR U5648 ( .A(x[536]), .B(y[536]), .Z(n1820) );
  XOR U5649 ( .A(x[534]), .B(y[534]), .Z(n1817) );
  XNOR U5650 ( .A(x[836]), .B(y[836]), .Z(n1818) );
  XOR U5651 ( .A(n1820), .B(n1819), .Z(n4568) );
  XOR U5652 ( .A(n4569), .B(n4568), .Z(n1446) );
  XOR U5653 ( .A(x[524]), .B(y[524]), .Z(n1508) );
  XOR U5654 ( .A(x[514]), .B(y[514]), .Z(n1505) );
  XNOR U5655 ( .A(x[518]), .B(y[518]), .Z(n1506) );
  XOR U5656 ( .A(n1508), .B(n1507), .Z(n4559) );
  XOR U5657 ( .A(x[1575]), .B(y[1575]), .Z(n3889) );
  XOR U5658 ( .A(x[377]), .B(y[377]), .Z(n3886) );
  XNOR U5659 ( .A(x[1577]), .B(y[1577]), .Z(n3887) );
  XNOR U5660 ( .A(n3886), .B(n3887), .Z(n3888) );
  XOR U5661 ( .A(n3889), .B(n3888), .Z(n4558) );
  XOR U5662 ( .A(n4559), .B(n4558), .Z(n4561) );
  XOR U5663 ( .A(x[512]), .B(y[512]), .Z(n4490) );
  XOR U5664 ( .A(x[510]), .B(y[510]), .Z(n4488) );
  XNOR U5665 ( .A(x[822]), .B(y[822]), .Z(n4489) );
  XOR U5666 ( .A(n4488), .B(n4489), .Z(n4491) );
  XNOR U5667 ( .A(n4490), .B(n4491), .Z(n4560) );
  XOR U5668 ( .A(n4561), .B(n4560), .Z(n1444) );
  XOR U5669 ( .A(x[508]), .B(y[508]), .Z(n4496) );
  XOR U5670 ( .A(x[504]), .B(y[504]), .Z(n4494) );
  XNOR U5671 ( .A(x[818]), .B(y[818]), .Z(n4495) );
  XOR U5672 ( .A(n4494), .B(n4495), .Z(n4497) );
  XNOR U5673 ( .A(n4496), .B(n4497), .Z(n3618) );
  XOR U5674 ( .A(x[859]), .B(y[859]), .Z(n2028) );
  XOR U5675 ( .A(x[466]), .B(y[466]), .Z(n2026) );
  XNOR U5676 ( .A(x[861]), .B(y[861]), .Z(n2027) );
  XOR U5677 ( .A(n2026), .B(n2027), .Z(n2029) );
  XOR U5678 ( .A(n2028), .B(n2029), .Z(n3619) );
  XNOR U5679 ( .A(n3618), .B(n3619), .Z(n3621) );
  XOR U5680 ( .A(x[502]), .B(y[502]), .Z(n1373) );
  XOR U5681 ( .A(x[492]), .B(y[492]), .Z(n1371) );
  XNOR U5682 ( .A(x[496]), .B(y[496]), .Z(n1372) );
  XOR U5683 ( .A(n1371), .B(n1372), .Z(n1374) );
  XNOR U5684 ( .A(n1373), .B(n1374), .Z(n3620) );
  XNOR U5685 ( .A(n3621), .B(n3620), .Z(n1443) );
  XNOR U5686 ( .A(n1444), .B(n1443), .Z(n1445) );
  XOR U5687 ( .A(n1446), .B(n1445), .Z(n5117) );
  XNOR U5688 ( .A(n5116), .B(n5117), .Z(n5119) );
  XOR U5689 ( .A(x[490]), .B(y[490]), .Z(n1379) );
  XOR U5690 ( .A(x[484]), .B(y[484]), .Z(n1377) );
  XNOR U5691 ( .A(x[488]), .B(y[488]), .Z(n1378) );
  XOR U5692 ( .A(n1377), .B(n1378), .Z(n1380) );
  XNOR U5693 ( .A(n1379), .B(n1380), .Z(n4563) );
  XOR U5694 ( .A(x[1571]), .B(y[1571]), .Z(n3923) );
  XOR U5695 ( .A(x[20]), .B(y[20]), .Z(n3920) );
  XNOR U5696 ( .A(x[1573]), .B(y[1573]), .Z(n3921) );
  XNOR U5697 ( .A(n3920), .B(n3921), .Z(n3922) );
  XOR U5698 ( .A(n3923), .B(n3922), .Z(n4562) );
  XOR U5699 ( .A(n4563), .B(n4562), .Z(n4565) );
  XOR U5700 ( .A(x[482]), .B(y[482]), .Z(n2128) );
  XOR U5701 ( .A(x[478]), .B(y[478]), .Z(n2126) );
  XNOR U5702 ( .A(x[804]), .B(y[804]), .Z(n2127) );
  XOR U5703 ( .A(n2126), .B(n2127), .Z(n2129) );
  XNOR U5704 ( .A(n2128), .B(n2129), .Z(n4564) );
  XOR U5705 ( .A(n4565), .B(n4564), .Z(n1440) );
  XOR U5706 ( .A(x[468]), .B(y[468]), .Z(n1974) );
  XOR U5707 ( .A(x[462]), .B(y[462]), .Z(n1972) );
  XNOR U5708 ( .A(x[464]), .B(y[464]), .Z(n1973) );
  XOR U5709 ( .A(n1972), .B(n1973), .Z(n1975) );
  XNOR U5710 ( .A(n1974), .B(n1975), .Z(n4526) );
  XOR U5711 ( .A(x[867]), .B(y[867]), .Z(n2040) );
  XOR U5712 ( .A(x[460]), .B(y[460]), .Z(n2038) );
  XNOR U5713 ( .A(x[869]), .B(y[869]), .Z(n2039) );
  XOR U5714 ( .A(n2038), .B(n2039), .Z(n2041) );
  XOR U5715 ( .A(n2040), .B(n2041), .Z(n4527) );
  XNOR U5716 ( .A(n4526), .B(n4527), .Z(n4529) );
  XOR U5717 ( .A(x[448]), .B(y[448]), .Z(n4509) );
  XOR U5718 ( .A(x[444]), .B(y[444]), .Z(n4507) );
  XOR U5719 ( .A(x[786]), .B(y[786]), .Z(n4506) );
  XOR U5720 ( .A(n4507), .B(n4506), .Z(n4508) );
  XOR U5721 ( .A(n4509), .B(n4508), .Z(n4528) );
  XOR U5722 ( .A(n4529), .B(n4528), .Z(n1438) );
  XOR U5723 ( .A(x[442]), .B(y[442]), .Z(n4513) );
  XOR U5724 ( .A(x[438]), .B(y[438]), .Z(n4511) );
  XOR U5725 ( .A(x[782]), .B(y[782]), .Z(n4510) );
  XOR U5726 ( .A(n4511), .B(n4510), .Z(n4512) );
  XOR U5727 ( .A(n4513), .B(n4512), .Z(n4660) );
  XOR U5728 ( .A(x[1567]), .B(y[1567]), .Z(n3014) );
  XOR U5729 ( .A(x[371]), .B(y[371]), .Z(n3012) );
  XNOR U5730 ( .A(x[1569]), .B(y[1569]), .Z(n3013) );
  XOR U5731 ( .A(n3012), .B(n3013), .Z(n3015) );
  XOR U5732 ( .A(n3014), .B(n3015), .Z(n4661) );
  XNOR U5733 ( .A(n4660), .B(n4661), .Z(n4663) );
  XOR U5734 ( .A(x[436]), .B(y[436]), .Z(n4460) );
  XOR U5735 ( .A(x[430]), .B(y[430]), .Z(n4458) );
  XNOR U5736 ( .A(x[434]), .B(y[434]), .Z(n4459) );
  XOR U5737 ( .A(n4458), .B(n4459), .Z(n4461) );
  XNOR U5738 ( .A(n4460), .B(n4461), .Z(n4662) );
  XNOR U5739 ( .A(n4663), .B(n4662), .Z(n1437) );
  XNOR U5740 ( .A(n1438), .B(n1437), .Z(n1439) );
  XNOR U5741 ( .A(n1440), .B(n1439), .Z(n5118) );
  XOR U5742 ( .A(n5119), .B(n5118), .Z(n5105) );
  XOR U5743 ( .A(x[654]), .B(y[654]), .Z(n2938) );
  XOR U5744 ( .A(x[650]), .B(y[650]), .Z(n2936) );
  XNOR U5745 ( .A(x[1460]), .B(y[1460]), .Z(n2937) );
  XOR U5746 ( .A(n2936), .B(n2937), .Z(n2939) );
  XNOR U5747 ( .A(n2938), .B(n2939), .Z(n3984) );
  XOR U5748 ( .A(x[827]), .B(y[827]), .Z(n2276) );
  XOR U5749 ( .A(x[486]), .B(y[486]), .Z(n2274) );
  XNOR U5750 ( .A(x[829]), .B(y[829]), .Z(n2275) );
  XOR U5751 ( .A(n2274), .B(n2275), .Z(n2277) );
  XOR U5752 ( .A(n2276), .B(n2277), .Z(n3985) );
  XNOR U5753 ( .A(n3984), .B(n3985), .Z(n3987) );
  XOR U5754 ( .A(x[648]), .B(y[648]), .Z(n2944) );
  XOR U5755 ( .A(x[644]), .B(y[644]), .Z(n2942) );
  XNOR U5756 ( .A(x[1082]), .B(y[1082]), .Z(n2943) );
  XOR U5757 ( .A(n2942), .B(n2943), .Z(n2945) );
  XNOR U5758 ( .A(n2944), .B(n2945), .Z(n3986) );
  XOR U5759 ( .A(n3987), .B(n3986), .Z(n4432) );
  XOR U5760 ( .A(x[642]), .B(y[642]), .Z(n4590) );
  XOR U5761 ( .A(x[638]), .B(y[638]), .Z(n4588) );
  XNOR U5762 ( .A(x[1462]), .B(y[1462]), .Z(n4589) );
  XOR U5763 ( .A(n4588), .B(n4589), .Z(n4591) );
  XNOR U5764 ( .A(n4590), .B(n4591), .Z(n4129) );
  XOR U5765 ( .A(x[1587]), .B(y[1587]), .Z(n3699) );
  XOR U5766 ( .A(x[1589]), .B(y[1589]), .Z(n3697) );
  XOR U5767 ( .A(x[1591]), .B(y[1591]), .Z(n3696) );
  XOR U5768 ( .A(n3697), .B(n3696), .Z(n3698) );
  XOR U5769 ( .A(n3699), .B(n3698), .Z(n4128) );
  XOR U5770 ( .A(n4129), .B(n4128), .Z(n4131) );
  XOR U5771 ( .A(x[636]), .B(y[636]), .Z(n4596) );
  XOR U5772 ( .A(x[632]), .B(y[632]), .Z(n4594) );
  XNOR U5773 ( .A(x[1078]), .B(y[1078]), .Z(n4595) );
  XOR U5774 ( .A(n4594), .B(n4595), .Z(n4597) );
  XNOR U5775 ( .A(n4596), .B(n4597), .Z(n4130) );
  XOR U5776 ( .A(n4131), .B(n4130), .Z(n4431) );
  XOR U5777 ( .A(x[628]), .B(y[628]), .Z(n4608) );
  XOR U5778 ( .A(x[624]), .B(y[624]), .Z(n4606) );
  XNOR U5779 ( .A(x[1464]), .B(y[1464]), .Z(n4607) );
  XOR U5780 ( .A(n4606), .B(n4607), .Z(n4609) );
  XNOR U5781 ( .A(n4608), .B(n4609), .Z(n1223) );
  XOR U5782 ( .A(x[835]), .B(y[835]), .Z(n2288) );
  XOR U5783 ( .A(x[480]), .B(y[480]), .Z(n2286) );
  XNOR U5784 ( .A(x[837]), .B(y[837]), .Z(n2287) );
  XOR U5785 ( .A(n2286), .B(n2287), .Z(n2289) );
  XOR U5786 ( .A(n2288), .B(n2289), .Z(n1224) );
  XNOR U5787 ( .A(n1223), .B(n1224), .Z(n1226) );
  XOR U5788 ( .A(x[622]), .B(y[622]), .Z(n4614) );
  XOR U5789 ( .A(x[618]), .B(y[618]), .Z(n4612) );
  XNOR U5790 ( .A(x[1074]), .B(y[1074]), .Z(n4613) );
  XOR U5791 ( .A(n4612), .B(n4613), .Z(n4615) );
  XNOR U5792 ( .A(n4614), .B(n4615), .Z(n1225) );
  XNOR U5793 ( .A(n1226), .B(n1225), .Z(n4430) );
  XOR U5794 ( .A(n4431), .B(n4430), .Z(n4433) );
  XOR U5795 ( .A(n4432), .B(n4433), .Z(n5183) );
  XOR U5796 ( .A(x[684]), .B(y[684]), .Z(n4311) );
  XOR U5797 ( .A(x[682]), .B(y[682]), .Z(n4309) );
  XOR U5798 ( .A(x[1094]), .B(y[1094]), .Z(n4308) );
  XOR U5799 ( .A(n4309), .B(n4308), .Z(n4310) );
  XOR U5800 ( .A(n4311), .B(n4310), .Z(n2637) );
  XOR U5801 ( .A(x[595]), .B(y[595]), .Z(n1882) );
  XOR U5802 ( .A(x[597]), .B(y[597]), .Z(n1881) );
  XOR U5803 ( .A(n1882), .B(n1881), .Z(n945) );
  XOR U5804 ( .A(x[589]), .B(y[589]), .Z(n942) );
  XNOR U5805 ( .A(x[1597]), .B(y[1597]), .Z(n943) );
  XNOR U5806 ( .A(n942), .B(n943), .Z(n944) );
  XOR U5807 ( .A(n945), .B(n944), .Z(n2635) );
  XOR U5808 ( .A(x[688]), .B(y[688]), .Z(n4307) );
  XOR U5809 ( .A(x[686]), .B(y[686]), .Z(n4305) );
  XOR U5810 ( .A(x[1454]), .B(y[1454]), .Z(n4304) );
  XOR U5811 ( .A(n4305), .B(n4304), .Z(n4306) );
  XNOR U5812 ( .A(n4307), .B(n4306), .Z(n2634) );
  XNOR U5813 ( .A(n2635), .B(n2634), .Z(n2636) );
  XNOR U5814 ( .A(n2637), .B(n2636), .Z(n2927) );
  XOR U5815 ( .A(x[680]), .B(y[680]), .Z(n4339) );
  XOR U5816 ( .A(x[676]), .B(y[676]), .Z(n4337) );
  XOR U5817 ( .A(x[1456]), .B(y[1456]), .Z(n4336) );
  XOR U5818 ( .A(n4337), .B(n4336), .Z(n4338) );
  XOR U5819 ( .A(n4339), .B(n4338), .Z(n2598) );
  XOR U5820 ( .A(x[819]), .B(y[819]), .Z(n2282) );
  XOR U5821 ( .A(x[172]), .B(y[172]), .Z(n2280) );
  XNOR U5822 ( .A(x[821]), .B(y[821]), .Z(n2281) );
  XOR U5823 ( .A(n2280), .B(n2281), .Z(n2283) );
  XOR U5824 ( .A(n2282), .B(n2283), .Z(n2599) );
  XNOR U5825 ( .A(n2598), .B(n2599), .Z(n2601) );
  XOR U5826 ( .A(x[672]), .B(y[672]), .Z(n4343) );
  XOR U5827 ( .A(x[670]), .B(y[670]), .Z(n4341) );
  XOR U5828 ( .A(x[1090]), .B(y[1090]), .Z(n4340) );
  XOR U5829 ( .A(n4341), .B(n4340), .Z(n4342) );
  XOR U5830 ( .A(n4343), .B(n4342), .Z(n2600) );
  XOR U5831 ( .A(n2601), .B(n2600), .Z(n2925) );
  XOR U5832 ( .A(x[668]), .B(y[668]), .Z(n4353) );
  XOR U5833 ( .A(x[664]), .B(y[664]), .Z(n4351) );
  XOR U5834 ( .A(x[1458]), .B(y[1458]), .Z(n4350) );
  XOR U5835 ( .A(n4351), .B(n4350), .Z(n4352) );
  XOR U5836 ( .A(n4353), .B(n4352), .Z(n2610) );
  XOR U5837 ( .A(x[1593]), .B(y[1593]), .Z(n3632) );
  XOR U5838 ( .A(x[587]), .B(y[587]), .Z(n3630) );
  XNOR U5839 ( .A(x[1595]), .B(y[1595]), .Z(n3631) );
  XOR U5840 ( .A(n3630), .B(n3631), .Z(n3633) );
  XOR U5841 ( .A(n3632), .B(n3633), .Z(n2611) );
  XNOR U5842 ( .A(n2610), .B(n2611), .Z(n2613) );
  XOR U5843 ( .A(x[662]), .B(y[662]), .Z(n4357) );
  XOR U5844 ( .A(x[658]), .B(y[658]), .Z(n4355) );
  XOR U5845 ( .A(x[1086]), .B(y[1086]), .Z(n4354) );
  XOR U5846 ( .A(n4355), .B(n4354), .Z(n4356) );
  XOR U5847 ( .A(n4357), .B(n4356), .Z(n2612) );
  XNOR U5848 ( .A(n2613), .B(n2612), .Z(n2924) );
  XNOR U5849 ( .A(n2925), .B(n2924), .Z(n2926) );
  XOR U5850 ( .A(n2927), .B(n2926), .Z(n5181) );
  XOR U5851 ( .A(x[724]), .B(y[724]), .Z(n4228) );
  XOR U5852 ( .A(x[722]), .B(y[722]), .Z(n4226) );
  XNOR U5853 ( .A(x[1110]), .B(y[1110]), .Z(n4227) );
  XOR U5854 ( .A(n4226), .B(n4227), .Z(n4229) );
  XNOR U5855 ( .A(n4228), .B(n4229), .Z(n2617) );
  XOR U5856 ( .A(x[720]), .B(y[720]), .Z(n4245) );
  XOR U5857 ( .A(x[718]), .B(y[718]), .Z(n4242) );
  XNOR U5858 ( .A(x[1448]), .B(y[1448]), .Z(n4243) );
  XNOR U5859 ( .A(n4242), .B(n4243), .Z(n4244) );
  XOR U5860 ( .A(n4245), .B(n4244), .Z(n2616) );
  XOR U5861 ( .A(n2617), .B(n2616), .Z(n2619) );
  XOR U5862 ( .A(x[716]), .B(y[716]), .Z(n4251) );
  XOR U5863 ( .A(x[712]), .B(y[712]), .Z(n4248) );
  XNOR U5864 ( .A(x[1106]), .B(y[1106]), .Z(n4249) );
  XNOR U5865 ( .A(n4248), .B(n4249), .Z(n4250) );
  XOR U5866 ( .A(n4251), .B(n4250), .Z(n2618) );
  XOR U5867 ( .A(n2619), .B(n2618), .Z(n2871) );
  XOR U5868 ( .A(x[708]), .B(y[708]), .Z(n4263) );
  XOR U5869 ( .A(x[706]), .B(y[706]), .Z(n4261) );
  XOR U5870 ( .A(x[1450]), .B(y[1450]), .Z(n4260) );
  XOR U5871 ( .A(n4261), .B(n4260), .Z(n4262) );
  XOR U5872 ( .A(n4263), .B(n4262), .Z(n2605) );
  XOR U5873 ( .A(x[591]), .B(y[591]), .Z(n1037) );
  XOR U5874 ( .A(x[599]), .B(y[599]), .Z(n1035) );
  XOR U5875 ( .A(x[1599]), .B(y[1599]), .Z(n1034) );
  XOR U5876 ( .A(n1035), .B(n1034), .Z(n1036) );
  XOR U5877 ( .A(n1037), .B(n1036), .Z(n2604) );
  XOR U5878 ( .A(n2605), .B(n2604), .Z(n2607) );
  XOR U5879 ( .A(x[704]), .B(y[704]), .Z(n4267) );
  XOR U5880 ( .A(x[702]), .B(y[702]), .Z(n4265) );
  XOR U5881 ( .A(x[1102]), .B(y[1102]), .Z(n4264) );
  XOR U5882 ( .A(n4265), .B(n4264), .Z(n4266) );
  XOR U5883 ( .A(n4267), .B(n4266), .Z(n2606) );
  XOR U5884 ( .A(n2607), .B(n2606), .Z(n2869) );
  XOR U5885 ( .A(x[700]), .B(y[700]), .Z(n4295) );
  XOR U5886 ( .A(x[698]), .B(y[698]), .Z(n4293) );
  XOR U5887 ( .A(x[1452]), .B(y[1452]), .Z(n4292) );
  XOR U5888 ( .A(n4293), .B(n4292), .Z(n4294) );
  XOR U5889 ( .A(n4295), .B(n4294), .Z(n2647) );
  XOR U5890 ( .A(x[811]), .B(y[811]), .Z(n4445) );
  XOR U5891 ( .A(x[178]), .B(y[178]), .Z(n4443) );
  XOR U5892 ( .A(x[813]), .B(y[813]), .Z(n4442) );
  XOR U5893 ( .A(n4443), .B(n4442), .Z(n4444) );
  XOR U5894 ( .A(n4445), .B(n4444), .Z(n2646) );
  XOR U5895 ( .A(n2647), .B(n2646), .Z(n2649) );
  XOR U5896 ( .A(x[694]), .B(y[694]), .Z(n4299) );
  XOR U5897 ( .A(x[690]), .B(y[690]), .Z(n4297) );
  XOR U5898 ( .A(x[1098]), .B(y[1098]), .Z(n4296) );
  XOR U5899 ( .A(n4297), .B(n4296), .Z(n4298) );
  XOR U5900 ( .A(n4299), .B(n4298), .Z(n2648) );
  XOR U5901 ( .A(n2649), .B(n2648), .Z(n2868) );
  XOR U5902 ( .A(n2869), .B(n2868), .Z(n2870) );
  XOR U5903 ( .A(n2871), .B(n2870), .Z(n5180) );
  XNOR U5904 ( .A(n5181), .B(n5180), .Z(n5182) );
  XNOR U5905 ( .A(n5183), .B(n5182), .Z(n5104) );
  XNOR U5906 ( .A(n5105), .B(n5104), .Z(n5107) );
  XOR U5907 ( .A(x[760]), .B(y[760]), .Z(n3042) );
  XOR U5908 ( .A(x[758]), .B(y[758]), .Z(n3040) );
  XNOR U5909 ( .A(x[1440]), .B(y[1440]), .Z(n3041) );
  XOR U5910 ( .A(n3040), .B(n3041), .Z(n3043) );
  XNOR U5911 ( .A(n3042), .B(n3043), .Z(n2629) );
  XOR U5912 ( .A(x[309]), .B(y[309]), .Z(n3169) );
  XOR U5913 ( .A(x[313]), .B(y[313]), .Z(n3166) );
  XNOR U5914 ( .A(x[317]), .B(y[317]), .Z(n3167) );
  XNOR U5915 ( .A(n3166), .B(n3167), .Z(n3168) );
  XOR U5916 ( .A(n3169), .B(n3168), .Z(n2628) );
  XOR U5917 ( .A(n2629), .B(n2628), .Z(n2631) );
  XOR U5918 ( .A(x[756]), .B(y[756]), .Z(n3048) );
  XOR U5919 ( .A(x[754]), .B(y[754]), .Z(n3046) );
  XNOR U5920 ( .A(x[1122]), .B(y[1122]), .Z(n3047) );
  XOR U5921 ( .A(n3046), .B(n3047), .Z(n3049) );
  XNOR U5922 ( .A(n3048), .B(n3049), .Z(n2630) );
  XOR U5923 ( .A(n2631), .B(n2630), .Z(n2920) );
  XOR U5924 ( .A(x[730]), .B(y[730]), .Z(n4222) );
  XOR U5925 ( .A(x[726]), .B(y[726]), .Z(n4220) );
  XNOR U5926 ( .A(x[1446]), .B(y[1446]), .Z(n4221) );
  XOR U5927 ( .A(n4220), .B(n4221), .Z(n4223) );
  XNOR U5928 ( .A(n4222), .B(n4223), .Z(n1118) );
  XOR U5929 ( .A(x[740]), .B(y[740]), .Z(n4182) );
  XOR U5930 ( .A(x[738]), .B(y[738]), .Z(n4180) );
  XNOR U5931 ( .A(x[1444]), .B(y[1444]), .Z(n4181) );
  XOR U5932 ( .A(n4180), .B(n4181), .Z(n4183) );
  XNOR U5933 ( .A(n4182), .B(n4183), .Z(n1115) );
  XOR U5934 ( .A(x[736]), .B(y[736]), .Z(n4188) );
  XOR U5935 ( .A(x[734]), .B(y[734]), .Z(n4186) );
  XNOR U5936 ( .A(x[1114]), .B(y[1114]), .Z(n4187) );
  XOR U5937 ( .A(n4186), .B(n4187), .Z(n4189) );
  XOR U5938 ( .A(n4188), .B(n4189), .Z(n1116) );
  XNOR U5939 ( .A(n1115), .B(n1116), .Z(n1117) );
  XOR U5940 ( .A(n1118), .B(n1117), .Z(n2919) );
  XOR U5941 ( .A(x[752]), .B(y[752]), .Z(n3060) );
  XOR U5942 ( .A(x[748]), .B(y[748]), .Z(n3058) );
  XNOR U5943 ( .A(x[1442]), .B(y[1442]), .Z(n3059) );
  XOR U5944 ( .A(n3058), .B(n3059), .Z(n3061) );
  XNOR U5945 ( .A(n3060), .B(n3061), .Z(n2623) );
  XOR U5946 ( .A(x[329]), .B(y[329]), .Z(n3175) );
  XOR U5947 ( .A(x[331]), .B(y[331]), .Z(n3172) );
  XNOR U5948 ( .A(x[332]), .B(y[332]), .Z(n3173) );
  XNOR U5949 ( .A(n3172), .B(n3173), .Z(n3174) );
  XOR U5950 ( .A(n3175), .B(n3174), .Z(n2622) );
  XOR U5951 ( .A(n2623), .B(n2622), .Z(n2625) );
  XOR U5952 ( .A(x[744]), .B(y[744]), .Z(n3066) );
  XOR U5953 ( .A(x[742]), .B(y[742]), .Z(n3064) );
  XNOR U5954 ( .A(x[1118]), .B(y[1118]), .Z(n3065) );
  XOR U5955 ( .A(n3064), .B(n3065), .Z(n3067) );
  XNOR U5956 ( .A(n3066), .B(n3067), .Z(n2624) );
  XNOR U5957 ( .A(n2625), .B(n2624), .Z(n2918) );
  XOR U5958 ( .A(n2919), .B(n2918), .Z(n2921) );
  XOR U5959 ( .A(n2920), .B(n2921), .Z(n5125) );
  XOR U5960 ( .A(x[792]), .B(y[792]), .Z(n3559) );
  XOR U5961 ( .A(x[790]), .B(y[790]), .Z(n3556) );
  XNOR U5962 ( .A(x[1434]), .B(y[1434]), .Z(n3557) );
  XOR U5963 ( .A(n3559), .B(n3558), .Z(n4544) );
  XOR U5964 ( .A(x[788]), .B(y[788]), .Z(n2412) );
  XOR U5965 ( .A(x[784]), .B(y[784]), .Z(n2410) );
  XNOR U5966 ( .A(x[1134]), .B(y[1134]), .Z(n2411) );
  XOR U5967 ( .A(n2410), .B(n2411), .Z(n2413) );
  XOR U5968 ( .A(n2412), .B(n2413), .Z(n4545) );
  XNOR U5969 ( .A(n4544), .B(n4545), .Z(n4547) );
  XOR U5970 ( .A(x[780]), .B(y[780]), .Z(n2464) );
  XOR U5971 ( .A(x[778]), .B(y[778]), .Z(n2462) );
  XNOR U5972 ( .A(x[1436]), .B(y[1436]), .Z(n2463) );
  XOR U5973 ( .A(n2462), .B(n2463), .Z(n2465) );
  XNOR U5974 ( .A(n2464), .B(n2465), .Z(n4546) );
  XOR U5975 ( .A(n4547), .B(n4546), .Z(n4478) );
  XOR U5976 ( .A(x[576]), .B(y[576]), .Z(n1871) );
  XOR U5977 ( .A(x[574]), .B(y[574]), .Z(n1869) );
  XNOR U5978 ( .A(x[858]), .B(y[858]), .Z(n1870) );
  XOR U5979 ( .A(n1869), .B(n1870), .Z(n1872) );
  XNOR U5980 ( .A(n1871), .B(n1872), .Z(n1918) );
  XOR U5981 ( .A(x[1340]), .B(y[1340]), .Z(n1877) );
  XOR U5982 ( .A(x[1334]), .B(y[1334]), .Z(n1875) );
  XNOR U5983 ( .A(x[1346]), .B(y[1346]), .Z(n1876) );
  XOR U5984 ( .A(n1875), .B(n1876), .Z(n1878) );
  XOR U5985 ( .A(n1877), .B(n1878), .Z(n1919) );
  XNOR U5986 ( .A(n1918), .B(n1919), .Z(n1921) );
  XOR U5987 ( .A(x[572]), .B(y[572]), .Z(n4448) );
  XOR U5988 ( .A(x[570]), .B(y[570]), .Z(n4446) );
  XNOR U5989 ( .A(x[854]), .B(y[854]), .Z(n4447) );
  XOR U5990 ( .A(n4446), .B(n4447), .Z(n4449) );
  XNOR U5991 ( .A(n4448), .B(n4449), .Z(n1920) );
  XOR U5992 ( .A(n1921), .B(n1920), .Z(n4477) );
  XOR U5993 ( .A(x[776]), .B(y[776]), .Z(n4080) );
  XOR U5994 ( .A(x[774]), .B(y[774]), .Z(n4078) );
  XNOR U5995 ( .A(x[1130]), .B(y[1130]), .Z(n4079) );
  XOR U5996 ( .A(n4078), .B(n4079), .Z(n4081) );
  XNOR U5997 ( .A(n4080), .B(n4081), .Z(n2640) );
  XOR U5998 ( .A(x[772]), .B(y[772]), .Z(n4090) );
  XOR U5999 ( .A(x[770]), .B(y[770]), .Z(n4088) );
  XNOR U6000 ( .A(x[1438]), .B(y[1438]), .Z(n4089) );
  XOR U6001 ( .A(n4088), .B(n4089), .Z(n4091) );
  XOR U6002 ( .A(n4090), .B(n4091), .Z(n2641) );
  XNOR U6003 ( .A(n2640), .B(n2641), .Z(n2643) );
  XOR U6004 ( .A(x[766]), .B(y[766]), .Z(n4096) );
  XOR U6005 ( .A(x[762]), .B(y[762]), .Z(n4094) );
  XNOR U6006 ( .A(x[1126]), .B(y[1126]), .Z(n4095) );
  XOR U6007 ( .A(n4094), .B(n4095), .Z(n4097) );
  XNOR U6008 ( .A(n4096), .B(n4097), .Z(n2642) );
  XNOR U6009 ( .A(n2643), .B(n2642), .Z(n4476) );
  XOR U6010 ( .A(n4477), .B(n4476), .Z(n4479) );
  XOR U6011 ( .A(n4478), .B(n4479), .Z(n5123) );
  XOR U6012 ( .A(x[812]), .B(y[812]), .Z(n1000) );
  XOR U6013 ( .A(x[810]), .B(y[810]), .Z(n998) );
  XNOR U6014 ( .A(x[1430]), .B(y[1430]), .Z(n999) );
  XOR U6015 ( .A(n998), .B(n999), .Z(n1001) );
  XNOR U6016 ( .A(n1000), .B(n1001), .Z(n1214) );
  XOR U6017 ( .A(x[241]), .B(y[241]), .Z(n3437) );
  XOR U6018 ( .A(x[243]), .B(y[243]), .Z(n3434) );
  XNOR U6019 ( .A(x[428]), .B(y[428]), .Z(n3435) );
  XOR U6020 ( .A(n3437), .B(n3436), .Z(n1213) );
  XOR U6021 ( .A(n1214), .B(n1213), .Z(n1216) );
  XOR U6022 ( .A(x[808]), .B(y[808]), .Z(n1006) );
  XOR U6023 ( .A(x[806]), .B(y[806]), .Z(n1004) );
  XNOR U6024 ( .A(x[1142]), .B(y[1142]), .Z(n1005) );
  XOR U6025 ( .A(n1004), .B(n1005), .Z(n1007) );
  XNOR U6026 ( .A(n1006), .B(n1007), .Z(n1215) );
  XOR U6027 ( .A(n1216), .B(n1215), .Z(n4426) );
  XOR U6028 ( .A(x[802]), .B(y[802]), .Z(n4074) );
  XOR U6029 ( .A(x[798]), .B(y[798]), .Z(n4072) );
  XNOR U6030 ( .A(x[1432]), .B(y[1432]), .Z(n4073) );
  XOR U6031 ( .A(n4072), .B(n4073), .Z(n4075) );
  XNOR U6032 ( .A(n4074), .B(n4075), .Z(n4538) );
  XOR U6033 ( .A(x[257]), .B(y[257]), .Z(n3414) );
  XOR U6034 ( .A(x[259]), .B(y[259]), .Z(n3412) );
  XNOR U6035 ( .A(x[263]), .B(y[263]), .Z(n3413) );
  XOR U6036 ( .A(n3412), .B(n3413), .Z(n3415) );
  XOR U6037 ( .A(n3414), .B(n3415), .Z(n4539) );
  XNOR U6038 ( .A(n4538), .B(n4539), .Z(n4541) );
  XOR U6039 ( .A(x[796]), .B(y[796]), .Z(n3515) );
  XOR U6040 ( .A(x[794]), .B(y[794]), .Z(n3513) );
  XOR U6041 ( .A(x[1138]), .B(y[1138]), .Z(n3512) );
  XOR U6042 ( .A(n3513), .B(n3512), .Z(n3514) );
  XOR U6043 ( .A(n3515), .B(n3514), .Z(n4540) );
  XOR U6044 ( .A(n4541), .B(n4540), .Z(n4425) );
  XOR U6045 ( .A(x[1350]), .B(y[1350]), .Z(n1905) );
  XOR U6046 ( .A(x[1344]), .B(y[1344]), .Z(n1903) );
  XOR U6047 ( .A(x[1348]), .B(y[1348]), .Z(n1902) );
  XOR U6048 ( .A(n1903), .B(n1902), .Z(n1904) );
  XOR U6049 ( .A(n1905), .B(n1904), .Z(n4941) );
  XOR U6050 ( .A(x[1352]), .B(y[1352]), .Z(n1901) );
  XOR U6051 ( .A(x[1332]), .B(y[1332]), .Z(n1899) );
  XOR U6052 ( .A(x[1336]), .B(y[1336]), .Z(n1898) );
  XOR U6053 ( .A(n1899), .B(n1898), .Z(n1900) );
  XOR U6054 ( .A(n1901), .B(n1900), .Z(n4940) );
  XOR U6055 ( .A(n4941), .B(n4940), .Z(n4943) );
  XOR U6056 ( .A(x[1330]), .B(y[1330]), .Z(n1909) );
  XOR U6057 ( .A(x[1328]), .B(y[1328]), .Z(n1907) );
  XOR U6058 ( .A(x[1338]), .B(y[1338]), .Z(n1906) );
  XOR U6059 ( .A(n1907), .B(n1906), .Z(n1908) );
  XOR U6060 ( .A(n1909), .B(n1908), .Z(n4942) );
  XNOR U6061 ( .A(n4943), .B(n4942), .Z(n4424) );
  XOR U6062 ( .A(n4425), .B(n4424), .Z(n4427) );
  XNOR U6063 ( .A(n4426), .B(n4427), .Z(n5122) );
  XNOR U6064 ( .A(n5123), .B(n5122), .Z(n5124) );
  XNOR U6065 ( .A(n5125), .B(n5124), .Z(n5106) );
  XOR U6066 ( .A(n5107), .B(n5106), .Z(n1342) );
  XOR U6067 ( .A(x[1144]), .B(y[1144]), .Z(n3534) );
  XOR U6068 ( .A(x[1136]), .B(y[1136]), .Z(n3532) );
  XNOR U6069 ( .A(x[1140]), .B(y[1140]), .Z(n3533) );
  XOR U6070 ( .A(n3532), .B(n3533), .Z(n3535) );
  XNOR U6071 ( .A(n3534), .B(n3535), .Z(n4817) );
  XOR U6072 ( .A(x[1132]), .B(y[1132]), .Z(n3529) );
  XOR U6073 ( .A(x[1124]), .B(y[1124]), .Z(n3526) );
  XNOR U6074 ( .A(x[1128]), .B(y[1128]), .Z(n3527) );
  XNOR U6075 ( .A(n3526), .B(n3527), .Z(n3528) );
  XOR U6076 ( .A(n3529), .B(n3528), .Z(n4816) );
  XOR U6077 ( .A(n4817), .B(n4816), .Z(n4819) );
  XOR U6078 ( .A(x[1120]), .B(y[1120]), .Z(n3541) );
  XOR U6079 ( .A(x[1112]), .B(y[1112]), .Z(n3538) );
  XNOR U6080 ( .A(x[1116]), .B(y[1116]), .Z(n3539) );
  XNOR U6081 ( .A(n3538), .B(n3539), .Z(n3540) );
  XOR U6082 ( .A(n3541), .B(n3540), .Z(n4818) );
  XOR U6083 ( .A(n4819), .B(n4818), .Z(n1526) );
  XOR U6084 ( .A(x[1192]), .B(y[1192]), .Z(n3507) );
  XOR U6085 ( .A(x[1184]), .B(y[1184]), .Z(n3505) );
  XOR U6086 ( .A(x[1188]), .B(y[1188]), .Z(n3504) );
  XOR U6087 ( .A(n3505), .B(n3504), .Z(n3506) );
  XOR U6088 ( .A(n3507), .B(n3506), .Z(n2265) );
  XOR U6089 ( .A(x[276]), .B(y[276]), .Z(n4367) );
  XOR U6090 ( .A(x[270]), .B(y[270]), .Z(n4365) );
  XOR U6091 ( .A(x[272]), .B(y[272]), .Z(n4364) );
  XOR U6092 ( .A(n4365), .B(n4364), .Z(n4366) );
  XOR U6093 ( .A(n4367), .B(n4366), .Z(n2264) );
  XOR U6094 ( .A(n2265), .B(n2264), .Z(n2267) );
  XOR U6095 ( .A(x[1180]), .B(y[1180]), .Z(n3511) );
  XOR U6096 ( .A(x[1172]), .B(y[1172]), .Z(n3509) );
  XOR U6097 ( .A(x[1176]), .B(y[1176]), .Z(n3508) );
  XOR U6098 ( .A(n3509), .B(n3508), .Z(n3510) );
  XOR U6099 ( .A(n3511), .B(n3510), .Z(n2266) );
  XOR U6100 ( .A(n2267), .B(n2266), .Z(n1524) );
  XOR U6101 ( .A(x[1108]), .B(y[1108]), .Z(n3581) );
  XOR U6102 ( .A(x[1100]), .B(y[1100]), .Z(n3579) );
  XOR U6103 ( .A(x[1104]), .B(y[1104]), .Z(n3578) );
  XOR U6104 ( .A(n3579), .B(n3578), .Z(n3580) );
  XOR U6105 ( .A(n3581), .B(n3580), .Z(n2077) );
  XOR U6106 ( .A(x[1096]), .B(y[1096]), .Z(n3577) );
  XOR U6107 ( .A(x[1088]), .B(y[1088]), .Z(n3575) );
  XOR U6108 ( .A(x[1092]), .B(y[1092]), .Z(n3574) );
  XOR U6109 ( .A(n3575), .B(n3574), .Z(n3576) );
  XOR U6110 ( .A(n3577), .B(n3576), .Z(n2076) );
  XOR U6111 ( .A(n2077), .B(n2076), .Z(n2079) );
  XOR U6112 ( .A(x[1084]), .B(y[1084]), .Z(n3585) );
  XOR U6113 ( .A(x[1076]), .B(y[1076]), .Z(n3583) );
  XOR U6114 ( .A(x[1080]), .B(y[1080]), .Z(n3582) );
  XOR U6115 ( .A(n3583), .B(n3582), .Z(n3584) );
  XOR U6116 ( .A(n3585), .B(n3584), .Z(n2078) );
  XNOR U6117 ( .A(n2079), .B(n2078), .Z(n1523) );
  XNOR U6118 ( .A(n1524), .B(n1523), .Z(n1525) );
  XNOR U6119 ( .A(n1526), .B(n1525), .Z(n1756) );
  XOR U6120 ( .A(x[1010]), .B(y[1010]), .Z(n2400) );
  XOR U6121 ( .A(x[1006]), .B(y[1006]), .Z(n2398) );
  XNOR U6122 ( .A(x[1008]), .B(y[1008]), .Z(n2399) );
  XOR U6123 ( .A(n2398), .B(n2399), .Z(n2401) );
  XNOR U6124 ( .A(n2400), .B(n2401), .Z(n1538) );
  XOR U6125 ( .A(x[52]), .B(y[52]), .Z(n4109) );
  XOR U6126 ( .A(x[44]), .B(y[44]), .Z(n4107) );
  XOR U6127 ( .A(x[630]), .B(y[630]), .Z(n4106) );
  XOR U6128 ( .A(n4107), .B(n4106), .Z(n4108) );
  XOR U6129 ( .A(n4109), .B(n4108), .Z(n1537) );
  XOR U6130 ( .A(n1538), .B(n1537), .Z(n1539) );
  XOR U6131 ( .A(x[1004]), .B(y[1004]), .Z(n2406) );
  XOR U6132 ( .A(x[1000]), .B(y[1000]), .Z(n2404) );
  XNOR U6133 ( .A(x[1002]), .B(y[1002]), .Z(n2405) );
  XOR U6134 ( .A(n2404), .B(n2405), .Z(n2407) );
  XOR U6135 ( .A(n2406), .B(n2407), .Z(n1540) );
  XOR U6136 ( .A(n1539), .B(n1540), .Z(n1575) );
  XOR U6137 ( .A(x[1264]), .B(y[1264]), .Z(n4970) );
  XOR U6138 ( .A(x[1262]), .B(y[1262]), .Z(n4968) );
  XNOR U6139 ( .A(x[1390]), .B(y[1390]), .Z(n4969) );
  XOR U6140 ( .A(n4968), .B(n4969), .Z(n4971) );
  XNOR U6141 ( .A(n4970), .B(n4971), .Z(n2552) );
  XOR U6142 ( .A(x[1396]), .B(y[1396]), .Z(n4964) );
  XOR U6143 ( .A(x[1260]), .B(y[1260]), .Z(n4962) );
  XNOR U6144 ( .A(x[1394]), .B(y[1394]), .Z(n4963) );
  XOR U6145 ( .A(n4962), .B(n4963), .Z(n4965) );
  XOR U6146 ( .A(n4964), .B(n4965), .Z(n2553) );
  XNOR U6147 ( .A(n2552), .B(n2553), .Z(n2554) );
  XOR U6148 ( .A(x[1400]), .B(y[1400]), .Z(n4976) );
  XOR U6149 ( .A(x[1258]), .B(y[1258]), .Z(n4974) );
  XNOR U6150 ( .A(x[1398]), .B(y[1398]), .Z(n4975) );
  XOR U6151 ( .A(n4974), .B(n4975), .Z(n4977) );
  XOR U6152 ( .A(n4976), .B(n4977), .Z(n2555) );
  XOR U6153 ( .A(n2554), .B(n2555), .Z(n1573) );
  XOR U6154 ( .A(x[998]), .B(y[998]), .Z(n2434) );
  XOR U6155 ( .A(x[994]), .B(y[994]), .Z(n2432) );
  XNOR U6156 ( .A(x[996]), .B(y[996]), .Z(n2433) );
  XOR U6157 ( .A(n2432), .B(n2433), .Z(n2435) );
  XNOR U6158 ( .A(n2434), .B(n2435), .Z(n1495) );
  XOR U6159 ( .A(x[30]), .B(y[30]), .Z(n4112) );
  XOR U6160 ( .A(x[22]), .B(y[22]), .Z(n4110) );
  XNOR U6161 ( .A(x[24]), .B(y[24]), .Z(n4111) );
  XOR U6162 ( .A(n4110), .B(n4111), .Z(n4113) );
  XOR U6163 ( .A(n4112), .B(n4113), .Z(n1496) );
  XNOR U6164 ( .A(n1495), .B(n1496), .Z(n1498) );
  XOR U6165 ( .A(x[992]), .B(y[992]), .Z(n2440) );
  XOR U6166 ( .A(x[988]), .B(y[988]), .Z(n2438) );
  XNOR U6167 ( .A(x[990]), .B(y[990]), .Z(n2439) );
  XOR U6168 ( .A(n2438), .B(n2439), .Z(n2441) );
  XNOR U6169 ( .A(n2440), .B(n2441), .Z(n1497) );
  XNOR U6170 ( .A(n1498), .B(n1497), .Z(n1574) );
  XOR U6171 ( .A(n1573), .B(n1574), .Z(n1576) );
  XOR U6172 ( .A(n1575), .B(n1576), .Z(n1755) );
  XOR U6173 ( .A(n1756), .B(n1755), .Z(n1758) );
  XOR U6174 ( .A(x[986]), .B(y[986]), .Z(n2452) );
  XOR U6175 ( .A(x[982]), .B(y[982]), .Z(n2450) );
  XNOR U6176 ( .A(x[984]), .B(y[984]), .Z(n2451) );
  XOR U6177 ( .A(n2450), .B(n2451), .Z(n2453) );
  XNOR U6178 ( .A(n2452), .B(n2453), .Z(n1459) );
  XOR U6179 ( .A(x[980]), .B(y[980]), .Z(n2446) );
  XOR U6180 ( .A(x[976]), .B(y[976]), .Z(n2444) );
  XNOR U6181 ( .A(x[978]), .B(y[978]), .Z(n2445) );
  XOR U6182 ( .A(n2444), .B(n2445), .Z(n2447) );
  XOR U6183 ( .A(n2446), .B(n2447), .Z(n1460) );
  XNOR U6184 ( .A(n1459), .B(n1460), .Z(n1461) );
  XOR U6185 ( .A(x[974]), .B(y[974]), .Z(n2458) );
  XOR U6186 ( .A(x[970]), .B(y[970]), .Z(n2456) );
  XNOR U6187 ( .A(x[972]), .B(y[972]), .Z(n2457) );
  XOR U6188 ( .A(n2456), .B(n2457), .Z(n2459) );
  XOR U6189 ( .A(n2458), .B(n2459), .Z(n1462) );
  XOR U6190 ( .A(n1461), .B(n1462), .Z(n1549) );
  XOR U6191 ( .A(x[1272]), .B(y[1272]), .Z(n5090) );
  XOR U6192 ( .A(x[1270]), .B(y[1270]), .Z(n5088) );
  XNOR U6193 ( .A(x[1302]), .B(y[1302]), .Z(n5089) );
  XOR U6194 ( .A(n5088), .B(n5089), .Z(n5091) );
  XNOR U6195 ( .A(n5090), .B(n5091), .Z(n1103) );
  XOR U6196 ( .A(x[1268]), .B(y[1268]), .Z(n5084) );
  XOR U6197 ( .A(x[1304]), .B(y[1304]), .Z(n5082) );
  XNOR U6198 ( .A(x[1388]), .B(y[1388]), .Z(n5083) );
  XOR U6199 ( .A(n5082), .B(n5083), .Z(n5085) );
  XOR U6200 ( .A(n5084), .B(n5085), .Z(n1104) );
  XNOR U6201 ( .A(n1103), .B(n1104), .Z(n1105) );
  XOR U6202 ( .A(x[1266]), .B(y[1266]), .Z(n5096) );
  XOR U6203 ( .A(x[1306]), .B(y[1306]), .Z(n5094) );
  XNOR U6204 ( .A(x[1392]), .B(y[1392]), .Z(n5095) );
  XOR U6205 ( .A(n5094), .B(n5095), .Z(n5097) );
  XOR U6206 ( .A(n5096), .B(n5097), .Z(n1106) );
  XOR U6207 ( .A(n1105), .B(n1106), .Z(n1547) );
  XOR U6208 ( .A(x[968]), .B(y[968]), .Z(n1319) );
  XOR U6209 ( .A(x[964]), .B(y[964]), .Z(n1317) );
  XNOR U6210 ( .A(x[966]), .B(y[966]), .Z(n1318) );
  XOR U6211 ( .A(n1317), .B(n1318), .Z(n1320) );
  XNOR U6212 ( .A(n1319), .B(n1320), .Z(n1419) );
  XOR U6213 ( .A(x[962]), .B(y[962]), .Z(n1313) );
  XOR U6214 ( .A(x[958]), .B(y[958]), .Z(n1311) );
  XNOR U6215 ( .A(x[960]), .B(y[960]), .Z(n1312) );
  XOR U6216 ( .A(n1311), .B(n1312), .Z(n1314) );
  XOR U6217 ( .A(n1313), .B(n1314), .Z(n1420) );
  XNOR U6218 ( .A(n1419), .B(n1420), .Z(n1422) );
  XOR U6219 ( .A(x[956]), .B(y[956]), .Z(n1325) );
  XOR U6220 ( .A(x[952]), .B(y[952]), .Z(n1323) );
  XNOR U6221 ( .A(x[954]), .B(y[954]), .Z(n1324) );
  XOR U6222 ( .A(n1323), .B(n1324), .Z(n1326) );
  XNOR U6223 ( .A(n1325), .B(n1326), .Z(n1421) );
  XNOR U6224 ( .A(n1422), .B(n1421), .Z(n1548) );
  XOR U6225 ( .A(n1547), .B(n1548), .Z(n1550) );
  XOR U6226 ( .A(n1549), .B(n1550), .Z(n1757) );
  XOR U6227 ( .A(n1758), .B(n1757), .Z(n1341) );
  XNOR U6228 ( .A(n1342), .B(n1341), .Z(n1343) );
  XOR U6229 ( .A(n1344), .B(n1343), .Z(n920) );
  XNOR U6230 ( .A(n921), .B(n920), .Z(o[0]) );
  NANDN U6231 ( .A(n919), .B(n918), .Z(n923) );
  NAND U6232 ( .A(n921), .B(n920), .Z(n922) );
  AND U6233 ( .A(n923), .B(n922), .Z(n6930) );
  NANDN U6234 ( .A(n925), .B(n924), .Z(n929) );
  NANDN U6235 ( .A(n927), .B(n926), .Z(n928) );
  AND U6236 ( .A(n929), .B(n928), .Z(n6505) );
  NANDN U6237 ( .A(n931), .B(n930), .Z(n935) );
  NANDN U6238 ( .A(n933), .B(n932), .Z(n934) );
  NAND U6239 ( .A(n935), .B(n934), .Z(n6506) );
  XNOR U6240 ( .A(n6505), .B(n6506), .Z(n6508) );
  NANDN U6241 ( .A(n937), .B(n936), .Z(n941) );
  NANDN U6242 ( .A(n939), .B(n938), .Z(n940) );
  AND U6243 ( .A(n941), .B(n940), .Z(n6507) );
  XOR U6244 ( .A(n6508), .B(n6507), .Z(n7238) );
  NANDN U6245 ( .A(n943), .B(n942), .Z(n947) );
  NAND U6246 ( .A(n945), .B(n944), .Z(n946) );
  AND U6247 ( .A(n947), .B(n946), .Z(n6798) );
  NANDN U6248 ( .A(n949), .B(n948), .Z(n953) );
  NANDN U6249 ( .A(n951), .B(n950), .Z(n952) );
  AND U6250 ( .A(n953), .B(n952), .Z(n6797) );
  XOR U6251 ( .A(n6798), .B(n6797), .Z(n6800) );
  NANDN U6252 ( .A(n955), .B(n954), .Z(n959) );
  NANDN U6253 ( .A(n957), .B(n956), .Z(n958) );
  AND U6254 ( .A(n959), .B(n958), .Z(n6799) );
  XOR U6255 ( .A(n6800), .B(n6799), .Z(n7236) );
  NANDN U6256 ( .A(n961), .B(n960), .Z(n965) );
  NANDN U6257 ( .A(n963), .B(n962), .Z(n964) );
  AND U6258 ( .A(n965), .B(n964), .Z(n5928) );
  NANDN U6259 ( .A(n967), .B(n966), .Z(n971) );
  NANDN U6260 ( .A(n969), .B(n968), .Z(n970) );
  NAND U6261 ( .A(n971), .B(n970), .Z(n5929) );
  XNOR U6262 ( .A(n5928), .B(n5929), .Z(n5931) );
  NANDN U6263 ( .A(n973), .B(n972), .Z(n977) );
  NANDN U6264 ( .A(n975), .B(n974), .Z(n976) );
  AND U6265 ( .A(n977), .B(n976), .Z(n5930) );
  XNOR U6266 ( .A(n5931), .B(n5930), .Z(n7235) );
  XNOR U6267 ( .A(n7236), .B(n7235), .Z(n7237) );
  XNOR U6268 ( .A(n7238), .B(n7237), .Z(n7184) );
  NANDN U6269 ( .A(n979), .B(n978), .Z(n983) );
  NANDN U6270 ( .A(n981), .B(n980), .Z(n982) );
  AND U6271 ( .A(n983), .B(n982), .Z(n6328) );
  XOR U6272 ( .A(n6328), .B(n6327), .Z(n6330) );
  XOR U6273 ( .A(n6330), .B(n6329), .Z(n7225) );
  NANDN U6274 ( .A(n993), .B(n992), .Z(n997) );
  NANDN U6275 ( .A(n995), .B(n994), .Z(n996) );
  AND U6276 ( .A(n997), .B(n996), .Z(n6394) );
  NANDN U6277 ( .A(n999), .B(n998), .Z(n1003) );
  NANDN U6278 ( .A(n1001), .B(n1000), .Z(n1002) );
  AND U6279 ( .A(n1003), .B(n1002), .Z(n6393) );
  XOR U6280 ( .A(n6394), .B(n6393), .Z(n6396) );
  NANDN U6281 ( .A(n1005), .B(n1004), .Z(n1009) );
  NANDN U6282 ( .A(n1007), .B(n1006), .Z(n1008) );
  AND U6283 ( .A(n1009), .B(n1008), .Z(n6395) );
  XOR U6284 ( .A(n6396), .B(n6395), .Z(n7224) );
  NANDN U6285 ( .A(n1011), .B(n1010), .Z(n1015) );
  NANDN U6286 ( .A(n1013), .B(n1012), .Z(n1014) );
  AND U6287 ( .A(n1015), .B(n1014), .Z(n5922) );
  NANDN U6288 ( .A(n1017), .B(n1016), .Z(n1021) );
  NANDN U6289 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U6290 ( .A(n1021), .B(n1020), .Z(n5923) );
  XNOR U6291 ( .A(n5922), .B(n5923), .Z(n5925) );
  NANDN U6292 ( .A(n1023), .B(n1022), .Z(n1027) );
  NANDN U6293 ( .A(n1025), .B(n1024), .Z(n1026) );
  AND U6294 ( .A(n1027), .B(n1026), .Z(n5924) );
  XNOR U6295 ( .A(n5925), .B(n5924), .Z(n7223) );
  XOR U6296 ( .A(n7224), .B(n7223), .Z(n7226) );
  XOR U6297 ( .A(n7225), .B(n7226), .Z(n7183) );
  XOR U6298 ( .A(n7184), .B(n7183), .Z(n7185) );
  NANDN U6299 ( .A(n1029), .B(n1028), .Z(n1033) );
  NAND U6300 ( .A(n1031), .B(n1030), .Z(n1032) );
  NAND U6301 ( .A(n1033), .B(n1032), .Z(n7373) );
  NANDN U6302 ( .A(n1039), .B(n1038), .Z(n1043) );
  NANDN U6303 ( .A(n1041), .B(n1040), .Z(n1042) );
  NAND U6304 ( .A(n1043), .B(n1042), .Z(n6848) );
  XNOR U6305 ( .A(n6847), .B(n6848), .Z(n6849) );
  NANDN U6306 ( .A(n1045), .B(n1044), .Z(n1049) );
  NAND U6307 ( .A(n1047), .B(n1046), .Z(n1048) );
  NAND U6308 ( .A(n1049), .B(n1048), .Z(n6850) );
  XOR U6309 ( .A(n6849), .B(n6850), .Z(n7371) );
  NAND U6310 ( .A(n1055), .B(n1054), .Z(n1060) );
  IV U6311 ( .A(n1056), .Z(n1058) );
  NANDN U6312 ( .A(n1058), .B(n1057), .Z(n1059) );
  NAND U6313 ( .A(n1060), .B(n1059), .Z(n5949) );
  XNOR U6314 ( .A(n5948), .B(n5949), .Z(n5950) );
  XOR U6315 ( .A(n5950), .B(n5951), .Z(n7372) );
  XNOR U6316 ( .A(n7371), .B(n7372), .Z(n7374) );
  XOR U6317 ( .A(n7373), .B(n7374), .Z(n7186) );
  XOR U6318 ( .A(n7185), .B(n7186), .Z(n6869) );
  NANDN U6319 ( .A(n1066), .B(n1065), .Z(n1070) );
  NAND U6320 ( .A(n1068), .B(n1067), .Z(n1069) );
  NAND U6321 ( .A(n1070), .B(n1069), .Z(n6867) );
  NANDN U6322 ( .A(n1072), .B(n1071), .Z(n1076) );
  NANDN U6323 ( .A(n1074), .B(n1073), .Z(n1075) );
  AND U6324 ( .A(n1076), .B(n1075), .Z(n6695) );
  NANDN U6325 ( .A(n1078), .B(n1077), .Z(n1082) );
  NANDN U6326 ( .A(n1080), .B(n1079), .Z(n1081) );
  NAND U6327 ( .A(n1082), .B(n1081), .Z(n6696) );
  XNOR U6328 ( .A(n6695), .B(n6696), .Z(n6698) );
  NANDN U6329 ( .A(n1084), .B(n1083), .Z(n1088) );
  NANDN U6330 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U6331 ( .A(n1088), .B(n1087), .Z(n6697) );
  XOR U6332 ( .A(n6698), .B(n6697), .Z(n5919) );
  NANDN U6333 ( .A(n1090), .B(n1089), .Z(n1094) );
  NANDN U6334 ( .A(n1092), .B(n1091), .Z(n1093) );
  AND U6335 ( .A(n1094), .B(n1093), .Z(n6331) );
  XNOR U6336 ( .A(n6331), .B(n6332), .Z(n6334) );
  XOR U6337 ( .A(n6334), .B(n6333), .Z(n5917) );
  NANDN U6338 ( .A(n1104), .B(n1103), .Z(n1108) );
  NANDN U6339 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U6340 ( .A(n1108), .B(n1107), .Z(n5916) );
  XNOR U6341 ( .A(n5917), .B(n5916), .Z(n5918) );
  XNOR U6342 ( .A(n5919), .B(n5918), .Z(n6898) );
  NANDN U6343 ( .A(n1110), .B(n1109), .Z(n1114) );
  OR U6344 ( .A(n1112), .B(n1111), .Z(n1113) );
  NAND U6345 ( .A(n1114), .B(n1113), .Z(n6895) );
  NANDN U6346 ( .A(n1116), .B(n1115), .Z(n1120) );
  NAND U6347 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U6348 ( .A(n1120), .B(n1119), .Z(n6896) );
  XOR U6349 ( .A(n6895), .B(n6896), .Z(n6897) );
  XNOR U6350 ( .A(n6898), .B(n6897), .Z(n6868) );
  XOR U6351 ( .A(n6867), .B(n6868), .Z(n6870) );
  XOR U6352 ( .A(n6869), .B(n6870), .Z(n7042) );
  NANDN U6353 ( .A(n1122), .B(n1121), .Z(n1126) );
  NAND U6354 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U6355 ( .A(n1126), .B(n1125), .Z(n7040) );
  NAND U6356 ( .A(n1128), .B(n1127), .Z(n1132) );
  NAND U6357 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U6358 ( .A(n1132), .B(n1131), .Z(n7039) );
  XNOR U6359 ( .A(n7040), .B(n7039), .Z(n7041) );
  XOR U6360 ( .A(n7042), .B(n7041), .Z(n7035) );
  NANDN U6361 ( .A(n1138), .B(n1137), .Z(n1142) );
  NANDN U6362 ( .A(n1140), .B(n1139), .Z(n1141) );
  AND U6363 ( .A(n1142), .B(n1141), .Z(n6511) );
  NANDN U6364 ( .A(n1144), .B(n1143), .Z(n1148) );
  NANDN U6365 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U6366 ( .A(n1148), .B(n1147), .Z(n6512) );
  XNOR U6367 ( .A(n6511), .B(n6512), .Z(n6514) );
  NANDN U6368 ( .A(n1150), .B(n1149), .Z(n1154) );
  NANDN U6369 ( .A(n1152), .B(n1151), .Z(n1153) );
  AND U6370 ( .A(n1154), .B(n1153), .Z(n6513) );
  XOR U6371 ( .A(n6514), .B(n6513), .Z(n6726) );
  XNOR U6372 ( .A(n5605), .B(n5606), .Z(n5608) );
  NANDN U6373 ( .A(n1164), .B(n1163), .Z(n1168) );
  NANDN U6374 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U6375 ( .A(n1168), .B(n1167), .Z(n5607) );
  XOR U6376 ( .A(n5608), .B(n5607), .Z(n6724) );
  XNOR U6377 ( .A(n6724), .B(n6723), .Z(n6725) );
  XNOR U6378 ( .A(n6726), .B(n6725), .Z(n7379) );
  XNOR U6379 ( .A(n7380), .B(n7379), .Z(n7382) );
  NANDN U6380 ( .A(n1174), .B(n1173), .Z(n1178) );
  NANDN U6381 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U6382 ( .A(n1178), .B(n1177), .Z(n6481) );
  NANDN U6383 ( .A(n1180), .B(n1179), .Z(n1184) );
  NANDN U6384 ( .A(n1182), .B(n1181), .Z(n1183) );
  NAND U6385 ( .A(n1184), .B(n1183), .Z(n6482) );
  XNOR U6386 ( .A(n6481), .B(n6482), .Z(n6484) );
  NANDN U6387 ( .A(n1186), .B(n1185), .Z(n1190) );
  NANDN U6388 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U6389 ( .A(n1190), .B(n1189), .Z(n6483) );
  XOR U6390 ( .A(n6484), .B(n6483), .Z(n7162) );
  NANDN U6391 ( .A(n1196), .B(n1195), .Z(n1200) );
  NANDN U6392 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U6393 ( .A(n1200), .B(n1199), .Z(n6468) );
  XNOR U6394 ( .A(n6467), .B(n6468), .Z(n6470) );
  NANDN U6395 ( .A(n1202), .B(n1201), .Z(n1206) );
  NANDN U6396 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U6397 ( .A(n1206), .B(n1205), .Z(n6469) );
  XOR U6398 ( .A(n6470), .B(n6469), .Z(n7160) );
  NANDN U6399 ( .A(n1208), .B(n1207), .Z(n1212) );
  NAND U6400 ( .A(n1210), .B(n1209), .Z(n1211) );
  NAND U6401 ( .A(n1212), .B(n1211), .Z(n7159) );
  XNOR U6402 ( .A(n7160), .B(n7159), .Z(n7161) );
  XNOR U6403 ( .A(n7162), .B(n7161), .Z(n7381) );
  XOR U6404 ( .A(n7382), .B(n7381), .Z(n6891) );
  NANDN U6405 ( .A(n1218), .B(n1217), .Z(n1222) );
  NAND U6406 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U6407 ( .A(n1222), .B(n1221), .Z(n7386) );
  NANDN U6408 ( .A(n1224), .B(n1223), .Z(n1228) );
  NAND U6409 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U6410 ( .A(n1228), .B(n1227), .Z(n7385) );
  XNOR U6411 ( .A(n7386), .B(n7385), .Z(n7387) );
  XNOR U6412 ( .A(n7388), .B(n7387), .Z(n7431) );
  NANDN U6413 ( .A(n1230), .B(n1229), .Z(n1234) );
  NANDN U6414 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U6415 ( .A(n1234), .B(n1233), .Z(n6683) );
  NANDN U6416 ( .A(n1236), .B(n1235), .Z(n1240) );
  NANDN U6417 ( .A(n1238), .B(n1237), .Z(n1239) );
  NAND U6418 ( .A(n1240), .B(n1239), .Z(n6684) );
  XNOR U6419 ( .A(n6683), .B(n6684), .Z(n6686) );
  NANDN U6420 ( .A(n1242), .B(n1241), .Z(n1246) );
  NANDN U6421 ( .A(n1244), .B(n1243), .Z(n1245) );
  AND U6422 ( .A(n1246), .B(n1245), .Z(n6685) );
  XOR U6423 ( .A(n6686), .B(n6685), .Z(n7428) );
  NANDN U6424 ( .A(n1248), .B(n1247), .Z(n1252) );
  NANDN U6425 ( .A(n1250), .B(n1249), .Z(n1251) );
  AND U6426 ( .A(n1252), .B(n1251), .Z(n6241) );
  NANDN U6427 ( .A(n1254), .B(n1253), .Z(n1258) );
  NANDN U6428 ( .A(n1256), .B(n1255), .Z(n1257) );
  NAND U6429 ( .A(n1258), .B(n1257), .Z(n6242) );
  XNOR U6430 ( .A(n6241), .B(n6242), .Z(n6244) );
  NANDN U6431 ( .A(n1260), .B(n1259), .Z(n1264) );
  NANDN U6432 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U6433 ( .A(n1264), .B(n1263), .Z(n6243) );
  XOR U6434 ( .A(n6244), .B(n6243), .Z(n7426) );
  NANDN U6435 ( .A(n1266), .B(n1265), .Z(n1270) );
  NANDN U6436 ( .A(n1268), .B(n1267), .Z(n1269) );
  AND U6437 ( .A(n1270), .B(n1269), .Z(n6499) );
  NANDN U6438 ( .A(n1272), .B(n1271), .Z(n1276) );
  NANDN U6439 ( .A(n1274), .B(n1273), .Z(n1275) );
  NAND U6440 ( .A(n1276), .B(n1275), .Z(n6500) );
  XNOR U6441 ( .A(n6499), .B(n6500), .Z(n6502) );
  NANDN U6442 ( .A(n1278), .B(n1277), .Z(n1282) );
  NANDN U6443 ( .A(n1280), .B(n1279), .Z(n1281) );
  AND U6444 ( .A(n1282), .B(n1281), .Z(n6501) );
  XNOR U6445 ( .A(n6502), .B(n6501), .Z(n7425) );
  XNOR U6446 ( .A(n7426), .B(n7425), .Z(n7427) );
  XOR U6447 ( .A(n7428), .B(n7427), .Z(n7432) );
  XNOR U6448 ( .A(n7431), .B(n7432), .Z(n7434) );
  XNOR U6449 ( .A(n5954), .B(n5955), .Z(n5957) );
  XOR U6450 ( .A(n5957), .B(n5956), .Z(n7418) );
  NANDN U6451 ( .A(n1300), .B(n1299), .Z(n1304) );
  NANDN U6452 ( .A(n1302), .B(n1301), .Z(n1303) );
  NAND U6453 ( .A(n1304), .B(n1303), .Z(n6802) );
  XNOR U6454 ( .A(n6801), .B(n6802), .Z(n6804) );
  NANDN U6455 ( .A(n1306), .B(n1305), .Z(n1310) );
  NANDN U6456 ( .A(n1308), .B(n1307), .Z(n1309) );
  AND U6457 ( .A(n1310), .B(n1309), .Z(n6803) );
  XOR U6458 ( .A(n6804), .B(n6803), .Z(n7416) );
  NANDN U6459 ( .A(n1312), .B(n1311), .Z(n1316) );
  NANDN U6460 ( .A(n1314), .B(n1313), .Z(n1315) );
  AND U6461 ( .A(n1316), .B(n1315), .Z(n5599) );
  NANDN U6462 ( .A(n1318), .B(n1317), .Z(n1322) );
  NANDN U6463 ( .A(n1320), .B(n1319), .Z(n1321) );
  NAND U6464 ( .A(n1322), .B(n1321), .Z(n5600) );
  XNOR U6465 ( .A(n5599), .B(n5600), .Z(n5602) );
  NANDN U6466 ( .A(n1324), .B(n1323), .Z(n1328) );
  NANDN U6467 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U6468 ( .A(n1328), .B(n1327), .Z(n5601) );
  XNOR U6469 ( .A(n5602), .B(n5601), .Z(n7415) );
  XNOR U6470 ( .A(n7416), .B(n7415), .Z(n7417) );
  XNOR U6471 ( .A(n7418), .B(n7417), .Z(n7433) );
  XOR U6472 ( .A(n7434), .B(n7433), .Z(n6890) );
  NANDN U6473 ( .A(n1330), .B(n1329), .Z(n1334) );
  NANDN U6474 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U6475 ( .A(n1334), .B(n1333), .Z(n6889) );
  XOR U6476 ( .A(n6890), .B(n6889), .Z(n6892) );
  XOR U6477 ( .A(n6891), .B(n6892), .Z(n7034) );
  NANDN U6478 ( .A(n1336), .B(n1335), .Z(n1340) );
  OR U6479 ( .A(n1338), .B(n1337), .Z(n1339) );
  AND U6480 ( .A(n1340), .B(n1339), .Z(n7033) );
  XOR U6481 ( .A(n7034), .B(n7033), .Z(n7036) );
  XOR U6482 ( .A(n7035), .B(n7036), .Z(n5287) );
  NANDN U6483 ( .A(n1342), .B(n1341), .Z(n1346) );
  NAND U6484 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U6485 ( .A(n1346), .B(n1345), .Z(n5286) );
  XNOR U6486 ( .A(n5287), .B(n5286), .Z(n5288) );
  NANDN U6487 ( .A(n1348), .B(n1347), .Z(n1352) );
  OR U6488 ( .A(n1350), .B(n1349), .Z(n1351) );
  NAND U6489 ( .A(n1352), .B(n1351), .Z(n5289) );
  XNOR U6490 ( .A(n5288), .B(n5289), .Z(n6929) );
  XNOR U6491 ( .A(n6930), .B(n6929), .Z(n6932) );
  NANDN U6492 ( .A(n1354), .B(n1353), .Z(n1358) );
  OR U6493 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U6494 ( .A(n1358), .B(n1357), .Z(n6620) );
  NANDN U6495 ( .A(n1360), .B(n1359), .Z(n1364) );
  NANDN U6496 ( .A(n1362), .B(n1361), .Z(n1363) );
  AND U6497 ( .A(n1364), .B(n1363), .Z(n6617) );
  NANDN U6498 ( .A(n1366), .B(n1365), .Z(n1370) );
  NAND U6499 ( .A(n1368), .B(n1367), .Z(n1369) );
  AND U6500 ( .A(n1370), .B(n1369), .Z(n6634) );
  NANDN U6501 ( .A(n1372), .B(n1371), .Z(n1376) );
  NANDN U6502 ( .A(n1374), .B(n1373), .Z(n1375) );
  AND U6503 ( .A(n1376), .B(n1375), .Z(n6633) );
  XOR U6504 ( .A(n6634), .B(n6633), .Z(n6636) );
  NANDN U6505 ( .A(n1378), .B(n1377), .Z(n1382) );
  NANDN U6506 ( .A(n1380), .B(n1379), .Z(n1381) );
  AND U6507 ( .A(n1382), .B(n1381), .Z(n6635) );
  XOR U6508 ( .A(n6636), .B(n6635), .Z(n6238) );
  NANDN U6509 ( .A(n1384), .B(n1383), .Z(n1388) );
  NANDN U6510 ( .A(n1386), .B(n1385), .Z(n1387) );
  AND U6511 ( .A(n1388), .B(n1387), .Z(n6033) );
  NANDN U6512 ( .A(n1390), .B(n1389), .Z(n1394) );
  NANDN U6513 ( .A(n1392), .B(n1391), .Z(n1393) );
  AND U6514 ( .A(n1394), .B(n1393), .Z(n6032) );
  XOR U6515 ( .A(n6033), .B(n6032), .Z(n6035) );
  XOR U6516 ( .A(n6035), .B(n6034), .Z(n6236) );
  XNOR U6517 ( .A(n6236), .B(n6235), .Z(n6237) );
  XOR U6518 ( .A(n6238), .B(n6237), .Z(n6618) );
  XNOR U6519 ( .A(n6617), .B(n6618), .Z(n6619) );
  XOR U6520 ( .A(n6620), .B(n6619), .Z(n7404) );
  NANDN U6521 ( .A(n1404), .B(n1403), .Z(n1408) );
  OR U6522 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U6523 ( .A(n1408), .B(n1407), .Z(n6586) );
  NANDN U6524 ( .A(n1414), .B(n1413), .Z(n1418) );
  NAND U6525 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U6526 ( .A(n1418), .B(n1417), .Z(n5732) );
  NANDN U6527 ( .A(n1420), .B(n1419), .Z(n1424) );
  NAND U6528 ( .A(n1422), .B(n1421), .Z(n1423) );
  NAND U6529 ( .A(n1424), .B(n1423), .Z(n5731) );
  XOR U6530 ( .A(n5732), .B(n5731), .Z(n5734) );
  XOR U6531 ( .A(n5733), .B(n5734), .Z(n6584) );
  NANDN U6532 ( .A(n1426), .B(n1425), .Z(n1430) );
  OR U6533 ( .A(n1428), .B(n1427), .Z(n1429) );
  NAND U6534 ( .A(n1430), .B(n1429), .Z(n6583) );
  XNOR U6535 ( .A(n6584), .B(n6583), .Z(n6585) );
  XNOR U6536 ( .A(n6586), .B(n6585), .Z(n7403) );
  NAND U6537 ( .A(n1432), .B(n1431), .Z(n1436) );
  NAND U6538 ( .A(n1434), .B(n1433), .Z(n1435) );
  NAND U6539 ( .A(n1436), .B(n1435), .Z(n7406) );
  NANDN U6540 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U6541 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U6542 ( .A(n1442), .B(n1441), .Z(n7048) );
  NANDN U6543 ( .A(n1444), .B(n1443), .Z(n1448) );
  NANDN U6544 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U6545 ( .A(n1448), .B(n1447), .Z(n7045) );
  NANDN U6546 ( .A(n1450), .B(n1449), .Z(n1454) );
  NAND U6547 ( .A(n1452), .B(n1451), .Z(n1453) );
  AND U6548 ( .A(n1454), .B(n1453), .Z(n5740) );
  NANDN U6549 ( .A(n1460), .B(n1459), .Z(n1464) );
  NANDN U6550 ( .A(n1462), .B(n1461), .Z(n1463) );
  NAND U6551 ( .A(n1464), .B(n1463), .Z(n5737) );
  XNOR U6552 ( .A(n5738), .B(n5737), .Z(n5739) );
  XOR U6553 ( .A(n5740), .B(n5739), .Z(n7046) );
  XNOR U6554 ( .A(n7045), .B(n7046), .Z(n7047) );
  XOR U6555 ( .A(n7048), .B(n7047), .Z(n5417) );
  NANDN U6556 ( .A(n1466), .B(n1465), .Z(n1470) );
  NANDN U6557 ( .A(n1468), .B(n1467), .Z(n1469) );
  AND U6558 ( .A(n1470), .B(n1469), .Z(n7054) );
  NANDN U6559 ( .A(n1472), .B(n1471), .Z(n1476) );
  NANDN U6560 ( .A(n1474), .B(n1473), .Z(n1475) );
  AND U6561 ( .A(n1476), .B(n1475), .Z(n7051) );
  NANDN U6562 ( .A(n1478), .B(n1477), .Z(n1482) );
  NAND U6563 ( .A(n1480), .B(n1479), .Z(n1481) );
  AND U6564 ( .A(n1482), .B(n1481), .Z(n6069) );
  NANDN U6565 ( .A(n1484), .B(n1483), .Z(n1488) );
  NANDN U6566 ( .A(n1486), .B(n1485), .Z(n1487) );
  NAND U6567 ( .A(n1488), .B(n1487), .Z(n6070) );
  NANDN U6568 ( .A(n1490), .B(n1489), .Z(n1494) );
  NAND U6569 ( .A(n1492), .B(n1491), .Z(n1493) );
  AND U6570 ( .A(n1494), .B(n1493), .Z(n6071) );
  XOR U6571 ( .A(n6072), .B(n6071), .Z(n5567) );
  NANDN U6572 ( .A(n1496), .B(n1495), .Z(n1500) );
  NAND U6573 ( .A(n1498), .B(n1497), .Z(n1499) );
  AND U6574 ( .A(n1500), .B(n1499), .Z(n5565) );
  NANDN U6575 ( .A(n1506), .B(n1505), .Z(n1510) );
  NAND U6576 ( .A(n1508), .B(n1507), .Z(n1509) );
  NAND U6577 ( .A(n1510), .B(n1509), .Z(n5833) );
  NANDN U6578 ( .A(n1512), .B(n1511), .Z(n1516) );
  NANDN U6579 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U6580 ( .A(n1516), .B(n1515), .Z(n5834) );
  XNOR U6581 ( .A(n5835), .B(n5834), .Z(n5564) );
  XNOR U6582 ( .A(n5565), .B(n5564), .Z(n5566) );
  XOR U6583 ( .A(n5567), .B(n5566), .Z(n7052) );
  XNOR U6584 ( .A(n7051), .B(n7052), .Z(n7053) );
  XOR U6585 ( .A(n7054), .B(n7053), .Z(n5415) );
  NANDN U6586 ( .A(n1518), .B(n1517), .Z(n1522) );
  NANDN U6587 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U6588 ( .A(n1522), .B(n1521), .Z(n6950) );
  NANDN U6589 ( .A(n1524), .B(n1523), .Z(n1528) );
  NANDN U6590 ( .A(n1526), .B(n1525), .Z(n1527) );
  AND U6591 ( .A(n1528), .B(n1527), .Z(n6947) );
  XNOR U6592 ( .A(n7206), .B(n7205), .Z(n7207) );
  XOR U6593 ( .A(n7208), .B(n7207), .Z(n6948) );
  XNOR U6594 ( .A(n6947), .B(n6948), .Z(n6949) );
  XNOR U6595 ( .A(n6950), .B(n6949), .Z(n5414) );
  XNOR U6596 ( .A(n5415), .B(n5414), .Z(n5416) );
  XOR U6597 ( .A(n5417), .B(n5416), .Z(n6820) );
  XNOR U6598 ( .A(n6819), .B(n6820), .Z(n6821) );
  NANDN U6599 ( .A(n1542), .B(n1541), .Z(n1546) );
  OR U6600 ( .A(n1544), .B(n1543), .Z(n1545) );
  AND U6601 ( .A(n1546), .B(n1545), .Z(n6956) );
  NANDN U6602 ( .A(n1552), .B(n1551), .Z(n1556) );
  NANDN U6603 ( .A(n1554), .B(n1553), .Z(n1555) );
  AND U6604 ( .A(n1556), .B(n1555), .Z(n5728) );
  NANDN U6605 ( .A(n1562), .B(n1561), .Z(n1566) );
  NAND U6606 ( .A(n1564), .B(n1563), .Z(n1565) );
  NAND U6607 ( .A(n1566), .B(n1565), .Z(n5725) );
  XNOR U6608 ( .A(n5726), .B(n5725), .Z(n5727) );
  XOR U6609 ( .A(n5728), .B(n5727), .Z(n6954) );
  XNOR U6610 ( .A(n6953), .B(n6954), .Z(n6955) );
  XOR U6611 ( .A(n6956), .B(n6955), .Z(n5423) );
  NANDN U6612 ( .A(n1568), .B(n1567), .Z(n1572) );
  NANDN U6613 ( .A(n1570), .B(n1569), .Z(n1571) );
  AND U6614 ( .A(n1572), .B(n1571), .Z(n7008) );
  NANDN U6615 ( .A(n1582), .B(n1581), .Z(n1586) );
  NANDN U6616 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U6617 ( .A(n1586), .B(n1585), .Z(n7135) );
  XOR U6618 ( .A(n7136), .B(n7135), .Z(n7138) );
  NANDN U6619 ( .A(n1588), .B(n1587), .Z(n1592) );
  NANDN U6620 ( .A(n1590), .B(n1589), .Z(n1591) );
  AND U6621 ( .A(n1592), .B(n1591), .Z(n7137) );
  XOR U6622 ( .A(n7138), .B(n7137), .Z(n5704) );
  NANDN U6623 ( .A(n1594), .B(n1593), .Z(n1598) );
  NANDN U6624 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U6625 ( .A(n1598), .B(n1597), .Z(n5851) );
  NANDN U6626 ( .A(n1600), .B(n1599), .Z(n1604) );
  NANDN U6627 ( .A(n1602), .B(n1601), .Z(n1603) );
  AND U6628 ( .A(n1604), .B(n1603), .Z(n5850) );
  XOR U6629 ( .A(n5851), .B(n5850), .Z(n5853) );
  NANDN U6630 ( .A(n1606), .B(n1605), .Z(n1610) );
  NANDN U6631 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U6632 ( .A(n1610), .B(n1609), .Z(n5852) );
  XOR U6633 ( .A(n5853), .B(n5852), .Z(n5702) );
  XNOR U6634 ( .A(n5702), .B(n5701), .Z(n5703) );
  XOR U6635 ( .A(n5704), .B(n5703), .Z(n7006) );
  XNOR U6636 ( .A(n7005), .B(n7006), .Z(n7007) );
  XOR U6637 ( .A(n7008), .B(n7007), .Z(n5421) );
  NANDN U6638 ( .A(n1616), .B(n1615), .Z(n1620) );
  NANDN U6639 ( .A(n1618), .B(n1617), .Z(n1619) );
  AND U6640 ( .A(n1620), .B(n1619), .Z(n7014) );
  NANDN U6641 ( .A(n1622), .B(n1621), .Z(n1626) );
  OR U6642 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U6643 ( .A(n1626), .B(n1625), .Z(n7011) );
  XNOR U6644 ( .A(n5696), .B(n5695), .Z(n5697) );
  XOR U6645 ( .A(n5698), .B(n5697), .Z(n7012) );
  XNOR U6646 ( .A(n7011), .B(n7012), .Z(n7013) );
  XNOR U6647 ( .A(n7014), .B(n7013), .Z(n5420) );
  XNOR U6648 ( .A(n5421), .B(n5420), .Z(n5422) );
  XOR U6649 ( .A(n5423), .B(n5422), .Z(n6822) );
  XNOR U6650 ( .A(n6821), .B(n6822), .Z(n7439) );
  NANDN U6651 ( .A(n1644), .B(n1643), .Z(n1648) );
  NAND U6652 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U6653 ( .A(n1648), .B(n1647), .Z(n5839) );
  NANDN U6654 ( .A(n1650), .B(n1649), .Z(n1654) );
  NANDN U6655 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U6656 ( .A(n1654), .B(n1653), .Z(n5840) );
  XOR U6657 ( .A(n5841), .B(n5840), .Z(n5435) );
  NANDN U6658 ( .A(n1656), .B(n1655), .Z(n1660) );
  NANDN U6659 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U6660 ( .A(n1660), .B(n1659), .Z(n6089) );
  NANDN U6661 ( .A(n1662), .B(n1661), .Z(n1666) );
  NANDN U6662 ( .A(n1664), .B(n1663), .Z(n1665) );
  NAND U6663 ( .A(n1666), .B(n1665), .Z(n6090) );
  NANDN U6664 ( .A(n1668), .B(n1667), .Z(n1672) );
  NANDN U6665 ( .A(n1670), .B(n1669), .Z(n1671) );
  AND U6666 ( .A(n1672), .B(n1671), .Z(n6091) );
  XOR U6667 ( .A(n6092), .B(n6091), .Z(n5433) );
  NANDN U6668 ( .A(n1674), .B(n1673), .Z(n1678) );
  NAND U6669 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U6670 ( .A(n1678), .B(n1677), .Z(n5432) );
  XNOR U6671 ( .A(n5433), .B(n5432), .Z(n5434) );
  XNOR U6672 ( .A(n5435), .B(n5434), .Z(n6305) );
  NANDN U6673 ( .A(n1680), .B(n1679), .Z(n1684) );
  NANDN U6674 ( .A(n1682), .B(n1681), .Z(n1683) );
  AND U6675 ( .A(n1684), .B(n1683), .Z(n6229) );
  NANDN U6676 ( .A(n1686), .B(n1685), .Z(n1690) );
  NAND U6677 ( .A(n1688), .B(n1687), .Z(n1689) );
  NAND U6678 ( .A(n1690), .B(n1689), .Z(n6230) );
  XNOR U6679 ( .A(n6229), .B(n6230), .Z(n6232) );
  NANDN U6680 ( .A(n1692), .B(n1691), .Z(n1696) );
  NANDN U6681 ( .A(n1694), .B(n1693), .Z(n1695) );
  AND U6682 ( .A(n1696), .B(n1695), .Z(n6231) );
  XOR U6683 ( .A(n6232), .B(n6231), .Z(n5967) );
  NANDN U6684 ( .A(n1702), .B(n1701), .Z(n1706) );
  NAND U6685 ( .A(n1704), .B(n1703), .Z(n1705) );
  NAND U6686 ( .A(n1706), .B(n1705), .Z(n6776) );
  XNOR U6687 ( .A(n6775), .B(n6776), .Z(n6778) );
  XOR U6688 ( .A(n6778), .B(n6777), .Z(n5965) );
  NANDN U6689 ( .A(n1712), .B(n1711), .Z(n1716) );
  NAND U6690 ( .A(n1714), .B(n1713), .Z(n1715) );
  NAND U6691 ( .A(n1716), .B(n1715), .Z(n5964) );
  XNOR U6692 ( .A(n5965), .B(n5964), .Z(n5966) );
  XOR U6693 ( .A(n5967), .B(n5966), .Z(n6306) );
  XNOR U6694 ( .A(n6305), .B(n6306), .Z(n6308) );
  NANDN U6695 ( .A(n1718), .B(n1717), .Z(n1722) );
  NANDN U6696 ( .A(n1720), .B(n1719), .Z(n1721) );
  AND U6697 ( .A(n1722), .B(n1721), .Z(n6013) );
  NANDN U6698 ( .A(n1724), .B(n1723), .Z(n1728) );
  NANDN U6699 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U6700 ( .A(n1728), .B(n1727), .Z(n6012) );
  XOR U6701 ( .A(n6013), .B(n6012), .Z(n6015) );
  NANDN U6702 ( .A(n1730), .B(n1729), .Z(n1734) );
  NANDN U6703 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U6704 ( .A(n1734), .B(n1733), .Z(n6014) );
  XOR U6705 ( .A(n6015), .B(n6014), .Z(n6029) );
  NANDN U6706 ( .A(n1736), .B(n1735), .Z(n1740) );
  NANDN U6707 ( .A(n1738), .B(n1737), .Z(n1739) );
  AND U6708 ( .A(n1740), .B(n1739), .Z(n6748) );
  XOR U6709 ( .A(n6748), .B(n6747), .Z(n6750) );
  NANDN U6710 ( .A(n1746), .B(n1745), .Z(n1750) );
  NANDN U6711 ( .A(n1748), .B(n1747), .Z(n1749) );
  AND U6712 ( .A(n1750), .B(n1749), .Z(n6749) );
  XOR U6713 ( .A(n6750), .B(n6749), .Z(n6027) );
  XNOR U6714 ( .A(n6027), .B(n6026), .Z(n6028) );
  XNOR U6715 ( .A(n6029), .B(n6028), .Z(n6307) );
  XOR U6716 ( .A(n6308), .B(n6307), .Z(n7062) );
  XNOR U6717 ( .A(n7062), .B(n7061), .Z(n7064) );
  NANDN U6718 ( .A(n1760), .B(n1759), .Z(n1764) );
  NANDN U6719 ( .A(n1762), .B(n1761), .Z(n1763) );
  AND U6720 ( .A(n1764), .B(n1763), .Z(n6568) );
  NANDN U6721 ( .A(n1766), .B(n1765), .Z(n1770) );
  OR U6722 ( .A(n1768), .B(n1767), .Z(n1769) );
  AND U6723 ( .A(n1770), .B(n1769), .Z(n6566) );
  NANDN U6724 ( .A(n1772), .B(n1771), .Z(n1776) );
  OR U6725 ( .A(n1774), .B(n1773), .Z(n1775) );
  NAND U6726 ( .A(n1776), .B(n1775), .Z(n6565) );
  XNOR U6727 ( .A(n6566), .B(n6565), .Z(n6567) );
  XNOR U6728 ( .A(n6568), .B(n6567), .Z(n7063) );
  XOR U6729 ( .A(n7064), .B(n7063), .Z(n6878) );
  NANDN U6730 ( .A(n1778), .B(n1777), .Z(n1782) );
  NANDN U6731 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U6732 ( .A(n1782), .B(n1781), .Z(n6017) );
  NANDN U6733 ( .A(n1784), .B(n1783), .Z(n1788) );
  NAND U6734 ( .A(n1786), .B(n1785), .Z(n1787) );
  NAND U6735 ( .A(n1788), .B(n1787), .Z(n5942) );
  NANDN U6736 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U6737 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U6738 ( .A(n1794), .B(n1793), .Z(n6289) );
  NANDN U6739 ( .A(n1796), .B(n1795), .Z(n1800) );
  NAND U6740 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U6741 ( .A(n1800), .B(n1799), .Z(n6290) );
  XNOR U6742 ( .A(n6289), .B(n6290), .Z(n6291) );
  NANDN U6743 ( .A(n1802), .B(n1801), .Z(n1806) );
  NANDN U6744 ( .A(n1804), .B(n1803), .Z(n1805) );
  NAND U6745 ( .A(n1806), .B(n1805), .Z(n6292) );
  XOR U6746 ( .A(n6291), .B(n6292), .Z(n5940) );
  XOR U6747 ( .A(n5940), .B(n5941), .Z(n5943) );
  XOR U6748 ( .A(n5942), .B(n5943), .Z(n6016) );
  XOR U6749 ( .A(n6017), .B(n6016), .Z(n6019) );
  NANDN U6750 ( .A(n1812), .B(n1811), .Z(n1816) );
  NAND U6751 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U6752 ( .A(n1816), .B(n1815), .Z(n6433) );
  NANDN U6753 ( .A(n1818), .B(n1817), .Z(n1822) );
  NAND U6754 ( .A(n1820), .B(n1819), .Z(n1821) );
  AND U6755 ( .A(n1822), .B(n1821), .Z(n5845) );
  NANDN U6756 ( .A(n1824), .B(n1823), .Z(n1828) );
  NANDN U6757 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U6758 ( .A(n1828), .B(n1827), .Z(n5844) );
  XOR U6759 ( .A(n5845), .B(n5844), .Z(n5847) );
  NANDN U6760 ( .A(n1830), .B(n1829), .Z(n1834) );
  NANDN U6761 ( .A(n1832), .B(n1831), .Z(n1833) );
  AND U6762 ( .A(n1834), .B(n1833), .Z(n5846) );
  XOR U6763 ( .A(n5847), .B(n5846), .Z(n6432) );
  NANDN U6764 ( .A(n1836), .B(n1835), .Z(n1840) );
  NANDN U6765 ( .A(n1838), .B(n1837), .Z(n1839) );
  AND U6766 ( .A(n1840), .B(n1839), .Z(n5585) );
  NANDN U6767 ( .A(n1842), .B(n1841), .Z(n1846) );
  NANDN U6768 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U6769 ( .A(n1846), .B(n1845), .Z(n5584) );
  XOR U6770 ( .A(n5585), .B(n5584), .Z(n5587) );
  NANDN U6771 ( .A(n1848), .B(n1847), .Z(n1852) );
  NANDN U6772 ( .A(n1850), .B(n1849), .Z(n1851) );
  AND U6773 ( .A(n1852), .B(n1851), .Z(n5586) );
  XNOR U6774 ( .A(n5587), .B(n5586), .Z(n6431) );
  XNOR U6775 ( .A(n6432), .B(n6431), .Z(n6434) );
  XOR U6776 ( .A(n6433), .B(n6434), .Z(n6018) );
  XOR U6777 ( .A(n6019), .B(n6018), .Z(n6937) );
  NANDN U6778 ( .A(n1854), .B(n1853), .Z(n1858) );
  NAND U6779 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U6780 ( .A(n1858), .B(n1857), .Z(n6047) );
  XNOR U6781 ( .A(n6047), .B(n6046), .Z(n6049) );
  NANDN U6782 ( .A(n1864), .B(n1863), .Z(n1868) );
  NANDN U6783 ( .A(n1866), .B(n1865), .Z(n1867) );
  NAND U6784 ( .A(n1868), .B(n1867), .Z(n6056) );
  NANDN U6785 ( .A(n1870), .B(n1869), .Z(n1874) );
  NANDN U6786 ( .A(n1872), .B(n1871), .Z(n1873) );
  NAND U6787 ( .A(n1874), .B(n1873), .Z(n6057) );
  XOR U6788 ( .A(n6056), .B(n6057), .Z(n6058) );
  NANDN U6789 ( .A(n1876), .B(n1875), .Z(n1880) );
  NANDN U6790 ( .A(n1878), .B(n1877), .Z(n1879) );
  NAND U6791 ( .A(n1880), .B(n1879), .Z(n6060) );
  XNOR U6792 ( .A(n6060), .B(n6062), .Z(n6059) );
  XNOR U6793 ( .A(n6058), .B(n6059), .Z(n6048) );
  XOR U6794 ( .A(n6049), .B(n6048), .Z(n6735) );
  NAND U6795 ( .A(n1888), .B(n1887), .Z(n1893) );
  IV U6796 ( .A(n1889), .Z(n1891) );
  NANDN U6797 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U6798 ( .A(n1893), .B(n1892), .Z(n6064) );
  XNOR U6799 ( .A(n6063), .B(n6064), .Z(n6065) );
  XNOR U6800 ( .A(n6065), .B(n6066), .Z(n6733) );
  XNOR U6801 ( .A(n6083), .B(n6084), .Z(n6085) );
  XOR U6802 ( .A(n6085), .B(n6086), .Z(n6734) );
  XOR U6803 ( .A(n6733), .B(n6734), .Z(n6736) );
  XOR U6804 ( .A(n6735), .B(n6736), .Z(n5972) );
  NANDN U6805 ( .A(n1919), .B(n1918), .Z(n1923) );
  NAND U6806 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U6807 ( .A(n1923), .B(n1922), .Z(n7267) );
  XOR U6808 ( .A(n7268), .B(n7267), .Z(n7270) );
  XNOR U6809 ( .A(n7269), .B(n7270), .Z(n5970) );
  NANDN U6810 ( .A(n1925), .B(n1924), .Z(n1929) );
  NANDN U6811 ( .A(n1927), .B(n1926), .Z(n1928) );
  AND U6812 ( .A(n1929), .B(n1928), .Z(n6857) );
  NANDN U6813 ( .A(n1931), .B(n1930), .Z(n1935) );
  NAND U6814 ( .A(n1933), .B(n1932), .Z(n1934) );
  NAND U6815 ( .A(n1935), .B(n1934), .Z(n6858) );
  XNOR U6816 ( .A(n6857), .B(n6858), .Z(n6860) );
  NANDN U6817 ( .A(n1937), .B(n1936), .Z(n1941) );
  NANDN U6818 ( .A(n1939), .B(n1938), .Z(n1940) );
  AND U6819 ( .A(n1941), .B(n1940), .Z(n6859) );
  XOR U6820 ( .A(n6860), .B(n6859), .Z(n7308) );
  NANDN U6821 ( .A(n1943), .B(n1942), .Z(n1947) );
  NANDN U6822 ( .A(n1945), .B(n1944), .Z(n1946) );
  AND U6823 ( .A(n1947), .B(n1946), .Z(n6917) );
  NANDN U6824 ( .A(n1949), .B(n1948), .Z(n1953) );
  NANDN U6825 ( .A(n1951), .B(n1950), .Z(n1952) );
  NAND U6826 ( .A(n1953), .B(n1952), .Z(n6918) );
  XNOR U6827 ( .A(n6917), .B(n6918), .Z(n6920) );
  NANDN U6828 ( .A(n1955), .B(n1954), .Z(n1959) );
  NANDN U6829 ( .A(n1957), .B(n1956), .Z(n1958) );
  AND U6830 ( .A(n1959), .B(n1958), .Z(n6919) );
  XOR U6831 ( .A(n6920), .B(n6919), .Z(n7306) );
  NANDN U6832 ( .A(n1961), .B(n1960), .Z(n1965) );
  NANDN U6833 ( .A(n1963), .B(n1962), .Z(n1964) );
  NAND U6834 ( .A(n1965), .B(n1964), .Z(n7305) );
  XNOR U6835 ( .A(n7306), .B(n7305), .Z(n7307) );
  XOR U6836 ( .A(n7308), .B(n7307), .Z(n5971) );
  XOR U6837 ( .A(n5970), .B(n5971), .Z(n5973) );
  XOR U6838 ( .A(n5972), .B(n5973), .Z(n6936) );
  NANDN U6839 ( .A(n1967), .B(n1966), .Z(n1971) );
  NAND U6840 ( .A(n1969), .B(n1968), .Z(n1970) );
  AND U6841 ( .A(n1971), .B(n1970), .Z(n6838) );
  NANDN U6842 ( .A(n1973), .B(n1972), .Z(n1977) );
  NANDN U6843 ( .A(n1975), .B(n1974), .Z(n1976) );
  AND U6844 ( .A(n1977), .B(n1976), .Z(n5988) );
  XNOR U6845 ( .A(n5988), .B(n5989), .Z(n5991) );
  XOR U6846 ( .A(n5991), .B(n5990), .Z(n6836) );
  XNOR U6847 ( .A(n6836), .B(n6835), .Z(n6837) );
  XNOR U6848 ( .A(n6838), .B(n6837), .Z(n6866) );
  NANDN U6849 ( .A(n1995), .B(n1994), .Z(n1999) );
  NANDN U6850 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U6851 ( .A(n1999), .B(n1998), .Z(n5999) );
  XOR U6852 ( .A(n5999), .B(n5998), .Z(n6001) );
  NANDN U6853 ( .A(n2005), .B(n2004), .Z(n2009) );
  NANDN U6854 ( .A(n2007), .B(n2006), .Z(n2008) );
  AND U6855 ( .A(n2009), .B(n2008), .Z(n6000) );
  XOR U6856 ( .A(n6001), .B(n6000), .Z(n5983) );
  XNOR U6857 ( .A(n5983), .B(n5982), .Z(n5984) );
  XNOR U6858 ( .A(n5985), .B(n5984), .Z(n6864) );
  NANDN U6859 ( .A(n2015), .B(n2014), .Z(n2019) );
  NAND U6860 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U6861 ( .A(n2019), .B(n2018), .Z(n6157) );
  NANDN U6862 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U6863 ( .A(n2023), .B(n2022), .Z(n2024) );
  NAND U6864 ( .A(n2025), .B(n2024), .Z(n6158) );
  XNOR U6865 ( .A(n6157), .B(n6158), .Z(n6159) );
  NANDN U6866 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U6867 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U6868 ( .A(n2031), .B(n2030), .Z(n6160) );
  XOR U6869 ( .A(n6159), .B(n6160), .Z(n6411) );
  NANDN U6870 ( .A(n2033), .B(n2032), .Z(n2037) );
  NAND U6871 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U6872 ( .A(n2037), .B(n2036), .Z(n6253) );
  NANDN U6873 ( .A(n2039), .B(n2038), .Z(n2043) );
  NANDN U6874 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U6875 ( .A(n2043), .B(n2042), .Z(n6254) );
  XNOR U6876 ( .A(n6253), .B(n6254), .Z(n6255) );
  NANDN U6877 ( .A(n2045), .B(n2044), .Z(n2049) );
  NANDN U6878 ( .A(n2047), .B(n2046), .Z(n2048) );
  NAND U6879 ( .A(n2049), .B(n2048), .Z(n6256) );
  XOR U6880 ( .A(n6255), .B(n6256), .Z(n6409) );
  XOR U6881 ( .A(n6409), .B(n6410), .Z(n6412) );
  XOR U6882 ( .A(n6411), .B(n6412), .Z(n6863) );
  XOR U6883 ( .A(n6864), .B(n6863), .Z(n6865) );
  XNOR U6884 ( .A(n6866), .B(n6865), .Z(n6935) );
  XOR U6885 ( .A(n6936), .B(n6935), .Z(n6938) );
  XNOR U6886 ( .A(n6937), .B(n6938), .Z(n6877) );
  XNOR U6887 ( .A(n6878), .B(n6877), .Z(n6880) );
  NANDN U6888 ( .A(n2055), .B(n2054), .Z(n2059) );
  NAND U6889 ( .A(n2057), .B(n2056), .Z(n2058) );
  AND U6890 ( .A(n2059), .B(n2058), .Z(n6602) );
  NANDN U6891 ( .A(n2061), .B(n2060), .Z(n2065) );
  NANDN U6892 ( .A(n2063), .B(n2062), .Z(n2064) );
  AND U6893 ( .A(n2065), .B(n2064), .Z(n6600) );
  NANDN U6894 ( .A(n2067), .B(n2066), .Z(n2071) );
  NAND U6895 ( .A(n2069), .B(n2068), .Z(n2070) );
  AND U6896 ( .A(n2071), .B(n2070), .Z(n6844) );
  XNOR U6897 ( .A(n6842), .B(n6841), .Z(n6843) );
  XNOR U6898 ( .A(n6844), .B(n6843), .Z(n6539) );
  NANDN U6899 ( .A(n2081), .B(n2080), .Z(n2085) );
  NANDN U6900 ( .A(n2083), .B(n2082), .Z(n2084) );
  AND U6901 ( .A(n2085), .B(n2084), .Z(n6314) );
  NANDN U6902 ( .A(n2087), .B(n2086), .Z(n2091) );
  NANDN U6903 ( .A(n2089), .B(n2088), .Z(n2090) );
  AND U6904 ( .A(n2091), .B(n2090), .Z(n5665) );
  NANDN U6905 ( .A(n2093), .B(n2092), .Z(n2097) );
  NANDN U6906 ( .A(n2095), .B(n2094), .Z(n2096) );
  NAND U6907 ( .A(n2097), .B(n2096), .Z(n5666) );
  XNOR U6908 ( .A(n5665), .B(n5666), .Z(n5668) );
  NANDN U6909 ( .A(n2099), .B(n2098), .Z(n2103) );
  NAND U6910 ( .A(n2101), .B(n2100), .Z(n2102) );
  AND U6911 ( .A(n2103), .B(n2102), .Z(n5667) );
  XOR U6912 ( .A(n5668), .B(n5667), .Z(n6312) );
  XNOR U6913 ( .A(n6312), .B(n6311), .Z(n6313) );
  XOR U6914 ( .A(n6314), .B(n6313), .Z(n6540) );
  XNOR U6915 ( .A(n6539), .B(n6540), .Z(n6541) );
  NANDN U6916 ( .A(n2109), .B(n2108), .Z(n2113) );
  NANDN U6917 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U6918 ( .A(n2113), .B(n2112), .Z(n5618) );
  NANDN U6919 ( .A(n2115), .B(n2114), .Z(n2119) );
  NANDN U6920 ( .A(n2117), .B(n2116), .Z(n2118) );
  AND U6921 ( .A(n2119), .B(n2118), .Z(n5617) );
  XOR U6922 ( .A(n5618), .B(n5617), .Z(n5620) );
  NANDN U6923 ( .A(n2121), .B(n2120), .Z(n2125) );
  NANDN U6924 ( .A(n2123), .B(n2122), .Z(n2124) );
  AND U6925 ( .A(n2125), .B(n2124), .Z(n5619) );
  XOR U6926 ( .A(n5620), .B(n5619), .Z(n6274) );
  NANDN U6927 ( .A(n2127), .B(n2126), .Z(n2131) );
  NANDN U6928 ( .A(n2129), .B(n2128), .Z(n2130) );
  AND U6929 ( .A(n2131), .B(n2130), .Z(n5995) );
  NANDN U6930 ( .A(n2133), .B(n2132), .Z(n2137) );
  NANDN U6931 ( .A(n2135), .B(n2134), .Z(n2136) );
  AND U6932 ( .A(n2137), .B(n2136), .Z(n5994) );
  XOR U6933 ( .A(n5995), .B(n5994), .Z(n5997) );
  NANDN U6934 ( .A(n2139), .B(n2138), .Z(n2143) );
  NANDN U6935 ( .A(n2141), .B(n2140), .Z(n2142) );
  AND U6936 ( .A(n2143), .B(n2142), .Z(n5996) );
  XOR U6937 ( .A(n5997), .B(n5996), .Z(n6272) );
  NANDN U6938 ( .A(n2145), .B(n2144), .Z(n2149) );
  NANDN U6939 ( .A(n2147), .B(n2146), .Z(n2148) );
  AND U6940 ( .A(n2149), .B(n2148), .Z(n5577) );
  NANDN U6941 ( .A(n2151), .B(n2150), .Z(n2155) );
  NANDN U6942 ( .A(n2153), .B(n2152), .Z(n2154) );
  AND U6943 ( .A(n2155), .B(n2154), .Z(n5576) );
  XOR U6944 ( .A(n5577), .B(n5576), .Z(n5579) );
  NANDN U6945 ( .A(n2157), .B(n2156), .Z(n2161) );
  NANDN U6946 ( .A(n2159), .B(n2158), .Z(n2160) );
  AND U6947 ( .A(n2161), .B(n2160), .Z(n5578) );
  XNOR U6948 ( .A(n5579), .B(n5578), .Z(n6271) );
  XNOR U6949 ( .A(n6272), .B(n6271), .Z(n6273) );
  XOR U6950 ( .A(n6274), .B(n6273), .Z(n6542) );
  XNOR U6951 ( .A(n6541), .B(n6542), .Z(n6599) );
  XOR U6952 ( .A(n6602), .B(n6601), .Z(n6879) );
  XOR U6953 ( .A(n6880), .B(n6879), .Z(n7438) );
  NANDN U6954 ( .A(n2163), .B(n2162), .Z(n2167) );
  NANDN U6955 ( .A(n2165), .B(n2164), .Z(n2166) );
  AND U6956 ( .A(n2167), .B(n2166), .Z(n6549) );
  XNOR U6957 ( .A(n5719), .B(n5720), .Z(n5722) );
  NANDN U6958 ( .A(n2177), .B(n2176), .Z(n2181) );
  NANDN U6959 ( .A(n2179), .B(n2178), .Z(n2180) );
  AND U6960 ( .A(n2181), .B(n2180), .Z(n5721) );
  XOR U6961 ( .A(n5722), .B(n5721), .Z(n6680) );
  NANDN U6962 ( .A(n2183), .B(n2182), .Z(n2187) );
  NANDN U6963 ( .A(n2185), .B(n2184), .Z(n2186) );
  AND U6964 ( .A(n2187), .B(n2186), .Z(n5689) );
  NANDN U6965 ( .A(n2189), .B(n2188), .Z(n2193) );
  NANDN U6966 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U6967 ( .A(n2193), .B(n2192), .Z(n5690) );
  XNOR U6968 ( .A(n5689), .B(n5690), .Z(n5692) );
  NANDN U6969 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U6970 ( .A(n2197), .B(n2196), .Z(n2198) );
  AND U6971 ( .A(n2199), .B(n2198), .Z(n5691) );
  XOR U6972 ( .A(n5692), .B(n5691), .Z(n6678) );
  XNOR U6973 ( .A(n6678), .B(n6677), .Z(n6679) );
  XOR U6974 ( .A(n6680), .B(n6679), .Z(n6550) );
  XNOR U6975 ( .A(n6549), .B(n6550), .Z(n6551) );
  NANDN U6976 ( .A(n2205), .B(n2204), .Z(n2209) );
  NANDN U6977 ( .A(n2207), .B(n2206), .Z(n2208) );
  AND U6978 ( .A(n2209), .B(n2208), .Z(n5769) );
  NANDN U6979 ( .A(n2211), .B(n2210), .Z(n2215) );
  NANDN U6980 ( .A(n2213), .B(n2212), .Z(n2214) );
  AND U6981 ( .A(n2215), .B(n2214), .Z(n5768) );
  XOR U6982 ( .A(n5769), .B(n5768), .Z(n5771) );
  NANDN U6983 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U6984 ( .A(n2219), .B(n2218), .Z(n2220) );
  AND U6985 ( .A(n2221), .B(n2220), .Z(n5770) );
  XOR U6986 ( .A(n5771), .B(n5770), .Z(n6674) );
  NANDN U6987 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U6988 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U6989 ( .A(n2227), .B(n2226), .Z(n5755) );
  NANDN U6990 ( .A(n2229), .B(n2228), .Z(n2233) );
  NANDN U6991 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U6992 ( .A(n2233), .B(n2232), .Z(n5754) );
  XOR U6993 ( .A(n5755), .B(n5754), .Z(n5757) );
  XOR U6994 ( .A(n5757), .B(n5756), .Z(n6672) );
  XNOR U6995 ( .A(n6672), .B(n6671), .Z(n6673) );
  XOR U6996 ( .A(n6674), .B(n6673), .Z(n6552) );
  XNOR U6997 ( .A(n6551), .B(n6552), .Z(n7076) );
  NANDN U6998 ( .A(n2243), .B(n2242), .Z(n2247) );
  NANDN U6999 ( .A(n2245), .B(n2244), .Z(n2246) );
  AND U7000 ( .A(n2247), .B(n2246), .Z(n5765) );
  NANDN U7001 ( .A(n2249), .B(n2248), .Z(n2253) );
  NAND U7002 ( .A(n2251), .B(n2250), .Z(n2252) );
  AND U7003 ( .A(n2253), .B(n2252), .Z(n5764) );
  XOR U7004 ( .A(n5765), .B(n5764), .Z(n5767) );
  XOR U7005 ( .A(n5767), .B(n5766), .Z(n7244) );
  NANDN U7006 ( .A(n2259), .B(n2258), .Z(n2263) );
  NAND U7007 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U7008 ( .A(n2263), .B(n2262), .Z(n7242) );
  XNOR U7009 ( .A(n7242), .B(n7241), .Z(n7243) );
  XOR U7010 ( .A(n7244), .B(n7243), .Z(n6557) );
  NANDN U7011 ( .A(n2269), .B(n2268), .Z(n2273) );
  NANDN U7012 ( .A(n2271), .B(n2270), .Z(n2272) );
  AND U7013 ( .A(n2273), .B(n2272), .Z(n6556) );
  NANDN U7014 ( .A(n2275), .B(n2274), .Z(n2279) );
  NANDN U7015 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U7016 ( .A(n2279), .B(n2278), .Z(n6187) );
  NANDN U7017 ( .A(n2281), .B(n2280), .Z(n2285) );
  NANDN U7018 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U7019 ( .A(n2285), .B(n2284), .Z(n6188) );
  XNOR U7020 ( .A(n6187), .B(n6188), .Z(n6190) );
  NANDN U7021 ( .A(n2287), .B(n2286), .Z(n2291) );
  NANDN U7022 ( .A(n2289), .B(n2288), .Z(n2290) );
  AND U7023 ( .A(n2291), .B(n2290), .Z(n6189) );
  XOR U7024 ( .A(n6190), .B(n6189), .Z(n6320) );
  NANDN U7025 ( .A(n2293), .B(n2292), .Z(n2297) );
  NAND U7026 ( .A(n2295), .B(n2294), .Z(n2296) );
  AND U7027 ( .A(n2297), .B(n2296), .Z(n6318) );
  NANDN U7028 ( .A(n2299), .B(n2298), .Z(n2303) );
  NAND U7029 ( .A(n2301), .B(n2300), .Z(n2302) );
  NAND U7030 ( .A(n2303), .B(n2302), .Z(n6317) );
  XNOR U7031 ( .A(n6318), .B(n6317), .Z(n6319) );
  XOR U7032 ( .A(n6320), .B(n6319), .Z(n6555) );
  XOR U7033 ( .A(n6556), .B(n6555), .Z(n6558) );
  XOR U7034 ( .A(n6557), .B(n6558), .Z(n7073) );
  NANDN U7035 ( .A(n2305), .B(n2304), .Z(n2309) );
  NANDN U7036 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U7037 ( .A(n2309), .B(n2308), .Z(n7074) );
  XOR U7038 ( .A(n7073), .B(n7074), .Z(n7075) );
  XOR U7039 ( .A(n7076), .B(n7075), .Z(n6268) );
  NANDN U7040 ( .A(n2311), .B(n2310), .Z(n2315) );
  OR U7041 ( .A(n2313), .B(n2312), .Z(n2314) );
  AND U7042 ( .A(n2315), .B(n2314), .Z(n6266) );
  NANDN U7043 ( .A(n2317), .B(n2316), .Z(n2321) );
  NAND U7044 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U7045 ( .A(n2321), .B(n2320), .Z(n7001) );
  NANDN U7046 ( .A(n2323), .B(n2322), .Z(n2327) );
  NANDN U7047 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U7048 ( .A(n2327), .B(n2326), .Z(n5318) );
  NANDN U7049 ( .A(n2329), .B(n2328), .Z(n2333) );
  NANDN U7050 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U7051 ( .A(n2333), .B(n2332), .Z(n5319) );
  XNOR U7052 ( .A(n5318), .B(n5319), .Z(n5321) );
  NANDN U7053 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U7054 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U7055 ( .A(n2339), .B(n2338), .Z(n5794) );
  NANDN U7056 ( .A(n2341), .B(n2340), .Z(n2345) );
  NANDN U7057 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U7058 ( .A(n2345), .B(n2344), .Z(n5795) );
  XNOR U7059 ( .A(n5794), .B(n5795), .Z(n5796) );
  NANDN U7060 ( .A(n2347), .B(n2346), .Z(n2351) );
  NANDN U7061 ( .A(n2349), .B(n2348), .Z(n2350) );
  NAND U7062 ( .A(n2351), .B(n2350), .Z(n5797) );
  XOR U7063 ( .A(n5796), .B(n5797), .Z(n6339) );
  NANDN U7064 ( .A(n2357), .B(n2356), .Z(n2361) );
  NANDN U7065 ( .A(n2359), .B(n2358), .Z(n2360) );
  AND U7066 ( .A(n2361), .B(n2360), .Z(n5804) );
  NANDN U7067 ( .A(n2363), .B(n2362), .Z(n2367) );
  NANDN U7068 ( .A(n2365), .B(n2364), .Z(n2366) );
  NAND U7069 ( .A(n2367), .B(n2366), .Z(n5805) );
  XNOR U7070 ( .A(n5804), .B(n5805), .Z(n5807) );
  NANDN U7071 ( .A(n2369), .B(n2368), .Z(n2373) );
  NANDN U7072 ( .A(n2371), .B(n2370), .Z(n2372) );
  AND U7073 ( .A(n2373), .B(n2372), .Z(n5806) );
  XNOR U7074 ( .A(n5807), .B(n5806), .Z(n6338) );
  XOR U7075 ( .A(n6337), .B(n6338), .Z(n6340) );
  XOR U7076 ( .A(n6339), .B(n6340), .Z(n5320) );
  XOR U7077 ( .A(n5321), .B(n5320), .Z(n7000) );
  NANDN U7078 ( .A(n2375), .B(n2374), .Z(n2379) );
  NAND U7079 ( .A(n2377), .B(n2376), .Z(n2378) );
  NAND U7080 ( .A(n2379), .B(n2378), .Z(n6999) );
  XOR U7081 ( .A(n7000), .B(n6999), .Z(n7002) );
  XOR U7082 ( .A(n7001), .B(n7002), .Z(n6265) );
  XOR U7083 ( .A(n6266), .B(n6265), .Z(n6267) );
  XOR U7084 ( .A(n7438), .B(n7437), .Z(n7440) );
  XOR U7085 ( .A(n7439), .B(n7440), .Z(n7444) );
  NANDN U7086 ( .A(n2381), .B(n2380), .Z(n2385) );
  NAND U7087 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U7088 ( .A(n2385), .B(n2384), .Z(n6827) );
  NANDN U7089 ( .A(n2387), .B(n2386), .Z(n2391) );
  NANDN U7090 ( .A(n2389), .B(n2388), .Z(n2390) );
  AND U7091 ( .A(n2391), .B(n2390), .Z(n6136) );
  NANDN U7092 ( .A(n2393), .B(n2392), .Z(n2397) );
  NANDN U7093 ( .A(n2395), .B(n2394), .Z(n2396) );
  AND U7094 ( .A(n2397), .B(n2396), .Z(n6455) );
  NANDN U7095 ( .A(n2399), .B(n2398), .Z(n2403) );
  NANDN U7096 ( .A(n2401), .B(n2400), .Z(n2402) );
  NAND U7097 ( .A(n2403), .B(n2402), .Z(n6456) );
  XNOR U7098 ( .A(n6455), .B(n6456), .Z(n6457) );
  NANDN U7099 ( .A(n2405), .B(n2404), .Z(n2409) );
  NANDN U7100 ( .A(n2407), .B(n2406), .Z(n2408) );
  NAND U7101 ( .A(n2409), .B(n2408), .Z(n6458) );
  XOR U7102 ( .A(n6457), .B(n6458), .Z(n7377) );
  NANDN U7103 ( .A(n2411), .B(n2410), .Z(n2415) );
  NANDN U7104 ( .A(n2413), .B(n2412), .Z(n2414) );
  AND U7105 ( .A(n2415), .B(n2414), .Z(n6914) );
  XOR U7106 ( .A(n6914), .B(n6913), .Z(n6916) );
  NANDN U7107 ( .A(n2421), .B(n2420), .Z(n2425) );
  NANDN U7108 ( .A(n2423), .B(n2422), .Z(n2424) );
  AND U7109 ( .A(n2425), .B(n2424), .Z(n6915) );
  XOR U7110 ( .A(n6916), .B(n6915), .Z(n7376) );
  NANDN U7111 ( .A(n2427), .B(n2426), .Z(n2431) );
  NANDN U7112 ( .A(n2429), .B(n2428), .Z(n2430) );
  AND U7113 ( .A(n2431), .B(n2430), .Z(n6461) );
  NANDN U7114 ( .A(n2433), .B(n2432), .Z(n2437) );
  NANDN U7115 ( .A(n2435), .B(n2434), .Z(n2436) );
  NAND U7116 ( .A(n2437), .B(n2436), .Z(n6462) );
  XNOR U7117 ( .A(n6461), .B(n6462), .Z(n6464) );
  NANDN U7118 ( .A(n2439), .B(n2438), .Z(n2443) );
  NANDN U7119 ( .A(n2441), .B(n2440), .Z(n2442) );
  AND U7120 ( .A(n2443), .B(n2442), .Z(n6463) );
  XNOR U7121 ( .A(n6464), .B(n6463), .Z(n7375) );
  XNOR U7122 ( .A(n7376), .B(n7375), .Z(n7378) );
  XOR U7123 ( .A(n7377), .B(n7378), .Z(n6133) );
  NANDN U7124 ( .A(n2445), .B(n2444), .Z(n2449) );
  NANDN U7125 ( .A(n2447), .B(n2446), .Z(n2448) );
  AND U7126 ( .A(n2449), .B(n2448), .Z(n6478) );
  NANDN U7127 ( .A(n2451), .B(n2450), .Z(n2455) );
  NANDN U7128 ( .A(n2453), .B(n2452), .Z(n2454) );
  AND U7129 ( .A(n2455), .B(n2454), .Z(n6477) );
  XOR U7130 ( .A(n6478), .B(n6477), .Z(n6480) );
  NANDN U7131 ( .A(n2457), .B(n2456), .Z(n2461) );
  NANDN U7132 ( .A(n2459), .B(n2458), .Z(n2460) );
  AND U7133 ( .A(n2461), .B(n2460), .Z(n6479) );
  XOR U7134 ( .A(n6480), .B(n6479), .Z(n5389) );
  NANDN U7135 ( .A(n2463), .B(n2462), .Z(n2467) );
  NANDN U7136 ( .A(n2465), .B(n2464), .Z(n2466) );
  AND U7137 ( .A(n2467), .B(n2466), .Z(n6910) );
  NANDN U7138 ( .A(n2469), .B(n2468), .Z(n2473) );
  NANDN U7139 ( .A(n2471), .B(n2470), .Z(n2472) );
  AND U7140 ( .A(n2473), .B(n2472), .Z(n6909) );
  XOR U7141 ( .A(n6910), .B(n6909), .Z(n6912) );
  NANDN U7142 ( .A(n2475), .B(n2474), .Z(n2479) );
  NANDN U7143 ( .A(n2477), .B(n2476), .Z(n2478) );
  AND U7144 ( .A(n2479), .B(n2478), .Z(n6911) );
  XOR U7145 ( .A(n6912), .B(n6911), .Z(n5387) );
  XNOR U7146 ( .A(n5387), .B(n5386), .Z(n5388) );
  XOR U7147 ( .A(n5389), .B(n5388), .Z(n6134) );
  XNOR U7148 ( .A(n6133), .B(n6134), .Z(n6135) );
  XOR U7149 ( .A(n6136), .B(n6135), .Z(n6826) );
  NANDN U7150 ( .A(n2485), .B(n2484), .Z(n2489) );
  OR U7151 ( .A(n2487), .B(n2486), .Z(n2488) );
  AND U7152 ( .A(n2489), .B(n2488), .Z(n6825) );
  XOR U7153 ( .A(n6826), .B(n6825), .Z(n6828) );
  XOR U7154 ( .A(n6827), .B(n6828), .Z(n5301) );
  NANDN U7155 ( .A(n2491), .B(n2490), .Z(n2495) );
  NANDN U7156 ( .A(n2493), .B(n2492), .Z(n2494) );
  AND U7157 ( .A(n2495), .B(n2494), .Z(n5299) );
  NANDN U7158 ( .A(n2497), .B(n2496), .Z(n2501) );
  NAND U7159 ( .A(n2499), .B(n2498), .Z(n2500) );
  AND U7160 ( .A(n2501), .B(n2500), .Z(n6126) );
  NANDN U7161 ( .A(n2507), .B(n2506), .Z(n2511) );
  NANDN U7162 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U7163 ( .A(n2511), .B(n2510), .Z(n6451) );
  XOR U7164 ( .A(n6452), .B(n6451), .Z(n6454) );
  XOR U7165 ( .A(n6454), .B(n6453), .Z(n6124) );
  XNOR U7166 ( .A(n6124), .B(n6123), .Z(n6125) );
  XNOR U7167 ( .A(n6126), .B(n6125), .Z(n7187) );
  NANDN U7168 ( .A(n2521), .B(n2520), .Z(n2525) );
  NANDN U7169 ( .A(n2523), .B(n2522), .Z(n2524) );
  AND U7170 ( .A(n2525), .B(n2524), .Z(n6353) );
  NANDN U7171 ( .A(n2527), .B(n2526), .Z(n2531) );
  NAND U7172 ( .A(n2529), .B(n2528), .Z(n2530) );
  NAND U7173 ( .A(n2531), .B(n2530), .Z(n6354) );
  NANDN U7174 ( .A(n2533), .B(n2532), .Z(n2537) );
  NANDN U7175 ( .A(n2535), .B(n2534), .Z(n2536) );
  AND U7176 ( .A(n2537), .B(n2536), .Z(n6355) );
  XOR U7177 ( .A(n6356), .B(n6355), .Z(n6490) );
  XNOR U7178 ( .A(n6403), .B(n6404), .Z(n6406) );
  NANDN U7179 ( .A(n2547), .B(n2546), .Z(n2551) );
  NANDN U7180 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U7181 ( .A(n2551), .B(n2550), .Z(n6405) );
  XOR U7182 ( .A(n6406), .B(n6405), .Z(n6488) );
  NANDN U7183 ( .A(n2553), .B(n2552), .Z(n2557) );
  NANDN U7184 ( .A(n2555), .B(n2554), .Z(n2556) );
  NAND U7185 ( .A(n2557), .B(n2556), .Z(n6487) );
  XNOR U7186 ( .A(n6488), .B(n6487), .Z(n6489) );
  XOR U7187 ( .A(n6490), .B(n6489), .Z(n7188) );
  XNOR U7188 ( .A(n7187), .B(n7188), .Z(n7190) );
  NANDN U7189 ( .A(n2559), .B(n2558), .Z(n2563) );
  NANDN U7190 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U7191 ( .A(n2563), .B(n2562), .Z(n5961) );
  NANDN U7192 ( .A(n2565), .B(n2564), .Z(n2569) );
  NANDN U7193 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U7194 ( .A(n2569), .B(n2568), .Z(n5960) );
  XOR U7195 ( .A(n5961), .B(n5960), .Z(n5963) );
  NANDN U7196 ( .A(n2571), .B(n2570), .Z(n2575) );
  NANDN U7197 ( .A(n2573), .B(n2572), .Z(n2574) );
  AND U7198 ( .A(n2575), .B(n2574), .Z(n5962) );
  XOR U7199 ( .A(n5963), .B(n5962), .Z(n5515) );
  NANDN U7200 ( .A(n2577), .B(n2576), .Z(n2581) );
  NANDN U7201 ( .A(n2579), .B(n2578), .Z(n2580) );
  AND U7202 ( .A(n2581), .B(n2580), .Z(n5934) );
  NANDN U7203 ( .A(n2583), .B(n2582), .Z(n2587) );
  NANDN U7204 ( .A(n2585), .B(n2584), .Z(n2586) );
  NAND U7205 ( .A(n2587), .B(n2586), .Z(n5935) );
  XNOR U7206 ( .A(n5934), .B(n5935), .Z(n5937) );
  NANDN U7207 ( .A(n2589), .B(n2588), .Z(n2593) );
  NANDN U7208 ( .A(n2591), .B(n2590), .Z(n2592) );
  AND U7209 ( .A(n2593), .B(n2592), .Z(n5936) );
  XOR U7210 ( .A(n5937), .B(n5936), .Z(n5513) );
  XNOR U7211 ( .A(n5513), .B(n5512), .Z(n5514) );
  XNOR U7212 ( .A(n5515), .B(n5514), .Z(n7189) );
  XOR U7213 ( .A(n7190), .B(n7189), .Z(n6885) );
  NANDN U7214 ( .A(n2599), .B(n2598), .Z(n2603) );
  NAND U7215 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U7216 ( .A(n2603), .B(n2602), .Z(n7150) );
  NAND U7217 ( .A(n2605), .B(n2604), .Z(n2609) );
  NAND U7218 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U7219 ( .A(n2609), .B(n2608), .Z(n7148) );
  NANDN U7220 ( .A(n2611), .B(n2610), .Z(n2615) );
  NAND U7221 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U7222 ( .A(n2615), .B(n2614), .Z(n7147) );
  XNOR U7223 ( .A(n7148), .B(n7147), .Z(n7149) );
  XNOR U7224 ( .A(n7150), .B(n7149), .Z(n7412) );
  NAND U7225 ( .A(n2617), .B(n2616), .Z(n2621) );
  NAND U7226 ( .A(n2619), .B(n2618), .Z(n2620) );
  AND U7227 ( .A(n2621), .B(n2620), .Z(n7126) );
  NAND U7228 ( .A(n2623), .B(n2622), .Z(n2627) );
  NAND U7229 ( .A(n2625), .B(n2624), .Z(n2626) );
  AND U7230 ( .A(n2627), .B(n2626), .Z(n7124) );
  NAND U7231 ( .A(n2629), .B(n2628), .Z(n2633) );
  NAND U7232 ( .A(n2631), .B(n2630), .Z(n2632) );
  NAND U7233 ( .A(n2633), .B(n2632), .Z(n7123) );
  XNOR U7234 ( .A(n7124), .B(n7123), .Z(n7125) );
  XNOR U7235 ( .A(n7126), .B(n7125), .Z(n7409) );
  NANDN U7236 ( .A(n2635), .B(n2634), .Z(n2639) );
  NANDN U7237 ( .A(n2637), .B(n2636), .Z(n2638) );
  AND U7238 ( .A(n2639), .B(n2638), .Z(n7155) );
  NANDN U7239 ( .A(n2641), .B(n2640), .Z(n2645) );
  NAND U7240 ( .A(n2643), .B(n2642), .Z(n2644) );
  AND U7241 ( .A(n2645), .B(n2644), .Z(n7154) );
  NAND U7242 ( .A(n2647), .B(n2646), .Z(n2651) );
  NAND U7243 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U7244 ( .A(n2651), .B(n2650), .Z(n7153) );
  XOR U7245 ( .A(n7154), .B(n7153), .Z(n7156) );
  XOR U7246 ( .A(n7155), .B(n7156), .Z(n7410) );
  XNOR U7247 ( .A(n7409), .B(n7410), .Z(n7411) );
  XOR U7248 ( .A(n7412), .B(n7411), .Z(n6884) );
  NANDN U7249 ( .A(n2653), .B(n2652), .Z(n2657) );
  NAND U7250 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U7251 ( .A(n2657), .B(n2656), .Z(n6883) );
  XOR U7252 ( .A(n6884), .B(n6883), .Z(n6886) );
  XNOR U7253 ( .A(n6885), .B(n6886), .Z(n5298) );
  XNOR U7254 ( .A(n5299), .B(n5298), .Z(n5300) );
  XOR U7255 ( .A(n5301), .B(n5300), .Z(n5294) );
  NANDN U7256 ( .A(n2659), .B(n2658), .Z(n2663) );
  NANDN U7257 ( .A(n2661), .B(n2660), .Z(n2662) );
  AND U7258 ( .A(n2663), .B(n2662), .Z(n5818) );
  NANDN U7259 ( .A(n2665), .B(n2664), .Z(n2669) );
  NAND U7260 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U7261 ( .A(n2669), .B(n2668), .Z(n5357) );
  NANDN U7262 ( .A(n2671), .B(n2670), .Z(n2675) );
  NANDN U7263 ( .A(n2673), .B(n2672), .Z(n2674) );
  AND U7264 ( .A(n2675), .B(n2674), .Z(n7285) );
  NANDN U7265 ( .A(n2677), .B(n2676), .Z(n2681) );
  NANDN U7266 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U7267 ( .A(n2681), .B(n2680), .Z(n7286) );
  XNOR U7268 ( .A(n7285), .B(n7286), .Z(n7288) );
  NANDN U7269 ( .A(n2683), .B(n2682), .Z(n2687) );
  NANDN U7270 ( .A(n2685), .B(n2684), .Z(n2686) );
  AND U7271 ( .A(n2687), .B(n2686), .Z(n7287) );
  XOR U7272 ( .A(n7288), .B(n7287), .Z(n5355) );
  NANDN U7273 ( .A(n2689), .B(n2688), .Z(n2693) );
  NAND U7274 ( .A(n2691), .B(n2690), .Z(n2692) );
  NAND U7275 ( .A(n2693), .B(n2692), .Z(n5354) );
  XNOR U7276 ( .A(n5355), .B(n5354), .Z(n5356) );
  XNOR U7277 ( .A(n5357), .B(n5356), .Z(n7017) );
  NANDN U7278 ( .A(n2695), .B(n2694), .Z(n2699) );
  NAND U7279 ( .A(n2697), .B(n2696), .Z(n2698) );
  AND U7280 ( .A(n2699), .B(n2698), .Z(n7354) );
  NANDN U7281 ( .A(n2701), .B(n2700), .Z(n2705) );
  NANDN U7282 ( .A(n2703), .B(n2702), .Z(n2704) );
  AND U7283 ( .A(n2705), .B(n2704), .Z(n7302) );
  NANDN U7284 ( .A(n2707), .B(n2706), .Z(n2711) );
  NANDN U7285 ( .A(n2709), .B(n2708), .Z(n2710) );
  AND U7286 ( .A(n2711), .B(n2710), .Z(n7301) );
  XOR U7287 ( .A(n7302), .B(n7301), .Z(n7304) );
  XOR U7288 ( .A(n7304), .B(n7303), .Z(n7352) );
  NANDN U7289 ( .A(n2717), .B(n2716), .Z(n2721) );
  NAND U7290 ( .A(n2719), .B(n2718), .Z(n2720) );
  NAND U7291 ( .A(n2721), .B(n2720), .Z(n7351) );
  XNOR U7292 ( .A(n7352), .B(n7351), .Z(n7353) );
  XOR U7293 ( .A(n7354), .B(n7353), .Z(n7018) );
  XNOR U7294 ( .A(n7017), .B(n7018), .Z(n7020) );
  NANDN U7295 ( .A(n2727), .B(n2726), .Z(n2731) );
  NANDN U7296 ( .A(n2729), .B(n2728), .Z(n2730) );
  AND U7297 ( .A(n2731), .B(n2730), .Z(n5885) );
  NANDN U7298 ( .A(n2733), .B(n2732), .Z(n2737) );
  NANDN U7299 ( .A(n2735), .B(n2734), .Z(n2736) );
  AND U7300 ( .A(n2737), .B(n2736), .Z(n5884) );
  XOR U7301 ( .A(n5885), .B(n5884), .Z(n5887) );
  NANDN U7302 ( .A(n2739), .B(n2738), .Z(n2743) );
  NANDN U7303 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U7304 ( .A(n2743), .B(n2742), .Z(n5886) );
  XOR U7305 ( .A(n5887), .B(n5886), .Z(n5381) );
  XNOR U7306 ( .A(n5381), .B(n5380), .Z(n5382) );
  XNOR U7307 ( .A(n5383), .B(n5382), .Z(n7019) );
  XOR U7308 ( .A(n7020), .B(n7019), .Z(n5978) );
  NANDN U7309 ( .A(n2753), .B(n2752), .Z(n2757) );
  OR U7310 ( .A(n2755), .B(n2754), .Z(n2756) );
  AND U7311 ( .A(n2757), .B(n2756), .Z(n6959) );
  NANDN U7312 ( .A(n2759), .B(n2758), .Z(n2763) );
  NAND U7313 ( .A(n2761), .B(n2760), .Z(n2762) );
  AND U7314 ( .A(n2763), .B(n2762), .Z(n7232) );
  NANDN U7315 ( .A(n2765), .B(n2764), .Z(n2769) );
  NANDN U7316 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U7317 ( .A(n2769), .B(n2768), .Z(n7260) );
  NANDN U7318 ( .A(n2771), .B(n2770), .Z(n2775) );
  NANDN U7319 ( .A(n2773), .B(n2772), .Z(n2774) );
  AND U7320 ( .A(n2775), .B(n2774), .Z(n7259) );
  XOR U7321 ( .A(n7260), .B(n7259), .Z(n7262) );
  NANDN U7322 ( .A(n2777), .B(n2776), .Z(n2781) );
  NANDN U7323 ( .A(n2779), .B(n2778), .Z(n2780) );
  AND U7324 ( .A(n2781), .B(n2780), .Z(n7261) );
  XOR U7325 ( .A(n7262), .B(n7261), .Z(n7230) );
  NANDN U7326 ( .A(n2783), .B(n2782), .Z(n2787) );
  NAND U7327 ( .A(n2785), .B(n2784), .Z(n2786) );
  NAND U7328 ( .A(n2787), .B(n2786), .Z(n7229) );
  XNOR U7329 ( .A(n7230), .B(n7229), .Z(n7231) );
  XOR U7330 ( .A(n7232), .B(n7231), .Z(n6960) );
  XNOR U7331 ( .A(n6959), .B(n6960), .Z(n6961) );
  XOR U7332 ( .A(n6962), .B(n6961), .Z(n5977) );
  NANDN U7333 ( .A(n2789), .B(n2788), .Z(n2793) );
  NAND U7334 ( .A(n2791), .B(n2790), .Z(n2792) );
  NAND U7335 ( .A(n2793), .B(n2792), .Z(n7369) );
  XNOR U7336 ( .A(n7319), .B(n7320), .Z(n7321) );
  NANDN U7337 ( .A(n2803), .B(n2802), .Z(n2807) );
  NANDN U7338 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U7339 ( .A(n2807), .B(n2806), .Z(n7322) );
  XOR U7340 ( .A(n7321), .B(n7322), .Z(n7367) );
  NANDN U7341 ( .A(n2809), .B(n2808), .Z(n2813) );
  NAND U7342 ( .A(n2811), .B(n2810), .Z(n2812) );
  NAND U7343 ( .A(n2813), .B(n2812), .Z(n7368) );
  XOR U7344 ( .A(n7367), .B(n7368), .Z(n7370) );
  XOR U7345 ( .A(n7369), .B(n7370), .Z(n7058) );
  NANDN U7346 ( .A(n2819), .B(n2818), .Z(n2823) );
  NANDN U7347 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U7348 ( .A(n2823), .B(n2822), .Z(n5530) );
  NANDN U7349 ( .A(n2825), .B(n2824), .Z(n2829) );
  NANDN U7350 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U7351 ( .A(n2829), .B(n2828), .Z(n5531) );
  XNOR U7352 ( .A(n5530), .B(n5531), .Z(n5532) );
  NANDN U7353 ( .A(n2831), .B(n2830), .Z(n2835) );
  NANDN U7354 ( .A(n2833), .B(n2832), .Z(n2834) );
  NAND U7355 ( .A(n2835), .B(n2834), .Z(n5533) );
  XOR U7356 ( .A(n5532), .B(n5533), .Z(n7421) );
  NANDN U7357 ( .A(n2837), .B(n2836), .Z(n2841) );
  NAND U7358 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U7359 ( .A(n2841), .B(n2840), .Z(n7422) );
  XOR U7360 ( .A(n7421), .B(n7422), .Z(n7424) );
  XOR U7361 ( .A(n7423), .B(n7424), .Z(n7057) );
  XOR U7362 ( .A(n7058), .B(n7057), .Z(n7060) );
  NANDN U7363 ( .A(n2843), .B(n2842), .Z(n2847) );
  NAND U7364 ( .A(n2845), .B(n2844), .Z(n2846) );
  AND U7365 ( .A(n2847), .B(n2846), .Z(n5592) );
  NANDN U7366 ( .A(n2853), .B(n2852), .Z(n2857) );
  NANDN U7367 ( .A(n2855), .B(n2854), .Z(n2856) );
  AND U7368 ( .A(n2857), .B(n2856), .Z(n5902) );
  XOR U7369 ( .A(n5903), .B(n5902), .Z(n5905) );
  XOR U7370 ( .A(n5905), .B(n5904), .Z(n5590) );
  NANDN U7371 ( .A(n2863), .B(n2862), .Z(n2867) );
  NAND U7372 ( .A(n2865), .B(n2864), .Z(n2866) );
  NAND U7373 ( .A(n2867), .B(n2866), .Z(n5589) );
  XNOR U7374 ( .A(n5590), .B(n5589), .Z(n5591) );
  XNOR U7375 ( .A(n5592), .B(n5591), .Z(n7059) );
  XNOR U7376 ( .A(n7060), .B(n7059), .Z(n5976) );
  XOR U7377 ( .A(n5977), .B(n5976), .Z(n5979) );
  XOR U7378 ( .A(n5978), .B(n5979), .Z(n5817) );
  OR U7379 ( .A(n2869), .B(n2868), .Z(n2873) );
  NANDN U7380 ( .A(n2871), .B(n2870), .Z(n2872) );
  NAND U7381 ( .A(n2873), .B(n2872), .Z(n6573) );
  NANDN U7382 ( .A(n2875), .B(n2874), .Z(n2879) );
  NANDN U7383 ( .A(n2877), .B(n2876), .Z(n2878) );
  AND U7384 ( .A(n2879), .B(n2878), .Z(n5482) );
  NANDN U7385 ( .A(n2881), .B(n2880), .Z(n2885) );
  NANDN U7386 ( .A(n2883), .B(n2882), .Z(n2884) );
  NAND U7387 ( .A(n2885), .B(n2884), .Z(n5483) );
  XNOR U7388 ( .A(n5482), .B(n5483), .Z(n5485) );
  NANDN U7389 ( .A(n2887), .B(n2886), .Z(n2891) );
  NANDN U7390 ( .A(n2889), .B(n2888), .Z(n2890) );
  AND U7391 ( .A(n2891), .B(n2890), .Z(n5484) );
  XOR U7392 ( .A(n5485), .B(n5484), .Z(n6208) );
  NANDN U7393 ( .A(n2893), .B(n2892), .Z(n2897) );
  NANDN U7394 ( .A(n2895), .B(n2894), .Z(n2896) );
  AND U7395 ( .A(n2897), .B(n2896), .Z(n7312) );
  NANDN U7396 ( .A(n2899), .B(n2898), .Z(n2903) );
  NANDN U7397 ( .A(n2901), .B(n2900), .Z(n2902) );
  AND U7398 ( .A(n2903), .B(n2902), .Z(n7311) );
  XOR U7399 ( .A(n7312), .B(n7311), .Z(n7314) );
  NANDN U7400 ( .A(n2905), .B(n2904), .Z(n2909) );
  NANDN U7401 ( .A(n2907), .B(n2906), .Z(n2908) );
  AND U7402 ( .A(n2909), .B(n2908), .Z(n7313) );
  XOR U7403 ( .A(n7314), .B(n7313), .Z(n6206) );
  XNOR U7404 ( .A(n6206), .B(n6205), .Z(n6207) );
  XNOR U7405 ( .A(n6208), .B(n6207), .Z(n6572) );
  XOR U7406 ( .A(n6572), .B(n6571), .Z(n6574) );
  XOR U7407 ( .A(n6573), .B(n6574), .Z(n6129) );
  NANDN U7408 ( .A(n2919), .B(n2918), .Z(n2923) );
  OR U7409 ( .A(n2921), .B(n2920), .Z(n2922) );
  AND U7410 ( .A(n2923), .B(n2922), .Z(n6591) );
  NANDN U7411 ( .A(n2925), .B(n2924), .Z(n2929) );
  NAND U7412 ( .A(n2927), .B(n2926), .Z(n2928) );
  AND U7413 ( .A(n2929), .B(n2928), .Z(n6590) );
  NANDN U7414 ( .A(n2931), .B(n2930), .Z(n2935) );
  NANDN U7415 ( .A(n2933), .B(n2932), .Z(n2934) );
  AND U7416 ( .A(n2935), .B(n2934), .Z(n5500) );
  NANDN U7417 ( .A(n2937), .B(n2936), .Z(n2941) );
  NANDN U7418 ( .A(n2939), .B(n2938), .Z(n2940) );
  NAND U7419 ( .A(n2941), .B(n2940), .Z(n5501) );
  XNOR U7420 ( .A(n5500), .B(n5501), .Z(n5503) );
  NANDN U7421 ( .A(n2943), .B(n2942), .Z(n2947) );
  NANDN U7422 ( .A(n2945), .B(n2944), .Z(n2946) );
  AND U7423 ( .A(n2947), .B(n2946), .Z(n5502) );
  XOR U7424 ( .A(n5503), .B(n5502), .Z(n6214) );
  NANDN U7425 ( .A(n2949), .B(n2948), .Z(n2953) );
  NANDN U7426 ( .A(n2951), .B(n2950), .Z(n2952) );
  AND U7427 ( .A(n2953), .B(n2952), .Z(n7316) );
  NANDN U7428 ( .A(n2955), .B(n2954), .Z(n2959) );
  NANDN U7429 ( .A(n2957), .B(n2956), .Z(n2958) );
  AND U7430 ( .A(n2959), .B(n2958), .Z(n7315) );
  XOR U7431 ( .A(n7316), .B(n7315), .Z(n7318) );
  NANDN U7432 ( .A(n2961), .B(n2960), .Z(n2965) );
  NANDN U7433 ( .A(n2963), .B(n2962), .Z(n2964) );
  AND U7434 ( .A(n2965), .B(n2964), .Z(n7317) );
  XOR U7435 ( .A(n7318), .B(n7317), .Z(n6212) );
  NANDN U7436 ( .A(n2967), .B(n2966), .Z(n2971) );
  NAND U7437 ( .A(n2969), .B(n2968), .Z(n2970) );
  NAND U7438 ( .A(n2971), .B(n2970), .Z(n6211) );
  XNOR U7439 ( .A(n6212), .B(n6211), .Z(n6213) );
  XOR U7440 ( .A(n6214), .B(n6213), .Z(n6589) );
  XOR U7441 ( .A(n6590), .B(n6589), .Z(n6592) );
  XNOR U7442 ( .A(n6591), .B(n6592), .Z(n6130) );
  XOR U7443 ( .A(n6129), .B(n6130), .Z(n6132) );
  NANDN U7444 ( .A(n2973), .B(n2972), .Z(n2977) );
  NAND U7445 ( .A(n2975), .B(n2974), .Z(n2976) );
  AND U7446 ( .A(n2977), .B(n2976), .Z(n5488) );
  NANDN U7447 ( .A(n2979), .B(n2978), .Z(n2983) );
  NANDN U7448 ( .A(n2981), .B(n2980), .Z(n2982) );
  NAND U7449 ( .A(n2983), .B(n2982), .Z(n5489) );
  XNOR U7450 ( .A(n5488), .B(n5489), .Z(n5491) );
  NANDN U7451 ( .A(n2985), .B(n2984), .Z(n2989) );
  NANDN U7452 ( .A(n2987), .B(n2986), .Z(n2988) );
  AND U7453 ( .A(n2989), .B(n2988), .Z(n5490) );
  XOR U7454 ( .A(n5491), .B(n5490), .Z(n5761) );
  XOR U7455 ( .A(n5907), .B(n5906), .Z(n5909) );
  XOR U7456 ( .A(n5909), .B(n5908), .Z(n5759) );
  NANDN U7457 ( .A(n3003), .B(n3002), .Z(n3007) );
  NANDN U7458 ( .A(n3005), .B(n3004), .Z(n3006) );
  NAND U7459 ( .A(n3007), .B(n3006), .Z(n5758) );
  XNOR U7460 ( .A(n5759), .B(n5758), .Z(n5760) );
  XNOR U7461 ( .A(n5761), .B(n5760), .Z(n6598) );
  NANDN U7462 ( .A(n3013), .B(n3012), .Z(n3017) );
  NANDN U7463 ( .A(n3015), .B(n3014), .Z(n3016) );
  AND U7464 ( .A(n3017), .B(n3016), .Z(n5653) );
  NANDN U7465 ( .A(n3019), .B(n3018), .Z(n3023) );
  NANDN U7466 ( .A(n3021), .B(n3020), .Z(n3022) );
  NAND U7467 ( .A(n3023), .B(n3022), .Z(n5654) );
  XNOR U7468 ( .A(n5653), .B(n5654), .Z(n5656) );
  NANDN U7469 ( .A(n3025), .B(n3024), .Z(n3029) );
  NAND U7470 ( .A(n3027), .B(n3026), .Z(n3028) );
  AND U7471 ( .A(n3029), .B(n3028), .Z(n5655) );
  XOR U7472 ( .A(n5656), .B(n5655), .Z(n5783) );
  XNOR U7473 ( .A(n5783), .B(n5782), .Z(n5784) );
  XNOR U7474 ( .A(n5785), .B(n5784), .Z(n6596) );
  NANDN U7475 ( .A(n3035), .B(n3034), .Z(n3039) );
  NAND U7476 ( .A(n3037), .B(n3036), .Z(n3038) );
  AND U7477 ( .A(n3039), .B(n3038), .Z(n5713) );
  NANDN U7478 ( .A(n3041), .B(n3040), .Z(n3045) );
  NANDN U7479 ( .A(n3043), .B(n3042), .Z(n3044) );
  NAND U7480 ( .A(n3045), .B(n3044), .Z(n5714) );
  XNOR U7481 ( .A(n5713), .B(n5714), .Z(n5716) );
  NANDN U7482 ( .A(n3047), .B(n3046), .Z(n3051) );
  NANDN U7483 ( .A(n3049), .B(n3048), .Z(n3050) );
  AND U7484 ( .A(n3051), .B(n3050), .Z(n5715) );
  XOR U7485 ( .A(n5716), .B(n5715), .Z(n5779) );
  NANDN U7486 ( .A(n3053), .B(n3052), .Z(n3057) );
  NAND U7487 ( .A(n3055), .B(n3054), .Z(n3056) );
  AND U7488 ( .A(n3057), .B(n3056), .Z(n5677) );
  NANDN U7489 ( .A(n3059), .B(n3058), .Z(n3063) );
  NANDN U7490 ( .A(n3061), .B(n3060), .Z(n3062) );
  NAND U7491 ( .A(n3063), .B(n3062), .Z(n5678) );
  XNOR U7492 ( .A(n5677), .B(n5678), .Z(n5680) );
  NANDN U7493 ( .A(n3065), .B(n3064), .Z(n3069) );
  NANDN U7494 ( .A(n3067), .B(n3066), .Z(n3068) );
  AND U7495 ( .A(n3069), .B(n3068), .Z(n5679) );
  XOR U7496 ( .A(n5680), .B(n5679), .Z(n5777) );
  NANDN U7497 ( .A(n3071), .B(n3070), .Z(n3075) );
  NANDN U7498 ( .A(n3073), .B(n3072), .Z(n3074) );
  AND U7499 ( .A(n3075), .B(n3074), .Z(n5506) );
  NANDN U7500 ( .A(n3077), .B(n3076), .Z(n3081) );
  NANDN U7501 ( .A(n3079), .B(n3078), .Z(n3080) );
  NAND U7502 ( .A(n3081), .B(n3080), .Z(n5507) );
  XNOR U7503 ( .A(n5506), .B(n5507), .Z(n5509) );
  NANDN U7504 ( .A(n3083), .B(n3082), .Z(n3087) );
  NANDN U7505 ( .A(n3085), .B(n3084), .Z(n3086) );
  AND U7506 ( .A(n3087), .B(n3086), .Z(n5508) );
  XNOR U7507 ( .A(n5509), .B(n5508), .Z(n5776) );
  XNOR U7508 ( .A(n5777), .B(n5776), .Z(n5778) );
  XNOR U7509 ( .A(n5779), .B(n5778), .Z(n6595) );
  XOR U7510 ( .A(n6596), .B(n6595), .Z(n6597) );
  XOR U7511 ( .A(n6598), .B(n6597), .Z(n6131) );
  XOR U7512 ( .A(n6132), .B(n6131), .Z(n5816) );
  XOR U7513 ( .A(n5817), .B(n5816), .Z(n5819) );
  XOR U7514 ( .A(n5818), .B(n5819), .Z(n5293) );
  NANDN U7515 ( .A(n3101), .B(n3100), .Z(n3105) );
  NANDN U7516 ( .A(n3103), .B(n3102), .Z(n3104) );
  AND U7517 ( .A(n3105), .B(n3104), .Z(n7273) );
  NANDN U7518 ( .A(n3107), .B(n3106), .Z(n3111) );
  NANDN U7519 ( .A(n3109), .B(n3108), .Z(n3110) );
  NAND U7520 ( .A(n3111), .B(n3110), .Z(n7274) );
  XNOR U7521 ( .A(n7273), .B(n7274), .Z(n7276) );
  NANDN U7522 ( .A(n3113), .B(n3112), .Z(n3117) );
  NANDN U7523 ( .A(n3115), .B(n3114), .Z(n3116) );
  AND U7524 ( .A(n3117), .B(n3116), .Z(n7275) );
  XOR U7525 ( .A(n7276), .B(n7275), .Z(n5309) );
  NAND U7526 ( .A(n3119), .B(n3118), .Z(n3123) );
  NAND U7527 ( .A(n3121), .B(n3120), .Z(n3122) );
  NAND U7528 ( .A(n3123), .B(n3122), .Z(n5308) );
  XNOR U7529 ( .A(n5309), .B(n5308), .Z(n5310) );
  XOR U7530 ( .A(n5311), .B(n5310), .Z(n6990) );
  XOR U7531 ( .A(n6989), .B(n6990), .Z(n6992) );
  XNOR U7532 ( .A(n6991), .B(n6992), .Z(n5823) );
  NANDN U7533 ( .A(n3125), .B(n3124), .Z(n3129) );
  NAND U7534 ( .A(n3127), .B(n3126), .Z(n3128) );
  NAND U7535 ( .A(n3129), .B(n3128), .Z(n5366) );
  NANDN U7536 ( .A(n3131), .B(n3130), .Z(n3135) );
  NANDN U7537 ( .A(n3133), .B(n3132), .Z(n3134) );
  AND U7538 ( .A(n3135), .B(n3134), .Z(n7279) );
  NANDN U7539 ( .A(n3137), .B(n3136), .Z(n3141) );
  NANDN U7540 ( .A(n3139), .B(n3138), .Z(n3140) );
  NAND U7541 ( .A(n3141), .B(n3140), .Z(n7280) );
  XNOR U7542 ( .A(n7279), .B(n7280), .Z(n7281) );
  NANDN U7543 ( .A(n3143), .B(n3142), .Z(n3147) );
  NANDN U7544 ( .A(n3145), .B(n3144), .Z(n3146) );
  NAND U7545 ( .A(n3147), .B(n3146), .Z(n7282) );
  XOR U7546 ( .A(n7281), .B(n7282), .Z(n5364) );
  NANDN U7547 ( .A(n3149), .B(n3148), .Z(n3153) );
  NAND U7548 ( .A(n3151), .B(n3150), .Z(n3152) );
  NAND U7549 ( .A(n3153), .B(n3152), .Z(n5365) );
  XOR U7550 ( .A(n5364), .B(n5365), .Z(n5367) );
  XOR U7551 ( .A(n5366), .B(n5367), .Z(n6548) );
  NANDN U7552 ( .A(n3155), .B(n3154), .Z(n3159) );
  NAND U7553 ( .A(n3157), .B(n3156), .Z(n3158) );
  NAND U7554 ( .A(n3159), .B(n3158), .Z(n5344) );
  NANDN U7555 ( .A(n3161), .B(n3160), .Z(n3165) );
  NANDN U7556 ( .A(n3163), .B(n3162), .Z(n3164) );
  AND U7557 ( .A(n3165), .B(n3164), .Z(n7253) );
  NANDN U7558 ( .A(n3167), .B(n3166), .Z(n3171) );
  NAND U7559 ( .A(n3169), .B(n3168), .Z(n3170) );
  NAND U7560 ( .A(n3171), .B(n3170), .Z(n7254) );
  XNOR U7561 ( .A(n7253), .B(n7254), .Z(n7255) );
  NANDN U7562 ( .A(n3173), .B(n3172), .Z(n3177) );
  NAND U7563 ( .A(n3175), .B(n3174), .Z(n3176) );
  NAND U7564 ( .A(n3177), .B(n3176), .Z(n7256) );
  XOR U7565 ( .A(n7255), .B(n7256), .Z(n5342) );
  NANDN U7566 ( .A(n3179), .B(n3178), .Z(n3183) );
  NAND U7567 ( .A(n3181), .B(n3180), .Z(n3182) );
  NAND U7568 ( .A(n3183), .B(n3182), .Z(n5343) );
  XOR U7569 ( .A(n5342), .B(n5343), .Z(n5345) );
  XOR U7570 ( .A(n5344), .B(n5345), .Z(n6546) );
  NANDN U7571 ( .A(n3185), .B(n3184), .Z(n3189) );
  NAND U7572 ( .A(n3187), .B(n3186), .Z(n3188) );
  NAND U7573 ( .A(n3189), .B(n3188), .Z(n7097) );
  NANDN U7574 ( .A(n3191), .B(n3190), .Z(n3195) );
  NANDN U7575 ( .A(n3193), .B(n3192), .Z(n3194) );
  AND U7576 ( .A(n3195), .B(n3194), .Z(n7295) );
  NANDN U7577 ( .A(n3197), .B(n3196), .Z(n3201) );
  NANDN U7578 ( .A(n3199), .B(n3198), .Z(n3200) );
  NAND U7579 ( .A(n3201), .B(n3200), .Z(n7296) );
  XNOR U7580 ( .A(n7295), .B(n7296), .Z(n7297) );
  NANDN U7581 ( .A(n3203), .B(n3202), .Z(n3207) );
  NANDN U7582 ( .A(n3205), .B(n3204), .Z(n3206) );
  NAND U7583 ( .A(n3207), .B(n3206), .Z(n7298) );
  XOR U7584 ( .A(n7297), .B(n7298), .Z(n7095) );
  NANDN U7585 ( .A(n3209), .B(n3208), .Z(n3213) );
  NAND U7586 ( .A(n3211), .B(n3210), .Z(n3212) );
  NAND U7587 ( .A(n3213), .B(n3212), .Z(n7096) );
  XOR U7588 ( .A(n7095), .B(n7096), .Z(n7098) );
  XOR U7589 ( .A(n7097), .B(n7098), .Z(n6545) );
  XOR U7590 ( .A(n6546), .B(n6545), .Z(n6547) );
  XOR U7591 ( .A(n6548), .B(n6547), .Z(n5822) );
  XOR U7592 ( .A(n5823), .B(n5822), .Z(n5825) );
  NANDN U7593 ( .A(n3215), .B(n3214), .Z(n3219) );
  NANDN U7594 ( .A(n3217), .B(n3216), .Z(n3218) );
  AND U7595 ( .A(n3219), .B(n3218), .Z(n5611) );
  NANDN U7596 ( .A(n3221), .B(n3220), .Z(n3225) );
  NANDN U7597 ( .A(n3223), .B(n3222), .Z(n3224) );
  NAND U7598 ( .A(n3225), .B(n3224), .Z(n5612) );
  XNOR U7599 ( .A(n5611), .B(n5612), .Z(n5613) );
  NANDN U7600 ( .A(n3227), .B(n3226), .Z(n3231) );
  NANDN U7601 ( .A(n3229), .B(n3228), .Z(n3230) );
  NAND U7602 ( .A(n3231), .B(n3230), .Z(n5614) );
  XOR U7603 ( .A(n5613), .B(n5614), .Z(n5348) );
  NANDN U7604 ( .A(n3233), .B(n3232), .Z(n3237) );
  NANDN U7605 ( .A(n3235), .B(n3234), .Z(n3236) );
  AND U7606 ( .A(n3237), .B(n3236), .Z(n5631) );
  NANDN U7607 ( .A(n3239), .B(n3238), .Z(n3243) );
  NANDN U7608 ( .A(n3241), .B(n3240), .Z(n3242) );
  NAND U7609 ( .A(n3243), .B(n3242), .Z(n5632) );
  XNOR U7610 ( .A(n5631), .B(n5632), .Z(n5633) );
  NANDN U7611 ( .A(n3245), .B(n3244), .Z(n3249) );
  NANDN U7612 ( .A(n3247), .B(n3246), .Z(n3248) );
  NAND U7613 ( .A(n3249), .B(n3248), .Z(n5634) );
  XOR U7614 ( .A(n5633), .B(n5634), .Z(n5346) );
  NANDN U7615 ( .A(n3251), .B(n3250), .Z(n3255) );
  NAND U7616 ( .A(n3253), .B(n3252), .Z(n3254) );
  NAND U7617 ( .A(n3255), .B(n3254), .Z(n5347) );
  XOR U7618 ( .A(n5346), .B(n5347), .Z(n5349) );
  XOR U7619 ( .A(n5348), .B(n5349), .Z(n6564) );
  NANDN U7620 ( .A(n3257), .B(n3256), .Z(n3261) );
  NANDN U7621 ( .A(n3259), .B(n3258), .Z(n3260) );
  AND U7622 ( .A(n3261), .B(n3260), .Z(n5625) );
  NANDN U7623 ( .A(n3263), .B(n3262), .Z(n3267) );
  NANDN U7624 ( .A(n3265), .B(n3264), .Z(n3266) );
  NAND U7625 ( .A(n3267), .B(n3266), .Z(n5626) );
  XNOR U7626 ( .A(n5625), .B(n5626), .Z(n5627) );
  NANDN U7627 ( .A(n3269), .B(n3268), .Z(n3273) );
  NANDN U7628 ( .A(n3271), .B(n3270), .Z(n3272) );
  NAND U7629 ( .A(n3273), .B(n3272), .Z(n5628) );
  XOR U7630 ( .A(n5627), .B(n5628), .Z(n5352) );
  NANDN U7631 ( .A(n3275), .B(n3274), .Z(n3279) );
  NANDN U7632 ( .A(n3277), .B(n3276), .Z(n3278) );
  AND U7633 ( .A(n3279), .B(n3278), .Z(n5464) );
  NANDN U7634 ( .A(n3281), .B(n3280), .Z(n3285) );
  NANDN U7635 ( .A(n3283), .B(n3282), .Z(n3284) );
  NAND U7636 ( .A(n3285), .B(n3284), .Z(n5465) );
  XNOR U7637 ( .A(n5464), .B(n5465), .Z(n5466) );
  NANDN U7638 ( .A(n3287), .B(n3286), .Z(n3291) );
  NANDN U7639 ( .A(n3289), .B(n3288), .Z(n3290) );
  NAND U7640 ( .A(n3291), .B(n3290), .Z(n5467) );
  XOR U7641 ( .A(n5466), .B(n5467), .Z(n5350) );
  NANDN U7642 ( .A(n3293), .B(n3292), .Z(n3297) );
  NAND U7643 ( .A(n3295), .B(n3294), .Z(n3296) );
  NAND U7644 ( .A(n3297), .B(n3296), .Z(n5351) );
  XOR U7645 ( .A(n5350), .B(n5351), .Z(n5353) );
  XOR U7646 ( .A(n5352), .B(n5353), .Z(n6562) );
  NANDN U7647 ( .A(n3299), .B(n3298), .Z(n3303) );
  NANDN U7648 ( .A(n3301), .B(n3300), .Z(n3302) );
  AND U7649 ( .A(n3303), .B(n3302), .Z(n5458) );
  NANDN U7650 ( .A(n3305), .B(n3304), .Z(n3309) );
  NANDN U7651 ( .A(n3307), .B(n3306), .Z(n3308) );
  NAND U7652 ( .A(n3309), .B(n3308), .Z(n5459) );
  XNOR U7653 ( .A(n5458), .B(n5459), .Z(n5460) );
  NANDN U7654 ( .A(n3311), .B(n3310), .Z(n3315) );
  NANDN U7655 ( .A(n3313), .B(n3312), .Z(n3314) );
  NAND U7656 ( .A(n3315), .B(n3314), .Z(n5461) );
  XOR U7657 ( .A(n5460), .B(n5461), .Z(n7079) );
  NANDN U7658 ( .A(n3317), .B(n3316), .Z(n3321) );
  NAND U7659 ( .A(n3319), .B(n3318), .Z(n3320) );
  NAND U7660 ( .A(n3321), .B(n3320), .Z(n7078) );
  NANDN U7661 ( .A(n3323), .B(n3322), .Z(n3327) );
  NANDN U7662 ( .A(n3325), .B(n3324), .Z(n3326) );
  AND U7663 ( .A(n3327), .B(n3326), .Z(n5476) );
  NANDN U7664 ( .A(n3329), .B(n3328), .Z(n3333) );
  NANDN U7665 ( .A(n3331), .B(n3330), .Z(n3332) );
  NAND U7666 ( .A(n3333), .B(n3332), .Z(n5477) );
  XNOR U7667 ( .A(n5476), .B(n5477), .Z(n5479) );
  NANDN U7668 ( .A(n3335), .B(n3334), .Z(n3339) );
  NANDN U7669 ( .A(n3337), .B(n3336), .Z(n3338) );
  AND U7670 ( .A(n3339), .B(n3338), .Z(n5478) );
  XNOR U7671 ( .A(n5479), .B(n5478), .Z(n7077) );
  XOR U7672 ( .A(n7078), .B(n7077), .Z(n7080) );
  XOR U7673 ( .A(n7079), .B(n7080), .Z(n6561) );
  XOR U7674 ( .A(n6562), .B(n6561), .Z(n6563) );
  XOR U7675 ( .A(n6564), .B(n6563), .Z(n5824) );
  XOR U7676 ( .A(n5825), .B(n5824), .Z(n7070) );
  NANDN U7677 ( .A(n3341), .B(n3340), .Z(n3345) );
  NANDN U7678 ( .A(n3343), .B(n3342), .Z(n3344) );
  AND U7679 ( .A(n3345), .B(n3344), .Z(n5596) );
  NANDN U7680 ( .A(n3347), .B(n3346), .Z(n3351) );
  NANDN U7681 ( .A(n3349), .B(n3348), .Z(n3350) );
  AND U7682 ( .A(n3351), .B(n3350), .Z(n5595) );
  XOR U7683 ( .A(n5596), .B(n5595), .Z(n5598) );
  NANDN U7684 ( .A(n3353), .B(n3352), .Z(n3357) );
  NANDN U7685 ( .A(n3355), .B(n3354), .Z(n3356) );
  AND U7686 ( .A(n3357), .B(n3356), .Z(n5597) );
  XOR U7687 ( .A(n5598), .B(n5597), .Z(n5377) );
  NANDN U7688 ( .A(n3359), .B(n3358), .Z(n3363) );
  NANDN U7689 ( .A(n3361), .B(n3360), .Z(n3362) );
  AND U7690 ( .A(n3363), .B(n3362), .Z(n6425) );
  NANDN U7691 ( .A(n3365), .B(n3364), .Z(n3369) );
  NAND U7692 ( .A(n3367), .B(n3366), .Z(n3368) );
  AND U7693 ( .A(n3369), .B(n3368), .Z(n6426) );
  XOR U7694 ( .A(n6425), .B(n6426), .Z(n6428) );
  NANDN U7695 ( .A(n3371), .B(n3370), .Z(n3375) );
  NANDN U7696 ( .A(n3373), .B(n3372), .Z(n3374) );
  AND U7697 ( .A(n3375), .B(n3374), .Z(n6427) );
  XOR U7698 ( .A(n6428), .B(n6427), .Z(n5375) );
  NANDN U7699 ( .A(n3377), .B(n3376), .Z(n3381) );
  NANDN U7700 ( .A(n3379), .B(n3378), .Z(n3380) );
  AND U7701 ( .A(n3381), .B(n3380), .Z(n6474) );
  NANDN U7702 ( .A(n3383), .B(n3382), .Z(n3387) );
  NANDN U7703 ( .A(n3385), .B(n3384), .Z(n3386) );
  AND U7704 ( .A(n3387), .B(n3386), .Z(n6473) );
  XOR U7705 ( .A(n6474), .B(n6473), .Z(n6476) );
  NANDN U7706 ( .A(n3389), .B(n3388), .Z(n3393) );
  NANDN U7707 ( .A(n3391), .B(n3390), .Z(n3392) );
  AND U7708 ( .A(n3393), .B(n3392), .Z(n6475) );
  XNOR U7709 ( .A(n6476), .B(n6475), .Z(n5374) );
  XNOR U7710 ( .A(n5375), .B(n5374), .Z(n5376) );
  XNOR U7711 ( .A(n5377), .B(n5376), .Z(n6199) );
  NANDN U7712 ( .A(n3395), .B(n3394), .Z(n3399) );
  NANDN U7713 ( .A(n3397), .B(n3396), .Z(n3398) );
  AND U7714 ( .A(n3399), .B(n3398), .Z(n6448) );
  NANDN U7715 ( .A(n3401), .B(n3400), .Z(n3405) );
  NANDN U7716 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U7717 ( .A(n3405), .B(n3404), .Z(n6447) );
  XOR U7718 ( .A(n6448), .B(n6447), .Z(n6450) );
  NANDN U7719 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U7720 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U7721 ( .A(n3411), .B(n3410), .Z(n6449) );
  XOR U7722 ( .A(n6450), .B(n6449), .Z(n7360) );
  NANDN U7723 ( .A(n3413), .B(n3412), .Z(n3417) );
  NANDN U7724 ( .A(n3415), .B(n3414), .Z(n3416) );
  AND U7725 ( .A(n3417), .B(n3416), .Z(n6854) );
  XOR U7726 ( .A(n6854), .B(n6853), .Z(n6856) );
  XOR U7727 ( .A(n6856), .B(n6855), .Z(n7358) );
  XNOR U7728 ( .A(n7358), .B(n7357), .Z(n7359) );
  XOR U7729 ( .A(n7360), .B(n7359), .Z(n6200) );
  XNOR U7730 ( .A(n6199), .B(n6200), .Z(n6201) );
  NANDN U7731 ( .A(n3435), .B(n3434), .Z(n3439) );
  NAND U7732 ( .A(n3437), .B(n3436), .Z(n3438) );
  AND U7733 ( .A(n3439), .B(n3438), .Z(n6342) );
  NAND U7734 ( .A(n3441), .B(n3440), .Z(n3445) );
  NAND U7735 ( .A(n3443), .B(n3442), .Z(n3444) );
  AND U7736 ( .A(n3445), .B(n3444), .Z(n6341) );
  XOR U7737 ( .A(n6342), .B(n6341), .Z(n6344) );
  NAND U7738 ( .A(n3447), .B(n3446), .Z(n3451) );
  NAND U7739 ( .A(n3449), .B(n3448), .Z(n3450) );
  AND U7740 ( .A(n3451), .B(n3450), .Z(n6343) );
  XOR U7741 ( .A(n6344), .B(n6343), .Z(n7346) );
  NANDN U7742 ( .A(n3453), .B(n3452), .Z(n3457) );
  NANDN U7743 ( .A(n3455), .B(n3454), .Z(n3456) );
  AND U7744 ( .A(n3457), .B(n3456), .Z(n6658) );
  NANDN U7745 ( .A(n3459), .B(n3458), .Z(n3463) );
  NANDN U7746 ( .A(n3461), .B(n3460), .Z(n3462) );
  AND U7747 ( .A(n3463), .B(n3462), .Z(n6657) );
  XOR U7748 ( .A(n6658), .B(n6657), .Z(n6660) );
  NANDN U7749 ( .A(n3465), .B(n3464), .Z(n3469) );
  NANDN U7750 ( .A(n3467), .B(n3466), .Z(n3468) );
  AND U7751 ( .A(n3469), .B(n3468), .Z(n6659) );
  XNOR U7752 ( .A(n6660), .B(n6659), .Z(n7345) );
  XNOR U7753 ( .A(n7346), .B(n7345), .Z(n7347) );
  XOR U7754 ( .A(n7348), .B(n7347), .Z(n6202) );
  XOR U7755 ( .A(n6201), .B(n6202), .Z(n6371) );
  XNOR U7756 ( .A(n6111), .B(n6112), .Z(n6113) );
  XOR U7757 ( .A(n6113), .B(n6114), .Z(n5400) );
  XNOR U7758 ( .A(n6441), .B(n6442), .Z(n6443) );
  XOR U7759 ( .A(n6443), .B(n6444), .Z(n5399) );
  NANDN U7760 ( .A(n3495), .B(n3494), .Z(n3499) );
  NAND U7761 ( .A(n3497), .B(n3496), .Z(n3498) );
  NAND U7762 ( .A(n3499), .B(n3498), .Z(n5398) );
  XOR U7763 ( .A(n5399), .B(n5398), .Z(n5401) );
  XOR U7764 ( .A(n5400), .B(n5401), .Z(n6832) );
  XNOR U7765 ( .A(n6105), .B(n6106), .Z(n6107) );
  XOR U7766 ( .A(n6107), .B(n6108), .Z(n5394) );
  NANDN U7767 ( .A(n3517), .B(n3516), .Z(n3521) );
  NANDN U7768 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U7769 ( .A(n3521), .B(n3520), .Z(n6398) );
  XNOR U7770 ( .A(n6397), .B(n6398), .Z(n6399) );
  XOR U7771 ( .A(n6399), .B(n6400), .Z(n5393) );
  NANDN U7772 ( .A(n3527), .B(n3526), .Z(n3531) );
  NAND U7773 ( .A(n3529), .B(n3528), .Z(n3530) );
  AND U7774 ( .A(n3531), .B(n3530), .Z(n6647) );
  NANDN U7775 ( .A(n3533), .B(n3532), .Z(n3537) );
  NANDN U7776 ( .A(n3535), .B(n3534), .Z(n3536) );
  NAND U7777 ( .A(n3537), .B(n3536), .Z(n6648) );
  XNOR U7778 ( .A(n6647), .B(n6648), .Z(n6650) );
  NANDN U7779 ( .A(n3539), .B(n3538), .Z(n3543) );
  NAND U7780 ( .A(n3541), .B(n3540), .Z(n3542) );
  AND U7781 ( .A(n3543), .B(n3542), .Z(n6649) );
  XNOR U7782 ( .A(n6650), .B(n6649), .Z(n5392) );
  XOR U7783 ( .A(n5393), .B(n5392), .Z(n5395) );
  XOR U7784 ( .A(n5394), .B(n5395), .Z(n6831) );
  XOR U7785 ( .A(n6832), .B(n6831), .Z(n6834) );
  XNOR U7786 ( .A(n6661), .B(n6662), .Z(n6663) );
  XOR U7787 ( .A(n6663), .B(n6664), .Z(n5330) );
  NANDN U7788 ( .A(n3557), .B(n3556), .Z(n3561) );
  NAND U7789 ( .A(n3559), .B(n3558), .Z(n3560) );
  AND U7790 ( .A(n3561), .B(n3560), .Z(n6347) );
  NAND U7791 ( .A(n3563), .B(n3562), .Z(n3567) );
  NAND U7792 ( .A(n3565), .B(n3564), .Z(n3566) );
  NAND U7793 ( .A(n3567), .B(n3566), .Z(n6348) );
  XNOR U7794 ( .A(n6347), .B(n6348), .Z(n6349) );
  NAND U7795 ( .A(n3569), .B(n3568), .Z(n3573) );
  NAND U7796 ( .A(n3571), .B(n3570), .Z(n3572) );
  NAND U7797 ( .A(n3573), .B(n3572), .Z(n6350) );
  XOR U7798 ( .A(n6349), .B(n6350), .Z(n5329) );
  XNOR U7799 ( .A(n6641), .B(n6642), .Z(n6644) );
  XNOR U7800 ( .A(n6644), .B(n6643), .Z(n5328) );
  XOR U7801 ( .A(n5329), .B(n5328), .Z(n5331) );
  XOR U7802 ( .A(n5330), .B(n5331), .Z(n6833) );
  XOR U7803 ( .A(n6834), .B(n6833), .Z(n6370) );
  NANDN U7804 ( .A(n3591), .B(n3590), .Z(n3595) );
  NANDN U7805 ( .A(n3593), .B(n3592), .Z(n3594) );
  NAND U7806 ( .A(n3595), .B(n3594), .Z(n6708) );
  XNOR U7807 ( .A(n6707), .B(n6708), .Z(n6709) );
  NANDN U7808 ( .A(n3597), .B(n3596), .Z(n3601) );
  NANDN U7809 ( .A(n3599), .B(n3598), .Z(n3600) );
  NAND U7810 ( .A(n3601), .B(n3600), .Z(n6710) );
  XOR U7811 ( .A(n6709), .B(n6710), .Z(n5336) );
  NANDN U7812 ( .A(n3607), .B(n3606), .Z(n3611) );
  NANDN U7813 ( .A(n3609), .B(n3608), .Z(n3610) );
  NAND U7814 ( .A(n3611), .B(n3610), .Z(n6003) );
  XNOR U7815 ( .A(n6002), .B(n6003), .Z(n6004) );
  NANDN U7816 ( .A(n3613), .B(n3612), .Z(n3617) );
  NANDN U7817 ( .A(n3615), .B(n3614), .Z(n3616) );
  NAND U7818 ( .A(n3617), .B(n3616), .Z(n6005) );
  XOR U7819 ( .A(n6004), .B(n6005), .Z(n5334) );
  NANDN U7820 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U7821 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U7822 ( .A(n3623), .B(n3622), .Z(n5335) );
  XOR U7823 ( .A(n5334), .B(n5335), .Z(n5337) );
  XOR U7824 ( .A(n5336), .B(n5337), .Z(n6302) );
  NANDN U7825 ( .A(n3625), .B(n3624), .Z(n3629) );
  NAND U7826 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U7827 ( .A(n3629), .B(n3628), .Z(n5316) );
  NANDN U7828 ( .A(n3631), .B(n3630), .Z(n3635) );
  NANDN U7829 ( .A(n3633), .B(n3632), .Z(n3634) );
  AND U7830 ( .A(n3635), .B(n3634), .Z(n6277) );
  NANDN U7831 ( .A(n3637), .B(n3636), .Z(n3641) );
  NANDN U7832 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U7833 ( .A(n3641), .B(n3640), .Z(n6278) );
  XNOR U7834 ( .A(n6277), .B(n6278), .Z(n6279) );
  NANDN U7835 ( .A(n3643), .B(n3642), .Z(n3647) );
  NANDN U7836 ( .A(n3645), .B(n3644), .Z(n3646) );
  NAND U7837 ( .A(n3647), .B(n3646), .Z(n6280) );
  XOR U7838 ( .A(n6279), .B(n6280), .Z(n5314) );
  NANDN U7839 ( .A(n3649), .B(n3648), .Z(n3653) );
  NANDN U7840 ( .A(n3651), .B(n3650), .Z(n3652) );
  NAND U7841 ( .A(n3653), .B(n3652), .Z(n5315) );
  XOR U7842 ( .A(n5314), .B(n5315), .Z(n5317) );
  XOR U7843 ( .A(n5316), .B(n5317), .Z(n6301) );
  XOR U7844 ( .A(n6302), .B(n6301), .Z(n6304) );
  NANDN U7845 ( .A(n3655), .B(n3654), .Z(n3659) );
  NANDN U7846 ( .A(n3657), .B(n3656), .Z(n3658) );
  NAND U7847 ( .A(n3659), .B(n3658), .Z(n5326) );
  NANDN U7848 ( .A(n3661), .B(n3660), .Z(n3665) );
  NANDN U7849 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U7850 ( .A(n3665), .B(n3664), .Z(n6283) );
  NANDN U7851 ( .A(n3667), .B(n3666), .Z(n3671) );
  NAND U7852 ( .A(n3669), .B(n3668), .Z(n3670) );
  NAND U7853 ( .A(n3671), .B(n3670), .Z(n6284) );
  XNOR U7854 ( .A(n6283), .B(n6284), .Z(n6285) );
  NANDN U7855 ( .A(n3673), .B(n3672), .Z(n3677) );
  NAND U7856 ( .A(n3675), .B(n3674), .Z(n3676) );
  NAND U7857 ( .A(n3677), .B(n3676), .Z(n6286) );
  XOR U7858 ( .A(n6285), .B(n6286), .Z(n5324) );
  NANDN U7859 ( .A(n3679), .B(n3678), .Z(n3683) );
  NANDN U7860 ( .A(n3681), .B(n3680), .Z(n3682) );
  NAND U7861 ( .A(n3683), .B(n3682), .Z(n5325) );
  XOR U7862 ( .A(n5324), .B(n5325), .Z(n5327) );
  XOR U7863 ( .A(n5326), .B(n5327), .Z(n6303) );
  XNOR U7864 ( .A(n6304), .B(n6303), .Z(n6369) );
  XOR U7865 ( .A(n6371), .B(n6372), .Z(n7067) );
  NANDN U7866 ( .A(n3685), .B(n3684), .Z(n3689) );
  NANDN U7867 ( .A(n3687), .B(n3686), .Z(n3688) );
  AND U7868 ( .A(n3689), .B(n3688), .Z(n6790) );
  NANDN U7869 ( .A(n3691), .B(n3690), .Z(n3695) );
  NANDN U7870 ( .A(n3693), .B(n3692), .Z(n3694) );
  NAND U7871 ( .A(n3695), .B(n3694), .Z(n5406) );
  XNOR U7872 ( .A(n6769), .B(n6770), .Z(n6771) );
  XOR U7873 ( .A(n6771), .B(n6772), .Z(n5404) );
  NANDN U7874 ( .A(n3709), .B(n3708), .Z(n3713) );
  NANDN U7875 ( .A(n3711), .B(n3710), .Z(n3712) );
  NAND U7876 ( .A(n3713), .B(n3712), .Z(n5405) );
  XOR U7877 ( .A(n5404), .B(n5405), .Z(n5407) );
  XOR U7878 ( .A(n5406), .B(n5407), .Z(n6788) );
  NANDN U7879 ( .A(n3715), .B(n3714), .Z(n3719) );
  NAND U7880 ( .A(n3717), .B(n3716), .Z(n3718) );
  NAND U7881 ( .A(n3719), .B(n3718), .Z(n5306) );
  NANDN U7882 ( .A(n3721), .B(n3720), .Z(n3725) );
  NANDN U7883 ( .A(n3723), .B(n3722), .Z(n3724) );
  AND U7884 ( .A(n3725), .B(n3724), .Z(n6247) );
  NANDN U7885 ( .A(n3727), .B(n3726), .Z(n3731) );
  NANDN U7886 ( .A(n3729), .B(n3728), .Z(n3730) );
  NAND U7887 ( .A(n3731), .B(n3730), .Z(n6248) );
  XNOR U7888 ( .A(n6247), .B(n6248), .Z(n6249) );
  NANDN U7889 ( .A(n3733), .B(n3732), .Z(n3737) );
  NANDN U7890 ( .A(n3735), .B(n3734), .Z(n3736) );
  NAND U7891 ( .A(n3737), .B(n3736), .Z(n6250) );
  XOR U7892 ( .A(n6249), .B(n6250), .Z(n5304) );
  NANDN U7893 ( .A(n3739), .B(n3738), .Z(n3743) );
  NAND U7894 ( .A(n3741), .B(n3740), .Z(n3742) );
  NAND U7895 ( .A(n3743), .B(n3742), .Z(n5305) );
  XOR U7896 ( .A(n5304), .B(n5305), .Z(n5307) );
  XOR U7897 ( .A(n5306), .B(n5307), .Z(n6787) );
  XOR U7898 ( .A(n6788), .B(n6787), .Z(n6789) );
  XOR U7899 ( .A(n6790), .B(n6789), .Z(n6438) );
  NANDN U7900 ( .A(n3745), .B(n3744), .Z(n3749) );
  NANDN U7901 ( .A(n3747), .B(n3746), .Z(n3748) );
  NAND U7902 ( .A(n3749), .B(n3748), .Z(n5362) );
  NANDN U7903 ( .A(n3751), .B(n3750), .Z(n3755) );
  NAND U7904 ( .A(n3753), .B(n3752), .Z(n3754) );
  AND U7905 ( .A(n3755), .B(n3754), .Z(n6763) );
  XNOR U7906 ( .A(n6763), .B(n6764), .Z(n6765) );
  XOR U7907 ( .A(n6765), .B(n6766), .Z(n5360) );
  NANDN U7908 ( .A(n3765), .B(n3764), .Z(n3769) );
  NANDN U7909 ( .A(n3767), .B(n3766), .Z(n3768) );
  NAND U7910 ( .A(n3769), .B(n3768), .Z(n5361) );
  XOR U7911 ( .A(n5360), .B(n5361), .Z(n5363) );
  XOR U7912 ( .A(n5362), .B(n5363), .Z(n6730) );
  NANDN U7913 ( .A(n3771), .B(n3770), .Z(n3775) );
  NAND U7914 ( .A(n3773), .B(n3772), .Z(n3774) );
  NAND U7915 ( .A(n3775), .B(n3774), .Z(n7105) );
  NANDN U7916 ( .A(n3777), .B(n3776), .Z(n3781) );
  NANDN U7917 ( .A(n3779), .B(n3778), .Z(n3780) );
  AND U7918 ( .A(n3781), .B(n3780), .Z(n6223) );
  NANDN U7919 ( .A(n3783), .B(n3782), .Z(n3787) );
  NANDN U7920 ( .A(n3785), .B(n3784), .Z(n3786) );
  NAND U7921 ( .A(n3787), .B(n3786), .Z(n6224) );
  XNOR U7922 ( .A(n6223), .B(n6224), .Z(n6225) );
  NANDN U7923 ( .A(n3789), .B(n3788), .Z(n3793) );
  NANDN U7924 ( .A(n3791), .B(n3790), .Z(n3792) );
  NAND U7925 ( .A(n3793), .B(n3792), .Z(n6226) );
  XOR U7926 ( .A(n6225), .B(n6226), .Z(n7103) );
  NANDN U7927 ( .A(n3795), .B(n3794), .Z(n3799) );
  NAND U7928 ( .A(n3797), .B(n3796), .Z(n3798) );
  NAND U7929 ( .A(n3799), .B(n3798), .Z(n7104) );
  XOR U7930 ( .A(n7103), .B(n7104), .Z(n7106) );
  XOR U7931 ( .A(n7105), .B(n7106), .Z(n6729) );
  XOR U7932 ( .A(n6730), .B(n6729), .Z(n6732) );
  NANDN U7933 ( .A(n3801), .B(n3800), .Z(n3805) );
  NAND U7934 ( .A(n3803), .B(n3802), .Z(n3804) );
  NAND U7935 ( .A(n3805), .B(n3804), .Z(n7093) );
  NANDN U7936 ( .A(n3807), .B(n3806), .Z(n3811) );
  NAND U7937 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U7938 ( .A(n3811), .B(n3810), .Z(n6217) );
  NANDN U7939 ( .A(n3813), .B(n3812), .Z(n3817) );
  NANDN U7940 ( .A(n3815), .B(n3814), .Z(n3816) );
  NAND U7941 ( .A(n3817), .B(n3816), .Z(n6218) );
  XNOR U7942 ( .A(n6217), .B(n6218), .Z(n6219) );
  NANDN U7943 ( .A(n3819), .B(n3818), .Z(n3823) );
  NANDN U7944 ( .A(n3821), .B(n3820), .Z(n3822) );
  NAND U7945 ( .A(n3823), .B(n3822), .Z(n6220) );
  XOR U7946 ( .A(n6219), .B(n6220), .Z(n7091) );
  NANDN U7947 ( .A(n3825), .B(n3824), .Z(n3829) );
  NAND U7948 ( .A(n3827), .B(n3826), .Z(n3828) );
  NAND U7949 ( .A(n3829), .B(n3828), .Z(n7092) );
  XOR U7950 ( .A(n7091), .B(n7092), .Z(n7094) );
  XOR U7951 ( .A(n7093), .B(n7094), .Z(n6731) );
  XOR U7952 ( .A(n6732), .B(n6731), .Z(n6436) );
  NANDN U7953 ( .A(n3831), .B(n3830), .Z(n3835) );
  NANDN U7954 ( .A(n3833), .B(n3832), .Z(n3834) );
  AND U7955 ( .A(n3835), .B(n3834), .Z(n5446) );
  NANDN U7956 ( .A(n3837), .B(n3836), .Z(n3841) );
  NANDN U7957 ( .A(n3839), .B(n3838), .Z(n3840) );
  NAND U7958 ( .A(n3841), .B(n3840), .Z(n5447) );
  XNOR U7959 ( .A(n5446), .B(n5447), .Z(n5448) );
  NANDN U7960 ( .A(n3843), .B(n3842), .Z(n3847) );
  NANDN U7961 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U7962 ( .A(n3847), .B(n3846), .Z(n5449) );
  XOR U7963 ( .A(n5448), .B(n5449), .Z(n7101) );
  NANDN U7964 ( .A(n3849), .B(n3848), .Z(n3853) );
  NANDN U7965 ( .A(n3851), .B(n3850), .Z(n3852) );
  AND U7966 ( .A(n3853), .B(n3852), .Z(n5524) );
  NANDN U7967 ( .A(n3855), .B(n3854), .Z(n3859) );
  NANDN U7968 ( .A(n3857), .B(n3856), .Z(n3858) );
  NAND U7969 ( .A(n3859), .B(n3858), .Z(n5525) );
  XNOR U7970 ( .A(n5524), .B(n5525), .Z(n5526) );
  NANDN U7971 ( .A(n3861), .B(n3860), .Z(n3865) );
  NANDN U7972 ( .A(n3863), .B(n3862), .Z(n3864) );
  NAND U7973 ( .A(n3865), .B(n3864), .Z(n5527) );
  XOR U7974 ( .A(n5526), .B(n5527), .Z(n7099) );
  NANDN U7975 ( .A(n3867), .B(n3866), .Z(n3871) );
  NAND U7976 ( .A(n3869), .B(n3868), .Z(n3870) );
  NAND U7977 ( .A(n3871), .B(n3870), .Z(n7100) );
  XOR U7978 ( .A(n7099), .B(n7100), .Z(n7102) );
  XOR U7979 ( .A(n7101), .B(n7102), .Z(n6626) );
  NANDN U7980 ( .A(n3877), .B(n3876), .Z(n3881) );
  NAND U7981 ( .A(n3879), .B(n3878), .Z(n3880) );
  NAND U7982 ( .A(n3881), .B(n3880), .Z(n6146) );
  XNOR U7983 ( .A(n6145), .B(n6146), .Z(n6147) );
  XOR U7984 ( .A(n6147), .B(n6148), .Z(n7089) );
  NANDN U7985 ( .A(n3887), .B(n3886), .Z(n3891) );
  NAND U7986 ( .A(n3889), .B(n3888), .Z(n3890) );
  AND U7987 ( .A(n3891), .B(n3890), .Z(n6151) );
  XNOR U7988 ( .A(n6151), .B(n6152), .Z(n6153) );
  NANDN U7989 ( .A(n3897), .B(n3896), .Z(n3901) );
  NANDN U7990 ( .A(n3899), .B(n3898), .Z(n3900) );
  NAND U7991 ( .A(n3901), .B(n3900), .Z(n6154) );
  XOR U7992 ( .A(n6153), .B(n6154), .Z(n7087) );
  NANDN U7993 ( .A(n3903), .B(n3902), .Z(n3907) );
  NAND U7994 ( .A(n3905), .B(n3904), .Z(n3906) );
  NAND U7995 ( .A(n3907), .B(n3906), .Z(n7088) );
  XOR U7996 ( .A(n7087), .B(n7088), .Z(n7090) );
  XOR U7997 ( .A(n7089), .B(n7090), .Z(n6624) );
  XNOR U7998 ( .A(n5892), .B(n5893), .Z(n5894) );
  XOR U7999 ( .A(n5894), .B(n5895), .Z(n7085) );
  NANDN U8000 ( .A(n3921), .B(n3920), .Z(n3925) );
  NAND U8001 ( .A(n3923), .B(n3922), .Z(n3924) );
  AND U8002 ( .A(n3925), .B(n3924), .Z(n6175) );
  NANDN U8003 ( .A(n3927), .B(n3926), .Z(n3931) );
  NANDN U8004 ( .A(n3929), .B(n3928), .Z(n3930) );
  NAND U8005 ( .A(n3931), .B(n3930), .Z(n6176) );
  XNOR U8006 ( .A(n6175), .B(n6176), .Z(n6177) );
  NANDN U8007 ( .A(n3933), .B(n3932), .Z(n3937) );
  NANDN U8008 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U8009 ( .A(n3937), .B(n3936), .Z(n6178) );
  XOR U8010 ( .A(n6177), .B(n6178), .Z(n7083) );
  NANDN U8011 ( .A(n3939), .B(n3938), .Z(n3943) );
  NAND U8012 ( .A(n3941), .B(n3940), .Z(n3942) );
  NAND U8013 ( .A(n3943), .B(n3942), .Z(n7084) );
  XOR U8014 ( .A(n7083), .B(n7084), .Z(n7086) );
  XOR U8015 ( .A(n7085), .B(n7086), .Z(n6623) );
  XOR U8016 ( .A(n6624), .B(n6623), .Z(n6625) );
  XNOR U8017 ( .A(n6626), .B(n6625), .Z(n6435) );
  XNOR U8018 ( .A(n6436), .B(n6435), .Z(n6437) );
  XOR U8019 ( .A(n6438), .B(n6437), .Z(n7068) );
  XNOR U8020 ( .A(n7067), .B(n7068), .Z(n7069) );
  XNOR U8021 ( .A(n7070), .B(n7069), .Z(n5292) );
  XOR U8022 ( .A(n5293), .B(n5292), .Z(n5295) );
  XOR U8023 ( .A(n5294), .B(n5295), .Z(n7443) );
  XOR U8024 ( .A(n7444), .B(n7443), .Z(n7446) );
  NANDN U8025 ( .A(n3945), .B(n3944), .Z(n3949) );
  NANDN U8026 ( .A(n3947), .B(n3946), .Z(n3948) );
  AND U8027 ( .A(n3949), .B(n3948), .Z(n7213) );
  NANDN U8028 ( .A(n3955), .B(n3954), .Z(n3959) );
  NANDN U8029 ( .A(n3957), .B(n3956), .Z(n3958) );
  AND U8030 ( .A(n3959), .B(n3958), .Z(n6323) );
  XOR U8031 ( .A(n6324), .B(n6323), .Z(n6326) );
  NANDN U8032 ( .A(n3961), .B(n3960), .Z(n3965) );
  NANDN U8033 ( .A(n3963), .B(n3962), .Z(n3964) );
  AND U8034 ( .A(n3965), .B(n3964), .Z(n6325) );
  XOR U8035 ( .A(n6326), .B(n6325), .Z(n7195) );
  NANDN U8036 ( .A(n3967), .B(n3966), .Z(n3971) );
  NANDN U8037 ( .A(n3969), .B(n3968), .Z(n3970) );
  AND U8038 ( .A(n3971), .B(n3970), .Z(n6689) );
  NANDN U8039 ( .A(n3973), .B(n3972), .Z(n3977) );
  NANDN U8040 ( .A(n3975), .B(n3974), .Z(n3976) );
  NAND U8041 ( .A(n3977), .B(n3976), .Z(n6690) );
  XNOR U8042 ( .A(n6689), .B(n6690), .Z(n6692) );
  NANDN U8043 ( .A(n3979), .B(n3978), .Z(n3983) );
  NANDN U8044 ( .A(n3981), .B(n3980), .Z(n3982) );
  AND U8045 ( .A(n3983), .B(n3982), .Z(n6691) );
  XOR U8046 ( .A(n6692), .B(n6691), .Z(n7194) );
  NANDN U8047 ( .A(n3985), .B(n3984), .Z(n3989) );
  NAND U8048 ( .A(n3987), .B(n3986), .Z(n3988) );
  NAND U8049 ( .A(n3989), .B(n3988), .Z(n7193) );
  XOR U8050 ( .A(n7194), .B(n7193), .Z(n7196) );
  XOR U8051 ( .A(n7195), .B(n7196), .Z(n7212) );
  OR U8052 ( .A(n3991), .B(n3990), .Z(n3995) );
  NANDN U8053 ( .A(n3993), .B(n3992), .Z(n3994) );
  NAND U8054 ( .A(n3995), .B(n3994), .Z(n7211) );
  XOR U8055 ( .A(n7212), .B(n7211), .Z(n7214) );
  XOR U8056 ( .A(n7213), .B(n7214), .Z(n7118) );
  NANDN U8057 ( .A(n3997), .B(n3996), .Z(n4001) );
  OR U8058 ( .A(n3999), .B(n3998), .Z(n4000) );
  AND U8059 ( .A(n4001), .B(n4000), .Z(n6611) );
  XOR U8060 ( .A(n7144), .B(n7143), .Z(n7146) );
  NANDN U8061 ( .A(n4011), .B(n4010), .Z(n4015) );
  NANDN U8062 ( .A(n4013), .B(n4012), .Z(n4014) );
  AND U8063 ( .A(n4015), .B(n4014), .Z(n7145) );
  XOR U8064 ( .A(n7146), .B(n7145), .Z(n5545) );
  XNOR U8065 ( .A(n7333), .B(n7334), .Z(n7336) );
  XOR U8066 ( .A(n7336), .B(n7335), .Z(n5543) );
  XNOR U8067 ( .A(n5543), .B(n5542), .Z(n5544) );
  XOR U8068 ( .A(n5545), .B(n5544), .Z(n6612) );
  XNOR U8069 ( .A(n6611), .B(n6612), .Z(n6613) );
  NANDN U8070 ( .A(n4037), .B(n4036), .Z(n4041) );
  NANDN U8071 ( .A(n4039), .B(n4038), .Z(n4040) );
  AND U8072 ( .A(n4041), .B(n4040), .Z(n6181) );
  NANDN U8073 ( .A(n4043), .B(n4042), .Z(n4047) );
  NANDN U8074 ( .A(n4045), .B(n4044), .Z(n4046) );
  NAND U8075 ( .A(n4047), .B(n4046), .Z(n6182) );
  XNOR U8076 ( .A(n6181), .B(n6182), .Z(n6184) );
  NANDN U8077 ( .A(n4049), .B(n4048), .Z(n4053) );
  NANDN U8078 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U8079 ( .A(n4053), .B(n4052), .Z(n6183) );
  XOR U8080 ( .A(n6184), .B(n6183), .Z(n5571) );
  XNOR U8081 ( .A(n5571), .B(n5570), .Z(n5572) );
  XOR U8082 ( .A(n5573), .B(n5572), .Z(n6614) );
  XNOR U8083 ( .A(n6613), .B(n6614), .Z(n7117) );
  XNOR U8084 ( .A(n7118), .B(n7117), .Z(n7120) );
  NANDN U8085 ( .A(n4067), .B(n4066), .Z(n4071) );
  NANDN U8086 ( .A(n4069), .B(n4068), .Z(n4070) );
  AND U8087 ( .A(n4071), .B(n4070), .Z(n5659) );
  NANDN U8088 ( .A(n4073), .B(n4072), .Z(n4077) );
  NANDN U8089 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U8090 ( .A(n4077), .B(n4076), .Z(n5660) );
  XNOR U8091 ( .A(n5659), .B(n5660), .Z(n5662) );
  NANDN U8092 ( .A(n4079), .B(n4078), .Z(n4083) );
  NANDN U8093 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U8094 ( .A(n4083), .B(n4082), .Z(n5661) );
  XOR U8095 ( .A(n5662), .B(n5661), .Z(n5791) );
  NANDN U8096 ( .A(n4089), .B(n4088), .Z(n4093) );
  NANDN U8097 ( .A(n4091), .B(n4090), .Z(n4092) );
  NAND U8098 ( .A(n4093), .B(n4092), .Z(n5684) );
  XNOR U8099 ( .A(n5683), .B(n5684), .Z(n5686) );
  NANDN U8100 ( .A(n4095), .B(n4094), .Z(n4099) );
  NANDN U8101 ( .A(n4097), .B(n4096), .Z(n4098) );
  AND U8102 ( .A(n4099), .B(n4098), .Z(n5685) );
  XOR U8103 ( .A(n5686), .B(n5685), .Z(n5789) );
  NANDN U8104 ( .A(n4101), .B(n4100), .Z(n4105) );
  NANDN U8105 ( .A(n4103), .B(n4102), .Z(n4104) );
  AND U8106 ( .A(n4105), .B(n4104), .Z(n5911) );
  XOR U8107 ( .A(n5911), .B(n5910), .Z(n5913) );
  NANDN U8108 ( .A(n4111), .B(n4110), .Z(n4115) );
  NANDN U8109 ( .A(n4113), .B(n4112), .Z(n4114) );
  AND U8110 ( .A(n4115), .B(n4114), .Z(n5912) );
  XNOR U8111 ( .A(n5913), .B(n5912), .Z(n5788) );
  XNOR U8112 ( .A(n5789), .B(n5788), .Z(n5790) );
  XOR U8113 ( .A(n5791), .B(n5790), .Z(n6606) );
  XOR U8114 ( .A(n6605), .B(n6606), .Z(n6608) );
  XNOR U8115 ( .A(n6607), .B(n6608), .Z(n7119) );
  XOR U8116 ( .A(n7120), .B(n7119), .Z(n7030) );
  NANDN U8117 ( .A(n4117), .B(n4116), .Z(n4121) );
  NAND U8118 ( .A(n4119), .B(n4118), .Z(n4120) );
  AND U8119 ( .A(n4121), .B(n4120), .Z(n7202) );
  NANDN U8120 ( .A(n4123), .B(n4122), .Z(n4127) );
  NAND U8121 ( .A(n4125), .B(n4124), .Z(n4126) );
  AND U8122 ( .A(n4127), .B(n4126), .Z(n7200) );
  XNOR U8123 ( .A(n7200), .B(n7199), .Z(n7201) );
  XNOR U8124 ( .A(n7202), .B(n7201), .Z(n5368) );
  XNOR U8125 ( .A(n5878), .B(n5879), .Z(n5881) );
  XOR U8126 ( .A(n5881), .B(n5880), .Z(n5455) );
  NANDN U8127 ( .A(n4149), .B(n4148), .Z(n4153) );
  NAND U8128 ( .A(n4151), .B(n4150), .Z(n4152) );
  NAND U8129 ( .A(n4153), .B(n4152), .Z(n5857) );
  NANDN U8130 ( .A(n4155), .B(n4154), .Z(n4159) );
  NANDN U8131 ( .A(n4157), .B(n4156), .Z(n4158) );
  AND U8132 ( .A(n4159), .B(n4158), .Z(n5858) );
  XOR U8133 ( .A(n5859), .B(n5858), .Z(n5453) );
  XNOR U8134 ( .A(n5453), .B(n5452), .Z(n5454) );
  XOR U8135 ( .A(n5455), .B(n5454), .Z(n5369) );
  XNOR U8136 ( .A(n5368), .B(n5369), .Z(n5370) );
  NANDN U8137 ( .A(n4165), .B(n4164), .Z(n4169) );
  OR U8138 ( .A(n4167), .B(n4166), .Z(n4168) );
  NAND U8139 ( .A(n4169), .B(n4168), .Z(n5371) );
  XNOR U8140 ( .A(n5370), .B(n5371), .Z(n5426) );
  NANDN U8141 ( .A(n4175), .B(n4174), .Z(n4179) );
  NANDN U8142 ( .A(n4177), .B(n4176), .Z(n4178) );
  AND U8143 ( .A(n4179), .B(n4178), .Z(n5707) );
  NANDN U8144 ( .A(n4181), .B(n4180), .Z(n4185) );
  NANDN U8145 ( .A(n4183), .B(n4182), .Z(n4184) );
  NAND U8146 ( .A(n4185), .B(n4184), .Z(n5708) );
  XNOR U8147 ( .A(n5707), .B(n5708), .Z(n5710) );
  NANDN U8148 ( .A(n4187), .B(n4186), .Z(n4191) );
  NANDN U8149 ( .A(n4189), .B(n4188), .Z(n4190) );
  AND U8150 ( .A(n4191), .B(n4190), .Z(n5709) );
  XOR U8151 ( .A(n5710), .B(n5709), .Z(n5642) );
  NANDN U8152 ( .A(n4193), .B(n4192), .Z(n4197) );
  NAND U8153 ( .A(n4195), .B(n4194), .Z(n4196) );
  NAND U8154 ( .A(n4197), .B(n4196), .Z(n5641) );
  XNOR U8155 ( .A(n5642), .B(n5641), .Z(n5643) );
  XNOR U8156 ( .A(n5644), .B(n5643), .Z(n6527) );
  NANDN U8157 ( .A(n4199), .B(n4198), .Z(n4203) );
  NANDN U8158 ( .A(n4201), .B(n4200), .Z(n4202) );
  AND U8159 ( .A(n4203), .B(n4202), .Z(n7326) );
  NANDN U8160 ( .A(n4205), .B(n4204), .Z(n4209) );
  NANDN U8161 ( .A(n4207), .B(n4206), .Z(n4208) );
  AND U8162 ( .A(n4209), .B(n4208), .Z(n7325) );
  XOR U8163 ( .A(n7326), .B(n7325), .Z(n7328) );
  NANDN U8164 ( .A(n4211), .B(n4210), .Z(n4215) );
  NANDN U8165 ( .A(n4213), .B(n4212), .Z(n4214) );
  AND U8166 ( .A(n4215), .B(n4214), .Z(n7327) );
  XOR U8167 ( .A(n7328), .B(n7327), .Z(n6196) );
  NANDN U8168 ( .A(n4221), .B(n4220), .Z(n4225) );
  NANDN U8169 ( .A(n4223), .B(n4222), .Z(n4224) );
  AND U8170 ( .A(n4225), .B(n4224), .Z(n5750) );
  XOR U8171 ( .A(n5751), .B(n5750), .Z(n5753) );
  NANDN U8172 ( .A(n4227), .B(n4226), .Z(n4231) );
  NANDN U8173 ( .A(n4229), .B(n4228), .Z(n4230) );
  AND U8174 ( .A(n4231), .B(n4230), .Z(n5752) );
  XOR U8175 ( .A(n5753), .B(n5752), .Z(n6194) );
  XNOR U8176 ( .A(n6194), .B(n6193), .Z(n6195) );
  XOR U8177 ( .A(n6196), .B(n6195), .Z(n6528) );
  XNOR U8178 ( .A(n6527), .B(n6528), .Z(n6529) );
  NANDN U8179 ( .A(n4237), .B(n4236), .Z(n4241) );
  NANDN U8180 ( .A(n4239), .B(n4238), .Z(n4240) );
  AND U8181 ( .A(n4241), .B(n4240), .Z(n5744) );
  NANDN U8182 ( .A(n4243), .B(n4242), .Z(n4247) );
  NAND U8183 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U8184 ( .A(n4247), .B(n4246), .Z(n5743) );
  XOR U8185 ( .A(n5744), .B(n5743), .Z(n5747) );
  NANDN U8186 ( .A(n4249), .B(n4248), .Z(n4253) );
  NAND U8187 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U8188 ( .A(n4253), .B(n4252), .Z(n5746) );
  XOR U8189 ( .A(n5747), .B(n5746), .Z(n6172) );
  NANDN U8190 ( .A(n4255), .B(n4254), .Z(n4259) );
  NANDN U8191 ( .A(n4257), .B(n4256), .Z(n4258) );
  AND U8192 ( .A(n4259), .B(n4258), .Z(n5773) );
  XOR U8193 ( .A(n5773), .B(n5772), .Z(n5775) );
  XOR U8194 ( .A(n5775), .B(n5774), .Z(n6170) );
  NANDN U8195 ( .A(n4269), .B(n4268), .Z(n4273) );
  NANDN U8196 ( .A(n4271), .B(n4270), .Z(n4272) );
  AND U8197 ( .A(n4273), .B(n4272), .Z(n7330) );
  NANDN U8198 ( .A(n4275), .B(n4274), .Z(n4279) );
  NANDN U8199 ( .A(n4277), .B(n4276), .Z(n4278) );
  AND U8200 ( .A(n4279), .B(n4278), .Z(n7329) );
  XOR U8201 ( .A(n7330), .B(n7329), .Z(n7332) );
  NANDN U8202 ( .A(n4281), .B(n4280), .Z(n4285) );
  NANDN U8203 ( .A(n4283), .B(n4282), .Z(n4284) );
  AND U8204 ( .A(n4285), .B(n4284), .Z(n7331) );
  XNOR U8205 ( .A(n7332), .B(n7331), .Z(n6169) );
  XNOR U8206 ( .A(n6170), .B(n6169), .Z(n6171) );
  XOR U8207 ( .A(n6172), .B(n6171), .Z(n6530) );
  XOR U8208 ( .A(n6529), .B(n6530), .Z(n5427) );
  XNOR U8209 ( .A(n5426), .B(n5427), .Z(n5429) );
  NANDN U8210 ( .A(n4287), .B(n4286), .Z(n4291) );
  NAND U8211 ( .A(n4289), .B(n4288), .Z(n4290) );
  AND U8212 ( .A(n4291), .B(n4290), .Z(n5801) );
  XOR U8213 ( .A(n5801), .B(n5800), .Z(n5803) );
  XOR U8214 ( .A(n5803), .B(n5802), .Z(n6166) );
  XOR U8215 ( .A(n5561), .B(n5560), .Z(n5563) );
  XOR U8216 ( .A(n5563), .B(n5562), .Z(n6164) );
  NAND U8217 ( .A(n4313), .B(n4312), .Z(n4317) );
  NAND U8218 ( .A(n4315), .B(n4314), .Z(n4316) );
  AND U8219 ( .A(n4317), .B(n4316), .Z(n6414) );
  NANDN U8220 ( .A(n4319), .B(n4318), .Z(n4323) );
  NANDN U8221 ( .A(n4321), .B(n4320), .Z(n4322) );
  AND U8222 ( .A(n4323), .B(n4322), .Z(n6413) );
  XOR U8223 ( .A(n6414), .B(n6413), .Z(n6416) );
  NANDN U8224 ( .A(n4325), .B(n4324), .Z(n4329) );
  NANDN U8225 ( .A(n4327), .B(n4326), .Z(n4328) );
  AND U8226 ( .A(n4329), .B(n4328), .Z(n6415) );
  XNOR U8227 ( .A(n6416), .B(n6415), .Z(n6163) );
  XNOR U8228 ( .A(n6164), .B(n6163), .Z(n6165) );
  XNOR U8229 ( .A(n6166), .B(n6165), .Z(n6521) );
  NANDN U8230 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U8231 ( .A(n4333), .B(n4332), .Z(n4334) );
  AND U8232 ( .A(n4335), .B(n4334), .Z(n5581) );
  XOR U8233 ( .A(n5581), .B(n5580), .Z(n5583) );
  XOR U8234 ( .A(n5583), .B(n5582), .Z(n6142) );
  NANDN U8235 ( .A(n4345), .B(n4344), .Z(n4349) );
  NAND U8236 ( .A(n4347), .B(n4346), .Z(n4348) );
  AND U8237 ( .A(n4349), .B(n4348), .Z(n5622) );
  XOR U8238 ( .A(n5622), .B(n5621), .Z(n5624) );
  XOR U8239 ( .A(n5624), .B(n5623), .Z(n6140) );
  NANDN U8240 ( .A(n4359), .B(n4358), .Z(n4363) );
  NANDN U8241 ( .A(n4361), .B(n4360), .Z(n4362) );
  AND U8242 ( .A(n4363), .B(n4362), .Z(n5899) );
  XOR U8243 ( .A(n5899), .B(n5898), .Z(n5901) );
  NANDN U8244 ( .A(n4369), .B(n4368), .Z(n4373) );
  NAND U8245 ( .A(n4371), .B(n4370), .Z(n4372) );
  AND U8246 ( .A(n4373), .B(n4372), .Z(n5900) );
  XNOR U8247 ( .A(n5901), .B(n5900), .Z(n6139) );
  XNOR U8248 ( .A(n6140), .B(n6139), .Z(n6141) );
  XOR U8249 ( .A(n6142), .B(n6141), .Z(n6522) );
  XNOR U8250 ( .A(n6521), .B(n6522), .Z(n6523) );
  NANDN U8251 ( .A(n4375), .B(n4374), .Z(n4379) );
  NANDN U8252 ( .A(n4377), .B(n4376), .Z(n4378) );
  AND U8253 ( .A(n4379), .B(n4378), .Z(n5638) );
  NANDN U8254 ( .A(n4381), .B(n4380), .Z(n4385) );
  NANDN U8255 ( .A(n4383), .B(n4382), .Z(n4384) );
  AND U8256 ( .A(n4385), .B(n4384), .Z(n5637) );
  XOR U8257 ( .A(n5638), .B(n5637), .Z(n5640) );
  NANDN U8258 ( .A(n4387), .B(n4386), .Z(n4391) );
  NANDN U8259 ( .A(n4389), .B(n4388), .Z(n4390) );
  AND U8260 ( .A(n4391), .B(n4390), .Z(n5639) );
  XOR U8261 ( .A(n5640), .B(n5639), .Z(n5650) );
  NANDN U8262 ( .A(n4393), .B(n4392), .Z(n4397) );
  NANDN U8263 ( .A(n4395), .B(n4394), .Z(n4396) );
  AND U8264 ( .A(n4397), .B(n4396), .Z(n5470) );
  NANDN U8265 ( .A(n4399), .B(n4398), .Z(n4403) );
  NANDN U8266 ( .A(n4401), .B(n4400), .Z(n4402) );
  NAND U8267 ( .A(n4403), .B(n4402), .Z(n5471) );
  XNOR U8268 ( .A(n5470), .B(n5471), .Z(n5473) );
  NANDN U8269 ( .A(n4405), .B(n4404), .Z(n4409) );
  NANDN U8270 ( .A(n4407), .B(n4406), .Z(n4408) );
  AND U8271 ( .A(n4409), .B(n4408), .Z(n5472) );
  XOR U8272 ( .A(n5473), .B(n5472), .Z(n5648) );
  NANDN U8273 ( .A(n4411), .B(n4410), .Z(n4415) );
  NANDN U8274 ( .A(n4413), .B(n4412), .Z(n4414) );
  AND U8275 ( .A(n4415), .B(n4414), .Z(n5889) );
  XOR U8276 ( .A(n5889), .B(n5888), .Z(n5891) );
  XNOR U8277 ( .A(n5891), .B(n5890), .Z(n5647) );
  XNOR U8278 ( .A(n5648), .B(n5647), .Z(n5649) );
  XOR U8279 ( .A(n5650), .B(n5649), .Z(n6524) );
  XNOR U8280 ( .A(n6523), .B(n6524), .Z(n5428) );
  XOR U8281 ( .A(n5429), .B(n5428), .Z(n7028) );
  NANDN U8282 ( .A(n4425), .B(n4424), .Z(n4429) );
  OR U8283 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U8284 ( .A(n4429), .B(n4428), .Z(n6535) );
  NANDN U8285 ( .A(n4431), .B(n4430), .Z(n4435) );
  OR U8286 ( .A(n4433), .B(n4432), .Z(n4434) );
  AND U8287 ( .A(n4435), .B(n4434), .Z(n6534) );
  NANDN U8288 ( .A(n4437), .B(n4436), .Z(n4441) );
  NANDN U8289 ( .A(n4439), .B(n4438), .Z(n4440) );
  AND U8290 ( .A(n4441), .B(n4440), .Z(n5862) );
  NANDN U8291 ( .A(n4447), .B(n4446), .Z(n4451) );
  NANDN U8292 ( .A(n4449), .B(n4448), .Z(n4450) );
  AND U8293 ( .A(n4451), .B(n4450), .Z(n5864) );
  XOR U8294 ( .A(n5865), .B(n5864), .Z(n6783) );
  NANDN U8295 ( .A(n4453), .B(n4452), .Z(n4457) );
  NANDN U8296 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U8297 ( .A(n4457), .B(n4456), .Z(n7247) );
  NANDN U8298 ( .A(n4459), .B(n4458), .Z(n4463) );
  NANDN U8299 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U8300 ( .A(n4463), .B(n4462), .Z(n7248) );
  XNOR U8301 ( .A(n7247), .B(n7248), .Z(n7250) );
  NANDN U8302 ( .A(n4465), .B(n4464), .Z(n4469) );
  NANDN U8303 ( .A(n4467), .B(n4466), .Z(n4468) );
  AND U8304 ( .A(n4469), .B(n4468), .Z(n7249) );
  XOR U8305 ( .A(n7250), .B(n7249), .Z(n6782) );
  NANDN U8306 ( .A(n4471), .B(n4470), .Z(n4475) );
  NAND U8307 ( .A(n4473), .B(n4472), .Z(n4474) );
  NAND U8308 ( .A(n4475), .B(n4474), .Z(n6781) );
  XOR U8309 ( .A(n6782), .B(n6781), .Z(n6784) );
  XNOR U8310 ( .A(n6783), .B(n6784), .Z(n6533) );
  XOR U8311 ( .A(n6534), .B(n6533), .Z(n6536) );
  XOR U8312 ( .A(n6535), .B(n6536), .Z(n5812) );
  NANDN U8313 ( .A(n4477), .B(n4476), .Z(n4481) );
  OR U8314 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U8315 ( .A(n4481), .B(n4480), .Z(n6579) );
  NANDN U8316 ( .A(n4483), .B(n4482), .Z(n4487) );
  NANDN U8317 ( .A(n4485), .B(n4484), .Z(n4486) );
  AND U8318 ( .A(n4487), .B(n4486), .Z(n5518) );
  NANDN U8319 ( .A(n4489), .B(n4488), .Z(n4493) );
  NANDN U8320 ( .A(n4491), .B(n4490), .Z(n4492) );
  NAND U8321 ( .A(n4493), .B(n4492), .Z(n5519) );
  XNOR U8322 ( .A(n5518), .B(n5519), .Z(n5521) );
  NANDN U8323 ( .A(n4495), .B(n4494), .Z(n4499) );
  NANDN U8324 ( .A(n4497), .B(n4496), .Z(n4498) );
  AND U8325 ( .A(n4499), .B(n4498), .Z(n5520) );
  XOR U8326 ( .A(n5521), .B(n5520), .Z(n6759) );
  NANDN U8327 ( .A(n4501), .B(n4500), .Z(n4505) );
  NANDN U8328 ( .A(n4503), .B(n4502), .Z(n4504) );
  AND U8329 ( .A(n4505), .B(n4504), .Z(n6714) );
  XOR U8330 ( .A(n6714), .B(n6713), .Z(n6716) );
  XOR U8331 ( .A(n6716), .B(n6715), .Z(n6758) );
  NANDN U8332 ( .A(n4515), .B(n4514), .Z(n4519) );
  NAND U8333 ( .A(n4517), .B(n4516), .Z(n4518) );
  NAND U8334 ( .A(n4519), .B(n4518), .Z(n6757) );
  XOR U8335 ( .A(n6758), .B(n6757), .Z(n6760) );
  XOR U8336 ( .A(n6759), .B(n6760), .Z(n6578) );
  NANDN U8337 ( .A(n4521), .B(n4520), .Z(n4525) );
  OR U8338 ( .A(n4523), .B(n4522), .Z(n4524) );
  NAND U8339 ( .A(n4525), .B(n4524), .Z(n6577) );
  XOR U8340 ( .A(n6578), .B(n6577), .Z(n6580) );
  XOR U8341 ( .A(n6579), .B(n6580), .Z(n5811) );
  NANDN U8342 ( .A(n4527), .B(n4526), .Z(n4531) );
  NAND U8343 ( .A(n4529), .B(n4528), .Z(n4530) );
  AND U8344 ( .A(n4531), .B(n4530), .Z(n7400) );
  NANDN U8345 ( .A(n4533), .B(n4532), .Z(n4537) );
  NAND U8346 ( .A(n4535), .B(n4534), .Z(n4536) );
  AND U8347 ( .A(n4537), .B(n4536), .Z(n7398) );
  NANDN U8348 ( .A(n4539), .B(n4538), .Z(n4543) );
  NAND U8349 ( .A(n4541), .B(n4540), .Z(n4542) );
  NAND U8350 ( .A(n4543), .B(n4542), .Z(n7397) );
  XNOR U8351 ( .A(n7398), .B(n7397), .Z(n7399) );
  XNOR U8352 ( .A(n7400), .B(n7399), .Z(n7219) );
  NANDN U8353 ( .A(n4545), .B(n4544), .Z(n4549) );
  NAND U8354 ( .A(n4547), .B(n4546), .Z(n4548) );
  AND U8355 ( .A(n4549), .B(n4548), .Z(n7180) );
  XNOR U8356 ( .A(n7178), .B(n7177), .Z(n7179) );
  XNOR U8357 ( .A(n7180), .B(n7179), .Z(n7217) );
  XNOR U8358 ( .A(n7166), .B(n7165), .Z(n7167) );
  XOR U8359 ( .A(n7168), .B(n7167), .Z(n7218) );
  XOR U8360 ( .A(n7217), .B(n7218), .Z(n7220) );
  XNOR U8361 ( .A(n7219), .B(n7220), .Z(n5810) );
  XOR U8362 ( .A(n5811), .B(n5810), .Z(n5813) );
  XNOR U8363 ( .A(n5812), .B(n5813), .Z(n7027) );
  NANDN U8364 ( .A(n4571), .B(n4570), .Z(n4575) );
  NANDN U8365 ( .A(n4573), .B(n4572), .Z(n4574) );
  AND U8366 ( .A(n4575), .B(n4574), .Z(n6980) );
  NANDN U8367 ( .A(n4577), .B(n4576), .Z(n4581) );
  NANDN U8368 ( .A(n4579), .B(n4578), .Z(n4580) );
  AND U8369 ( .A(n4581), .B(n4580), .Z(n6977) );
  NANDN U8370 ( .A(n4583), .B(n4582), .Z(n4587) );
  NANDN U8371 ( .A(n4585), .B(n4584), .Z(n4586) );
  AND U8372 ( .A(n4587), .B(n4586), .Z(n5494) );
  NANDN U8373 ( .A(n4589), .B(n4588), .Z(n4593) );
  NANDN U8374 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U8375 ( .A(n4593), .B(n4592), .Z(n5495) );
  XNOR U8376 ( .A(n5494), .B(n5495), .Z(n5497) );
  NANDN U8377 ( .A(n4595), .B(n4594), .Z(n4599) );
  NANDN U8378 ( .A(n4597), .B(n4596), .Z(n4598) );
  AND U8379 ( .A(n4599), .B(n4598), .Z(n5496) );
  XOR U8380 ( .A(n5497), .B(n5496), .Z(n5674) );
  NANDN U8381 ( .A(n4601), .B(n4600), .Z(n4605) );
  NANDN U8382 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U8383 ( .A(n4605), .B(n4604), .Z(n7140) );
  NANDN U8384 ( .A(n4607), .B(n4606), .Z(n4611) );
  NANDN U8385 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U8386 ( .A(n4611), .B(n4610), .Z(n7139) );
  XOR U8387 ( .A(n7140), .B(n7139), .Z(n7142) );
  NANDN U8388 ( .A(n4613), .B(n4612), .Z(n4617) );
  NANDN U8389 ( .A(n4615), .B(n4614), .Z(n4616) );
  AND U8390 ( .A(n4617), .B(n4616), .Z(n7141) );
  XOR U8391 ( .A(n7142), .B(n7141), .Z(n5672) );
  NANDN U8392 ( .A(n4619), .B(n4618), .Z(n4623) );
  NAND U8393 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U8394 ( .A(n4623), .B(n4622), .Z(n5671) );
  XNOR U8395 ( .A(n5672), .B(n5671), .Z(n5673) );
  XOR U8396 ( .A(n5674), .B(n5673), .Z(n6978) );
  XNOR U8397 ( .A(n6977), .B(n6978), .Z(n6979) );
  XOR U8398 ( .A(n6980), .B(n6979), .Z(n5410) );
  NANDN U8399 ( .A(n4625), .B(n4624), .Z(n4629) );
  NANDN U8400 ( .A(n4627), .B(n4626), .Z(n4628) );
  AND U8401 ( .A(n4629), .B(n4628), .Z(n6986) );
  NANDN U8402 ( .A(n4631), .B(n4630), .Z(n4635) );
  NANDN U8403 ( .A(n4633), .B(n4632), .Z(n4634) );
  AND U8404 ( .A(n4635), .B(n4634), .Z(n6983) );
  NANDN U8405 ( .A(n4637), .B(n4636), .Z(n4641) );
  NAND U8406 ( .A(n4639), .B(n4638), .Z(n4640) );
  AND U8407 ( .A(n4641), .B(n4640), .Z(n7394) );
  NANDN U8408 ( .A(n4643), .B(n4642), .Z(n4647) );
  NANDN U8409 ( .A(n4645), .B(n4644), .Z(n4646) );
  AND U8410 ( .A(n4647), .B(n4646), .Z(n6036) );
  NANDN U8411 ( .A(n4649), .B(n4648), .Z(n4653) );
  NANDN U8412 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U8413 ( .A(n4653), .B(n4652), .Z(n6037) );
  XNOR U8414 ( .A(n6036), .B(n6037), .Z(n6039) );
  NANDN U8415 ( .A(n4655), .B(n4654), .Z(n4659) );
  NANDN U8416 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U8417 ( .A(n4659), .B(n4658), .Z(n6038) );
  XOR U8418 ( .A(n6039), .B(n6038), .Z(n7392) );
  NANDN U8419 ( .A(n4661), .B(n4660), .Z(n4665) );
  NAND U8420 ( .A(n4663), .B(n4662), .Z(n4664) );
  NAND U8421 ( .A(n4665), .B(n4664), .Z(n7391) );
  XNOR U8422 ( .A(n7392), .B(n7391), .Z(n7393) );
  XOR U8423 ( .A(n7394), .B(n7393), .Z(n6984) );
  XNOR U8424 ( .A(n6983), .B(n6984), .Z(n6985) );
  XOR U8425 ( .A(n6986), .B(n6985), .Z(n5409) );
  NANDN U8426 ( .A(n4667), .B(n4666), .Z(n4671) );
  OR U8427 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U8428 ( .A(n4671), .B(n4670), .Z(n6926) );
  NANDN U8429 ( .A(n4685), .B(n4684), .Z(n4689) );
  NANDN U8430 ( .A(n4687), .B(n4686), .Z(n4688) );
  NAND U8431 ( .A(n4689), .B(n4688), .Z(n6628) );
  XNOR U8432 ( .A(n6627), .B(n6628), .Z(n6630) );
  NANDN U8433 ( .A(n4691), .B(n4690), .Z(n4695) );
  NANDN U8434 ( .A(n4693), .B(n4692), .Z(n4694) );
  AND U8435 ( .A(n4695), .B(n4694), .Z(n6629) );
  XOR U8436 ( .A(n6630), .B(n6629), .Z(n7172) );
  XOR U8437 ( .A(n7172), .B(n7171), .Z(n7174) );
  XNOR U8438 ( .A(n7173), .B(n7174), .Z(n6923) );
  XNOR U8439 ( .A(n6924), .B(n6923), .Z(n6925) );
  XNOR U8440 ( .A(n6926), .B(n6925), .Z(n5408) );
  XOR U8441 ( .A(n5409), .B(n5408), .Z(n5411) );
  XOR U8442 ( .A(n5410), .B(n5411), .Z(n6872) );
  NANDN U8443 ( .A(n4701), .B(n4700), .Z(n4705) );
  NANDN U8444 ( .A(n4703), .B(n4702), .Z(n4704) );
  AND U8445 ( .A(n4705), .B(n4704), .Z(n7110) );
  OR U8446 ( .A(n4707), .B(n4706), .Z(n4711) );
  NANDN U8447 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U8448 ( .A(n4711), .B(n4710), .Z(n6382) );
  NANDN U8449 ( .A(n4713), .B(n4712), .Z(n4717) );
  NANDN U8450 ( .A(n4715), .B(n4714), .Z(n4716) );
  AND U8451 ( .A(n4717), .B(n4716), .Z(n5443) );
  NANDN U8452 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U8453 ( .A(n4721), .B(n4720), .Z(n4722) );
  AND U8454 ( .A(n4723), .B(n4722), .Z(n5442) );
  XOR U8455 ( .A(n5443), .B(n5442), .Z(n5445) );
  XOR U8456 ( .A(n5445), .B(n5444), .Z(n6262) );
  NANDN U8457 ( .A(n4733), .B(n4732), .Z(n4737) );
  NANDN U8458 ( .A(n4735), .B(n4734), .Z(n4736) );
  AND U8459 ( .A(n4737), .B(n4736), .Z(n5438) );
  XOR U8460 ( .A(n5439), .B(n5438), .Z(n5441) );
  NANDN U8461 ( .A(n4739), .B(n4738), .Z(n4743) );
  NANDN U8462 ( .A(n4741), .B(n4740), .Z(n4742) );
  AND U8463 ( .A(n4743), .B(n4742), .Z(n5440) );
  XOR U8464 ( .A(n5441), .B(n5440), .Z(n6260) );
  NANDN U8465 ( .A(n4745), .B(n4744), .Z(n4749) );
  NANDN U8466 ( .A(n4747), .B(n4746), .Z(n4748) );
  AND U8467 ( .A(n4749), .B(n4748), .Z(n7292) );
  NANDN U8468 ( .A(n4751), .B(n4750), .Z(n4755) );
  NANDN U8469 ( .A(n4753), .B(n4752), .Z(n4754) );
  AND U8470 ( .A(n4755), .B(n4754), .Z(n7291) );
  XOR U8471 ( .A(n7292), .B(n7291), .Z(n7294) );
  XNOR U8472 ( .A(n7294), .B(n7293), .Z(n6259) );
  XNOR U8473 ( .A(n6260), .B(n6259), .Z(n6261) );
  XNOR U8474 ( .A(n6262), .B(n6261), .Z(n6381) );
  XOR U8475 ( .A(n6382), .B(n6381), .Z(n6383) );
  XOR U8476 ( .A(n6668), .B(n6667), .Z(n6670) );
  XOR U8477 ( .A(n6670), .B(n6669), .Z(n6102) );
  XOR U8478 ( .A(n6654), .B(n6653), .Z(n6656) );
  XOR U8479 ( .A(n6656), .B(n6655), .Z(n6100) );
  XNOR U8480 ( .A(n6100), .B(n6099), .Z(n6101) );
  XOR U8481 ( .A(n6102), .B(n6101), .Z(n6384) );
  XNOR U8482 ( .A(n6383), .B(n6384), .Z(n7107) );
  XNOR U8483 ( .A(n6117), .B(n6118), .Z(n6120) );
  NANDN U8484 ( .A(n4797), .B(n4796), .Z(n4801) );
  NANDN U8485 ( .A(n4799), .B(n4798), .Z(n4800) );
  AND U8486 ( .A(n4801), .B(n4800), .Z(n6119) );
  XOR U8487 ( .A(n6120), .B(n6119), .Z(n6704) );
  NANDN U8488 ( .A(n4807), .B(n4806), .Z(n4811) );
  NAND U8489 ( .A(n4809), .B(n4808), .Z(n4810) );
  NAND U8490 ( .A(n4811), .B(n4810), .Z(n6701) );
  XNOR U8491 ( .A(n6702), .B(n6701), .Z(n6703) );
  XNOR U8492 ( .A(n6704), .B(n6703), .Z(n6365) );
  XNOR U8493 ( .A(n6900), .B(n6899), .Z(n6901) );
  XNOR U8494 ( .A(n6902), .B(n6901), .Z(n6363) );
  NANDN U8495 ( .A(n4829), .B(n4828), .Z(n4833) );
  NANDN U8496 ( .A(n4831), .B(n4830), .Z(n4832) );
  AND U8497 ( .A(n4833), .B(n4832), .Z(n6009) );
  NANDN U8498 ( .A(n4835), .B(n4834), .Z(n4839) );
  NANDN U8499 ( .A(n4837), .B(n4836), .Z(n4838) );
  AND U8500 ( .A(n4839), .B(n4838), .Z(n6008) );
  XOR U8501 ( .A(n6009), .B(n6008), .Z(n6011) );
  NANDN U8502 ( .A(n4841), .B(n4840), .Z(n4845) );
  NANDN U8503 ( .A(n4843), .B(n4842), .Z(n4844) );
  AND U8504 ( .A(n4845), .B(n4844), .Z(n6010) );
  XOR U8505 ( .A(n6011), .B(n6010), .Z(n6296) );
  XNOR U8506 ( .A(n6296), .B(n6295), .Z(n6297) );
  XOR U8507 ( .A(n6298), .B(n6297), .Z(n6364) );
  XOR U8508 ( .A(n6363), .B(n6364), .Z(n6366) );
  XOR U8509 ( .A(n6365), .B(n6366), .Z(n7108) );
  XNOR U8510 ( .A(n7107), .B(n7108), .Z(n7109) );
  XNOR U8511 ( .A(n7110), .B(n7109), .Z(n6871) );
  XNOR U8512 ( .A(n6872), .B(n6871), .Z(n6874) );
  NANDN U8513 ( .A(n4851), .B(n4850), .Z(n4855) );
  NAND U8514 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U8515 ( .A(n4855), .B(n4854), .Z(n6391) );
  NANDN U8516 ( .A(n4857), .B(n4856), .Z(n4861) );
  NANDN U8517 ( .A(n4859), .B(n4858), .Z(n4860) );
  AND U8518 ( .A(n4861), .B(n4860), .Z(n5875) );
  NANDN U8519 ( .A(n4863), .B(n4862), .Z(n4867) );
  NANDN U8520 ( .A(n4865), .B(n4864), .Z(n4866) );
  AND U8521 ( .A(n4867), .B(n4866), .Z(n5874) );
  XOR U8522 ( .A(n5875), .B(n5874), .Z(n5877) );
  NANDN U8523 ( .A(n4869), .B(n4868), .Z(n4873) );
  NANDN U8524 ( .A(n4871), .B(n4870), .Z(n4872) );
  AND U8525 ( .A(n4873), .B(n4872), .Z(n5876) );
  XOR U8526 ( .A(n5877), .B(n5876), .Z(n6390) );
  NANDN U8527 ( .A(n4875), .B(n4874), .Z(n4879) );
  NAND U8528 ( .A(n4877), .B(n4876), .Z(n4878) );
  NAND U8529 ( .A(n4879), .B(n4878), .Z(n6389) );
  XNOR U8530 ( .A(n6390), .B(n6389), .Z(n6392) );
  XOR U8531 ( .A(n6391), .B(n6392), .Z(n6096) );
  NANDN U8532 ( .A(n4881), .B(n4880), .Z(n4885) );
  NANDN U8533 ( .A(n4883), .B(n4882), .Z(n4884) );
  AND U8534 ( .A(n4885), .B(n4884), .Z(n6807) );
  NANDN U8535 ( .A(n4887), .B(n4886), .Z(n4891) );
  NANDN U8536 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U8537 ( .A(n4891), .B(n4890), .Z(n6808) );
  XNOR U8538 ( .A(n6807), .B(n6808), .Z(n6809) );
  NANDN U8539 ( .A(n4893), .B(n4892), .Z(n4897) );
  NANDN U8540 ( .A(n4895), .B(n4894), .Z(n4896) );
  NAND U8541 ( .A(n4897), .B(n4896), .Z(n6810) );
  XOR U8542 ( .A(n6809), .B(n6810), .Z(n5946) );
  NANDN U8543 ( .A(n4903), .B(n4902), .Z(n4907) );
  NAND U8544 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U8545 ( .A(n4907), .B(n4906), .Z(n5945) );
  XOR U8546 ( .A(n5944), .B(n5945), .Z(n5947) );
  XOR U8547 ( .A(n5946), .B(n5947), .Z(n6095) );
  XOR U8548 ( .A(n6096), .B(n6095), .Z(n6097) );
  NAND U8549 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U8550 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U8551 ( .A(n4913), .B(n4912), .Z(n6076) );
  NAND U8552 ( .A(n4915), .B(n4914), .Z(n4919) );
  NAND U8553 ( .A(n4917), .B(n4916), .Z(n4918) );
  AND U8554 ( .A(n4919), .B(n4918), .Z(n6075) );
  XOR U8555 ( .A(n6076), .B(n6075), .Z(n6078) );
  NAND U8556 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U8557 ( .A(n4923), .B(n4922), .Z(n4924) );
  AND U8558 ( .A(n4925), .B(n4924), .Z(n6077) );
  XOR U8559 ( .A(n6078), .B(n6077), .Z(n6754) );
  XOR U8560 ( .A(n6053), .B(n6052), .Z(n6055) );
  NANDN U8561 ( .A(n4935), .B(n4934), .Z(n4939) );
  NANDN U8562 ( .A(n4937), .B(n4936), .Z(n4938) );
  AND U8563 ( .A(n4939), .B(n4938), .Z(n6054) );
  XOR U8564 ( .A(n6055), .B(n6054), .Z(n6752) );
  XNOR U8565 ( .A(n6752), .B(n6751), .Z(n6753) );
  XOR U8566 ( .A(n6754), .B(n6753), .Z(n6098) );
  XNOR U8567 ( .A(n6097), .B(n6098), .Z(n6995) );
  XNOR U8568 ( .A(n5537), .B(n5536), .Z(n5538) );
  XNOR U8569 ( .A(n5539), .B(n5538), .Z(n5826) );
  NANDN U8570 ( .A(n4957), .B(n4956), .Z(n4961) );
  NAND U8571 ( .A(n4959), .B(n4958), .Z(n4960) );
  AND U8572 ( .A(n4961), .B(n4960), .Z(n6816) );
  NANDN U8573 ( .A(n4963), .B(n4962), .Z(n4967) );
  NANDN U8574 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U8575 ( .A(n4967), .B(n4966), .Z(n6740) );
  NANDN U8576 ( .A(n4969), .B(n4968), .Z(n4973) );
  NANDN U8577 ( .A(n4971), .B(n4970), .Z(n4972) );
  AND U8578 ( .A(n4973), .B(n4972), .Z(n6739) );
  XOR U8579 ( .A(n6740), .B(n6739), .Z(n6742) );
  NANDN U8580 ( .A(n4975), .B(n4974), .Z(n4979) );
  NANDN U8581 ( .A(n4977), .B(n4976), .Z(n4978) );
  AND U8582 ( .A(n4979), .B(n4978), .Z(n6741) );
  XOR U8583 ( .A(n6742), .B(n6741), .Z(n6814) );
  NANDN U8584 ( .A(n4981), .B(n4980), .Z(n4985) );
  NAND U8585 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U8586 ( .A(n4985), .B(n4984), .Z(n6813) );
  XNOR U8587 ( .A(n6814), .B(n6813), .Z(n6815) );
  XOR U8588 ( .A(n6816), .B(n6815), .Z(n5827) );
  XNOR U8589 ( .A(n5826), .B(n5827), .Z(n5828) );
  NANDN U8590 ( .A(n4987), .B(n4986), .Z(n4991) );
  NANDN U8591 ( .A(n4989), .B(n4988), .Z(n4990) );
  AND U8592 ( .A(n4991), .B(n4990), .Z(n6496) );
  NANDN U8593 ( .A(n4993), .B(n4992), .Z(n4997) );
  NANDN U8594 ( .A(n4995), .B(n4994), .Z(n4996) );
  AND U8595 ( .A(n4997), .B(n4996), .Z(n6419) );
  NAND U8596 ( .A(n4999), .B(n4998), .Z(n5003) );
  NAND U8597 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U8598 ( .A(n5003), .B(n5002), .Z(n6420) );
  NAND U8599 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U8600 ( .A(n5007), .B(n5006), .Z(n5008) );
  AND U8601 ( .A(n5009), .B(n5008), .Z(n6421) );
  XOR U8602 ( .A(n6422), .B(n6421), .Z(n6494) );
  NANDN U8603 ( .A(n5011), .B(n5010), .Z(n5015) );
  NAND U8604 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U8605 ( .A(n5015), .B(n5014), .Z(n6493) );
  XNOR U8606 ( .A(n6494), .B(n6493), .Z(n6495) );
  XOR U8607 ( .A(n6496), .B(n6495), .Z(n5829) );
  XOR U8608 ( .A(n5828), .B(n5829), .Z(n6996) );
  XNOR U8609 ( .A(n6995), .B(n6996), .Z(n6998) );
  NANDN U8610 ( .A(n5017), .B(n5016), .Z(n5021) );
  NANDN U8611 ( .A(n5019), .B(n5018), .Z(n5020) );
  AND U8612 ( .A(n5021), .B(n5020), .Z(n6043) );
  NANDN U8613 ( .A(n5023), .B(n5022), .Z(n5027) );
  NANDN U8614 ( .A(n5025), .B(n5024), .Z(n5026) );
  AND U8615 ( .A(n5027), .B(n5026), .Z(n6042) );
  XOR U8616 ( .A(n6043), .B(n6042), .Z(n6045) );
  XOR U8617 ( .A(n6045), .B(n6044), .Z(n6023) );
  NANDN U8618 ( .A(n5033), .B(n5032), .Z(n5037) );
  NANDN U8619 ( .A(n5035), .B(n5034), .Z(n5036) );
  AND U8620 ( .A(n5037), .B(n5036), .Z(n6638) );
  NANDN U8621 ( .A(n5039), .B(n5038), .Z(n5043) );
  NANDN U8622 ( .A(n5041), .B(n5040), .Z(n5042) );
  AND U8623 ( .A(n5043), .B(n5042), .Z(n6637) );
  XOR U8624 ( .A(n6638), .B(n6637), .Z(n6640) );
  NANDN U8625 ( .A(n5045), .B(n5044), .Z(n5049) );
  NANDN U8626 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U8627 ( .A(n5049), .B(n5048), .Z(n6639) );
  XOR U8628 ( .A(n6640), .B(n6639), .Z(n6021) );
  XNOR U8629 ( .A(n6021), .B(n6020), .Z(n6022) );
  XNOR U8630 ( .A(n6023), .B(n6022), .Z(n6520) );
  NANDN U8631 ( .A(n5055), .B(n5054), .Z(n5059) );
  NAND U8632 ( .A(n5057), .B(n5056), .Z(n5058) );
  AND U8633 ( .A(n5059), .B(n5058), .Z(n7132) );
  XNOR U8634 ( .A(n6717), .B(n6718), .Z(n6720) );
  XOR U8635 ( .A(n6720), .B(n6719), .Z(n7130) );
  XNOR U8636 ( .A(n7130), .B(n7129), .Z(n7131) );
  XNOR U8637 ( .A(n7132), .B(n7131), .Z(n6518) );
  NANDN U8638 ( .A(n5077), .B(n5076), .Z(n5081) );
  NAND U8639 ( .A(n5079), .B(n5078), .Z(n5080) );
  AND U8640 ( .A(n5081), .B(n5080), .Z(n6794) );
  NANDN U8641 ( .A(n5083), .B(n5082), .Z(n5087) );
  NANDN U8642 ( .A(n5085), .B(n5084), .Z(n5086) );
  AND U8643 ( .A(n5087), .B(n5086), .Z(n6744) );
  NANDN U8644 ( .A(n5089), .B(n5088), .Z(n5093) );
  NANDN U8645 ( .A(n5091), .B(n5090), .Z(n5092) );
  AND U8646 ( .A(n5093), .B(n5092), .Z(n6743) );
  XOR U8647 ( .A(n6744), .B(n6743), .Z(n6746) );
  NANDN U8648 ( .A(n5095), .B(n5094), .Z(n5099) );
  NANDN U8649 ( .A(n5097), .B(n5096), .Z(n5098) );
  AND U8650 ( .A(n5099), .B(n5098), .Z(n6745) );
  XOR U8651 ( .A(n6746), .B(n6745), .Z(n6792) );
  XNOR U8652 ( .A(n6792), .B(n6791), .Z(n6793) );
  XNOR U8653 ( .A(n6794), .B(n6793), .Z(n6517) );
  XOR U8654 ( .A(n6518), .B(n6517), .Z(n6519) );
  XOR U8655 ( .A(n6520), .B(n6519), .Z(n6997) );
  XOR U8656 ( .A(n6998), .B(n6997), .Z(n6873) );
  XOR U8657 ( .A(n6874), .B(n6873), .Z(n7023) );
  XOR U8658 ( .A(n7024), .B(n7023), .Z(n7026) );
  NANDN U8659 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U8660 ( .A(n5107), .B(n5106), .Z(n5108) );
  AND U8661 ( .A(n5109), .B(n5108), .Z(n7114) );
  NANDN U8662 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U8663 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U8664 ( .A(n5115), .B(n5114), .Z(n7113) );
  XNOR U8665 ( .A(n7114), .B(n7113), .Z(n7116) );
  NANDN U8666 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U8667 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U8668 ( .A(n5121), .B(n5120), .Z(n6943) );
  NANDN U8669 ( .A(n5123), .B(n5122), .Z(n5127) );
  NANDN U8670 ( .A(n5125), .B(n5124), .Z(n5126) );
  AND U8671 ( .A(n5127), .B(n5126), .Z(n6942) );
  NANDN U8672 ( .A(n5129), .B(n5128), .Z(n5133) );
  NANDN U8673 ( .A(n5131), .B(n5130), .Z(n5132) );
  AND U8674 ( .A(n5133), .B(n5132), .Z(n7364) );
  NAND U8675 ( .A(n5135), .B(n5134), .Z(n5139) );
  NAND U8676 ( .A(n5137), .B(n5136), .Z(n5138) );
  NAND U8677 ( .A(n5139), .B(n5138), .Z(n7265) );
  NANDN U8678 ( .A(n5141), .B(n5140), .Z(n5145) );
  NAND U8679 ( .A(n5143), .B(n5142), .Z(n5144) );
  AND U8680 ( .A(n5145), .B(n5144), .Z(n6080) );
  NANDN U8681 ( .A(n5147), .B(n5146), .Z(n5151) );
  NAND U8682 ( .A(n5149), .B(n5148), .Z(n5150) );
  AND U8683 ( .A(n5151), .B(n5150), .Z(n6079) );
  XOR U8684 ( .A(n6080), .B(n6079), .Z(n6082) );
  NANDN U8685 ( .A(n5153), .B(n5152), .Z(n5157) );
  NAND U8686 ( .A(n5155), .B(n5154), .Z(n5156) );
  AND U8687 ( .A(n5157), .B(n5156), .Z(n6081) );
  XOR U8688 ( .A(n6082), .B(n6081), .Z(n7264) );
  NAND U8689 ( .A(n5159), .B(n5158), .Z(n5163) );
  NAND U8690 ( .A(n5161), .B(n5160), .Z(n5162) );
  NAND U8691 ( .A(n5163), .B(n5162), .Z(n7263) );
  XNOR U8692 ( .A(n7264), .B(n7263), .Z(n7266) );
  XOR U8693 ( .A(n7265), .B(n7266), .Z(n7363) );
  XOR U8694 ( .A(n7364), .B(n7363), .Z(n7366) );
  NANDN U8695 ( .A(n5165), .B(n5164), .Z(n5169) );
  NAND U8696 ( .A(n5167), .B(n5166), .Z(n5168) );
  NAND U8697 ( .A(n5169), .B(n5168), .Z(n6907) );
  NANDN U8698 ( .A(n5175), .B(n5174), .Z(n5179) );
  NANDN U8699 ( .A(n5177), .B(n5176), .Z(n5178) );
  NAND U8700 ( .A(n5179), .B(n5178), .Z(n6906) );
  XOR U8701 ( .A(n6905), .B(n6906), .Z(n6908) );
  XOR U8702 ( .A(n6907), .B(n6908), .Z(n7365) );
  XOR U8703 ( .A(n7366), .B(n7365), .Z(n6941) );
  XOR U8704 ( .A(n6942), .B(n6941), .Z(n6944) );
  XNOR U8705 ( .A(n6943), .B(n6944), .Z(n6376) );
  NANDN U8706 ( .A(n5181), .B(n5180), .Z(n5185) );
  NANDN U8707 ( .A(n5183), .B(n5182), .Z(n5184) );
  AND U8708 ( .A(n5185), .B(n5184), .Z(n6973) );
  NANDN U8709 ( .A(n5191), .B(n5190), .Z(n5195) );
  NANDN U8710 ( .A(n5193), .B(n5192), .Z(n5194) );
  AND U8711 ( .A(n5195), .B(n5194), .Z(n7341) );
  NANDN U8712 ( .A(n5197), .B(n5196), .Z(n5201) );
  NANDN U8713 ( .A(n5199), .B(n5198), .Z(n5200) );
  AND U8714 ( .A(n5201), .B(n5200), .Z(n7339) );
  NANDN U8715 ( .A(n5203), .B(n5202), .Z(n5207) );
  NANDN U8716 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U8717 ( .A(n5207), .B(n5206), .Z(n7340) );
  XOR U8718 ( .A(n7339), .B(n7340), .Z(n7342) );
  XOR U8719 ( .A(n7341), .B(n7342), .Z(n6972) );
  XOR U8720 ( .A(n6971), .B(n6972), .Z(n6974) );
  XOR U8721 ( .A(n6973), .B(n6974), .Z(n6375) );
  XOR U8722 ( .A(n6376), .B(n6375), .Z(n6378) );
  NANDN U8723 ( .A(n5209), .B(n5208), .Z(n5213) );
  OR U8724 ( .A(n5211), .B(n5210), .Z(n5212) );
  AND U8725 ( .A(n5213), .B(n5212), .Z(n6967) );
  NANDN U8726 ( .A(n5219), .B(n5218), .Z(n5223) );
  NANDN U8727 ( .A(n5221), .B(n5220), .Z(n5222) );
  AND U8728 ( .A(n5223), .B(n5222), .Z(n5339) );
  XNOR U8729 ( .A(n5868), .B(n5869), .Z(n5870) );
  XOR U8730 ( .A(n5870), .B(n5871), .Z(n6385) );
  NANDN U8731 ( .A(n5241), .B(n5240), .Z(n5245) );
  NAND U8732 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U8733 ( .A(n5245), .B(n5244), .Z(n6386) );
  XOR U8734 ( .A(n6385), .B(n6386), .Z(n6388) );
  XOR U8735 ( .A(n6387), .B(n6388), .Z(n5338) );
  XOR U8736 ( .A(n5339), .B(n5338), .Z(n5341) );
  NANDN U8737 ( .A(n5247), .B(n5246), .Z(n5251) );
  NANDN U8738 ( .A(n5249), .B(n5248), .Z(n5250) );
  AND U8739 ( .A(n5251), .B(n5250), .Z(n5548) );
  NANDN U8740 ( .A(n5253), .B(n5252), .Z(n5257) );
  NANDN U8741 ( .A(n5255), .B(n5254), .Z(n5256) );
  NAND U8742 ( .A(n5257), .B(n5256), .Z(n5549) );
  XNOR U8743 ( .A(n5548), .B(n5549), .Z(n5550) );
  NANDN U8744 ( .A(n5259), .B(n5258), .Z(n5263) );
  NANDN U8745 ( .A(n5261), .B(n5260), .Z(n5262) );
  NAND U8746 ( .A(n5263), .B(n5262), .Z(n5551) );
  XOR U8747 ( .A(n5550), .B(n5551), .Z(n6361) );
  NANDN U8748 ( .A(n5265), .B(n5264), .Z(n5269) );
  NANDN U8749 ( .A(n5267), .B(n5266), .Z(n5268) );
  AND U8750 ( .A(n5269), .B(n5268), .Z(n5554) );
  NANDN U8751 ( .A(n5271), .B(n5270), .Z(n5275) );
  NANDN U8752 ( .A(n5273), .B(n5272), .Z(n5274) );
  NAND U8753 ( .A(n5275), .B(n5274), .Z(n5555) );
  XNOR U8754 ( .A(n5554), .B(n5555), .Z(n5556) );
  NANDN U8755 ( .A(n5277), .B(n5276), .Z(n5281) );
  NANDN U8756 ( .A(n5279), .B(n5278), .Z(n5280) );
  NAND U8757 ( .A(n5281), .B(n5280), .Z(n5557) );
  XOR U8758 ( .A(n5556), .B(n5557), .Z(n6359) );
  XOR U8759 ( .A(n6359), .B(n6360), .Z(n6362) );
  XOR U8760 ( .A(n6361), .B(n6362), .Z(n5340) );
  XOR U8761 ( .A(n5341), .B(n5340), .Z(n6965) );
  XOR U8762 ( .A(n6966), .B(n6965), .Z(n6968) );
  XOR U8763 ( .A(n6967), .B(n6968), .Z(n6377) );
  XOR U8764 ( .A(n6378), .B(n6377), .Z(n7115) );
  XOR U8765 ( .A(n7116), .B(n7115), .Z(n7025) );
  XOR U8766 ( .A(n7026), .B(n7025), .Z(n7445) );
  XNOR U8767 ( .A(n7446), .B(n7445), .Z(n6931) );
  XNOR U8768 ( .A(n6932), .B(n6931), .Z(o[1]) );
  NANDN U8769 ( .A(n5287), .B(n5286), .Z(n5291) );
  NANDN U8770 ( .A(n5289), .B(n5288), .Z(n5290) );
  AND U8771 ( .A(n5291), .B(n5290), .Z(n8366) );
  NANDN U8772 ( .A(n5293), .B(n5292), .Z(n5297) );
  NANDN U8773 ( .A(n5295), .B(n5294), .Z(n5296) );
  AND U8774 ( .A(n5297), .B(n5296), .Z(n8364) );
  NANDN U8775 ( .A(n5299), .B(n5298), .Z(n5303) );
  NANDN U8776 ( .A(n5301), .B(n5300), .Z(n5302) );
  AND U8777 ( .A(n5303), .B(n5302), .Z(n8382) );
  NANDN U8778 ( .A(n5309), .B(n5308), .Z(n5313) );
  NANDN U8779 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U8780 ( .A(n5313), .B(n5312), .Z(n8301) );
  XOR U8781 ( .A(n8302), .B(n8301), .Z(n8304) );
  XOR U8782 ( .A(n8304), .B(n8303), .Z(n8407) );
  NANDN U8783 ( .A(n5319), .B(n5318), .Z(n5323) );
  NAND U8784 ( .A(n5321), .B(n5320), .Z(n5322) );
  AND U8785 ( .A(n5323), .B(n5322), .Z(n8406) );
  NAND U8786 ( .A(n5329), .B(n5328), .Z(n5333) );
  NAND U8787 ( .A(n5331), .B(n5330), .Z(n5332) );
  AND U8788 ( .A(n5333), .B(n5332), .Z(n8291) );
  XOR U8789 ( .A(n8292), .B(n8291), .Z(n8294) );
  XNOR U8790 ( .A(n8294), .B(n8293), .Z(n8405) );
  XOR U8791 ( .A(n8406), .B(n8405), .Z(n8408) );
  XOR U8792 ( .A(n8407), .B(n8408), .Z(n7857) );
  XNOR U8793 ( .A(n8049), .B(n8050), .Z(n8052) );
  XOR U8794 ( .A(n8052), .B(n8051), .Z(n8471) );
  NANDN U8795 ( .A(n5355), .B(n5354), .Z(n5359) );
  NANDN U8796 ( .A(n5357), .B(n5356), .Z(n5358) );
  AND U8797 ( .A(n5359), .B(n5358), .Z(n8074) );
  XOR U8798 ( .A(n8074), .B(n8073), .Z(n8076) );
  XNOR U8799 ( .A(n8076), .B(n8075), .Z(n8470) );
  XOR U8800 ( .A(n8471), .B(n8470), .Z(n8473) );
  XOR U8801 ( .A(n8472), .B(n8473), .Z(n7856) );
  NANDN U8802 ( .A(n5369), .B(n5368), .Z(n5373) );
  NANDN U8803 ( .A(n5371), .B(n5370), .Z(n5372) );
  AND U8804 ( .A(n5373), .B(n5372), .Z(n7939) );
  NANDN U8805 ( .A(n5375), .B(n5374), .Z(n5379) );
  NANDN U8806 ( .A(n5377), .B(n5376), .Z(n5378) );
  AND U8807 ( .A(n5379), .B(n5378), .Z(n8216) );
  NANDN U8808 ( .A(n5381), .B(n5380), .Z(n5385) );
  NANDN U8809 ( .A(n5383), .B(n5382), .Z(n5384) );
  AND U8810 ( .A(n5385), .B(n5384), .Z(n8213) );
  NANDN U8811 ( .A(n5387), .B(n5386), .Z(n5391) );
  NANDN U8812 ( .A(n5389), .B(n5388), .Z(n5390) );
  NAND U8813 ( .A(n5391), .B(n5390), .Z(n8214) );
  XNOR U8814 ( .A(n8213), .B(n8214), .Z(n8215) );
  XOR U8815 ( .A(n8216), .B(n8215), .Z(n7938) );
  NAND U8816 ( .A(n5393), .B(n5392), .Z(n5397) );
  NAND U8817 ( .A(n5395), .B(n5394), .Z(n5396) );
  AND U8818 ( .A(n5397), .B(n5396), .Z(n8016) );
  NAND U8819 ( .A(n5399), .B(n5398), .Z(n5403) );
  NAND U8820 ( .A(n5401), .B(n5400), .Z(n5402) );
  AND U8821 ( .A(n5403), .B(n5402), .Z(n8013) );
  XNOR U8822 ( .A(n8013), .B(n8014), .Z(n8015) );
  XNOR U8823 ( .A(n8016), .B(n8015), .Z(n7937) );
  XOR U8824 ( .A(n7938), .B(n7937), .Z(n7940) );
  XNOR U8825 ( .A(n7939), .B(n7940), .Z(n7855) );
  XOR U8826 ( .A(n7856), .B(n7855), .Z(n7858) );
  XNOR U8827 ( .A(n7857), .B(n7858), .Z(n8381) );
  XNOR U8828 ( .A(n8382), .B(n8381), .Z(n8383) );
  NANDN U8829 ( .A(n5409), .B(n5408), .Z(n5413) );
  OR U8830 ( .A(n5411), .B(n5410), .Z(n5412) );
  AND U8831 ( .A(n5413), .B(n5412), .Z(n8191) );
  NANDN U8832 ( .A(n5415), .B(n5414), .Z(n5419) );
  NANDN U8833 ( .A(n5417), .B(n5416), .Z(n5418) );
  AND U8834 ( .A(n5419), .B(n5418), .Z(n8189) );
  NANDN U8835 ( .A(n5421), .B(n5420), .Z(n5425) );
  NANDN U8836 ( .A(n5423), .B(n5422), .Z(n5424) );
  NAND U8837 ( .A(n5425), .B(n5424), .Z(n8190) );
  XOR U8838 ( .A(n8189), .B(n8190), .Z(n8192) );
  XOR U8839 ( .A(n8191), .B(n8192), .Z(n8384) );
  XNOR U8840 ( .A(n8383), .B(n8384), .Z(n8363) );
  XOR U8841 ( .A(n8364), .B(n8363), .Z(n8365) );
  XOR U8842 ( .A(n8366), .B(n8365), .Z(n7805) );
  NANDN U8843 ( .A(n5427), .B(n5426), .Z(n5431) );
  NAND U8844 ( .A(n5429), .B(n5428), .Z(n5430) );
  NAND U8845 ( .A(n5431), .B(n5430), .Z(n8357) );
  NANDN U8846 ( .A(n5433), .B(n5432), .Z(n5437) );
  NANDN U8847 ( .A(n5435), .B(n5434), .Z(n5436) );
  AND U8848 ( .A(n5437), .B(n5436), .Z(n7827) );
  NANDN U8849 ( .A(n5447), .B(n5446), .Z(n5451) );
  NANDN U8850 ( .A(n5449), .B(n5448), .Z(n5450) );
  NAND U8851 ( .A(n5451), .B(n5450), .Z(n8019) );
  XNOR U8852 ( .A(n8020), .B(n8019), .Z(n8021) );
  XOR U8853 ( .A(n8022), .B(n8021), .Z(n7828) );
  XNOR U8854 ( .A(n7827), .B(n7828), .Z(n7830) );
  NANDN U8855 ( .A(n5453), .B(n5452), .Z(n5457) );
  NANDN U8856 ( .A(n5455), .B(n5454), .Z(n5456) );
  AND U8857 ( .A(n5457), .B(n5456), .Z(n7829) );
  XOR U8858 ( .A(n7830), .B(n7829), .Z(n7840) );
  NANDN U8859 ( .A(n5459), .B(n5458), .Z(n5463) );
  NANDN U8860 ( .A(n5461), .B(n5460), .Z(n5462) );
  NAND U8861 ( .A(n5463), .B(n5462), .Z(n7473) );
  NANDN U8862 ( .A(n5465), .B(n5464), .Z(n5469) );
  NANDN U8863 ( .A(n5467), .B(n5466), .Z(n5468) );
  NAND U8864 ( .A(n5469), .B(n5468), .Z(n7471) );
  NANDN U8865 ( .A(n5471), .B(n5470), .Z(n5475) );
  NAND U8866 ( .A(n5473), .B(n5472), .Z(n5474) );
  NAND U8867 ( .A(n5475), .B(n5474), .Z(n7472) );
  XOR U8868 ( .A(n7471), .B(n7472), .Z(n7474) );
  XOR U8869 ( .A(n7473), .B(n7474), .Z(n8100) );
  NANDN U8870 ( .A(n5477), .B(n5476), .Z(n5481) );
  NAND U8871 ( .A(n5479), .B(n5478), .Z(n5480) );
  NAND U8872 ( .A(n5481), .B(n5480), .Z(n7635) );
  NANDN U8873 ( .A(n5483), .B(n5482), .Z(n5487) );
  NAND U8874 ( .A(n5485), .B(n5484), .Z(n5486) );
  NAND U8875 ( .A(n5487), .B(n5486), .Z(n7633) );
  NANDN U8876 ( .A(n5489), .B(n5488), .Z(n5493) );
  NAND U8877 ( .A(n5491), .B(n5490), .Z(n5492) );
  NAND U8878 ( .A(n5493), .B(n5492), .Z(n7634) );
  XOR U8879 ( .A(n7633), .B(n7634), .Z(n7636) );
  XOR U8880 ( .A(n7635), .B(n7636), .Z(n8099) );
  XOR U8881 ( .A(n8100), .B(n8099), .Z(n8102) );
  NANDN U8882 ( .A(n5495), .B(n5494), .Z(n5499) );
  NAND U8883 ( .A(n5497), .B(n5496), .Z(n5498) );
  NAND U8884 ( .A(n5499), .B(n5498), .Z(n7545) );
  NANDN U8885 ( .A(n5501), .B(n5500), .Z(n5505) );
  NAND U8886 ( .A(n5503), .B(n5502), .Z(n5504) );
  NAND U8887 ( .A(n5505), .B(n5504), .Z(n7543) );
  NANDN U8888 ( .A(n5507), .B(n5506), .Z(n5511) );
  NAND U8889 ( .A(n5509), .B(n5508), .Z(n5510) );
  NAND U8890 ( .A(n5511), .B(n5510), .Z(n7544) );
  XOR U8891 ( .A(n7543), .B(n7544), .Z(n7546) );
  XOR U8892 ( .A(n7545), .B(n7546), .Z(n8101) );
  XOR U8893 ( .A(n8102), .B(n8101), .Z(n7838) );
  NANDN U8894 ( .A(n5513), .B(n5512), .Z(n5517) );
  NANDN U8895 ( .A(n5515), .B(n5514), .Z(n5516) );
  AND U8896 ( .A(n5517), .B(n5516), .Z(n8104) );
  NANDN U8897 ( .A(n5519), .B(n5518), .Z(n5523) );
  NAND U8898 ( .A(n5521), .B(n5520), .Z(n5522) );
  NAND U8899 ( .A(n5523), .B(n5522), .Z(n7469) );
  NANDN U8900 ( .A(n5525), .B(n5524), .Z(n5529) );
  NANDN U8901 ( .A(n5527), .B(n5526), .Z(n5528) );
  NAND U8902 ( .A(n5529), .B(n5528), .Z(n7467) );
  NANDN U8903 ( .A(n5531), .B(n5530), .Z(n5535) );
  NANDN U8904 ( .A(n5533), .B(n5532), .Z(n5534) );
  NAND U8905 ( .A(n5535), .B(n5534), .Z(n7468) );
  XOR U8906 ( .A(n7467), .B(n7468), .Z(n7470) );
  XOR U8907 ( .A(n7469), .B(n7470), .Z(n8103) );
  XOR U8908 ( .A(n8104), .B(n8103), .Z(n8106) );
  NANDN U8909 ( .A(n5537), .B(n5536), .Z(n5541) );
  NANDN U8910 ( .A(n5539), .B(n5538), .Z(n5540) );
  AND U8911 ( .A(n5541), .B(n5540), .Z(n8105) );
  XNOR U8912 ( .A(n8106), .B(n8105), .Z(n7837) );
  XNOR U8913 ( .A(n7838), .B(n7837), .Z(n7839) );
  XNOR U8914 ( .A(n7840), .B(n7839), .Z(n8358) );
  XOR U8915 ( .A(n8357), .B(n8358), .Z(n8360) );
  NANDN U8916 ( .A(n5543), .B(n5542), .Z(n5547) );
  NANDN U8917 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U8918 ( .A(n5547), .B(n5546), .Z(n8327) );
  NANDN U8919 ( .A(n5549), .B(n5548), .Z(n5553) );
  NANDN U8920 ( .A(n5551), .B(n5550), .Z(n5552) );
  NAND U8921 ( .A(n5553), .B(n5552), .Z(n7519) );
  NANDN U8922 ( .A(n5555), .B(n5554), .Z(n5559) );
  NANDN U8923 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U8924 ( .A(n5559), .B(n5558), .Z(n7517) );
  XNOR U8925 ( .A(n7517), .B(n7518), .Z(n7520) );
  XOR U8926 ( .A(n7519), .B(n7520), .Z(n8328) );
  XNOR U8927 ( .A(n8327), .B(n8328), .Z(n8330) );
  NANDN U8928 ( .A(n5565), .B(n5564), .Z(n5569) );
  NANDN U8929 ( .A(n5567), .B(n5566), .Z(n5568) );
  AND U8930 ( .A(n5569), .B(n5568), .Z(n8329) );
  XOR U8931 ( .A(n8330), .B(n8329), .Z(n7820) );
  NANDN U8932 ( .A(n5571), .B(n5570), .Z(n5575) );
  NANDN U8933 ( .A(n5573), .B(n5572), .Z(n5574) );
  AND U8934 ( .A(n5575), .B(n5574), .Z(n8064) );
  IV U8935 ( .A(n7998), .Z(n5588) );
  XOR U8936 ( .A(n5588), .B(n7997), .Z(n8063) );
  XOR U8937 ( .A(n8064), .B(n8063), .Z(n8066) );
  NANDN U8938 ( .A(n5590), .B(n5589), .Z(n5594) );
  NANDN U8939 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U8940 ( .A(n5594), .B(n5593), .Z(n8065) );
  XOR U8941 ( .A(n8066), .B(n8065), .Z(n7818) );
  NANDN U8942 ( .A(n5600), .B(n5599), .Z(n5604) );
  NAND U8943 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U8944 ( .A(n5604), .B(n5603), .Z(n8264) );
  NANDN U8945 ( .A(n5606), .B(n5605), .Z(n5610) );
  NAND U8946 ( .A(n5608), .B(n5607), .Z(n5609) );
  NAND U8947 ( .A(n5610), .B(n5609), .Z(n8263) );
  XNOR U8948 ( .A(n8264), .B(n8263), .Z(n8265) );
  XNOR U8949 ( .A(n8266), .B(n8265), .Z(n7824) );
  NANDN U8950 ( .A(n5612), .B(n5611), .Z(n5616) );
  NANDN U8951 ( .A(n5614), .B(n5613), .Z(n5615) );
  NAND U8952 ( .A(n5616), .B(n5615), .Z(n7515) );
  XOR U8953 ( .A(n7513), .B(n7514), .Z(n7516) );
  XOR U8954 ( .A(n7515), .B(n7516), .Z(n7823) );
  XOR U8955 ( .A(n7824), .B(n7823), .Z(n7826) );
  NANDN U8956 ( .A(n5626), .B(n5625), .Z(n5630) );
  NANDN U8957 ( .A(n5628), .B(n5627), .Z(n5629) );
  AND U8958 ( .A(n5630), .B(n5629), .Z(n7620) );
  NANDN U8959 ( .A(n5632), .B(n5631), .Z(n5636) );
  NANDN U8960 ( .A(n5634), .B(n5633), .Z(n5635) );
  AND U8961 ( .A(n5636), .B(n5635), .Z(n7618) );
  XNOR U8962 ( .A(n7618), .B(n7617), .Z(n7619) );
  XNOR U8963 ( .A(n7620), .B(n7619), .Z(n7825) );
  XNOR U8964 ( .A(n7826), .B(n7825), .Z(n7817) );
  XNOR U8965 ( .A(n7818), .B(n7817), .Z(n7819) );
  XNOR U8966 ( .A(n7820), .B(n7819), .Z(n8359) );
  XOR U8967 ( .A(n8360), .B(n8359), .Z(n7788) );
  NANDN U8968 ( .A(n5642), .B(n5641), .Z(n5646) );
  NANDN U8969 ( .A(n5644), .B(n5643), .Z(n5645) );
  AND U8970 ( .A(n5646), .B(n5645), .Z(n7932) );
  NANDN U8971 ( .A(n5648), .B(n5647), .Z(n5652) );
  NANDN U8972 ( .A(n5650), .B(n5649), .Z(n5651) );
  AND U8973 ( .A(n5652), .B(n5651), .Z(n7930) );
  NANDN U8974 ( .A(n5654), .B(n5653), .Z(n5658) );
  NAND U8975 ( .A(n5656), .B(n5655), .Z(n5657) );
  AND U8976 ( .A(n5658), .B(n5657), .Z(n8227) );
  NANDN U8977 ( .A(n5660), .B(n5659), .Z(n5664) );
  NAND U8978 ( .A(n5662), .B(n5661), .Z(n5663) );
  AND U8979 ( .A(n5664), .B(n5663), .Z(n8226) );
  NANDN U8980 ( .A(n5666), .B(n5665), .Z(n5670) );
  NAND U8981 ( .A(n5668), .B(n5667), .Z(n5669) );
  NAND U8982 ( .A(n5670), .B(n5669), .Z(n8225) );
  XOR U8983 ( .A(n8226), .B(n8225), .Z(n8228) );
  XOR U8984 ( .A(n8227), .B(n8228), .Z(n7929) );
  XOR U8985 ( .A(n7930), .B(n7929), .Z(n7931) );
  XOR U8986 ( .A(n7932), .B(n7931), .Z(n7899) );
  NANDN U8987 ( .A(n5672), .B(n5671), .Z(n5676) );
  NANDN U8988 ( .A(n5674), .B(n5673), .Z(n5675) );
  AND U8989 ( .A(n5676), .B(n5675), .Z(n7926) );
  NANDN U8990 ( .A(n5678), .B(n5677), .Z(n5682) );
  NAND U8991 ( .A(n5680), .B(n5679), .Z(n5681) );
  AND U8992 ( .A(n5682), .B(n5681), .Z(n8500) );
  NANDN U8993 ( .A(n5684), .B(n5683), .Z(n5688) );
  NAND U8994 ( .A(n5686), .B(n5685), .Z(n5687) );
  AND U8995 ( .A(n5688), .B(n5687), .Z(n8499) );
  NANDN U8996 ( .A(n5690), .B(n5689), .Z(n5694) );
  NAND U8997 ( .A(n5692), .B(n5691), .Z(n5693) );
  NAND U8998 ( .A(n5694), .B(n5693), .Z(n8498) );
  XOR U8999 ( .A(n8499), .B(n8498), .Z(n8501) );
  XOR U9000 ( .A(n8500), .B(n8501), .Z(n7925) );
  XOR U9001 ( .A(n7926), .B(n7925), .Z(n7928) );
  NANDN U9002 ( .A(n5696), .B(n5695), .Z(n5700) );
  NANDN U9003 ( .A(n5698), .B(n5697), .Z(n5699) );
  AND U9004 ( .A(n5700), .B(n5699), .Z(n7927) );
  XOR U9005 ( .A(n7928), .B(n7927), .Z(n7898) );
  NANDN U9006 ( .A(n5702), .B(n5701), .Z(n5706) );
  NANDN U9007 ( .A(n5704), .B(n5703), .Z(n5705) );
  AND U9008 ( .A(n5706), .B(n5705), .Z(n8060) );
  NANDN U9009 ( .A(n5708), .B(n5707), .Z(n5712) );
  NAND U9010 ( .A(n5710), .B(n5709), .Z(n5711) );
  AND U9011 ( .A(n5712), .B(n5711), .Z(n8494) );
  NANDN U9012 ( .A(n5714), .B(n5713), .Z(n5718) );
  NAND U9013 ( .A(n5716), .B(n5715), .Z(n5717) );
  AND U9014 ( .A(n5718), .B(n5717), .Z(n8493) );
  NANDN U9015 ( .A(n5720), .B(n5719), .Z(n5724) );
  NAND U9016 ( .A(n5722), .B(n5721), .Z(n5723) );
  NAND U9017 ( .A(n5724), .B(n5723), .Z(n8492) );
  XOR U9018 ( .A(n8493), .B(n8492), .Z(n8495) );
  XOR U9019 ( .A(n8494), .B(n8495), .Z(n8059) );
  XOR U9020 ( .A(n8060), .B(n8059), .Z(n8062) );
  NANDN U9021 ( .A(n5726), .B(n5725), .Z(n5730) );
  NANDN U9022 ( .A(n5728), .B(n5727), .Z(n5729) );
  AND U9023 ( .A(n5730), .B(n5729), .Z(n8061) );
  XNOR U9024 ( .A(n8062), .B(n8061), .Z(n7897) );
  XOR U9025 ( .A(n7898), .B(n7897), .Z(n7900) );
  XOR U9026 ( .A(n7899), .B(n7900), .Z(n7846) );
  NANDN U9027 ( .A(n5732), .B(n5731), .Z(n5736) );
  OR U9028 ( .A(n5734), .B(n5733), .Z(n5735) );
  AND U9029 ( .A(n5736), .B(n5735), .Z(n7936) );
  NANDN U9030 ( .A(n5738), .B(n5737), .Z(n5742) );
  NANDN U9031 ( .A(n5740), .B(n5739), .Z(n5741) );
  AND U9032 ( .A(n5742), .B(n5741), .Z(n7934) );
  IV U9033 ( .A(n5743), .Z(n5745) );
  NANDN U9034 ( .A(n5745), .B(n5744), .Z(n5749) );
  NAND U9035 ( .A(n5747), .B(n5746), .Z(n5748) );
  NAND U9036 ( .A(n5749), .B(n5748), .Z(n8453) );
  XOR U9037 ( .A(n8451), .B(n8452), .Z(n8454) );
  XOR U9038 ( .A(n8453), .B(n8454), .Z(n7933) );
  XOR U9039 ( .A(n7934), .B(n7933), .Z(n7935) );
  XOR U9040 ( .A(n7936), .B(n7935), .Z(n7749) );
  NANDN U9041 ( .A(n5759), .B(n5758), .Z(n5763) );
  NANDN U9042 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U9043 ( .A(n5763), .B(n5762), .Z(n7966) );
  XOR U9044 ( .A(n8459), .B(n8460), .Z(n8462) );
  XOR U9045 ( .A(n8461), .B(n8462), .Z(n7965) );
  XOR U9046 ( .A(n7966), .B(n7965), .Z(n7968) );
  NANDN U9047 ( .A(n5777), .B(n5776), .Z(n5781) );
  NANDN U9048 ( .A(n5779), .B(n5778), .Z(n5780) );
  AND U9049 ( .A(n5781), .B(n5780), .Z(n7967) );
  XOR U9050 ( .A(n7968), .B(n7967), .Z(n7748) );
  NANDN U9051 ( .A(n5783), .B(n5782), .Z(n5787) );
  NANDN U9052 ( .A(n5785), .B(n5784), .Z(n5786) );
  AND U9053 ( .A(n5787), .B(n5786), .Z(n8058) );
  NANDN U9054 ( .A(n5789), .B(n5788), .Z(n5793) );
  NANDN U9055 ( .A(n5791), .B(n5790), .Z(n5792) );
  AND U9056 ( .A(n5793), .B(n5792), .Z(n8056) );
  NANDN U9057 ( .A(n5795), .B(n5794), .Z(n5799) );
  NANDN U9058 ( .A(n5797), .B(n5796), .Z(n5798) );
  AND U9059 ( .A(n5799), .B(n5798), .Z(n7674) );
  NANDN U9060 ( .A(n5805), .B(n5804), .Z(n5809) );
  NAND U9061 ( .A(n5807), .B(n5806), .Z(n5808) );
  NAND U9062 ( .A(n5809), .B(n5808), .Z(n7671) );
  XOR U9063 ( .A(n8056), .B(n8055), .Z(n8057) );
  XNOR U9064 ( .A(n8058), .B(n8057), .Z(n7747) );
  XOR U9065 ( .A(n7748), .B(n7747), .Z(n7750) );
  XOR U9066 ( .A(n7749), .B(n7750), .Z(n7844) );
  NANDN U9067 ( .A(n5811), .B(n5810), .Z(n5815) );
  OR U9068 ( .A(n5813), .B(n5812), .Z(n5814) );
  AND U9069 ( .A(n5815), .B(n5814), .Z(n7843) );
  XNOR U9070 ( .A(n7844), .B(n7843), .Z(n7845) );
  XNOR U9071 ( .A(n7846), .B(n7845), .Z(n7787) );
  XNOR U9072 ( .A(n7788), .B(n7787), .Z(n7790) );
  NANDN U9073 ( .A(n5817), .B(n5816), .Z(n5821) );
  OR U9074 ( .A(n5819), .B(n5818), .Z(n5820) );
  AND U9075 ( .A(n5821), .B(n5820), .Z(n7789) );
  XOR U9076 ( .A(n7790), .B(n7789), .Z(n8372) );
  NANDN U9077 ( .A(n5827), .B(n5826), .Z(n5831) );
  NANDN U9078 ( .A(n5829), .B(n5828), .Z(n5830) );
  AND U9079 ( .A(n5831), .B(n5830), .Z(n8288) );
  NANDN U9080 ( .A(n5833), .B(n5832), .Z(n5837) );
  NAND U9081 ( .A(n5835), .B(n5834), .Z(n5836) );
  AND U9082 ( .A(n5837), .B(n5836), .Z(n8004) );
  NANDN U9083 ( .A(n5839), .B(n5838), .Z(n5843) );
  NAND U9084 ( .A(n5841), .B(n5840), .Z(n5842) );
  AND U9085 ( .A(n5843), .B(n5842), .Z(n8002) );
  NAND U9086 ( .A(n5845), .B(n5844), .Z(n5849) );
  NAND U9087 ( .A(n5847), .B(n5846), .Z(n5848) );
  NAND U9088 ( .A(n5849), .B(n5848), .Z(n8001) );
  XNOR U9089 ( .A(n8002), .B(n8001), .Z(n8003) );
  XNOR U9090 ( .A(n8004), .B(n8003), .Z(n7659) );
  NAND U9091 ( .A(n5851), .B(n5850), .Z(n5855) );
  NAND U9092 ( .A(n5853), .B(n5852), .Z(n5854) );
  AND U9093 ( .A(n5855), .B(n5854), .Z(n8010) );
  NANDN U9094 ( .A(n5857), .B(n5856), .Z(n5861) );
  NAND U9095 ( .A(n5859), .B(n5858), .Z(n5860) );
  AND U9096 ( .A(n5861), .B(n5860), .Z(n8008) );
  NANDN U9097 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U9098 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U9099 ( .A(n5867), .B(n5866), .Z(n8007) );
  XNOR U9100 ( .A(n8008), .B(n8007), .Z(n8009) );
  XOR U9101 ( .A(n8010), .B(n8009), .Z(n7660) );
  XNOR U9102 ( .A(n7659), .B(n7660), .Z(n7662) );
  NANDN U9103 ( .A(n5869), .B(n5868), .Z(n5873) );
  NANDN U9104 ( .A(n5871), .B(n5870), .Z(n5872) );
  AND U9105 ( .A(n5873), .B(n5872), .Z(n7626) );
  NANDN U9106 ( .A(n5879), .B(n5878), .Z(n5883) );
  NAND U9107 ( .A(n5881), .B(n5880), .Z(n5882) );
  NAND U9108 ( .A(n5883), .B(n5882), .Z(n7623) );
  XNOR U9109 ( .A(n7624), .B(n7623), .Z(n7625) );
  XNOR U9110 ( .A(n7626), .B(n7625), .Z(n7661) );
  XNOR U9111 ( .A(n7662), .B(n7661), .Z(n8287) );
  XNOR U9112 ( .A(n8288), .B(n8287), .Z(n8290) );
  NANDN U9113 ( .A(n5893), .B(n5892), .Z(n5897) );
  NANDN U9114 ( .A(n5895), .B(n5894), .Z(n5896) );
  NAND U9115 ( .A(n5897), .B(n5896), .Z(n7595) );
  XNOR U9116 ( .A(n7596), .B(n7595), .Z(n7597) );
  XOR U9117 ( .A(n7598), .B(n7597), .Z(n8257) );
  XNOR U9118 ( .A(n7548), .B(n7547), .Z(n7549) );
  XOR U9119 ( .A(n7550), .B(n7549), .Z(n8255) );
  NAND U9120 ( .A(n5911), .B(n5910), .Z(n5915) );
  NAND U9121 ( .A(n5913), .B(n5912), .Z(n5914) );
  AND U9122 ( .A(n5915), .B(n5914), .Z(n8256) );
  XOR U9123 ( .A(n8255), .B(n8256), .Z(n8258) );
  XOR U9124 ( .A(n8257), .B(n8258), .Z(n8289) );
  XOR U9125 ( .A(n8290), .B(n8289), .Z(n7455) );
  XNOR U9126 ( .A(n7456), .B(n7455), .Z(n7458) );
  NANDN U9127 ( .A(n5917), .B(n5916), .Z(n5921) );
  NANDN U9128 ( .A(n5919), .B(n5918), .Z(n5920) );
  AND U9129 ( .A(n5921), .B(n5920), .Z(n7579) );
  NANDN U9130 ( .A(n5923), .B(n5922), .Z(n5927) );
  NAND U9131 ( .A(n5925), .B(n5924), .Z(n5926) );
  AND U9132 ( .A(n5927), .B(n5926), .Z(n8204) );
  NANDN U9133 ( .A(n5929), .B(n5928), .Z(n5933) );
  NAND U9134 ( .A(n5931), .B(n5930), .Z(n5932) );
  AND U9135 ( .A(n5933), .B(n5932), .Z(n8202) );
  NANDN U9136 ( .A(n5935), .B(n5934), .Z(n5939) );
  NAND U9137 ( .A(n5937), .B(n5936), .Z(n5938) );
  NAND U9138 ( .A(n5939), .B(n5938), .Z(n8201) );
  XNOR U9139 ( .A(n8202), .B(n8201), .Z(n8203) );
  XOR U9140 ( .A(n8204), .B(n8203), .Z(n7580) );
  XNOR U9141 ( .A(n7579), .B(n7580), .Z(n7582) );
  XOR U9142 ( .A(n7582), .B(n7581), .Z(n8284) );
  NANDN U9143 ( .A(n5949), .B(n5948), .Z(n5953) );
  NANDN U9144 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U9145 ( .A(n5953), .B(n5952), .Z(n7573) );
  NANDN U9146 ( .A(n5955), .B(n5954), .Z(n5959) );
  NAND U9147 ( .A(n5957), .B(n5956), .Z(n5958) );
  NAND U9148 ( .A(n5959), .B(n5958), .Z(n7571) );
  XOR U9149 ( .A(n7571), .B(n7572), .Z(n7574) );
  XOR U9150 ( .A(n7573), .B(n7574), .Z(n7575) );
  XOR U9151 ( .A(n7576), .B(n7575), .Z(n7578) );
  NANDN U9152 ( .A(n5965), .B(n5964), .Z(n5969) );
  NANDN U9153 ( .A(n5967), .B(n5966), .Z(n5968) );
  AND U9154 ( .A(n5969), .B(n5968), .Z(n7577) );
  XOR U9155 ( .A(n7578), .B(n7577), .Z(n8282) );
  NANDN U9156 ( .A(n5971), .B(n5970), .Z(n5975) );
  OR U9157 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U9158 ( .A(n5975), .B(n5974), .Z(n8281) );
  XNOR U9159 ( .A(n8282), .B(n8281), .Z(n8283) );
  XNOR U9160 ( .A(n8284), .B(n8283), .Z(n7457) );
  XOR U9161 ( .A(n7458), .B(n7457), .Z(n7795) );
  NANDN U9162 ( .A(n5977), .B(n5976), .Z(n5981) );
  OR U9163 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U9164 ( .A(n5981), .B(n5980), .Z(n8123) );
  NANDN U9165 ( .A(n5983), .B(n5982), .Z(n5987) );
  NANDN U9166 ( .A(n5985), .B(n5984), .Z(n5986) );
  AND U9167 ( .A(n5987), .B(n5986), .Z(n8148) );
  NANDN U9168 ( .A(n5989), .B(n5988), .Z(n5993) );
  NAND U9169 ( .A(n5991), .B(n5990), .Z(n5992) );
  NAND U9170 ( .A(n5993), .B(n5992), .Z(n7631) );
  XOR U9171 ( .A(n7629), .B(n7630), .Z(n7632) );
  XOR U9172 ( .A(n7631), .B(n7632), .Z(n8145) );
  NANDN U9173 ( .A(n6003), .B(n6002), .Z(n6007) );
  NANDN U9174 ( .A(n6005), .B(n6004), .Z(n6006) );
  NAND U9175 ( .A(n6007), .B(n6006), .Z(n7639) );
  XNOR U9176 ( .A(n7637), .B(n7638), .Z(n7640) );
  XOR U9177 ( .A(n7639), .B(n7640), .Z(n8146) );
  XNOR U9178 ( .A(n8145), .B(n8146), .Z(n8147) );
  XOR U9179 ( .A(n8148), .B(n8147), .Z(n7992) );
  NANDN U9180 ( .A(n6021), .B(n6020), .Z(n6025) );
  NANDN U9181 ( .A(n6023), .B(n6022), .Z(n6024) );
  AND U9182 ( .A(n6025), .B(n6024), .Z(n7650) );
  NANDN U9183 ( .A(n6027), .B(n6026), .Z(n6031) );
  NANDN U9184 ( .A(n6029), .B(n6028), .Z(n6030) );
  AND U9185 ( .A(n6031), .B(n6030), .Z(n7647) );
  NANDN U9186 ( .A(n6037), .B(n6036), .Z(n6041) );
  NAND U9187 ( .A(n6039), .B(n6038), .Z(n6040) );
  NAND U9188 ( .A(n6041), .B(n6040), .Z(n7553) );
  XNOR U9189 ( .A(n7553), .B(n7554), .Z(n7556) );
  XOR U9190 ( .A(n7555), .B(n7556), .Z(n7648) );
  XNOR U9191 ( .A(n7647), .B(n7648), .Z(n7649) );
  XNOR U9192 ( .A(n7650), .B(n7649), .Z(n7989) );
  XNOR U9193 ( .A(n7990), .B(n7989), .Z(n7991) );
  XOR U9194 ( .A(n7992), .B(n7991), .Z(n8124) );
  XNOR U9195 ( .A(n8123), .B(n8124), .Z(n8126) );
  NANDN U9196 ( .A(n6047), .B(n6046), .Z(n6051) );
  NAND U9197 ( .A(n6049), .B(n6048), .Z(n6050) );
  AND U9198 ( .A(n6051), .B(n6050), .Z(n8457) );
  XNOR U9199 ( .A(n8456), .B(n8455), .Z(n8458) );
  XNOR U9200 ( .A(n8457), .B(n8458), .Z(n8238) );
  IV U9201 ( .A(n6060), .Z(n6061) );
  ANDN U9202 ( .B(n6062), .A(n6061), .Z(n8450) );
  NANDN U9203 ( .A(n6064), .B(n6063), .Z(n6068) );
  NANDN U9204 ( .A(n6066), .B(n6065), .Z(n6067) );
  AND U9205 ( .A(n6068), .B(n6067), .Z(n8449) );
  XOR U9206 ( .A(n8450), .B(n8449), .Z(n7679) );
  NANDN U9207 ( .A(n6070), .B(n6069), .Z(n6074) );
  NAND U9208 ( .A(n6072), .B(n6071), .Z(n6073) );
  NAND U9209 ( .A(n6074), .B(n6073), .Z(n7677) );
  XNOR U9210 ( .A(n7677), .B(n7678), .Z(n7680) );
  XOR U9211 ( .A(n7679), .B(n7680), .Z(n8237) );
  XOR U9212 ( .A(n8238), .B(n8237), .Z(n8240) );
  NANDN U9213 ( .A(n6084), .B(n6083), .Z(n6088) );
  NANDN U9214 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U9215 ( .A(n6088), .B(n6087), .Z(n7681) );
  NANDN U9216 ( .A(n6090), .B(n6089), .Z(n6094) );
  NAND U9217 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U9218 ( .A(n6094), .B(n6093), .Z(n7682) );
  XOR U9219 ( .A(n7681), .B(n7682), .Z(n7684) );
  XOR U9220 ( .A(n7683), .B(n7684), .Z(n8239) );
  XOR U9221 ( .A(n8240), .B(n8239), .Z(n7894) );
  NANDN U9222 ( .A(n6100), .B(n6099), .Z(n6104) );
  NANDN U9223 ( .A(n6102), .B(n6101), .Z(n6103) );
  AND U9224 ( .A(n6104), .B(n6103), .Z(n8139) );
  NANDN U9225 ( .A(n6106), .B(n6105), .Z(n6110) );
  NANDN U9226 ( .A(n6108), .B(n6107), .Z(n6109) );
  NAND U9227 ( .A(n6110), .B(n6109), .Z(n8187) );
  NANDN U9228 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U9229 ( .A(n6114), .B(n6113), .Z(n6115) );
  NAND U9230 ( .A(n6116), .B(n6115), .Z(n8185) );
  NANDN U9231 ( .A(n6118), .B(n6117), .Z(n6122) );
  NAND U9232 ( .A(n6120), .B(n6119), .Z(n6121) );
  NAND U9233 ( .A(n6122), .B(n6121), .Z(n8186) );
  XNOR U9234 ( .A(n8185), .B(n8186), .Z(n8188) );
  XOR U9235 ( .A(n8187), .B(n8188), .Z(n8140) );
  XNOR U9236 ( .A(n8139), .B(n8140), .Z(n8142) );
  NANDN U9237 ( .A(n6124), .B(n6123), .Z(n6128) );
  NANDN U9238 ( .A(n6126), .B(n6125), .Z(n6127) );
  AND U9239 ( .A(n6128), .B(n6127), .Z(n8141) );
  XNOR U9240 ( .A(n8142), .B(n8141), .Z(n7891) );
  XNOR U9241 ( .A(n7892), .B(n7891), .Z(n7893) );
  XNOR U9242 ( .A(n7894), .B(n7893), .Z(n8125) );
  XOR U9243 ( .A(n8126), .B(n8125), .Z(n7794) );
  NANDN U9244 ( .A(n6134), .B(n6133), .Z(n6138) );
  NAND U9245 ( .A(n6136), .B(n6135), .Z(n6137) );
  AND U9246 ( .A(n6138), .B(n6137), .Z(n7986) );
  NANDN U9247 ( .A(n6140), .B(n6139), .Z(n6144) );
  NANDN U9248 ( .A(n6142), .B(n6141), .Z(n6143) );
  AND U9249 ( .A(n6144), .B(n6143), .Z(n8321) );
  NANDN U9250 ( .A(n6146), .B(n6145), .Z(n6150) );
  NANDN U9251 ( .A(n6148), .B(n6147), .Z(n6149) );
  NAND U9252 ( .A(n6150), .B(n6149), .Z(n8271) );
  NANDN U9253 ( .A(n6152), .B(n6151), .Z(n6156) );
  NANDN U9254 ( .A(n6154), .B(n6153), .Z(n6155) );
  NAND U9255 ( .A(n6156), .B(n6155), .Z(n8269) );
  NANDN U9256 ( .A(n6158), .B(n6157), .Z(n6162) );
  NANDN U9257 ( .A(n6160), .B(n6159), .Z(n6161) );
  NAND U9258 ( .A(n6162), .B(n6161), .Z(n8270) );
  XNOR U9259 ( .A(n8269), .B(n8270), .Z(n8272) );
  XOR U9260 ( .A(n8271), .B(n8272), .Z(n8322) );
  XNOR U9261 ( .A(n8321), .B(n8322), .Z(n8324) );
  NANDN U9262 ( .A(n6164), .B(n6163), .Z(n6168) );
  NANDN U9263 ( .A(n6166), .B(n6165), .Z(n6167) );
  AND U9264 ( .A(n6168), .B(n6167), .Z(n8323) );
  XOR U9265 ( .A(n8324), .B(n8323), .Z(n7984) );
  NANDN U9266 ( .A(n6170), .B(n6169), .Z(n6174) );
  NANDN U9267 ( .A(n6172), .B(n6171), .Z(n6173) );
  AND U9268 ( .A(n6174), .B(n6173), .Z(n8318) );
  NANDN U9269 ( .A(n6176), .B(n6175), .Z(n6180) );
  NANDN U9270 ( .A(n6178), .B(n6177), .Z(n6179) );
  AND U9271 ( .A(n6180), .B(n6179), .Z(n8233) );
  NANDN U9272 ( .A(n6182), .B(n6181), .Z(n6186) );
  NAND U9273 ( .A(n6184), .B(n6183), .Z(n6185) );
  AND U9274 ( .A(n6186), .B(n6185), .Z(n8232) );
  NANDN U9275 ( .A(n6188), .B(n6187), .Z(n6192) );
  NAND U9276 ( .A(n6190), .B(n6189), .Z(n6191) );
  NAND U9277 ( .A(n6192), .B(n6191), .Z(n8231) );
  XOR U9278 ( .A(n8232), .B(n8231), .Z(n8234) );
  XOR U9279 ( .A(n8233), .B(n8234), .Z(n8317) );
  XOR U9280 ( .A(n8318), .B(n8317), .Z(n8320) );
  NANDN U9281 ( .A(n6194), .B(n6193), .Z(n6198) );
  NANDN U9282 ( .A(n6196), .B(n6195), .Z(n6197) );
  AND U9283 ( .A(n6198), .B(n6197), .Z(n8319) );
  XNOR U9284 ( .A(n8320), .B(n8319), .Z(n7983) );
  XNOR U9285 ( .A(n7984), .B(n7983), .Z(n7985) );
  XNOR U9286 ( .A(n7986), .B(n7985), .Z(n8117) );
  XNOR U9287 ( .A(n8118), .B(n8117), .Z(n8120) );
  NANDN U9288 ( .A(n6200), .B(n6199), .Z(n6204) );
  NANDN U9289 ( .A(n6202), .B(n6201), .Z(n6203) );
  AND U9290 ( .A(n6204), .B(n6203), .Z(n8114) );
  NANDN U9291 ( .A(n6206), .B(n6205), .Z(n6210) );
  NANDN U9292 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U9293 ( .A(n6210), .B(n6209), .Z(n7964) );
  NANDN U9294 ( .A(n6212), .B(n6211), .Z(n6216) );
  NANDN U9295 ( .A(n6214), .B(n6213), .Z(n6215) );
  AND U9296 ( .A(n6216), .B(n6215), .Z(n7962) );
  NANDN U9297 ( .A(n6218), .B(n6217), .Z(n6222) );
  NANDN U9298 ( .A(n6220), .B(n6219), .Z(n6221) );
  AND U9299 ( .A(n6222), .B(n6221), .Z(n8209) );
  NANDN U9300 ( .A(n6224), .B(n6223), .Z(n6228) );
  NANDN U9301 ( .A(n6226), .B(n6225), .Z(n6227) );
  AND U9302 ( .A(n6228), .B(n6227), .Z(n8208) );
  NANDN U9303 ( .A(n6230), .B(n6229), .Z(n6234) );
  NAND U9304 ( .A(n6232), .B(n6231), .Z(n6233) );
  NAND U9305 ( .A(n6234), .B(n6233), .Z(n8207) );
  XOR U9306 ( .A(n8208), .B(n8207), .Z(n8210) );
  XOR U9307 ( .A(n8209), .B(n8210), .Z(n7961) );
  XOR U9308 ( .A(n7962), .B(n7961), .Z(n7963) );
  XOR U9309 ( .A(n7964), .B(n7963), .Z(n8112) );
  NANDN U9310 ( .A(n6236), .B(n6235), .Z(n6240) );
  NANDN U9311 ( .A(n6238), .B(n6237), .Z(n6239) );
  AND U9312 ( .A(n6240), .B(n6239), .Z(n7955) );
  NANDN U9313 ( .A(n6242), .B(n6241), .Z(n6246) );
  NAND U9314 ( .A(n6244), .B(n6243), .Z(n6245) );
  NAND U9315 ( .A(n6246), .B(n6245), .Z(n8275) );
  NANDN U9316 ( .A(n6248), .B(n6247), .Z(n6252) );
  NANDN U9317 ( .A(n6250), .B(n6249), .Z(n6251) );
  NAND U9318 ( .A(n6252), .B(n6251), .Z(n8273) );
  NANDN U9319 ( .A(n6254), .B(n6253), .Z(n6258) );
  NANDN U9320 ( .A(n6256), .B(n6255), .Z(n6257) );
  NAND U9321 ( .A(n6258), .B(n6257), .Z(n8274) );
  XNOR U9322 ( .A(n8273), .B(n8274), .Z(n8276) );
  XOR U9323 ( .A(n8275), .B(n8276), .Z(n7956) );
  XNOR U9324 ( .A(n7955), .B(n7956), .Z(n7958) );
  NANDN U9325 ( .A(n6260), .B(n6259), .Z(n6264) );
  NANDN U9326 ( .A(n6262), .B(n6261), .Z(n6263) );
  AND U9327 ( .A(n6264), .B(n6263), .Z(n7957) );
  XNOR U9328 ( .A(n7958), .B(n7957), .Z(n8111) );
  XNOR U9329 ( .A(n8112), .B(n8111), .Z(n8113) );
  XNOR U9330 ( .A(n8114), .B(n8113), .Z(n8119) );
  XNOR U9331 ( .A(n8120), .B(n8119), .Z(n7793) );
  XOR U9332 ( .A(n7794), .B(n7793), .Z(n7796) );
  XOR U9333 ( .A(n7795), .B(n7796), .Z(n8370) );
  NAND U9334 ( .A(n6266), .B(n6265), .Z(n6270) );
  NANDN U9335 ( .A(n6268), .B(n6267), .Z(n6269) );
  AND U9336 ( .A(n6270), .B(n6269), .Z(n8519) );
  NANDN U9337 ( .A(n6272), .B(n6271), .Z(n6276) );
  NANDN U9338 ( .A(n6274), .B(n6273), .Z(n6275) );
  AND U9339 ( .A(n6276), .B(n6275), .Z(n8108) );
  NANDN U9340 ( .A(n6278), .B(n6277), .Z(n6282) );
  NANDN U9341 ( .A(n6280), .B(n6279), .Z(n6281) );
  NAND U9342 ( .A(n6282), .B(n6281), .Z(n7565) );
  NANDN U9343 ( .A(n6284), .B(n6283), .Z(n6288) );
  NANDN U9344 ( .A(n6286), .B(n6285), .Z(n6287) );
  NAND U9345 ( .A(n6288), .B(n6287), .Z(n7563) );
  NANDN U9346 ( .A(n6290), .B(n6289), .Z(n6294) );
  NANDN U9347 ( .A(n6292), .B(n6291), .Z(n6293) );
  NAND U9348 ( .A(n6294), .B(n6293), .Z(n7564) );
  XOR U9349 ( .A(n7563), .B(n7564), .Z(n7566) );
  XOR U9350 ( .A(n7565), .B(n7566), .Z(n8107) );
  XOR U9351 ( .A(n8108), .B(n8107), .Z(n8110) );
  NANDN U9352 ( .A(n6296), .B(n6295), .Z(n6300) );
  NANDN U9353 ( .A(n6298), .B(n6297), .Z(n6299) );
  AND U9354 ( .A(n6300), .B(n6299), .Z(n8109) );
  XOR U9355 ( .A(n8110), .B(n8109), .Z(n7725) );
  NANDN U9356 ( .A(n6306), .B(n6305), .Z(n6310) );
  NAND U9357 ( .A(n6308), .B(n6307), .Z(n6309) );
  NAND U9358 ( .A(n6310), .B(n6309), .Z(n7723) );
  XOR U9359 ( .A(n7724), .B(n7723), .Z(n7726) );
  XOR U9360 ( .A(n7725), .B(n7726), .Z(n8308) );
  NANDN U9361 ( .A(n6312), .B(n6311), .Z(n6316) );
  NANDN U9362 ( .A(n6314), .B(n6313), .Z(n6315) );
  AND U9363 ( .A(n6316), .B(n6315), .Z(n7560) );
  NANDN U9364 ( .A(n6318), .B(n6317), .Z(n6322) );
  NANDN U9365 ( .A(n6320), .B(n6319), .Z(n6321) );
  AND U9366 ( .A(n6322), .B(n6321), .Z(n7557) );
  NANDN U9367 ( .A(n6332), .B(n6331), .Z(n6336) );
  NAND U9368 ( .A(n6334), .B(n6333), .Z(n6335) );
  NAND U9369 ( .A(n6336), .B(n6335), .Z(n8421) );
  XNOR U9370 ( .A(n8422), .B(n8421), .Z(n8423) );
  XOR U9371 ( .A(n8424), .B(n8423), .Z(n7558) );
  XNOR U9372 ( .A(n7557), .B(n7558), .Z(n7559) );
  XOR U9373 ( .A(n7560), .B(n7559), .Z(n7767) );
  NAND U9374 ( .A(n6342), .B(n6341), .Z(n6346) );
  NAND U9375 ( .A(n6344), .B(n6343), .Z(n6345) );
  AND U9376 ( .A(n6346), .B(n6345), .Z(n8446) );
  NANDN U9377 ( .A(n6348), .B(n6347), .Z(n6352) );
  NANDN U9378 ( .A(n6350), .B(n6349), .Z(n6351) );
  AND U9379 ( .A(n6352), .B(n6351), .Z(n8444) );
  NANDN U9380 ( .A(n6354), .B(n6353), .Z(n6358) );
  NAND U9381 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U9382 ( .A(n6358), .B(n6357), .Z(n8443) );
  XNOR U9383 ( .A(n8444), .B(n8443), .Z(n8445) );
  XNOR U9384 ( .A(n8446), .B(n8445), .Z(n8083) );
  XOR U9385 ( .A(n8084), .B(n8083), .Z(n8086) );
  XOR U9386 ( .A(n8086), .B(n8085), .Z(n7766) );
  NANDN U9387 ( .A(n6364), .B(n6363), .Z(n6368) );
  NANDN U9388 ( .A(n6366), .B(n6365), .Z(n6367) );
  NAND U9389 ( .A(n6368), .B(n6367), .Z(n7765) );
  XOR U9390 ( .A(n7766), .B(n7765), .Z(n7768) );
  XOR U9391 ( .A(n7767), .B(n7768), .Z(n8306) );
  NANDN U9392 ( .A(n6370), .B(n6369), .Z(n6374) );
  NAND U9393 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U9394 ( .A(n6374), .B(n6373), .Z(n8305) );
  XNOR U9395 ( .A(n8306), .B(n8305), .Z(n8307) );
  XOR U9396 ( .A(n8308), .B(n8307), .Z(n8517) );
  NAND U9397 ( .A(n6376), .B(n6375), .Z(n6380) );
  NAND U9398 ( .A(n6378), .B(n6377), .Z(n6379) );
  NAND U9399 ( .A(n6380), .B(n6379), .Z(n8516) );
  XOR U9400 ( .A(n8517), .B(n8516), .Z(n8518) );
  XOR U9401 ( .A(n8519), .B(n8518), .Z(n8369) );
  XNOR U9402 ( .A(n8370), .B(n8369), .Z(n8371) );
  XNOR U9403 ( .A(n8372), .B(n8371), .Z(n7806) );
  XOR U9404 ( .A(n7805), .B(n7806), .Z(n7808) );
  NANDN U9405 ( .A(n6398), .B(n6397), .Z(n6402) );
  NANDN U9406 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U9407 ( .A(n6402), .B(n6401), .Z(n8242) );
  NANDN U9408 ( .A(n6404), .B(n6403), .Z(n6408) );
  NAND U9409 ( .A(n6406), .B(n6405), .Z(n6407) );
  NAND U9410 ( .A(n6408), .B(n6407), .Z(n8241) );
  XNOR U9411 ( .A(n8242), .B(n8241), .Z(n8243) );
  XOR U9412 ( .A(n8244), .B(n8243), .Z(n7500) );
  XOR U9413 ( .A(n7499), .B(n7500), .Z(n7502) );
  XOR U9414 ( .A(n7501), .B(n7502), .Z(n8068) );
  XNOR U9415 ( .A(n8067), .B(n8068), .Z(n8070) );
  NAND U9416 ( .A(n6414), .B(n6413), .Z(n6418) );
  NAND U9417 ( .A(n6416), .B(n6415), .Z(n6417) );
  AND U9418 ( .A(n6418), .B(n6417), .Z(n8440) );
  NANDN U9419 ( .A(n6420), .B(n6419), .Z(n6424) );
  NAND U9420 ( .A(n6422), .B(n6421), .Z(n6423) );
  AND U9421 ( .A(n6424), .B(n6423), .Z(n8438) );
  NAND U9422 ( .A(n6426), .B(n6425), .Z(n6430) );
  NAND U9423 ( .A(n6428), .B(n6427), .Z(n6429) );
  NAND U9424 ( .A(n6430), .B(n6429), .Z(n8437) );
  XOR U9425 ( .A(n8260), .B(n8259), .Z(n8261) );
  XNOR U9426 ( .A(n8261), .B(n8262), .Z(n8069) );
  XOR U9427 ( .A(n8070), .B(n8069), .Z(n7869) );
  NANDN U9428 ( .A(n6436), .B(n6435), .Z(n6440) );
  NANDN U9429 ( .A(n6438), .B(n6437), .Z(n6439) );
  AND U9430 ( .A(n6440), .B(n6439), .Z(n7867) );
  NANDN U9431 ( .A(n6442), .B(n6441), .Z(n6446) );
  NANDN U9432 ( .A(n6444), .B(n6443), .Z(n6445) );
  NAND U9433 ( .A(n6446), .B(n6445), .Z(n7511) );
  XOR U9434 ( .A(n7509), .B(n7510), .Z(n7512) );
  XOR U9435 ( .A(n7511), .B(n7512), .Z(n8161) );
  NANDN U9436 ( .A(n6456), .B(n6455), .Z(n6460) );
  NANDN U9437 ( .A(n6458), .B(n6457), .Z(n6459) );
  AND U9438 ( .A(n6460), .B(n6459), .Z(n8489) );
  NANDN U9439 ( .A(n6462), .B(n6461), .Z(n6466) );
  NAND U9440 ( .A(n6464), .B(n6463), .Z(n6465) );
  AND U9441 ( .A(n6466), .B(n6465), .Z(n8487) );
  NANDN U9442 ( .A(n6468), .B(n6467), .Z(n6472) );
  NAND U9443 ( .A(n6470), .B(n6469), .Z(n6471) );
  NAND U9444 ( .A(n6472), .B(n6471), .Z(n8486) );
  XNOR U9445 ( .A(n8487), .B(n8486), .Z(n8488) );
  XOR U9446 ( .A(n8489), .B(n8488), .Z(n8162) );
  XNOR U9447 ( .A(n8161), .B(n8162), .Z(n8164) );
  NANDN U9448 ( .A(n6482), .B(n6481), .Z(n6486) );
  NAND U9449 ( .A(n6484), .B(n6483), .Z(n6485) );
  NAND U9450 ( .A(n6486), .B(n6485), .Z(n8219) );
  XNOR U9451 ( .A(n8220), .B(n8219), .Z(n8221) );
  XNOR U9452 ( .A(n8222), .B(n8221), .Z(n8163) );
  XOR U9453 ( .A(n8164), .B(n8163), .Z(n8090) );
  NANDN U9454 ( .A(n6488), .B(n6487), .Z(n6492) );
  NANDN U9455 ( .A(n6490), .B(n6489), .Z(n6491) );
  AND U9456 ( .A(n6492), .B(n6491), .Z(n7478) );
  NANDN U9457 ( .A(n6494), .B(n6493), .Z(n6498) );
  NANDN U9458 ( .A(n6496), .B(n6495), .Z(n6497) );
  AND U9459 ( .A(n6498), .B(n6497), .Z(n7475) );
  NANDN U9460 ( .A(n6500), .B(n6499), .Z(n6504) );
  NAND U9461 ( .A(n6502), .B(n6501), .Z(n6503) );
  AND U9462 ( .A(n6504), .B(n6503), .Z(n8198) );
  NANDN U9463 ( .A(n6506), .B(n6505), .Z(n6510) );
  NAND U9464 ( .A(n6508), .B(n6507), .Z(n6509) );
  AND U9465 ( .A(n6510), .B(n6509), .Z(n8196) );
  NANDN U9466 ( .A(n6512), .B(n6511), .Z(n6516) );
  NAND U9467 ( .A(n6514), .B(n6513), .Z(n6515) );
  NAND U9468 ( .A(n6516), .B(n6515), .Z(n8195) );
  XNOR U9469 ( .A(n8196), .B(n8195), .Z(n8197) );
  XOR U9470 ( .A(n8198), .B(n8197), .Z(n7476) );
  XNOR U9471 ( .A(n7475), .B(n7476), .Z(n7477) );
  XOR U9472 ( .A(n7478), .B(n7477), .Z(n8088) );
  XNOR U9473 ( .A(n8088), .B(n8087), .Z(n8089) );
  XOR U9474 ( .A(n8090), .B(n8089), .Z(n7868) );
  XOR U9475 ( .A(n7867), .B(n7868), .Z(n7870) );
  XOR U9476 ( .A(n7869), .B(n7870), .Z(n8396) );
  NANDN U9477 ( .A(n6522), .B(n6521), .Z(n6526) );
  NANDN U9478 ( .A(n6524), .B(n6523), .Z(n6525) );
  NAND U9479 ( .A(n6526), .B(n6525), .Z(n7523) );
  NANDN U9480 ( .A(n6528), .B(n6527), .Z(n6532) );
  NANDN U9481 ( .A(n6530), .B(n6529), .Z(n6531) );
  NAND U9482 ( .A(n6532), .B(n6531), .Z(n7521) );
  NANDN U9483 ( .A(n6534), .B(n6533), .Z(n6538) );
  OR U9484 ( .A(n6536), .B(n6535), .Z(n6537) );
  AND U9485 ( .A(n6538), .B(n6537), .Z(n7522) );
  XOR U9486 ( .A(n7521), .B(n7522), .Z(n7524) );
  XOR U9487 ( .A(n7523), .B(n7524), .Z(n7614) );
  NANDN U9488 ( .A(n6540), .B(n6539), .Z(n6544) );
  NANDN U9489 ( .A(n6542), .B(n6541), .Z(n6543) );
  NAND U9490 ( .A(n6544), .B(n6543), .Z(n7779) );
  NANDN U9491 ( .A(n6550), .B(n6549), .Z(n6554) );
  NANDN U9492 ( .A(n6552), .B(n6551), .Z(n6553) );
  NAND U9493 ( .A(n6554), .B(n6553), .Z(n7778) );
  XOR U9494 ( .A(n7777), .B(n7778), .Z(n7780) );
  XOR U9495 ( .A(n7779), .B(n7780), .Z(n7613) );
  XOR U9496 ( .A(n7614), .B(n7613), .Z(n7616) );
  NANDN U9497 ( .A(n6556), .B(n6555), .Z(n6560) );
  NANDN U9498 ( .A(n6558), .B(n6557), .Z(n6559) );
  AND U9499 ( .A(n6560), .B(n6559), .Z(n7719) );
  NANDN U9500 ( .A(n6566), .B(n6565), .Z(n6570) );
  NANDN U9501 ( .A(n6568), .B(n6567), .Z(n6569) );
  AND U9502 ( .A(n6570), .B(n6569), .Z(n7717) );
  XOR U9503 ( .A(n7718), .B(n7717), .Z(n7720) );
  XNOR U9504 ( .A(n7719), .B(n7720), .Z(n7615) );
  XOR U9505 ( .A(n7616), .B(n7615), .Z(n8394) );
  NANDN U9506 ( .A(n6572), .B(n6571), .Z(n6576) );
  NANDN U9507 ( .A(n6574), .B(n6573), .Z(n6575) );
  AND U9508 ( .A(n6576), .B(n6575), .Z(n7920) );
  NANDN U9509 ( .A(n6578), .B(n6577), .Z(n6582) );
  OR U9510 ( .A(n6580), .B(n6579), .Z(n6581) );
  NAND U9511 ( .A(n6582), .B(n6581), .Z(n7919) );
  XNOR U9512 ( .A(n7920), .B(n7919), .Z(n7921) );
  NANDN U9513 ( .A(n6584), .B(n6583), .Z(n6588) );
  NANDN U9514 ( .A(n6586), .B(n6585), .Z(n6587) );
  AND U9515 ( .A(n6588), .B(n6587), .Z(n7604) );
  NANDN U9516 ( .A(n6590), .B(n6589), .Z(n6594) );
  OR U9517 ( .A(n6592), .B(n6591), .Z(n6593) );
  AND U9518 ( .A(n6594), .B(n6593), .Z(n7602) );
  XNOR U9519 ( .A(n7604), .B(n7603), .Z(n7922) );
  XNOR U9520 ( .A(n7921), .B(n7922), .Z(n8313) );
  NANDN U9521 ( .A(n6600), .B(n6599), .Z(n6604) );
  NAND U9522 ( .A(n6602), .B(n6601), .Z(n6603) );
  NAND U9523 ( .A(n6604), .B(n6603), .Z(n8311) );
  NANDN U9524 ( .A(n6606), .B(n6605), .Z(n6610) );
  NANDN U9525 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U9526 ( .A(n6610), .B(n6609), .Z(n7655) );
  NANDN U9527 ( .A(n6612), .B(n6611), .Z(n6616) );
  NANDN U9528 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U9529 ( .A(n6616), .B(n6615), .Z(n7654) );
  NANDN U9530 ( .A(n6618), .B(n6617), .Z(n6622) );
  NAND U9531 ( .A(n6620), .B(n6619), .Z(n6621) );
  NAND U9532 ( .A(n6622), .B(n6621), .Z(n7653) );
  XOR U9533 ( .A(n7654), .B(n7653), .Z(n7656) );
  XOR U9534 ( .A(n7655), .B(n7656), .Z(n8312) );
  XNOR U9535 ( .A(n8311), .B(n8312), .Z(n8314) );
  XOR U9536 ( .A(n8313), .B(n8314), .Z(n8393) );
  NANDN U9537 ( .A(n6628), .B(n6627), .Z(n6632) );
  NAND U9538 ( .A(n6630), .B(n6629), .Z(n6631) );
  AND U9539 ( .A(n6632), .B(n6631), .Z(n7644) );
  XNOR U9540 ( .A(n7642), .B(n7641), .Z(n7643) );
  XNOR U9541 ( .A(n7644), .B(n7643), .Z(n8167) );
  NANDN U9542 ( .A(n6642), .B(n6641), .Z(n6646) );
  NAND U9543 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U9544 ( .A(n6646), .B(n6645), .Z(n7592) );
  NANDN U9545 ( .A(n6648), .B(n6647), .Z(n6652) );
  NAND U9546 ( .A(n6650), .B(n6649), .Z(n6651) );
  AND U9547 ( .A(n6652), .B(n6651), .Z(n7590) );
  XNOR U9548 ( .A(n7590), .B(n7589), .Z(n7591) );
  XOR U9549 ( .A(n7592), .B(n7591), .Z(n8168) );
  XNOR U9550 ( .A(n8167), .B(n8168), .Z(n8169) );
  NANDN U9551 ( .A(n6662), .B(n6661), .Z(n6666) );
  NANDN U9552 ( .A(n6664), .B(n6663), .Z(n6665) );
  AND U9553 ( .A(n6666), .B(n6665), .Z(n7462) );
  XNOR U9554 ( .A(n7462), .B(n7461), .Z(n7463) );
  XOR U9555 ( .A(n7464), .B(n7463), .Z(n8170) );
  XOR U9556 ( .A(n8169), .B(n8170), .Z(n7712) );
  XNOR U9557 ( .A(n7711), .B(n7712), .Z(n7714) );
  NANDN U9558 ( .A(n6672), .B(n6671), .Z(n6676) );
  NANDN U9559 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U9560 ( .A(n6676), .B(n6675), .Z(n8479) );
  NANDN U9561 ( .A(n6678), .B(n6677), .Z(n6682) );
  NANDN U9562 ( .A(n6680), .B(n6679), .Z(n6681) );
  AND U9563 ( .A(n6682), .B(n6681), .Z(n8477) );
  NANDN U9564 ( .A(n6684), .B(n6683), .Z(n6688) );
  NAND U9565 ( .A(n6686), .B(n6685), .Z(n6687) );
  NAND U9566 ( .A(n6688), .B(n6687), .Z(n8429) );
  NANDN U9567 ( .A(n6690), .B(n6689), .Z(n6694) );
  NAND U9568 ( .A(n6692), .B(n6691), .Z(n6693) );
  NAND U9569 ( .A(n6694), .B(n6693), .Z(n8427) );
  NANDN U9570 ( .A(n6696), .B(n6695), .Z(n6700) );
  NAND U9571 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U9572 ( .A(n6700), .B(n6699), .Z(n8428) );
  XOR U9573 ( .A(n8427), .B(n8428), .Z(n8430) );
  XOR U9574 ( .A(n8429), .B(n8430), .Z(n8476) );
  XOR U9575 ( .A(n8477), .B(n8476), .Z(n8478) );
  XOR U9576 ( .A(n8479), .B(n8478), .Z(n7713) );
  XOR U9577 ( .A(n7714), .B(n7713), .Z(n7608) );
  NANDN U9578 ( .A(n6702), .B(n6701), .Z(n6706) );
  NANDN U9579 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U9580 ( .A(n6706), .B(n6705), .Z(n8130) );
  NANDN U9581 ( .A(n6708), .B(n6707), .Z(n6712) );
  NANDN U9582 ( .A(n6710), .B(n6709), .Z(n6711) );
  AND U9583 ( .A(n6712), .B(n6711), .Z(n8175) );
  NANDN U9584 ( .A(n6718), .B(n6717), .Z(n6722) );
  NAND U9585 ( .A(n6720), .B(n6719), .Z(n6721) );
  NAND U9586 ( .A(n6722), .B(n6721), .Z(n8173) );
  XOR U9587 ( .A(n8174), .B(n8173), .Z(n8176) );
  XOR U9588 ( .A(n8175), .B(n8176), .Z(n8129) );
  XOR U9589 ( .A(n8130), .B(n8129), .Z(n8132) );
  NANDN U9590 ( .A(n6724), .B(n6723), .Z(n6728) );
  NANDN U9591 ( .A(n6726), .B(n6725), .Z(n6727) );
  AND U9592 ( .A(n6728), .B(n6727), .Z(n8131) );
  XOR U9593 ( .A(n8132), .B(n8131), .Z(n7732) );
  NANDN U9594 ( .A(n6734), .B(n6733), .Z(n6738) );
  OR U9595 ( .A(n6736), .B(n6735), .Z(n6737) );
  NAND U9596 ( .A(n6738), .B(n6737), .Z(n8151) );
  XNOR U9597 ( .A(n8032), .B(n8031), .Z(n8033) );
  XNOR U9598 ( .A(n8034), .B(n8033), .Z(n8152) );
  XOR U9599 ( .A(n8151), .B(n8152), .Z(n8154) );
  NANDN U9600 ( .A(n6752), .B(n6751), .Z(n6756) );
  NANDN U9601 ( .A(n6754), .B(n6753), .Z(n6755) );
  AND U9602 ( .A(n6756), .B(n6755), .Z(n8153) );
  XNOR U9603 ( .A(n8154), .B(n8153), .Z(n7729) );
  XNOR U9604 ( .A(n7730), .B(n7729), .Z(n7731) );
  XNOR U9605 ( .A(n7732), .B(n7731), .Z(n7607) );
  XNOR U9606 ( .A(n7608), .B(n7607), .Z(n7609) );
  NANDN U9607 ( .A(n6758), .B(n6757), .Z(n6762) );
  OR U9608 ( .A(n6760), .B(n6759), .Z(n6761) );
  AND U9609 ( .A(n6762), .B(n6761), .Z(n7834) );
  NANDN U9610 ( .A(n6764), .B(n6763), .Z(n6768) );
  NANDN U9611 ( .A(n6766), .B(n6765), .Z(n6767) );
  NAND U9612 ( .A(n6768), .B(n6767), .Z(n7569) );
  NANDN U9613 ( .A(n6770), .B(n6769), .Z(n6774) );
  NANDN U9614 ( .A(n6772), .B(n6771), .Z(n6773) );
  NAND U9615 ( .A(n6774), .B(n6773), .Z(n7567) );
  NANDN U9616 ( .A(n6776), .B(n6775), .Z(n6780) );
  NAND U9617 ( .A(n6778), .B(n6777), .Z(n6779) );
  NAND U9618 ( .A(n6780), .B(n6779), .Z(n7568) );
  XOR U9619 ( .A(n7567), .B(n7568), .Z(n7570) );
  XOR U9620 ( .A(n7569), .B(n7570), .Z(n7833) );
  XOR U9621 ( .A(n7834), .B(n7833), .Z(n7836) );
  NANDN U9622 ( .A(n6782), .B(n6781), .Z(n6786) );
  OR U9623 ( .A(n6784), .B(n6783), .Z(n6785) );
  AND U9624 ( .A(n6786), .B(n6785), .Z(n7835) );
  XOR U9625 ( .A(n7836), .B(n7835), .Z(n7738) );
  NANDN U9626 ( .A(n6792), .B(n6791), .Z(n6796) );
  NANDN U9627 ( .A(n6794), .B(n6793), .Z(n6795) );
  AND U9628 ( .A(n6796), .B(n6795), .Z(n7980) );
  NANDN U9629 ( .A(n6802), .B(n6801), .Z(n6806) );
  NAND U9630 ( .A(n6804), .B(n6803), .Z(n6805) );
  NAND U9631 ( .A(n6806), .B(n6805), .Z(n8247) );
  NANDN U9632 ( .A(n6808), .B(n6807), .Z(n6812) );
  NANDN U9633 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U9634 ( .A(n6812), .B(n6811), .Z(n8248) );
  XOR U9635 ( .A(n8247), .B(n8248), .Z(n8250) );
  XOR U9636 ( .A(n8249), .B(n8250), .Z(n7979) );
  XOR U9637 ( .A(n7980), .B(n7979), .Z(n7982) );
  NANDN U9638 ( .A(n6814), .B(n6813), .Z(n6818) );
  NANDN U9639 ( .A(n6816), .B(n6815), .Z(n6817) );
  AND U9640 ( .A(n6818), .B(n6817), .Z(n7981) );
  XNOR U9641 ( .A(n7982), .B(n7981), .Z(n7735) );
  XNOR U9642 ( .A(n7736), .B(n7735), .Z(n7737) );
  XOR U9643 ( .A(n7738), .B(n7737), .Z(n7610) );
  XNOR U9644 ( .A(n7609), .B(n7610), .Z(n7695) );
  NANDN U9645 ( .A(n6820), .B(n6819), .Z(n6824) );
  NANDN U9646 ( .A(n6822), .B(n6821), .Z(n6823) );
  NAND U9647 ( .A(n6824), .B(n6823), .Z(n7696) );
  XNOR U9648 ( .A(n7695), .B(n7696), .Z(n7697) );
  NANDN U9649 ( .A(n6826), .B(n6825), .Z(n6830) );
  OR U9650 ( .A(n6828), .B(n6827), .Z(n6829) );
  AND U9651 ( .A(n6830), .B(n6829), .Z(n7539) );
  NANDN U9652 ( .A(n6836), .B(n6835), .Z(n6840) );
  NANDN U9653 ( .A(n6838), .B(n6837), .Z(n6839) );
  AND U9654 ( .A(n6840), .B(n6839), .Z(n7912) );
  NANDN U9655 ( .A(n6842), .B(n6841), .Z(n6846) );
  NANDN U9656 ( .A(n6844), .B(n6843), .Z(n6845) );
  AND U9657 ( .A(n6846), .B(n6845), .Z(n7910) );
  NANDN U9658 ( .A(n6848), .B(n6847), .Z(n6852) );
  NANDN U9659 ( .A(n6850), .B(n6849), .Z(n6851) );
  NAND U9660 ( .A(n6852), .B(n6851), .Z(n8253) );
  NANDN U9661 ( .A(n6858), .B(n6857), .Z(n6862) );
  NAND U9662 ( .A(n6860), .B(n6859), .Z(n6861) );
  NAND U9663 ( .A(n6862), .B(n6861), .Z(n8252) );
  XOR U9664 ( .A(n8251), .B(n8252), .Z(n8254) );
  XOR U9665 ( .A(n8253), .B(n8254), .Z(n7909) );
  XOR U9666 ( .A(n7910), .B(n7909), .Z(n7911) );
  XOR U9667 ( .A(n7912), .B(n7911), .Z(n7706) );
  XNOR U9668 ( .A(n7706), .B(n7705), .Z(n7707) );
  XNOR U9669 ( .A(n7708), .B(n7707), .Z(n7537) );
  XOR U9670 ( .A(n7537), .B(n7538), .Z(n7540) );
  XOR U9671 ( .A(n7539), .B(n7540), .Z(n7698) );
  XNOR U9672 ( .A(n7697), .B(n7698), .Z(n7799) );
  XOR U9673 ( .A(n7800), .B(n7799), .Z(n7801) );
  NANDN U9674 ( .A(n6872), .B(n6871), .Z(n6876) );
  NAND U9675 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U9676 ( .A(n6876), .B(n6875), .Z(n7784) );
  NANDN U9677 ( .A(n6878), .B(n6877), .Z(n6882) );
  NAND U9678 ( .A(n6880), .B(n6879), .Z(n6881) );
  AND U9679 ( .A(n6882), .B(n6881), .Z(n7782) );
  NANDN U9680 ( .A(n6884), .B(n6883), .Z(n6888) );
  OR U9681 ( .A(n6886), .B(n6885), .Z(n6887) );
  AND U9682 ( .A(n6888), .B(n6887), .Z(n7533) );
  NANDN U9683 ( .A(n6890), .B(n6889), .Z(n6894) );
  OR U9684 ( .A(n6892), .B(n6891), .Z(n6893) );
  AND U9685 ( .A(n6894), .B(n6893), .Z(n7531) );
  NANDN U9686 ( .A(n6900), .B(n6899), .Z(n6904) );
  NANDN U9687 ( .A(n6902), .B(n6901), .Z(n6903) );
  AND U9688 ( .A(n6904), .B(n6903), .Z(n8298) );
  NANDN U9689 ( .A(n6918), .B(n6917), .Z(n6922) );
  NAND U9690 ( .A(n6920), .B(n6919), .Z(n6921) );
  NAND U9691 ( .A(n6922), .B(n6921), .Z(n8431) );
  XNOR U9692 ( .A(n8432), .B(n8431), .Z(n8433) );
  XOR U9693 ( .A(n8434), .B(n8433), .Z(n8296) );
  XNOR U9694 ( .A(n8295), .B(n8296), .Z(n8297) );
  XOR U9695 ( .A(n8298), .B(n8297), .Z(n7772) );
  NANDN U9696 ( .A(n6924), .B(n6923), .Z(n6928) );
  NANDN U9697 ( .A(n6926), .B(n6925), .Z(n6927) );
  AND U9698 ( .A(n6928), .B(n6927), .Z(n7771) );
  XOR U9699 ( .A(n7772), .B(n7771), .Z(n7774) );
  XOR U9700 ( .A(n7773), .B(n7774), .Z(n7532) );
  XOR U9701 ( .A(n7531), .B(n7532), .Z(n7534) );
  XNOR U9702 ( .A(n7533), .B(n7534), .Z(n7781) );
  XNOR U9703 ( .A(n7782), .B(n7781), .Z(n7783) );
  XOR U9704 ( .A(n7784), .B(n7783), .Z(n7802) );
  XNOR U9705 ( .A(n7801), .B(n7802), .Z(n7807) );
  XOR U9706 ( .A(n7808), .B(n7807), .Z(n7450) );
  NANDN U9707 ( .A(n6930), .B(n6929), .Z(n6934) );
  NAND U9708 ( .A(n6932), .B(n6931), .Z(n6933) );
  NAND U9709 ( .A(n6934), .B(n6933), .Z(n7449) );
  XNOR U9710 ( .A(n7450), .B(n7449), .Z(n7452) );
  NANDN U9711 ( .A(n6936), .B(n6935), .Z(n6940) );
  OR U9712 ( .A(n6938), .B(n6937), .Z(n6939) );
  AND U9713 ( .A(n6940), .B(n6939), .Z(n7744) );
  NANDN U9714 ( .A(n6942), .B(n6941), .Z(n6946) );
  NANDN U9715 ( .A(n6944), .B(n6943), .Z(n6945) );
  AND U9716 ( .A(n6946), .B(n6945), .Z(n7742) );
  NANDN U9717 ( .A(n6948), .B(n6947), .Z(n6952) );
  NAND U9718 ( .A(n6950), .B(n6949), .Z(n6951) );
  AND U9719 ( .A(n6952), .B(n6951), .Z(n8418) );
  NANDN U9720 ( .A(n6954), .B(n6953), .Z(n6958) );
  NAND U9721 ( .A(n6956), .B(n6955), .Z(n6957) );
  AND U9722 ( .A(n6958), .B(n6957), .Z(n8416) );
  NANDN U9723 ( .A(n6960), .B(n6959), .Z(n6964) );
  NAND U9724 ( .A(n6962), .B(n6961), .Z(n6963) );
  NAND U9725 ( .A(n6964), .B(n6963), .Z(n8415) );
  XNOR U9726 ( .A(n8416), .B(n8415), .Z(n8417) );
  XNOR U9727 ( .A(n8418), .B(n8417), .Z(n7741) );
  XNOR U9728 ( .A(n7742), .B(n7741), .Z(n7743) );
  XOR U9729 ( .A(n7744), .B(n7743), .Z(n8390) );
  NANDN U9730 ( .A(n6966), .B(n6965), .Z(n6970) );
  OR U9731 ( .A(n6968), .B(n6967), .Z(n6969) );
  AND U9732 ( .A(n6970), .B(n6969), .Z(n8506) );
  NANDN U9733 ( .A(n6972), .B(n6971), .Z(n6976) );
  OR U9734 ( .A(n6974), .B(n6973), .Z(n6975) );
  AND U9735 ( .A(n6976), .B(n6975), .Z(n8505) );
  NANDN U9736 ( .A(n6978), .B(n6977), .Z(n6982) );
  NAND U9737 ( .A(n6980), .B(n6979), .Z(n6981) );
  AND U9738 ( .A(n6982), .B(n6981), .Z(n7762) );
  NANDN U9739 ( .A(n6984), .B(n6983), .Z(n6988) );
  NAND U9740 ( .A(n6986), .B(n6985), .Z(n6987) );
  AND U9741 ( .A(n6988), .B(n6987), .Z(n7760) );
  NANDN U9742 ( .A(n6990), .B(n6989), .Z(n6994) );
  NANDN U9743 ( .A(n6992), .B(n6991), .Z(n6993) );
  NAND U9744 ( .A(n6994), .B(n6993), .Z(n7759) );
  XNOR U9745 ( .A(n7760), .B(n7759), .Z(n7761) );
  XNOR U9746 ( .A(n7762), .B(n7761), .Z(n8504) );
  XOR U9747 ( .A(n8505), .B(n8504), .Z(n8507) );
  XOR U9748 ( .A(n8506), .B(n8507), .Z(n8388) );
  NANDN U9749 ( .A(n7000), .B(n6999), .Z(n7004) );
  OR U9750 ( .A(n7002), .B(n7001), .Z(n7003) );
  AND U9751 ( .A(n7004), .B(n7003), .Z(n7525) );
  NANDN U9752 ( .A(n7006), .B(n7005), .Z(n7010) );
  NAND U9753 ( .A(n7008), .B(n7007), .Z(n7009) );
  AND U9754 ( .A(n7010), .B(n7009), .Z(n7756) );
  NANDN U9755 ( .A(n7012), .B(n7011), .Z(n7016) );
  NAND U9756 ( .A(n7014), .B(n7013), .Z(n7015) );
  AND U9757 ( .A(n7016), .B(n7015), .Z(n7754) );
  NANDN U9758 ( .A(n7018), .B(n7017), .Z(n7022) );
  NAND U9759 ( .A(n7020), .B(n7019), .Z(n7021) );
  NAND U9760 ( .A(n7022), .B(n7021), .Z(n7753) );
  XNOR U9761 ( .A(n7754), .B(n7753), .Z(n7755) );
  XOR U9762 ( .A(n7756), .B(n7755), .Z(n7526) );
  XOR U9763 ( .A(n7525), .B(n7526), .Z(n7528) );
  XNOR U9764 ( .A(n7527), .B(n7528), .Z(n8387) );
  XOR U9765 ( .A(n7692), .B(n7691), .Z(n7694) );
  NANDN U9766 ( .A(n7028), .B(n7027), .Z(n7032) );
  NANDN U9767 ( .A(n7030), .B(n7029), .Z(n7031) );
  AND U9768 ( .A(n7032), .B(n7031), .Z(n8513) );
  NANDN U9769 ( .A(n7034), .B(n7033), .Z(n7038) );
  OR U9770 ( .A(n7036), .B(n7035), .Z(n7037) );
  AND U9771 ( .A(n7038), .B(n7037), .Z(n8511) );
  NANDN U9772 ( .A(n7040), .B(n7039), .Z(n7044) );
  NAND U9773 ( .A(n7042), .B(n7041), .Z(n7043) );
  AND U9774 ( .A(n7044), .B(n7043), .Z(n7704) );
  NANDN U9775 ( .A(n7046), .B(n7045), .Z(n7050) );
  NAND U9776 ( .A(n7048), .B(n7047), .Z(n7049) );
  NAND U9777 ( .A(n7050), .B(n7049), .Z(n8413) );
  NANDN U9778 ( .A(n7052), .B(n7051), .Z(n7056) );
  NAND U9779 ( .A(n7054), .B(n7053), .Z(n7055) );
  NAND U9780 ( .A(n7056), .B(n7055), .Z(n8411) );
  XNOR U9781 ( .A(n8411), .B(n8412), .Z(n8414) );
  XOR U9782 ( .A(n8413), .B(n8414), .Z(n7701) );
  NANDN U9783 ( .A(n7062), .B(n7061), .Z(n7066) );
  NAND U9784 ( .A(n7064), .B(n7063), .Z(n7065) );
  NAND U9785 ( .A(n7066), .B(n7065), .Z(n7702) );
  XOR U9786 ( .A(n7701), .B(n7702), .Z(n7703) );
  XOR U9787 ( .A(n7704), .B(n7703), .Z(n8510) );
  XOR U9788 ( .A(n8513), .B(n8512), .Z(n7693) );
  XOR U9789 ( .A(n7694), .B(n7693), .Z(n8378) );
  NANDN U9790 ( .A(n7068), .B(n7067), .Z(n7072) );
  NANDN U9791 ( .A(n7070), .B(n7069), .Z(n7071) );
  AND U9792 ( .A(n7072), .B(n7071), .Z(n8400) );
  NAND U9793 ( .A(n7078), .B(n7077), .Z(n7082) );
  NAND U9794 ( .A(n7080), .B(n7079), .Z(n7081) );
  AND U9795 ( .A(n7082), .B(n7081), .Z(n7885) );
  XOR U9796 ( .A(n8037), .B(n8038), .Z(n8040) );
  XOR U9797 ( .A(n8039), .B(n8040), .Z(n7886) );
  XNOR U9798 ( .A(n7885), .B(n7886), .Z(n7887) );
  XOR U9799 ( .A(n8077), .B(n8078), .Z(n8080) );
  XOR U9800 ( .A(n8079), .B(n8080), .Z(n7888) );
  XOR U9801 ( .A(n7887), .B(n7888), .Z(n7812) );
  XNOR U9802 ( .A(n7811), .B(n7812), .Z(n7813) );
  NANDN U9803 ( .A(n7108), .B(n7107), .Z(n7112) );
  NANDN U9804 ( .A(n7110), .B(n7109), .Z(n7111) );
  NAND U9805 ( .A(n7112), .B(n7111), .Z(n7814) );
  XNOR U9806 ( .A(n7813), .B(n7814), .Z(n8399) );
  XOR U9807 ( .A(n8402), .B(n8401), .Z(n7688) );
  NANDN U9808 ( .A(n7118), .B(n7117), .Z(n7122) );
  NAND U9809 ( .A(n7120), .B(n7119), .Z(n7121) );
  NAND U9810 ( .A(n7122), .B(n7121), .Z(n8351) );
  NANDN U9811 ( .A(n7124), .B(n7123), .Z(n7128) );
  NANDN U9812 ( .A(n7126), .B(n7125), .Z(n7127) );
  AND U9813 ( .A(n7128), .B(n7127), .Z(n8158) );
  NANDN U9814 ( .A(n7130), .B(n7129), .Z(n7134) );
  NANDN U9815 ( .A(n7132), .B(n7131), .Z(n7133) );
  AND U9816 ( .A(n7134), .B(n7133), .Z(n8155) );
  XNOR U9817 ( .A(n8180), .B(n8179), .Z(n8181) );
  XOR U9818 ( .A(n8182), .B(n8181), .Z(n8156) );
  XNOR U9819 ( .A(n8155), .B(n8156), .Z(n8157) );
  XOR U9820 ( .A(n8158), .B(n8157), .Z(n7952) );
  NANDN U9821 ( .A(n7148), .B(n7147), .Z(n7152) );
  NANDN U9822 ( .A(n7150), .B(n7149), .Z(n7151) );
  AND U9823 ( .A(n7152), .B(n7151), .Z(n7976) );
  NANDN U9824 ( .A(n7154), .B(n7153), .Z(n7158) );
  NANDN U9825 ( .A(n7156), .B(n7155), .Z(n7157) );
  AND U9826 ( .A(n7158), .B(n7157), .Z(n7973) );
  NANDN U9827 ( .A(n7160), .B(n7159), .Z(n7164) );
  NANDN U9828 ( .A(n7162), .B(n7161), .Z(n7163) );
  NAND U9829 ( .A(n7164), .B(n7163), .Z(n7974) );
  XNOR U9830 ( .A(n7973), .B(n7974), .Z(n7975) );
  XOR U9831 ( .A(n7976), .B(n7975), .Z(n7950) );
  NANDN U9832 ( .A(n7166), .B(n7165), .Z(n7170) );
  NANDN U9833 ( .A(n7168), .B(n7167), .Z(n7169) );
  AND U9834 ( .A(n7170), .B(n7169), .Z(n8136) );
  NANDN U9835 ( .A(n7172), .B(n7171), .Z(n7176) );
  OR U9836 ( .A(n7174), .B(n7173), .Z(n7175) );
  AND U9837 ( .A(n7176), .B(n7175), .Z(n8133) );
  NANDN U9838 ( .A(n7178), .B(n7177), .Z(n7182) );
  NANDN U9839 ( .A(n7180), .B(n7179), .Z(n7181) );
  NAND U9840 ( .A(n7182), .B(n7181), .Z(n8134) );
  XNOR U9841 ( .A(n8133), .B(n8134), .Z(n8135) );
  XNOR U9842 ( .A(n8136), .B(n8135), .Z(n7949) );
  XNOR U9843 ( .A(n7950), .B(n7949), .Z(n7951) );
  XNOR U9844 ( .A(n7952), .B(n7951), .Z(n8352) );
  XOR U9845 ( .A(n8351), .B(n8352), .Z(n8354) );
  NANDN U9846 ( .A(n7188), .B(n7187), .Z(n7192) );
  NAND U9847 ( .A(n7190), .B(n7189), .Z(n7191) );
  AND U9848 ( .A(n7192), .B(n7191), .Z(n8334) );
  NANDN U9849 ( .A(n7194), .B(n7193), .Z(n7198) );
  OR U9850 ( .A(n7196), .B(n7195), .Z(n7197) );
  AND U9851 ( .A(n7198), .B(n7197), .Z(n7916) );
  NANDN U9852 ( .A(n7200), .B(n7199), .Z(n7204) );
  NANDN U9853 ( .A(n7202), .B(n7201), .Z(n7203) );
  AND U9854 ( .A(n7204), .B(n7203), .Z(n7913) );
  NANDN U9855 ( .A(n7206), .B(n7205), .Z(n7210) );
  NANDN U9856 ( .A(n7208), .B(n7207), .Z(n7209) );
  NAND U9857 ( .A(n7210), .B(n7209), .Z(n7914) );
  XNOR U9858 ( .A(n7913), .B(n7914), .Z(n7915) );
  XNOR U9859 ( .A(n7916), .B(n7915), .Z(n8333) );
  XNOR U9860 ( .A(n8334), .B(n8333), .Z(n8335) );
  XNOR U9861 ( .A(n8336), .B(n8335), .Z(n8353) );
  XOR U9862 ( .A(n8354), .B(n8353), .Z(n7864) );
  NANDN U9863 ( .A(n7212), .B(n7211), .Z(n7216) );
  OR U9864 ( .A(n7214), .B(n7213), .Z(n7215) );
  AND U9865 ( .A(n7216), .B(n7215), .Z(n7875) );
  NANDN U9866 ( .A(n7218), .B(n7217), .Z(n7222) );
  NANDN U9867 ( .A(n7220), .B(n7219), .Z(n7221) );
  AND U9868 ( .A(n7222), .B(n7221), .Z(n7873) );
  NANDN U9869 ( .A(n7224), .B(n7223), .Z(n7228) );
  OR U9870 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U9871 ( .A(n7228), .B(n7227), .Z(n8482) );
  NANDN U9872 ( .A(n7230), .B(n7229), .Z(n7234) );
  NANDN U9873 ( .A(n7232), .B(n7231), .Z(n7233) );
  AND U9874 ( .A(n7234), .B(n7233), .Z(n8480) );
  NANDN U9875 ( .A(n7236), .B(n7235), .Z(n7240) );
  NANDN U9876 ( .A(n7238), .B(n7237), .Z(n7239) );
  NAND U9877 ( .A(n7240), .B(n7239), .Z(n8481) );
  XOR U9878 ( .A(n8480), .B(n8481), .Z(n8483) );
  XOR U9879 ( .A(n8482), .B(n8483), .Z(n7874) );
  XOR U9880 ( .A(n7873), .B(n7874), .Z(n7876) );
  XOR U9881 ( .A(n7875), .B(n7876), .Z(n7851) );
  NANDN U9882 ( .A(n7242), .B(n7241), .Z(n7246) );
  NANDN U9883 ( .A(n7244), .B(n7243), .Z(n7245) );
  AND U9884 ( .A(n7246), .B(n7245), .Z(n7970) );
  NANDN U9885 ( .A(n7248), .B(n7247), .Z(n7252) );
  NAND U9886 ( .A(n7250), .B(n7249), .Z(n7251) );
  NAND U9887 ( .A(n7252), .B(n7251), .Z(n7587) );
  NANDN U9888 ( .A(n7254), .B(n7253), .Z(n7258) );
  NANDN U9889 ( .A(n7256), .B(n7255), .Z(n7257) );
  NAND U9890 ( .A(n7258), .B(n7257), .Z(n7585) );
  XOR U9891 ( .A(n7585), .B(n7586), .Z(n7588) );
  XOR U9892 ( .A(n7587), .B(n7588), .Z(n7969) );
  XOR U9893 ( .A(n7970), .B(n7969), .Z(n7972) );
  XOR U9894 ( .A(n7972), .B(n7971), .Z(n7946) );
  NANDN U9895 ( .A(n7268), .B(n7267), .Z(n7272) );
  NANDN U9896 ( .A(n7270), .B(n7269), .Z(n7271) );
  AND U9897 ( .A(n7272), .B(n7271), .Z(n7665) );
  NANDN U9898 ( .A(n7274), .B(n7273), .Z(n7278) );
  NAND U9899 ( .A(n7276), .B(n7275), .Z(n7277) );
  AND U9900 ( .A(n7278), .B(n7277), .Z(n7496) );
  NANDN U9901 ( .A(n7280), .B(n7279), .Z(n7284) );
  NANDN U9902 ( .A(n7282), .B(n7281), .Z(n7283) );
  AND U9903 ( .A(n7284), .B(n7283), .Z(n7494) );
  NANDN U9904 ( .A(n7286), .B(n7285), .Z(n7290) );
  NAND U9905 ( .A(n7288), .B(n7287), .Z(n7289) );
  NAND U9906 ( .A(n7290), .B(n7289), .Z(n7493) );
  XNOR U9907 ( .A(n7494), .B(n7493), .Z(n7495) );
  XOR U9908 ( .A(n7496), .B(n7495), .Z(n7666) );
  XNOR U9909 ( .A(n7665), .B(n7666), .Z(n7668) );
  NANDN U9910 ( .A(n7296), .B(n7295), .Z(n7300) );
  NANDN U9911 ( .A(n7298), .B(n7297), .Z(n7299) );
  AND U9912 ( .A(n7300), .B(n7299), .Z(n7482) );
  XNOR U9913 ( .A(n7482), .B(n7481), .Z(n7483) );
  XNOR U9914 ( .A(n7484), .B(n7483), .Z(n7667) );
  XOR U9915 ( .A(n7668), .B(n7667), .Z(n7944) );
  NANDN U9916 ( .A(n7306), .B(n7305), .Z(n7310) );
  NANDN U9917 ( .A(n7308), .B(n7307), .Z(n7309) );
  AND U9918 ( .A(n7310), .B(n7309), .Z(n8464) );
  NANDN U9919 ( .A(n7320), .B(n7319), .Z(n7324) );
  NANDN U9920 ( .A(n7322), .B(n7321), .Z(n7323) );
  NAND U9921 ( .A(n7324), .B(n7323), .Z(n7487) );
  XNOR U9922 ( .A(n7488), .B(n7487), .Z(n7489) );
  XOR U9923 ( .A(n7490), .B(n7489), .Z(n8465) );
  XNOR U9924 ( .A(n8464), .B(n8465), .Z(n8467) );
  NANDN U9925 ( .A(n7334), .B(n7333), .Z(n7338) );
  NAND U9926 ( .A(n7336), .B(n7335), .Z(n7337) );
  NAND U9927 ( .A(n7338), .B(n7337), .Z(n8025) );
  XNOR U9928 ( .A(n8026), .B(n8025), .Z(n8027) );
  XNOR U9929 ( .A(n8028), .B(n8027), .Z(n8466) );
  XNOR U9930 ( .A(n8467), .B(n8466), .Z(n7943) );
  XNOR U9931 ( .A(n7944), .B(n7943), .Z(n7945) );
  XNOR U9932 ( .A(n7946), .B(n7945), .Z(n7849) );
  NANDN U9933 ( .A(n7340), .B(n7339), .Z(n7344) );
  NANDN U9934 ( .A(n7342), .B(n7341), .Z(n7343) );
  AND U9935 ( .A(n7344), .B(n7343), .Z(n8096) );
  NANDN U9936 ( .A(n7346), .B(n7345), .Z(n7350) );
  NANDN U9937 ( .A(n7348), .B(n7347), .Z(n7349) );
  AND U9938 ( .A(n7350), .B(n7349), .Z(n7508) );
  NANDN U9939 ( .A(n7352), .B(n7351), .Z(n7356) );
  NANDN U9940 ( .A(n7354), .B(n7353), .Z(n7355) );
  AND U9941 ( .A(n7356), .B(n7355), .Z(n7506) );
  NANDN U9942 ( .A(n7358), .B(n7357), .Z(n7362) );
  NANDN U9943 ( .A(n7360), .B(n7359), .Z(n7361) );
  AND U9944 ( .A(n7362), .B(n7361), .Z(n7505) );
  XOR U9945 ( .A(n7506), .B(n7505), .Z(n7507) );
  XOR U9946 ( .A(n7508), .B(n7507), .Z(n8094) );
  XNOR U9947 ( .A(n8094), .B(n8093), .Z(n8095) );
  XOR U9948 ( .A(n8096), .B(n8095), .Z(n7850) );
  XOR U9949 ( .A(n7849), .B(n7850), .Z(n7852) );
  XOR U9950 ( .A(n7851), .B(n7852), .Z(n7862) );
  XOR U9951 ( .A(n8278), .B(n8277), .Z(n8280) );
  XOR U9952 ( .A(n8280), .B(n8279), .Z(n8342) );
  NANDN U9953 ( .A(n7380), .B(n7379), .Z(n7384) );
  NAND U9954 ( .A(n7382), .B(n7381), .Z(n7383) );
  AND U9955 ( .A(n7384), .B(n7383), .Z(n8340) );
  NANDN U9956 ( .A(n7386), .B(n7385), .Z(n7390) );
  NANDN U9957 ( .A(n7388), .B(n7387), .Z(n7389) );
  AND U9958 ( .A(n7390), .B(n7389), .Z(n7906) );
  NANDN U9959 ( .A(n7392), .B(n7391), .Z(n7396) );
  NANDN U9960 ( .A(n7394), .B(n7393), .Z(n7395) );
  AND U9961 ( .A(n7396), .B(n7395), .Z(n7904) );
  NANDN U9962 ( .A(n7398), .B(n7397), .Z(n7402) );
  NANDN U9963 ( .A(n7400), .B(n7399), .Z(n7401) );
  NAND U9964 ( .A(n7402), .B(n7401), .Z(n7903) );
  XNOR U9965 ( .A(n7904), .B(n7903), .Z(n7905) );
  XNOR U9966 ( .A(n7906), .B(n7905), .Z(n8339) );
  XNOR U9967 ( .A(n8340), .B(n8339), .Z(n8341) );
  XOR U9968 ( .A(n8342), .B(n8341), .Z(n8347) );
  NANDN U9969 ( .A(n7404), .B(n7403), .Z(n7408) );
  NANDN U9970 ( .A(n7406), .B(n7405), .Z(n7407) );
  NAND U9971 ( .A(n7408), .B(n7407), .Z(n8345) );
  NANDN U9972 ( .A(n7410), .B(n7409), .Z(n7414) );
  NAND U9973 ( .A(n7412), .B(n7411), .Z(n7413) );
  AND U9974 ( .A(n7414), .B(n7413), .Z(n7879) );
  NANDN U9975 ( .A(n7416), .B(n7415), .Z(n7420) );
  NANDN U9976 ( .A(n7418), .B(n7417), .Z(n7419) );
  AND U9977 ( .A(n7420), .B(n7419), .Z(n8045) );
  NANDN U9978 ( .A(n7426), .B(n7425), .Z(n7430) );
  NANDN U9979 ( .A(n7428), .B(n7427), .Z(n7429) );
  NAND U9980 ( .A(n7430), .B(n7429), .Z(n8044) );
  XOR U9981 ( .A(n8043), .B(n8044), .Z(n8046) );
  XOR U9982 ( .A(n8045), .B(n8046), .Z(n7880) );
  XNOR U9983 ( .A(n7879), .B(n7880), .Z(n7881) );
  NANDN U9984 ( .A(n7432), .B(n7431), .Z(n7436) );
  NAND U9985 ( .A(n7434), .B(n7433), .Z(n7435) );
  NAND U9986 ( .A(n7436), .B(n7435), .Z(n7882) );
  XNOR U9987 ( .A(n7881), .B(n7882), .Z(n8346) );
  XOR U9988 ( .A(n8345), .B(n8346), .Z(n8348) );
  XOR U9989 ( .A(n8347), .B(n8348), .Z(n7861) );
  NANDN U9990 ( .A(n7438), .B(n7437), .Z(n7442) );
  NANDN U9991 ( .A(n7440), .B(n7439), .Z(n7441) );
  AND U9992 ( .A(n7442), .B(n7441), .Z(n7685) );
  XOR U9993 ( .A(n7686), .B(n7685), .Z(n7687) );
  XOR U9994 ( .A(n7688), .B(n7687), .Z(n8375) );
  NAND U9995 ( .A(n7444), .B(n7443), .Z(n7448) );
  NAND U9996 ( .A(n7446), .B(n7445), .Z(n7447) );
  AND U9997 ( .A(n7448), .B(n7447), .Z(n8376) );
  XOR U9998 ( .A(n8375), .B(n8376), .Z(n8377) );
  XNOR U9999 ( .A(n7452), .B(n7451), .Z(o[2]) );
  NANDN U10000 ( .A(n7450), .B(n7449), .Z(n7454) );
  NAND U10001 ( .A(n7452), .B(n7451), .Z(n7453) );
  AND U10002 ( .A(n7454), .B(n7453), .Z(n9056) );
  NANDN U10003 ( .A(n7456), .B(n7455), .Z(n7460) );
  NAND U10004 ( .A(n7458), .B(n7457), .Z(n7459) );
  AND U10005 ( .A(n7460), .B(n7459), .Z(n8845) );
  NANDN U10006 ( .A(n7462), .B(n7461), .Z(n7466) );
  NANDN U10007 ( .A(n7464), .B(n7463), .Z(n7465) );
  AND U10008 ( .A(n7466), .B(n7465), .Z(n9021) );
  XOR U10009 ( .A(n9021), .B(n9020), .Z(n9023) );
  XOR U10010 ( .A(n9023), .B(n9022), .Z(n8554) );
  NANDN U10011 ( .A(n7476), .B(n7475), .Z(n7480) );
  NAND U10012 ( .A(n7478), .B(n7477), .Z(n7479) );
  AND U10013 ( .A(n7480), .B(n7479), .Z(n8553) );
  NANDN U10014 ( .A(n7482), .B(n7481), .Z(n7486) );
  NANDN U10015 ( .A(n7484), .B(n7483), .Z(n7485) );
  AND U10016 ( .A(n7486), .B(n7485), .Z(n9027) );
  NANDN U10017 ( .A(n7488), .B(n7487), .Z(n7492) );
  NANDN U10018 ( .A(n7490), .B(n7489), .Z(n7491) );
  AND U10019 ( .A(n7492), .B(n7491), .Z(n9025) );
  NANDN U10020 ( .A(n7494), .B(n7493), .Z(n7498) );
  NANDN U10021 ( .A(n7496), .B(n7495), .Z(n7497) );
  AND U10022 ( .A(n7498), .B(n7497), .Z(n9024) );
  XOR U10023 ( .A(n9025), .B(n9024), .Z(n9026) );
  XNOR U10024 ( .A(n9027), .B(n9026), .Z(n8552) );
  XOR U10025 ( .A(n8553), .B(n8552), .Z(n8555) );
  XOR U10026 ( .A(n8554), .B(n8555), .Z(n8753) );
  NANDN U10027 ( .A(n7500), .B(n7499), .Z(n7504) );
  NANDN U10028 ( .A(n7502), .B(n7501), .Z(n7503) );
  NAND U10029 ( .A(n7504), .B(n7503), .Z(n8998) );
  XOR U10030 ( .A(n8961), .B(n8960), .Z(n8963) );
  XOR U10031 ( .A(n8963), .B(n8962), .Z(n8997) );
  XOR U10032 ( .A(n8996), .B(n8997), .Z(n8999) );
  XOR U10033 ( .A(n8998), .B(n8999), .Z(n8750) );
  XOR U10034 ( .A(n8750), .B(n8751), .Z(n8752) );
  XOR U10035 ( .A(n8753), .B(n8752), .Z(n8842) );
  NANDN U10036 ( .A(n7526), .B(n7525), .Z(n7530) );
  OR U10037 ( .A(n7528), .B(n7527), .Z(n7529) );
  AND U10038 ( .A(n7530), .B(n7529), .Z(n8843) );
  XOR U10039 ( .A(n8842), .B(n8843), .Z(n8844) );
  XOR U10040 ( .A(n8845), .B(n8844), .Z(n8541) );
  NANDN U10041 ( .A(n7532), .B(n7531), .Z(n7536) );
  NANDN U10042 ( .A(n7534), .B(n7533), .Z(n7535) );
  AND U10043 ( .A(n7536), .B(n7535), .Z(n8879) );
  NANDN U10044 ( .A(n7538), .B(n7537), .Z(n7542) );
  NANDN U10045 ( .A(n7540), .B(n7539), .Z(n7541) );
  AND U10046 ( .A(n7542), .B(n7541), .Z(n8877) );
  NANDN U10047 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U10048 ( .A(n7550), .B(n7549), .Z(n7551) );
  NAND U10049 ( .A(n7552), .B(n7551), .Z(n8571) );
  XNOR U10050 ( .A(n8570), .B(n8571), .Z(n8573) );
  XOR U10051 ( .A(n8573), .B(n8572), .Z(n8596) );
  NANDN U10052 ( .A(n7558), .B(n7557), .Z(n7562) );
  NAND U10053 ( .A(n7560), .B(n7559), .Z(n7561) );
  AND U10054 ( .A(n7562), .B(n7561), .Z(n8595) );
  XOR U10055 ( .A(n9029), .B(n9028), .Z(n9032) );
  XNOR U10056 ( .A(n9032), .B(n9031), .Z(n8594) );
  XOR U10057 ( .A(n8595), .B(n8594), .Z(n8597) );
  XOR U10058 ( .A(n8596), .B(n8597), .Z(n8757) );
  NANDN U10059 ( .A(n7580), .B(n7579), .Z(n7584) );
  NAND U10060 ( .A(n7582), .B(n7581), .Z(n7583) );
  AND U10061 ( .A(n7584), .B(n7583), .Z(n8589) );
  NANDN U10062 ( .A(n7590), .B(n7589), .Z(n7594) );
  NANDN U10063 ( .A(n7592), .B(n7591), .Z(n7593) );
  AND U10064 ( .A(n7594), .B(n7593), .Z(n8952) );
  XOR U10065 ( .A(n8953), .B(n8952), .Z(n8955) );
  NANDN U10066 ( .A(n7596), .B(n7595), .Z(n7600) );
  NANDN U10067 ( .A(n7598), .B(n7597), .Z(n7599) );
  AND U10068 ( .A(n7600), .B(n7599), .Z(n8954) );
  XNOR U10069 ( .A(n8955), .B(n8954), .Z(n8588) );
  XOR U10070 ( .A(n8589), .B(n8588), .Z(n8591) );
  XOR U10071 ( .A(n8590), .B(n8591), .Z(n8755) );
  NANDN U10072 ( .A(n7602), .B(n7601), .Z(n7606) );
  NANDN U10073 ( .A(n7604), .B(n7603), .Z(n7605) );
  AND U10074 ( .A(n7606), .B(n7605), .Z(n8754) );
  XNOR U10075 ( .A(n8755), .B(n8754), .Z(n8756) );
  XNOR U10076 ( .A(n8757), .B(n8756), .Z(n8876) );
  XNOR U10077 ( .A(n8877), .B(n8876), .Z(n8878) );
  XNOR U10078 ( .A(n8879), .B(n8878), .Z(n8540) );
  XNOR U10079 ( .A(n8541), .B(n8540), .Z(n8542) );
  NANDN U10080 ( .A(n7608), .B(n7607), .Z(n7612) );
  NANDN U10081 ( .A(n7610), .B(n7609), .Z(n7611) );
  AND U10082 ( .A(n7612), .B(n7611), .Z(n8731) );
  NANDN U10083 ( .A(n7618), .B(n7617), .Z(n7622) );
  NANDN U10084 ( .A(n7620), .B(n7619), .Z(n7621) );
  AND U10085 ( .A(n7622), .B(n7621), .Z(n8800) );
  NANDN U10086 ( .A(n7624), .B(n7623), .Z(n7628) );
  NANDN U10087 ( .A(n7626), .B(n7625), .Z(n7627) );
  NAND U10088 ( .A(n7628), .B(n7627), .Z(n8801) );
  XNOR U10089 ( .A(n8800), .B(n8801), .Z(n8802) );
  XOR U10090 ( .A(n8802), .B(n8803), .Z(n8938) );
  XNOR U10091 ( .A(n8576), .B(n8577), .Z(n8578) );
  NANDN U10092 ( .A(n7642), .B(n7641), .Z(n7646) );
  NANDN U10093 ( .A(n7644), .B(n7643), .Z(n7645) );
  NAND U10094 ( .A(n7646), .B(n7645), .Z(n8579) );
  XOR U10095 ( .A(n8578), .B(n8579), .Z(n8936) );
  NANDN U10096 ( .A(n7648), .B(n7647), .Z(n7652) );
  NAND U10097 ( .A(n7650), .B(n7649), .Z(n7651) );
  NAND U10098 ( .A(n7652), .B(n7651), .Z(n8937) );
  XOR U10099 ( .A(n8936), .B(n8937), .Z(n8939) );
  XOR U10100 ( .A(n8938), .B(n8939), .Z(n8933) );
  NANDN U10101 ( .A(n7654), .B(n7653), .Z(n7658) );
  OR U10102 ( .A(n7656), .B(n7655), .Z(n7657) );
  AND U10103 ( .A(n7658), .B(n7657), .Z(n8932) );
  XOR U10104 ( .A(n8933), .B(n8932), .Z(n8935) );
  NANDN U10105 ( .A(n7660), .B(n7659), .Z(n7664) );
  NAND U10106 ( .A(n7662), .B(n7661), .Z(n7663) );
  NAND U10107 ( .A(n7664), .B(n7663), .Z(n8950) );
  NANDN U10108 ( .A(n7666), .B(n7665), .Z(n7670) );
  NAND U10109 ( .A(n7668), .B(n7667), .Z(n7669) );
  NAND U10110 ( .A(n7670), .B(n7669), .Z(n8948) );
  NANDN U10111 ( .A(n7672), .B(n7671), .Z(n7676) );
  NANDN U10112 ( .A(n7674), .B(n7673), .Z(n7675) );
  AND U10113 ( .A(n7676), .B(n7675), .Z(n8812) );
  XNOR U10114 ( .A(n8812), .B(n8813), .Z(n8815) );
  XNOR U10115 ( .A(n8815), .B(n8814), .Z(n8949) );
  XOR U10116 ( .A(n8948), .B(n8949), .Z(n8951) );
  XOR U10117 ( .A(n8950), .B(n8951), .Z(n8934) );
  XNOR U10118 ( .A(n8935), .B(n8934), .Z(n8728) );
  XNOR U10119 ( .A(n8729), .B(n8728), .Z(n8730) );
  XOR U10120 ( .A(n8731), .B(n8730), .Z(n8543) );
  XNOR U10121 ( .A(n8542), .B(n8543), .Z(n8673) );
  NAND U10122 ( .A(n7686), .B(n7685), .Z(n7690) );
  NANDN U10123 ( .A(n7688), .B(n7687), .Z(n7689) );
  AND U10124 ( .A(n7690), .B(n7689), .Z(n8671) );
  XNOR U10125 ( .A(n8671), .B(n8670), .Z(n8672) );
  XOR U10126 ( .A(n8673), .B(n8672), .Z(n8529) );
  NANDN U10127 ( .A(n7696), .B(n7695), .Z(n7700) );
  NANDN U10128 ( .A(n7698), .B(n7697), .Z(n7699) );
  AND U10129 ( .A(n7700), .B(n7699), .Z(n8761) );
  NANDN U10130 ( .A(n7706), .B(n7705), .Z(n7710) );
  NANDN U10131 ( .A(n7708), .B(n7707), .Z(n7709) );
  AND U10132 ( .A(n7710), .B(n7709), .Z(n8891) );
  NANDN U10133 ( .A(n7712), .B(n7711), .Z(n7716) );
  NAND U10134 ( .A(n7714), .B(n7713), .Z(n7715) );
  NAND U10135 ( .A(n7716), .B(n7715), .Z(n8888) );
  NANDN U10136 ( .A(n7718), .B(n7717), .Z(n7722) );
  NANDN U10137 ( .A(n7720), .B(n7719), .Z(n7721) );
  AND U10138 ( .A(n7722), .B(n7721), .Z(n8889) );
  XOR U10139 ( .A(n8888), .B(n8889), .Z(n8890) );
  XOR U10140 ( .A(n8891), .B(n8890), .Z(n8723) );
  NANDN U10141 ( .A(n7724), .B(n7723), .Z(n7728) );
  OR U10142 ( .A(n7726), .B(n7725), .Z(n7727) );
  NAND U10143 ( .A(n7728), .B(n7727), .Z(n8702) );
  NANDN U10144 ( .A(n7730), .B(n7729), .Z(n7734) );
  NANDN U10145 ( .A(n7732), .B(n7731), .Z(n7733) );
  NAND U10146 ( .A(n7734), .B(n7733), .Z(n8700) );
  NANDN U10147 ( .A(n7736), .B(n7735), .Z(n7740) );
  NANDN U10148 ( .A(n7738), .B(n7737), .Z(n7739) );
  NAND U10149 ( .A(n7740), .B(n7739), .Z(n8701) );
  XOR U10150 ( .A(n8700), .B(n8701), .Z(n8703) );
  XOR U10151 ( .A(n8702), .B(n8703), .Z(n8722) );
  XOR U10152 ( .A(n8723), .B(n8722), .Z(n8725) );
  XNOR U10153 ( .A(n8724), .B(n8725), .Z(n8760) );
  NANDN U10154 ( .A(n7742), .B(n7741), .Z(n7746) );
  NAND U10155 ( .A(n7744), .B(n7743), .Z(n7745) );
  AND U10156 ( .A(n7746), .B(n7745), .Z(n8855) );
  NANDN U10157 ( .A(n7748), .B(n7747), .Z(n7752) );
  OR U10158 ( .A(n7750), .B(n7749), .Z(n7751) );
  AND U10159 ( .A(n7752), .B(n7751), .Z(n8710) );
  NANDN U10160 ( .A(n7754), .B(n7753), .Z(n7758) );
  NANDN U10161 ( .A(n7756), .B(n7755), .Z(n7757) );
  NAND U10162 ( .A(n7758), .B(n7757), .Z(n8711) );
  XNOR U10163 ( .A(n8710), .B(n8711), .Z(n8713) );
  NANDN U10164 ( .A(n7760), .B(n7759), .Z(n7764) );
  NANDN U10165 ( .A(n7762), .B(n7761), .Z(n7763) );
  AND U10166 ( .A(n7764), .B(n7763), .Z(n8712) );
  XOR U10167 ( .A(n8713), .B(n8712), .Z(n8853) );
  NANDN U10168 ( .A(n7766), .B(n7765), .Z(n7770) );
  OR U10169 ( .A(n7768), .B(n7767), .Z(n7769) );
  AND U10170 ( .A(n7770), .B(n7769), .Z(n8882) );
  NANDN U10171 ( .A(n7772), .B(n7771), .Z(n7776) );
  NANDN U10172 ( .A(n7774), .B(n7773), .Z(n7775) );
  NAND U10173 ( .A(n7776), .B(n7775), .Z(n8883) );
  XNOR U10174 ( .A(n8882), .B(n8883), .Z(n8885) );
  XNOR U10175 ( .A(n8885), .B(n8884), .Z(n8852) );
  XNOR U10176 ( .A(n8853), .B(n8852), .Z(n8854) );
  XNOR U10177 ( .A(n8855), .B(n8854), .Z(n8762) );
  XOR U10178 ( .A(n8763), .B(n8762), .Z(n8537) );
  NANDN U10179 ( .A(n7782), .B(n7781), .Z(n7786) );
  NANDN U10180 ( .A(n7784), .B(n7783), .Z(n7785) );
  AND U10181 ( .A(n7786), .B(n7785), .Z(n8683) );
  NANDN U10182 ( .A(n7788), .B(n7787), .Z(n7792) );
  NAND U10183 ( .A(n7790), .B(n7789), .Z(n7791) );
  AND U10184 ( .A(n7792), .B(n7791), .Z(n8682) );
  NANDN U10185 ( .A(n7794), .B(n7793), .Z(n7798) );
  OR U10186 ( .A(n7796), .B(n7795), .Z(n7797) );
  AND U10187 ( .A(n7798), .B(n7797), .Z(n8684) );
  XOR U10188 ( .A(n8685), .B(n8684), .Z(n8535) );
  NAND U10189 ( .A(n7800), .B(n7799), .Z(n7804) );
  NANDN U10190 ( .A(n7802), .B(n7801), .Z(n7803) );
  AND U10191 ( .A(n7804), .B(n7803), .Z(n8534) );
  XNOR U10192 ( .A(n8535), .B(n8534), .Z(n8536) );
  XNOR U10193 ( .A(n8537), .B(n8536), .Z(n8528) );
  NAND U10194 ( .A(n7806), .B(n7805), .Z(n7810) );
  NAND U10195 ( .A(n7808), .B(n7807), .Z(n7809) );
  AND U10196 ( .A(n7810), .B(n7809), .Z(n8530) );
  XOR U10197 ( .A(n8531), .B(n8530), .Z(n9055) );
  XNOR U10198 ( .A(n9056), .B(n9055), .Z(n9058) );
  NANDN U10199 ( .A(n7812), .B(n7811), .Z(n7816) );
  NANDN U10200 ( .A(n7814), .B(n7813), .Z(n7815) );
  NAND U10201 ( .A(n7816), .B(n7815), .Z(n8982) );
  NANDN U10202 ( .A(n7818), .B(n7817), .Z(n7822) );
  NANDN U10203 ( .A(n7820), .B(n7819), .Z(n7821) );
  AND U10204 ( .A(n7822), .B(n7821), .Z(n8603) );
  NANDN U10205 ( .A(n7828), .B(n7827), .Z(n7832) );
  NAND U10206 ( .A(n7830), .B(n7829), .Z(n7831) );
  NAND U10207 ( .A(n7832), .B(n7831), .Z(n8656) );
  XNOR U10208 ( .A(n8656), .B(n8657), .Z(n8659) );
  XOR U10209 ( .A(n8658), .B(n8659), .Z(n8600) );
  NANDN U10210 ( .A(n7838), .B(n7837), .Z(n7842) );
  NANDN U10211 ( .A(n7840), .B(n7839), .Z(n7841) );
  NAND U10212 ( .A(n7842), .B(n7841), .Z(n8601) );
  XOR U10213 ( .A(n8600), .B(n8601), .Z(n8602) );
  XOR U10214 ( .A(n8603), .B(n8602), .Z(n8981) );
  NANDN U10215 ( .A(n7844), .B(n7843), .Z(n7848) );
  NANDN U10216 ( .A(n7846), .B(n7845), .Z(n7847) );
  NAND U10217 ( .A(n7848), .B(n7847), .Z(n8980) );
  XNOR U10218 ( .A(n8981), .B(n8980), .Z(n8983) );
  NANDN U10219 ( .A(n7850), .B(n7849), .Z(n7854) );
  OR U10220 ( .A(n7852), .B(n7851), .Z(n7853) );
  AND U10221 ( .A(n7854), .B(n7853), .Z(n8871) );
  NANDN U10222 ( .A(n7856), .B(n7855), .Z(n7860) );
  OR U10223 ( .A(n7858), .B(n7857), .Z(n7859) );
  AND U10224 ( .A(n7860), .B(n7859), .Z(n8870) );
  XNOR U10225 ( .A(n8871), .B(n8870), .Z(n8872) );
  XOR U10226 ( .A(n8873), .B(n8872), .Z(n8719) );
  NANDN U10227 ( .A(n7862), .B(n7861), .Z(n7866) );
  NANDN U10228 ( .A(n7864), .B(n7863), .Z(n7865) );
  AND U10229 ( .A(n7866), .B(n7865), .Z(n8716) );
  NANDN U10230 ( .A(n7868), .B(n7867), .Z(n7872) );
  OR U10231 ( .A(n7870), .B(n7869), .Z(n7871) );
  AND U10232 ( .A(n7872), .B(n7871), .Z(n8975) );
  NANDN U10233 ( .A(n7874), .B(n7873), .Z(n7878) );
  OR U10234 ( .A(n7876), .B(n7875), .Z(n7877) );
  AND U10235 ( .A(n7878), .B(n7877), .Z(n8970) );
  NANDN U10236 ( .A(n7880), .B(n7879), .Z(n7884) );
  NANDN U10237 ( .A(n7882), .B(n7881), .Z(n7883) );
  AND U10238 ( .A(n7884), .B(n7883), .Z(n8969) );
  NANDN U10239 ( .A(n7886), .B(n7885), .Z(n7890) );
  NANDN U10240 ( .A(n7888), .B(n7887), .Z(n7889) );
  NAND U10241 ( .A(n7890), .B(n7889), .Z(n8968) );
  XOR U10242 ( .A(n8969), .B(n8968), .Z(n8971) );
  XNOR U10243 ( .A(n8970), .B(n8971), .Z(n8974) );
  XNOR U10244 ( .A(n8975), .B(n8974), .Z(n8976) );
  NANDN U10245 ( .A(n7892), .B(n7891), .Z(n7896) );
  NANDN U10246 ( .A(n7894), .B(n7893), .Z(n7895) );
  AND U10247 ( .A(n7896), .B(n7895), .Z(n8839) );
  NANDN U10248 ( .A(n7898), .B(n7897), .Z(n7902) );
  OR U10249 ( .A(n7900), .B(n7899), .Z(n7901) );
  AND U10250 ( .A(n7902), .B(n7901), .Z(n8837) );
  NANDN U10251 ( .A(n7904), .B(n7903), .Z(n7908) );
  NANDN U10252 ( .A(n7906), .B(n7905), .Z(n7907) );
  AND U10253 ( .A(n7908), .B(n7907), .Z(n8781) );
  NANDN U10254 ( .A(n7914), .B(n7913), .Z(n7918) );
  NAND U10255 ( .A(n7916), .B(n7915), .Z(n7917) );
  NAND U10256 ( .A(n7918), .B(n7917), .Z(n8779) );
  XOR U10257 ( .A(n8778), .B(n8779), .Z(n8780) );
  XNOR U10258 ( .A(n8781), .B(n8780), .Z(n8836) );
  XNOR U10259 ( .A(n8837), .B(n8836), .Z(n8838) );
  XOR U10260 ( .A(n8839), .B(n8838), .Z(n8977) );
  XOR U10261 ( .A(n8976), .B(n8977), .Z(n8717) );
  XNOR U10262 ( .A(n8716), .B(n8717), .Z(n8718) );
  XOR U10263 ( .A(n8719), .B(n8718), .Z(n8899) );
  NANDN U10264 ( .A(n7920), .B(n7919), .Z(n7924) );
  NAND U10265 ( .A(n7922), .B(n7921), .Z(n7923) );
  AND U10266 ( .A(n7924), .B(n7923), .Z(n9046) );
  XOR U10267 ( .A(n8783), .B(n8782), .Z(n8785) );
  XOR U10268 ( .A(n8784), .B(n8785), .Z(n9044) );
  NANDN U10269 ( .A(n7938), .B(n7937), .Z(n7942) );
  OR U10270 ( .A(n7940), .B(n7939), .Z(n7941) );
  NAND U10271 ( .A(n7942), .B(n7941), .Z(n9043) );
  XNOR U10272 ( .A(n9044), .B(n9043), .Z(n9045) );
  XOR U10273 ( .A(n9046), .B(n9045), .Z(n8774) );
  NANDN U10274 ( .A(n7944), .B(n7943), .Z(n7948) );
  NANDN U10275 ( .A(n7946), .B(n7945), .Z(n7947) );
  AND U10276 ( .A(n7948), .B(n7947), .Z(n8666) );
  NANDN U10277 ( .A(n7950), .B(n7949), .Z(n7954) );
  NANDN U10278 ( .A(n7952), .B(n7951), .Z(n7953) );
  AND U10279 ( .A(n7954), .B(n7953), .Z(n8665) );
  NANDN U10280 ( .A(n7956), .B(n7955), .Z(n7960) );
  NAND U10281 ( .A(n7958), .B(n7957), .Z(n7959) );
  AND U10282 ( .A(n7960), .B(n7959), .Z(n8832) );
  XOR U10283 ( .A(n8831), .B(n8830), .Z(n8833) );
  XNOR U10284 ( .A(n8832), .B(n8833), .Z(n8664) );
  XOR U10285 ( .A(n8665), .B(n8664), .Z(n8667) );
  XOR U10286 ( .A(n8666), .B(n8667), .Z(n8773) );
  NANDN U10287 ( .A(n7974), .B(n7973), .Z(n7978) );
  NAND U10288 ( .A(n7976), .B(n7975), .Z(n7977) );
  NAND U10289 ( .A(n7978), .B(n7977), .Z(n8944) );
  XOR U10290 ( .A(n8944), .B(n8945), .Z(n8947) );
  XOR U10291 ( .A(n8946), .B(n8947), .Z(n8604) );
  NANDN U10292 ( .A(n7984), .B(n7983), .Z(n7988) );
  NANDN U10293 ( .A(n7986), .B(n7985), .Z(n7987) );
  NAND U10294 ( .A(n7988), .B(n7987), .Z(n8605) );
  XNOR U10295 ( .A(n8604), .B(n8605), .Z(n8606) );
  NANDN U10296 ( .A(n7990), .B(n7989), .Z(n7994) );
  NANDN U10297 ( .A(n7992), .B(n7991), .Z(n7993) );
  NAND U10298 ( .A(n7994), .B(n7993), .Z(n8607) );
  XNOR U10299 ( .A(n8606), .B(n8607), .Z(n8772) );
  XOR U10300 ( .A(n8773), .B(n8772), .Z(n8775) );
  XOR U10301 ( .A(n8774), .B(n8775), .Z(n8547) );
  NANDN U10302 ( .A(n7996), .B(n7995), .Z(n8000) );
  NANDN U10303 ( .A(n7998), .B(n7997), .Z(n7999) );
  AND U10304 ( .A(n8000), .B(n7999), .Z(n8818) );
  NANDN U10305 ( .A(n8002), .B(n8001), .Z(n8006) );
  NANDN U10306 ( .A(n8004), .B(n8003), .Z(n8005) );
  NAND U10307 ( .A(n8006), .B(n8005), .Z(n8819) );
  XNOR U10308 ( .A(n8818), .B(n8819), .Z(n8820) );
  NANDN U10309 ( .A(n8008), .B(n8007), .Z(n8012) );
  NANDN U10310 ( .A(n8010), .B(n8009), .Z(n8011) );
  NAND U10311 ( .A(n8012), .B(n8011), .Z(n8821) );
  XNOR U10312 ( .A(n8820), .B(n8821), .Z(n9010) );
  NANDN U10313 ( .A(n8014), .B(n8013), .Z(n8018) );
  NAND U10314 ( .A(n8016), .B(n8015), .Z(n8017) );
  NAND U10315 ( .A(n8018), .B(n8017), .Z(n9008) );
  NANDN U10316 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U10317 ( .A(n8022), .B(n8021), .Z(n8023) );
  AND U10318 ( .A(n8024), .B(n8023), .Z(n8794) );
  NANDN U10319 ( .A(n8026), .B(n8025), .Z(n8030) );
  NANDN U10320 ( .A(n8028), .B(n8027), .Z(n8029) );
  NAND U10321 ( .A(n8030), .B(n8029), .Z(n8795) );
  XNOR U10322 ( .A(n8794), .B(n8795), .Z(n8796) );
  NANDN U10323 ( .A(n8032), .B(n8031), .Z(n8036) );
  NANDN U10324 ( .A(n8034), .B(n8033), .Z(n8035) );
  NAND U10325 ( .A(n8036), .B(n8035), .Z(n8797) );
  XOR U10326 ( .A(n8796), .B(n8797), .Z(n9009) );
  XNOR U10327 ( .A(n9008), .B(n9009), .Z(n9011) );
  XOR U10328 ( .A(n9010), .B(n9011), .Z(n8737) );
  NANDN U10329 ( .A(n8038), .B(n8037), .Z(n8042) );
  NANDN U10330 ( .A(n8040), .B(n8039), .Z(n8041) );
  NAND U10331 ( .A(n8042), .B(n8041), .Z(n8994) );
  NANDN U10332 ( .A(n8044), .B(n8043), .Z(n8048) );
  NANDN U10333 ( .A(n8046), .B(n8045), .Z(n8047) );
  NAND U10334 ( .A(n8048), .B(n8047), .Z(n8992) );
  NANDN U10335 ( .A(n8050), .B(n8049), .Z(n8054) );
  NAND U10336 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U10337 ( .A(n8054), .B(n8053), .Z(n8993) );
  XNOR U10338 ( .A(n8992), .B(n8993), .Z(n8995) );
  XOR U10339 ( .A(n8994), .B(n8995), .Z(n8734) );
  XOR U10340 ( .A(n8789), .B(n8788), .Z(n8791) );
  XNOR U10341 ( .A(n8790), .B(n8791), .Z(n8735) );
  XOR U10342 ( .A(n8734), .B(n8735), .Z(n8736) );
  XOR U10343 ( .A(n8737), .B(n8736), .Z(n8848) );
  NANDN U10344 ( .A(n8068), .B(n8067), .Z(n8072) );
  NAND U10345 ( .A(n8070), .B(n8069), .Z(n8071) );
  AND U10346 ( .A(n8072), .B(n8071), .Z(n8895) );
  NANDN U10347 ( .A(n8078), .B(n8077), .Z(n8082) );
  NANDN U10348 ( .A(n8080), .B(n8079), .Z(n8081) );
  AND U10349 ( .A(n8082), .B(n8081), .Z(n9003) );
  XNOR U10350 ( .A(n9003), .B(n9002), .Z(n9004) );
  XOR U10351 ( .A(n9005), .B(n9004), .Z(n8893) );
  NANDN U10352 ( .A(n8088), .B(n8087), .Z(n8092) );
  NANDN U10353 ( .A(n8090), .B(n8089), .Z(n8091) );
  NAND U10354 ( .A(n8092), .B(n8091), .Z(n8892) );
  XOR U10355 ( .A(n8893), .B(n8892), .Z(n8894) );
  XOR U10356 ( .A(n8895), .B(n8894), .Z(n8847) );
  NANDN U10357 ( .A(n8094), .B(n8093), .Z(n8098) );
  NANDN U10358 ( .A(n8096), .B(n8095), .Z(n8097) );
  AND U10359 ( .A(n8098), .B(n8097), .Z(n8628) );
  XNOR U10360 ( .A(n8617), .B(n8616), .Z(n8618) );
  XOR U10361 ( .A(n8619), .B(n8618), .Z(n8629) );
  XNOR U10362 ( .A(n8628), .B(n8629), .Z(n8630) );
  NANDN U10363 ( .A(n8112), .B(n8111), .Z(n8116) );
  NANDN U10364 ( .A(n8114), .B(n8113), .Z(n8115) );
  NAND U10365 ( .A(n8116), .B(n8115), .Z(n8631) );
  XNOR U10366 ( .A(n8630), .B(n8631), .Z(n8846) );
  XOR U10367 ( .A(n8847), .B(n8846), .Z(n8849) );
  XOR U10368 ( .A(n8848), .B(n8849), .Z(n8546) );
  XNOR U10369 ( .A(n8547), .B(n8546), .Z(n8549) );
  NANDN U10370 ( .A(n8118), .B(n8117), .Z(n8122) );
  NAND U10371 ( .A(n8120), .B(n8119), .Z(n8121) );
  AND U10372 ( .A(n8122), .B(n8121), .Z(n8691) );
  NANDN U10373 ( .A(n8124), .B(n8123), .Z(n8128) );
  NAND U10374 ( .A(n8126), .B(n8125), .Z(n8127) );
  AND U10375 ( .A(n8128), .B(n8127), .Z(n8689) );
  NANDN U10376 ( .A(n8134), .B(n8133), .Z(n8138) );
  NAND U10377 ( .A(n8136), .B(n8135), .Z(n8137) );
  NAND U10378 ( .A(n8138), .B(n8137), .Z(n8660) );
  NANDN U10379 ( .A(n8140), .B(n8139), .Z(n8144) );
  NAND U10380 ( .A(n8142), .B(n8141), .Z(n8143) );
  NAND U10381 ( .A(n8144), .B(n8143), .Z(n8661) );
  XOR U10382 ( .A(n8660), .B(n8661), .Z(n8663) );
  XOR U10383 ( .A(n8662), .B(n8663), .Z(n8925) );
  NANDN U10384 ( .A(n8146), .B(n8145), .Z(n8150) );
  NAND U10385 ( .A(n8148), .B(n8147), .Z(n8149) );
  NAND U10386 ( .A(n8150), .B(n8149), .Z(n8942) );
  NANDN U10387 ( .A(n8156), .B(n8155), .Z(n8160) );
  NAND U10388 ( .A(n8158), .B(n8157), .Z(n8159) );
  NAND U10389 ( .A(n8160), .B(n8159), .Z(n8941) );
  XOR U10390 ( .A(n8940), .B(n8941), .Z(n8943) );
  XOR U10391 ( .A(n8942), .B(n8943), .Z(n8923) );
  NANDN U10392 ( .A(n8162), .B(n8161), .Z(n8166) );
  NAND U10393 ( .A(n8164), .B(n8163), .Z(n8165) );
  AND U10394 ( .A(n8166), .B(n8165), .Z(n8560) );
  NANDN U10395 ( .A(n8168), .B(n8167), .Z(n8172) );
  NANDN U10396 ( .A(n8170), .B(n8169), .Z(n8171) );
  AND U10397 ( .A(n8172), .B(n8171), .Z(n8559) );
  NANDN U10398 ( .A(n8174), .B(n8173), .Z(n8178) );
  OR U10399 ( .A(n8176), .B(n8175), .Z(n8177) );
  AND U10400 ( .A(n8178), .B(n8177), .Z(n8959) );
  NANDN U10401 ( .A(n8180), .B(n8179), .Z(n8184) );
  NANDN U10402 ( .A(n8182), .B(n8181), .Z(n8183) );
  AND U10403 ( .A(n8184), .B(n8183), .Z(n8957) );
  XOR U10404 ( .A(n8957), .B(n8956), .Z(n8958) );
  XNOR U10405 ( .A(n8959), .B(n8958), .Z(n8558) );
  XOR U10406 ( .A(n8559), .B(n8558), .Z(n8561) );
  XNOR U10407 ( .A(n8560), .B(n8561), .Z(n8922) );
  XNOR U10408 ( .A(n8923), .B(n8922), .Z(n8924) );
  XNOR U10409 ( .A(n8925), .B(n8924), .Z(n8688) );
  XNOR U10410 ( .A(n8689), .B(n8688), .Z(n8690) );
  XNOR U10411 ( .A(n8691), .B(n8690), .Z(n8548) );
  XOR U10412 ( .A(n8549), .B(n8548), .Z(n8898) );
  XOR U10413 ( .A(n8899), .B(n8898), .Z(n8901) );
  NANDN U10414 ( .A(n8190), .B(n8189), .Z(n8194) );
  NANDN U10415 ( .A(n8192), .B(n8191), .Z(n8193) );
  AND U10416 ( .A(n8194), .B(n8193), .Z(n8859) );
  NANDN U10417 ( .A(n8196), .B(n8195), .Z(n8200) );
  NANDN U10418 ( .A(n8198), .B(n8197), .Z(n8199) );
  AND U10419 ( .A(n8200), .B(n8199), .Z(n9040) );
  NANDN U10420 ( .A(n8202), .B(n8201), .Z(n8206) );
  NANDN U10421 ( .A(n8204), .B(n8203), .Z(n8205) );
  AND U10422 ( .A(n8206), .B(n8205), .Z(n9039) );
  XOR U10423 ( .A(n9040), .B(n9039), .Z(n9042) );
  NANDN U10424 ( .A(n8208), .B(n8207), .Z(n8212) );
  OR U10425 ( .A(n8210), .B(n8209), .Z(n8211) );
  AND U10426 ( .A(n8212), .B(n8211), .Z(n9041) );
  XOR U10427 ( .A(n9042), .B(n9041), .Z(n8612) );
  NANDN U10428 ( .A(n8214), .B(n8213), .Z(n8218) );
  NAND U10429 ( .A(n8216), .B(n8215), .Z(n8217) );
  AND U10430 ( .A(n8218), .B(n8217), .Z(n8611) );
  NANDN U10431 ( .A(n8220), .B(n8219), .Z(n8224) );
  NANDN U10432 ( .A(n8222), .B(n8221), .Z(n8223) );
  AND U10433 ( .A(n8224), .B(n8223), .Z(n8649) );
  NANDN U10434 ( .A(n8226), .B(n8225), .Z(n8230) );
  OR U10435 ( .A(n8228), .B(n8227), .Z(n8229) );
  AND U10436 ( .A(n8230), .B(n8229), .Z(n8648) );
  XOR U10437 ( .A(n8649), .B(n8648), .Z(n8651) );
  NANDN U10438 ( .A(n8232), .B(n8231), .Z(n8236) );
  OR U10439 ( .A(n8234), .B(n8233), .Z(n8235) );
  AND U10440 ( .A(n8236), .B(n8235), .Z(n8650) );
  XNOR U10441 ( .A(n8651), .B(n8650), .Z(n8610) );
  XOR U10442 ( .A(n8611), .B(n8610), .Z(n8613) );
  XOR U10443 ( .A(n8612), .B(n8613), .Z(n8931) );
  NANDN U10444 ( .A(n8242), .B(n8241), .Z(n8246) );
  NANDN U10445 ( .A(n8244), .B(n8243), .Z(n8245) );
  AND U10446 ( .A(n8246), .B(n8245), .Z(n8582) );
  XNOR U10447 ( .A(n8582), .B(n8583), .Z(n8584) );
  XOR U10448 ( .A(n8584), .B(n8585), .Z(n8965) );
  XNOR U10449 ( .A(n8965), .B(n8964), .Z(n8967) );
  XOR U10450 ( .A(n8966), .B(n8967), .Z(n8928) );
  NANDN U10451 ( .A(n8264), .B(n8263), .Z(n8268) );
  NANDN U10452 ( .A(n8266), .B(n8265), .Z(n8267) );
  AND U10453 ( .A(n8268), .B(n8267), .Z(n8806) );
  XNOR U10454 ( .A(n8806), .B(n8807), .Z(n8809) );
  XOR U10455 ( .A(n8809), .B(n8808), .Z(n8987) );
  XOR U10456 ( .A(n8987), .B(n8986), .Z(n8989) );
  XNOR U10457 ( .A(n8988), .B(n8989), .Z(n8929) );
  XOR U10458 ( .A(n8928), .B(n8929), .Z(n8930) );
  XNOR U10459 ( .A(n8931), .B(n8930), .Z(n8858) );
  XNOR U10460 ( .A(n8859), .B(n8858), .Z(n8861) );
  NANDN U10461 ( .A(n8282), .B(n8281), .Z(n8286) );
  NANDN U10462 ( .A(n8284), .B(n8283), .Z(n8285) );
  AND U10463 ( .A(n8286), .B(n8285), .Z(n8707) );
  NANDN U10464 ( .A(n8296), .B(n8295), .Z(n8300) );
  NAND U10465 ( .A(n8298), .B(n8297), .Z(n8299) );
  NAND U10466 ( .A(n8300), .B(n8299), .Z(n9012) );
  XNOR U10467 ( .A(n9012), .B(n9013), .Z(n9015) );
  XOR U10468 ( .A(n9014), .B(n9015), .Z(n8704) );
  XNOR U10469 ( .A(n8705), .B(n8704), .Z(n8706) );
  XNOR U10470 ( .A(n8707), .B(n8706), .Z(n8860) );
  XOR U10471 ( .A(n8861), .B(n8860), .Z(n8769) );
  NANDN U10472 ( .A(n8306), .B(n8305), .Z(n8310) );
  NANDN U10473 ( .A(n8308), .B(n8307), .Z(n8309) );
  AND U10474 ( .A(n8310), .B(n8309), .Z(n9052) );
  NAND U10475 ( .A(n8312), .B(n8311), .Z(n8316) );
  NANDN U10476 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U10477 ( .A(n8316), .B(n8315), .Z(n9050) );
  NANDN U10478 ( .A(n8322), .B(n8321), .Z(n8326) );
  NAND U10479 ( .A(n8324), .B(n8323), .Z(n8325) );
  AND U10480 ( .A(n8326), .B(n8325), .Z(n8565) );
  NANDN U10481 ( .A(n8328), .B(n8327), .Z(n8332) );
  NAND U10482 ( .A(n8330), .B(n8329), .Z(n8331) );
  NAND U10483 ( .A(n8332), .B(n8331), .Z(n8564) );
  XNOR U10484 ( .A(n8565), .B(n8564), .Z(n8566) );
  XNOR U10485 ( .A(n8567), .B(n8566), .Z(n8634) );
  NANDN U10486 ( .A(n8334), .B(n8333), .Z(n8338) );
  NANDN U10487 ( .A(n8336), .B(n8335), .Z(n8337) );
  NAND U10488 ( .A(n8338), .B(n8337), .Z(n8635) );
  XNOR U10489 ( .A(n8634), .B(n8635), .Z(n8637) );
  NANDN U10490 ( .A(n8340), .B(n8339), .Z(n8344) );
  NANDN U10491 ( .A(n8342), .B(n8341), .Z(n8343) );
  AND U10492 ( .A(n8344), .B(n8343), .Z(n8636) );
  XNOR U10493 ( .A(n8637), .B(n8636), .Z(n9049) );
  XOR U10494 ( .A(n9052), .B(n9051), .Z(n8767) );
  NAND U10495 ( .A(n8346), .B(n8345), .Z(n8350) );
  NAND U10496 ( .A(n8348), .B(n8347), .Z(n8349) );
  AND U10497 ( .A(n8350), .B(n8349), .Z(n8919) );
  NAND U10498 ( .A(n8352), .B(n8351), .Z(n8356) );
  NAND U10499 ( .A(n8354), .B(n8353), .Z(n8355) );
  AND U10500 ( .A(n8356), .B(n8355), .Z(n8917) );
  NAND U10501 ( .A(n8358), .B(n8357), .Z(n8362) );
  NAND U10502 ( .A(n8360), .B(n8359), .Z(n8361) );
  NAND U10503 ( .A(n8362), .B(n8361), .Z(n8916) );
  XNOR U10504 ( .A(n8919), .B(n8918), .Z(n8766) );
  XNOR U10505 ( .A(n8767), .B(n8766), .Z(n8768) );
  XOR U10506 ( .A(n8769), .B(n8768), .Z(n8900) );
  XOR U10507 ( .A(n8901), .B(n8900), .Z(n8907) );
  NAND U10508 ( .A(n8364), .B(n8363), .Z(n8368) );
  NAND U10509 ( .A(n8366), .B(n8365), .Z(n8367) );
  AND U10510 ( .A(n8368), .B(n8367), .Z(n8904) );
  NANDN U10511 ( .A(n8370), .B(n8369), .Z(n8374) );
  NANDN U10512 ( .A(n8372), .B(n8371), .Z(n8373) );
  NAND U10513 ( .A(n8374), .B(n8373), .Z(n8905) );
  XNOR U10514 ( .A(n8904), .B(n8905), .Z(n8906) );
  XNOR U10515 ( .A(n8907), .B(n8906), .Z(n8525) );
  NAND U10516 ( .A(n8376), .B(n8375), .Z(n8380) );
  NANDN U10517 ( .A(n8378), .B(n8377), .Z(n8379) );
  AND U10518 ( .A(n8380), .B(n8379), .Z(n8523) );
  NANDN U10519 ( .A(n8382), .B(n8381), .Z(n8386) );
  NANDN U10520 ( .A(n8384), .B(n8383), .Z(n8385) );
  AND U10521 ( .A(n8386), .B(n8385), .Z(n8677) );
  NANDN U10522 ( .A(n8388), .B(n8387), .Z(n8392) );
  NANDN U10523 ( .A(n8390), .B(n8389), .Z(n8391) );
  AND U10524 ( .A(n8392), .B(n8391), .Z(n8676) );
  XNOR U10525 ( .A(n8677), .B(n8676), .Z(n8679) );
  NANDN U10526 ( .A(n8394), .B(n8393), .Z(n8398) );
  NANDN U10527 ( .A(n8396), .B(n8395), .Z(n8397) );
  AND U10528 ( .A(n8398), .B(n8397), .Z(n8678) );
  XOR U10529 ( .A(n8679), .B(n8678), .Z(n8913) );
  NANDN U10530 ( .A(n8400), .B(n8399), .Z(n8404) );
  NAND U10531 ( .A(n8402), .B(n8401), .Z(n8403) );
  AND U10532 ( .A(n8404), .B(n8403), .Z(n8865) );
  NANDN U10533 ( .A(n8406), .B(n8405), .Z(n8410) );
  OR U10534 ( .A(n8408), .B(n8407), .Z(n8409) );
  AND U10535 ( .A(n8410), .B(n8409), .Z(n8738) );
  XNOR U10536 ( .A(n8738), .B(n8739), .Z(n8740) );
  NANDN U10537 ( .A(n8416), .B(n8415), .Z(n8420) );
  NANDN U10538 ( .A(n8418), .B(n8417), .Z(n8419) );
  NAND U10539 ( .A(n8420), .B(n8419), .Z(n8741) );
  XNOR U10540 ( .A(n8740), .B(n8741), .Z(n8694) );
  NANDN U10541 ( .A(n8422), .B(n8421), .Z(n8426) );
  NANDN U10542 ( .A(n8424), .B(n8423), .Z(n8425) );
  AND U10543 ( .A(n8426), .B(n8425), .Z(n8653) );
  XOR U10544 ( .A(n8653), .B(n8652), .Z(n8655) );
  NANDN U10545 ( .A(n8432), .B(n8431), .Z(n8436) );
  NANDN U10546 ( .A(n8434), .B(n8433), .Z(n8435) );
  AND U10547 ( .A(n8436), .B(n8435), .Z(n8654) );
  XOR U10548 ( .A(n8655), .B(n8654), .Z(n8827) );
  NANDN U10549 ( .A(n8438), .B(n8437), .Z(n8442) );
  NANDN U10550 ( .A(n8440), .B(n8439), .Z(n8441) );
  AND U10551 ( .A(n8442), .B(n8441), .Z(n8825) );
  NANDN U10552 ( .A(n8444), .B(n8443), .Z(n8448) );
  NANDN U10553 ( .A(n8446), .B(n8445), .Z(n8447) );
  NAND U10554 ( .A(n8448), .B(n8447), .Z(n8824) );
  XOR U10555 ( .A(n8641), .B(n8640), .Z(n8644) );
  XOR U10556 ( .A(n8643), .B(n9168), .Z(n8463) );
  XOR U10557 ( .A(n8644), .B(n8463), .Z(n9017) );
  NANDN U10558 ( .A(n8465), .B(n8464), .Z(n8469) );
  NAND U10559 ( .A(n8467), .B(n8466), .Z(n8468) );
  AND U10560 ( .A(n8469), .B(n8468), .Z(n9016) );
  XNOR U10561 ( .A(n9017), .B(n9016), .Z(n9019) );
  XOR U10562 ( .A(n9018), .B(n9019), .Z(n8745) );
  NANDN U10563 ( .A(n8471), .B(n8470), .Z(n8475) );
  OR U10564 ( .A(n8473), .B(n8472), .Z(n8474) );
  AND U10565 ( .A(n8475), .B(n8474), .Z(n8744) );
  XNOR U10566 ( .A(n8745), .B(n8744), .Z(n8746) );
  NANDN U10567 ( .A(n8481), .B(n8480), .Z(n8485) );
  NANDN U10568 ( .A(n8483), .B(n8482), .Z(n8484) );
  AND U10569 ( .A(n8485), .B(n8484), .Z(n8623) );
  NANDN U10570 ( .A(n8487), .B(n8486), .Z(n8491) );
  NANDN U10571 ( .A(n8489), .B(n8488), .Z(n8490) );
  AND U10572 ( .A(n8491), .B(n8490), .Z(n9036) );
  NANDN U10573 ( .A(n8493), .B(n8492), .Z(n8497) );
  OR U10574 ( .A(n8495), .B(n8494), .Z(n8496) );
  AND U10575 ( .A(n8497), .B(n8496), .Z(n9035) );
  XOR U10576 ( .A(n9036), .B(n9035), .Z(n9038) );
  NANDN U10577 ( .A(n8499), .B(n8498), .Z(n8503) );
  OR U10578 ( .A(n8501), .B(n8500), .Z(n8502) );
  AND U10579 ( .A(n8503), .B(n8502), .Z(n9037) );
  XNOR U10580 ( .A(n9038), .B(n9037), .Z(n8622) );
  XNOR U10581 ( .A(n8623), .B(n8622), .Z(n8624) );
  XOR U10582 ( .A(n8625), .B(n8624), .Z(n8747) );
  XOR U10583 ( .A(n8746), .B(n8747), .Z(n8695) );
  XNOR U10584 ( .A(n8694), .B(n8695), .Z(n8696) );
  NANDN U10585 ( .A(n8505), .B(n8504), .Z(n8509) );
  OR U10586 ( .A(n8507), .B(n8506), .Z(n8508) );
  NAND U10587 ( .A(n8509), .B(n8508), .Z(n8697) );
  XNOR U10588 ( .A(n8696), .B(n8697), .Z(n8864) );
  XNOR U10589 ( .A(n8865), .B(n8864), .Z(n8866) );
  NANDN U10590 ( .A(n8511), .B(n8510), .Z(n8515) );
  NAND U10591 ( .A(n8513), .B(n8512), .Z(n8514) );
  NAND U10592 ( .A(n8515), .B(n8514), .Z(n8867) );
  XNOR U10593 ( .A(n8866), .B(n8867), .Z(n8910) );
  NAND U10594 ( .A(n8517), .B(n8516), .Z(n8521) );
  NAND U10595 ( .A(n8519), .B(n8518), .Z(n8520) );
  NAND U10596 ( .A(n8521), .B(n8520), .Z(n8911) );
  XNOR U10597 ( .A(n8910), .B(n8911), .Z(n8912) );
  XOR U10598 ( .A(n8913), .B(n8912), .Z(n8522) );
  XOR U10599 ( .A(n8523), .B(n8522), .Z(n8524) );
  XOR U10600 ( .A(n8525), .B(n8524), .Z(n9057) );
  XNOR U10601 ( .A(n9058), .B(n9057), .Z(o[3]) );
  NAND U10602 ( .A(n8523), .B(n8522), .Z(n8527) );
  NANDN U10603 ( .A(n8525), .B(n8524), .Z(n8526) );
  AND U10604 ( .A(n8527), .B(n8526), .Z(n9064) );
  NANDN U10605 ( .A(n8529), .B(n8528), .Z(n8533) );
  NAND U10606 ( .A(n8531), .B(n8530), .Z(n8532) );
  NAND U10607 ( .A(n8533), .B(n8532), .Z(n9062) );
  NANDN U10608 ( .A(n8535), .B(n8534), .Z(n8539) );
  NANDN U10609 ( .A(n8537), .B(n8536), .Z(n8538) );
  AND U10610 ( .A(n8539), .B(n8538), .Z(n9310) );
  NANDN U10611 ( .A(n8541), .B(n8540), .Z(n8545) );
  NANDN U10612 ( .A(n8543), .B(n8542), .Z(n8544) );
  AND U10613 ( .A(n8545), .B(n8544), .Z(n9127) );
  NANDN U10614 ( .A(n8547), .B(n8546), .Z(n8551) );
  NAND U10615 ( .A(n8549), .B(n8548), .Z(n8550) );
  AND U10616 ( .A(n8551), .B(n8550), .Z(n9125) );
  NANDN U10617 ( .A(n8553), .B(n8552), .Z(n8557) );
  OR U10618 ( .A(n8555), .B(n8554), .Z(n8556) );
  NAND U10619 ( .A(n8557), .B(n8556), .Z(n9230) );
  NANDN U10620 ( .A(n8559), .B(n8558), .Z(n8563) );
  OR U10621 ( .A(n8561), .B(n8560), .Z(n8562) );
  NAND U10622 ( .A(n8563), .B(n8562), .Z(n9228) );
  NANDN U10623 ( .A(n8565), .B(n8564), .Z(n8569) );
  NANDN U10624 ( .A(n8567), .B(n8566), .Z(n8568) );
  NAND U10625 ( .A(n8569), .B(n8568), .Z(n9229) );
  XOR U10626 ( .A(n9228), .B(n9229), .Z(n9231) );
  XOR U10627 ( .A(n9230), .B(n9231), .Z(n9285) );
  NANDN U10628 ( .A(n8571), .B(n8570), .Z(n8575) );
  NAND U10629 ( .A(n8573), .B(n8572), .Z(n8574) );
  NAND U10630 ( .A(n8575), .B(n8574), .Z(n9192) );
  NANDN U10631 ( .A(n8577), .B(n8576), .Z(n8581) );
  NANDN U10632 ( .A(n8579), .B(n8578), .Z(n8580) );
  NAND U10633 ( .A(n8581), .B(n8580), .Z(n9190) );
  NANDN U10634 ( .A(n8583), .B(n8582), .Z(n8587) );
  NANDN U10635 ( .A(n8585), .B(n8584), .Z(n8586) );
  NAND U10636 ( .A(n8587), .B(n8586), .Z(n9191) );
  XOR U10637 ( .A(n9190), .B(n9191), .Z(n9193) );
  XOR U10638 ( .A(n9192), .B(n9193), .Z(n9153) );
  NANDN U10639 ( .A(n8589), .B(n8588), .Z(n8593) );
  OR U10640 ( .A(n8591), .B(n8590), .Z(n8592) );
  AND U10641 ( .A(n8593), .B(n8592), .Z(n9152) );
  XOR U10642 ( .A(n9153), .B(n9152), .Z(n9155) );
  NANDN U10643 ( .A(n8595), .B(n8594), .Z(n8599) );
  OR U10644 ( .A(n8597), .B(n8596), .Z(n8598) );
  AND U10645 ( .A(n8599), .B(n8598), .Z(n9154) );
  XOR U10646 ( .A(n9155), .B(n9154), .Z(n9283) );
  XNOR U10647 ( .A(n9283), .B(n9282), .Z(n9284) );
  XOR U10648 ( .A(n9285), .B(n9284), .Z(n9083) );
  NANDN U10649 ( .A(n8605), .B(n8604), .Z(n8609) );
  NANDN U10650 ( .A(n8607), .B(n8606), .Z(n8608) );
  AND U10651 ( .A(n8609), .B(n8608), .Z(n9272) );
  NANDN U10652 ( .A(n8611), .B(n8610), .Z(n8615) );
  OR U10653 ( .A(n8613), .B(n8612), .Z(n8614) );
  AND U10654 ( .A(n8615), .B(n8614), .Z(n9239) );
  NANDN U10655 ( .A(n8617), .B(n8616), .Z(n8621) );
  NANDN U10656 ( .A(n8619), .B(n8618), .Z(n8620) );
  AND U10657 ( .A(n8621), .B(n8620), .Z(n9237) );
  NANDN U10658 ( .A(n8623), .B(n8622), .Z(n8627) );
  NANDN U10659 ( .A(n8625), .B(n8624), .Z(n8626) );
  AND U10660 ( .A(n8627), .B(n8626), .Z(n9236) );
  XOR U10661 ( .A(n9237), .B(n9236), .Z(n9238) );
  XOR U10662 ( .A(n9239), .B(n9238), .Z(n9271) );
  NANDN U10663 ( .A(n8629), .B(n8628), .Z(n8633) );
  NANDN U10664 ( .A(n8631), .B(n8630), .Z(n8632) );
  NAND U10665 ( .A(n8633), .B(n8632), .Z(n9270) );
  XOR U10666 ( .A(n9271), .B(n9270), .Z(n9273) );
  XOR U10667 ( .A(n9272), .B(n9273), .Z(n9081) );
  NANDN U10668 ( .A(n8635), .B(n8634), .Z(n8639) );
  NAND U10669 ( .A(n8637), .B(n8636), .Z(n8638) );
  AND U10670 ( .A(n8639), .B(n8638), .Z(n9199) );
  NOR U10671 ( .A(n8643), .B(n9168), .Z(n8642) );
  XNOR U10672 ( .A(n9171), .B(n8642), .Z(n8647) );
  IV U10673 ( .A(n8643), .Z(n9169) );
  XNOR U10674 ( .A(n9169), .B(n9168), .Z(n8645) );
  NAND U10675 ( .A(n8645), .B(n8644), .Z(n8646) );
  NAND U10676 ( .A(n8647), .B(n8646), .Z(n9181) );
  XOR U10677 ( .A(n9179), .B(n9178), .Z(n9180) );
  XOR U10678 ( .A(n9181), .B(n9180), .Z(n9220) );
  XOR U10679 ( .A(n9220), .B(n9221), .Z(n9223) );
  XNOR U10680 ( .A(n9223), .B(n9222), .Z(n9198) );
  XNOR U10681 ( .A(n9199), .B(n9198), .Z(n9201) );
  NANDN U10682 ( .A(n8665), .B(n8664), .Z(n8669) );
  OR U10683 ( .A(n8667), .B(n8666), .Z(n8668) );
  AND U10684 ( .A(n8669), .B(n8668), .Z(n9200) );
  XNOR U10685 ( .A(n9201), .B(n9200), .Z(n9080) );
  XNOR U10686 ( .A(n9081), .B(n9080), .Z(n9082) );
  XNOR U10687 ( .A(n9083), .B(n9082), .Z(n9124) );
  XOR U10688 ( .A(n9127), .B(n9126), .Z(n9309) );
  XNOR U10689 ( .A(n9310), .B(n9309), .Z(n9312) );
  NANDN U10690 ( .A(n8671), .B(n8670), .Z(n8675) );
  NAND U10691 ( .A(n8673), .B(n8672), .Z(n8674) );
  AND U10692 ( .A(n8675), .B(n8674), .Z(n9311) );
  XOR U10693 ( .A(n9312), .B(n9311), .Z(n9063) );
  XNOR U10694 ( .A(n9062), .B(n9063), .Z(n9065) );
  NANDN U10695 ( .A(n8677), .B(n8676), .Z(n8681) );
  NAND U10696 ( .A(n8679), .B(n8678), .Z(n8680) );
  AND U10697 ( .A(n8681), .B(n8680), .Z(n9075) );
  NANDN U10698 ( .A(n8683), .B(n8682), .Z(n8687) );
  NAND U10699 ( .A(n8685), .B(n8684), .Z(n8686) );
  NAND U10700 ( .A(n8687), .B(n8686), .Z(n9074) );
  NANDN U10701 ( .A(n8689), .B(n8688), .Z(n8693) );
  NANDN U10702 ( .A(n8691), .B(n8690), .Z(n8692) );
  AND U10703 ( .A(n8693), .B(n8692), .Z(n9260) );
  NANDN U10704 ( .A(n8695), .B(n8694), .Z(n8699) );
  NANDN U10705 ( .A(n8697), .B(n8696), .Z(n8698) );
  AND U10706 ( .A(n8699), .B(n8698), .Z(n9259) );
  NANDN U10707 ( .A(n8705), .B(n8704), .Z(n8709) );
  NANDN U10708 ( .A(n8707), .B(n8706), .Z(n8708) );
  AND U10709 ( .A(n8709), .B(n8708), .Z(n9093) );
  NANDN U10710 ( .A(n8711), .B(n8710), .Z(n8715) );
  NAND U10711 ( .A(n8713), .B(n8712), .Z(n8714) );
  NAND U10712 ( .A(n8715), .B(n8714), .Z(n9092) );
  XOR U10713 ( .A(n9093), .B(n9092), .Z(n9094) );
  XOR U10714 ( .A(n9095), .B(n9094), .Z(n9258) );
  XOR U10715 ( .A(n9259), .B(n9258), .Z(n9261) );
  XOR U10716 ( .A(n9260), .B(n9261), .Z(n9290) );
  NANDN U10717 ( .A(n8717), .B(n8716), .Z(n8721) );
  NAND U10718 ( .A(n8719), .B(n8718), .Z(n8720) );
  NAND U10719 ( .A(n8721), .B(n8720), .Z(n9288) );
  NANDN U10720 ( .A(n8723), .B(n8722), .Z(n8727) );
  NANDN U10721 ( .A(n8725), .B(n8724), .Z(n8726) );
  AND U10722 ( .A(n8727), .B(n8726), .Z(n9265) );
  NANDN U10723 ( .A(n8729), .B(n8728), .Z(n8733) );
  NANDN U10724 ( .A(n8731), .B(n8730), .Z(n8732) );
  NAND U10725 ( .A(n8733), .B(n8732), .Z(n9264) );
  XNOR U10726 ( .A(n9265), .B(n9264), .Z(n9266) );
  NANDN U10727 ( .A(n8739), .B(n8738), .Z(n8743) );
  NANDN U10728 ( .A(n8741), .B(n8740), .Z(n8742) );
  NAND U10729 ( .A(n8743), .B(n8742), .Z(n9086) );
  XOR U10730 ( .A(n9087), .B(n9086), .Z(n9089) );
  NANDN U10731 ( .A(n8745), .B(n8744), .Z(n8749) );
  NANDN U10732 ( .A(n8747), .B(n8746), .Z(n8748) );
  NAND U10733 ( .A(n8749), .B(n8748), .Z(n9088) );
  XOR U10734 ( .A(n9089), .B(n9088), .Z(n9139) );
  NANDN U10735 ( .A(n8755), .B(n8754), .Z(n8759) );
  NANDN U10736 ( .A(n8757), .B(n8756), .Z(n8758) );
  NAND U10737 ( .A(n8759), .B(n8758), .Z(n9137) );
  XOR U10738 ( .A(n9136), .B(n9137), .Z(n9138) );
  XOR U10739 ( .A(n9139), .B(n9138), .Z(n9267) );
  XNOR U10740 ( .A(n9266), .B(n9267), .Z(n9289) );
  XOR U10741 ( .A(n9288), .B(n9289), .Z(n9291) );
  XOR U10742 ( .A(n9290), .B(n9291), .Z(n9076) );
  XOR U10743 ( .A(n9077), .B(n9076), .Z(n9318) );
  NANDN U10744 ( .A(n8761), .B(n8760), .Z(n8765) );
  NAND U10745 ( .A(n8763), .B(n8762), .Z(n8764) );
  AND U10746 ( .A(n8765), .B(n8764), .Z(n9133) );
  NANDN U10747 ( .A(n8767), .B(n8766), .Z(n8771) );
  NANDN U10748 ( .A(n8769), .B(n8768), .Z(n8770) );
  AND U10749 ( .A(n8771), .B(n8770), .Z(n9130) );
  NANDN U10750 ( .A(n8773), .B(n8772), .Z(n8777) );
  OR U10751 ( .A(n8775), .B(n8774), .Z(n8776) );
  AND U10752 ( .A(n8777), .B(n8776), .Z(n9114) );
  NANDN U10753 ( .A(n8783), .B(n8782), .Z(n8787) );
  OR U10754 ( .A(n8785), .B(n8784), .Z(n8786) );
  NAND U10755 ( .A(n8787), .B(n8786), .Z(n9224) );
  NANDN U10756 ( .A(n8789), .B(n8788), .Z(n8793) );
  OR U10757 ( .A(n8791), .B(n8790), .Z(n8792) );
  NAND U10758 ( .A(n8793), .B(n8792), .Z(n9225) );
  XOR U10759 ( .A(n9224), .B(n9225), .Z(n9227) );
  XOR U10760 ( .A(n9226), .B(n9227), .Z(n9279) );
  NANDN U10761 ( .A(n8795), .B(n8794), .Z(n8799) );
  NANDN U10762 ( .A(n8797), .B(n8796), .Z(n8798) );
  NAND U10763 ( .A(n8799), .B(n8798), .Z(n9184) );
  NANDN U10764 ( .A(n8801), .B(n8800), .Z(n8805) );
  NANDN U10765 ( .A(n8803), .B(n8802), .Z(n8804) );
  NAND U10766 ( .A(n8805), .B(n8804), .Z(n9182) );
  NANDN U10767 ( .A(n8807), .B(n8806), .Z(n8811) );
  NAND U10768 ( .A(n8809), .B(n8808), .Z(n8810) );
  NAND U10769 ( .A(n8811), .B(n8810), .Z(n9183) );
  XOR U10770 ( .A(n9182), .B(n9183), .Z(n9185) );
  XOR U10771 ( .A(n9184), .B(n9185), .Z(n9213) );
  NANDN U10772 ( .A(n8813), .B(n8812), .Z(n8817) );
  NAND U10773 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U10774 ( .A(n8817), .B(n8816), .Z(n9163) );
  NANDN U10775 ( .A(n8819), .B(n8818), .Z(n8823) );
  NANDN U10776 ( .A(n8821), .B(n8820), .Z(n8822) );
  NAND U10777 ( .A(n8823), .B(n8822), .Z(n9162) );
  XOR U10778 ( .A(n9163), .B(n9162), .Z(n9165) );
  NANDN U10779 ( .A(n8825), .B(n8824), .Z(n8829) );
  NANDN U10780 ( .A(n8827), .B(n8826), .Z(n8828) );
  AND U10781 ( .A(n8829), .B(n8828), .Z(n9164) );
  XOR U10782 ( .A(n9165), .B(n9164), .Z(n9211) );
  NANDN U10783 ( .A(n8831), .B(n8830), .Z(n8835) );
  OR U10784 ( .A(n8833), .B(n8832), .Z(n8834) );
  AND U10785 ( .A(n8835), .B(n8834), .Z(n9210) );
  XOR U10786 ( .A(n9211), .B(n9210), .Z(n9212) );
  XOR U10787 ( .A(n9213), .B(n9212), .Z(n9277) );
  NANDN U10788 ( .A(n8837), .B(n8836), .Z(n8841) );
  NANDN U10789 ( .A(n8839), .B(n8838), .Z(n8840) );
  AND U10790 ( .A(n8841), .B(n8840), .Z(n9276) );
  XNOR U10791 ( .A(n9277), .B(n9276), .Z(n9278) );
  XOR U10792 ( .A(n9279), .B(n9278), .Z(n9113) );
  XOR U10793 ( .A(n9113), .B(n9112), .Z(n9115) );
  XOR U10794 ( .A(n9114), .B(n9115), .Z(n9131) );
  NANDN U10795 ( .A(n8847), .B(n8846), .Z(n8851) );
  NANDN U10796 ( .A(n8849), .B(n8848), .Z(n8850) );
  AND U10797 ( .A(n8851), .B(n8850), .Z(n9119) );
  NANDN U10798 ( .A(n8853), .B(n8852), .Z(n8857) );
  NANDN U10799 ( .A(n8855), .B(n8854), .Z(n8856) );
  AND U10800 ( .A(n8857), .B(n8856), .Z(n9118) );
  XNOR U10801 ( .A(n9119), .B(n9118), .Z(n9120) );
  NANDN U10802 ( .A(n8859), .B(n8858), .Z(n8863) );
  NAND U10803 ( .A(n8861), .B(n8860), .Z(n8862) );
  NAND U10804 ( .A(n8863), .B(n8862), .Z(n9121) );
  XNOR U10805 ( .A(n9120), .B(n9121), .Z(n9297) );
  NANDN U10806 ( .A(n8865), .B(n8864), .Z(n8869) );
  NANDN U10807 ( .A(n8867), .B(n8866), .Z(n8868) );
  AND U10808 ( .A(n8869), .B(n8868), .Z(n9295) );
  NANDN U10809 ( .A(n8871), .B(n8870), .Z(n8875) );
  NAND U10810 ( .A(n8873), .B(n8872), .Z(n8874) );
  AND U10811 ( .A(n8875), .B(n8874), .Z(n9104) );
  NANDN U10812 ( .A(n8877), .B(n8876), .Z(n8881) );
  NANDN U10813 ( .A(n8879), .B(n8878), .Z(n8880) );
  AND U10814 ( .A(n8881), .B(n8880), .Z(n9102) );
  NANDN U10815 ( .A(n8883), .B(n8882), .Z(n8887) );
  NAND U10816 ( .A(n8885), .B(n8884), .Z(n8886) );
  AND U10817 ( .A(n8887), .B(n8886), .Z(n9249) );
  NAND U10818 ( .A(n8893), .B(n8892), .Z(n8897) );
  NAND U10819 ( .A(n8895), .B(n8894), .Z(n8896) );
  AND U10820 ( .A(n8897), .B(n8896), .Z(n9246) );
  XNOR U10821 ( .A(n9247), .B(n9246), .Z(n9248) );
  XOR U10822 ( .A(n9249), .B(n9248), .Z(n9103) );
  XOR U10823 ( .A(n9102), .B(n9103), .Z(n9105) );
  XNOR U10824 ( .A(n9104), .B(n9105), .Z(n9294) );
  XOR U10825 ( .A(n9297), .B(n9296), .Z(n9316) );
  XOR U10826 ( .A(n9315), .B(n9316), .Z(n9317) );
  XNOR U10827 ( .A(n9318), .B(n9317), .Z(n9071) );
  NAND U10828 ( .A(n8899), .B(n8898), .Z(n8903) );
  NAND U10829 ( .A(n8901), .B(n8900), .Z(n8902) );
  AND U10830 ( .A(n8903), .B(n8902), .Z(n9069) );
  NANDN U10831 ( .A(n8905), .B(n8904), .Z(n8909) );
  NANDN U10832 ( .A(n8907), .B(n8906), .Z(n8908) );
  AND U10833 ( .A(n8909), .B(n8908), .Z(n9324) );
  NANDN U10834 ( .A(n8911), .B(n8910), .Z(n8915) );
  NANDN U10835 ( .A(n8913), .B(n8912), .Z(n8914) );
  AND U10836 ( .A(n8915), .B(n8914), .Z(n9322) );
  NANDN U10837 ( .A(n8917), .B(n8916), .Z(n8921) );
  NAND U10838 ( .A(n8919), .B(n8918), .Z(n8920) );
  AND U10839 ( .A(n8921), .B(n8920), .Z(n9253) );
  NANDN U10840 ( .A(n8923), .B(n8922), .Z(n8927) );
  NANDN U10841 ( .A(n8925), .B(n8924), .Z(n8926) );
  AND U10842 ( .A(n8927), .B(n8926), .Z(n9099) );
  XNOR U10843 ( .A(n9097), .B(n9096), .Z(n9098) );
  XNOR U10844 ( .A(n9099), .B(n9098), .Z(n9252) );
  XOR U10845 ( .A(n9141), .B(n9140), .Z(n9143) );
  XOR U10846 ( .A(n9142), .B(n9143), .Z(n9159) );
  XOR U10847 ( .A(n9173), .B(n9172), .Z(n9175) );
  XOR U10848 ( .A(n9174), .B(n9175), .Z(n9147) );
  XOR U10849 ( .A(n9147), .B(n9146), .Z(n9149) );
  XOR U10850 ( .A(n9148), .B(n9149), .Z(n9157) );
  NANDN U10851 ( .A(n8969), .B(n8968), .Z(n8973) );
  OR U10852 ( .A(n8971), .B(n8970), .Z(n8972) );
  AND U10853 ( .A(n8973), .B(n8972), .Z(n9156) );
  XNOR U10854 ( .A(n9157), .B(n9156), .Z(n9158) );
  XNOR U10855 ( .A(n9159), .B(n9158), .Z(n9254) );
  XOR U10856 ( .A(n9255), .B(n9254), .Z(n9303) );
  NANDN U10857 ( .A(n8975), .B(n8974), .Z(n8979) );
  NANDN U10858 ( .A(n8977), .B(n8976), .Z(n8978) );
  AND U10859 ( .A(n8979), .B(n8978), .Z(n9111) );
  NAND U10860 ( .A(n8981), .B(n8980), .Z(n8985) );
  NANDN U10861 ( .A(n8983), .B(n8982), .Z(n8984) );
  AND U10862 ( .A(n8985), .B(n8984), .Z(n9109) );
  NANDN U10863 ( .A(n8987), .B(n8986), .Z(n8991) );
  OR U10864 ( .A(n8989), .B(n8988), .Z(n8990) );
  AND U10865 ( .A(n8991), .B(n8990), .Z(n9233) );
  XOR U10866 ( .A(n9233), .B(n9232), .Z(n9235) );
  NANDN U10867 ( .A(n8997), .B(n8996), .Z(n9001) );
  NANDN U10868 ( .A(n8999), .B(n8998), .Z(n9000) );
  AND U10869 ( .A(n9001), .B(n9000), .Z(n9234) );
  XOR U10870 ( .A(n9235), .B(n9234), .Z(n9207) );
  NANDN U10871 ( .A(n9003), .B(n9002), .Z(n9007) );
  NANDN U10872 ( .A(n9005), .B(n9004), .Z(n9006) );
  AND U10873 ( .A(n9007), .B(n9006), .Z(n9205) );
  XNOR U10874 ( .A(n9205), .B(n9204), .Z(n9206) );
  XOR U10875 ( .A(n9207), .B(n9206), .Z(n9243) );
  XNOR U10876 ( .A(n9215), .B(n9214), .Z(n9217) );
  IV U10877 ( .A(n9028), .Z(n9030) );
  NANDN U10878 ( .A(n9030), .B(n9029), .Z(n9034) );
  NAND U10879 ( .A(n9032), .B(n9031), .Z(n9033) );
  NAND U10880 ( .A(n9034), .B(n9033), .Z(n9195) );
  XOR U10881 ( .A(n9194), .B(n9195), .Z(n9197) );
  XOR U10882 ( .A(n9196), .B(n9197), .Z(n9189) );
  XOR U10883 ( .A(n9187), .B(n9186), .Z(n9188) );
  XNOR U10884 ( .A(n9189), .B(n9188), .Z(n9216) );
  XOR U10885 ( .A(n9217), .B(n9216), .Z(n9241) );
  NANDN U10886 ( .A(n9044), .B(n9043), .Z(n9048) );
  NAND U10887 ( .A(n9046), .B(n9045), .Z(n9047) );
  NAND U10888 ( .A(n9048), .B(n9047), .Z(n9240) );
  XNOR U10889 ( .A(n9241), .B(n9240), .Z(n9242) );
  XOR U10890 ( .A(n9243), .B(n9242), .Z(n9108) );
  XOR U10891 ( .A(n9109), .B(n9108), .Z(n9110) );
  XOR U10892 ( .A(n9111), .B(n9110), .Z(n9300) );
  NANDN U10893 ( .A(n9050), .B(n9049), .Z(n9054) );
  NAND U10894 ( .A(n9052), .B(n9051), .Z(n9053) );
  AND U10895 ( .A(n9054), .B(n9053), .Z(n9301) );
  XOR U10896 ( .A(n9300), .B(n9301), .Z(n9302) );
  XNOR U10897 ( .A(n9322), .B(n9321), .Z(n9323) );
  XNOR U10898 ( .A(n9324), .B(n9323), .Z(n9068) );
  XOR U10899 ( .A(n9069), .B(n9068), .Z(n9070) );
  XOR U10900 ( .A(n9071), .B(n9070), .Z(n9307) );
  NANDN U10901 ( .A(n9056), .B(n9055), .Z(n9060) );
  NAND U10902 ( .A(n9058), .B(n9057), .Z(n9059) );
  AND U10903 ( .A(n9060), .B(n9059), .Z(n9306) );
  XNOR U10904 ( .A(n9307), .B(n9306), .Z(n9061) );
  XNOR U10905 ( .A(n9308), .B(n9061), .Z(o[4]) );
  NAND U10906 ( .A(n9063), .B(n9062), .Z(n9067) );
  NANDN U10907 ( .A(n9065), .B(n9064), .Z(n9066) );
  NAND U10908 ( .A(n9067), .B(n9066), .Z(n9330) );
  NAND U10909 ( .A(n9069), .B(n9068), .Z(n9073) );
  NAND U10910 ( .A(n9071), .B(n9070), .Z(n9072) );
  NAND U10911 ( .A(n9073), .B(n9072), .Z(n9328) );
  NANDN U10912 ( .A(n9075), .B(n9074), .Z(n9079) );
  NAND U10913 ( .A(n9077), .B(n9076), .Z(n9078) );
  AND U10914 ( .A(n9079), .B(n9078), .Z(n9456) );
  NANDN U10915 ( .A(n9081), .B(n9080), .Z(n9085) );
  NANDN U10916 ( .A(n9083), .B(n9082), .Z(n9084) );
  AND U10917 ( .A(n9085), .B(n9084), .Z(n9443) );
  NAND U10918 ( .A(n9087), .B(n9086), .Z(n9091) );
  NAND U10919 ( .A(n9089), .B(n9088), .Z(n9090) );
  AND U10920 ( .A(n9091), .B(n9090), .Z(n9401) );
  NANDN U10921 ( .A(n9097), .B(n9096), .Z(n9101) );
  NANDN U10922 ( .A(n9099), .B(n9098), .Z(n9100) );
  AND U10923 ( .A(n9101), .B(n9100), .Z(n9399) );
  XOR U10924 ( .A(n9400), .B(n9399), .Z(n9402) );
  XOR U10925 ( .A(n9401), .B(n9402), .Z(n9442) );
  NANDN U10926 ( .A(n9103), .B(n9102), .Z(n9107) );
  NANDN U10927 ( .A(n9105), .B(n9104), .Z(n9106) );
  AND U10928 ( .A(n9107), .B(n9106), .Z(n9441) );
  XOR U10929 ( .A(n9442), .B(n9441), .Z(n9444) );
  XOR U10930 ( .A(n9443), .B(n9444), .Z(n9454) );
  NANDN U10931 ( .A(n9113), .B(n9112), .Z(n9117) );
  NANDN U10932 ( .A(n9115), .B(n9114), .Z(n9116) );
  AND U10933 ( .A(n9117), .B(n9116), .Z(n9448) );
  NANDN U10934 ( .A(n9119), .B(n9118), .Z(n9123) );
  NANDN U10935 ( .A(n9121), .B(n9120), .Z(n9122) );
  AND U10936 ( .A(n9123), .B(n9122), .Z(n9447) );
  XOR U10937 ( .A(n9448), .B(n9447), .Z(n9450) );
  XNOR U10938 ( .A(n9449), .B(n9450), .Z(n9453) );
  XNOR U10939 ( .A(n9456), .B(n9455), .Z(n9348) );
  NANDN U10940 ( .A(n9125), .B(n9124), .Z(n9129) );
  NANDN U10941 ( .A(n9127), .B(n9126), .Z(n9128) );
  NAND U10942 ( .A(n9129), .B(n9128), .Z(n9347) );
  NANDN U10943 ( .A(n9131), .B(n9130), .Z(n9135) );
  NANDN U10944 ( .A(n9133), .B(n9132), .Z(n9134) );
  NAND U10945 ( .A(n9135), .B(n9134), .Z(n9346) );
  XNOR U10946 ( .A(n9347), .B(n9346), .Z(n9349) );
  NANDN U10947 ( .A(n9141), .B(n9140), .Z(n9145) );
  OR U10948 ( .A(n9143), .B(n9142), .Z(n9144) );
  AND U10949 ( .A(n9145), .B(n9144), .Z(n9419) );
  NANDN U10950 ( .A(n9147), .B(n9146), .Z(n9151) );
  OR U10951 ( .A(n9149), .B(n9148), .Z(n9150) );
  AND U10952 ( .A(n9151), .B(n9150), .Z(n9418) );
  XOR U10953 ( .A(n9418), .B(n9417), .Z(n9420) );
  XOR U10954 ( .A(n9419), .B(n9420), .Z(n9430) );
  NANDN U10955 ( .A(n9157), .B(n9156), .Z(n9161) );
  NANDN U10956 ( .A(n9159), .B(n9158), .Z(n9160) );
  NAND U10957 ( .A(n9161), .B(n9160), .Z(n9429) );
  XOR U10958 ( .A(n9430), .B(n9429), .Z(n9432) );
  XOR U10959 ( .A(n9431), .B(n9432), .Z(n9438) );
  NAND U10960 ( .A(n9163), .B(n9162), .Z(n9167) );
  NAND U10961 ( .A(n9165), .B(n9164), .Z(n9166) );
  AND U10962 ( .A(n9167), .B(n9166), .Z(n9414) );
  ANDN U10963 ( .B(n9169), .A(n9168), .Z(n9170) );
  AND U10964 ( .A(n9171), .B(n9170), .Z(n9390) );
  NANDN U10965 ( .A(n9173), .B(n9172), .Z(n9177) );
  OR U10966 ( .A(n9175), .B(n9174), .Z(n9176) );
  NAND U10967 ( .A(n9177), .B(n9176), .Z(n9389) );
  XOR U10968 ( .A(n9390), .B(n9389), .Z(n9387) );
  XNOR U10969 ( .A(n9386), .B(n9385), .Z(n9388) );
  XOR U10970 ( .A(n9387), .B(n9388), .Z(n9413) );
  XOR U10971 ( .A(n9414), .B(n9413), .Z(n9416) );
  XOR U10972 ( .A(n9392), .B(n9391), .Z(n9394) );
  XOR U10973 ( .A(n9393), .B(n9394), .Z(n9415) );
  XOR U10974 ( .A(n9416), .B(n9415), .Z(n9375) );
  NANDN U10975 ( .A(n9199), .B(n9198), .Z(n9203) );
  NAND U10976 ( .A(n9201), .B(n9200), .Z(n9202) );
  AND U10977 ( .A(n9203), .B(n9202), .Z(n9373) );
  NANDN U10978 ( .A(n9205), .B(n9204), .Z(n9209) );
  NANDN U10979 ( .A(n9207), .B(n9206), .Z(n9208) );
  AND U10980 ( .A(n9209), .B(n9208), .Z(n9411) );
  NANDN U10981 ( .A(n9215), .B(n9214), .Z(n9219) );
  NAND U10982 ( .A(n9217), .B(n9216), .Z(n9218) );
  AND U10983 ( .A(n9219), .B(n9218), .Z(n9409) );
  XNOR U10984 ( .A(n9410), .B(n9409), .Z(n9412) );
  XOR U10985 ( .A(n9411), .B(n9412), .Z(n9374) );
  XOR U10986 ( .A(n9373), .B(n9374), .Z(n9376) );
  XOR U10987 ( .A(n9375), .B(n9376), .Z(n9436) );
  XOR U10988 ( .A(n9395), .B(n9396), .Z(n9398) );
  XOR U10989 ( .A(n9398), .B(n9397), .Z(n9381) );
  XOR U10990 ( .A(n9379), .B(n9380), .Z(n9382) );
  XOR U10991 ( .A(n9381), .B(n9382), .Z(n9425) );
  NANDN U10992 ( .A(n9241), .B(n9240), .Z(n9245) );
  NAND U10993 ( .A(n9243), .B(n9242), .Z(n9244) );
  AND U10994 ( .A(n9245), .B(n9244), .Z(n9424) );
  NANDN U10995 ( .A(n9247), .B(n9246), .Z(n9251) );
  NANDN U10996 ( .A(n9249), .B(n9248), .Z(n9250) );
  AND U10997 ( .A(n9251), .B(n9250), .Z(n9423) );
  XOR U10998 ( .A(n9424), .B(n9423), .Z(n9426) );
  XNOR U10999 ( .A(n9425), .B(n9426), .Z(n9435) );
  XNOR U11000 ( .A(n9436), .B(n9435), .Z(n9437) );
  XOR U11001 ( .A(n9438), .B(n9437), .Z(n9342) );
  NANDN U11002 ( .A(n9253), .B(n9252), .Z(n9257) );
  NAND U11003 ( .A(n9255), .B(n9254), .Z(n9256) );
  NAND U11004 ( .A(n9257), .B(n9256), .Z(n9340) );
  NANDN U11005 ( .A(n9259), .B(n9258), .Z(n9263) );
  NANDN U11006 ( .A(n9261), .B(n9260), .Z(n9262) );
  AND U11007 ( .A(n9263), .B(n9262), .Z(n9370) );
  NANDN U11008 ( .A(n9265), .B(n9264), .Z(n9269) );
  NANDN U11009 ( .A(n9267), .B(n9266), .Z(n9268) );
  AND U11010 ( .A(n9269), .B(n9268), .Z(n9368) );
  NANDN U11011 ( .A(n9271), .B(n9270), .Z(n9275) );
  OR U11012 ( .A(n9273), .B(n9272), .Z(n9274) );
  AND U11013 ( .A(n9275), .B(n9274), .Z(n9408) );
  NANDN U11014 ( .A(n9277), .B(n9276), .Z(n9281) );
  NAND U11015 ( .A(n9279), .B(n9278), .Z(n9280) );
  AND U11016 ( .A(n9281), .B(n9280), .Z(n9406) );
  NANDN U11017 ( .A(n9283), .B(n9282), .Z(n9287) );
  NAND U11018 ( .A(n9285), .B(n9284), .Z(n9286) );
  AND U11019 ( .A(n9287), .B(n9286), .Z(n9405) );
  XOR U11020 ( .A(n9406), .B(n9405), .Z(n9407) );
  XOR U11021 ( .A(n9408), .B(n9407), .Z(n9367) );
  XNOR U11022 ( .A(n9368), .B(n9367), .Z(n9369) );
  XOR U11023 ( .A(n9370), .B(n9369), .Z(n9341) );
  XNOR U11024 ( .A(n9340), .B(n9341), .Z(n9343) );
  NAND U11025 ( .A(n9289), .B(n9288), .Z(n9293) );
  NAND U11026 ( .A(n9291), .B(n9290), .Z(n9292) );
  NAND U11027 ( .A(n9293), .B(n9292), .Z(n9354) );
  NANDN U11028 ( .A(n9295), .B(n9294), .Z(n9299) );
  NAND U11029 ( .A(n9297), .B(n9296), .Z(n9298) );
  AND U11030 ( .A(n9299), .B(n9298), .Z(n9353) );
  NAND U11031 ( .A(n9301), .B(n9300), .Z(n9305) );
  NANDN U11032 ( .A(n9303), .B(n9302), .Z(n9304) );
  AND U11033 ( .A(n9305), .B(n9304), .Z(n9352) );
  XOR U11034 ( .A(n9353), .B(n9352), .Z(n9355) );
  XNOR U11035 ( .A(n9354), .B(n9355), .Z(n9361) );
  XOR U11036 ( .A(n9362), .B(n9361), .Z(n9364) );
  XNOR U11037 ( .A(n9363), .B(n9364), .Z(n9329) );
  XOR U11038 ( .A(n9330), .B(n9331), .Z(n9360) );
  NANDN U11039 ( .A(n9310), .B(n9309), .Z(n9314) );
  NAND U11040 ( .A(n9312), .B(n9311), .Z(n9313) );
  AND U11041 ( .A(n9314), .B(n9313), .Z(n9335) );
  NAND U11042 ( .A(n9316), .B(n9315), .Z(n9320) );
  NANDN U11043 ( .A(n9318), .B(n9317), .Z(n9319) );
  AND U11044 ( .A(n9320), .B(n9319), .Z(n9334) );
  XOR U11045 ( .A(n9335), .B(n9334), .Z(n9337) );
  NANDN U11046 ( .A(n9322), .B(n9321), .Z(n9326) );
  NANDN U11047 ( .A(n9324), .B(n9323), .Z(n9325) );
  AND U11048 ( .A(n9326), .B(n9325), .Z(n9336) );
  XOR U11049 ( .A(n9337), .B(n9336), .Z(n9358) );
  XOR U11050 ( .A(n9359), .B(n9358), .Z(n9327) );
  XNOR U11051 ( .A(n9360), .B(n9327), .Z(o[5]) );
  NANDN U11052 ( .A(n9329), .B(n9328), .Z(n9333) );
  NANDN U11053 ( .A(n9331), .B(n9330), .Z(n9332) );
  NAND U11054 ( .A(n9333), .B(n9332), .Z(n9462) );
  NAND U11055 ( .A(n9335), .B(n9334), .Z(n9339) );
  NAND U11056 ( .A(n9337), .B(n9336), .Z(n9338) );
  AND U11057 ( .A(n9339), .B(n9338), .Z(n9461) );
  NAND U11058 ( .A(n9341), .B(n9340), .Z(n9345) );
  NANDN U11059 ( .A(n9343), .B(n9342), .Z(n9344) );
  AND U11060 ( .A(n9345), .B(n9344), .Z(n9520) );
  NAND U11061 ( .A(n9347), .B(n9346), .Z(n9351) );
  NANDN U11062 ( .A(n9349), .B(n9348), .Z(n9350) );
  AND U11063 ( .A(n9351), .B(n9350), .Z(n9517) );
  NAND U11064 ( .A(n9353), .B(n9352), .Z(n9357) );
  NAND U11065 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U11066 ( .A(n9357), .B(n9356), .Z(n9518) );
  XOR U11067 ( .A(n9520), .B(n9519), .Z(n9460) );
  XOR U11068 ( .A(n9461), .B(n9460), .Z(n9463) );
  XNOR U11069 ( .A(n9462), .B(n9463), .Z(n9525) );
  NAND U11070 ( .A(n9362), .B(n9361), .Z(n9366) );
  NAND U11071 ( .A(n9364), .B(n9363), .Z(n9365) );
  AND U11072 ( .A(n9366), .B(n9365), .Z(n9469) );
  NANDN U11073 ( .A(n9368), .B(n9367), .Z(n9372) );
  NAND U11074 ( .A(n9370), .B(n9369), .Z(n9371) );
  NAND U11075 ( .A(n9372), .B(n9371), .Z(n9472) );
  NANDN U11076 ( .A(n9374), .B(n9373), .Z(n9378) );
  OR U11077 ( .A(n9376), .B(n9375), .Z(n9377) );
  NAND U11078 ( .A(n9378), .B(n9377), .Z(n9499) );
  NANDN U11079 ( .A(n9380), .B(n9379), .Z(n9384) );
  OR U11080 ( .A(n9382), .B(n9381), .Z(n9383) );
  AND U11081 ( .A(n9384), .B(n9383), .Z(n9488) );
  AND U11082 ( .A(n9390), .B(n9389), .Z(n9493) );
  XNOR U11083 ( .A(n9493), .B(n9492), .Z(n9494) );
  XOR U11084 ( .A(n9495), .B(n9494), .Z(n9487) );
  XOR U11085 ( .A(n9487), .B(n9486), .Z(n9489) );
  XNOR U11086 ( .A(n9488), .B(n9489), .Z(n9498) );
  XOR U11087 ( .A(n9499), .B(n9498), .Z(n9500) );
  NANDN U11088 ( .A(n9400), .B(n9399), .Z(n9404) );
  OR U11089 ( .A(n9402), .B(n9401), .Z(n9403) );
  AND U11090 ( .A(n9404), .B(n9403), .Z(n9501) );
  XOR U11091 ( .A(n9500), .B(n9501), .Z(n9506) );
  XOR U11092 ( .A(n9480), .B(n9481), .Z(n9483) );
  NANDN U11093 ( .A(n9418), .B(n9417), .Z(n9422) );
  OR U11094 ( .A(n9420), .B(n9419), .Z(n9421) );
  AND U11095 ( .A(n9422), .B(n9421), .Z(n9482) );
  XOR U11096 ( .A(n9483), .B(n9482), .Z(n9477) );
  NANDN U11097 ( .A(n9424), .B(n9423), .Z(n9428) );
  OR U11098 ( .A(n9426), .B(n9425), .Z(n9427) );
  AND U11099 ( .A(n9428), .B(n9427), .Z(n9476) );
  XNOR U11100 ( .A(n9477), .B(n9476), .Z(n9479) );
  NANDN U11101 ( .A(n9430), .B(n9429), .Z(n9434) );
  OR U11102 ( .A(n9432), .B(n9431), .Z(n9433) );
  AND U11103 ( .A(n9434), .B(n9433), .Z(n9478) );
  XOR U11104 ( .A(n9479), .B(n9478), .Z(n9505) );
  XOR U11105 ( .A(n9504), .B(n9505), .Z(n9507) );
  XNOR U11106 ( .A(n9506), .B(n9507), .Z(n9473) );
  XOR U11107 ( .A(n9472), .B(n9473), .Z(n9475) );
  NANDN U11108 ( .A(n9436), .B(n9435), .Z(n9440) );
  NANDN U11109 ( .A(n9438), .B(n9437), .Z(n9439) );
  AND U11110 ( .A(n9440), .B(n9439), .Z(n9513) );
  NANDN U11111 ( .A(n9442), .B(n9441), .Z(n9446) );
  OR U11112 ( .A(n9444), .B(n9443), .Z(n9445) );
  NAND U11113 ( .A(n9446), .B(n9445), .Z(n9510) );
  NANDN U11114 ( .A(n9448), .B(n9447), .Z(n9452) );
  OR U11115 ( .A(n9450), .B(n9449), .Z(n9451) );
  NAND U11116 ( .A(n9452), .B(n9451), .Z(n9511) );
  XNOR U11117 ( .A(n9510), .B(n9511), .Z(n9514) );
  XNOR U11118 ( .A(n9513), .B(n9514), .Z(n9474) );
  XOR U11119 ( .A(n9475), .B(n9474), .Z(n9467) );
  NANDN U11120 ( .A(n9454), .B(n9453), .Z(n9458) );
  NAND U11121 ( .A(n9456), .B(n9455), .Z(n9457) );
  NAND U11122 ( .A(n9458), .B(n9457), .Z(n9466) );
  XNOR U11123 ( .A(n9524), .B(n9523), .Z(n9459) );
  XNOR U11124 ( .A(n9525), .B(n9459), .Z(o[6]) );
  NAND U11125 ( .A(n9461), .B(n9460), .Z(n9465) );
  NAND U11126 ( .A(n9463), .B(n9462), .Z(n9464) );
  AND U11127 ( .A(n9465), .B(n9464), .Z(n9547) );
  NANDN U11128 ( .A(n9467), .B(n9466), .Z(n9471) );
  NANDN U11129 ( .A(n9469), .B(n9468), .Z(n9470) );
  AND U11130 ( .A(n9471), .B(n9470), .Z(n9550) );
  NAND U11131 ( .A(n9481), .B(n9480), .Z(n9485) );
  NAND U11132 ( .A(n9483), .B(n9482), .Z(n9484) );
  NAND U11133 ( .A(n9485), .B(n9484), .Z(n9540) );
  NANDN U11134 ( .A(n9487), .B(n9486), .Z(n9491) );
  NANDN U11135 ( .A(n9489), .B(n9488), .Z(n9490) );
  NAND U11136 ( .A(n9491), .B(n9490), .Z(n9535) );
  NANDN U11137 ( .A(n9493), .B(n9492), .Z(n9497) );
  NAND U11138 ( .A(n9495), .B(n9494), .Z(n9496) );
  NAND U11139 ( .A(n9497), .B(n9496), .Z(n9536) );
  XOR U11140 ( .A(n9535), .B(n9536), .Z(n9539) );
  XOR U11141 ( .A(n9540), .B(n9539), .Z(n9537) );
  XOR U11142 ( .A(n9538), .B(n9537), .Z(n9533) );
  NAND U11143 ( .A(n9499), .B(n9498), .Z(n9503) );
  NAND U11144 ( .A(n9501), .B(n9500), .Z(n9502) );
  AND U11145 ( .A(n9503), .B(n9502), .Z(n9532) );
  NANDN U11146 ( .A(n9505), .B(n9504), .Z(n9509) );
  NANDN U11147 ( .A(n9507), .B(n9506), .Z(n9508) );
  AND U11148 ( .A(n9509), .B(n9508), .Z(n9531) );
  XOR U11149 ( .A(n9532), .B(n9531), .Z(n9534) );
  XOR U11150 ( .A(n9533), .B(n9534), .Z(n9528) );
  IV U11151 ( .A(n9510), .Z(n9512) );
  NANDN U11152 ( .A(n9512), .B(n9511), .Z(n9516) );
  NANDN U11153 ( .A(n9514), .B(n9513), .Z(n9515) );
  AND U11154 ( .A(n9516), .B(n9515), .Z(n9527) );
  XOR U11155 ( .A(n9528), .B(n9527), .Z(n9529) );
  XOR U11156 ( .A(n9530), .B(n9529), .Z(n9549) );
  NANDN U11157 ( .A(n9518), .B(n9517), .Z(n9522) );
  NAND U11158 ( .A(n9520), .B(n9519), .Z(n9521) );
  AND U11159 ( .A(n9522), .B(n9521), .Z(n9548) );
  XNOR U11160 ( .A(n9550), .B(n9551), .Z(n9546) );
  XNOR U11161 ( .A(n9546), .B(n9545), .Z(n9526) );
  XNOR U11162 ( .A(n9547), .B(n9526), .Z(o[7]) );
  IV U11163 ( .A(n9542), .Z(n9559) );
  ANDN U11164 ( .B(n9538), .A(n9537), .Z(n9558) );
  XOR U11165 ( .A(n9559), .B(n9558), .Z(n9544) );
  ANDN U11166 ( .B(n9540), .A(n9539), .Z(n9541) );
  NANDN U11167 ( .A(n9542), .B(n9541), .Z(n9543) );
  NAND U11168 ( .A(n9544), .B(n9543), .Z(n9561) );
  XOR U11169 ( .A(n9560), .B(n9561), .Z(n9563) );
  XOR U11170 ( .A(n9562), .B(n9563), .Z(n9557) );
  NANDN U11171 ( .A(n9549), .B(n9548), .Z(n9553) );
  NANDN U11172 ( .A(n9551), .B(n9550), .Z(n9552) );
  AND U11173 ( .A(n9553), .B(n9552), .Z(n9555) );
  XOR U11174 ( .A(n9556), .B(n9555), .Z(n9554) );
  XNOR U11175 ( .A(n9557), .B(n9554), .Z(o[8]) );
  NANDN U11176 ( .A(n9559), .B(n9558), .Z(n9567) );
  XNOR U11177 ( .A(n9566), .B(n9567), .Z(n9565) );
  XOR U11178 ( .A(n9565), .B(n9564), .Z(o[9]) );
endmodule

