
module modexp_1_N_N4_CC1 ( clk, rst, m, e, n, c );
  input [3:0] m;
  input [3:0] e;
  input [3:0] n;
  output [3:0] c;
  input clk, rst;
  wire   \cin[1][3] , \cin[1][2] , \cin[1][1] ,
         \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 , n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554;
  assign \cin[1][3]  = m[3];
  assign \cin[1][2]  = m[2];
  assign \cin[1][1]  = m[1];
  assign \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4  = m[0];

  NANDN U778 ( .A(n810), .B(n[1]), .Z(n494) );
  NAND U779 ( .A(n810), .B(n792), .Z(n495) );
  NANDN U780 ( .A(n807), .B(n495), .Z(n496) );
  NAND U781 ( .A(n494), .B(n496), .Z(n814) );
  XOR U782 ( .A(\cin[1][3] ), .B(n1103), .Z(n497) );
  ANDN U783 ( .B(n497), .A(n1100), .Z(n498) );
  NAND U784 ( .A(n1103), .B(\cin[1][3] ), .Z(n499) );
  NANDN U785 ( .A(n498), .B(n499), .Z(n500) );
  ANDN U786 ( .B(n500), .A(n1349), .Z(n1129) );
  XOR U787 ( .A(n[2]), .B(n1678), .Z(n501) );
  ANDN U788 ( .B(n501), .A(n1707), .Z(n502) );
  XNOR U789 ( .A(n1679), .B(n502), .Z(n1697) );
  XNOR U790 ( .A(\cin[1][3] ), .B(n1289), .Z(n503) );
  AND U791 ( .A(n1286), .B(n503), .Z(n504) );
  NANDN U792 ( .A(n1289), .B(\cin[1][3] ), .Z(n505) );
  NANDN U793 ( .A(n504), .B(n505), .Z(n506) );
  AND U794 ( .A(n1294), .B(n506), .Z(n1301) );
  NAND U795 ( .A(n[0]), .B(n2314), .Z(n507) );
  ANDN U796 ( .B(n2292), .A(n[0]), .Z(n508) );
  XNOR U797 ( .A(n2291), .B(n507), .Z(n509) );
  NANDN U798 ( .A(n508), .B(n509), .Z(n2302) );
  XOR U799 ( .A(\cin[1][3] ), .B(n2333), .Z(n510) );
  ANDN U800 ( .B(n510), .A(n2330), .Z(n511) );
  NAND U801 ( .A(n2333), .B(\cin[1][3] ), .Z(n512) );
  NANDN U802 ( .A(n511), .B(n512), .Z(n513) );
  ANDN U803 ( .B(n513), .A(n2536), .Z(n2357) );
  OR U804 ( .A(n1632), .B(n2233), .Z(n514) );
  NANDN U805 ( .A(n[1]), .B(n1653), .Z(n515) );
  AND U806 ( .A(n514), .B(n515), .Z(n516) );
  NAND U807 ( .A(n1648), .B(n[2]), .Z(n517) );
  ANDN U808 ( .B(n517), .A(n1630), .Z(n518) );
  XOR U809 ( .A(n1648), .B(n[2]), .Z(n519) );
  NAND U810 ( .A(n519), .B(n516), .Z(n520) );
  AND U811 ( .A(n518), .B(n520), .Z(n521) );
  ANDN U812 ( .B(n1631), .A(n1636), .Z(n522) );
  ANDN U813 ( .B(n522), .A(n521), .Z(n523) );
  NANDN U814 ( .A(n1639), .B(n523), .Z(n1651) );
  NANDN U815 ( .A(n2167), .B(n[3]), .Z(n524) );
  XNOR U816 ( .A(n2167), .B(n[3]), .Z(n525) );
  NAND U817 ( .A(n2164), .B(n525), .Z(n526) );
  NAND U818 ( .A(n524), .B(n526), .Z(n527) );
  XNOR U819 ( .A(n2161), .B(n527), .Z(n528) );
  NAND U820 ( .A(n2178), .B(n528), .Z(n2220) );
  XNOR U821 ( .A(n2224), .B(n2223), .Z(n529) );
  ANDN U822 ( .B(n529), .A(n2235), .Z(n530) );
  XNOR U823 ( .A(n2225), .B(n530), .Z(n2264) );
  NAND U824 ( .A(n2488), .B(n2500), .Z(n531) );
  NANDN U825 ( .A(n[1]), .B(n2517), .Z(n532) );
  NAND U826 ( .A(n531), .B(n532), .Z(n533) );
  NAND U827 ( .A(n2522), .B(n533), .Z(n534) );
  XOR U828 ( .A(n2522), .B(n533), .Z(n535) );
  NAND U829 ( .A(n535), .B(n793), .Z(n536) );
  NAND U830 ( .A(n534), .B(n536), .Z(n537) );
  ANDN U831 ( .B(n537), .A(n2501), .Z(n538) );
  ANDN U832 ( .B(n2504), .A(n2509), .Z(n539) );
  ANDN U833 ( .B(n539), .A(n538), .Z(n540) );
  ANDN U834 ( .B(n540), .A(n2502), .Z(n2520) );
  XOR U835 ( .A(n[2]), .B(n820), .Z(n541) );
  NANDN U836 ( .A(n823), .B(n541), .Z(n542) );
  NAND U837 ( .A(n[2]), .B(n820), .Z(n543) );
  AND U838 ( .A(n542), .B(n543), .Z(n831) );
  NAND U839 ( .A(n1676), .B(n[1]), .Z(n544) );
  XOR U840 ( .A(n1676), .B(n[1]), .Z(n545) );
  NAND U841 ( .A(n545), .B(n1677), .Z(n546) );
  NAND U842 ( .A(n544), .B(n546), .Z(n1678) );
  NOR U843 ( .A(n[1]), .B(n1014), .Z(n547) );
  OR U844 ( .A(n2488), .B(n1026), .Z(n548) );
  AND U845 ( .A(n547), .B(n548), .Z(n549) );
  OR U846 ( .A(n1015), .B(n549), .Z(n550) );
  ANDN U847 ( .B(n550), .A(n1018), .Z(n551) );
  ANDN U848 ( .B(n1021), .A(n1017), .Z(n552) );
  ANDN U849 ( .B(n552), .A(n1022), .Z(n553) );
  NANDN U850 ( .A(n551), .B(n553), .Z(n1033) );
  ANDN U851 ( .B(n2191), .A(n2051), .Z(n2053) );
  XOR U852 ( .A(n[2]), .B(n2286), .Z(n554) );
  NAND U853 ( .A(n2287), .B(n554), .Z(n555) );
  XNOR U854 ( .A(\cin[1][2] ), .B(n555), .Z(n556) );
  NAND U855 ( .A(\cin[1][2] ), .B(n2552), .Z(n557) );
  AND U856 ( .A(n556), .B(n557), .Z(n2316) );
  ANDN U857 ( .B(n[0]), .A(n2102), .Z(n2103) );
  ANDN U858 ( .B(n[0]), .A(n1655), .Z(n1779) );
  OR U859 ( .A(n2235), .B(n2233), .Z(n558) );
  NANDN U860 ( .A(n[1]), .B(n2249), .Z(n559) );
  AND U861 ( .A(n558), .B(n559), .Z(n560) );
  NAND U862 ( .A(n2256), .B(n[2]), .Z(n561) );
  ANDN U863 ( .B(n561), .A(n2239), .Z(n562) );
  XOR U864 ( .A(n2256), .B(n[2]), .Z(n563) );
  NAND U865 ( .A(n563), .B(n560), .Z(n564) );
  AND U866 ( .A(n562), .B(n564), .Z(n565) );
  AND U867 ( .A(n2245), .B(n2243), .Z(n566) );
  ANDN U868 ( .B(n566), .A(n565), .Z(n567) );
  NANDN U869 ( .A(n2241), .B(n567), .Z(n2262) );
  ANDN U870 ( .B(n[0]), .A(n2524), .Z(n2529) );
  OR U871 ( .A(n[0]), .B(n871), .Z(n568) );
  NANDN U872 ( .A(n[1]), .B(n876), .Z(n569) );
  AND U873 ( .A(n568), .B(n569), .Z(n570) );
  NANDN U874 ( .A(n570), .B(n849), .Z(n571) );
  NANDN U875 ( .A(n850), .B(n571), .Z(n572) );
  NAND U876 ( .A(n852), .B(n572), .Z(n573) );
  NANDN U877 ( .A(n862), .B(n863), .Z(n574) );
  OR U878 ( .A(n573), .B(n857), .Z(n575) );
  ANDN U879 ( .B(n575), .A(n574), .Z(n576) );
  XOR U880 ( .A(n573), .B(n857), .Z(n577) );
  NANDN U881 ( .A(n[3]), .B(n577), .Z(n578) );
  NAND U882 ( .A(n576), .B(n578), .Z(n874) );
  NAND U883 ( .A(n[0]), .B(n1429), .Z(n579) );
  XNOR U884 ( .A(n1416), .B(n579), .Z(n580) );
  NANDN U885 ( .A(n[0]), .B(n1415), .Z(n581) );
  NAND U886 ( .A(n580), .B(n581), .Z(n1430) );
  XNOR U887 ( .A(\cin[1][3] ), .B(n1007), .Z(n582) );
  AND U888 ( .A(n1004), .B(n582), .Z(n583) );
  NANDN U889 ( .A(n1007), .B(\cin[1][3] ), .Z(n584) );
  NANDN U890 ( .A(n583), .B(n584), .Z(n585) );
  AND U891 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .B(
        n585), .Z(n1003) );
  NAND U892 ( .A(n[2]), .B(n1678), .Z(n586) );
  ANDN U893 ( .B(n586), .A(n[3]), .Z(n587) );
  XOR U894 ( .A(n[2]), .B(n1678), .Z(n588) );
  NAND U895 ( .A(n588), .B(n1679), .Z(n589) );
  AND U896 ( .A(n587), .B(n589), .Z(n590) );
  AND U897 ( .A(\cin[1][3] ), .B(n1975), .Z(n591) );
  NANDN U898 ( .A(n590), .B(n2275), .Z(n592) );
  AND U899 ( .A(n591), .B(n592), .Z(n1712) );
  XNOR U900 ( .A(n1026), .B(n[1]), .Z(n593) );
  NANDN U901 ( .A(n2276), .B(n593), .Z(n594) );
  NANDN U902 ( .A(n1026), .B(n[1]), .Z(n595) );
  AND U903 ( .A(n594), .B(n595), .Z(n1027) );
  ANDN U904 ( .B(n1532), .A(n1531), .Z(n596) );
  XNOR U905 ( .A(n1530), .B(n596), .Z(n597) );
  NANDN U906 ( .A(n1529), .B(n1528), .Z(n598) );
  ANDN U907 ( .B(n598), .A(n1521), .Z(n599) );
  XNOR U908 ( .A(n597), .B(n599), .Z(n1559) );
  NANDN U909 ( .A(n[1]), .B(n1329), .Z(n600) );
  NANDN U910 ( .A(n1310), .B(n2488), .Z(n601) );
  AND U911 ( .A(n600), .B(n601), .Z(n602) );
  NOR U912 ( .A(n1312), .B(n1317), .Z(n603) );
  OR U913 ( .A(n1313), .B(n602), .Z(n604) );
  AND U914 ( .A(n603), .B(n604), .Z(n605) );
  ANDN U915 ( .B(n1319), .A(n1320), .Z(n606) );
  OR U916 ( .A(n605), .B(n1315), .Z(n607) );
  NAND U917 ( .A(n606), .B(n607), .Z(n1332) );
  OR U918 ( .A(n[3]), .B(n2026), .Z(n608) );
  NAND U919 ( .A(n2014), .B(n608), .Z(n609) );
  AND U920 ( .A(n2191), .B(n609), .Z(n2024) );
  XOR U921 ( .A(n[2]), .B(n2111), .Z(n610) );
  NANDN U922 ( .A(n2114), .B(n610), .Z(n611) );
  NAND U923 ( .A(n[2]), .B(n2111), .Z(n612) );
  AND U924 ( .A(n611), .B(n612), .Z(n2124) );
  XOR U925 ( .A(n[2]), .B(n2312), .Z(n613) );
  NANDN U926 ( .A(n2316), .B(n613), .Z(n614) );
  NAND U927 ( .A(n[2]), .B(n2312), .Z(n615) );
  AND U928 ( .A(n614), .B(n615), .Z(n2324) );
  NOR U929 ( .A(n1832), .B(n1887), .Z(n1863) );
  NANDN U930 ( .A(n1913), .B(n[1]), .Z(n1917) );
  XNOR U931 ( .A(\cin[1][3] ), .B(n1891), .Z(n616) );
  AND U932 ( .A(n1888), .B(n616), .Z(n617) );
  NANDN U933 ( .A(n1891), .B(\cin[1][3] ), .Z(n618) );
  NANDN U934 ( .A(n617), .B(n618), .Z(n619) );
  AND U935 ( .A(n1950), .B(n619), .Z(n1905) );
  ANDN U936 ( .B(n[0]), .A(n1946), .Z(n1960) );
  XOR U937 ( .A(n[1]), .B(n2455), .Z(n620) );
  NANDN U938 ( .A(n2458), .B(n620), .Z(n621) );
  NAND U939 ( .A(n[1]), .B(n2455), .Z(n622) );
  AND U940 ( .A(n621), .B(n622), .Z(n2451) );
  NANDN U941 ( .A(n2270), .B(n2268), .Z(n623) );
  ANDN U942 ( .B(n623), .A(n2269), .Z(n624) );
  XNOR U943 ( .A(n2268), .B(n2270), .Z(n625) );
  NANDN U944 ( .A(n[3]), .B(n625), .Z(n626) );
  NAND U945 ( .A(n624), .B(n626), .Z(n2368) );
  NAND U946 ( .A(n2518), .B(n2522), .Z(n627) );
  XOR U947 ( .A(n2518), .B(n2522), .Z(n628) );
  NANDN U948 ( .A(n[2]), .B(n628), .Z(n629) );
  NAND U949 ( .A(n627), .B(n629), .Z(n2510) );
  NAND U950 ( .A(n[1]), .B(n2529), .Z(n630) );
  XOR U951 ( .A(n[1]), .B(n2529), .Z(n631) );
  NANDN U952 ( .A(n2532), .B(n631), .Z(n632) );
  NAND U953 ( .A(n630), .B(n632), .Z(n2537) );
  OR U954 ( .A(n839), .B(\cin[1][2] ), .Z(n633) );
  ANDN U955 ( .B(\cin[1][3] ), .A(n839), .Z(n634) );
  XNOR U956 ( .A(n836), .B(n634), .Z(n635) );
  NAND U957 ( .A(\cin[1][2] ), .B(n635), .Z(n636) );
  NAND U958 ( .A(n633), .B(n636), .Z(n857) );
  NAND U959 ( .A(n[2]), .B(n1076), .Z(n637) );
  XOR U960 ( .A(n[2]), .B(n1076), .Z(n638) );
  NANDN U961 ( .A(n1079), .B(n638), .Z(n639) );
  NAND U962 ( .A(n637), .B(n639), .Z(n1095) );
  NANDN U963 ( .A(n1144), .B(n[1]), .Z(n1122) );
  XOR U964 ( .A(n[1]), .B(n989), .Z(n640) );
  NAND U965 ( .A(n640), .B(n992), .Z(n641) );
  NAND U966 ( .A(n[1]), .B(n989), .Z(n642) );
  AND U967 ( .A(n641), .B(n642), .Z(n983) );
  NAND U968 ( .A(n1429), .B(n[2]), .Z(n643) );
  AND U969 ( .A(n1426), .B(n643), .Z(n1447) );
  ANDN U970 ( .B(n[0]), .A(n1487), .Z(n1494) );
  XOR U971 ( .A(n[2]), .B(n1693), .Z(n644) );
  NANDN U972 ( .A(n1697), .B(n644), .Z(n645) );
  NAND U973 ( .A(n[2]), .B(n1693), .Z(n646) );
  AND U974 ( .A(n645), .B(n646), .Z(n1708) );
  ANDN U975 ( .B(n1003), .A(n1002), .Z(n647) );
  XNOR U976 ( .A(n1001), .B(n647), .Z(n648) );
  NAND U977 ( .A(n1000), .B(n999), .Z(n649) );
  ANDN U978 ( .B(n649), .A(n986), .Z(n650) );
  XNOR U979 ( .A(n648), .B(n650), .Z(n1022) );
  NOR U980 ( .A(n792), .B(n1751), .Z(n1732) );
  XOR U981 ( .A(n[1]), .B(n1180), .Z(n651) );
  NANDN U982 ( .A(n1184), .B(n651), .Z(n652) );
  NAND U983 ( .A(n[1]), .B(n1180), .Z(n653) );
  AND U984 ( .A(n652), .B(n653), .Z(n1090) );
  XOR U985 ( .A(n[2]), .B(n1763), .Z(n654) );
  NAND U986 ( .A(n654), .B(n1766), .Z(n655) );
  NAND U987 ( .A(n[2]), .B(n1763), .Z(n656) );
  AND U988 ( .A(n655), .B(n656), .Z(n1792) );
  NAND U989 ( .A(n[1]), .B(n1342), .Z(n657) );
  XOR U990 ( .A(n[1]), .B(n1342), .Z(n658) );
  NANDN U991 ( .A(n1345), .B(n658), .Z(n659) );
  NAND U992 ( .A(n657), .B(n659), .Z(n1351) );
  NAND U993 ( .A(n[2]), .B(n1603), .Z(n660) );
  ANDN U994 ( .B(n660), .A(n1579), .Z(n1602) );
  XOR U995 ( .A(n2031), .B(n2030), .Z(n2036) );
  XOR U996 ( .A(n[1]), .B(n2103), .Z(n661) );
  NANDN U997 ( .A(n2125), .B(n661), .Z(n662) );
  XNOR U998 ( .A(n2104), .B(n662), .Z(n2118) );
  NAND U999 ( .A(n[1]), .B(n2362), .Z(n663) );
  XOR U1000 ( .A(n[1]), .B(n2362), .Z(n664) );
  NANDN U1001 ( .A(n2365), .B(n664), .Z(n665) );
  NAND U1002 ( .A(n663), .B(n665), .Z(n2375) );
  XOR U1003 ( .A(n[2]), .B(n2350), .Z(n666) );
  NANDN U1004 ( .A(n2349), .B(n666), .Z(n667) );
  NAND U1005 ( .A(n[2]), .B(n2350), .Z(n668) );
  AND U1006 ( .A(n667), .B(n668), .Z(n2354) );
  OR U1007 ( .A(n[3]), .B(n1836), .Z(n669) );
  ANDN U1008 ( .B(n669), .A(n1838), .Z(n670) );
  XOR U1009 ( .A(n[3]), .B(n1836), .Z(n671) );
  NANDN U1010 ( .A(n1833), .B(n671), .Z(n672) );
  NAND U1011 ( .A(n670), .B(n672), .Z(n673) );
  XNOR U1012 ( .A(n1831), .B(n673), .Z(n1887) );
  XOR U1013 ( .A(n[2]), .B(n1664), .Z(n674) );
  NAND U1014 ( .A(n[2]), .B(n1664), .Z(n675) );
  NANDN U1015 ( .A(n1662), .B(n674), .Z(n676) );
  NAND U1016 ( .A(n675), .B(n676), .Z(n677) );
  OR U1017 ( .A(n677), .B(n1658), .Z(n678) );
  AND U1018 ( .A(n1656), .B(n678), .Z(n679) );
  XOR U1019 ( .A(n677), .B(n1658), .Z(n680) );
  NANDN U1020 ( .A(n[3]), .B(n680), .Z(n681) );
  NAND U1021 ( .A(n679), .B(n681), .Z(n1781) );
  NAND U1022 ( .A(n[1]), .B(n1960), .Z(n682) );
  XOR U1023 ( .A(n[1]), .B(n1960), .Z(n683) );
  NANDN U1024 ( .A(n1962), .B(n683), .Z(n684) );
  NAND U1025 ( .A(n682), .B(n684), .Z(n1971) );
  ANDN U1026 ( .B(n[0]), .A(n2197), .Z(n2192) );
  NAND U1027 ( .A(n2210), .B(n[2]), .Z(n685) );
  AND U1028 ( .A(n2189), .B(n685), .Z(n2209) );
  XOR U1029 ( .A(n2451), .B(n2454), .Z(n686) );
  NANDN U1030 ( .A(n[2]), .B(n686), .Z(n687) );
  NAND U1031 ( .A(n2451), .B(n2454), .Z(n688) );
  AND U1032 ( .A(n687), .B(n688), .Z(n2474) );
  NANDN U1033 ( .A(n[3]), .B(n2545), .Z(n689) );
  ANDN U1034 ( .B(n689), .A(n2548), .Z(n690) );
  XNOR U1035 ( .A(n2545), .B(n[3]), .Z(n691) );
  NAND U1036 ( .A(n691), .B(n2546), .Z(n692) );
  NAND U1037 ( .A(n690), .B(n692), .Z(n2539) );
  XNOR U1038 ( .A(n2270), .B(n2268), .Z(n693) );
  XNOR U1039 ( .A(n[3]), .B(n693), .Z(n694) );
  NANDN U1040 ( .A(n2269), .B(n2270), .Z(n695) );
  NAND U1041 ( .A(n694), .B(n695), .Z(n2552) );
  NAND U1042 ( .A(n[2]), .B(n840), .Z(n696) );
  ANDN U1043 ( .B(n696), .A(n[3]), .Z(n697) );
  XOR U1044 ( .A(n[2]), .B(n840), .Z(n698) );
  NAND U1045 ( .A(n698), .B(n814), .Z(n699) );
  AND U1046 ( .A(n697), .B(n699), .Z(n700) );
  OR U1047 ( .A(n815), .B(n700), .Z(n701) );
  AND U1048 ( .A(\cin[1][3] ), .B(n701), .Z(n835) );
  NAND U1049 ( .A(n[1]), .B(n1080), .Z(n702) );
  XOR U1050 ( .A(n[1]), .B(n1080), .Z(n703) );
  NANDN U1051 ( .A(n1083), .B(n703), .Z(n704) );
  NAND U1052 ( .A(n702), .B(n704), .Z(n1076) );
  ANDN U1053 ( .B(n[3]), .A(n909), .Z(n907) );
  NAND U1054 ( .A(n1388), .B(n[1]), .Z(n705) );
  XOR U1055 ( .A(n1388), .B(n[1]), .Z(n706) );
  NAND U1056 ( .A(n706), .B(n1389), .Z(n707) );
  NAND U1057 ( .A(n705), .B(n707), .Z(n1393) );
  XNOR U1058 ( .A(\cin[1][3] ), .B(n915), .Z(n708) );
  AND U1059 ( .A(n912), .B(n708), .Z(n709) );
  NANDN U1060 ( .A(n915), .B(\cin[1][3] ), .Z(n710) );
  NANDN U1061 ( .A(n709), .B(n710), .Z(n711) );
  AND U1062 ( .A(\cin[1][1] ), .B(n711), .Z(n932) );
  OR U1063 ( .A(n1131), .B(n1126), .Z(n712) );
  ANDN U1064 ( .B(n712), .A(n1127), .Z(n713) );
  XNOR U1065 ( .A(n1129), .B(n1128), .Z(n714) );
  XNOR U1066 ( .A(n713), .B(n714), .Z(n715) );
  NAND U1067 ( .A(n715), .B(n1146), .Z(n1217) );
  ANDN U1068 ( .B(n[0]), .A(n995), .Z(n989) );
  NAND U1069 ( .A(n1266), .B(n[1]), .Z(n716) );
  XOR U1070 ( .A(n1266), .B(n[1]), .Z(n717) );
  NAND U1071 ( .A(n717), .B(n1269), .Z(n718) );
  NAND U1072 ( .A(n716), .B(n718), .Z(n1265) );
  XOR U1073 ( .A(n[2]), .B(n1247), .Z(n719) );
  NANDN U1074 ( .A(n1244), .B(n719), .Z(n720) );
  NAND U1075 ( .A(n[2]), .B(n1247), .Z(n721) );
  AND U1076 ( .A(n720), .B(n721), .Z(n1239) );
  XOR U1077 ( .A(n[1]), .B(n1676), .Z(n722) );
  ANDN U1078 ( .B(n722), .A(n1707), .Z(n723) );
  XNOR U1079 ( .A(n1677), .B(n723), .Z(n1686) );
  XOR U1080 ( .A(n[1]), .B(n1494), .Z(n724) );
  NANDN U1081 ( .A(n1497), .B(n724), .Z(n725) );
  NAND U1082 ( .A(n[1]), .B(n1494), .Z(n726) );
  AND U1083 ( .A(n725), .B(n726), .Z(n1489) );
  NAND U1084 ( .A(n1483), .B(n[3]), .Z(n727) );
  XOR U1085 ( .A(n1483), .B(n[3]), .Z(n728) );
  NANDN U1086 ( .A(n1479), .B(n728), .Z(n729) );
  NAND U1087 ( .A(n727), .B(n729), .Z(n730) );
  XNOR U1088 ( .A(n730), .B(n1466), .Z(n731) );
  XNOR U1089 ( .A(n1465), .B(n731), .Z(n732) );
  NANDN U1090 ( .A(n1481), .B(n730), .Z(n733) );
  NAND U1091 ( .A(n732), .B(n733), .Z(n1530) );
  ANDN U1092 ( .B(\cin[1][1] ), .A(n1720), .Z(n1699) );
  NAND U1093 ( .A(n1093), .B(n[2]), .Z(n734) );
  XOR U1094 ( .A(n1093), .B(n[2]), .Z(n735) );
  NANDN U1095 ( .A(n1090), .B(n735), .Z(n736) );
  NAND U1096 ( .A(n734), .B(n736), .Z(n1043) );
  XOR U1097 ( .A(n1713), .B(n1714), .Z(n1757) );
  NAND U1098 ( .A(n2044), .B(n2016), .Z(n737) );
  XOR U1099 ( .A(n2044), .B(n2016), .Z(n738) );
  NANDN U1100 ( .A(n[1]), .B(n738), .Z(n739) );
  NAND U1101 ( .A(n737), .B(n739), .Z(n740) );
  OR U1102 ( .A(n740), .B(n2001), .Z(n741) );
  NANDN U1103 ( .A(n2000), .B(n741), .Z(n742) );
  NAND U1104 ( .A(n2025), .B(n742), .Z(n2014) );
  AND U1105 ( .A(n1033), .B(n[0]), .Z(n743) );
  XNOR U1106 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n743), .Z(n1041) );
  NAND U1107 ( .A(n[1]), .B(n1767), .Z(n744) );
  XOR U1108 ( .A(n[1]), .B(n1767), .Z(n745) );
  NANDN U1109 ( .A(n1770), .B(n745), .Z(n746) );
  NAND U1110 ( .A(n744), .B(n746), .Z(n1763) );
  NAND U1111 ( .A(n[1]), .B(n2279), .Z(n747) );
  XOR U1112 ( .A(n[1]), .B(n2279), .Z(n748) );
  NANDN U1113 ( .A(n2282), .B(n748), .Z(n749) );
  NAND U1114 ( .A(n747), .B(n749), .Z(n2286) );
  NAND U1115 ( .A(n1358), .B(n[2]), .Z(n750) );
  XOR U1116 ( .A(n1358), .B(n[2]), .Z(n751) );
  NAND U1117 ( .A(n751), .B(n1351), .Z(n752) );
  NAND U1118 ( .A(n750), .B(n752), .Z(n753) );
  OR U1119 ( .A(n753), .B(n1366), .Z(n754) );
  AND U1120 ( .A(n1364), .B(n754), .Z(n755) );
  XOR U1121 ( .A(n753), .B(n1366), .Z(n756) );
  NANDN U1122 ( .A(n[3]), .B(n756), .Z(n757) );
  NAND U1123 ( .A(n755), .B(n757), .Z(n1367) );
  XOR U1124 ( .A(n1610), .B(n1609), .Z(n1616) );
  NAND U1125 ( .A(n[1]), .B(n1870), .Z(n758) );
  XOR U1126 ( .A(n[1]), .B(n1870), .Z(n759) );
  NANDN U1127 ( .A(n1873), .B(n759), .Z(n760) );
  NAND U1128 ( .A(n758), .B(n760), .Z(n1856) );
  NANDN U1129 ( .A(n2071), .B(n2072), .Z(n761) );
  ANDN U1130 ( .B(n761), .A(n2153), .Z(n2129) );
  XOR U1131 ( .A(n[2]), .B(n1648), .Z(n762) );
  NANDN U1132 ( .A(n1645), .B(n762), .Z(n763) );
  NAND U1133 ( .A(n[2]), .B(n1648), .Z(n764) );
  AND U1134 ( .A(n763), .B(n764), .Z(n1641) );
  ANDN U1135 ( .B(n2198), .A(n2106), .Z(n2116) );
  NAND U1136 ( .A(n2103), .B(n[1]), .Z(n765) );
  XOR U1137 ( .A(n2103), .B(n[1]), .Z(n766) );
  NAND U1138 ( .A(n766), .B(n2104), .Z(n767) );
  NAND U1139 ( .A(n765), .B(n767), .Z(n2111) );
  NAND U1140 ( .A(n2375), .B(n[2]), .Z(n768) );
  XOR U1141 ( .A(n2375), .B(n[2]), .Z(n769) );
  NAND U1142 ( .A(n769), .B(n2378), .Z(n770) );
  NAND U1143 ( .A(n768), .B(n770), .Z(n2395) );
  XOR U1144 ( .A(n[1]), .B(n1779), .Z(n771) );
  NAND U1145 ( .A(n771), .B(n1783), .Z(n772) );
  NAND U1146 ( .A(n[1]), .B(n1779), .Z(n773) );
  AND U1147 ( .A(n772), .B(n773), .Z(n1662) );
  XOR U1148 ( .A(n1881), .B(n1880), .Z(n1906) );
  XOR U1149 ( .A(n[1]), .B(n2192), .Z(n774) );
  NAND U1150 ( .A(n774), .B(n2195), .Z(n775) );
  NAND U1151 ( .A(n[1]), .B(n2192), .Z(n776) );
  AND U1152 ( .A(n775), .B(n776), .Z(n2186) );
  XOR U1153 ( .A(n2355), .B(n2354), .Z(n777) );
  NANDN U1154 ( .A(n[3]), .B(n777), .Z(n778) );
  NAND U1155 ( .A(n2355), .B(n2354), .Z(n779) );
  AND U1156 ( .A(n778), .B(n779), .Z(n780) );
  XOR U1157 ( .A(n2356), .B(n2357), .Z(n781) );
  XNOR U1158 ( .A(n780), .B(n781), .Z(n782) );
  NANDN U1159 ( .A(n2358), .B(n782), .Z(n2403) );
  NANDN U1160 ( .A(n2449), .B(n[1]), .Z(n2423) );
  AND U1161 ( .A(n1931), .B(n[0]), .Z(n783) );
  XNOR U1162 ( .A(n1910), .B(n783), .Z(n1946) );
  XOR U1163 ( .A(n2212), .B(n2211), .Z(n2218) );
  XOR U1164 ( .A(n[2]), .B(n2256), .Z(n784) );
  NANDN U1165 ( .A(n2253), .B(n784), .Z(n785) );
  NAND U1166 ( .A(n[2]), .B(n2256), .Z(n786) );
  AND U1167 ( .A(n785), .B(n786), .Z(n2260) );
  NANDN U1168 ( .A(n2517), .B(n[1]), .Z(n2500) );
  XOR U1169 ( .A(\cin[1][3] ), .B(n2493), .Z(n787) );
  NAND U1170 ( .A(n2494), .B(n787), .Z(n788) );
  XNOR U1171 ( .A(n2495), .B(n788), .Z(n2513) );
  XOR U1172 ( .A(n[2]), .B(n2537), .Z(n789) );
  NANDN U1173 ( .A(n2541), .B(n789), .Z(n790) );
  NAND U1174 ( .A(n[2]), .B(n2537), .Z(n791) );
  AND U1175 ( .A(n790), .B(n791), .Z(n2545) );
  IV U1176 ( .A(n[1]), .Z(n792) );
  IV U1177 ( .A(n[2]), .Z(n793) );
  IV U1178 ( .A(n[3]), .Z(n794) );
  OR U1179 ( .A(e[2]), .B(e[3]), .Z(n1949) );
  AND U1180 ( .A(e[1]), .B(n1949), .Z(n1992) );
  NANDN U1181 ( .A(e[2]), .B(e[3]), .Z(n1356) );
  NAND U1182 ( .A(\cin[1][2] ), .B(\cin[1][3] ), .Z(n840) );
  AND U1183 ( .A(\cin[1][3] ), .B(n794), .Z(n1068) );
  OR U1184 ( .A(\cin[1][1] ), .B(n792), .Z(n795) );
  ANDN U1185 ( .B(n[2]), .A(\cin[1][2] ), .Z(n1067) );
  ANDN U1186 ( .B(n795), .A(n1067), .Z(n798) );
  ANDN U1187 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n[0]), .Z(n2488) );
  XOR U1188 ( .A(n792), .B(\cin[1][1] ), .Z(n796) );
  NANDN U1189 ( .A(n2488), .B(n796), .Z(n797) );
  NAND U1190 ( .A(n798), .B(n797), .Z(n1052) );
  NANDN U1191 ( .A(n[2]), .B(\cin[1][2] ), .Z(n2271) );
  NAND U1192 ( .A(n1052), .B(n2271), .Z(n799) );
  NAND U1193 ( .A(\cin[1][3] ), .B(n799), .Z(n800) );
  NANDN U1194 ( .A(n1068), .B(n800), .Z(n816) );
  NAND U1195 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[1][3] ), .Z(n801) );
  NAND U1196 ( .A(n[0]), .B(n801), .Z(n807) );
  AND U1197 ( .A(\cin[1][1] ), .B(\cin[1][3] ), .Z(n810) );
  XOR U1198 ( .A(n[2]), .B(n814), .Z(n802) );
  NAND U1199 ( .A(n816), .B(n802), .Z(n803) );
  XOR U1200 ( .A(n840), .B(n803), .Z(n823) );
  IV U1201 ( .A(n816), .Z(n815) );
  NANDN U1202 ( .A(n815), .B(n[0]), .Z(n804) );
  XNOR U1203 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n804), .Z(n806) );
  NANDN U1204 ( .A(\cin[1][3] ), .B(n815), .Z(n805) );
  NAND U1205 ( .A(n806), .B(n805), .Z(n830) );
  NAND U1206 ( .A(n[0]), .B(n830), .Z(n824) );
  NANDN U1207 ( .A(n[1]), .B(n824), .Z(n813) );
  NOR U1208 ( .A(n792), .B(n824), .Z(n811) );
  XOR U1209 ( .A(n792), .B(n807), .Z(n808) );
  NAND U1210 ( .A(n816), .B(n808), .Z(n809) );
  XNOR U1211 ( .A(n810), .B(n809), .Z(n827) );
  NANDN U1212 ( .A(n811), .B(n827), .Z(n812) );
  AND U1213 ( .A(n813), .B(n812), .Z(n820) );
  NANDN U1214 ( .A(n[3]), .B(n831), .Z(n819) );
  OR U1215 ( .A(n831), .B(n816), .Z(n817) );
  NAND U1216 ( .A(n835), .B(n817), .Z(n818) );
  AND U1217 ( .A(n819), .B(n818), .Z(n828) );
  XOR U1218 ( .A(n[2]), .B(n820), .Z(n821) );
  NANDN U1219 ( .A(n828), .B(n821), .Z(n822) );
  XNOR U1220 ( .A(n823), .B(n822), .Z(n839) );
  XOR U1221 ( .A(n792), .B(n824), .Z(n825) );
  NANDN U1222 ( .A(n828), .B(n825), .Z(n826) );
  XNOR U1223 ( .A(n827), .B(n826), .Z(n845) );
  ANDN U1224 ( .B(n[0]), .A(n828), .Z(n829) );
  XNOR U1225 ( .A(n830), .B(n829), .Z(n846) );
  NAND U1226 ( .A(\cin[1][1] ), .B(n846), .Z(n843) );
  NANDN U1227 ( .A(n845), .B(n843), .Z(n836) );
  XNOR U1228 ( .A(n[3]), .B(n831), .Z(n833) );
  OR U1229 ( .A(n831), .B(\cin[1][3] ), .Z(n832) );
  NAND U1230 ( .A(n833), .B(n832), .Z(n834) );
  AND U1231 ( .A(n835), .B(n834), .Z(n862) );
  ANDN U1232 ( .B(\cin[1][3] ), .A(n839), .Z(n837) );
  AND U1233 ( .A(n837), .B(n836), .Z(n838) );
  NAND U1234 ( .A(\cin[1][2] ), .B(n838), .Z(n842) );
  NANDN U1235 ( .A(n840), .B(n839), .Z(n841) );
  AND U1236 ( .A(n842), .B(n841), .Z(n863) );
  NAND U1237 ( .A(n843), .B(\cin[1][2] ), .Z(n844) );
  XOR U1238 ( .A(n845), .B(n844), .Z(n869) );
  NAND U1239 ( .A(n[2]), .B(n869), .Z(n852) );
  NOR U1240 ( .A(n[2]), .B(n869), .Z(n850) );
  AND U1241 ( .A(\cin[1][2] ), .B(\cin[1][1] ), .Z(n892) );
  XOR U1242 ( .A(n846), .B(n892), .Z(n876) );
  OR U1243 ( .A(n876), .B(n792), .Z(n849) );
  NAND U1244 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[1][2] ), .Z(n871) );
  AND U1245 ( .A(n[0]), .B(n871), .Z(n872) );
  XNOR U1246 ( .A(n[1]), .B(n876), .Z(n847) );
  NAND U1247 ( .A(n872), .B(n847), .Z(n848) );
  AND U1248 ( .A(n849), .B(n848), .Z(n866) );
  OR U1249 ( .A(n850), .B(n866), .Z(n851) );
  AND U1250 ( .A(n852), .B(n851), .Z(n854) );
  NANDN U1251 ( .A(n[3]), .B(n854), .Z(n853) );
  AND U1252 ( .A(n874), .B(n853), .Z(n859) );
  ANDN U1253 ( .B(n[3]), .A(n854), .Z(n856) );
  ANDN U1254 ( .B(n859), .A(n856), .Z(n855) );
  XNOR U1255 ( .A(n857), .B(n855), .Z(n909) );
  NANDN U1256 ( .A(n[3]), .B(n909), .Z(n865) );
  XNOR U1257 ( .A(n862), .B(n863), .Z(n861) );
  OR U1258 ( .A(n857), .B(n856), .Z(n858) );
  NAND U1259 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U1260 ( .A(n861), .B(n860), .Z(n934) );
  NANDN U1261 ( .A(n863), .B(n862), .Z(n864) );
  NANDN U1262 ( .A(n934), .B(n864), .Z(n906) );
  ANDN U1263 ( .B(n865), .A(n906), .Z(n885) );
  XNOR U1264 ( .A(n[2]), .B(n866), .Z(n867) );
  NAND U1265 ( .A(n874), .B(n867), .Z(n868) );
  XNOR U1266 ( .A(n869), .B(n868), .Z(n886) );
  AND U1267 ( .A(n886), .B(n[2]), .Z(n883) );
  NANDN U1268 ( .A(n885), .B(n883), .Z(n888) );
  NAND U1269 ( .A(n874), .B(n[0]), .Z(n870) );
  XNOR U1270 ( .A(n871), .B(n870), .Z(n891) );
  NAND U1271 ( .A(n[0]), .B(n891), .Z(n893) );
  NANDN U1272 ( .A(n[1]), .B(n893), .Z(n879) );
  NOR U1273 ( .A(n792), .B(n893), .Z(n877) );
  XOR U1274 ( .A(n[1]), .B(n872), .Z(n873) );
  NAND U1275 ( .A(n874), .B(n873), .Z(n875) );
  XNOR U1276 ( .A(n876), .B(n875), .Z(n897) );
  NANDN U1277 ( .A(n877), .B(n897), .Z(n878) );
  AND U1278 ( .A(n879), .B(n878), .Z(n889) );
  OR U1279 ( .A(n886), .B(n[2]), .Z(n880) );
  NAND U1280 ( .A(n889), .B(n880), .Z(n881) );
  ANDN U1281 ( .B(n881), .A(n907), .Z(n882) );
  NANDN U1282 ( .A(n883), .B(n882), .Z(n884) );
  NAND U1283 ( .A(n885), .B(n884), .Z(n895) );
  IV U1284 ( .A(n895), .Z(n908) );
  NANDN U1285 ( .A(n908), .B(n[2]), .Z(n887) );
  ANDN U1286 ( .B(n887), .A(n886), .Z(n905) );
  ANDN U1287 ( .B(n888), .A(n905), .Z(n903) );
  NAND U1288 ( .A(n895), .B(n889), .Z(n902) );
  XNOR U1289 ( .A(n903), .B(n902), .Z(n915) );
  NAND U1290 ( .A(n895), .B(n[0]), .Z(n890) );
  XNOR U1291 ( .A(n891), .B(n890), .Z(n916) );
  IV U1292 ( .A(n916), .Z(n920) );
  AND U1293 ( .A(n892), .B(n920), .Z(n901) );
  XOR U1294 ( .A(n792), .B(n893), .Z(n894) );
  NAND U1295 ( .A(n895), .B(n894), .Z(n896) );
  XNOR U1296 ( .A(n897), .B(n896), .Z(n919) );
  AND U1297 ( .A(\cin[1][1] ), .B(n920), .Z(n898) );
  OR U1298 ( .A(\cin[1][2] ), .B(n898), .Z(n899) );
  NAND U1299 ( .A(n919), .B(n899), .Z(n900) );
  NANDN U1300 ( .A(n901), .B(n900), .Z(n912) );
  NAND U1301 ( .A(n903), .B(n902), .Z(n904) );
  NANDN U1302 ( .A(n905), .B(n904), .Z(n927) );
  NAND U1303 ( .A(n907), .B(n906), .Z(n911) );
  NANDN U1304 ( .A(n908), .B(n[3]), .Z(n910) );
  AND U1305 ( .A(n910), .B(n909), .Z(n930) );
  ANDN U1306 ( .B(n911), .A(n930), .Z(n928) );
  XOR U1307 ( .A(n927), .B(n928), .Z(n931) );
  XOR U1308 ( .A(n932), .B(n931), .Z(n948) );
  XOR U1309 ( .A(n912), .B(\cin[1][3] ), .Z(n913) );
  NAND U1310 ( .A(\cin[1][1] ), .B(n913), .Z(n914) );
  XNOR U1311 ( .A(n915), .B(n914), .Z(n955) );
  NAND U1312 ( .A(n[3]), .B(n955), .Z(n943) );
  NOR U1313 ( .A(n[3]), .B(n955), .Z(n945) );
  XNOR U1314 ( .A(\cin[1][2] ), .B(n916), .Z(n917) );
  NAND U1315 ( .A(\cin[1][1] ), .B(n917), .Z(n918) );
  XNOR U1316 ( .A(n919), .B(n918), .Z(n961) );
  ANDN U1317 ( .B(n[2]), .A(n961), .Z(n941) );
  XOR U1318 ( .A(\cin[1][1] ), .B(n920), .Z(n969) );
  NANDN U1319 ( .A(n969), .B(n[1]), .Z(n923) );
  NAND U1320 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(\cin[1][1] ), .Z(n964) );
  AND U1321 ( .A(n[0]), .B(n964), .Z(n965) );
  XNOR U1322 ( .A(n[1]), .B(n969), .Z(n921) );
  NAND U1323 ( .A(n965), .B(n921), .Z(n922) );
  AND U1324 ( .A(n923), .B(n922), .Z(n958) );
  NANDN U1325 ( .A(n941), .B(n958), .Z(n924) );
  AND U1326 ( .A(n961), .B(n793), .Z(n938) );
  ANDN U1327 ( .B(n924), .A(n938), .Z(n952) );
  NANDN U1328 ( .A(n945), .B(n952), .Z(n925) );
  AND U1329 ( .A(n943), .B(n925), .Z(n926) );
  XNOR U1330 ( .A(n948), .B(n926), .Z(n950) );
  AND U1331 ( .A(n928), .B(n927), .Z(n929) );
  NOR U1332 ( .A(n930), .B(n929), .Z(n936) );
  AND U1333 ( .A(n932), .B(n931), .Z(n933) );
  XNOR U1334 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U1335 ( .A(n936), .B(n935), .Z(n951) );
  ANDN U1336 ( .B(n969), .A(n[1]), .Z(n940) );
  IV U1337 ( .A(n964), .Z(n1009) );
  ANDN U1338 ( .B(n1009), .A(n[0]), .Z(n937) );
  NOR U1339 ( .A(n938), .B(n937), .Z(n939) );
  NANDN U1340 ( .A(n940), .B(n939), .Z(n942) );
  ANDN U1341 ( .B(n942), .A(n941), .Z(n944) );
  NAND U1342 ( .A(n944), .B(n943), .Z(n946) );
  ANDN U1343 ( .B(n946), .A(n945), .Z(n947) );
  NANDN U1344 ( .A(n951), .B(n947), .Z(n949) );
  NOR U1345 ( .A(n949), .B(n948), .Z(n967) );
  ANDN U1346 ( .B(n950), .A(n967), .Z(n1001) );
  NOR U1347 ( .A(n1001), .B(n951), .Z(n957) );
  XOR U1348 ( .A(n[3]), .B(n952), .Z(n953) );
  NANDN U1349 ( .A(n967), .B(n953), .Z(n954) );
  XNOR U1350 ( .A(n955), .B(n954), .Z(n974) );
  AND U1351 ( .A(n974), .B(n[3]), .Z(n962) );
  NANDN U1352 ( .A(n957), .B(n962), .Z(n976) );
  OR U1353 ( .A(n974), .B(n[3]), .Z(n956) );
  AND U1354 ( .A(n957), .B(n956), .Z(n981) );
  XNOR U1355 ( .A(n[2]), .B(n958), .Z(n959) );
  NANDN U1356 ( .A(n967), .B(n959), .Z(n960) );
  XNOR U1357 ( .A(n961), .B(n960), .Z(n979) );
  ANDN U1358 ( .B(n[2]), .A(n979), .Z(n980) );
  NOR U1359 ( .A(n980), .B(n962), .Z(n972) );
  NANDN U1360 ( .A(n967), .B(n[0]), .Z(n963) );
  XOR U1361 ( .A(n964), .B(n963), .Z(n995) );
  XOR U1362 ( .A(n965), .B(n[1]), .Z(n966) );
  NANDN U1363 ( .A(n967), .B(n966), .Z(n968) );
  XOR U1364 ( .A(n969), .B(n968), .Z(n992) );
  NANDN U1365 ( .A(n[2]), .B(n979), .Z(n970) );
  NANDN U1366 ( .A(n983), .B(n970), .Z(n971) );
  NAND U1367 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1368 ( .A(n981), .B(n973), .Z(n993) );
  IV U1369 ( .A(n993), .Z(n977) );
  NANDN U1370 ( .A(n977), .B(n[3]), .Z(n975) );
  ANDN U1371 ( .B(n975), .A(n974), .Z(n986) );
  ANDN U1372 ( .B(n976), .A(n986), .Z(n1000) );
  NANDN U1373 ( .A(n977), .B(n[2]), .Z(n978) );
  AND U1374 ( .A(n979), .B(n978), .Z(n985) );
  NANDN U1375 ( .A(n981), .B(n980), .Z(n982) );
  ANDN U1376 ( .B(n982), .A(n985), .Z(n988) );
  NANDN U1377 ( .A(n983), .B(n993), .Z(n987) );
  NAND U1378 ( .A(n988), .B(n987), .Z(n984) );
  NANDN U1379 ( .A(n985), .B(n984), .Z(n999) );
  XNOR U1380 ( .A(n988), .B(n987), .Z(n1007) );
  XOR U1381 ( .A(n[1]), .B(n989), .Z(n990) );
  NAND U1382 ( .A(n993), .B(n990), .Z(n991) );
  XNOR U1383 ( .A(n992), .B(n991), .Z(n1013) );
  NANDN U1384 ( .A(n1013), .B(\cin[1][2] ), .Z(n998) );
  XNOR U1385 ( .A(\cin[1][2] ), .B(n1013), .Z(n996) );
  NAND U1386 ( .A(n993), .B(n[0]), .Z(n994) );
  XNOR U1387 ( .A(n995), .B(n994), .Z(n1008) );
  AND U1388 ( .A(\cin[1][1] ), .B(n1008), .Z(n1010) );
  NAND U1389 ( .A(n996), .B(n1010), .Z(n997) );
  NAND U1390 ( .A(n998), .B(n997), .Z(n1004) );
  XNOR U1391 ( .A(n1000), .B(n999), .Z(n1002) );
  XOR U1392 ( .A(n1003), .B(n1002), .Z(n1021) );
  XOR U1393 ( .A(n1004), .B(\cin[1][3] ), .Z(n1005) );
  NAND U1394 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1005), .Z(n1006) );
  XNOR U1395 ( .A(n1007), .B(n1006), .Z(n1035) );
  NOR U1396 ( .A(n[3]), .B(n1035), .Z(n1017) );
  XOR U1397 ( .A(n1009), .B(n1008), .Z(n1026) );
  XOR U1398 ( .A(\cin[1][2] ), .B(n1010), .Z(n1011) );
  NAND U1399 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1011), .Z(n1012) );
  XNOR U1400 ( .A(n1013), .B(n1012), .Z(n1030) );
  AND U1401 ( .A(n1030), .B(n[2]), .Z(n1014) );
  ANDN U1402 ( .B(n793), .A(n1030), .Z(n1015) );
  AND U1403 ( .A(n1035), .B(n[3]), .Z(n1018) );
  NANDN U1404 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n[0]), .Z(n2276) );
  NANDN U1405 ( .A(n1014), .B(n1027), .Z(n1016) );
  ANDN U1406 ( .B(n1016), .A(n1015), .Z(n1031) );
  NANDN U1407 ( .A(n1017), .B(n1031), .Z(n1019) );
  ANDN U1408 ( .B(n1019), .A(n1018), .Z(n1020) );
  NANDN U1409 ( .A(n1021), .B(n1020), .Z(n1023) );
  ANDN U1410 ( .B(n1023), .A(n1022), .Z(n1045) );
  XOR U1411 ( .A(n2276), .B(n792), .Z(n1024) );
  NAND U1412 ( .A(n1033), .B(n1024), .Z(n1025) );
  XNOR U1413 ( .A(n1026), .B(n1025), .Z(n1184) );
  AND U1414 ( .A(n[0]), .B(n1041), .Z(n1180) );
  XNOR U1415 ( .A(n[2]), .B(n1027), .Z(n1028) );
  NAND U1416 ( .A(n1033), .B(n1028), .Z(n1029) );
  XNOR U1417 ( .A(n1030), .B(n1029), .Z(n1093) );
  NAND U1418 ( .A(n[3]), .B(n1043), .Z(n1038) );
  ANDN U1419 ( .B(n794), .A(n1043), .Z(n1036) );
  XOR U1420 ( .A(n[3]), .B(n1031), .Z(n1032) );
  NAND U1421 ( .A(n1033), .B(n1032), .Z(n1034) );
  XNOR U1422 ( .A(n1035), .B(n1034), .Z(n1046) );
  NANDN U1423 ( .A(n1036), .B(n1046), .Z(n1037) );
  NAND U1424 ( .A(n1038), .B(n1037), .Z(n1039) );
  AND U1425 ( .A(n1045), .B(n1039), .Z(n1181) );
  NANDN U1426 ( .A(n1181), .B(n[0]), .Z(n1040) );
  XOR U1427 ( .A(n1041), .B(n1040), .Z(n1294) );
  NANDN U1428 ( .A(n1356), .B(n1294), .Z(n1042) );
  ANDN U1429 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(e[3]), .Z(n1951) );
  ANDN U1430 ( .B(n1042), .A(n1951), .Z(n1339) );
  AND U1431 ( .A(e[2]), .B(e[3]), .Z(n1374) );
  NAND U1432 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1294), .Z(n1308) );
  XOR U1433 ( .A(n[3]), .B(n1043), .Z(n1044) );
  XNOR U1434 ( .A(n1046), .B(n1044), .Z(n1048) );
  NAND U1435 ( .A(n1046), .B(n1045), .Z(n1047) );
  NAND U1436 ( .A(n1048), .B(n1047), .Z(n1355) );
  NANDN U1437 ( .A(n1355), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1058)
         );
  NAND U1438 ( .A(n[0]), .B(n1058), .Z(n1062) );
  NANDN U1439 ( .A(n[1]), .B(n1062), .Z(n1051) );
  NOR U1440 ( .A(n792), .B(n1062), .Z(n1049) );
  NANDN U1441 ( .A(n1355), .B(\cin[1][1] ), .Z(n1066) );
  OR U1442 ( .A(n1049), .B(n1066), .Z(n1050) );
  AND U1443 ( .A(n1051), .B(n1050), .Z(n1069) );
  XNOR U1444 ( .A(n[2]), .B(n1069), .Z(n1055) );
  NANDN U1445 ( .A(\cin[1][3] ), .B(n[3]), .Z(n1054) );
  ANDN U1446 ( .B(n2271), .A(n1068), .Z(n1053) );
  AND U1447 ( .A(n1053), .B(n1052), .Z(n1072) );
  ANDN U1448 ( .B(n1054), .A(n1072), .Z(n2275) );
  NANDN U1449 ( .A(n1055), .B(n2275), .Z(n1056) );
  XNOR U1450 ( .A(\cin[1][2] ), .B(n1056), .Z(n1057) );
  ANDN U1451 ( .B(n1057), .A(n1355), .Z(n1079) );
  ANDN U1452 ( .B(n2275), .A(n1355), .Z(n1064) );
  AND U1453 ( .A(n[0]), .B(n1064), .Z(n1059) );
  NAND U1454 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1059), .Z(n1061) );
  NANDN U1455 ( .A(n1059), .B(n1058), .Z(n1060) );
  AND U1456 ( .A(n1061), .B(n1060), .Z(n1086) );
  ANDN U1457 ( .B(n[0]), .A(n1086), .Z(n1080) );
  XOR U1458 ( .A(n792), .B(n1062), .Z(n1063) );
  NAND U1459 ( .A(n1064), .B(n1063), .Z(n1065) );
  XOR U1460 ( .A(n1066), .B(n1065), .Z(n1083) );
  ANDN U1461 ( .B(n1068), .A(n1067), .Z(n2274) );
  NAND U1462 ( .A(n1069), .B(n2271), .Z(n1070) );
  ANDN U1463 ( .B(n1070), .A(n1355), .Z(n1071) );
  NAND U1464 ( .A(n2274), .B(n1071), .Z(n1094) );
  NAND U1465 ( .A(n1095), .B(n1094), .Z(n1075) );
  AND U1466 ( .A(\cin[1][3] ), .B(n1072), .Z(n2288) );
  NANDN U1467 ( .A(n1355), .B(n2288), .Z(n1073) );
  AND U1468 ( .A(n1094), .B(n1073), .Z(n1098) );
  NAND U1469 ( .A(n[3]), .B(n1098), .Z(n1074) );
  AND U1470 ( .A(n1075), .B(n1074), .Z(n1084) );
  XOR U1471 ( .A(n[2]), .B(n1076), .Z(n1077) );
  NAND U1472 ( .A(n1084), .B(n1077), .Z(n1078) );
  XNOR U1473 ( .A(n1079), .B(n1078), .Z(n1103) );
  XOR U1474 ( .A(n[1]), .B(n1080), .Z(n1081) );
  NAND U1475 ( .A(n1084), .B(n1081), .Z(n1082) );
  XNOR U1476 ( .A(n1083), .B(n1082), .Z(n1111) );
  NAND U1477 ( .A(\cin[1][2] ), .B(n1111), .Z(n1089) );
  XOR U1478 ( .A(\cin[1][2] ), .B(n1111), .Z(n1087) );
  NAND U1479 ( .A(n1084), .B(n[0]), .Z(n1085) );
  XNOR U1480 ( .A(n1086), .B(n1085), .Z(n1105) );
  AND U1481 ( .A(\cin[1][1] ), .B(n1105), .Z(n1108) );
  NAND U1482 ( .A(n1087), .B(n1108), .Z(n1088) );
  AND U1483 ( .A(n1089), .B(n1088), .Z(n1100) );
  XNOR U1484 ( .A(n[2]), .B(n1090), .Z(n1091) );
  NANDN U1485 ( .A(n1181), .B(n1091), .Z(n1092) );
  XNOR U1486 ( .A(n1093), .B(n1092), .Z(n1349) );
  NANDN U1487 ( .A(n1094), .B(n1095), .Z(n1097) );
  NANDN U1488 ( .A(n1095), .B(n[3]), .Z(n1096) );
  AND U1489 ( .A(n1097), .B(n1096), .Z(n1099) );
  ANDN U1490 ( .B(n1099), .A(n1098), .Z(n1128) );
  NAND U1491 ( .A(n1129), .B(n1128), .Z(n1130) );
  OR U1492 ( .A(n1129), .B(n1128), .Z(n1119) );
  XNOR U1493 ( .A(\cin[1][3] ), .B(n1100), .Z(n1101) );
  ANDN U1494 ( .B(n1101), .A(n1349), .Z(n1102) );
  XNOR U1495 ( .A(n1103), .B(n1102), .Z(n1134) );
  AND U1496 ( .A(n1134), .B(n[3]), .Z(n1126) );
  NANDN U1497 ( .A(n1349), .B(\cin[1][1] ), .Z(n1104) );
  XNOR U1498 ( .A(n1105), .B(n1104), .Z(n1144) );
  ANDN U1499 ( .B(n1144), .A(n[1]), .Z(n1106) );
  ANDN U1500 ( .B(n2488), .A(n1349), .Z(n1158) );
  OR U1501 ( .A(n1106), .B(n1158), .Z(n1107) );
  AND U1502 ( .A(n1122), .B(n1107), .Z(n1112) );
  XOR U1503 ( .A(\cin[1][2] ), .B(n1108), .Z(n1109) );
  NANDN U1504 ( .A(n1349), .B(n1109), .Z(n1110) );
  XNOR U1505 ( .A(n1111), .B(n1110), .Z(n1139) );
  NAND U1506 ( .A(n1112), .B(n1139), .Z(n1115) );
  XOR U1507 ( .A(n1112), .B(n1139), .Z(n1113) );
  NAND U1508 ( .A(n793), .B(n1113), .Z(n1114) );
  NAND U1509 ( .A(n1115), .B(n1114), .Z(n1116) );
  NANDN U1510 ( .A(n1126), .B(n1116), .Z(n1117) );
  NOR U1511 ( .A(n[3]), .B(n1134), .Z(n1127) );
  ANDN U1512 ( .B(n1117), .A(n1127), .Z(n1118) );
  NANDN U1513 ( .A(n1119), .B(n1118), .Z(n1146) );
  XNOR U1514 ( .A(n[1]), .B(n1144), .Z(n1120) );
  NANDN U1515 ( .A(n1349), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1145)
         );
  AND U1516 ( .A(n[0]), .B(n1145), .Z(n1141) );
  NAND U1517 ( .A(n1120), .B(n1141), .Z(n1121) );
  AND U1518 ( .A(n1122), .B(n1121), .Z(n1136) );
  NANDN U1519 ( .A(n[2]), .B(n1136), .Z(n1125) );
  NOR U1520 ( .A(n793), .B(n1136), .Z(n1123) );
  NANDN U1521 ( .A(n1123), .B(n1139), .Z(n1124) );
  AND U1522 ( .A(n1125), .B(n1124), .Z(n1131) );
  AND U1523 ( .A(n1130), .B(n1217), .Z(n1187) );
  XOR U1524 ( .A(n[3]), .B(n1131), .Z(n1132) );
  NAND U1525 ( .A(n1146), .B(n1132), .Z(n1133) );
  XNOR U1526 ( .A(n1134), .B(n1133), .Z(n1189) );
  OR U1527 ( .A(n1189), .B(n[3]), .Z(n1135) );
  AND U1528 ( .A(n1187), .B(n1135), .Z(n1165) );
  XOR U1529 ( .A(n793), .B(n1136), .Z(n1137) );
  AND U1530 ( .A(n1137), .B(n1146), .Z(n1138) );
  XNOR U1531 ( .A(n1139), .B(n1138), .Z(n1166) );
  NAND U1532 ( .A(n[2]), .B(n1166), .Z(n1140) );
  AND U1533 ( .A(n1189), .B(n[3]), .Z(n1186) );
  ANDN U1534 ( .B(n1140), .A(n1186), .Z(n1156) );
  XOR U1535 ( .A(n[2]), .B(n1166), .Z(n1154) );
  XOR U1536 ( .A(n1141), .B(n[1]), .Z(n1142) );
  NAND U1537 ( .A(n1146), .B(n1142), .Z(n1143) );
  XNOR U1538 ( .A(n1144), .B(n1143), .Z(n1161) );
  XOR U1539 ( .A(n1161), .B(n792), .Z(n1150) );
  XNOR U1540 ( .A(n1146), .B(n1145), .Z(n1148) );
  NANDN U1541 ( .A(n[0]), .B(n1146), .Z(n1147) );
  NAND U1542 ( .A(n1148), .B(n1147), .Z(n1159) );
  NAND U1543 ( .A(n[0]), .B(n1159), .Z(n1149) );
  NAND U1544 ( .A(n1150), .B(n1149), .Z(n1152) );
  NAND U1545 ( .A(n792), .B(n1161), .Z(n1151) );
  AND U1546 ( .A(n1152), .B(n1151), .Z(n1153) );
  NAND U1547 ( .A(n1154), .B(n1153), .Z(n1155) );
  NAND U1548 ( .A(n1156), .B(n1155), .Z(n1157) );
  AND U1549 ( .A(n1165), .B(n1157), .Z(n1188) );
  ANDN U1550 ( .B(n[1]), .A(n1188), .Z(n1160) );
  NANDN U1551 ( .A(n1160), .B(n1161), .Z(n1163) );
  ANDN U1552 ( .B(n[0]), .A(n1188), .Z(n1173) );
  ANDN U1553 ( .B(n1159), .A(n1158), .Z(n1172) );
  AND U1554 ( .A(n1173), .B(n1172), .Z(n1171) );
  XNOR U1555 ( .A(n1161), .B(n1160), .Z(n1170) );
  NANDN U1556 ( .A(n1171), .B(n1170), .Z(n1162) );
  NAND U1557 ( .A(n1163), .B(n1162), .Z(n1192) );
  NANDN U1558 ( .A(n793), .B(n1166), .Z(n1164) );
  OR U1559 ( .A(n1165), .B(n1164), .Z(n1168) );
  NANDN U1560 ( .A(n1188), .B(n[2]), .Z(n1167) );
  ANDN U1561 ( .B(n1167), .A(n1166), .Z(n1195) );
  ANDN U1562 ( .B(n1168), .A(n1195), .Z(n1193) );
  XNOR U1563 ( .A(n1192), .B(n1193), .Z(n1169) );
  IV U1564 ( .A(n1169), .Z(n1199) );
  AND U1565 ( .A(\cin[1][3] ), .B(n1199), .Z(n1179) );
  XNOR U1566 ( .A(\cin[1][3] ), .B(n1169), .Z(n1177) );
  XOR U1567 ( .A(n1171), .B(n1170), .Z(n1208) );
  NANDN U1568 ( .A(n1208), .B(\cin[1][2] ), .Z(n1176) );
  XNOR U1569 ( .A(\cin[1][2] ), .B(n1208), .Z(n1174) );
  XOR U1570 ( .A(n1173), .B(n1172), .Z(n1201) );
  ANDN U1571 ( .B(\cin[1][1] ), .A(n1201), .Z(n1205) );
  NAND U1572 ( .A(n1174), .B(n1205), .Z(n1175) );
  AND U1573 ( .A(n1176), .B(n1175), .Z(n1196) );
  ANDN U1574 ( .B(n1177), .A(n1196), .Z(n1178) );
  OR U1575 ( .A(n1179), .B(n1178), .Z(n1185) );
  XOR U1576 ( .A(n[1]), .B(n1180), .Z(n1182) );
  ANDN U1577 ( .B(n1182), .A(n1181), .Z(n1183) );
  XNOR U1578 ( .A(n1184), .B(n1183), .Z(n1340) );
  ANDN U1579 ( .B(n1185), .A(n1340), .Z(n1214) );
  NANDN U1580 ( .A(n1187), .B(n1186), .Z(n1191) );
  NANDN U1581 ( .A(n1188), .B(n[3]), .Z(n1190) );
  ANDN U1582 ( .B(n1190), .A(n1189), .Z(n1213) );
  ANDN U1583 ( .B(n1191), .A(n1213), .Z(n1211) );
  NAND U1584 ( .A(n1193), .B(n1192), .Z(n1194) );
  NANDN U1585 ( .A(n1195), .B(n1194), .Z(n1210) );
  XOR U1586 ( .A(n1211), .B(n1210), .Z(n1215) );
  XOR U1587 ( .A(n1214), .B(n1215), .Z(n1237) );
  XNOR U1588 ( .A(\cin[1][3] ), .B(n1196), .Z(n1197) );
  ANDN U1589 ( .B(n1197), .A(n1340), .Z(n1198) );
  XNOR U1590 ( .A(n1199), .B(n1198), .Z(n1242) );
  AND U1591 ( .A(n1242), .B(n[3]), .Z(n1226) );
  NOR U1592 ( .A(n[3]), .B(n1242), .Z(n1220) );
  NANDN U1593 ( .A(n1340), .B(\cin[1][1] ), .Z(n1200) );
  XNOR U1594 ( .A(n1201), .B(n1200), .Z(n1255) );
  NAND U1595 ( .A(n[1]), .B(n1255), .Z(n1225) );
  NANDN U1596 ( .A(n1340), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1202)
         );
  AND U1597 ( .A(n[0]), .B(n1202), .Z(n1251) );
  IV U1598 ( .A(n1255), .Z(n1221) );
  XNOR U1599 ( .A(n[1]), .B(n1221), .Z(n1203) );
  NAND U1600 ( .A(n1251), .B(n1203), .Z(n1204) );
  AND U1601 ( .A(n1225), .B(n1204), .Z(n1244) );
  XOR U1602 ( .A(\cin[1][2] ), .B(n1205), .Z(n1206) );
  NANDN U1603 ( .A(n1340), .B(n1206), .Z(n1207) );
  XNOR U1604 ( .A(n1208), .B(n1207), .Z(n1247) );
  OR U1605 ( .A(n1220), .B(n1239), .Z(n1209) );
  NANDN U1606 ( .A(n1226), .B(n1209), .Z(n1235) );
  AND U1607 ( .A(n1211), .B(n1210), .Z(n1212) );
  NOR U1608 ( .A(n1213), .B(n1212), .Z(n1219) );
  AND U1609 ( .A(n1215), .B(n1214), .Z(n1216) );
  XOR U1610 ( .A(n1217), .B(n1216), .Z(n1218) );
  XNOR U1611 ( .A(n1219), .B(n1218), .Z(n1238) );
  NOR U1612 ( .A(n1220), .B(n1238), .Z(n1233) );
  NANDN U1613 ( .A(n1340), .B(n2488), .Z(n1223) );
  NANDN U1614 ( .A(n[1]), .B(n1221), .Z(n1222) );
  NAND U1615 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U1616 ( .A(n1225), .B(n1224), .Z(n1228) );
  NAND U1617 ( .A(n[2]), .B(n1228), .Z(n1227) );
  ANDN U1618 ( .B(n1227), .A(n1226), .Z(n1231) );
  XOR U1619 ( .A(n1228), .B(n[2]), .Z(n1229) );
  NAND U1620 ( .A(n1229), .B(n1247), .Z(n1230) );
  AND U1621 ( .A(n1231), .B(n1230), .Z(n1232) );
  ANDN U1622 ( .B(n1233), .A(n1232), .Z(n1234) );
  ANDN U1623 ( .B(n1234), .A(n1237), .Z(n1248) );
  IV U1624 ( .A(n1248), .Z(n1253) );
  AND U1625 ( .A(n1235), .B(n1253), .Z(n1236) );
  XNOR U1626 ( .A(n1237), .B(n1236), .Z(n1304) );
  ANDN U1627 ( .B(n1304), .A(n1238), .Z(n1277) );
  XNOR U1628 ( .A(n[3]), .B(n1239), .Z(n1240) );
  NAND U1629 ( .A(n1253), .B(n1240), .Z(n1241) );
  XNOR U1630 ( .A(n1242), .B(n1241), .Z(n1279) );
  OR U1631 ( .A(n1279), .B(n[3]), .Z(n1243) );
  AND U1632 ( .A(n1277), .B(n1243), .Z(n1261) );
  XNOR U1633 ( .A(n[2]), .B(n1244), .Z(n1245) );
  NAND U1634 ( .A(n1253), .B(n1245), .Z(n1246) );
  XNOR U1635 ( .A(n1247), .B(n1246), .Z(n1262) );
  AND U1636 ( .A(n1262), .B(n[2]), .Z(n1257) );
  NANDN U1637 ( .A(n1261), .B(n1257), .Z(n1264) );
  AND U1638 ( .A(n1279), .B(n[3]), .Z(n1276) );
  ANDN U1639 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n1340), .Z(n1250) );
  ANDN U1640 ( .B(n[0]), .A(n1248), .Z(n1249) );
  XOR U1641 ( .A(n1250), .B(n1249), .Z(n1272) );
  ANDN U1642 ( .B(n[0]), .A(n1272), .Z(n1266) );
  XOR U1643 ( .A(n[1]), .B(n1251), .Z(n1252) );
  NAND U1644 ( .A(n1253), .B(n1252), .Z(n1254) );
  XNOR U1645 ( .A(n1255), .B(n1254), .Z(n1269) );
  OR U1646 ( .A(n1262), .B(n[2]), .Z(n1256) );
  NAND U1647 ( .A(n1265), .B(n1256), .Z(n1258) );
  ANDN U1648 ( .B(n1258), .A(n1257), .Z(n1259) );
  NANDN U1649 ( .A(n1276), .B(n1259), .Z(n1260) );
  NAND U1650 ( .A(n1261), .B(n1260), .Z(n1270) );
  IV U1651 ( .A(n1270), .Z(n1278) );
  NANDN U1652 ( .A(n1278), .B(n[2]), .Z(n1263) );
  ANDN U1653 ( .B(n1263), .A(n1262), .Z(n1285) );
  ANDN U1654 ( .B(n1264), .A(n1285), .Z(n1283) );
  NAND U1655 ( .A(n1270), .B(n1265), .Z(n1282) );
  XNOR U1656 ( .A(n1283), .B(n1282), .Z(n1289) );
  XOR U1657 ( .A(n[1]), .B(n1266), .Z(n1267) );
  NAND U1658 ( .A(n1270), .B(n1267), .Z(n1268) );
  XNOR U1659 ( .A(n1269), .B(n1268), .Z(n1293) );
  NANDN U1660 ( .A(n1293), .B(\cin[1][2] ), .Z(n1275) );
  XNOR U1661 ( .A(\cin[1][2] ), .B(n1293), .Z(n1273) );
  NAND U1662 ( .A(n1270), .B(n[0]), .Z(n1271) );
  XOR U1663 ( .A(n1272), .B(n1271), .Z(n1296) );
  ANDN U1664 ( .B(\cin[1][1] ), .A(n1296), .Z(n1290) );
  NAND U1665 ( .A(n1273), .B(n1290), .Z(n1274) );
  NAND U1666 ( .A(n1275), .B(n1274), .Z(n1286) );
  NANDN U1667 ( .A(n1277), .B(n1276), .Z(n1281) );
  NANDN U1668 ( .A(n1278), .B(n[3]), .Z(n1280) );
  ANDN U1669 ( .B(n1280), .A(n1279), .Z(n1300) );
  ANDN U1670 ( .B(n1281), .A(n1300), .Z(n1298) );
  NAND U1671 ( .A(n1283), .B(n1282), .Z(n1284) );
  NANDN U1672 ( .A(n1285), .B(n1284), .Z(n1297) );
  XOR U1673 ( .A(n1298), .B(n1297), .Z(n1302) );
  XNOR U1674 ( .A(n1301), .B(n1302), .Z(n1319) );
  XOR U1675 ( .A(n1286), .B(\cin[1][3] ), .Z(n1287) );
  NAND U1676 ( .A(n1294), .B(n1287), .Z(n1288) );
  XNOR U1677 ( .A(n1289), .B(n1288), .Z(n1334) );
  AND U1678 ( .A(n1334), .B(n[3]), .Z(n1315) );
  NOR U1679 ( .A(n[3]), .B(n1334), .Z(n1317) );
  XOR U1680 ( .A(\cin[1][2] ), .B(n1290), .Z(n1291) );
  NAND U1681 ( .A(n1294), .B(n1291), .Z(n1292) );
  XNOR U1682 ( .A(n1293), .B(n1292), .Z(n1325) );
  NOR U1683 ( .A(n[2]), .B(n1325), .Z(n1312) );
  NAND U1684 ( .A(n1294), .B(\cin[1][1] ), .Z(n1295) );
  XOR U1685 ( .A(n1296), .B(n1295), .Z(n1329) );
  ANDN U1686 ( .B(n[1]), .A(n1329), .Z(n1310) );
  AND U1687 ( .A(n1325), .B(n[2]), .Z(n1313) );
  AND U1688 ( .A(n1298), .B(n1297), .Z(n1299) );
  NOR U1689 ( .A(n1300), .B(n1299), .Z(n1306) );
  AND U1690 ( .A(n1302), .B(n1301), .Z(n1303) );
  XOR U1691 ( .A(n1304), .B(n1303), .Z(n1305) );
  XNOR U1692 ( .A(n1306), .B(n1305), .Z(n1320) );
  NAND U1693 ( .A(n1332), .B(n[0]), .Z(n1307) );
  XOR U1694 ( .A(n1308), .B(n1307), .Z(n1336) );
  XNOR U1695 ( .A(n[1]), .B(n1329), .Z(n1309) );
  AND U1696 ( .A(n[0]), .B(n1308), .Z(n1326) );
  NAND U1697 ( .A(n1309), .B(n1326), .Z(n1311) );
  ANDN U1698 ( .B(n1311), .A(n1310), .Z(n1322) );
  OR U1699 ( .A(n1312), .B(n1322), .Z(n1314) );
  ANDN U1700 ( .B(n1314), .A(n1313), .Z(n1330) );
  NANDN U1701 ( .A(n1315), .B(n1330), .Z(n1316) );
  NANDN U1702 ( .A(n1317), .B(n1316), .Z(n1318) );
  NANDN U1703 ( .A(n1319), .B(n1318), .Z(n1321) );
  ANDN U1704 ( .B(n1321), .A(n1320), .Z(n1364) );
  XNOR U1705 ( .A(n[2]), .B(n1322), .Z(n1323) );
  NAND U1706 ( .A(n1332), .B(n1323), .Z(n1324) );
  XNOR U1707 ( .A(n1325), .B(n1324), .Z(n1358) );
  ANDN U1708 ( .B(n[0]), .A(n1336), .Z(n1342) );
  XOR U1709 ( .A(n[1]), .B(n1326), .Z(n1327) );
  NAND U1710 ( .A(n1332), .B(n1327), .Z(n1328) );
  XNOR U1711 ( .A(n1329), .B(n1328), .Z(n1345) );
  XNOR U1712 ( .A(n[3]), .B(n1330), .Z(n1331) );
  NAND U1713 ( .A(n1332), .B(n1331), .Z(n1333) );
  XNOR U1714 ( .A(n1334), .B(n1333), .Z(n1366) );
  AND U1715 ( .A(n[0]), .B(n1367), .Z(n1335) );
  XOR U1716 ( .A(n1336), .B(n1335), .Z(n1337) );
  NAND U1717 ( .A(n1374), .B(n1337), .Z(n1338) );
  NAND U1718 ( .A(n1339), .B(n1338), .Z(n1626) );
  IV U1719 ( .A(n1626), .Z(n1632) );
  OR U1720 ( .A(n1340), .B(n1356), .Z(n1341) );
  ANDN U1721 ( .B(\cin[1][1] ), .A(e[3]), .Z(n1957) );
  ANDN U1722 ( .B(n1341), .A(n1957), .Z(n1348) );
  XOR U1723 ( .A(n1342), .B(n[1]), .Z(n1343) );
  AND U1724 ( .A(n1367), .B(n1343), .Z(n1344) );
  XOR U1725 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U1726 ( .A(n1374), .B(n1346), .Z(n1347) );
  NAND U1727 ( .A(n1348), .B(n1347), .Z(n1591) );
  IV U1728 ( .A(n1591), .Z(n1488) );
  OR U1729 ( .A(n1349), .B(n1356), .Z(n1350) );
  ANDN U1730 ( .B(\cin[1][2] ), .A(e[3]), .Z(n1968) );
  ANDN U1731 ( .B(n1350), .A(n1968), .Z(n1354) );
  NAND U1732 ( .A(n1351), .B(n1367), .Z(n1359) );
  XNOR U1733 ( .A(n1358), .B(n1359), .Z(n1361) );
  AND U1734 ( .A(n1367), .B(n[2]), .Z(n1360) );
  XNOR U1735 ( .A(n1361), .B(n1360), .Z(n1352) );
  NAND U1736 ( .A(n1374), .B(n1352), .Z(n1353) );
  NAND U1737 ( .A(n1354), .B(n1353), .Z(n1624) );
  AND U1738 ( .A(n1624), .B(n1626), .Z(n1458) );
  OR U1739 ( .A(n1356), .B(n1355), .Z(n1357) );
  ANDN U1740 ( .B(\cin[1][3] ), .A(e[3]), .Z(n1977) );
  ANDN U1741 ( .B(n1357), .A(n1977), .Z(n1376) );
  NANDN U1742 ( .A(n1359), .B(n1358), .Z(n1363) );
  NAND U1743 ( .A(n1361), .B(n1360), .Z(n1362) );
  AND U1744 ( .A(n1363), .B(n1362), .Z(n1372) );
  NANDN U1745 ( .A(n1364), .B(n[3]), .Z(n1365) );
  NAND U1746 ( .A(n1366), .B(n1365), .Z(n1370) );
  ANDN U1747 ( .B(n1367), .A(n1366), .Z(n1368) );
  NAND U1748 ( .A(n[3]), .B(n1368), .Z(n1369) );
  NAND U1749 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U1750 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1751 ( .A(n1374), .B(n1373), .Z(n1375) );
  NAND U1752 ( .A(n1376), .B(n1375), .Z(n1605) );
  ANDN U1753 ( .B(n1605), .A(n1488), .Z(n1387) );
  AND U1754 ( .A(n1624), .B(n1605), .Z(n1396) );
  ANDN U1755 ( .B(n[2]), .A(n1396), .Z(n1390) );
  IV U1756 ( .A(n1387), .Z(n1389) );
  NAND U1757 ( .A(n[1]), .B(n1389), .Z(n1380) );
  NANDN U1758 ( .A(n[1]), .B(n1387), .Z(n1378) );
  ANDN U1759 ( .B(n1605), .A(n1632), .Z(n1415) );
  IV U1760 ( .A(n1415), .Z(n1397) );
  OR U1761 ( .A(n[0]), .B(n1397), .Z(n1377) );
  NAND U1762 ( .A(n1378), .B(n1377), .Z(n1379) );
  NAND U1763 ( .A(n1380), .B(n1379), .Z(n1381) );
  NANDN U1764 ( .A(n[2]), .B(n1396), .Z(n1392) );
  NAND U1765 ( .A(n1381), .B(n1392), .Z(n1382) );
  NANDN U1766 ( .A(n1390), .B(n1382), .Z(n1384) );
  NANDN U1767 ( .A(n[3]), .B(n1605), .Z(n1383) );
  AND U1768 ( .A(n1384), .B(n1383), .Z(n1406) );
  AND U1769 ( .A(n[0]), .B(n1397), .Z(n1388) );
  XOR U1770 ( .A(n[1]), .B(n1388), .Z(n1385) );
  NANDN U1771 ( .A(n1406), .B(n1385), .Z(n1386) );
  XNOR U1772 ( .A(n1387), .B(n1386), .Z(n1414) );
  OR U1773 ( .A(n1390), .B(n1393), .Z(n1391) );
  AND U1774 ( .A(n1392), .B(n1391), .Z(n1404) );
  OR U1775 ( .A(n1404), .B(n[3]), .Z(n1425) );
  XOR U1776 ( .A(n[2]), .B(n1393), .Z(n1394) );
  NANDN U1777 ( .A(n1406), .B(n1394), .Z(n1395) );
  XNOR U1778 ( .A(n1396), .B(n1395), .Z(n1426) );
  ANDN U1779 ( .B(n1426), .A(n[2]), .Z(n1403) );
  XNOR U1780 ( .A(n1415), .B(n1406), .Z(n1399) );
  NANDN U1781 ( .A(n[0]), .B(n1397), .Z(n1398) );
  NAND U1782 ( .A(n1399), .B(n1398), .Z(n1416) );
  NAND U1783 ( .A(n[0]), .B(n1416), .Z(n1411) );
  NANDN U1784 ( .A(n[1]), .B(n1411), .Z(n1402) );
  NOR U1785 ( .A(n792), .B(n1411), .Z(n1400) );
  NANDN U1786 ( .A(n1400), .B(n1414), .Z(n1401) );
  AND U1787 ( .A(n1402), .B(n1401), .Z(n1428) );
  NANDN U1788 ( .A(n1403), .B(n1428), .Z(n1409) );
  XOR U1789 ( .A(n1404), .B(n[3]), .Z(n1405) );
  NANDN U1790 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U1791 ( .A(n1407), .B(n1605), .Z(n1444) );
  NANDN U1792 ( .A(n1444), .B(n[3]), .Z(n1408) );
  AND U1793 ( .A(n1409), .B(n1408), .Z(n1410) );
  NANDN U1794 ( .A(n1426), .B(n[2]), .Z(n1424) );
  NAND U1795 ( .A(n1410), .B(n1424), .Z(n1442) );
  NAND U1796 ( .A(n1425), .B(n1442), .Z(n1429) );
  XOR U1797 ( .A(n792), .B(n1411), .Z(n1412) );
  NAND U1798 ( .A(n1429), .B(n1412), .Z(n1413) );
  XNOR U1799 ( .A(n1414), .B(n1413), .Z(n1433) );
  NAND U1800 ( .A(n1591), .B(n1430), .Z(n1417) );
  NAND U1801 ( .A(n1624), .B(n1417), .Z(n1418) );
  XNOR U1802 ( .A(n1433), .B(n1418), .Z(n1471) );
  ANDN U1803 ( .B(n[2]), .A(n1471), .Z(n1463) );
  ANDN U1804 ( .B(n1471), .A(n[2]), .Z(n1462) );
  ANDN U1805 ( .B(n1458), .A(n[0]), .Z(n1419) );
  AND U1806 ( .A(n1624), .B(n1591), .Z(n1431) );
  XOR U1807 ( .A(n1431), .B(n1430), .Z(n1475) );
  OR U1808 ( .A(n1475), .B(n792), .Z(n1461) );
  NAND U1809 ( .A(n1419), .B(n1461), .Z(n1421) );
  ANDN U1810 ( .B(n1475), .A(n[1]), .Z(n1420) );
  ANDN U1811 ( .B(n1421), .A(n1420), .Z(n1422) );
  NANDN U1812 ( .A(n1462), .B(n1422), .Z(n1423) );
  NANDN U1813 ( .A(n1463), .B(n1423), .Z(n1453) );
  OR U1814 ( .A(n1425), .B(n1424), .Z(n1427) );
  ANDN U1815 ( .B(n1427), .A(n1447), .Z(n1446) );
  NAND U1816 ( .A(n1429), .B(n1428), .Z(n1445) );
  XOR U1817 ( .A(n1446), .B(n1445), .Z(n1440) );
  OR U1818 ( .A(n1624), .B(n1440), .Z(n1436) );
  IV U1819 ( .A(n1605), .Z(n1581) );
  NOR U1820 ( .A(n1581), .B(n1440), .Z(n1438) );
  NAND U1821 ( .A(n1431), .B(n1430), .Z(n1432) );
  NANDN U1822 ( .A(n1433), .B(n1432), .Z(n1437) );
  XNOR U1823 ( .A(n1438), .B(n1437), .Z(n1434) );
  NAND U1824 ( .A(n1624), .B(n1434), .Z(n1435) );
  NAND U1825 ( .A(n1436), .B(n1435), .Z(n1483) );
  OR U1826 ( .A(n1453), .B(n1483), .Z(n1452) );
  AND U1827 ( .A(n1438), .B(n1437), .Z(n1439) );
  OR U1828 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1829 ( .A(n1624), .B(n1441), .Z(n1466) );
  NANDN U1830 ( .A(n1442), .B(n[3]), .Z(n1443) );
  AND U1831 ( .A(n1444), .B(n1443), .Z(n1450) );
  AND U1832 ( .A(n1446), .B(n1445), .Z(n1448) );
  NOR U1833 ( .A(n1448), .B(n1447), .Z(n1449) );
  XOR U1834 ( .A(n1450), .B(n1449), .Z(n1465) );
  OR U1835 ( .A(n1466), .B(n1465), .Z(n1451) );
  ANDN U1836 ( .B(n1452), .A(n1451), .Z(n1456) );
  XOR U1837 ( .A(n1453), .B(n1483), .Z(n1454) );
  NANDN U1838 ( .A(n[3]), .B(n1454), .Z(n1455) );
  NAND U1839 ( .A(n1456), .B(n1455), .Z(n1481) );
  NAND U1840 ( .A(n1481), .B(n[0]), .Z(n1457) );
  XNOR U1841 ( .A(n1458), .B(n1457), .Z(n1487) );
  XNOR U1842 ( .A(n[1]), .B(n1475), .Z(n1459) );
  ANDN U1843 ( .B(n[0]), .A(n1458), .Z(n1472) );
  NAND U1844 ( .A(n1459), .B(n1472), .Z(n1460) );
  NAND U1845 ( .A(n1461), .B(n1460), .Z(n1468) );
  NANDN U1846 ( .A(n1462), .B(n1468), .Z(n1464) );
  ANDN U1847 ( .B(n1464), .A(n1463), .Z(n1479) );
  NAND U1848 ( .A(n1466), .B(n1465), .Z(n1467) );
  AND U1849 ( .A(n1530), .B(n1467), .Z(n1517) );
  XOR U1850 ( .A(n[2]), .B(n1468), .Z(n1469) );
  AND U1851 ( .A(n1469), .B(n1481), .Z(n1470) );
  XOR U1852 ( .A(n1471), .B(n1470), .Z(n1492) );
  OR U1853 ( .A(n1492), .B(n793), .Z(n1478) );
  XOR U1854 ( .A(n[1]), .B(n1472), .Z(n1473) );
  NAND U1855 ( .A(n1481), .B(n1473), .Z(n1474) );
  XNOR U1856 ( .A(n1475), .B(n1474), .Z(n1497) );
  XOR U1857 ( .A(n1492), .B(n793), .Z(n1476) );
  NANDN U1858 ( .A(n1489), .B(n1476), .Z(n1477) );
  NAND U1859 ( .A(n1478), .B(n1477), .Z(n1520) );
  XNOR U1860 ( .A(n[3]), .B(n1479), .Z(n1480) );
  NAND U1861 ( .A(n1481), .B(n1480), .Z(n1482) );
  XNOR U1862 ( .A(n1483), .B(n1482), .Z(n1514) );
  AND U1863 ( .A(n1514), .B(n[3]), .Z(n1516) );
  OR U1864 ( .A(n1520), .B(n1516), .Z(n1484) );
  AND U1865 ( .A(n1517), .B(n1484), .Z(n1513) );
  OR U1866 ( .A(n1514), .B(n[3]), .Z(n1485) );
  NAND U1867 ( .A(n1513), .B(n1485), .Z(n1519) );
  NAND U1868 ( .A(n1519), .B(n[0]), .Z(n1486) );
  XOR U1869 ( .A(n1487), .B(n1486), .Z(n1504) );
  IV U1870 ( .A(n1504), .Z(n1493) );
  XNOR U1871 ( .A(n1488), .B(n1493), .Z(n1545) );
  XNOR U1872 ( .A(n[2]), .B(n1489), .Z(n1490) );
  NAND U1873 ( .A(n1519), .B(n1490), .Z(n1491) );
  XNOR U1874 ( .A(n1492), .B(n1491), .Z(n1522) );
  AND U1875 ( .A(n1591), .B(n1493), .Z(n1498) );
  XOR U1876 ( .A(n[1]), .B(n1494), .Z(n1495) );
  NAND U1877 ( .A(n1519), .B(n1495), .Z(n1496) );
  XNOR U1878 ( .A(n1497), .B(n1496), .Z(n1507) );
  NAND U1879 ( .A(n1498), .B(n1507), .Z(n1501) );
  XOR U1880 ( .A(n1498), .B(n1507), .Z(n1499) );
  NAND U1881 ( .A(n1499), .B(n1624), .Z(n1500) );
  AND U1882 ( .A(n1501), .B(n1500), .Z(n1523) );
  XOR U1883 ( .A(n1581), .B(n1523), .Z(n1502) );
  NAND U1884 ( .A(n1591), .B(n1502), .Z(n1503) );
  XNOR U1885 ( .A(n1522), .B(n1503), .Z(n1563) );
  ANDN U1886 ( .B(n[3]), .A(n1563), .Z(n1553) );
  XNOR U1887 ( .A(n1624), .B(n1504), .Z(n1505) );
  AND U1888 ( .A(n1505), .B(n1591), .Z(n1506) );
  XNOR U1889 ( .A(n1507), .B(n1506), .Z(n1570) );
  AND U1890 ( .A(n1570), .B(n[2]), .Z(n1550) );
  NOR U1891 ( .A(n1553), .B(n1550), .Z(n1512) );
  NANDN U1892 ( .A(n1545), .B(n[1]), .Z(n1549) );
  ANDN U1893 ( .B(n1545), .A(n[1]), .Z(n1508) );
  ANDN U1894 ( .B(n1591), .A(n1632), .Z(n1622) );
  ANDN U1895 ( .B(n1622), .A(n[0]), .Z(n1587) );
  OR U1896 ( .A(n1508), .B(n1587), .Z(n1509) );
  AND U1897 ( .A(n1549), .B(n1509), .Z(n1510) );
  NOR U1898 ( .A(n[2]), .B(n1570), .Z(n1551) );
  OR U1899 ( .A(n1510), .B(n1551), .Z(n1511) );
  AND U1900 ( .A(n1512), .B(n1511), .Z(n1535) );
  OR U1901 ( .A(n1513), .B(n794), .Z(n1515) );
  ANDN U1902 ( .B(n1515), .A(n1514), .Z(n1521) );
  NANDN U1903 ( .A(n1517), .B(n1516), .Z(n1518) );
  ANDN U1904 ( .B(n1518), .A(n1521), .Z(n1528) );
  AND U1905 ( .A(n1520), .B(n1519), .Z(n1529) );
  AND U1906 ( .A(n1522), .B(n1605), .Z(n1526) );
  XNOR U1907 ( .A(n1581), .B(n1522), .Z(n1524) );
  ANDN U1908 ( .B(n1524), .A(n1523), .Z(n1525) );
  OR U1909 ( .A(n1526), .B(n1525), .Z(n1527) );
  AND U1910 ( .A(n1527), .B(n1591), .Z(n1532) );
  XOR U1911 ( .A(n1529), .B(n1528), .Z(n1531) );
  XNOR U1912 ( .A(n1532), .B(n1531), .Z(n1557) );
  ANDN U1913 ( .B(n1559), .A(n1557), .Z(n1533) );
  ANDN U1914 ( .B(n1563), .A(n[3]), .Z(n1554) );
  ANDN U1915 ( .B(n1533), .A(n1554), .Z(n1534) );
  NANDN U1916 ( .A(n1535), .B(n1534), .Z(n1568) );
  IV U1917 ( .A(n1622), .Z(n1538) );
  AND U1918 ( .A(n[0]), .B(n1538), .Z(n1547) );
  XOR U1919 ( .A(n[1]), .B(n1547), .Z(n1536) );
  NAND U1920 ( .A(n1568), .B(n1536), .Z(n1537) );
  XOR U1921 ( .A(n1545), .B(n1537), .Z(n1583) );
  NAND U1922 ( .A(n[1]), .B(n1583), .Z(n1544) );
  XNOR U1923 ( .A(n1538), .B(n1568), .Z(n1540) );
  NANDN U1924 ( .A(n[0]), .B(n1538), .Z(n1539) );
  NAND U1925 ( .A(n1540), .B(n1539), .Z(n1588) );
  NOR U1926 ( .A(n[1]), .B(n1583), .Z(n1541) );
  ANDN U1927 ( .B(n1588), .A(n1541), .Z(n1542) );
  NAND U1928 ( .A(n[0]), .B(n1542), .Z(n1543) );
  NAND U1929 ( .A(n1544), .B(n1543), .Z(n1576) );
  XNOR U1930 ( .A(n[1]), .B(n1545), .Z(n1546) );
  NAND U1931 ( .A(n1547), .B(n1546), .Z(n1548) );
  AND U1932 ( .A(n1549), .B(n1548), .Z(n1566) );
  NANDN U1933 ( .A(n1550), .B(n1566), .Z(n1552) );
  ANDN U1934 ( .B(n1552), .A(n1551), .Z(n1560) );
  OR U1935 ( .A(n1553), .B(n1560), .Z(n1555) );
  ANDN U1936 ( .B(n1555), .A(n1554), .Z(n1556) );
  XOR U1937 ( .A(n1557), .B(n1556), .Z(n1558) );
  AND U1938 ( .A(n1568), .B(n1558), .Z(n1618) );
  ANDN U1939 ( .B(n1559), .A(n1618), .Z(n1565) );
  XOR U1940 ( .A(n[3]), .B(n1560), .Z(n1561) );
  NAND U1941 ( .A(n1568), .B(n1561), .Z(n1562) );
  XNOR U1942 ( .A(n1563), .B(n1562), .Z(n1611) );
  NANDN U1943 ( .A(n[3]), .B(n1611), .Z(n1564) );
  AND U1944 ( .A(n1565), .B(n1564), .Z(n1578) );
  XNOR U1945 ( .A(n[2]), .B(n1566), .Z(n1567) );
  NAND U1946 ( .A(n1568), .B(n1567), .Z(n1569) );
  XNOR U1947 ( .A(n1570), .B(n1569), .Z(n1579) );
  NAND U1948 ( .A(n[2]), .B(n1579), .Z(n1577) );
  NOR U1949 ( .A(n[2]), .B(n1579), .Z(n1571) );
  NANDN U1950 ( .A(n1571), .B(n1576), .Z(n1572) );
  AND U1951 ( .A(n1577), .B(n1572), .Z(n1574) );
  NANDN U1952 ( .A(n1611), .B(n[3]), .Z(n1573) );
  NAND U1953 ( .A(n1574), .B(n1573), .Z(n1575) );
  NAND U1954 ( .A(n1578), .B(n1575), .Z(n1603) );
  AND U1955 ( .A(n1576), .B(n1603), .Z(n1600) );
  OR U1956 ( .A(n1578), .B(n1577), .Z(n1580) );
  ANDN U1957 ( .B(n1580), .A(n1602), .Z(n1599) );
  XNOR U1958 ( .A(n1600), .B(n1599), .Z(n1608) );
  AND U1959 ( .A(n1608), .B(n1605), .Z(n1597) );
  XNOR U1960 ( .A(n1581), .B(n1608), .Z(n1595) );
  AND U1961 ( .A(n[1]), .B(n1603), .Z(n1585) );
  AND U1962 ( .A(n[0]), .B(n1603), .Z(n1586) );
  AND U1963 ( .A(n1588), .B(n1586), .Z(n1582) );
  XNOR U1964 ( .A(n1583), .B(n1582), .Z(n1584) );
  XNOR U1965 ( .A(n1585), .B(n1584), .Z(n1628) );
  NANDN U1966 ( .A(n1628), .B(n1624), .Z(n1594) );
  XNOR U1967 ( .A(n1628), .B(n1624), .Z(n1592) );
  XOR U1968 ( .A(n1588), .B(n1586), .Z(n1590) );
  NAND U1969 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U1970 ( .A(n1590), .B(n1589), .Z(n1621) );
  AND U1971 ( .A(n1621), .B(n1591), .Z(n1623) );
  NAND U1972 ( .A(n1592), .B(n1623), .Z(n1593) );
  AND U1973 ( .A(n1594), .B(n1593), .Z(n1604) );
  ANDN U1974 ( .B(n1595), .A(n1604), .Z(n1596) );
  OR U1975 ( .A(n1597), .B(n1596), .Z(n1598) );
  AND U1976 ( .A(n1598), .B(n1626), .Z(n1615) );
  NANDN U1977 ( .A(n1600), .B(n1599), .Z(n1601) );
  NANDN U1978 ( .A(n1602), .B(n1601), .Z(n1610) );
  ANDN U1979 ( .B(n1603), .A(n794), .Z(n1612) );
  XNOR U1980 ( .A(n1611), .B(n1612), .Z(n1609) );
  XNOR U1981 ( .A(n1615), .B(n1616), .Z(n1631) );
  XNOR U1982 ( .A(n1605), .B(n1604), .Z(n1606) );
  ANDN U1983 ( .B(n1606), .A(n1632), .Z(n1607) );
  XNOR U1984 ( .A(n1608), .B(n1607), .Z(n1644) );
  NOR U1985 ( .A(n[3]), .B(n1644), .Z(n1636) );
  NAND U1986 ( .A(n1610), .B(n1609), .Z(n1614) );
  NANDN U1987 ( .A(n1612), .B(n1611), .Z(n1613) );
  AND U1988 ( .A(n1614), .B(n1613), .Z(n1620) );
  AND U1989 ( .A(n1616), .B(n1615), .Z(n1617) );
  XNOR U1990 ( .A(n1618), .B(n1617), .Z(n1619) );
  XNOR U1991 ( .A(n1620), .B(n1619), .Z(n1639) );
  XOR U1992 ( .A(n1622), .B(n1621), .Z(n1653) );
  OR U1993 ( .A(n[0]), .B(n[1]), .Z(n2233) );
  AND U1994 ( .A(n1644), .B(n[3]), .Z(n1630) );
  XOR U1995 ( .A(n1624), .B(n1623), .Z(n1625) );
  NAND U1996 ( .A(n1626), .B(n1625), .Z(n1627) );
  XNOR U1997 ( .A(n1628), .B(n1627), .Z(n1648) );
  NAND U1998 ( .A(n1651), .B(n[0]), .Z(n1629) );
  XOR U1999 ( .A(n1632), .B(n1629), .Z(n1655) );
  NOR U2000 ( .A(n1631), .B(n1630), .Z(n1638) );
  NANDN U2001 ( .A(n1653), .B(n[1]), .Z(n1635) );
  XNOR U2002 ( .A(n[1]), .B(n1653), .Z(n1633) );
  AND U2003 ( .A(n[0]), .B(n1632), .Z(n1649) );
  NAND U2004 ( .A(n1633), .B(n1649), .Z(n1634) );
  AND U2005 ( .A(n1635), .B(n1634), .Z(n1645) );
  OR U2006 ( .A(n1636), .B(n1641), .Z(n1637) );
  NAND U2007 ( .A(n1638), .B(n1637), .Z(n1640) );
  ANDN U2008 ( .B(n1640), .A(n1639), .Z(n1656) );
  XNOR U2009 ( .A(n[3]), .B(n1641), .Z(n1642) );
  NAND U2010 ( .A(n1651), .B(n1642), .Z(n1643) );
  XNOR U2011 ( .A(n1644), .B(n1643), .Z(n1658) );
  XNOR U2012 ( .A(n[2]), .B(n1645), .Z(n1646) );
  NAND U2013 ( .A(n1651), .B(n1646), .Z(n1647) );
  XNOR U2014 ( .A(n1648), .B(n1647), .Z(n1664) );
  XOR U2015 ( .A(n[1]), .B(n1649), .Z(n1650) );
  NAND U2016 ( .A(n1651), .B(n1650), .Z(n1652) );
  XOR U2017 ( .A(n1653), .B(n1652), .Z(n1783) );
  NAND U2018 ( .A(n1781), .B(n[0]), .Z(n1654) );
  XNOR U2019 ( .A(n1655), .B(n1654), .Z(n1950) );
  NAND U2020 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1950), .Z(n1910) );
  NANDN U2021 ( .A(n1656), .B(n[3]), .Z(n1657) );
  NAND U2022 ( .A(n1658), .B(n1657), .Z(n1661) );
  ANDN U2023 ( .B(n1781), .A(n1658), .Z(n1659) );
  NAND U2024 ( .A(n[3]), .B(n1659), .Z(n1660) );
  NAND U2025 ( .A(n1661), .B(n1660), .Z(n1668) );
  ANDN U2026 ( .B(n1781), .A(n1662), .Z(n1663) );
  XOR U2027 ( .A(n1664), .B(n1663), .Z(n1690) );
  AND U2028 ( .A(n1781), .B(n[2]), .Z(n1689) );
  NAND U2029 ( .A(n1690), .B(n1689), .Z(n1666) );
  NAND U2030 ( .A(n1664), .B(n1663), .Z(n1665) );
  NAND U2031 ( .A(n1666), .B(n1665), .Z(n1667) );
  XNOR U2032 ( .A(n1668), .B(n1667), .Z(n1975) );
  NAND U2033 ( .A(\cin[1][1] ), .B(n1975), .Z(n1677) );
  NAND U2034 ( .A(n2275), .B(n1975), .Z(n1707) );
  NAND U2035 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1975), .Z(n1669) );
  AND U2036 ( .A(n[0]), .B(n1669), .Z(n1676) );
  ANDN U2037 ( .B(n[0]), .A(n1707), .Z(n1670) );
  NAND U2038 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n1670), .Z(n1672) );
  NANDN U2039 ( .A(n1670), .B(n1669), .Z(n1671) );
  NAND U2040 ( .A(n1672), .B(n1671), .Z(n1688) );
  NAND U2041 ( .A(n[0]), .B(n1688), .Z(n1683) );
  NANDN U2042 ( .A(n[1]), .B(n1683), .Z(n1675) );
  NOR U2043 ( .A(n792), .B(n1683), .Z(n1673) );
  NANDN U2044 ( .A(n1673), .B(n1686), .Z(n1674) );
  AND U2045 ( .A(n1675), .B(n1674), .Z(n1693) );
  NAND U2046 ( .A(\cin[1][2] ), .B(n1975), .Z(n1679) );
  NANDN U2047 ( .A(n1707), .B(n1712), .Z(n1680) );
  NANDN U2048 ( .A(n1708), .B(n1680), .Z(n1682) );
  NANDN U2049 ( .A(n1712), .B(n[3]), .Z(n1681) );
  NAND U2050 ( .A(n1682), .B(n1681), .Z(n1695) );
  XOR U2051 ( .A(n792), .B(n1683), .Z(n1684) );
  NANDN U2052 ( .A(n1695), .B(n1684), .Z(n1685) );
  XNOR U2053 ( .A(n1686), .B(n1685), .Z(n1698) );
  NANDN U2054 ( .A(n1695), .B(n[0]), .Z(n1687) );
  XNOR U2055 ( .A(n1688), .B(n1687), .Z(n1720) );
  XOR U2056 ( .A(\cin[1][2] ), .B(n1699), .Z(n1691) );
  XNOR U2057 ( .A(n1690), .B(n1689), .Z(n1967) );
  IV U2058 ( .A(n1967), .Z(n1744) );
  ANDN U2059 ( .B(n1691), .A(n1744), .Z(n1692) );
  XNOR U2060 ( .A(n1698), .B(n1692), .Z(n1736) );
  XOR U2061 ( .A(n1693), .B(n[2]), .Z(n1694) );
  NANDN U2062 ( .A(n1695), .B(n1694), .Z(n1696) );
  XNOR U2063 ( .A(n1697), .B(n1696), .Z(n1718) );
  AND U2064 ( .A(\cin[1][3] ), .B(n1718), .Z(n1705) );
  XOR U2065 ( .A(\cin[1][3] ), .B(n1718), .Z(n1703) );
  NAND U2066 ( .A(\cin[1][2] ), .B(n1698), .Z(n1702) );
  XOR U2067 ( .A(\cin[1][2] ), .B(n1698), .Z(n1700) );
  NAND U2068 ( .A(n1700), .B(n1699), .Z(n1701) );
  AND U2069 ( .A(n1702), .B(n1701), .Z(n1715) );
  ANDN U2070 ( .B(n1703), .A(n1715), .Z(n1704) );
  OR U2071 ( .A(n1705), .B(n1704), .Z(n1706) );
  AND U2072 ( .A(n1706), .B(n1967), .Z(n1714) );
  OR U2073 ( .A(n1707), .B(n1708), .Z(n1710) );
  NAND U2074 ( .A(n[3]), .B(n1708), .Z(n1709) );
  AND U2075 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U2076 ( .A(n1712), .B(n1711), .Z(n1713) );
  AND U2077 ( .A(n1714), .B(n1713), .Z(n1760) );
  XNOR U2078 ( .A(\cin[1][3] ), .B(n1715), .Z(n1716) );
  NAND U2079 ( .A(n1967), .B(n1716), .Z(n1717) );
  XNOR U2080 ( .A(n1718), .B(n1717), .Z(n1743) );
  ANDN U2081 ( .B(n1743), .A(n[3]), .Z(n1753) );
  NOR U2082 ( .A(n1760), .B(n1753), .Z(n1728) );
  NANDN U2083 ( .A(n1743), .B(n[3]), .Z(n1755) );
  AND U2084 ( .A(n1736), .B(n[2]), .Z(n1738) );
  ANDN U2085 ( .B(n1755), .A(n1738), .Z(n1726) );
  NOR U2086 ( .A(n[2]), .B(n1736), .Z(n1739) );
  NAND U2087 ( .A(n1967), .B(\cin[1][1] ), .Z(n1719) );
  XOR U2088 ( .A(n1720), .B(n1719), .Z(n1751) );
  NANDN U2089 ( .A(n[1]), .B(n1751), .Z(n1723) );
  NAND U2090 ( .A(n1967), .B(n2488), .Z(n1721) );
  OR U2091 ( .A(n1721), .B(n1732), .Z(n1722) );
  AND U2092 ( .A(n1723), .B(n1722), .Z(n1724) );
  NANDN U2093 ( .A(n1739), .B(n1724), .Z(n1725) );
  AND U2094 ( .A(n1726), .B(n1725), .Z(n1727) );
  ANDN U2095 ( .B(n1728), .A(n1727), .Z(n1729) );
  NANDN U2096 ( .A(n1757), .B(n1729), .Z(n1749) );
  NAND U2097 ( .A(n1967), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1730)
         );
  AND U2098 ( .A(n[0]), .B(n1730), .Z(n1747) );
  XNOR U2099 ( .A(n[1]), .B(n1751), .Z(n1731) );
  NAND U2100 ( .A(n1747), .B(n1731), .Z(n1733) );
  ANDN U2101 ( .B(n1733), .A(n1732), .Z(n1737) );
  XNOR U2102 ( .A(n[2]), .B(n1737), .Z(n1734) );
  NAND U2103 ( .A(n1749), .B(n1734), .Z(n1735) );
  XNOR U2104 ( .A(n1736), .B(n1735), .Z(n1766) );
  NANDN U2105 ( .A(n1738), .B(n1737), .Z(n1740) );
  ANDN U2106 ( .B(n1740), .A(n1739), .Z(n1752) );
  XOR U2107 ( .A(n[3]), .B(n1752), .Z(n1741) );
  NAND U2108 ( .A(n1749), .B(n1741), .Z(n1742) );
  XNOR U2109 ( .A(n1743), .B(n1742), .Z(n1789) );
  ANDN U2110 ( .B(n[3]), .A(n1789), .Z(n1785) );
  IV U2111 ( .A(n1749), .Z(n1759) );
  ANDN U2112 ( .B(n[0]), .A(n1759), .Z(n1746) );
  ANDN U2113 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n1744), .Z(n1745) );
  XOR U2114 ( .A(n1746), .B(n1745), .Z(n1772) );
  ANDN U2115 ( .B(n[0]), .A(n1772), .Z(n1767) );
  XOR U2116 ( .A(n[1]), .B(n1747), .Z(n1748) );
  NAND U2117 ( .A(n1749), .B(n1748), .Z(n1750) );
  XNOR U2118 ( .A(n1751), .B(n1750), .Z(n1770) );
  NANDN U2119 ( .A(n1785), .B(n1792), .Z(n1762) );
  NANDN U2120 ( .A(n1753), .B(n1752), .Z(n1754) );
  AND U2121 ( .A(n1755), .B(n1754), .Z(n1756) );
  XNOR U2122 ( .A(n1757), .B(n1756), .Z(n1758) );
  NANDN U2123 ( .A(n1759), .B(n1758), .Z(n1819) );
  ANDN U2124 ( .B(n1819), .A(n1760), .Z(n1786) );
  NANDN U2125 ( .A(n[3]), .B(n1789), .Z(n1761) );
  NAND U2126 ( .A(n1786), .B(n1761), .Z(n1791) );
  ANDN U2127 ( .B(n1762), .A(n1791), .Z(n1787) );
  XOR U2128 ( .A(n1763), .B(n[2]), .Z(n1764) );
  NANDN U2129 ( .A(n1787), .B(n1764), .Z(n1765) );
  XNOR U2130 ( .A(n1766), .B(n1765), .Z(n1796) );
  ANDN U2131 ( .B(\cin[1][3] ), .A(n1796), .Z(n1778) );
  XNOR U2132 ( .A(\cin[1][3] ), .B(n1796), .Z(n1776) );
  XOR U2133 ( .A(n1767), .B(n[1]), .Z(n1768) );
  NANDN U2134 ( .A(n1787), .B(n1768), .Z(n1769) );
  XNOR U2135 ( .A(n1770), .B(n1769), .Z(n1800) );
  NAND U2136 ( .A(\cin[1][2] ), .B(n1800), .Z(n1775) );
  XOR U2137 ( .A(\cin[1][2] ), .B(n1800), .Z(n1773) );
  NANDN U2138 ( .A(n1787), .B(n[0]), .Z(n1771) );
  XOR U2139 ( .A(n1772), .B(n1771), .Z(n1802) );
  ANDN U2140 ( .B(\cin[1][1] ), .A(n1802), .Z(n1797) );
  NAND U2141 ( .A(n1773), .B(n1797), .Z(n1774) );
  AND U2142 ( .A(n1775), .B(n1774), .Z(n1793) );
  ANDN U2143 ( .B(n1776), .A(n1793), .Z(n1777) );
  OR U2144 ( .A(n1778), .B(n1777), .Z(n1784) );
  XOR U2145 ( .A(n[1]), .B(n1779), .Z(n1780) );
  NAND U2146 ( .A(n1781), .B(n1780), .Z(n1782) );
  XNOR U2147 ( .A(n1783), .B(n1782), .Z(n1956) );
  ANDN U2148 ( .B(n1784), .A(n1956), .Z(n1817) );
  NANDN U2149 ( .A(n1786), .B(n1785), .Z(n1790) );
  NANDN U2150 ( .A(n1787), .B(n[3]), .Z(n1788) );
  AND U2151 ( .A(n1789), .B(n1788), .Z(n1815) );
  ANDN U2152 ( .B(n1790), .A(n1815), .Z(n1813) );
  NANDN U2153 ( .A(n1792), .B(n1791), .Z(n1812) );
  XOR U2154 ( .A(n1813), .B(n1812), .Z(n1816) );
  XOR U2155 ( .A(n1817), .B(n1816), .Z(n1831) );
  XNOR U2156 ( .A(\cin[1][3] ), .B(n1793), .Z(n1794) );
  NANDN U2157 ( .A(n1956), .B(n1794), .Z(n1795) );
  XNOR U2158 ( .A(n1796), .B(n1795), .Z(n1836) );
  XOR U2159 ( .A(\cin[1][2] ), .B(n1797), .Z(n1798) );
  ANDN U2160 ( .B(n1798), .A(n1956), .Z(n1799) );
  XNOR U2161 ( .A(n1800), .B(n1799), .Z(n1849) );
  AND U2162 ( .A(n1849), .B(n[2]), .Z(n1828) );
  NANDN U2163 ( .A(n1956), .B(\cin[1][1] ), .Z(n1801) );
  XOR U2164 ( .A(n1802), .B(n1801), .Z(n1844) );
  ANDN U2165 ( .B(n1844), .A(n[1]), .Z(n1806) );
  ANDN U2166 ( .B(n2488), .A(n1956), .Z(n1803) );
  OR U2167 ( .A(n1844), .B(n792), .Z(n1827) );
  NAND U2168 ( .A(n1803), .B(n1827), .Z(n1804) );
  ANDN U2169 ( .B(n793), .A(n1849), .Z(n1829) );
  ANDN U2170 ( .B(n1804), .A(n1829), .Z(n1805) );
  NANDN U2171 ( .A(n1806), .B(n1805), .Z(n1807) );
  NANDN U2172 ( .A(n1828), .B(n1807), .Z(n1808) );
  NAND U2173 ( .A(n1836), .B(n1808), .Z(n1811) );
  XOR U2174 ( .A(n1836), .B(n1808), .Z(n1809) );
  NAND U2175 ( .A(n[3]), .B(n1809), .Z(n1810) );
  NAND U2176 ( .A(n1811), .B(n1810), .Z(n1822) );
  AND U2177 ( .A(n1813), .B(n1812), .Z(n1814) );
  NOR U2178 ( .A(n1815), .B(n1814), .Z(n1821) );
  AND U2179 ( .A(n1817), .B(n1816), .Z(n1818) );
  XOR U2180 ( .A(n1819), .B(n1818), .Z(n1820) );
  XNOR U2181 ( .A(n1821), .B(n1820), .Z(n1832) );
  ANDN U2182 ( .B(n1822), .A(n1832), .Z(n1823) );
  NANDN U2183 ( .A(n1831), .B(n1823), .Z(n1847) );
  IV U2184 ( .A(n1847), .Z(n1838) );
  XNOR U2185 ( .A(n[1]), .B(n1844), .Z(n1825) );
  NANDN U2186 ( .A(n1956), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n1824)
         );
  AND U2187 ( .A(n[0]), .B(n1824), .Z(n1841) );
  NAND U2188 ( .A(n1825), .B(n1841), .Z(n1826) );
  AND U2189 ( .A(n1827), .B(n1826), .Z(n1845) );
  NANDN U2190 ( .A(n1828), .B(n1845), .Z(n1830) );
  ANDN U2191 ( .B(n1830), .A(n1829), .Z(n1833) );
  XOR U2192 ( .A(n[3]), .B(n1833), .Z(n1834) );
  NAND U2193 ( .A(n1847), .B(n1834), .Z(n1835) );
  XNOR U2194 ( .A(n1836), .B(n1835), .Z(n1865) );
  OR U2195 ( .A(n1865), .B(n[3]), .Z(n1837) );
  AND U2196 ( .A(n1863), .B(n1837), .Z(n1858) );
  AND U2197 ( .A(n1865), .B(n[3]), .Z(n1862) );
  ANDN U2198 ( .B(n[0]), .A(n1838), .Z(n1840) );
  ANDN U2199 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n1956), .Z(n1839) );
  XOR U2200 ( .A(n1840), .B(n1839), .Z(n1876) );
  ANDN U2201 ( .B(n[0]), .A(n1876), .Z(n1870) );
  XOR U2202 ( .A(n1841), .B(n[1]), .Z(n1842) );
  NAND U2203 ( .A(n1847), .B(n1842), .Z(n1843) );
  XNOR U2204 ( .A(n1844), .B(n1843), .Z(n1873) );
  XNOR U2205 ( .A(n[2]), .B(n1845), .Z(n1846) );
  NAND U2206 ( .A(n1847), .B(n1846), .Z(n1848) );
  XNOR U2207 ( .A(n1849), .B(n1848), .Z(n1854) );
  OR U2208 ( .A(n1854), .B(n[2]), .Z(n1850) );
  NAND U2209 ( .A(n1856), .B(n1850), .Z(n1851) );
  AND U2210 ( .A(n1854), .B(n[2]), .Z(n1857) );
  ANDN U2211 ( .B(n1851), .A(n1857), .Z(n1852) );
  NANDN U2212 ( .A(n1862), .B(n1852), .Z(n1853) );
  AND U2213 ( .A(n1858), .B(n1853), .Z(n1864) );
  NANDN U2214 ( .A(n1864), .B(n[2]), .Z(n1855) );
  ANDN U2215 ( .B(n1855), .A(n1854), .Z(n1861) );
  IV U2216 ( .A(n1864), .Z(n1874) );
  AND U2217 ( .A(n1856), .B(n1874), .Z(n1869) );
  NANDN U2218 ( .A(n1858), .B(n1857), .Z(n1859) );
  ANDN U2219 ( .B(n1859), .A(n1861), .Z(n1868) );
  NANDN U2220 ( .A(n1869), .B(n1868), .Z(n1860) );
  NANDN U2221 ( .A(n1861), .B(n1860), .Z(n1881) );
  NANDN U2222 ( .A(n1863), .B(n1862), .Z(n1867) );
  NANDN U2223 ( .A(n1864), .B(n[3]), .Z(n1866) );
  ANDN U2224 ( .B(n1866), .A(n1865), .Z(n1883) );
  ANDN U2225 ( .B(n1867), .A(n1883), .Z(n1880) );
  XOR U2226 ( .A(n1869), .B(n1868), .Z(n1891) );
  XOR U2227 ( .A(n[1]), .B(n1870), .Z(n1871) );
  NAND U2228 ( .A(n1874), .B(n1871), .Z(n1872) );
  XNOR U2229 ( .A(n1873), .B(n1872), .Z(n1895) );
  NAND U2230 ( .A(\cin[1][2] ), .B(n1895), .Z(n1879) );
  XOR U2231 ( .A(\cin[1][2] ), .B(n1895), .Z(n1877) );
  NAND U2232 ( .A(n1874), .B(n[0]), .Z(n1875) );
  XNOR U2233 ( .A(n1876), .B(n1875), .Z(n1898) );
  AND U2234 ( .A(\cin[1][1] ), .B(n1898), .Z(n1892) );
  NAND U2235 ( .A(n1877), .B(n1892), .Z(n1878) );
  NAND U2236 ( .A(n1879), .B(n1878), .Z(n1888) );
  AND U2237 ( .A(n1906), .B(n1905), .Z(n1885) );
  NAND U2238 ( .A(n1881), .B(n1880), .Z(n1882) );
  NANDN U2239 ( .A(n1883), .B(n1882), .Z(n1884) );
  XNOR U2240 ( .A(n1885), .B(n1884), .Z(n1886) );
  XNOR U2241 ( .A(n1887), .B(n1886), .Z(n1923) );
  XOR U2242 ( .A(n1888), .B(\cin[1][3] ), .Z(n1889) );
  NAND U2243 ( .A(n1950), .B(n1889), .Z(n1890) );
  XNOR U2244 ( .A(n1891), .B(n1890), .Z(n1933) );
  ANDN U2245 ( .B(n794), .A(n1933), .Z(n1941) );
  ANDN U2246 ( .B(n1923), .A(n1941), .Z(n1909) );
  XOR U2247 ( .A(\cin[1][2] ), .B(n1892), .Z(n1893) );
  NAND U2248 ( .A(n1950), .B(n1893), .Z(n1894) );
  XNOR U2249 ( .A(n1895), .B(n1894), .Z(n1927) );
  OR U2250 ( .A(n1927), .B(n793), .Z(n1896) );
  AND U2251 ( .A(n1933), .B(n[3]), .Z(n1939) );
  ANDN U2252 ( .B(n1896), .A(n1939), .Z(n1904) );
  NAND U2253 ( .A(n1950), .B(\cin[1][1] ), .Z(n1897) );
  XNOR U2254 ( .A(n1898), .B(n1897), .Z(n1913) );
  ANDN U2255 ( .B(n1913), .A(n[1]), .Z(n1899) );
  OR U2256 ( .A(n1899), .B(n2488), .Z(n1900) );
  AND U2257 ( .A(n1917), .B(n1900), .Z(n1902) );
  XOR U2258 ( .A(n793), .B(n1927), .Z(n1901) );
  NANDN U2259 ( .A(n1902), .B(n1901), .Z(n1903) );
  NAND U2260 ( .A(n1904), .B(n1903), .Z(n1907) );
  XNOR U2261 ( .A(n1906), .B(n1905), .Z(n1938) );
  AND U2262 ( .A(n1907), .B(n1938), .Z(n1908) );
  NAND U2263 ( .A(n1909), .B(n1908), .Z(n1931) );
  AND U2264 ( .A(n[0]), .B(n1910), .Z(n1914) );
  XOR U2265 ( .A(n1914), .B(n[1]), .Z(n1911) );
  NAND U2266 ( .A(n1931), .B(n1911), .Z(n1912) );
  XNOR U2267 ( .A(n1913), .B(n1912), .Z(n1962) );
  NAND U2268 ( .A(n[2]), .B(n1971), .Z(n1922) );
  XNOR U2269 ( .A(n[1]), .B(n1913), .Z(n1915) );
  NAND U2270 ( .A(n1915), .B(n1914), .Z(n1916) );
  NAND U2271 ( .A(n1917), .B(n1916), .Z(n1925) );
  XOR U2272 ( .A(n[2]), .B(n1925), .Z(n1918) );
  AND U2273 ( .A(n1931), .B(n1918), .Z(n1919) );
  XOR U2274 ( .A(n1927), .B(n1919), .Z(n1983) );
  XOR U2275 ( .A(n1971), .B(n[2]), .Z(n1920) );
  NANDN U2276 ( .A(n1983), .B(n1920), .Z(n1921) );
  NAND U2277 ( .A(n1922), .B(n1921), .Z(n1934) );
  OR U2278 ( .A(n1934), .B(n[3]), .Z(n1924) );
  AND U2279 ( .A(n1924), .B(n1923), .Z(n1937) );
  NAND U2280 ( .A(n[2]), .B(n1925), .Z(n1929) );
  ANDN U2281 ( .B(n793), .A(n1925), .Z(n1926) );
  OR U2282 ( .A(n1927), .B(n1926), .Z(n1928) );
  AND U2283 ( .A(n1929), .B(n1928), .Z(n1940) );
  XNOR U2284 ( .A(n[3]), .B(n1940), .Z(n1930) );
  NAND U2285 ( .A(n1931), .B(n1930), .Z(n1932) );
  XNOR U2286 ( .A(n1933), .B(n1932), .Z(n1989) );
  XOR U2287 ( .A(n1934), .B(n[3]), .Z(n1935) );
  NANDN U2288 ( .A(n1989), .B(n1935), .Z(n1936) );
  NAND U2289 ( .A(n1937), .B(n1936), .Z(n1945) );
  NOR U2290 ( .A(n1939), .B(n1938), .Z(n1943) );
  OR U2291 ( .A(n1941), .B(n1940), .Z(n1942) );
  NAND U2292 ( .A(n1943), .B(n1942), .Z(n1944) );
  NANDN U2293 ( .A(n1945), .B(n1944), .Z(n1986) );
  AND U2294 ( .A(n[0]), .B(n1986), .Z(n1947) );
  XOR U2295 ( .A(n1947), .B(n1946), .Z(n1948) );
  NAND U2296 ( .A(n1992), .B(n1948), .Z(n1955) );
  ANDN U2297 ( .B(n1949), .A(e[1]), .Z(n1976) );
  NAND U2298 ( .A(n1976), .B(n1950), .Z(n1953) );
  NANDN U2299 ( .A(e[2]), .B(n1951), .Z(n1952) );
  NAND U2300 ( .A(n1953), .B(n1952), .Z(n1954) );
  ANDN U2301 ( .B(n1955), .A(n1954), .Z(n2235) );
  NANDN U2302 ( .A(n1956), .B(n1976), .Z(n1959) );
  NANDN U2303 ( .A(e[2]), .B(n1957), .Z(n1958) );
  NAND U2304 ( .A(n1959), .B(n1958), .Z(n1966) );
  XOR U2305 ( .A(n1960), .B(n[1]), .Z(n1961) );
  AND U2306 ( .A(n1986), .B(n1961), .Z(n1963) );
  XOR U2307 ( .A(n1963), .B(n1962), .Z(n1964) );
  NAND U2308 ( .A(n1992), .B(n1964), .Z(n1965) );
  NANDN U2309 ( .A(n1966), .B(n1965), .Z(n2198) );
  NAND U2310 ( .A(n1967), .B(n1976), .Z(n1970) );
  NANDN U2311 ( .A(e[2]), .B(n1968), .Z(n1969) );
  NAND U2312 ( .A(n1970), .B(n1969), .Z(n1974) );
  AND U2313 ( .A(n1986), .B(n[2]), .Z(n1980) );
  AND U2314 ( .A(n1971), .B(n1986), .Z(n1982) );
  XNOR U2315 ( .A(n1983), .B(n1982), .Z(n1981) );
  XNOR U2316 ( .A(n1980), .B(n1981), .Z(n1972) );
  NAND U2317 ( .A(n1992), .B(n1972), .Z(n1973) );
  NANDN U2318 ( .A(n1974), .B(n1973), .Z(n2227) );
  ANDN U2319 ( .B(n2227), .A(n2235), .Z(n2073) );
  NAND U2320 ( .A(n1976), .B(n1975), .Z(n1979) );
  NANDN U2321 ( .A(e[2]), .B(n1977), .Z(n1978) );
  NAND U2322 ( .A(n1979), .B(n1978), .Z(n1994) );
  NAND U2323 ( .A(n1981), .B(n1980), .Z(n1985) );
  NANDN U2324 ( .A(n1983), .B(n1982), .Z(n1984) );
  AND U2325 ( .A(n1985), .B(n1984), .Z(n1988) );
  NAND U2326 ( .A(n[3]), .B(n1986), .Z(n1987) );
  XNOR U2327 ( .A(n1988), .B(n1987), .Z(n1990) );
  XOR U2328 ( .A(n1990), .B(n1989), .Z(n1991) );
  NAND U2329 ( .A(n1992), .B(n1991), .Z(n1993) );
  NANDN U2330 ( .A(n1994), .B(n1993), .Z(n2191) );
  NANDN U2331 ( .A(n[3]), .B(n2191), .Z(n2025) );
  AND U2332 ( .A(n2227), .B(n2191), .Z(n2006) );
  ANDN U2333 ( .B(n[2]), .A(n2006), .Z(n2000) );
  IV U2334 ( .A(n2198), .Z(n2107) );
  ANDN U2335 ( .B(n2191), .A(n2107), .Z(n2016) );
  ANDN U2336 ( .B(n2191), .A(n2235), .Z(n1995) );
  ANDN U2337 ( .B(n1995), .A(n[0]), .Z(n2044) );
  AND U2338 ( .A(n2006), .B(n793), .Z(n2001) );
  IV U2339 ( .A(n1995), .Z(n2009) );
  AND U2340 ( .A(n[0]), .B(n2009), .Z(n2012) );
  OR U2341 ( .A(n2012), .B(n[1]), .Z(n1999) );
  AND U2342 ( .A(n2012), .B(n[1]), .Z(n1997) );
  IV U2343 ( .A(n2016), .Z(n1996) );
  OR U2344 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U2345 ( .A(n1999), .B(n1998), .Z(n2003) );
  OR U2346 ( .A(n2000), .B(n2003), .Z(n2002) );
  ANDN U2347 ( .B(n2002), .A(n2001), .Z(n2026) );
  XOR U2348 ( .A(n[2]), .B(n2003), .Z(n2004) );
  AND U2349 ( .A(n2004), .B(n2014), .Z(n2005) );
  XNOR U2350 ( .A(n2006), .B(n2005), .Z(n2031) );
  NAND U2351 ( .A(n[2]), .B(n2031), .Z(n2008) );
  NOR U2352 ( .A(n794), .B(n2024), .Z(n2007) );
  ANDN U2353 ( .B(n2008), .A(n2007), .Z(n2022) );
  XOR U2354 ( .A(n[2]), .B(n2031), .Z(n2020) );
  XNOR U2355 ( .A(n2009), .B(n2014), .Z(n2011) );
  NANDN U2356 ( .A(n[0]), .B(n2009), .Z(n2010) );
  NAND U2357 ( .A(n2011), .B(n2010), .Z(n2045) );
  NAND U2358 ( .A(n[0]), .B(n2045), .Z(n2038) );
  NANDN U2359 ( .A(n[1]), .B(n2038), .Z(n2019) );
  NOR U2360 ( .A(n792), .B(n2038), .Z(n2017) );
  XOR U2361 ( .A(n[1]), .B(n2012), .Z(n2013) );
  NAND U2362 ( .A(n2014), .B(n2013), .Z(n2015) );
  XNOR U2363 ( .A(n2016), .B(n2015), .Z(n2041) );
  NANDN U2364 ( .A(n2017), .B(n2041), .Z(n2018) );
  AND U2365 ( .A(n2019), .B(n2018), .Z(n2029) );
  NAND U2366 ( .A(n2020), .B(n2029), .Z(n2021) );
  NAND U2367 ( .A(n2022), .B(n2021), .Z(n2028) );
  NANDN U2368 ( .A(n2028), .B(n[3]), .Z(n2023) );
  AND U2369 ( .A(n2024), .B(n2023), .Z(n2035) );
  OR U2370 ( .A(n2026), .B(n2025), .Z(n2027) );
  AND U2371 ( .A(n2028), .B(n2027), .Z(n2042) );
  ANDN U2372 ( .B(n2029), .A(n2042), .Z(n2037) );
  ANDN U2373 ( .B(n[2]), .A(n2042), .Z(n2030) );
  NANDN U2374 ( .A(n2037), .B(n2036), .Z(n2033) );
  NOR U2375 ( .A(n2031), .B(n2030), .Z(n2032) );
  ANDN U2376 ( .B(n2033), .A(n2032), .Z(n2034) );
  XNOR U2377 ( .A(n2035), .B(n2034), .Z(n2071) );
  XNOR U2378 ( .A(n2037), .B(n2036), .Z(n2051) );
  IV U2379 ( .A(n2227), .Z(n2117) );
  XOR U2380 ( .A(n2038), .B(n792), .Z(n2039) );
  NANDN U2381 ( .A(n2042), .B(n2039), .Z(n2040) );
  XNOR U2382 ( .A(n2041), .B(n2040), .Z(n2059) );
  NANDN U2383 ( .A(n2117), .B(n2059), .Z(n2048) );
  NANDN U2384 ( .A(n2042), .B(n[0]), .Z(n2043) );
  XNOR U2385 ( .A(n2045), .B(n2043), .Z(n2047) );
  NAND U2386 ( .A(n2045), .B(n2044), .Z(n2046) );
  NAND U2387 ( .A(n2047), .B(n2046), .Z(n2060) );
  AND U2388 ( .A(n2060), .B(n2198), .Z(n2057) );
  ANDN U2389 ( .B(n2048), .A(n2057), .Z(n2052) );
  ANDN U2390 ( .B(n2053), .A(n2052), .Z(n2049) );
  OR U2391 ( .A(n2049), .B(n2051), .Z(n2050) );
  AND U2392 ( .A(n2050), .B(n2227), .Z(n2072) );
  ANDN U2393 ( .B(n2071), .A(n2072), .Z(n2069) );
  NANDN U2394 ( .A(n2227), .B(n2051), .Z(n2056) );
  XNOR U2395 ( .A(n2053), .B(n2052), .Z(n2054) );
  NAND U2396 ( .A(n2227), .B(n2054), .Z(n2055) );
  AND U2397 ( .A(n2056), .B(n2055), .Z(n2089) );
  ANDN U2398 ( .B(n2089), .A(n794), .Z(n2081) );
  NOR U2399 ( .A(n[3]), .B(n2089), .Z(n2080) );
  NOR U2400 ( .A(n2117), .B(n2057), .Z(n2058) );
  XOR U2401 ( .A(n2059), .B(n2058), .Z(n2099) );
  NOR U2402 ( .A(n793), .B(n2099), .Z(n2078) );
  AND U2403 ( .A(n2198), .B(n2227), .Z(n2105) );
  XOR U2404 ( .A(n2105), .B(n2060), .Z(n2094) );
  ANDN U2405 ( .B(n[1]), .A(n2094), .Z(n2075) );
  NANDN U2406 ( .A(n[1]), .B(n2094), .Z(n2062) );
  NANDN U2407 ( .A(n[0]), .B(n2073), .Z(n2061) );
  NAND U2408 ( .A(n2062), .B(n2061), .Z(n2063) );
  NANDN U2409 ( .A(n2075), .B(n2063), .Z(n2064) );
  ANDN U2410 ( .B(n2099), .A(n[2]), .Z(n2077) );
  ANDN U2411 ( .B(n2064), .A(n2077), .Z(n2065) );
  OR U2412 ( .A(n2078), .B(n2065), .Z(n2066) );
  NANDN U2413 ( .A(n2080), .B(n2066), .Z(n2067) );
  NANDN U2414 ( .A(n2081), .B(n2067), .Z(n2068) );
  AND U2415 ( .A(n2069), .B(n2068), .Z(n2097) );
  NANDN U2416 ( .A(n2097), .B(n[0]), .Z(n2070) );
  XNOR U2417 ( .A(n2073), .B(n2070), .Z(n2102) );
  XNOR U2418 ( .A(n2072), .B(n2071), .Z(n2084) );
  ANDN U2419 ( .B(n[0]), .A(n2073), .Z(n2091) );
  XNOR U2420 ( .A(n[1]), .B(n2094), .Z(n2074) );
  NAND U2421 ( .A(n2091), .B(n2074), .Z(n2076) );
  ANDN U2422 ( .B(n2076), .A(n2075), .Z(n2095) );
  OR U2423 ( .A(n2077), .B(n2095), .Z(n2079) );
  ANDN U2424 ( .B(n2079), .A(n2078), .Z(n2086) );
  OR U2425 ( .A(n2080), .B(n2086), .Z(n2082) );
  ANDN U2426 ( .B(n2082), .A(n2081), .Z(n2083) );
  XNOR U2427 ( .A(n2084), .B(n2083), .Z(n2085) );
  ANDN U2428 ( .B(n2085), .A(n2097), .Z(n2153) );
  XNOR U2429 ( .A(n[3]), .B(n2086), .Z(n2087) );
  NANDN U2430 ( .A(n2097), .B(n2087), .Z(n2088) );
  XNOR U2431 ( .A(n2089), .B(n2088), .Z(n2127) );
  OR U2432 ( .A(n2127), .B(n[3]), .Z(n2090) );
  AND U2433 ( .A(n2129), .B(n2090), .Z(n2123) );
  AND U2434 ( .A(n2127), .B(n[3]), .Z(n2128) );
  XOR U2435 ( .A(n[1]), .B(n2091), .Z(n2092) );
  NANDN U2436 ( .A(n2097), .B(n2092), .Z(n2093) );
  XOR U2437 ( .A(n2094), .B(n2093), .Z(n2104) );
  XNOR U2438 ( .A(n[2]), .B(n2095), .Z(n2096) );
  NANDN U2439 ( .A(n2097), .B(n2096), .Z(n2098) );
  XNOR U2440 ( .A(n2099), .B(n2098), .Z(n2114) );
  NANDN U2441 ( .A(n2128), .B(n2124), .Z(n2100) );
  AND U2442 ( .A(n2123), .B(n2100), .Z(n2125) );
  NANDN U2443 ( .A(n2125), .B(n[0]), .Z(n2101) );
  XOR U2444 ( .A(n2102), .B(n2101), .Z(n2106) );
  XNOR U2445 ( .A(n2105), .B(n2118), .Z(n2115) );
  XOR U2446 ( .A(n2116), .B(n2115), .Z(n2173) );
  ANDN U2447 ( .B(n[2]), .A(n2173), .Z(n2144) );
  XNOR U2448 ( .A(n2107), .B(n2106), .Z(n2180) );
  NAND U2449 ( .A(n[1]), .B(n2180), .Z(n2141) );
  IV U2450 ( .A(n2180), .Z(n2137) );
  XNOR U2451 ( .A(n[1]), .B(n2137), .Z(n2108) );
  ANDN U2452 ( .B(n2198), .A(n2235), .Z(n2232) );
  IV U2453 ( .A(n2232), .Z(n2175) );
  AND U2454 ( .A(n[0]), .B(n2175), .Z(n2176) );
  NAND U2455 ( .A(n2108), .B(n2176), .Z(n2109) );
  AND U2456 ( .A(n2141), .B(n2109), .Z(n2170) );
  NANDN U2457 ( .A(n2144), .B(n2170), .Z(n2110) );
  AND U2458 ( .A(n2173), .B(n793), .Z(n2143) );
  ANDN U2459 ( .B(n2110), .A(n2143), .Z(n2164) );
  XOR U2460 ( .A(n2111), .B(n[2]), .Z(n2112) );
  NANDN U2461 ( .A(n2125), .B(n2112), .Z(n2113) );
  XNOR U2462 ( .A(n2114), .B(n2113), .Z(n2131) );
  IV U2463 ( .A(n2191), .Z(n2224) );
  NAND U2464 ( .A(n2116), .B(n2115), .Z(n2120) );
  OR U2465 ( .A(n2118), .B(n2117), .Z(n2119) );
  AND U2466 ( .A(n2120), .B(n2119), .Z(n2132) );
  XOR U2467 ( .A(n2224), .B(n2132), .Z(n2121) );
  NAND U2468 ( .A(n2198), .B(n2121), .Z(n2122) );
  XNOR U2469 ( .A(n2131), .B(n2122), .Z(n2167) );
  NOR U2470 ( .A(n2124), .B(n2123), .Z(n2147) );
  NANDN U2471 ( .A(n2125), .B(n[3]), .Z(n2126) );
  NANDN U2472 ( .A(n2127), .B(n2126), .Z(n2148) );
  NANDN U2473 ( .A(n2129), .B(n2128), .Z(n2130) );
  AND U2474 ( .A(n2148), .B(n2130), .Z(n2146) );
  XNOR U2475 ( .A(n2147), .B(n2146), .Z(n2151) );
  AND U2476 ( .A(n2131), .B(n2191), .Z(n2135) );
  XNOR U2477 ( .A(n2224), .B(n2131), .Z(n2133) );
  ANDN U2478 ( .B(n2133), .A(n2132), .Z(n2134) );
  OR U2479 ( .A(n2135), .B(n2134), .Z(n2136) );
  AND U2480 ( .A(n2136), .B(n2198), .Z(n2150) );
  XNOR U2481 ( .A(n2151), .B(n2150), .Z(n2161) );
  ANDN U2482 ( .B(n2137), .A(n[1]), .Z(n2139) );
  ANDN U2483 ( .B(n2232), .A(n[0]), .Z(n2138) );
  OR U2484 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U2485 ( .A(n2141), .B(n2140), .Z(n2142) );
  NANDN U2486 ( .A(n2143), .B(n2142), .Z(n2145) );
  ANDN U2487 ( .B(n2145), .A(n2144), .Z(n2157) );
  NAND U2488 ( .A(n794), .B(n2157), .Z(n2156) );
  NANDN U2489 ( .A(n2147), .B(n2146), .Z(n2149) );
  AND U2490 ( .A(n2149), .B(n2148), .Z(n2155) );
  AND U2491 ( .A(n2151), .B(n2150), .Z(n2152) );
  XNOR U2492 ( .A(n2153), .B(n2152), .Z(n2154) );
  XNOR U2493 ( .A(n2155), .B(n2154), .Z(n2163) );
  ANDN U2494 ( .B(n2156), .A(n2163), .Z(n2160) );
  XOR U2495 ( .A(n2157), .B(n794), .Z(n2158) );
  NAND U2496 ( .A(n2158), .B(n2167), .Z(n2159) );
  NAND U2497 ( .A(n2160), .B(n2159), .Z(n2162) );
  NANDN U2498 ( .A(n2162), .B(n2161), .Z(n2178) );
  ANDN U2499 ( .B(n2220), .A(n2163), .Z(n2169) );
  XOR U2500 ( .A(n[3]), .B(n2164), .Z(n2165) );
  NAND U2501 ( .A(n2178), .B(n2165), .Z(n2166) );
  XNOR U2502 ( .A(n2167), .B(n2166), .Z(n2213) );
  NANDN U2503 ( .A(n[3]), .B(n2213), .Z(n2168) );
  AND U2504 ( .A(n2169), .B(n2168), .Z(n2188) );
  XNOR U2505 ( .A(n[2]), .B(n2170), .Z(n2171) );
  NAND U2506 ( .A(n2178), .B(n2171), .Z(n2172) );
  XNOR U2507 ( .A(n2173), .B(n2172), .Z(n2189) );
  NANDN U2508 ( .A(n2189), .B(n[2]), .Z(n2187) );
  ANDN U2509 ( .B(n2189), .A(n[2]), .Z(n2181) );
  NAND U2510 ( .A(n2178), .B(n[0]), .Z(n2174) );
  XOR U2511 ( .A(n2175), .B(n2174), .Z(n2197) );
  XOR U2512 ( .A(n2176), .B(n[1]), .Z(n2177) );
  NAND U2513 ( .A(n2178), .B(n2177), .Z(n2179) );
  XNOR U2514 ( .A(n2180), .B(n2179), .Z(n2195) );
  OR U2515 ( .A(n2181), .B(n2186), .Z(n2182) );
  AND U2516 ( .A(n2187), .B(n2182), .Z(n2184) );
  NANDN U2517 ( .A(n2213), .B(n[3]), .Z(n2183) );
  NAND U2518 ( .A(n2184), .B(n2183), .Z(n2185) );
  NAND U2519 ( .A(n2188), .B(n2185), .Z(n2210) );
  ANDN U2520 ( .B(n2210), .A(n2186), .Z(n2207) );
  OR U2521 ( .A(n2188), .B(n2187), .Z(n2190) );
  ANDN U2522 ( .B(n2190), .A(n2209), .Z(n2206) );
  XNOR U2523 ( .A(n2207), .B(n2206), .Z(n2225) );
  AND U2524 ( .A(n2225), .B(n2191), .Z(n2204) );
  XNOR U2525 ( .A(n2224), .B(n2225), .Z(n2202) );
  XOR U2526 ( .A(n[1]), .B(n2192), .Z(n2193) );
  NAND U2527 ( .A(n2210), .B(n2193), .Z(n2194) );
  XNOR U2528 ( .A(n2195), .B(n2194), .Z(n2230) );
  NANDN U2529 ( .A(n2230), .B(n2227), .Z(n2201) );
  XNOR U2530 ( .A(n2230), .B(n2227), .Z(n2199) );
  NAND U2531 ( .A(n2210), .B(n[0]), .Z(n2196) );
  XNOR U2532 ( .A(n2197), .B(n2196), .Z(n2231) );
  AND U2533 ( .A(n2231), .B(n2198), .Z(n2226) );
  NAND U2534 ( .A(n2199), .B(n2226), .Z(n2200) );
  NAND U2535 ( .A(n2201), .B(n2200), .Z(n2223) );
  AND U2536 ( .A(n2202), .B(n2223), .Z(n2203) );
  OR U2537 ( .A(n2204), .B(n2203), .Z(n2205) );
  ANDN U2538 ( .B(n2205), .A(n2235), .Z(n2217) );
  NANDN U2539 ( .A(n2207), .B(n2206), .Z(n2208) );
  NANDN U2540 ( .A(n2209), .B(n2208), .Z(n2212) );
  ANDN U2541 ( .B(n2210), .A(n794), .Z(n2214) );
  XNOR U2542 ( .A(n2213), .B(n2214), .Z(n2211) );
  XNOR U2543 ( .A(n2217), .B(n2218), .Z(n2243) );
  NAND U2544 ( .A(n2212), .B(n2211), .Z(n2216) );
  NANDN U2545 ( .A(n2214), .B(n2213), .Z(n2215) );
  AND U2546 ( .A(n2216), .B(n2215), .Z(n2222) );
  AND U2547 ( .A(n2218), .B(n2217), .Z(n2219) );
  XNOR U2548 ( .A(n2220), .B(n2219), .Z(n2221) );
  XNOR U2549 ( .A(n2222), .B(n2221), .Z(n2245) );
  NOR U2550 ( .A(n[3]), .B(n2264), .Z(n2241) );
  XOR U2551 ( .A(n2227), .B(n2226), .Z(n2228) );
  NANDN U2552 ( .A(n2235), .B(n2228), .Z(n2229) );
  XNOR U2553 ( .A(n2230), .B(n2229), .Z(n2256) );
  AND U2554 ( .A(n2264), .B(n[3]), .Z(n2239) );
  XOR U2555 ( .A(n2232), .B(n2231), .Z(n2249) );
  NAND U2556 ( .A(n2262), .B(n[0]), .Z(n2234) );
  XNOR U2557 ( .A(n2235), .B(n2234), .Z(n2266) );
  NANDN U2558 ( .A(n2249), .B(n[1]), .Z(n2238) );
  XNOR U2559 ( .A(n[1]), .B(n2249), .Z(n2236) );
  AND U2560 ( .A(n[0]), .B(n2235), .Z(n2246) );
  NAND U2561 ( .A(n2236), .B(n2246), .Z(n2237) );
  AND U2562 ( .A(n2238), .B(n2237), .Z(n2253) );
  NANDN U2563 ( .A(n2239), .B(n2260), .Z(n2240) );
  NANDN U2564 ( .A(n2241), .B(n2240), .Z(n2242) );
  NANDN U2565 ( .A(n2243), .B(n2242), .Z(n2244) );
  NAND U2566 ( .A(n2245), .B(n2244), .Z(n2269) );
  AND U2567 ( .A(n[0]), .B(n2266), .Z(n2366) );
  NAND U2568 ( .A(n[1]), .B(n2366), .Z(n2252) );
  XOR U2569 ( .A(n[1]), .B(n2246), .Z(n2247) );
  NAND U2570 ( .A(n2262), .B(n2247), .Z(n2248) );
  XOR U2571 ( .A(n2249), .B(n2248), .Z(n2370) );
  NANDN U2572 ( .A(n2366), .B(n792), .Z(n2250) );
  NAND U2573 ( .A(n2370), .B(n2250), .Z(n2251) );
  AND U2574 ( .A(n2252), .B(n2251), .Z(n2293) );
  XNOR U2575 ( .A(n[2]), .B(n2253), .Z(n2254) );
  NAND U2576 ( .A(n2262), .B(n2254), .Z(n2255) );
  XNOR U2577 ( .A(n2256), .B(n2255), .Z(n2296) );
  XOR U2578 ( .A(n[2]), .B(n2296), .Z(n2257) );
  NANDN U2579 ( .A(n2293), .B(n2257), .Z(n2259) );
  NAND U2580 ( .A(n[2]), .B(n2296), .Z(n2258) );
  AND U2581 ( .A(n2259), .B(n2258), .Z(n2268) );
  XNOR U2582 ( .A(n[3]), .B(n2260), .Z(n2261) );
  NAND U2583 ( .A(n2262), .B(n2261), .Z(n2263) );
  XNOR U2584 ( .A(n2264), .B(n2263), .Z(n2270) );
  NAND U2585 ( .A(n2368), .B(n[0]), .Z(n2265) );
  XNOR U2586 ( .A(n2266), .B(n2265), .Z(n2267) );
  OR U2587 ( .A(e[0]), .B(n2267), .Z(n2527) );
  IV U2588 ( .A(n2267), .Z(n2494) );
  AND U2589 ( .A(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .B(n2494), .Z(n2497) );
  ANDN U2590 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n2552), .Z(n2292) );
  ANDN U2591 ( .B(n[0]), .A(n2292), .Z(n2279) );
  ANDN U2592 ( .B(\cin[1][1] ), .A(n2552), .Z(n2282) );
  NAND U2593 ( .A(n2286), .B(n2271), .Z(n2272) );
  ANDN U2594 ( .B(n2272), .A(n2552), .Z(n2273) );
  AND U2595 ( .A(n2274), .B(n2273), .Z(n2322) );
  ANDN U2596 ( .B(n2275), .A(n2552), .Z(n2287) );
  NAND U2597 ( .A(n2276), .B(n2287), .Z(n2278) );
  OR U2598 ( .A(n2287), .B(n2292), .Z(n2277) );
  NAND U2599 ( .A(n2278), .B(n2277), .Z(n2291) );
  NAND U2600 ( .A(n[0]), .B(n2291), .Z(n2298) );
  NANDN U2601 ( .A(n[1]), .B(n2298), .Z(n2285) );
  NOR U2602 ( .A(n792), .B(n2298), .Z(n2283) );
  XOR U2603 ( .A(n[1]), .B(n2279), .Z(n2280) );
  NAND U2604 ( .A(n2287), .B(n2280), .Z(n2281) );
  XNOR U2605 ( .A(n2282), .B(n2281), .Z(n2301) );
  NANDN U2606 ( .A(n2283), .B(n2301), .Z(n2284) );
  AND U2607 ( .A(n2285), .B(n2284), .Z(n2312) );
  NANDN U2608 ( .A(n2552), .B(n2288), .Z(n2323) );
  NANDN U2609 ( .A(n794), .B(n2323), .Z(n2289) );
  NAND U2610 ( .A(n2324), .B(n2289), .Z(n2290) );
  NANDN U2611 ( .A(n2322), .B(n2290), .Z(n2314) );
  XNOR U2612 ( .A(n[2]), .B(n2293), .Z(n2294) );
  NAND U2613 ( .A(n2368), .B(n2294), .Z(n2295) );
  XNOR U2614 ( .A(n2296), .B(n2295), .Z(n2536) );
  ANDN U2615 ( .B(\cin[1][1] ), .A(n2536), .Z(n2297) );
  XOR U2616 ( .A(n2302), .B(n2297), .Z(n2342) );
  XOR U2617 ( .A(n792), .B(n2298), .Z(n2299) );
  NAND U2618 ( .A(n2314), .B(n2299), .Z(n2300) );
  XNOR U2619 ( .A(n2301), .B(n2300), .Z(n2317) );
  AND U2620 ( .A(\cin[1][1] ), .B(n2302), .Z(n2318) );
  XOR U2621 ( .A(\cin[1][2] ), .B(n2318), .Z(n2303) );
  ANDN U2622 ( .B(n2303), .A(n2536), .Z(n2304) );
  XNOR U2623 ( .A(n2317), .B(n2304), .Z(n2350) );
  XOR U2624 ( .A(n[2]), .B(n2350), .Z(n2309) );
  OR U2625 ( .A(n2342), .B(n792), .Z(n2346) );
  NANDN U2626 ( .A(n2536), .B(n2488), .Z(n2306) );
  NANDN U2627 ( .A(n[1]), .B(n2342), .Z(n2305) );
  NAND U2628 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U2629 ( .A(n2346), .B(n2307), .Z(n2308) );
  NAND U2630 ( .A(n2309), .B(n2308), .Z(n2311) );
  NAND U2631 ( .A(n[2]), .B(n2350), .Z(n2310) );
  AND U2632 ( .A(n2311), .B(n2310), .Z(n2329) );
  NAND U2633 ( .A(n794), .B(n2329), .Z(n2328) );
  XOR U2634 ( .A(n[2]), .B(n2312), .Z(n2313) );
  NAND U2635 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U2636 ( .A(n2316), .B(n2315), .Z(n2333) );
  NAND U2637 ( .A(\cin[1][2] ), .B(n2317), .Z(n2321) );
  XOR U2638 ( .A(\cin[1][2] ), .B(n2317), .Z(n2319) );
  NAND U2639 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2640 ( .A(n2321), .B(n2320), .Z(n2330) );
  XNOR U2641 ( .A(n2322), .B(n2324), .Z(n2326) );
  NANDN U2642 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U2643 ( .A(n2326), .B(n2325), .Z(n2356) );
  NANDN U2644 ( .A(n2357), .B(n2356), .Z(n2327) );
  ANDN U2645 ( .B(n2328), .A(n2327), .Z(n2336) );
  XOR U2646 ( .A(n794), .B(n2329), .Z(n2334) );
  XNOR U2647 ( .A(\cin[1][3] ), .B(n2330), .Z(n2331) );
  NANDN U2648 ( .A(n2536), .B(n2331), .Z(n2332) );
  XNOR U2649 ( .A(n2333), .B(n2332), .Z(n2355) );
  NAND U2650 ( .A(n2334), .B(n2355), .Z(n2335) );
  NAND U2651 ( .A(n2336), .B(n2335), .Z(n2352) );
  NANDN U2652 ( .A(n2536), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n2337)
         );
  AND U2653 ( .A(n[0]), .B(n2337), .Z(n2343) );
  XOR U2654 ( .A(n[1]), .B(n2343), .Z(n2338) );
  NAND U2655 ( .A(n2352), .B(n2338), .Z(n2339) );
  XNOR U2656 ( .A(n2342), .B(n2339), .Z(n2365) );
  IV U2657 ( .A(n2352), .Z(n2358) );
  ANDN U2658 ( .B(n[0]), .A(n2358), .Z(n2341) );
  ANDN U2659 ( .B(\MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), 
        .A(n2536), .Z(n2340) );
  XOR U2660 ( .A(n2341), .B(n2340), .Z(n2372) );
  ANDN U2661 ( .B(n[0]), .A(n2372), .Z(n2362) );
  XNOR U2662 ( .A(n[1]), .B(n2342), .Z(n2344) );
  NAND U2663 ( .A(n2344), .B(n2343), .Z(n2345) );
  AND U2664 ( .A(n2346), .B(n2345), .Z(n2349) );
  XNOR U2665 ( .A(n[2]), .B(n2349), .Z(n2347) );
  NAND U2666 ( .A(n2352), .B(n2347), .Z(n2348) );
  XNOR U2667 ( .A(n2350), .B(n2348), .Z(n2378) );
  XNOR U2668 ( .A(n[3]), .B(n2354), .Z(n2351) );
  NAND U2669 ( .A(n2352), .B(n2351), .Z(n2353) );
  XNOR U2670 ( .A(n2355), .B(n2353), .Z(n2392) );
  ANDN U2671 ( .B(n[3]), .A(n2392), .Z(n2388) );
  OR U2672 ( .A(n2395), .B(n2388), .Z(n2361) );
  NANDN U2673 ( .A(n2356), .B(n2357), .Z(n2359) );
  AND U2674 ( .A(n2359), .B(n2403), .Z(n2389) );
  NANDN U2675 ( .A(n[3]), .B(n2392), .Z(n2360) );
  NAND U2676 ( .A(n2389), .B(n2360), .Z(n2394) );
  ANDN U2677 ( .B(n2361), .A(n2394), .Z(n2390) );
  XOR U2678 ( .A(n2362), .B(n[1]), .Z(n2363) );
  NANDN U2679 ( .A(n2390), .B(n2363), .Z(n2364) );
  XNOR U2680 ( .A(n2365), .B(n2364), .Z(n2379) );
  XOR U2681 ( .A(n[1]), .B(n2366), .Z(n2367) );
  NAND U2682 ( .A(n2368), .B(n2367), .Z(n2369) );
  XNOR U2683 ( .A(n2370), .B(n2369), .Z(n2528) );
  NANDN U2684 ( .A(n2390), .B(n[0]), .Z(n2371) );
  XNOR U2685 ( .A(n2372), .B(n2371), .Z(n2411) );
  AND U2686 ( .A(\cin[1][1] ), .B(n2411), .Z(n2380) );
  XOR U2687 ( .A(n2380), .B(\cin[1][2] ), .Z(n2373) );
  NANDN U2688 ( .A(n2528), .B(n2373), .Z(n2374) );
  XNOR U2689 ( .A(n2379), .B(n2374), .Z(n2426) );
  XOR U2690 ( .A(n2375), .B(n[2]), .Z(n2376) );
  NANDN U2691 ( .A(n2390), .B(n2376), .Z(n2377) );
  XNOR U2692 ( .A(n2378), .B(n2377), .Z(n2409) );
  ANDN U2693 ( .B(\cin[1][3] ), .A(n2409), .Z(n2386) );
  XNOR U2694 ( .A(\cin[1][3] ), .B(n2409), .Z(n2384) );
  NAND U2695 ( .A(\cin[1][2] ), .B(n2379), .Z(n2383) );
  XOR U2696 ( .A(\cin[1][2] ), .B(n2379), .Z(n2381) );
  NAND U2697 ( .A(n2381), .B(n2380), .Z(n2382) );
  NAND U2698 ( .A(n2383), .B(n2382), .Z(n2406) );
  AND U2699 ( .A(n2384), .B(n2406), .Z(n2385) );
  OR U2700 ( .A(n2386), .B(n2385), .Z(n2387) );
  ANDN U2701 ( .B(n2387), .A(n2528), .Z(n2400) );
  NANDN U2702 ( .A(n2389), .B(n2388), .Z(n2393) );
  NANDN U2703 ( .A(n2390), .B(n[3]), .Z(n2391) );
  AND U2704 ( .A(n2392), .B(n2391), .Z(n2399) );
  ANDN U2705 ( .B(n2393), .A(n2399), .Z(n2397) );
  NAND U2706 ( .A(n2395), .B(n2394), .Z(n2396) );
  XOR U2707 ( .A(n2397), .B(n2396), .Z(n2401) );
  XOR U2708 ( .A(n2400), .B(n2401), .Z(n2435) );
  AND U2709 ( .A(n2397), .B(n2396), .Z(n2398) );
  NOR U2710 ( .A(n2399), .B(n2398), .Z(n2405) );
  AND U2711 ( .A(n2401), .B(n2400), .Z(n2402) );
  XOR U2712 ( .A(n2403), .B(n2402), .Z(n2404) );
  XNOR U2713 ( .A(n2405), .B(n2404), .Z(n2437) );
  NOR U2714 ( .A(n2435), .B(n2437), .Z(n2419) );
  XOR U2715 ( .A(n2406), .B(\cin[1][3] ), .Z(n2407) );
  NANDN U2716 ( .A(n2528), .B(n2407), .Z(n2408) );
  XNOR U2717 ( .A(n2409), .B(n2408), .Z(n2441) );
  NAND U2718 ( .A(n[3]), .B(n2441), .Z(n2433) );
  ANDN U2719 ( .B(n[2]), .A(n2426), .Z(n2428) );
  ANDN U2720 ( .B(n2433), .A(n2428), .Z(n2417) );
  NANDN U2721 ( .A(n2528), .B(\cin[1][1] ), .Z(n2410) );
  XNOR U2722 ( .A(n2411), .B(n2410), .Z(n2449) );
  ANDN U2723 ( .B(n2449), .A(n[1]), .Z(n2413) );
  NANDN U2724 ( .A(n2528), .B(n2488), .Z(n2412) );
  NANDN U2725 ( .A(n2413), .B(n2412), .Z(n2414) );
  AND U2726 ( .A(n2423), .B(n2414), .Z(n2415) );
  ANDN U2727 ( .B(n2426), .A(n[2]), .Z(n2429) );
  OR U2728 ( .A(n2415), .B(n2429), .Z(n2416) );
  AND U2729 ( .A(n2417), .B(n2416), .Z(n2418) );
  ANDN U2730 ( .B(n2419), .A(n2418), .Z(n2420) );
  NOR U2731 ( .A(n[3]), .B(n2441), .Z(n2431) );
  ANDN U2732 ( .B(n2420), .A(n2431), .Z(n2447) );
  XNOR U2733 ( .A(n[1]), .B(n2449), .Z(n2421) );
  NANDN U2734 ( .A(n2528), .B(
        \MODMULT2[3].modmult_2/MODMULT_STEP[1].modmult_step_/N4 ), .Z(n2444)
         );
  AND U2735 ( .A(n[0]), .B(n2444), .Z(n2445) );
  NAND U2736 ( .A(n2421), .B(n2445), .Z(n2422) );
  NAND U2737 ( .A(n2423), .B(n2422), .Z(n2427) );
  XNOR U2738 ( .A(n793), .B(n2427), .Z(n2424) );
  NANDN U2739 ( .A(n2447), .B(n2424), .Z(n2425) );
  XNOR U2740 ( .A(n2426), .B(n2425), .Z(n2454) );
  OR U2741 ( .A(n2428), .B(n2427), .Z(n2430) );
  ANDN U2742 ( .B(n2430), .A(n2429), .Z(n2438) );
  NANDN U2743 ( .A(n2431), .B(n2438), .Z(n2432) );
  AND U2744 ( .A(n2433), .B(n2432), .Z(n2434) );
  XNOR U2745 ( .A(n2435), .B(n2434), .Z(n2436) );
  ANDN U2746 ( .B(n2436), .A(n2447), .Z(n2483) );
  NOR U2747 ( .A(n2483), .B(n2437), .Z(n2469) );
  XOR U2748 ( .A(n[3]), .B(n2438), .Z(n2439) );
  NANDN U2749 ( .A(n2447), .B(n2439), .Z(n2440) );
  XNOR U2750 ( .A(n2441), .B(n2440), .Z(n2472) );
  OR U2751 ( .A(n2472), .B(n[3]), .Z(n2442) );
  AND U2752 ( .A(n2469), .B(n2442), .Z(n2475) );
  NANDN U2753 ( .A(n2447), .B(n[0]), .Z(n2443) );
  XOR U2754 ( .A(n2444), .B(n2443), .Z(n2460) );
  ANDN U2755 ( .B(n[0]), .A(n2460), .Z(n2455) );
  XOR U2756 ( .A(n2445), .B(n[1]), .Z(n2446) );
  NANDN U2757 ( .A(n2447), .B(n2446), .Z(n2448) );
  XNOR U2758 ( .A(n2449), .B(n2448), .Z(n2458) );
  AND U2759 ( .A(n2472), .B(n[3]), .Z(n2468) );
  OR U2760 ( .A(n2474), .B(n2468), .Z(n2450) );
  AND U2761 ( .A(n2475), .B(n2450), .Z(n2470) );
  XNOR U2762 ( .A(n2451), .B(n[2]), .Z(n2452) );
  NANDN U2763 ( .A(n2470), .B(n2452), .Z(n2453) );
  XNOR U2764 ( .A(n2454), .B(n2453), .Z(n2495) );
  AND U2765 ( .A(\cin[1][3] ), .B(n2495), .Z(n2466) );
  XOR U2766 ( .A(\cin[1][3] ), .B(n2495), .Z(n2464) );
  XOR U2767 ( .A(n2455), .B(n[1]), .Z(n2456) );
  NANDN U2768 ( .A(n2470), .B(n2456), .Z(n2457) );
  XNOR U2769 ( .A(n2458), .B(n2457), .Z(n2492) );
  NAND U2770 ( .A(\cin[1][2] ), .B(n2492), .Z(n2463) );
  XOR U2771 ( .A(\cin[1][2] ), .B(n2492), .Z(n2461) );
  NANDN U2772 ( .A(n2470), .B(n[0]), .Z(n2459) );
  XNOR U2773 ( .A(n2460), .B(n2459), .Z(n2487) );
  AND U2774 ( .A(\cin[1][1] ), .B(n2487), .Z(n2489) );
  NAND U2775 ( .A(n2461), .B(n2489), .Z(n2462) );
  NAND U2776 ( .A(n2463), .B(n2462), .Z(n2493) );
  AND U2777 ( .A(n2464), .B(n2493), .Z(n2465) );
  OR U2778 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2779 ( .A(n2467), .B(n2494), .Z(n2480) );
  NANDN U2780 ( .A(n2469), .B(n2468), .Z(n2473) );
  NANDN U2781 ( .A(n2470), .B(n[3]), .Z(n2471) );
  NANDN U2782 ( .A(n2472), .B(n2471), .Z(n2478) );
  AND U2783 ( .A(n2473), .B(n2478), .Z(n2477) );
  NANDN U2784 ( .A(n2475), .B(n2474), .Z(n2476) );
  XOR U2785 ( .A(n2477), .B(n2476), .Z(n2481) );
  XNOR U2786 ( .A(n2480), .B(n2481), .Z(n2504) );
  NAND U2787 ( .A(n2477), .B(n2476), .Z(n2479) );
  AND U2788 ( .A(n2479), .B(n2478), .Z(n2485) );
  AND U2789 ( .A(n2481), .B(n2480), .Z(n2482) );
  XNOR U2790 ( .A(n2483), .B(n2482), .Z(n2484) );
  XNOR U2791 ( .A(n2485), .B(n2484), .Z(n2509) );
  NAND U2792 ( .A(n2494), .B(\cin[1][1] ), .Z(n2486) );
  XNOR U2793 ( .A(n2487), .B(n2486), .Z(n2517) );
  XOR U2794 ( .A(\cin[1][2] ), .B(n2489), .Z(n2490) );
  NAND U2795 ( .A(n2494), .B(n2490), .Z(n2491) );
  XNOR U2796 ( .A(n2492), .B(n2491), .Z(n2522) );
  ANDN U2797 ( .B(n[3]), .A(n2513), .Z(n2501) );
  ANDN U2798 ( .B(n2513), .A(n[3]), .Z(n2502) );
  NANDN U2799 ( .A(n2520), .B(n[0]), .Z(n2496) );
  XNOR U2800 ( .A(n2497), .B(n2496), .Z(n2524) );
  XNOR U2801 ( .A(n[1]), .B(n2517), .Z(n2498) );
  ANDN U2802 ( .B(n[0]), .A(n2497), .Z(n2514) );
  NAND U2803 ( .A(n2498), .B(n2514), .Z(n2499) );
  AND U2804 ( .A(n2500), .B(n2499), .Z(n2518) );
  NANDN U2805 ( .A(n2501), .B(n2510), .Z(n2503) );
  ANDN U2806 ( .B(n2503), .A(n2502), .Z(n2505) );
  XNOR U2807 ( .A(n2505), .B(n2504), .Z(n2507) );
  NAND U2808 ( .A(n2505), .B(n2520), .Z(n2506) );
  NAND U2809 ( .A(n2507), .B(n2506), .Z(n2508) );
  NANDN U2810 ( .A(n2509), .B(n2508), .Z(n2548) );
  XNOR U2811 ( .A(n[3]), .B(n2510), .Z(n2511) );
  NANDN U2812 ( .A(n2520), .B(n2511), .Z(n2512) );
  XNOR U2813 ( .A(n2513), .B(n2512), .Z(n2546) );
  XOR U2814 ( .A(n[1]), .B(n2514), .Z(n2515) );
  NANDN U2815 ( .A(n2520), .B(n2515), .Z(n2516) );
  XNOR U2816 ( .A(n2517), .B(n2516), .Z(n2532) );
  XNOR U2817 ( .A(n[2]), .B(n2518), .Z(n2519) );
  NANDN U2818 ( .A(n2520), .B(n2519), .Z(n2521) );
  XNOR U2819 ( .A(n2522), .B(n2521), .Z(n2541) );
  AND U2820 ( .A(n[0]), .B(n2539), .Z(n2523) );
  XOR U2821 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U2822 ( .A(e[0]), .B(n2525), .Z(n2526) );
  NAND U2823 ( .A(n2527), .B(n2526), .Z(c[0]) );
  OR U2824 ( .A(n2528), .B(e[0]), .Z(n2535) );
  XOR U2825 ( .A(n2529), .B(n[1]), .Z(n2530) );
  AND U2826 ( .A(n2539), .B(n2530), .Z(n2531) );
  XOR U2827 ( .A(n2532), .B(n2531), .Z(n2533) );
  NAND U2828 ( .A(e[0]), .B(n2533), .Z(n2534) );
  NAND U2829 ( .A(n2535), .B(n2534), .Z(c[1]) );
  OR U2830 ( .A(n2536), .B(e[0]), .Z(n2544) );
  XOR U2831 ( .A(n2537), .B(n[2]), .Z(n2538) );
  AND U2832 ( .A(n2539), .B(n2538), .Z(n2540) );
  XOR U2833 ( .A(n2541), .B(n2540), .Z(n2542) );
  NAND U2834 ( .A(e[0]), .B(n2542), .Z(n2543) );
  NAND U2835 ( .A(n2544), .B(n2543), .Z(c[2]) );
  XNOR U2836 ( .A(n[3]), .B(n2545), .Z(n2547) );
  XOR U2837 ( .A(n2546), .B(n2547), .Z(n2550) );
  NANDN U2838 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U2839 ( .A(n2550), .B(n2549), .Z(n2551) );
  NANDN U2840 ( .A(n2551), .B(e[0]), .Z(n2554) );
  OR U2841 ( .A(e[0]), .B(n2552), .Z(n2553) );
  NAND U2842 ( .A(n2554), .B(n2553), .Z(c[3]) );
endmodule

