
module hamming_N1600_CC4 ( clk, rst, x, y, o );
  input [399:0] x;
  input [399:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  OR U403 ( .A(n886), .B(n887), .Z(n1) );
  NANDN U404 ( .A(n889), .B(n888), .Z(n2) );
  NAND U405 ( .A(n1), .B(n2), .Z(n1857) );
  OR U406 ( .A(n469), .B(n470), .Z(n3) );
  NANDN U407 ( .A(n472), .B(n471), .Z(n4) );
  NAND U408 ( .A(n3), .B(n4), .Z(n1456) );
  OR U409 ( .A(n1322), .B(n1323), .Z(n5) );
  NANDN U410 ( .A(n1325), .B(n1324), .Z(n6) );
  AND U411 ( .A(n5), .B(n6), .Z(n1726) );
  NANDN U412 ( .A(n989), .B(n988), .Z(n7) );
  NANDN U413 ( .A(n986), .B(n987), .Z(n8) );
  AND U414 ( .A(n7), .B(n8), .Z(n1609) );
  OR U415 ( .A(n678), .B(n679), .Z(n9) );
  NANDN U416 ( .A(n681), .B(n680), .Z(n10) );
  NAND U417 ( .A(n9), .B(n10), .Z(n1597) );
  OR U418 ( .A(n1732), .B(n1733), .Z(n11) );
  NANDN U419 ( .A(n1735), .B(n1734), .Z(n12) );
  NAND U420 ( .A(n11), .B(n12), .Z(n2065) );
  OR U421 ( .A(n1618), .B(n1619), .Z(n13) );
  OR U422 ( .A(n1616), .B(n1617), .Z(n14) );
  AND U423 ( .A(n13), .B(n14), .Z(n2130) );
  OR U424 ( .A(n1600), .B(n1601), .Z(n15) );
  NANDN U425 ( .A(n1603), .B(n1602), .Z(n16) );
  NAND U426 ( .A(n15), .B(n16), .Z(n2071) );
  OR U427 ( .A(n2216), .B(n2217), .Z(n17) );
  NAND U428 ( .A(n2219), .B(n2218), .Z(n18) );
  NAND U429 ( .A(n17), .B(n18), .Z(n2337) );
  OR U430 ( .A(n2164), .B(n2165), .Z(n19) );
  NANDN U431 ( .A(n2166), .B(n2167), .Z(n20) );
  NAND U432 ( .A(n19), .B(n20), .Z(n2318) );
  OR U433 ( .A(n2244), .B(n2245), .Z(n21) );
  NANDN U434 ( .A(n2243), .B(n2242), .Z(n22) );
  NAND U435 ( .A(n21), .B(n22), .Z(n2300) );
  OR U436 ( .A(n942), .B(n943), .Z(n23) );
  NANDN U437 ( .A(n945), .B(n944), .Z(n24) );
  AND U438 ( .A(n23), .B(n24), .Z(n1580) );
  OR U439 ( .A(n808), .B(n809), .Z(n25) );
  NANDN U440 ( .A(n811), .B(n810), .Z(n26) );
  NAND U441 ( .A(n25), .B(n26), .Z(n1741) );
  OR U442 ( .A(n531), .B(n532), .Z(n27) );
  NANDN U443 ( .A(n534), .B(n533), .Z(n28) );
  NAND U444 ( .A(n27), .B(n28), .Z(n1402) );
  OR U445 ( .A(n882), .B(n883), .Z(n29) );
  NANDN U446 ( .A(n885), .B(n884), .Z(n30) );
  NAND U447 ( .A(n29), .B(n30), .Z(n1858) );
  OR U448 ( .A(n473), .B(n474), .Z(n31) );
  NANDN U449 ( .A(n476), .B(n475), .Z(n32) );
  NAND U450 ( .A(n31), .B(n32), .Z(n1458) );
  OR U451 ( .A(n1318), .B(n1319), .Z(n33) );
  NANDN U452 ( .A(n1321), .B(n1320), .Z(n34) );
  NAND U453 ( .A(n33), .B(n34), .Z(n1727) );
  OR U454 ( .A(n564), .B(n565), .Z(n35) );
  NANDN U455 ( .A(n567), .B(n566), .Z(n36) );
  AND U456 ( .A(n35), .B(n36), .Z(n1789) );
  OR U457 ( .A(n550), .B(n551), .Z(n37) );
  NANDN U458 ( .A(n553), .B(n552), .Z(n38) );
  AND U459 ( .A(n37), .B(n38), .Z(n1769) );
  OR U460 ( .A(n439), .B(n440), .Z(n39) );
  NANDN U461 ( .A(n442), .B(n441), .Z(n40) );
  NAND U462 ( .A(n39), .B(n40), .Z(n1476) );
  OR U463 ( .A(n682), .B(n683), .Z(n41) );
  NANDN U464 ( .A(n685), .B(n684), .Z(n42) );
  NAND U465 ( .A(n41), .B(n42), .Z(n1596) );
  OR U466 ( .A(n1407), .B(n1406), .Z(n43) );
  NAND U467 ( .A(n1408), .B(n1409), .Z(n44) );
  AND U468 ( .A(n43), .B(n44), .Z(n1999) );
  OR U469 ( .A(n1854), .B(n1853), .Z(n45) );
  NAND U470 ( .A(n1855), .B(n1856), .Z(n46) );
  AND U471 ( .A(n45), .B(n46), .Z(n1946) );
  OR U472 ( .A(n1460), .B(n1461), .Z(n47) );
  NANDN U473 ( .A(n1462), .B(n1463), .Z(n48) );
  AND U474 ( .A(n47), .B(n48), .Z(n1940) );
  OR U475 ( .A(n1472), .B(n1473), .Z(n49) );
  NANDN U476 ( .A(n1474), .B(n1475), .Z(n50) );
  AND U477 ( .A(n49), .B(n50), .Z(n1936) );
  OR U478 ( .A(n1736), .B(n1737), .Z(n51) );
  NANDN U479 ( .A(n1739), .B(n1738), .Z(n52) );
  AND U480 ( .A(n51), .B(n52), .Z(n2066) );
  OR U481 ( .A(n1785), .B(n1786), .Z(n53) );
  NANDN U482 ( .A(n1788), .B(n1787), .Z(n54) );
  NAND U483 ( .A(n53), .B(n54), .Z(n2059) );
  OR U484 ( .A(n1765), .B(n1766), .Z(n55) );
  NANDN U485 ( .A(n1768), .B(n1767), .Z(n56) );
  NAND U486 ( .A(n55), .B(n56), .Z(n2053) );
  XOR U487 ( .A(n2006), .B(n2007), .Z(n1982) );
  OR U488 ( .A(n1604), .B(n1605), .Z(n57) );
  NANDN U489 ( .A(n1607), .B(n1606), .Z(n58) );
  AND U490 ( .A(n57), .B(n58), .Z(n2072) );
  OR U491 ( .A(n2129), .B(n2130), .Z(n59) );
  NANDN U492 ( .A(n2131), .B(n2132), .Z(n60) );
  NAND U493 ( .A(n59), .B(n60), .Z(n2209) );
  OR U494 ( .A(n1909), .B(n1910), .Z(n61) );
  NANDN U495 ( .A(n1912), .B(n1911), .Z(n62) );
  AND U496 ( .A(n61), .B(n62), .Z(n2198) );
  OR U497 ( .A(n2030), .B(n2031), .Z(n63) );
  NANDN U498 ( .A(n2032), .B(n2033), .Z(n64) );
  AND U499 ( .A(n63), .B(n64), .Z(n2233) );
  OR U500 ( .A(n2314), .B(n2313), .Z(n65) );
  NAND U501 ( .A(n2315), .B(n2316), .Z(n66) );
  AND U502 ( .A(n65), .B(n66), .Z(n2352) );
  OR U503 ( .A(n2362), .B(n2363), .Z(n67) );
  OR U504 ( .A(n2360), .B(n2361), .Z(n68) );
  AND U505 ( .A(n67), .B(n68), .Z(n2375) );
  OR U506 ( .A(n2356), .B(n2357), .Z(n69) );
  NAND U507 ( .A(n2359), .B(n2358), .Z(n70) );
  NAND U508 ( .A(n69), .B(n70), .Z(n2385) );
  OR U509 ( .A(n1298), .B(n1299), .Z(n71) );
  NANDN U510 ( .A(n1301), .B(n1300), .Z(n72) );
  NAND U511 ( .A(n71), .B(n72), .Z(n1565) );
  OR U512 ( .A(n453), .B(n454), .Z(n73) );
  NANDN U513 ( .A(n456), .B(n455), .Z(n74) );
  NAND U514 ( .A(n73), .B(n74), .Z(n1422) );
  OR U515 ( .A(n670), .B(n671), .Z(n75) );
  NANDN U516 ( .A(n673), .B(n672), .Z(n76) );
  AND U517 ( .A(n75), .B(n76), .Z(n1534) );
  OR U518 ( .A(n946), .B(n947), .Z(n77) );
  NANDN U519 ( .A(n949), .B(n948), .Z(n78) );
  NAND U520 ( .A(n77), .B(n78), .Z(n1583) );
  OR U521 ( .A(n578), .B(n579), .Z(n79) );
  NANDN U522 ( .A(n581), .B(n580), .Z(n80) );
  AND U523 ( .A(n79), .B(n80), .Z(n1835) );
  OR U524 ( .A(n924), .B(n925), .Z(n81) );
  NANDN U525 ( .A(n927), .B(n926), .Z(n82) );
  NAND U526 ( .A(n81), .B(n82), .Z(n1751) );
  OR U527 ( .A(n828), .B(n829), .Z(n83) );
  NANDN U528 ( .A(n831), .B(n830), .Z(n84) );
  NAND U529 ( .A(n83), .B(n84), .Z(n1407) );
  OR U530 ( .A(n481), .B(n482), .Z(n85) );
  NANDN U531 ( .A(n484), .B(n483), .Z(n86) );
  NAND U532 ( .A(n85), .B(n86), .Z(n1460) );
  OR U533 ( .A(n708), .B(n709), .Z(n87) );
  NANDN U534 ( .A(n711), .B(n710), .Z(n88) );
  NAND U535 ( .A(n87), .B(n88), .Z(n1733) );
  OR U536 ( .A(n738), .B(n739), .Z(n89) );
  NANDN U537 ( .A(n741), .B(n740), .Z(n90) );
  NAND U538 ( .A(n89), .B(n90), .Z(n1766) );
  OR U539 ( .A(n435), .B(n436), .Z(n91) );
  NANDN U540 ( .A(n438), .B(n437), .Z(n92) );
  NAND U541 ( .A(n91), .B(n92), .Z(n1477) );
  OR U542 ( .A(n982), .B(n983), .Z(n93) );
  NANDN U543 ( .A(n985), .B(n984), .Z(n94) );
  AND U544 ( .A(n93), .B(n94), .Z(n1608) );
  NANDN U545 ( .A(n1095), .B(n1094), .Z(n95) );
  NANDN U546 ( .A(n1092), .B(n1093), .Z(n96) );
  AND U547 ( .A(n95), .B(n96), .Z(n1685) );
  OR U548 ( .A(n1426), .B(n1427), .Z(n97) );
  NANDN U549 ( .A(n1429), .B(n1428), .Z(n98) );
  AND U550 ( .A(n97), .B(n98), .Z(n2017) );
  OR U551 ( .A(n1858), .B(n1857), .Z(n99) );
  NAND U552 ( .A(n1859), .B(n1860), .Z(n100) );
  AND U553 ( .A(n99), .B(n100), .Z(n1943) );
  OR U554 ( .A(n1456), .B(n1457), .Z(n101) );
  NANDN U555 ( .A(n1458), .B(n1459), .Z(n102) );
  AND U556 ( .A(n101), .B(n102), .Z(n1939) );
  OR U557 ( .A(n1468), .B(n1469), .Z(n103) );
  NANDN U558 ( .A(n1470), .B(n1471), .Z(n104) );
  AND U559 ( .A(n103), .B(n104), .Z(n1935) );
  XNOR U560 ( .A(n2059), .B(n2060), .Z(n2061) );
  OR U561 ( .A(n1761), .B(n1762), .Z(n105) );
  NANDN U562 ( .A(n1764), .B(n1763), .Z(n106) );
  NAND U563 ( .A(n105), .B(n106), .Z(n2055) );
  OR U564 ( .A(n1612), .B(n1613), .Z(n107) );
  NANDN U565 ( .A(n1615), .B(n1614), .Z(n108) );
  AND U566 ( .A(n107), .B(n108), .Z(n2129) );
  NANDN U567 ( .A(n1652), .B(n1653), .Z(n109) );
  NANDN U568 ( .A(n1650), .B(n1651), .Z(n110) );
  NAND U569 ( .A(n109), .B(n110), .Z(n1949) );
  NANDN U570 ( .A(n1820), .B(n1819), .Z(n111) );
  NANDN U571 ( .A(n1821), .B(n1822), .Z(n112) );
  NAND U572 ( .A(n111), .B(n112), .Z(n2107) );
  OR U573 ( .A(n1927), .B(n1928), .Z(n113) );
  OR U574 ( .A(n1926), .B(n1925), .Z(n114) );
  NAND U575 ( .A(n113), .B(n114), .Z(n2218) );
  OR U576 ( .A(n2139), .B(n2140), .Z(n115) );
  NANDN U577 ( .A(n2142), .B(n2141), .Z(n116) );
  AND U578 ( .A(n115), .B(n116), .Z(n2211) );
  NANDN U579 ( .A(n2097), .B(n2098), .Z(n117) );
  NANDN U580 ( .A(n2096), .B(n2095), .Z(n118) );
  AND U581 ( .A(n117), .B(n118), .Z(n2164) );
  NANDN U582 ( .A(n426), .B(n425), .Z(n119) );
  NANDN U583 ( .A(n427), .B(n428), .Z(n120) );
  NAND U584 ( .A(n119), .B(n120), .Z(n1523) );
  OR U585 ( .A(n1905), .B(n1906), .Z(n121) );
  NANDN U586 ( .A(n1907), .B(n1908), .Z(n122) );
  NAND U587 ( .A(n121), .B(n122), .Z(n2201) );
  OR U588 ( .A(n1953), .B(n1954), .Z(n123) );
  NAND U589 ( .A(n1956), .B(n1955), .Z(n124) );
  NAND U590 ( .A(n123), .B(n124), .Z(n2151) );
  OR U591 ( .A(n2214), .B(n2215), .Z(n125) );
  NANDN U592 ( .A(n2212), .B(n2213), .Z(n126) );
  AND U593 ( .A(n125), .B(n126), .Z(n2336) );
  OR U594 ( .A(n2300), .B(n2299), .Z(n127) );
  NAND U595 ( .A(n2301), .B(n2302), .Z(n128) );
  AND U596 ( .A(n127), .B(n128), .Z(n2358) );
  NAND U597 ( .A(n2351), .B(n2349), .Z(n129) );
  XOR U598 ( .A(n2349), .B(n2351), .Z(n130) );
  NANDN U599 ( .A(n2350), .B(n130), .Z(n131) );
  NAND U600 ( .A(n129), .B(n131), .Z(n2381) );
  OR U601 ( .A(n2354), .B(n2355), .Z(n132) );
  NANDN U602 ( .A(n2352), .B(n2353), .Z(n133) );
  AND U603 ( .A(n132), .B(n133), .Z(n2386) );
  OR U604 ( .A(n1308), .B(n1309), .Z(n134) );
  NANDN U605 ( .A(n1311), .B(n1310), .Z(n135) );
  NAND U606 ( .A(n134), .B(n135), .Z(n1567) );
  OR U607 ( .A(n457), .B(n458), .Z(n136) );
  NANDN U608 ( .A(n460), .B(n459), .Z(n137) );
  NAND U609 ( .A(n136), .B(n137), .Z(n1424) );
  OR U610 ( .A(n1136), .B(n1137), .Z(n138) );
  NANDN U611 ( .A(n1139), .B(n1138), .Z(n139) );
  NAND U612 ( .A(n138), .B(n139), .Z(n1417) );
  OR U613 ( .A(n1188), .B(n1189), .Z(n140) );
  NANDN U614 ( .A(n1191), .B(n1190), .Z(n141) );
  NAND U615 ( .A(n140), .B(n141), .Z(n1439) );
  OR U616 ( .A(n674), .B(n675), .Z(n142) );
  NANDN U617 ( .A(n677), .B(n676), .Z(n143) );
  NAND U618 ( .A(n142), .B(n143), .Z(n1537) );
  OR U619 ( .A(n768), .B(n769), .Z(n144) );
  NANDN U620 ( .A(n771), .B(n770), .Z(n145) );
  NAND U621 ( .A(n144), .B(n145), .Z(n1577) );
  OR U622 ( .A(n954), .B(n955), .Z(n146) );
  NANDN U623 ( .A(n957), .B(n956), .Z(n147) );
  AND U624 ( .A(n146), .B(n147), .Z(n1847) );
  XOR U625 ( .A(n1749), .B(n1750), .Z(n1752) );
  OR U626 ( .A(n832), .B(n833), .Z(n148) );
  NANDN U627 ( .A(n835), .B(n834), .Z(n149) );
  NAND U628 ( .A(n148), .B(n149), .Z(n1406) );
  OR U629 ( .A(n527), .B(n528), .Z(n150) );
  NANDN U630 ( .A(n530), .B(n529), .Z(n151) );
  NAND U631 ( .A(n150), .B(n151), .Z(n1403) );
  OR U632 ( .A(n890), .B(n891), .Z(n152) );
  NANDN U633 ( .A(n893), .B(n892), .Z(n153) );
  AND U634 ( .A(n152), .B(n153), .Z(n1859) );
  OR U635 ( .A(n1326), .B(n1327), .Z(n154) );
  NANDN U636 ( .A(n1329), .B(n1328), .Z(n155) );
  AND U637 ( .A(n154), .B(n155), .Z(n1729) );
  OR U638 ( .A(n978), .B(n979), .Z(n156) );
  NANDN U639 ( .A(n981), .B(n980), .Z(n157) );
  AND U640 ( .A(n156), .B(n157), .Z(n1397) );
  NANDN U641 ( .A(n1021), .B(n1020), .Z(n158) );
  NANDN U642 ( .A(n1022), .B(n1023), .Z(n159) );
  NAND U643 ( .A(n158), .B(n159), .Z(n1613) );
  OR U644 ( .A(n990), .B(n991), .Z(n160) );
  NANDN U645 ( .A(n993), .B(n992), .Z(n161) );
  AND U646 ( .A(n160), .B(n161), .Z(n1610) );
  NANDN U647 ( .A(n1045), .B(n1044), .Z(n162) );
  NANDN U648 ( .A(n1046), .B(n1047), .Z(n163) );
  NAND U649 ( .A(n162), .B(n163), .Z(n1714) );
  OR U650 ( .A(n391), .B(n392), .Z(n164) );
  NANDN U651 ( .A(n394), .B(n393), .Z(n165) );
  AND U652 ( .A(n164), .B(n165), .Z(n1594) );
  OR U653 ( .A(n443), .B(n444), .Z(n166) );
  NANDN U654 ( .A(n446), .B(n445), .Z(n167) );
  NAND U655 ( .A(n166), .B(n167), .Z(n1478) );
  NANDN U656 ( .A(n463), .B(n464), .Z(n168) );
  NANDN U657 ( .A(n462), .B(n461), .Z(n169) );
  AND U658 ( .A(n168), .B(n169), .Z(n1354) );
  OR U659 ( .A(n686), .B(n687), .Z(n170) );
  NANDN U660 ( .A(n689), .B(n688), .Z(n171) );
  NAND U661 ( .A(n170), .B(n171), .Z(n1599) );
  NANDN U662 ( .A(n1013), .B(n1012), .Z(n172) );
  NANDN U663 ( .A(n1010), .B(n1011), .Z(n173) );
  AND U664 ( .A(n172), .B(n173), .Z(n1691) );
  OR U665 ( .A(n1088), .B(n1089), .Z(n174) );
  NANDN U666 ( .A(n1091), .B(n1090), .Z(n175) );
  NAND U667 ( .A(n174), .B(n175), .Z(n1684) );
  XNOR U668 ( .A(n2034), .B(n2035), .Z(n2036) );
  OR U669 ( .A(n1862), .B(n1861), .Z(n176) );
  NAND U670 ( .A(n1863), .B(n1864), .Z(n177) );
  AND U671 ( .A(n176), .B(n177), .Z(n1944) );
  OR U672 ( .A(n1464), .B(n1465), .Z(n178) );
  NAND U673 ( .A(n1467), .B(n1466), .Z(n179) );
  NAND U674 ( .A(n178), .B(n179), .Z(n1937) );
  XOR U675 ( .A(n2065), .B(n2066), .Z(n2068) );
  OR U676 ( .A(n1781), .B(n1782), .Z(n180) );
  NANDN U677 ( .A(n1784), .B(n1783), .Z(n181) );
  NAND U678 ( .A(n180), .B(n181), .Z(n2062) );
  XOR U679 ( .A(n2053), .B(n2054), .Z(n2056) );
  XNOR U680 ( .A(n2089), .B(n2090), .Z(n2091) );
  XNOR U681 ( .A(n2099), .B(n2100), .Z(n2101) );
  NANDN U682 ( .A(n1702), .B(n1703), .Z(n182) );
  NANDN U683 ( .A(n1705), .B(n1704), .Z(n183) );
  NAND U684 ( .A(n182), .B(n183), .Z(n2024) );
  OR U685 ( .A(n387), .B(n388), .Z(n184) );
  NANDN U686 ( .A(n389), .B(n390), .Z(n185) );
  AND U687 ( .A(n184), .B(n185), .Z(n1650) );
  XNOR U688 ( .A(n2071), .B(n2072), .Z(n2073) );
  OR U689 ( .A(n1939), .B(n1940), .Z(n186) );
  NAND U690 ( .A(n1942), .B(n1941), .Z(n187) );
  NAND U691 ( .A(n186), .B(n187), .Z(n2193) );
  NANDN U692 ( .A(n2108), .B(n2107), .Z(n188) );
  NANDN U693 ( .A(n2105), .B(n2106), .Z(n189) );
  AND U694 ( .A(n188), .B(n189), .Z(n2156) );
  XOR U695 ( .A(oglobal[3]), .B(n2184), .Z(n190) );
  NANDN U696 ( .A(n2185), .B(n190), .Z(n191) );
  NAND U697 ( .A(oglobal[3]), .B(n2184), .Z(n192) );
  AND U698 ( .A(n191), .B(n192), .Z(n2329) );
  XOR U699 ( .A(n2176), .B(n2174), .Z(n193) );
  NAND U700 ( .A(n193), .B(n2175), .Z(n194) );
  NAND U701 ( .A(n2176), .B(n2174), .Z(n195) );
  AND U702 ( .A(n194), .B(n195), .Z(n2323) );
  OR U703 ( .A(n2209), .B(n2208), .Z(n196) );
  NAND U704 ( .A(n2210), .B(n2211), .Z(n197) );
  AND U705 ( .A(n196), .B(n197), .Z(n2339) );
  XNOR U706 ( .A(n2317), .B(n2318), .Z(n2319) );
  XOR U707 ( .A(n2110), .B(n2109), .Z(n2111) );
  XOR U708 ( .A(n2226), .B(n2227), .Z(n2229) );
  OR U709 ( .A(n2150), .B(n2151), .Z(n198) );
  NANDN U710 ( .A(n2153), .B(n2152), .Z(n199) );
  AND U711 ( .A(n198), .B(n199), .Z(n2313) );
  OR U712 ( .A(n1889), .B(n1890), .Z(n200) );
  NANDN U713 ( .A(n1892), .B(n1891), .Z(n201) );
  NAND U714 ( .A(n200), .B(n201), .Z(n2272) );
  OR U715 ( .A(n2311), .B(n2312), .Z(n202) );
  OR U716 ( .A(n2310), .B(n2309), .Z(n203) );
  NAND U717 ( .A(n202), .B(n203), .Z(n2355) );
  XOR U718 ( .A(n2389), .B(n2391), .Z(n204) );
  NANDN U719 ( .A(n2390), .B(n204), .Z(n205) );
  NAND U720 ( .A(n2389), .B(n2391), .Z(n206) );
  AND U721 ( .A(n205), .B(n206), .Z(n2397) );
  XOR U722 ( .A(n858), .B(n859), .Z(n861) );
  XNOR U723 ( .A(n1564), .B(n1565), .Z(n1566) );
  OR U724 ( .A(n319), .B(n320), .Z(n207) );
  NANDN U725 ( .A(n322), .B(n321), .Z(n208) );
  NAND U726 ( .A(n207), .B(n208), .Z(n1553) );
  XNOR U727 ( .A(n1416), .B(n1417), .Z(n1418) );
  OR U728 ( .A(n1270), .B(n1271), .Z(n209) );
  NANDN U729 ( .A(n1273), .B(n1272), .Z(n210) );
  NAND U730 ( .A(n209), .B(n210), .Z(n1431) );
  OR U731 ( .A(n722), .B(n723), .Z(n211) );
  NANDN U732 ( .A(n725), .B(n724), .Z(n212) );
  NAND U733 ( .A(n211), .B(n212), .Z(n1547) );
  OR U734 ( .A(n666), .B(n667), .Z(n213) );
  NANDN U735 ( .A(n669), .B(n668), .Z(n214) );
  NAND U736 ( .A(n213), .B(n214), .Z(n1535) );
  OR U737 ( .A(n938), .B(n939), .Z(n215) );
  NANDN U738 ( .A(n941), .B(n940), .Z(n216) );
  NAND U739 ( .A(n215), .B(n216), .Z(n1581) );
  XNOR U740 ( .A(n1586), .B(n1587), .Z(n1588) );
  OR U741 ( .A(n950), .B(n951), .Z(n217) );
  NANDN U742 ( .A(n953), .B(n952), .Z(n218) );
  NAND U743 ( .A(n217), .B(n218), .Z(n1848) );
  OR U744 ( .A(n574), .B(n575), .Z(n219) );
  NANDN U745 ( .A(n577), .B(n576), .Z(n220) );
  NAND U746 ( .A(n219), .B(n220), .Z(n1836) );
  OR U747 ( .A(n934), .B(n935), .Z(n221) );
  NANDN U748 ( .A(n937), .B(n936), .Z(n222) );
  AND U749 ( .A(n221), .B(n222), .Z(n1750) );
  OR U750 ( .A(n836), .B(n837), .Z(n223) );
  NANDN U751 ( .A(n839), .B(n838), .Z(n224) );
  AND U752 ( .A(n223), .B(n224), .Z(n1408) );
  OR U753 ( .A(n477), .B(n478), .Z(n225) );
  NANDN U754 ( .A(n480), .B(n479), .Z(n226) );
  NAND U755 ( .A(n225), .B(n226), .Z(n1461) );
  OR U756 ( .A(n465), .B(n466), .Z(n227) );
  NANDN U757 ( .A(n468), .B(n467), .Z(n228) );
  NAND U758 ( .A(n227), .B(n228), .Z(n1457) );
  OR U759 ( .A(n718), .B(n719), .Z(n229) );
  NANDN U760 ( .A(n721), .B(n720), .Z(n230) );
  NAND U761 ( .A(n229), .B(n230), .Z(n1735) );
  XNOR U762 ( .A(n1726), .B(n1727), .Z(n1728) );
  OR U763 ( .A(n560), .B(n561), .Z(n231) );
  NANDN U764 ( .A(n563), .B(n562), .Z(n232) );
  NAND U765 ( .A(n231), .B(n232), .Z(n1790) );
  OR U766 ( .A(n742), .B(n743), .Z(n233) );
  NANDN U767 ( .A(n745), .B(n744), .Z(n234) );
  NAND U768 ( .A(n233), .B(n234), .Z(n1765) );
  OR U769 ( .A(n546), .B(n547), .Z(n235) );
  NANDN U770 ( .A(n549), .B(n548), .Z(n236) );
  NAND U771 ( .A(n235), .B(n236), .Z(n1770) );
  OR U772 ( .A(n974), .B(n975), .Z(n237) );
  NANDN U773 ( .A(n977), .B(n976), .Z(n238) );
  NAND U774 ( .A(n237), .B(n238), .Z(n1396) );
  NANDN U775 ( .A(n1025), .B(n1024), .Z(n239) );
  NANDN U776 ( .A(n1026), .B(n1027), .Z(n240) );
  NAND U777 ( .A(n239), .B(n240), .Z(n1615) );
  XOR U778 ( .A(n1706), .B(n1707), .Z(n1709) );
  NANDN U779 ( .A(n1041), .B(n1040), .Z(n241) );
  NANDN U780 ( .A(n1042), .B(n1043), .Z(n242) );
  NAND U781 ( .A(n241), .B(n242), .Z(n1702) );
  OR U782 ( .A(n347), .B(n348), .Z(n243) );
  NANDN U783 ( .A(n350), .B(n349), .Z(n244) );
  AND U784 ( .A(n243), .B(n244), .Z(n1618) );
  OR U785 ( .A(n1102), .B(n1103), .Z(n245) );
  NANDN U786 ( .A(n1105), .B(n1104), .Z(n246) );
  NAND U787 ( .A(n245), .B(n246), .Z(n1832) );
  OR U788 ( .A(n764), .B(n765), .Z(n247) );
  NANDN U789 ( .A(n767), .B(n766), .Z(n248) );
  NAND U790 ( .A(n247), .B(n248), .Z(n1603) );
  OR U791 ( .A(n1000), .B(n1001), .Z(n249) );
  NANDN U792 ( .A(n1003), .B(n1002), .Z(n250) );
  NAND U793 ( .A(n249), .B(n250), .Z(n1693) );
  OR U794 ( .A(n1084), .B(n1085), .Z(n251) );
  NANDN U795 ( .A(n1087), .B(n1086), .Z(n252) );
  NAND U796 ( .A(n251), .B(n252), .Z(n1687) );
  NANDN U797 ( .A(n825), .B(n824), .Z(n253) );
  NANDN U798 ( .A(n826), .B(n827), .Z(n254) );
  NAND U799 ( .A(n253), .B(n254), .Z(n1493) );
  OR U800 ( .A(n1422), .B(n1423), .Z(n255) );
  NANDN U801 ( .A(n1424), .B(n1425), .Z(n256) );
  AND U802 ( .A(n255), .B(n256), .Z(n2018) );
  NANDN U803 ( .A(n1442), .B(n1443), .Z(n257) );
  NANDN U804 ( .A(n1445), .B(n1444), .Z(n258) );
  NAND U805 ( .A(n257), .B(n258), .Z(n2047) );
  OR U806 ( .A(n1576), .B(n1577), .Z(n259) );
  NANDN U807 ( .A(n1579), .B(n1578), .Z(n260) );
  NAND U808 ( .A(n259), .B(n260), .Z(n2037) );
  OR U809 ( .A(n1740), .B(n1741), .Z(n261) );
  NAND U810 ( .A(n1743), .B(n1742), .Z(n262) );
  NAND U811 ( .A(n261), .B(n262), .Z(n1996) );
  OR U812 ( .A(n1402), .B(n1403), .Z(n263) );
  NANDN U813 ( .A(n1404), .B(n1405), .Z(n264) );
  NAND U814 ( .A(n263), .B(n264), .Z(n2001) );
  OR U815 ( .A(n1452), .B(n1453), .Z(n265) );
  NANDN U816 ( .A(n1455), .B(n1454), .Z(n266) );
  NAND U817 ( .A(n265), .B(n266), .Z(n1941) );
  OR U818 ( .A(n1476), .B(n1477), .Z(n267) );
  NANDN U819 ( .A(n1478), .B(n1479), .Z(n268) );
  NAND U820 ( .A(n267), .B(n268), .Z(n1930) );
  XOR U821 ( .A(n1945), .B(n1946), .Z(n1984) );
  OR U822 ( .A(n1608), .B(n1609), .Z(n269) );
  NANDN U823 ( .A(n1610), .B(n1611), .Z(n270) );
  AND U824 ( .A(n269), .B(n270), .Z(n2131) );
  NANDN U825 ( .A(n1592), .B(n1593), .Z(n271) );
  NANDN U826 ( .A(n1594), .B(n1595), .Z(n272) );
  AND U827 ( .A(n271), .B(n272), .Z(n2139) );
  NANDN U828 ( .A(n1715), .B(n1714), .Z(n273) );
  NANDN U829 ( .A(n1712), .B(n1713), .Z(n274) );
  AND U830 ( .A(n273), .B(n274), .Z(n2027) );
  XOR U831 ( .A(n1655), .B(n1654), .Z(n1656) );
  OR U832 ( .A(n1596), .B(n1597), .Z(n275) );
  NANDN U833 ( .A(n1599), .B(n1598), .Z(n276) );
  NAND U834 ( .A(n275), .B(n276), .Z(n2074) );
  OR U835 ( .A(n1722), .B(n1723), .Z(n277) );
  NANDN U836 ( .A(n1725), .B(n1724), .Z(n278) );
  NAND U837 ( .A(n277), .B(n278), .Z(n1894) );
  OR U838 ( .A(n1935), .B(n1936), .Z(n279) );
  NAND U839 ( .A(n1938), .B(n1937), .Z(n280) );
  NAND U840 ( .A(n279), .B(n280), .Z(n2195) );
  XOR U841 ( .A(n2188), .B(n2189), .Z(n2169) );
  OR U842 ( .A(n2127), .B(n2128), .Z(n281) );
  OR U843 ( .A(n2126), .B(n2125), .Z(n282) );
  NAND U844 ( .A(n281), .B(n282), .Z(n2202) );
  OR U845 ( .A(n1951), .B(n1952), .Z(n283) );
  NANDN U846 ( .A(n1949), .B(n1950), .Z(n284) );
  AND U847 ( .A(n283), .B(n284), .Z(n2150) );
  XNOR U848 ( .A(n2325), .B(n2326), .Z(n2333) );
  OR U849 ( .A(n970), .B(n971), .Z(n285) );
  NANDN U850 ( .A(n972), .B(n973), .Z(n286) );
  NAND U851 ( .A(n285), .B(n286), .Z(n1796) );
  OR U852 ( .A(n1921), .B(n1922), .Z(n287) );
  NAND U853 ( .A(n1924), .B(n1923), .Z(n288) );
  NAND U854 ( .A(n287), .B(n288), .Z(n2227) );
  OR U855 ( .A(n2117), .B(n2118), .Z(n289) );
  NANDN U856 ( .A(n2116), .B(n2115), .Z(n290) );
  NAND U857 ( .A(n289), .B(n290), .Z(n2223) );
  OR U858 ( .A(n2198), .B(n2199), .Z(n291) );
  NANDN U859 ( .A(n2201), .B(n2200), .Z(n292) );
  NAND U860 ( .A(n291), .B(n292), .Z(n2295) );
  XOR U861 ( .A(n2338), .B(n2339), .Z(n2288) );
  NANDN U862 ( .A(n2238), .B(n2239), .Z(n293) );
  NANDN U863 ( .A(n2240), .B(n2241), .Z(n294) );
  AND U864 ( .A(n293), .B(n294), .Z(n2299) );
  NANDN U865 ( .A(n2154), .B(n2155), .Z(n295) );
  NANDN U866 ( .A(n2157), .B(n2156), .Z(n296) );
  NAND U867 ( .A(n295), .B(n296), .Z(n2314) );
  OR U868 ( .A(n2271), .B(n2272), .Z(n297) );
  NANDN U869 ( .A(n2274), .B(n2273), .Z(n298) );
  AND U870 ( .A(n297), .B(n298), .Z(n2281) );
  XNOR U871 ( .A(n2345), .B(n2346), .Z(n2350) );
  OR U872 ( .A(n2386), .B(n2387), .Z(n299) );
  OR U873 ( .A(n2385), .B(n2384), .Z(n300) );
  NAND U874 ( .A(n299), .B(n300), .Z(n2389) );
  XNOR U875 ( .A(x[330]), .B(y[330]), .Z(n1143) );
  XNOR U876 ( .A(x[33]), .B(y[33]), .Z(n1141) );
  XNOR U877 ( .A(x[332]), .B(y[332]), .Z(n1140) );
  XNOR U878 ( .A(n1141), .B(n1140), .Z(n1142) );
  XNOR U879 ( .A(n1143), .B(n1142), .Z(n1047) );
  XNOR U880 ( .A(x[374]), .B(y[374]), .Z(n557) );
  XNOR U881 ( .A(x[376]), .B(y[376]), .Z(n555) );
  XNOR U882 ( .A(x[395]), .B(y[395]), .Z(n554) );
  XNOR U883 ( .A(n555), .B(n554), .Z(n556) );
  XNOR U884 ( .A(n557), .B(n556), .Z(n1044) );
  XNOR U885 ( .A(x[326]), .B(y[326]), .Z(n1149) );
  XNOR U886 ( .A(x[328]), .B(y[328]), .Z(n1147) );
  XNOR U887 ( .A(x[383]), .B(y[383]), .Z(n1146) );
  XNOR U888 ( .A(n1147), .B(n1146), .Z(n1148) );
  XOR U889 ( .A(n1149), .B(n1148), .Z(n1045) );
  XOR U890 ( .A(n1044), .B(n1045), .Z(n1046) );
  XNOR U891 ( .A(n1047), .B(n1046), .Z(n1073) );
  XNOR U892 ( .A(x[350]), .B(y[350]), .Z(n354) );
  XNOR U893 ( .A(x[352]), .B(y[352]), .Z(n352) );
  XNOR U894 ( .A(x[389]), .B(y[389]), .Z(n351) );
  XNOR U895 ( .A(n352), .B(n351), .Z(n353) );
  XNOR U896 ( .A(n354), .B(n353), .Z(n464) );
  XNOR U897 ( .A(x[346]), .B(y[346]), .Z(n398) );
  XNOR U898 ( .A(x[25]), .B(y[25]), .Z(n396) );
  XNOR U899 ( .A(x[348]), .B(y[348]), .Z(n395) );
  XNOR U900 ( .A(n396), .B(n395), .Z(n397) );
  XNOR U901 ( .A(n398), .B(n397), .Z(n461) );
  XNOR U902 ( .A(x[358]), .B(y[358]), .Z(n1195) );
  XNOR U903 ( .A(x[360]), .B(y[360]), .Z(n1193) );
  XNOR U904 ( .A(x[391]), .B(y[391]), .Z(n1192) );
  XNOR U905 ( .A(n1193), .B(n1192), .Z(n1194) );
  XOR U906 ( .A(n1195), .B(n1194), .Z(n462) );
  XOR U907 ( .A(n461), .B(n462), .Z(n463) );
  XNOR U908 ( .A(n464), .B(n463), .Z(n1072) );
  XNOR U909 ( .A(n1073), .B(n1072), .Z(n1075) );
  XNOR U910 ( .A(x[322]), .B(y[322]), .Z(n1277) );
  XNOR U911 ( .A(x[37]), .B(y[37]), .Z(n1275) );
  XNOR U912 ( .A(x[324]), .B(y[324]), .Z(n1274) );
  XNOR U913 ( .A(n1275), .B(n1274), .Z(n1276) );
  XNOR U914 ( .A(n1277), .B(n1276), .Z(n1043) );
  XNOR U915 ( .A(x[378]), .B(y[378]), .Z(n494) );
  XNOR U916 ( .A(x[9]), .B(y[9]), .Z(n492) );
  XNOR U917 ( .A(x[380]), .B(y[380]), .Z(n491) );
  XNOR U918 ( .A(n492), .B(n491), .Z(n493) );
  XNOR U919 ( .A(n494), .B(n493), .Z(n1040) );
  XNOR U920 ( .A(x[318]), .B(y[318]), .Z(n1283) );
  XNOR U921 ( .A(x[320]), .B(y[320]), .Z(n1281) );
  XNOR U922 ( .A(x[381]), .B(y[381]), .Z(n1280) );
  XNOR U923 ( .A(n1281), .B(n1280), .Z(n1282) );
  XOR U924 ( .A(n1283), .B(n1282), .Z(n1041) );
  XOR U925 ( .A(n1040), .B(n1041), .Z(n1042) );
  XNOR U926 ( .A(n1043), .B(n1042), .Z(n1074) );
  XOR U927 ( .A(n1075), .B(n1074), .Z(n422) );
  XNOR U928 ( .A(x[338]), .B(y[338]), .Z(n1109) );
  XNOR U929 ( .A(x[29]), .B(y[29]), .Z(n1107) );
  XNOR U930 ( .A(x[340]), .B(y[340]), .Z(n1106) );
  XNOR U931 ( .A(n1107), .B(n1106), .Z(n1108) );
  XNOR U932 ( .A(n1109), .B(n1108), .Z(n897) );
  XNOR U933 ( .A(x[370]), .B(y[370]), .Z(n585) );
  XNOR U934 ( .A(x[13]), .B(y[13]), .Z(n583) );
  XNOR U935 ( .A(x[372]), .B(y[372]), .Z(n582) );
  XNOR U936 ( .A(n583), .B(n582), .Z(n584) );
  XNOR U937 ( .A(n585), .B(n584), .Z(n894) );
  XNOR U938 ( .A(x[334]), .B(y[334]), .Z(n1305) );
  XNOR U939 ( .A(x[336]), .B(y[336]), .Z(n1303) );
  XNOR U940 ( .A(x[385]), .B(y[385]), .Z(n1302) );
  XNOR U941 ( .A(n1303), .B(n1302), .Z(n1304) );
  XOR U942 ( .A(n1305), .B(n1304), .Z(n895) );
  XNOR U943 ( .A(n894), .B(n895), .Z(n896) );
  XOR U944 ( .A(n897), .B(n896), .Z(n1339) );
  XNOR U945 ( .A(x[342]), .B(y[342]), .Z(n1231) );
  XNOR U946 ( .A(x[344]), .B(y[344]), .Z(n1229) );
  XNOR U947 ( .A(x[387]), .B(y[387]), .Z(n1228) );
  XNOR U948 ( .A(n1229), .B(n1228), .Z(n1230) );
  XNOR U949 ( .A(n1231), .B(n1230), .Z(n543) );
  XNOR U950 ( .A(x[366]), .B(y[366]), .Z(n571) );
  XNOR U951 ( .A(x[368]), .B(y[368]), .Z(n569) );
  XNOR U952 ( .A(x[393]), .B(y[393]), .Z(n568) );
  XNOR U953 ( .A(n569), .B(n568), .Z(n570) );
  XNOR U954 ( .A(n571), .B(n570), .Z(n540) );
  XNOR U955 ( .A(x[362]), .B(y[362]), .Z(n1161) );
  XNOR U956 ( .A(x[17]), .B(y[17]), .Z(n1159) );
  XNOR U957 ( .A(x[364]), .B(y[364]), .Z(n1158) );
  XNOR U958 ( .A(n1159), .B(n1158), .Z(n1160) );
  XOR U959 ( .A(n1161), .B(n1160), .Z(n541) );
  XNOR U960 ( .A(n540), .B(n541), .Z(n542) );
  XOR U961 ( .A(n543), .B(n542), .Z(n1336) );
  XNOR U962 ( .A(x[354]), .B(y[354]), .Z(n322) );
  XNOR U963 ( .A(x[21]), .B(y[21]), .Z(n320) );
  XNOR U964 ( .A(x[356]), .B(y[356]), .Z(n319) );
  XOR U965 ( .A(n320), .B(n319), .Z(n321) );
  XOR U966 ( .A(n322), .B(n321), .Z(n1337) );
  XOR U967 ( .A(n1336), .B(n1337), .Z(n1338) );
  XNOR U968 ( .A(n1339), .B(n1338), .Z(n419) );
  XNOR U969 ( .A(x[294]), .B(y[294]), .Z(n1329) );
  XNOR U970 ( .A(x[296]), .B(y[296]), .Z(n1327) );
  XNOR U971 ( .A(x[375]), .B(y[375]), .Z(n1326) );
  XOR U972 ( .A(n1327), .B(n1326), .Z(n1328) );
  XOR U973 ( .A(n1329), .B(n1328), .Z(n1084) );
  XNOR U974 ( .A(x[390]), .B(y[390]), .Z(n831) );
  XNOR U975 ( .A(x[392]), .B(y[392]), .Z(n829) );
  XNOR U976 ( .A(x[399]), .B(y[399]), .Z(n828) );
  XOR U977 ( .A(n829), .B(n828), .Z(n830) );
  XOR U978 ( .A(n831), .B(n830), .Z(n1085) );
  XOR U979 ( .A(n1084), .B(n1085), .Z(n1086) );
  XNOR U980 ( .A(x[298]), .B(y[298]), .Z(n1191) );
  XNOR U981 ( .A(x[49]), .B(y[49]), .Z(n1189) );
  XNOR U982 ( .A(x[300]), .B(y[300]), .Z(n1188) );
  XOR U983 ( .A(n1189), .B(n1188), .Z(n1190) );
  XOR U984 ( .A(n1191), .B(n1190), .Z(n1087) );
  XNOR U985 ( .A(n1086), .B(n1087), .Z(n996) );
  XNOR U986 ( .A(x[302]), .B(y[302]), .Z(n1273) );
  XNOR U987 ( .A(x[304]), .B(y[304]), .Z(n1271) );
  XNOR U988 ( .A(x[377]), .B(y[377]), .Z(n1270) );
  XOR U989 ( .A(n1271), .B(n1270), .Z(n1272) );
  XOR U990 ( .A(n1273), .B(n1272), .Z(n1088) );
  XNOR U991 ( .A(x[386]), .B(y[386]), .Z(n811) );
  XNOR U992 ( .A(x[5]), .B(y[5]), .Z(n809) );
  XNOR U993 ( .A(x[388]), .B(y[388]), .Z(n808) );
  XOR U994 ( .A(n809), .B(n808), .Z(n810) );
  XOR U995 ( .A(n811), .B(n810), .Z(n1089) );
  XOR U996 ( .A(n1088), .B(n1089), .Z(n1090) );
  XNOR U997 ( .A(x[306]), .B(y[306]), .Z(n1321) );
  XNOR U998 ( .A(x[45]), .B(y[45]), .Z(n1319) );
  XNOR U999 ( .A(x[308]), .B(y[308]), .Z(n1318) );
  XOR U1000 ( .A(n1319), .B(n1318), .Z(n1320) );
  XOR U1001 ( .A(n1321), .B(n1320), .Z(n1091) );
  XNOR U1002 ( .A(n1090), .B(n1091), .Z(n994) );
  XNOR U1003 ( .A(x[310]), .B(y[310]), .Z(n1185) );
  XNOR U1004 ( .A(x[312]), .B(y[312]), .Z(n1183) );
  XNOR U1005 ( .A(x[379]), .B(y[379]), .Z(n1182) );
  XNOR U1006 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U1007 ( .A(n1185), .B(n1184), .Z(n1029) );
  XNOR U1008 ( .A(x[382]), .B(y[382]), .Z(n627) );
  XNOR U1009 ( .A(x[384]), .B(y[384]), .Z(n625) );
  XNOR U1010 ( .A(x[397]), .B(y[397]), .Z(n624) );
  XNOR U1011 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1012 ( .A(n627), .B(n626), .Z(n1028) );
  XOR U1013 ( .A(n1029), .B(n1028), .Z(n1030) );
  XNOR U1014 ( .A(x[314]), .B(y[314]), .Z(n1179) );
  XNOR U1015 ( .A(x[41]), .B(y[41]), .Z(n1177) );
  XNOR U1016 ( .A(x[316]), .B(y[316]), .Z(n1176) );
  XNOR U1017 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U1018 ( .A(n1179), .B(n1178), .Z(n1031) );
  XNOR U1019 ( .A(n1030), .B(n1031), .Z(n995) );
  XNOR U1020 ( .A(n994), .B(n995), .Z(n997) );
  XNOR U1021 ( .A(n996), .B(n997), .Z(n420) );
  XOR U1022 ( .A(n419), .B(n420), .Z(n421) );
  XOR U1023 ( .A(n422), .B(n421), .Z(n1342) );
  XNOR U1024 ( .A(x[36]), .B(y[36]), .Z(n805) );
  XNOR U1025 ( .A(x[38]), .B(y[38]), .Z(n802) );
  XNOR U1026 ( .A(x[40]), .B(y[40]), .Z(n803) );
  XOR U1027 ( .A(n802), .B(n803), .Z(n804) );
  XNOR U1028 ( .A(n805), .B(n804), .Z(n371) );
  XNOR U1029 ( .A(x[30]), .B(y[30]), .Z(n799) );
  XNOR U1030 ( .A(x[32]), .B(y[32]), .Z(n796) );
  XNOR U1031 ( .A(x[34]), .B(y[34]), .Z(n797) );
  XOR U1032 ( .A(n796), .B(n797), .Z(n798) );
  XNOR U1033 ( .A(n799), .B(n798), .Z(n369) );
  XNOR U1034 ( .A(x[24]), .B(y[24]), .Z(n793) );
  XNOR U1035 ( .A(x[26]), .B(y[26]), .Z(n790) );
  XNOR U1036 ( .A(x[28]), .B(y[28]), .Z(n791) );
  XOR U1037 ( .A(n790), .B(n791), .Z(n792) );
  XNOR U1038 ( .A(n793), .B(n792), .Z(n370) );
  XNOR U1039 ( .A(n369), .B(n370), .Z(n372) );
  XNOR U1040 ( .A(n371), .B(n372), .Z(n342) );
  XNOR U1041 ( .A(x[54]), .B(y[54]), .Z(n855) );
  XNOR U1042 ( .A(x[56]), .B(y[56]), .Z(n852) );
  XNOR U1043 ( .A(x[58]), .B(y[58]), .Z(n853) );
  XOR U1044 ( .A(n852), .B(n853), .Z(n854) );
  XNOR U1045 ( .A(n855), .B(n854), .Z(n415) );
  XNOR U1046 ( .A(x[48]), .B(y[48]), .Z(n843) );
  XNOR U1047 ( .A(x[50]), .B(y[50]), .Z(n840) );
  XNOR U1048 ( .A(x[52]), .B(y[52]), .Z(n841) );
  XOR U1049 ( .A(n840), .B(n841), .Z(n842) );
  XNOR U1050 ( .A(n843), .B(n842), .Z(n413) );
  XNOR U1051 ( .A(x[42]), .B(y[42]), .Z(n849) );
  XNOR U1052 ( .A(x[44]), .B(y[44]), .Z(n846) );
  XNOR U1053 ( .A(x[46]), .B(y[46]), .Z(n847) );
  XOR U1054 ( .A(n846), .B(n847), .Z(n848) );
  XNOR U1055 ( .A(n849), .B(n848), .Z(n414) );
  XNOR U1056 ( .A(n413), .B(n414), .Z(n416) );
  XNOR U1057 ( .A(n415), .B(n416), .Z(n341) );
  XOR U1058 ( .A(n342), .B(n341), .Z(n343) );
  XNOR U1059 ( .A(x[18]), .B(y[18]), .Z(n893) );
  XNOR U1060 ( .A(x[20]), .B(y[20]), .Z(n891) );
  XNOR U1061 ( .A(x[22]), .B(y[22]), .Z(n890) );
  XOR U1062 ( .A(n891), .B(n890), .Z(n892) );
  XOR U1063 ( .A(n893), .B(n892), .Z(n1249) );
  XNOR U1064 ( .A(x[12]), .B(y[12]), .Z(n885) );
  XNOR U1065 ( .A(x[14]), .B(y[14]), .Z(n883) );
  XNOR U1066 ( .A(x[16]), .B(y[16]), .Z(n882) );
  XOR U1067 ( .A(n883), .B(n882), .Z(n884) );
  XOR U1068 ( .A(n885), .B(n884), .Z(n1246) );
  XNOR U1069 ( .A(x[6]), .B(y[6]), .Z(n889) );
  XNOR U1070 ( .A(x[8]), .B(y[8]), .Z(n887) );
  XNOR U1071 ( .A(x[10]), .B(y[10]), .Z(n886) );
  XOR U1072 ( .A(n887), .B(n886), .Z(n888) );
  XNOR U1073 ( .A(n889), .B(n888), .Z(n1247) );
  XNOR U1074 ( .A(n1246), .B(n1247), .Z(n1248) );
  XNOR U1075 ( .A(n1249), .B(n1248), .Z(n344) );
  XOR U1076 ( .A(n343), .B(n344), .Z(n787) );
  XNOR U1077 ( .A(x[245]), .B(y[245]), .Z(n663) );
  XNOR U1078 ( .A(x[243]), .B(y[243]), .Z(n661) );
  XNOR U1079 ( .A(x[323]), .B(y[323]), .Z(n660) );
  XNOR U1080 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U1081 ( .A(n663), .B(n662), .Z(n1287) );
  XNOR U1082 ( .A(x[241]), .B(y[241]), .Z(n699) );
  XNOR U1083 ( .A(x[239]), .B(y[239]), .Z(n697) );
  XNOR U1084 ( .A(x[325]), .B(y[325]), .Z(n696) );
  XNOR U1085 ( .A(n697), .B(n696), .Z(n698) );
  XNOR U1086 ( .A(n699), .B(n698), .Z(n1286) );
  XOR U1087 ( .A(n1287), .B(n1286), .Z(n1288) );
  XNOR U1088 ( .A(x[237]), .B(y[237]), .Z(n693) );
  XNOR U1089 ( .A(x[235]), .B(y[235]), .Z(n691) );
  XNOR U1090 ( .A(x[327]), .B(y[327]), .Z(n690) );
  XNOR U1091 ( .A(n691), .B(n690), .Z(n692) );
  XNOR U1092 ( .A(n693), .B(n692), .Z(n1289) );
  XOR U1093 ( .A(n1288), .B(n1289), .Z(n389) );
  XNOR U1094 ( .A(x[261]), .B(y[261]), .Z(n741) );
  XNOR U1095 ( .A(x[259]), .B(y[259]), .Z(n739) );
  XNOR U1096 ( .A(x[315]), .B(y[315]), .Z(n738) );
  XOR U1097 ( .A(n739), .B(n738), .Z(n740) );
  XOR U1098 ( .A(n741), .B(n740), .Z(n338) );
  XNOR U1099 ( .A(x[265]), .B(y[265]), .Z(n745) );
  XNOR U1100 ( .A(x[263]), .B(y[263]), .Z(n743) );
  XNOR U1101 ( .A(x[313]), .B(y[313]), .Z(n742) );
  XOR U1102 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U1103 ( .A(n745), .B(n744), .Z(n336) );
  XNOR U1104 ( .A(x[269]), .B(y[269]), .Z(n721) );
  XNOR U1105 ( .A(x[267]), .B(y[267]), .Z(n719) );
  XNOR U1106 ( .A(x[311]), .B(y[311]), .Z(n718) );
  XOR U1107 ( .A(n719), .B(n718), .Z(n720) );
  XOR U1108 ( .A(n721), .B(n720), .Z(n335) );
  XNOR U1109 ( .A(n336), .B(n335), .Z(n337) );
  XOR U1110 ( .A(n338), .B(n337), .Z(n387) );
  XNOR U1111 ( .A(x[257]), .B(y[257]), .Z(n749) );
  XNOR U1112 ( .A(x[255]), .B(y[255]), .Z(n747) );
  XNOR U1113 ( .A(x[317]), .B(y[317]), .Z(n746) );
  XNOR U1114 ( .A(n747), .B(n746), .Z(n748) );
  XNOR U1115 ( .A(n749), .B(n748), .Z(n1125) );
  XNOR U1116 ( .A(x[253]), .B(y[253]), .Z(n657) );
  XNOR U1117 ( .A(x[251]), .B(y[251]), .Z(n655) );
  XNOR U1118 ( .A(x[319]), .B(y[319]), .Z(n654) );
  XNOR U1119 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1120 ( .A(n657), .B(n656), .Z(n1124) );
  XOR U1121 ( .A(n1125), .B(n1124), .Z(n1126) );
  XNOR U1122 ( .A(x[249]), .B(y[249]), .Z(n651) );
  XNOR U1123 ( .A(x[247]), .B(y[247]), .Z(n649) );
  XNOR U1124 ( .A(x[321]), .B(y[321]), .Z(n648) );
  XNOR U1125 ( .A(n649), .B(n648), .Z(n650) );
  XNOR U1126 ( .A(n651), .B(n650), .Z(n1127) );
  XOR U1127 ( .A(n1126), .B(n1127), .Z(n388) );
  XOR U1128 ( .A(n387), .B(n388), .Z(n390) );
  XNOR U1129 ( .A(n389), .B(n390), .Z(n784) );
  XNOR U1130 ( .A(x[91]), .B(y[91]), .Z(n488) );
  XNOR U1131 ( .A(x[83]), .B(y[83]), .Z(n485) );
  XNOR U1132 ( .A(x[87]), .B(y[87]), .Z(n486) );
  XOR U1133 ( .A(n485), .B(n486), .Z(n487) );
  XOR U1134 ( .A(n488), .B(n487), .Z(n391) );
  XNOR U1135 ( .A(x[79]), .B(y[79]), .Z(n609) );
  XNOR U1136 ( .A(x[71]), .B(y[71]), .Z(n606) );
  XNOR U1137 ( .A(x[75]), .B(y[75]), .Z(n607) );
  XOR U1138 ( .A(n606), .B(n607), .Z(n608) );
  XOR U1139 ( .A(n609), .B(n608), .Z(n392) );
  XOR U1140 ( .A(n391), .B(n392), .Z(n393) );
  XNOR U1141 ( .A(x[67]), .B(y[67]), .Z(n621) );
  XNOR U1142 ( .A(x[59]), .B(y[59]), .Z(n618) );
  XNOR U1143 ( .A(x[63]), .B(y[63]), .Z(n619) );
  XOR U1144 ( .A(n618), .B(n619), .Z(n620) );
  XOR U1145 ( .A(n621), .B(n620), .Z(n394) );
  XNOR U1146 ( .A(n393), .B(n394), .Z(n644) );
  XNOR U1147 ( .A(x[55]), .B(y[55]), .Z(n1063) );
  XNOR U1148 ( .A(x[47]), .B(y[47]), .Z(n1060) );
  XNOR U1149 ( .A(x[51]), .B(y[51]), .Z(n1061) );
  XOR U1150 ( .A(n1060), .B(n1061), .Z(n1062) );
  XOR U1151 ( .A(n1063), .B(n1062), .Z(n1225) );
  XNOR U1152 ( .A(x[43]), .B(y[43]), .Z(n1057) );
  XNOR U1153 ( .A(x[35]), .B(y[35]), .Z(n1054) );
  XNOR U1154 ( .A(x[39]), .B(y[39]), .Z(n1055) );
  XOR U1155 ( .A(n1054), .B(n1055), .Z(n1056) );
  XOR U1156 ( .A(n1057), .B(n1056), .Z(n1222) );
  XNOR U1157 ( .A(x[31]), .B(y[31]), .Z(n1069) );
  XNOR U1158 ( .A(x[23]), .B(y[23]), .Z(n1066) );
  XNOR U1159 ( .A(x[27]), .B(y[27]), .Z(n1067) );
  XOR U1160 ( .A(n1066), .B(n1067), .Z(n1068) );
  XNOR U1161 ( .A(n1069), .B(n1068), .Z(n1223) );
  XNOR U1162 ( .A(n1222), .B(n1223), .Z(n1224) );
  XNOR U1163 ( .A(n1225), .B(n1224), .Z(n643) );
  XNOR U1164 ( .A(x[19]), .B(y[19]), .Z(n873) );
  XNOR U1165 ( .A(x[11]), .B(y[11]), .Z(n870) );
  XNOR U1166 ( .A(x[15]), .B(y[15]), .Z(n871) );
  XOR U1167 ( .A(n870), .B(n871), .Z(n872) );
  XOR U1168 ( .A(n873), .B(n872), .Z(n1102) );
  XNOR U1169 ( .A(x[7]), .B(y[7]), .Z(n867) );
  XNOR U1170 ( .A(x[1]), .B(y[1]), .Z(n864) );
  XNOR U1171 ( .A(x[3]), .B(y[3]), .Z(n865) );
  XOR U1172 ( .A(n864), .B(n865), .Z(n866) );
  XOR U1173 ( .A(n867), .B(n866), .Z(n1103) );
  XOR U1174 ( .A(n1102), .B(n1103), .Z(n1104) );
  XNOR U1175 ( .A(x[0]), .B(y[0]), .Z(n879) );
  XNOR U1176 ( .A(x[2]), .B(y[2]), .Z(n876) );
  XNOR U1177 ( .A(x[4]), .B(y[4]), .Z(n877) );
  XOR U1178 ( .A(n876), .B(n877), .Z(n878) );
  XOR U1179 ( .A(n879), .B(n878), .Z(n1105) );
  XNOR U1180 ( .A(n1104), .B(n1105), .Z(n642) );
  XOR U1181 ( .A(n643), .B(n642), .Z(n645) );
  XOR U1182 ( .A(n644), .B(n645), .Z(n785) );
  XOR U1183 ( .A(n784), .B(n785), .Z(n786) );
  XNOR U1184 ( .A(n787), .B(n786), .Z(n1343) );
  XNOR U1185 ( .A(n1342), .B(n1343), .Z(n1344) );
  XNOR U1186 ( .A(x[155]), .B(y[155]), .Z(n771) );
  XNOR U1187 ( .A(x[151]), .B(y[151]), .Z(n769) );
  XNOR U1188 ( .A(x[153]), .B(y[153]), .Z(n768) );
  XOR U1189 ( .A(n769), .B(n768), .Z(n770) );
  XNOR U1190 ( .A(n771), .B(n770), .Z(n1314) );
  XNOR U1191 ( .A(x[161]), .B(y[161]), .Z(n673) );
  XNOR U1192 ( .A(x[157]), .B(y[157]), .Z(n671) );
  XNOR U1193 ( .A(x[159]), .B(y[159]), .Z(n670) );
  XOR U1194 ( .A(n671), .B(n670), .Z(n672) );
  XNOR U1195 ( .A(n673), .B(n672), .Z(n1312) );
  XNOR U1196 ( .A(x[167]), .B(y[167]), .Z(n949) );
  XNOR U1197 ( .A(x[163]), .B(y[163]), .Z(n947) );
  XNOR U1198 ( .A(x[165]), .B(y[165]), .Z(n946) );
  XOR U1199 ( .A(n947), .B(n946), .Z(n948) );
  XNOR U1200 ( .A(n949), .B(n948), .Z(n1313) );
  XNOR U1201 ( .A(n1312), .B(n1313), .Z(n1315) );
  XNOR U1202 ( .A(n1314), .B(n1315), .Z(n310) );
  XNOR U1203 ( .A(x[149]), .B(y[149]), .Z(n725) );
  XNOR U1204 ( .A(x[145]), .B(y[145]), .Z(n723) );
  XNOR U1205 ( .A(x[147]), .B(y[147]), .Z(n722) );
  XOR U1206 ( .A(n723), .B(n722), .Z(n724) );
  XOR U1207 ( .A(n725), .B(n724), .Z(n1259) );
  XNOR U1208 ( .A(x[143]), .B(y[143]), .Z(n669) );
  XNOR U1209 ( .A(x[139]), .B(y[139]), .Z(n667) );
  XNOR U1210 ( .A(x[141]), .B(y[141]), .Z(n666) );
  XOR U1211 ( .A(n667), .B(n666), .Z(n668) );
  XNOR U1212 ( .A(n669), .B(n668), .Z(n1258) );
  XNOR U1213 ( .A(n1259), .B(n1258), .Z(n1261) );
  XNOR U1214 ( .A(x[137]), .B(y[137]), .Z(n957) );
  XNOR U1215 ( .A(x[131]), .B(y[131]), .Z(n955) );
  XNOR U1216 ( .A(x[135]), .B(y[135]), .Z(n954) );
  XOR U1217 ( .A(n955), .B(n954), .Z(n956) );
  XNOR U1218 ( .A(n957), .B(n956), .Z(n1260) );
  XOR U1219 ( .A(n1261), .B(n1260), .Z(n308) );
  XNOR U1220 ( .A(x[127]), .B(y[127]), .Z(n450) );
  XNOR U1221 ( .A(x[119]), .B(y[119]), .Z(n447) );
  XNOR U1222 ( .A(x[123]), .B(y[123]), .Z(n448) );
  XOR U1223 ( .A(n447), .B(n448), .Z(n449) );
  XOR U1224 ( .A(n450), .B(n449), .Z(n1131) );
  XNOR U1225 ( .A(x[115]), .B(y[115]), .Z(n961) );
  XNOR U1226 ( .A(x[107]), .B(y[107]), .Z(n958) );
  XNOR U1227 ( .A(x[111]), .B(y[111]), .Z(n959) );
  XOR U1228 ( .A(n958), .B(n959), .Z(n960) );
  XNOR U1229 ( .A(n961), .B(n960), .Z(n1130) );
  XNOR U1230 ( .A(n1131), .B(n1130), .Z(n1133) );
  XNOR U1231 ( .A(x[103]), .B(y[103]), .Z(n615) );
  XNOR U1232 ( .A(x[95]), .B(y[95]), .Z(n612) );
  XNOR U1233 ( .A(x[99]), .B(y[99]), .Z(n613) );
  XOR U1234 ( .A(n612), .B(n613), .Z(n614) );
  XNOR U1235 ( .A(n615), .B(n614), .Z(n1132) );
  XOR U1236 ( .A(n1133), .B(n1132), .Z(n307) );
  XOR U1237 ( .A(n308), .B(n307), .Z(n309) );
  XOR U1238 ( .A(n310), .B(n309), .Z(n428) );
  XNOR U1239 ( .A(x[233]), .B(y[233]), .Z(n705) );
  XNOR U1240 ( .A(x[231]), .B(y[231]), .Z(n703) );
  XNOR U1241 ( .A(x[329]), .B(y[329]), .Z(n702) );
  XNOR U1242 ( .A(n703), .B(n702), .Z(n704) );
  XNOR U1243 ( .A(n705), .B(n704), .Z(n1293) );
  XNOR U1244 ( .A(x[229]), .B(y[229]), .Z(n597) );
  XNOR U1245 ( .A(x[227]), .B(y[227]), .Z(n595) );
  XNOR U1246 ( .A(x[331]), .B(y[331]), .Z(n594) );
  XNOR U1247 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U1248 ( .A(n597), .B(n596), .Z(n1292) );
  XOR U1249 ( .A(n1293), .B(n1292), .Z(n1294) );
  XNOR U1250 ( .A(x[225]), .B(y[225]), .Z(n591) );
  XNOR U1251 ( .A(x[223]), .B(y[223]), .Z(n589) );
  XNOR U1252 ( .A(x[333]), .B(y[333]), .Z(n588) );
  XNOR U1253 ( .A(n589), .B(n588), .Z(n590) );
  XNOR U1254 ( .A(n591), .B(n590), .Z(n1295) );
  XOR U1255 ( .A(n1294), .B(n1295), .Z(n378) );
  XNOR U1256 ( .A(x[215]), .B(y[215]), .Z(n761) );
  XNOR U1257 ( .A(x[211]), .B(y[211]), .Z(n758) );
  XNOR U1258 ( .A(x[213]), .B(y[213]), .Z(n759) );
  XOR U1259 ( .A(n758), .B(n759), .Z(n760) );
  XOR U1260 ( .A(n761), .B(n760), .Z(n1153) );
  XNOR U1261 ( .A(x[209]), .B(y[209]), .Z(n755) );
  XNOR U1262 ( .A(x[205]), .B(y[205]), .Z(n752) );
  XNOR U1263 ( .A(x[207]), .B(y[207]), .Z(n753) );
  XOR U1264 ( .A(n752), .B(n753), .Z(n754) );
  XNOR U1265 ( .A(n755), .B(n754), .Z(n1152) );
  XNOR U1266 ( .A(n1153), .B(n1152), .Z(n1155) );
  XNOR U1267 ( .A(x[221]), .B(y[221]), .Z(n603) );
  XNOR U1268 ( .A(x[217]), .B(y[217]), .Z(n600) );
  XNOR U1269 ( .A(x[219]), .B(y[219]), .Z(n601) );
  XOR U1270 ( .A(n600), .B(n601), .Z(n602) );
  XNOR U1271 ( .A(n603), .B(n602), .Z(n1154) );
  XOR U1272 ( .A(n1155), .B(n1154), .Z(n375) );
  XNOR U1273 ( .A(x[275]), .B(y[275]), .Z(n937) );
  XNOR U1274 ( .A(x[289]), .B(y[289]), .Z(n935) );
  XNOR U1275 ( .A(x[301]), .B(y[301]), .Z(n934) );
  XOR U1276 ( .A(n935), .B(n934), .Z(n936) );
  XNOR U1277 ( .A(n937), .B(n936), .Z(n315) );
  XNOR U1278 ( .A(x[273]), .B(y[273]), .Z(n711) );
  XNOR U1279 ( .A(x[271]), .B(y[271]), .Z(n709) );
  XNOR U1280 ( .A(x[309]), .B(y[309]), .Z(n708) );
  XOR U1281 ( .A(n709), .B(n708), .Z(n710) );
  XNOR U1282 ( .A(n711), .B(n710), .Z(n313) );
  XNOR U1283 ( .A(x[283]), .B(y[283]), .Z(n925) );
  XNOR U1284 ( .A(x[285]), .B(y[285]), .Z(n924) );
  XOR U1285 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U1286 ( .A(x[277]), .B(y[277]), .Z(n909) );
  XNOR U1287 ( .A(x[279]), .B(y[279]), .Z(n907) );
  XNOR U1288 ( .A(x[293]), .B(y[293]), .Z(n906) );
  XNOR U1289 ( .A(n907), .B(n906), .Z(n908) );
  XNOR U1290 ( .A(n909), .B(n908), .Z(n927) );
  XNOR U1291 ( .A(n926), .B(n927), .Z(n314) );
  XNOR U1292 ( .A(n313), .B(n314), .Z(n316) );
  XNOR U1293 ( .A(n315), .B(n316), .Z(n376) );
  XOR U1294 ( .A(n375), .B(n376), .Z(n377) );
  XNOR U1295 ( .A(n378), .B(n377), .Z(n425) );
  XNOR U1296 ( .A(x[203]), .B(y[203]), .Z(n767) );
  XNOR U1297 ( .A(x[199]), .B(y[199]), .Z(n765) );
  XNOR U1298 ( .A(x[201]), .B(y[201]), .Z(n764) );
  XOR U1299 ( .A(n765), .B(n764), .Z(n766) );
  XOR U1300 ( .A(n767), .B(n766), .Z(n1265) );
  XNOR U1301 ( .A(x[197]), .B(y[197]), .Z(n685) );
  XNOR U1302 ( .A(x[193]), .B(y[193]), .Z(n683) );
  XNOR U1303 ( .A(x[195]), .B(y[195]), .Z(n682) );
  XOR U1304 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U1305 ( .A(n685), .B(n684), .Z(n1264) );
  XNOR U1306 ( .A(n1265), .B(n1264), .Z(n1267) );
  XNOR U1307 ( .A(x[191]), .B(y[191]), .Z(n681) );
  XNOR U1308 ( .A(x[187]), .B(y[187]), .Z(n679) );
  XNOR U1309 ( .A(x[189]), .B(y[189]), .Z(n678) );
  XOR U1310 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U1311 ( .A(n681), .B(n680), .Z(n1266) );
  XOR U1312 ( .A(n1267), .B(n1266), .Z(n303) );
  XNOR U1313 ( .A(x[173]), .B(y[173]), .Z(n941) );
  XNOR U1314 ( .A(x[169]), .B(y[169]), .Z(n939) );
  XNOR U1315 ( .A(x[171]), .B(y[171]), .Z(n938) );
  XOR U1316 ( .A(n939), .B(n938), .Z(n940) );
  XOR U1317 ( .A(n941), .B(n940), .Z(n1331) );
  XNOR U1318 ( .A(x[179]), .B(y[179]), .Z(n945) );
  XNOR U1319 ( .A(x[175]), .B(y[175]), .Z(n943) );
  XNOR U1320 ( .A(x[177]), .B(y[177]), .Z(n942) );
  XOR U1321 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U1322 ( .A(n945), .B(n944), .Z(n1330) );
  XNOR U1323 ( .A(n1331), .B(n1330), .Z(n1333) );
  XNOR U1324 ( .A(x[185]), .B(y[185]), .Z(n689) );
  XNOR U1325 ( .A(x[181]), .B(y[181]), .Z(n687) );
  XNOR U1326 ( .A(x[183]), .B(y[183]), .Z(n686) );
  XOR U1327 ( .A(n687), .B(n686), .Z(n688) );
  XNOR U1328 ( .A(n689), .B(n688), .Z(n1332) );
  XOR U1329 ( .A(n1333), .B(n1332), .Z(n302) );
  XNOR U1330 ( .A(x[303]), .B(y[303]), .Z(n715) );
  XNOR U1331 ( .A(x[305]), .B(y[305]), .Z(n713) );
  XNOR U1332 ( .A(x[307]), .B(y[307]), .Z(n712) );
  XNOR U1333 ( .A(n713), .B(n712), .Z(n714) );
  XNOR U1334 ( .A(n715), .B(n714), .Z(n827) );
  XNOR U1335 ( .A(x[287]), .B(y[287]), .Z(n931) );
  XNOR U1336 ( .A(x[281]), .B(y[281]), .Z(n929) );
  XNOR U1337 ( .A(x[291]), .B(y[291]), .Z(n928) );
  XNOR U1338 ( .A(n929), .B(n928), .Z(n930) );
  XNOR U1339 ( .A(n931), .B(n930), .Z(n824) );
  XNOR U1340 ( .A(x[295]), .B(y[295]), .Z(n915) );
  XNOR U1341 ( .A(x[297]), .B(y[297]), .Z(n913) );
  XNOR U1342 ( .A(x[299]), .B(y[299]), .Z(n912) );
  XNOR U1343 ( .A(n913), .B(n912), .Z(n914) );
  XOR U1344 ( .A(n915), .B(n914), .Z(n825) );
  XOR U1345 ( .A(n824), .B(n825), .Z(n826) );
  XNOR U1346 ( .A(n827), .B(n826), .Z(n301) );
  XOR U1347 ( .A(n302), .B(n301), .Z(n304) );
  XOR U1348 ( .A(n303), .B(n304), .Z(n426) );
  XOR U1349 ( .A(n425), .B(n426), .Z(n427) );
  XOR U1350 ( .A(n428), .B(n427), .Z(n1099) );
  XNOR U1351 ( .A(x[266]), .B(y[266]), .Z(n1243) );
  XNOR U1352 ( .A(x[65]), .B(y[65]), .Z(n1240) );
  XNOR U1353 ( .A(x[268]), .B(y[268]), .Z(n1241) );
  XOR U1354 ( .A(n1240), .B(n1241), .Z(n1242) );
  XOR U1355 ( .A(n1243), .B(n1242), .Z(n982) );
  XNOR U1356 ( .A(x[270]), .B(y[270]), .Z(n1115) );
  XNOR U1357 ( .A(x[272]), .B(y[272]), .Z(n1112) );
  XNOR U1358 ( .A(x[369]), .B(y[369]), .Z(n1113) );
  XOR U1359 ( .A(n1112), .B(n1113), .Z(n1114) );
  XOR U1360 ( .A(n1115), .B(n1114), .Z(n983) );
  XOR U1361 ( .A(n982), .B(n983), .Z(n984) );
  XNOR U1362 ( .A(x[274]), .B(y[274]), .Z(n1121) );
  XNOR U1363 ( .A(x[61]), .B(y[61]), .Z(n1118) );
  XNOR U1364 ( .A(x[276]), .B(y[276]), .Z(n1119) );
  XOR U1365 ( .A(n1118), .B(n1119), .Z(n1120) );
  XOR U1366 ( .A(n1121), .B(n1120), .Z(n985) );
  XNOR U1367 ( .A(n984), .B(n985), .Z(n1081) );
  XNOR U1368 ( .A(x[394]), .B(y[394]), .Z(n537) );
  XOR U1369 ( .A(x[396]), .B(y[396]), .Z(n535) );
  XNOR U1370 ( .A(oglobal[0]), .B(n535), .Z(n536) );
  XOR U1371 ( .A(n537), .B(n536), .Z(n1004) );
  XNOR U1372 ( .A(x[286]), .B(y[286]), .Z(n1139) );
  XNOR U1373 ( .A(x[288]), .B(y[288]), .Z(n1137) );
  XNOR U1374 ( .A(x[373]), .B(y[373]), .Z(n1136) );
  XOR U1375 ( .A(n1137), .B(n1136), .Z(n1138) );
  XOR U1376 ( .A(n1139), .B(n1138), .Z(n1005) );
  XNOR U1377 ( .A(n1004), .B(n1005), .Z(n1006) );
  XNOR U1378 ( .A(x[290]), .B(y[290]), .Z(n1301) );
  XNOR U1379 ( .A(x[53]), .B(y[53]), .Z(n1299) );
  XNOR U1380 ( .A(x[292]), .B(y[292]), .Z(n1298) );
  XOR U1381 ( .A(n1299), .B(n1298), .Z(n1300) );
  XOR U1382 ( .A(n1301), .B(n1300), .Z(n1007) );
  XNOR U1383 ( .A(n1006), .B(n1007), .Z(n1078) );
  XNOR U1384 ( .A(x[278]), .B(y[278]), .Z(n1311) );
  XNOR U1385 ( .A(x[280]), .B(y[280]), .Z(n1309) );
  XNOR U1386 ( .A(x[371]), .B(y[371]), .Z(n1308) );
  XOR U1387 ( .A(n1309), .B(n1308), .Z(n1310) );
  XOR U1388 ( .A(n1311), .B(n1310), .Z(n1000) );
  XNOR U1389 ( .A(x[194]), .B(y[194]), .Z(n476) );
  XNOR U1390 ( .A(x[196]), .B(y[196]), .Z(n474) );
  XNOR U1391 ( .A(x[398]), .B(y[398]), .Z(n473) );
  XOR U1392 ( .A(n474), .B(n473), .Z(n475) );
  XOR U1393 ( .A(n476), .B(n475), .Z(n1001) );
  XOR U1394 ( .A(n1000), .B(n1001), .Z(n1002) );
  XNOR U1395 ( .A(x[282]), .B(y[282]), .Z(n1325) );
  XNOR U1396 ( .A(x[57]), .B(y[57]), .Z(n1323) );
  XNOR U1397 ( .A(x[284]), .B(y[284]), .Z(n1322) );
  XOR U1398 ( .A(n1323), .B(n1322), .Z(n1324) );
  XOR U1399 ( .A(n1325), .B(n1324), .Z(n1003) );
  XNOR U1400 ( .A(n1002), .B(n1003), .Z(n1079) );
  XOR U1401 ( .A(n1078), .B(n1079), .Z(n1080) );
  XNOR U1402 ( .A(n1081), .B(n1080), .Z(n432) );
  XNOR U1403 ( .A(x[190]), .B(y[190]), .Z(n775) );
  XNOR U1404 ( .A(x[101]), .B(y[101]), .Z(n772) );
  XNOR U1405 ( .A(x[192]), .B(y[192]), .Z(n773) );
  XOR U1406 ( .A(n772), .B(n773), .Z(n774) );
  XOR U1407 ( .A(n775), .B(n774), .Z(n990) );
  XNOR U1408 ( .A(x[198]), .B(y[198]), .Z(n781) );
  XNOR U1409 ( .A(x[200]), .B(y[200]), .Z(n778) );
  XNOR U1410 ( .A(x[351]), .B(y[351]), .Z(n779) );
  XOR U1411 ( .A(n778), .B(n779), .Z(n780) );
  XOR U1412 ( .A(n781), .B(n780), .Z(n991) );
  XOR U1413 ( .A(n990), .B(n991), .Z(n992) );
  XNOR U1414 ( .A(x[202]), .B(y[202]), .Z(n729) );
  XNOR U1415 ( .A(x[97]), .B(y[97]), .Z(n726) );
  XNOR U1416 ( .A(x[204]), .B(y[204]), .Z(n727) );
  XOR U1417 ( .A(n726), .B(n727), .Z(n728) );
  XOR U1418 ( .A(n729), .B(n728), .Z(n993) );
  XNOR U1419 ( .A(n992), .B(n993), .Z(n1255) );
  XNOR U1420 ( .A(x[206]), .B(y[206]), .Z(n460) );
  XNOR U1421 ( .A(x[208]), .B(y[208]), .Z(n458) );
  XNOR U1422 ( .A(x[353]), .B(y[353]), .Z(n457) );
  XOR U1423 ( .A(n458), .B(n457), .Z(n459) );
  XOR U1424 ( .A(n460), .B(n459), .Z(n974) );
  XNOR U1425 ( .A(x[210]), .B(y[210]), .Z(n677) );
  XNOR U1426 ( .A(x[93]), .B(y[93]), .Z(n675) );
  XNOR U1427 ( .A(x[212]), .B(y[212]), .Z(n674) );
  XOR U1428 ( .A(n675), .B(n674), .Z(n676) );
  XOR U1429 ( .A(n677), .B(n676), .Z(n975) );
  XOR U1430 ( .A(n974), .B(n975), .Z(n976) );
  XNOR U1431 ( .A(x[214]), .B(y[214]), .Z(n456) );
  XNOR U1432 ( .A(x[216]), .B(y[216]), .Z(n454) );
  XNOR U1433 ( .A(x[355]), .B(y[355]), .Z(n453) );
  XOR U1434 ( .A(n454), .B(n453), .Z(n455) );
  XOR U1435 ( .A(n456), .B(n455), .Z(n977) );
  XNOR U1436 ( .A(n976), .B(n977), .Z(n1252) );
  XNOR U1437 ( .A(x[218]), .B(y[218]), .Z(n953) );
  XNOR U1438 ( .A(x[89]), .B(y[89]), .Z(n951) );
  XNOR U1439 ( .A(x[220]), .B(y[220]), .Z(n950) );
  XOR U1440 ( .A(n951), .B(n950), .Z(n952) );
  XOR U1441 ( .A(n953), .B(n952), .Z(n978) );
  XNOR U1442 ( .A(x[222]), .B(y[222]), .Z(n484) );
  XNOR U1443 ( .A(x[224]), .B(y[224]), .Z(n482) );
  XNOR U1444 ( .A(x[357]), .B(y[357]), .Z(n481) );
  XOR U1445 ( .A(n482), .B(n481), .Z(n483) );
  XOR U1446 ( .A(n484), .B(n483), .Z(n979) );
  XOR U1447 ( .A(n978), .B(n979), .Z(n980) );
  XNOR U1448 ( .A(x[226]), .B(y[226]), .Z(n480) );
  XNOR U1449 ( .A(x[85]), .B(y[85]), .Z(n478) );
  XNOR U1450 ( .A(x[228]), .B(y[228]), .Z(n477) );
  XOR U1451 ( .A(n478), .B(n477), .Z(n479) );
  XOR U1452 ( .A(n480), .B(n479), .Z(n981) );
  XNOR U1453 ( .A(n980), .B(n981), .Z(n1253) );
  XOR U1454 ( .A(n1252), .B(n1253), .Z(n1254) );
  XNOR U1455 ( .A(n1255), .B(n1254), .Z(n430) );
  XNOR U1456 ( .A(x[230]), .B(y[230]), .Z(n1201) );
  XNOR U1457 ( .A(x[232]), .B(y[232]), .Z(n1199) );
  XNOR U1458 ( .A(x[359]), .B(y[359]), .Z(n1198) );
  XNOR U1459 ( .A(n1199), .B(n1198), .Z(n1200) );
  XNOR U1460 ( .A(n1201), .B(n1200), .Z(n1015) );
  XNOR U1461 ( .A(x[234]), .B(y[234]), .Z(n1207) );
  XNOR U1462 ( .A(x[81]), .B(y[81]), .Z(n1205) );
  XNOR U1463 ( .A(x[236]), .B(y[236]), .Z(n1204) );
  XNOR U1464 ( .A(n1205), .B(n1204), .Z(n1206) );
  XNOR U1465 ( .A(n1207), .B(n1206), .Z(n1014) );
  XOR U1466 ( .A(n1015), .B(n1014), .Z(n1016) );
  XNOR U1467 ( .A(x[238]), .B(y[238]), .Z(n326) );
  XNOR U1468 ( .A(x[240]), .B(y[240]), .Z(n324) );
  XNOR U1469 ( .A(x[361]), .B(y[361]), .Z(n323) );
  XNOR U1470 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U1471 ( .A(n326), .B(n325), .Z(n1017) );
  XNOR U1472 ( .A(n1016), .B(n1017), .Z(n901) );
  XNOR U1473 ( .A(x[250]), .B(y[250]), .Z(n366) );
  XNOR U1474 ( .A(x[73]), .B(y[73]), .Z(n364) );
  XNOR U1475 ( .A(x[252]), .B(y[252]), .Z(n363) );
  XNOR U1476 ( .A(n364), .B(n363), .Z(n365) );
  XNOR U1477 ( .A(n366), .B(n365), .Z(n1027) );
  XNOR U1478 ( .A(x[246]), .B(y[246]), .Z(n360) );
  XNOR U1479 ( .A(x[248]), .B(y[248]), .Z(n358) );
  XNOR U1480 ( .A(x[363]), .B(y[363]), .Z(n357) );
  XNOR U1481 ( .A(n358), .B(n357), .Z(n359) );
  XNOR U1482 ( .A(n360), .B(n359), .Z(n1024) );
  XNOR U1483 ( .A(x[242]), .B(y[242]), .Z(n332) );
  XNOR U1484 ( .A(x[77]), .B(y[77]), .Z(n330) );
  XNOR U1485 ( .A(x[244]), .B(y[244]), .Z(n329) );
  XNOR U1486 ( .A(n330), .B(n329), .Z(n331) );
  XOR U1487 ( .A(n332), .B(n331), .Z(n1025) );
  XOR U1488 ( .A(n1024), .B(n1025), .Z(n1026) );
  XNOR U1489 ( .A(n1027), .B(n1026), .Z(n900) );
  XOR U1490 ( .A(n901), .B(n900), .Z(n903) );
  XNOR U1491 ( .A(x[262]), .B(y[262]), .Z(n1237) );
  XNOR U1492 ( .A(x[264]), .B(y[264]), .Z(n1235) );
  XNOR U1493 ( .A(x[367]), .B(y[367]), .Z(n1234) );
  XNOR U1494 ( .A(n1235), .B(n1234), .Z(n1236) );
  XNOR U1495 ( .A(n1237), .B(n1236), .Z(n1023) );
  XNOR U1496 ( .A(x[258]), .B(y[258]), .Z(n410) );
  XNOR U1497 ( .A(x[69]), .B(y[69]), .Z(n408) );
  XNOR U1498 ( .A(x[260]), .B(y[260]), .Z(n407) );
  XNOR U1499 ( .A(n408), .B(n407), .Z(n409) );
  XNOR U1500 ( .A(n410), .B(n409), .Z(n1020) );
  XNOR U1501 ( .A(x[254]), .B(y[254]), .Z(n404) );
  XNOR U1502 ( .A(x[256]), .B(y[256]), .Z(n402) );
  XNOR U1503 ( .A(x[365]), .B(y[365]), .Z(n401) );
  XNOR U1504 ( .A(n402), .B(n401), .Z(n403) );
  XOR U1505 ( .A(n404), .B(n403), .Z(n1021) );
  XOR U1506 ( .A(n1020), .B(n1021), .Z(n1022) );
  XNOR U1507 ( .A(n1023), .B(n1022), .Z(n902) );
  XNOR U1508 ( .A(n903), .B(n902), .Z(n429) );
  XOR U1509 ( .A(n430), .B(n429), .Z(n431) );
  XNOR U1510 ( .A(n432), .B(n431), .Z(n1097) );
  XNOR U1511 ( .A(x[142]), .B(y[142]), .Z(n639) );
  XNOR U1512 ( .A(x[125]), .B(y[125]), .Z(n637) );
  XNOR U1513 ( .A(x[144]), .B(y[144]), .Z(n636) );
  XNOR U1514 ( .A(n637), .B(n636), .Z(n638) );
  XNOR U1515 ( .A(n639), .B(n638), .Z(n1035) );
  XNOR U1516 ( .A(x[146]), .B(y[146]), .Z(n506) );
  XNOR U1517 ( .A(x[148]), .B(y[148]), .Z(n504) );
  XNOR U1518 ( .A(x[339]), .B(y[339]), .Z(n503) );
  XNOR U1519 ( .A(n504), .B(n503), .Z(n505) );
  XNOR U1520 ( .A(n506), .B(n505), .Z(n1034) );
  XOR U1521 ( .A(n1035), .B(n1034), .Z(n1036) );
  XNOR U1522 ( .A(x[150]), .B(y[150]), .Z(n500) );
  XNOR U1523 ( .A(x[121]), .B(y[121]), .Z(n498) );
  XNOR U1524 ( .A(x[152]), .B(y[152]), .Z(n497) );
  XNOR U1525 ( .A(n498), .B(n497), .Z(n499) );
  XNOR U1526 ( .A(n500), .B(n499), .Z(n1037) );
  XOR U1527 ( .A(n1036), .B(n1037), .Z(n1217) );
  XNOR U1528 ( .A(x[138]), .B(y[138]), .Z(n633) );
  XNOR U1529 ( .A(x[140]), .B(y[140]), .Z(n631) );
  XNOR U1530 ( .A(x[337]), .B(y[337]), .Z(n630) );
  XNOR U1531 ( .A(n631), .B(n630), .Z(n632) );
  XNOR U1532 ( .A(n633), .B(n632), .Z(n1050) );
  XNOR U1533 ( .A(x[134]), .B(y[134]), .Z(n821) );
  XNOR U1534 ( .A(x[129]), .B(y[129]), .Z(n819) );
  XNOR U1535 ( .A(x[136]), .B(y[136]), .Z(n818) );
  XNOR U1536 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U1537 ( .A(n821), .B(n820), .Z(n1048) );
  XNOR U1538 ( .A(x[130]), .B(y[130]), .Z(n815) );
  XNOR U1539 ( .A(x[132]), .B(y[132]), .Z(n813) );
  XNOR U1540 ( .A(x[335]), .B(y[335]), .Z(n812) );
  XNOR U1541 ( .A(n813), .B(n812), .Z(n814) );
  XOR U1542 ( .A(n815), .B(n814), .Z(n1049) );
  XOR U1543 ( .A(n1048), .B(n1049), .Z(n1051) );
  XNOR U1544 ( .A(n1050), .B(n1051), .Z(n1216) );
  XNOR U1545 ( .A(n1217), .B(n1216), .Z(n1219) );
  XNOR U1546 ( .A(x[126]), .B(y[126]), .Z(n839) );
  XNOR U1547 ( .A(x[128]), .B(y[128]), .Z(n837) );
  XNOR U1548 ( .A(x[133]), .B(y[133]), .Z(n836) );
  XOR U1549 ( .A(n837), .B(n836), .Z(n838) );
  XOR U1550 ( .A(n839), .B(n838), .Z(n921) );
  XNOR U1551 ( .A(x[120]), .B(y[120]), .Z(n835) );
  XNOR U1552 ( .A(x[122]), .B(y[122]), .Z(n833) );
  XNOR U1553 ( .A(x[124]), .B(y[124]), .Z(n832) );
  XOR U1554 ( .A(n833), .B(n832), .Z(n834) );
  XOR U1555 ( .A(n835), .B(n834), .Z(n918) );
  XNOR U1556 ( .A(x[114]), .B(y[114]), .Z(n534) );
  XNOR U1557 ( .A(x[116]), .B(y[116]), .Z(n532) );
  XNOR U1558 ( .A(x[118]), .B(y[118]), .Z(n531) );
  XOR U1559 ( .A(n532), .B(n531), .Z(n533) );
  XNOR U1560 ( .A(n534), .B(n533), .Z(n919) );
  XNOR U1561 ( .A(n918), .B(n919), .Z(n920) );
  XOR U1562 ( .A(n921), .B(n920), .Z(n1218) );
  XOR U1563 ( .A(n1219), .B(n1218), .Z(n972) );
  XNOR U1564 ( .A(x[154]), .B(y[154]), .Z(n549) );
  XNOR U1565 ( .A(x[156]), .B(y[156]), .Z(n547) );
  XNOR U1566 ( .A(x[341]), .B(y[341]), .Z(n546) );
  XOR U1567 ( .A(n547), .B(n546), .Z(n548) );
  XOR U1568 ( .A(n549), .B(n548), .Z(n1092) );
  XNOR U1569 ( .A(x[158]), .B(y[158]), .Z(n553) );
  XNOR U1570 ( .A(x[117]), .B(y[117]), .Z(n551) );
  XNOR U1571 ( .A(x[160]), .B(y[160]), .Z(n550) );
  XOR U1572 ( .A(n551), .B(n550), .Z(n552) );
  XNOR U1573 ( .A(n553), .B(n552), .Z(n1093) );
  XOR U1574 ( .A(n1092), .B(n1093), .Z(n1095) );
  XNOR U1575 ( .A(x[162]), .B(y[162]), .Z(n577) );
  XNOR U1576 ( .A(x[164]), .B(y[164]), .Z(n575) );
  XNOR U1577 ( .A(x[343]), .B(y[343]), .Z(n574) );
  XOR U1578 ( .A(n575), .B(n574), .Z(n576) );
  XNOR U1579 ( .A(n577), .B(n576), .Z(n1094) );
  XOR U1580 ( .A(n1095), .B(n1094), .Z(n384) );
  XNOR U1581 ( .A(x[178]), .B(y[178]), .Z(n1167) );
  XNOR U1582 ( .A(x[180]), .B(y[180]), .Z(n1164) );
  XNOR U1583 ( .A(x[347]), .B(y[347]), .Z(n1165) );
  XOR U1584 ( .A(n1164), .B(n1165), .Z(n1166) );
  XOR U1585 ( .A(n1167), .B(n1166), .Z(n986) );
  XNOR U1586 ( .A(x[182]), .B(y[182]), .Z(n1173) );
  XNOR U1587 ( .A(x[105]), .B(y[105]), .Z(n1170) );
  XNOR U1588 ( .A(x[184]), .B(y[184]), .Z(n1171) );
  XOR U1589 ( .A(n1170), .B(n1171), .Z(n1172) );
  XNOR U1590 ( .A(n1173), .B(n1172), .Z(n987) );
  XOR U1591 ( .A(n986), .B(n987), .Z(n989) );
  XNOR U1592 ( .A(x[186]), .B(y[186]), .Z(n735) );
  XNOR U1593 ( .A(x[188]), .B(y[188]), .Z(n732) );
  XNOR U1594 ( .A(x[349]), .B(y[349]), .Z(n733) );
  XOR U1595 ( .A(n732), .B(n733), .Z(n734) );
  XNOR U1596 ( .A(n735), .B(n734), .Z(n988) );
  XOR U1597 ( .A(n989), .B(n988), .Z(n381) );
  XNOR U1598 ( .A(x[166]), .B(y[166]), .Z(n581) );
  XNOR U1599 ( .A(x[113]), .B(y[113]), .Z(n579) );
  XNOR U1600 ( .A(x[168]), .B(y[168]), .Z(n578) );
  XOR U1601 ( .A(n579), .B(n578), .Z(n580) );
  XOR U1602 ( .A(n581), .B(n580), .Z(n1010) );
  XNOR U1603 ( .A(x[170]), .B(y[170]), .Z(n563) );
  XNOR U1604 ( .A(x[172]), .B(y[172]), .Z(n561) );
  XNOR U1605 ( .A(x[345]), .B(y[345]), .Z(n560) );
  XOR U1606 ( .A(n561), .B(n560), .Z(n562) );
  XNOR U1607 ( .A(n563), .B(n562), .Z(n1011) );
  XOR U1608 ( .A(n1010), .B(n1011), .Z(n1013) );
  XNOR U1609 ( .A(x[174]), .B(y[174]), .Z(n567) );
  XNOR U1610 ( .A(x[109]), .B(y[109]), .Z(n565) );
  XNOR U1611 ( .A(x[176]), .B(y[176]), .Z(n564) );
  XOR U1612 ( .A(n565), .B(n564), .Z(n566) );
  XNOR U1613 ( .A(n567), .B(n566), .Z(n1012) );
  XOR U1614 ( .A(n1013), .B(n1012), .Z(n382) );
  XOR U1615 ( .A(n381), .B(n382), .Z(n383) );
  XNOR U1616 ( .A(n384), .B(n383), .Z(n970) );
  XNOR U1617 ( .A(x[108]), .B(y[108]), .Z(n530) );
  XNOR U1618 ( .A(x[110]), .B(y[110]), .Z(n528) );
  XNOR U1619 ( .A(x[112]), .B(y[112]), .Z(n527) );
  XOR U1620 ( .A(n528), .B(n527), .Z(n529) );
  XOR U1621 ( .A(n530), .B(n529), .Z(n967) );
  XNOR U1622 ( .A(x[102]), .B(y[102]), .Z(n472) );
  XNOR U1623 ( .A(x[104]), .B(y[104]), .Z(n470) );
  XNOR U1624 ( .A(x[106]), .B(y[106]), .Z(n469) );
  XOR U1625 ( .A(n470), .B(n469), .Z(n471) );
  XOR U1626 ( .A(n472), .B(n471), .Z(n964) );
  XNOR U1627 ( .A(x[96]), .B(y[96]), .Z(n468) );
  XNOR U1628 ( .A(x[98]), .B(y[98]), .Z(n466) );
  XNOR U1629 ( .A(x[100]), .B(y[100]), .Z(n465) );
  XOR U1630 ( .A(n466), .B(n465), .Z(n467) );
  XNOR U1631 ( .A(n468), .B(n467), .Z(n965) );
  XNOR U1632 ( .A(n964), .B(n965), .Z(n966) );
  XNOR U1633 ( .A(n967), .B(n966), .Z(n1213) );
  XNOR U1634 ( .A(x[90]), .B(y[90]), .Z(n446) );
  XNOR U1635 ( .A(x[92]), .B(y[92]), .Z(n444) );
  XNOR U1636 ( .A(x[94]), .B(y[94]), .Z(n443) );
  XOR U1637 ( .A(n444), .B(n443), .Z(n445) );
  XOR U1638 ( .A(n446), .B(n445), .Z(n860) );
  XNOR U1639 ( .A(x[78]), .B(y[78]), .Z(n442) );
  XNOR U1640 ( .A(x[80]), .B(y[80]), .Z(n440) );
  XNOR U1641 ( .A(x[82]), .B(y[82]), .Z(n439) );
  XOR U1642 ( .A(n440), .B(n439), .Z(n441) );
  XOR U1643 ( .A(n442), .B(n441), .Z(n858) );
  XNOR U1644 ( .A(x[84]), .B(y[84]), .Z(n438) );
  XNOR U1645 ( .A(x[86]), .B(y[86]), .Z(n436) );
  XNOR U1646 ( .A(x[88]), .B(y[88]), .Z(n435) );
  XOR U1647 ( .A(n436), .B(n435), .Z(n437) );
  XNOR U1648 ( .A(n438), .B(n437), .Z(n859) );
  XOR U1649 ( .A(n860), .B(n861), .Z(n1211) );
  XNOR U1650 ( .A(x[60]), .B(y[60]), .Z(n512) );
  XNOR U1651 ( .A(x[62]), .B(y[62]), .Z(n509) );
  XNOR U1652 ( .A(x[64]), .B(y[64]), .Z(n510) );
  XOR U1653 ( .A(n509), .B(n510), .Z(n511) );
  XOR U1654 ( .A(n512), .B(n511), .Z(n347) );
  XNOR U1655 ( .A(x[72]), .B(y[72]), .Z(n518) );
  XNOR U1656 ( .A(x[74]), .B(y[74]), .Z(n515) );
  XNOR U1657 ( .A(x[76]), .B(y[76]), .Z(n516) );
  XOR U1658 ( .A(n515), .B(n516), .Z(n517) );
  XOR U1659 ( .A(n518), .B(n517), .Z(n348) );
  XOR U1660 ( .A(n347), .B(n348), .Z(n349) );
  XNOR U1661 ( .A(x[66]), .B(y[66]), .Z(n524) );
  XNOR U1662 ( .A(x[68]), .B(y[68]), .Z(n521) );
  XNOR U1663 ( .A(x[70]), .B(y[70]), .Z(n522) );
  XOR U1664 ( .A(n521), .B(n522), .Z(n523) );
  XOR U1665 ( .A(n524), .B(n523), .Z(n350) );
  XNOR U1666 ( .A(n349), .B(n350), .Z(n1210) );
  XOR U1667 ( .A(n1211), .B(n1210), .Z(n1212) );
  XOR U1668 ( .A(n1213), .B(n1212), .Z(n971) );
  XOR U1669 ( .A(n970), .B(n971), .Z(n973) );
  XNOR U1670 ( .A(n972), .B(n973), .Z(n1096) );
  XNOR U1671 ( .A(n1097), .B(n1096), .Z(n1098) );
  XOR U1672 ( .A(n1099), .B(n1098), .Z(n1345) );
  XNOR U1673 ( .A(n1344), .B(n1345), .Z(o[0]) );
  NANDN U1674 ( .A(n302), .B(n301), .Z(n306) );
  OR U1675 ( .A(n304), .B(n303), .Z(n305) );
  AND U1676 ( .A(n306), .B(n305), .Z(n1725) );
  OR U1677 ( .A(n308), .B(n307), .Z(n312) );
  NANDN U1678 ( .A(n310), .B(n309), .Z(n311) );
  AND U1679 ( .A(n312), .B(n311), .Z(n1722) );
  OR U1680 ( .A(n314), .B(n313), .Z(n318) );
  OR U1681 ( .A(n316), .B(n315), .Z(n317) );
  NAND U1682 ( .A(n318), .B(n317), .Z(n1699) );
  OR U1683 ( .A(n324), .B(n323), .Z(n328) );
  OR U1684 ( .A(n326), .B(n325), .Z(n327) );
  AND U1685 ( .A(n328), .B(n327), .Z(n1552) );
  XNOR U1686 ( .A(n1553), .B(n1552), .Z(n1554) );
  OR U1687 ( .A(n330), .B(n329), .Z(n334) );
  OR U1688 ( .A(n332), .B(n331), .Z(n333) );
  AND U1689 ( .A(n334), .B(n333), .Z(n1555) );
  XOR U1690 ( .A(n1554), .B(n1555), .Z(n1696) );
  NANDN U1691 ( .A(n336), .B(n335), .Z(n340) );
  NAND U1692 ( .A(n338), .B(n337), .Z(n339) );
  NAND U1693 ( .A(n340), .B(n339), .Z(n1697) );
  XNOR U1694 ( .A(n1696), .B(n1697), .Z(n1698) );
  XOR U1695 ( .A(n1699), .B(n1698), .Z(n1723) );
  XOR U1696 ( .A(n1722), .B(n1723), .Z(n1724) );
  XNOR U1697 ( .A(n1725), .B(n1724), .Z(n1867) );
  OR U1698 ( .A(n342), .B(n341), .Z(n346) );
  NANDN U1699 ( .A(n344), .B(n343), .Z(n345) );
  NAND U1700 ( .A(n346), .B(n345), .Z(n1681) );
  OR U1701 ( .A(n352), .B(n351), .Z(n356) );
  OR U1702 ( .A(n354), .B(n353), .Z(n355) );
  NAND U1703 ( .A(n356), .B(n355), .Z(n1587) );
  OR U1704 ( .A(n358), .B(n357), .Z(n362) );
  OR U1705 ( .A(n360), .B(n359), .Z(n361) );
  AND U1706 ( .A(n362), .B(n361), .Z(n1586) );
  OR U1707 ( .A(n364), .B(n363), .Z(n368) );
  OR U1708 ( .A(n366), .B(n365), .Z(n367) );
  AND U1709 ( .A(n368), .B(n367), .Z(n1589) );
  XOR U1710 ( .A(n1588), .B(n1589), .Z(n1616) );
  OR U1711 ( .A(n370), .B(n369), .Z(n374) );
  OR U1712 ( .A(n372), .B(n371), .Z(n373) );
  NAND U1713 ( .A(n374), .B(n373), .Z(n1617) );
  XNOR U1714 ( .A(n1616), .B(n1617), .Z(n1619) );
  XOR U1715 ( .A(n1618), .B(n1619), .Z(n1678) );
  OR U1716 ( .A(n376), .B(n375), .Z(n380) );
  NAND U1717 ( .A(n378), .B(n377), .Z(n379) );
  NAND U1718 ( .A(n380), .B(n379), .Z(n1679) );
  XNOR U1719 ( .A(n1678), .B(n1679), .Z(n1680) );
  XNOR U1720 ( .A(n1681), .B(n1680), .Z(n1865) );
  OR U1721 ( .A(n382), .B(n381), .Z(n386) );
  NANDN U1722 ( .A(n384), .B(n383), .Z(n385) );
  AND U1723 ( .A(n386), .B(n385), .Z(n1652) );
  OR U1724 ( .A(n396), .B(n395), .Z(n400) );
  OR U1725 ( .A(n398), .B(n397), .Z(n399) );
  NAND U1726 ( .A(n400), .B(n399), .Z(n1541) );
  OR U1727 ( .A(n402), .B(n401), .Z(n406) );
  OR U1728 ( .A(n404), .B(n403), .Z(n405) );
  AND U1729 ( .A(n406), .B(n405), .Z(n1540) );
  XNOR U1730 ( .A(n1541), .B(n1540), .Z(n1542) );
  OR U1731 ( .A(n408), .B(n407), .Z(n412) );
  OR U1732 ( .A(n410), .B(n409), .Z(n411) );
  NAND U1733 ( .A(n412), .B(n411), .Z(n1543) );
  XOR U1734 ( .A(n1542), .B(n1543), .Z(n1593) );
  OR U1735 ( .A(n414), .B(n413), .Z(n418) );
  OR U1736 ( .A(n416), .B(n415), .Z(n417) );
  NAND U1737 ( .A(n418), .B(n417), .Z(n1592) );
  XNOR U1738 ( .A(n1593), .B(n1592), .Z(n1595) );
  XNOR U1739 ( .A(n1594), .B(n1595), .Z(n1651) );
  XNOR U1740 ( .A(n1650), .B(n1651), .Z(n1653) );
  XNOR U1741 ( .A(n1652), .B(n1653), .Z(n1866) );
  XOR U1742 ( .A(n1865), .B(n1866), .Z(n1868) );
  XOR U1743 ( .A(n1867), .B(n1868), .Z(n1662) );
  OR U1744 ( .A(n420), .B(n419), .Z(n424) );
  NANDN U1745 ( .A(n422), .B(n421), .Z(n423) );
  NAND U1746 ( .A(n424), .B(n423), .Z(n1522) );
  XNOR U1747 ( .A(n1522), .B(n1523), .Z(n1524) );
  OR U1748 ( .A(n430), .B(n429), .Z(n434) );
  NANDN U1749 ( .A(n432), .B(n431), .Z(n433) );
  AND U1750 ( .A(n434), .B(n433), .Z(n1525) );
  XOR U1751 ( .A(n1524), .B(n1525), .Z(n1661) );
  XOR U1752 ( .A(n1477), .B(n1476), .Z(n1479) );
  XOR U1753 ( .A(n1479), .B(n1478), .Z(n1356) );
  OR U1754 ( .A(n448), .B(n447), .Z(n452) );
  NANDN U1755 ( .A(n450), .B(n449), .Z(n451) );
  NAND U1756 ( .A(n452), .B(n451), .Z(n1423) );
  XOR U1757 ( .A(n1423), .B(n1422), .Z(n1425) );
  XOR U1758 ( .A(n1425), .B(n1424), .Z(n1355) );
  XNOR U1759 ( .A(n1355), .B(n1354), .Z(n1357) );
  XNOR U1760 ( .A(n1356), .B(n1357), .Z(n1816) );
  XOR U1761 ( .A(n1457), .B(n1456), .Z(n1459) );
  XOR U1762 ( .A(n1459), .B(n1458), .Z(n1362) );
  XOR U1763 ( .A(n1461), .B(n1460), .Z(n1463) );
  OR U1764 ( .A(n486), .B(n485), .Z(n490) );
  NANDN U1765 ( .A(n488), .B(n487), .Z(n489) );
  NAND U1766 ( .A(n490), .B(n489), .Z(n1462) );
  XOR U1767 ( .A(n1463), .B(n1462), .Z(n1361) );
  OR U1768 ( .A(n492), .B(n491), .Z(n496) );
  OR U1769 ( .A(n494), .B(n493), .Z(n495) );
  NAND U1770 ( .A(n496), .B(n495), .Z(n1444) );
  OR U1771 ( .A(n498), .B(n497), .Z(n502) );
  OR U1772 ( .A(n500), .B(n499), .Z(n501) );
  AND U1773 ( .A(n502), .B(n501), .Z(n1442) );
  OR U1774 ( .A(n504), .B(n503), .Z(n508) );
  OR U1775 ( .A(n506), .B(n505), .Z(n507) );
  NAND U1776 ( .A(n508), .B(n507), .Z(n1443) );
  XOR U1777 ( .A(n1442), .B(n1443), .Z(n1445) );
  XNOR U1778 ( .A(n1444), .B(n1445), .Z(n1360) );
  XNOR U1779 ( .A(n1361), .B(n1360), .Z(n1363) );
  XNOR U1780 ( .A(n1362), .B(n1363), .Z(n1814) );
  OR U1781 ( .A(n510), .B(n509), .Z(n514) );
  NANDN U1782 ( .A(n512), .B(n511), .Z(n513) );
  NAND U1783 ( .A(n514), .B(n513), .Z(n1473) );
  OR U1784 ( .A(n516), .B(n515), .Z(n520) );
  NANDN U1785 ( .A(n518), .B(n517), .Z(n519) );
  NAND U1786 ( .A(n520), .B(n519), .Z(n1472) );
  XOR U1787 ( .A(n1473), .B(n1472), .Z(n1475) );
  OR U1788 ( .A(n522), .B(n521), .Z(n526) );
  NANDN U1789 ( .A(n524), .B(n523), .Z(n525) );
  NAND U1790 ( .A(n526), .B(n525), .Z(n1474) );
  XOR U1791 ( .A(n1475), .B(n1474), .Z(n1368) );
  XOR U1792 ( .A(n1403), .B(n1402), .Z(n1405) );
  NAND U1793 ( .A(n535), .B(oglobal[0]), .Z(n539) );
  OR U1794 ( .A(n537), .B(n536), .Z(n538) );
  NAND U1795 ( .A(n539), .B(n538), .Z(n1404) );
  XOR U1796 ( .A(n1405), .B(n1404), .Z(n1367) );
  NANDN U1797 ( .A(n541), .B(n540), .Z(n545) );
  NAND U1798 ( .A(n543), .B(n542), .Z(n544) );
  AND U1799 ( .A(n545), .B(n544), .Z(n1366) );
  XNOR U1800 ( .A(n1367), .B(n1366), .Z(n1369) );
  XNOR U1801 ( .A(n1368), .B(n1369), .Z(n1813) );
  XOR U1802 ( .A(n1814), .B(n1813), .Z(n1815) );
  XNOR U1803 ( .A(n1816), .B(n1815), .Z(n1531) );
  XNOR U1804 ( .A(n1770), .B(n1769), .Z(n1771) );
  OR U1805 ( .A(n555), .B(n554), .Z(n559) );
  OR U1806 ( .A(n557), .B(n556), .Z(n558) );
  AND U1807 ( .A(n559), .B(n558), .Z(n1772) );
  XOR U1808 ( .A(n1771), .B(n1772), .Z(n1381) );
  XNOR U1809 ( .A(n1790), .B(n1789), .Z(n1791) );
  OR U1810 ( .A(n569), .B(n568), .Z(n573) );
  OR U1811 ( .A(n571), .B(n570), .Z(n572) );
  AND U1812 ( .A(n573), .B(n572), .Z(n1792) );
  XOR U1813 ( .A(n1791), .B(n1792), .Z(n1378) );
  XNOR U1814 ( .A(n1836), .B(n1835), .Z(n1837) );
  OR U1815 ( .A(n583), .B(n582), .Z(n587) );
  OR U1816 ( .A(n585), .B(n584), .Z(n586) );
  AND U1817 ( .A(n587), .B(n586), .Z(n1838) );
  XOR U1818 ( .A(n1837), .B(n1838), .Z(n1379) );
  XOR U1819 ( .A(n1378), .B(n1379), .Z(n1380) );
  XNOR U1820 ( .A(n1381), .B(n1380), .Z(n1824) );
  OR U1821 ( .A(n589), .B(n588), .Z(n593) );
  OR U1822 ( .A(n591), .B(n590), .Z(n592) );
  NAND U1823 ( .A(n593), .B(n592), .Z(n1782) );
  OR U1824 ( .A(n595), .B(n594), .Z(n599) );
  OR U1825 ( .A(n597), .B(n596), .Z(n598) );
  NAND U1826 ( .A(n599), .B(n598), .Z(n1781) );
  XOR U1827 ( .A(n1782), .B(n1781), .Z(n1783) );
  OR U1828 ( .A(n601), .B(n600), .Z(n605) );
  NANDN U1829 ( .A(n603), .B(n602), .Z(n604) );
  NAND U1830 ( .A(n605), .B(n604), .Z(n1784) );
  XNOR U1831 ( .A(n1783), .B(n1784), .Z(n1483) );
  OR U1832 ( .A(n607), .B(n606), .Z(n611) );
  NANDN U1833 ( .A(n609), .B(n608), .Z(n610) );
  NAND U1834 ( .A(n611), .B(n610), .Z(n1453) );
  OR U1835 ( .A(n613), .B(n612), .Z(n617) );
  NANDN U1836 ( .A(n615), .B(n614), .Z(n616) );
  NAND U1837 ( .A(n617), .B(n616), .Z(n1452) );
  XOR U1838 ( .A(n1453), .B(n1452), .Z(n1454) );
  OR U1839 ( .A(n619), .B(n618), .Z(n623) );
  NANDN U1840 ( .A(n621), .B(n620), .Z(n622) );
  NAND U1841 ( .A(n623), .B(n622), .Z(n1455) );
  XNOR U1842 ( .A(n1454), .B(n1455), .Z(n1481) );
  OR U1843 ( .A(n625), .B(n624), .Z(n629) );
  OR U1844 ( .A(n627), .B(n626), .Z(n628) );
  NAND U1845 ( .A(n629), .B(n628), .Z(n1737) );
  OR U1846 ( .A(n631), .B(n630), .Z(n635) );
  OR U1847 ( .A(n633), .B(n632), .Z(n634) );
  NAND U1848 ( .A(n635), .B(n634), .Z(n1736) );
  XOR U1849 ( .A(n1737), .B(n1736), .Z(n1738) );
  OR U1850 ( .A(n637), .B(n636), .Z(n641) );
  OR U1851 ( .A(n639), .B(n638), .Z(n640) );
  NAND U1852 ( .A(n641), .B(n640), .Z(n1739) );
  XNOR U1853 ( .A(n1738), .B(n1739), .Z(n1480) );
  XOR U1854 ( .A(n1481), .B(n1480), .Z(n1482) );
  XNOR U1855 ( .A(n1483), .B(n1482), .Z(n1823) );
  XOR U1856 ( .A(n1824), .B(n1823), .Z(n1825) );
  NAND U1857 ( .A(n643), .B(n642), .Z(n647) );
  NAND U1858 ( .A(n645), .B(n644), .Z(n646) );
  NAND U1859 ( .A(n647), .B(n646), .Z(n1826) );
  XOR U1860 ( .A(n1825), .B(n1826), .Z(n1528) );
  OR U1861 ( .A(n649), .B(n648), .Z(n653) );
  OR U1862 ( .A(n651), .B(n650), .Z(n652) );
  NAND U1863 ( .A(n653), .B(n652), .Z(n1762) );
  OR U1864 ( .A(n655), .B(n654), .Z(n659) );
  OR U1865 ( .A(n657), .B(n656), .Z(n658) );
  NAND U1866 ( .A(n659), .B(n658), .Z(n1761) );
  XOR U1867 ( .A(n1762), .B(n1761), .Z(n1763) );
  OR U1868 ( .A(n661), .B(n660), .Z(n665) );
  OR U1869 ( .A(n663), .B(n662), .Z(n664) );
  NAND U1870 ( .A(n665), .B(n664), .Z(n1764) );
  XNOR U1871 ( .A(n1763), .B(n1764), .Z(n1501) );
  XNOR U1872 ( .A(n1535), .B(n1534), .Z(n1536) );
  XOR U1873 ( .A(n1536), .B(n1537), .Z(n1498) );
  XOR U1874 ( .A(n1597), .B(n1596), .Z(n1598) );
  XNOR U1875 ( .A(n1598), .B(n1599), .Z(n1499) );
  XNOR U1876 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U1877 ( .A(n1501), .B(n1500), .Z(n1639) );
  OR U1878 ( .A(n691), .B(n690), .Z(n695) );
  OR U1879 ( .A(n693), .B(n692), .Z(n694) );
  NAND U1880 ( .A(n695), .B(n694), .Z(n1786) );
  OR U1881 ( .A(n697), .B(n696), .Z(n701) );
  OR U1882 ( .A(n699), .B(n698), .Z(n700) );
  NAND U1883 ( .A(n701), .B(n700), .Z(n1785) );
  XOR U1884 ( .A(n1786), .B(n1785), .Z(n1787) );
  OR U1885 ( .A(n703), .B(n702), .Z(n707) );
  OR U1886 ( .A(n705), .B(n704), .Z(n706) );
  NAND U1887 ( .A(n707), .B(n706), .Z(n1788) );
  XNOR U1888 ( .A(n1787), .B(n1788), .Z(n1519) );
  OR U1889 ( .A(n713), .B(n712), .Z(n717) );
  OR U1890 ( .A(n715), .B(n714), .Z(n716) );
  NAND U1891 ( .A(n717), .B(n716), .Z(n1732) );
  XOR U1892 ( .A(n1733), .B(n1732), .Z(n1734) );
  XNOR U1893 ( .A(n1734), .B(n1735), .Z(n1517) );
  OR U1894 ( .A(n727), .B(n726), .Z(n731) );
  NANDN U1895 ( .A(n729), .B(n728), .Z(n730) );
  AND U1896 ( .A(n731), .B(n730), .Z(n1546) );
  XNOR U1897 ( .A(n1547), .B(n1546), .Z(n1548) );
  OR U1898 ( .A(n733), .B(n732), .Z(n737) );
  NANDN U1899 ( .A(n735), .B(n734), .Z(n736) );
  NAND U1900 ( .A(n737), .B(n736), .Z(n1549) );
  XNOR U1901 ( .A(n1548), .B(n1549), .Z(n1516) );
  XOR U1902 ( .A(n1517), .B(n1516), .Z(n1518) );
  XNOR U1903 ( .A(n1519), .B(n1518), .Z(n1638) );
  XNOR U1904 ( .A(n1639), .B(n1638), .Z(n1641) );
  XOR U1905 ( .A(n1766), .B(n1765), .Z(n1767) );
  OR U1906 ( .A(n747), .B(n746), .Z(n751) );
  OR U1907 ( .A(n749), .B(n748), .Z(n750) );
  NAND U1908 ( .A(n751), .B(n750), .Z(n1768) );
  XNOR U1909 ( .A(n1767), .B(n1768), .Z(n1507) );
  OR U1910 ( .A(n753), .B(n752), .Z(n757) );
  NANDN U1911 ( .A(n755), .B(n754), .Z(n756) );
  NAND U1912 ( .A(n757), .B(n756), .Z(n1601) );
  OR U1913 ( .A(n759), .B(n758), .Z(n763) );
  NANDN U1914 ( .A(n761), .B(n760), .Z(n762) );
  NAND U1915 ( .A(n763), .B(n762), .Z(n1600) );
  XOR U1916 ( .A(n1601), .B(n1600), .Z(n1602) );
  XNOR U1917 ( .A(n1602), .B(n1603), .Z(n1505) );
  OR U1918 ( .A(n773), .B(n772), .Z(n777) );
  NANDN U1919 ( .A(n775), .B(n774), .Z(n776) );
  NAND U1920 ( .A(n777), .B(n776), .Z(n1576) );
  XOR U1921 ( .A(n1577), .B(n1576), .Z(n1578) );
  OR U1922 ( .A(n779), .B(n778), .Z(n783) );
  NANDN U1923 ( .A(n781), .B(n780), .Z(n782) );
  NAND U1924 ( .A(n783), .B(n782), .Z(n1579) );
  XNOR U1925 ( .A(n1578), .B(n1579), .Z(n1504) );
  XOR U1926 ( .A(n1505), .B(n1504), .Z(n1506) );
  XNOR U1927 ( .A(n1507), .B(n1506), .Z(n1640) );
  XOR U1928 ( .A(n1641), .B(n1640), .Z(n1529) );
  XNOR U1929 ( .A(n1528), .B(n1529), .Z(n1530) );
  XNOR U1930 ( .A(n1531), .B(n1530), .Z(n1660) );
  XOR U1931 ( .A(n1661), .B(n1660), .Z(n1663) );
  XNOR U1932 ( .A(n1662), .B(n1663), .Z(n1351) );
  NAND U1933 ( .A(n785), .B(n784), .Z(n789) );
  NAND U1934 ( .A(n787), .B(n786), .Z(n788) );
  NAND U1935 ( .A(n789), .B(n788), .Z(n1669) );
  OR U1936 ( .A(n791), .B(n790), .Z(n795) );
  NANDN U1937 ( .A(n793), .B(n792), .Z(n794) );
  NAND U1938 ( .A(n795), .B(n794), .Z(n1854) );
  OR U1939 ( .A(n797), .B(n796), .Z(n801) );
  NANDN U1940 ( .A(n799), .B(n798), .Z(n800) );
  NAND U1941 ( .A(n801), .B(n800), .Z(n1853) );
  XOR U1942 ( .A(n1854), .B(n1853), .Z(n1856) );
  OR U1943 ( .A(n803), .B(n802), .Z(n807) );
  NANDN U1944 ( .A(n805), .B(n804), .Z(n806) );
  AND U1945 ( .A(n807), .B(n806), .Z(n1855) );
  XOR U1946 ( .A(n1856), .B(n1855), .Z(n1494) );
  OR U1947 ( .A(n813), .B(n812), .Z(n817) );
  OR U1948 ( .A(n815), .B(n814), .Z(n816) );
  NAND U1949 ( .A(n817), .B(n816), .Z(n1740) );
  XOR U1950 ( .A(n1741), .B(n1740), .Z(n1743) );
  OR U1951 ( .A(n819), .B(n818), .Z(n823) );
  OR U1952 ( .A(n821), .B(n820), .Z(n822) );
  AND U1953 ( .A(n823), .B(n822), .Z(n1742) );
  XOR U1954 ( .A(n1743), .B(n1742), .Z(n1492) );
  XNOR U1955 ( .A(n1492), .B(n1493), .Z(n1495) );
  XNOR U1956 ( .A(n1494), .B(n1495), .Z(n1802) );
  XOR U1957 ( .A(n1407), .B(n1406), .Z(n1409) );
  XOR U1958 ( .A(n1409), .B(n1408), .Z(n1488) );
  OR U1959 ( .A(n841), .B(n840), .Z(n845) );
  NANDN U1960 ( .A(n843), .B(n842), .Z(n844) );
  NAND U1961 ( .A(n845), .B(n844), .Z(n1862) );
  OR U1962 ( .A(n847), .B(n846), .Z(n851) );
  NANDN U1963 ( .A(n849), .B(n848), .Z(n850) );
  NAND U1964 ( .A(n851), .B(n850), .Z(n1861) );
  XOR U1965 ( .A(n1862), .B(n1861), .Z(n1864) );
  OR U1966 ( .A(n853), .B(n852), .Z(n857) );
  NANDN U1967 ( .A(n855), .B(n854), .Z(n856) );
  AND U1968 ( .A(n857), .B(n856), .Z(n1863) );
  XOR U1969 ( .A(n1864), .B(n1863), .Z(n1486) );
  NANDN U1970 ( .A(n859), .B(n858), .Z(n863) );
  NANDN U1971 ( .A(n861), .B(n860), .Z(n862) );
  NAND U1972 ( .A(n863), .B(n862), .Z(n1487) );
  XNOR U1973 ( .A(n1486), .B(n1487), .Z(n1489) );
  XNOR U1974 ( .A(n1488), .B(n1489), .Z(n1801) );
  XOR U1975 ( .A(n1802), .B(n1801), .Z(n1803) );
  OR U1976 ( .A(n865), .B(n864), .Z(n869) );
  NANDN U1977 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1978 ( .A(n869), .B(n868), .Z(n1465) );
  OR U1979 ( .A(n871), .B(n870), .Z(n875) );
  NANDN U1980 ( .A(n873), .B(n872), .Z(n874) );
  NAND U1981 ( .A(n875), .B(n874), .Z(n1464) );
  XOR U1982 ( .A(n1465), .B(n1464), .Z(n1467) );
  OR U1983 ( .A(n877), .B(n876), .Z(n881) );
  NANDN U1984 ( .A(n879), .B(n878), .Z(n880) );
  AND U1985 ( .A(n881), .B(n880), .Z(n1466) );
  XOR U1986 ( .A(n1467), .B(n1466), .Z(n1512) );
  XOR U1987 ( .A(n1858), .B(n1857), .Z(n1860) );
  XOR U1988 ( .A(n1860), .B(n1859), .Z(n1510) );
  NANDN U1989 ( .A(n895), .B(n894), .Z(n899) );
  NAND U1990 ( .A(n897), .B(n896), .Z(n898) );
  NAND U1991 ( .A(n899), .B(n898), .Z(n1511) );
  XNOR U1992 ( .A(n1510), .B(n1511), .Z(n1513) );
  XNOR U1993 ( .A(n1512), .B(n1513), .Z(n1804) );
  XNOR U1994 ( .A(n1803), .B(n1804), .Z(n1667) );
  NANDN U1995 ( .A(n901), .B(n900), .Z(n905) );
  NANDN U1996 ( .A(n903), .B(n902), .Z(n904) );
  NAND U1997 ( .A(n905), .B(n904), .Z(n1657) );
  OR U1998 ( .A(n907), .B(n906), .Z(n911) );
  OR U1999 ( .A(n909), .B(n908), .Z(n910) );
  NAND U2000 ( .A(n911), .B(n910), .Z(n1744) );
  XOR U2001 ( .A(oglobal[1]), .B(n1744), .Z(n1745) );
  OR U2002 ( .A(n913), .B(n912), .Z(n917) );
  OR U2003 ( .A(n915), .B(n914), .Z(n916) );
  NAND U2004 ( .A(n917), .B(n916), .Z(n1746) );
  XOR U2005 ( .A(n1745), .B(n1746), .Z(n1384) );
  NANDN U2006 ( .A(n919), .B(n918), .Z(n923) );
  NAND U2007 ( .A(n921), .B(n920), .Z(n922) );
  NAND U2008 ( .A(n923), .B(n922), .Z(n1385) );
  XNOR U2009 ( .A(n1384), .B(n1385), .Z(n1386) );
  OR U2010 ( .A(n929), .B(n928), .Z(n933) );
  OR U2011 ( .A(n931), .B(n930), .Z(n932) );
  NAND U2012 ( .A(n933), .B(n932), .Z(n1749) );
  XOR U2013 ( .A(n1751), .B(n1752), .Z(n1387) );
  XNOR U2014 ( .A(n1386), .B(n1387), .Z(n1655) );
  XNOR U2015 ( .A(n1581), .B(n1580), .Z(n1582) );
  XOR U2016 ( .A(n1582), .B(n1583), .Z(n1375) );
  XNOR U2017 ( .A(n1848), .B(n1847), .Z(n1849) );
  OR U2018 ( .A(n959), .B(n958), .Z(n963) );
  NANDN U2019 ( .A(n961), .B(n960), .Z(n962) );
  NAND U2020 ( .A(n963), .B(n962), .Z(n1850) );
  XOR U2021 ( .A(n1849), .B(n1850), .Z(n1372) );
  NANDN U2022 ( .A(n965), .B(n964), .Z(n969) );
  NAND U2023 ( .A(n967), .B(n966), .Z(n968) );
  NAND U2024 ( .A(n969), .B(n968), .Z(n1373) );
  XNOR U2025 ( .A(n1372), .B(n1373), .Z(n1374) );
  XOR U2026 ( .A(n1375), .B(n1374), .Z(n1654) );
  XOR U2027 ( .A(n1657), .B(n1656), .Z(n1666) );
  XNOR U2028 ( .A(n1667), .B(n1666), .Z(n1668) );
  XNOR U2029 ( .A(n1669), .B(n1668), .Z(n1797) );
  XNOR U2030 ( .A(n1396), .B(n1397), .Z(n1398) );
  XOR U2031 ( .A(n1608), .B(n1609), .Z(n1611) );
  XOR U2032 ( .A(n1611), .B(n1610), .Z(n1399) );
  XOR U2033 ( .A(n1398), .B(n1399), .Z(n1629) );
  OR U2034 ( .A(n995), .B(n994), .Z(n999) );
  OR U2035 ( .A(n997), .B(n996), .Z(n998) );
  NAND U2036 ( .A(n999), .B(n998), .Z(n1626) );
  NANDN U2037 ( .A(n1005), .B(n1004), .Z(n1009) );
  NANDN U2038 ( .A(n1007), .B(n1006), .Z(n1008) );
  NAND U2039 ( .A(n1009), .B(n1008), .Z(n1690) );
  XNOR U2040 ( .A(n1690), .B(n1691), .Z(n1692) );
  XOR U2041 ( .A(n1693), .B(n1692), .Z(n1627) );
  XNOR U2042 ( .A(n1626), .B(n1627), .Z(n1628) );
  XOR U2043 ( .A(n1629), .B(n1628), .Z(n1675) );
  OR U2044 ( .A(n1015), .B(n1014), .Z(n1019) );
  NANDN U2045 ( .A(n1017), .B(n1016), .Z(n1018) );
  AND U2046 ( .A(n1019), .B(n1018), .Z(n1612) );
  XOR U2047 ( .A(n1612), .B(n1613), .Z(n1614) );
  XNOR U2048 ( .A(n1614), .B(n1615), .Z(n1809) );
  OR U2049 ( .A(n1029), .B(n1028), .Z(n1033) );
  NANDN U2050 ( .A(n1031), .B(n1030), .Z(n1032) );
  NAND U2051 ( .A(n1033), .B(n1032), .Z(n1704) );
  OR U2052 ( .A(n1035), .B(n1034), .Z(n1039) );
  NANDN U2053 ( .A(n1037), .B(n1036), .Z(n1038) );
  NAND U2054 ( .A(n1039), .B(n1038), .Z(n1703) );
  XOR U2055 ( .A(n1703), .B(n1702), .Z(n1705) );
  XOR U2056 ( .A(n1704), .B(n1705), .Z(n1808) );
  NANDN U2057 ( .A(n1049), .B(n1048), .Z(n1053) );
  NANDN U2058 ( .A(n1051), .B(n1050), .Z(n1052) );
  NAND U2059 ( .A(n1053), .B(n1052), .Z(n1713) );
  OR U2060 ( .A(n1055), .B(n1054), .Z(n1059) );
  NANDN U2061 ( .A(n1057), .B(n1056), .Z(n1058) );
  NAND U2062 ( .A(n1059), .B(n1058), .Z(n1469) );
  OR U2063 ( .A(n1061), .B(n1060), .Z(n1065) );
  NANDN U2064 ( .A(n1063), .B(n1062), .Z(n1064) );
  NAND U2065 ( .A(n1065), .B(n1064), .Z(n1468) );
  XOR U2066 ( .A(n1469), .B(n1468), .Z(n1471) );
  OR U2067 ( .A(n1067), .B(n1066), .Z(n1071) );
  NANDN U2068 ( .A(n1069), .B(n1068), .Z(n1070) );
  NAND U2069 ( .A(n1071), .B(n1070), .Z(n1470) );
  XOR U2070 ( .A(n1471), .B(n1470), .Z(n1712) );
  XOR U2071 ( .A(n1713), .B(n1712), .Z(n1715) );
  XNOR U2072 ( .A(n1714), .B(n1715), .Z(n1807) );
  XNOR U2073 ( .A(n1808), .B(n1807), .Z(n1810) );
  XOR U2074 ( .A(n1809), .B(n1810), .Z(n1672) );
  NAND U2075 ( .A(n1073), .B(n1072), .Z(n1077) );
  NANDN U2076 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U2077 ( .A(n1077), .B(n1076), .Z(n1647) );
  OR U2078 ( .A(n1079), .B(n1078), .Z(n1083) );
  NANDN U2079 ( .A(n1081), .B(n1080), .Z(n1082) );
  NAND U2080 ( .A(n1083), .B(n1082), .Z(n1644) );
  XNOR U2081 ( .A(n1684), .B(n1685), .Z(n1686) );
  XOR U2082 ( .A(n1687), .B(n1686), .Z(n1645) );
  XNOR U2083 ( .A(n1644), .B(n1645), .Z(n1646) );
  XOR U2084 ( .A(n1647), .B(n1646), .Z(n1673) );
  XOR U2085 ( .A(n1672), .B(n1673), .Z(n1674) );
  XNOR U2086 ( .A(n1675), .B(n1674), .Z(n1795) );
  XOR U2087 ( .A(n1796), .B(n1795), .Z(n1798) );
  XNOR U2088 ( .A(n1797), .B(n1798), .Z(n1873) );
  NANDN U2089 ( .A(n1097), .B(n1096), .Z(n1101) );
  NAND U2090 ( .A(n1099), .B(n1098), .Z(n1100) );
  NAND U2091 ( .A(n1101), .B(n1100), .Z(n1871) );
  OR U2092 ( .A(n1107), .B(n1106), .Z(n1111) );
  OR U2093 ( .A(n1109), .B(n1108), .Z(n1110) );
  NAND U2094 ( .A(n1111), .B(n1110), .Z(n1427) );
  OR U2095 ( .A(n1113), .B(n1112), .Z(n1117) );
  NANDN U2096 ( .A(n1115), .B(n1114), .Z(n1116) );
  NAND U2097 ( .A(n1117), .B(n1116), .Z(n1426) );
  XOR U2098 ( .A(n1427), .B(n1426), .Z(n1428) );
  OR U2099 ( .A(n1119), .B(n1118), .Z(n1123) );
  NANDN U2100 ( .A(n1121), .B(n1120), .Z(n1122) );
  NAND U2101 ( .A(n1123), .B(n1122), .Z(n1429) );
  XNOR U2102 ( .A(n1428), .B(n1429), .Z(n1830) );
  OR U2103 ( .A(n1125), .B(n1124), .Z(n1129) );
  NANDN U2104 ( .A(n1127), .B(n1126), .Z(n1128) );
  AND U2105 ( .A(n1129), .B(n1128), .Z(n1829) );
  XOR U2106 ( .A(n1830), .B(n1829), .Z(n1831) );
  XOR U2107 ( .A(n1832), .B(n1831), .Z(n1635) );
  NANDN U2108 ( .A(n1131), .B(n1130), .Z(n1135) );
  NAND U2109 ( .A(n1133), .B(n1132), .Z(n1134) );
  NAND U2110 ( .A(n1135), .B(n1134), .Z(n1777) );
  OR U2111 ( .A(n1141), .B(n1140), .Z(n1145) );
  OR U2112 ( .A(n1143), .B(n1142), .Z(n1144) );
  AND U2113 ( .A(n1145), .B(n1144), .Z(n1416) );
  OR U2114 ( .A(n1147), .B(n1146), .Z(n1151) );
  OR U2115 ( .A(n1149), .B(n1148), .Z(n1150) );
  AND U2116 ( .A(n1151), .B(n1150), .Z(n1419) );
  XOR U2117 ( .A(n1418), .B(n1419), .Z(n1775) );
  NANDN U2118 ( .A(n1153), .B(n1152), .Z(n1157) );
  NAND U2119 ( .A(n1155), .B(n1154), .Z(n1156) );
  AND U2120 ( .A(n1157), .B(n1156), .Z(n1776) );
  XNOR U2121 ( .A(n1775), .B(n1776), .Z(n1778) );
  XNOR U2122 ( .A(n1777), .B(n1778), .Z(n1633) );
  OR U2123 ( .A(n1159), .B(n1158), .Z(n1163) );
  OR U2124 ( .A(n1161), .B(n1160), .Z(n1162) );
  NAND U2125 ( .A(n1163), .B(n1162), .Z(n1842) );
  OR U2126 ( .A(n1165), .B(n1164), .Z(n1169) );
  NANDN U2127 ( .A(n1167), .B(n1166), .Z(n1168) );
  AND U2128 ( .A(n1169), .B(n1168), .Z(n1841) );
  XNOR U2129 ( .A(n1842), .B(n1841), .Z(n1843) );
  OR U2130 ( .A(n1171), .B(n1170), .Z(n1175) );
  NANDN U2131 ( .A(n1173), .B(n1172), .Z(n1174) );
  NAND U2132 ( .A(n1175), .B(n1174), .Z(n1844) );
  XOR U2133 ( .A(n1843), .B(n1844), .Z(n1708) );
  OR U2134 ( .A(n1177), .B(n1176), .Z(n1181) );
  OR U2135 ( .A(n1179), .B(n1178), .Z(n1180) );
  NAND U2136 ( .A(n1181), .B(n1180), .Z(n1437) );
  OR U2137 ( .A(n1183), .B(n1182), .Z(n1187) );
  OR U2138 ( .A(n1185), .B(n1184), .Z(n1186) );
  AND U2139 ( .A(n1187), .B(n1186), .Z(n1436) );
  XNOR U2140 ( .A(n1437), .B(n1436), .Z(n1438) );
  XOR U2141 ( .A(n1438), .B(n1439), .Z(n1706) );
  OR U2142 ( .A(n1193), .B(n1192), .Z(n1197) );
  OR U2143 ( .A(n1195), .B(n1194), .Z(n1196) );
  NAND U2144 ( .A(n1197), .B(n1196), .Z(n1605) );
  OR U2145 ( .A(n1199), .B(n1198), .Z(n1203) );
  OR U2146 ( .A(n1201), .B(n1200), .Z(n1202) );
  NAND U2147 ( .A(n1203), .B(n1202), .Z(n1604) );
  XOR U2148 ( .A(n1605), .B(n1604), .Z(n1606) );
  OR U2149 ( .A(n1205), .B(n1204), .Z(n1209) );
  OR U2150 ( .A(n1207), .B(n1206), .Z(n1208) );
  NAND U2151 ( .A(n1209), .B(n1208), .Z(n1607) );
  XNOR U2152 ( .A(n1606), .B(n1607), .Z(n1707) );
  XOR U2153 ( .A(n1708), .B(n1709), .Z(n1632) );
  XOR U2154 ( .A(n1633), .B(n1632), .Z(n1634) );
  XOR U2155 ( .A(n1635), .B(n1634), .Z(n1393) );
  NAND U2156 ( .A(n1211), .B(n1210), .Z(n1215) );
  NAND U2157 ( .A(n1213), .B(n1212), .Z(n1214) );
  NAND U2158 ( .A(n1215), .B(n1214), .Z(n1390) );
  NAND U2159 ( .A(n1217), .B(n1216), .Z(n1221) );
  NANDN U2160 ( .A(n1219), .B(n1218), .Z(n1220) );
  NAND U2161 ( .A(n1221), .B(n1220), .Z(n1391) );
  XNOR U2162 ( .A(n1390), .B(n1391), .Z(n1392) );
  XOR U2163 ( .A(n1393), .B(n1392), .Z(n1719) );
  NANDN U2164 ( .A(n1223), .B(n1222), .Z(n1227) );
  NAND U2165 ( .A(n1225), .B(n1224), .Z(n1226) );
  NAND U2166 ( .A(n1227), .B(n1226), .Z(n1573) );
  OR U2167 ( .A(n1229), .B(n1228), .Z(n1233) );
  OR U2168 ( .A(n1231), .B(n1230), .Z(n1232) );
  NAND U2169 ( .A(n1233), .B(n1232), .Z(n1559) );
  OR U2170 ( .A(n1235), .B(n1234), .Z(n1239) );
  OR U2171 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U2172 ( .A(n1239), .B(n1238), .Z(n1558) );
  XNOR U2173 ( .A(n1559), .B(n1558), .Z(n1560) );
  OR U2174 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U2175 ( .A(n1243), .B(n1242), .Z(n1244) );
  NAND U2176 ( .A(n1245), .B(n1244), .Z(n1561) );
  XOR U2177 ( .A(n1560), .B(n1561), .Z(n1570) );
  NANDN U2178 ( .A(n1247), .B(n1246), .Z(n1251) );
  NAND U2179 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U2180 ( .A(n1251), .B(n1250), .Z(n1571) );
  XNOR U2181 ( .A(n1570), .B(n1571), .Z(n1572) );
  XNOR U2182 ( .A(n1573), .B(n1572), .Z(n1620) );
  OR U2183 ( .A(n1253), .B(n1252), .Z(n1257) );
  NANDN U2184 ( .A(n1255), .B(n1254), .Z(n1256) );
  AND U2185 ( .A(n1257), .B(n1256), .Z(n1621) );
  XNOR U2186 ( .A(n1620), .B(n1621), .Z(n1623) );
  NANDN U2187 ( .A(n1259), .B(n1258), .Z(n1263) );
  NAND U2188 ( .A(n1261), .B(n1260), .Z(n1262) );
  NAND U2189 ( .A(n1263), .B(n1262), .Z(n1413) );
  NANDN U2190 ( .A(n1265), .B(n1264), .Z(n1269) );
  NAND U2191 ( .A(n1267), .B(n1266), .Z(n1268) );
  NAND U2192 ( .A(n1269), .B(n1268), .Z(n1410) );
  OR U2193 ( .A(n1275), .B(n1274), .Z(n1279) );
  OR U2194 ( .A(n1277), .B(n1276), .Z(n1278) );
  AND U2195 ( .A(n1279), .B(n1278), .Z(n1430) );
  XNOR U2196 ( .A(n1431), .B(n1430), .Z(n1432) );
  OR U2197 ( .A(n1281), .B(n1280), .Z(n1285) );
  OR U2198 ( .A(n1283), .B(n1282), .Z(n1284) );
  NAND U2199 ( .A(n1285), .B(n1284), .Z(n1433) );
  XNOR U2200 ( .A(n1432), .B(n1433), .Z(n1411) );
  XNOR U2201 ( .A(n1410), .B(n1411), .Z(n1412) );
  XOR U2202 ( .A(n1413), .B(n1412), .Z(n1622) );
  XOR U2203 ( .A(n1623), .B(n1622), .Z(n1717) );
  OR U2204 ( .A(n1287), .B(n1286), .Z(n1291) );
  NANDN U2205 ( .A(n1289), .B(n1288), .Z(n1290) );
  NAND U2206 ( .A(n1291), .B(n1290), .Z(n1449) );
  OR U2207 ( .A(n1293), .B(n1292), .Z(n1297) );
  NANDN U2208 ( .A(n1295), .B(n1294), .Z(n1296) );
  NAND U2209 ( .A(n1297), .B(n1296), .Z(n1446) );
  OR U2210 ( .A(n1303), .B(n1302), .Z(n1307) );
  OR U2211 ( .A(n1305), .B(n1304), .Z(n1306) );
  AND U2212 ( .A(n1307), .B(n1306), .Z(n1564) );
  XNOR U2213 ( .A(n1566), .B(n1567), .Z(n1447) );
  XNOR U2214 ( .A(n1446), .B(n1447), .Z(n1448) );
  XNOR U2215 ( .A(n1449), .B(n1448), .Z(n1822) );
  OR U2216 ( .A(n1313), .B(n1312), .Z(n1317) );
  OR U2217 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U2218 ( .A(n1317), .B(n1316), .Z(n1758) );
  XOR U2219 ( .A(n1728), .B(n1729), .Z(n1755) );
  NANDN U2220 ( .A(n1331), .B(n1330), .Z(n1335) );
  NAND U2221 ( .A(n1333), .B(n1332), .Z(n1334) );
  AND U2222 ( .A(n1335), .B(n1334), .Z(n1756) );
  XNOR U2223 ( .A(n1755), .B(n1756), .Z(n1757) );
  XNOR U2224 ( .A(n1758), .B(n1757), .Z(n1819) );
  OR U2225 ( .A(n1337), .B(n1336), .Z(n1341) );
  NANDN U2226 ( .A(n1339), .B(n1338), .Z(n1340) );
  NAND U2227 ( .A(n1341), .B(n1340), .Z(n1820) );
  XOR U2228 ( .A(n1819), .B(n1820), .Z(n1821) );
  XNOR U2229 ( .A(n1822), .B(n1821), .Z(n1716) );
  XOR U2230 ( .A(n1717), .B(n1716), .Z(n1718) );
  XOR U2231 ( .A(n1719), .B(n1718), .Z(n1872) );
  XNOR U2232 ( .A(n1871), .B(n1872), .Z(n1874) );
  XNOR U2233 ( .A(n1873), .B(n1874), .Z(n1349) );
  NANDN U2234 ( .A(n1343), .B(n1342), .Z(n1347) );
  NANDN U2235 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U2236 ( .A(n1347), .B(n1346), .Z(n1348) );
  XOR U2237 ( .A(n1349), .B(n1348), .Z(n1350) );
  XNOR U2238 ( .A(n1351), .B(n1350), .Z(o[1]) );
  OR U2239 ( .A(n1349), .B(n1348), .Z(n1353) );
  NANDN U2240 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U2241 ( .A(n1353), .B(n1352), .Z(n1878) );
  NAND U2242 ( .A(n1355), .B(n1354), .Z(n1359) );
  NANDN U2243 ( .A(n1357), .B(n1356), .Z(n1358) );
  NAND U2244 ( .A(n1359), .B(n1358), .Z(n2092) );
  NAND U2245 ( .A(n1361), .B(n1360), .Z(n1365) );
  NANDN U2246 ( .A(n1363), .B(n1362), .Z(n1364) );
  NAND U2247 ( .A(n1365), .B(n1364), .Z(n2089) );
  NAND U2248 ( .A(n1367), .B(n1366), .Z(n1371) );
  NANDN U2249 ( .A(n1369), .B(n1368), .Z(n1370) );
  AND U2250 ( .A(n1371), .B(n1370), .Z(n2090) );
  XOR U2251 ( .A(n2092), .B(n2091), .Z(n2125) );
  NANDN U2252 ( .A(n1373), .B(n1372), .Z(n1377) );
  NAND U2253 ( .A(n1375), .B(n1374), .Z(n1376) );
  NAND U2254 ( .A(n1377), .B(n1376), .Z(n2102) );
  OR U2255 ( .A(n1379), .B(n1378), .Z(n1383) );
  NANDN U2256 ( .A(n1381), .B(n1380), .Z(n1382) );
  NAND U2257 ( .A(n1383), .B(n1382), .Z(n2099) );
  NANDN U2258 ( .A(n1385), .B(n1384), .Z(n1389) );
  NANDN U2259 ( .A(n1387), .B(n1386), .Z(n1388) );
  AND U2260 ( .A(n1389), .B(n1388), .Z(n2100) );
  XOR U2261 ( .A(n2102), .B(n2101), .Z(n2126) );
  XNOR U2262 ( .A(n2125), .B(n2126), .Z(n2128) );
  NANDN U2263 ( .A(n1391), .B(n1390), .Z(n1395) );
  NANDN U2264 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U2265 ( .A(n1395), .B(n1394), .Z(n2127) );
  XOR U2266 ( .A(n2128), .B(n2127), .Z(n1964) );
  NANDN U2267 ( .A(n1397), .B(n1396), .Z(n1401) );
  NANDN U2268 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U2269 ( .A(n1401), .B(n1400), .Z(n1927) );
  XOR U2270 ( .A(oglobal[2]), .B(n1999), .Z(n2000) );
  XOR U2271 ( .A(n2001), .B(n2000), .Z(n1925) );
  NANDN U2272 ( .A(n1411), .B(n1410), .Z(n1415) );
  NAND U2273 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U2274 ( .A(n1415), .B(n1414), .Z(n1926) );
  XNOR U2275 ( .A(n1925), .B(n1926), .Z(n1928) );
  XOR U2276 ( .A(n1927), .B(n1928), .Z(n2122) );
  NANDN U2277 ( .A(n1417), .B(n1416), .Z(n1421) );
  NAND U2278 ( .A(n1419), .B(n1418), .Z(n1420) );
  AND U2279 ( .A(n1421), .B(n1420), .Z(n2019) );
  XNOR U2280 ( .A(n2018), .B(n2017), .Z(n2020) );
  XNOR U2281 ( .A(n2019), .B(n2020), .Z(n1990) );
  NANDN U2282 ( .A(n1431), .B(n1430), .Z(n1435) );
  NANDN U2283 ( .A(n1433), .B(n1432), .Z(n1434) );
  AND U2284 ( .A(n1435), .B(n1434), .Z(n2048) );
  NANDN U2285 ( .A(n1437), .B(n1436), .Z(n1441) );
  NANDN U2286 ( .A(n1439), .B(n1438), .Z(n1440) );
  AND U2287 ( .A(n1441), .B(n1440), .Z(n2046) );
  XNOR U2288 ( .A(n2046), .B(n2047), .Z(n2049) );
  XNOR U2289 ( .A(n2048), .B(n2049), .Z(n1987) );
  NANDN U2290 ( .A(n1447), .B(n1446), .Z(n1451) );
  NAND U2291 ( .A(n1449), .B(n1448), .Z(n1450) );
  AND U2292 ( .A(n1451), .B(n1450), .Z(n1988) );
  XNOR U2293 ( .A(n1987), .B(n1988), .Z(n1989) );
  XOR U2294 ( .A(n1990), .B(n1989), .Z(n2120) );
  XOR U2295 ( .A(n1939), .B(n1940), .Z(n1942) );
  XOR U2296 ( .A(n1941), .B(n1942), .Z(n1931) );
  XOR U2297 ( .A(n1935), .B(n1936), .Z(n1938) );
  XOR U2298 ( .A(n1937), .B(n1938), .Z(n1929) );
  XNOR U2299 ( .A(n1929), .B(n1930), .Z(n1932) );
  XNOR U2300 ( .A(n1931), .B(n1932), .Z(n2119) );
  XNOR U2301 ( .A(n2120), .B(n2119), .Z(n2121) );
  XNOR U2302 ( .A(n2122), .B(n2121), .Z(n1963) );
  XNOR U2303 ( .A(n1964), .B(n1963), .Z(n1966) );
  OR U2304 ( .A(n1481), .B(n1480), .Z(n1485) );
  NANDN U2305 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U2306 ( .A(n1485), .B(n1484), .Z(n1906) );
  OR U2307 ( .A(n1487), .B(n1486), .Z(n1491) );
  OR U2308 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U2309 ( .A(n1491), .B(n1490), .Z(n1905) );
  XOR U2310 ( .A(n1906), .B(n1905), .Z(n1908) );
  OR U2311 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U2312 ( .A(n1495), .B(n1494), .Z(n1496) );
  NAND U2313 ( .A(n1497), .B(n1496), .Z(n1907) );
  XOR U2314 ( .A(n1908), .B(n1907), .Z(n2032) );
  NANDN U2315 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U2316 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U2317 ( .A(n1503), .B(n1502), .Z(n2030) );
  OR U2318 ( .A(n1505), .B(n1504), .Z(n1509) );
  NANDN U2319 ( .A(n1507), .B(n1506), .Z(n1508) );
  NAND U2320 ( .A(n1509), .B(n1508), .Z(n1915) );
  OR U2321 ( .A(n1511), .B(n1510), .Z(n1515) );
  OR U2322 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND U2323 ( .A(n1515), .B(n1514), .Z(n1913) );
  XOR U2324 ( .A(n1915), .B(n1913), .Z(n1917) );
  OR U2325 ( .A(n1517), .B(n1516), .Z(n1521) );
  NANDN U2326 ( .A(n1519), .B(n1518), .Z(n1520) );
  NAND U2327 ( .A(n1521), .B(n1520), .Z(n1916) );
  XOR U2328 ( .A(n1917), .B(n1916), .Z(n2031) );
  XOR U2329 ( .A(n2030), .B(n2031), .Z(n2033) );
  XNOR U2330 ( .A(n2032), .B(n2033), .Z(n1965) );
  XNOR U2331 ( .A(n1966), .B(n1965), .Z(n2110) );
  NANDN U2332 ( .A(n1523), .B(n1522), .Z(n1527) );
  NAND U2333 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U2334 ( .A(n1527), .B(n1526), .Z(n2117) );
  NANDN U2335 ( .A(n1529), .B(n1528), .Z(n1533) );
  NANDN U2336 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U2337 ( .A(n1533), .B(n1532), .Z(n2116) );
  NANDN U2338 ( .A(n1535), .B(n1534), .Z(n1539) );
  NANDN U2339 ( .A(n1537), .B(n1536), .Z(n1538) );
  AND U2340 ( .A(n1539), .B(n1538), .Z(n2042) );
  NANDN U2341 ( .A(n1541), .B(n1540), .Z(n1545) );
  NANDN U2342 ( .A(n1543), .B(n1542), .Z(n1544) );
  AND U2343 ( .A(n1545), .B(n1544), .Z(n2041) );
  NANDN U2344 ( .A(n1547), .B(n1546), .Z(n1551) );
  NANDN U2345 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U2346 ( .A(n1551), .B(n1550), .Z(n2040) );
  XNOR U2347 ( .A(n2041), .B(n2040), .Z(n2043) );
  XNOR U2348 ( .A(n2042), .B(n2043), .Z(n1978) );
  NANDN U2349 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U2350 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U2351 ( .A(n1557), .B(n1556), .Z(n2013) );
  NANDN U2352 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U2353 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U2354 ( .A(n1563), .B(n1562), .Z(n2012) );
  NANDN U2355 ( .A(n1565), .B(n1564), .Z(n1569) );
  NANDN U2356 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U2357 ( .A(n1569), .B(n1568), .Z(n2011) );
  XNOR U2358 ( .A(n2012), .B(n2011), .Z(n2014) );
  XNOR U2359 ( .A(n2013), .B(n2014), .Z(n1975) );
  NANDN U2360 ( .A(n1571), .B(n1570), .Z(n1575) );
  NANDN U2361 ( .A(n1573), .B(n1572), .Z(n1574) );
  AND U2362 ( .A(n1575), .B(n1574), .Z(n1976) );
  XNOR U2363 ( .A(n1975), .B(n1976), .Z(n1977) );
  XOR U2364 ( .A(n1978), .B(n1977), .Z(n1902) );
  NANDN U2365 ( .A(n1581), .B(n1580), .Z(n1585) );
  NANDN U2366 ( .A(n1583), .B(n1582), .Z(n1584) );
  NAND U2367 ( .A(n1585), .B(n1584), .Z(n2034) );
  NANDN U2368 ( .A(n1587), .B(n1586), .Z(n1591) );
  NAND U2369 ( .A(n1589), .B(n1588), .Z(n1590) );
  AND U2370 ( .A(n1591), .B(n1590), .Z(n2035) );
  XOR U2371 ( .A(n2037), .B(n2036), .Z(n2142) );
  XOR U2372 ( .A(n2074), .B(n2073), .Z(n2140) );
  XOR U2373 ( .A(n2139), .B(n2140), .Z(n2141) );
  XOR U2374 ( .A(n2142), .B(n2141), .Z(n1899) );
  XOR U2375 ( .A(n2129), .B(n2130), .Z(n2132) );
  XOR U2376 ( .A(n2131), .B(n2132), .Z(n1900) );
  XOR U2377 ( .A(n1899), .B(n1900), .Z(n1901) );
  XNOR U2378 ( .A(n1902), .B(n1901), .Z(n2115) );
  XOR U2379 ( .A(n2116), .B(n2115), .Z(n2118) );
  XOR U2380 ( .A(n2117), .B(n2118), .Z(n2109) );
  NAND U2381 ( .A(n1621), .B(n1620), .Z(n1625) );
  NANDN U2382 ( .A(n1623), .B(n1622), .Z(n1624) );
  NAND U2383 ( .A(n1625), .B(n1624), .Z(n1955) );
  NANDN U2384 ( .A(n1627), .B(n1626), .Z(n1631) );
  NAND U2385 ( .A(n1629), .B(n1628), .Z(n1630) );
  NAND U2386 ( .A(n1631), .B(n1630), .Z(n1954) );
  NANDN U2387 ( .A(n1633), .B(n1632), .Z(n1637) );
  OR U2388 ( .A(n1635), .B(n1634), .Z(n1636) );
  NAND U2389 ( .A(n1637), .B(n1636), .Z(n1953) );
  XOR U2390 ( .A(n1954), .B(n1953), .Z(n1956) );
  XOR U2391 ( .A(n1955), .B(n1956), .Z(n2146) );
  NAND U2392 ( .A(n1639), .B(n1638), .Z(n1643) );
  NANDN U2393 ( .A(n1641), .B(n1640), .Z(n1642) );
  NAND U2394 ( .A(n1643), .B(n1642), .Z(n1952) );
  NANDN U2395 ( .A(n1645), .B(n1644), .Z(n1649) );
  NAND U2396 ( .A(n1647), .B(n1646), .Z(n1648) );
  NAND U2397 ( .A(n1649), .B(n1648), .Z(n1950) );
  XOR U2398 ( .A(n1950), .B(n1949), .Z(n1951) );
  XOR U2399 ( .A(n1952), .B(n1951), .Z(n2143) );
  NAND U2400 ( .A(n1655), .B(n1654), .Z(n1659) );
  NANDN U2401 ( .A(n1657), .B(n1656), .Z(n1658) );
  NAND U2402 ( .A(n1659), .B(n1658), .Z(n2144) );
  XNOR U2403 ( .A(n2143), .B(n2144), .Z(n2145) );
  XOR U2404 ( .A(n2146), .B(n2145), .Z(n2112) );
  XNOR U2405 ( .A(n2111), .B(n2112), .Z(n1885) );
  NANDN U2406 ( .A(n1661), .B(n1660), .Z(n1665) );
  OR U2407 ( .A(n1663), .B(n1662), .Z(n1664) );
  NAND U2408 ( .A(n1665), .B(n1664), .Z(n1884) );
  NANDN U2409 ( .A(n1667), .B(n1666), .Z(n1671) );
  NANDN U2410 ( .A(n1669), .B(n1668), .Z(n1670) );
  AND U2411 ( .A(n1671), .B(n1670), .Z(n1921) );
  OR U2412 ( .A(n1673), .B(n1672), .Z(n1677) );
  NANDN U2413 ( .A(n1675), .B(n1674), .Z(n1676) );
  NAND U2414 ( .A(n1677), .B(n1676), .Z(n1922) );
  XOR U2415 ( .A(n1921), .B(n1922), .Z(n1924) );
  NANDN U2416 ( .A(n1679), .B(n1678), .Z(n1683) );
  NANDN U2417 ( .A(n1681), .B(n1680), .Z(n1682) );
  NAND U2418 ( .A(n1683), .B(n1682), .Z(n2084) );
  NANDN U2419 ( .A(n1685), .B(n1684), .Z(n1689) );
  NAND U2420 ( .A(n1687), .B(n1686), .Z(n1688) );
  AND U2421 ( .A(n1689), .B(n1688), .Z(n1912) );
  NANDN U2422 ( .A(n1691), .B(n1690), .Z(n1695) );
  NAND U2423 ( .A(n1693), .B(n1692), .Z(n1694) );
  AND U2424 ( .A(n1695), .B(n1694), .Z(n1909) );
  OR U2425 ( .A(n1697), .B(n1696), .Z(n1701) );
  OR U2426 ( .A(n1699), .B(n1698), .Z(n1700) );
  AND U2427 ( .A(n1701), .B(n1700), .Z(n1910) );
  XOR U2428 ( .A(n1909), .B(n1910), .Z(n1911) );
  XNOR U2429 ( .A(n1912), .B(n1911), .Z(n2083) );
  XNOR U2430 ( .A(n2084), .B(n2083), .Z(n2086) );
  NANDN U2431 ( .A(n1707), .B(n1706), .Z(n1711) );
  NANDN U2432 ( .A(n1709), .B(n1708), .Z(n1710) );
  AND U2433 ( .A(n1711), .B(n1710), .Z(n2025) );
  XNOR U2434 ( .A(n2024), .B(n2025), .Z(n2026) );
  XOR U2435 ( .A(n2026), .B(n2027), .Z(n2085) );
  XOR U2436 ( .A(n2086), .B(n2085), .Z(n1959) );
  NAND U2437 ( .A(n1717), .B(n1716), .Z(n1721) );
  NAND U2438 ( .A(n1719), .B(n1718), .Z(n1720) );
  NAND U2439 ( .A(n1721), .B(n1720), .Z(n1957) );
  NANDN U2440 ( .A(n1727), .B(n1726), .Z(n1731) );
  NAND U2441 ( .A(n1729), .B(n1728), .Z(n1730) );
  NAND U2442 ( .A(n1731), .B(n1730), .Z(n2067) );
  XOR U2443 ( .A(n2067), .B(n2068), .Z(n2098) );
  OR U2444 ( .A(oglobal[1]), .B(n1744), .Z(n1748) );
  NANDN U2445 ( .A(n1746), .B(n1745), .Z(n1747) );
  NAND U2446 ( .A(n1748), .B(n1747), .Z(n1993) );
  NANDN U2447 ( .A(n1750), .B(n1749), .Z(n1754) );
  NANDN U2448 ( .A(n1752), .B(n1751), .Z(n1753) );
  NAND U2449 ( .A(n1754), .B(n1753), .Z(n1994) );
  XNOR U2450 ( .A(n1993), .B(n1994), .Z(n1995) );
  XNOR U2451 ( .A(n1996), .B(n1995), .Z(n2095) );
  OR U2452 ( .A(n1756), .B(n1755), .Z(n1760) );
  OR U2453 ( .A(n1758), .B(n1757), .Z(n1759) );
  AND U2454 ( .A(n1760), .B(n1759), .Z(n2096) );
  XOR U2455 ( .A(n2095), .B(n2096), .Z(n2097) );
  XNOR U2456 ( .A(n2098), .B(n2097), .Z(n1893) );
  XOR U2457 ( .A(n1894), .B(n1893), .Z(n1896) );
  NANDN U2458 ( .A(n1770), .B(n1769), .Z(n1774) );
  NAND U2459 ( .A(n1772), .B(n1771), .Z(n1773) );
  AND U2460 ( .A(n1774), .B(n1773), .Z(n2054) );
  XOR U2461 ( .A(n2055), .B(n2056), .Z(n2136) );
  OR U2462 ( .A(n1776), .B(n1775), .Z(n1780) );
  NANDN U2463 ( .A(n1778), .B(n1777), .Z(n1779) );
  NAND U2464 ( .A(n1780), .B(n1779), .Z(n2133) );
  NANDN U2465 ( .A(n1790), .B(n1789), .Z(n1794) );
  NAND U2466 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2467 ( .A(n1794), .B(n1793), .Z(n2060) );
  XOR U2468 ( .A(n2062), .B(n2061), .Z(n2134) );
  XNOR U2469 ( .A(n2133), .B(n2134), .Z(n2135) );
  XOR U2470 ( .A(n2136), .B(n2135), .Z(n1895) );
  XNOR U2471 ( .A(n1896), .B(n1895), .Z(n1958) );
  XOR U2472 ( .A(n1957), .B(n1958), .Z(n1960) );
  XNOR U2473 ( .A(n1959), .B(n1960), .Z(n1923) );
  XNOR U2474 ( .A(n1924), .B(n1923), .Z(n1883) );
  XNOR U2475 ( .A(n1884), .B(n1883), .Z(n1886) );
  XOR U2476 ( .A(n1885), .B(n1886), .Z(n1877) );
  XOR U2477 ( .A(n1878), .B(n1877), .Z(n1879) );
  NANDN U2478 ( .A(n1796), .B(n1795), .Z(n1800) );
  OR U2479 ( .A(n1798), .B(n1797), .Z(n1799) );
  AND U2480 ( .A(n1800), .B(n1799), .Z(n1889) );
  OR U2481 ( .A(n1802), .B(n1801), .Z(n1806) );
  NANDN U2482 ( .A(n1804), .B(n1803), .Z(n1805) );
  NAND U2483 ( .A(n1806), .B(n1805), .Z(n1972) );
  NAND U2484 ( .A(n1808), .B(n1807), .Z(n1812) );
  OR U2485 ( .A(n1810), .B(n1809), .Z(n1811) );
  NAND U2486 ( .A(n1812), .B(n1811), .Z(n1969) );
  OR U2487 ( .A(n1814), .B(n1813), .Z(n1818) );
  NANDN U2488 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2489 ( .A(n1818), .B(n1817), .Z(n1970) );
  XNOR U2490 ( .A(n1969), .B(n1970), .Z(n1971) );
  XOR U2491 ( .A(n1972), .B(n1971), .Z(n2080) );
  OR U2492 ( .A(n1824), .B(n1823), .Z(n1828) );
  NANDN U2493 ( .A(n1826), .B(n1825), .Z(n1827) );
  NAND U2494 ( .A(n1828), .B(n1827), .Z(n2106) );
  OR U2495 ( .A(n1830), .B(n1829), .Z(n1834) );
  NAND U2496 ( .A(n1832), .B(n1831), .Z(n1833) );
  NAND U2497 ( .A(n1834), .B(n1833), .Z(n1981) );
  NANDN U2498 ( .A(n1836), .B(n1835), .Z(n1840) );
  NAND U2499 ( .A(n1838), .B(n1837), .Z(n1839) );
  AND U2500 ( .A(n1840), .B(n1839), .Z(n2007) );
  NANDN U2501 ( .A(n1842), .B(n1841), .Z(n1846) );
  NANDN U2502 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U2503 ( .A(n1846), .B(n1845), .Z(n2004) );
  NANDN U2504 ( .A(n1848), .B(n1847), .Z(n1852) );
  NANDN U2505 ( .A(n1850), .B(n1849), .Z(n1851) );
  AND U2506 ( .A(n1852), .B(n1851), .Z(n2005) );
  XOR U2507 ( .A(n2004), .B(n2005), .Z(n2006) );
  XOR U2508 ( .A(n1981), .B(n1982), .Z(n1983) );
  XOR U2509 ( .A(n1943), .B(n1944), .Z(n1945) );
  XOR U2510 ( .A(n1983), .B(n1984), .Z(n2105) );
  XOR U2511 ( .A(n2106), .B(n2105), .Z(n2108) );
  XOR U2512 ( .A(n2107), .B(n2108), .Z(n2077) );
  OR U2513 ( .A(n1866), .B(n1865), .Z(n1870) );
  NAND U2514 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U2515 ( .A(n1870), .B(n1869), .Z(n2078) );
  XNOR U2516 ( .A(n2077), .B(n2078), .Z(n2079) );
  XNOR U2517 ( .A(n2080), .B(n2079), .Z(n1890) );
  XOR U2518 ( .A(n1889), .B(n1890), .Z(n1891) );
  NAND U2519 ( .A(n1872), .B(n1871), .Z(n1876) );
  NANDN U2520 ( .A(n1874), .B(n1873), .Z(n1875) );
  NAND U2521 ( .A(n1876), .B(n1875), .Z(n1892) );
  XNOR U2522 ( .A(n1891), .B(n1892), .Z(n1880) );
  XOR U2523 ( .A(n1879), .B(n1880), .Z(o[2]) );
  OR U2524 ( .A(n1878), .B(n1877), .Z(n1882) );
  NANDN U2525 ( .A(n1880), .B(n1879), .Z(n1881) );
  AND U2526 ( .A(n1882), .B(n1881), .Z(n2265) );
  IV U2527 ( .A(n2265), .Z(n2264) );
  OR U2528 ( .A(n1884), .B(n1883), .Z(n1888) );
  NANDN U2529 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2530 ( .A(n1888), .B(n1887), .Z(n2271) );
  XOR U2531 ( .A(n2271), .B(n2272), .Z(n2273) );
  NANDN U2532 ( .A(n1894), .B(n1893), .Z(n1898) );
  NANDN U2533 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2534 ( .A(n1898), .B(n1897), .Z(n2244) );
  NAND U2535 ( .A(n1900), .B(n1899), .Z(n1904) );
  NANDN U2536 ( .A(n1902), .B(n1901), .Z(n1903) );
  NAND U2537 ( .A(n1904), .B(n1903), .Z(n2243) );
  IV U2538 ( .A(n1913), .Z(n1914) );
  NANDN U2539 ( .A(n1915), .B(n1914), .Z(n1920) );
  IV U2540 ( .A(n1916), .Z(n1918) );
  NAND U2541 ( .A(n1918), .B(n1917), .Z(n1919) );
  NAND U2542 ( .A(n1920), .B(n1919), .Z(n2199) );
  XOR U2543 ( .A(n2198), .B(n2199), .Z(n2200) );
  XNOR U2544 ( .A(n2201), .B(n2200), .Z(n2242) );
  XOR U2545 ( .A(n2243), .B(n2242), .Z(n2245) );
  XOR U2546 ( .A(n2244), .B(n2245), .Z(n2226) );
  OR U2547 ( .A(n1930), .B(n1929), .Z(n1934) );
  OR U2548 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2549 ( .A(n1934), .B(n1933), .Z(n2216) );
  OR U2550 ( .A(n1944), .B(n1943), .Z(n1948) );
  NANDN U2551 ( .A(n1946), .B(n1945), .Z(n1947) );
  NAND U2552 ( .A(n1948), .B(n1947), .Z(n2192) );
  XNOR U2553 ( .A(n2193), .B(n2192), .Z(n2194) );
  XNOR U2554 ( .A(n2195), .B(n2194), .Z(n2217) );
  XOR U2555 ( .A(n2216), .B(n2217), .Z(n2219) );
  XOR U2556 ( .A(n2218), .B(n2219), .Z(n2153) );
  XOR U2557 ( .A(n2150), .B(n2151), .Z(n2152) );
  XOR U2558 ( .A(n2153), .B(n2152), .Z(n2228) );
  XOR U2559 ( .A(n2229), .B(n2228), .Z(n2255) );
  NANDN U2560 ( .A(n1958), .B(n1957), .Z(n1962) );
  NANDN U2561 ( .A(n1960), .B(n1959), .Z(n1961) );
  AND U2562 ( .A(n1962), .B(n1961), .Z(n2253) );
  NAND U2563 ( .A(n1964), .B(n1963), .Z(n1968) );
  NANDN U2564 ( .A(n1966), .B(n1965), .Z(n1967) );
  NAND U2565 ( .A(n1968), .B(n1967), .Z(n2252) );
  XNOR U2566 ( .A(n2253), .B(n2252), .Z(n2254) );
  XNOR U2567 ( .A(n2255), .B(n2254), .Z(n2274) );
  XOR U2568 ( .A(n2273), .B(n2274), .Z(n2268) );
  NANDN U2569 ( .A(n1970), .B(n1969), .Z(n1974) );
  NANDN U2570 ( .A(n1972), .B(n1971), .Z(n1973) );
  AND U2571 ( .A(n1974), .B(n1973), .Z(n2238) );
  NANDN U2572 ( .A(n1976), .B(n1975), .Z(n1980) );
  NAND U2573 ( .A(n1978), .B(n1977), .Z(n1979) );
  NAND U2574 ( .A(n1980), .B(n1979), .Z(n2215) );
  OR U2575 ( .A(n1982), .B(n1981), .Z(n1986) );
  NANDN U2576 ( .A(n1984), .B(n1983), .Z(n1985) );
  NAND U2577 ( .A(n1986), .B(n1985), .Z(n2213) );
  NANDN U2578 ( .A(n1988), .B(n1987), .Z(n1992) );
  NAND U2579 ( .A(n1990), .B(n1989), .Z(n1991) );
  NAND U2580 ( .A(n1992), .B(n1991), .Z(n2212) );
  XOR U2581 ( .A(n2213), .B(n2212), .Z(n2214) );
  XOR U2582 ( .A(n2215), .B(n2214), .Z(n2239) );
  XOR U2583 ( .A(n2238), .B(n2239), .Z(n2240) );
  NANDN U2584 ( .A(n1994), .B(n1993), .Z(n1998) );
  NAND U2585 ( .A(n1996), .B(n1995), .Z(n1997) );
  NAND U2586 ( .A(n1998), .B(n1997), .Z(n2176) );
  OR U2587 ( .A(oglobal[2]), .B(n1999), .Z(n2003) );
  NAND U2588 ( .A(n2001), .B(n2000), .Z(n2002) );
  NAND U2589 ( .A(n2003), .B(n2002), .Z(n2175) );
  OR U2590 ( .A(n2005), .B(n2004), .Z(n2009) );
  NANDN U2591 ( .A(n2007), .B(n2006), .Z(n2008) );
  NAND U2592 ( .A(n2009), .B(n2008), .Z(n2174) );
  XNOR U2593 ( .A(n2175), .B(n2174), .Z(n2010) );
  XNOR U2594 ( .A(n2176), .B(n2010), .Z(n2161) );
  OR U2595 ( .A(n2012), .B(n2011), .Z(n2016) );
  OR U2596 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2597 ( .A(n2016), .B(n2015), .Z(n2185) );
  OR U2598 ( .A(n2018), .B(n2017), .Z(n2022) );
  OR U2599 ( .A(n2020), .B(n2019), .Z(n2021) );
  AND U2600 ( .A(n2022), .B(n2021), .Z(n2184) );
  XNOR U2601 ( .A(oglobal[3]), .B(n2184), .Z(n2023) );
  XNOR U2602 ( .A(n2185), .B(n2023), .Z(n2159) );
  NANDN U2603 ( .A(n2025), .B(n2024), .Z(n2029) );
  NAND U2604 ( .A(n2027), .B(n2026), .Z(n2028) );
  AND U2605 ( .A(n2029), .B(n2028), .Z(n2158) );
  XNOR U2606 ( .A(n2159), .B(n2158), .Z(n2160) );
  XNOR U2607 ( .A(n2161), .B(n2160), .Z(n2234) );
  NANDN U2608 ( .A(n2035), .B(n2034), .Z(n2039) );
  NAND U2609 ( .A(n2037), .B(n2036), .Z(n2038) );
  NAND U2610 ( .A(n2039), .B(n2038), .Z(n2178) );
  OR U2611 ( .A(n2041), .B(n2040), .Z(n2045) );
  OR U2612 ( .A(n2043), .B(n2042), .Z(n2044) );
  NAND U2613 ( .A(n2045), .B(n2044), .Z(n2180) );
  OR U2614 ( .A(n2047), .B(n2046), .Z(n2051) );
  OR U2615 ( .A(n2049), .B(n2048), .Z(n2050) );
  NAND U2616 ( .A(n2051), .B(n2050), .Z(n2177) );
  IV U2617 ( .A(n2177), .Z(n2179) );
  XOR U2618 ( .A(n2180), .B(n2179), .Z(n2052) );
  XOR U2619 ( .A(n2178), .B(n2052), .Z(n2170) );
  NANDN U2620 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U2621 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U2622 ( .A(n2058), .B(n2057), .Z(n2189) );
  NANDN U2623 ( .A(n2060), .B(n2059), .Z(n2064) );
  NAND U2624 ( .A(n2062), .B(n2061), .Z(n2063) );
  AND U2625 ( .A(n2064), .B(n2063), .Z(n2186) );
  NANDN U2626 ( .A(n2066), .B(n2065), .Z(n2070) );
  NANDN U2627 ( .A(n2068), .B(n2067), .Z(n2069) );
  AND U2628 ( .A(n2070), .B(n2069), .Z(n2187) );
  XOR U2629 ( .A(n2186), .B(n2187), .Z(n2188) );
  NANDN U2630 ( .A(n2072), .B(n2071), .Z(n2076) );
  NAND U2631 ( .A(n2074), .B(n2073), .Z(n2075) );
  AND U2632 ( .A(n2076), .B(n2075), .Z(n2168) );
  XNOR U2633 ( .A(n2169), .B(n2168), .Z(n2171) );
  XOR U2634 ( .A(n2170), .B(n2171), .Z(n2232) );
  XOR U2635 ( .A(n2233), .B(n2232), .Z(n2235) );
  XNOR U2636 ( .A(n2234), .B(n2235), .Z(n2241) );
  XOR U2637 ( .A(n2240), .B(n2241), .Z(n2248) );
  NANDN U2638 ( .A(n2078), .B(n2077), .Z(n2082) );
  NAND U2639 ( .A(n2080), .B(n2079), .Z(n2081) );
  NAND U2640 ( .A(n2082), .B(n2081), .Z(n2246) );
  NAND U2641 ( .A(n2084), .B(n2083), .Z(n2088) );
  NANDN U2642 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U2643 ( .A(n2088), .B(n2087), .Z(n2155) );
  NANDN U2644 ( .A(n2090), .B(n2089), .Z(n2094) );
  NAND U2645 ( .A(n2092), .B(n2091), .Z(n2093) );
  AND U2646 ( .A(n2094), .B(n2093), .Z(n2166) );
  NANDN U2647 ( .A(n2100), .B(n2099), .Z(n2104) );
  NAND U2648 ( .A(n2102), .B(n2101), .Z(n2103) );
  AND U2649 ( .A(n2104), .B(n2103), .Z(n2165) );
  XOR U2650 ( .A(n2164), .B(n2165), .Z(n2167) );
  XOR U2651 ( .A(n2166), .B(n2167), .Z(n2154) );
  XOR U2652 ( .A(n2155), .B(n2154), .Z(n2157) );
  XOR U2653 ( .A(n2157), .B(n2156), .Z(n2247) );
  XNOR U2654 ( .A(n2246), .B(n2247), .Z(n2249) );
  XNOR U2655 ( .A(n2248), .B(n2249), .Z(n2261) );
  NAND U2656 ( .A(n2110), .B(n2109), .Z(n2114) );
  NANDN U2657 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U2658 ( .A(n2114), .B(n2113), .Z(n2259) );
  NANDN U2659 ( .A(n2120), .B(n2119), .Z(n2124) );
  NANDN U2660 ( .A(n2122), .B(n2121), .Z(n2123) );
  NAND U2661 ( .A(n2124), .B(n2123), .Z(n2204) );
  NANDN U2662 ( .A(n2134), .B(n2133), .Z(n2138) );
  NAND U2663 ( .A(n2136), .B(n2135), .Z(n2137) );
  NAND U2664 ( .A(n2138), .B(n2137), .Z(n2208) );
  XOR U2665 ( .A(n2209), .B(n2208), .Z(n2210) );
  XNOR U2666 ( .A(n2210), .B(n2211), .Z(n2203) );
  XNOR U2667 ( .A(n2202), .B(n2203), .Z(n2205) );
  XOR U2668 ( .A(n2204), .B(n2205), .Z(n2220) );
  NANDN U2669 ( .A(n2144), .B(n2143), .Z(n2148) );
  NANDN U2670 ( .A(n2146), .B(n2145), .Z(n2147) );
  NAND U2671 ( .A(n2148), .B(n2147), .Z(n2221) );
  XNOR U2672 ( .A(n2220), .B(n2221), .Z(n2222) );
  XNOR U2673 ( .A(n2223), .B(n2222), .Z(n2258) );
  XNOR U2674 ( .A(n2259), .B(n2258), .Z(n2260) );
  XNOR U2675 ( .A(n2261), .B(n2260), .Z(n2266) );
  XNOR U2676 ( .A(n2268), .B(n2266), .Z(n2149) );
  XNOR U2677 ( .A(n2264), .B(n2149), .Z(o[3]) );
  XOR U2678 ( .A(n2313), .B(n2314), .Z(n2316) );
  OR U2679 ( .A(n2159), .B(n2158), .Z(n2163) );
  OR U2680 ( .A(n2161), .B(n2160), .Z(n2162) );
  NAND U2681 ( .A(n2163), .B(n2162), .Z(n2320) );
  NAND U2682 ( .A(n2169), .B(n2168), .Z(n2173) );
  NANDN U2683 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2684 ( .A(n2173), .B(n2172), .Z(n2294) );
  NAND U2685 ( .A(n2177), .B(n2178), .Z(n2183) );
  ANDN U2686 ( .B(n2179), .A(n2178), .Z(n2181) );
  NANDN U2687 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U2688 ( .A(n2183), .B(n2182), .Z(n2324) );
  XOR U2689 ( .A(n2323), .B(n2324), .Z(n2326) );
  XNOR U2690 ( .A(n2329), .B(oglobal[4]), .Z(n2325) );
  OR U2691 ( .A(n2187), .B(n2186), .Z(n2191) );
  NANDN U2692 ( .A(n2189), .B(n2188), .Z(n2190) );
  AND U2693 ( .A(n2191), .B(n2190), .Z(n2330) );
  OR U2694 ( .A(n2193), .B(n2192), .Z(n2197) );
  OR U2695 ( .A(n2195), .B(n2194), .Z(n2196) );
  NAND U2696 ( .A(n2197), .B(n2196), .Z(n2331) );
  XNOR U2697 ( .A(n2330), .B(n2331), .Z(n2332) );
  XNOR U2698 ( .A(n2333), .B(n2332), .Z(n2293) );
  XNOR U2699 ( .A(n2294), .B(n2293), .Z(n2296) );
  XOR U2700 ( .A(n2296), .B(n2295), .Z(n2317) );
  XOR U2701 ( .A(n2320), .B(n2319), .Z(n2290) );
  NANDN U2702 ( .A(n2203), .B(n2202), .Z(n2207) );
  NAND U2703 ( .A(n2205), .B(n2204), .Z(n2206) );
  NAND U2704 ( .A(n2207), .B(n2206), .Z(n2287) );
  XOR U2705 ( .A(n2336), .B(n2337), .Z(n2338) );
  XOR U2706 ( .A(n2287), .B(n2288), .Z(n2289) );
  XOR U2707 ( .A(n2290), .B(n2289), .Z(n2315) );
  XNOR U2708 ( .A(n2316), .B(n2315), .Z(n2306) );
  OR U2709 ( .A(n2221), .B(n2220), .Z(n2225) );
  OR U2710 ( .A(n2223), .B(n2222), .Z(n2224) );
  NAND U2711 ( .A(n2225), .B(n2224), .Z(n2304) );
  NANDN U2712 ( .A(n2227), .B(n2226), .Z(n2231) );
  NANDN U2713 ( .A(n2229), .B(n2228), .Z(n2230) );
  NAND U2714 ( .A(n2231), .B(n2230), .Z(n2303) );
  XNOR U2715 ( .A(n2304), .B(n2303), .Z(n2305) );
  XNOR U2716 ( .A(n2306), .B(n2305), .Z(n2275) );
  NANDN U2717 ( .A(n2233), .B(n2232), .Z(n2237) );
  NANDN U2718 ( .A(n2235), .B(n2234), .Z(n2236) );
  NAND U2719 ( .A(n2237), .B(n2236), .Z(n2301) );
  XOR U2720 ( .A(n2299), .B(n2300), .Z(n2302) );
  XOR U2721 ( .A(n2301), .B(n2302), .Z(n2309) );
  NANDN U2722 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2723 ( .A(n2249), .B(n2248), .Z(n2250) );
  AND U2724 ( .A(n2251), .B(n2250), .Z(n2310) );
  XNOR U2725 ( .A(n2309), .B(n2310), .Z(n2312) );
  NANDN U2726 ( .A(n2253), .B(n2252), .Z(n2257) );
  NAND U2727 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2728 ( .A(n2257), .B(n2256), .Z(n2311) );
  XOR U2729 ( .A(n2312), .B(n2311), .Z(n2276) );
  XNOR U2730 ( .A(n2275), .B(n2276), .Z(n2278) );
  OR U2731 ( .A(n2259), .B(n2258), .Z(n2263) );
  OR U2732 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U2733 ( .A(n2263), .B(n2262), .Z(n2277) );
  XOR U2734 ( .A(n2278), .B(n2277), .Z(n2283) );
  NAND U2735 ( .A(n2264), .B(n2266), .Z(n2270) );
  NANDN U2736 ( .A(n2266), .B(n2265), .Z(n2267) );
  NANDN U2737 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U2738 ( .A(n2270), .B(n2269), .Z(n2282) );
  XNOR U2739 ( .A(n2282), .B(n2281), .Z(n2284) );
  XOR U2740 ( .A(n2283), .B(n2284), .Z(o[4]) );
  NAND U2741 ( .A(n2276), .B(n2275), .Z(n2280) );
  OR U2742 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U2743 ( .A(n2280), .B(n2279), .Z(n2351) );
  NANDN U2744 ( .A(n2282), .B(n2281), .Z(n2286) );
  NAND U2745 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U2746 ( .A(n2286), .B(n2285), .Z(n2349) );
  NANDN U2747 ( .A(n2288), .B(n2287), .Z(n2292) );
  OR U2748 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U2749 ( .A(n2292), .B(n2291), .Z(n2357) );
  OR U2750 ( .A(n2294), .B(n2293), .Z(n2298) );
  OR U2751 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2752 ( .A(n2298), .B(n2297), .Z(n2356) );
  XOR U2753 ( .A(n2357), .B(n2356), .Z(n2359) );
  XOR U2754 ( .A(n2359), .B(n2358), .Z(n2343) );
  OR U2755 ( .A(n2304), .B(n2303), .Z(n2308) );
  OR U2756 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2757 ( .A(n2308), .B(n2307), .Z(n2344) );
  XNOR U2758 ( .A(n2343), .B(n2344), .Z(n2346) );
  NANDN U2759 ( .A(n2318), .B(n2317), .Z(n2322) );
  NANDN U2760 ( .A(n2320), .B(n2319), .Z(n2321) );
  AND U2761 ( .A(n2322), .B(n2321), .Z(n2362) );
  NANDN U2762 ( .A(n2324), .B(n2323), .Z(n2328) );
  NANDN U2763 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U2764 ( .A(n2328), .B(n2327), .Z(n2365) );
  NANDN U2765 ( .A(n2329), .B(oglobal[4]), .Z(n2364) );
  XOR U2766 ( .A(oglobal[5]), .B(n2364), .Z(n2366) );
  XNOR U2767 ( .A(n2365), .B(n2366), .Z(n2368) );
  OR U2768 ( .A(n2331), .B(n2330), .Z(n2335) );
  OR U2769 ( .A(n2333), .B(n2332), .Z(n2334) );
  NAND U2770 ( .A(n2335), .B(n2334), .Z(n2367) );
  XOR U2771 ( .A(n2368), .B(n2367), .Z(n2360) );
  OR U2772 ( .A(n2337), .B(n2336), .Z(n2341) );
  NANDN U2773 ( .A(n2339), .B(n2338), .Z(n2340) );
  AND U2774 ( .A(n2341), .B(n2340), .Z(n2361) );
  XNOR U2775 ( .A(n2360), .B(n2361), .Z(n2363) );
  XOR U2776 ( .A(n2362), .B(n2363), .Z(n2353) );
  XOR U2777 ( .A(n2352), .B(n2353), .Z(n2354) );
  XOR U2778 ( .A(n2355), .B(n2354), .Z(n2345) );
  XNOR U2779 ( .A(n2349), .B(n2350), .Z(n2342) );
  XOR U2780 ( .A(n2351), .B(n2342), .Z(o[5]) );
  OR U2781 ( .A(n2344), .B(n2343), .Z(n2348) );
  NANDN U2782 ( .A(n2346), .B(n2345), .Z(n2347) );
  AND U2783 ( .A(n2348), .B(n2347), .Z(n2379) );
  NANDN U2784 ( .A(n2364), .B(oglobal[5]), .Z(n2371) );
  XOR U2785 ( .A(oglobal[6]), .B(n2371), .Z(n2372) );
  OR U2786 ( .A(n2366), .B(n2365), .Z(n2370) );
  OR U2787 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U2788 ( .A(n2370), .B(n2369), .Z(n2373) );
  XNOR U2789 ( .A(n2372), .B(n2373), .Z(n2374) );
  XOR U2790 ( .A(n2375), .B(n2374), .Z(n2384) );
  XNOR U2791 ( .A(n2385), .B(n2384), .Z(n2387) );
  XOR U2792 ( .A(n2386), .B(n2387), .Z(n2380) );
  XNOR U2793 ( .A(n2381), .B(n2380), .Z(n2378) );
  XOR U2794 ( .A(n2379), .B(n2378), .Z(o[6]) );
  NANDN U2795 ( .A(n2371), .B(oglobal[6]), .Z(n2392) );
  XOR U2796 ( .A(oglobal[7]), .B(n2392), .Z(n2394) );
  NANDN U2797 ( .A(n2373), .B(n2372), .Z(n2377) );
  NANDN U2798 ( .A(n2375), .B(n2374), .Z(n2376) );
  NAND U2799 ( .A(n2377), .B(n2376), .Z(n2393) );
  XNOR U2800 ( .A(n2394), .B(n2393), .Z(n2391) );
  NANDN U2801 ( .A(n2379), .B(n2378), .Z(n2383) );
  NANDN U2802 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U2803 ( .A(n2383), .B(n2382), .Z(n2390) );
  XOR U2804 ( .A(n2390), .B(n2389), .Z(n2388) );
  XOR U2805 ( .A(n2391), .B(n2388), .Z(o[7]) );
  XNOR U2806 ( .A(n2397), .B(oglobal[8]), .Z(n2399) );
  NANDN U2807 ( .A(n2392), .B(oglobal[7]), .Z(n2396) );
  OR U2808 ( .A(n2394), .B(n2393), .Z(n2395) );
  AND U2809 ( .A(n2396), .B(n2395), .Z(n2398) );
  XOR U2810 ( .A(n2399), .B(n2398), .Z(o[8]) );
  NAND U2811 ( .A(n2397), .B(oglobal[8]), .Z(n2401) );
  OR U2812 ( .A(n2399), .B(n2398), .Z(n2400) );
  NAND U2813 ( .A(n2401), .B(n2400), .Z(n2402) );
  XOR U2814 ( .A(n2402), .B(oglobal[9]), .Z(o[9]) );
  NAND U2815 ( .A(oglobal[9]), .B(n2402), .Z(n2403) );
  XNOR U2816 ( .A(oglobal[10]), .B(n2403), .Z(o[10]) );
endmodule

