
module hamming_N1600_CC16 ( clk, rst, x, y, o );
  input [99:0] x;
  input [99:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U103 ( .A(n334), .B(n333), .Z(n1) );
  NAND U104 ( .A(n331), .B(n332), .Z(n2) );
  NAND U105 ( .A(n1), .B(n2), .Z(n494) );
  XOR U106 ( .A(n518), .B(oglobal[1]), .Z(n3) );
  NANDN U107 ( .A(n519), .B(n3), .Z(n4) );
  NAND U108 ( .A(n518), .B(oglobal[1]), .Z(n5) );
  AND U109 ( .A(n4), .B(n5), .Z(n560) );
  XOR U110 ( .A(n544), .B(n542), .Z(n6) );
  NANDN U111 ( .A(n543), .B(n6), .Z(n7) );
  NAND U112 ( .A(n544), .B(n542), .Z(n8) );
  AND U113 ( .A(n7), .B(n8), .Z(n575) );
  NAND U114 ( .A(n438), .B(n439), .Z(n9) );
  XOR U115 ( .A(n438), .B(n439), .Z(n10) );
  NANDN U116 ( .A(n437), .B(n10), .Z(n11) );
  NAND U117 ( .A(n9), .B(n11), .Z(n584) );
  NAND U118 ( .A(n578), .B(n580), .Z(n12) );
  XOR U119 ( .A(n578), .B(n580), .Z(n13) );
  NAND U120 ( .A(n13), .B(n579), .Z(n14) );
  NAND U121 ( .A(n12), .B(n14), .Z(n626) );
  NAND U122 ( .A(n571), .B(n573), .Z(n15) );
  XOR U123 ( .A(n571), .B(n573), .Z(n16) );
  NAND U124 ( .A(n16), .B(n572), .Z(n17) );
  NAND U125 ( .A(n15), .B(n17), .Z(n632) );
  NAND U126 ( .A(n330), .B(n329), .Z(n18) );
  NAND U127 ( .A(n327), .B(n328), .Z(n19) );
  AND U128 ( .A(n18), .B(n19), .Z(n493) );
  NAND U129 ( .A(n179), .B(n178), .Z(n20) );
  NAND U130 ( .A(n176), .B(n177), .Z(n21) );
  NAND U131 ( .A(n20), .B(n21), .Z(n503) );
  XOR U132 ( .A(n306), .B(n304), .Z(n22) );
  NANDN U133 ( .A(n305), .B(n22), .Z(n23) );
  NAND U134 ( .A(n306), .B(n304), .Z(n24) );
  AND U135 ( .A(n23), .B(n24), .Z(n524) );
  NAND U136 ( .A(n513), .B(n514), .Z(n25) );
  XOR U137 ( .A(n513), .B(n514), .Z(n26) );
  NANDN U138 ( .A(n512), .B(n26), .Z(n27) );
  NAND U139 ( .A(n25), .B(n27), .Z(n555) );
  NAND U140 ( .A(n516), .B(n517), .Z(n28) );
  XOR U141 ( .A(n516), .B(n517), .Z(n29) );
  NANDN U142 ( .A(n515), .B(n29), .Z(n30) );
  NAND U143 ( .A(n28), .B(n30), .Z(n561) );
  XOR U144 ( .A(n466), .B(n467), .Z(n31) );
  NANDN U145 ( .A(n468), .B(n31), .Z(n32) );
  NAND U146 ( .A(n466), .B(n467), .Z(n33) );
  AND U147 ( .A(n32), .B(n33), .Z(n557) );
  XOR U148 ( .A(n477), .B(n478), .Z(n34) );
  NANDN U149 ( .A(n479), .B(n34), .Z(n35) );
  NAND U150 ( .A(n477), .B(n478), .Z(n36) );
  AND U151 ( .A(n35), .B(n36), .Z(n569) );
  XOR U152 ( .A(n501), .B(n499), .Z(n37) );
  NANDN U153 ( .A(n500), .B(n37), .Z(n38) );
  NAND U154 ( .A(n501), .B(n499), .Z(n39) );
  AND U155 ( .A(n38), .B(n39), .Z(n563) );
  XNOR U156 ( .A(n455), .B(n454), .Z(n457) );
  NAND U157 ( .A(n441), .B(n442), .Z(n40) );
  XOR U158 ( .A(n441), .B(n442), .Z(n41) );
  NANDN U159 ( .A(n440), .B(n41), .Z(n42) );
  NAND U160 ( .A(n40), .B(n42), .Z(n586) );
  NAND U161 ( .A(n576), .B(n577), .Z(n43) );
  XOR U162 ( .A(n576), .B(n577), .Z(n44) );
  NANDN U163 ( .A(n575), .B(n44), .Z(n45) );
  NAND U164 ( .A(n43), .B(n45), .Z(n628) );
  NAND U165 ( .A(n162), .B(n163), .Z(n46) );
  XOR U166 ( .A(n162), .B(n163), .Z(n47) );
  NANDN U167 ( .A(n161), .B(n47), .Z(n48) );
  NAND U168 ( .A(n46), .B(n48), .Z(n439) );
  XOR U169 ( .A(n633), .B(n631), .Z(n49) );
  NANDN U170 ( .A(n632), .B(n49), .Z(n50) );
  NAND U171 ( .A(n633), .B(n631), .Z(n51) );
  AND U172 ( .A(n50), .B(n51), .Z(n642) );
  NAND U173 ( .A(n638), .B(n639), .Z(n52) );
  XOR U174 ( .A(n638), .B(n639), .Z(n53) );
  NAND U175 ( .A(n53), .B(n637), .Z(n54) );
  NAND U176 ( .A(n52), .B(n54), .Z(n655) );
  NAND U177 ( .A(n350), .B(n349), .Z(n55) );
  NAND U178 ( .A(n347), .B(n348), .Z(n56) );
  AND U179 ( .A(n55), .B(n56), .Z(n460) );
  NAND U180 ( .A(n464), .B(n465), .Z(n57) );
  XOR U181 ( .A(n464), .B(n465), .Z(n58) );
  NANDN U182 ( .A(n463), .B(n58), .Z(n59) );
  NAND U183 ( .A(n57), .B(n59), .Z(n558) );
  NAND U184 ( .A(n509), .B(n511), .Z(n60) );
  XOR U185 ( .A(n509), .B(n511), .Z(n61) );
  NAND U186 ( .A(n61), .B(n510), .Z(n62) );
  NAND U187 ( .A(n60), .B(n62), .Z(n583) );
  XOR U188 ( .A(n523), .B(n521), .Z(n63) );
  NANDN U189 ( .A(n522), .B(n63), .Z(n64) );
  NAND U190 ( .A(n523), .B(n521), .Z(n65) );
  AND U191 ( .A(n64), .B(n65), .Z(n580) );
  NAND U192 ( .A(n541), .B(n538), .Z(n66) );
  NANDN U193 ( .A(n541), .B(n540), .Z(n67) );
  NANDN U194 ( .A(n539), .B(n67), .Z(n68) );
  NAND U195 ( .A(n66), .B(n68), .Z(n577) );
  XOR U196 ( .A(n561), .B(n559), .Z(n69) );
  NANDN U197 ( .A(n560), .B(n69), .Z(n70) );
  NAND U198 ( .A(n561), .B(n559), .Z(n71) );
  AND U199 ( .A(n70), .B(n71), .Z(n618) );
  NAND U200 ( .A(n564), .B(n565), .Z(n72) );
  XOR U201 ( .A(n564), .B(n565), .Z(n73) );
  NANDN U202 ( .A(n563), .B(n73), .Z(n74) );
  NAND U203 ( .A(n72), .B(n74), .Z(n615) );
  NAND U204 ( .A(n444), .B(n445), .Z(n75) );
  XOR U205 ( .A(n444), .B(n445), .Z(n76) );
  NANDN U206 ( .A(n443), .B(n76), .Z(n77) );
  NAND U207 ( .A(n75), .B(n77), .Z(n585) );
  NAND U208 ( .A(n159), .B(n160), .Z(n78) );
  XOR U209 ( .A(n159), .B(n160), .Z(n79) );
  NANDN U210 ( .A(n158), .B(n79), .Z(n80) );
  NAND U211 ( .A(n78), .B(n80), .Z(n438) );
  XOR U212 ( .A(n642), .B(n640), .Z(n81) );
  NANDN U213 ( .A(n641), .B(n81), .Z(n82) );
  NAND U214 ( .A(n642), .B(n640), .Z(n83) );
  AND U215 ( .A(n82), .B(n83), .Z(n652) );
  NAND U216 ( .A(n556), .B(n558), .Z(n84) );
  XOR U217 ( .A(n556), .B(n558), .Z(n85) );
  NAND U218 ( .A(n85), .B(n557), .Z(n86) );
  NAND U219 ( .A(n84), .B(n86), .Z(n621) );
  NAND U220 ( .A(n569), .B(n568), .Z(n87) );
  NAND U221 ( .A(n566), .B(n567), .Z(n88) );
  NAND U222 ( .A(n87), .B(n88), .Z(n614) );
  XNOR U223 ( .A(n443), .B(n444), .Z(n89) );
  XNOR U224 ( .A(n445), .B(n89), .Z(n454) );
  NAND U225 ( .A(n582), .B(n583), .Z(n90) );
  XOR U226 ( .A(n582), .B(n583), .Z(n91) );
  NANDN U227 ( .A(n581), .B(n91), .Z(n92) );
  NAND U228 ( .A(n90), .B(n92), .Z(n625) );
  NAND U229 ( .A(n553), .B(n554), .Z(n93) );
  XOR U230 ( .A(n553), .B(n554), .Z(n94) );
  NANDN U231 ( .A(n552), .B(n94), .Z(n95) );
  NAND U232 ( .A(n93), .B(n95), .Z(n633) );
  XOR U233 ( .A(n166), .B(n164), .Z(n96) );
  XNOR U234 ( .A(n167), .B(n96), .Z(n412) );
  NANDN U235 ( .A(n547), .B(n550), .Z(n97) );
  OR U236 ( .A(n550), .B(n549), .Z(n98) );
  NANDN U237 ( .A(n548), .B(n98), .Z(n99) );
  NAND U238 ( .A(n97), .B(n99), .Z(n590) );
  NAND U239 ( .A(n584), .B(n586), .Z(n100) );
  XOR U240 ( .A(n584), .B(n586), .Z(n101) );
  NAND U241 ( .A(n101), .B(n585), .Z(n102) );
  NAND U242 ( .A(n100), .B(n102), .Z(n611) );
  NAND U243 ( .A(n651), .B(n653), .Z(n103) );
  XOR U244 ( .A(n651), .B(n653), .Z(n104) );
  NAND U245 ( .A(n104), .B(n652), .Z(n105) );
  NAND U246 ( .A(n103), .B(n105), .Z(n661) );
  NAND U247 ( .A(n310), .B(n309), .Z(n106) );
  NAND U248 ( .A(n307), .B(n308), .Z(n107) );
  NAND U249 ( .A(n106), .B(n107), .Z(n501) );
  NAND U250 ( .A(n175), .B(n174), .Z(n108) );
  NAND U251 ( .A(n172), .B(n173), .Z(n109) );
  AND U252 ( .A(n108), .B(n109), .Z(n504) );
  NAND U253 ( .A(n302), .B(n303), .Z(n110) );
  XOR U254 ( .A(n302), .B(n303), .Z(n111) );
  NANDN U255 ( .A(n301), .B(n111), .Z(n112) );
  NAND U256 ( .A(n110), .B(n112), .Z(n525) );
  NAND U257 ( .A(n325), .B(n326), .Z(n113) );
  XOR U258 ( .A(n325), .B(n326), .Z(n114) );
  NANDN U259 ( .A(n324), .B(n114), .Z(n115) );
  NAND U260 ( .A(n113), .B(n115), .Z(n533) );
  XOR U261 ( .A(n260), .B(n261), .Z(n116) );
  NANDN U262 ( .A(n262), .B(n116), .Z(n117) );
  NAND U263 ( .A(n260), .B(n261), .Z(n118) );
  AND U264 ( .A(n117), .B(n118), .Z(n474) );
  NAND U265 ( .A(n461), .B(n462), .Z(n119) );
  XOR U266 ( .A(n461), .B(n462), .Z(n120) );
  NANDN U267 ( .A(n460), .B(n120), .Z(n121) );
  NAND U268 ( .A(n119), .B(n121), .Z(n556) );
  NAND U269 ( .A(n230), .B(n231), .Z(n122) );
  XOR U270 ( .A(n230), .B(n231), .Z(n123) );
  NANDN U271 ( .A(n229), .B(n123), .Z(n124) );
  NAND U272 ( .A(n122), .B(n124), .Z(n539) );
  XOR U273 ( .A(n206), .B(n207), .Z(n125) );
  NANDN U274 ( .A(n208), .B(n125), .Z(n126) );
  NAND U275 ( .A(n206), .B(n207), .Z(n127) );
  AND U276 ( .A(n126), .B(n127), .Z(n542) );
  XOR U277 ( .A(n582), .B(n581), .Z(n128) );
  XNOR U278 ( .A(n583), .B(n128), .Z(n579) );
  AND U279 ( .A(n613), .B(oglobal[3]), .Z(n636) );
  NAND U280 ( .A(n615), .B(n614), .Z(n129) );
  XOR U281 ( .A(n615), .B(n614), .Z(n130) );
  NANDN U282 ( .A(n616), .B(n130), .Z(n131) );
  NAND U283 ( .A(n129), .B(n131), .Z(n639) );
  XOR U284 ( .A(n155), .B(n156), .Z(n132) );
  NANDN U285 ( .A(n157), .B(n132), .Z(n133) );
  NAND U286 ( .A(n155), .B(n156), .Z(n134) );
  AND U287 ( .A(n133), .B(n134), .Z(n449) );
  XOR U288 ( .A(n590), .B(n588), .Z(n135) );
  XNOR U289 ( .A(n591), .B(n135), .Z(n598) );
  NAND U290 ( .A(n611), .B(n612), .Z(n136) );
  XOR U291 ( .A(n611), .B(n612), .Z(n137) );
  NANDN U292 ( .A(n610), .B(n137), .Z(n138) );
  NAND U293 ( .A(n136), .B(n138), .Z(n647) );
  XOR U294 ( .A(oglobal[6]), .B(n660), .Z(n139) );
  NANDN U295 ( .A(n661), .B(n139), .Z(n140) );
  NAND U296 ( .A(oglobal[6]), .B(n660), .Z(n141) );
  AND U297 ( .A(n140), .B(n141), .Z(n662) );
  XOR U298 ( .A(x[53]), .B(y[53]), .Z(n213) );
  XOR U299 ( .A(x[51]), .B(y[51]), .Z(n210) );
  XOR U300 ( .A(x[49]), .B(y[49]), .Z(n211) );
  XOR U301 ( .A(n210), .B(n211), .Z(n212) );
  XOR U302 ( .A(n213), .B(n212), .Z(n325) );
  XOR U303 ( .A(x[47]), .B(y[47]), .Z(n225) );
  XOR U304 ( .A(x[45]), .B(y[45]), .Z(n222) );
  XOR U305 ( .A(x[43]), .B(y[43]), .Z(n223) );
  XOR U306 ( .A(n222), .B(n223), .Z(n224) );
  XOR U307 ( .A(n225), .B(n224), .Z(n326) );
  XOR U308 ( .A(x[57]), .B(y[57]), .Z(n361) );
  XOR U309 ( .A(x[99]), .B(y[99]), .Z(n359) );
  XNOR U310 ( .A(x[55]), .B(y[55]), .Z(n360) );
  XOR U311 ( .A(n359), .B(n360), .Z(n362) );
  XOR U312 ( .A(n361), .B(n362), .Z(n324) );
  XOR U313 ( .A(n326), .B(n324), .Z(n142) );
  XOR U314 ( .A(n325), .B(n142), .Z(n160) );
  XOR U315 ( .A(x[17]), .B(y[17]), .Z(n391) );
  XOR U316 ( .A(x[15]), .B(y[15]), .Z(n389) );
  XNOR U317 ( .A(x[13]), .B(y[13]), .Z(n390) );
  XOR U318 ( .A(n389), .B(n390), .Z(n392) );
  XOR U319 ( .A(n391), .B(n392), .Z(n261) );
  XOR U320 ( .A(x[11]), .B(y[11]), .Z(n397) );
  XOR U321 ( .A(x[9]), .B(y[9]), .Z(n395) );
  XNOR U322 ( .A(x[7]), .B(y[7]), .Z(n396) );
  XOR U323 ( .A(n395), .B(n396), .Z(n398) );
  XNOR U324 ( .A(n397), .B(n398), .Z(n262) );
  XOR U325 ( .A(x[23]), .B(y[23]), .Z(n195) );
  XOR U326 ( .A(x[21]), .B(y[21]), .Z(n193) );
  XNOR U327 ( .A(x[19]), .B(y[19]), .Z(n194) );
  XOR U328 ( .A(n193), .B(n194), .Z(n196) );
  XOR U329 ( .A(n195), .B(n196), .Z(n260) );
  XOR U330 ( .A(n262), .B(n260), .Z(n143) );
  XNOR U331 ( .A(n261), .B(n143), .Z(n159) );
  XOR U332 ( .A(x[35]), .B(y[35]), .Z(n189) );
  XOR U333 ( .A(x[33]), .B(y[33]), .Z(n187) );
  XNOR U334 ( .A(x[31]), .B(y[31]), .Z(n188) );
  XOR U335 ( .A(n187), .B(n188), .Z(n190) );
  XOR U336 ( .A(n189), .B(n190), .Z(n254) );
  XOR U337 ( .A(x[29]), .B(y[29]), .Z(n201) );
  XOR U338 ( .A(x[27]), .B(y[27]), .Z(n199) );
  XNOR U339 ( .A(x[25]), .B(y[25]), .Z(n200) );
  XOR U340 ( .A(n199), .B(n200), .Z(n202) );
  XNOR U341 ( .A(n201), .B(n202), .Z(n257) );
  XOR U342 ( .A(x[41]), .B(y[41]), .Z(n218) );
  XOR U343 ( .A(x[39]), .B(y[39]), .Z(n216) );
  XNOR U344 ( .A(x[37]), .B(y[37]), .Z(n217) );
  XOR U345 ( .A(n216), .B(n217), .Z(n219) );
  XOR U346 ( .A(n218), .B(n219), .Z(n253) );
  XOR U347 ( .A(n257), .B(n253), .Z(n144) );
  XOR U348 ( .A(n254), .B(n144), .Z(n158) );
  XOR U349 ( .A(n159), .B(n158), .Z(n145) );
  XNOR U350 ( .A(n160), .B(n145), .Z(n157) );
  XOR U351 ( .A(x[0]), .B(y[0]), .Z(n292) );
  XOR U352 ( .A(x[2]), .B(y[2]), .Z(n290) );
  XOR U353 ( .A(x[4]), .B(y[4]), .Z(n289) );
  XOR U354 ( .A(n290), .B(n289), .Z(n291) );
  XNOR U355 ( .A(n292), .B(n291), .Z(n303) );
  XOR U356 ( .A(x[5]), .B(y[5]), .Z(n286) );
  XOR U357 ( .A(x[1]), .B(y[1]), .Z(n284) );
  XOR U358 ( .A(x[3]), .B(y[3]), .Z(n283) );
  XOR U359 ( .A(n284), .B(n283), .Z(n285) );
  XNOR U360 ( .A(n286), .B(n285), .Z(n302) );
  XOR U361 ( .A(x[6]), .B(y[6]), .Z(n278) );
  XOR U362 ( .A(x[10]), .B(y[10]), .Z(n276) );
  XOR U363 ( .A(x[8]), .B(y[8]), .Z(n275) );
  XOR U364 ( .A(n276), .B(n275), .Z(n277) );
  XOR U365 ( .A(n278), .B(n277), .Z(n301) );
  XOR U366 ( .A(n302), .B(n301), .Z(n146) );
  XNOR U367 ( .A(n303), .B(n146), .Z(n163) );
  XOR U368 ( .A(x[90]), .B(y[90]), .Z(n297) );
  XNOR U369 ( .A(x[92]), .B(y[92]), .Z(n295) );
  XNOR U370 ( .A(oglobal[0]), .B(n295), .Z(n296) );
  XNOR U371 ( .A(n297), .B(n296), .Z(n231) );
  XOR U372 ( .A(x[78]), .B(y[78]), .Z(n314) );
  XOR U373 ( .A(x[82]), .B(y[82]), .Z(n311) );
  XNOR U374 ( .A(x[80]), .B(y[80]), .Z(n312) );
  XNOR U375 ( .A(n311), .B(n312), .Z(n313) );
  XNOR U376 ( .A(n314), .B(n313), .Z(n230) );
  XOR U377 ( .A(x[84]), .B(y[84]), .Z(n272) );
  XOR U378 ( .A(x[88]), .B(y[88]), .Z(n269) );
  XNOR U379 ( .A(x[86]), .B(y[86]), .Z(n270) );
  XNOR U380 ( .A(n269), .B(n270), .Z(n271) );
  XOR U381 ( .A(n272), .B(n271), .Z(n229) );
  XOR U382 ( .A(n230), .B(n229), .Z(n147) );
  XNOR U383 ( .A(n231), .B(n147), .Z(n162) );
  XOR U384 ( .A(x[18]), .B(y[18]), .Z(n319) );
  XOR U385 ( .A(x[22]), .B(y[22]), .Z(n318) );
  XOR U386 ( .A(x[20]), .B(y[20]), .Z(n317) );
  XNOR U387 ( .A(n318), .B(n317), .Z(n320) );
  XNOR U388 ( .A(n319), .B(n320), .Z(n430) );
  XOR U389 ( .A(x[12]), .B(y[12]), .Z(n266) );
  XOR U390 ( .A(x[16]), .B(y[16]), .Z(n264) );
  XOR U391 ( .A(x[14]), .B(y[14]), .Z(n263) );
  XOR U392 ( .A(n264), .B(n263), .Z(n265) );
  XOR U393 ( .A(n266), .B(n265), .Z(n429) );
  XOR U394 ( .A(x[24]), .B(y[24]), .Z(n310) );
  XOR U395 ( .A(x[28]), .B(y[28]), .Z(n308) );
  XOR U396 ( .A(x[26]), .B(y[26]), .Z(n307) );
  XOR U397 ( .A(n308), .B(n307), .Z(n309) );
  XOR U398 ( .A(n310), .B(n309), .Z(n428) );
  XNOR U399 ( .A(n429), .B(n428), .Z(n148) );
  XNOR U400 ( .A(n430), .B(n148), .Z(n161) );
  XOR U401 ( .A(n162), .B(n161), .Z(n149) );
  XOR U402 ( .A(n163), .B(n149), .Z(n155) );
  XOR U403 ( .A(x[54]), .B(y[54]), .Z(n330) );
  XOR U404 ( .A(x[58]), .B(y[58]), .Z(n328) );
  XOR U405 ( .A(x[56]), .B(y[56]), .Z(n327) );
  XOR U406 ( .A(n328), .B(n327), .Z(n329) );
  XOR U407 ( .A(n330), .B(n329), .Z(n421) );
  XOR U408 ( .A(x[60]), .B(y[60]), .Z(n175) );
  XOR U409 ( .A(x[64]), .B(y[64]), .Z(n173) );
  XOR U410 ( .A(x[62]), .B(y[62]), .Z(n172) );
  XOR U411 ( .A(n173), .B(n172), .Z(n174) );
  XOR U412 ( .A(n175), .B(n174), .Z(n425) );
  XOR U413 ( .A(x[48]), .B(y[48]), .Z(n334) );
  XOR U414 ( .A(x[52]), .B(y[52]), .Z(n332) );
  XOR U415 ( .A(x[50]), .B(y[50]), .Z(n331) );
  XOR U416 ( .A(n332), .B(n331), .Z(n333) );
  XOR U417 ( .A(n334), .B(n333), .Z(n423) );
  XNOR U418 ( .A(n425), .B(n423), .Z(n150) );
  XOR U419 ( .A(n421), .B(n150), .Z(n167) );
  XOR U420 ( .A(x[42]), .B(y[42]), .Z(n182) );
  XOR U421 ( .A(x[46]), .B(y[46]), .Z(n180) );
  XNOR U422 ( .A(x[44]), .B(y[44]), .Z(n181) );
  XOR U423 ( .A(n180), .B(n181), .Z(n183) );
  XOR U424 ( .A(n182), .B(n183), .Z(n247) );
  XOR U425 ( .A(x[36]), .B(y[36]), .Z(n344) );
  XOR U426 ( .A(x[40]), .B(y[40]), .Z(n341) );
  XNOR U427 ( .A(x[38]), .B(y[38]), .Z(n342) );
  XNOR U428 ( .A(n341), .B(n342), .Z(n343) );
  XNOR U429 ( .A(n344), .B(n343), .Z(n246) );
  XOR U430 ( .A(n247), .B(n246), .Z(n249) );
  XOR U431 ( .A(x[30]), .B(y[30]), .Z(n337) );
  XOR U432 ( .A(x[34]), .B(y[34]), .Z(n335) );
  XNOR U433 ( .A(x[32]), .B(y[32]), .Z(n336) );
  XOR U434 ( .A(n335), .B(n336), .Z(n338) );
  XOR U435 ( .A(n337), .B(n338), .Z(n248) );
  XOR U436 ( .A(n249), .B(n248), .Z(n165) );
  IV U437 ( .A(n165), .Z(n164) );
  XOR U438 ( .A(x[94]), .B(y[94]), .Z(n404) );
  XOR U439 ( .A(x[98]), .B(y[98]), .Z(n401) );
  XOR U440 ( .A(x[96]), .B(y[96]), .Z(n402) );
  XOR U441 ( .A(n401), .B(n402), .Z(n403) );
  XOR U442 ( .A(n404), .B(n403), .Z(n415) );
  XOR U443 ( .A(x[72]), .B(y[72]), .Z(n350) );
  XOR U444 ( .A(x[76]), .B(y[76]), .Z(n348) );
  XOR U445 ( .A(x[74]), .B(y[74]), .Z(n347) );
  XOR U446 ( .A(n348), .B(n347), .Z(n349) );
  XOR U447 ( .A(n350), .B(n349), .Z(n418) );
  XOR U448 ( .A(x[66]), .B(y[66]), .Z(n179) );
  XOR U449 ( .A(x[70]), .B(y[70]), .Z(n177) );
  XOR U450 ( .A(x[68]), .B(y[68]), .Z(n176) );
  XOR U451 ( .A(n177), .B(n176), .Z(n178) );
  XOR U452 ( .A(n179), .B(n178), .Z(n416) );
  XNOR U453 ( .A(n418), .B(n416), .Z(n151) );
  XNOR U454 ( .A(n415), .B(n151), .Z(n166) );
  XOR U455 ( .A(x[61]), .B(y[61]), .Z(n368) );
  XOR U456 ( .A(x[97]), .B(y[97]), .Z(n365) );
  XOR U457 ( .A(x[59]), .B(y[59]), .Z(n366) );
  XOR U458 ( .A(n365), .B(n366), .Z(n367) );
  XOR U459 ( .A(n368), .B(n367), .Z(n306) );
  XOR U460 ( .A(x[77]), .B(y[77]), .Z(n235) );
  XOR U461 ( .A(x[89]), .B(y[89]), .Z(n233) );
  XOR U462 ( .A(x[75]), .B(y[75]), .Z(n232) );
  XOR U463 ( .A(n233), .B(n232), .Z(n234) );
  XOR U464 ( .A(n235), .B(n234), .Z(n380) );
  XOR U465 ( .A(x[85]), .B(y[85]), .Z(n377) );
  XOR U466 ( .A(x[83]), .B(y[83]), .Z(n378) );
  XOR U467 ( .A(n377), .B(n378), .Z(n379) );
  XNOR U468 ( .A(n380), .B(n379), .Z(n305) );
  XOR U469 ( .A(x[69]), .B(y[69]), .Z(n386) );
  XOR U470 ( .A(x[93]), .B(y[93]), .Z(n383) );
  XOR U471 ( .A(x[67]), .B(y[67]), .Z(n384) );
  XOR U472 ( .A(n383), .B(n384), .Z(n385) );
  XOR U473 ( .A(n386), .B(n385), .Z(n304) );
  XOR U474 ( .A(n305), .B(n304), .Z(n152) );
  XNOR U475 ( .A(n306), .B(n152), .Z(n410) );
  XOR U476 ( .A(x[81]), .B(y[81]), .Z(n373) );
  XOR U477 ( .A(x[87]), .B(y[87]), .Z(n371) );
  XNOR U478 ( .A(x[79]), .B(y[79]), .Z(n372) );
  XOR U479 ( .A(n371), .B(n372), .Z(n374) );
  XOR U480 ( .A(n373), .B(n374), .Z(n207) );
  XOR U481 ( .A(x[65]), .B(y[65]), .Z(n355) );
  XOR U482 ( .A(x[95]), .B(y[95]), .Z(n353) );
  XNOR U483 ( .A(x[63]), .B(y[63]), .Z(n354) );
  XOR U484 ( .A(n353), .B(n354), .Z(n356) );
  XNOR U485 ( .A(n355), .B(n356), .Z(n208) );
  XOR U486 ( .A(x[73]), .B(y[73]), .Z(n240) );
  XOR U487 ( .A(x[91]), .B(y[91]), .Z(n238) );
  XNOR U488 ( .A(x[71]), .B(y[71]), .Z(n239) );
  XOR U489 ( .A(n238), .B(n239), .Z(n241) );
  XOR U490 ( .A(n240), .B(n241), .Z(n206) );
  XOR U491 ( .A(n208), .B(n206), .Z(n153) );
  XOR U492 ( .A(n207), .B(n153), .Z(n409) );
  XOR U493 ( .A(n410), .B(n409), .Z(n411) );
  XOR U494 ( .A(n412), .B(n411), .Z(n156) );
  XOR U495 ( .A(n155), .B(n156), .Z(n154) );
  XNOR U496 ( .A(n157), .B(n154), .Z(o[0]) );
  OR U497 ( .A(n166), .B(n164), .Z(n170) );
  ANDN U498 ( .B(n166), .A(n165), .Z(n168) );
  NANDN U499 ( .A(n168), .B(n167), .Z(n169) );
  AND U500 ( .A(n170), .B(n169), .Z(n437) );
  XOR U501 ( .A(n439), .B(n437), .Z(n171) );
  XNOR U502 ( .A(n438), .B(n171), .Z(n451) );
  NANDN U503 ( .A(n181), .B(n180), .Z(n185) );
  NANDN U504 ( .A(n183), .B(n182), .Z(n184) );
  AND U505 ( .A(n185), .B(n184), .Z(n502) );
  XOR U506 ( .A(n503), .B(n502), .Z(n186) );
  XOR U507 ( .A(n504), .B(n186), .Z(n544) );
  NANDN U508 ( .A(n188), .B(n187), .Z(n192) );
  NANDN U509 ( .A(n190), .B(n189), .Z(n191) );
  NAND U510 ( .A(n192), .B(n191), .Z(n464) );
  NANDN U511 ( .A(n194), .B(n193), .Z(n198) );
  NANDN U512 ( .A(n196), .B(n195), .Z(n197) );
  NAND U513 ( .A(n198), .B(n197), .Z(n465) );
  NANDN U514 ( .A(n200), .B(n199), .Z(n204) );
  NANDN U515 ( .A(n202), .B(n201), .Z(n203) );
  AND U516 ( .A(n204), .B(n203), .Z(n463) );
  XOR U517 ( .A(n465), .B(n463), .Z(n205) );
  XOR U518 ( .A(n464), .B(n205), .Z(n543) );
  XNOR U519 ( .A(n543), .B(n542), .Z(n209) );
  XNOR U520 ( .A(n544), .B(n209), .Z(n550) );
  NAND U521 ( .A(n211), .B(n210), .Z(n215) );
  NAND U522 ( .A(n213), .B(n212), .Z(n214) );
  AND U523 ( .A(n215), .B(n214), .Z(n466) );
  NANDN U524 ( .A(n217), .B(n216), .Z(n221) );
  NANDN U525 ( .A(n219), .B(n218), .Z(n220) );
  NAND U526 ( .A(n221), .B(n220), .Z(n468) );
  NAND U527 ( .A(n223), .B(n222), .Z(n227) );
  NAND U528 ( .A(n225), .B(n224), .Z(n226) );
  AND U529 ( .A(n227), .B(n226), .Z(n467) );
  XOR U530 ( .A(n468), .B(n467), .Z(n228) );
  XOR U531 ( .A(n466), .B(n228), .Z(n541) );
  NAND U532 ( .A(n233), .B(n232), .Z(n237) );
  NAND U533 ( .A(n235), .B(n234), .Z(n236) );
  AND U534 ( .A(n237), .B(n236), .Z(n519) );
  NANDN U535 ( .A(n239), .B(n238), .Z(n243) );
  NANDN U536 ( .A(n241), .B(n240), .Z(n242) );
  NAND U537 ( .A(n243), .B(n242), .Z(n518) );
  XOR U538 ( .A(n518), .B(oglobal[1]), .Z(n244) );
  XOR U539 ( .A(n519), .B(n244), .Z(n540) );
  IV U540 ( .A(n540), .Z(n538) );
  XOR U541 ( .A(n539), .B(n538), .Z(n245) );
  XOR U542 ( .A(n541), .B(n245), .Z(n549) );
  IV U543 ( .A(n549), .Z(n547) );
  NAND U544 ( .A(n247), .B(n246), .Z(n251) );
  NAND U545 ( .A(n249), .B(n248), .Z(n250) );
  AND U546 ( .A(n251), .B(n250), .Z(n548) );
  XOR U547 ( .A(n547), .B(n548), .Z(n252) );
  XOR U548 ( .A(n550), .B(n252), .Z(n455) );
  IV U549 ( .A(n253), .Z(n255) );
  NANDN U550 ( .A(n255), .B(n254), .Z(n259) );
  ANDN U551 ( .B(n255), .A(n254), .Z(n256) );
  OR U552 ( .A(n257), .B(n256), .Z(n258) );
  AND U553 ( .A(n259), .B(n258), .Z(n472) );
  NAND U554 ( .A(n264), .B(n263), .Z(n268) );
  NAND U555 ( .A(n266), .B(n265), .Z(n267) );
  NAND U556 ( .A(n268), .B(n267), .Z(n517) );
  NANDN U557 ( .A(n270), .B(n269), .Z(n274) );
  NAND U558 ( .A(n272), .B(n271), .Z(n273) );
  NAND U559 ( .A(n274), .B(n273), .Z(n516) );
  NAND U560 ( .A(n276), .B(n275), .Z(n280) );
  NAND U561 ( .A(n278), .B(n277), .Z(n279) );
  AND U562 ( .A(n280), .B(n279), .Z(n515) );
  XOR U563 ( .A(n516), .B(n515), .Z(n281) );
  XOR U564 ( .A(n517), .B(n281), .Z(n471) );
  IV U565 ( .A(n471), .Z(n470) );
  XOR U566 ( .A(n474), .B(n470), .Z(n282) );
  XNOR U567 ( .A(n472), .B(n282), .Z(n445) );
  NAND U568 ( .A(n284), .B(n283), .Z(n288) );
  NAND U569 ( .A(n286), .B(n285), .Z(n287) );
  AND U570 ( .A(n288), .B(n287), .Z(n513) );
  NAND U571 ( .A(n290), .B(n289), .Z(n294) );
  NAND U572 ( .A(n292), .B(n291), .Z(n293) );
  AND U573 ( .A(n294), .B(n293), .Z(n514) );
  NANDN U574 ( .A(n295), .B(oglobal[0]), .Z(n299) );
  NAND U575 ( .A(n297), .B(n296), .Z(n298) );
  NAND U576 ( .A(n299), .B(n298), .Z(n512) );
  XOR U577 ( .A(n514), .B(n512), .Z(n300) );
  XOR U578 ( .A(n513), .B(n300), .Z(n526) );
  XNOR U579 ( .A(n525), .B(n524), .Z(n527) );
  XOR U580 ( .A(n526), .B(n527), .Z(n444) );
  NANDN U581 ( .A(n312), .B(n311), .Z(n316) );
  NAND U582 ( .A(n314), .B(n313), .Z(n315) );
  AND U583 ( .A(n316), .B(n315), .Z(n500) );
  NAND U584 ( .A(n318), .B(n317), .Z(n322) );
  NANDN U585 ( .A(n320), .B(n319), .Z(n321) );
  NAND U586 ( .A(n322), .B(n321), .Z(n499) );
  XOR U587 ( .A(n500), .B(n499), .Z(n323) );
  XNOR U588 ( .A(n501), .B(n323), .Z(n534) );
  XNOR U589 ( .A(n493), .B(n494), .Z(n496) );
  NANDN U590 ( .A(n336), .B(n335), .Z(n340) );
  NANDN U591 ( .A(n338), .B(n337), .Z(n339) );
  NAND U592 ( .A(n340), .B(n339), .Z(n461) );
  NANDN U593 ( .A(n342), .B(n341), .Z(n346) );
  NAND U594 ( .A(n344), .B(n343), .Z(n345) );
  NAND U595 ( .A(n346), .B(n345), .Z(n462) );
  XOR U596 ( .A(n462), .B(n460), .Z(n351) );
  XOR U597 ( .A(n461), .B(n351), .Z(n495) );
  XOR U598 ( .A(n496), .B(n495), .Z(n532) );
  IV U599 ( .A(n532), .Z(n531) );
  XOR U600 ( .A(n533), .B(n531), .Z(n352) );
  XOR U601 ( .A(n534), .B(n352), .Z(n443) );
  NANDN U602 ( .A(n354), .B(n353), .Z(n358) );
  NANDN U603 ( .A(n356), .B(n355), .Z(n357) );
  AND U604 ( .A(n358), .B(n357), .Z(n487) );
  NANDN U605 ( .A(n360), .B(n359), .Z(n364) );
  NANDN U606 ( .A(n362), .B(n361), .Z(n363) );
  AND U607 ( .A(n364), .B(n363), .Z(n486) );
  XOR U608 ( .A(n487), .B(n486), .Z(n489) );
  NAND U609 ( .A(n366), .B(n365), .Z(n370) );
  NAND U610 ( .A(n368), .B(n367), .Z(n369) );
  AND U611 ( .A(n370), .B(n369), .Z(n488) );
  XOR U612 ( .A(n489), .B(n488), .Z(n523) );
  NANDN U613 ( .A(n372), .B(n371), .Z(n376) );
  NANDN U614 ( .A(n374), .B(n373), .Z(n375) );
  AND U615 ( .A(n376), .B(n375), .Z(n481) );
  NAND U616 ( .A(n378), .B(n377), .Z(n382) );
  NAND U617 ( .A(n380), .B(n379), .Z(n381) );
  AND U618 ( .A(n382), .B(n381), .Z(n480) );
  XOR U619 ( .A(n481), .B(n480), .Z(n483) );
  NAND U620 ( .A(n384), .B(n383), .Z(n388) );
  NAND U621 ( .A(n386), .B(n385), .Z(n387) );
  AND U622 ( .A(n388), .B(n387), .Z(n482) );
  XNOR U623 ( .A(n483), .B(n482), .Z(n522) );
  NANDN U624 ( .A(n390), .B(n389), .Z(n394) );
  NANDN U625 ( .A(n392), .B(n391), .Z(n393) );
  AND U626 ( .A(n394), .B(n393), .Z(n477) );
  NANDN U627 ( .A(n396), .B(n395), .Z(n400) );
  NANDN U628 ( .A(n398), .B(n397), .Z(n399) );
  NAND U629 ( .A(n400), .B(n399), .Z(n479) );
  NAND U630 ( .A(n402), .B(n401), .Z(n406) );
  NAND U631 ( .A(n404), .B(n403), .Z(n405) );
  AND U632 ( .A(n406), .B(n405), .Z(n478) );
  XOR U633 ( .A(n479), .B(n478), .Z(n407) );
  XNOR U634 ( .A(n477), .B(n407), .Z(n521) );
  XOR U635 ( .A(n522), .B(n521), .Z(n408) );
  XNOR U636 ( .A(n523), .B(n408), .Z(n442) );
  NAND U637 ( .A(n410), .B(n409), .Z(n414) );
  NAND U638 ( .A(n412), .B(n411), .Z(n413) );
  NAND U639 ( .A(n414), .B(n413), .Z(n440) );
  OR U640 ( .A(n416), .B(n415), .Z(n420) );
  AND U641 ( .A(n416), .B(n415), .Z(n417) );
  OR U642 ( .A(n418), .B(n417), .Z(n419) );
  AND U643 ( .A(n420), .B(n419), .Z(n509) );
  IV U644 ( .A(n421), .Z(n422) );
  NANDN U645 ( .A(n423), .B(n422), .Z(n427) );
  ANDN U646 ( .B(n423), .A(n422), .Z(n424) );
  OR U647 ( .A(n425), .B(n424), .Z(n426) );
  AND U648 ( .A(n427), .B(n426), .Z(n511) );
  OR U649 ( .A(n429), .B(n428), .Z(n433) );
  AND U650 ( .A(n429), .B(n428), .Z(n431) );
  OR U651 ( .A(n431), .B(n430), .Z(n432) );
  AND U652 ( .A(n433), .B(n432), .Z(n510) );
  XOR U653 ( .A(n511), .B(n510), .Z(n434) );
  XNOR U654 ( .A(n509), .B(n434), .Z(n441) );
  XNOR U655 ( .A(n440), .B(n441), .Z(n435) );
  XNOR U656 ( .A(n442), .B(n435), .Z(n456) );
  XOR U657 ( .A(n457), .B(n456), .Z(n448) );
  IV U658 ( .A(n448), .Z(n447) );
  XOR U659 ( .A(n451), .B(n447), .Z(n436) );
  XNOR U660 ( .A(n449), .B(n436), .Z(o[1]) );
  XNOR U661 ( .A(n586), .B(n585), .Z(n446) );
  XOR U662 ( .A(n584), .B(n446), .Z(n596) );
  IV U663 ( .A(n596), .Z(n595) );
  OR U664 ( .A(n449), .B(n447), .Z(n453) );
  ANDN U665 ( .B(n449), .A(n448), .Z(n450) );
  OR U666 ( .A(n451), .B(n450), .Z(n452) );
  AND U667 ( .A(n453), .B(n452), .Z(n597) );
  NANDN U668 ( .A(n455), .B(n454), .Z(n459) );
  NAND U669 ( .A(n457), .B(n456), .Z(n458) );
  NAND U670 ( .A(n459), .B(n458), .Z(n589) );
  IV U671 ( .A(n589), .Z(n588) );
  XOR U672 ( .A(n558), .B(n557), .Z(n469) );
  XOR U673 ( .A(n556), .B(n469), .Z(n571) );
  OR U674 ( .A(n472), .B(n470), .Z(n476) );
  ANDN U675 ( .B(n472), .A(n471), .Z(n473) );
  OR U676 ( .A(n474), .B(n473), .Z(n475) );
  AND U677 ( .A(n476), .B(n475), .Z(n573) );
  NAND U678 ( .A(n481), .B(n480), .Z(n485) );
  NAND U679 ( .A(n483), .B(n482), .Z(n484) );
  AND U680 ( .A(n485), .B(n484), .Z(n567) );
  NAND U681 ( .A(n487), .B(n486), .Z(n491) );
  NAND U682 ( .A(n489), .B(n488), .Z(n490) );
  AND U683 ( .A(n491), .B(n490), .Z(n566) );
  XOR U684 ( .A(n567), .B(n566), .Z(n568) );
  XOR U685 ( .A(n569), .B(n568), .Z(n572) );
  XNOR U686 ( .A(n573), .B(n572), .Z(n492) );
  XOR U687 ( .A(n571), .B(n492), .Z(n554) );
  NANDN U688 ( .A(n494), .B(n493), .Z(n498) );
  NAND U689 ( .A(n496), .B(n495), .Z(n497) );
  AND U690 ( .A(n498), .B(n497), .Z(n565) );
  NANDN U691 ( .A(n503), .B(n502), .Z(n507) );
  ANDN U692 ( .B(n503), .A(n502), .Z(n505) );
  NANDN U693 ( .A(n505), .B(n504), .Z(n506) );
  AND U694 ( .A(n507), .B(n506), .Z(n564) );
  XNOR U695 ( .A(n563), .B(n564), .Z(n508) );
  XNOR U696 ( .A(n565), .B(n508), .Z(n581) );
  XNOR U697 ( .A(n555), .B(oglobal[2]), .Z(n559) );
  XNOR U698 ( .A(n561), .B(n560), .Z(n520) );
  XOR U699 ( .A(n559), .B(n520), .Z(n582) );
  OR U700 ( .A(n525), .B(n524), .Z(n529) );
  NANDN U701 ( .A(n527), .B(n526), .Z(n528) );
  NAND U702 ( .A(n529), .B(n528), .Z(n578) );
  XOR U703 ( .A(n580), .B(n578), .Z(n530) );
  XNOR U704 ( .A(n579), .B(n530), .Z(n553) );
  OR U705 ( .A(n533), .B(n531), .Z(n537) );
  ANDN U706 ( .B(n533), .A(n532), .Z(n535) );
  OR U707 ( .A(n535), .B(n534), .Z(n536) );
  AND U708 ( .A(n537), .B(n536), .Z(n576) );
  XNOR U709 ( .A(n577), .B(n575), .Z(n545) );
  XOR U710 ( .A(n576), .B(n545), .Z(n552) );
  XOR U711 ( .A(n553), .B(n552), .Z(n546) );
  XOR U712 ( .A(n554), .B(n546), .Z(n591) );
  XNOR U713 ( .A(n597), .B(n598), .Z(n551) );
  XOR U714 ( .A(n595), .B(n551), .Z(o[2]) );
  ANDN U715 ( .B(oglobal[2]), .A(n555), .Z(n613) );
  XOR U716 ( .A(oglobal[3]), .B(n613), .Z(n617) );
  IV U717 ( .A(n617), .Z(n619) );
  XNOR U718 ( .A(n621), .B(n618), .Z(n562) );
  XOR U719 ( .A(n619), .B(n562), .Z(n616) );
  XOR U720 ( .A(n615), .B(n614), .Z(n570) );
  XOR U721 ( .A(n616), .B(n570), .Z(n631) );
  XOR U722 ( .A(n631), .B(n632), .Z(n574) );
  XNOR U723 ( .A(n633), .B(n574), .Z(n612) );
  XOR U724 ( .A(n626), .B(n625), .Z(n627) );
  XOR U725 ( .A(n628), .B(n627), .Z(n610) );
  XOR U726 ( .A(n610), .B(n611), .Z(n587) );
  XOR U727 ( .A(n612), .B(n587), .Z(n604) );
  IV U728 ( .A(n604), .Z(n603) );
  OR U729 ( .A(n590), .B(n588), .Z(n594) );
  ANDN U730 ( .B(n590), .A(n589), .Z(n592) );
  NANDN U731 ( .A(n592), .B(n591), .Z(n593) );
  AND U732 ( .A(n594), .B(n593), .Z(n607) );
  OR U733 ( .A(n597), .B(n595), .Z(n601) );
  ANDN U734 ( .B(n597), .A(n596), .Z(n599) );
  OR U735 ( .A(n599), .B(n598), .Z(n600) );
  AND U736 ( .A(n601), .B(n600), .Z(n605) );
  XNOR U737 ( .A(n607), .B(n605), .Z(n602) );
  XOR U738 ( .A(n603), .B(n602), .Z(o[3]) );
  OR U739 ( .A(n605), .B(n603), .Z(n609) );
  ANDN U740 ( .B(n605), .A(n604), .Z(n606) );
  OR U741 ( .A(n607), .B(n606), .Z(n608) );
  AND U742 ( .A(n609), .B(n608), .Z(n645) );
  XOR U743 ( .A(n636), .B(oglobal[4]), .Z(n638) );
  NANDN U744 ( .A(n617), .B(n618), .Z(n623) );
  NOR U745 ( .A(n619), .B(n618), .Z(n620) );
  OR U746 ( .A(n621), .B(n620), .Z(n622) );
  AND U747 ( .A(n623), .B(n622), .Z(n637) );
  XNOR U748 ( .A(n639), .B(n637), .Z(n624) );
  XOR U749 ( .A(n638), .B(n624), .Z(n641) );
  OR U750 ( .A(n626), .B(n625), .Z(n630) );
  NANDN U751 ( .A(n628), .B(n627), .Z(n629) );
  AND U752 ( .A(n630), .B(n629), .Z(n640) );
  XNOR U753 ( .A(n640), .B(n642), .Z(n634) );
  XOR U754 ( .A(n641), .B(n634), .Z(n644) );
  IV U755 ( .A(n644), .Z(n643) );
  XOR U756 ( .A(n647), .B(n643), .Z(n635) );
  XNOR U757 ( .A(n645), .B(n635), .Z(o[4]) );
  AND U758 ( .A(n636), .B(oglobal[4]), .Z(n654) );
  XOR U759 ( .A(oglobal[5]), .B(n654), .Z(n656) );
  XNOR U760 ( .A(n656), .B(n655), .Z(n653) );
  OR U761 ( .A(n645), .B(n643), .Z(n649) );
  ANDN U762 ( .B(n645), .A(n644), .Z(n646) );
  OR U763 ( .A(n647), .B(n646), .Z(n648) );
  AND U764 ( .A(n649), .B(n648), .Z(n651) );
  XOR U765 ( .A(n652), .B(n651), .Z(n650) );
  XNOR U766 ( .A(n653), .B(n650), .Z(o[5]) );
  NAND U767 ( .A(n654), .B(oglobal[5]), .Z(n658) );
  NAND U768 ( .A(n656), .B(n655), .Z(n657) );
  NAND U769 ( .A(n658), .B(n657), .Z(n660) );
  XOR U770 ( .A(n661), .B(n660), .Z(n659) );
  XNOR U771 ( .A(oglobal[6]), .B(n659), .Z(o[6]) );
  XNOR U772 ( .A(n662), .B(oglobal[7]), .Z(o[7]) );
  ANDN U773 ( .B(oglobal[7]), .A(n662), .Z(n663) );
  XOR U774 ( .A(n663), .B(oglobal[8]), .Z(o[8]) );
  NAND U775 ( .A(n663), .B(oglobal[8]), .Z(n664) );
  XNOR U776 ( .A(oglobal[9]), .B(n664), .Z(o[9]) );
  NANDN U777 ( .A(n664), .B(oglobal[9]), .Z(n665) );
  XNOR U778 ( .A(oglobal[10]), .B(n665), .Z(o[10]) );
endmodule

