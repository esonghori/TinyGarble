
module mult_N128_CC2 ( clk, rst, a, b, c );
  input [127:0] a;
  input [63:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471;
  wire   [255:0] sreg;

  DFF \sreg_reg[191]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U67 ( .A(n13834), .B(n13833), .Z(n13840) );
  NAND U68 ( .A(n12695), .B(n12694), .Z(n1) );
  XOR U69 ( .A(n12694), .B(n12695), .Z(n2) );
  NANDN U70 ( .A(n12696), .B(n2), .Z(n3) );
  NAND U71 ( .A(n1), .B(n3), .Z(n12985) );
  NAND U72 ( .A(n13551), .B(n13549), .Z(n4) );
  XOR U73 ( .A(n13549), .B(n13551), .Z(n5) );
  NANDN U74 ( .A(n13550), .B(n5), .Z(n6) );
  NAND U75 ( .A(n4), .B(n6), .Z(n13844) );
  OR U76 ( .A(n33753), .B(n33754), .Z(n7) );
  NAND U77 ( .A(n33751), .B(n33752), .Z(n8) );
  AND U78 ( .A(n7), .B(n8), .Z(n33764) );
  NAND U79 ( .A(n38052), .B(n38053), .Z(n9) );
  NANDN U80 ( .A(n38051), .B(n38050), .Z(n10) );
  NAND U81 ( .A(n9), .B(n10), .Z(n38059) );
  OR U82 ( .A(n38182), .B(n38183), .Z(n11) );
  NANDN U83 ( .A(n38185), .B(n38184), .Z(n12) );
  NAND U84 ( .A(n11), .B(n12), .Z(n38218) );
  NAND U85 ( .A(n9713), .B(n9714), .Z(n13) );
  NANDN U86 ( .A(n9712), .B(n9711), .Z(n14) );
  NAND U87 ( .A(n13), .B(n14), .Z(n10076) );
  NAND U88 ( .A(n15219), .B(n15218), .Z(n15) );
  NANDN U89 ( .A(n15217), .B(n15216), .Z(n16) );
  AND U90 ( .A(n15), .B(n16), .Z(n15383) );
  NAND U91 ( .A(n8208), .B(n8207), .Z(n17) );
  NANDN U92 ( .A(n8206), .B(n8205), .Z(n18) );
  AND U93 ( .A(n17), .B(n18), .Z(n8402) );
  OR U94 ( .A(n16021), .B(n16022), .Z(n19) );
  NANDN U95 ( .A(n16024), .B(n16023), .Z(n20) );
  AND U96 ( .A(n19), .B(n20), .Z(n16145) );
  OR U97 ( .A(n20907), .B(n20908), .Z(n21) );
  NANDN U98 ( .A(n20910), .B(n20909), .Z(n22) );
  AND U99 ( .A(n21), .B(n22), .Z(n21278) );
  OR U100 ( .A(n23210), .B(n23211), .Z(n23) );
  NANDN U101 ( .A(n23213), .B(n23212), .Z(n24) );
  AND U102 ( .A(n23), .B(n24), .Z(n23573) );
  NAND U103 ( .A(n26925), .B(n26926), .Z(n25) );
  NANDN U104 ( .A(n26924), .B(n26923), .Z(n26) );
  NAND U105 ( .A(n25), .B(n26), .Z(n27191) );
  NAND U106 ( .A(n4536), .B(n4537), .Z(n27) );
  NANDN U107 ( .A(n4535), .B(n4534), .Z(n28) );
  NAND U108 ( .A(n27), .B(n28), .Z(n4626) );
  XNOR U109 ( .A(n7007), .B(n7008), .Z(n7010) );
  NAND U110 ( .A(n8409), .B(n8408), .Z(n29) );
  NANDN U111 ( .A(n8407), .B(n8406), .Z(n30) );
  AND U112 ( .A(n29), .B(n30), .Z(n8598) );
  NAND U113 ( .A(n12966), .B(n12965), .Z(n31) );
  NANDN U114 ( .A(n12964), .B(n12963), .Z(n32) );
  AND U115 ( .A(n31), .B(n32), .Z(n13255) );
  XNOR U116 ( .A(n14379), .B(n14378), .Z(n14380) );
  NANDN U117 ( .A(n14397), .B(n14396), .Z(n33) );
  NANDN U118 ( .A(n14395), .B(n14394), .Z(n34) );
  AND U119 ( .A(n33), .B(n34), .Z(n14425) );
  NAND U120 ( .A(n16157), .B(n16156), .Z(n35) );
  NANDN U121 ( .A(n16155), .B(n16154), .Z(n36) );
  AND U122 ( .A(n35), .B(n36), .Z(n16677) );
  NAND U123 ( .A(n21578), .B(n21579), .Z(n37) );
  NANDN U124 ( .A(n21577), .B(n21576), .Z(n38) );
  NAND U125 ( .A(n37), .B(n38), .Z(n21608) );
  NAND U126 ( .A(n22475), .B(n22476), .Z(n39) );
  NANDN U127 ( .A(n22474), .B(n22473), .Z(n40) );
  NAND U128 ( .A(n39), .B(n40), .Z(n23003) );
  NAND U129 ( .A(n25494), .B(n25493), .Z(n41) );
  NAND U130 ( .A(n25491), .B(n25492), .Z(n42) );
  NAND U131 ( .A(n41), .B(n42), .Z(n25889) );
  XNOR U132 ( .A(n26754), .B(n26753), .Z(n26755) );
  XNOR U133 ( .A(n27306), .B(n27305), .Z(n27307) );
  NAND U134 ( .A(n27692), .B(n27693), .Z(n43) );
  NANDN U135 ( .A(n27691), .B(n27690), .Z(n44) );
  NAND U136 ( .A(n43), .B(n44), .Z(n27943) );
  NAND U137 ( .A(n27709), .B(n27710), .Z(n45) );
  NANDN U138 ( .A(n27712), .B(n27711), .Z(n46) );
  NAND U139 ( .A(n45), .B(n46), .Z(n27957) );
  XNOR U140 ( .A(n33004), .B(n33003), .Z(n32999) );
  NAND U141 ( .A(n2974), .B(n2975), .Z(n47) );
  NANDN U142 ( .A(n2977), .B(n2976), .Z(n48) );
  NAND U143 ( .A(n47), .B(n48), .Z(n3129) );
  NAND U144 ( .A(n6543), .B(n6544), .Z(n49) );
  NANDN U145 ( .A(n6542), .B(n6541), .Z(n50) );
  NAND U146 ( .A(n49), .B(n50), .Z(n6679) );
  XNOR U147 ( .A(n11266), .B(n11265), .Z(n11272) );
  NAND U148 ( .A(n27857), .B(n27858), .Z(n51) );
  NANDN U149 ( .A(n27856), .B(n27855), .Z(n52) );
  NAND U150 ( .A(n51), .B(n52), .Z(n28183) );
  NAND U151 ( .A(n27976), .B(n27977), .Z(n53) );
  NANDN U152 ( .A(n27975), .B(n27974), .Z(n54) );
  NAND U153 ( .A(n53), .B(n54), .Z(n28210) );
  XNOR U154 ( .A(n29303), .B(n29304), .Z(n29306) );
  NANDN U155 ( .A(n34116), .B(n34115), .Z(n55) );
  NANDN U156 ( .A(n34118), .B(n34117), .Z(n56) );
  NAND U157 ( .A(n55), .B(n56), .Z(n34233) );
  XNOR U158 ( .A(n34243), .B(n34244), .Z(n34176) );
  OR U159 ( .A(n36953), .B(n36954), .Z(n57) );
  NAND U160 ( .A(n36952), .B(n36951), .Z(n58) );
  NAND U161 ( .A(n57), .B(n58), .Z(n37002) );
  NAND U162 ( .A(n1982), .B(n1983), .Z(n59) );
  NANDN U163 ( .A(n1981), .B(n1980), .Z(n60) );
  NAND U164 ( .A(n59), .B(n60), .Z(n2009) );
  NANDN U165 ( .A(n23589), .B(n23588), .Z(n61) );
  NANDN U166 ( .A(n23591), .B(n23590), .Z(n62) );
  NAND U167 ( .A(n61), .B(n62), .Z(n23886) );
  XNOR U168 ( .A(n28753), .B(n28754), .Z(n28756) );
  NANDN U169 ( .A(n34934), .B(n34933), .Z(n63) );
  NANDN U170 ( .A(n34936), .B(n34935), .Z(n64) );
  NAND U171 ( .A(n63), .B(n64), .Z(n35105) );
  NAND U172 ( .A(n12987), .B(n12988), .Z(n65) );
  NANDN U173 ( .A(n12986), .B(n12985), .Z(n66) );
  NAND U174 ( .A(n65), .B(n66), .Z(n12995) );
  NAND U175 ( .A(n13845), .B(n13846), .Z(n67) );
  NANDN U176 ( .A(n13844), .B(n13843), .Z(n68) );
  NAND U177 ( .A(n67), .B(n68), .Z(n13853) );
  NAND U178 ( .A(n29349), .B(n29350), .Z(n69) );
  NANDN U179 ( .A(n29348), .B(n29347), .Z(n70) );
  NAND U180 ( .A(n69), .B(n70), .Z(n29619) );
  NAND U181 ( .A(n35146), .B(n35145), .Z(n71) );
  NANDN U182 ( .A(n35144), .B(n35143), .Z(n72) );
  NAND U183 ( .A(n71), .B(n72), .Z(n35413) );
  NAND U184 ( .A(n35724), .B(n35725), .Z(n73) );
  NANDN U185 ( .A(n35723), .B(n35722), .Z(n74) );
  NAND U186 ( .A(n73), .B(n74), .Z(n35898) );
  XNOR U187 ( .A(n38156), .B(n38157), .Z(n38149) );
  NAND U188 ( .A(n38147), .B(n38146), .Z(n75) );
  NANDN U189 ( .A(n38145), .B(n38144), .Z(n76) );
  AND U190 ( .A(n75), .B(n76), .Z(n38183) );
  NAND U191 ( .A(n32669), .B(n32668), .Z(n77) );
  NANDN U192 ( .A(n32667), .B(n32666), .Z(n78) );
  AND U193 ( .A(n77), .B(n78), .Z(n32675) );
  NAND U194 ( .A(n36220), .B(n36221), .Z(n79) );
  NANDN U195 ( .A(n36219), .B(n36218), .Z(n80) );
  NAND U196 ( .A(n79), .B(n80), .Z(n36476) );
  NAND U197 ( .A(n37997), .B(n37998), .Z(n81) );
  NANDN U198 ( .A(n37996), .B(n37995), .Z(n82) );
  NAND U199 ( .A(n81), .B(n82), .Z(n38112) );
  XOR U200 ( .A(n33957), .B(n33955), .Z(n83) );
  NAND U201 ( .A(n83), .B(n33956), .Z(n84) );
  NAND U202 ( .A(n33957), .B(n33955), .Z(n85) );
  AND U203 ( .A(n84), .B(n85), .Z(n33961) );
  XOR U204 ( .A(n38263), .B(n38262), .Z(n86) );
  NAND U205 ( .A(n86), .B(n38261), .Z(n87) );
  NAND U206 ( .A(n38263), .B(n38262), .Z(n88) );
  AND U207 ( .A(n87), .B(n88), .Z(n38270) );
  XOR U208 ( .A(n38385), .B(n38384), .Z(n89) );
  NANDN U209 ( .A(n38383), .B(n89), .Z(n90) );
  NAND U210 ( .A(n38385), .B(n38384), .Z(n91) );
  AND U211 ( .A(n90), .B(n91), .Z(n38416) );
  XNOR U212 ( .A(n12895), .B(n12896), .Z(n12898) );
  XNOR U213 ( .A(n18912), .B(n18913), .Z(n18915) );
  XNOR U214 ( .A(n19763), .B(n19764), .Z(n19766) );
  XNOR U215 ( .A(n24095), .B(n24096), .Z(n24098) );
  XNOR U216 ( .A(n24583), .B(n24584), .Z(n24586) );
  XNOR U217 ( .A(n25940), .B(n25941), .Z(n25943) );
  NAND U218 ( .A(n9772), .B(n9771), .Z(n92) );
  NANDN U219 ( .A(n9770), .B(n9769), .Z(n93) );
  AND U220 ( .A(n92), .B(n93), .Z(n10024) );
  XNOR U221 ( .A(n10541), .B(n10540), .Z(n10542) );
  NAND U222 ( .A(n12915), .B(n12916), .Z(n94) );
  NANDN U223 ( .A(n12914), .B(n12913), .Z(n95) );
  NAND U224 ( .A(n94), .B(n95), .Z(n13119) );
  NAND U225 ( .A(n13345), .B(n13344), .Z(n96) );
  NANDN U226 ( .A(n13343), .B(n13342), .Z(n97) );
  AND U227 ( .A(n96), .B(n97), .Z(n13634) );
  NAND U228 ( .A(n15336), .B(n15337), .Z(n98) );
  NANDN U229 ( .A(n15339), .B(n15338), .Z(n99) );
  NAND U230 ( .A(n98), .B(n99), .Z(n15608) );
  NAND U231 ( .A(n17527), .B(n17528), .Z(n100) );
  NANDN U232 ( .A(n17530), .B(n17529), .Z(n101) );
  NAND U233 ( .A(n100), .B(n101), .Z(n17607) );
  NAND U234 ( .A(n18489), .B(n18488), .Z(n102) );
  NANDN U235 ( .A(n18487), .B(n18486), .Z(n103) );
  AND U236 ( .A(n102), .B(n103), .Z(n18961) );
  NAND U237 ( .A(n22356), .B(n22355), .Z(n104) );
  NANDN U238 ( .A(n22354), .B(n22353), .Z(n105) );
  AND U239 ( .A(n104), .B(n105), .Z(n22701) );
  NAND U240 ( .A(n24847), .B(n24846), .Z(n106) );
  NANDN U241 ( .A(n24845), .B(n24844), .Z(n107) );
  AND U242 ( .A(n106), .B(n107), .Z(n25297) );
  NAND U243 ( .A(n26406), .B(n26407), .Z(n108) );
  NANDN U244 ( .A(n26409), .B(n26408), .Z(n109) );
  NAND U245 ( .A(n108), .B(n109), .Z(n26613) );
  NANDN U246 ( .A(n986), .B(b[40]), .Z(n110) );
  AND U247 ( .A(b[41]), .B(n110), .Z(n111) );
  XNOR U248 ( .A(b[40]), .B(n986), .Z(n112) );
  NAND U249 ( .A(n112), .B(b[39]), .Z(n113) );
  NAND U250 ( .A(n111), .B(n113), .Z(n5009) );
  XNOR U251 ( .A(n6023), .B(n6024), .Z(n6026) );
  OR U252 ( .A(n6196), .B(n6197), .Z(n6451) );
  NAND U253 ( .A(n7126), .B(n7127), .Z(n114) );
  NANDN U254 ( .A(n7125), .B(n7124), .Z(n115) );
  NAND U255 ( .A(n114), .B(n115), .Z(n7365) );
  XNOR U256 ( .A(n8362), .B(n8363), .Z(n8365) );
  XOR U257 ( .A(n8332), .B(n8333), .Z(n8334) );
  NAND U258 ( .A(n9534), .B(n9535), .Z(n116) );
  NANDN U259 ( .A(n9533), .B(n9532), .Z(n117) );
  NAND U260 ( .A(n116), .B(n117), .Z(n9637) );
  NAND U261 ( .A(n10337), .B(n10338), .Z(n118) );
  NANDN U262 ( .A(n10336), .B(n10335), .Z(n119) );
  NAND U263 ( .A(n118), .B(n119), .Z(n10695) );
  NAND U264 ( .A(n10757), .B(n10756), .Z(n120) );
  NANDN U265 ( .A(n10755), .B(n10754), .Z(n121) );
  AND U266 ( .A(n120), .B(n121), .Z(n11015) );
  OR U267 ( .A(n11052), .B(n11053), .Z(n122) );
  NANDN U268 ( .A(n11055), .B(n11054), .Z(n123) );
  AND U269 ( .A(n122), .B(n123), .Z(n11542) );
  OR U270 ( .A(n11510), .B(n11511), .Z(n124) );
  NANDN U271 ( .A(n11513), .B(n11512), .Z(n125) );
  AND U272 ( .A(n124), .B(n125), .Z(n11815) );
  OR U273 ( .A(n12635), .B(n12636), .Z(n126) );
  NANDN U274 ( .A(n12638), .B(n12637), .Z(n127) );
  AND U275 ( .A(n126), .B(n127), .Z(n12954) );
  OR U276 ( .A(n12876), .B(n12877), .Z(n128) );
  NANDN U277 ( .A(n12879), .B(n12878), .Z(n129) );
  AND U278 ( .A(n128), .B(n129), .Z(n13243) );
  OR U279 ( .A(n14066), .B(n14067), .Z(n130) );
  NANDN U280 ( .A(n14069), .B(n14068), .Z(n131) );
  AND U281 ( .A(n130), .B(n131), .Z(n14384) );
  OR U282 ( .A(n14326), .B(n14327), .Z(n132) );
  NANDN U283 ( .A(n14329), .B(n14328), .Z(n133) );
  NAND U284 ( .A(n132), .B(n133), .Z(n14670) );
  NAND U285 ( .A(n14548), .B(n14547), .Z(n134) );
  NANDN U286 ( .A(n14546), .B(n14545), .Z(n135) );
  AND U287 ( .A(n134), .B(n135), .Z(n14713) );
  OR U288 ( .A(n14445), .B(n14446), .Z(n136) );
  NAND U289 ( .A(n14443), .B(n14444), .Z(n137) );
  AND U290 ( .A(n136), .B(n137), .Z(n14948) );
  OR U291 ( .A(n14789), .B(n14790), .Z(n138) );
  NANDN U292 ( .A(n14792), .B(n14791), .Z(n139) );
  AND U293 ( .A(n138), .B(n139), .Z(n15249) );
  OR U294 ( .A(n16309), .B(n16310), .Z(n140) );
  NANDN U295 ( .A(n16312), .B(n16311), .Z(n141) );
  AND U296 ( .A(n140), .B(n141), .Z(n16660) );
  OR U297 ( .A(n16443), .B(n16444), .Z(n142) );
  NAND U298 ( .A(n16441), .B(n16442), .Z(n143) );
  AND U299 ( .A(n142), .B(n143), .Z(n16956) );
  OR U300 ( .A(n16797), .B(n16798), .Z(n144) );
  NANDN U301 ( .A(n16800), .B(n16799), .Z(n145) );
  AND U302 ( .A(n144), .B(n145), .Z(n17260) );
  OR U303 ( .A(n17775), .B(n17776), .Z(n146) );
  NANDN U304 ( .A(n17778), .B(n17777), .Z(n147) );
  NAND U305 ( .A(n146), .B(n147), .Z(n17888) );
  OR U306 ( .A(n22381), .B(n22382), .Z(n148) );
  NANDN U307 ( .A(n22384), .B(n22383), .Z(n149) );
  AND U308 ( .A(n148), .B(n149), .Z(n22463) );
  OR U309 ( .A(n22789), .B(n22790), .Z(n150) );
  NANDN U310 ( .A(n22792), .B(n22791), .Z(n151) );
  AND U311 ( .A(n150), .B(n151), .Z(n23272) );
  OR U312 ( .A(n25882), .B(n25883), .Z(n152) );
  NANDN U313 ( .A(n25885), .B(n25884), .Z(n153) );
  AND U314 ( .A(n152), .B(n153), .Z(n26022) );
  XNOR U315 ( .A(n27299), .B(n27300), .Z(n27302) );
  NAND U316 ( .A(n27506), .B(n27507), .Z(n154) );
  NANDN U317 ( .A(n27505), .B(n27504), .Z(n155) );
  NAND U318 ( .A(n154), .B(n155), .Z(n27645) );
  XOR U319 ( .A(n30267), .B(n30268), .Z(n30217) );
  NAND U320 ( .A(n2739), .B(n2738), .Z(n156) );
  NANDN U321 ( .A(n2737), .B(n2736), .Z(n157) );
  AND U322 ( .A(n156), .B(n157), .Z(n2835) );
  NAND U323 ( .A(n4131), .B(n4132), .Z(n158) );
  NANDN U324 ( .A(n4134), .B(n4133), .Z(n159) );
  NAND U325 ( .A(n158), .B(n159), .Z(n4325) );
  NAND U326 ( .A(n5176), .B(n5177), .Z(n160) );
  NANDN U327 ( .A(n5175), .B(n5174), .Z(n161) );
  NAND U328 ( .A(n160), .B(n161), .Z(n5511) );
  XOR U329 ( .A(n7001), .B(n7002), .Z(n7003) );
  NAND U330 ( .A(n6413), .B(n6414), .Z(n162) );
  NANDN U331 ( .A(n6412), .B(n6411), .Z(n163) );
  NAND U332 ( .A(n162), .B(n163), .Z(n6669) );
  NAND U333 ( .A(n7120), .B(n7121), .Z(n164) );
  NANDN U334 ( .A(n7123), .B(n7122), .Z(n165) );
  NAND U335 ( .A(n164), .B(n165), .Z(n7288) );
  OR U336 ( .A(n7090), .B(n7089), .Z(n166) );
  NAND U337 ( .A(n7092), .B(n7091), .Z(n167) );
  NAND U338 ( .A(n166), .B(n167), .Z(n7282) );
  NAND U339 ( .A(n7377), .B(n7376), .Z(n168) );
  NANDN U340 ( .A(n7375), .B(n7374), .Z(n169) );
  AND U341 ( .A(n168), .B(n169), .Z(n7651) );
  XNOR U342 ( .A(n7536), .B(n7537), .Z(n7647) );
  NANDN U343 ( .A(n7782), .B(n7781), .Z(n170) );
  NANDN U344 ( .A(n7780), .B(n7779), .Z(n171) );
  AND U345 ( .A(n170), .B(n171), .Z(n8216) );
  NAND U346 ( .A(n8404), .B(n8405), .Z(n172) );
  NANDN U347 ( .A(n8403), .B(n8402), .Z(n173) );
  NAND U348 ( .A(n172), .B(n173), .Z(n8597) );
  NAND U349 ( .A(n11316), .B(n11317), .Z(n174) );
  NANDN U350 ( .A(n11315), .B(n11314), .Z(n175) );
  NAND U351 ( .A(n174), .B(n175), .Z(n11583) );
  NAND U352 ( .A(n11830), .B(n11829), .Z(n176) );
  NANDN U353 ( .A(n11828), .B(n11827), .Z(n177) );
  AND U354 ( .A(n176), .B(n177), .Z(n12115) );
  NANDN U355 ( .A(n11883), .B(n11882), .Z(n178) );
  NANDN U356 ( .A(n11881), .B(n11880), .Z(n179) );
  AND U357 ( .A(n178), .B(n179), .Z(n12406) );
  XNOR U358 ( .A(n12689), .B(n12688), .Z(n12690) );
  NAND U359 ( .A(n12681), .B(n12680), .Z(n180) );
  NANDN U360 ( .A(n12679), .B(n12678), .Z(n181) );
  NAND U361 ( .A(n180), .B(n181), .Z(n12725) );
  NANDN U362 ( .A(n12960), .B(n12959), .Z(n182) );
  NANDN U363 ( .A(n12962), .B(n12961), .Z(n183) );
  NAND U364 ( .A(n182), .B(n183), .Z(n13256) );
  XOR U365 ( .A(n13543), .B(n13544), .Z(n13545) );
  NANDN U366 ( .A(n13830), .B(n13829), .Z(n184) );
  NANDN U367 ( .A(n13828), .B(n13827), .Z(n185) );
  AND U368 ( .A(n184), .B(n185), .Z(n14112) );
  NAND U369 ( .A(n13995), .B(n13994), .Z(n186) );
  NAND U370 ( .A(n13992), .B(n13993), .Z(n187) );
  NAND U371 ( .A(n186), .B(n187), .Z(n14381) );
  NAND U372 ( .A(n14392), .B(n14393), .Z(n188) );
  NANDN U373 ( .A(n14391), .B(n14390), .Z(n189) );
  NAND U374 ( .A(n188), .B(n189), .Z(n14426) );
  XOR U375 ( .A(n14930), .B(n14931), .Z(n14932) );
  XOR U376 ( .A(n15506), .B(n15507), .Z(n15508) );
  NAND U377 ( .A(n15261), .B(n15260), .Z(n190) );
  NAND U378 ( .A(n15258), .B(n15259), .Z(n191) );
  NAND U379 ( .A(n190), .B(n191), .Z(n15531) );
  NAND U380 ( .A(n15828), .B(n15829), .Z(n192) );
  NANDN U381 ( .A(n15827), .B(n15826), .Z(n193) );
  NAND U382 ( .A(n192), .B(n193), .Z(n15868) );
  NANDN U383 ( .A(n16151), .B(n16150), .Z(n194) );
  NANDN U384 ( .A(n16153), .B(n16152), .Z(n195) );
  NAND U385 ( .A(n194), .B(n195), .Z(n16676) );
  XOR U386 ( .A(n16938), .B(n16939), .Z(n16940) );
  NANDN U387 ( .A(n17275), .B(n17274), .Z(n196) );
  NANDN U388 ( .A(n17273), .B(n17272), .Z(n197) );
  AND U389 ( .A(n196), .B(n197), .Z(n17543) );
  XOR U390 ( .A(n18409), .B(n18410), .Z(n18411) );
  NANDN U391 ( .A(n18400), .B(n18399), .Z(n198) );
  NANDN U392 ( .A(n18402), .B(n18401), .Z(n199) );
  NAND U393 ( .A(n198), .B(n199), .Z(n18690) );
  NANDN U394 ( .A(n19264), .B(n19263), .Z(n200) );
  NANDN U395 ( .A(n19262), .B(n19261), .Z(n201) );
  AND U396 ( .A(n200), .B(n201), .Z(n19304) );
  NAND U397 ( .A(n20126), .B(n20125), .Z(n202) );
  NANDN U398 ( .A(n20124), .B(n20123), .Z(n203) );
  AND U399 ( .A(n202), .B(n203), .Z(n20422) );
  XNOR U400 ( .A(n21273), .B(n21272), .Z(n21274) );
  NANDN U401 ( .A(n21293), .B(n21292), .Z(n204) );
  NANDN U402 ( .A(n21291), .B(n21290), .Z(n205) );
  AND U403 ( .A(n204), .B(n205), .Z(n21324) );
  NANDN U404 ( .A(n21573), .B(n21572), .Z(n206) );
  NANDN U405 ( .A(n21575), .B(n21574), .Z(n207) );
  NAND U406 ( .A(n206), .B(n207), .Z(n21607) );
  NAND U407 ( .A(n21860), .B(n21859), .Z(n208) );
  NANDN U408 ( .A(n21858), .B(n21857), .Z(n209) );
  AND U409 ( .A(n208), .B(n209), .Z(n22138) );
  NAND U410 ( .A(n22130), .B(n22129), .Z(n210) );
  NANDN U411 ( .A(n22128), .B(n22127), .Z(n211) );
  AND U412 ( .A(n210), .B(n211), .Z(n22179) );
  NAND U413 ( .A(n22427), .B(n22426), .Z(n212) );
  NANDN U414 ( .A(n22425), .B(n22424), .Z(n213) );
  NAND U415 ( .A(n212), .B(n213), .Z(n22712) );
  NANDN U416 ( .A(n22470), .B(n22469), .Z(n214) );
  NANDN U417 ( .A(n22472), .B(n22471), .Z(n215) );
  NAND U418 ( .A(n214), .B(n215), .Z(n23002) );
  XNOR U419 ( .A(n23567), .B(n23566), .Z(n23568) );
  NANDN U420 ( .A(n23579), .B(n23578), .Z(n216) );
  NANDN U421 ( .A(n23581), .B(n23580), .Z(n217) );
  NAND U422 ( .A(n216), .B(n217), .Z(n23862) );
  XNOR U423 ( .A(n24428), .B(n24427), .Z(n24429) );
  NANDN U424 ( .A(n24440), .B(n24439), .Z(n218) );
  NANDN U425 ( .A(n24442), .B(n24441), .Z(n219) );
  NAND U426 ( .A(n218), .B(n219), .Z(n24478) );
  NAND U427 ( .A(n25026), .B(n25025), .Z(n220) );
  NANDN U428 ( .A(n25024), .B(n25023), .Z(n221) );
  AND U429 ( .A(n220), .B(n221), .Z(n25329) );
  XNOR U430 ( .A(n26217), .B(n26218), .Z(n26220) );
  NAND U431 ( .A(n26359), .B(n26360), .Z(n222) );
  NANDN U432 ( .A(n26358), .B(n26357), .Z(n223) );
  NAND U433 ( .A(n222), .B(n223), .Z(n26756) );
  NAND U434 ( .A(n26805), .B(n26804), .Z(n224) );
  NANDN U435 ( .A(n26803), .B(n26802), .Z(n225) );
  AND U436 ( .A(n224), .B(n225), .Z(n27308) );
  NAND U437 ( .A(n27169), .B(n27168), .Z(n226) );
  NAND U438 ( .A(n27166), .B(n27167), .Z(n227) );
  NAND U439 ( .A(n226), .B(n227), .Z(n27592) );
  NAND U440 ( .A(n28227), .B(n28228), .Z(n228) );
  NANDN U441 ( .A(n28226), .B(n28225), .Z(n229) );
  NAND U442 ( .A(n228), .B(n229), .Z(n28565) );
  NAND U443 ( .A(n28889), .B(n28890), .Z(n230) );
  NANDN U444 ( .A(n28888), .B(n28887), .Z(n231) );
  NAND U445 ( .A(n230), .B(n231), .Z(n29134) );
  NANDN U446 ( .A(n30941), .B(n30940), .Z(n232) );
  NANDN U447 ( .A(n30943), .B(n30942), .Z(n233) );
  NAND U448 ( .A(n232), .B(n233), .Z(n31105) );
  NAND U449 ( .A(n32256), .B(n32257), .Z(n234) );
  NANDN U450 ( .A(n32255), .B(n32254), .Z(n235) );
  NAND U451 ( .A(n234), .B(n235), .Z(n32576) );
  XNOR U452 ( .A(n32701), .B(n32700), .Z(n32686) );
  XNOR U453 ( .A(n33148), .B(n33149), .Z(n33168) );
  XNOR U454 ( .A(n33649), .B(n33650), .Z(n33652) );
  NANDN U455 ( .A(n971), .B(a[0]), .Z(n236) );
  ANDN U456 ( .B(n236), .A(n972), .Z(n237) );
  XNOR U457 ( .A(a[0]), .B(n971), .Z(n238) );
  NAND U458 ( .A(n238), .B(b[14]), .Z(n239) );
  NAND U459 ( .A(n237), .B(n239), .Z(n1619) );
  NAND U460 ( .A(n2961), .B(n2962), .Z(n240) );
  NANDN U461 ( .A(n2964), .B(n2963), .Z(n241) );
  NAND U462 ( .A(n240), .B(n241), .Z(n3125) );
  NAND U463 ( .A(n3222), .B(n3221), .Z(n242) );
  NANDN U464 ( .A(n3220), .B(n3219), .Z(n243) );
  AND U465 ( .A(n242), .B(n243), .Z(n3346) );
  NAND U466 ( .A(n3482), .B(n3481), .Z(n244) );
  NANDN U467 ( .A(n3480), .B(n3479), .Z(n245) );
  NAND U468 ( .A(n244), .B(n245), .Z(n3625) );
  NAND U469 ( .A(n5268), .B(n5269), .Z(n246) );
  NANDN U470 ( .A(n5267), .B(n5266), .Z(n247) );
  NAND U471 ( .A(n246), .B(n247), .Z(n5526) );
  NAND U472 ( .A(n5057), .B(n5056), .Z(n248) );
  NANDN U473 ( .A(n5055), .B(n5054), .Z(n249) );
  AND U474 ( .A(n248), .B(n249), .Z(n5255) );
  NAND U475 ( .A(n6087), .B(n6088), .Z(n250) );
  NANDN U476 ( .A(n6086), .B(n6085), .Z(n251) );
  NAND U477 ( .A(n250), .B(n251), .Z(n6184) );
  XNOR U478 ( .A(n7067), .B(n7068), .Z(n7062) );
  NANDN U479 ( .A(n7379), .B(n7378), .Z(n252) );
  NANDN U480 ( .A(n7381), .B(n7380), .Z(n253) );
  NAND U481 ( .A(n252), .B(n253), .Z(n7724) );
  NAND U482 ( .A(n9572), .B(n9571), .Z(n254) );
  NANDN U483 ( .A(n9570), .B(n9569), .Z(n255) );
  AND U484 ( .A(n254), .B(n255), .Z(n9606) );
  XNOR U485 ( .A(n11263), .B(n11264), .Z(n11266) );
  NAND U486 ( .A(n11866), .B(n11867), .Z(n256) );
  NANDN U487 ( .A(n11865), .B(n11864), .Z(n257) );
  NAND U488 ( .A(n256), .B(n257), .Z(n12413) );
  XOR U489 ( .A(n13550), .B(n13549), .Z(n258) );
  XNOR U490 ( .A(n13551), .B(n258), .Z(n13555) );
  NAND U491 ( .A(n16160), .B(n16161), .Z(n259) );
  NANDN U492 ( .A(n16159), .B(n16158), .Z(n260) );
  NAND U493 ( .A(n259), .B(n260), .Z(n16689) );
  NAND U494 ( .A(n18745), .B(n18744), .Z(n261) );
  NAND U495 ( .A(n18742), .B(n18743), .Z(n262) );
  AND U496 ( .A(n261), .B(n262), .Z(n19278) );
  NAND U497 ( .A(n25662), .B(n25661), .Z(n263) );
  NANDN U498 ( .A(n25660), .B(n25659), .Z(n264) );
  AND U499 ( .A(n263), .B(n264), .Z(n26186) );
  XOR U500 ( .A(n27949), .B(n27948), .Z(n28181) );
  NAND U501 ( .A(n27935), .B(n27934), .Z(n265) );
  NANDN U502 ( .A(n27933), .B(n27932), .Z(n266) );
  NAND U503 ( .A(n265), .B(n266), .Z(n28455) );
  NANDN U504 ( .A(n29152), .B(n29151), .Z(n267) );
  NANDN U505 ( .A(n29154), .B(n29153), .Z(n268) );
  NAND U506 ( .A(n267), .B(n268), .Z(n29589) );
  XNOR U507 ( .A(n30415), .B(n30416), .Z(n30402) );
  NAND U508 ( .A(n30842), .B(n30841), .Z(n269) );
  NANDN U509 ( .A(n30840), .B(n30839), .Z(n270) );
  AND U510 ( .A(n269), .B(n270), .Z(n31057) );
  NAND U511 ( .A(n32868), .B(n32869), .Z(n271) );
  NANDN U512 ( .A(n32867), .B(n32866), .Z(n272) );
  NAND U513 ( .A(n271), .B(n272), .Z(n33091) );
  NANDN U514 ( .A(n32839), .B(n32838), .Z(n273) );
  NANDN U515 ( .A(n32841), .B(n32840), .Z(n274) );
  NAND U516 ( .A(n273), .B(n274), .Z(n32923) );
  NAND U517 ( .A(n32994), .B(n32995), .Z(n275) );
  NANDN U518 ( .A(n32993), .B(n32992), .Z(n276) );
  NAND U519 ( .A(n275), .B(n276), .Z(n33195) );
  NANDN U520 ( .A(n32935), .B(n32934), .Z(n277) );
  NANDN U521 ( .A(n32937), .B(n32936), .Z(n278) );
  NAND U522 ( .A(n277), .B(n278), .Z(n33204) );
  NAND U523 ( .A(n36594), .B(n36593), .Z(n279) );
  NANDN U524 ( .A(n36592), .B(n36591), .Z(n280) );
  NAND U525 ( .A(n279), .B(n280), .Z(n36702) );
  NAND U526 ( .A(n36941), .B(n36940), .Z(n281) );
  NANDN U527 ( .A(n36939), .B(n36938), .Z(n282) );
  NAND U528 ( .A(n281), .B(n282), .Z(n37003) );
  NAND U529 ( .A(n36937), .B(n36936), .Z(n283) );
  NANDN U530 ( .A(n36935), .B(n36934), .Z(n284) );
  AND U531 ( .A(n283), .B(n284), .Z(n37012) );
  XOR U532 ( .A(n37046), .B(n37047), .Z(n37050) );
  OR U533 ( .A(n3128), .B(n3129), .Z(n285) );
  NANDN U534 ( .A(n3131), .B(n3130), .Z(n286) );
  NAND U535 ( .A(n285), .B(n286), .Z(n3296) );
  NAND U536 ( .A(n4099), .B(n4098), .Z(n287) );
  NANDN U537 ( .A(n4097), .B(n4096), .Z(n288) );
  AND U538 ( .A(n287), .B(n288), .Z(n4400) );
  NAND U539 ( .A(n4612), .B(n4613), .Z(n289) );
  NANDN U540 ( .A(n4611), .B(n4610), .Z(n290) );
  NAND U541 ( .A(n289), .B(n290), .Z(n4784) );
  NANDN U542 ( .A(n6680), .B(n6679), .Z(n291) );
  NANDN U543 ( .A(n6682), .B(n6681), .Z(n292) );
  NAND U544 ( .A(n291), .B(n292), .Z(n6822) );
  OR U545 ( .A(n9295), .B(n9296), .Z(n293) );
  NAND U546 ( .A(n9293), .B(n9294), .Z(n294) );
  AND U547 ( .A(n293), .B(n294), .Z(n9319) );
  NAND U548 ( .A(n9517), .B(n9516), .Z(n295) );
  NANDN U549 ( .A(n9519), .B(n9518), .Z(n296) );
  NAND U550 ( .A(n295), .B(n296), .Z(n9602) );
  NANDN U551 ( .A(n16975), .B(n16974), .Z(n297) );
  NANDN U552 ( .A(n16977), .B(n16976), .Z(n298) );
  NAND U553 ( .A(n297), .B(n298), .Z(n17001) );
  NAND U554 ( .A(n17874), .B(n17875), .Z(n299) );
  NANDN U555 ( .A(n17873), .B(n17872), .Z(n300) );
  NAND U556 ( .A(n299), .B(n300), .Z(n18149) );
  NAND U557 ( .A(n27892), .B(n27891), .Z(n301) );
  NAND U558 ( .A(n27890), .B(n27889), .Z(n302) );
  AND U559 ( .A(n301), .B(n302), .Z(n27921) );
  NAND U560 ( .A(n28212), .B(n28211), .Z(n303) );
  NAND U561 ( .A(n28209), .B(n28210), .Z(n304) );
  NAND U562 ( .A(n303), .B(n304), .Z(n28495) );
  NAND U563 ( .A(n28453), .B(n28452), .Z(n305) );
  NANDN U564 ( .A(n28451), .B(n28450), .Z(n306) );
  AND U565 ( .A(n305), .B(n306), .Z(n28488) );
  NAND U566 ( .A(n29645), .B(n29644), .Z(n307) );
  NAND U567 ( .A(n29642), .B(n29643), .Z(n308) );
  NAND U568 ( .A(n307), .B(n308), .Z(n30145) );
  NAND U569 ( .A(n30428), .B(n30427), .Z(n309) );
  NAND U570 ( .A(n30426), .B(n30425), .Z(n310) );
  AND U571 ( .A(n309), .B(n310), .Z(n30691) );
  XNOR U572 ( .A(n31403), .B(n31402), .Z(n31234) );
  NANDN U573 ( .A(n31767), .B(n31766), .Z(n311) );
  NANDN U574 ( .A(n31765), .B(n31764), .Z(n312) );
  AND U575 ( .A(n311), .B(n312), .Z(n32051) );
  NANDN U576 ( .A(n33404), .B(n33403), .Z(n313) );
  NANDN U577 ( .A(n33406), .B(n33405), .Z(n314) );
  NAND U578 ( .A(n313), .B(n314), .Z(n33563) );
  NAND U579 ( .A(n34234), .B(n34233), .Z(n315) );
  NANDN U580 ( .A(n34232), .B(n34231), .Z(n316) );
  NAND U581 ( .A(n315), .B(n316), .Z(n34531) );
  NANDN U582 ( .A(n34174), .B(n34173), .Z(n317) );
  NANDN U583 ( .A(n34176), .B(n34175), .Z(n318) );
  NAND U584 ( .A(n317), .B(n318), .Z(n34360) );
  NAND U585 ( .A(n34788), .B(n34789), .Z(n319) );
  NANDN U586 ( .A(n34787), .B(n34786), .Z(n320) );
  NAND U587 ( .A(n319), .B(n320), .Z(n35023) );
  NAND U588 ( .A(n35042), .B(n35041), .Z(n321) );
  NANDN U589 ( .A(n35040), .B(n35039), .Z(n322) );
  NAND U590 ( .A(n321), .B(n322), .Z(n35137) );
  NAND U591 ( .A(n37010), .B(n37009), .Z(n323) );
  NANDN U592 ( .A(n37008), .B(n37007), .Z(n324) );
  AND U593 ( .A(n323), .B(n324), .Z(n37099) );
  XNOR U594 ( .A(n37186), .B(n37187), .Z(n37189) );
  NAND U595 ( .A(n37283), .B(n37284), .Z(n325) );
  NANDN U596 ( .A(n37282), .B(n37281), .Z(n326) );
  NAND U597 ( .A(n325), .B(n326), .Z(n37393) );
  NAND U598 ( .A(n37343), .B(n37342), .Z(n327) );
  NAND U599 ( .A(n37341), .B(n37340), .Z(n328) );
  NAND U600 ( .A(n327), .B(n328), .Z(n37489) );
  NAND U601 ( .A(n4954), .B(n4953), .Z(n329) );
  NAND U602 ( .A(n4952), .B(n4951), .Z(n330) );
  NAND U603 ( .A(n329), .B(n330), .Z(n5139) );
  NAND U604 ( .A(n24173), .B(n24174), .Z(n331) );
  NANDN U605 ( .A(n24172), .B(n24171), .Z(n332) );
  NAND U606 ( .A(n331), .B(n332), .Z(n24181) );
  NANDN U607 ( .A(n27624), .B(n27623), .Z(n333) );
  NANDN U608 ( .A(n27626), .B(n27625), .Z(n334) );
  NAND U609 ( .A(n333), .B(n334), .Z(n27633) );
  NAND U610 ( .A(n27907), .B(n27908), .Z(n335) );
  NANDN U611 ( .A(n27906), .B(n27905), .Z(n336) );
  NAND U612 ( .A(n335), .B(n336), .Z(n27915) );
  XNOR U613 ( .A(n29054), .B(n29055), .Z(n29057) );
  NAND U614 ( .A(n31965), .B(n31964), .Z(n337) );
  NANDN U615 ( .A(n31963), .B(n31962), .Z(n338) );
  AND U616 ( .A(n337), .B(n338), .Z(n31978) );
  NAND U617 ( .A(n35105), .B(n35104), .Z(n339) );
  NAND U618 ( .A(n35103), .B(n35102), .Z(n340) );
  AND U619 ( .A(n339), .B(n340), .Z(n35262) );
  NAND U620 ( .A(n35926), .B(n35927), .Z(n341) );
  NANDN U621 ( .A(n35925), .B(n35924), .Z(n342) );
  NAND U622 ( .A(n341), .B(n342), .Z(n36196) );
  NAND U623 ( .A(n38072), .B(n38071), .Z(n343) );
  NANDN U624 ( .A(n38070), .B(n38069), .Z(n344) );
  AND U625 ( .A(n343), .B(n344), .Z(n38157) );
  OR U626 ( .A(n38117), .B(n38118), .Z(n345) );
  NANDN U627 ( .A(n38120), .B(n38119), .Z(n346) );
  NAND U628 ( .A(n345), .B(n346), .Z(n38184) );
  ANDN U629 ( .B(n1022), .A(n1021), .Z(n1042) );
  OR U630 ( .A(n2107), .B(n2108), .Z(n347) );
  NAND U631 ( .A(n2106), .B(n2105), .Z(n348) );
  NAND U632 ( .A(n347), .B(n348), .Z(n2194) );
  NAND U633 ( .A(n12716), .B(n12717), .Z(n349) );
  NANDN U634 ( .A(n12715), .B(n12714), .Z(n350) );
  NAND U635 ( .A(n349), .B(n350), .Z(n12997) );
  NAND U636 ( .A(n13571), .B(n13572), .Z(n351) );
  NANDN U637 ( .A(n13570), .B(n13569), .Z(n352) );
  NAND U638 ( .A(n351), .B(n352), .Z(n13855) );
  NAND U639 ( .A(n14423), .B(n14424), .Z(n353) );
  NANDN U640 ( .A(n14422), .B(n14421), .Z(n354) );
  NAND U641 ( .A(n353), .B(n354), .Z(n14706) );
  NAND U642 ( .A(n21605), .B(n21606), .Z(n355) );
  NANDN U643 ( .A(n21604), .B(n21603), .Z(n356) );
  NAND U644 ( .A(n355), .B(n356), .Z(n21887) );
  NAND U645 ( .A(n23611), .B(n23612), .Z(n357) );
  NANDN U646 ( .A(n23610), .B(n23609), .Z(n358) );
  NAND U647 ( .A(n357), .B(n358), .Z(n23900) );
  NAND U648 ( .A(n35901), .B(n35900), .Z(n359) );
  NANDN U649 ( .A(n35899), .B(n35898), .Z(n360) );
  AND U650 ( .A(n359), .B(n360), .Z(n36050) );
  NAND U651 ( .A(n36597), .B(n36598), .Z(n361) );
  NANDN U652 ( .A(n36596), .B(n36595), .Z(n362) );
  NAND U653 ( .A(n361), .B(n362), .Z(n36602) );
  NANDN U654 ( .A(n37195), .B(n37194), .Z(n363) );
  NANDN U655 ( .A(n37193), .B(n37192), .Z(n364) );
  AND U656 ( .A(n363), .B(n364), .Z(n37199) );
  NANDN U657 ( .A(n37671), .B(n37670), .Z(n365) );
  NANDN U658 ( .A(n37669), .B(n37668), .Z(n366) );
  AND U659 ( .A(n365), .B(n366), .Z(n37763) );
  NAND U660 ( .A(n1916), .B(n1917), .Z(n367) );
  NANDN U661 ( .A(n1915), .B(n1914), .Z(n368) );
  NAND U662 ( .A(n367), .B(n368), .Z(n1999) );
  NAND U663 ( .A(n4602), .B(n4603), .Z(n369) );
  NANDN U664 ( .A(n4601), .B(n4600), .Z(n370) );
  NAND U665 ( .A(n369), .B(n370), .Z(n4775) );
  NAND U666 ( .A(n5344), .B(n5345), .Z(n371) );
  NANDN U667 ( .A(n5343), .B(n5342), .Z(n372) );
  NAND U668 ( .A(n371), .B(n372), .Z(n5535) );
  XOR U669 ( .A(n29895), .B(n29894), .Z(n373) );
  NANDN U670 ( .A(n29893), .B(n373), .Z(n374) );
  NAND U671 ( .A(n29895), .B(n29894), .Z(n375) );
  AND U672 ( .A(n374), .B(n375), .Z(n30172) );
  NAND U673 ( .A(n31227), .B(n31225), .Z(n376) );
  NANDN U674 ( .A(n31227), .B(n31224), .Z(n377) );
  NANDN U675 ( .A(n31226), .B(n377), .Z(n378) );
  NAND U676 ( .A(n376), .B(n378), .Z(n31487) );
  XOR U677 ( .A(n32449), .B(n32448), .Z(n379) );
  NANDN U678 ( .A(n32447), .B(n379), .Z(n380) );
  NAND U679 ( .A(n32449), .B(n32448), .Z(n381) );
  AND U680 ( .A(n380), .B(n381), .Z(n32676) );
  NAND U681 ( .A(n33766), .B(n33767), .Z(n382) );
  NANDN U682 ( .A(n33765), .B(n33764), .Z(n383) );
  NAND U683 ( .A(n382), .B(n383), .Z(n33960) );
  NAND U684 ( .A(n36346), .B(n36345), .Z(n384) );
  XOR U685 ( .A(n36345), .B(n36346), .Z(n385) );
  NAND U686 ( .A(n385), .B(n36344), .Z(n386) );
  NAND U687 ( .A(n384), .B(n386), .Z(n36484) );
  XOR U688 ( .A(n37994), .B(n37993), .Z(n387) );
  NANDN U689 ( .A(n37992), .B(n387), .Z(n388) );
  NAND U690 ( .A(n37994), .B(n37993), .Z(n389) );
  AND U691 ( .A(n388), .B(n389), .Z(n38060) );
  NAND U692 ( .A(n38112), .B(n38111), .Z(n390) );
  NANDN U693 ( .A(n38110), .B(n38109), .Z(n391) );
  AND U694 ( .A(n390), .B(n391), .Z(n38115) );
  XOR U695 ( .A(n38271), .B(n38270), .Z(n392) );
  NANDN U696 ( .A(n38269), .B(n392), .Z(n393) );
  NAND U697 ( .A(n38271), .B(n38270), .Z(n394) );
  AND U698 ( .A(n393), .B(n394), .Z(n38308) );
  NAND U699 ( .A(n38416), .B(n38414), .Z(n395) );
  XOR U700 ( .A(n38414), .B(n38416), .Z(n396) );
  NANDN U701 ( .A(n38415), .B(n396), .Z(n397) );
  NAND U702 ( .A(n395), .B(n397), .Z(n38455) );
  XNOR U703 ( .A(n14320), .B(n14321), .Z(n14323) );
  XNOR U704 ( .A(n20023), .B(n20024), .Z(n20026) );
  XOR U705 ( .A(n20261), .B(n20262), .Z(n20263) );
  XOR U706 ( .A(n23180), .B(n23181), .Z(n23182) );
  XNOR U707 ( .A(n24367), .B(n24368), .Z(n24370) );
  XOR U708 ( .A(n24899), .B(n24900), .Z(n24901) );
  XOR U709 ( .A(n26606), .B(n26607), .Z(n26608) );
  NAND U710 ( .A(n9649), .B(n9650), .Z(n398) );
  NANDN U711 ( .A(n9648), .B(n9647), .Z(n399) );
  NAND U712 ( .A(n398), .B(n399), .Z(n10048) );
  NAND U713 ( .A(n11071), .B(n11072), .Z(n400) );
  NANDN U714 ( .A(n11074), .B(n11073), .Z(n401) );
  NAND U715 ( .A(n400), .B(n401), .Z(n11331) );
  NAND U716 ( .A(n11114), .B(n11113), .Z(n402) );
  NANDN U717 ( .A(n11112), .B(n11111), .Z(n403) );
  AND U718 ( .A(n402), .B(n403), .Z(n11481) );
  NAND U719 ( .A(n11479), .B(n11478), .Z(n404) );
  NANDN U720 ( .A(n11477), .B(n11476), .Z(n405) );
  AND U721 ( .A(n404), .B(n405), .Z(n11804) );
  NAND U722 ( .A(n11344), .B(n11345), .Z(n406) );
  NANDN U723 ( .A(n11343), .B(n11342), .Z(n407) );
  NAND U724 ( .A(n406), .B(n407), .Z(n11606) );
  NAND U725 ( .A(n12071), .B(n12072), .Z(n408) );
  NANDN U726 ( .A(n12070), .B(n12069), .Z(n409) );
  NAND U727 ( .A(n408), .B(n409), .Z(n12328) );
  NAND U728 ( .A(n12023), .B(n12024), .Z(n410) );
  NANDN U729 ( .A(n12026), .B(n12025), .Z(n411) );
  NAND U730 ( .A(n410), .B(n411), .Z(n12157) );
  NAND U731 ( .A(n12475), .B(n12476), .Z(n412) );
  NANDN U732 ( .A(n12474), .B(n12473), .Z(n413) );
  NAND U733 ( .A(n412), .B(n413), .Z(n12750) );
  NAND U734 ( .A(n12604), .B(n12603), .Z(n414) );
  NANDN U735 ( .A(n12602), .B(n12601), .Z(n415) );
  AND U736 ( .A(n414), .B(n415), .Z(n12908) );
  NAND U737 ( .A(n12756), .B(n12757), .Z(n416) );
  NANDN U738 ( .A(n12755), .B(n12754), .Z(n417) );
  NAND U739 ( .A(n416), .B(n417), .Z(n13019) );
  NAND U740 ( .A(n13654), .B(n13655), .Z(n418) );
  NANDN U741 ( .A(n13657), .B(n13656), .Z(n419) );
  NAND U742 ( .A(n418), .B(n419), .Z(n13875) );
  NAND U743 ( .A(n14041), .B(n14040), .Z(n420) );
  NANDN U744 ( .A(n14039), .B(n14038), .Z(n421) );
  AND U745 ( .A(n420), .B(n421), .Z(n14331) );
  NAND U746 ( .A(n14461), .B(n14462), .Z(n422) );
  NANDN U747 ( .A(n14460), .B(n14459), .Z(n423) );
  NAND U748 ( .A(n422), .B(n423), .Z(n14835) );
  NAND U749 ( .A(n14758), .B(n14757), .Z(n424) );
  NANDN U750 ( .A(n14756), .B(n14755), .Z(n425) );
  AND U751 ( .A(n424), .B(n425), .Z(n15227) );
  NAND U752 ( .A(n14840), .B(n14841), .Z(n426) );
  NANDN U753 ( .A(n14839), .B(n14838), .Z(n427) );
  NAND U754 ( .A(n426), .B(n427), .Z(n15022) );
  NAND U755 ( .A(n15045), .B(n15046), .Z(n428) );
  NANDN U756 ( .A(n15044), .B(n15043), .Z(n429) );
  NAND U757 ( .A(n428), .B(n429), .Z(n15408) );
  NAND U758 ( .A(n15622), .B(n15623), .Z(n430) );
  NANDN U759 ( .A(n15621), .B(n15620), .Z(n431) );
  NAND U760 ( .A(n430), .B(n431), .Z(n15893) );
  NAND U761 ( .A(n16188), .B(n16189), .Z(n432) );
  NANDN U762 ( .A(n16187), .B(n16186), .Z(n433) );
  NAND U763 ( .A(n432), .B(n433), .Z(n16432) );
  NAND U764 ( .A(n16766), .B(n16765), .Z(n434) );
  NANDN U765 ( .A(n16764), .B(n16763), .Z(n435) );
  AND U766 ( .A(n434), .B(n435), .Z(n17198) );
  NAND U767 ( .A(n16848), .B(n16849), .Z(n436) );
  NANDN U768 ( .A(n16847), .B(n16846), .Z(n437) );
  NAND U769 ( .A(n436), .B(n437), .Z(n17051) );
  NAND U770 ( .A(n17928), .B(n17929), .Z(n438) );
  NANDN U771 ( .A(n17927), .B(n17926), .Z(n439) );
  NAND U772 ( .A(n438), .B(n439), .Z(n18188) );
  NAND U773 ( .A(n18193), .B(n18194), .Z(n440) );
  NANDN U774 ( .A(n18192), .B(n18191), .Z(n441) );
  NAND U775 ( .A(n440), .B(n441), .Z(n18565) );
  NAND U776 ( .A(n18571), .B(n18572), .Z(n442) );
  NANDN U777 ( .A(n18570), .B(n18569), .Z(n443) );
  NAND U778 ( .A(n442), .B(n443), .Z(n18767) );
  NAND U779 ( .A(n18772), .B(n18773), .Z(n444) );
  NANDN U780 ( .A(n18771), .B(n18770), .Z(n445) );
  NAND U781 ( .A(n444), .B(n445), .Z(n19044) );
  NAND U782 ( .A(n19379), .B(n19380), .Z(n446) );
  NANDN U783 ( .A(n19382), .B(n19381), .Z(n447) );
  NAND U784 ( .A(n446), .B(n447), .Z(n19611) );
  NAND U785 ( .A(n19624), .B(n19625), .Z(n448) );
  NANDN U786 ( .A(n19623), .B(n19622), .Z(n449) );
  NAND U787 ( .A(n448), .B(n449), .Z(n19905) );
  NAND U788 ( .A(n20787), .B(n20788), .Z(n450) );
  NANDN U789 ( .A(n20786), .B(n20785), .Z(n451) );
  NAND U790 ( .A(n450), .B(n451), .Z(n21067) );
  NAND U791 ( .A(n20965), .B(n20964), .Z(n452) );
  NANDN U792 ( .A(n20963), .B(n20962), .Z(n453) );
  AND U793 ( .A(n452), .B(n453), .Z(n21172) );
  NAND U794 ( .A(n21262), .B(n21263), .Z(n454) );
  NANDN U795 ( .A(n21265), .B(n21264), .Z(n455) );
  NAND U796 ( .A(n454), .B(n455), .Z(n21342) );
  NAND U797 ( .A(n21216), .B(n21215), .Z(n456) );
  NANDN U798 ( .A(n21214), .B(n21213), .Z(n457) );
  AND U799 ( .A(n456), .B(n457), .Z(n21513) );
  NAND U800 ( .A(n21361), .B(n21362), .Z(n458) );
  NANDN U801 ( .A(n21360), .B(n21359), .Z(n459) );
  NAND U802 ( .A(n458), .B(n459), .Z(n21637) );
  NAND U803 ( .A(n21826), .B(n21825), .Z(n460) );
  NANDN U804 ( .A(n21824), .B(n21823), .Z(n461) );
  AND U805 ( .A(n460), .B(n461), .Z(n22106) );
  NAND U806 ( .A(n21783), .B(n21784), .Z(n462) );
  NANDN U807 ( .A(n21786), .B(n21785), .Z(n463) );
  NAND U808 ( .A(n462), .B(n463), .Z(n21895) );
  NAND U809 ( .A(n22214), .B(n22215), .Z(n464) );
  NANDN U810 ( .A(n22213), .B(n22212), .Z(n465) );
  NAND U811 ( .A(n464), .B(n465), .Z(n22504) );
  NAND U812 ( .A(n23528), .B(n23529), .Z(n466) );
  NANDN U813 ( .A(n23527), .B(n23526), .Z(n467) );
  NAND U814 ( .A(n466), .B(n467), .Z(n23695) );
  NAND U815 ( .A(n23367), .B(n23368), .Z(n468) );
  NANDN U816 ( .A(n23366), .B(n23365), .Z(n469) );
  NAND U817 ( .A(n468), .B(n469), .Z(n23765) );
  NAND U818 ( .A(n23731), .B(n23730), .Z(n470) );
  NANDN U819 ( .A(n23729), .B(n23728), .Z(n471) );
  AND U820 ( .A(n470), .B(n471), .Z(n24035) );
  NAND U821 ( .A(n23939), .B(n23940), .Z(n472) );
  NANDN U822 ( .A(n23938), .B(n23937), .Z(n473) );
  NAND U823 ( .A(n472), .B(n473), .Z(n24219) );
  NAND U824 ( .A(n24079), .B(n24078), .Z(n474) );
  NANDN U825 ( .A(n24077), .B(n24076), .Z(n475) );
  AND U826 ( .A(n474), .B(n475), .Z(n24416) );
  NAND U827 ( .A(n24639), .B(n24640), .Z(n476) );
  NANDN U828 ( .A(n24638), .B(n24637), .Z(n477) );
  NAND U829 ( .A(n476), .B(n477), .Z(n24926) );
  NAND U830 ( .A(n25401), .B(n25402), .Z(n478) );
  NANDN U831 ( .A(n25400), .B(n25399), .Z(n479) );
  NAND U832 ( .A(n478), .B(n479), .Z(n25775) );
  NAND U833 ( .A(n25765), .B(n25764), .Z(n480) );
  NANDN U834 ( .A(n25763), .B(n25762), .Z(n481) );
  AND U835 ( .A(n480), .B(n481), .Z(n26017) );
  NAND U836 ( .A(n25798), .B(n25799), .Z(n482) );
  NANDN U837 ( .A(n25797), .B(n25796), .Z(n483) );
  NAND U838 ( .A(n482), .B(n483), .Z(n26049) );
  NAND U839 ( .A(n26054), .B(n26055), .Z(n484) );
  NANDN U840 ( .A(n26053), .B(n26052), .Z(n485) );
  NAND U841 ( .A(n484), .B(n485), .Z(n26260) );
  NAND U842 ( .A(n26550), .B(n26549), .Z(n486) );
  NANDN U843 ( .A(n26548), .B(n26547), .Z(n487) );
  AND U844 ( .A(n486), .B(n487), .Z(n26864) );
  XNOR U845 ( .A(n6117), .B(n6118), .Z(n6120) );
  XOR U846 ( .A(n6129), .B(n6130), .Z(n6131) );
  XOR U847 ( .A(n6123), .B(n6124), .Z(n6125) );
  XNOR U848 ( .A(n6740), .B(n6741), .Z(n6792) );
  XNOR U849 ( .A(n6460), .B(n6461), .Z(n6463) );
  NAND U850 ( .A(n7704), .B(n7703), .Z(n488) );
  NANDN U851 ( .A(n7702), .B(n7701), .Z(n489) );
  AND U852 ( .A(n488), .B(n489), .Z(n7767) );
  XNOR U853 ( .A(n7848), .B(n7849), .Z(n7841) );
  NAND U854 ( .A(n9396), .B(n9397), .Z(n490) );
  NANDN U855 ( .A(n9395), .B(n9394), .Z(n491) );
  NAND U856 ( .A(n490), .B(n491), .Z(n9780) );
  NANDN U857 ( .A(n9417), .B(n9416), .Z(n492) );
  NANDN U858 ( .A(n9419), .B(n9418), .Z(n493) );
  NAND U859 ( .A(n492), .B(n493), .Z(n9773) );
  NANDN U860 ( .A(n9822), .B(n9821), .Z(n494) );
  NANDN U861 ( .A(n9824), .B(n9823), .Z(n495) );
  NAND U862 ( .A(n494), .B(n495), .Z(n10043) );
  NAND U863 ( .A(n10016), .B(n10017), .Z(n496) );
  NANDN U864 ( .A(n10015), .B(n10014), .Z(n497) );
  NAND U865 ( .A(n496), .B(n497), .Z(n10176) );
  NAND U866 ( .A(n10068), .B(n10069), .Z(n498) );
  NANDN U867 ( .A(n10067), .B(n10066), .Z(n499) );
  NAND U868 ( .A(n498), .B(n499), .Z(n10397) );
  NAND U869 ( .A(n10280), .B(n10281), .Z(n500) );
  NANDN U870 ( .A(n10279), .B(n10278), .Z(n501) );
  NAND U871 ( .A(n500), .B(n501), .Z(n10658) );
  NAND U872 ( .A(n10897), .B(n10896), .Z(n502) );
  NANDN U873 ( .A(n10895), .B(n10894), .Z(n503) );
  AND U874 ( .A(n502), .B(n503), .Z(n11007) );
  OR U875 ( .A(n12331), .B(n12332), .Z(n504) );
  NANDN U876 ( .A(n12334), .B(n12333), .Z(n505) );
  AND U877 ( .A(n504), .B(n505), .Z(n12683) );
  XOR U878 ( .A(n13531), .B(n13532), .Z(n13533) );
  OR U879 ( .A(n13376), .B(n13377), .Z(n506) );
  NANDN U880 ( .A(n13379), .B(n13378), .Z(n507) );
  AND U881 ( .A(n506), .B(n507), .Z(n13818) );
  XOR U882 ( .A(n14948), .B(n14949), .Z(n14950) );
  XNOR U883 ( .A(n15524), .B(n15525), .Z(n15527) );
  OR U884 ( .A(n15789), .B(n15790), .Z(n508) );
  NANDN U885 ( .A(n15792), .B(n15791), .Z(n509) );
  AND U886 ( .A(n508), .B(n509), .Z(n16100) );
  XNOR U887 ( .A(n16956), .B(n16957), .Z(n16959) );
  OR U888 ( .A(n17508), .B(n17509), .Z(n510) );
  NANDN U889 ( .A(n17511), .B(n17510), .Z(n511) );
  AND U890 ( .A(n510), .B(n511), .Z(n17578) );
  OR U891 ( .A(n18025), .B(n18026), .Z(n512) );
  NANDN U892 ( .A(n18028), .B(n18027), .Z(n513) );
  AND U893 ( .A(n512), .B(n513), .Z(n18404) );
  NAND U894 ( .A(n18658), .B(n18657), .Z(n514) );
  NANDN U895 ( .A(n18656), .B(n18655), .Z(n515) );
  AND U896 ( .A(n514), .B(n515), .Z(n18863) );
  OR U897 ( .A(n18514), .B(n18515), .Z(n516) );
  NANDN U898 ( .A(n18517), .B(n18516), .Z(n517) );
  AND U899 ( .A(n516), .B(n517), .Z(n18979) );
  OR U900 ( .A(n18893), .B(n18894), .Z(n518) );
  NANDN U901 ( .A(n18896), .B(n18895), .Z(n519) );
  AND U902 ( .A(n518), .B(n519), .Z(n19251) );
  XOR U903 ( .A(n19547), .B(n19548), .Z(n19549) );
  OR U904 ( .A(n19407), .B(n19408), .Z(n520) );
  NANDN U905 ( .A(n19410), .B(n19409), .Z(n521) );
  AND U906 ( .A(n520), .B(n521), .Z(n19824) );
  OR U907 ( .A(n19744), .B(n19745), .Z(n522) );
  NANDN U908 ( .A(n19747), .B(n19746), .Z(n523) );
  AND U909 ( .A(n522), .B(n523), .Z(n20113) );
  XOR U910 ( .A(n20404), .B(n20405), .Z(n20406) );
  XNOR U911 ( .A(n20708), .B(n20709), .Z(n20711) );
  XOR U912 ( .A(n20990), .B(n20991), .Z(n20992) );
  OR U913 ( .A(n21508), .B(n21509), .Z(n524) );
  NANDN U914 ( .A(n21511), .B(n21510), .Z(n525) );
  NAND U915 ( .A(n524), .B(n525), .Z(n21851) );
  OR U916 ( .A(n21764), .B(n21765), .Z(n526) );
  NANDN U917 ( .A(n21767), .B(n21766), .Z(n527) );
  AND U918 ( .A(n526), .B(n527), .Z(n22117) );
  OR U919 ( .A(n23667), .B(n23668), .Z(n528) );
  NANDN U920 ( .A(n23670), .B(n23669), .Z(n529) );
  AND U921 ( .A(n528), .B(n529), .Z(n24138) );
  XOR U922 ( .A(n24502), .B(n24503), .Z(n24504) );
  XNOR U923 ( .A(n24792), .B(n24793), .Z(n24795) );
  XOR U924 ( .A(n25320), .B(n25321), .Z(n25322) );
  XNOR U925 ( .A(n25363), .B(n25364), .Z(n25366) );
  XNOR U926 ( .A(n26162), .B(n26163), .Z(n26165) );
  OR U927 ( .A(n25970), .B(n25971), .Z(n530) );
  NANDN U928 ( .A(n25973), .B(n25972), .Z(n531) );
  AND U929 ( .A(n530), .B(n531), .Z(n26224) );
  XOR U930 ( .A(n26747), .B(n26748), .Z(n26749) );
  OR U931 ( .A(n26587), .B(n26588), .Z(n532) );
  NANDN U932 ( .A(n26590), .B(n26589), .Z(n533) );
  AND U933 ( .A(n532), .B(n533), .Z(n27027) );
  NAND U934 ( .A(n27159), .B(n27158), .Z(n534) );
  NANDN U935 ( .A(n27157), .B(n27156), .Z(n535) );
  AND U936 ( .A(n534), .B(n535), .Z(n27499) );
  XNOR U937 ( .A(n28144), .B(n28145), .Z(n28147) );
  XNOR U938 ( .A(n28271), .B(n28272), .Z(n28274) );
  XNOR U939 ( .A(n32559), .B(n32560), .Z(n32562) );
  XNOR U940 ( .A(n2162), .B(n2163), .Z(n2165) );
  XOR U941 ( .A(n3159), .B(n3160), .Z(n3161) );
  NAND U942 ( .A(n3264), .B(n3263), .Z(n536) );
  NANDN U943 ( .A(n3262), .B(n3261), .Z(n537) );
  AND U944 ( .A(n536), .B(n537), .Z(n3387) );
  NAND U945 ( .A(n4129), .B(n4130), .Z(n538) );
  NANDN U946 ( .A(n4128), .B(n4127), .Z(n539) );
  NAND U947 ( .A(n538), .B(n539), .Z(n4324) );
  XNOR U948 ( .A(n5380), .B(n5381), .Z(n5383) );
  NAND U949 ( .A(n5806), .B(n5807), .Z(n540) );
  NANDN U950 ( .A(n5805), .B(n5804), .Z(n541) );
  NAND U951 ( .A(n540), .B(n541), .Z(n6137) );
  NAND U952 ( .A(n5552), .B(n5553), .Z(n542) );
  NANDN U953 ( .A(n5551), .B(n5550), .Z(n543) );
  NAND U954 ( .A(n542), .B(n543), .Z(n5771) );
  NANDN U955 ( .A(n6256), .B(n6255), .Z(n544) );
  NANDN U956 ( .A(n6258), .B(n6257), .Z(n545) );
  NAND U957 ( .A(n544), .B(n545), .Z(n6542) );
  NAND U958 ( .A(n6327), .B(n6328), .Z(n546) );
  NANDN U959 ( .A(n6326), .B(n6325), .Z(n547) );
  NAND U960 ( .A(n546), .B(n547), .Z(n6536) );
  XNOR U961 ( .A(n6275), .B(n6274), .Z(n6276) );
  XOR U962 ( .A(n6353), .B(n6354), .Z(n6355) );
  NAND U963 ( .A(n6624), .B(n6625), .Z(n548) );
  NANDN U964 ( .A(n6627), .B(n6626), .Z(n549) );
  NAND U965 ( .A(n548), .B(n549), .Z(n7022) );
  NANDN U966 ( .A(n6416), .B(n6415), .Z(n550) );
  NANDN U967 ( .A(n6418), .B(n6417), .Z(n551) );
  NAND U968 ( .A(n550), .B(n551), .Z(n6668) );
  XNOR U969 ( .A(n7010), .B(n7009), .Z(n6839) );
  NAND U970 ( .A(n7243), .B(n7244), .Z(n552) );
  NANDN U971 ( .A(n7242), .B(n7241), .Z(n553) );
  NAND U972 ( .A(n552), .B(n553), .Z(n7357) );
  NAND U973 ( .A(n8127), .B(n8126), .Z(n554) );
  NANDN U974 ( .A(n8125), .B(n8124), .Z(n555) );
  AND U975 ( .A(n554), .B(n555), .Z(n8480) );
  XNOR U976 ( .A(n8215), .B(n8216), .Z(n8218) );
  NAND U977 ( .A(n7852), .B(n7853), .Z(n556) );
  NANDN U978 ( .A(n7855), .B(n7854), .Z(n557) );
  AND U979 ( .A(n556), .B(n557), .Z(n8209) );
  NAND U980 ( .A(n8400), .B(n8401), .Z(n558) );
  NANDN U981 ( .A(n8399), .B(n8398), .Z(n559) );
  NAND U982 ( .A(n558), .B(n559), .Z(n8600) );
  XOR U983 ( .A(n8581), .B(n8582), .Z(n8585) );
  NAND U984 ( .A(n8578), .B(n8577), .Z(n560) );
  NANDN U985 ( .A(n8576), .B(n8575), .Z(n561) );
  AND U986 ( .A(n560), .B(n561), .Z(n8908) );
  NAND U987 ( .A(n10701), .B(n10702), .Z(n562) );
  NANDN U988 ( .A(n10700), .B(n10699), .Z(n563) );
  NAND U989 ( .A(n562), .B(n563), .Z(n10967) );
  NAND U990 ( .A(n10988), .B(n10987), .Z(n564) );
  NANDN U991 ( .A(n10986), .B(n10985), .Z(n565) );
  AND U992 ( .A(n564), .B(n565), .Z(n11252) );
  NANDN U993 ( .A(n11013), .B(n11012), .Z(n566) );
  NANDN U994 ( .A(n11015), .B(n11014), .Z(n567) );
  NAND U995 ( .A(n566), .B(n567), .Z(n11302) );
  XOR U996 ( .A(n11535), .B(n11536), .Z(n11537) );
  NAND U997 ( .A(n11547), .B(n11548), .Z(n568) );
  NANDN U998 ( .A(n11550), .B(n11549), .Z(n569) );
  NAND U999 ( .A(n568), .B(n569), .Z(n11574) );
  NANDN U1000 ( .A(n12378), .B(n12377), .Z(n570) );
  NANDN U1001 ( .A(n12380), .B(n12379), .Z(n571) );
  NAND U1002 ( .A(n570), .B(n571), .Z(n12442) );
  XNOR U1003 ( .A(n13228), .B(n13227), .Z(n13229) );
  NANDN U1004 ( .A(n13234), .B(n13233), .Z(n572) );
  NANDN U1005 ( .A(n13236), .B(n13235), .Z(n573) );
  NAND U1006 ( .A(n572), .B(n573), .Z(n13293) );
  NAND U1007 ( .A(n13825), .B(n13826), .Z(n574) );
  NANDN U1008 ( .A(n13824), .B(n13823), .Z(n575) );
  NAND U1009 ( .A(n574), .B(n575), .Z(n14111) );
  NAND U1010 ( .A(n14097), .B(n14098), .Z(n576) );
  NANDN U1011 ( .A(n14100), .B(n14099), .Z(n577) );
  NAND U1012 ( .A(n576), .B(n577), .Z(n14140) );
  NANDN U1013 ( .A(n14679), .B(n14678), .Z(n578) );
  NANDN U1014 ( .A(n14677), .B(n14676), .Z(n579) );
  AND U1015 ( .A(n578), .B(n579), .Z(n14955) );
  NANDN U1016 ( .A(n15255), .B(n15254), .Z(n580) );
  NANDN U1017 ( .A(n15257), .B(n15256), .Z(n581) );
  NAND U1018 ( .A(n580), .B(n581), .Z(n15530) );
  NANDN U1019 ( .A(n15833), .B(n15832), .Z(n582) );
  NANDN U1020 ( .A(n15831), .B(n15830), .Z(n583) );
  AND U1021 ( .A(n582), .B(n583), .Z(n15867) );
  XOR U1022 ( .A(n16107), .B(n16106), .Z(n584) );
  NANDN U1023 ( .A(n16108), .B(n584), .Z(n585) );
  NAND U1024 ( .A(n16107), .B(n16106), .Z(n586) );
  AND U1025 ( .A(n585), .B(n586), .Z(n16395) );
  NANDN U1026 ( .A(n16673), .B(n16672), .Z(n587) );
  NANDN U1027 ( .A(n16675), .B(n16674), .Z(n588) );
  NAND U1028 ( .A(n587), .B(n588), .Z(n16971) );
  NANDN U1029 ( .A(n17312), .B(n17311), .Z(n589) );
  NANDN U1030 ( .A(n17310), .B(n17309), .Z(n590) );
  AND U1031 ( .A(n589), .B(n590), .Z(n17831) );
  NAND U1032 ( .A(n17587), .B(n17586), .Z(n591) );
  NANDN U1033 ( .A(n17585), .B(n17584), .Z(n592) );
  NAND U1034 ( .A(n591), .B(n592), .Z(n18128) );
  NAND U1035 ( .A(n17897), .B(n17896), .Z(n593) );
  NANDN U1036 ( .A(n17895), .B(n17894), .Z(n594) );
  AND U1037 ( .A(n593), .B(n594), .Z(n18156) );
  XNOR U1038 ( .A(n18678), .B(n18677), .Z(n18679) );
  NANDN U1039 ( .A(n18993), .B(n18992), .Z(n595) );
  NANDN U1040 ( .A(n18991), .B(n18990), .Z(n596) );
  AND U1041 ( .A(n595), .B(n596), .Z(n19012) );
  NAND U1042 ( .A(n19259), .B(n19260), .Z(n597) );
  NANDN U1043 ( .A(n19258), .B(n19257), .Z(n598) );
  NAND U1044 ( .A(n597), .B(n598), .Z(n19305) );
  NANDN U1045 ( .A(n19830), .B(n19829), .Z(n599) );
  NANDN U1046 ( .A(n19832), .B(n19831), .Z(n600) );
  NAND U1047 ( .A(n599), .B(n600), .Z(n19879) );
  NAND U1048 ( .A(n20121), .B(n20122), .Z(n601) );
  NANDN U1049 ( .A(n20120), .B(n20119), .Z(n602) );
  NAND U1050 ( .A(n601), .B(n602), .Z(n20423) );
  NAND U1051 ( .A(n20576), .B(n20577), .Z(n603) );
  NANDN U1052 ( .A(n20575), .B(n20574), .Z(n604) );
  NAND U1053 ( .A(n603), .B(n604), .Z(n21005) );
  NANDN U1054 ( .A(n22124), .B(n22123), .Z(n605) );
  NANDN U1055 ( .A(n22126), .B(n22125), .Z(n606) );
  NAND U1056 ( .A(n605), .B(n606), .Z(n22178) );
  NAND U1057 ( .A(n23287), .B(n23286), .Z(n607) );
  NANDN U1058 ( .A(n23285), .B(n23284), .Z(n608) );
  AND U1059 ( .A(n607), .B(n608), .Z(n23335) );
  NANDN U1060 ( .A(n24152), .B(n24151), .Z(n609) );
  NANDN U1061 ( .A(n24150), .B(n24149), .Z(n610) );
  AND U1062 ( .A(n609), .B(n610), .Z(n24192) );
  NAND U1063 ( .A(n25201), .B(n25202), .Z(n611) );
  NANDN U1064 ( .A(n25200), .B(n25199), .Z(n612) );
  NAND U1065 ( .A(n611), .B(n612), .Z(n25350) );
  NAND U1066 ( .A(n25361), .B(n25362), .Z(n613) );
  NANDN U1067 ( .A(n25360), .B(n25359), .Z(n614) );
  NAND U1068 ( .A(n613), .B(n614), .Z(n25654) );
  NANDN U1069 ( .A(n26238), .B(n26237), .Z(n615) );
  NANDN U1070 ( .A(n26236), .B(n26235), .Z(n616) );
  AND U1071 ( .A(n615), .B(n616), .Z(n26763) );
  NAND U1072 ( .A(n27032), .B(n27033), .Z(n617) );
  NANDN U1073 ( .A(n27035), .B(n27034), .Z(n618) );
  NAND U1074 ( .A(n617), .B(n618), .Z(n27311) );
  NAND U1075 ( .A(n27067), .B(n27068), .Z(n619) );
  NANDN U1076 ( .A(n27066), .B(n27065), .Z(n620) );
  NAND U1077 ( .A(n619), .B(n620), .Z(n27355) );
  NAND U1078 ( .A(n27496), .B(n27497), .Z(n621) );
  NANDN U1079 ( .A(n27495), .B(n27494), .Z(n622) );
  NAND U1080 ( .A(n621), .B(n622), .Z(n27865) );
  XOR U1081 ( .A(n28741), .B(n28742), .Z(n28743) );
  NAND U1082 ( .A(n28570), .B(n28571), .Z(n623) );
  NANDN U1083 ( .A(n28569), .B(n28568), .Z(n624) );
  NAND U1084 ( .A(n623), .B(n624), .Z(n28797) );
  XOR U1085 ( .A(n29858), .B(b[1]), .Z(n625) );
  NAND U1086 ( .A(n625), .B(n29108), .Z(n626) );
  NAND U1087 ( .A(n29858), .B(b[1]), .Z(n627) );
  AND U1088 ( .A(n626), .B(n627), .Z(n29472) );
  NAND U1089 ( .A(n29224), .B(n29225), .Z(n628) );
  NANDN U1090 ( .A(n29227), .B(n29226), .Z(n629) );
  NAND U1091 ( .A(n628), .B(n629), .Z(n29579) );
  XNOR U1092 ( .A(n29708), .B(n29709), .Z(n29711) );
  NAND U1093 ( .A(n29704), .B(n29705), .Z(n630) );
  NANDN U1094 ( .A(n29707), .B(n29706), .Z(n631) );
  AND U1095 ( .A(n630), .B(n631), .Z(n30107) );
  XNOR U1096 ( .A(n29994), .B(n29995), .Z(n29997) );
  OR U1097 ( .A(n30267), .B(n30268), .Z(n632) );
  NANDN U1098 ( .A(n30266), .B(n30265), .Z(n633) );
  NAND U1099 ( .A(n632), .B(n633), .Z(n30599) );
  NAND U1100 ( .A(n32287), .B(n32288), .Z(n634) );
  NANDN U1101 ( .A(n32286), .B(n32285), .Z(n635) );
  NAND U1102 ( .A(n634), .B(n635), .Z(n32505) );
  XNOR U1103 ( .A(n32698), .B(n32699), .Z(n32701) );
  XNOR U1104 ( .A(n32736), .B(n32737), .Z(n32711) );
  XNOR U1105 ( .A(n32740), .B(n32741), .Z(n32743) );
  XOR U1106 ( .A(n33152), .B(n33002), .Z(n33003) );
  XNOR U1107 ( .A(n33652), .B(n33651), .Z(n33645) );
  NAND U1108 ( .A(n33909), .B(n33910), .Z(n636) );
  NANDN U1109 ( .A(n33912), .B(n33911), .Z(n637) );
  NAND U1110 ( .A(n636), .B(n637), .Z(n34121) );
  XOR U1111 ( .A(n34865), .B(n34866), .Z(n34867) );
  OR U1112 ( .A(n35185), .B(n35186), .Z(n638) );
  NANDN U1113 ( .A(n35184), .B(n35183), .Z(n639) );
  AND U1114 ( .A(n638), .B(n639), .Z(n35329) );
  NAND U1115 ( .A(n2061), .B(n2062), .Z(n640) );
  NANDN U1116 ( .A(n2060), .B(n2059), .Z(n641) );
  NAND U1117 ( .A(n640), .B(n641), .Z(n2128) );
  NAND U1118 ( .A(n1962), .B(n1963), .Z(n642) );
  NANDN U1119 ( .A(n1961), .B(n1960), .Z(n643) );
  NAND U1120 ( .A(n642), .B(n643), .Z(n2039) );
  NAND U1121 ( .A(n2264), .B(n2265), .Z(n644) );
  NANDN U1122 ( .A(n2263), .B(n2262), .Z(n645) );
  NAND U1123 ( .A(n644), .B(n645), .Z(n2390) );
  NAND U1124 ( .A(n2442), .B(n2443), .Z(n646) );
  NANDN U1125 ( .A(n2445), .B(n2444), .Z(n647) );
  NAND U1126 ( .A(n646), .B(n647), .Z(n2630) );
  XOR U1127 ( .A(n2792), .B(n2793), .Z(n2794) );
  XOR U1128 ( .A(n3201), .B(n3202), .Z(n3203) );
  XOR U1129 ( .A(n4072), .B(n4073), .Z(n4074) );
  NAND U1130 ( .A(n3842), .B(n3843), .Z(n648) );
  NANDN U1131 ( .A(n3841), .B(n3840), .Z(n649) );
  NAND U1132 ( .A(n648), .B(n649), .Z(n4063) );
  NANDN U1133 ( .A(n4154), .B(n4153), .Z(n650) );
  NANDN U1134 ( .A(n4156), .B(n4155), .Z(n651) );
  NAND U1135 ( .A(n650), .B(n651), .Z(n4267) );
  NANDN U1136 ( .A(n4589), .B(n4588), .Z(n652) );
  NANDN U1137 ( .A(n4587), .B(n4586), .Z(n653) );
  AND U1138 ( .A(n652), .B(n653), .Z(n4623) );
  XNOR U1139 ( .A(n4616), .B(n4617), .Z(n4613) );
  NAND U1140 ( .A(n4322), .B(n4323), .Z(n654) );
  NANDN U1141 ( .A(n4321), .B(n4320), .Z(n655) );
  NAND U1142 ( .A(n654), .B(n655), .Z(n4445) );
  XNOR U1143 ( .A(n4977), .B(n4978), .Z(n5035) );
  XOR U1144 ( .A(n4906), .B(n4907), .Z(n4908) );
  NAND U1145 ( .A(n5272), .B(n5273), .Z(n656) );
  NANDN U1146 ( .A(n5271), .B(n5270), .Z(n657) );
  NAND U1147 ( .A(n656), .B(n657), .Z(n5367) );
  NAND U1148 ( .A(n5318), .B(n5319), .Z(n658) );
  NANDN U1149 ( .A(n5317), .B(n5316), .Z(n659) );
  NAND U1150 ( .A(n658), .B(n659), .Z(n5523) );
  NAND U1151 ( .A(n5046), .B(n5047), .Z(n660) );
  NANDN U1152 ( .A(n5045), .B(n5044), .Z(n661) );
  NAND U1153 ( .A(n660), .B(n661), .Z(n5257) );
  NAND U1154 ( .A(n5591), .B(n5592), .Z(n662) );
  NANDN U1155 ( .A(n5590), .B(n5589), .Z(n663) );
  NAND U1156 ( .A(n662), .B(n663), .Z(n5766) );
  NAND U1157 ( .A(n5372), .B(n5373), .Z(n664) );
  NANDN U1158 ( .A(n5371), .B(n5370), .Z(n665) );
  NAND U1159 ( .A(n664), .B(n665), .Z(n5547) );
  NAND U1160 ( .A(n6097), .B(n6098), .Z(n666) );
  NANDN U1161 ( .A(n6096), .B(n6095), .Z(n667) );
  NAND U1162 ( .A(n666), .B(n667), .Z(n6286) );
  NAND U1163 ( .A(n6525), .B(n6526), .Z(n668) );
  NANDN U1164 ( .A(n6528), .B(n6527), .Z(n669) );
  NAND U1165 ( .A(n668), .B(n669), .Z(n6797) );
  OR U1166 ( .A(n6949), .B(n6950), .Z(n670) );
  NANDN U1167 ( .A(n6952), .B(n6951), .Z(n671) );
  AND U1168 ( .A(n670), .B(n671), .Z(n7072) );
  NAND U1169 ( .A(n6704), .B(n6703), .Z(n672) );
  NANDN U1170 ( .A(n6702), .B(n6701), .Z(n673) );
  AND U1171 ( .A(n672), .B(n673), .Z(n7028) );
  NANDN U1172 ( .A(n7881), .B(n7880), .Z(n674) );
  NANDN U1173 ( .A(n7883), .B(n7882), .Z(n675) );
  NAND U1174 ( .A(n674), .B(n675), .Z(n8223) );
  XNOR U1175 ( .A(n7963), .B(n7964), .Z(n7966) );
  XOR U1176 ( .A(n12121), .B(n12122), .Z(n12123) );
  NANDN U1177 ( .A(n12446), .B(n12445), .Z(n676) );
  NANDN U1178 ( .A(n12448), .B(n12447), .Z(n677) );
  NAND U1179 ( .A(n676), .B(n677), .Z(n12980) );
  XOR U1180 ( .A(n12973), .B(n12974), .Z(n12975) );
  XOR U1181 ( .A(n13261), .B(n13262), .Z(n13263) );
  NAND U1182 ( .A(n13298), .B(n13299), .Z(n678) );
  NANDN U1183 ( .A(n13297), .B(n13296), .Z(n679) );
  NAND U1184 ( .A(n678), .B(n679), .Z(n13838) );
  XOR U1185 ( .A(n13831), .B(n13832), .Z(n13833) );
  NAND U1186 ( .A(n14109), .B(n14110), .Z(n680) );
  NANDN U1187 ( .A(n14108), .B(n14107), .Z(n681) );
  NAND U1188 ( .A(n680), .B(n681), .Z(n14399) );
  NAND U1189 ( .A(n14148), .B(n14149), .Z(n682) );
  NANDN U1190 ( .A(n14147), .B(n14146), .Z(n683) );
  NAND U1191 ( .A(n682), .B(n683), .Z(n14687) );
  XOR U1192 ( .A(n14680), .B(n14681), .Z(n14682) );
  NAND U1193 ( .A(n14663), .B(n14662), .Z(n684) );
  NAND U1194 ( .A(n14661), .B(n14660), .Z(n685) );
  NAND U1195 ( .A(n684), .B(n685), .Z(n14966) );
  XNOR U1196 ( .A(n15001), .B(n15002), .Z(n15004) );
  NAND U1197 ( .A(n15247), .B(n15246), .Z(n686) );
  NAND U1198 ( .A(n15245), .B(n15244), .Z(n687) );
  NAND U1199 ( .A(n686), .B(n687), .Z(n15542) );
  XNOR U1200 ( .A(n15577), .B(n15578), .Z(n15580) );
  NAND U1201 ( .A(n15837), .B(n15836), .Z(n688) );
  NANDN U1202 ( .A(n15835), .B(n15834), .Z(n689) );
  AND U1203 ( .A(n688), .B(n689), .Z(n16122) );
  NAND U1204 ( .A(n16659), .B(n16658), .Z(n690) );
  NAND U1205 ( .A(n16656), .B(n16657), .Z(n691) );
  NAND U1206 ( .A(n690), .B(n691), .Z(n16975) );
  XNOR U1207 ( .A(n17013), .B(n17014), .Z(n17016) );
  XNOR U1208 ( .A(n17549), .B(n17550), .Z(n17552) );
  NAND U1209 ( .A(n17829), .B(n17830), .Z(n692) );
  NANDN U1210 ( .A(n17828), .B(n17827), .Z(n693) );
  NAND U1211 ( .A(n692), .B(n693), .Z(n17873) );
  NAND U1212 ( .A(n17901), .B(n17900), .Z(n694) );
  NAND U1213 ( .A(n17898), .B(n17899), .Z(n695) );
  NAND U1214 ( .A(n694), .B(n695), .Z(n18416) );
  XOR U1215 ( .A(n18695), .B(n18696), .Z(n18697) );
  XNOR U1216 ( .A(n19273), .B(n19274), .Z(n19280) );
  NAND U1217 ( .A(n19556), .B(n19555), .Z(n696) );
  NAND U1218 ( .A(n19554), .B(n19553), .Z(n697) );
  AND U1219 ( .A(n696), .B(n697), .Z(n19846) );
  XOR U1220 ( .A(n21580), .B(n21581), .Z(n21582) );
  XOR U1221 ( .A(n21861), .B(n21862), .Z(n21863) );
  NANDN U1222 ( .A(n21614), .B(n21613), .Z(n698) );
  NANDN U1223 ( .A(n21616), .B(n21615), .Z(n699) );
  NAND U1224 ( .A(n698), .B(n699), .Z(n22156) );
  XOR U1225 ( .A(n22149), .B(n22150), .Z(n22151) );
  NAND U1226 ( .A(n22186), .B(n22187), .Z(n700) );
  NANDN U1227 ( .A(n22185), .B(n22184), .Z(n701) );
  NAND U1228 ( .A(n700), .B(n701), .Z(n22731) );
  XOR U1229 ( .A(n22724), .B(n22725), .Z(n22726) );
  NAND U1230 ( .A(n23001), .B(n23000), .Z(n702) );
  NANDN U1231 ( .A(n22999), .B(n22998), .Z(n703) );
  AND U1232 ( .A(n702), .B(n703), .Z(n23300) );
  NAND U1233 ( .A(n23271), .B(n23270), .Z(n704) );
  NAND U1234 ( .A(n23268), .B(n23269), .Z(n705) );
  NAND U1235 ( .A(n704), .B(n705), .Z(n23589) );
  XOR U1236 ( .A(n23874), .B(n23875), .Z(n23876) );
  XOR U1237 ( .A(n24741), .B(n24742), .Z(n24743) );
  NAND U1238 ( .A(n24801), .B(n24800), .Z(n706) );
  NANDN U1239 ( .A(n24799), .B(n24798), .Z(n707) );
  AND U1240 ( .A(n706), .B(n707), .Z(n25069) );
  NAND U1241 ( .A(n25328), .B(n25329), .Z(n708) );
  NANDN U1242 ( .A(n25327), .B(n25326), .Z(n709) );
  NAND U1243 ( .A(n708), .B(n709), .Z(n25612) );
  NAND U1244 ( .A(n25889), .B(n25888), .Z(n710) );
  NAND U1245 ( .A(n25887), .B(n25886), .Z(n711) );
  NAND U1246 ( .A(n710), .B(n711), .Z(n26180) );
  NAND U1247 ( .A(n26210), .B(n26209), .Z(n712) );
  NAND U1248 ( .A(n26208), .B(n26207), .Z(n713) );
  NAND U1249 ( .A(n712), .B(n713), .Z(n26499) );
  NAND U1250 ( .A(n26761), .B(n26762), .Z(n714) );
  NANDN U1251 ( .A(n26760), .B(n26759), .Z(n715) );
  NAND U1252 ( .A(n714), .B(n715), .Z(n27049) );
  XOR U1253 ( .A(n27042), .B(n27043), .Z(n27044) );
  XOR U1254 ( .A(n27611), .B(n27612), .Z(n27613) );
  NAND U1255 ( .A(n27597), .B(n27598), .Z(n716) );
  NANDN U1256 ( .A(n27596), .B(n27595), .Z(n717) );
  NAND U1257 ( .A(n716), .B(n717), .Z(n27886) );
  NAND U1258 ( .A(n27954), .B(n27955), .Z(n718) );
  NANDN U1259 ( .A(n27953), .B(n27952), .Z(n719) );
  NAND U1260 ( .A(n718), .B(n719), .Z(n28463) );
  NAND U1261 ( .A(n27945), .B(n27944), .Z(n720) );
  NANDN U1262 ( .A(n27943), .B(n27942), .Z(n721) );
  AND U1263 ( .A(n720), .B(n721), .Z(n28457) );
  NAND U1264 ( .A(n28127), .B(n28128), .Z(n722) );
  NANDN U1265 ( .A(n28126), .B(n28125), .Z(n723) );
  NAND U1266 ( .A(n722), .B(n723), .Z(n28451) );
  NAND U1267 ( .A(n28893), .B(n28894), .Z(n724) );
  NANDN U1268 ( .A(n28892), .B(n28891), .Z(n725) );
  NAND U1269 ( .A(n724), .B(n725), .Z(n29142) );
  XOR U1270 ( .A(n29018), .B(n29019), .Z(n29020) );
  NAND U1271 ( .A(n28611), .B(n28610), .Z(n726) );
  NAND U1272 ( .A(n28609), .B(n28608), .Z(n727) );
  NAND U1273 ( .A(n726), .B(n727), .Z(n28784) );
  NAND U1274 ( .A(n30473), .B(n30474), .Z(n728) );
  NANDN U1275 ( .A(n30472), .B(n30471), .Z(n729) );
  NAND U1276 ( .A(n728), .B(n729), .Z(n30740) );
  NAND U1277 ( .A(n30477), .B(n30478), .Z(n730) );
  NANDN U1278 ( .A(n30476), .B(n30475), .Z(n731) );
  NAND U1279 ( .A(n730), .B(n731), .Z(n30794) );
  NAND U1280 ( .A(n30747), .B(n30748), .Z(n732) );
  NANDN U1281 ( .A(n30746), .B(n30745), .Z(n733) );
  NAND U1282 ( .A(n732), .B(n733), .Z(n31071) );
  XNOR U1283 ( .A(n31056), .B(n31057), .Z(n31059) );
  XNOR U1284 ( .A(n31406), .B(n31407), .Z(n31409) );
  XOR U1285 ( .A(n31816), .B(n31817), .Z(n31818) );
  NAND U1286 ( .A(n31586), .B(n31585), .Z(n734) );
  NANDN U1287 ( .A(n31584), .B(n31583), .Z(n735) );
  AND U1288 ( .A(n734), .B(n735), .Z(n31765) );
  NAND U1289 ( .A(n32512), .B(n32513), .Z(n736) );
  NANDN U1290 ( .A(n32511), .B(n32510), .Z(n737) );
  NAND U1291 ( .A(n736), .B(n737), .Z(n32681) );
  XNOR U1292 ( .A(n32876), .B(n32877), .Z(n32879) );
  NAND U1293 ( .A(n32825), .B(n32826), .Z(n738) );
  NANDN U1294 ( .A(n32828), .B(n32827), .Z(n739) );
  NAND U1295 ( .A(n738), .B(n739), .Z(n32925) );
  XNOR U1296 ( .A(n33307), .B(n33308), .Z(n33310) );
  XOR U1297 ( .A(n33319), .B(n33320), .Z(n33321) );
  XNOR U1298 ( .A(n33933), .B(n33934), .Z(n33831) );
  XOR U1299 ( .A(n34197), .B(n34198), .Z(n34317) );
  XNOR U1300 ( .A(n34373), .B(n34374), .Z(n34392) );
  NAND U1301 ( .A(n36242), .B(n36243), .Z(n740) );
  NANDN U1302 ( .A(n36241), .B(n36240), .Z(n741) );
  NAND U1303 ( .A(n740), .B(n741), .Z(n36360) );
  NANDN U1304 ( .A(n36532), .B(n36531), .Z(n742) );
  NANDN U1305 ( .A(n36534), .B(n36533), .Z(n743) );
  NAND U1306 ( .A(n742), .B(n743), .Z(n36715) );
  NANDN U1307 ( .A(n36588), .B(n36587), .Z(n744) );
  NANDN U1308 ( .A(n36590), .B(n36589), .Z(n745) );
  NAND U1309 ( .A(n744), .B(n745), .Z(n36703) );
  NAND U1310 ( .A(n1625), .B(n1626), .Z(n746) );
  NANDN U1311 ( .A(n1628), .B(n1627), .Z(n747) );
  NAND U1312 ( .A(n746), .B(n747), .Z(n1671) );
  NAND U1313 ( .A(n1537), .B(n1536), .Z(n748) );
  NANDN U1314 ( .A(n1535), .B(n1534), .Z(n749) );
  AND U1315 ( .A(n748), .B(n749), .Z(n1642) );
  NAND U1316 ( .A(n1804), .B(n1803), .Z(n750) );
  NANDN U1317 ( .A(n1802), .B(n1801), .Z(n751) );
  AND U1318 ( .A(n750), .B(n751), .Z(n1888) );
  XOR U1319 ( .A(n2430), .B(n2431), .Z(n2432) );
  NAND U1320 ( .A(n2239), .B(n2238), .Z(n752) );
  NANDN U1321 ( .A(n2237), .B(n2236), .Z(n753) );
  AND U1322 ( .A(n752), .B(n753), .Z(n2395) );
  NANDN U1323 ( .A(n2889), .B(n2888), .Z(n754) );
  NANDN U1324 ( .A(n2887), .B(n2886), .Z(n755) );
  AND U1325 ( .A(n754), .B(n755), .Z(n2920) );
  NAND U1326 ( .A(n3126), .B(n3127), .Z(n756) );
  NANDN U1327 ( .A(n3125), .B(n3124), .Z(n757) );
  NAND U1328 ( .A(n756), .B(n757), .Z(n3297) );
  NAND U1329 ( .A(n3576), .B(n3577), .Z(n758) );
  NANDN U1330 ( .A(n3575), .B(n3574), .Z(n759) );
  NAND U1331 ( .A(n758), .B(n759), .Z(n3751) );
  NANDN U1332 ( .A(n5927), .B(n5926), .Z(n760) );
  NANDN U1333 ( .A(n5925), .B(n5924), .Z(n761) );
  AND U1334 ( .A(n760), .B(n761), .Z(n5959) );
  XOR U1335 ( .A(n7500), .B(n7501), .Z(n7502) );
  NAND U1336 ( .A(n7733), .B(n7734), .Z(n762) );
  NANDN U1337 ( .A(n7736), .B(n7735), .Z(n763) );
  NAND U1338 ( .A(n762), .B(n763), .Z(n7981) );
  OR U1339 ( .A(n7725), .B(n7726), .Z(n764) );
  NAND U1340 ( .A(n7724), .B(n7723), .Z(n765) );
  NAND U1341 ( .A(n764), .B(n765), .Z(n7976) );
  NANDN U1342 ( .A(n8270), .B(n8269), .Z(n766) );
  NANDN U1343 ( .A(n8272), .B(n8271), .Z(n767) );
  NAND U1344 ( .A(n766), .B(n767), .Z(n8759) );
  NANDN U1345 ( .A(n12413), .B(n12412), .Z(n768) );
  NANDN U1346 ( .A(n12415), .B(n12414), .Z(n769) );
  NAND U1347 ( .A(n768), .B(n769), .Z(n12703) );
  NAND U1348 ( .A(n16691), .B(n16690), .Z(n770) );
  NANDN U1349 ( .A(n16689), .B(n16688), .Z(n771) );
  AND U1350 ( .A(n770), .B(n771), .Z(n16984) );
  NAND U1351 ( .A(n23017), .B(n23016), .Z(n772) );
  NANDN U1352 ( .A(n23015), .B(n23014), .Z(n773) );
  AND U1353 ( .A(n772), .B(n773), .Z(n23312) );
  XNOR U1354 ( .A(n27928), .B(n27929), .Z(n27923) );
  NAND U1355 ( .A(n28443), .B(n28442), .Z(n774) );
  NANDN U1356 ( .A(n28441), .B(n28440), .Z(n775) );
  NAND U1357 ( .A(n774), .B(n775), .Z(n28490) );
  XNOR U1358 ( .A(n28778), .B(n28779), .Z(n28780) );
  OR U1359 ( .A(n28792), .B(n28793), .Z(n776) );
  NAND U1360 ( .A(n28791), .B(n28790), .Z(n777) );
  NAND U1361 ( .A(n776), .B(n777), .Z(n29148) );
  NAND U1362 ( .A(n29594), .B(n29595), .Z(n778) );
  NANDN U1363 ( .A(n29593), .B(n29592), .Z(n779) );
  NAND U1364 ( .A(n778), .B(n779), .Z(n29625) );
  NAND U1365 ( .A(n29585), .B(n29584), .Z(n780) );
  NANDN U1366 ( .A(n29583), .B(n29582), .Z(n781) );
  AND U1367 ( .A(n780), .B(n781), .Z(n29637) );
  XNOR U1368 ( .A(n31400), .B(n31401), .Z(n31403) );
  NAND U1369 ( .A(n31511), .B(n31512), .Z(n782) );
  NANDN U1370 ( .A(n31510), .B(n31509), .Z(n783) );
  NAND U1371 ( .A(n782), .B(n783), .Z(n31746) );
  XOR U1372 ( .A(n32242), .B(n32243), .Z(n32244) );
  XOR U1373 ( .A(n33128), .B(n33129), .Z(n33130) );
  XNOR U1374 ( .A(n33140), .B(n33141), .Z(n33143) );
  NANDN U1375 ( .A(n33382), .B(n33381), .Z(n784) );
  NANDN U1376 ( .A(n33384), .B(n33383), .Z(n785) );
  NAND U1377 ( .A(n784), .B(n785), .Z(n33565) );
  NAND U1378 ( .A(n34327), .B(n34328), .Z(n786) );
  NANDN U1379 ( .A(n34330), .B(n34329), .Z(n787) );
  NAND U1380 ( .A(n786), .B(n787), .Z(n34534) );
  NANDN U1381 ( .A(n35036), .B(n35035), .Z(n788) );
  NANDN U1382 ( .A(n35038), .B(n35037), .Z(n789) );
  NAND U1383 ( .A(n788), .B(n789), .Z(n35140) );
  NAND U1384 ( .A(n35115), .B(n35114), .Z(n790) );
  NANDN U1385 ( .A(n35113), .B(n35112), .Z(n791) );
  NAND U1386 ( .A(n790), .B(n791), .Z(n35400) );
  XNOR U1387 ( .A(n35888), .B(n35889), .Z(n35758) );
  NANDN U1388 ( .A(n35464), .B(n35463), .Z(n792) );
  NANDN U1389 ( .A(n35466), .B(n35465), .Z(n793) );
  NAND U1390 ( .A(n792), .B(n793), .Z(n35723) );
  NAND U1391 ( .A(n35591), .B(n35590), .Z(n794) );
  NANDN U1392 ( .A(n35589), .B(n35588), .Z(n795) );
  AND U1393 ( .A(n794), .B(n795), .Z(n35719) );
  NAND U1394 ( .A(n36523), .B(n36524), .Z(n796) );
  NANDN U1395 ( .A(n36522), .B(n36521), .Z(n797) );
  NAND U1396 ( .A(n796), .B(n797), .Z(n36610) );
  XNOR U1397 ( .A(n37100), .B(n37101), .Z(n37093) );
  NAND U1398 ( .A(n37224), .B(n37225), .Z(n798) );
  NANDN U1399 ( .A(n37223), .B(n37222), .Z(n799) );
  NAND U1400 ( .A(n798), .B(n799), .Z(n37398) );
  NAND U1401 ( .A(n37577), .B(n37578), .Z(n800) );
  NANDN U1402 ( .A(n37576), .B(n37575), .Z(n801) );
  NAND U1403 ( .A(n800), .B(n801), .Z(n37663) );
  XOR U1404 ( .A(n38287), .B(n38288), .Z(n38289) );
  NAND U1405 ( .A(n1116), .B(n1117), .Z(n802) );
  NANDN U1406 ( .A(n1115), .B(n1114), .Z(n803) );
  NAND U1407 ( .A(n802), .B(n803), .Z(n1150) );
  NANDN U1408 ( .A(n1394), .B(n1393), .Z(n804) );
  NANDN U1409 ( .A(n1396), .B(n1395), .Z(n805) );
  NAND U1410 ( .A(n804), .B(n805), .Z(n1504) );
  NAND U1411 ( .A(n1650), .B(n1649), .Z(n806) );
  NANDN U1412 ( .A(n1648), .B(n1647), .Z(n807) );
  AND U1413 ( .A(n806), .B(n807), .Z(n1658) );
  NAND U1414 ( .A(n1897), .B(n1896), .Z(n808) );
  NANDN U1415 ( .A(n1895), .B(n1894), .Z(n809) );
  AND U1416 ( .A(n808), .B(n809), .Z(n1990) );
  NAND U1417 ( .A(n3167), .B(n3168), .Z(n810) );
  NANDN U1418 ( .A(n3166), .B(n3165), .Z(n811) );
  NAND U1419 ( .A(n810), .B(n811), .Z(n3304) );
  NAND U1420 ( .A(n3331), .B(n3332), .Z(n812) );
  NANDN U1421 ( .A(n3330), .B(n3329), .Z(n813) );
  NAND U1422 ( .A(n812), .B(n813), .Z(n3461) );
  NAND U1423 ( .A(n3776), .B(n3775), .Z(n814) );
  NAND U1424 ( .A(n3773), .B(n3774), .Z(n815) );
  NAND U1425 ( .A(n814), .B(n815), .Z(n3932) );
  NAND U1426 ( .A(n6361), .B(n6362), .Z(n816) );
  NANDN U1427 ( .A(n6360), .B(n6359), .Z(n817) );
  NAND U1428 ( .A(n816), .B(n817), .Z(n6580) );
  OR U1429 ( .A(n6823), .B(n6824), .Z(n818) );
  NAND U1430 ( .A(n6822), .B(n6821), .Z(n819) );
  NAND U1431 ( .A(n818), .B(n819), .Z(n7053) );
  NAND U1432 ( .A(n9603), .B(n9604), .Z(n820) );
  NANDN U1433 ( .A(n9602), .B(n9601), .Z(n821) );
  NAND U1434 ( .A(n820), .B(n821), .Z(n9855) );
  NAND U1435 ( .A(n11277), .B(n11278), .Z(n822) );
  NANDN U1436 ( .A(n11276), .B(n11275), .Z(n823) );
  NAND U1437 ( .A(n822), .B(n823), .Z(n11285) );
  NANDN U1438 ( .A(n19858), .B(n19857), .Z(n824) );
  NANDN U1439 ( .A(n19860), .B(n19859), .Z(n825) );
  NAND U1440 ( .A(n824), .B(n825), .Z(n19867) );
  NANDN U1441 ( .A(n21021), .B(n21020), .Z(n826) );
  NANDN U1442 ( .A(n21023), .B(n21022), .Z(n827) );
  NAND U1443 ( .A(n826), .B(n827), .Z(n21030) );
  NAND U1444 ( .A(n26195), .B(n26194), .Z(n828) );
  NANDN U1445 ( .A(n26193), .B(n26192), .Z(n829) );
  AND U1446 ( .A(n828), .B(n829), .Z(n26202) );
  NAND U1447 ( .A(n29598), .B(n29599), .Z(n830) );
  NANDN U1448 ( .A(n29597), .B(n29596), .Z(n831) );
  NAND U1449 ( .A(n830), .B(n831), .Z(n29620) );
  NAND U1450 ( .A(n29660), .B(n29661), .Z(n832) );
  NANDN U1451 ( .A(n29659), .B(n29658), .Z(n833) );
  NAND U1452 ( .A(n832), .B(n833), .Z(n30149) );
  NAND U1453 ( .A(n30190), .B(n30191), .Z(n834) );
  NANDN U1454 ( .A(n30189), .B(n30188), .Z(n835) );
  NAND U1455 ( .A(n834), .B(n835), .Z(n30696) );
  NAND U1456 ( .A(n33970), .B(n33971), .Z(n836) );
  NANDN U1457 ( .A(n33969), .B(n33968), .Z(n837) );
  NAND U1458 ( .A(n836), .B(n837), .Z(n34340) );
  NAND U1459 ( .A(n34145), .B(n34146), .Z(n838) );
  NANDN U1460 ( .A(n34144), .B(n34143), .Z(n839) );
  NAND U1461 ( .A(n838), .B(n839), .Z(n34164) );
  NAND U1462 ( .A(n34532), .B(n34533), .Z(n840) );
  NANDN U1463 ( .A(n34531), .B(n34530), .Z(n841) );
  NAND U1464 ( .A(n840), .B(n841), .Z(n34719) );
  NAND U1465 ( .A(n35021), .B(n35022), .Z(n842) );
  NANDN U1466 ( .A(n35020), .B(n35019), .Z(n843) );
  NAND U1467 ( .A(n842), .B(n843), .Z(n35091) );
  NANDN U1468 ( .A(n35733), .B(n35732), .Z(n844) );
  NANDN U1469 ( .A(n35735), .B(n35734), .Z(n845) );
  NAND U1470 ( .A(n844), .B(n845), .Z(n35900) );
  NANDN U1471 ( .A(n35929), .B(n35928), .Z(n846) );
  NANDN U1472 ( .A(n35931), .B(n35930), .Z(n847) );
  NAND U1473 ( .A(n846), .B(n847), .Z(n36061) );
  NAND U1474 ( .A(n37184), .B(n37185), .Z(n848) );
  NANDN U1475 ( .A(n37183), .B(n37182), .Z(n849) );
  NAND U1476 ( .A(n848), .B(n849), .Z(n37204) );
  NAND U1477 ( .A(n37490), .B(n37491), .Z(n850) );
  NANDN U1478 ( .A(n37489), .B(n37488), .Z(n851) );
  NAND U1479 ( .A(n850), .B(n851), .Z(n37507) );
  XNOR U1480 ( .A(n37852), .B(n37853), .Z(n37857) );
  NAND U1481 ( .A(n37913), .B(n37912), .Z(n852) );
  NANDN U1482 ( .A(n37911), .B(n37910), .Z(n853) );
  AND U1483 ( .A(n852), .B(n853), .Z(n37928) );
  NAND U1484 ( .A(n38121), .B(n38122), .Z(n854) );
  NANDN U1485 ( .A(n38124), .B(n38123), .Z(n855) );
  NAND U1486 ( .A(n854), .B(n855), .Z(n38179) );
  NANDN U1487 ( .A(n4424), .B(n4423), .Z(n856) );
  NANDN U1488 ( .A(n4426), .B(n4425), .Z(n857) );
  NAND U1489 ( .A(n856), .B(n857), .Z(n4601) );
  NAND U1490 ( .A(n9318), .B(n9317), .Z(n858) );
  NAND U1491 ( .A(n9315), .B(n9316), .Z(n859) );
  NAND U1492 ( .A(n858), .B(n859), .Z(n9583) );
  NAND U1493 ( .A(n10716), .B(n10717), .Z(n860) );
  NANDN U1494 ( .A(n10715), .B(n10714), .Z(n861) );
  NAND U1495 ( .A(n860), .B(n861), .Z(n11003) );
  NAND U1496 ( .A(n11862), .B(n11863), .Z(n862) );
  NANDN U1497 ( .A(n11861), .B(n11860), .Z(n863) );
  NAND U1498 ( .A(n862), .B(n863), .Z(n12147) );
  NAND U1499 ( .A(n12996), .B(n12997), .Z(n864) );
  NANDN U1500 ( .A(n12995), .B(n12994), .Z(n865) );
  NAND U1501 ( .A(n864), .B(n865), .Z(n13287) );
  NAND U1502 ( .A(n13854), .B(n13855), .Z(n866) );
  NANDN U1503 ( .A(n13853), .B(n13852), .Z(n867) );
  NAND U1504 ( .A(n866), .B(n867), .Z(n14137) );
  NAND U1505 ( .A(n14705), .B(n14706), .Z(n868) );
  NANDN U1506 ( .A(n14704), .B(n14703), .Z(n869) );
  NAND U1507 ( .A(n868), .B(n869), .Z(n14992) );
  NAND U1508 ( .A(n17289), .B(n17290), .Z(n870) );
  NANDN U1509 ( .A(n17288), .B(n17287), .Z(n871) );
  NAND U1510 ( .A(n870), .B(n871), .Z(n17575) );
  NAND U1511 ( .A(n18147), .B(n18148), .Z(n872) );
  NANDN U1512 ( .A(n18146), .B(n18145), .Z(n873) );
  NAND U1513 ( .A(n872), .B(n873), .Z(n18435) );
  NAND U1514 ( .A(n19296), .B(n19297), .Z(n874) );
  NANDN U1515 ( .A(n19295), .B(n19294), .Z(n875) );
  NAND U1516 ( .A(n874), .B(n875), .Z(n19583) );
  NAND U1517 ( .A(n21886), .B(n21887), .Z(n876) );
  NANDN U1518 ( .A(n21885), .B(n21884), .Z(n877) );
  NAND U1519 ( .A(n876), .B(n877), .Z(n22175) );
  NAND U1520 ( .A(n23899), .B(n23900), .Z(n878) );
  NANDN U1521 ( .A(n23898), .B(n23897), .Z(n879) );
  NAND U1522 ( .A(n878), .B(n879), .Z(n24183) );
  NAND U1523 ( .A(n24766), .B(n24767), .Z(n880) );
  NANDN U1524 ( .A(n24765), .B(n24764), .Z(n881) );
  NAND U1525 ( .A(n880), .B(n881), .Z(n25053) );
  NAND U1526 ( .A(n26776), .B(n26777), .Z(n882) );
  NANDN U1527 ( .A(n26775), .B(n26774), .Z(n883) );
  NAND U1528 ( .A(n882), .B(n883), .Z(n27062) );
  NAND U1529 ( .A(n27634), .B(n27635), .Z(n884) );
  NANDN U1530 ( .A(n27633), .B(n27632), .Z(n885) );
  NAND U1531 ( .A(n884), .B(n885), .Z(n27917) );
  NAND U1532 ( .A(n31968), .B(n31969), .Z(n886) );
  NANDN U1533 ( .A(n31967), .B(n31966), .Z(n887) );
  NAND U1534 ( .A(n886), .B(n887), .Z(n31980) );
  NAND U1535 ( .A(n32201), .B(n32200), .Z(n888) );
  NANDN U1536 ( .A(n32199), .B(n32198), .Z(n889) );
  AND U1537 ( .A(n888), .B(n889), .Z(n32441) );
  OR U1538 ( .A(n35262), .B(n35263), .Z(n890) );
  NANDN U1539 ( .A(n35265), .B(n35264), .Z(n891) );
  AND U1540 ( .A(n890), .B(n891), .Z(n35435) );
  NAND U1541 ( .A(n36068), .B(n36069), .Z(n892) );
  NANDN U1542 ( .A(n36067), .B(n36066), .Z(n893) );
  NAND U1543 ( .A(n892), .B(n893), .Z(n36336) );
  NAND U1544 ( .A(n1032), .B(n1031), .Z(n894) );
  XOR U1545 ( .A(n1031), .B(n1032), .Z(n895) );
  NANDN U1546 ( .A(n1033), .B(n895), .Z(n896) );
  NAND U1547 ( .A(n894), .B(n896), .Z(n1043) );
  NAND U1548 ( .A(n1232), .B(n1233), .Z(n897) );
  NANDN U1549 ( .A(n1231), .B(n1230), .Z(n898) );
  NAND U1550 ( .A(n897), .B(n898), .Z(n1272) );
  NAND U1551 ( .A(n2103), .B(n2104), .Z(n899) );
  NANDN U1552 ( .A(n2102), .B(n2101), .Z(n900) );
  NAND U1553 ( .A(n899), .B(n900), .Z(n2197) );
  NAND U1554 ( .A(n2536), .B(n2537), .Z(n901) );
  NANDN U1555 ( .A(n2535), .B(n2534), .Z(n902) );
  NAND U1556 ( .A(n901), .B(n902), .Z(n2650) );
  NAND U1557 ( .A(n4256), .B(n4257), .Z(n903) );
  NANDN U1558 ( .A(n4255), .B(n4254), .Z(n904) );
  NAND U1559 ( .A(n903), .B(n904), .Z(n4420) );
  NAND U1560 ( .A(n4967), .B(n4968), .Z(n905) );
  NANDN U1561 ( .A(n4966), .B(n4965), .Z(n906) );
  NAND U1562 ( .A(n905), .B(n906), .Z(n5147) );
  NAND U1563 ( .A(n5745), .B(n5746), .Z(n907) );
  NANDN U1564 ( .A(n5744), .B(n5743), .Z(n908) );
  NAND U1565 ( .A(n907), .B(n908), .Z(n5943) );
  NAND U1566 ( .A(n8005), .B(n8006), .Z(n909) );
  NANDN U1567 ( .A(n8004), .B(n8003), .Z(n910) );
  NAND U1568 ( .A(n909), .B(n910), .Z(n8248) );
  NAND U1569 ( .A(n28486), .B(n28485), .Z(n911) );
  NAND U1570 ( .A(n28483), .B(n28484), .Z(n912) );
  NAND U1571 ( .A(n911), .B(n912), .Z(n28775) );
  NAND U1572 ( .A(n29340), .B(n29339), .Z(n913) );
  XOR U1573 ( .A(n29339), .B(n29340), .Z(n914) );
  NAND U1574 ( .A(n914), .B(n29338), .Z(n915) );
  NAND U1575 ( .A(n913), .B(n915), .Z(n29615) );
  NAND U1576 ( .A(n30446), .B(n30444), .Z(n916) );
  XOR U1577 ( .A(n30444), .B(n30446), .Z(n917) );
  NANDN U1578 ( .A(n30445), .B(n917), .Z(n918) );
  NAND U1579 ( .A(n916), .B(n918), .Z(n30705) );
  NAND U1580 ( .A(n31733), .B(n31731), .Z(n919) );
  XOR U1581 ( .A(n31731), .B(n31733), .Z(n920) );
  NANDN U1582 ( .A(n31732), .B(n920), .Z(n921) );
  NAND U1583 ( .A(n919), .B(n921), .Z(n31973) );
  XOR U1584 ( .A(n32903), .B(n32902), .Z(n922) );
  NANDN U1585 ( .A(n32901), .B(n922), .Z(n923) );
  NAND U1586 ( .A(n32903), .B(n32902), .Z(n924) );
  AND U1587 ( .A(n923), .B(n924), .Z(n33118) );
  NAND U1588 ( .A(n33961), .B(n33959), .Z(n925) );
  XOR U1589 ( .A(n33959), .B(n33961), .Z(n926) );
  NANDN U1590 ( .A(n33960), .B(n926), .Z(n927) );
  NAND U1591 ( .A(n925), .B(n927), .Z(n34157) );
  XOR U1592 ( .A(n36059), .B(n36058), .Z(n928) );
  NANDN U1593 ( .A(n36057), .B(n928), .Z(n929) );
  NAND U1594 ( .A(n36059), .B(n36058), .Z(n930) );
  AND U1595 ( .A(n929), .B(n930), .Z(n36208) );
  NAND U1596 ( .A(n36484), .B(n36483), .Z(n931) );
  XOR U1597 ( .A(n36483), .B(n36484), .Z(n932) );
  NAND U1598 ( .A(n932), .B(n36482), .Z(n933) );
  NAND U1599 ( .A(n931), .B(n933), .Z(n36603) );
  NAND U1600 ( .A(n37091), .B(n37089), .Z(n934) );
  XOR U1601 ( .A(n37089), .B(n37091), .Z(n935) );
  NANDN U1602 ( .A(n37090), .B(n935), .Z(n936) );
  NAND U1603 ( .A(n934), .B(n936), .Z(n37200) );
  XOR U1604 ( .A(n37771), .B(n37770), .Z(n937) );
  NANDN U1605 ( .A(n37769), .B(n937), .Z(n938) );
  NAND U1606 ( .A(n37771), .B(n37770), .Z(n939) );
  AND U1607 ( .A(n938), .B(n939), .Z(n37846) );
  NAND U1608 ( .A(n38116), .B(n38115), .Z(n940) );
  XOR U1609 ( .A(n38115), .B(n38116), .Z(n941) );
  NAND U1610 ( .A(n941), .B(n38114), .Z(n942) );
  NAND U1611 ( .A(n940), .B(n942), .Z(n38172) );
  NANDN U1612 ( .A(n38215), .B(n38214), .Z(n943) );
  NANDN U1613 ( .A(n38213), .B(n38212), .Z(n944) );
  AND U1614 ( .A(n943), .B(n944), .Z(n38262) );
  NAND U1615 ( .A(n38308), .B(n38307), .Z(n945) );
  XOR U1616 ( .A(n38307), .B(n38308), .Z(n946) );
  NAND U1617 ( .A(n946), .B(n38306), .Z(n947) );
  NAND U1618 ( .A(n945), .B(n947), .Z(n38350) );
  NAND U1619 ( .A(n38389), .B(n38388), .Z(n948) );
  NANDN U1620 ( .A(n38387), .B(n38386), .Z(n949) );
  AND U1621 ( .A(n948), .B(n949), .Z(n38414) );
  OR U1622 ( .A(n985), .B(n38461), .Z(n950) );
  NANDN U1623 ( .A(n38462), .B(n950), .Z(n951) );
  ANDN U1624 ( .B(n951), .A(n38463), .Z(n952) );
  NANDN U1625 ( .A(n38465), .B(n38464), .Z(n953) );
  XNOR U1626 ( .A(n38465), .B(n38464), .Z(n954) );
  NAND U1627 ( .A(n954), .B(n38466), .Z(n955) );
  NAND U1628 ( .A(n953), .B(n955), .Z(n956) );
  XNOR U1629 ( .A(n952), .B(n956), .Z(n957) );
  NAND U1630 ( .A(n38468), .B(n38467), .Z(n958) );
  XOR U1631 ( .A(n38468), .B(n38467), .Z(n959) );
  NAND U1632 ( .A(n959), .B(n38469), .Z(n960) );
  AND U1633 ( .A(n958), .B(n960), .Z(n961) );
  XNOR U1634 ( .A(n957), .B(n961), .Z(n962) );
  NANDN U1635 ( .A(n38470), .B(n38471), .Z(n963) );
  XNOR U1636 ( .A(n962), .B(n963), .Z(c[255]) );
  XOR U1637 ( .A(b[55]), .B(b[56]), .Z(n964) );
  IV U1638 ( .A(n964), .Z(n965) );
  IV U1639 ( .A(b[0]), .Z(n966) );
  IV U1640 ( .A(b[3]), .Z(n967) );
  IV U1641 ( .A(b[5]), .Z(n968) );
  IV U1642 ( .A(b[9]), .Z(n969) );
  IV U1643 ( .A(b[11]), .Z(n970) );
  IV U1644 ( .A(b[13]), .Z(n971) );
  IV U1645 ( .A(b[15]), .Z(n972) );
  IV U1646 ( .A(b[31]), .Z(n973) );
  IV U1647 ( .A(b[33]), .Z(n974) );
  IV U1648 ( .A(b[37]), .Z(n975) );
  IV U1649 ( .A(b[39]), .Z(n976) );
  IV U1650 ( .A(b[43]), .Z(n977) );
  IV U1651 ( .A(b[47]), .Z(n978) );
  IV U1652 ( .A(b[49]), .Z(n979) );
  IV U1653 ( .A(b[51]), .Z(n980) );
  IV U1654 ( .A(b[53]), .Z(n981) );
  IV U1655 ( .A(b[55]), .Z(n982) );
  IV U1656 ( .A(b[57]), .Z(n983) );
  IV U1657 ( .A(b[61]), .Z(n984) );
  IV U1658 ( .A(b[63]), .Z(n985) );
  IV U1659 ( .A(a[0]), .Z(n986) );
  IV U1660 ( .A(a[126]), .Z(n987) );
  NANDN U1661 ( .A(n966), .B(a[0]), .Z(n989) );
  XNOR U1662 ( .A(n989), .B(sreg[64]), .Z(c[64]) );
  NANDN U1663 ( .A(n966), .B(a[1]), .Z(n994) );
  IV U1664 ( .A(b[1]), .Z(n29232) );
  NANDN U1665 ( .A(n29232), .B(a[0]), .Z(n988) );
  XOR U1666 ( .A(n994), .B(n988), .Z(n997) );
  XNOR U1667 ( .A(sreg[65]), .B(n997), .Z(n999) );
  NANDN U1668 ( .A(n989), .B(sreg[64]), .Z(n998) );
  XOR U1669 ( .A(n999), .B(n998), .Z(c[65]) );
  NANDN U1670 ( .A(n966), .B(a[2]), .Z(n990) );
  XOR U1671 ( .A(n29232), .B(n990), .Z(n992) );
  IV U1672 ( .A(a[1]), .Z(n10457) );
  NANDN U1673 ( .A(n10457), .B(n966), .Z(n991) );
  AND U1674 ( .A(n992), .B(n991), .Z(n1014) );
  NANDN U1675 ( .A(n986), .B(b[2]), .Z(n993) );
  XOR U1676 ( .A(n29232), .B(n993), .Z(n996) );
  OR U1677 ( .A(n994), .B(a[0]), .Z(n995) );
  AND U1678 ( .A(n996), .B(n995), .Z(n1013) );
  XNOR U1679 ( .A(n1014), .B(n1013), .Z(n1018) );
  NAND U1680 ( .A(n997), .B(sreg[65]), .Z(n1001) );
  OR U1681 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1682 ( .A(n1001), .B(n1000), .Z(n1016) );
  XNOR U1683 ( .A(n1016), .B(sreg[66]), .Z(n1017) );
  XOR U1684 ( .A(n1018), .B(n1017), .Z(c[66]) );
  XNOR U1685 ( .A(n967), .B(a[0]), .Z(n1004) );
  XNOR U1686 ( .A(n967), .B(b[1]), .Z(n1002) );
  XNOR U1687 ( .A(n967), .B(b[2]), .Z(n1027) );
  AND U1688 ( .A(n1002), .B(n1027), .Z(n1003) );
  NAND U1689 ( .A(n1004), .B(n1003), .Z(n1006) );
  XOR U1690 ( .A(b[3]), .B(n10457), .Z(n1028) );
  XNOR U1691 ( .A(n29232), .B(b[2]), .Z(n28939) );
  NANDN U1692 ( .A(n1028), .B(n28939), .Z(n1005) );
  AND U1693 ( .A(n1006), .B(n1005), .Z(n1021) );
  NANDN U1694 ( .A(n966), .B(a[3]), .Z(n1007) );
  XOR U1695 ( .A(n29232), .B(n1007), .Z(n1009) );
  IV U1696 ( .A(a[2]), .Z(n10363) );
  NANDN U1697 ( .A(n10363), .B(n966), .Z(n1008) );
  AND U1698 ( .A(n1009), .B(n1008), .Z(n1022) );
  XOR U1699 ( .A(n1021), .B(n1022), .Z(n1032) );
  ANDN U1700 ( .B(n986), .A(n967), .Z(n1010) );
  NAND U1701 ( .A(n1010), .B(n28939), .Z(n1012) );
  NOR U1702 ( .A(n967), .B(b[2]), .Z(n29370) );
  AND U1703 ( .A(b[3]), .B(n29232), .Z(n29371) );
  NAND U1704 ( .A(n29370), .B(n29371), .Z(n1011) );
  AND U1705 ( .A(n1012), .B(n1011), .Z(n1031) );
  AND U1706 ( .A(n1014), .B(n1013), .Z(n1033) );
  XNOR U1707 ( .A(n1031), .B(n1033), .Z(n1015) );
  XNOR U1708 ( .A(n1032), .B(n1015), .Z(n1035) );
  XNOR U1709 ( .A(sreg[67]), .B(n1035), .Z(n1037) );
  NAND U1710 ( .A(n1016), .B(sreg[66]), .Z(n1020) );
  OR U1711 ( .A(n1018), .B(n1017), .Z(n1019) );
  AND U1712 ( .A(n1020), .B(n1019), .Z(n1036) );
  XOR U1713 ( .A(n1037), .B(n1036), .Z(c[67]) );
  IV U1714 ( .A(n1042), .Z(n1040) );
  XNOR U1715 ( .A(b[3]), .B(b[4]), .Z(n29363) );
  NOR U1716 ( .A(n986), .B(n29363), .Z(n1064) );
  NANDN U1717 ( .A(n966), .B(a[4]), .Z(n1023) );
  XOR U1718 ( .A(n29232), .B(n1023), .Z(n1025) );
  IV U1719 ( .A(a[3]), .Z(n10524) );
  NANDN U1720 ( .A(n10524), .B(n966), .Z(n1024) );
  AND U1721 ( .A(n1025), .B(n1024), .Z(n1062) );
  XOR U1722 ( .A(b[3]), .B(n10363), .Z(n1058) );
  NANDN U1723 ( .A(n1058), .B(n28939), .Z(n1030) );
  XNOR U1724 ( .A(n29232), .B(b[3]), .Z(n1026) );
  AND U1725 ( .A(n1027), .B(n1026), .Z(n28938) );
  NANDN U1726 ( .A(n1028), .B(n28938), .Z(n1029) );
  AND U1727 ( .A(n1030), .B(n1029), .Z(n1061) );
  XNOR U1728 ( .A(n1062), .B(n1061), .Z(n1063) );
  XOR U1729 ( .A(n1064), .B(n1063), .Z(n1041) );
  XNOR U1730 ( .A(n1041), .B(n1043), .Z(n1034) );
  XNOR U1731 ( .A(n1040), .B(n1034), .Z(n1068) );
  NAND U1732 ( .A(sreg[67]), .B(n1035), .Z(n1039) );
  OR U1733 ( .A(n1037), .B(n1036), .Z(n1038) );
  NAND U1734 ( .A(n1039), .B(n1038), .Z(n1067) );
  XNOR U1735 ( .A(n1067), .B(sreg[68]), .Z(n1069) );
  XNOR U1736 ( .A(n1068), .B(n1069), .Z(c[68]) );
  NANDN U1737 ( .A(n1040), .B(n1041), .Z(n1046) );
  NOR U1738 ( .A(n1042), .B(n1041), .Z(n1044) );
  OR U1739 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1740 ( .A(n1046), .B(n1045), .Z(n1074) );
  NANDN U1741 ( .A(n966), .B(a[5]), .Z(n1047) );
  XOR U1742 ( .A(n29232), .B(n1047), .Z(n1049) );
  IV U1743 ( .A(a[4]), .Z(n10854) );
  NANDN U1744 ( .A(n10854), .B(n966), .Z(n1048) );
  AND U1745 ( .A(n1049), .B(n1048), .Z(n1079) );
  XNOR U1746 ( .A(n968), .B(a[0]), .Z(n1052) );
  XNOR U1747 ( .A(n968), .B(b[3]), .Z(n1087) );
  IV U1748 ( .A(b[4]), .Z(n30042) );
  XOR U1749 ( .A(n968), .B(n30042), .Z(n1050) );
  AND U1750 ( .A(n1087), .B(n1050), .Z(n1051) );
  NAND U1751 ( .A(n1052), .B(n1051), .Z(n1054) );
  XOR U1752 ( .A(n968), .B(a[1]), .Z(n1088) );
  OR U1753 ( .A(n1088), .B(n29363), .Z(n1053) );
  AND U1754 ( .A(n1054), .B(n1053), .Z(n1078) );
  XNOR U1755 ( .A(n1079), .B(n1078), .Z(n1094) );
  ANDN U1756 ( .B(n30042), .A(b[3]), .Z(n1055) );
  NANDN U1757 ( .A(n968), .B(n1055), .Z(n1057) );
  ANDN U1758 ( .B(b[5]), .A(n29363), .Z(n29866) );
  NANDN U1759 ( .A(a[0]), .B(n29866), .Z(n1056) );
  NAND U1760 ( .A(n1057), .B(n1056), .Z(n1092) );
  XNOR U1761 ( .A(n967), .B(a[3]), .Z(n1080) );
  NAND U1762 ( .A(n1080), .B(n28939), .Z(n1060) );
  NANDN U1763 ( .A(n1058), .B(n28938), .Z(n1059) );
  AND U1764 ( .A(n1060), .B(n1059), .Z(n1091) );
  XNOR U1765 ( .A(n1092), .B(n1091), .Z(n1093) );
  XNOR U1766 ( .A(n1094), .B(n1093), .Z(n1072) );
  NANDN U1767 ( .A(n1062), .B(n1061), .Z(n1066) );
  NANDN U1768 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1769 ( .A(n1066), .B(n1065), .Z(n1073) );
  XOR U1770 ( .A(n1072), .B(n1073), .Z(n1075) );
  XOR U1771 ( .A(n1074), .B(n1075), .Z(n1097) );
  XNOR U1772 ( .A(sreg[69]), .B(n1097), .Z(n1099) );
  NAND U1773 ( .A(n1067), .B(sreg[68]), .Z(n1071) );
  NANDN U1774 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1775 ( .A(n1071), .B(n1070), .Z(n1098) );
  XOR U1776 ( .A(n1099), .B(n1098), .Z(c[69]) );
  OR U1777 ( .A(n1073), .B(n1072), .Z(n1077) );
  NAND U1778 ( .A(n1075), .B(n1074), .Z(n1076) );
  NAND U1779 ( .A(n1077), .B(n1076), .Z(n1105) );
  ANDN U1780 ( .B(n1079), .A(n1078), .Z(n1111) );
  XNOR U1781 ( .A(n967), .B(a[4]), .Z(n1118) );
  NAND U1782 ( .A(n1118), .B(n28939), .Z(n1082) );
  NAND U1783 ( .A(n1080), .B(n28938), .Z(n1081) );
  NAND U1784 ( .A(n1082), .B(n1081), .Z(n1117) );
  XOR U1785 ( .A(b[6]), .B(b[5]), .Z(n29949) );
  NANDN U1786 ( .A(n986), .B(n29949), .Z(n1115) );
  NANDN U1787 ( .A(n966), .B(a[6]), .Z(n1083) );
  XOR U1788 ( .A(n29232), .B(n1083), .Z(n1085) );
  IV U1789 ( .A(a[5]), .Z(n11202) );
  NANDN U1790 ( .A(n11202), .B(n966), .Z(n1084) );
  AND U1791 ( .A(n1085), .B(n1084), .Z(n1114) );
  XNOR U1792 ( .A(n1115), .B(n1114), .Z(n1116) );
  XNOR U1793 ( .A(n1117), .B(n1116), .Z(n1108) );
  XNOR U1794 ( .A(n968), .B(b[4]), .Z(n1086) );
  AND U1795 ( .A(n1087), .B(n1086), .Z(n29864) );
  NANDN U1796 ( .A(n1088), .B(n29864), .Z(n1090) );
  XNOR U1797 ( .A(n968), .B(a[2]), .Z(n1121) );
  NANDN U1798 ( .A(n29363), .B(n1121), .Z(n1089) );
  NAND U1799 ( .A(n1090), .B(n1089), .Z(n1109) );
  XNOR U1800 ( .A(n1108), .B(n1109), .Z(n1110) );
  XOR U1801 ( .A(n1111), .B(n1110), .Z(n1102) );
  NANDN U1802 ( .A(n1092), .B(n1091), .Z(n1096) );
  NANDN U1803 ( .A(n1094), .B(n1093), .Z(n1095) );
  NAND U1804 ( .A(n1096), .B(n1095), .Z(n1103) );
  XNOR U1805 ( .A(n1102), .B(n1103), .Z(n1104) );
  XNOR U1806 ( .A(n1105), .B(n1104), .Z(n1135) );
  NAND U1807 ( .A(sreg[69]), .B(n1097), .Z(n1101) );
  OR U1808 ( .A(n1099), .B(n1098), .Z(n1100) );
  NAND U1809 ( .A(n1101), .B(n1100), .Z(n1133) );
  XNOR U1810 ( .A(n1133), .B(sreg[70]), .Z(n1134) );
  XOR U1811 ( .A(n1135), .B(n1134), .Z(c[70]) );
  NANDN U1812 ( .A(n1103), .B(n1102), .Z(n1107) );
  NAND U1813 ( .A(n1105), .B(n1104), .Z(n1106) );
  NAND U1814 ( .A(n1107), .B(n1106), .Z(n1146) );
  NANDN U1815 ( .A(n1109), .B(n1108), .Z(n1113) );
  NANDN U1816 ( .A(n1111), .B(n1110), .Z(n1112) );
  NAND U1817 ( .A(n1113), .B(n1112), .Z(n1144) );
  XNOR U1818 ( .A(n967), .B(a[5]), .Z(n1166) );
  NAND U1819 ( .A(n1166), .B(n28939), .Z(n1120) );
  NAND U1820 ( .A(n1118), .B(n28938), .Z(n1119) );
  AND U1821 ( .A(n1120), .B(n1119), .Z(n1149) );
  XNOR U1822 ( .A(n1150), .B(n1149), .Z(n1151) );
  XOR U1823 ( .A(n968), .B(n10524), .Z(n1174) );
  NANDN U1824 ( .A(n29363), .B(n1174), .Z(n1123) );
  NAND U1825 ( .A(n1121), .B(n29864), .Z(n1122) );
  NAND U1826 ( .A(n1123), .B(n1122), .Z(n1170) );
  IV U1827 ( .A(b[7]), .Z(n31123) );
  XNOR U1828 ( .A(n31123), .B(b[5]), .Z(n1161) );
  XNOR U1829 ( .A(n31123), .B(a[0]), .Z(n1124) );
  NAND U1830 ( .A(n1161), .B(n1124), .Z(n1125) );
  XNOR U1831 ( .A(n31123), .B(b[6]), .Z(n1162) );
  NANDN U1832 ( .A(n1125), .B(n1162), .Z(n1127) );
  XOR U1833 ( .A(n31123), .B(n10457), .Z(n1163) );
  NAND U1834 ( .A(n1163), .B(n29949), .Z(n1126) );
  NAND U1835 ( .A(n1127), .B(n1126), .Z(n1169) );
  XOR U1836 ( .A(n1170), .B(n1169), .Z(n1158) );
  ANDN U1837 ( .B(n968), .A(b[6]), .Z(n1128) );
  OR U1838 ( .A(n1128), .B(n986), .Z(n1129) );
  NANDN U1839 ( .A(n968), .B(b[6]), .Z(n30374) );
  ANDN U1840 ( .B(n30374), .A(n31123), .Z(n30751) );
  AND U1841 ( .A(n1129), .B(n30751), .Z(n1156) );
  NANDN U1842 ( .A(n966), .B(a[7]), .Z(n1130) );
  XOR U1843 ( .A(n29232), .B(n1130), .Z(n1132) );
  IV U1844 ( .A(a[6]), .Z(n11406) );
  NANDN U1845 ( .A(n11406), .B(n966), .Z(n1131) );
  AND U1846 ( .A(n1132), .B(n1131), .Z(n1155) );
  XOR U1847 ( .A(n1156), .B(n1155), .Z(n1157) );
  XOR U1848 ( .A(n1158), .B(n1157), .Z(n1152) );
  XNOR U1849 ( .A(n1151), .B(n1152), .Z(n1143) );
  XNOR U1850 ( .A(n1144), .B(n1143), .Z(n1145) );
  XNOR U1851 ( .A(n1146), .B(n1145), .Z(n1138) );
  XNOR U1852 ( .A(n1138), .B(sreg[71]), .Z(n1140) );
  NAND U1853 ( .A(n1133), .B(sreg[70]), .Z(n1137) );
  OR U1854 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1855 ( .A(n1137), .B(n1136), .Z(n1139) );
  XOR U1856 ( .A(n1140), .B(n1139), .Z(c[71]) );
  NAND U1857 ( .A(n1138), .B(sreg[71]), .Z(n1142) );
  OR U1858 ( .A(n1140), .B(n1139), .Z(n1141) );
  NAND U1859 ( .A(n1142), .B(n1141), .Z(n1220) );
  XNOR U1860 ( .A(n1220), .B(sreg[72]), .Z(n1222) );
  NAND U1861 ( .A(n1144), .B(n1143), .Z(n1148) );
  OR U1862 ( .A(n1146), .B(n1145), .Z(n1147) );
  NAND U1863 ( .A(n1148), .B(n1147), .Z(n1180) );
  NANDN U1864 ( .A(n1150), .B(n1149), .Z(n1154) );
  NANDN U1865 ( .A(n1152), .B(n1151), .Z(n1153) );
  NAND U1866 ( .A(n1154), .B(n1153), .Z(n1177) );
  OR U1867 ( .A(n1156), .B(n1155), .Z(n1160) );
  NANDN U1868 ( .A(n1158), .B(n1157), .Z(n1159) );
  NAND U1869 ( .A(n1160), .B(n1159), .Z(n1217) );
  XOR U1870 ( .A(n31123), .B(n10363), .Z(n1195) );
  NAND U1871 ( .A(n1195), .B(n29949), .Z(n1165) );
  AND U1872 ( .A(n1162), .B(n1161), .Z(n29948) );
  NAND U1873 ( .A(n29948), .B(n1163), .Z(n1164) );
  NAND U1874 ( .A(n1165), .B(n1164), .Z(n1183) );
  XOR U1875 ( .A(b[3]), .B(n11406), .Z(n1192) );
  NANDN U1876 ( .A(n1192), .B(n28939), .Z(n1168) );
  NAND U1877 ( .A(n1166), .B(n28938), .Z(n1167) );
  AND U1878 ( .A(n1168), .B(n1167), .Z(n1184) );
  XNOR U1879 ( .A(n1183), .B(n1184), .Z(n1185) );
  NAND U1880 ( .A(n1170), .B(n1169), .Z(n1186) );
  XOR U1881 ( .A(n1185), .B(n1186), .Z(n1214) );
  XNOR U1882 ( .A(n31123), .B(b[8]), .Z(n30509) );
  NAND U1883 ( .A(a[0]), .B(n30509), .Z(n1211) );
  NANDN U1884 ( .A(n966), .B(a[8]), .Z(n1171) );
  XOR U1885 ( .A(n29232), .B(n1171), .Z(n1173) );
  IV U1886 ( .A(a[7]), .Z(n11694) );
  NANDN U1887 ( .A(n11694), .B(n966), .Z(n1172) );
  AND U1888 ( .A(n1173), .B(n1172), .Z(n1209) );
  NAND U1889 ( .A(n29864), .B(n1174), .Z(n1176) );
  XNOR U1890 ( .A(n968), .B(a[4]), .Z(n1205) );
  NANDN U1891 ( .A(n29363), .B(n1205), .Z(n1175) );
  AND U1892 ( .A(n1176), .B(n1175), .Z(n1208) );
  XNOR U1893 ( .A(n1209), .B(n1208), .Z(n1210) );
  XNOR U1894 ( .A(n1211), .B(n1210), .Z(n1215) );
  XNOR U1895 ( .A(n1214), .B(n1215), .Z(n1216) );
  XNOR U1896 ( .A(n1217), .B(n1216), .Z(n1178) );
  XNOR U1897 ( .A(n1177), .B(n1178), .Z(n1179) );
  XOR U1898 ( .A(n1180), .B(n1179), .Z(n1221) );
  XOR U1899 ( .A(n1222), .B(n1221), .Z(c[72]) );
  NANDN U1900 ( .A(n1178), .B(n1177), .Z(n1182) );
  NAND U1901 ( .A(n1180), .B(n1179), .Z(n1181) );
  NAND U1902 ( .A(n1182), .B(n1181), .Z(n1233) );
  NANDN U1903 ( .A(n1184), .B(n1183), .Z(n1188) );
  NANDN U1904 ( .A(n1186), .B(n1185), .Z(n1187) );
  NAND U1905 ( .A(n1188), .B(n1187), .Z(n1237) );
  NANDN U1906 ( .A(n966), .B(a[9]), .Z(n1189) );
  XOR U1907 ( .A(n29232), .B(n1189), .Z(n1191) );
  IV U1908 ( .A(a[8]), .Z(n11986) );
  NANDN U1909 ( .A(n11986), .B(n966), .Z(n1190) );
  AND U1910 ( .A(n1191), .B(n1190), .Z(n1247) );
  XOR U1911 ( .A(b[3]), .B(n11694), .Z(n1260) );
  NANDN U1912 ( .A(n1260), .B(n28939), .Z(n1194) );
  NANDN U1913 ( .A(n1192), .B(n28938), .Z(n1193) );
  AND U1914 ( .A(n1194), .B(n1193), .Z(n1246) );
  XNOR U1915 ( .A(n1247), .B(n1246), .Z(n1248) );
  XNOR U1916 ( .A(n31123), .B(a[3]), .Z(n1266) );
  NAND U1917 ( .A(n1266), .B(n29949), .Z(n1197) );
  NAND U1918 ( .A(n29948), .B(n1195), .Z(n1196) );
  NAND U1919 ( .A(n1197), .B(n1196), .Z(n1252) );
  XOR U1920 ( .A(n969), .B(n10457), .Z(n1254) );
  NAND U1921 ( .A(n30509), .B(n1254), .Z(n1201) );
  XNOR U1922 ( .A(n969), .B(a[0]), .Z(n1312) );
  XNOR U1923 ( .A(n969), .B(b[7]), .Z(n1199) );
  XNOR U1924 ( .A(n969), .B(b[8]), .Z(n1198) );
  AND U1925 ( .A(n1199), .B(n1198), .Z(n30846) );
  NAND U1926 ( .A(n1312), .B(n30846), .Z(n1200) );
  AND U1927 ( .A(n1201), .B(n1200), .Z(n1253) );
  XNOR U1928 ( .A(n1252), .B(n1253), .Z(n1243) );
  NOR U1929 ( .A(b[7]), .B(b[8]), .Z(n1202) );
  NANDN U1930 ( .A(n969), .B(n1202), .Z(n1204) );
  ANDN U1931 ( .B(n30509), .A(n969), .Z(n30849) );
  NANDN U1932 ( .A(a[0]), .B(n30849), .Z(n1203) );
  NAND U1933 ( .A(n1204), .B(n1203), .Z(n1241) );
  XOR U1934 ( .A(n968), .B(n11202), .Z(n1257) );
  NANDN U1935 ( .A(n29363), .B(n1257), .Z(n1207) );
  NAND U1936 ( .A(n1205), .B(n29864), .Z(n1206) );
  NAND U1937 ( .A(n1207), .B(n1206), .Z(n1240) );
  XOR U1938 ( .A(n1241), .B(n1240), .Z(n1242) );
  XOR U1939 ( .A(n1243), .B(n1242), .Z(n1249) );
  XOR U1940 ( .A(n1248), .B(n1249), .Z(n1234) );
  NANDN U1941 ( .A(n1209), .B(n1208), .Z(n1213) );
  NAND U1942 ( .A(n1211), .B(n1210), .Z(n1212) );
  NAND U1943 ( .A(n1213), .B(n1212), .Z(n1235) );
  XNOR U1944 ( .A(n1234), .B(n1235), .Z(n1236) );
  XNOR U1945 ( .A(n1237), .B(n1236), .Z(n1230) );
  NANDN U1946 ( .A(n1215), .B(n1214), .Z(n1219) );
  NAND U1947 ( .A(n1217), .B(n1216), .Z(n1218) );
  AND U1948 ( .A(n1219), .B(n1218), .Z(n1231) );
  XNOR U1949 ( .A(n1230), .B(n1231), .Z(n1232) );
  XNOR U1950 ( .A(n1233), .B(n1232), .Z(n1225) );
  XNOR U1951 ( .A(n1225), .B(sreg[73]), .Z(n1227) );
  NAND U1952 ( .A(n1220), .B(sreg[72]), .Z(n1224) );
  OR U1953 ( .A(n1222), .B(n1221), .Z(n1223) );
  AND U1954 ( .A(n1224), .B(n1223), .Z(n1226) );
  XOR U1955 ( .A(n1227), .B(n1226), .Z(c[73]) );
  NAND U1956 ( .A(n1225), .B(sreg[73]), .Z(n1229) );
  OR U1957 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1958 ( .A(n1229), .B(n1228), .Z(n1321) );
  XNOR U1959 ( .A(n1321), .B(sreg[74]), .Z(n1323) );
  NANDN U1960 ( .A(n1235), .B(n1234), .Z(n1239) );
  NAND U1961 ( .A(n1237), .B(n1236), .Z(n1238) );
  NAND U1962 ( .A(n1239), .B(n1238), .Z(n1270) );
  OR U1963 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U1964 ( .A(n1243), .B(n1242), .Z(n1244) );
  NAND U1965 ( .A(n1245), .B(n1244), .Z(n1277) );
  NANDN U1966 ( .A(n1247), .B(n1246), .Z(n1251) );
  NANDN U1967 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U1968 ( .A(n1251), .B(n1250), .Z(n1276) );
  NANDN U1969 ( .A(n1253), .B(n1252), .Z(n1296) );
  NAND U1970 ( .A(n30846), .B(n1254), .Z(n1256) );
  XNOR U1971 ( .A(n969), .B(a[2]), .Z(n1307) );
  NAND U1972 ( .A(n30509), .B(n1307), .Z(n1255) );
  NAND U1973 ( .A(n1256), .B(n1255), .Z(n1294) );
  NAND U1974 ( .A(n29864), .B(n1257), .Z(n1259) );
  XOR U1975 ( .A(n968), .B(n11406), .Z(n1318) );
  NANDN U1976 ( .A(n29363), .B(n1318), .Z(n1258) );
  AND U1977 ( .A(n1259), .B(n1258), .Z(n1293) );
  XNOR U1978 ( .A(n1294), .B(n1293), .Z(n1295) );
  XNOR U1979 ( .A(n1296), .B(n1295), .Z(n1282) );
  XNOR U1980 ( .A(n967), .B(a[8]), .Z(n1304) );
  NAND U1981 ( .A(n1304), .B(n28939), .Z(n1262) );
  NANDN U1982 ( .A(n1260), .B(n28938), .Z(n1261) );
  AND U1983 ( .A(n1262), .B(n1261), .Z(n1281) );
  XNOR U1984 ( .A(n1282), .B(n1281), .Z(n1283) );
  XOR U1985 ( .A(n969), .B(b[10]), .Z(n31369) );
  NOR U1986 ( .A(n986), .B(n31369), .Z(n1290) );
  NANDN U1987 ( .A(n966), .B(a[10]), .Z(n1263) );
  XOR U1988 ( .A(n29232), .B(n1263), .Z(n1265) );
  IV U1989 ( .A(a[9]), .Z(n12258) );
  NANDN U1990 ( .A(n12258), .B(n966), .Z(n1264) );
  AND U1991 ( .A(n1265), .B(n1264), .Z(n1288) );
  XOR U1992 ( .A(b[7]), .B(n10854), .Z(n1299) );
  NANDN U1993 ( .A(n1299), .B(n29949), .Z(n1268) );
  NAND U1994 ( .A(n1266), .B(n29948), .Z(n1267) );
  AND U1995 ( .A(n1268), .B(n1267), .Z(n1287) );
  XNOR U1996 ( .A(n1288), .B(n1287), .Z(n1289) );
  XOR U1997 ( .A(n1290), .B(n1289), .Z(n1284) );
  XNOR U1998 ( .A(n1283), .B(n1284), .Z(n1275) );
  XNOR U1999 ( .A(n1276), .B(n1275), .Z(n1278) );
  XNOR U2000 ( .A(n1277), .B(n1278), .Z(n1269) );
  XNOR U2001 ( .A(n1270), .B(n1269), .Z(n1271) );
  XOR U2002 ( .A(n1272), .B(n1271), .Z(n1322) );
  XOR U2003 ( .A(n1323), .B(n1322), .Z(c[74]) );
  NANDN U2004 ( .A(n1270), .B(n1269), .Z(n1274) );
  NAND U2005 ( .A(n1272), .B(n1271), .Z(n1273) );
  NAND U2006 ( .A(n1274), .B(n1273), .Z(n1334) );
  NAND U2007 ( .A(n1276), .B(n1275), .Z(n1280) );
  NANDN U2008 ( .A(n1278), .B(n1277), .Z(n1279) );
  NAND U2009 ( .A(n1280), .B(n1279), .Z(n1332) );
  NANDN U2010 ( .A(n1282), .B(n1281), .Z(n1286) );
  NANDN U2011 ( .A(n1284), .B(n1283), .Z(n1285) );
  NAND U2012 ( .A(n1286), .B(n1285), .Z(n1339) );
  NANDN U2013 ( .A(n1288), .B(n1287), .Z(n1292) );
  NANDN U2014 ( .A(n1290), .B(n1289), .Z(n1291) );
  NAND U2015 ( .A(n1292), .B(n1291), .Z(n1338) );
  NANDN U2016 ( .A(n1294), .B(n1293), .Z(n1298) );
  NAND U2017 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U2018 ( .A(n1298), .B(n1297), .Z(n1375) );
  XOR U2019 ( .A(b[7]), .B(n11202), .Z(n1357) );
  NANDN U2020 ( .A(n1357), .B(n29949), .Z(n1301) );
  NANDN U2021 ( .A(n1299), .B(n29948), .Z(n1300) );
  NAND U2022 ( .A(n1301), .B(n1300), .Z(n1346) );
  NOR U2023 ( .A(b[9]), .B(b[10]), .Z(n1302) );
  OR U2024 ( .A(n1302), .B(n986), .Z(n1303) );
  NANDN U2025 ( .A(n969), .B(b[10]), .Z(n31367) );
  ANDN U2026 ( .B(n31367), .A(n970), .Z(n31890) );
  NAND U2027 ( .A(n1303), .B(n31890), .Z(n1343) );
  XOR U2028 ( .A(b[3]), .B(n12258), .Z(n1360) );
  NANDN U2029 ( .A(n1360), .B(n28939), .Z(n1306) );
  NAND U2030 ( .A(n1304), .B(n28938), .Z(n1305) );
  NAND U2031 ( .A(n1306), .B(n1305), .Z(n1344) );
  XOR U2032 ( .A(n1343), .B(n1344), .Z(n1345) );
  XNOR U2033 ( .A(n1346), .B(n1345), .Z(n1376) );
  XNOR U2034 ( .A(n1375), .B(n1376), .Z(n1377) );
  XOR U2035 ( .A(b[9]), .B(n10524), .Z(n1366) );
  NANDN U2036 ( .A(n1366), .B(n30509), .Z(n1309) );
  NAND U2037 ( .A(n1307), .B(n30846), .Z(n1308) );
  NAND U2038 ( .A(n1309), .B(n1308), .Z(n1356) );
  XNOR U2039 ( .A(n970), .B(b[9]), .Z(n1311) );
  XNOR U2040 ( .A(n970), .B(b[10]), .Z(n1310) );
  AND U2041 ( .A(n1311), .B(n1310), .Z(n31119) );
  NANDN U2042 ( .A(n1312), .B(n31119), .Z(n1314) );
  XOR U2043 ( .A(b[11]), .B(n10457), .Z(n1352) );
  OR U2044 ( .A(n1352), .B(n31369), .Z(n1313) );
  NAND U2045 ( .A(n1314), .B(n1313), .Z(n1355) );
  XNOR U2046 ( .A(n1356), .B(n1355), .Z(n1372) );
  NANDN U2047 ( .A(n966), .B(a[11]), .Z(n1315) );
  XOR U2048 ( .A(n29232), .B(n1315), .Z(n1317) );
  IV U2049 ( .A(a[10]), .Z(n12555) );
  NANDN U2050 ( .A(n12555), .B(n966), .Z(n1316) );
  AND U2051 ( .A(n1317), .B(n1316), .Z(n1370) );
  NAND U2052 ( .A(n29864), .B(n1318), .Z(n1320) );
  XOR U2053 ( .A(n968), .B(n11694), .Z(n1349) );
  NANDN U2054 ( .A(n29363), .B(n1349), .Z(n1319) );
  AND U2055 ( .A(n1320), .B(n1319), .Z(n1369) );
  XNOR U2056 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U2057 ( .A(n1372), .B(n1371), .Z(n1378) );
  XOR U2058 ( .A(n1377), .B(n1378), .Z(n1337) );
  XNOR U2059 ( .A(n1338), .B(n1337), .Z(n1340) );
  XNOR U2060 ( .A(n1339), .B(n1340), .Z(n1331) );
  XOR U2061 ( .A(n1332), .B(n1331), .Z(n1333) );
  XNOR U2062 ( .A(n1334), .B(n1333), .Z(n1326) );
  XNOR U2063 ( .A(n1326), .B(sreg[75]), .Z(n1328) );
  NAND U2064 ( .A(n1321), .B(sreg[74]), .Z(n1325) );
  OR U2065 ( .A(n1323), .B(n1322), .Z(n1324) );
  AND U2066 ( .A(n1325), .B(n1324), .Z(n1327) );
  XOR U2067 ( .A(n1328), .B(n1327), .Z(c[75]) );
  NAND U2068 ( .A(n1326), .B(sreg[75]), .Z(n1330) );
  OR U2069 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U2070 ( .A(n1330), .B(n1329), .Z(n1441) );
  XNOR U2071 ( .A(n1441), .B(sreg[76]), .Z(n1443) );
  NAND U2072 ( .A(n1332), .B(n1331), .Z(n1336) );
  NAND U2073 ( .A(n1334), .B(n1333), .Z(n1335) );
  NAND U2074 ( .A(n1336), .B(n1335), .Z(n1384) );
  NAND U2075 ( .A(n1338), .B(n1337), .Z(n1342) );
  NANDN U2076 ( .A(n1340), .B(n1339), .Z(n1341) );
  NAND U2077 ( .A(n1342), .B(n1341), .Z(n1381) );
  NANDN U2078 ( .A(n1344), .B(n1343), .Z(n1348) );
  OR U2079 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U2080 ( .A(n1348), .B(n1347), .Z(n1390) );
  NAND U2081 ( .A(n29864), .B(n1349), .Z(n1351) );
  XOR U2082 ( .A(n968), .B(n11986), .Z(n1424) );
  NANDN U2083 ( .A(n29363), .B(n1424), .Z(n1350) );
  NAND U2084 ( .A(n1351), .B(n1350), .Z(n1394) );
  XOR U2085 ( .A(b[11]), .B(n10363), .Z(n1427) );
  OR U2086 ( .A(n1427), .B(n31369), .Z(n1354) );
  NANDN U2087 ( .A(n1352), .B(n31119), .Z(n1353) );
  AND U2088 ( .A(n1354), .B(n1353), .Z(n1393) );
  XNOR U2089 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U2090 ( .A(n1356), .B(n1355), .Z(n1406) );
  XOR U2091 ( .A(b[7]), .B(n11406), .Z(n1438) );
  NANDN U2092 ( .A(n1438), .B(n29949), .Z(n1359) );
  NANDN U2093 ( .A(n1357), .B(n29948), .Z(n1358) );
  NAND U2094 ( .A(n1359), .B(n1358), .Z(n1404) );
  XNOR U2095 ( .A(n967), .B(a[10]), .Z(n1418) );
  NAND U2096 ( .A(n1418), .B(n28939), .Z(n1362) );
  NANDN U2097 ( .A(n1360), .B(n28938), .Z(n1361) );
  AND U2098 ( .A(n1362), .B(n1361), .Z(n1403) );
  XNOR U2099 ( .A(n1404), .B(n1403), .Z(n1405) );
  XNOR U2100 ( .A(n1406), .B(n1405), .Z(n1396) );
  XNOR U2101 ( .A(n1395), .B(n1396), .Z(n1399) );
  XOR U2102 ( .A(n970), .B(b[12]), .Z(n31550) );
  NOR U2103 ( .A(n986), .B(n31550), .Z(n1412) );
  NANDN U2104 ( .A(n966), .B(a[12]), .Z(n1363) );
  XOR U2105 ( .A(n29232), .B(n1363), .Z(n1365) );
  IV U2106 ( .A(a[11]), .Z(n12830) );
  NANDN U2107 ( .A(n12830), .B(n966), .Z(n1364) );
  AND U2108 ( .A(n1365), .B(n1364), .Z(n1410) );
  NANDN U2109 ( .A(n1366), .B(n30846), .Z(n1368) );
  XNOR U2110 ( .A(n969), .B(a[4]), .Z(n1421) );
  NAND U2111 ( .A(n30509), .B(n1421), .Z(n1367) );
  AND U2112 ( .A(n1368), .B(n1367), .Z(n1409) );
  XNOR U2113 ( .A(n1410), .B(n1409), .Z(n1411) );
  XOR U2114 ( .A(n1412), .B(n1411), .Z(n1397) );
  NANDN U2115 ( .A(n1370), .B(n1369), .Z(n1374) );
  NAND U2116 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U2117 ( .A(n1374), .B(n1373), .Z(n1398) );
  XOR U2118 ( .A(n1397), .B(n1398), .Z(n1400) );
  XOR U2119 ( .A(n1399), .B(n1400), .Z(n1388) );
  NANDN U2120 ( .A(n1376), .B(n1375), .Z(n1380) );
  NAND U2121 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U2122 ( .A(n1380), .B(n1379), .Z(n1387) );
  XOR U2123 ( .A(n1388), .B(n1387), .Z(n1389) );
  XNOR U2124 ( .A(n1390), .B(n1389), .Z(n1382) );
  XNOR U2125 ( .A(n1381), .B(n1382), .Z(n1383) );
  XOR U2126 ( .A(n1384), .B(n1383), .Z(n1442) );
  XOR U2127 ( .A(n1443), .B(n1442), .Z(c[76]) );
  NANDN U2128 ( .A(n1382), .B(n1381), .Z(n1386) );
  NAND U2129 ( .A(n1384), .B(n1383), .Z(n1385) );
  NAND U2130 ( .A(n1386), .B(n1385), .Z(n1454) );
  OR U2131 ( .A(n1388), .B(n1387), .Z(n1392) );
  NAND U2132 ( .A(n1390), .B(n1389), .Z(n1391) );
  NAND U2133 ( .A(n1392), .B(n1391), .Z(n1452) );
  NANDN U2134 ( .A(n1398), .B(n1397), .Z(n1402) );
  OR U2135 ( .A(n1400), .B(n1399), .Z(n1401) );
  NAND U2136 ( .A(n1402), .B(n1401), .Z(n1505) );
  XNOR U2137 ( .A(n1504), .B(n1505), .Z(n1506) );
  NANDN U2138 ( .A(n1404), .B(n1403), .Z(n1408) );
  NAND U2139 ( .A(n1406), .B(n1405), .Z(n1407) );
  NAND U2140 ( .A(n1408), .B(n1407), .Z(n1498) );
  NANDN U2141 ( .A(n1410), .B(n1409), .Z(n1414) );
  NANDN U2142 ( .A(n1412), .B(n1411), .Z(n1413) );
  AND U2143 ( .A(n1414), .B(n1413), .Z(n1499) );
  XNOR U2144 ( .A(n1498), .B(n1499), .Z(n1500) );
  NOR U2145 ( .A(b[11]), .B(b[12]), .Z(n1415) );
  NANDN U2146 ( .A(n971), .B(n1415), .Z(n1417) );
  ANDN U2147 ( .B(b[13]), .A(n31550), .Z(n31877) );
  NANDN U2148 ( .A(a[0]), .B(n31877), .Z(n1416) );
  NAND U2149 ( .A(n1417), .B(n1416), .Z(n1468) );
  XOR U2150 ( .A(n967), .B(n12830), .Z(n1463) );
  NAND U2151 ( .A(n28939), .B(n1463), .Z(n1420) );
  NAND U2152 ( .A(n1418), .B(n28938), .Z(n1419) );
  NAND U2153 ( .A(n1420), .B(n1419), .Z(n1466) );
  XOR U2154 ( .A(b[9]), .B(n11202), .Z(n1480) );
  NANDN U2155 ( .A(n1480), .B(n30509), .Z(n1423) );
  NAND U2156 ( .A(n1421), .B(n30846), .Z(n1422) );
  AND U2157 ( .A(n1423), .B(n1422), .Z(n1467) );
  XNOR U2158 ( .A(n1466), .B(n1467), .Z(n1469) );
  XOR U2159 ( .A(n1468), .B(n1469), .Z(n1492) );
  NAND U2160 ( .A(n29864), .B(n1424), .Z(n1426) );
  XNOR U2161 ( .A(n968), .B(a[9]), .Z(n1460) );
  NANDN U2162 ( .A(n29363), .B(n1460), .Z(n1425) );
  NAND U2163 ( .A(n1426), .B(n1425), .Z(n1493) );
  XOR U2164 ( .A(n1492), .B(n1493), .Z(n1494) );
  XOR U2165 ( .A(b[11]), .B(n10524), .Z(n1475) );
  OR U2166 ( .A(n1475), .B(n31369), .Z(n1429) );
  NANDN U2167 ( .A(n1427), .B(n31119), .Z(n1428) );
  NAND U2168 ( .A(n1429), .B(n1428), .Z(n1479) );
  XOR U2169 ( .A(n971), .B(n10457), .Z(n1483) );
  ANDN U2170 ( .B(n1483), .A(n31550), .Z(n1434) );
  XNOR U2171 ( .A(n971), .B(a[0]), .Z(n1432) );
  XNOR U2172 ( .A(n971), .B(b[11]), .Z(n1431) );
  XNOR U2173 ( .A(n971), .B(b[12]), .Z(n1430) );
  AND U2174 ( .A(n1431), .B(n1430), .Z(n31874) );
  NAND U2175 ( .A(n1432), .B(n31874), .Z(n1433) );
  NANDN U2176 ( .A(n1434), .B(n1433), .Z(n1478) );
  XNOR U2177 ( .A(n1479), .B(n1478), .Z(n1489) );
  NANDN U2178 ( .A(n966), .B(a[13]), .Z(n1435) );
  XOR U2179 ( .A(n29232), .B(n1435), .Z(n1437) );
  IV U2180 ( .A(a[12]), .Z(n13106) );
  NANDN U2181 ( .A(n13106), .B(n966), .Z(n1436) );
  AND U2182 ( .A(n1437), .B(n1436), .Z(n1487) );
  XOR U2183 ( .A(b[7]), .B(n11694), .Z(n1457) );
  NANDN U2184 ( .A(n1457), .B(n29949), .Z(n1440) );
  NANDN U2185 ( .A(n1438), .B(n29948), .Z(n1439) );
  AND U2186 ( .A(n1440), .B(n1439), .Z(n1486) );
  XNOR U2187 ( .A(n1487), .B(n1486), .Z(n1488) );
  XOR U2188 ( .A(n1489), .B(n1488), .Z(n1495) );
  XOR U2189 ( .A(n1494), .B(n1495), .Z(n1501) );
  XOR U2190 ( .A(n1500), .B(n1501), .Z(n1507) );
  XOR U2191 ( .A(n1506), .B(n1507), .Z(n1451) );
  XOR U2192 ( .A(n1452), .B(n1451), .Z(n1453) );
  XNOR U2193 ( .A(n1454), .B(n1453), .Z(n1446) );
  XNOR U2194 ( .A(n1446), .B(sreg[77]), .Z(n1448) );
  NAND U2195 ( .A(n1441), .B(sreg[76]), .Z(n1445) );
  OR U2196 ( .A(n1443), .B(n1442), .Z(n1444) );
  AND U2197 ( .A(n1445), .B(n1444), .Z(n1447) );
  XOR U2198 ( .A(n1448), .B(n1447), .Z(c[77]) );
  NAND U2199 ( .A(n1446), .B(sreg[77]), .Z(n1450) );
  OR U2200 ( .A(n1448), .B(n1447), .Z(n1449) );
  NAND U2201 ( .A(n1450), .B(n1449), .Z(n1577) );
  XNOR U2202 ( .A(n1577), .B(sreg[78]), .Z(n1579) );
  NAND U2203 ( .A(n1452), .B(n1451), .Z(n1456) );
  NAND U2204 ( .A(n1454), .B(n1453), .Z(n1455) );
  NAND U2205 ( .A(n1456), .B(n1455), .Z(n1513) );
  XOR U2206 ( .A(b[7]), .B(n11986), .Z(n1568) );
  NANDN U2207 ( .A(n1568), .B(n29949), .Z(n1459) );
  NANDN U2208 ( .A(n1457), .B(n29948), .Z(n1458) );
  AND U2209 ( .A(n1459), .B(n1458), .Z(n1538) );
  XOR U2210 ( .A(n968), .B(n12555), .Z(n1562) );
  NANDN U2211 ( .A(n29363), .B(n1562), .Z(n1462) );
  NAND U2212 ( .A(n1460), .B(n29864), .Z(n1461) );
  AND U2213 ( .A(n1462), .B(n1461), .Z(n1539) );
  XOR U2214 ( .A(n1538), .B(n1539), .Z(n1540) );
  XOR U2215 ( .A(b[3]), .B(n13106), .Z(n1565) );
  NANDN U2216 ( .A(n1565), .B(n28939), .Z(n1465) );
  NAND U2217 ( .A(n1463), .B(n28938), .Z(n1464) );
  AND U2218 ( .A(n1465), .B(n1464), .Z(n1541) );
  XNOR U2219 ( .A(n1540), .B(n1541), .Z(n1528) );
  NANDN U2220 ( .A(n1467), .B(n1466), .Z(n1471) );
  NAND U2221 ( .A(n1469), .B(n1468), .Z(n1470) );
  NAND U2222 ( .A(n1471), .B(n1470), .Z(n1529) );
  XOR U2223 ( .A(n1528), .B(n1529), .Z(n1530) );
  NANDN U2224 ( .A(n966), .B(a[14]), .Z(n1472) );
  XOR U2225 ( .A(n29232), .B(n1472), .Z(n1474) );
  IV U2226 ( .A(a[13]), .Z(n13509) );
  NANDN U2227 ( .A(n13509), .B(n966), .Z(n1473) );
  AND U2228 ( .A(n1474), .B(n1473), .Z(n1523) );
  XOR U2229 ( .A(b[11]), .B(n10854), .Z(n1559) );
  OR U2230 ( .A(n1559), .B(n31369), .Z(n1477) );
  NANDN U2231 ( .A(n1475), .B(n31119), .Z(n1476) );
  NAND U2232 ( .A(n1477), .B(n1476), .Z(n1522) );
  XOR U2233 ( .A(n1523), .B(n1522), .Z(n1524) );
  XOR U2234 ( .A(b[13]), .B(b[14]), .Z(n1550) );
  AND U2235 ( .A(a[0]), .B(n1550), .Z(n1525) );
  XOR U2236 ( .A(n1524), .B(n1525), .Z(n1531) );
  XOR U2237 ( .A(n1530), .B(n1531), .Z(n1574) );
  NAND U2238 ( .A(n1479), .B(n1478), .Z(n1536) );
  NANDN U2239 ( .A(n1480), .B(n30846), .Z(n1482) );
  XOR U2240 ( .A(n969), .B(n11406), .Z(n1556) );
  NAND U2241 ( .A(n30509), .B(n1556), .Z(n1481) );
  NAND U2242 ( .A(n1482), .B(n1481), .Z(n1535) );
  NAND U2243 ( .A(n31874), .B(n1483), .Z(n1485) );
  XNOR U2244 ( .A(n971), .B(a[2]), .Z(n1544) );
  NANDN U2245 ( .A(n31550), .B(n1544), .Z(n1484) );
  AND U2246 ( .A(n1485), .B(n1484), .Z(n1534) );
  XNOR U2247 ( .A(n1535), .B(n1534), .Z(n1537) );
  XNOR U2248 ( .A(n1536), .B(n1537), .Z(n1571) );
  NANDN U2249 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U2250 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U2251 ( .A(n1491), .B(n1490), .Z(n1572) );
  XNOR U2252 ( .A(n1571), .B(n1572), .Z(n1573) );
  XNOR U2253 ( .A(n1574), .B(n1573), .Z(n1517) );
  OR U2254 ( .A(n1493), .B(n1492), .Z(n1497) );
  NAND U2255 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U2256 ( .A(n1497), .B(n1496), .Z(n1516) );
  XNOR U2257 ( .A(n1517), .B(n1516), .Z(n1518) );
  NANDN U2258 ( .A(n1499), .B(n1498), .Z(n1503) );
  NAND U2259 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U2260 ( .A(n1503), .B(n1502), .Z(n1519) );
  XOR U2261 ( .A(n1518), .B(n1519), .Z(n1510) );
  NANDN U2262 ( .A(n1505), .B(n1504), .Z(n1509) );
  NAND U2263 ( .A(n1507), .B(n1506), .Z(n1508) );
  AND U2264 ( .A(n1509), .B(n1508), .Z(n1511) );
  XNOR U2265 ( .A(n1510), .B(n1511), .Z(n1512) );
  XOR U2266 ( .A(n1513), .B(n1512), .Z(n1578) );
  XOR U2267 ( .A(n1579), .B(n1578), .Z(c[78]) );
  NANDN U2268 ( .A(n1511), .B(n1510), .Z(n1515) );
  NAND U2269 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND U2270 ( .A(n1515), .B(n1514), .Z(n1590) );
  NANDN U2271 ( .A(n1517), .B(n1516), .Z(n1521) );
  NANDN U2272 ( .A(n1519), .B(n1518), .Z(n1520) );
  NAND U2273 ( .A(n1521), .B(n1520), .Z(n1587) );
  OR U2274 ( .A(n1523), .B(n1522), .Z(n1527) );
  NANDN U2275 ( .A(n1525), .B(n1524), .Z(n1526) );
  NAND U2276 ( .A(n1527), .B(n1526), .Z(n1644) );
  OR U2277 ( .A(n1529), .B(n1528), .Z(n1533) );
  NANDN U2278 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U2279 ( .A(n1533), .B(n1532), .Z(n1641) );
  XNOR U2280 ( .A(n1641), .B(n1642), .Z(n1643) );
  XNOR U2281 ( .A(n1644), .B(n1643), .Z(n1596) );
  OR U2282 ( .A(n1539), .B(n1538), .Z(n1543) );
  NANDN U2283 ( .A(n1541), .B(n1540), .Z(n1542) );
  NAND U2284 ( .A(n1543), .B(n1542), .Z(n1648) );
  XOR U2285 ( .A(b[13]), .B(n10524), .Z(n1632) );
  OR U2286 ( .A(n1632), .B(n31550), .Z(n1546) );
  NAND U2287 ( .A(n1544), .B(n31874), .Z(n1545) );
  NAND U2288 ( .A(n1546), .B(n1545), .Z(n1612) );
  XNOR U2289 ( .A(n972), .B(a[0]), .Z(n1549) );
  XNOR U2290 ( .A(n972), .B(b[13]), .Z(n1548) );
  XNOR U2291 ( .A(n972), .B(b[14]), .Z(n1547) );
  AND U2292 ( .A(n1548), .B(n1547), .Z(n32011) );
  NAND U2293 ( .A(n1549), .B(n32011), .Z(n1552) );
  IV U2294 ( .A(n1550), .Z(n32010) );
  XNOR U2295 ( .A(n972), .B(a[1]), .Z(n1605) );
  NANDN U2296 ( .A(n32010), .B(n1605), .Z(n1551) );
  NAND U2297 ( .A(n1552), .B(n1551), .Z(n1611) );
  XNOR U2298 ( .A(n1612), .B(n1611), .Z(n1638) );
  NANDN U2299 ( .A(n966), .B(a[15]), .Z(n1553) );
  XOR U2300 ( .A(n29232), .B(n1553), .Z(n1555) );
  IV U2301 ( .A(a[14]), .Z(n14210) );
  NANDN U2302 ( .A(n14210), .B(n966), .Z(n1554) );
  AND U2303 ( .A(n1555), .B(n1554), .Z(n1636) );
  NAND U2304 ( .A(n30846), .B(n1556), .Z(n1558) );
  XOR U2305 ( .A(n969), .B(n11694), .Z(n1613) );
  NAND U2306 ( .A(n30509), .B(n1613), .Z(n1557) );
  AND U2307 ( .A(n1558), .B(n1557), .Z(n1635) );
  XNOR U2308 ( .A(n1636), .B(n1635), .Z(n1637) );
  XOR U2309 ( .A(n1638), .B(n1637), .Z(n1647) );
  XNOR U2310 ( .A(n1648), .B(n1647), .Z(n1649) );
  XNOR U2311 ( .A(n970), .B(a[5]), .Z(n1602) );
  NANDN U2312 ( .A(n31369), .B(n1602), .Z(n1561) );
  NANDN U2313 ( .A(n1559), .B(n31119), .Z(n1560) );
  NAND U2314 ( .A(n1561), .B(n1560), .Z(n1627) );
  NAND U2315 ( .A(n29864), .B(n1562), .Z(n1564) );
  XNOR U2316 ( .A(n968), .B(a[11]), .Z(n1599) );
  NANDN U2317 ( .A(n29363), .B(n1599), .Z(n1563) );
  NAND U2318 ( .A(n1564), .B(n1563), .Z(n1625) );
  XOR U2319 ( .A(b[3]), .B(n13509), .Z(n1616) );
  NANDN U2320 ( .A(n1616), .B(n28939), .Z(n1567) );
  NANDN U2321 ( .A(n1565), .B(n28938), .Z(n1566) );
  NAND U2322 ( .A(n1567), .B(n1566), .Z(n1626) );
  XNOR U2323 ( .A(n1625), .B(n1626), .Z(n1628) );
  XOR U2324 ( .A(n1627), .B(n1628), .Z(n1622) );
  XOR U2325 ( .A(b[7]), .B(n12258), .Z(n1608) );
  NANDN U2326 ( .A(n1608), .B(n29949), .Z(n1570) );
  NANDN U2327 ( .A(n1568), .B(n29948), .Z(n1569) );
  NAND U2328 ( .A(n1570), .B(n1569), .Z(n1620) );
  XNOR U2329 ( .A(n1619), .B(n1620), .Z(n1621) );
  XOR U2330 ( .A(n1622), .B(n1621), .Z(n1650) );
  XOR U2331 ( .A(n1649), .B(n1650), .Z(n1593) );
  NANDN U2332 ( .A(n1572), .B(n1571), .Z(n1576) );
  NAND U2333 ( .A(n1574), .B(n1573), .Z(n1575) );
  AND U2334 ( .A(n1576), .B(n1575), .Z(n1594) );
  XOR U2335 ( .A(n1593), .B(n1594), .Z(n1595) );
  XOR U2336 ( .A(n1596), .B(n1595), .Z(n1588) );
  XOR U2337 ( .A(n1587), .B(n1588), .Z(n1589) );
  XNOR U2338 ( .A(n1590), .B(n1589), .Z(n1582) );
  XNOR U2339 ( .A(n1582), .B(sreg[79]), .Z(n1584) );
  NAND U2340 ( .A(n1577), .B(sreg[78]), .Z(n1581) );
  OR U2341 ( .A(n1579), .B(n1578), .Z(n1580) );
  AND U2342 ( .A(n1581), .B(n1580), .Z(n1583) );
  XOR U2343 ( .A(n1584), .B(n1583), .Z(c[79]) );
  NAND U2344 ( .A(n1582), .B(sreg[79]), .Z(n1586) );
  OR U2345 ( .A(n1584), .B(n1583), .Z(n1585) );
  NAND U2346 ( .A(n1586), .B(n1585), .Z(n1730) );
  XNOR U2347 ( .A(n1730), .B(sreg[80]), .Z(n1732) );
  OR U2348 ( .A(n1588), .B(n1587), .Z(n1592) );
  NAND U2349 ( .A(n1590), .B(n1589), .Z(n1591) );
  NAND U2350 ( .A(n1592), .B(n1591), .Z(n1654) );
  NAND U2351 ( .A(n1594), .B(n1593), .Z(n1598) );
  NANDN U2352 ( .A(n1596), .B(n1595), .Z(n1597) );
  NAND U2353 ( .A(n1598), .B(n1597), .Z(n1651) );
  XOR U2354 ( .A(b[5]), .B(n13106), .Z(n1700) );
  OR U2355 ( .A(n1700), .B(n29363), .Z(n1601) );
  NAND U2356 ( .A(n1599), .B(n29864), .Z(n1600) );
  NAND U2357 ( .A(n1601), .B(n1600), .Z(n1727) );
  XOR U2358 ( .A(b[11]), .B(n11406), .Z(n1712) );
  OR U2359 ( .A(n1712), .B(n31369), .Z(n1604) );
  NAND U2360 ( .A(n1602), .B(n31119), .Z(n1603) );
  NAND U2361 ( .A(n1604), .B(n1603), .Z(n1724) );
  XOR U2362 ( .A(b[15]), .B(n10363), .Z(n1686) );
  OR U2363 ( .A(n1686), .B(n32010), .Z(n1607) );
  NAND U2364 ( .A(n1605), .B(n32011), .Z(n1606) );
  AND U2365 ( .A(n1607), .B(n1606), .Z(n1725) );
  XNOR U2366 ( .A(n1724), .B(n1725), .Z(n1726) );
  XNOR U2367 ( .A(n1727), .B(n1726), .Z(n1703) );
  XNOR U2368 ( .A(n31123), .B(a[10]), .Z(n1709) );
  NAND U2369 ( .A(n1709), .B(n29949), .Z(n1610) );
  NANDN U2370 ( .A(n1608), .B(n29948), .Z(n1609) );
  NAND U2371 ( .A(n1610), .B(n1609), .Z(n1704) );
  XOR U2372 ( .A(n1703), .B(n1704), .Z(n1706) );
  NAND U2373 ( .A(n1612), .B(n1611), .Z(n1721) );
  NAND U2374 ( .A(n30846), .B(n1613), .Z(n1615) );
  XOR U2375 ( .A(n969), .B(n11986), .Z(n1683) );
  NAND U2376 ( .A(n30509), .B(n1683), .Z(n1614) );
  NAND U2377 ( .A(n1615), .B(n1614), .Z(n1719) );
  XOR U2378 ( .A(b[3]), .B(n14210), .Z(n1697) );
  NANDN U2379 ( .A(n1697), .B(n28939), .Z(n1618) );
  NANDN U2380 ( .A(n1616), .B(n28938), .Z(n1617) );
  AND U2381 ( .A(n1618), .B(n1617), .Z(n1718) );
  XNOR U2382 ( .A(n1719), .B(n1718), .Z(n1720) );
  XNOR U2383 ( .A(n1721), .B(n1720), .Z(n1705) );
  XNOR U2384 ( .A(n1706), .B(n1705), .Z(n1663) );
  NANDN U2385 ( .A(n1620), .B(n1619), .Z(n1624) );
  NAND U2386 ( .A(n1622), .B(n1621), .Z(n1623) );
  NAND U2387 ( .A(n1624), .B(n1623), .Z(n1664) );
  XNOR U2388 ( .A(n1663), .B(n1664), .Z(n1665) );
  NANDN U2389 ( .A(n966), .B(a[16]), .Z(n1629) );
  XOR U2390 ( .A(n29232), .B(n1629), .Z(n1631) );
  IV U2391 ( .A(a[15]), .Z(n13976) );
  NANDN U2392 ( .A(n13976), .B(n966), .Z(n1630) );
  AND U2393 ( .A(n1631), .B(n1630), .Z(n1677) );
  XOR U2394 ( .A(n971), .B(n10854), .Z(n1715) );
  NANDN U2395 ( .A(n31550), .B(n1715), .Z(n1634) );
  NANDN U2396 ( .A(n1632), .B(n31874), .Z(n1633) );
  NAND U2397 ( .A(n1634), .B(n1633), .Z(n1675) );
  XOR U2398 ( .A(b[16]), .B(b[15]), .Z(n32543) );
  NANDN U2399 ( .A(n986), .B(n32543), .Z(n1676) );
  XNOR U2400 ( .A(n1675), .B(n1676), .Z(n1678) );
  XOR U2401 ( .A(n1677), .B(n1678), .Z(n1669) );
  NANDN U2402 ( .A(n1636), .B(n1635), .Z(n1640) );
  NAND U2403 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U2404 ( .A(n1640), .B(n1639), .Z(n1670) );
  XNOR U2405 ( .A(n1669), .B(n1670), .Z(n1672) );
  XOR U2406 ( .A(n1671), .B(n1672), .Z(n1666) );
  XOR U2407 ( .A(n1665), .B(n1666), .Z(n1660) );
  NANDN U2408 ( .A(n1642), .B(n1641), .Z(n1646) );
  NAND U2409 ( .A(n1644), .B(n1643), .Z(n1645) );
  NAND U2410 ( .A(n1646), .B(n1645), .Z(n1657) );
  XNOR U2411 ( .A(n1657), .B(n1658), .Z(n1659) );
  XNOR U2412 ( .A(n1660), .B(n1659), .Z(n1652) );
  XNOR U2413 ( .A(n1651), .B(n1652), .Z(n1653) );
  XOR U2414 ( .A(n1654), .B(n1653), .Z(n1731) );
  XOR U2415 ( .A(n1732), .B(n1731), .Z(c[80]) );
  NANDN U2416 ( .A(n1652), .B(n1651), .Z(n1656) );
  NAND U2417 ( .A(n1654), .B(n1653), .Z(n1655) );
  NAND U2418 ( .A(n1656), .B(n1655), .Z(n1743) );
  NANDN U2419 ( .A(n1658), .B(n1657), .Z(n1662) );
  NAND U2420 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U2421 ( .A(n1662), .B(n1661), .Z(n1741) );
  NANDN U2422 ( .A(n1664), .B(n1663), .Z(n1668) );
  NANDN U2423 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U2424 ( .A(n1668), .B(n1667), .Z(n1747) );
  NAND U2425 ( .A(n1670), .B(n1669), .Z(n1674) );
  NANDN U2426 ( .A(n1672), .B(n1671), .Z(n1673) );
  AND U2427 ( .A(n1674), .B(n1673), .Z(n1746) );
  XNOR U2428 ( .A(n1747), .B(n1746), .Z(n1748) );
  NANDN U2429 ( .A(n1676), .B(n1675), .Z(n1680) );
  NAND U2430 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U2431 ( .A(n1680), .B(n1679), .Z(n1798) );
  ANDN U2432 ( .B(n972), .A(b[16]), .Z(n1681) );
  OR U2433 ( .A(n1681), .B(n986), .Z(n1682) );
  NANDN U2434 ( .A(n972), .B(b[16]), .Z(n32809) );
  AND U2435 ( .A(n32809), .B(b[17]), .Z(n33153) );
  AND U2436 ( .A(n1682), .B(n33153), .Z(n1759) );
  NAND U2437 ( .A(n30846), .B(n1683), .Z(n1685) );
  XNOR U2438 ( .A(n969), .B(a[9]), .Z(n1783) );
  NAND U2439 ( .A(n30509), .B(n1783), .Z(n1684) );
  NAND U2440 ( .A(n1685), .B(n1684), .Z(n1758) );
  XOR U2441 ( .A(n1759), .B(n1758), .Z(n1760) );
  XOR U2442 ( .A(b[15]), .B(n10524), .Z(n1777) );
  OR U2443 ( .A(n1777), .B(n32010), .Z(n1688) );
  NANDN U2444 ( .A(n1686), .B(n32011), .Z(n1687) );
  NAND U2445 ( .A(n1688), .B(n1687), .Z(n1765) );
  XOR U2446 ( .A(n986), .B(b[16]), .Z(n1689) );
  XOR U2447 ( .A(b[16]), .B(n972), .Z(n32811) );
  NAND U2448 ( .A(n1689), .B(n32811), .Z(n1691) );
  XNOR U2449 ( .A(b[17]), .B(b[16]), .Z(n1690) );
  OR U2450 ( .A(n1691), .B(n1690), .Z(n1693) );
  XNOR U2451 ( .A(b[17]), .B(a[1]), .Z(n1768) );
  NANDN U2452 ( .A(n1768), .B(n32543), .Z(n1692) );
  NAND U2453 ( .A(n1693), .B(n1692), .Z(n1764) );
  XOR U2454 ( .A(n1765), .B(n1764), .Z(n1761) );
  XOR U2455 ( .A(n1760), .B(n1761), .Z(n1795) );
  NANDN U2456 ( .A(n966), .B(a[17]), .Z(n1694) );
  XOR U2457 ( .A(n29232), .B(n1694), .Z(n1696) );
  IV U2458 ( .A(a[16]), .Z(n14259) );
  NANDN U2459 ( .A(n14259), .B(n966), .Z(n1695) );
  AND U2460 ( .A(n1696), .B(n1695), .Z(n1803) );
  XNOR U2461 ( .A(n967), .B(a[15]), .Z(n1780) );
  NAND U2462 ( .A(n1780), .B(n28939), .Z(n1699) );
  NANDN U2463 ( .A(n1697), .B(n28938), .Z(n1698) );
  NAND U2464 ( .A(n1699), .B(n1698), .Z(n1801) );
  XOR U2465 ( .A(n968), .B(n13509), .Z(n1789) );
  NANDN U2466 ( .A(n29363), .B(n1789), .Z(n1702) );
  NANDN U2467 ( .A(n1700), .B(n29864), .Z(n1701) );
  AND U2468 ( .A(n1702), .B(n1701), .Z(n1802) );
  XNOR U2469 ( .A(n1801), .B(n1802), .Z(n1804) );
  XNOR U2470 ( .A(n1803), .B(n1804), .Z(n1796) );
  XNOR U2471 ( .A(n1795), .B(n1796), .Z(n1797) );
  XNOR U2472 ( .A(n1798), .B(n1797), .Z(n1813) );
  NANDN U2473 ( .A(n1704), .B(n1703), .Z(n1708) );
  OR U2474 ( .A(n1706), .B(n1705), .Z(n1707) );
  NAND U2475 ( .A(n1708), .B(n1707), .Z(n1812) );
  XOR U2476 ( .A(b[7]), .B(n12830), .Z(n1792) );
  NANDN U2477 ( .A(n1792), .B(n29949), .Z(n1711) );
  NAND U2478 ( .A(n1709), .B(n29948), .Z(n1710) );
  NAND U2479 ( .A(n1711), .B(n1710), .Z(n1755) );
  XOR U2480 ( .A(b[11]), .B(n11694), .Z(n1771) );
  OR U2481 ( .A(n1771), .B(n31369), .Z(n1714) );
  NANDN U2482 ( .A(n1712), .B(n31119), .Z(n1713) );
  NAND U2483 ( .A(n1714), .B(n1713), .Z(n1752) );
  XOR U2484 ( .A(b[13]), .B(n11202), .Z(n1786) );
  OR U2485 ( .A(n1786), .B(n31550), .Z(n1717) );
  NAND U2486 ( .A(n1715), .B(n31874), .Z(n1716) );
  AND U2487 ( .A(n1717), .B(n1716), .Z(n1753) );
  XNOR U2488 ( .A(n1752), .B(n1753), .Z(n1754) );
  XNOR U2489 ( .A(n1755), .B(n1754), .Z(n1808) );
  NANDN U2490 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U2491 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2492 ( .A(n1723), .B(n1722), .Z(n1805) );
  NANDN U2493 ( .A(n1725), .B(n1724), .Z(n1729) );
  NAND U2494 ( .A(n1727), .B(n1726), .Z(n1728) );
  NAND U2495 ( .A(n1729), .B(n1728), .Z(n1806) );
  XNOR U2496 ( .A(n1805), .B(n1806), .Z(n1807) );
  XOR U2497 ( .A(n1808), .B(n1807), .Z(n1811) );
  XNOR U2498 ( .A(n1812), .B(n1811), .Z(n1814) );
  XOR U2499 ( .A(n1813), .B(n1814), .Z(n1749) );
  XNOR U2500 ( .A(n1748), .B(n1749), .Z(n1740) );
  XOR U2501 ( .A(n1741), .B(n1740), .Z(n1742) );
  XNOR U2502 ( .A(n1743), .B(n1742), .Z(n1735) );
  XNOR U2503 ( .A(n1735), .B(sreg[81]), .Z(n1737) );
  NAND U2504 ( .A(n1730), .B(sreg[80]), .Z(n1734) );
  OR U2505 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U2506 ( .A(n1734), .B(n1733), .Z(n1736) );
  XOR U2507 ( .A(n1737), .B(n1736), .Z(c[81]) );
  NAND U2508 ( .A(n1735), .B(sreg[81]), .Z(n1739) );
  OR U2509 ( .A(n1737), .B(n1736), .Z(n1738) );
  NAND U2510 ( .A(n1739), .B(n1738), .Z(n1904) );
  XNOR U2511 ( .A(n1904), .B(sreg[82]), .Z(n1906) );
  NAND U2512 ( .A(n1741), .B(n1740), .Z(n1745) );
  NAND U2513 ( .A(n1743), .B(n1742), .Z(n1744) );
  NAND U2514 ( .A(n1745), .B(n1744), .Z(n1820) );
  NANDN U2515 ( .A(n1747), .B(n1746), .Z(n1751) );
  NANDN U2516 ( .A(n1749), .B(n1748), .Z(n1750) );
  NAND U2517 ( .A(n1751), .B(n1750), .Z(n1817) );
  NANDN U2518 ( .A(n1753), .B(n1752), .Z(n1757) );
  NAND U2519 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U2520 ( .A(n1757), .B(n1756), .Z(n1895) );
  OR U2521 ( .A(n1759), .B(n1758), .Z(n1763) );
  NANDN U2522 ( .A(n1761), .B(n1760), .Z(n1762) );
  NAND U2523 ( .A(n1763), .B(n1762), .Z(n1823) );
  NAND U2524 ( .A(n1765), .B(n1764), .Z(n1852) );
  XNOR U2525 ( .A(b[17]), .B(n10363), .Z(n1836) );
  NAND U2526 ( .A(n1836), .B(n32543), .Z(n1770) );
  XOR U2527 ( .A(b[17]), .B(b[16]), .Z(n1767) );
  XNOR U2528 ( .A(b[17]), .B(n972), .Z(n1766) );
  AND U2529 ( .A(n1767), .B(n1766), .Z(n32541) );
  NANDN U2530 ( .A(n1768), .B(n32541), .Z(n1769) );
  NAND U2531 ( .A(n1770), .B(n1769), .Z(n1850) );
  XNOR U2532 ( .A(n970), .B(a[8]), .Z(n1870) );
  NANDN U2533 ( .A(n31369), .B(n1870), .Z(n1773) );
  NANDN U2534 ( .A(n1771), .B(n31119), .Z(n1772) );
  AND U2535 ( .A(n1773), .B(n1772), .Z(n1849) );
  XNOR U2536 ( .A(n1850), .B(n1849), .Z(n1851) );
  XNOR U2537 ( .A(n1852), .B(n1851), .Z(n1824) );
  XNOR U2538 ( .A(n1823), .B(n1824), .Z(n1825) );
  NANDN U2539 ( .A(n966), .B(a[18]), .Z(n1774) );
  XOR U2540 ( .A(n29232), .B(n1774), .Z(n1776) );
  IV U2541 ( .A(a[17]), .Z(n14514) );
  NANDN U2542 ( .A(n14514), .B(n966), .Z(n1775) );
  AND U2543 ( .A(n1776), .B(n1775), .Z(n1883) );
  XOR U2544 ( .A(b[15]), .B(n10854), .Z(n1867) );
  OR U2545 ( .A(n1867), .B(n32010), .Z(n1779) );
  NANDN U2546 ( .A(n1777), .B(n32011), .Z(n1778) );
  NAND U2547 ( .A(n1779), .B(n1778), .Z(n1882) );
  XOR U2548 ( .A(n1883), .B(n1882), .Z(n1884) );
  XOR U2549 ( .A(b[17]), .B(b[18]), .Z(n1830) );
  AND U2550 ( .A(a[0]), .B(n1830), .Z(n1885) );
  XOR U2551 ( .A(n1884), .B(n1885), .Z(n1826) );
  XNOR U2552 ( .A(n1825), .B(n1826), .Z(n1894) );
  XNOR U2553 ( .A(n1895), .B(n1894), .Z(n1897) );
  XOR U2554 ( .A(n967), .B(n14259), .Z(n1876) );
  NAND U2555 ( .A(n1876), .B(n28939), .Z(n1782) );
  NAND U2556 ( .A(n1780), .B(n28938), .Z(n1781) );
  NAND U2557 ( .A(n1782), .B(n1781), .Z(n1846) );
  XOR U2558 ( .A(n969), .B(n12555), .Z(n1833) );
  NAND U2559 ( .A(n30509), .B(n1833), .Z(n1785) );
  NAND U2560 ( .A(n1783), .B(n30846), .Z(n1784) );
  NAND U2561 ( .A(n1785), .B(n1784), .Z(n1843) );
  XOR U2562 ( .A(b[13]), .B(n11406), .Z(n1864) );
  OR U2563 ( .A(n1864), .B(n31550), .Z(n1788) );
  NANDN U2564 ( .A(n1786), .B(n31874), .Z(n1787) );
  AND U2565 ( .A(n1788), .B(n1787), .Z(n1844) );
  XNOR U2566 ( .A(n1843), .B(n1844), .Z(n1845) );
  XNOR U2567 ( .A(n1846), .B(n1845), .Z(n1858) );
  NAND U2568 ( .A(n29864), .B(n1789), .Z(n1791) );
  XNOR U2569 ( .A(n968), .B(a[14]), .Z(n1861) );
  NANDN U2570 ( .A(n29363), .B(n1861), .Z(n1790) );
  NAND U2571 ( .A(n1791), .B(n1790), .Z(n1856) );
  XOR U2572 ( .A(b[7]), .B(n13106), .Z(n1879) );
  NANDN U2573 ( .A(n1879), .B(n29949), .Z(n1794) );
  NANDN U2574 ( .A(n1792), .B(n29948), .Z(n1793) );
  AND U2575 ( .A(n1794), .B(n1793), .Z(n1855) );
  XNOR U2576 ( .A(n1856), .B(n1855), .Z(n1857) );
  XOR U2577 ( .A(n1858), .B(n1857), .Z(n1896) );
  XNOR U2578 ( .A(n1897), .B(n1896), .Z(n1891) );
  NANDN U2579 ( .A(n1796), .B(n1795), .Z(n1800) );
  NAND U2580 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U2581 ( .A(n1800), .B(n1799), .Z(n1889) );
  XNOR U2582 ( .A(n1889), .B(n1888), .Z(n1890) );
  XOR U2583 ( .A(n1891), .B(n1890), .Z(n1898) );
  NANDN U2584 ( .A(n1806), .B(n1805), .Z(n1810) );
  NAND U2585 ( .A(n1808), .B(n1807), .Z(n1809) );
  NAND U2586 ( .A(n1810), .B(n1809), .Z(n1899) );
  XNOR U2587 ( .A(n1898), .B(n1899), .Z(n1900) );
  NAND U2588 ( .A(n1812), .B(n1811), .Z(n1816) );
  NANDN U2589 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U2590 ( .A(n1816), .B(n1815), .Z(n1901) );
  XNOR U2591 ( .A(n1900), .B(n1901), .Z(n1818) );
  XNOR U2592 ( .A(n1817), .B(n1818), .Z(n1819) );
  XOR U2593 ( .A(n1820), .B(n1819), .Z(n1905) );
  XOR U2594 ( .A(n1906), .B(n1905), .Z(c[82]) );
  NANDN U2595 ( .A(n1818), .B(n1817), .Z(n1822) );
  NAND U2596 ( .A(n1820), .B(n1819), .Z(n1821) );
  NAND U2597 ( .A(n1822), .B(n1821), .Z(n1917) );
  NANDN U2598 ( .A(n1824), .B(n1823), .Z(n1828) );
  NANDN U2599 ( .A(n1826), .B(n1825), .Z(n1827) );
  NAND U2600 ( .A(n1828), .B(n1827), .Z(n1918) );
  IV U2601 ( .A(b[19]), .Z(n33020) );
  OR U2602 ( .A(b[17]), .B(n33020), .Z(n1829) );
  OR U2603 ( .A(n1829), .B(b[18]), .Z(n1832) );
  IV U2604 ( .A(n1830), .Z(n33021) );
  ANDN U2605 ( .B(b[19]), .A(n33021), .Z(n33284) );
  NANDN U2606 ( .A(a[0]), .B(n33284), .Z(n1831) );
  NAND U2607 ( .A(n1832), .B(n1831), .Z(n1925) );
  NAND U2608 ( .A(n30846), .B(n1833), .Z(n1835) );
  XNOR U2609 ( .A(n969), .B(a[11]), .Z(n1957) );
  NAND U2610 ( .A(n30509), .B(n1957), .Z(n1834) );
  AND U2611 ( .A(n1835), .B(n1834), .Z(n1924) );
  XNOR U2612 ( .A(n1925), .B(n1924), .Z(n1926) );
  XNOR U2613 ( .A(b[17]), .B(n10524), .Z(n1948) );
  NAND U2614 ( .A(n1948), .B(n32543), .Z(n1838) );
  NAND U2615 ( .A(n1836), .B(n32541), .Z(n1837) );
  NAND U2616 ( .A(n1838), .B(n1837), .Z(n1965) );
  XNOR U2617 ( .A(n33020), .B(b[17]), .Z(n1967) );
  XNOR U2618 ( .A(n33020), .B(a[0]), .Z(n1839) );
  NAND U2619 ( .A(n1967), .B(n1839), .Z(n1840) );
  XNOR U2620 ( .A(n33020), .B(b[18]), .Z(n1966) );
  NANDN U2621 ( .A(n1840), .B(n1966), .Z(n1842) );
  XOR U2622 ( .A(b[19]), .B(n10457), .Z(n1968) );
  OR U2623 ( .A(n1968), .B(n33021), .Z(n1841) );
  NAND U2624 ( .A(n1842), .B(n1841), .Z(n1964) );
  XOR U2625 ( .A(n1965), .B(n1964), .Z(n1927) );
  XOR U2626 ( .A(n1926), .B(n1927), .Z(n1974) );
  NANDN U2627 ( .A(n1844), .B(n1843), .Z(n1848) );
  NAND U2628 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U2629 ( .A(n1848), .B(n1847), .Z(n1975) );
  XNOR U2630 ( .A(n1974), .B(n1975), .Z(n1976) );
  NANDN U2631 ( .A(n1850), .B(n1849), .Z(n1854) );
  NAND U2632 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U2633 ( .A(n1854), .B(n1853), .Z(n1977) );
  XNOR U2634 ( .A(n1976), .B(n1977), .Z(n1919) );
  XNOR U2635 ( .A(n1918), .B(n1919), .Z(n1920) );
  NANDN U2636 ( .A(n1856), .B(n1855), .Z(n1860) );
  NAND U2637 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2638 ( .A(n1860), .B(n1859), .Z(n1985) );
  XOR U2639 ( .A(b[5]), .B(n13976), .Z(n1933) );
  OR U2640 ( .A(n1933), .B(n29363), .Z(n1863) );
  NAND U2641 ( .A(n1861), .B(n29864), .Z(n1862) );
  NAND U2642 ( .A(n1863), .B(n1862), .Z(n1942) );
  XOR U2643 ( .A(b[13]), .B(n11694), .Z(n1954) );
  OR U2644 ( .A(n1954), .B(n31550), .Z(n1866) );
  NANDN U2645 ( .A(n1864), .B(n31874), .Z(n1865) );
  NAND U2646 ( .A(n1866), .B(n1865), .Z(n1939) );
  XOR U2647 ( .A(b[15]), .B(n11202), .Z(n1951) );
  OR U2648 ( .A(n1951), .B(n32010), .Z(n1869) );
  NANDN U2649 ( .A(n1867), .B(n32011), .Z(n1868) );
  AND U2650 ( .A(n1869), .B(n1868), .Z(n1940) );
  XNOR U2651 ( .A(n1939), .B(n1940), .Z(n1941) );
  XNOR U2652 ( .A(n1942), .B(n1941), .Z(n1983) );
  XOR U2653 ( .A(b[11]), .B(n12258), .Z(n1971) );
  OR U2654 ( .A(n1971), .B(n31369), .Z(n1872) );
  NAND U2655 ( .A(n1870), .B(n31119), .Z(n1871) );
  NAND U2656 ( .A(n1872), .B(n1871), .Z(n1963) );
  NANDN U2657 ( .A(n966), .B(a[19]), .Z(n1873) );
  XOR U2658 ( .A(n29232), .B(n1873), .Z(n1875) );
  IV U2659 ( .A(a[18]), .Z(n14905) );
  NANDN U2660 ( .A(n14905), .B(n966), .Z(n1874) );
  AND U2661 ( .A(n1875), .B(n1874), .Z(n1960) );
  XOR U2662 ( .A(n967), .B(n14514), .Z(n1936) );
  NAND U2663 ( .A(n28939), .B(n1936), .Z(n1878) );
  NAND U2664 ( .A(n28938), .B(n1876), .Z(n1877) );
  AND U2665 ( .A(n1878), .B(n1877), .Z(n1961) );
  XNOR U2666 ( .A(n1960), .B(n1961), .Z(n1962) );
  XNOR U2667 ( .A(n1963), .B(n1962), .Z(n1980) );
  XOR U2668 ( .A(b[7]), .B(n13509), .Z(n1930) );
  NANDN U2669 ( .A(n1930), .B(n29949), .Z(n1881) );
  NANDN U2670 ( .A(n1879), .B(n29948), .Z(n1880) );
  NAND U2671 ( .A(n1881), .B(n1880), .Z(n1981) );
  XNOR U2672 ( .A(n1980), .B(n1981), .Z(n1982) );
  XOR U2673 ( .A(n1983), .B(n1982), .Z(n1984) );
  XOR U2674 ( .A(n1985), .B(n1984), .Z(n1987) );
  OR U2675 ( .A(n1883), .B(n1882), .Z(n1887) );
  NANDN U2676 ( .A(n1885), .B(n1884), .Z(n1886) );
  AND U2677 ( .A(n1887), .B(n1886), .Z(n1986) );
  XNOR U2678 ( .A(n1987), .B(n1986), .Z(n1921) );
  XOR U2679 ( .A(n1920), .B(n1921), .Z(n1993) );
  NANDN U2680 ( .A(n1889), .B(n1888), .Z(n1893) );
  NANDN U2681 ( .A(n1891), .B(n1890), .Z(n1892) );
  NAND U2682 ( .A(n1893), .B(n1892), .Z(n1991) );
  XNOR U2683 ( .A(n1991), .B(n1990), .Z(n1992) );
  XNOR U2684 ( .A(n1993), .B(n1992), .Z(n1914) );
  NANDN U2685 ( .A(n1899), .B(n1898), .Z(n1903) );
  NANDN U2686 ( .A(n1901), .B(n1900), .Z(n1902) );
  NAND U2687 ( .A(n1903), .B(n1902), .Z(n1915) );
  XNOR U2688 ( .A(n1914), .B(n1915), .Z(n1916) );
  XNOR U2689 ( .A(n1917), .B(n1916), .Z(n1909) );
  XNOR U2690 ( .A(n1909), .B(sreg[83]), .Z(n1911) );
  NAND U2691 ( .A(n1904), .B(sreg[82]), .Z(n1908) );
  OR U2692 ( .A(n1906), .B(n1905), .Z(n1907) );
  AND U2693 ( .A(n1908), .B(n1907), .Z(n1910) );
  XOR U2694 ( .A(n1911), .B(n1910), .Z(c[83]) );
  NAND U2695 ( .A(n1909), .B(sreg[83]), .Z(n1913) );
  OR U2696 ( .A(n1911), .B(n1910), .Z(n1912) );
  NAND U2697 ( .A(n1913), .B(n1912), .Z(n2091) );
  XNOR U2698 ( .A(n2091), .B(sreg[84]), .Z(n2093) );
  NANDN U2699 ( .A(n1919), .B(n1918), .Z(n1923) );
  NANDN U2700 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U2701 ( .A(n1923), .B(n1922), .Z(n2003) );
  NANDN U2702 ( .A(n1925), .B(n1924), .Z(n1929) );
  NANDN U2703 ( .A(n1927), .B(n1926), .Z(n1928) );
  NAND U2704 ( .A(n1929), .B(n1928), .Z(n2015) );
  XOR U2705 ( .A(b[7]), .B(n14210), .Z(n2056) );
  NANDN U2706 ( .A(n2056), .B(n29949), .Z(n1932) );
  NANDN U2707 ( .A(n1930), .B(n29948), .Z(n1931) );
  AND U2708 ( .A(n1932), .B(n1931), .Z(n2026) );
  XOR U2709 ( .A(n968), .B(n14259), .Z(n2053) );
  NANDN U2710 ( .A(n29363), .B(n2053), .Z(n1935) );
  NANDN U2711 ( .A(n1933), .B(n29864), .Z(n1934) );
  AND U2712 ( .A(n1935), .B(n1934), .Z(n2027) );
  XOR U2713 ( .A(n2026), .B(n2027), .Z(n2028) );
  XOR U2714 ( .A(n967), .B(n14905), .Z(n2088) );
  NAND U2715 ( .A(n2088), .B(n28939), .Z(n1938) );
  NAND U2716 ( .A(n1936), .B(n28938), .Z(n1937) );
  AND U2717 ( .A(n1938), .B(n1937), .Z(n2029) );
  XNOR U2718 ( .A(n2028), .B(n2029), .Z(n2020) );
  NANDN U2719 ( .A(n1940), .B(n1939), .Z(n1944) );
  NAND U2720 ( .A(n1942), .B(n1941), .Z(n1943) );
  NAND U2721 ( .A(n1944), .B(n1943), .Z(n2021) );
  XOR U2722 ( .A(n2020), .B(n2021), .Z(n2022) );
  XOR U2723 ( .A(n33020), .B(b[20]), .Z(n33634) );
  NOR U2724 ( .A(n986), .B(n33634), .Z(n2066) );
  NANDN U2725 ( .A(n966), .B(a[20]), .Z(n1945) );
  XOR U2726 ( .A(n29232), .B(n1945), .Z(n1947) );
  IV U2727 ( .A(a[19]), .Z(n15113) );
  NANDN U2728 ( .A(n15113), .B(n966), .Z(n1946) );
  AND U2729 ( .A(n1947), .B(n1946), .Z(n2064) );
  XNOR U2730 ( .A(b[17]), .B(n10854), .Z(n2050) );
  NAND U2731 ( .A(n2050), .B(n32543), .Z(n1950) );
  NAND U2732 ( .A(n1948), .B(n32541), .Z(n1949) );
  AND U2733 ( .A(n1950), .B(n1949), .Z(n2063) );
  XNOR U2734 ( .A(n2064), .B(n2063), .Z(n2065) );
  XOR U2735 ( .A(n2066), .B(n2065), .Z(n2023) );
  XNOR U2736 ( .A(n2022), .B(n2023), .Z(n2014) );
  XNOR U2737 ( .A(n2015), .B(n2014), .Z(n2017) );
  NANDN U2738 ( .A(n1951), .B(n32011), .Z(n1953) );
  XNOR U2739 ( .A(n972), .B(a[6]), .Z(n2044) );
  NANDN U2740 ( .A(n32010), .B(n2044), .Z(n1952) );
  AND U2741 ( .A(n1953), .B(n1952), .Z(n2032) );
  XOR U2742 ( .A(b[13]), .B(n11986), .Z(n2047) );
  OR U2743 ( .A(n2047), .B(n31550), .Z(n1956) );
  NANDN U2744 ( .A(n1954), .B(n31874), .Z(n1955) );
  AND U2745 ( .A(n1956), .B(n1955), .Z(n2033) );
  XOR U2746 ( .A(n2032), .B(n2033), .Z(n2034) );
  XOR U2747 ( .A(b[9]), .B(n13106), .Z(n2082) );
  NANDN U2748 ( .A(n2082), .B(n30509), .Z(n1959) );
  NAND U2749 ( .A(n1957), .B(n30846), .Z(n1958) );
  AND U2750 ( .A(n1959), .B(n1958), .Z(n2035) );
  XNOR U2751 ( .A(n2034), .B(n2035), .Z(n2038) );
  XOR U2752 ( .A(n2038), .B(n2039), .Z(n2040) );
  NAND U2753 ( .A(n1965), .B(n1964), .Z(n2061) );
  AND U2754 ( .A(n1967), .B(n1966), .Z(n33283) );
  NANDN U2755 ( .A(n1968), .B(n33283), .Z(n1970) );
  XNOR U2756 ( .A(n33020), .B(a[2]), .Z(n2069) );
  NANDN U2757 ( .A(n33021), .B(n2069), .Z(n1969) );
  NAND U2758 ( .A(n1970), .B(n1969), .Z(n2060) );
  XOR U2759 ( .A(b[11]), .B(n12555), .Z(n2079) );
  OR U2760 ( .A(n2079), .B(n31369), .Z(n1973) );
  NANDN U2761 ( .A(n1971), .B(n31119), .Z(n1972) );
  AND U2762 ( .A(n1973), .B(n1972), .Z(n2059) );
  XNOR U2763 ( .A(n2060), .B(n2059), .Z(n2062) );
  XNOR U2764 ( .A(n2061), .B(n2062), .Z(n2041) );
  XNOR U2765 ( .A(n2040), .B(n2041), .Z(n2016) );
  XOR U2766 ( .A(n2017), .B(n2016), .Z(n2011) );
  NANDN U2767 ( .A(n1975), .B(n1974), .Z(n1979) );
  NANDN U2768 ( .A(n1977), .B(n1976), .Z(n1978) );
  NAND U2769 ( .A(n1979), .B(n1978), .Z(n2008) );
  XNOR U2770 ( .A(n2008), .B(n2009), .Z(n2010) );
  XOR U2771 ( .A(n2011), .B(n2010), .Z(n2002) );
  XOR U2772 ( .A(n2003), .B(n2002), .Z(n2005) );
  NANDN U2773 ( .A(n1985), .B(n1984), .Z(n1989) );
  OR U2774 ( .A(n1987), .B(n1986), .Z(n1988) );
  NAND U2775 ( .A(n1989), .B(n1988), .Z(n2004) );
  XNOR U2776 ( .A(n2005), .B(n2004), .Z(n1996) );
  NANDN U2777 ( .A(n1991), .B(n1990), .Z(n1995) );
  NAND U2778 ( .A(n1993), .B(n1992), .Z(n1994) );
  NAND U2779 ( .A(n1995), .B(n1994), .Z(n1997) );
  XNOR U2780 ( .A(n1996), .B(n1997), .Z(n1998) );
  XOR U2781 ( .A(n1999), .B(n1998), .Z(n2092) );
  XOR U2782 ( .A(n2093), .B(n2092), .Z(c[84]) );
  NANDN U2783 ( .A(n1997), .B(n1996), .Z(n2001) );
  NAND U2784 ( .A(n1999), .B(n1998), .Z(n2000) );
  NAND U2785 ( .A(n2001), .B(n2000), .Z(n2104) );
  NANDN U2786 ( .A(n2003), .B(n2002), .Z(n2007) );
  OR U2787 ( .A(n2005), .B(n2004), .Z(n2006) );
  NAND U2788 ( .A(n2007), .B(n2006), .Z(n2102) );
  NANDN U2789 ( .A(n2009), .B(n2008), .Z(n2013) );
  NAND U2790 ( .A(n2011), .B(n2010), .Z(n2012) );
  NAND U2791 ( .A(n2013), .B(n2012), .Z(n2107) );
  NAND U2792 ( .A(n2015), .B(n2014), .Z(n2019) );
  NANDN U2793 ( .A(n2017), .B(n2016), .Z(n2018) );
  NAND U2794 ( .A(n2019), .B(n2018), .Z(n2106) );
  OR U2795 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U2796 ( .A(n2023), .B(n2022), .Z(n2024) );
  NAND U2797 ( .A(n2025), .B(n2024), .Z(n2112) );
  OR U2798 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U2799 ( .A(n2029), .B(n2028), .Z(n2030) );
  AND U2800 ( .A(n2031), .B(n2030), .Z(n2109) );
  OR U2801 ( .A(n2033), .B(n2032), .Z(n2037) );
  NANDN U2802 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U2803 ( .A(n2037), .B(n2036), .Z(n2110) );
  XOR U2804 ( .A(n2109), .B(n2110), .Z(n2111) );
  XNOR U2805 ( .A(n2112), .B(n2111), .Z(n2118) );
  OR U2806 ( .A(n2039), .B(n2038), .Z(n2043) );
  NANDN U2807 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2808 ( .A(n2043), .B(n2042), .Z(n2115) );
  XOR U2809 ( .A(b[15]), .B(n11694), .Z(n2139) );
  OR U2810 ( .A(n2139), .B(n32010), .Z(n2046) );
  NAND U2811 ( .A(n2044), .B(n32011), .Z(n2045) );
  NAND U2812 ( .A(n2046), .B(n2045), .Z(n2164) );
  XOR U2813 ( .A(n971), .B(n12258), .Z(n2188) );
  NANDN U2814 ( .A(n31550), .B(n2188), .Z(n2049) );
  NANDN U2815 ( .A(n2047), .B(n31874), .Z(n2048) );
  AND U2816 ( .A(n2049), .B(n2048), .Z(n2162) );
  XNOR U2817 ( .A(b[17]), .B(a[5]), .Z(n2151) );
  NANDN U2818 ( .A(n2151), .B(n32543), .Z(n2052) );
  NAND U2819 ( .A(n2050), .B(n32541), .Z(n2051) );
  AND U2820 ( .A(n2052), .B(n2051), .Z(n2163) );
  XOR U2821 ( .A(n2164), .B(n2165), .Z(n2136) );
  NAND U2822 ( .A(n29864), .B(n2053), .Z(n2055) );
  XNOR U2823 ( .A(n968), .B(a[17]), .Z(n2145) );
  NANDN U2824 ( .A(n29363), .B(n2145), .Z(n2054) );
  NAND U2825 ( .A(n2055), .B(n2054), .Z(n2134) );
  XNOR U2826 ( .A(n31123), .B(a[15]), .Z(n2142) );
  NAND U2827 ( .A(n2142), .B(n29949), .Z(n2058) );
  NANDN U2828 ( .A(n2056), .B(n29948), .Z(n2057) );
  AND U2829 ( .A(n2058), .B(n2057), .Z(n2133) );
  XNOR U2830 ( .A(n2134), .B(n2133), .Z(n2135) );
  XOR U2831 ( .A(n2136), .B(n2135), .Z(n2127) );
  XOR U2832 ( .A(n2127), .B(n2128), .Z(n2129) );
  NANDN U2833 ( .A(n2064), .B(n2063), .Z(n2068) );
  NANDN U2834 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U2835 ( .A(n2068), .B(n2067), .Z(n2124) );
  NAND U2836 ( .A(n2069), .B(n33283), .Z(n2071) );
  XNOR U2837 ( .A(n33020), .B(a[3]), .Z(n2177) );
  NANDN U2838 ( .A(n33021), .B(n2177), .Z(n2070) );
  NAND U2839 ( .A(n2071), .B(n2070), .Z(n2187) );
  XOR U2840 ( .A(n986), .B(b[19]), .Z(n2072) );
  NAND U2841 ( .A(n2072), .B(n33634), .Z(n2074) );
  XNOR U2842 ( .A(b[21]), .B(b[20]), .Z(n2073) );
  OR U2843 ( .A(n2074), .B(n2073), .Z(n2076) );
  XNOR U2844 ( .A(b[21]), .B(a[1]), .Z(n2156) );
  OR U2845 ( .A(n2156), .B(n33634), .Z(n2075) );
  NAND U2846 ( .A(n2076), .B(n2075), .Z(n2186) );
  XOR U2847 ( .A(n2187), .B(n2186), .Z(n2182) );
  NANDN U2848 ( .A(n33020), .B(b[20]), .Z(n33632) );
  NAND U2849 ( .A(n33632), .B(b[21]), .Z(n33984) );
  NOR U2850 ( .A(b[19]), .B(b[20]), .Z(n2077) );
  OR U2851 ( .A(n2077), .B(n986), .Z(n2078) );
  NANDN U2852 ( .A(n33984), .B(n2078), .Z(n2180) );
  XOR U2853 ( .A(b[11]), .B(n12830), .Z(n2159) );
  OR U2854 ( .A(n2159), .B(n31369), .Z(n2081) );
  NANDN U2855 ( .A(n2079), .B(n31119), .Z(n2080) );
  NAND U2856 ( .A(n2081), .B(n2080), .Z(n2181) );
  XOR U2857 ( .A(n2180), .B(n2181), .Z(n2183) );
  XNOR U2858 ( .A(n2182), .B(n2183), .Z(n2121) );
  XOR U2859 ( .A(b[9]), .B(n13509), .Z(n2148) );
  NANDN U2860 ( .A(n2148), .B(n30509), .Z(n2084) );
  NANDN U2861 ( .A(n2082), .B(n30846), .Z(n2083) );
  NAND U2862 ( .A(n2084), .B(n2083), .Z(n2171) );
  NANDN U2863 ( .A(n966), .B(a[21]), .Z(n2085) );
  XOR U2864 ( .A(n29232), .B(n2085), .Z(n2087) );
  IV U2865 ( .A(a[20]), .Z(n15484) );
  NANDN U2866 ( .A(n15484), .B(n966), .Z(n2086) );
  AND U2867 ( .A(n2087), .B(n2086), .Z(n2168) );
  XOR U2868 ( .A(b[3]), .B(n15113), .Z(n2191) );
  NANDN U2869 ( .A(n2191), .B(n28939), .Z(n2090) );
  NAND U2870 ( .A(n28938), .B(n2088), .Z(n2089) );
  AND U2871 ( .A(n2090), .B(n2089), .Z(n2169) );
  XNOR U2872 ( .A(n2168), .B(n2169), .Z(n2170) );
  XNOR U2873 ( .A(n2171), .B(n2170), .Z(n2122) );
  XOR U2874 ( .A(n2121), .B(n2122), .Z(n2123) );
  XNOR U2875 ( .A(n2124), .B(n2123), .Z(n2130) );
  XNOR U2876 ( .A(n2129), .B(n2130), .Z(n2116) );
  XNOR U2877 ( .A(n2115), .B(n2116), .Z(n2117) );
  XNOR U2878 ( .A(n2118), .B(n2117), .Z(n2105) );
  XNOR U2879 ( .A(n2106), .B(n2105), .Z(n2108) );
  XOR U2880 ( .A(n2107), .B(n2108), .Z(n2101) );
  XNOR U2881 ( .A(n2102), .B(n2101), .Z(n2103) );
  XNOR U2882 ( .A(n2104), .B(n2103), .Z(n2096) );
  XNOR U2883 ( .A(n2096), .B(sreg[85]), .Z(n2098) );
  NAND U2884 ( .A(n2091), .B(sreg[84]), .Z(n2095) );
  OR U2885 ( .A(n2093), .B(n2092), .Z(n2094) );
  AND U2886 ( .A(n2095), .B(n2094), .Z(n2097) );
  XOR U2887 ( .A(n2098), .B(n2097), .Z(c[85]) );
  NAND U2888 ( .A(n2096), .B(sreg[85]), .Z(n2100) );
  OR U2889 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2890 ( .A(n2100), .B(n2099), .Z(n2296) );
  XNOR U2891 ( .A(n2296), .B(sreg[86]), .Z(n2298) );
  OR U2892 ( .A(n2110), .B(n2109), .Z(n2114) );
  NANDN U2893 ( .A(n2112), .B(n2111), .Z(n2113) );
  NAND U2894 ( .A(n2114), .B(n2113), .Z(n2203) );
  NANDN U2895 ( .A(n2116), .B(n2115), .Z(n2120) );
  NANDN U2896 ( .A(n2118), .B(n2117), .Z(n2119) );
  NAND U2897 ( .A(n2120), .B(n2119), .Z(n2201) );
  NANDN U2898 ( .A(n2122), .B(n2121), .Z(n2126) );
  OR U2899 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U2900 ( .A(n2126), .B(n2125), .Z(n2208) );
  OR U2901 ( .A(n2128), .B(n2127), .Z(n2132) );
  NANDN U2902 ( .A(n2130), .B(n2129), .Z(n2131) );
  NAND U2903 ( .A(n2132), .B(n2131), .Z(n2207) );
  NANDN U2904 ( .A(n2134), .B(n2133), .Z(n2138) );
  NAND U2905 ( .A(n2136), .B(n2135), .Z(n2137) );
  NAND U2906 ( .A(n2138), .B(n2137), .Z(n2285) );
  XOR U2907 ( .A(b[15]), .B(n11986), .Z(n2218) );
  OR U2908 ( .A(n2218), .B(n32010), .Z(n2141) );
  NANDN U2909 ( .A(n2139), .B(n32011), .Z(n2140) );
  NAND U2910 ( .A(n2141), .B(n2140), .Z(n2275) );
  XOR U2911 ( .A(n31123), .B(n14259), .Z(n2253) );
  NAND U2912 ( .A(n2253), .B(n29949), .Z(n2144) );
  NAND U2913 ( .A(n2142), .B(n29948), .Z(n2143) );
  NAND U2914 ( .A(n2144), .B(n2143), .Z(n2272) );
  XOR U2915 ( .A(b[5]), .B(n14905), .Z(n2259) );
  OR U2916 ( .A(n2259), .B(n29363), .Z(n2147) );
  NAND U2917 ( .A(n2145), .B(n29864), .Z(n2146) );
  AND U2918 ( .A(n2147), .B(n2146), .Z(n2273) );
  XNOR U2919 ( .A(n2272), .B(n2273), .Z(n2274) );
  XNOR U2920 ( .A(n2275), .B(n2274), .Z(n2239) );
  XOR U2921 ( .A(b[9]), .B(n14210), .Z(n2256) );
  NANDN U2922 ( .A(n2256), .B(n30509), .Z(n2150) );
  NANDN U2923 ( .A(n2148), .B(n30846), .Z(n2149) );
  NAND U2924 ( .A(n2150), .B(n2149), .Z(n2269) );
  XNOR U2925 ( .A(b[17]), .B(a[6]), .Z(n2221) );
  NANDN U2926 ( .A(n2221), .B(n32543), .Z(n2153) );
  NANDN U2927 ( .A(n2151), .B(n32541), .Z(n2152) );
  NAND U2928 ( .A(n2153), .B(n2152), .Z(n2266) );
  XNOR U2929 ( .A(b[21]), .B(a[2]), .Z(n2240) );
  OR U2930 ( .A(n2240), .B(n33634), .Z(n2158) );
  XNOR U2931 ( .A(b[21]), .B(n33020), .Z(n2155) );
  XOR U2932 ( .A(b[21]), .B(b[20]), .Z(n2154) );
  AND U2933 ( .A(n2155), .B(n2154), .Z(n33464) );
  NANDN U2934 ( .A(n2156), .B(n33464), .Z(n2157) );
  AND U2935 ( .A(n2158), .B(n2157), .Z(n2267) );
  XNOR U2936 ( .A(n2266), .B(n2267), .Z(n2268) );
  XNOR U2937 ( .A(n2269), .B(n2268), .Z(n2236) );
  XOR U2938 ( .A(b[11]), .B(n13106), .Z(n2250) );
  OR U2939 ( .A(n2250), .B(n31369), .Z(n2161) );
  NANDN U2940 ( .A(n2159), .B(n31119), .Z(n2160) );
  NAND U2941 ( .A(n2161), .B(n2160), .Z(n2237) );
  XNOR U2942 ( .A(n2236), .B(n2237), .Z(n2238) );
  XOR U2943 ( .A(n2239), .B(n2238), .Z(n2290) );
  OR U2944 ( .A(n2163), .B(n2162), .Z(n2167) );
  NANDN U2945 ( .A(n2165), .B(n2164), .Z(n2166) );
  NAND U2946 ( .A(n2167), .B(n2166), .Z(n2291) );
  XOR U2947 ( .A(n2290), .B(n2291), .Z(n2293) );
  NANDN U2948 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2949 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2950 ( .A(n2173), .B(n2172), .Z(n2292) );
  XOR U2951 ( .A(n2293), .B(n2292), .Z(n2284) );
  XNOR U2952 ( .A(n2285), .B(n2284), .Z(n2287) );
  XNOR U2953 ( .A(b[21]), .B(b[22]), .Z(n33867) );
  NANDN U2954 ( .A(n33867), .B(a[0]), .Z(n2233) );
  NANDN U2955 ( .A(n966), .B(a[22]), .Z(n2174) );
  XOR U2956 ( .A(n29232), .B(n2174), .Z(n2176) );
  IV U2957 ( .A(a[21]), .Z(n16220) );
  NANDN U2958 ( .A(n16220), .B(n966), .Z(n2175) );
  AND U2959 ( .A(n2176), .B(n2175), .Z(n2231) );
  NAND U2960 ( .A(n2177), .B(n33283), .Z(n2179) );
  XNOR U2961 ( .A(n33020), .B(a[4]), .Z(n2224) );
  NANDN U2962 ( .A(n33021), .B(n2224), .Z(n2178) );
  AND U2963 ( .A(n2179), .B(n2178), .Z(n2230) );
  XNOR U2964 ( .A(n2231), .B(n2230), .Z(n2232) );
  XNOR U2965 ( .A(n2233), .B(n2232), .Z(n2281) );
  NANDN U2966 ( .A(n2181), .B(n2180), .Z(n2185) );
  OR U2967 ( .A(n2183), .B(n2182), .Z(n2184) );
  AND U2968 ( .A(n2185), .B(n2184), .Z(n2278) );
  NAND U2969 ( .A(n2187), .B(n2186), .Z(n2264) );
  NAND U2970 ( .A(n31874), .B(n2188), .Z(n2190) );
  XNOR U2971 ( .A(n971), .B(a[10]), .Z(n2227) );
  NANDN U2972 ( .A(n31550), .B(n2227), .Z(n2189) );
  NAND U2973 ( .A(n2190), .B(n2189), .Z(n2263) );
  XOR U2974 ( .A(b[3]), .B(n15484), .Z(n2215) );
  NANDN U2975 ( .A(n2215), .B(n28939), .Z(n2193) );
  NANDN U2976 ( .A(n2191), .B(n28938), .Z(n2192) );
  AND U2977 ( .A(n2193), .B(n2192), .Z(n2262) );
  XNOR U2978 ( .A(n2263), .B(n2262), .Z(n2265) );
  XNOR U2979 ( .A(n2264), .B(n2265), .Z(n2279) );
  XNOR U2980 ( .A(n2278), .B(n2279), .Z(n2280) );
  XNOR U2981 ( .A(n2281), .B(n2280), .Z(n2286) );
  XOR U2982 ( .A(n2287), .B(n2286), .Z(n2206) );
  XOR U2983 ( .A(n2207), .B(n2206), .Z(n2209) );
  XOR U2984 ( .A(n2208), .B(n2209), .Z(n2200) );
  XOR U2985 ( .A(n2201), .B(n2200), .Z(n2202) );
  XOR U2986 ( .A(n2203), .B(n2202), .Z(n2195) );
  XNOR U2987 ( .A(n2194), .B(n2195), .Z(n2196) );
  XOR U2988 ( .A(n2197), .B(n2196), .Z(n2297) );
  XOR U2989 ( .A(n2298), .B(n2297), .Z(c[86]) );
  NANDN U2990 ( .A(n2195), .B(n2194), .Z(n2199) );
  NAND U2991 ( .A(n2197), .B(n2196), .Z(n2198) );
  NAND U2992 ( .A(n2199), .B(n2198), .Z(n2309) );
  NAND U2993 ( .A(n2201), .B(n2200), .Z(n2205) );
  NANDN U2994 ( .A(n2203), .B(n2202), .Z(n2204) );
  NAND U2995 ( .A(n2205), .B(n2204), .Z(n2306) );
  NANDN U2996 ( .A(n2207), .B(n2206), .Z(n2211) );
  OR U2997 ( .A(n2209), .B(n2208), .Z(n2210) );
  NAND U2998 ( .A(n2211), .B(n2210), .Z(n2409) );
  IV U2999 ( .A(b[23]), .Z(n34510) );
  OR U3000 ( .A(b[21]), .B(n34510), .Z(n2212) );
  OR U3001 ( .A(b[22]), .B(n2212), .Z(n2214) );
  ANDN U3002 ( .B(b[23]), .A(n33867), .Z(n34046) );
  NANDN U3003 ( .A(a[0]), .B(n34046), .Z(n2213) );
  NAND U3004 ( .A(n2214), .B(n2213), .Z(n2371) );
  XOR U3005 ( .A(b[3]), .B(n16220), .Z(n2332) );
  NANDN U3006 ( .A(n2332), .B(n28939), .Z(n2217) );
  NANDN U3007 ( .A(n2215), .B(n28938), .Z(n2216) );
  AND U3008 ( .A(n2217), .B(n2216), .Z(n2370) );
  XNOR U3009 ( .A(n2371), .B(n2370), .Z(n2372) );
  NANDN U3010 ( .A(n2218), .B(n32011), .Z(n2220) );
  XOR U3011 ( .A(b[15]), .B(n12258), .Z(n2364) );
  OR U3012 ( .A(n2364), .B(n32010), .Z(n2219) );
  NAND U3013 ( .A(n2220), .B(n2219), .Z(n2373) );
  XOR U3014 ( .A(n2372), .B(n2373), .Z(n2312) );
  XNOR U3015 ( .A(b[17]), .B(a[7]), .Z(n2350) );
  NANDN U3016 ( .A(n2350), .B(n32543), .Z(n2223) );
  NANDN U3017 ( .A(n2221), .B(n32541), .Z(n2222) );
  NAND U3018 ( .A(n2223), .B(n2222), .Z(n2327) );
  NAND U3019 ( .A(n2224), .B(n33283), .Z(n2226) );
  XOR U3020 ( .A(b[19]), .B(n11202), .Z(n2356) );
  OR U3021 ( .A(n2356), .B(n33021), .Z(n2225) );
  NAND U3022 ( .A(n2226), .B(n2225), .Z(n2324) );
  XOR U3023 ( .A(n971), .B(n12830), .Z(n2335) );
  NANDN U3024 ( .A(n31550), .B(n2335), .Z(n2229) );
  NAND U3025 ( .A(n2227), .B(n31874), .Z(n2228) );
  AND U3026 ( .A(n2229), .B(n2228), .Z(n2325) );
  XNOR U3027 ( .A(n2324), .B(n2325), .Z(n2326) );
  XNOR U3028 ( .A(n2327), .B(n2326), .Z(n2313) );
  XNOR U3029 ( .A(n2312), .B(n2313), .Z(n2314) );
  NANDN U3030 ( .A(n2231), .B(n2230), .Z(n2235) );
  NAND U3031 ( .A(n2233), .B(n2232), .Z(n2234) );
  NAND U3032 ( .A(n2235), .B(n2234), .Z(n2315) );
  XOR U3033 ( .A(n2314), .B(n2315), .Z(n2394) );
  XNOR U3034 ( .A(n2394), .B(n2395), .Z(n2396) );
  XNOR U3035 ( .A(b[21]), .B(a[3]), .Z(n2341) );
  OR U3036 ( .A(n2341), .B(n33634), .Z(n2242) );
  NANDN U3037 ( .A(n2240), .B(n33464), .Z(n2241) );
  NAND U3038 ( .A(n2242), .B(n2241), .Z(n2331) );
  XNOR U3039 ( .A(n34510), .B(b[21]), .Z(n2359) );
  XNOR U3040 ( .A(n34510), .B(a[0]), .Z(n2243) );
  NAND U3041 ( .A(n2359), .B(n2243), .Z(n2244) );
  XNOR U3042 ( .A(n34510), .B(b[22]), .Z(n2360) );
  NANDN U3043 ( .A(n2244), .B(n2360), .Z(n2246) );
  XOR U3044 ( .A(n34510), .B(n10457), .Z(n2361) );
  NANDN U3045 ( .A(n33867), .B(n2361), .Z(n2245) );
  NAND U3046 ( .A(n2246), .B(n2245), .Z(n2330) );
  XNOR U3047 ( .A(n2331), .B(n2330), .Z(n2321) );
  NANDN U3048 ( .A(n966), .B(a[23]), .Z(n2247) );
  XOR U3049 ( .A(n29232), .B(n2247), .Z(n2249) );
  IV U3050 ( .A(a[22]), .Z(n15963) );
  NANDN U3051 ( .A(n15963), .B(n966), .Z(n2248) );
  AND U3052 ( .A(n2249), .B(n2248), .Z(n2319) );
  XOR U3053 ( .A(b[11]), .B(n13509), .Z(n2367) );
  OR U3054 ( .A(n2367), .B(n31369), .Z(n2252) );
  NANDN U3055 ( .A(n2250), .B(n31119), .Z(n2251) );
  AND U3056 ( .A(n2252), .B(n2251), .Z(n2318) );
  XNOR U3057 ( .A(n2319), .B(n2318), .Z(n2320) );
  XOR U3058 ( .A(n2321), .B(n2320), .Z(n2388) );
  XOR U3059 ( .A(n31123), .B(n14514), .Z(n2344) );
  NAND U3060 ( .A(n2344), .B(n29949), .Z(n2255) );
  NAND U3061 ( .A(n29948), .B(n2253), .Z(n2254) );
  NAND U3062 ( .A(n2255), .B(n2254), .Z(n2379) );
  XOR U3063 ( .A(n969), .B(n13976), .Z(n2353) );
  NAND U3064 ( .A(n30509), .B(n2353), .Z(n2258) );
  NANDN U3065 ( .A(n2256), .B(n30846), .Z(n2257) );
  NAND U3066 ( .A(n2258), .B(n2257), .Z(n2376) );
  XOR U3067 ( .A(b[5]), .B(n15113), .Z(n2347) );
  OR U3068 ( .A(n2347), .B(n29363), .Z(n2261) );
  NANDN U3069 ( .A(n2259), .B(n29864), .Z(n2260) );
  AND U3070 ( .A(n2261), .B(n2260), .Z(n2377) );
  XNOR U3071 ( .A(n2376), .B(n2377), .Z(n2378) );
  XNOR U3072 ( .A(n2379), .B(n2378), .Z(n2389) );
  XNOR U3073 ( .A(n2388), .B(n2389), .Z(n2391) );
  XNOR U3074 ( .A(n2391), .B(n2390), .Z(n2385) );
  NANDN U3075 ( .A(n2267), .B(n2266), .Z(n2271) );
  NAND U3076 ( .A(n2269), .B(n2268), .Z(n2270) );
  NAND U3077 ( .A(n2271), .B(n2270), .Z(n2383) );
  NANDN U3078 ( .A(n2273), .B(n2272), .Z(n2277) );
  NAND U3079 ( .A(n2275), .B(n2274), .Z(n2276) );
  AND U3080 ( .A(n2277), .B(n2276), .Z(n2382) );
  XNOR U3081 ( .A(n2383), .B(n2382), .Z(n2384) );
  XOR U3082 ( .A(n2385), .B(n2384), .Z(n2397) );
  XOR U3083 ( .A(n2396), .B(n2397), .Z(n2406) );
  OR U3084 ( .A(n2279), .B(n2278), .Z(n2283) );
  OR U3085 ( .A(n2281), .B(n2280), .Z(n2282) );
  NAND U3086 ( .A(n2283), .B(n2282), .Z(n2403) );
  NAND U3087 ( .A(n2285), .B(n2284), .Z(n2289) );
  OR U3088 ( .A(n2287), .B(n2286), .Z(n2288) );
  NAND U3089 ( .A(n2289), .B(n2288), .Z(n2400) );
  NANDN U3090 ( .A(n2291), .B(n2290), .Z(n2295) );
  OR U3091 ( .A(n2293), .B(n2292), .Z(n2294) );
  AND U3092 ( .A(n2295), .B(n2294), .Z(n2401) );
  XNOR U3093 ( .A(n2400), .B(n2401), .Z(n2402) );
  XOR U3094 ( .A(n2403), .B(n2402), .Z(n2407) );
  XOR U3095 ( .A(n2406), .B(n2407), .Z(n2408) );
  XNOR U3096 ( .A(n2409), .B(n2408), .Z(n2307) );
  XNOR U3097 ( .A(n2306), .B(n2307), .Z(n2308) );
  XNOR U3098 ( .A(n2309), .B(n2308), .Z(n2301) );
  XNOR U3099 ( .A(n2301), .B(sreg[87]), .Z(n2303) );
  NAND U3100 ( .A(n2296), .B(sreg[86]), .Z(n2300) );
  OR U3101 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U3102 ( .A(n2300), .B(n2299), .Z(n2302) );
  XOR U3103 ( .A(n2303), .B(n2302), .Z(c[87]) );
  NAND U3104 ( .A(n2301), .B(sreg[87]), .Z(n2305) );
  OR U3105 ( .A(n2303), .B(n2302), .Z(n2304) );
  NAND U3106 ( .A(n2305), .B(n2304), .Z(n2524) );
  XNOR U3107 ( .A(n2524), .B(sreg[88]), .Z(n2526) );
  NANDN U3108 ( .A(n2307), .B(n2306), .Z(n2311) );
  NAND U3109 ( .A(n2309), .B(n2308), .Z(n2310) );
  NAND U3110 ( .A(n2311), .B(n2310), .Z(n2415) );
  NANDN U3111 ( .A(n2313), .B(n2312), .Z(n2317) );
  NANDN U3112 ( .A(n2315), .B(n2314), .Z(n2316) );
  NAND U3113 ( .A(n2317), .B(n2316), .Z(n2427) );
  NANDN U3114 ( .A(n2319), .B(n2318), .Z(n2323) );
  NAND U3115 ( .A(n2321), .B(n2320), .Z(n2322) );
  NAND U3116 ( .A(n2323), .B(n2322), .Z(n2512) );
  NANDN U3117 ( .A(n2325), .B(n2324), .Z(n2329) );
  NAND U3118 ( .A(n2327), .B(n2326), .Z(n2328) );
  NAND U3119 ( .A(n2329), .B(n2328), .Z(n2513) );
  XNOR U3120 ( .A(n2512), .B(n2513), .Z(n2514) );
  NAND U3121 ( .A(n2331), .B(n2330), .Z(n2439) );
  XOR U3122 ( .A(b[3]), .B(n15963), .Z(n2454) );
  NANDN U3123 ( .A(n2454), .B(n28939), .Z(n2334) );
  NANDN U3124 ( .A(n2332), .B(n28938), .Z(n2333) );
  NAND U3125 ( .A(n2334), .B(n2333), .Z(n2437) );
  NAND U3126 ( .A(n31874), .B(n2335), .Z(n2337) );
  XOR U3127 ( .A(n971), .B(n13106), .Z(n2470) );
  NANDN U3128 ( .A(n31550), .B(n2470), .Z(n2336) );
  AND U3129 ( .A(n2337), .B(n2336), .Z(n2436) );
  XNOR U3130 ( .A(n2437), .B(n2436), .Z(n2438) );
  XNOR U3131 ( .A(n2439), .B(n2438), .Z(n2515) );
  XNOR U3132 ( .A(n2514), .B(n2515), .Z(n2430) );
  XNOR U3133 ( .A(b[24]), .B(b[23]), .Z(n34219) );
  NANDN U3134 ( .A(n34219), .B(a[0]), .Z(n2449) );
  NANDN U3135 ( .A(n966), .B(a[24]), .Z(n2338) );
  XOR U3136 ( .A(n29232), .B(n2338), .Z(n2340) );
  IV U3137 ( .A(a[23]), .Z(n16269) );
  NANDN U3138 ( .A(n16269), .B(n966), .Z(n2339) );
  AND U3139 ( .A(n2340), .B(n2339), .Z(n2447) );
  XNOR U3140 ( .A(b[21]), .B(n10854), .Z(n2497) );
  NANDN U3141 ( .A(n33634), .B(n2497), .Z(n2343) );
  NANDN U3142 ( .A(n2341), .B(n33464), .Z(n2342) );
  AND U3143 ( .A(n2343), .B(n2342), .Z(n2446) );
  XNOR U3144 ( .A(n2447), .B(n2446), .Z(n2448) );
  XOR U3145 ( .A(n2449), .B(n2448), .Z(n2473) );
  XOR U3146 ( .A(n31123), .B(n14905), .Z(n2485) );
  NAND U3147 ( .A(n2485), .B(n29949), .Z(n2346) );
  NAND U3148 ( .A(n29948), .B(n2344), .Z(n2345) );
  NAND U3149 ( .A(n2346), .B(n2345), .Z(n2482) );
  XOR U3150 ( .A(b[5]), .B(n15484), .Z(n2488) );
  OR U3151 ( .A(n2488), .B(n29363), .Z(n2349) );
  NANDN U3152 ( .A(n2347), .B(n29864), .Z(n2348) );
  NAND U3153 ( .A(n2349), .B(n2348), .Z(n2479) );
  XNOR U3154 ( .A(b[17]), .B(a[8]), .Z(n2491) );
  NANDN U3155 ( .A(n2491), .B(n32543), .Z(n2352) );
  NANDN U3156 ( .A(n2350), .B(n32541), .Z(n2351) );
  AND U3157 ( .A(n2352), .B(n2351), .Z(n2480) );
  XNOR U3158 ( .A(n2479), .B(n2480), .Z(n2481) );
  XNOR U3159 ( .A(n2482), .B(n2481), .Z(n2474) );
  XNOR U3160 ( .A(n2473), .B(n2474), .Z(n2476) );
  NAND U3161 ( .A(n30846), .B(n2353), .Z(n2355) );
  XNOR U3162 ( .A(n969), .B(a[16]), .Z(n2500) );
  NAND U3163 ( .A(n30509), .B(n2500), .Z(n2354) );
  NAND U3164 ( .A(n2355), .B(n2354), .Z(n2444) );
  NANDN U3165 ( .A(n2356), .B(n33283), .Z(n2358) );
  XNOR U3166 ( .A(n33020), .B(a[6]), .Z(n2494) );
  NANDN U3167 ( .A(n33021), .B(n2494), .Z(n2357) );
  NAND U3168 ( .A(n2358), .B(n2357), .Z(n2442) );
  AND U3169 ( .A(n2360), .B(n2359), .Z(n34044) );
  NAND U3170 ( .A(n2361), .B(n34044), .Z(n2363) );
  XNOR U3171 ( .A(n34510), .B(a[2]), .Z(n2460) );
  NANDN U3172 ( .A(n33867), .B(n2460), .Z(n2362) );
  NAND U3173 ( .A(n2363), .B(n2362), .Z(n2443) );
  XNOR U3174 ( .A(n2442), .B(n2443), .Z(n2445) );
  XOR U3175 ( .A(n2444), .B(n2445), .Z(n2509) );
  NANDN U3176 ( .A(n2364), .B(n32011), .Z(n2366) );
  XOR U3177 ( .A(b[15]), .B(n12555), .Z(n2457) );
  OR U3178 ( .A(n2457), .B(n32010), .Z(n2365) );
  NAND U3179 ( .A(n2366), .B(n2365), .Z(n2507) );
  XOR U3180 ( .A(b[11]), .B(n14210), .Z(n2503) );
  OR U3181 ( .A(n2503), .B(n31369), .Z(n2369) );
  NANDN U3182 ( .A(n2367), .B(n31119), .Z(n2368) );
  AND U3183 ( .A(n2369), .B(n2368), .Z(n2506) );
  XNOR U3184 ( .A(n2507), .B(n2506), .Z(n2508) );
  XOR U3185 ( .A(n2509), .B(n2508), .Z(n2475) );
  XNOR U3186 ( .A(n2476), .B(n2475), .Z(n2521) );
  NANDN U3187 ( .A(n2371), .B(n2370), .Z(n2375) );
  NANDN U3188 ( .A(n2373), .B(n2372), .Z(n2374) );
  NAND U3189 ( .A(n2375), .B(n2374), .Z(n2518) );
  NANDN U3190 ( .A(n2377), .B(n2376), .Z(n2381) );
  NAND U3191 ( .A(n2379), .B(n2378), .Z(n2380) );
  NAND U3192 ( .A(n2381), .B(n2380), .Z(n2519) );
  XNOR U3193 ( .A(n2518), .B(n2519), .Z(n2520) );
  XOR U3194 ( .A(n2521), .B(n2520), .Z(n2431) );
  NANDN U3195 ( .A(n2383), .B(n2382), .Z(n2387) );
  NAND U3196 ( .A(n2385), .B(n2384), .Z(n2386) );
  NAND U3197 ( .A(n2387), .B(n2386), .Z(n2433) );
  XOR U3198 ( .A(n2432), .B(n2433), .Z(n2424) );
  OR U3199 ( .A(n2389), .B(n2388), .Z(n2393) );
  OR U3200 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U3201 ( .A(n2393), .B(n2392), .Z(n2425) );
  XNOR U3202 ( .A(n2424), .B(n2425), .Z(n2426) );
  XOR U3203 ( .A(n2427), .B(n2426), .Z(n2418) );
  NANDN U3204 ( .A(n2395), .B(n2394), .Z(n2399) );
  NAND U3205 ( .A(n2397), .B(n2396), .Z(n2398) );
  NAND U3206 ( .A(n2399), .B(n2398), .Z(n2419) );
  XNOR U3207 ( .A(n2418), .B(n2419), .Z(n2420) );
  NANDN U3208 ( .A(n2401), .B(n2400), .Z(n2405) );
  NAND U3209 ( .A(n2403), .B(n2402), .Z(n2404) );
  NAND U3210 ( .A(n2405), .B(n2404), .Z(n2421) );
  XOR U3211 ( .A(n2420), .B(n2421), .Z(n2412) );
  NAND U3212 ( .A(n2407), .B(n2406), .Z(n2411) );
  NAND U3213 ( .A(n2409), .B(n2408), .Z(n2410) );
  AND U3214 ( .A(n2411), .B(n2410), .Z(n2413) );
  XNOR U3215 ( .A(n2412), .B(n2413), .Z(n2414) );
  XOR U3216 ( .A(n2415), .B(n2414), .Z(n2525) );
  XOR U3217 ( .A(n2526), .B(n2525), .Z(c[88]) );
  NANDN U3218 ( .A(n2413), .B(n2412), .Z(n2417) );
  NAND U3219 ( .A(n2415), .B(n2414), .Z(n2416) );
  NAND U3220 ( .A(n2417), .B(n2416), .Z(n2537) );
  NANDN U3221 ( .A(n2419), .B(n2418), .Z(n2423) );
  NANDN U3222 ( .A(n2421), .B(n2420), .Z(n2422) );
  NAND U3223 ( .A(n2423), .B(n2422), .Z(n2535) );
  NANDN U3224 ( .A(n2425), .B(n2424), .Z(n2429) );
  NANDN U3225 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U3226 ( .A(n2429), .B(n2428), .Z(n2538) );
  OR U3227 ( .A(n2431), .B(n2430), .Z(n2435) );
  NANDN U3228 ( .A(n2433), .B(n2432), .Z(n2434) );
  NAND U3229 ( .A(n2435), .B(n2434), .Z(n2539) );
  XNOR U3230 ( .A(n2538), .B(n2539), .Z(n2540) );
  NANDN U3231 ( .A(n2437), .B(n2436), .Z(n2441) );
  NAND U3232 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U3233 ( .A(n2441), .B(n2440), .Z(n2629) );
  XNOR U3234 ( .A(n2629), .B(n2630), .Z(n2631) );
  NANDN U3235 ( .A(n2447), .B(n2446), .Z(n2451) );
  NAND U3236 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U3237 ( .A(n2451), .B(n2450), .Z(n2623) );
  NANDN U3238 ( .A(n34510), .B(b[24]), .Z(n34509) );
  NAND U3239 ( .A(n34509), .B(b[25]), .Z(n34814) );
  ANDN U3240 ( .B(n34510), .A(b[24]), .Z(n2452) );
  OR U3241 ( .A(n2452), .B(n986), .Z(n2453) );
  NANDN U3242 ( .A(n34814), .B(n2453), .Z(n2611) );
  XOR U3243 ( .A(b[3]), .B(n16269), .Z(n2582) );
  NANDN U3244 ( .A(n2582), .B(n28939), .Z(n2456) );
  NANDN U3245 ( .A(n2454), .B(n28938), .Z(n2455) );
  NAND U3246 ( .A(n2456), .B(n2455), .Z(n2612) );
  XNOR U3247 ( .A(n2611), .B(n2612), .Z(n2613) );
  NANDN U3248 ( .A(n2457), .B(n32011), .Z(n2459) );
  XOR U3249 ( .A(b[15]), .B(n12830), .Z(n2579) );
  OR U3250 ( .A(n2579), .B(n32010), .Z(n2458) );
  AND U3251 ( .A(n2459), .B(n2458), .Z(n2614) );
  XNOR U3252 ( .A(n2613), .B(n2614), .Z(n2624) );
  XNOR U3253 ( .A(n2623), .B(n2624), .Z(n2625) );
  NAND U3254 ( .A(n2460), .B(n34044), .Z(n2462) );
  XNOR U3255 ( .A(n34510), .B(a[3]), .Z(n2568) );
  NANDN U3256 ( .A(n33867), .B(n2568), .Z(n2461) );
  NAND U3257 ( .A(n2462), .B(n2461), .Z(n2578) );
  XNOR U3258 ( .A(b[25]), .B(n34510), .Z(n2604) );
  XNOR U3259 ( .A(b[25]), .B(n986), .Z(n2463) );
  NAND U3260 ( .A(n2604), .B(n2463), .Z(n2464) );
  XNOR U3261 ( .A(b[25]), .B(b[24]), .Z(n2603) );
  OR U3262 ( .A(n2464), .B(n2603), .Z(n2466) );
  XNOR U3263 ( .A(b[25]), .B(a[1]), .Z(n2605) );
  OR U3264 ( .A(n2605), .B(n34219), .Z(n2465) );
  NAND U3265 ( .A(n2466), .B(n2465), .Z(n2577) );
  XNOR U3266 ( .A(n2578), .B(n2577), .Z(n2620) );
  NANDN U3267 ( .A(n966), .B(a[25]), .Z(n2467) );
  XOR U3268 ( .A(n29232), .B(n2467), .Z(n2469) );
  IV U3269 ( .A(a[24]), .Z(n16508) );
  NANDN U3270 ( .A(n16508), .B(n966), .Z(n2468) );
  AND U3271 ( .A(n2469), .B(n2468), .Z(n2618) );
  NAND U3272 ( .A(n31874), .B(n2470), .Z(n2472) );
  XNOR U3273 ( .A(n971), .B(a[13]), .Z(n2588) );
  NANDN U3274 ( .A(n31550), .B(n2588), .Z(n2471) );
  AND U3275 ( .A(n2472), .B(n2471), .Z(n2617) );
  XNOR U3276 ( .A(n2618), .B(n2617), .Z(n2619) );
  XOR U3277 ( .A(n2620), .B(n2619), .Z(n2626) );
  XOR U3278 ( .A(n2625), .B(n2626), .Z(n2632) );
  XOR U3279 ( .A(n2631), .B(n2632), .Z(n2641) );
  OR U3280 ( .A(n2474), .B(n2473), .Z(n2478) );
  OR U3281 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U3282 ( .A(n2478), .B(n2477), .Z(n2642) );
  XNOR U3283 ( .A(n2641), .B(n2642), .Z(n2644) );
  NANDN U3284 ( .A(n2480), .B(n2479), .Z(n2484) );
  NAND U3285 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3286 ( .A(n2484), .B(n2483), .Z(n2635) );
  XOR U3287 ( .A(n31123), .B(n15113), .Z(n2556) );
  NAND U3288 ( .A(n2556), .B(n29949), .Z(n2487) );
  NAND U3289 ( .A(n29948), .B(n2485), .Z(n2486) );
  NAND U3290 ( .A(n2487), .B(n2486), .Z(n2574) );
  XOR U3291 ( .A(b[5]), .B(n16220), .Z(n2585) );
  OR U3292 ( .A(n2585), .B(n29363), .Z(n2490) );
  NANDN U3293 ( .A(n2488), .B(n29864), .Z(n2489) );
  NAND U3294 ( .A(n2490), .B(n2489), .Z(n2571) );
  XNOR U3295 ( .A(b[17]), .B(a[9]), .Z(n2608) );
  NANDN U3296 ( .A(n2608), .B(n32543), .Z(n2493) );
  NANDN U3297 ( .A(n2491), .B(n32541), .Z(n2492) );
  AND U3298 ( .A(n2493), .B(n2492), .Z(n2572) );
  XNOR U3299 ( .A(n2571), .B(n2572), .Z(n2573) );
  XNOR U3300 ( .A(n2574), .B(n2573), .Z(n2597) );
  NAND U3301 ( .A(n2494), .B(n33283), .Z(n2496) );
  XOR U3302 ( .A(n33020), .B(n11694), .Z(n2591) );
  NANDN U3303 ( .A(n33021), .B(n2591), .Z(n2495) );
  NAND U3304 ( .A(n2496), .B(n2495), .Z(n2553) );
  XNOR U3305 ( .A(b[21]), .B(a[5]), .Z(n2600) );
  OR U3306 ( .A(n2600), .B(n33634), .Z(n2499) );
  NAND U3307 ( .A(n2497), .B(n33464), .Z(n2498) );
  NAND U3308 ( .A(n2499), .B(n2498), .Z(n2550) );
  XOR U3309 ( .A(b[9]), .B(n14514), .Z(n2559) );
  NANDN U3310 ( .A(n2559), .B(n30509), .Z(n2502) );
  NAND U3311 ( .A(n2500), .B(n30846), .Z(n2501) );
  AND U3312 ( .A(n2502), .B(n2501), .Z(n2551) );
  XNOR U3313 ( .A(n2550), .B(n2551), .Z(n2552) );
  XNOR U3314 ( .A(n2553), .B(n2552), .Z(n2594) );
  XNOR U3315 ( .A(n970), .B(a[15]), .Z(n2562) );
  NANDN U3316 ( .A(n31369), .B(n2562), .Z(n2505) );
  NANDN U3317 ( .A(n2503), .B(n31119), .Z(n2504) );
  NAND U3318 ( .A(n2505), .B(n2504), .Z(n2595) );
  XNOR U3319 ( .A(n2594), .B(n2595), .Z(n2596) );
  XOR U3320 ( .A(n2597), .B(n2596), .Z(n2636) );
  XNOR U3321 ( .A(n2635), .B(n2636), .Z(n2637) );
  NANDN U3322 ( .A(n2507), .B(n2506), .Z(n2511) );
  NAND U3323 ( .A(n2509), .B(n2508), .Z(n2510) );
  AND U3324 ( .A(n2511), .B(n2510), .Z(n2638) );
  XNOR U3325 ( .A(n2637), .B(n2638), .Z(n2643) );
  XNOR U3326 ( .A(n2644), .B(n2643), .Z(n2547) );
  NANDN U3327 ( .A(n2513), .B(n2512), .Z(n2517) );
  NANDN U3328 ( .A(n2515), .B(n2514), .Z(n2516) );
  NAND U3329 ( .A(n2517), .B(n2516), .Z(n2544) );
  NANDN U3330 ( .A(n2519), .B(n2518), .Z(n2523) );
  NAND U3331 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U3332 ( .A(n2523), .B(n2522), .Z(n2545) );
  XNOR U3333 ( .A(n2544), .B(n2545), .Z(n2546) );
  XOR U3334 ( .A(n2547), .B(n2546), .Z(n2541) );
  XOR U3335 ( .A(n2540), .B(n2541), .Z(n2534) );
  XNOR U3336 ( .A(n2535), .B(n2534), .Z(n2536) );
  XNOR U3337 ( .A(n2537), .B(n2536), .Z(n2529) );
  XNOR U3338 ( .A(n2529), .B(sreg[89]), .Z(n2531) );
  NAND U3339 ( .A(n2524), .B(sreg[88]), .Z(n2528) );
  OR U3340 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U3341 ( .A(n2528), .B(n2527), .Z(n2530) );
  XOR U3342 ( .A(n2531), .B(n2530), .Z(c[89]) );
  NAND U3343 ( .A(n2529), .B(sreg[89]), .Z(n2533) );
  OR U3344 ( .A(n2531), .B(n2530), .Z(n2532) );
  NAND U3345 ( .A(n2533), .B(n2532), .Z(n2770) );
  XNOR U3346 ( .A(n2770), .B(sreg[90]), .Z(n2772) );
  NANDN U3347 ( .A(n2539), .B(n2538), .Z(n2543) );
  NAND U3348 ( .A(n2541), .B(n2540), .Z(n2542) );
  NAND U3349 ( .A(n2543), .B(n2542), .Z(n2648) );
  NANDN U3350 ( .A(n2545), .B(n2544), .Z(n2549) );
  NAND U3351 ( .A(n2547), .B(n2546), .Z(n2548) );
  NAND U3352 ( .A(n2549), .B(n2548), .Z(n2765) );
  NANDN U3353 ( .A(n2551), .B(n2550), .Z(n2555) );
  NAND U3354 ( .A(n2553), .B(n2552), .Z(n2554) );
  NAND U3355 ( .A(n2555), .B(n2554), .Z(n2661) );
  XOR U3356 ( .A(n31123), .B(n15484), .Z(n2730) );
  NAND U3357 ( .A(n2730), .B(n29949), .Z(n2558) );
  NAND U3358 ( .A(n29948), .B(n2556), .Z(n2557) );
  NAND U3359 ( .A(n2558), .B(n2557), .Z(n2749) );
  XOR U3360 ( .A(b[9]), .B(n14905), .Z(n2677) );
  NANDN U3361 ( .A(n2677), .B(n30509), .Z(n2561) );
  NANDN U3362 ( .A(n2559), .B(n30846), .Z(n2560) );
  NAND U3363 ( .A(n2561), .B(n2560), .Z(n2746) );
  XOR U3364 ( .A(b[11]), .B(n14259), .Z(n2686) );
  OR U3365 ( .A(n2686), .B(n31369), .Z(n2564) );
  NAND U3366 ( .A(n2562), .B(n31119), .Z(n2563) );
  AND U3367 ( .A(n2564), .B(n2563), .Z(n2747) );
  XNOR U3368 ( .A(n2746), .B(n2747), .Z(n2748) );
  XNOR U3369 ( .A(n2749), .B(n2748), .Z(n2659) );
  XOR U3370 ( .A(b[25]), .B(b[26]), .Z(n34618) );
  NAND U3371 ( .A(a[0]), .B(n34618), .Z(n2704) );
  NANDN U3372 ( .A(n966), .B(a[26]), .Z(n2565) );
  XOR U3373 ( .A(n29232), .B(n2565), .Z(n2567) );
  IV U3374 ( .A(a[25]), .Z(n16916) );
  NANDN U3375 ( .A(n16916), .B(n966), .Z(n2566) );
  AND U3376 ( .A(n2567), .B(n2566), .Z(n2702) );
  NAND U3377 ( .A(n2568), .B(n34044), .Z(n2570) );
  XNOR U3378 ( .A(n34510), .B(a[4]), .Z(n2683) );
  NANDN U3379 ( .A(n33867), .B(n2683), .Z(n2569) );
  AND U3380 ( .A(n2570), .B(n2569), .Z(n2701) );
  XNOR U3381 ( .A(n2702), .B(n2701), .Z(n2703) );
  XNOR U3382 ( .A(n2704), .B(n2703), .Z(n2660) );
  XOR U3383 ( .A(n2659), .B(n2660), .Z(n2662) );
  XOR U3384 ( .A(n2661), .B(n2662), .Z(n2754) );
  NANDN U3385 ( .A(n2572), .B(n2571), .Z(n2576) );
  NAND U3386 ( .A(n2574), .B(n2573), .Z(n2575) );
  NAND U3387 ( .A(n2576), .B(n2575), .Z(n2674) );
  NAND U3388 ( .A(n2578), .B(n2577), .Z(n2738) );
  NANDN U3389 ( .A(n2579), .B(n32011), .Z(n2581) );
  XOR U3390 ( .A(b[15]), .B(n13106), .Z(n2698) );
  OR U3391 ( .A(n2698), .B(n32010), .Z(n2580) );
  NAND U3392 ( .A(n2581), .B(n2580), .Z(n2737) );
  XOR U3393 ( .A(b[3]), .B(n16508), .Z(n2695) );
  NANDN U3394 ( .A(n2695), .B(n28939), .Z(n2584) );
  NANDN U3395 ( .A(n2582), .B(n28938), .Z(n2583) );
  AND U3396 ( .A(n2584), .B(n2583), .Z(n2736) );
  XNOR U3397 ( .A(n2737), .B(n2736), .Z(n2739) );
  XNOR U3398 ( .A(n2738), .B(n2739), .Z(n2671) );
  XOR U3399 ( .A(b[5]), .B(n15963), .Z(n2733) );
  OR U3400 ( .A(n2733), .B(n29363), .Z(n2587) );
  NANDN U3401 ( .A(n2585), .B(n29864), .Z(n2586) );
  NAND U3402 ( .A(n2587), .B(n2586), .Z(n2710) );
  XOR U3403 ( .A(n971), .B(n14210), .Z(n2724) );
  NANDN U3404 ( .A(n31550), .B(n2724), .Z(n2590) );
  NAND U3405 ( .A(n2588), .B(n31874), .Z(n2589) );
  NAND U3406 ( .A(n2590), .B(n2589), .Z(n2707) );
  NAND U3407 ( .A(n33283), .B(n2591), .Z(n2593) );
  XOR U3408 ( .A(n33020), .B(n11986), .Z(n2727) );
  NANDN U3409 ( .A(n33021), .B(n2727), .Z(n2592) );
  AND U3410 ( .A(n2593), .B(n2592), .Z(n2708) );
  XNOR U3411 ( .A(n2707), .B(n2708), .Z(n2709) );
  XNOR U3412 ( .A(n2710), .B(n2709), .Z(n2672) );
  XNOR U3413 ( .A(n2671), .B(n2672), .Z(n2673) );
  XOR U3414 ( .A(n2674), .B(n2673), .Z(n2752) );
  NANDN U3415 ( .A(n2595), .B(n2594), .Z(n2599) );
  NAND U3416 ( .A(n2597), .B(n2596), .Z(n2598) );
  AND U3417 ( .A(n2599), .B(n2598), .Z(n2753) );
  XNOR U3418 ( .A(n2752), .B(n2753), .Z(n2755) );
  XNOR U3419 ( .A(n2754), .B(n2755), .Z(n2656) );
  XNOR U3420 ( .A(b[21]), .B(a[6]), .Z(n2680) );
  OR U3421 ( .A(n2680), .B(n33634), .Z(n2602) );
  NANDN U3422 ( .A(n2600), .B(n33464), .Z(n2601) );
  NAND U3423 ( .A(n2602), .B(n2601), .Z(n2743) );
  XNOR U3424 ( .A(b[25]), .B(n10363), .Z(n2713) );
  NANDN U3425 ( .A(n34219), .B(n2713), .Z(n2607) );
  ANDN U3426 ( .B(n2604), .A(n2603), .Z(n34217) );
  NANDN U3427 ( .A(n2605), .B(n34217), .Z(n2606) );
  NAND U3428 ( .A(n2607), .B(n2606), .Z(n2740) );
  XNOR U3429 ( .A(b[17]), .B(a[10]), .Z(n2689) );
  NANDN U3430 ( .A(n2689), .B(n32543), .Z(n2610) );
  NANDN U3431 ( .A(n2608), .B(n32541), .Z(n2609) );
  AND U3432 ( .A(n2610), .B(n2609), .Z(n2741) );
  XNOR U3433 ( .A(n2740), .B(n2741), .Z(n2742) );
  XNOR U3434 ( .A(n2743), .B(n2742), .Z(n2668) );
  NANDN U3435 ( .A(n2612), .B(n2611), .Z(n2616) );
  NAND U3436 ( .A(n2614), .B(n2613), .Z(n2615) );
  NAND U3437 ( .A(n2616), .B(n2615), .Z(n2665) );
  NANDN U3438 ( .A(n2618), .B(n2617), .Z(n2622) );
  NAND U3439 ( .A(n2620), .B(n2619), .Z(n2621) );
  AND U3440 ( .A(n2622), .B(n2621), .Z(n2666) );
  XNOR U3441 ( .A(n2665), .B(n2666), .Z(n2667) );
  XOR U3442 ( .A(n2668), .B(n2667), .Z(n2653) );
  NANDN U3443 ( .A(n2624), .B(n2623), .Z(n2628) );
  NAND U3444 ( .A(n2626), .B(n2625), .Z(n2627) );
  NAND U3445 ( .A(n2628), .B(n2627), .Z(n2654) );
  XOR U3446 ( .A(n2653), .B(n2654), .Z(n2655) );
  XNOR U3447 ( .A(n2656), .B(n2655), .Z(n2761) );
  NANDN U3448 ( .A(n2630), .B(n2629), .Z(n2634) );
  NAND U3449 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U3450 ( .A(n2634), .B(n2633), .Z(n2758) );
  NANDN U3451 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U3452 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U3453 ( .A(n2640), .B(n2639), .Z(n2759) );
  XNOR U3454 ( .A(n2758), .B(n2759), .Z(n2760) );
  XNOR U3455 ( .A(n2761), .B(n2760), .Z(n2764) );
  XNOR U3456 ( .A(n2765), .B(n2764), .Z(n2767) );
  OR U3457 ( .A(n2642), .B(n2641), .Z(n2646) );
  OR U3458 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U3459 ( .A(n2646), .B(n2645), .Z(n2766) );
  XNOR U3460 ( .A(n2767), .B(n2766), .Z(n2647) );
  XOR U3461 ( .A(n2648), .B(n2647), .Z(n2649) );
  XOR U3462 ( .A(n2650), .B(n2649), .Z(n2771) );
  XOR U3463 ( .A(n2772), .B(n2771), .Z(c[90]) );
  NAND U3464 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U3465 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U3466 ( .A(n2652), .B(n2651), .Z(n2783) );
  OR U3467 ( .A(n2654), .B(n2653), .Z(n2658) );
  NANDN U3468 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U3469 ( .A(n2658), .B(n2657), .Z(n2899) );
  NANDN U3470 ( .A(n2660), .B(n2659), .Z(n2664) );
  OR U3471 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U3472 ( .A(n2664), .B(n2663), .Z(n2893) );
  NANDN U3473 ( .A(n2666), .B(n2665), .Z(n2670) );
  NAND U3474 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U3475 ( .A(n2670), .B(n2669), .Z(n2890) );
  NANDN U3476 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U3477 ( .A(n2674), .B(n2673), .Z(n2675) );
  NAND U3478 ( .A(n2676), .B(n2675), .Z(n2891) );
  XNOR U3479 ( .A(n2890), .B(n2891), .Z(n2892) );
  XNOR U3480 ( .A(n2893), .B(n2892), .Z(n2896) );
  XOR U3481 ( .A(b[9]), .B(n15113), .Z(n2856) );
  NANDN U3482 ( .A(n2856), .B(n30509), .Z(n2679) );
  NANDN U3483 ( .A(n2677), .B(n30846), .Z(n2678) );
  NAND U3484 ( .A(n2679), .B(n2678), .Z(n2877) );
  XNOR U3485 ( .A(b[21]), .B(n11694), .Z(n2853) );
  NANDN U3486 ( .A(n33634), .B(n2853), .Z(n2682) );
  NANDN U3487 ( .A(n2680), .B(n33464), .Z(n2681) );
  NAND U3488 ( .A(n2682), .B(n2681), .Z(n2874) );
  NAND U3489 ( .A(n2683), .B(n34044), .Z(n2685) );
  XNOR U3490 ( .A(n34510), .B(a[5]), .Z(n2865) );
  NANDN U3491 ( .A(n33867), .B(n2865), .Z(n2684) );
  AND U3492 ( .A(n2685), .B(n2684), .Z(n2875) );
  XNOR U3493 ( .A(n2874), .B(n2875), .Z(n2876) );
  XNOR U3494 ( .A(n2877), .B(n2876), .Z(n2801) );
  XNOR U3495 ( .A(n970), .B(a[17]), .Z(n2841) );
  NANDN U3496 ( .A(n31369), .B(n2841), .Z(n2688) );
  NANDN U3497 ( .A(n2686), .B(n31119), .Z(n2687) );
  NAND U3498 ( .A(n2688), .B(n2687), .Z(n2799) );
  XNOR U3499 ( .A(b[17]), .B(n12830), .Z(n2844) );
  NAND U3500 ( .A(n2844), .B(n32543), .Z(n2691) );
  NANDN U3501 ( .A(n2689), .B(n32541), .Z(n2690) );
  AND U3502 ( .A(n2691), .B(n2690), .Z(n2798) );
  XNOR U3503 ( .A(n2799), .B(n2798), .Z(n2800) );
  XOR U3504 ( .A(n2801), .B(n2800), .Z(n2795) );
  IV U3505 ( .A(b[27]), .Z(n35375) );
  OR U3506 ( .A(b[25]), .B(n35375), .Z(n2692) );
  OR U3507 ( .A(n2692), .B(b[26]), .Z(n2694) );
  ANDN U3508 ( .B(n34618), .A(n35375), .Z(n34849) );
  NANDN U3509 ( .A(a[0]), .B(n34849), .Z(n2693) );
  NAND U3510 ( .A(n2694), .B(n2693), .Z(n2805) );
  XOR U3511 ( .A(b[3]), .B(n16916), .Z(n2862) );
  NANDN U3512 ( .A(n2862), .B(n28939), .Z(n2697) );
  NANDN U3513 ( .A(n2695), .B(n28938), .Z(n2696) );
  AND U3514 ( .A(n2697), .B(n2696), .Z(n2804) );
  XNOR U3515 ( .A(n2805), .B(n2804), .Z(n2806) );
  NANDN U3516 ( .A(n2698), .B(n32011), .Z(n2700) );
  XOR U3517 ( .A(b[15]), .B(n13509), .Z(n2812) );
  OR U3518 ( .A(n2812), .B(n32010), .Z(n2699) );
  NAND U3519 ( .A(n2700), .B(n2699), .Z(n2807) );
  XNOR U3520 ( .A(n2806), .B(n2807), .Z(n2792) );
  NANDN U3521 ( .A(n2702), .B(n2701), .Z(n2706) );
  NAND U3522 ( .A(n2704), .B(n2703), .Z(n2705) );
  NAND U3523 ( .A(n2706), .B(n2705), .Z(n2793) );
  XNOR U3524 ( .A(n2795), .B(n2794), .Z(n2880) );
  NANDN U3525 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U3526 ( .A(n2710), .B(n2709), .Z(n2711) );
  NAND U3527 ( .A(n2712), .B(n2711), .Z(n2881) );
  XOR U3528 ( .A(n2880), .B(n2881), .Z(n2882) );
  XNOR U3529 ( .A(b[25]), .B(n10524), .Z(n2823) );
  NANDN U3530 ( .A(n34219), .B(n2823), .Z(n2715) );
  NAND U3531 ( .A(n34217), .B(n2713), .Z(n2714) );
  NAND U3532 ( .A(n2715), .B(n2714), .Z(n2811) );
  XNOR U3533 ( .A(n35375), .B(a[0]), .Z(n2718) );
  XNOR U3534 ( .A(n35375), .B(b[25]), .Z(n2816) );
  XOR U3535 ( .A(b[27]), .B(b[26]), .Z(n2716) );
  AND U3536 ( .A(n2816), .B(n2716), .Z(n2717) );
  NAND U3537 ( .A(n2718), .B(n2717), .Z(n2720) );
  XOR U3538 ( .A(b[27]), .B(n10457), .Z(n2817) );
  NANDN U3539 ( .A(n2817), .B(n34618), .Z(n2719) );
  NAND U3540 ( .A(n2720), .B(n2719), .Z(n2810) );
  XNOR U3541 ( .A(n2811), .B(n2810), .Z(n2871) );
  NANDN U3542 ( .A(n966), .B(a[27]), .Z(n2721) );
  XOR U3543 ( .A(n29232), .B(n2721), .Z(n2723) );
  IV U3544 ( .A(a[26]), .Z(n17133) );
  NANDN U3545 ( .A(n17133), .B(n966), .Z(n2722) );
  AND U3546 ( .A(n2723), .B(n2722), .Z(n2869) );
  NAND U3547 ( .A(n31874), .B(n2724), .Z(n2726) );
  XOR U3548 ( .A(n971), .B(n13976), .Z(n2859) );
  NANDN U3549 ( .A(n31550), .B(n2859), .Z(n2725) );
  AND U3550 ( .A(n2726), .B(n2725), .Z(n2868) );
  XNOR U3551 ( .A(n2869), .B(n2868), .Z(n2870) );
  XOR U3552 ( .A(n2871), .B(n2870), .Z(n2832) );
  NAND U3553 ( .A(n33283), .B(n2727), .Z(n2729) );
  XNOR U3554 ( .A(n33020), .B(a[9]), .Z(n2850) );
  NANDN U3555 ( .A(n33021), .B(n2850), .Z(n2728) );
  NAND U3556 ( .A(n2729), .B(n2728), .Z(n2829) );
  XOR U3557 ( .A(n31123), .B(n16220), .Z(n2838) );
  NAND U3558 ( .A(n2838), .B(n29949), .Z(n2732) );
  NAND U3559 ( .A(n29948), .B(n2730), .Z(n2731) );
  NAND U3560 ( .A(n2732), .B(n2731), .Z(n2826) );
  XOR U3561 ( .A(n968), .B(n16269), .Z(n2847) );
  NANDN U3562 ( .A(n29363), .B(n2847), .Z(n2735) );
  NANDN U3563 ( .A(n2733), .B(n29864), .Z(n2734) );
  AND U3564 ( .A(n2735), .B(n2734), .Z(n2827) );
  XNOR U3565 ( .A(n2826), .B(n2827), .Z(n2828) );
  XNOR U3566 ( .A(n2829), .B(n2828), .Z(n2833) );
  XOR U3567 ( .A(n2832), .B(n2833), .Z(n2834) );
  XOR U3568 ( .A(n2834), .B(n2835), .Z(n2889) );
  NANDN U3569 ( .A(n2741), .B(n2740), .Z(n2745) );
  NAND U3570 ( .A(n2743), .B(n2742), .Z(n2744) );
  NAND U3571 ( .A(n2745), .B(n2744), .Z(n2887) );
  NANDN U3572 ( .A(n2747), .B(n2746), .Z(n2751) );
  NAND U3573 ( .A(n2749), .B(n2748), .Z(n2750) );
  AND U3574 ( .A(n2751), .B(n2750), .Z(n2886) );
  XNOR U3575 ( .A(n2887), .B(n2886), .Z(n2888) );
  XOR U3576 ( .A(n2889), .B(n2888), .Z(n2883) );
  XNOR U3577 ( .A(n2882), .B(n2883), .Z(n2897) );
  XNOR U3578 ( .A(n2896), .B(n2897), .Z(n2898) );
  XNOR U3579 ( .A(n2899), .B(n2898), .Z(n2787) );
  OR U3580 ( .A(n2753), .B(n2752), .Z(n2757) );
  NANDN U3581 ( .A(n2755), .B(n2754), .Z(n2756) );
  AND U3582 ( .A(n2757), .B(n2756), .Z(n2786) );
  XNOR U3583 ( .A(n2787), .B(n2786), .Z(n2788) );
  NANDN U3584 ( .A(n2759), .B(n2758), .Z(n2763) );
  NANDN U3585 ( .A(n2761), .B(n2760), .Z(n2762) );
  NAND U3586 ( .A(n2763), .B(n2762), .Z(n2789) );
  XOR U3587 ( .A(n2788), .B(n2789), .Z(n2780) );
  NAND U3588 ( .A(n2765), .B(n2764), .Z(n2769) );
  NANDN U3589 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U3590 ( .A(n2769), .B(n2768), .Z(n2781) );
  XNOR U3591 ( .A(n2780), .B(n2781), .Z(n2782) );
  XNOR U3592 ( .A(n2783), .B(n2782), .Z(n2775) );
  XNOR U3593 ( .A(n2775), .B(sreg[91]), .Z(n2777) );
  NAND U3594 ( .A(n2770), .B(sreg[90]), .Z(n2774) );
  OR U3595 ( .A(n2772), .B(n2771), .Z(n2773) );
  AND U3596 ( .A(n2774), .B(n2773), .Z(n2776) );
  XOR U3597 ( .A(n2777), .B(n2776), .Z(c[91]) );
  NAND U3598 ( .A(n2775), .B(sreg[91]), .Z(n2779) );
  OR U3599 ( .A(n2777), .B(n2776), .Z(n2778) );
  NAND U3600 ( .A(n2779), .B(n2778), .Z(n3032) );
  XNOR U3601 ( .A(n3032), .B(sreg[92]), .Z(n3034) );
  NANDN U3602 ( .A(n2781), .B(n2780), .Z(n2785) );
  NAND U3603 ( .A(n2783), .B(n2782), .Z(n2784) );
  NAND U3604 ( .A(n2785), .B(n2784), .Z(n2905) );
  NANDN U3605 ( .A(n2787), .B(n2786), .Z(n2791) );
  NANDN U3606 ( .A(n2789), .B(n2788), .Z(n2790) );
  NAND U3607 ( .A(n2791), .B(n2790), .Z(n2903) );
  OR U3608 ( .A(n2793), .B(n2792), .Z(n2797) );
  NANDN U3609 ( .A(n2795), .B(n2794), .Z(n2796) );
  NAND U3610 ( .A(n2797), .B(n2796), .Z(n2914) );
  NANDN U3611 ( .A(n2799), .B(n2798), .Z(n2803) );
  NAND U3612 ( .A(n2801), .B(n2800), .Z(n2802) );
  NAND U3613 ( .A(n2803), .B(n2802), .Z(n2929) );
  NANDN U3614 ( .A(n2805), .B(n2804), .Z(n2809) );
  NANDN U3615 ( .A(n2807), .B(n2806), .Z(n2808) );
  NAND U3616 ( .A(n2809), .B(n2808), .Z(n2926) );
  NAND U3617 ( .A(n2811), .B(n2810), .Z(n2958) );
  NANDN U3618 ( .A(n2812), .B(n32011), .Z(n2814) );
  XOR U3619 ( .A(b[15]), .B(n14210), .Z(n2935) );
  OR U3620 ( .A(n2935), .B(n32010), .Z(n2813) );
  NAND U3621 ( .A(n2814), .B(n2813), .Z(n2956) );
  XOR U3622 ( .A(n35375), .B(b[26]), .Z(n2815) );
  ANDN U3623 ( .B(n2816), .A(n2815), .Z(n34848) );
  NANDN U3624 ( .A(n2817), .B(n34848), .Z(n2819) );
  XNOR U3625 ( .A(n35375), .B(a[2]), .Z(n2938) );
  NAND U3626 ( .A(n34618), .B(n2938), .Z(n2818) );
  AND U3627 ( .A(n2819), .B(n2818), .Z(n2955) );
  XNOR U3628 ( .A(n2956), .B(n2955), .Z(n2957) );
  XNOR U3629 ( .A(n2958), .B(n2957), .Z(n3026) );
  XOR U3630 ( .A(n35375), .B(b[28]), .Z(n34968) );
  NOR U3631 ( .A(n986), .B(n34968), .Z(n3005) );
  NANDN U3632 ( .A(n966), .B(a[28]), .Z(n2820) );
  XOR U3633 ( .A(n29232), .B(n2820), .Z(n2822) );
  IV U3634 ( .A(a[27]), .Z(n17960) );
  NANDN U3635 ( .A(n17960), .B(n966), .Z(n2821) );
  AND U3636 ( .A(n2822), .B(n2821), .Z(n3003) );
  XNOR U3637 ( .A(b[25]), .B(n10854), .Z(n2996) );
  NANDN U3638 ( .A(n34219), .B(n2996), .Z(n2825) );
  NAND U3639 ( .A(n2823), .B(n34217), .Z(n2824) );
  AND U3640 ( .A(n2825), .B(n2824), .Z(n3002) );
  XNOR U3641 ( .A(n3003), .B(n3002), .Z(n3004) );
  XOR U3642 ( .A(n3005), .B(n3004), .Z(n3027) );
  XOR U3643 ( .A(n3026), .B(n3027), .Z(n3028) );
  NANDN U3644 ( .A(n2827), .B(n2826), .Z(n2831) );
  NAND U3645 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U3646 ( .A(n2831), .B(n2830), .Z(n3029) );
  XNOR U3647 ( .A(n3028), .B(n3029), .Z(n2927) );
  XNOR U3648 ( .A(n2926), .B(n2927), .Z(n2928) );
  XOR U3649 ( .A(n2929), .B(n2928), .Z(n2915) );
  XNOR U3650 ( .A(n2914), .B(n2915), .Z(n2916) );
  OR U3651 ( .A(n2833), .B(n2832), .Z(n2837) );
  NAND U3652 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U3653 ( .A(n2837), .B(n2836), .Z(n3011) );
  XOR U3654 ( .A(n31123), .B(n15963), .Z(n2981) );
  NAND U3655 ( .A(n2981), .B(n29949), .Z(n2840) );
  NAND U3656 ( .A(n29948), .B(n2838), .Z(n2839) );
  NAND U3657 ( .A(n2840), .B(n2839), .Z(n2990) );
  XOR U3658 ( .A(b[11]), .B(n14905), .Z(n2952) );
  OR U3659 ( .A(n2952), .B(n31369), .Z(n2843) );
  NAND U3660 ( .A(n2841), .B(n31119), .Z(n2842) );
  NAND U3661 ( .A(n2843), .B(n2842), .Z(n2987) );
  XNOR U3662 ( .A(b[17]), .B(a[12]), .Z(n2971) );
  NANDN U3663 ( .A(n2971), .B(n32543), .Z(n2846) );
  NAND U3664 ( .A(n2844), .B(n32541), .Z(n2845) );
  AND U3665 ( .A(n2846), .B(n2845), .Z(n2988) );
  XNOR U3666 ( .A(n2987), .B(n2988), .Z(n2989) );
  XNOR U3667 ( .A(n2990), .B(n2989), .Z(n3017) );
  NAND U3668 ( .A(n29864), .B(n2847), .Z(n2849) );
  XNOR U3669 ( .A(n968), .B(a[24]), .Z(n2965) );
  NANDN U3670 ( .A(n29363), .B(n2965), .Z(n2848) );
  NAND U3671 ( .A(n2849), .B(n2848), .Z(n2976) );
  NAND U3672 ( .A(n2850), .B(n33283), .Z(n2852) );
  XNOR U3673 ( .A(n33020), .B(a[10]), .Z(n2949) );
  NANDN U3674 ( .A(n33021), .B(n2949), .Z(n2851) );
  NAND U3675 ( .A(n2852), .B(n2851), .Z(n2974) );
  XNOR U3676 ( .A(b[21]), .B(a[8]), .Z(n2984) );
  OR U3677 ( .A(n2984), .B(n33634), .Z(n2855) );
  NAND U3678 ( .A(n2853), .B(n33464), .Z(n2854) );
  NAND U3679 ( .A(n2855), .B(n2854), .Z(n2975) );
  XNOR U3680 ( .A(n2974), .B(n2975), .Z(n2977) );
  XOR U3681 ( .A(n2976), .B(n2977), .Z(n3014) );
  NANDN U3682 ( .A(n2856), .B(n30846), .Z(n2858) );
  XNOR U3683 ( .A(n969), .B(a[20]), .Z(n2999) );
  NAND U3684 ( .A(n30509), .B(n2999), .Z(n2857) );
  NAND U3685 ( .A(n2858), .B(n2857), .Z(n3015) );
  XNOR U3686 ( .A(n3014), .B(n3015), .Z(n3016) );
  XOR U3687 ( .A(n3017), .B(n3016), .Z(n3009) );
  NAND U3688 ( .A(n31874), .B(n2859), .Z(n2861) );
  XNOR U3689 ( .A(n971), .B(a[16]), .Z(n2946) );
  NANDN U3690 ( .A(n31550), .B(n2946), .Z(n2860) );
  NAND U3691 ( .A(n2861), .B(n2860), .Z(n2963) );
  XNOR U3692 ( .A(n967), .B(a[26]), .Z(n2968) );
  NAND U3693 ( .A(n2968), .B(n28939), .Z(n2864) );
  NANDN U3694 ( .A(n2862), .B(n28938), .Z(n2863) );
  NAND U3695 ( .A(n2864), .B(n2863), .Z(n2961) );
  NAND U3696 ( .A(n2865), .B(n34044), .Z(n2867) );
  XNOR U3697 ( .A(n34510), .B(a[6]), .Z(n2993) );
  NANDN U3698 ( .A(n33867), .B(n2993), .Z(n2866) );
  NAND U3699 ( .A(n2867), .B(n2866), .Z(n2962) );
  XNOR U3700 ( .A(n2961), .B(n2962), .Z(n2964) );
  XOR U3701 ( .A(n2963), .B(n2964), .Z(n3023) );
  NANDN U3702 ( .A(n2869), .B(n2868), .Z(n2873) );
  NAND U3703 ( .A(n2871), .B(n2870), .Z(n2872) );
  NAND U3704 ( .A(n2873), .B(n2872), .Z(n3020) );
  NANDN U3705 ( .A(n2875), .B(n2874), .Z(n2879) );
  NAND U3706 ( .A(n2877), .B(n2876), .Z(n2878) );
  NAND U3707 ( .A(n2879), .B(n2878), .Z(n3021) );
  XNOR U3708 ( .A(n3020), .B(n3021), .Z(n3022) );
  XOR U3709 ( .A(n3023), .B(n3022), .Z(n3008) );
  XOR U3710 ( .A(n3009), .B(n3008), .Z(n3010) );
  XNOR U3711 ( .A(n3011), .B(n3010), .Z(n2917) );
  XOR U3712 ( .A(n2916), .B(n2917), .Z(n2911) );
  OR U3713 ( .A(n2881), .B(n2880), .Z(n2885) );
  NANDN U3714 ( .A(n2883), .B(n2882), .Z(n2884) );
  NAND U3715 ( .A(n2885), .B(n2884), .Z(n2921) );
  XNOR U3716 ( .A(n2921), .B(n2920), .Z(n2922) );
  NANDN U3717 ( .A(n2891), .B(n2890), .Z(n2895) );
  NAND U3718 ( .A(n2893), .B(n2892), .Z(n2894) );
  NAND U3719 ( .A(n2895), .B(n2894), .Z(n2923) );
  XOR U3720 ( .A(n2922), .B(n2923), .Z(n2908) );
  NANDN U3721 ( .A(n2897), .B(n2896), .Z(n2901) );
  NAND U3722 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U3723 ( .A(n2901), .B(n2900), .Z(n2909) );
  XNOR U3724 ( .A(n2908), .B(n2909), .Z(n2910) );
  XOR U3725 ( .A(n2911), .B(n2910), .Z(n2902) );
  XNOR U3726 ( .A(n2903), .B(n2902), .Z(n2904) );
  XOR U3727 ( .A(n2905), .B(n2904), .Z(n3033) );
  XOR U3728 ( .A(n3034), .B(n3033), .Z(c[92]) );
  NANDN U3729 ( .A(n2903), .B(n2902), .Z(n2907) );
  NAND U3730 ( .A(n2905), .B(n2904), .Z(n2906) );
  NAND U3731 ( .A(n2907), .B(n2906), .Z(n3045) );
  NANDN U3732 ( .A(n2909), .B(n2908), .Z(n2913) );
  NAND U3733 ( .A(n2911), .B(n2910), .Z(n2912) );
  NAND U3734 ( .A(n2913), .B(n2912), .Z(n3043) );
  NANDN U3735 ( .A(n2915), .B(n2914), .Z(n2919) );
  NANDN U3736 ( .A(n2917), .B(n2916), .Z(n2918) );
  NAND U3737 ( .A(n2919), .B(n2918), .Z(n3049) );
  NANDN U3738 ( .A(n2921), .B(n2920), .Z(n2925) );
  NANDN U3739 ( .A(n2923), .B(n2922), .Z(n2924) );
  AND U3740 ( .A(n2925), .B(n2924), .Z(n3048) );
  XNOR U3741 ( .A(n3049), .B(n3048), .Z(n3050) );
  NANDN U3742 ( .A(n2927), .B(n2926), .Z(n2931) );
  NAND U3743 ( .A(n2929), .B(n2928), .Z(n2930) );
  NAND U3744 ( .A(n2931), .B(n2930), .Z(n3056) );
  NANDN U3745 ( .A(n966), .B(a[29]), .Z(n2932) );
  XOR U3746 ( .A(n29232), .B(n2932), .Z(n2934) );
  IV U3747 ( .A(a[28]), .Z(n17702) );
  NANDN U3748 ( .A(n17702), .B(n966), .Z(n2933) );
  AND U3749 ( .A(n2934), .B(n2933), .Z(n3107) );
  NANDN U3750 ( .A(n2935), .B(n32011), .Z(n2937) );
  XNOR U3751 ( .A(n972), .B(a[15]), .Z(n3097) );
  NANDN U3752 ( .A(n32010), .B(n3097), .Z(n2936) );
  AND U3753 ( .A(n2937), .B(n2936), .Z(n3106) );
  XNOR U3754 ( .A(n3107), .B(n3106), .Z(n3108) );
  NAND U3755 ( .A(n2938), .B(n34848), .Z(n2940) );
  XNOR U3756 ( .A(n35375), .B(a[3]), .Z(n3141) );
  NAND U3757 ( .A(n34618), .B(n3141), .Z(n2939) );
  NAND U3758 ( .A(n2940), .B(n2939), .Z(n3088) );
  IV U3759 ( .A(b[29]), .Z(n35540) );
  XNOR U3760 ( .A(n35540), .B(b[27]), .Z(n2942) );
  XNOR U3761 ( .A(n35540), .B(a[0]), .Z(n2941) );
  NAND U3762 ( .A(n2942), .B(n2941), .Z(n2943) );
  XOR U3763 ( .A(b[29]), .B(b[28]), .Z(n3092) );
  NANDN U3764 ( .A(n2943), .B(n3092), .Z(n2945) );
  XOR U3765 ( .A(b[29]), .B(n10457), .Z(n3094) );
  OR U3766 ( .A(n3094), .B(n34968), .Z(n2944) );
  NAND U3767 ( .A(n2945), .B(n2944), .Z(n3087) );
  XOR U3768 ( .A(n3088), .B(n3087), .Z(n3109) );
  XOR U3769 ( .A(n3108), .B(n3109), .Z(n3118) );
  XOR U3770 ( .A(b[13]), .B(n14514), .Z(n3075) );
  OR U3771 ( .A(n3075), .B(n31550), .Z(n2948) );
  NAND U3772 ( .A(n2946), .B(n31874), .Z(n2947) );
  NAND U3773 ( .A(n2948), .B(n2947), .Z(n3115) );
  NAND U3774 ( .A(n2949), .B(n33283), .Z(n2951) );
  XOR U3775 ( .A(n33020), .B(n12830), .Z(n3078) );
  NANDN U3776 ( .A(n33021), .B(n3078), .Z(n2950) );
  NAND U3777 ( .A(n2951), .B(n2950), .Z(n3112) );
  XOR U3778 ( .A(b[11]), .B(n15113), .Z(n3081) );
  OR U3779 ( .A(n3081), .B(n31369), .Z(n2954) );
  NANDN U3780 ( .A(n2952), .B(n31119), .Z(n2953) );
  AND U3781 ( .A(n2954), .B(n2953), .Z(n3113) );
  XNOR U3782 ( .A(n3112), .B(n3113), .Z(n3114) );
  XNOR U3783 ( .A(n3115), .B(n3114), .Z(n3119) );
  XNOR U3784 ( .A(n3118), .B(n3119), .Z(n3120) );
  NANDN U3785 ( .A(n2956), .B(n2955), .Z(n2960) );
  NAND U3786 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U3787 ( .A(n2960), .B(n2959), .Z(n3121) );
  XOR U3788 ( .A(n3120), .B(n3121), .Z(n3127) );
  XOR U3789 ( .A(b[5]), .B(n16916), .Z(n3100) );
  OR U3790 ( .A(n3100), .B(n29363), .Z(n2967) );
  NAND U3791 ( .A(n2965), .B(n29864), .Z(n2966) );
  NAND U3792 ( .A(n2967), .B(n2966), .Z(n3135) );
  XOR U3793 ( .A(n967), .B(n17960), .Z(n3103) );
  NAND U3794 ( .A(n3103), .B(n28939), .Z(n2970) );
  NAND U3795 ( .A(n2968), .B(n28938), .Z(n2969) );
  NAND U3796 ( .A(n2970), .B(n2969), .Z(n3132) );
  XNOR U3797 ( .A(b[17]), .B(a[13]), .Z(n3089) );
  NANDN U3798 ( .A(n3089), .B(n32543), .Z(n2973) );
  NANDN U3799 ( .A(n2971), .B(n32541), .Z(n2972) );
  AND U3800 ( .A(n2973), .B(n2972), .Z(n3133) );
  XNOR U3801 ( .A(n3132), .B(n3133), .Z(n3134) );
  XOR U3802 ( .A(n3135), .B(n3134), .Z(n3128) );
  XNOR U3803 ( .A(n3128), .B(n3129), .Z(n3131) );
  OR U3804 ( .A(b[28]), .B(n35540), .Z(n2978) );
  OR U3805 ( .A(n2978), .B(b[27]), .Z(n2980) );
  ANDN U3806 ( .B(b[29]), .A(n34968), .Z(n35189) );
  NANDN U3807 ( .A(a[0]), .B(n35189), .Z(n2979) );
  NAND U3808 ( .A(n2980), .B(n2979), .Z(n3154) );
  XNOR U3809 ( .A(n31123), .B(a[23]), .Z(n3072) );
  NAND U3810 ( .A(n3072), .B(n29949), .Z(n2983) );
  NAND U3811 ( .A(n2981), .B(n29948), .Z(n2982) );
  AND U3812 ( .A(n2983), .B(n2982), .Z(n3153) );
  XNOR U3813 ( .A(n3154), .B(n3153), .Z(n3155) );
  XNOR U3814 ( .A(b[21]), .B(n12258), .Z(n3144) );
  NANDN U3815 ( .A(n33634), .B(n3144), .Z(n2986) );
  NANDN U3816 ( .A(n2984), .B(n33464), .Z(n2985) );
  NAND U3817 ( .A(n2986), .B(n2985), .Z(n3156) );
  XNOR U3818 ( .A(n3155), .B(n3156), .Z(n3130) );
  XNOR U3819 ( .A(n3131), .B(n3130), .Z(n3124) );
  XNOR U3820 ( .A(n3125), .B(n3124), .Z(n3126) );
  XNOR U3821 ( .A(n3127), .B(n3126), .Z(n3054) );
  NANDN U3822 ( .A(n2988), .B(n2987), .Z(n2992) );
  NAND U3823 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U3824 ( .A(n2992), .B(n2991), .Z(n3069) );
  NAND U3825 ( .A(n2993), .B(n34044), .Z(n2995) );
  XOR U3826 ( .A(n34510), .B(n11694), .Z(n3147) );
  NANDN U3827 ( .A(n33867), .B(n3147), .Z(n2994) );
  NAND U3828 ( .A(n2995), .B(n2994), .Z(n3162) );
  XNOR U3829 ( .A(b[25]), .B(n11202), .Z(n3150) );
  NANDN U3830 ( .A(n34219), .B(n3150), .Z(n2998) );
  NAND U3831 ( .A(n2996), .B(n34217), .Z(n2997) );
  AND U3832 ( .A(n2998), .B(n2997), .Z(n3159) );
  XOR U3833 ( .A(n969), .B(n16220), .Z(n3084) );
  NAND U3834 ( .A(n30509), .B(n3084), .Z(n3001) );
  NAND U3835 ( .A(n2999), .B(n30846), .Z(n3000) );
  AND U3836 ( .A(n3001), .B(n3000), .Z(n3160) );
  XNOR U3837 ( .A(n3162), .B(n3161), .Z(n3067) );
  NANDN U3838 ( .A(n3003), .B(n3002), .Z(n3007) );
  NANDN U3839 ( .A(n3005), .B(n3004), .Z(n3006) );
  AND U3840 ( .A(n3007), .B(n3006), .Z(n3066) );
  XNOR U3841 ( .A(n3067), .B(n3066), .Z(n3068) );
  XNOR U3842 ( .A(n3069), .B(n3068), .Z(n3055) );
  XOR U3843 ( .A(n3054), .B(n3055), .Z(n3057) );
  XNOR U3844 ( .A(n3056), .B(n3057), .Z(n3168) );
  OR U3845 ( .A(n3009), .B(n3008), .Z(n3013) );
  NAND U3846 ( .A(n3011), .B(n3010), .Z(n3012) );
  NAND U3847 ( .A(n3013), .B(n3012), .Z(n3166) );
  NANDN U3848 ( .A(n3015), .B(n3014), .Z(n3019) );
  NAND U3849 ( .A(n3017), .B(n3016), .Z(n3018) );
  NAND U3850 ( .A(n3019), .B(n3018), .Z(n3063) );
  NANDN U3851 ( .A(n3021), .B(n3020), .Z(n3025) );
  NAND U3852 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U3853 ( .A(n3025), .B(n3024), .Z(n3060) );
  OR U3854 ( .A(n3027), .B(n3026), .Z(n3031) );
  NAND U3855 ( .A(n3029), .B(n3028), .Z(n3030) );
  AND U3856 ( .A(n3031), .B(n3030), .Z(n3061) );
  XNOR U3857 ( .A(n3060), .B(n3061), .Z(n3062) );
  XOR U3858 ( .A(n3063), .B(n3062), .Z(n3165) );
  XNOR U3859 ( .A(n3166), .B(n3165), .Z(n3167) );
  XNOR U3860 ( .A(n3168), .B(n3167), .Z(n3051) );
  XNOR U3861 ( .A(n3050), .B(n3051), .Z(n3042) );
  XOR U3862 ( .A(n3043), .B(n3042), .Z(n3044) );
  XNOR U3863 ( .A(n3045), .B(n3044), .Z(n3037) );
  XNOR U3864 ( .A(n3037), .B(sreg[93]), .Z(n3039) );
  NAND U3865 ( .A(n3032), .B(sreg[92]), .Z(n3036) );
  OR U3866 ( .A(n3034), .B(n3033), .Z(n3035) );
  AND U3867 ( .A(n3036), .B(n3035), .Z(n3038) );
  XOR U3868 ( .A(n3039), .B(n3038), .Z(c[93]) );
  NAND U3869 ( .A(n3037), .B(sreg[93]), .Z(n3041) );
  OR U3870 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3871 ( .A(n3041), .B(n3040), .Z(n3307) );
  XNOR U3872 ( .A(n3307), .B(sreg[94]), .Z(n3309) );
  NAND U3873 ( .A(n3043), .B(n3042), .Z(n3047) );
  NAND U3874 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U3875 ( .A(n3047), .B(n3046), .Z(n3172) );
  NANDN U3876 ( .A(n3049), .B(n3048), .Z(n3053) );
  NANDN U3877 ( .A(n3051), .B(n3050), .Z(n3052) );
  NAND U3878 ( .A(n3053), .B(n3052), .Z(n3169) );
  NANDN U3879 ( .A(n3055), .B(n3054), .Z(n3059) );
  OR U3880 ( .A(n3057), .B(n3056), .Z(n3058) );
  NAND U3881 ( .A(n3059), .B(n3058), .Z(n3301) );
  NANDN U3882 ( .A(n3061), .B(n3060), .Z(n3065) );
  NAND U3883 ( .A(n3063), .B(n3062), .Z(n3064) );
  NAND U3884 ( .A(n3065), .B(n3064), .Z(n3289) );
  NANDN U3885 ( .A(n3067), .B(n3066), .Z(n3071) );
  NAND U3886 ( .A(n3069), .B(n3068), .Z(n3070) );
  NAND U3887 ( .A(n3071), .B(n3070), .Z(n3286) );
  XOR U3888 ( .A(n31123), .B(n16508), .Z(n3252) );
  NAND U3889 ( .A(n3252), .B(n29949), .Z(n3074) );
  NAND U3890 ( .A(n3072), .B(n29948), .Z(n3073) );
  NAND U3891 ( .A(n3074), .B(n3073), .Z(n3184) );
  XOR U3892 ( .A(b[13]), .B(n14905), .Z(n3226) );
  OR U3893 ( .A(n3226), .B(n31550), .Z(n3077) );
  NANDN U3894 ( .A(n3075), .B(n31874), .Z(n3076) );
  NAND U3895 ( .A(n3077), .B(n3076), .Z(n3181) );
  NAND U3896 ( .A(n33283), .B(n3078), .Z(n3080) );
  XOR U3897 ( .A(n33020), .B(n13106), .Z(n3258) );
  NANDN U3898 ( .A(n33021), .B(n3258), .Z(n3079) );
  AND U3899 ( .A(n3080), .B(n3079), .Z(n3182) );
  XNOR U3900 ( .A(n3181), .B(n3182), .Z(n3183) );
  XNOR U3901 ( .A(n3184), .B(n3183), .Z(n3280) );
  XOR U3902 ( .A(n970), .B(n15484), .Z(n3241) );
  NANDN U3903 ( .A(n31369), .B(n3241), .Z(n3083) );
  NANDN U3904 ( .A(n3081), .B(n31119), .Z(n3082) );
  NAND U3905 ( .A(n3083), .B(n3082), .Z(n3278) );
  NAND U3906 ( .A(n30846), .B(n3084), .Z(n3086) );
  XNOR U3907 ( .A(n969), .B(a[22]), .Z(n3223) );
  NAND U3908 ( .A(n30509), .B(n3223), .Z(n3085) );
  AND U3909 ( .A(n3086), .B(n3085), .Z(n3277) );
  XNOR U3910 ( .A(n3278), .B(n3277), .Z(n3279) );
  XOR U3911 ( .A(n3280), .B(n3279), .Z(n3215) );
  NAND U3912 ( .A(n3088), .B(n3087), .Z(n3263) );
  XNOR U3913 ( .A(b[17]), .B(a[14]), .Z(n3249) );
  NANDN U3914 ( .A(n3249), .B(n32543), .Z(n3091) );
  NANDN U3915 ( .A(n3089), .B(n32541), .Z(n3090) );
  NAND U3916 ( .A(n3091), .B(n3090), .Z(n3262) );
  XNOR U3917 ( .A(n35375), .B(b[29]), .Z(n3093) );
  AND U3918 ( .A(n3093), .B(n3092), .Z(n35188) );
  NANDN U3919 ( .A(n3094), .B(n35188), .Z(n3096) );
  XNOR U3920 ( .A(n35540), .B(a[2]), .Z(n3187) );
  NANDN U3921 ( .A(n34968), .B(n3187), .Z(n3095) );
  AND U3922 ( .A(n3096), .B(n3095), .Z(n3261) );
  XNOR U3923 ( .A(n3262), .B(n3261), .Z(n3264) );
  XNOR U3924 ( .A(n3263), .B(n3264), .Z(n3213) );
  XOR U3925 ( .A(b[15]), .B(n14259), .Z(n3198) );
  OR U3926 ( .A(n3198), .B(n32010), .Z(n3099) );
  NAND U3927 ( .A(n3097), .B(n32011), .Z(n3098) );
  NAND U3928 ( .A(n3099), .B(n3098), .Z(n3274) );
  XOR U3929 ( .A(b[5]), .B(n17133), .Z(n3255) );
  OR U3930 ( .A(n3255), .B(n29363), .Z(n3102) );
  NANDN U3931 ( .A(n3100), .B(n29864), .Z(n3101) );
  NAND U3932 ( .A(n3102), .B(n3101), .Z(n3271) );
  XOR U3933 ( .A(b[3]), .B(n17702), .Z(n3246) );
  NANDN U3934 ( .A(n3246), .B(n28939), .Z(n3105) );
  NAND U3935 ( .A(n28938), .B(n3103), .Z(n3104) );
  AND U3936 ( .A(n3105), .B(n3104), .Z(n3272) );
  XNOR U3937 ( .A(n3271), .B(n3272), .Z(n3273) );
  XNOR U3938 ( .A(n3274), .B(n3273), .Z(n3214) );
  XOR U3939 ( .A(n3213), .B(n3214), .Z(n3216) );
  XOR U3940 ( .A(n3215), .B(n3216), .Z(n3204) );
  NANDN U3941 ( .A(n3107), .B(n3106), .Z(n3111) );
  NANDN U3942 ( .A(n3109), .B(n3108), .Z(n3110) );
  AND U3943 ( .A(n3111), .B(n3110), .Z(n3201) );
  NANDN U3944 ( .A(n3113), .B(n3112), .Z(n3117) );
  NAND U3945 ( .A(n3115), .B(n3114), .Z(n3116) );
  NAND U3946 ( .A(n3117), .B(n3116), .Z(n3202) );
  XNOR U3947 ( .A(n3204), .B(n3203), .Z(n3284) );
  NANDN U3948 ( .A(n3119), .B(n3118), .Z(n3123) );
  NANDN U3949 ( .A(n3121), .B(n3120), .Z(n3122) );
  AND U3950 ( .A(n3123), .B(n3122), .Z(n3283) );
  XOR U3951 ( .A(n3284), .B(n3283), .Z(n3285) );
  XOR U3952 ( .A(n3286), .B(n3285), .Z(n3290) );
  XNOR U3953 ( .A(n3289), .B(n3290), .Z(n3291) );
  NANDN U3954 ( .A(n3133), .B(n3132), .Z(n3137) );
  NAND U3955 ( .A(n3135), .B(n3134), .Z(n3136) );
  NAND U3956 ( .A(n3137), .B(n3136), .Z(n3222) );
  XOR U3957 ( .A(b[29]), .B(b[30]), .Z(n35313) );
  AND U3958 ( .A(n35313), .B(a[0]), .Z(n3178) );
  NANDN U3959 ( .A(n966), .B(a[30]), .Z(n3138) );
  XOR U3960 ( .A(n29232), .B(n3138), .Z(n3140) );
  IV U3961 ( .A(a[29]), .Z(n18003) );
  NANDN U3962 ( .A(n18003), .B(n966), .Z(n3139) );
  AND U3963 ( .A(n3140), .B(n3139), .Z(n3176) );
  NAND U3964 ( .A(n3141), .B(n34848), .Z(n3143) );
  XNOR U3965 ( .A(n35375), .B(a[4]), .Z(n3232) );
  NAND U3966 ( .A(n34618), .B(n3232), .Z(n3142) );
  AND U3967 ( .A(n3143), .B(n3142), .Z(n3175) );
  XNOR U3968 ( .A(n3176), .B(n3175), .Z(n3177) );
  XOR U3969 ( .A(n3178), .B(n3177), .Z(n3219) );
  XNOR U3970 ( .A(b[21]), .B(a[10]), .Z(n3229) );
  OR U3971 ( .A(n3229), .B(n33634), .Z(n3146) );
  NAND U3972 ( .A(n3144), .B(n33464), .Z(n3145) );
  NAND U3973 ( .A(n3146), .B(n3145), .Z(n3268) );
  NAND U3974 ( .A(n34044), .B(n3147), .Z(n3149) );
  XOR U3975 ( .A(n34510), .B(n11986), .Z(n3235) );
  NANDN U3976 ( .A(n33867), .B(n3235), .Z(n3148) );
  NAND U3977 ( .A(n3149), .B(n3148), .Z(n3265) );
  XNOR U3978 ( .A(b[25]), .B(n11406), .Z(n3238) );
  NANDN U3979 ( .A(n34219), .B(n3238), .Z(n3152) );
  NAND U3980 ( .A(n34217), .B(n3150), .Z(n3151) );
  AND U3981 ( .A(n3152), .B(n3151), .Z(n3266) );
  XNOR U3982 ( .A(n3265), .B(n3266), .Z(n3267) );
  XNOR U3983 ( .A(n3268), .B(n3267), .Z(n3220) );
  XNOR U3984 ( .A(n3219), .B(n3220), .Z(n3221) );
  XNOR U3985 ( .A(n3222), .B(n3221), .Z(n3210) );
  NANDN U3986 ( .A(n3154), .B(n3153), .Z(n3158) );
  NANDN U3987 ( .A(n3156), .B(n3155), .Z(n3157) );
  NAND U3988 ( .A(n3158), .B(n3157), .Z(n3207) );
  OR U3989 ( .A(n3160), .B(n3159), .Z(n3164) );
  NAND U3990 ( .A(n3162), .B(n3161), .Z(n3163) );
  NAND U3991 ( .A(n3164), .B(n3163), .Z(n3208) );
  XNOR U3992 ( .A(n3207), .B(n3208), .Z(n3209) );
  XOR U3993 ( .A(n3210), .B(n3209), .Z(n3295) );
  XNOR U3994 ( .A(n3296), .B(n3295), .Z(n3298) );
  XOR U3995 ( .A(n3297), .B(n3298), .Z(n3292) );
  XNOR U3996 ( .A(n3291), .B(n3292), .Z(n3302) );
  XNOR U3997 ( .A(n3301), .B(n3302), .Z(n3303) );
  XNOR U3998 ( .A(n3303), .B(n3304), .Z(n3170) );
  XNOR U3999 ( .A(n3169), .B(n3170), .Z(n3171) );
  XOR U4000 ( .A(n3172), .B(n3171), .Z(n3308) );
  XOR U4001 ( .A(n3309), .B(n3308), .Z(c[94]) );
  NANDN U4002 ( .A(n3170), .B(n3169), .Z(n3174) );
  NAND U4003 ( .A(n3172), .B(n3171), .Z(n3173) );
  NAND U4004 ( .A(n3174), .B(n3173), .Z(n3320) );
  NANDN U4005 ( .A(n3176), .B(n3175), .Z(n3180) );
  NANDN U4006 ( .A(n3178), .B(n3177), .Z(n3179) );
  NAND U4007 ( .A(n3180), .B(n3179), .Z(n3390) );
  NANDN U4008 ( .A(n3182), .B(n3181), .Z(n3186) );
  NAND U4009 ( .A(n3184), .B(n3183), .Z(n3185) );
  NAND U4010 ( .A(n3186), .B(n3185), .Z(n3391) );
  XNOR U4011 ( .A(n3390), .B(n3391), .Z(n3392) );
  NAND U4012 ( .A(n3187), .B(n35188), .Z(n3189) );
  XOR U4013 ( .A(b[29]), .B(n10524), .Z(n3354) );
  OR U4014 ( .A(n3354), .B(n34968), .Z(n3188) );
  NAND U4015 ( .A(n3189), .B(n3188), .Z(n3418) );
  XOR U4016 ( .A(b[31]), .B(n10457), .Z(n3405) );
  ANDN U4017 ( .B(n35313), .A(n3405), .Z(n3194) );
  XNOR U4018 ( .A(n973), .B(a[0]), .Z(n3192) );
  XNOR U4019 ( .A(n973), .B(b[29]), .Z(n3191) );
  XNOR U4020 ( .A(n973), .B(b[30]), .Z(n3190) );
  AND U4021 ( .A(n3191), .B(n3190), .Z(n35311) );
  NAND U4022 ( .A(n3192), .B(n35311), .Z(n3193) );
  NANDN U4023 ( .A(n3194), .B(n3193), .Z(n3417) );
  XNOR U4024 ( .A(n3418), .B(n3417), .Z(n3381) );
  NANDN U4025 ( .A(n966), .B(a[31]), .Z(n3195) );
  XOR U4026 ( .A(n29232), .B(n3195), .Z(n3197) );
  IV U4027 ( .A(a[30]), .Z(n18804) );
  NANDN U4028 ( .A(n18804), .B(n966), .Z(n3196) );
  AND U4029 ( .A(n3197), .B(n3196), .Z(n3379) );
  NANDN U4030 ( .A(n3198), .B(n32011), .Z(n3200) );
  XNOR U4031 ( .A(n972), .B(a[17]), .Z(n3363) );
  NANDN U4032 ( .A(n32010), .B(n3363), .Z(n3199) );
  AND U4033 ( .A(n3200), .B(n3199), .Z(n3378) );
  XNOR U4034 ( .A(n3379), .B(n3378), .Z(n3380) );
  XOR U4035 ( .A(n3381), .B(n3380), .Z(n3393) );
  XOR U4036 ( .A(n3392), .B(n3393), .Z(n3334) );
  OR U4037 ( .A(n3202), .B(n3201), .Z(n3206) );
  NANDN U4038 ( .A(n3204), .B(n3203), .Z(n3205) );
  NAND U4039 ( .A(n3206), .B(n3205), .Z(n3333) );
  XOR U4040 ( .A(n3334), .B(n3333), .Z(n3335) );
  NANDN U4041 ( .A(n3208), .B(n3207), .Z(n3212) );
  NAND U4042 ( .A(n3210), .B(n3209), .Z(n3211) );
  NAND U4043 ( .A(n3212), .B(n3211), .Z(n3336) );
  XOR U4044 ( .A(n3335), .B(n3336), .Z(n3332) );
  NANDN U4045 ( .A(n3214), .B(n3213), .Z(n3218) );
  OR U4046 ( .A(n3216), .B(n3215), .Z(n3217) );
  NAND U4047 ( .A(n3218), .B(n3217), .Z(n3345) );
  XNOR U4048 ( .A(n3345), .B(n3346), .Z(n3347) );
  XOR U4049 ( .A(b[9]), .B(n16269), .Z(n3402) );
  NANDN U4050 ( .A(n3402), .B(n30509), .Z(n3225) );
  NAND U4051 ( .A(n3223), .B(n30846), .Z(n3224) );
  NAND U4052 ( .A(n3225), .B(n3224), .Z(n3369) );
  XOR U4053 ( .A(b[13]), .B(n15113), .Z(n3357) );
  OR U4054 ( .A(n3357), .B(n31550), .Z(n3228) );
  NANDN U4055 ( .A(n3226), .B(n31874), .Z(n3227) );
  NAND U4056 ( .A(n3228), .B(n3227), .Z(n3366) );
  XNOR U4057 ( .A(b[21]), .B(a[11]), .Z(n3360) );
  OR U4058 ( .A(n3360), .B(n33634), .Z(n3231) );
  NANDN U4059 ( .A(n3229), .B(n33464), .Z(n3230) );
  AND U4060 ( .A(n3231), .B(n3230), .Z(n3367) );
  XNOR U4061 ( .A(n3366), .B(n3367), .Z(n3368) );
  XNOR U4062 ( .A(n3369), .B(n3368), .Z(n3399) );
  NAND U4063 ( .A(n3232), .B(n34848), .Z(n3234) );
  XOR U4064 ( .A(n35375), .B(n11202), .Z(n3431) );
  NAND U4065 ( .A(n34618), .B(n3431), .Z(n3233) );
  NAND U4066 ( .A(n3234), .B(n3233), .Z(n3446) );
  NAND U4067 ( .A(n34044), .B(n3235), .Z(n3237) );
  XOR U4068 ( .A(n34510), .B(n12258), .Z(n3408) );
  NANDN U4069 ( .A(n33867), .B(n3408), .Z(n3236) );
  NAND U4070 ( .A(n3237), .B(n3236), .Z(n3443) );
  XNOR U4071 ( .A(b[25]), .B(n11694), .Z(n3428) );
  NANDN U4072 ( .A(n34219), .B(n3428), .Z(n3240) );
  NAND U4073 ( .A(n34217), .B(n3238), .Z(n3239) );
  AND U4074 ( .A(n3240), .B(n3239), .Z(n3444) );
  XNOR U4075 ( .A(n3443), .B(n3444), .Z(n3445) );
  XNOR U4076 ( .A(n3446), .B(n3445), .Z(n3396) );
  XNOR U4077 ( .A(n970), .B(a[21]), .Z(n3425) );
  NANDN U4078 ( .A(n31369), .B(n3425), .Z(n3243) );
  NAND U4079 ( .A(n31119), .B(n3241), .Z(n3242) );
  NAND U4080 ( .A(n3243), .B(n3242), .Z(n3397) );
  XNOR U4081 ( .A(n3396), .B(n3397), .Z(n3398) );
  XOR U4082 ( .A(n3399), .B(n3398), .Z(n3339) );
  NOR U4083 ( .A(b[29]), .B(b[30]), .Z(n3244) );
  OR U4084 ( .A(n3244), .B(n986), .Z(n3245) );
  NANDN U4085 ( .A(n35540), .B(b[30]), .Z(n35539) );
  AND U4086 ( .A(n35539), .B(b[31]), .Z(n35818) );
  IV U4087 ( .A(n35818), .Z(n35629) );
  ANDN U4088 ( .B(n3245), .A(n35629), .Z(n3373) );
  XNOR U4089 ( .A(n967), .B(a[29]), .Z(n3422) );
  NAND U4090 ( .A(n3422), .B(n28939), .Z(n3248) );
  NANDN U4091 ( .A(n3246), .B(n28938), .Z(n3247) );
  NAND U4092 ( .A(n3248), .B(n3247), .Z(n3372) );
  XOR U4093 ( .A(n3373), .B(n3372), .Z(n3374) );
  XNOR U4094 ( .A(b[17]), .B(a[15]), .Z(n3419) );
  NANDN U4095 ( .A(n3419), .B(n32543), .Z(n3251) );
  NANDN U4096 ( .A(n3249), .B(n32541), .Z(n3250) );
  NAND U4097 ( .A(n3251), .B(n3250), .Z(n3375) );
  XOR U4098 ( .A(n3374), .B(n3375), .Z(n3384) );
  XOR U4099 ( .A(n31123), .B(n16916), .Z(n3437) );
  NAND U4100 ( .A(n3437), .B(n29949), .Z(n3254) );
  NAND U4101 ( .A(n29948), .B(n3252), .Z(n3253) );
  NAND U4102 ( .A(n3254), .B(n3253), .Z(n3414) );
  XOR U4103 ( .A(b[5]), .B(n17960), .Z(n3440) );
  OR U4104 ( .A(n3440), .B(n29363), .Z(n3257) );
  NANDN U4105 ( .A(n3255), .B(n29864), .Z(n3256) );
  NAND U4106 ( .A(n3257), .B(n3256), .Z(n3411) );
  NAND U4107 ( .A(n33283), .B(n3258), .Z(n3260) );
  XOR U4108 ( .A(n33020), .B(n13509), .Z(n3434) );
  NANDN U4109 ( .A(n33021), .B(n3434), .Z(n3259) );
  AND U4110 ( .A(n3260), .B(n3259), .Z(n3412) );
  XNOR U4111 ( .A(n3411), .B(n3412), .Z(n3413) );
  XNOR U4112 ( .A(n3414), .B(n3413), .Z(n3385) );
  XNOR U4113 ( .A(n3384), .B(n3385), .Z(n3386) );
  XNOR U4114 ( .A(n3386), .B(n3387), .Z(n3340) );
  XNOR U4115 ( .A(n3339), .B(n3340), .Z(n3342) );
  NANDN U4116 ( .A(n3266), .B(n3265), .Z(n3270) );
  NAND U4117 ( .A(n3268), .B(n3267), .Z(n3269) );
  NAND U4118 ( .A(n3270), .B(n3269), .Z(n3449) );
  NANDN U4119 ( .A(n3272), .B(n3271), .Z(n3276) );
  NAND U4120 ( .A(n3274), .B(n3273), .Z(n3275) );
  AND U4121 ( .A(n3276), .B(n3275), .Z(n3450) );
  XNOR U4122 ( .A(n3449), .B(n3450), .Z(n3451) );
  NANDN U4123 ( .A(n3278), .B(n3277), .Z(n3282) );
  NAND U4124 ( .A(n3280), .B(n3279), .Z(n3281) );
  NAND U4125 ( .A(n3282), .B(n3281), .Z(n3452) );
  XOR U4126 ( .A(n3451), .B(n3452), .Z(n3341) );
  XOR U4127 ( .A(n3342), .B(n3341), .Z(n3348) );
  XNOR U4128 ( .A(n3347), .B(n3348), .Z(n3329) );
  OR U4129 ( .A(n3284), .B(n3283), .Z(n3288) );
  NAND U4130 ( .A(n3286), .B(n3285), .Z(n3287) );
  NAND U4131 ( .A(n3288), .B(n3287), .Z(n3330) );
  XNOR U4132 ( .A(n3329), .B(n3330), .Z(n3331) );
  XNOR U4133 ( .A(n3332), .B(n3331), .Z(n3326) );
  NANDN U4134 ( .A(n3290), .B(n3289), .Z(n3294) );
  NANDN U4135 ( .A(n3292), .B(n3291), .Z(n3293) );
  NAND U4136 ( .A(n3294), .B(n3293), .Z(n3324) );
  NAND U4137 ( .A(n3296), .B(n3295), .Z(n3300) );
  NANDN U4138 ( .A(n3298), .B(n3297), .Z(n3299) );
  AND U4139 ( .A(n3300), .B(n3299), .Z(n3323) );
  XNOR U4140 ( .A(n3324), .B(n3323), .Z(n3325) );
  XOR U4141 ( .A(n3326), .B(n3325), .Z(n3317) );
  NANDN U4142 ( .A(n3302), .B(n3301), .Z(n3306) );
  NANDN U4143 ( .A(n3304), .B(n3303), .Z(n3305) );
  NAND U4144 ( .A(n3306), .B(n3305), .Z(n3318) );
  XOR U4145 ( .A(n3317), .B(n3318), .Z(n3319) );
  XNOR U4146 ( .A(n3320), .B(n3319), .Z(n3312) );
  XNOR U4147 ( .A(n3312), .B(sreg[95]), .Z(n3314) );
  NAND U4148 ( .A(n3307), .B(sreg[94]), .Z(n3311) );
  OR U4149 ( .A(n3309), .B(n3308), .Z(n3310) );
  AND U4150 ( .A(n3311), .B(n3310), .Z(n3313) );
  XOR U4151 ( .A(n3314), .B(n3313), .Z(c[95]) );
  NAND U4152 ( .A(n3312), .B(sreg[95]), .Z(n3316) );
  OR U4153 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U4154 ( .A(n3316), .B(n3315), .Z(n3602) );
  XNOR U4155 ( .A(n3602), .B(sreg[96]), .Z(n3604) );
  OR U4156 ( .A(n3318), .B(n3317), .Z(n3322) );
  NAND U4157 ( .A(n3320), .B(n3319), .Z(n3321) );
  NAND U4158 ( .A(n3322), .B(n3321), .Z(n3458) );
  NANDN U4159 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U4160 ( .A(n3326), .B(n3325), .Z(n3327) );
  NAND U4161 ( .A(n3328), .B(n3327), .Z(n3456) );
  OR U4162 ( .A(n3334), .B(n3333), .Z(n3338) );
  NANDN U4163 ( .A(n3336), .B(n3335), .Z(n3337) );
  NAND U4164 ( .A(n3338), .B(n3337), .Z(n3462) );
  XNOR U4165 ( .A(n3461), .B(n3462), .Z(n3463) );
  OR U4166 ( .A(n3340), .B(n3339), .Z(n3344) );
  OR U4167 ( .A(n3342), .B(n3341), .Z(n3343) );
  NAND U4168 ( .A(n3344), .B(n3343), .Z(n3470) );
  NANDN U4169 ( .A(n3346), .B(n3345), .Z(n3350) );
  NAND U4170 ( .A(n3348), .B(n3347), .Z(n3349) );
  NAND U4171 ( .A(n3350), .B(n3349), .Z(n3467) );
  XNOR U4172 ( .A(n973), .B(b[32]), .Z(n35620) );
  NAND U4173 ( .A(a[0]), .B(n35620), .Z(n3559) );
  NANDN U4174 ( .A(n966), .B(a[32]), .Z(n3351) );
  XOR U4175 ( .A(n29232), .B(n3351), .Z(n3353) );
  IV U4176 ( .A(a[31]), .Z(n18639) );
  NANDN U4177 ( .A(n18639), .B(n966), .Z(n3352) );
  AND U4178 ( .A(n3353), .B(n3352), .Z(n3557) );
  NANDN U4179 ( .A(n3354), .B(n35188), .Z(n3356) );
  XOR U4180 ( .A(b[29]), .B(n10854), .Z(n3509) );
  OR U4181 ( .A(n3509), .B(n34968), .Z(n3355) );
  AND U4182 ( .A(n3356), .B(n3355), .Z(n3556) );
  XNOR U4183 ( .A(n3557), .B(n3556), .Z(n3558) );
  XOR U4184 ( .A(n3559), .B(n3558), .Z(n3568) );
  XOR U4185 ( .A(b[13]), .B(n15484), .Z(n3495) );
  OR U4186 ( .A(n3495), .B(n31550), .Z(n3359) );
  NANDN U4187 ( .A(n3357), .B(n31874), .Z(n3358) );
  NAND U4188 ( .A(n3359), .B(n3358), .Z(n3518) );
  XNOR U4189 ( .A(b[21]), .B(a[12]), .Z(n3547) );
  OR U4190 ( .A(n3547), .B(n33634), .Z(n3362) );
  NANDN U4191 ( .A(n3360), .B(n33464), .Z(n3361) );
  NAND U4192 ( .A(n3362), .B(n3361), .Z(n3515) );
  XOR U4193 ( .A(b[15]), .B(n14905), .Z(n3498) );
  OR U4194 ( .A(n3498), .B(n32010), .Z(n3365) );
  NAND U4195 ( .A(n3363), .B(n32011), .Z(n3364) );
  AND U4196 ( .A(n3365), .B(n3364), .Z(n3516) );
  XNOR U4197 ( .A(n3515), .B(n3516), .Z(n3517) );
  XNOR U4198 ( .A(n3518), .B(n3517), .Z(n3569) );
  XNOR U4199 ( .A(n3568), .B(n3569), .Z(n3571) );
  NANDN U4200 ( .A(n3367), .B(n3366), .Z(n3371) );
  NAND U4201 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U4202 ( .A(n3371), .B(n3370), .Z(n3570) );
  XNOR U4203 ( .A(n3571), .B(n3570), .Z(n3581) );
  OR U4204 ( .A(n3373), .B(n3372), .Z(n3377) );
  NANDN U4205 ( .A(n3375), .B(n3374), .Z(n3376) );
  NAND U4206 ( .A(n3377), .B(n3376), .Z(n3578) );
  NANDN U4207 ( .A(n3379), .B(n3378), .Z(n3383) );
  NAND U4208 ( .A(n3381), .B(n3380), .Z(n3382) );
  AND U4209 ( .A(n3383), .B(n3382), .Z(n3579) );
  XNOR U4210 ( .A(n3578), .B(n3579), .Z(n3580) );
  XOR U4211 ( .A(n3581), .B(n3580), .Z(n3597) );
  NANDN U4212 ( .A(n3385), .B(n3384), .Z(n3389) );
  NAND U4213 ( .A(n3387), .B(n3386), .Z(n3388) );
  AND U4214 ( .A(n3389), .B(n3388), .Z(n3596) );
  XOR U4215 ( .A(n3597), .B(n3596), .Z(n3598) );
  NANDN U4216 ( .A(n3391), .B(n3390), .Z(n3395) );
  NAND U4217 ( .A(n3393), .B(n3392), .Z(n3394) );
  NAND U4218 ( .A(n3395), .B(n3394), .Z(n3599) );
  XOR U4219 ( .A(n3598), .B(n3599), .Z(n3577) );
  NANDN U4220 ( .A(n3397), .B(n3396), .Z(n3401) );
  NAND U4221 ( .A(n3399), .B(n3398), .Z(n3400) );
  NAND U4222 ( .A(n3401), .B(n3400), .Z(n3476) );
  XOR U4223 ( .A(n969), .B(n16508), .Z(n3486) );
  NAND U4224 ( .A(n30509), .B(n3486), .Z(n3404) );
  NANDN U4225 ( .A(n3402), .B(n30846), .Z(n3403) );
  NAND U4226 ( .A(n3404), .B(n3403), .Z(n3565) );
  XOR U4227 ( .A(b[31]), .B(n10363), .Z(n3533) );
  NANDN U4228 ( .A(n3533), .B(n35313), .Z(n3407) );
  NANDN U4229 ( .A(n3405), .B(n35311), .Z(n3406) );
  NAND U4230 ( .A(n3407), .B(n3406), .Z(n3562) );
  NAND U4231 ( .A(n34044), .B(n3408), .Z(n3410) );
  XOR U4232 ( .A(n34510), .B(n12555), .Z(n3550) );
  NANDN U4233 ( .A(n33867), .B(n3550), .Z(n3409) );
  AND U4234 ( .A(n3410), .B(n3409), .Z(n3563) );
  XNOR U4235 ( .A(n3562), .B(n3563), .Z(n3564) );
  XNOR U4236 ( .A(n3565), .B(n3564), .Z(n3584) );
  NANDN U4237 ( .A(n3412), .B(n3411), .Z(n3416) );
  NAND U4238 ( .A(n3414), .B(n3413), .Z(n3415) );
  NAND U4239 ( .A(n3416), .B(n3415), .Z(n3585) );
  XNOR U4240 ( .A(n3584), .B(n3585), .Z(n3586) );
  NAND U4241 ( .A(n3418), .B(n3417), .Z(n3481) );
  XNOR U4242 ( .A(b[17]), .B(a[16]), .Z(n3544) );
  NANDN U4243 ( .A(n3544), .B(n32543), .Z(n3421) );
  NANDN U4244 ( .A(n3419), .B(n32541), .Z(n3420) );
  NAND U4245 ( .A(n3421), .B(n3420), .Z(n3480) );
  XOR U4246 ( .A(n967), .B(n18804), .Z(n3504) );
  NAND U4247 ( .A(n3504), .B(n28939), .Z(n3424) );
  NAND U4248 ( .A(n3422), .B(n28938), .Z(n3423) );
  AND U4249 ( .A(n3424), .B(n3423), .Z(n3479) );
  XNOR U4250 ( .A(n3480), .B(n3479), .Z(n3482) );
  XNOR U4251 ( .A(n3481), .B(n3482), .Z(n3587) );
  XNOR U4252 ( .A(n3586), .B(n3587), .Z(n3473) );
  XOR U4253 ( .A(b[11]), .B(n15963), .Z(n3492) );
  OR U4254 ( .A(n3492), .B(n31369), .Z(n3427) );
  NAND U4255 ( .A(n3425), .B(n31119), .Z(n3426) );
  NAND U4256 ( .A(n3427), .B(n3426), .Z(n3524) );
  XNOR U4257 ( .A(b[25]), .B(n11986), .Z(n3553) );
  NANDN U4258 ( .A(n34219), .B(n3553), .Z(n3430) );
  NAND U4259 ( .A(n34217), .B(n3428), .Z(n3429) );
  NAND U4260 ( .A(n3430), .B(n3429), .Z(n3521) );
  NAND U4261 ( .A(n34848), .B(n3431), .Z(n3433) );
  XOR U4262 ( .A(n35375), .B(n11406), .Z(n3501) );
  NAND U4263 ( .A(n34618), .B(n3501), .Z(n3432) );
  AND U4264 ( .A(n3433), .B(n3432), .Z(n3522) );
  XNOR U4265 ( .A(n3521), .B(n3522), .Z(n3523) );
  XNOR U4266 ( .A(n3524), .B(n3523), .Z(n3590) );
  NAND U4267 ( .A(n33283), .B(n3434), .Z(n3436) );
  XOR U4268 ( .A(n33020), .B(n14210), .Z(n3512) );
  NANDN U4269 ( .A(n33021), .B(n3512), .Z(n3435) );
  NAND U4270 ( .A(n3436), .B(n3435), .Z(n3530) );
  XNOR U4271 ( .A(n31123), .B(a[26]), .Z(n3483) );
  NAND U4272 ( .A(n3483), .B(n29949), .Z(n3439) );
  NAND U4273 ( .A(n29948), .B(n3437), .Z(n3438) );
  NAND U4274 ( .A(n3439), .B(n3438), .Z(n3527) );
  XOR U4275 ( .A(b[5]), .B(n17702), .Z(n3489) );
  OR U4276 ( .A(n3489), .B(n29363), .Z(n3442) );
  NANDN U4277 ( .A(n3440), .B(n29864), .Z(n3441) );
  AND U4278 ( .A(n3442), .B(n3441), .Z(n3528) );
  XNOR U4279 ( .A(n3527), .B(n3528), .Z(n3529) );
  XOR U4280 ( .A(n3530), .B(n3529), .Z(n3591) );
  XOR U4281 ( .A(n3590), .B(n3591), .Z(n3593) );
  NANDN U4282 ( .A(n3444), .B(n3443), .Z(n3448) );
  NAND U4283 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U4284 ( .A(n3448), .B(n3447), .Z(n3592) );
  XOR U4285 ( .A(n3593), .B(n3592), .Z(n3474) );
  XNOR U4286 ( .A(n3473), .B(n3474), .Z(n3475) );
  XNOR U4287 ( .A(n3476), .B(n3475), .Z(n3574) );
  NANDN U4288 ( .A(n3450), .B(n3449), .Z(n3454) );
  NANDN U4289 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U4290 ( .A(n3454), .B(n3453), .Z(n3575) );
  XNOR U4291 ( .A(n3574), .B(n3575), .Z(n3576) );
  XNOR U4292 ( .A(n3577), .B(n3576), .Z(n3468) );
  XOR U4293 ( .A(n3467), .B(n3468), .Z(n3469) );
  XOR U4294 ( .A(n3470), .B(n3469), .Z(n3464) );
  XNOR U4295 ( .A(n3463), .B(n3464), .Z(n3455) );
  XNOR U4296 ( .A(n3456), .B(n3455), .Z(n3457) );
  XOR U4297 ( .A(n3458), .B(n3457), .Z(n3603) );
  XOR U4298 ( .A(n3604), .B(n3603), .Z(c[96]) );
  NANDN U4299 ( .A(n3456), .B(n3455), .Z(n3460) );
  NAND U4300 ( .A(n3458), .B(n3457), .Z(n3459) );
  NAND U4301 ( .A(n3460), .B(n3459), .Z(n3615) );
  NANDN U4302 ( .A(n3462), .B(n3461), .Z(n3466) );
  NANDN U4303 ( .A(n3464), .B(n3463), .Z(n3465) );
  NAND U4304 ( .A(n3466), .B(n3465), .Z(n3612) );
  OR U4305 ( .A(n3468), .B(n3467), .Z(n3472) );
  NANDN U4306 ( .A(n3470), .B(n3469), .Z(n3471) );
  NAND U4307 ( .A(n3472), .B(n3471), .Z(n3621) );
  OR U4308 ( .A(n3474), .B(n3473), .Z(n3478) );
  OR U4309 ( .A(n3476), .B(n3475), .Z(n3477) );
  NAND U4310 ( .A(n3478), .B(n3477), .Z(n3758) );
  XNOR U4311 ( .A(n31123), .B(a[27]), .Z(n3678) );
  NAND U4312 ( .A(n3678), .B(n29949), .Z(n3485) );
  NAND U4313 ( .A(n3483), .B(n29948), .Z(n3484) );
  AND U4314 ( .A(n3485), .B(n3484), .Z(n3696) );
  NAND U4315 ( .A(n30846), .B(n3486), .Z(n3488) );
  XNOR U4316 ( .A(n969), .B(a[25]), .Z(n3651) );
  NAND U4317 ( .A(n30509), .B(n3651), .Z(n3487) );
  AND U4318 ( .A(n3488), .B(n3487), .Z(n3694) );
  XOR U4319 ( .A(b[5]), .B(n18003), .Z(n3672) );
  OR U4320 ( .A(n3672), .B(n29363), .Z(n3491) );
  NANDN U4321 ( .A(n3489), .B(n29864), .Z(n3490) );
  NAND U4322 ( .A(n3491), .B(n3490), .Z(n3722) );
  XOR U4323 ( .A(b[11]), .B(n16269), .Z(n3642) );
  OR U4324 ( .A(n3642), .B(n31369), .Z(n3494) );
  NANDN U4325 ( .A(n3492), .B(n31119), .Z(n3493) );
  NAND U4326 ( .A(n3494), .B(n3493), .Z(n3719) );
  XOR U4327 ( .A(b[13]), .B(n16220), .Z(n3645) );
  OR U4328 ( .A(n3645), .B(n31550), .Z(n3497) );
  NANDN U4329 ( .A(n3495), .B(n31874), .Z(n3496) );
  AND U4330 ( .A(n3497), .B(n3496), .Z(n3720) );
  XNOR U4331 ( .A(n3719), .B(n3720), .Z(n3721) );
  XOR U4332 ( .A(n3722), .B(n3721), .Z(n3693) );
  XNOR U4333 ( .A(n3694), .B(n3693), .Z(n3695) );
  XNOR U4334 ( .A(n3696), .B(n3695), .Z(n3633) );
  XOR U4335 ( .A(b[15]), .B(n15113), .Z(n3660) );
  OR U4336 ( .A(n3660), .B(n32010), .Z(n3500) );
  NANDN U4337 ( .A(n3498), .B(n32011), .Z(n3499) );
  NAND U4338 ( .A(n3500), .B(n3499), .Z(n3728) );
  NAND U4339 ( .A(n34848), .B(n3501), .Z(n3503) );
  XOR U4340 ( .A(n35375), .B(n11694), .Z(n3657) );
  NAND U4341 ( .A(n34618), .B(n3657), .Z(n3502) );
  NAND U4342 ( .A(n3503), .B(n3502), .Z(n3725) );
  XOR U4343 ( .A(b[3]), .B(n18639), .Z(n3710) );
  NANDN U4344 ( .A(n3710), .B(n28939), .Z(n3506) );
  NAND U4345 ( .A(n28938), .B(n3504), .Z(n3505) );
  AND U4346 ( .A(n3506), .B(n3505), .Z(n3726) );
  XNOR U4347 ( .A(n3725), .B(n3726), .Z(n3727) );
  XNOR U4348 ( .A(n3728), .B(n3727), .Z(n3631) );
  NOR U4349 ( .A(b[31]), .B(b[32]), .Z(n3507) );
  OR U4350 ( .A(n3507), .B(n986), .Z(n3508) );
  NANDN U4351 ( .A(n973), .B(b[32]), .Z(n35778) );
  AND U4352 ( .A(n35778), .B(b[33]), .Z(n36130) );
  AND U4353 ( .A(n3508), .B(n36130), .Z(n3663) );
  NANDN U4354 ( .A(n3509), .B(n35188), .Z(n3511) );
  XNOR U4355 ( .A(n35540), .B(a[5]), .Z(n3681) );
  NANDN U4356 ( .A(n34968), .B(n3681), .Z(n3510) );
  NAND U4357 ( .A(n3511), .B(n3510), .Z(n3664) );
  XNOR U4358 ( .A(n3663), .B(n3664), .Z(n3666) );
  NAND U4359 ( .A(n3512), .B(n33283), .Z(n3514) );
  XOR U4360 ( .A(b[19]), .B(n13976), .Z(n3707) );
  OR U4361 ( .A(n3707), .B(n33021), .Z(n3513) );
  NAND U4362 ( .A(n3514), .B(n3513), .Z(n3665) );
  XOR U4363 ( .A(n3666), .B(n3665), .Z(n3630) );
  XOR U4364 ( .A(n3631), .B(n3630), .Z(n3632) );
  XNOR U4365 ( .A(n3633), .B(n3632), .Z(n3739) );
  NANDN U4366 ( .A(n3516), .B(n3515), .Z(n3520) );
  NAND U4367 ( .A(n3518), .B(n3517), .Z(n3519) );
  NAND U4368 ( .A(n3520), .B(n3519), .Z(n3738) );
  NANDN U4369 ( .A(n3522), .B(n3521), .Z(n3526) );
  NAND U4370 ( .A(n3524), .B(n3523), .Z(n3525) );
  AND U4371 ( .A(n3526), .B(n3525), .Z(n3737) );
  XNOR U4372 ( .A(n3738), .B(n3737), .Z(n3740) );
  XOR U4373 ( .A(n3739), .B(n3740), .Z(n3624) );
  XNOR U4374 ( .A(n3625), .B(n3624), .Z(n3627) );
  NANDN U4375 ( .A(n3528), .B(n3527), .Z(n3532) );
  NAND U4376 ( .A(n3530), .B(n3529), .Z(n3531) );
  NAND U4377 ( .A(n3532), .B(n3531), .Z(n3639) );
  XNOR U4378 ( .A(n973), .B(a[3]), .Z(n3716) );
  NAND U4379 ( .A(n3716), .B(n35313), .Z(n3535) );
  NANDN U4380 ( .A(n3533), .B(n35311), .Z(n3534) );
  NAND U4381 ( .A(n3535), .B(n3534), .Z(n3706) );
  XNOR U4382 ( .A(n974), .B(a[0]), .Z(n3538) );
  XNOR U4383 ( .A(n974), .B(b[31]), .Z(n3537) );
  XNOR U4384 ( .A(n974), .B(b[32]), .Z(n3536) );
  AND U4385 ( .A(n3537), .B(n3536), .Z(n35621) );
  NAND U4386 ( .A(n3538), .B(n35621), .Z(n3540) );
  XOR U4387 ( .A(b[33]), .B(n10457), .Z(n3675) );
  NANDN U4388 ( .A(n3675), .B(n35620), .Z(n3539) );
  NAND U4389 ( .A(n3540), .B(n3539), .Z(n3705) );
  XNOR U4390 ( .A(n3706), .B(n3705), .Z(n3734) );
  NANDN U4391 ( .A(n966), .B(a[33]), .Z(n3541) );
  XOR U4392 ( .A(n29232), .B(n3541), .Z(n3543) );
  IV U4393 ( .A(a[32]), .Z(n18841) );
  NANDN U4394 ( .A(n18841), .B(n966), .Z(n3542) );
  AND U4395 ( .A(n3543), .B(n3542), .Z(n3732) );
  XNOR U4396 ( .A(b[17]), .B(n14514), .Z(n3684) );
  NAND U4397 ( .A(n3684), .B(n32543), .Z(n3546) );
  NANDN U4398 ( .A(n3544), .B(n32541), .Z(n3545) );
  AND U4399 ( .A(n3546), .B(n3545), .Z(n3731) );
  XNOR U4400 ( .A(n3732), .B(n3731), .Z(n3733) );
  XOR U4401 ( .A(n3734), .B(n3733), .Z(n3636) );
  XNOR U4402 ( .A(b[21]), .B(a[13]), .Z(n3669) );
  OR U4403 ( .A(n3669), .B(n33634), .Z(n3549) );
  NANDN U4404 ( .A(n3547), .B(n33464), .Z(n3548) );
  NAND U4405 ( .A(n3549), .B(n3548), .Z(n3690) );
  NAND U4406 ( .A(n34044), .B(n3550), .Z(n3552) );
  XOR U4407 ( .A(n34510), .B(n12830), .Z(n3648) );
  NANDN U4408 ( .A(n33867), .B(n3648), .Z(n3551) );
  NAND U4409 ( .A(n3552), .B(n3551), .Z(n3687) );
  XNOR U4410 ( .A(b[25]), .B(n12258), .Z(n3654) );
  NANDN U4411 ( .A(n34219), .B(n3654), .Z(n3555) );
  NAND U4412 ( .A(n34217), .B(n3553), .Z(n3554) );
  AND U4413 ( .A(n3555), .B(n3554), .Z(n3688) );
  XNOR U4414 ( .A(n3687), .B(n3688), .Z(n3689) );
  XNOR U4415 ( .A(n3690), .B(n3689), .Z(n3637) );
  XOR U4416 ( .A(n3636), .B(n3637), .Z(n3638) );
  XNOR U4417 ( .A(n3639), .B(n3638), .Z(n3746) );
  NANDN U4418 ( .A(n3557), .B(n3556), .Z(n3561) );
  NAND U4419 ( .A(n3559), .B(n3558), .Z(n3560) );
  NAND U4420 ( .A(n3561), .B(n3560), .Z(n3743) );
  NANDN U4421 ( .A(n3563), .B(n3562), .Z(n3567) );
  NAND U4422 ( .A(n3565), .B(n3564), .Z(n3566) );
  NAND U4423 ( .A(n3567), .B(n3566), .Z(n3744) );
  XNOR U4424 ( .A(n3743), .B(n3744), .Z(n3745) );
  XOR U4425 ( .A(n3746), .B(n3745), .Z(n3626) );
  XOR U4426 ( .A(n3627), .B(n3626), .Z(n3755) );
  OR U4427 ( .A(n3569), .B(n3568), .Z(n3573) );
  OR U4428 ( .A(n3571), .B(n3570), .Z(n3572) );
  AND U4429 ( .A(n3573), .B(n3572), .Z(n3756) );
  XNOR U4430 ( .A(n3755), .B(n3756), .Z(n3757) );
  XNOR U4431 ( .A(n3758), .B(n3757), .Z(n3618) );
  NANDN U4432 ( .A(n3579), .B(n3578), .Z(n3583) );
  NAND U4433 ( .A(n3581), .B(n3580), .Z(n3582) );
  NAND U4434 ( .A(n3583), .B(n3582), .Z(n3702) );
  NANDN U4435 ( .A(n3585), .B(n3584), .Z(n3589) );
  NANDN U4436 ( .A(n3587), .B(n3586), .Z(n3588) );
  NAND U4437 ( .A(n3589), .B(n3588), .Z(n3699) );
  NANDN U4438 ( .A(n3591), .B(n3590), .Z(n3595) );
  OR U4439 ( .A(n3593), .B(n3592), .Z(n3594) );
  AND U4440 ( .A(n3595), .B(n3594), .Z(n3700) );
  XNOR U4441 ( .A(n3699), .B(n3700), .Z(n3701) );
  XNOR U4442 ( .A(n3702), .B(n3701), .Z(n3749) );
  OR U4443 ( .A(n3597), .B(n3596), .Z(n3601) );
  NANDN U4444 ( .A(n3599), .B(n3598), .Z(n3600) );
  AND U4445 ( .A(n3601), .B(n3600), .Z(n3750) );
  XOR U4446 ( .A(n3749), .B(n3750), .Z(n3752) );
  XOR U4447 ( .A(n3751), .B(n3752), .Z(n3619) );
  XNOR U4448 ( .A(n3618), .B(n3619), .Z(n3620) );
  XNOR U4449 ( .A(n3621), .B(n3620), .Z(n3613) );
  XNOR U4450 ( .A(n3612), .B(n3613), .Z(n3614) );
  XNOR U4451 ( .A(n3615), .B(n3614), .Z(n3607) );
  XNOR U4452 ( .A(n3607), .B(sreg[97]), .Z(n3609) );
  NAND U4453 ( .A(n3602), .B(sreg[96]), .Z(n3606) );
  OR U4454 ( .A(n3604), .B(n3603), .Z(n3605) );
  AND U4455 ( .A(n3606), .B(n3605), .Z(n3608) );
  XOR U4456 ( .A(n3609), .B(n3608), .Z(c[97]) );
  NAND U4457 ( .A(n3607), .B(sreg[97]), .Z(n3611) );
  OR U4458 ( .A(n3609), .B(n3608), .Z(n3610) );
  NAND U4459 ( .A(n3611), .B(n3610), .Z(n3916) );
  XNOR U4460 ( .A(n3916), .B(sreg[98]), .Z(n3918) );
  NANDN U4461 ( .A(n3613), .B(n3612), .Z(n3617) );
  NAND U4462 ( .A(n3615), .B(n3614), .Z(n3616) );
  NAND U4463 ( .A(n3617), .B(n3616), .Z(n3764) );
  NANDN U4464 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U4465 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U4466 ( .A(n3623), .B(n3622), .Z(n3761) );
  NAND U4467 ( .A(n3625), .B(n3624), .Z(n3629) );
  NANDN U4468 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U4469 ( .A(n3629), .B(n3628), .Z(n3775) );
  NAND U4470 ( .A(n3631), .B(n3630), .Z(n3635) );
  NANDN U4471 ( .A(n3633), .B(n3632), .Z(n3634) );
  NAND U4472 ( .A(n3635), .B(n3634), .Z(n3786) );
  OR U4473 ( .A(n3637), .B(n3636), .Z(n3641) );
  NAND U4474 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U4475 ( .A(n3641), .B(n3640), .Z(n3783) );
  XOR U4476 ( .A(b[11]), .B(n16508), .Z(n3813) );
  OR U4477 ( .A(n3813), .B(n31369), .Z(n3644) );
  NANDN U4478 ( .A(n3642), .B(n31119), .Z(n3643) );
  NAND U4479 ( .A(n3644), .B(n3643), .Z(n3895) );
  XOR U4480 ( .A(b[13]), .B(n15963), .Z(n3819) );
  OR U4481 ( .A(n3819), .B(n31550), .Z(n3647) );
  NANDN U4482 ( .A(n3645), .B(n31874), .Z(n3646) );
  NAND U4483 ( .A(n3647), .B(n3646), .Z(n3892) );
  NAND U4484 ( .A(n34044), .B(n3648), .Z(n3650) );
  XOR U4485 ( .A(n34510), .B(n13106), .Z(n3850) );
  NANDN U4486 ( .A(n33867), .B(n3850), .Z(n3649) );
  AND U4487 ( .A(n3650), .B(n3649), .Z(n3893) );
  XNOR U4488 ( .A(n3892), .B(n3893), .Z(n3894) );
  XNOR U4489 ( .A(n3895), .B(n3894), .Z(n3798) );
  XOR U4490 ( .A(b[9]), .B(n17133), .Z(n3859) );
  NANDN U4491 ( .A(n3859), .B(n30509), .Z(n3653) );
  NAND U4492 ( .A(n3651), .B(n30846), .Z(n3652) );
  NAND U4493 ( .A(n3653), .B(n3652), .Z(n3865) );
  XNOR U4494 ( .A(b[25]), .B(n12555), .Z(n3853) );
  NANDN U4495 ( .A(n34219), .B(n3853), .Z(n3656) );
  NAND U4496 ( .A(n34217), .B(n3654), .Z(n3655) );
  NAND U4497 ( .A(n3656), .B(n3655), .Z(n3862) );
  NAND U4498 ( .A(n34848), .B(n3657), .Z(n3659) );
  XOR U4499 ( .A(n35375), .B(n11986), .Z(n3856) );
  NAND U4500 ( .A(n34618), .B(n3856), .Z(n3658) );
  AND U4501 ( .A(n3659), .B(n3658), .Z(n3863) );
  XNOR U4502 ( .A(n3862), .B(n3863), .Z(n3864) );
  XNOR U4503 ( .A(n3865), .B(n3864), .Z(n3795) );
  NANDN U4504 ( .A(n3660), .B(n32011), .Z(n3662) );
  XNOR U4505 ( .A(n972), .B(a[20]), .Z(n3816) );
  NANDN U4506 ( .A(n32010), .B(n3816), .Z(n3661) );
  NAND U4507 ( .A(n3662), .B(n3661), .Z(n3796) );
  XNOR U4508 ( .A(n3795), .B(n3796), .Z(n3797) );
  XOR U4509 ( .A(n3798), .B(n3797), .Z(n3784) );
  XNOR U4510 ( .A(n3783), .B(n3784), .Z(n3785) );
  XOR U4511 ( .A(n3786), .B(n3785), .Z(n3774) );
  OR U4512 ( .A(n3664), .B(n3663), .Z(n3668) );
  OR U4513 ( .A(n3666), .B(n3665), .Z(n3667) );
  NAND U4514 ( .A(n3668), .B(n3667), .Z(n3905) );
  XNOR U4515 ( .A(b[21]), .B(a[14]), .Z(n3874) );
  OR U4516 ( .A(n3874), .B(n33634), .Z(n3671) );
  NANDN U4517 ( .A(n3669), .B(n33464), .Z(n3670) );
  NAND U4518 ( .A(n3671), .B(n3670), .Z(n3871) );
  XOR U4519 ( .A(b[5]), .B(n18804), .Z(n3877) );
  OR U4520 ( .A(n3877), .B(n29363), .Z(n3674) );
  NANDN U4521 ( .A(n3672), .B(n29864), .Z(n3673) );
  NAND U4522 ( .A(n3674), .B(n3673), .Z(n3868) );
  XOR U4523 ( .A(b[33]), .B(n10363), .Z(n3801) );
  NANDN U4524 ( .A(n3801), .B(n35620), .Z(n3677) );
  NANDN U4525 ( .A(n3675), .B(n35621), .Z(n3676) );
  AND U4526 ( .A(n3677), .B(n3676), .Z(n3869) );
  XNOR U4527 ( .A(n3868), .B(n3869), .Z(n3870) );
  XNOR U4528 ( .A(n3871), .B(n3870), .Z(n3843) );
  XOR U4529 ( .A(n31123), .B(n17702), .Z(n3847) );
  NAND U4530 ( .A(n3847), .B(n29949), .Z(n3680) );
  NAND U4531 ( .A(n3678), .B(n29948), .Z(n3679) );
  NAND U4532 ( .A(n3680), .B(n3679), .Z(n3837) );
  NAND U4533 ( .A(n3681), .B(n35188), .Z(n3683) );
  XOR U4534 ( .A(b[29]), .B(n11406), .Z(n3844) );
  OR U4535 ( .A(n3844), .B(n34968), .Z(n3682) );
  NAND U4536 ( .A(n3683), .B(n3682), .Z(n3834) );
  XNOR U4537 ( .A(b[17]), .B(a[18]), .Z(n3886) );
  NANDN U4538 ( .A(n3886), .B(n32543), .Z(n3686) );
  NAND U4539 ( .A(n3684), .B(n32541), .Z(n3685) );
  AND U4540 ( .A(n3686), .B(n3685), .Z(n3835) );
  XNOR U4541 ( .A(n3834), .B(n3835), .Z(n3836) );
  XNOR U4542 ( .A(n3837), .B(n3836), .Z(n3840) );
  NANDN U4543 ( .A(n3688), .B(n3687), .Z(n3692) );
  NAND U4544 ( .A(n3690), .B(n3689), .Z(n3691) );
  NAND U4545 ( .A(n3692), .B(n3691), .Z(n3841) );
  XNOR U4546 ( .A(n3840), .B(n3841), .Z(n3842) );
  XOR U4547 ( .A(n3843), .B(n3842), .Z(n3904) );
  XNOR U4548 ( .A(n3905), .B(n3904), .Z(n3907) );
  NANDN U4549 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U4550 ( .A(n3696), .B(n3695), .Z(n3697) );
  NAND U4551 ( .A(n3698), .B(n3697), .Z(n3906) );
  XOR U4552 ( .A(n3907), .B(n3906), .Z(n3773) );
  XOR U4553 ( .A(n3774), .B(n3773), .Z(n3776) );
  XOR U4554 ( .A(n3775), .B(n3776), .Z(n3780) );
  NANDN U4555 ( .A(n3700), .B(n3699), .Z(n3704) );
  NAND U4556 ( .A(n3702), .B(n3701), .Z(n3703) );
  NAND U4557 ( .A(n3704), .B(n3703), .Z(n3778) );
  NAND U4558 ( .A(n3706), .B(n3705), .Z(n3825) );
  NANDN U4559 ( .A(n3707), .B(n33283), .Z(n3709) );
  XOR U4560 ( .A(b[19]), .B(n14259), .Z(n3810) );
  OR U4561 ( .A(n3810), .B(n33021), .Z(n3708) );
  NAND U4562 ( .A(n3709), .B(n3708), .Z(n3823) );
  XNOR U4563 ( .A(n967), .B(a[32]), .Z(n3880) );
  NAND U4564 ( .A(n3880), .B(n28939), .Z(n3712) );
  NANDN U4565 ( .A(n3710), .B(n28938), .Z(n3711) );
  AND U4566 ( .A(n3712), .B(n3711), .Z(n3822) );
  XNOR U4567 ( .A(n3823), .B(n3822), .Z(n3824) );
  XNOR U4568 ( .A(n3825), .B(n3824), .Z(n3899) );
  XNOR U4569 ( .A(n974), .B(b[34]), .Z(n35985) );
  NAND U4570 ( .A(a[0]), .B(n35985), .Z(n3831) );
  NANDN U4571 ( .A(n966), .B(a[34]), .Z(n3713) );
  XOR U4572 ( .A(n29232), .B(n3713), .Z(n3715) );
  IV U4573 ( .A(a[33]), .Z(n19656) );
  NANDN U4574 ( .A(n19656), .B(n966), .Z(n3714) );
  AND U4575 ( .A(n3715), .B(n3714), .Z(n3829) );
  NAND U4576 ( .A(n3716), .B(n35311), .Z(n3718) );
  XNOR U4577 ( .A(n973), .B(a[4]), .Z(n3883) );
  NAND U4578 ( .A(n3883), .B(n35313), .Z(n3717) );
  AND U4579 ( .A(n3718), .B(n3717), .Z(n3828) );
  XNOR U4580 ( .A(n3829), .B(n3828), .Z(n3830) );
  XNOR U4581 ( .A(n3831), .B(n3830), .Z(n3898) );
  XNOR U4582 ( .A(n3899), .B(n3898), .Z(n3901) );
  NANDN U4583 ( .A(n3720), .B(n3719), .Z(n3724) );
  NAND U4584 ( .A(n3722), .B(n3721), .Z(n3723) );
  NAND U4585 ( .A(n3724), .B(n3723), .Z(n3900) );
  XNOR U4586 ( .A(n3901), .B(n3900), .Z(n3792) );
  NANDN U4587 ( .A(n3726), .B(n3725), .Z(n3730) );
  NAND U4588 ( .A(n3728), .B(n3727), .Z(n3729) );
  NAND U4589 ( .A(n3730), .B(n3729), .Z(n3789) );
  NANDN U4590 ( .A(n3732), .B(n3731), .Z(n3736) );
  NAND U4591 ( .A(n3734), .B(n3733), .Z(n3735) );
  NAND U4592 ( .A(n3736), .B(n3735), .Z(n3790) );
  XNOR U4593 ( .A(n3789), .B(n3790), .Z(n3791) );
  XOR U4594 ( .A(n3792), .B(n3791), .Z(n3910) );
  NANDN U4595 ( .A(n3738), .B(n3737), .Z(n3742) );
  NAND U4596 ( .A(n3740), .B(n3739), .Z(n3741) );
  AND U4597 ( .A(n3742), .B(n3741), .Z(n3911) );
  XNOR U4598 ( .A(n3910), .B(n3911), .Z(n3913) );
  NANDN U4599 ( .A(n3744), .B(n3743), .Z(n3748) );
  NAND U4600 ( .A(n3746), .B(n3745), .Z(n3747) );
  AND U4601 ( .A(n3748), .B(n3747), .Z(n3912) );
  XNOR U4602 ( .A(n3913), .B(n3912), .Z(n3777) );
  XNOR U4603 ( .A(n3778), .B(n3777), .Z(n3779) );
  XNOR U4604 ( .A(n3780), .B(n3779), .Z(n3770) );
  NANDN U4605 ( .A(n3750), .B(n3749), .Z(n3754) );
  OR U4606 ( .A(n3752), .B(n3751), .Z(n3753) );
  NAND U4607 ( .A(n3754), .B(n3753), .Z(n3768) );
  NANDN U4608 ( .A(n3756), .B(n3755), .Z(n3760) );
  NAND U4609 ( .A(n3758), .B(n3757), .Z(n3759) );
  AND U4610 ( .A(n3760), .B(n3759), .Z(n3767) );
  XNOR U4611 ( .A(n3768), .B(n3767), .Z(n3769) );
  XOR U4612 ( .A(n3770), .B(n3769), .Z(n3762) );
  XNOR U4613 ( .A(n3761), .B(n3762), .Z(n3763) );
  XOR U4614 ( .A(n3764), .B(n3763), .Z(n3917) );
  XOR U4615 ( .A(n3918), .B(n3917), .Z(c[98]) );
  NANDN U4616 ( .A(n3762), .B(n3761), .Z(n3766) );
  NAND U4617 ( .A(n3764), .B(n3763), .Z(n3765) );
  NAND U4618 ( .A(n3766), .B(n3765), .Z(n3929) );
  NANDN U4619 ( .A(n3768), .B(n3767), .Z(n3772) );
  NANDN U4620 ( .A(n3770), .B(n3769), .Z(n3771) );
  NAND U4621 ( .A(n3772), .B(n3771), .Z(n3927) );
  NANDN U4622 ( .A(n3778), .B(n3777), .Z(n3782) );
  NANDN U4623 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4624 ( .A(n3782), .B(n3781), .Z(n3933) );
  XNOR U4625 ( .A(n3932), .B(n3933), .Z(n3934) );
  NANDN U4626 ( .A(n3784), .B(n3783), .Z(n3788) );
  NANDN U4627 ( .A(n3786), .B(n3785), .Z(n3787) );
  NAND U4628 ( .A(n3788), .B(n3787), .Z(n4081) );
  NANDN U4629 ( .A(n3790), .B(n3789), .Z(n3794) );
  NAND U4630 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U4631 ( .A(n3794), .B(n3793), .Z(n4069) );
  NANDN U4632 ( .A(n3796), .B(n3795), .Z(n3800) );
  NAND U4633 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U4634 ( .A(n3800), .B(n3799), .Z(n4066) );
  XOR U4635 ( .A(n974), .B(n10524), .Z(n3971) );
  NAND U4636 ( .A(n35620), .B(n3971), .Z(n3803) );
  NANDN U4637 ( .A(n3801), .B(n35621), .Z(n3802) );
  NAND U4638 ( .A(n3803), .B(n3802), .Z(n4008) );
  XNOR U4639 ( .A(b[35]), .B(n10457), .Z(n4042) );
  NAND U4640 ( .A(n35985), .B(n4042), .Z(n3807) );
  XNOR U4641 ( .A(b[35]), .B(n986), .Z(n4110) );
  XNOR U4642 ( .A(b[35]), .B(n974), .Z(n3805) );
  XOR U4643 ( .A(b[35]), .B(b[34]), .Z(n3804) );
  AND U4644 ( .A(n3805), .B(n3804), .Z(n35986) );
  NAND U4645 ( .A(n4110), .B(n35986), .Z(n3806) );
  NAND U4646 ( .A(n3807), .B(n3806), .Z(n4007) );
  XNOR U4647 ( .A(n4008), .B(n4007), .Z(n4033) );
  NANDN U4648 ( .A(n974), .B(b[34]), .Z(n36104) );
  NAND U4649 ( .A(n36104), .B(b[35]), .Z(n36383) );
  NOR U4650 ( .A(b[33]), .B(b[34]), .Z(n3808) );
  OR U4651 ( .A(n3808), .B(n986), .Z(n3809) );
  NANDN U4652 ( .A(n36383), .B(n3809), .Z(n4030) );
  NANDN U4653 ( .A(n3810), .B(n33283), .Z(n3812) );
  XNOR U4654 ( .A(n33020), .B(a[17]), .Z(n4015) );
  NANDN U4655 ( .A(n33021), .B(n4015), .Z(n3811) );
  NAND U4656 ( .A(n3812), .B(n3811), .Z(n4031) );
  XNOR U4657 ( .A(n4030), .B(n4031), .Z(n4032) );
  XOR U4658 ( .A(n4033), .B(n4032), .Z(n3983) );
  XOR U4659 ( .A(b[11]), .B(n16916), .Z(n4054) );
  OR U4660 ( .A(n4054), .B(n31369), .Z(n3815) );
  NANDN U4661 ( .A(n3813), .B(n31119), .Z(n3814) );
  NAND U4662 ( .A(n3815), .B(n3814), .Z(n3953) );
  XOR U4663 ( .A(b[15]), .B(n16220), .Z(n4045) );
  OR U4664 ( .A(n4045), .B(n32010), .Z(n3818) );
  NAND U4665 ( .A(n3816), .B(n32011), .Z(n3817) );
  NAND U4666 ( .A(n3818), .B(n3817), .Z(n3950) );
  XOR U4667 ( .A(n971), .B(n16269), .Z(n4057) );
  NANDN U4668 ( .A(n31550), .B(n4057), .Z(n3821) );
  NANDN U4669 ( .A(n3819), .B(n31874), .Z(n3820) );
  AND U4670 ( .A(n3821), .B(n3820), .Z(n3951) );
  XNOR U4671 ( .A(n3950), .B(n3951), .Z(n3952) );
  XNOR U4672 ( .A(n3953), .B(n3952), .Z(n3984) );
  XOR U4673 ( .A(n3983), .B(n3984), .Z(n3985) );
  NANDN U4674 ( .A(n3823), .B(n3822), .Z(n3827) );
  NAND U4675 ( .A(n3825), .B(n3824), .Z(n3826) );
  NAND U4676 ( .A(n3827), .B(n3826), .Z(n3986) );
  XOR U4677 ( .A(n3985), .B(n3986), .Z(n3947) );
  NANDN U4678 ( .A(n3829), .B(n3828), .Z(n3833) );
  NAND U4679 ( .A(n3831), .B(n3830), .Z(n3832) );
  NAND U4680 ( .A(n3833), .B(n3832), .Z(n3944) );
  NANDN U4681 ( .A(n3835), .B(n3834), .Z(n3839) );
  NAND U4682 ( .A(n3837), .B(n3836), .Z(n3838) );
  NAND U4683 ( .A(n3839), .B(n3838), .Z(n3945) );
  XNOR U4684 ( .A(n3944), .B(n3945), .Z(n3946) );
  XNOR U4685 ( .A(n3947), .B(n3946), .Z(n4067) );
  XNOR U4686 ( .A(n4066), .B(n4067), .Z(n4068) );
  XOR U4687 ( .A(n4069), .B(n4068), .Z(n4078) );
  NANDN U4688 ( .A(n3844), .B(n35188), .Z(n3846) );
  XNOR U4689 ( .A(n35540), .B(a[7]), .Z(n4018) );
  NANDN U4690 ( .A(n34968), .B(n4018), .Z(n3845) );
  AND U4691 ( .A(n3846), .B(n3845), .Z(n4024) );
  XOR U4692 ( .A(n31123), .B(n18003), .Z(n3974) );
  NAND U4693 ( .A(n3974), .B(n29949), .Z(n3849) );
  NAND U4694 ( .A(n29948), .B(n3847), .Z(n3848) );
  AND U4695 ( .A(n3849), .B(n3848), .Z(n4025) );
  XOR U4696 ( .A(n4024), .B(n4025), .Z(n4026) );
  NAND U4697 ( .A(n3850), .B(n34044), .Z(n3852) );
  XOR U4698 ( .A(n34510), .B(n13509), .Z(n4036) );
  NANDN U4699 ( .A(n33867), .B(n4036), .Z(n3851) );
  AND U4700 ( .A(n3852), .B(n3851), .Z(n4027) );
  XNOR U4701 ( .A(n4026), .B(n4027), .Z(n3997) );
  XNOR U4702 ( .A(b[25]), .B(n12830), .Z(n3977) );
  NANDN U4703 ( .A(n34219), .B(n3977), .Z(n3855) );
  NAND U4704 ( .A(n34217), .B(n3853), .Z(n3854) );
  NAND U4705 ( .A(n3855), .B(n3854), .Z(n4004) );
  NAND U4706 ( .A(n34848), .B(n3856), .Z(n3858) );
  XOR U4707 ( .A(n35375), .B(n12258), .Z(n3980) );
  NAND U4708 ( .A(n34618), .B(n3980), .Z(n3857) );
  NAND U4709 ( .A(n3858), .B(n3857), .Z(n4001) );
  XOR U4710 ( .A(n969), .B(n17960), .Z(n4051) );
  NAND U4711 ( .A(n30509), .B(n4051), .Z(n3861) );
  NANDN U4712 ( .A(n3859), .B(n30846), .Z(n3860) );
  AND U4713 ( .A(n3861), .B(n3860), .Z(n4002) );
  XNOR U4714 ( .A(n4001), .B(n4002), .Z(n4003) );
  XNOR U4715 ( .A(n4004), .B(n4003), .Z(n3995) );
  NANDN U4716 ( .A(n3863), .B(n3862), .Z(n3867) );
  NAND U4717 ( .A(n3865), .B(n3864), .Z(n3866) );
  NAND U4718 ( .A(n3867), .B(n3866), .Z(n3996) );
  XOR U4719 ( .A(n3995), .B(n3996), .Z(n3998) );
  XOR U4720 ( .A(n3997), .B(n3998), .Z(n4075) );
  NANDN U4721 ( .A(n3869), .B(n3868), .Z(n3873) );
  NAND U4722 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4723 ( .A(n3873), .B(n3872), .Z(n4072) );
  XNOR U4724 ( .A(b[21]), .B(a[15]), .Z(n4009) );
  OR U4725 ( .A(n4009), .B(n33634), .Z(n3876) );
  NANDN U4726 ( .A(n3874), .B(n33464), .Z(n3875) );
  NAND U4727 ( .A(n3876), .B(n3875), .Z(n3965) );
  XOR U4728 ( .A(b[5]), .B(n18639), .Z(n4039) );
  OR U4729 ( .A(n4039), .B(n29363), .Z(n3879) );
  NANDN U4730 ( .A(n3877), .B(n29864), .Z(n3878) );
  NAND U4731 ( .A(n3879), .B(n3878), .Z(n3962) );
  XOR U4732 ( .A(b[3]), .B(n19656), .Z(n4012) );
  NANDN U4733 ( .A(n4012), .B(n28939), .Z(n3882) );
  NAND U4734 ( .A(n3880), .B(n28938), .Z(n3881) );
  AND U4735 ( .A(n3882), .B(n3881), .Z(n3963) );
  XNOR U4736 ( .A(n3962), .B(n3963), .Z(n3964) );
  XNOR U4737 ( .A(n3965), .B(n3964), .Z(n3989) );
  XOR U4738 ( .A(b[31]), .B(n11202), .Z(n4021) );
  NANDN U4739 ( .A(n4021), .B(n35313), .Z(n3885) );
  NAND U4740 ( .A(n3883), .B(n35311), .Z(n3884) );
  NAND U4741 ( .A(n3885), .B(n3884), .Z(n3959) );
  XNOR U4742 ( .A(b[17]), .B(a[19]), .Z(n4048) );
  NANDN U4743 ( .A(n4048), .B(n32543), .Z(n3888) );
  NANDN U4744 ( .A(n3886), .B(n32541), .Z(n3887) );
  AND U4745 ( .A(n3888), .B(n3887), .Z(n3957) );
  NANDN U4746 ( .A(n966), .B(a[35]), .Z(n3889) );
  XOR U4747 ( .A(n29232), .B(n3889), .Z(n3891) );
  IV U4748 ( .A(a[34]), .Z(n19513) );
  NANDN U4749 ( .A(n19513), .B(n966), .Z(n3890) );
  AND U4750 ( .A(n3891), .B(n3890), .Z(n3956) );
  XNOR U4751 ( .A(n3957), .B(n3956), .Z(n3958) );
  XOR U4752 ( .A(n3959), .B(n3958), .Z(n3990) );
  XOR U4753 ( .A(n3989), .B(n3990), .Z(n3992) );
  NANDN U4754 ( .A(n3893), .B(n3892), .Z(n3897) );
  NAND U4755 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4756 ( .A(n3897), .B(n3896), .Z(n3991) );
  XOR U4757 ( .A(n3992), .B(n3991), .Z(n4073) );
  XNOR U4758 ( .A(n4075), .B(n4074), .Z(n4061) );
  OR U4759 ( .A(n3899), .B(n3898), .Z(n3903) );
  OR U4760 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4761 ( .A(n3903), .B(n3902), .Z(n4060) );
  XOR U4762 ( .A(n4061), .B(n4060), .Z(n4062) );
  XOR U4763 ( .A(n4063), .B(n4062), .Z(n4079) );
  XNOR U4764 ( .A(n4078), .B(n4079), .Z(n4080) );
  XNOR U4765 ( .A(n4081), .B(n4080), .Z(n3941) );
  NAND U4766 ( .A(n3905), .B(n3904), .Z(n3909) );
  OR U4767 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U4768 ( .A(n3909), .B(n3908), .Z(n3938) );
  NAND U4769 ( .A(n3911), .B(n3910), .Z(n3915) );
  NANDN U4770 ( .A(n3913), .B(n3912), .Z(n3914) );
  NAND U4771 ( .A(n3915), .B(n3914), .Z(n3939) );
  XNOR U4772 ( .A(n3938), .B(n3939), .Z(n3940) );
  XOR U4773 ( .A(n3941), .B(n3940), .Z(n3935) );
  XOR U4774 ( .A(n3934), .B(n3935), .Z(n3926) );
  XOR U4775 ( .A(n3927), .B(n3926), .Z(n3928) );
  XNOR U4776 ( .A(n3929), .B(n3928), .Z(n3921) );
  XNOR U4777 ( .A(n3921), .B(sreg[99]), .Z(n3923) );
  NAND U4778 ( .A(n3916), .B(sreg[98]), .Z(n3920) );
  OR U4779 ( .A(n3918), .B(n3917), .Z(n3919) );
  AND U4780 ( .A(n3920), .B(n3919), .Z(n3922) );
  XOR U4781 ( .A(n3923), .B(n3922), .Z(c[99]) );
  NAND U4782 ( .A(n3921), .B(sreg[99]), .Z(n3925) );
  OR U4783 ( .A(n3923), .B(n3922), .Z(n3924) );
  NAND U4784 ( .A(n3925), .B(n3924), .Z(n4244) );
  XNOR U4785 ( .A(n4244), .B(sreg[100]), .Z(n4246) );
  NAND U4786 ( .A(n3927), .B(n3926), .Z(n3931) );
  NAND U4787 ( .A(n3929), .B(n3928), .Z(n3930) );
  NAND U4788 ( .A(n3931), .B(n3930), .Z(n4087) );
  NANDN U4789 ( .A(n3933), .B(n3932), .Z(n3937) );
  NAND U4790 ( .A(n3935), .B(n3934), .Z(n3936) );
  NAND U4791 ( .A(n3937), .B(n3936), .Z(n4085) );
  NANDN U4792 ( .A(n3939), .B(n3938), .Z(n3943) );
  NAND U4793 ( .A(n3941), .B(n3940), .Z(n3942) );
  NAND U4794 ( .A(n3943), .B(n3942), .Z(n4240) );
  NANDN U4795 ( .A(n3945), .B(n3944), .Z(n3949) );
  NAND U4796 ( .A(n3947), .B(n3946), .Z(n3948) );
  NAND U4797 ( .A(n3949), .B(n3948), .Z(n4099) );
  NANDN U4798 ( .A(n3951), .B(n3950), .Z(n3955) );
  NAND U4799 ( .A(n3953), .B(n3952), .Z(n3954) );
  NAND U4800 ( .A(n3955), .B(n3954), .Z(n4135) );
  NANDN U4801 ( .A(n3957), .B(n3956), .Z(n3961) );
  NAND U4802 ( .A(n3959), .B(n3958), .Z(n3960) );
  AND U4803 ( .A(n3961), .B(n3960), .Z(n4136) );
  XNOR U4804 ( .A(n4135), .B(n4136), .Z(n4137) );
  NANDN U4805 ( .A(n3963), .B(n3962), .Z(n3967) );
  NAND U4806 ( .A(n3965), .B(n3964), .Z(n3966) );
  NAND U4807 ( .A(n3967), .B(n3966), .Z(n4155) );
  IV U4808 ( .A(a[36]), .Z(n19980) );
  NANDN U4809 ( .A(n19980), .B(b[0]), .Z(n3968) );
  XOR U4810 ( .A(n29232), .B(n3968), .Z(n3970) );
  IV U4811 ( .A(a[35]), .Z(n20315) );
  NANDN U4812 ( .A(n20315), .B(n966), .Z(n3969) );
  AND U4813 ( .A(n3970), .B(n3969), .Z(n4100) );
  XOR U4814 ( .A(b[33]), .B(n10854), .Z(n4181) );
  NANDN U4815 ( .A(n4181), .B(n35620), .Z(n3973) );
  NAND U4816 ( .A(n3971), .B(n35621), .Z(n3972) );
  AND U4817 ( .A(n3973), .B(n3972), .Z(n4101) );
  XOR U4818 ( .A(n4100), .B(n4101), .Z(n4102) );
  XOR U4819 ( .A(b[36]), .B(b[35]), .Z(n36311) );
  NANDN U4820 ( .A(n986), .B(n36311), .Z(n4113) );
  XOR U4821 ( .A(n4102), .B(n4113), .Z(n4153) );
  XOR U4822 ( .A(n31123), .B(n18804), .Z(n4121) );
  NAND U4823 ( .A(n4121), .B(n29949), .Z(n3976) );
  NAND U4824 ( .A(n29948), .B(n3974), .Z(n3975) );
  NAND U4825 ( .A(n3976), .B(n3975), .Z(n4196) );
  XNOR U4826 ( .A(b[25]), .B(n13106), .Z(n4211) );
  NANDN U4827 ( .A(n34219), .B(n4211), .Z(n3979) );
  NAND U4828 ( .A(n34217), .B(n3977), .Z(n3978) );
  NAND U4829 ( .A(n3979), .B(n3978), .Z(n4193) );
  NAND U4830 ( .A(n34848), .B(n3980), .Z(n3982) );
  XOR U4831 ( .A(n35375), .B(n12555), .Z(n4175) );
  NAND U4832 ( .A(n34618), .B(n4175), .Z(n3981) );
  AND U4833 ( .A(n3982), .B(n3981), .Z(n4194) );
  XNOR U4834 ( .A(n4193), .B(n4194), .Z(n4195) );
  XNOR U4835 ( .A(n4196), .B(n4195), .Z(n4154) );
  XOR U4836 ( .A(n4153), .B(n4154), .Z(n4156) );
  XNOR U4837 ( .A(n4155), .B(n4156), .Z(n4138) );
  XNOR U4838 ( .A(n4137), .B(n4138), .Z(n4096) );
  OR U4839 ( .A(n3984), .B(n3983), .Z(n3988) );
  NANDN U4840 ( .A(n3986), .B(n3985), .Z(n3987) );
  NAND U4841 ( .A(n3988), .B(n3987), .Z(n4097) );
  XNOR U4842 ( .A(n4096), .B(n4097), .Z(n4098) );
  XOR U4843 ( .A(n4099), .B(n4098), .Z(n4229) );
  NANDN U4844 ( .A(n3990), .B(n3989), .Z(n3994) );
  OR U4845 ( .A(n3992), .B(n3991), .Z(n3993) );
  NAND U4846 ( .A(n3994), .B(n3993), .Z(n4090) );
  NANDN U4847 ( .A(n3996), .B(n3995), .Z(n4000) );
  OR U4848 ( .A(n3998), .B(n3997), .Z(n3999) );
  AND U4849 ( .A(n4000), .B(n3999), .Z(n4091) );
  XNOR U4850 ( .A(n4090), .B(n4091), .Z(n4092) );
  NANDN U4851 ( .A(n4002), .B(n4001), .Z(n4006) );
  NAND U4852 ( .A(n4004), .B(n4003), .Z(n4005) );
  NAND U4853 ( .A(n4006), .B(n4005), .Z(n4223) );
  NAND U4854 ( .A(n4008), .B(n4007), .Z(n4129) );
  XNOR U4855 ( .A(b[21]), .B(n14259), .Z(n4208) );
  NANDN U4856 ( .A(n33634), .B(n4208), .Z(n4011) );
  NANDN U4857 ( .A(n4009), .B(n33464), .Z(n4010) );
  NAND U4858 ( .A(n4011), .B(n4010), .Z(n4128) );
  XOR U4859 ( .A(b[3]), .B(n19513), .Z(n4187) );
  NANDN U4860 ( .A(n4187), .B(n28939), .Z(n4014) );
  NANDN U4861 ( .A(n4012), .B(n28938), .Z(n4013) );
  AND U4862 ( .A(n4014), .B(n4013), .Z(n4127) );
  XNOR U4863 ( .A(n4128), .B(n4127), .Z(n4130) );
  XNOR U4864 ( .A(n4129), .B(n4130), .Z(n4220) );
  NAND U4865 ( .A(n4015), .B(n33283), .Z(n4017) );
  XOR U4866 ( .A(b[19]), .B(n14905), .Z(n4115) );
  OR U4867 ( .A(n4115), .B(n33021), .Z(n4016) );
  NAND U4868 ( .A(n4017), .B(n4016), .Z(n4160) );
  NAND U4869 ( .A(n4018), .B(n35188), .Z(n4020) );
  XOR U4870 ( .A(n35540), .B(n11986), .Z(n4199) );
  NANDN U4871 ( .A(n34968), .B(n4199), .Z(n4019) );
  NAND U4872 ( .A(n4020), .B(n4019), .Z(n4157) );
  XOR U4873 ( .A(b[31]), .B(n11406), .Z(n4202) );
  NANDN U4874 ( .A(n4202), .B(n35313), .Z(n4023) );
  NANDN U4875 ( .A(n4021), .B(n35311), .Z(n4022) );
  AND U4876 ( .A(n4023), .B(n4022), .Z(n4158) );
  XNOR U4877 ( .A(n4157), .B(n4158), .Z(n4159) );
  XNOR U4878 ( .A(n4160), .B(n4159), .Z(n4221) );
  XNOR U4879 ( .A(n4220), .B(n4221), .Z(n4222) );
  XOR U4880 ( .A(n4223), .B(n4222), .Z(n4150) );
  OR U4881 ( .A(n4025), .B(n4024), .Z(n4029) );
  NANDN U4882 ( .A(n4027), .B(n4026), .Z(n4028) );
  NAND U4883 ( .A(n4029), .B(n4028), .Z(n4148) );
  NANDN U4884 ( .A(n4031), .B(n4030), .Z(n4035) );
  NAND U4885 ( .A(n4033), .B(n4032), .Z(n4034) );
  NAND U4886 ( .A(n4035), .B(n4034), .Z(n4141) );
  NAND U4887 ( .A(n34044), .B(n4036), .Z(n4038) );
  XOR U4888 ( .A(n34510), .B(n14210), .Z(n4118) );
  NANDN U4889 ( .A(n33867), .B(n4118), .Z(n4037) );
  NAND U4890 ( .A(n4038), .B(n4037), .Z(n4166) );
  XOR U4891 ( .A(b[5]), .B(n18841), .Z(n4124) );
  OR U4892 ( .A(n4124), .B(n29363), .Z(n4041) );
  NANDN U4893 ( .A(n4039), .B(n29864), .Z(n4040) );
  NAND U4894 ( .A(n4041), .B(n4040), .Z(n4163) );
  XNOR U4895 ( .A(b[35]), .B(a[2]), .Z(n4105) );
  NANDN U4896 ( .A(n4105), .B(n35985), .Z(n4044) );
  NAND U4897 ( .A(n4042), .B(n35986), .Z(n4043) );
  AND U4898 ( .A(n4044), .B(n4043), .Z(n4164) );
  XNOR U4899 ( .A(n4163), .B(n4164), .Z(n4165) );
  XOR U4900 ( .A(n4166), .B(n4165), .Z(n4142) );
  XNOR U4901 ( .A(n4141), .B(n4142), .Z(n4143) );
  NANDN U4902 ( .A(n4045), .B(n32011), .Z(n4047) );
  XOR U4903 ( .A(b[15]), .B(n15963), .Z(n4217) );
  OR U4904 ( .A(n4217), .B(n32010), .Z(n4046) );
  NAND U4905 ( .A(n4047), .B(n4046), .Z(n4133) );
  XNOR U4906 ( .A(b[17]), .B(a[20]), .Z(n4184) );
  NANDN U4907 ( .A(n4184), .B(n32543), .Z(n4050) );
  NANDN U4908 ( .A(n4048), .B(n32541), .Z(n4049) );
  NAND U4909 ( .A(n4050), .B(n4049), .Z(n4131) );
  NAND U4910 ( .A(n30846), .B(n4051), .Z(n4053) );
  XNOR U4911 ( .A(n969), .B(a[28]), .Z(n4178) );
  NAND U4912 ( .A(n30509), .B(n4178), .Z(n4052) );
  NAND U4913 ( .A(n4053), .B(n4052), .Z(n4132) );
  XNOR U4914 ( .A(n4131), .B(n4132), .Z(n4134) );
  XOR U4915 ( .A(n4133), .B(n4134), .Z(n4172) );
  XNOR U4916 ( .A(n970), .B(a[26]), .Z(n4205) );
  NANDN U4917 ( .A(n31369), .B(n4205), .Z(n4056) );
  NANDN U4918 ( .A(n4054), .B(n31119), .Z(n4055) );
  NAND U4919 ( .A(n4056), .B(n4055), .Z(n4170) );
  NAND U4920 ( .A(n31874), .B(n4057), .Z(n4059) );
  XNOR U4921 ( .A(n971), .B(a[24]), .Z(n4214) );
  NANDN U4922 ( .A(n31550), .B(n4214), .Z(n4058) );
  AND U4923 ( .A(n4059), .B(n4058), .Z(n4169) );
  XNOR U4924 ( .A(n4170), .B(n4169), .Z(n4171) );
  XNOR U4925 ( .A(n4172), .B(n4171), .Z(n4144) );
  XOR U4926 ( .A(n4143), .B(n4144), .Z(n4147) );
  XOR U4927 ( .A(n4148), .B(n4147), .Z(n4149) );
  XOR U4928 ( .A(n4150), .B(n4149), .Z(n4093) );
  XOR U4929 ( .A(n4092), .B(n4093), .Z(n4227) );
  OR U4930 ( .A(n4061), .B(n4060), .Z(n4065) );
  NAND U4931 ( .A(n4063), .B(n4062), .Z(n4064) );
  AND U4932 ( .A(n4065), .B(n4064), .Z(n4226) );
  XNOR U4933 ( .A(n4227), .B(n4226), .Z(n4228) );
  XOR U4934 ( .A(n4229), .B(n4228), .Z(n4235) );
  NANDN U4935 ( .A(n4067), .B(n4066), .Z(n4071) );
  NANDN U4936 ( .A(n4069), .B(n4068), .Z(n4070) );
  NAND U4937 ( .A(n4071), .B(n4070), .Z(n4232) );
  OR U4938 ( .A(n4073), .B(n4072), .Z(n4077) );
  NANDN U4939 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U4940 ( .A(n4077), .B(n4076), .Z(n4233) );
  XNOR U4941 ( .A(n4232), .B(n4233), .Z(n4234) );
  XNOR U4942 ( .A(n4235), .B(n4234), .Z(n4238) );
  NANDN U4943 ( .A(n4079), .B(n4078), .Z(n4083) );
  NAND U4944 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U4945 ( .A(n4083), .B(n4082), .Z(n4239) );
  XNOR U4946 ( .A(n4238), .B(n4239), .Z(n4241) );
  XNOR U4947 ( .A(n4240), .B(n4241), .Z(n4084) );
  XOR U4948 ( .A(n4085), .B(n4084), .Z(n4086) );
  XOR U4949 ( .A(n4087), .B(n4086), .Z(n4245) );
  XOR U4950 ( .A(n4246), .B(n4245), .Z(c[100]) );
  NAND U4951 ( .A(n4085), .B(n4084), .Z(n4089) );
  NAND U4952 ( .A(n4087), .B(n4086), .Z(n4088) );
  NAND U4953 ( .A(n4089), .B(n4088), .Z(n4257) );
  NANDN U4954 ( .A(n4091), .B(n4090), .Z(n4095) );
  NANDN U4955 ( .A(n4093), .B(n4092), .Z(n4094) );
  NAND U4956 ( .A(n4095), .B(n4094), .Z(n4399) );
  XNOR U4957 ( .A(n4399), .B(n4400), .Z(n4401) );
  NANDN U4958 ( .A(n4101), .B(n4100), .Z(n4104) );
  OR U4959 ( .A(n4102), .B(n4113), .Z(n4103) );
  AND U4960 ( .A(n4104), .B(n4103), .Z(n4396) );
  XNOR U4961 ( .A(b[35]), .B(n10524), .Z(n4342) );
  NAND U4962 ( .A(n35985), .B(n4342), .Z(n4107) );
  NANDN U4963 ( .A(n4105), .B(n35986), .Z(n4106) );
  NAND U4964 ( .A(n4107), .B(n4106), .Z(n4292) );
  XNOR U4965 ( .A(n975), .B(b[35]), .Z(n4109) );
  XNOR U4966 ( .A(n975), .B(b[36]), .Z(n4108) );
  AND U4967 ( .A(n4109), .B(n4108), .Z(n36309) );
  NANDN U4968 ( .A(n4110), .B(n36309), .Z(n4112) );
  XOR U4969 ( .A(b[37]), .B(n10457), .Z(n4296) );
  NANDN U4970 ( .A(n4296), .B(n36311), .Z(n4111) );
  NAND U4971 ( .A(n4112), .B(n4111), .Z(n4291) );
  XNOR U4972 ( .A(n4292), .B(n4291), .Z(n4311) );
  NAND U4973 ( .A(b[36]), .B(b[35]), .Z(n36580) );
  ANDN U4974 ( .B(n36580), .A(n975), .Z(n4114) );
  AND U4975 ( .A(n4114), .B(n4113), .Z(n4309) );
  NANDN U4976 ( .A(n4115), .B(n33283), .Z(n4117) );
  XNOR U4977 ( .A(n33020), .B(a[19]), .Z(n4299) );
  NANDN U4978 ( .A(n33021), .B(n4299), .Z(n4116) );
  AND U4979 ( .A(n4117), .B(n4116), .Z(n4308) );
  XNOR U4980 ( .A(n4309), .B(n4308), .Z(n4310) );
  XOR U4981 ( .A(n4311), .B(n4310), .Z(n4394) );
  NAND U4982 ( .A(n34044), .B(n4118), .Z(n4120) );
  XOR U4983 ( .A(n34510), .B(n13976), .Z(n4282) );
  NANDN U4984 ( .A(n33867), .B(n4282), .Z(n4119) );
  NAND U4985 ( .A(n4120), .B(n4119), .Z(n4317) );
  XOR U4986 ( .A(n31123), .B(n18639), .Z(n4276) );
  NAND U4987 ( .A(n4276), .B(n29949), .Z(n4123) );
  NAND U4988 ( .A(n29948), .B(n4121), .Z(n4122) );
  NAND U4989 ( .A(n4123), .B(n4122), .Z(n4314) );
  XOR U4990 ( .A(b[5]), .B(n19656), .Z(n4369) );
  OR U4991 ( .A(n4369), .B(n29363), .Z(n4126) );
  NANDN U4992 ( .A(n4124), .B(n29864), .Z(n4125) );
  AND U4993 ( .A(n4126), .B(n4125), .Z(n4315) );
  XNOR U4994 ( .A(n4314), .B(n4315), .Z(n4316) );
  XNOR U4995 ( .A(n4317), .B(n4316), .Z(n4393) );
  XOR U4996 ( .A(n4394), .B(n4393), .Z(n4395) );
  XOR U4997 ( .A(n4396), .B(n4395), .Z(n4327) );
  XNOR U4998 ( .A(n4324), .B(n4325), .Z(n4326) );
  XOR U4999 ( .A(n4327), .B(n4326), .Z(n4259) );
  NANDN U5000 ( .A(n4136), .B(n4135), .Z(n4140) );
  NAND U5001 ( .A(n4138), .B(n4137), .Z(n4139) );
  AND U5002 ( .A(n4140), .B(n4139), .Z(n4258) );
  XOR U5003 ( .A(n4259), .B(n4258), .Z(n4260) );
  NANDN U5004 ( .A(n4142), .B(n4141), .Z(n4146) );
  NANDN U5005 ( .A(n4144), .B(n4143), .Z(n4145) );
  AND U5006 ( .A(n4146), .B(n4145), .Z(n4261) );
  XOR U5007 ( .A(n4260), .B(n4261), .Z(n4408) );
  OR U5008 ( .A(n4148), .B(n4147), .Z(n4152) );
  NANDN U5009 ( .A(n4150), .B(n4149), .Z(n4151) );
  AND U5010 ( .A(n4152), .B(n4151), .Z(n4405) );
  NANDN U5011 ( .A(n4158), .B(n4157), .Z(n4162) );
  NAND U5012 ( .A(n4160), .B(n4159), .Z(n4161) );
  NAND U5013 ( .A(n4162), .B(n4161), .Z(n4330) );
  NANDN U5014 ( .A(n4164), .B(n4163), .Z(n4168) );
  NAND U5015 ( .A(n4166), .B(n4165), .Z(n4167) );
  AND U5016 ( .A(n4168), .B(n4167), .Z(n4331) );
  XNOR U5017 ( .A(n4330), .B(n4331), .Z(n4332) );
  NANDN U5018 ( .A(n4170), .B(n4169), .Z(n4174) );
  NAND U5019 ( .A(n4172), .B(n4171), .Z(n4173) );
  NAND U5020 ( .A(n4174), .B(n4173), .Z(n4333) );
  XOR U5021 ( .A(n4332), .B(n4333), .Z(n4271) );
  NAND U5022 ( .A(n34848), .B(n4175), .Z(n4177) );
  XOR U5023 ( .A(n35375), .B(n12830), .Z(n4375) );
  NAND U5024 ( .A(n34618), .B(n4375), .Z(n4176) );
  NAND U5025 ( .A(n4177), .B(n4176), .Z(n4366) );
  XOR U5026 ( .A(b[9]), .B(n18003), .Z(n4348) );
  NANDN U5027 ( .A(n4348), .B(n30509), .Z(n4180) );
  NAND U5028 ( .A(n4178), .B(n30846), .Z(n4179) );
  NAND U5029 ( .A(n4180), .B(n4179), .Z(n4363) );
  XOR U5030 ( .A(b[33]), .B(n11202), .Z(n4305) );
  NANDN U5031 ( .A(n4305), .B(n35620), .Z(n4183) );
  NANDN U5032 ( .A(n4181), .B(n35621), .Z(n4182) );
  AND U5033 ( .A(n4183), .B(n4182), .Z(n4364) );
  XNOR U5034 ( .A(n4363), .B(n4364), .Z(n4365) );
  XNOR U5035 ( .A(n4366), .B(n4365), .Z(n4390) );
  XNOR U5036 ( .A(b[17]), .B(n16220), .Z(n4378) );
  NAND U5037 ( .A(n4378), .B(n32543), .Z(n4186) );
  NANDN U5038 ( .A(n4184), .B(n32541), .Z(n4185) );
  AND U5039 ( .A(n4186), .B(n4185), .Z(n4360) );
  XNOR U5040 ( .A(n967), .B(a[35]), .Z(n4384) );
  NAND U5041 ( .A(n4384), .B(n28939), .Z(n4189) );
  NANDN U5042 ( .A(n4187), .B(n28938), .Z(n4188) );
  AND U5043 ( .A(n4189), .B(n4188), .Z(n4358) );
  NANDN U5044 ( .A(n966), .B(a[37]), .Z(n4190) );
  XOR U5045 ( .A(n29232), .B(n4190), .Z(n4192) );
  NANDN U5046 ( .A(b[0]), .B(a[36]), .Z(n4191) );
  AND U5047 ( .A(n4192), .B(n4191), .Z(n4357) );
  XNOR U5048 ( .A(n4358), .B(n4357), .Z(n4359) );
  XNOR U5049 ( .A(n4360), .B(n4359), .Z(n4388) );
  NANDN U5050 ( .A(n4194), .B(n4193), .Z(n4198) );
  NAND U5051 ( .A(n4196), .B(n4195), .Z(n4197) );
  NAND U5052 ( .A(n4198), .B(n4197), .Z(n4387) );
  XOR U5053 ( .A(n4388), .B(n4387), .Z(n4389) );
  XOR U5054 ( .A(n4390), .B(n4389), .Z(n4270) );
  XNOR U5055 ( .A(n4271), .B(n4270), .Z(n4273) );
  NAND U5056 ( .A(n35188), .B(n4199), .Z(n4201) );
  XOR U5057 ( .A(n35540), .B(n12258), .Z(n4381) );
  NANDN U5058 ( .A(n34968), .B(n4381), .Z(n4200) );
  NAND U5059 ( .A(n4201), .B(n4200), .Z(n4288) );
  XOR U5060 ( .A(b[31]), .B(n11694), .Z(n4302) );
  NANDN U5061 ( .A(n4302), .B(n35313), .Z(n4204) );
  NANDN U5062 ( .A(n4202), .B(n35311), .Z(n4203) );
  NAND U5063 ( .A(n4204), .B(n4203), .Z(n4285) );
  XOR U5064 ( .A(b[11]), .B(n17960), .Z(n4354) );
  OR U5065 ( .A(n4354), .B(n31369), .Z(n4207) );
  NAND U5066 ( .A(n4205), .B(n31119), .Z(n4206) );
  AND U5067 ( .A(n4207), .B(n4206), .Z(n4286) );
  XNOR U5068 ( .A(n4285), .B(n4286), .Z(n4287) );
  XNOR U5069 ( .A(n4288), .B(n4287), .Z(n4323) );
  XNOR U5070 ( .A(b[21]), .B(a[17]), .Z(n4293) );
  OR U5071 ( .A(n4293), .B(n33634), .Z(n4210) );
  NAND U5072 ( .A(n4208), .B(n33464), .Z(n4209) );
  NAND U5073 ( .A(n4210), .B(n4209), .Z(n4339) );
  XNOR U5074 ( .A(b[25]), .B(n13509), .Z(n4372) );
  NANDN U5075 ( .A(n34219), .B(n4372), .Z(n4213) );
  NAND U5076 ( .A(n34217), .B(n4211), .Z(n4212) );
  NAND U5077 ( .A(n4213), .B(n4212), .Z(n4336) );
  XOR U5078 ( .A(b[13]), .B(n16916), .Z(n4351) );
  OR U5079 ( .A(n4351), .B(n31550), .Z(n4216) );
  NAND U5080 ( .A(n4214), .B(n31874), .Z(n4215) );
  AND U5081 ( .A(n4216), .B(n4215), .Z(n4337) );
  XNOR U5082 ( .A(n4336), .B(n4337), .Z(n4338) );
  XNOR U5083 ( .A(n4339), .B(n4338), .Z(n4320) );
  NANDN U5084 ( .A(n4217), .B(n32011), .Z(n4219) );
  XNOR U5085 ( .A(n972), .B(a[23]), .Z(n4279) );
  NANDN U5086 ( .A(n32010), .B(n4279), .Z(n4218) );
  NAND U5087 ( .A(n4219), .B(n4218), .Z(n4321) );
  XNOR U5088 ( .A(n4320), .B(n4321), .Z(n4322) );
  XOR U5089 ( .A(n4323), .B(n4322), .Z(n4272) );
  XOR U5090 ( .A(n4273), .B(n4272), .Z(n4264) );
  NANDN U5091 ( .A(n4221), .B(n4220), .Z(n4225) );
  NAND U5092 ( .A(n4223), .B(n4222), .Z(n4224) );
  AND U5093 ( .A(n4225), .B(n4224), .Z(n4265) );
  XNOR U5094 ( .A(n4264), .B(n4265), .Z(n4266) );
  XOR U5095 ( .A(n4267), .B(n4266), .Z(n4406) );
  XOR U5096 ( .A(n4405), .B(n4406), .Z(n4407) );
  XOR U5097 ( .A(n4408), .B(n4407), .Z(n4402) );
  XOR U5098 ( .A(n4401), .B(n4402), .Z(n4414) );
  NAND U5099 ( .A(n4227), .B(n4226), .Z(n4231) );
  OR U5100 ( .A(n4229), .B(n4228), .Z(n4230) );
  NAND U5101 ( .A(n4231), .B(n4230), .Z(n4411) );
  NANDN U5102 ( .A(n4233), .B(n4232), .Z(n4237) );
  NANDN U5103 ( .A(n4235), .B(n4234), .Z(n4236) );
  NAND U5104 ( .A(n4237), .B(n4236), .Z(n4412) );
  XNOR U5105 ( .A(n4411), .B(n4412), .Z(n4413) );
  XNOR U5106 ( .A(n4414), .B(n4413), .Z(n4254) );
  NAND U5107 ( .A(n4239), .B(n4238), .Z(n4243) );
  NANDN U5108 ( .A(n4241), .B(n4240), .Z(n4242) );
  AND U5109 ( .A(n4243), .B(n4242), .Z(n4255) );
  XNOR U5110 ( .A(n4254), .B(n4255), .Z(n4256) );
  XNOR U5111 ( .A(n4257), .B(n4256), .Z(n4249) );
  XNOR U5112 ( .A(n4249), .B(sreg[101]), .Z(n4251) );
  NAND U5113 ( .A(n4244), .B(sreg[100]), .Z(n4248) );
  OR U5114 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U5115 ( .A(n4248), .B(n4247), .Z(n4250) );
  XOR U5116 ( .A(n4251), .B(n4250), .Z(c[101]) );
  NAND U5117 ( .A(n4249), .B(sreg[101]), .Z(n4253) );
  OR U5118 ( .A(n4251), .B(n4250), .Z(n4252) );
  NAND U5119 ( .A(n4253), .B(n4252), .Z(n4590) );
  XNOR U5120 ( .A(n4590), .B(sreg[102]), .Z(n4592) );
  OR U5121 ( .A(n4259), .B(n4258), .Z(n4263) );
  NAND U5122 ( .A(n4261), .B(n4260), .Z(n4262) );
  NAND U5123 ( .A(n4263), .B(n4262), .Z(n4428) );
  NANDN U5124 ( .A(n4265), .B(n4264), .Z(n4269) );
  NAND U5125 ( .A(n4267), .B(n4266), .Z(n4268) );
  AND U5126 ( .A(n4269), .B(n4268), .Z(n4427) );
  XNOR U5127 ( .A(n4428), .B(n4427), .Z(n4429) );
  NAND U5128 ( .A(n4271), .B(n4270), .Z(n4275) );
  NANDN U5129 ( .A(n4273), .B(n4272), .Z(n4274) );
  NAND U5130 ( .A(n4275), .B(n4274), .Z(n4434) );
  XOR U5131 ( .A(n31123), .B(n18841), .Z(n4525) );
  NAND U5132 ( .A(n4525), .B(n29949), .Z(n4278) );
  NAND U5133 ( .A(n29948), .B(n4276), .Z(n4277) );
  NAND U5134 ( .A(n4278), .B(n4277), .Z(n4490) );
  XOR U5135 ( .A(b[15]), .B(n16508), .Z(n4568) );
  OR U5136 ( .A(n4568), .B(n32010), .Z(n4281) );
  NAND U5137 ( .A(n4279), .B(n32011), .Z(n4280) );
  NAND U5138 ( .A(n4281), .B(n4280), .Z(n4487) );
  NAND U5139 ( .A(n34044), .B(n4282), .Z(n4284) );
  XOR U5140 ( .A(b[23]), .B(n14259), .Z(n4577) );
  OR U5141 ( .A(n4577), .B(n33867), .Z(n4283) );
  AND U5142 ( .A(n4284), .B(n4283), .Z(n4488) );
  XNOR U5143 ( .A(n4487), .B(n4488), .Z(n4489) );
  XNOR U5144 ( .A(n4490), .B(n4489), .Z(n4586) );
  NANDN U5145 ( .A(n4286), .B(n4285), .Z(n4290) );
  NAND U5146 ( .A(n4288), .B(n4287), .Z(n4289) );
  NAND U5147 ( .A(n4290), .B(n4289), .Z(n4587) );
  XNOR U5148 ( .A(n4586), .B(n4587), .Z(n4588) );
  NAND U5149 ( .A(n4292), .B(n4291), .Z(n4536) );
  XNOR U5150 ( .A(b[21]), .B(a[18]), .Z(n4522) );
  OR U5151 ( .A(n4522), .B(n33634), .Z(n4295) );
  NANDN U5152 ( .A(n4293), .B(n33464), .Z(n4294) );
  NAND U5153 ( .A(n4295), .B(n4294), .Z(n4535) );
  NANDN U5154 ( .A(n4296), .B(n36309), .Z(n4298) );
  XNOR U5155 ( .A(n975), .B(a[2]), .Z(n4511) );
  NAND U5156 ( .A(n4511), .B(n36311), .Z(n4297) );
  AND U5157 ( .A(n4298), .B(n4297), .Z(n4534) );
  XNOR U5158 ( .A(n4535), .B(n4534), .Z(n4537) );
  XNOR U5159 ( .A(n4536), .B(n4537), .Z(n4589) );
  XNOR U5160 ( .A(n4588), .B(n4589), .Z(n4448) );
  NAND U5161 ( .A(n4299), .B(n33283), .Z(n4301) );
  XOR U5162 ( .A(b[19]), .B(n15484), .Z(n4562) );
  OR U5163 ( .A(n4562), .B(n33021), .Z(n4300) );
  NAND U5164 ( .A(n4301), .B(n4300), .Z(n4496) );
  XOR U5165 ( .A(b[31]), .B(n11986), .Z(n4481) );
  NANDN U5166 ( .A(n4481), .B(n35313), .Z(n4304) );
  NANDN U5167 ( .A(n4302), .B(n35311), .Z(n4303) );
  NAND U5168 ( .A(n4304), .B(n4303), .Z(n4493) );
  XOR U5169 ( .A(b[33]), .B(n11406), .Z(n4472) );
  NANDN U5170 ( .A(n4472), .B(n35620), .Z(n4307) );
  NANDN U5171 ( .A(n4305), .B(n35621), .Z(n4306) );
  AND U5172 ( .A(n4307), .B(n4306), .Z(n4494) );
  XNOR U5173 ( .A(n4493), .B(n4494), .Z(n4495) );
  XNOR U5174 ( .A(n4496), .B(n4495), .Z(n4466) );
  NANDN U5175 ( .A(n4309), .B(n4308), .Z(n4313) );
  NAND U5176 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND U5177 ( .A(n4313), .B(n4312), .Z(n4463) );
  NANDN U5178 ( .A(n4315), .B(n4314), .Z(n4319) );
  NAND U5179 ( .A(n4317), .B(n4316), .Z(n4318) );
  NAND U5180 ( .A(n4319), .B(n4318), .Z(n4464) );
  XNOR U5181 ( .A(n4463), .B(n4464), .Z(n4465) );
  XOR U5182 ( .A(n4466), .B(n4465), .Z(n4446) );
  XNOR U5183 ( .A(n4446), .B(n4445), .Z(n4447) );
  XOR U5184 ( .A(n4448), .B(n4447), .Z(n4460) );
  NANDN U5185 ( .A(n4325), .B(n4324), .Z(n4329) );
  NAND U5186 ( .A(n4327), .B(n4326), .Z(n4328) );
  NAND U5187 ( .A(n4329), .B(n4328), .Z(n4457) );
  NANDN U5188 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U5189 ( .A(n4333), .B(n4332), .Z(n4334) );
  NAND U5190 ( .A(n4335), .B(n4334), .Z(n4458) );
  XNOR U5191 ( .A(n4457), .B(n4458), .Z(n4459) );
  XNOR U5192 ( .A(n4460), .B(n4459), .Z(n4433) );
  XNOR U5193 ( .A(n4434), .B(n4433), .Z(n4435) );
  NANDN U5194 ( .A(n4337), .B(n4336), .Z(n4341) );
  NAND U5195 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND U5196 ( .A(n4341), .B(n4340), .Z(n4583) );
  XNOR U5197 ( .A(b[35]), .B(a[4]), .Z(n4475) );
  NANDN U5198 ( .A(n4475), .B(n35985), .Z(n4344) );
  NAND U5199 ( .A(n4342), .B(n35986), .Z(n4343) );
  AND U5200 ( .A(n4344), .B(n4343), .Z(n4551) );
  NANDN U5201 ( .A(n966), .B(a[38]), .Z(n4345) );
  XOR U5202 ( .A(n29232), .B(n4345), .Z(n4347) );
  IV U5203 ( .A(a[37]), .Z(n20352) );
  NANDN U5204 ( .A(n20352), .B(n966), .Z(n4346) );
  AND U5205 ( .A(n4347), .B(n4346), .Z(n4550) );
  XOR U5206 ( .A(n4551), .B(n4550), .Z(n4553) );
  XOR U5207 ( .A(b[37]), .B(b[38]), .Z(n36553) );
  NANDN U5208 ( .A(n986), .B(n36553), .Z(n4552) );
  XOR U5209 ( .A(n4553), .B(n4552), .Z(n4580) );
  XOR U5210 ( .A(n969), .B(n18804), .Z(n4556) );
  NAND U5211 ( .A(n30509), .B(n4556), .Z(n4350) );
  NANDN U5212 ( .A(n4348), .B(n30846), .Z(n4349) );
  NAND U5213 ( .A(n4350), .B(n4349), .Z(n4541) );
  XOR U5214 ( .A(n971), .B(n17133), .Z(n4565) );
  NANDN U5215 ( .A(n31550), .B(n4565), .Z(n4353) );
  NANDN U5216 ( .A(n4351), .B(n31874), .Z(n4352) );
  NAND U5217 ( .A(n4353), .B(n4352), .Z(n4538) );
  XOR U5218 ( .A(b[11]), .B(n17702), .Z(n4559) );
  OR U5219 ( .A(n4559), .B(n31369), .Z(n4356) );
  NANDN U5220 ( .A(n4354), .B(n31119), .Z(n4355) );
  AND U5221 ( .A(n4356), .B(n4355), .Z(n4539) );
  XNOR U5222 ( .A(n4538), .B(n4539), .Z(n4540) );
  XOR U5223 ( .A(n4541), .B(n4540), .Z(n4581) );
  XOR U5224 ( .A(n4580), .B(n4581), .Z(n4582) );
  XOR U5225 ( .A(n4583), .B(n4582), .Z(n4454) );
  NANDN U5226 ( .A(n4358), .B(n4357), .Z(n4362) );
  NANDN U5227 ( .A(n4360), .B(n4359), .Z(n4361) );
  NAND U5228 ( .A(n4362), .B(n4361), .Z(n4452) );
  NANDN U5229 ( .A(n4364), .B(n4363), .Z(n4368) );
  NAND U5230 ( .A(n4366), .B(n4365), .Z(n4367) );
  NAND U5231 ( .A(n4368), .B(n4367), .Z(n4546) );
  XOR U5232 ( .A(b[5]), .B(n19513), .Z(n4484) );
  OR U5233 ( .A(n4484), .B(n29363), .Z(n4371) );
  NANDN U5234 ( .A(n4369), .B(n29864), .Z(n4370) );
  NAND U5235 ( .A(n4371), .B(n4370), .Z(n4502) );
  XNOR U5236 ( .A(b[25]), .B(n14210), .Z(n4469) );
  NANDN U5237 ( .A(n34219), .B(n4469), .Z(n4374) );
  NAND U5238 ( .A(n34217), .B(n4372), .Z(n4373) );
  NAND U5239 ( .A(n4374), .B(n4373), .Z(n4499) );
  NAND U5240 ( .A(n34848), .B(n4375), .Z(n4377) );
  XOR U5241 ( .A(n35375), .B(n13106), .Z(n4528) );
  NAND U5242 ( .A(n34618), .B(n4528), .Z(n4376) );
  AND U5243 ( .A(n4377), .B(n4376), .Z(n4500) );
  XNOR U5244 ( .A(n4499), .B(n4500), .Z(n4501) );
  XNOR U5245 ( .A(n4502), .B(n4501), .Z(n4544) );
  XNOR U5246 ( .A(b[17]), .B(a[22]), .Z(n4478) );
  NANDN U5247 ( .A(n4478), .B(n32543), .Z(n4380) );
  NAND U5248 ( .A(n4378), .B(n32541), .Z(n4379) );
  NAND U5249 ( .A(n4380), .B(n4379), .Z(n4508) );
  NAND U5250 ( .A(n35188), .B(n4381), .Z(n4383) );
  XOR U5251 ( .A(n35540), .B(n12555), .Z(n4531) );
  NANDN U5252 ( .A(n34968), .B(n4531), .Z(n4382) );
  NAND U5253 ( .A(n4383), .B(n4382), .Z(n4505) );
  XOR U5254 ( .A(b[3]), .B(n19980), .Z(n4574) );
  NANDN U5255 ( .A(n4574), .B(n28939), .Z(n4386) );
  NAND U5256 ( .A(n4384), .B(n28938), .Z(n4385) );
  AND U5257 ( .A(n4386), .B(n4385), .Z(n4506) );
  XNOR U5258 ( .A(n4505), .B(n4506), .Z(n4507) );
  XOR U5259 ( .A(n4508), .B(n4507), .Z(n4545) );
  XOR U5260 ( .A(n4544), .B(n4545), .Z(n4547) );
  XNOR U5261 ( .A(n4546), .B(n4547), .Z(n4451) );
  XOR U5262 ( .A(n4452), .B(n4451), .Z(n4453) );
  XOR U5263 ( .A(n4454), .B(n4453), .Z(n4442) );
  OR U5264 ( .A(n4388), .B(n4387), .Z(n4392) );
  NAND U5265 ( .A(n4390), .B(n4389), .Z(n4391) );
  NAND U5266 ( .A(n4392), .B(n4391), .Z(n4439) );
  OR U5267 ( .A(n4394), .B(n4393), .Z(n4398) );
  NANDN U5268 ( .A(n4396), .B(n4395), .Z(n4397) );
  NAND U5269 ( .A(n4398), .B(n4397), .Z(n4440) );
  XNOR U5270 ( .A(n4439), .B(n4440), .Z(n4441) );
  XOR U5271 ( .A(n4442), .B(n4441), .Z(n4436) );
  XOR U5272 ( .A(n4435), .B(n4436), .Z(n4430) );
  XNOR U5273 ( .A(n4429), .B(n4430), .Z(n4423) );
  NANDN U5274 ( .A(n4400), .B(n4399), .Z(n4404) );
  NANDN U5275 ( .A(n4402), .B(n4401), .Z(n4403) );
  NAND U5276 ( .A(n4404), .B(n4403), .Z(n4424) );
  XNOR U5277 ( .A(n4423), .B(n4424), .Z(n4425) );
  OR U5278 ( .A(n4406), .B(n4405), .Z(n4410) );
  NANDN U5279 ( .A(n4408), .B(n4407), .Z(n4409) );
  NAND U5280 ( .A(n4410), .B(n4409), .Z(n4426) );
  XOR U5281 ( .A(n4425), .B(n4426), .Z(n4417) );
  NANDN U5282 ( .A(n4412), .B(n4411), .Z(n4416) );
  NAND U5283 ( .A(n4414), .B(n4413), .Z(n4415) );
  NAND U5284 ( .A(n4416), .B(n4415), .Z(n4418) );
  XNOR U5285 ( .A(n4417), .B(n4418), .Z(n4419) );
  XOR U5286 ( .A(n4420), .B(n4419), .Z(n4591) );
  XOR U5287 ( .A(n4592), .B(n4591), .Z(c[102]) );
  NANDN U5288 ( .A(n4418), .B(n4417), .Z(n4422) );
  NAND U5289 ( .A(n4420), .B(n4419), .Z(n4421) );
  NAND U5290 ( .A(n4422), .B(n4421), .Z(n4603) );
  NANDN U5291 ( .A(n4428), .B(n4427), .Z(n4432) );
  NAND U5292 ( .A(n4430), .B(n4429), .Z(n4431) );
  NAND U5293 ( .A(n4432), .B(n4431), .Z(n4769) );
  NAND U5294 ( .A(n4434), .B(n4433), .Z(n4438) );
  OR U5295 ( .A(n4436), .B(n4435), .Z(n4437) );
  NAND U5296 ( .A(n4438), .B(n4437), .Z(n4766) );
  NANDN U5297 ( .A(n4440), .B(n4439), .Z(n4444) );
  NANDN U5298 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U5299 ( .A(n4444), .B(n4443), .Z(n4760) );
  OR U5300 ( .A(n4446), .B(n4445), .Z(n4450) );
  OR U5301 ( .A(n4448), .B(n4447), .Z(n4449) );
  NAND U5302 ( .A(n4450), .B(n4449), .Z(n4761) );
  XOR U5303 ( .A(n4760), .B(n4761), .Z(n4762) );
  OR U5304 ( .A(n4452), .B(n4451), .Z(n4456) );
  NANDN U5305 ( .A(n4454), .B(n4453), .Z(n4455) );
  AND U5306 ( .A(n4456), .B(n4455), .Z(n4763) );
  XNOR U5307 ( .A(n4762), .B(n4763), .Z(n4604) );
  NANDN U5308 ( .A(n4458), .B(n4457), .Z(n4462) );
  NANDN U5309 ( .A(n4460), .B(n4459), .Z(n4461) );
  NAND U5310 ( .A(n4462), .B(n4461), .Z(n4605) );
  XOR U5311 ( .A(n4604), .B(n4605), .Z(n4606) );
  NANDN U5312 ( .A(n4464), .B(n4463), .Z(n4468) );
  NAND U5313 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U5314 ( .A(n4468), .B(n4467), .Z(n4616) );
  XNOR U5315 ( .A(b[25]), .B(n13976), .Z(n4676) );
  NANDN U5316 ( .A(n34219), .B(n4676), .Z(n4471) );
  NAND U5317 ( .A(n34217), .B(n4469), .Z(n4470) );
  NAND U5318 ( .A(n4471), .B(n4470), .Z(n4724) );
  XOR U5319 ( .A(b[33]), .B(n11694), .Z(n4685) );
  NANDN U5320 ( .A(n4685), .B(n35620), .Z(n4474) );
  NANDN U5321 ( .A(n4472), .B(n35621), .Z(n4473) );
  NAND U5322 ( .A(n4474), .B(n4473), .Z(n4721) );
  XNOR U5323 ( .A(b[35]), .B(a[5]), .Z(n4739) );
  NANDN U5324 ( .A(n4739), .B(n35985), .Z(n4477) );
  NANDN U5325 ( .A(n4475), .B(n35986), .Z(n4476) );
  AND U5326 ( .A(n4477), .B(n4476), .Z(n4722) );
  XNOR U5327 ( .A(n4721), .B(n4722), .Z(n4723) );
  XNOR U5328 ( .A(n4724), .B(n4723), .Z(n4635) );
  XNOR U5329 ( .A(b[17]), .B(a[23]), .Z(n4703) );
  NANDN U5330 ( .A(n4703), .B(n32543), .Z(n4480) );
  NANDN U5331 ( .A(n4478), .B(n32541), .Z(n4479) );
  NAND U5332 ( .A(n4480), .B(n4479), .Z(n4682) );
  XOR U5333 ( .A(b[31]), .B(n12258), .Z(n4691) );
  NANDN U5334 ( .A(n4691), .B(n35313), .Z(n4483) );
  NANDN U5335 ( .A(n4481), .B(n35311), .Z(n4482) );
  NAND U5336 ( .A(n4483), .B(n4482), .Z(n4679) );
  XOR U5337 ( .A(b[5]), .B(n20315), .Z(n4673) );
  OR U5338 ( .A(n4673), .B(n29363), .Z(n4486) );
  NANDN U5339 ( .A(n4484), .B(n29864), .Z(n4485) );
  AND U5340 ( .A(n4486), .B(n4485), .Z(n4680) );
  XNOR U5341 ( .A(n4679), .B(n4680), .Z(n4681) );
  XNOR U5342 ( .A(n4682), .B(n4681), .Z(n4632) );
  NANDN U5343 ( .A(n4488), .B(n4487), .Z(n4492) );
  NAND U5344 ( .A(n4490), .B(n4489), .Z(n4491) );
  NAND U5345 ( .A(n4492), .B(n4491), .Z(n4633) );
  XNOR U5346 ( .A(n4632), .B(n4633), .Z(n4634) );
  XOR U5347 ( .A(n4635), .B(n4634), .Z(n4667) );
  NANDN U5348 ( .A(n4494), .B(n4493), .Z(n4498) );
  NAND U5349 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U5350 ( .A(n4498), .B(n4497), .Z(n4664) );
  NANDN U5351 ( .A(n4500), .B(n4499), .Z(n4504) );
  NAND U5352 ( .A(n4502), .B(n4501), .Z(n4503) );
  AND U5353 ( .A(n4504), .B(n4503), .Z(n4665) );
  XNOR U5354 ( .A(n4664), .B(n4665), .Z(n4666) );
  XNOR U5355 ( .A(n4667), .B(n4666), .Z(n4615) );
  NANDN U5356 ( .A(n4506), .B(n4505), .Z(n4510) );
  NAND U5357 ( .A(n4508), .B(n4507), .Z(n4509) );
  NAND U5358 ( .A(n4510), .B(n4509), .Z(n4641) );
  XOR U5359 ( .A(b[37]), .B(n10524), .Z(n4661) );
  NANDN U5360 ( .A(n4661), .B(n36311), .Z(n4513) );
  NAND U5361 ( .A(n4511), .B(n36309), .Z(n4512) );
  NAND U5362 ( .A(n4513), .B(n4512), .Z(n4651) );
  XOR U5363 ( .A(b[39]), .B(n10457), .Z(n4670) );
  ANDN U5364 ( .B(n36553), .A(n4670), .Z(n4518) );
  XNOR U5365 ( .A(n976), .B(a[0]), .Z(n4516) );
  XNOR U5366 ( .A(n976), .B(b[37]), .Z(n4515) );
  XNOR U5367 ( .A(n976), .B(b[38]), .Z(n4514) );
  AND U5368 ( .A(n4515), .B(n4514), .Z(n36643) );
  NAND U5369 ( .A(n4516), .B(n36643), .Z(n4517) );
  NANDN U5370 ( .A(n4518), .B(n4517), .Z(n4650) );
  XNOR U5371 ( .A(n4651), .B(n4650), .Z(n4745) );
  NANDN U5372 ( .A(n966), .B(a[39]), .Z(n4519) );
  XOR U5373 ( .A(n29232), .B(n4519), .Z(n4521) );
  IV U5374 ( .A(a[38]), .Z(n20686) );
  NANDN U5375 ( .A(n20686), .B(n966), .Z(n4520) );
  AND U5376 ( .A(n4521), .B(n4520), .Z(n4743) );
  XNOR U5377 ( .A(b[21]), .B(n15113), .Z(n4733) );
  NANDN U5378 ( .A(n33634), .B(n4733), .Z(n4524) );
  NANDN U5379 ( .A(n4522), .B(n33464), .Z(n4523) );
  AND U5380 ( .A(n4524), .B(n4523), .Z(n4742) );
  XNOR U5381 ( .A(n4743), .B(n4742), .Z(n4744) );
  XOR U5382 ( .A(n4745), .B(n4744), .Z(n4638) );
  XOR U5383 ( .A(n31123), .B(n19656), .Z(n4736) );
  NAND U5384 ( .A(n4736), .B(n29949), .Z(n4527) );
  NAND U5385 ( .A(n29948), .B(n4525), .Z(n4526) );
  NAND U5386 ( .A(n4527), .B(n4526), .Z(n4655) );
  NAND U5387 ( .A(n34848), .B(n4528), .Z(n4530) );
  XOR U5388 ( .A(n35375), .B(n13509), .Z(n4712) );
  NAND U5389 ( .A(n34618), .B(n4712), .Z(n4529) );
  NAND U5390 ( .A(n4530), .B(n4529), .Z(n4652) );
  NAND U5391 ( .A(n35188), .B(n4531), .Z(n4533) );
  XOR U5392 ( .A(n35540), .B(n12830), .Z(n4688) );
  NANDN U5393 ( .A(n34968), .B(n4688), .Z(n4532) );
  AND U5394 ( .A(n4533), .B(n4532), .Z(n4653) );
  XNOR U5395 ( .A(n4652), .B(n4653), .Z(n4654) );
  XNOR U5396 ( .A(n4655), .B(n4654), .Z(n4639) );
  XOR U5397 ( .A(n4638), .B(n4639), .Z(n4640) );
  XNOR U5398 ( .A(n4641), .B(n4640), .Z(n4629) );
  NANDN U5399 ( .A(n4539), .B(n4538), .Z(n4543) );
  NAND U5400 ( .A(n4541), .B(n4540), .Z(n4542) );
  NAND U5401 ( .A(n4543), .B(n4542), .Z(n4627) );
  XNOR U5402 ( .A(n4626), .B(n4627), .Z(n4628) );
  XOR U5403 ( .A(n4629), .B(n4628), .Z(n4614) );
  XOR U5404 ( .A(n4615), .B(n4614), .Z(n4617) );
  NANDN U5405 ( .A(n4545), .B(n4544), .Z(n4549) );
  OR U5406 ( .A(n4547), .B(n4546), .Z(n4548) );
  NAND U5407 ( .A(n4549), .B(n4548), .Z(n4611) );
  NANDN U5408 ( .A(n4551), .B(n4550), .Z(n4555) );
  OR U5409 ( .A(n4553), .B(n4552), .Z(n4554) );
  NAND U5410 ( .A(n4555), .B(n4554), .Z(n4755) );
  NAND U5411 ( .A(n30846), .B(n4556), .Z(n4558) );
  XNOR U5412 ( .A(n969), .B(a[31]), .Z(n4715) );
  NAND U5413 ( .A(n30509), .B(n4715), .Z(n4557) );
  AND U5414 ( .A(n4558), .B(n4557), .Z(n4750) );
  XNOR U5415 ( .A(n970), .B(a[29]), .Z(n4700) );
  NANDN U5416 ( .A(n31369), .B(n4700), .Z(n4561) );
  NANDN U5417 ( .A(n4559), .B(n31119), .Z(n4560) );
  AND U5418 ( .A(n4561), .B(n4560), .Z(n4749) );
  NANDN U5419 ( .A(n4562), .B(n33283), .Z(n4564) );
  XNOR U5420 ( .A(n33020), .B(a[21]), .Z(n4709) );
  NANDN U5421 ( .A(n33021), .B(n4709), .Z(n4563) );
  AND U5422 ( .A(n4564), .B(n4563), .Z(n4748) );
  XNOR U5423 ( .A(n4749), .B(n4748), .Z(n4751) );
  XNOR U5424 ( .A(n4750), .B(n4751), .Z(n4697) );
  NAND U5425 ( .A(n31874), .B(n4565), .Z(n4567) );
  XNOR U5426 ( .A(n971), .B(a[27]), .Z(n4706) );
  NANDN U5427 ( .A(n31550), .B(n4706), .Z(n4566) );
  NAND U5428 ( .A(n4567), .B(n4566), .Z(n4695) );
  NANDN U5429 ( .A(n4568), .B(n32011), .Z(n4570) );
  XOR U5430 ( .A(b[15]), .B(n16916), .Z(n4718) );
  OR U5431 ( .A(n4718), .B(n32010), .Z(n4569) );
  AND U5432 ( .A(n4570), .B(n4569), .Z(n4694) );
  XNOR U5433 ( .A(n4695), .B(n4694), .Z(n4696) );
  XOR U5434 ( .A(n4697), .B(n4696), .Z(n4754) );
  XOR U5435 ( .A(n4755), .B(n4754), .Z(n4757) );
  NOR U5436 ( .A(b[37]), .B(b[38]), .Z(n4571) );
  NANDN U5437 ( .A(n976), .B(n4571), .Z(n4573) );
  ANDN U5438 ( .B(n36553), .A(n976), .Z(n36646) );
  NANDN U5439 ( .A(a[0]), .B(n36646), .Z(n4572) );
  NAND U5440 ( .A(n4573), .B(n4572), .Z(n4728) );
  XNOR U5441 ( .A(n967), .B(a[37]), .Z(n4644) );
  NAND U5442 ( .A(n4644), .B(n28939), .Z(n4576) );
  NANDN U5443 ( .A(n4574), .B(n28938), .Z(n4575) );
  AND U5444 ( .A(n4576), .B(n4575), .Z(n4727) );
  XNOR U5445 ( .A(n4728), .B(n4727), .Z(n4729) );
  NANDN U5446 ( .A(n4577), .B(n34044), .Z(n4579) );
  XNOR U5447 ( .A(n34510), .B(a[17]), .Z(n4647) );
  NANDN U5448 ( .A(n33867), .B(n4647), .Z(n4578) );
  AND U5449 ( .A(n4579), .B(n4578), .Z(n4730) );
  XNOR U5450 ( .A(n4729), .B(n4730), .Z(n4756) );
  XNOR U5451 ( .A(n4757), .B(n4756), .Z(n4620) );
  NAND U5452 ( .A(n4581), .B(n4580), .Z(n4585) );
  NAND U5453 ( .A(n4583), .B(n4582), .Z(n4584) );
  AND U5454 ( .A(n4585), .B(n4584), .Z(n4621) );
  XNOR U5455 ( .A(n4620), .B(n4621), .Z(n4622) );
  XOR U5456 ( .A(n4622), .B(n4623), .Z(n4610) );
  XNOR U5457 ( .A(n4611), .B(n4610), .Z(n4612) );
  XOR U5458 ( .A(n4613), .B(n4612), .Z(n4607) );
  XOR U5459 ( .A(n4606), .B(n4607), .Z(n4767) );
  XNOR U5460 ( .A(n4766), .B(n4767), .Z(n4768) );
  XOR U5461 ( .A(n4769), .B(n4768), .Z(n4600) );
  XNOR U5462 ( .A(n4601), .B(n4600), .Z(n4602) );
  XNOR U5463 ( .A(n4603), .B(n4602), .Z(n4595) );
  XNOR U5464 ( .A(n4595), .B(sreg[103]), .Z(n4597) );
  NAND U5465 ( .A(n4590), .B(sreg[102]), .Z(n4594) );
  OR U5466 ( .A(n4592), .B(n4591), .Z(n4593) );
  AND U5467 ( .A(n4594), .B(n4593), .Z(n4596) );
  XOR U5468 ( .A(n4597), .B(n4596), .Z(c[103]) );
  NAND U5469 ( .A(n4595), .B(sreg[103]), .Z(n4599) );
  OR U5470 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U5471 ( .A(n4599), .B(n4598), .Z(n4955) );
  XNOR U5472 ( .A(n4955), .B(sreg[104]), .Z(n4957) );
  OR U5473 ( .A(n4605), .B(n4604), .Z(n4609) );
  NAND U5474 ( .A(n4607), .B(n4606), .Z(n4608) );
  NAND U5475 ( .A(n4609), .B(n4608), .Z(n4779) );
  NANDN U5476 ( .A(n4615), .B(n4614), .Z(n4619) );
  OR U5477 ( .A(n4617), .B(n4616), .Z(n4618) );
  NAND U5478 ( .A(n4619), .B(n4618), .Z(n4785) );
  XNOR U5479 ( .A(n4784), .B(n4785), .Z(n4786) );
  NANDN U5480 ( .A(n4621), .B(n4620), .Z(n4625) );
  NAND U5481 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U5482 ( .A(n4625), .B(n4624), .Z(n4954) );
  NANDN U5483 ( .A(n4627), .B(n4626), .Z(n4631) );
  NAND U5484 ( .A(n4629), .B(n4628), .Z(n4630) );
  NAND U5485 ( .A(n4631), .B(n4630), .Z(n4903) );
  NANDN U5486 ( .A(n4633), .B(n4632), .Z(n4637) );
  NAND U5487 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U5488 ( .A(n4637), .B(n4636), .Z(n4906) );
  OR U5489 ( .A(n4639), .B(n4638), .Z(n4643) );
  NAND U5490 ( .A(n4641), .B(n4640), .Z(n4642) );
  NAND U5491 ( .A(n4643), .B(n4642), .Z(n4907) );
  XOR U5492 ( .A(n967), .B(n20686), .Z(n4823) );
  NAND U5493 ( .A(n4823), .B(n28939), .Z(n4646) );
  NAND U5494 ( .A(n4644), .B(n28938), .Z(n4645) );
  NAND U5495 ( .A(n4646), .B(n4645), .Z(n4870) );
  NAND U5496 ( .A(n4647), .B(n34044), .Z(n4649) );
  XOR U5497 ( .A(n34510), .B(n14905), .Z(n4832) );
  NANDN U5498 ( .A(n33867), .B(n4832), .Z(n4648) );
  AND U5499 ( .A(n4649), .B(n4648), .Z(n4871) );
  XNOR U5500 ( .A(n4870), .B(n4871), .Z(n4872) );
  NAND U5501 ( .A(n4651), .B(n4650), .Z(n4873) );
  XOR U5502 ( .A(n4872), .B(n4873), .Z(n4885) );
  NANDN U5503 ( .A(n4653), .B(n4652), .Z(n4657) );
  NAND U5504 ( .A(n4655), .B(n4654), .Z(n4656) );
  NAND U5505 ( .A(n4657), .B(n4656), .Z(n4882) );
  XOR U5506 ( .A(n976), .B(b[40]), .Z(n36905) );
  NOR U5507 ( .A(n986), .B(n36905), .Z(n4942) );
  NANDN U5508 ( .A(n966), .B(a[40]), .Z(n4658) );
  XOR U5509 ( .A(n29232), .B(n4658), .Z(n4660) );
  IV U5510 ( .A(a[39]), .Z(n20867) );
  NANDN U5511 ( .A(n20867), .B(n966), .Z(n4659) );
  AND U5512 ( .A(n4660), .B(n4659), .Z(n4940) );
  NANDN U5513 ( .A(n4661), .B(n36309), .Z(n4663) );
  XNOR U5514 ( .A(n975), .B(a[4]), .Z(n4829) );
  NAND U5515 ( .A(n4829), .B(n36311), .Z(n4662) );
  AND U5516 ( .A(n4663), .B(n4662), .Z(n4939) );
  XNOR U5517 ( .A(n4940), .B(n4939), .Z(n4941) );
  XOR U5518 ( .A(n4942), .B(n4941), .Z(n4883) );
  XOR U5519 ( .A(n4882), .B(n4883), .Z(n4884) );
  XNOR U5520 ( .A(n4885), .B(n4884), .Z(n4909) );
  XOR U5521 ( .A(n4908), .B(n4909), .Z(n4900) );
  NANDN U5522 ( .A(n4665), .B(n4664), .Z(n4669) );
  NANDN U5523 ( .A(n4667), .B(n4666), .Z(n4668) );
  AND U5524 ( .A(n4669), .B(n4668), .Z(n4901) );
  XNOR U5525 ( .A(n4900), .B(n4901), .Z(n4902) );
  XNOR U5526 ( .A(n4903), .B(n4902), .Z(n4951) );
  XOR U5527 ( .A(b[39]), .B(n10363), .Z(n4850) );
  NANDN U5528 ( .A(n4850), .B(n36553), .Z(n4672) );
  NANDN U5529 ( .A(n4670), .B(n36643), .Z(n4671) );
  NAND U5530 ( .A(n4672), .B(n4671), .Z(n4879) );
  XOR U5531 ( .A(b[5]), .B(n19980), .Z(n4811) );
  OR U5532 ( .A(n4811), .B(n29363), .Z(n4675) );
  NANDN U5533 ( .A(n4673), .B(n29864), .Z(n4674) );
  NAND U5534 ( .A(n4675), .B(n4674), .Z(n4876) );
  XNOR U5535 ( .A(b[25]), .B(n14259), .Z(n4805) );
  NANDN U5536 ( .A(n34219), .B(n4805), .Z(n4678) );
  NAND U5537 ( .A(n34217), .B(n4676), .Z(n4677) );
  AND U5538 ( .A(n4678), .B(n4677), .Z(n4877) );
  XNOR U5539 ( .A(n4876), .B(n4877), .Z(n4878) );
  XOR U5540 ( .A(n4879), .B(n4878), .Z(n4890) );
  NANDN U5541 ( .A(n4680), .B(n4679), .Z(n4684) );
  NAND U5542 ( .A(n4682), .B(n4681), .Z(n4683) );
  NAND U5543 ( .A(n4684), .B(n4683), .Z(n4889) );
  XOR U5544 ( .A(b[33]), .B(n11986), .Z(n4808) );
  NANDN U5545 ( .A(n4808), .B(n35620), .Z(n4687) );
  NANDN U5546 ( .A(n4685), .B(n35621), .Z(n4686) );
  NAND U5547 ( .A(n4687), .B(n4686), .Z(n4838) );
  NAND U5548 ( .A(n35188), .B(n4688), .Z(n4690) );
  XOR U5549 ( .A(n35540), .B(n13106), .Z(n4933) );
  NANDN U5550 ( .A(n34968), .B(n4933), .Z(n4689) );
  NAND U5551 ( .A(n4690), .B(n4689), .Z(n4835) );
  XOR U5552 ( .A(b[31]), .B(n12555), .Z(n4936) );
  NANDN U5553 ( .A(n4936), .B(n35313), .Z(n4693) );
  NANDN U5554 ( .A(n4691), .B(n35311), .Z(n4692) );
  AND U5555 ( .A(n4693), .B(n4692), .Z(n4836) );
  XNOR U5556 ( .A(n4835), .B(n4836), .Z(n4837) );
  XOR U5557 ( .A(n4838), .B(n4837), .Z(n4888) );
  XNOR U5558 ( .A(n4889), .B(n4888), .Z(n4891) );
  XNOR U5559 ( .A(n4890), .B(n4891), .Z(n4793) );
  NANDN U5560 ( .A(n4695), .B(n4694), .Z(n4699) );
  NAND U5561 ( .A(n4697), .B(n4696), .Z(n4698) );
  NAND U5562 ( .A(n4699), .B(n4698), .Z(n4791) );
  XOR U5563 ( .A(b[11]), .B(n18804), .Z(n4841) );
  OR U5564 ( .A(n4841), .B(n31369), .Z(n4702) );
  NAND U5565 ( .A(n4700), .B(n31119), .Z(n4701) );
  NAND U5566 ( .A(n4702), .B(n4701), .Z(n4948) );
  XNOR U5567 ( .A(b[17]), .B(a[24]), .Z(n4799) );
  NANDN U5568 ( .A(n4799), .B(n32543), .Z(n4705) );
  NANDN U5569 ( .A(n4703), .B(n32541), .Z(n4704) );
  NAND U5570 ( .A(n4705), .B(n4704), .Z(n4945) );
  XOR U5571 ( .A(b[13]), .B(n17702), .Z(n4847) );
  OR U5572 ( .A(n4847), .B(n31550), .Z(n4708) );
  NAND U5573 ( .A(n4706), .B(n31874), .Z(n4707) );
  AND U5574 ( .A(n4708), .B(n4707), .Z(n4946) );
  XNOR U5575 ( .A(n4945), .B(n4946), .Z(n4947) );
  XOR U5576 ( .A(n4948), .B(n4947), .Z(n4920) );
  NAND U5577 ( .A(n4709), .B(n33283), .Z(n4711) );
  XOR U5578 ( .A(n33020), .B(n15963), .Z(n4820) );
  NANDN U5579 ( .A(n33021), .B(n4820), .Z(n4710) );
  NAND U5580 ( .A(n4711), .B(n4710), .Z(n4867) );
  NAND U5581 ( .A(n34848), .B(n4712), .Z(n4714) );
  XOR U5582 ( .A(n35375), .B(n14210), .Z(n4802) );
  NAND U5583 ( .A(n34618), .B(n4802), .Z(n4713) );
  NAND U5584 ( .A(n4714), .B(n4713), .Z(n4864) );
  XOR U5585 ( .A(b[9]), .B(n18841), .Z(n4844) );
  NANDN U5586 ( .A(n4844), .B(n30509), .Z(n4717) );
  NAND U5587 ( .A(n4715), .B(n30846), .Z(n4716) );
  AND U5588 ( .A(n4717), .B(n4716), .Z(n4865) );
  XNOR U5589 ( .A(n4864), .B(n4865), .Z(n4866) );
  XOR U5590 ( .A(n4867), .B(n4866), .Z(n4918) );
  NANDN U5591 ( .A(n4718), .B(n32011), .Z(n4720) );
  XNOR U5592 ( .A(n972), .B(a[26]), .Z(n4930) );
  NANDN U5593 ( .A(n32010), .B(n4930), .Z(n4719) );
  NAND U5594 ( .A(n4720), .B(n4719), .Z(n4919) );
  XNOR U5595 ( .A(n4918), .B(n4919), .Z(n4921) );
  XNOR U5596 ( .A(n4920), .B(n4921), .Z(n4926) );
  NANDN U5597 ( .A(n4722), .B(n4721), .Z(n4726) );
  NAND U5598 ( .A(n4724), .B(n4723), .Z(n4725) );
  AND U5599 ( .A(n4726), .B(n4725), .Z(n4924) );
  NANDN U5600 ( .A(n4728), .B(n4727), .Z(n4732) );
  NAND U5601 ( .A(n4730), .B(n4729), .Z(n4731) );
  NAND U5602 ( .A(n4732), .B(n4731), .Z(n4925) );
  XNOR U5603 ( .A(n4924), .B(n4925), .Z(n4927) );
  XOR U5604 ( .A(n4926), .B(n4927), .Z(n4790) );
  XNOR U5605 ( .A(n4791), .B(n4790), .Z(n4792) );
  XNOR U5606 ( .A(n4793), .B(n4792), .Z(n4915) );
  XNOR U5607 ( .A(b[21]), .B(a[20]), .Z(n4861) );
  OR U5608 ( .A(n4861), .B(n33634), .Z(n4735) );
  NAND U5609 ( .A(n4733), .B(n33464), .Z(n4734) );
  NAND U5610 ( .A(n4735), .B(n4734), .Z(n4817) );
  XOR U5611 ( .A(n31123), .B(n19513), .Z(n4796) );
  NAND U5612 ( .A(n4796), .B(n29949), .Z(n4738) );
  NAND U5613 ( .A(n29948), .B(n4736), .Z(n4737) );
  NAND U5614 ( .A(n4738), .B(n4737), .Z(n4814) );
  XNOR U5615 ( .A(b[35]), .B(a[6]), .Z(n4826) );
  NANDN U5616 ( .A(n4826), .B(n35985), .Z(n4741) );
  NANDN U5617 ( .A(n4739), .B(n35986), .Z(n4740) );
  AND U5618 ( .A(n4741), .B(n4740), .Z(n4815) );
  XNOR U5619 ( .A(n4814), .B(n4815), .Z(n4816) );
  XNOR U5620 ( .A(n4817), .B(n4816), .Z(n4897) );
  NANDN U5621 ( .A(n4743), .B(n4742), .Z(n4747) );
  NAND U5622 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U5623 ( .A(n4747), .B(n4746), .Z(n4894) );
  OR U5624 ( .A(n4749), .B(n4748), .Z(n4753) );
  OR U5625 ( .A(n4751), .B(n4750), .Z(n4752) );
  NAND U5626 ( .A(n4753), .B(n4752), .Z(n4895) );
  XNOR U5627 ( .A(n4894), .B(n4895), .Z(n4896) );
  XOR U5628 ( .A(n4897), .B(n4896), .Z(n4912) );
  NANDN U5629 ( .A(n4755), .B(n4754), .Z(n4759) );
  OR U5630 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5631 ( .A(n4759), .B(n4758), .Z(n4913) );
  XOR U5632 ( .A(n4912), .B(n4913), .Z(n4914) );
  XOR U5633 ( .A(n4915), .B(n4914), .Z(n4952) );
  XOR U5634 ( .A(n4951), .B(n4952), .Z(n4953) );
  XOR U5635 ( .A(n4954), .B(n4953), .Z(n4787) );
  XOR U5636 ( .A(n4786), .B(n4787), .Z(n4778) );
  XNOR U5637 ( .A(n4779), .B(n4778), .Z(n4781) );
  OR U5638 ( .A(n4761), .B(n4760), .Z(n4765) );
  NANDN U5639 ( .A(n4763), .B(n4762), .Z(n4764) );
  NAND U5640 ( .A(n4765), .B(n4764), .Z(n4780) );
  XNOR U5641 ( .A(n4781), .B(n4780), .Z(n4772) );
  NANDN U5642 ( .A(n4767), .B(n4766), .Z(n4771) );
  NAND U5643 ( .A(n4769), .B(n4768), .Z(n4770) );
  AND U5644 ( .A(n4771), .B(n4770), .Z(n4773) );
  XNOR U5645 ( .A(n4772), .B(n4773), .Z(n4774) );
  XOR U5646 ( .A(n4775), .B(n4774), .Z(n4956) );
  XOR U5647 ( .A(n4957), .B(n4956), .Z(c[104]) );
  NANDN U5648 ( .A(n4773), .B(n4772), .Z(n4777) );
  NAND U5649 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U5650 ( .A(n4777), .B(n4776), .Z(n4968) );
  NAND U5651 ( .A(n4779), .B(n4778), .Z(n4783) );
  OR U5652 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U5653 ( .A(n4783), .B(n4782), .Z(n4966) );
  NANDN U5654 ( .A(n4785), .B(n4784), .Z(n4789) );
  NAND U5655 ( .A(n4787), .B(n4786), .Z(n4788) );
  NAND U5656 ( .A(n4789), .B(n4788), .Z(n5140) );
  NAND U5657 ( .A(n4791), .B(n4790), .Z(n4795) );
  OR U5658 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U5659 ( .A(n4795), .B(n4794), .Z(n5033) );
  XOR U5660 ( .A(n31123), .B(n20315), .Z(n5096) );
  NAND U5661 ( .A(n5096), .B(n29949), .Z(n4798) );
  NAND U5662 ( .A(n29948), .B(n4796), .Z(n4797) );
  NAND U5663 ( .A(n4798), .B(n4797), .Z(n5061) );
  XNOR U5664 ( .A(b[17]), .B(a[25]), .Z(n5114) );
  NANDN U5665 ( .A(n5114), .B(n32543), .Z(n4801) );
  NANDN U5666 ( .A(n4799), .B(n32541), .Z(n4800) );
  NAND U5667 ( .A(n4801), .B(n4800), .Z(n5058) );
  NAND U5668 ( .A(n34848), .B(n4802), .Z(n4804) );
  XOR U5669 ( .A(n35375), .B(n13976), .Z(n5093) );
  NAND U5670 ( .A(n34618), .B(n5093), .Z(n4803) );
  AND U5671 ( .A(n4804), .B(n4803), .Z(n5059) );
  XNOR U5672 ( .A(n5058), .B(n5059), .Z(n5060) );
  XNOR U5673 ( .A(n5061), .B(n5060), .Z(n5057) );
  XNOR U5674 ( .A(b[25]), .B(n14514), .Z(n5072) );
  NANDN U5675 ( .A(n34219), .B(n5072), .Z(n4807) );
  NAND U5676 ( .A(n34217), .B(n4805), .Z(n4806) );
  NAND U5677 ( .A(n4807), .B(n4806), .Z(n5084) );
  XOR U5678 ( .A(b[33]), .B(n12258), .Z(n5002) );
  NANDN U5679 ( .A(n5002), .B(n35620), .Z(n4810) );
  NANDN U5680 ( .A(n4808), .B(n35621), .Z(n4809) );
  NAND U5681 ( .A(n4810), .B(n4809), .Z(n5081) );
  XOR U5682 ( .A(b[5]), .B(n20352), .Z(n5075) );
  OR U5683 ( .A(n5075), .B(n29363), .Z(n4813) );
  NANDN U5684 ( .A(n4811), .B(n29864), .Z(n4812) );
  AND U5685 ( .A(n4813), .B(n4812), .Z(n5082) );
  XNOR U5686 ( .A(n5081), .B(n5082), .Z(n5083) );
  XNOR U5687 ( .A(n5084), .B(n5083), .Z(n5054) );
  NANDN U5688 ( .A(n4815), .B(n4814), .Z(n4819) );
  NAND U5689 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U5690 ( .A(n4819), .B(n4818), .Z(n5055) );
  XNOR U5691 ( .A(n5054), .B(n5055), .Z(n5056) );
  XOR U5692 ( .A(n5057), .B(n5056), .Z(n5038) );
  NAND U5693 ( .A(n33283), .B(n4820), .Z(n4822) );
  XOR U5694 ( .A(b[19]), .B(n16269), .Z(n5123) );
  OR U5695 ( .A(n5123), .B(n33021), .Z(n4821) );
  NAND U5696 ( .A(n4822), .B(n4821), .Z(n5017) );
  XOR U5697 ( .A(b[3]), .B(n20867), .Z(n5069) );
  NANDN U5698 ( .A(n5069), .B(n28939), .Z(n4825) );
  NAND U5699 ( .A(n28938), .B(n4823), .Z(n4824) );
  NAND U5700 ( .A(n4825), .B(n4824), .Z(n5014) );
  XNOR U5701 ( .A(b[35]), .B(a[7]), .Z(n5005) );
  NANDN U5702 ( .A(n5005), .B(n35985), .Z(n4828) );
  NANDN U5703 ( .A(n4826), .B(n35986), .Z(n4827) );
  AND U5704 ( .A(n4828), .B(n4827), .Z(n5015) );
  XNOR U5705 ( .A(n5014), .B(n5015), .Z(n5016) );
  XNOR U5706 ( .A(n5017), .B(n5016), .Z(n5047) );
  XOR U5707 ( .A(b[37]), .B(n11202), .Z(n5099) );
  NANDN U5708 ( .A(n5099), .B(n36311), .Z(n4831) );
  NAND U5709 ( .A(n4829), .B(n36309), .Z(n4830) );
  NAND U5710 ( .A(n4831), .B(n4830), .Z(n5011) );
  NAND U5711 ( .A(n34044), .B(n4832), .Z(n4834) );
  XOR U5712 ( .A(b[23]), .B(n15113), .Z(n5066) );
  OR U5713 ( .A(n5066), .B(n33867), .Z(n4833) );
  NAND U5714 ( .A(n4834), .B(n4833), .Z(n5008) );
  XNOR U5715 ( .A(n5008), .B(n5009), .Z(n5010) );
  XNOR U5716 ( .A(n5011), .B(n5010), .Z(n5044) );
  NANDN U5717 ( .A(n4836), .B(n4835), .Z(n4840) );
  NAND U5718 ( .A(n4838), .B(n4837), .Z(n4839) );
  NAND U5719 ( .A(n4840), .B(n4839), .Z(n5045) );
  XNOR U5720 ( .A(n5044), .B(n5045), .Z(n5046) );
  XOR U5721 ( .A(n5047), .B(n5046), .Z(n5039) );
  XOR U5722 ( .A(n5038), .B(n5039), .Z(n5040) );
  XOR U5723 ( .A(b[11]), .B(n18639), .Z(n5105) );
  OR U5724 ( .A(n5105), .B(n31369), .Z(n4843) );
  NANDN U5725 ( .A(n4841), .B(n31119), .Z(n4842) );
  NAND U5726 ( .A(n4843), .B(n4842), .Z(n5129) );
  XOR U5727 ( .A(b[9]), .B(n19656), .Z(n5108) );
  NANDN U5728 ( .A(n5108), .B(n30509), .Z(n4846) );
  NANDN U5729 ( .A(n4844), .B(n30846), .Z(n4845) );
  NAND U5730 ( .A(n4846), .B(n4845), .Z(n5126) );
  XOR U5731 ( .A(b[13]), .B(n18003), .Z(n4999) );
  OR U5732 ( .A(n4999), .B(n31550), .Z(n4849) );
  NANDN U5733 ( .A(n4847), .B(n31874), .Z(n4848) );
  AND U5734 ( .A(n4849), .B(n4848), .Z(n5127) );
  XNOR U5735 ( .A(n5126), .B(n5127), .Z(n5128) );
  XNOR U5736 ( .A(n5129), .B(n5128), .Z(n5021) );
  XOR U5737 ( .A(b[39]), .B(n10524), .Z(n4996) );
  NANDN U5738 ( .A(n4996), .B(n36553), .Z(n4852) );
  NANDN U5739 ( .A(n4850), .B(n36643), .Z(n4851) );
  NAND U5740 ( .A(n4852), .B(n4851), .Z(n5065) );
  XNOR U5741 ( .A(b[41]), .B(n10457), .Z(n5078) );
  ANDN U5742 ( .B(n5078), .A(n36905), .Z(n4857) );
  XNOR U5743 ( .A(b[41]), .B(n986), .Z(n4855) );
  XNOR U5744 ( .A(b[41]), .B(n976), .Z(n4854) );
  XOR U5745 ( .A(b[41]), .B(b[40]), .Z(n4853) );
  AND U5746 ( .A(n4854), .B(n4853), .Z(n36807) );
  NAND U5747 ( .A(n4855), .B(n36807), .Z(n4856) );
  NANDN U5748 ( .A(n4857), .B(n4856), .Z(n5064) );
  XNOR U5749 ( .A(n5065), .B(n5064), .Z(n5090) );
  NANDN U5750 ( .A(n966), .B(a[41]), .Z(n4858) );
  XOR U5751 ( .A(n29232), .B(n4858), .Z(n4860) );
  IV U5752 ( .A(a[40]), .Z(n21149) );
  NANDN U5753 ( .A(n21149), .B(n966), .Z(n4859) );
  AND U5754 ( .A(n4860), .B(n4859), .Z(n5088) );
  XNOR U5755 ( .A(b[21]), .B(a[21]), .Z(n5120) );
  OR U5756 ( .A(n5120), .B(n33634), .Z(n4863) );
  NANDN U5757 ( .A(n4861), .B(n33464), .Z(n4862) );
  AND U5758 ( .A(n4863), .B(n4862), .Z(n5087) );
  XNOR U5759 ( .A(n5088), .B(n5087), .Z(n5089) );
  XOR U5760 ( .A(n5090), .B(n5089), .Z(n5020) );
  XOR U5761 ( .A(n5021), .B(n5020), .Z(n5022) );
  NANDN U5762 ( .A(n4865), .B(n4864), .Z(n4869) );
  NAND U5763 ( .A(n4867), .B(n4866), .Z(n4868) );
  AND U5764 ( .A(n4869), .B(n4868), .Z(n5023) );
  XNOR U5765 ( .A(n5022), .B(n5023), .Z(n5051) );
  NANDN U5766 ( .A(n4871), .B(n4870), .Z(n4875) );
  NANDN U5767 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U5768 ( .A(n4875), .B(n4874), .Z(n5049) );
  NANDN U5769 ( .A(n4877), .B(n4876), .Z(n4881) );
  NAND U5770 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U5771 ( .A(n4881), .B(n4880), .Z(n5048) );
  XNOR U5772 ( .A(n5049), .B(n5048), .Z(n5050) );
  XOR U5773 ( .A(n5051), .B(n5050), .Z(n5041) );
  XNOR U5774 ( .A(n5040), .B(n5041), .Z(n5032) );
  XNOR U5775 ( .A(n5033), .B(n5032), .Z(n5034) );
  OR U5776 ( .A(n4883), .B(n4882), .Z(n4887) );
  NAND U5777 ( .A(n4885), .B(n4884), .Z(n4886) );
  AND U5778 ( .A(n4887), .B(n4886), .Z(n4978) );
  OR U5779 ( .A(n4889), .B(n4888), .Z(n4893) );
  OR U5780 ( .A(n4891), .B(n4890), .Z(n4892) );
  AND U5781 ( .A(n4893), .B(n4892), .Z(n4975) );
  NANDN U5782 ( .A(n4895), .B(n4894), .Z(n4899) );
  NAND U5783 ( .A(n4897), .B(n4896), .Z(n4898) );
  AND U5784 ( .A(n4899), .B(n4898), .Z(n4976) );
  XNOR U5785 ( .A(n4975), .B(n4976), .Z(n4977) );
  XNOR U5786 ( .A(n5034), .B(n5035), .Z(n5135) );
  NANDN U5787 ( .A(n4901), .B(n4900), .Z(n4905) );
  NANDN U5788 ( .A(n4903), .B(n4902), .Z(n4904) );
  NAND U5789 ( .A(n4905), .B(n4904), .Z(n5132) );
  OR U5790 ( .A(n4907), .B(n4906), .Z(n4911) );
  NANDN U5791 ( .A(n4909), .B(n4908), .Z(n4910) );
  NAND U5792 ( .A(n4911), .B(n4910), .Z(n4970) );
  OR U5793 ( .A(n4913), .B(n4912), .Z(n4917) );
  NAND U5794 ( .A(n4915), .B(n4914), .Z(n4916) );
  AND U5795 ( .A(n4917), .B(n4916), .Z(n4969) );
  XOR U5796 ( .A(n4970), .B(n4969), .Z(n4971) );
  OR U5797 ( .A(n4919), .B(n4918), .Z(n4923) );
  OR U5798 ( .A(n4921), .B(n4920), .Z(n4922) );
  NAND U5799 ( .A(n4923), .B(n4922), .Z(n4981) );
  OR U5800 ( .A(n4925), .B(n4924), .Z(n4929) );
  NANDN U5801 ( .A(n4927), .B(n4926), .Z(n4928) );
  NAND U5802 ( .A(n4929), .B(n4928), .Z(n4982) );
  XNOR U5803 ( .A(n4981), .B(n4982), .Z(n4983) );
  XOR U5804 ( .A(b[15]), .B(n17960), .Z(n5111) );
  OR U5805 ( .A(n5111), .B(n32010), .Z(n4932) );
  NAND U5806 ( .A(n4930), .B(n32011), .Z(n4931) );
  NAND U5807 ( .A(n4932), .B(n4931), .Z(n4990) );
  NAND U5808 ( .A(n35188), .B(n4933), .Z(n4935) );
  XOR U5809 ( .A(n35540), .B(n13509), .Z(n5102) );
  NANDN U5810 ( .A(n34968), .B(n5102), .Z(n4934) );
  NAND U5811 ( .A(n4935), .B(n4934), .Z(n4987) );
  XOR U5812 ( .A(b[31]), .B(n12830), .Z(n5117) );
  NANDN U5813 ( .A(n5117), .B(n35313), .Z(n4938) );
  NANDN U5814 ( .A(n4936), .B(n35311), .Z(n4937) );
  AND U5815 ( .A(n4938), .B(n4937), .Z(n4988) );
  XNOR U5816 ( .A(n4987), .B(n4988), .Z(n4989) );
  XNOR U5817 ( .A(n4990), .B(n4989), .Z(n5029) );
  NANDN U5818 ( .A(n4940), .B(n4939), .Z(n4944) );
  NANDN U5819 ( .A(n4942), .B(n4941), .Z(n4943) );
  NAND U5820 ( .A(n4944), .B(n4943), .Z(n5026) );
  NANDN U5821 ( .A(n4946), .B(n4945), .Z(n4950) );
  NAND U5822 ( .A(n4948), .B(n4947), .Z(n4949) );
  NAND U5823 ( .A(n4950), .B(n4949), .Z(n5027) );
  XNOR U5824 ( .A(n5026), .B(n5027), .Z(n5028) );
  XOR U5825 ( .A(n5029), .B(n5028), .Z(n4984) );
  XOR U5826 ( .A(n4983), .B(n4984), .Z(n4972) );
  XOR U5827 ( .A(n4971), .B(n4972), .Z(n5133) );
  XNOR U5828 ( .A(n5132), .B(n5133), .Z(n5134) );
  XNOR U5829 ( .A(n5135), .B(n5134), .Z(n5138) );
  XOR U5830 ( .A(n5138), .B(n5139), .Z(n5141) );
  XOR U5831 ( .A(n5140), .B(n5141), .Z(n4965) );
  XNOR U5832 ( .A(n4966), .B(n4965), .Z(n4967) );
  XNOR U5833 ( .A(n4968), .B(n4967), .Z(n4960) );
  XNOR U5834 ( .A(n4960), .B(sreg[105]), .Z(n4962) );
  NAND U5835 ( .A(n4955), .B(sreg[104]), .Z(n4959) );
  OR U5836 ( .A(n4957), .B(n4956), .Z(n4958) );
  AND U5837 ( .A(n4959), .B(n4958), .Z(n4961) );
  XOR U5838 ( .A(n4962), .B(n4961), .Z(c[105]) );
  NAND U5839 ( .A(n4960), .B(sreg[105]), .Z(n4964) );
  OR U5840 ( .A(n4962), .B(n4961), .Z(n4963) );
  NAND U5841 ( .A(n4964), .B(n4963), .Z(n5332) );
  XNOR U5842 ( .A(n5332), .B(sreg[106]), .Z(n5334) );
  OR U5843 ( .A(n4970), .B(n4969), .Z(n4974) );
  NANDN U5844 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5845 ( .A(n4974), .B(n4973), .Z(n5153) );
  OR U5846 ( .A(n4976), .B(n4975), .Z(n4980) );
  OR U5847 ( .A(n4978), .B(n4977), .Z(n4979) );
  AND U5848 ( .A(n4980), .B(n4979), .Z(n5162) );
  NANDN U5849 ( .A(n4982), .B(n4981), .Z(n4986) );
  NAND U5850 ( .A(n4984), .B(n4983), .Z(n4985) );
  AND U5851 ( .A(n4986), .B(n4985), .Z(n5163) );
  XOR U5852 ( .A(n5162), .B(n5163), .Z(n5164) );
  NANDN U5853 ( .A(n4988), .B(n4987), .Z(n4992) );
  NAND U5854 ( .A(n4990), .B(n4989), .Z(n4991) );
  NAND U5855 ( .A(n4992), .B(n4991), .Z(n5272) );
  NANDN U5856 ( .A(n966), .B(a[42]), .Z(n4993) );
  XOR U5857 ( .A(n29232), .B(n4993), .Z(n4995) );
  IV U5858 ( .A(a[41]), .Z(n21441) );
  NANDN U5859 ( .A(n21441), .B(n966), .Z(n4994) );
  AND U5860 ( .A(n4995), .B(n4994), .Z(n5209) );
  XOR U5861 ( .A(b[39]), .B(n10854), .Z(n5280) );
  NANDN U5862 ( .A(n5280), .B(n36553), .Z(n4998) );
  NANDN U5863 ( .A(n4996), .B(n36643), .Z(n4997) );
  NAND U5864 ( .A(n4998), .B(n4997), .Z(n5207) );
  XOR U5865 ( .A(b[41]), .B(b[42]), .Z(n37068) );
  NANDN U5866 ( .A(n986), .B(n37068), .Z(n5208) );
  XNOR U5867 ( .A(n5207), .B(n5208), .Z(n5210) );
  XOR U5868 ( .A(n5209), .B(n5210), .Z(n5270) );
  XOR U5869 ( .A(b[13]), .B(n18804), .Z(n5286) );
  OR U5870 ( .A(n5286), .B(n31550), .Z(n5001) );
  NANDN U5871 ( .A(n4999), .B(n31874), .Z(n5000) );
  NAND U5872 ( .A(n5001), .B(n5000), .Z(n5181) );
  XOR U5873 ( .A(b[33]), .B(n12555), .Z(n5245) );
  NANDN U5874 ( .A(n5245), .B(n35620), .Z(n5004) );
  NANDN U5875 ( .A(n5002), .B(n35621), .Z(n5003) );
  NAND U5876 ( .A(n5004), .B(n5003), .Z(n5178) );
  XNOR U5877 ( .A(b[35]), .B(a[8]), .Z(n5248) );
  NANDN U5878 ( .A(n5248), .B(n35985), .Z(n5007) );
  NANDN U5879 ( .A(n5005), .B(n35986), .Z(n5006) );
  AND U5880 ( .A(n5007), .B(n5006), .Z(n5179) );
  XNOR U5881 ( .A(n5178), .B(n5179), .Z(n5180) );
  XNOR U5882 ( .A(n5181), .B(n5180), .Z(n5271) );
  XNOR U5883 ( .A(n5270), .B(n5271), .Z(n5273) );
  XNOR U5884 ( .A(n5272), .B(n5273), .Z(n5323) );
  NANDN U5885 ( .A(n5009), .B(n5008), .Z(n5013) );
  NAND U5886 ( .A(n5011), .B(n5010), .Z(n5012) );
  NAND U5887 ( .A(n5013), .B(n5012), .Z(n5321) );
  NANDN U5888 ( .A(n5015), .B(n5014), .Z(n5019) );
  NAND U5889 ( .A(n5017), .B(n5016), .Z(n5018) );
  AND U5890 ( .A(n5019), .B(n5018), .Z(n5320) );
  XNOR U5891 ( .A(n5321), .B(n5320), .Z(n5322) );
  XOR U5892 ( .A(n5323), .B(n5322), .Z(n5168) );
  NAND U5893 ( .A(n5021), .B(n5020), .Z(n5025) );
  NAND U5894 ( .A(n5023), .B(n5022), .Z(n5024) );
  NAND U5895 ( .A(n5025), .B(n5024), .Z(n5169) );
  XOR U5896 ( .A(n5168), .B(n5169), .Z(n5170) );
  NANDN U5897 ( .A(n5027), .B(n5026), .Z(n5031) );
  NAND U5898 ( .A(n5029), .B(n5028), .Z(n5030) );
  AND U5899 ( .A(n5031), .B(n5030), .Z(n5171) );
  XOR U5900 ( .A(n5170), .B(n5171), .Z(n5165) );
  XOR U5901 ( .A(n5164), .B(n5165), .Z(n5159) );
  NAND U5902 ( .A(n5033), .B(n5032), .Z(n5037) );
  OR U5903 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U5904 ( .A(n5037), .B(n5036), .Z(n5156) );
  NAND U5905 ( .A(n5039), .B(n5038), .Z(n5043) );
  NANDN U5906 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5907 ( .A(n5043), .B(n5042), .Z(n5263) );
  NANDN U5908 ( .A(n5049), .B(n5048), .Z(n5053) );
  NANDN U5909 ( .A(n5051), .B(n5050), .Z(n5052) );
  NAND U5910 ( .A(n5053), .B(n5052), .Z(n5254) );
  XNOR U5911 ( .A(n5254), .B(n5255), .Z(n5256) );
  XNOR U5912 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U5913 ( .A(n5059), .B(n5058), .Z(n5063) );
  NAND U5914 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U5915 ( .A(n5063), .B(n5062), .Z(n5319) );
  NAND U5916 ( .A(n5065), .B(n5064), .Z(n5176) );
  NANDN U5917 ( .A(n5066), .B(n34044), .Z(n5068) );
  XOR U5918 ( .A(b[23]), .B(n15484), .Z(n5251) );
  OR U5919 ( .A(n5251), .B(n33867), .Z(n5067) );
  NAND U5920 ( .A(n5068), .B(n5067), .Z(n5175) );
  XNOR U5921 ( .A(n967), .B(a[40]), .Z(n5184) );
  NAND U5922 ( .A(n5184), .B(n28939), .Z(n5071) );
  NANDN U5923 ( .A(n5069), .B(n28938), .Z(n5070) );
  AND U5924 ( .A(n5071), .B(n5070), .Z(n5174) );
  XNOR U5925 ( .A(n5175), .B(n5174), .Z(n5177) );
  XNOR U5926 ( .A(n5176), .B(n5177), .Z(n5316) );
  XNOR U5927 ( .A(b[25]), .B(n14905), .Z(n5187) );
  NANDN U5928 ( .A(n34219), .B(n5187), .Z(n5074) );
  NAND U5929 ( .A(n34217), .B(n5072), .Z(n5073) );
  NAND U5930 ( .A(n5074), .B(n5073), .Z(n5277) );
  XOR U5931 ( .A(b[5]), .B(n20686), .Z(n5198) );
  OR U5932 ( .A(n5198), .B(n29363), .Z(n5077) );
  NANDN U5933 ( .A(n5075), .B(n29864), .Z(n5076) );
  NAND U5934 ( .A(n5077), .B(n5076), .Z(n5274) );
  XNOR U5935 ( .A(b[41]), .B(a[2]), .Z(n5219) );
  OR U5936 ( .A(n5219), .B(n36905), .Z(n5080) );
  NAND U5937 ( .A(n5078), .B(n36807), .Z(n5079) );
  AND U5938 ( .A(n5080), .B(n5079), .Z(n5275) );
  XNOR U5939 ( .A(n5274), .B(n5275), .Z(n5276) );
  XNOR U5940 ( .A(n5277), .B(n5276), .Z(n5317) );
  XNOR U5941 ( .A(n5316), .B(n5317), .Z(n5318) );
  XNOR U5942 ( .A(n5319), .B(n5318), .Z(n5266) );
  NANDN U5943 ( .A(n5082), .B(n5081), .Z(n5086) );
  NAND U5944 ( .A(n5084), .B(n5083), .Z(n5085) );
  NAND U5945 ( .A(n5086), .B(n5085), .Z(n5267) );
  XNOR U5946 ( .A(n5266), .B(n5267), .Z(n5268) );
  NANDN U5947 ( .A(n5088), .B(n5087), .Z(n5092) );
  NAND U5948 ( .A(n5090), .B(n5089), .Z(n5091) );
  NAND U5949 ( .A(n5092), .B(n5091), .Z(n5329) );
  NAND U5950 ( .A(n34848), .B(n5093), .Z(n5095) );
  XOR U5951 ( .A(n35375), .B(n14259), .Z(n5192) );
  NAND U5952 ( .A(n34618), .B(n5192), .Z(n5094) );
  NAND U5953 ( .A(n5095), .B(n5094), .Z(n5204) );
  XOR U5954 ( .A(n31123), .B(n19980), .Z(n5195) );
  NAND U5955 ( .A(n5195), .B(n29949), .Z(n5098) );
  NAND U5956 ( .A(n29948), .B(n5096), .Z(n5097) );
  NAND U5957 ( .A(n5098), .B(n5097), .Z(n5201) );
  XOR U5958 ( .A(b[37]), .B(n11406), .Z(n5283) );
  NANDN U5959 ( .A(n5283), .B(n36311), .Z(n5101) );
  NANDN U5960 ( .A(n5099), .B(n36309), .Z(n5100) );
  AND U5961 ( .A(n5101), .B(n5100), .Z(n5202) );
  XNOR U5962 ( .A(n5201), .B(n5202), .Z(n5203) );
  XOR U5963 ( .A(n5204), .B(n5203), .Z(n5312) );
  NAND U5964 ( .A(n35188), .B(n5102), .Z(n5104) );
  XOR U5965 ( .A(n35540), .B(n14210), .Z(n5289) );
  NANDN U5966 ( .A(n34968), .B(n5289), .Z(n5103) );
  NAND U5967 ( .A(n5104), .B(n5103), .Z(n5301) );
  XOR U5968 ( .A(b[11]), .B(n18841), .Z(n5292) );
  OR U5969 ( .A(n5292), .B(n31369), .Z(n5107) );
  NANDN U5970 ( .A(n5105), .B(n31119), .Z(n5106) );
  NAND U5971 ( .A(n5107), .B(n5106), .Z(n5298) );
  XOR U5972 ( .A(b[9]), .B(n19513), .Z(n5295) );
  NANDN U5973 ( .A(n5295), .B(n30509), .Z(n5110) );
  NANDN U5974 ( .A(n5108), .B(n30846), .Z(n5109) );
  AND U5975 ( .A(n5110), .B(n5109), .Z(n5299) );
  XNOR U5976 ( .A(n5298), .B(n5299), .Z(n5300) );
  XOR U5977 ( .A(n5301), .B(n5300), .Z(n5310) );
  NANDN U5978 ( .A(n5111), .B(n32011), .Z(n5113) );
  XNOR U5979 ( .A(n972), .B(a[28]), .Z(n5242) );
  NANDN U5980 ( .A(n32010), .B(n5242), .Z(n5112) );
  AND U5981 ( .A(n5113), .B(n5112), .Z(n5215) );
  XNOR U5982 ( .A(b[17]), .B(n17133), .Z(n5233) );
  NAND U5983 ( .A(n5233), .B(n32543), .Z(n5116) );
  NANDN U5984 ( .A(n5114), .B(n32541), .Z(n5115) );
  AND U5985 ( .A(n5116), .B(n5115), .Z(n5214) );
  NANDN U5986 ( .A(n5117), .B(n35311), .Z(n5119) );
  XNOR U5987 ( .A(n973), .B(a[12]), .Z(n5236) );
  NAND U5988 ( .A(n5236), .B(n35313), .Z(n5118) );
  AND U5989 ( .A(n5119), .B(n5118), .Z(n5213) );
  XNOR U5990 ( .A(n5214), .B(n5213), .Z(n5216) );
  XNOR U5991 ( .A(n5215), .B(n5216), .Z(n5307) );
  XNOR U5992 ( .A(b[21]), .B(a[22]), .Z(n5230) );
  OR U5993 ( .A(n5230), .B(n33634), .Z(n5122) );
  NANDN U5994 ( .A(n5120), .B(n33464), .Z(n5121) );
  NAND U5995 ( .A(n5122), .B(n5121), .Z(n5305) );
  NANDN U5996 ( .A(n5123), .B(n33283), .Z(n5125) );
  XNOR U5997 ( .A(n33020), .B(a[24]), .Z(n5239) );
  NANDN U5998 ( .A(n33021), .B(n5239), .Z(n5124) );
  AND U5999 ( .A(n5125), .B(n5124), .Z(n5304) );
  XNOR U6000 ( .A(n5305), .B(n5304), .Z(n5306) );
  XNOR U6001 ( .A(n5307), .B(n5306), .Z(n5311) );
  XNOR U6002 ( .A(n5310), .B(n5311), .Z(n5313) );
  XNOR U6003 ( .A(n5312), .B(n5313), .Z(n5327) );
  NANDN U6004 ( .A(n5127), .B(n5126), .Z(n5131) );
  NAND U6005 ( .A(n5129), .B(n5128), .Z(n5130) );
  AND U6006 ( .A(n5131), .B(n5130), .Z(n5326) );
  XNOR U6007 ( .A(n5327), .B(n5326), .Z(n5328) );
  XOR U6008 ( .A(n5329), .B(n5328), .Z(n5269) );
  XOR U6009 ( .A(n5268), .B(n5269), .Z(n5260) );
  XNOR U6010 ( .A(n5261), .B(n5260), .Z(n5262) );
  XNOR U6011 ( .A(n5263), .B(n5262), .Z(n5157) );
  XNOR U6012 ( .A(n5156), .B(n5157), .Z(n5158) );
  XOR U6013 ( .A(n5159), .B(n5158), .Z(n5150) );
  NANDN U6014 ( .A(n5133), .B(n5132), .Z(n5137) );
  NAND U6015 ( .A(n5135), .B(n5134), .Z(n5136) );
  AND U6016 ( .A(n5137), .B(n5136), .Z(n5151) );
  XNOR U6017 ( .A(n5150), .B(n5151), .Z(n5152) );
  XNOR U6018 ( .A(n5153), .B(n5152), .Z(n5144) );
  NANDN U6019 ( .A(n5139), .B(n5138), .Z(n5143) );
  OR U6020 ( .A(n5141), .B(n5140), .Z(n5142) );
  AND U6021 ( .A(n5143), .B(n5142), .Z(n5145) );
  XNOR U6022 ( .A(n5144), .B(n5145), .Z(n5146) );
  XOR U6023 ( .A(n5147), .B(n5146), .Z(n5333) );
  XOR U6024 ( .A(n5334), .B(n5333), .Z(c[106]) );
  NANDN U6025 ( .A(n5145), .B(n5144), .Z(n5149) );
  NAND U6026 ( .A(n5147), .B(n5146), .Z(n5148) );
  NAND U6027 ( .A(n5149), .B(n5148), .Z(n5345) );
  NANDN U6028 ( .A(n5151), .B(n5150), .Z(n5155) );
  NAND U6029 ( .A(n5153), .B(n5152), .Z(n5154) );
  NAND U6030 ( .A(n5155), .B(n5154), .Z(n5343) );
  NANDN U6031 ( .A(n5157), .B(n5156), .Z(n5161) );
  NANDN U6032 ( .A(n5159), .B(n5158), .Z(n5160) );
  NAND U6033 ( .A(n5161), .B(n5160), .Z(n5346) );
  OR U6034 ( .A(n5163), .B(n5162), .Z(n5167) );
  NANDN U6035 ( .A(n5165), .B(n5164), .Z(n5166) );
  AND U6036 ( .A(n5167), .B(n5166), .Z(n5347) );
  XNOR U6037 ( .A(n5346), .B(n5347), .Z(n5348) );
  OR U6038 ( .A(n5169), .B(n5168), .Z(n5173) );
  NAND U6039 ( .A(n5171), .B(n5170), .Z(n5172) );
  NAND U6040 ( .A(n5173), .B(n5172), .Z(n5359) );
  NANDN U6041 ( .A(n5179), .B(n5178), .Z(n5183) );
  NAND U6042 ( .A(n5181), .B(n5180), .Z(n5182) );
  AND U6043 ( .A(n5183), .B(n5182), .Z(n5381) );
  XOR U6044 ( .A(b[3]), .B(n21441), .Z(n5484) );
  NANDN U6045 ( .A(n5484), .B(n28939), .Z(n5186) );
  NAND U6046 ( .A(n5184), .B(n28938), .Z(n5185) );
  NAND U6047 ( .A(n5186), .B(n5185), .Z(n5434) );
  XNOR U6048 ( .A(b[25]), .B(n15113), .Z(n5410) );
  NANDN U6049 ( .A(n34219), .B(n5410), .Z(n5189) );
  NAND U6050 ( .A(n34217), .B(n5187), .Z(n5188) );
  AND U6051 ( .A(n5189), .B(n5188), .Z(n5435) );
  XNOR U6052 ( .A(n5434), .B(n5435), .Z(n5436) );
  OR U6053 ( .A(b[41]), .B(b[42]), .Z(n5190) );
  NANDN U6054 ( .A(n986), .B(n5190), .Z(n5191) );
  NAND U6055 ( .A(b[42]), .B(b[41]), .Z(n37134) );
  NAND U6056 ( .A(b[43]), .B(n37134), .Z(n37365) );
  ANDN U6057 ( .B(n5191), .A(n37365), .Z(n5437) );
  XNOR U6058 ( .A(n5436), .B(n5437), .Z(n5380) );
  NAND U6059 ( .A(n34848), .B(n5192), .Z(n5194) );
  XOR U6060 ( .A(n35375), .B(n14514), .Z(n5386) );
  NAND U6061 ( .A(n34618), .B(n5386), .Z(n5193) );
  NAND U6062 ( .A(n5194), .B(n5193), .Z(n5470) );
  XOR U6063 ( .A(n31123), .B(n20352), .Z(n5493) );
  NAND U6064 ( .A(n5493), .B(n29949), .Z(n5197) );
  NAND U6065 ( .A(n29948), .B(n5195), .Z(n5196) );
  NAND U6066 ( .A(n5197), .B(n5196), .Z(n5467) );
  XOR U6067 ( .A(b[5]), .B(n20867), .Z(n5389) );
  OR U6068 ( .A(n5389), .B(n29363), .Z(n5200) );
  NANDN U6069 ( .A(n5198), .B(n29864), .Z(n5199) );
  AND U6070 ( .A(n5200), .B(n5199), .Z(n5468) );
  XNOR U6071 ( .A(n5467), .B(n5468), .Z(n5469) );
  XNOR U6072 ( .A(n5470), .B(n5469), .Z(n5382) );
  XOR U6073 ( .A(n5383), .B(n5382), .Z(n5508) );
  NANDN U6074 ( .A(n5202), .B(n5201), .Z(n5206) );
  NAND U6075 ( .A(n5204), .B(n5203), .Z(n5205) );
  NAND U6076 ( .A(n5206), .B(n5205), .Z(n5509) );
  XOR U6077 ( .A(n5508), .B(n5509), .Z(n5510) );
  XNOR U6078 ( .A(n5511), .B(n5510), .Z(n5373) );
  NANDN U6079 ( .A(n5208), .B(n5207), .Z(n5212) );
  NAND U6080 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U6081 ( .A(n5212), .B(n5211), .Z(n5503) );
  OR U6082 ( .A(n5214), .B(n5213), .Z(n5218) );
  OR U6083 ( .A(n5216), .B(n5215), .Z(n5217) );
  AND U6084 ( .A(n5218), .B(n5217), .Z(n5502) );
  XNOR U6085 ( .A(n5503), .B(n5502), .Z(n5504) );
  XNOR U6086 ( .A(b[41]), .B(a[3]), .Z(n5458) );
  OR U6087 ( .A(n5458), .B(n36905), .Z(n5221) );
  NANDN U6088 ( .A(n5219), .B(n36807), .Z(n5220) );
  NAND U6089 ( .A(n5221), .B(n5220), .Z(n5480) );
  XNOR U6090 ( .A(n977), .B(a[0]), .Z(n5224) );
  XNOR U6091 ( .A(n977), .B(b[41]), .Z(n5223) );
  XNOR U6092 ( .A(n977), .B(b[42]), .Z(n5222) );
  AND U6093 ( .A(n5223), .B(n5222), .Z(n37069) );
  NAND U6094 ( .A(n5224), .B(n37069), .Z(n5226) );
  XNOR U6095 ( .A(n977), .B(a[1]), .Z(n5392) );
  NAND U6096 ( .A(n5392), .B(n37068), .Z(n5225) );
  NAND U6097 ( .A(n5226), .B(n5225), .Z(n5479) );
  XNOR U6098 ( .A(n5480), .B(n5479), .Z(n5464) );
  NANDN U6099 ( .A(n966), .B(a[43]), .Z(n5227) );
  XOR U6100 ( .A(n29232), .B(n5227), .Z(n5229) );
  IV U6101 ( .A(a[42]), .Z(n22246) );
  NANDN U6102 ( .A(n22246), .B(n966), .Z(n5228) );
  AND U6103 ( .A(n5229), .B(n5228), .Z(n5462) );
  XNOR U6104 ( .A(b[21]), .B(n16269), .Z(n5395) );
  NANDN U6105 ( .A(n33634), .B(n5395), .Z(n5232) );
  NANDN U6106 ( .A(n5230), .B(n33464), .Z(n5231) );
  AND U6107 ( .A(n5232), .B(n5231), .Z(n5461) );
  XNOR U6108 ( .A(n5462), .B(n5461), .Z(n5463) );
  XOR U6109 ( .A(n5464), .B(n5463), .Z(n5505) );
  XNOR U6110 ( .A(n5504), .B(n5505), .Z(n5370) );
  XNOR U6111 ( .A(b[17]), .B(a[27]), .Z(n5446) );
  NANDN U6112 ( .A(n5446), .B(n32543), .Z(n5235) );
  NAND U6113 ( .A(n5233), .B(n32541), .Z(n5234) );
  NAND U6114 ( .A(n5235), .B(n5234), .Z(n5443) );
  XOR U6115 ( .A(b[31]), .B(n13509), .Z(n5398) );
  NANDN U6116 ( .A(n5398), .B(n35313), .Z(n5238) );
  NAND U6117 ( .A(n5236), .B(n35311), .Z(n5237) );
  NAND U6118 ( .A(n5238), .B(n5237), .Z(n5440) );
  NAND U6119 ( .A(n5239), .B(n33283), .Z(n5241) );
  XOR U6120 ( .A(n33020), .B(n16916), .Z(n5449) );
  NANDN U6121 ( .A(n33021), .B(n5449), .Z(n5240) );
  AND U6122 ( .A(n5241), .B(n5240), .Z(n5441) );
  XNOR U6123 ( .A(n5440), .B(n5441), .Z(n5442) );
  XNOR U6124 ( .A(n5443), .B(n5442), .Z(n5499) );
  XOR U6125 ( .A(b[15]), .B(n18003), .Z(n5452) );
  OR U6126 ( .A(n5452), .B(n32010), .Z(n5244) );
  NAND U6127 ( .A(n5242), .B(n32011), .Z(n5243) );
  NAND U6128 ( .A(n5244), .B(n5243), .Z(n5407) );
  XOR U6129 ( .A(b[33]), .B(n12830), .Z(n5419) );
  NANDN U6130 ( .A(n5419), .B(n35620), .Z(n5247) );
  NANDN U6131 ( .A(n5245), .B(n35621), .Z(n5246) );
  NAND U6132 ( .A(n5247), .B(n5246), .Z(n5404) );
  XNOR U6133 ( .A(b[35]), .B(a[9]), .Z(n5422) );
  NANDN U6134 ( .A(n5422), .B(n35985), .Z(n5250) );
  NANDN U6135 ( .A(n5248), .B(n35986), .Z(n5249) );
  AND U6136 ( .A(n5250), .B(n5249), .Z(n5405) );
  XNOR U6137 ( .A(n5404), .B(n5405), .Z(n5406) );
  XNOR U6138 ( .A(n5407), .B(n5406), .Z(n5496) );
  NANDN U6139 ( .A(n5251), .B(n34044), .Z(n5253) );
  XOR U6140 ( .A(b[23]), .B(n16220), .Z(n5481) );
  OR U6141 ( .A(n5481), .B(n33867), .Z(n5252) );
  NAND U6142 ( .A(n5253), .B(n5252), .Z(n5497) );
  XNOR U6143 ( .A(n5496), .B(n5497), .Z(n5498) );
  XOR U6144 ( .A(n5499), .B(n5498), .Z(n5371) );
  XNOR U6145 ( .A(n5370), .B(n5371), .Z(n5372) );
  XOR U6146 ( .A(n5373), .B(n5372), .Z(n5358) );
  XNOR U6147 ( .A(n5359), .B(n5358), .Z(n5361) );
  NANDN U6148 ( .A(n5255), .B(n5254), .Z(n5259) );
  NAND U6149 ( .A(n5257), .B(n5256), .Z(n5258) );
  NAND U6150 ( .A(n5259), .B(n5258), .Z(n5360) );
  XNOR U6151 ( .A(n5361), .B(n5360), .Z(n5354) );
  NANDN U6152 ( .A(n5261), .B(n5260), .Z(n5265) );
  NAND U6153 ( .A(n5263), .B(n5262), .Z(n5264) );
  NAND U6154 ( .A(n5265), .B(n5264), .Z(n5353) );
  NANDN U6155 ( .A(n5275), .B(n5274), .Z(n5279) );
  NAND U6156 ( .A(n5277), .B(n5276), .Z(n5278) );
  NAND U6157 ( .A(n5279), .B(n5278), .Z(n5514) );
  XOR U6158 ( .A(b[39]), .B(n11202), .Z(n5490) );
  NANDN U6159 ( .A(n5490), .B(n36553), .Z(n5282) );
  NANDN U6160 ( .A(n5280), .B(n36643), .Z(n5281) );
  NAND U6161 ( .A(n5282), .B(n5281), .Z(n5476) );
  XOR U6162 ( .A(b[37]), .B(n11694), .Z(n5416) );
  NANDN U6163 ( .A(n5416), .B(n36311), .Z(n5285) );
  NANDN U6164 ( .A(n5283), .B(n36309), .Z(n5284) );
  NAND U6165 ( .A(n5285), .B(n5284), .Z(n5473) );
  XOR U6166 ( .A(b[13]), .B(n18639), .Z(n5401) );
  OR U6167 ( .A(n5401), .B(n31550), .Z(n5288) );
  NANDN U6168 ( .A(n5286), .B(n31874), .Z(n5287) );
  AND U6169 ( .A(n5288), .B(n5287), .Z(n5474) );
  XNOR U6170 ( .A(n5473), .B(n5474), .Z(n5475) );
  XOR U6171 ( .A(n5476), .B(n5475), .Z(n5374) );
  NAND U6172 ( .A(n35188), .B(n5289), .Z(n5291) );
  XOR U6173 ( .A(n35540), .B(n13976), .Z(n5487) );
  NANDN U6174 ( .A(n34968), .B(n5487), .Z(n5290) );
  NAND U6175 ( .A(n5291), .B(n5290), .Z(n5431) );
  XOR U6176 ( .A(b[11]), .B(n19656), .Z(n5425) );
  OR U6177 ( .A(n5425), .B(n31369), .Z(n5294) );
  NANDN U6178 ( .A(n5292), .B(n31119), .Z(n5293) );
  NAND U6179 ( .A(n5294), .B(n5293), .Z(n5428) );
  XOR U6180 ( .A(b[9]), .B(n20315), .Z(n5413) );
  NANDN U6181 ( .A(n5413), .B(n30509), .Z(n5297) );
  NANDN U6182 ( .A(n5295), .B(n30846), .Z(n5296) );
  AND U6183 ( .A(n5297), .B(n5296), .Z(n5429) );
  XNOR U6184 ( .A(n5428), .B(n5429), .Z(n5430) );
  XOR U6185 ( .A(n5431), .B(n5430), .Z(n5375) );
  XNOR U6186 ( .A(n5374), .B(n5375), .Z(n5377) );
  NANDN U6187 ( .A(n5299), .B(n5298), .Z(n5303) );
  NAND U6188 ( .A(n5301), .B(n5300), .Z(n5302) );
  NAND U6189 ( .A(n5303), .B(n5302), .Z(n5376) );
  XOR U6190 ( .A(n5377), .B(n5376), .Z(n5515) );
  XNOR U6191 ( .A(n5514), .B(n5515), .Z(n5516) );
  NANDN U6192 ( .A(n5305), .B(n5304), .Z(n5309) );
  NAND U6193 ( .A(n5307), .B(n5306), .Z(n5308) );
  AND U6194 ( .A(n5309), .B(n5308), .Z(n5517) );
  XOR U6195 ( .A(n5516), .B(n5517), .Z(n5365) );
  OR U6196 ( .A(n5311), .B(n5310), .Z(n5315) );
  OR U6197 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U6198 ( .A(n5315), .B(n5314), .Z(n5364) );
  XOR U6199 ( .A(n5365), .B(n5364), .Z(n5366) );
  XNOR U6200 ( .A(n5367), .B(n5366), .Z(n5527) );
  XNOR U6201 ( .A(n5526), .B(n5527), .Z(n5528) );
  NANDN U6202 ( .A(n5321), .B(n5320), .Z(n5325) );
  NAND U6203 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U6204 ( .A(n5325), .B(n5324), .Z(n5520) );
  NANDN U6205 ( .A(n5327), .B(n5326), .Z(n5331) );
  NAND U6206 ( .A(n5329), .B(n5328), .Z(n5330) );
  AND U6207 ( .A(n5331), .B(n5330), .Z(n5521) );
  XNOR U6208 ( .A(n5520), .B(n5521), .Z(n5522) );
  XOR U6209 ( .A(n5523), .B(n5522), .Z(n5529) );
  XNOR U6210 ( .A(n5528), .B(n5529), .Z(n5352) );
  XNOR U6211 ( .A(n5353), .B(n5352), .Z(n5355) );
  XNOR U6212 ( .A(n5354), .B(n5355), .Z(n5349) );
  XOR U6213 ( .A(n5348), .B(n5349), .Z(n5342) );
  XNOR U6214 ( .A(n5343), .B(n5342), .Z(n5344) );
  XNOR U6215 ( .A(n5345), .B(n5344), .Z(n5337) );
  XNOR U6216 ( .A(n5337), .B(sreg[107]), .Z(n5339) );
  NAND U6217 ( .A(n5332), .B(sreg[106]), .Z(n5336) );
  OR U6218 ( .A(n5334), .B(n5333), .Z(n5335) );
  AND U6219 ( .A(n5336), .B(n5335), .Z(n5338) );
  XOR U6220 ( .A(n5339), .B(n5338), .Z(c[107]) );
  NAND U6221 ( .A(n5337), .B(sreg[107]), .Z(n5341) );
  OR U6222 ( .A(n5339), .B(n5338), .Z(n5340) );
  NAND U6223 ( .A(n5341), .B(n5340), .Z(n5733) );
  XNOR U6224 ( .A(n5733), .B(sreg[108]), .Z(n5735) );
  NANDN U6225 ( .A(n5347), .B(n5346), .Z(n5351) );
  NAND U6226 ( .A(n5349), .B(n5348), .Z(n5350) );
  NAND U6227 ( .A(n5351), .B(n5350), .Z(n5532) );
  NAND U6228 ( .A(n5353), .B(n5352), .Z(n5357) );
  NANDN U6229 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U6230 ( .A(n5357), .B(n5356), .Z(n5730) );
  NAND U6231 ( .A(n5359), .B(n5358), .Z(n5363) );
  OR U6232 ( .A(n5361), .B(n5360), .Z(n5362) );
  NAND U6233 ( .A(n5363), .B(n5362), .Z(n5727) );
  NANDN U6234 ( .A(n5365), .B(n5364), .Z(n5369) );
  OR U6235 ( .A(n5367), .B(n5366), .Z(n5368) );
  NAND U6236 ( .A(n5369), .B(n5368), .Z(n5721) );
  OR U6237 ( .A(n5375), .B(n5374), .Z(n5379) );
  OR U6238 ( .A(n5377), .B(n5376), .Z(n5378) );
  NAND U6239 ( .A(n5379), .B(n5378), .Z(n5612) );
  OR U6240 ( .A(n5381), .B(n5380), .Z(n5385) );
  OR U6241 ( .A(n5383), .B(n5382), .Z(n5384) );
  AND U6242 ( .A(n5385), .B(n5384), .Z(n5611) );
  XOR U6243 ( .A(n5612), .B(n5611), .Z(n5613) );
  NAND U6244 ( .A(n34848), .B(n5386), .Z(n5388) );
  XOR U6245 ( .A(n35375), .B(n14905), .Z(n5673) );
  NAND U6246 ( .A(n34618), .B(n5673), .Z(n5387) );
  NAND U6247 ( .A(n5388), .B(n5387), .Z(n5563) );
  XOR U6248 ( .A(b[5]), .B(n21149), .Z(n5688) );
  OR U6249 ( .A(n5688), .B(n29363), .Z(n5391) );
  NANDN U6250 ( .A(n5389), .B(n29864), .Z(n5390) );
  NAND U6251 ( .A(n5391), .B(n5390), .Z(n5560) );
  XOR U6252 ( .A(b[43]), .B(n10363), .Z(n5575) );
  NANDN U6253 ( .A(n5575), .B(n37068), .Z(n5394) );
  NAND U6254 ( .A(n5392), .B(n37069), .Z(n5393) );
  AND U6255 ( .A(n5394), .B(n5393), .Z(n5561) );
  XNOR U6256 ( .A(n5560), .B(n5561), .Z(n5562) );
  XNOR U6257 ( .A(n5563), .B(n5562), .Z(n5592) );
  XNOR U6258 ( .A(b[21]), .B(a[24]), .Z(n5682) );
  OR U6259 ( .A(n5682), .B(n33634), .Z(n5397) );
  NAND U6260 ( .A(n5395), .B(n33464), .Z(n5396) );
  NAND U6261 ( .A(n5397), .B(n5396), .Z(n5670) );
  XOR U6262 ( .A(b[31]), .B(n14210), .Z(n5641) );
  NANDN U6263 ( .A(n5641), .B(n35313), .Z(n5400) );
  NANDN U6264 ( .A(n5398), .B(n35311), .Z(n5399) );
  NAND U6265 ( .A(n5400), .B(n5399), .Z(n5667) );
  XOR U6266 ( .A(b[13]), .B(n18841), .Z(n5566) );
  OR U6267 ( .A(n5566), .B(n31550), .Z(n5403) );
  NANDN U6268 ( .A(n5401), .B(n31874), .Z(n5402) );
  AND U6269 ( .A(n5403), .B(n5402), .Z(n5668) );
  XNOR U6270 ( .A(n5667), .B(n5668), .Z(n5669) );
  XNOR U6271 ( .A(n5670), .B(n5669), .Z(n5589) );
  NANDN U6272 ( .A(n5405), .B(n5404), .Z(n5409) );
  NAND U6273 ( .A(n5407), .B(n5406), .Z(n5408) );
  NAND U6274 ( .A(n5409), .B(n5408), .Z(n5590) );
  XNOR U6275 ( .A(n5589), .B(n5590), .Z(n5591) );
  XOR U6276 ( .A(n5592), .B(n5591), .Z(n5601) );
  XNOR U6277 ( .A(b[25]), .B(a[20]), .Z(n5664) );
  OR U6278 ( .A(n5664), .B(n34219), .Z(n5412) );
  NAND U6279 ( .A(n34217), .B(n5410), .Z(n5411) );
  NAND U6280 ( .A(n5412), .B(n5411), .Z(n5694) );
  XOR U6281 ( .A(b[9]), .B(n19980), .Z(n5638) );
  NANDN U6282 ( .A(n5638), .B(n30509), .Z(n5415) );
  NANDN U6283 ( .A(n5413), .B(n30846), .Z(n5414) );
  NAND U6284 ( .A(n5415), .B(n5414), .Z(n5691) );
  XOR U6285 ( .A(b[37]), .B(n11986), .Z(n5572) );
  NANDN U6286 ( .A(n5572), .B(n36311), .Z(n5418) );
  NANDN U6287 ( .A(n5416), .B(n36309), .Z(n5417) );
  AND U6288 ( .A(n5418), .B(n5417), .Z(n5692) );
  XNOR U6289 ( .A(n5691), .B(n5692), .Z(n5693) );
  XNOR U6290 ( .A(n5694), .B(n5693), .Z(n5617) );
  XOR U6291 ( .A(b[33]), .B(n13106), .Z(n5650) );
  NANDN U6292 ( .A(n5650), .B(n35620), .Z(n5421) );
  NANDN U6293 ( .A(n5419), .B(n35621), .Z(n5420) );
  NAND U6294 ( .A(n5421), .B(n5420), .Z(n5557) );
  XNOR U6295 ( .A(b[35]), .B(a[10]), .Z(n5569) );
  NANDN U6296 ( .A(n5569), .B(n35985), .Z(n5424) );
  NANDN U6297 ( .A(n5422), .B(n35986), .Z(n5423) );
  NAND U6298 ( .A(n5424), .B(n5423), .Z(n5554) );
  XOR U6299 ( .A(b[11]), .B(n19513), .Z(n5635) );
  OR U6300 ( .A(n5635), .B(n31369), .Z(n5427) );
  NANDN U6301 ( .A(n5425), .B(n31119), .Z(n5426) );
  AND U6302 ( .A(n5427), .B(n5426), .Z(n5555) );
  XNOR U6303 ( .A(n5554), .B(n5555), .Z(n5556) );
  XOR U6304 ( .A(n5557), .B(n5556), .Z(n5618) );
  XNOR U6305 ( .A(n5617), .B(n5618), .Z(n5619) );
  NANDN U6306 ( .A(n5429), .B(n5428), .Z(n5433) );
  NAND U6307 ( .A(n5431), .B(n5430), .Z(n5432) );
  AND U6308 ( .A(n5433), .B(n5432), .Z(n5620) );
  XNOR U6309 ( .A(n5619), .B(n5620), .Z(n5600) );
  NANDN U6310 ( .A(n5435), .B(n5434), .Z(n5439) );
  NAND U6311 ( .A(n5437), .B(n5436), .Z(n5438) );
  AND U6312 ( .A(n5439), .B(n5438), .Z(n5599) );
  XNOR U6313 ( .A(n5600), .B(n5599), .Z(n5602) );
  XOR U6314 ( .A(n5601), .B(n5602), .Z(n5614) );
  XNOR U6315 ( .A(n5613), .B(n5614), .Z(n5545) );
  NANDN U6316 ( .A(n5441), .B(n5440), .Z(n5445) );
  NAND U6317 ( .A(n5443), .B(n5442), .Z(n5444) );
  AND U6318 ( .A(n5445), .B(n5444), .Z(n5712) );
  XNOR U6319 ( .A(b[17]), .B(a[28]), .Z(n5647) );
  NANDN U6320 ( .A(n5647), .B(n32543), .Z(n5448) );
  NANDN U6321 ( .A(n5446), .B(n32541), .Z(n5447) );
  NAND U6322 ( .A(n5448), .B(n5447), .Z(n5632) );
  NAND U6323 ( .A(n33283), .B(n5449), .Z(n5451) );
  XOR U6324 ( .A(b[19]), .B(n17133), .Z(n5656) );
  OR U6325 ( .A(n5656), .B(n33021), .Z(n5450) );
  NAND U6326 ( .A(n5451), .B(n5450), .Z(n5629) );
  XOR U6327 ( .A(b[15]), .B(n18804), .Z(n5644) );
  OR U6328 ( .A(n5644), .B(n32010), .Z(n5454) );
  NANDN U6329 ( .A(n5452), .B(n32011), .Z(n5453) );
  AND U6330 ( .A(n5454), .B(n5453), .Z(n5630) );
  XNOR U6331 ( .A(n5629), .B(n5630), .Z(n5631) );
  XNOR U6332 ( .A(n5632), .B(n5631), .Z(n5710) );
  NANDN U6333 ( .A(n966), .B(a[44]), .Z(n5455) );
  XOR U6334 ( .A(n29232), .B(n5455), .Z(n5457) );
  IV U6335 ( .A(a[43]), .Z(n21996) );
  NANDN U6336 ( .A(n21996), .B(n966), .Z(n5456) );
  AND U6337 ( .A(n5457), .B(n5456), .Z(n5625) );
  XNOR U6338 ( .A(b[41]), .B(n10854), .Z(n5661) );
  NANDN U6339 ( .A(n36905), .B(n5661), .Z(n5460) );
  NANDN U6340 ( .A(n5458), .B(n36807), .Z(n5459) );
  NAND U6341 ( .A(n5460), .B(n5459), .Z(n5623) );
  XNOR U6342 ( .A(n977), .B(b[44]), .Z(n37261) );
  NANDN U6343 ( .A(n986), .B(n37261), .Z(n5624) );
  XNOR U6344 ( .A(n5623), .B(n5624), .Z(n5626) );
  XOR U6345 ( .A(n5625), .B(n5626), .Z(n5709) );
  XNOR U6346 ( .A(n5710), .B(n5709), .Z(n5711) );
  XOR U6347 ( .A(n5712), .B(n5711), .Z(n5596) );
  NANDN U6348 ( .A(n5462), .B(n5461), .Z(n5466) );
  NAND U6349 ( .A(n5464), .B(n5463), .Z(n5465) );
  NAND U6350 ( .A(n5466), .B(n5465), .Z(n5593) );
  NANDN U6351 ( .A(n5468), .B(n5467), .Z(n5472) );
  NAND U6352 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U6353 ( .A(n5472), .B(n5471), .Z(n5594) );
  XNOR U6354 ( .A(n5593), .B(n5594), .Z(n5595) );
  XOR U6355 ( .A(n5596), .B(n5595), .Z(n5608) );
  NANDN U6356 ( .A(n5474), .B(n5473), .Z(n5478) );
  NAND U6357 ( .A(n5476), .B(n5475), .Z(n5477) );
  NAND U6358 ( .A(n5478), .B(n5477), .Z(n5706) );
  NAND U6359 ( .A(n5480), .B(n5479), .Z(n5552) );
  NANDN U6360 ( .A(n5481), .B(n34044), .Z(n5483) );
  XOR U6361 ( .A(b[23]), .B(n15963), .Z(n5586) );
  OR U6362 ( .A(n5586), .B(n33867), .Z(n5482) );
  NAND U6363 ( .A(n5483), .B(n5482), .Z(n5551) );
  XNOR U6364 ( .A(n967), .B(a[42]), .Z(n5676) );
  NAND U6365 ( .A(n5676), .B(n28939), .Z(n5486) );
  NANDN U6366 ( .A(n5484), .B(n28938), .Z(n5485) );
  AND U6367 ( .A(n5486), .B(n5485), .Z(n5550) );
  XNOR U6368 ( .A(n5551), .B(n5550), .Z(n5553) );
  XNOR U6369 ( .A(n5552), .B(n5553), .Z(n5703) );
  NAND U6370 ( .A(n35188), .B(n5487), .Z(n5489) );
  XOR U6371 ( .A(b[29]), .B(n14259), .Z(n5653) );
  OR U6372 ( .A(n5653), .B(n34968), .Z(n5488) );
  NAND U6373 ( .A(n5489), .B(n5488), .Z(n5700) );
  XOR U6374 ( .A(b[39]), .B(n11406), .Z(n5679) );
  NANDN U6375 ( .A(n5679), .B(n36553), .Z(n5492) );
  NANDN U6376 ( .A(n5490), .B(n36643), .Z(n5491) );
  NAND U6377 ( .A(n5492), .B(n5491), .Z(n5697) );
  XOR U6378 ( .A(n31123), .B(n20686), .Z(n5685) );
  NAND U6379 ( .A(n5685), .B(n29949), .Z(n5495) );
  NAND U6380 ( .A(n29948), .B(n5493), .Z(n5494) );
  AND U6381 ( .A(n5495), .B(n5494), .Z(n5698) );
  XNOR U6382 ( .A(n5697), .B(n5698), .Z(n5699) );
  XNOR U6383 ( .A(n5700), .B(n5699), .Z(n5704) );
  XNOR U6384 ( .A(n5703), .B(n5704), .Z(n5705) );
  XNOR U6385 ( .A(n5706), .B(n5705), .Z(n5606) );
  NANDN U6386 ( .A(n5497), .B(n5496), .Z(n5501) );
  NAND U6387 ( .A(n5499), .B(n5498), .Z(n5500) );
  AND U6388 ( .A(n5501), .B(n5500), .Z(n5605) );
  XNOR U6389 ( .A(n5606), .B(n5605), .Z(n5607) );
  XNOR U6390 ( .A(n5608), .B(n5607), .Z(n5544) );
  XOR U6391 ( .A(n5545), .B(n5544), .Z(n5546) );
  XOR U6392 ( .A(n5547), .B(n5546), .Z(n5722) );
  XNOR U6393 ( .A(n5721), .B(n5722), .Z(n5723) );
  NANDN U6394 ( .A(n5503), .B(n5502), .Z(n5507) );
  NAND U6395 ( .A(n5505), .B(n5504), .Z(n5506) );
  NAND U6396 ( .A(n5507), .B(n5506), .Z(n5541) );
  OR U6397 ( .A(n5509), .B(n5508), .Z(n5513) );
  NAND U6398 ( .A(n5511), .B(n5510), .Z(n5512) );
  NAND U6399 ( .A(n5513), .B(n5512), .Z(n5538) );
  NANDN U6400 ( .A(n5515), .B(n5514), .Z(n5519) );
  NAND U6401 ( .A(n5517), .B(n5516), .Z(n5518) );
  NAND U6402 ( .A(n5519), .B(n5518), .Z(n5539) );
  XNOR U6403 ( .A(n5538), .B(n5539), .Z(n5540) );
  XNOR U6404 ( .A(n5541), .B(n5540), .Z(n5724) );
  XOR U6405 ( .A(n5723), .B(n5724), .Z(n5718) );
  NANDN U6406 ( .A(n5521), .B(n5520), .Z(n5525) );
  NANDN U6407 ( .A(n5523), .B(n5522), .Z(n5524) );
  NAND U6408 ( .A(n5525), .B(n5524), .Z(n5715) );
  NANDN U6409 ( .A(n5527), .B(n5526), .Z(n5531) );
  NANDN U6410 ( .A(n5529), .B(n5528), .Z(n5530) );
  AND U6411 ( .A(n5531), .B(n5530), .Z(n5716) );
  XNOR U6412 ( .A(n5715), .B(n5716), .Z(n5717) );
  XOR U6413 ( .A(n5718), .B(n5717), .Z(n5728) );
  XOR U6414 ( .A(n5727), .B(n5728), .Z(n5729) );
  XNOR U6415 ( .A(n5730), .B(n5729), .Z(n5533) );
  XNOR U6416 ( .A(n5532), .B(n5533), .Z(n5534) );
  XOR U6417 ( .A(n5535), .B(n5534), .Z(n5734) );
  XOR U6418 ( .A(n5735), .B(n5734), .Z(c[108]) );
  NANDN U6419 ( .A(n5533), .B(n5532), .Z(n5537) );
  NAND U6420 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U6421 ( .A(n5537), .B(n5536), .Z(n5746) );
  NANDN U6422 ( .A(n5539), .B(n5538), .Z(n5543) );
  NAND U6423 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U6424 ( .A(n5543), .B(n5542), .Z(n5753) );
  OR U6425 ( .A(n5545), .B(n5544), .Z(n5549) );
  NANDN U6426 ( .A(n5547), .B(n5546), .Z(n5548) );
  AND U6427 ( .A(n5549), .B(n5548), .Z(n5754) );
  XNOR U6428 ( .A(n5753), .B(n5754), .Z(n5755) );
  NANDN U6429 ( .A(n5555), .B(n5554), .Z(n5559) );
  NAND U6430 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U6431 ( .A(n5559), .B(n5558), .Z(n5772) );
  XNOR U6432 ( .A(n5771), .B(n5772), .Z(n5773) );
  NANDN U6433 ( .A(n5561), .B(n5560), .Z(n5565) );
  NAND U6434 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U6435 ( .A(n5565), .B(n5564), .Z(n5897) );
  XOR U6436 ( .A(n971), .B(n19656), .Z(n5817) );
  NANDN U6437 ( .A(n31550), .B(n5817), .Z(n5568) );
  NANDN U6438 ( .A(n5566), .B(n31874), .Z(n5567) );
  NAND U6439 ( .A(n5568), .B(n5567), .Z(n5921) );
  XNOR U6440 ( .A(b[35]), .B(a[11]), .Z(n5903) );
  NANDN U6441 ( .A(n5903), .B(n35985), .Z(n5571) );
  NANDN U6442 ( .A(n5569), .B(n35986), .Z(n5570) );
  NAND U6443 ( .A(n5571), .B(n5570), .Z(n5918) );
  XOR U6444 ( .A(b[37]), .B(n12258), .Z(n5906) );
  NANDN U6445 ( .A(n5906), .B(n36311), .Z(n5574) );
  NANDN U6446 ( .A(n5572), .B(n36309), .Z(n5573) );
  AND U6447 ( .A(n5574), .B(n5573), .Z(n5919) );
  XNOR U6448 ( .A(n5918), .B(n5919), .Z(n5920) );
  XNOR U6449 ( .A(n5921), .B(n5920), .Z(n5895) );
  XOR U6450 ( .A(b[43]), .B(n10524), .Z(n5792) );
  NANDN U6451 ( .A(n5792), .B(n37068), .Z(n5577) );
  NANDN U6452 ( .A(n5575), .B(n37069), .Z(n5576) );
  NAND U6453 ( .A(n5577), .B(n5576), .Z(n5869) );
  XNOR U6454 ( .A(b[45]), .B(a[1]), .Z(n5870) );
  ANDN U6455 ( .B(n37261), .A(n5870), .Z(n5582) );
  XNOR U6456 ( .A(b[45]), .B(n986), .Z(n5580) );
  XNOR U6457 ( .A(b[45]), .B(n977), .Z(n5579) );
  XOR U6458 ( .A(b[45]), .B(b[44]), .Z(n5578) );
  AND U6459 ( .A(n5579), .B(n5578), .Z(n37262) );
  NAND U6460 ( .A(n5580), .B(n37262), .Z(n5581) );
  NANDN U6461 ( .A(n5582), .B(n5581), .Z(n5868) );
  XNOR U6462 ( .A(n5869), .B(n5868), .Z(n5885) );
  NANDN U6463 ( .A(n966), .B(a[45]), .Z(n5583) );
  XOR U6464 ( .A(n29232), .B(n5583), .Z(n5585) );
  IV U6465 ( .A(a[44]), .Z(n22289) );
  NANDN U6466 ( .A(n22289), .B(n966), .Z(n5584) );
  AND U6467 ( .A(n5585), .B(n5584), .Z(n5883) );
  NANDN U6468 ( .A(n5586), .B(n34044), .Z(n5588) );
  XNOR U6469 ( .A(n34510), .B(a[23]), .Z(n5909) );
  NANDN U6470 ( .A(n33867), .B(n5909), .Z(n5587) );
  AND U6471 ( .A(n5588), .B(n5587), .Z(n5882) );
  XNOR U6472 ( .A(n5883), .B(n5882), .Z(n5884) );
  XOR U6473 ( .A(n5885), .B(n5884), .Z(n5894) );
  XOR U6474 ( .A(n5895), .B(n5894), .Z(n5896) );
  XOR U6475 ( .A(n5897), .B(n5896), .Z(n5774) );
  XOR U6476 ( .A(n5773), .B(n5774), .Z(n5768) );
  NANDN U6477 ( .A(n5594), .B(n5593), .Z(n5598) );
  NAND U6478 ( .A(n5596), .B(n5595), .Z(n5597) );
  AND U6479 ( .A(n5598), .B(n5597), .Z(n5765) );
  XNOR U6480 ( .A(n5766), .B(n5765), .Z(n5767) );
  XNOR U6481 ( .A(n5768), .B(n5767), .Z(n5934) );
  NANDN U6482 ( .A(n5600), .B(n5599), .Z(n5604) );
  NAND U6483 ( .A(n5602), .B(n5601), .Z(n5603) );
  AND U6484 ( .A(n5604), .B(n5603), .Z(n5935) );
  XNOR U6485 ( .A(n5934), .B(n5935), .Z(n5936) );
  NANDN U6486 ( .A(n5606), .B(n5605), .Z(n5610) );
  NANDN U6487 ( .A(n5608), .B(n5607), .Z(n5609) );
  AND U6488 ( .A(n5610), .B(n5609), .Z(n5937) );
  XNOR U6489 ( .A(n5936), .B(n5937), .Z(n5762) );
  OR U6490 ( .A(n5612), .B(n5611), .Z(n5616) );
  NANDN U6491 ( .A(n5614), .B(n5613), .Z(n5615) );
  NAND U6492 ( .A(n5616), .B(n5615), .Z(n5760) );
  NANDN U6493 ( .A(n5618), .B(n5617), .Z(n5622) );
  NAND U6494 ( .A(n5620), .B(n5619), .Z(n5621) );
  NAND U6495 ( .A(n5622), .B(n5621), .Z(n5927) );
  NANDN U6496 ( .A(n5624), .B(n5623), .Z(n5628) );
  NAND U6497 ( .A(n5626), .B(n5625), .Z(n5627) );
  NAND U6498 ( .A(n5628), .B(n5627), .Z(n5848) );
  NANDN U6499 ( .A(n5630), .B(n5629), .Z(n5634) );
  NAND U6500 ( .A(n5632), .B(n5631), .Z(n5633) );
  AND U6501 ( .A(n5634), .B(n5633), .Z(n5847) );
  XNOR U6502 ( .A(n5848), .B(n5847), .Z(n5849) );
  XOR U6503 ( .A(b[11]), .B(n20315), .Z(n5900) );
  OR U6504 ( .A(n5900), .B(n31369), .Z(n5637) );
  NANDN U6505 ( .A(n5635), .B(n31119), .Z(n5636) );
  NAND U6506 ( .A(n5637), .B(n5636), .Z(n5786) );
  XOR U6507 ( .A(b[9]), .B(n20352), .Z(n5798) );
  NANDN U6508 ( .A(n5798), .B(n30509), .Z(n5640) );
  NANDN U6509 ( .A(n5638), .B(n30846), .Z(n5639) );
  NAND U6510 ( .A(n5640), .B(n5639), .Z(n5783) );
  XOR U6511 ( .A(b[31]), .B(n13976), .Z(n5820) );
  NANDN U6512 ( .A(n5820), .B(n35313), .Z(n5643) );
  NANDN U6513 ( .A(n5641), .B(n35311), .Z(n5642) );
  AND U6514 ( .A(n5643), .B(n5642), .Z(n5784) );
  XNOR U6515 ( .A(n5783), .B(n5784), .Z(n5785) );
  XNOR U6516 ( .A(n5786), .B(n5785), .Z(n5836) );
  XOR U6517 ( .A(n972), .B(n18639), .Z(n5814) );
  NANDN U6518 ( .A(n32010), .B(n5814), .Z(n5646) );
  NANDN U6519 ( .A(n5644), .B(n32011), .Z(n5645) );
  NAND U6520 ( .A(n5646), .B(n5645), .Z(n5879) );
  XNOR U6521 ( .A(b[17]), .B(n18003), .Z(n5811) );
  NAND U6522 ( .A(n5811), .B(n32543), .Z(n5649) );
  NANDN U6523 ( .A(n5647), .B(n32541), .Z(n5648) );
  NAND U6524 ( .A(n5649), .B(n5648), .Z(n5876) );
  XOR U6525 ( .A(n974), .B(n13509), .Z(n5823) );
  NAND U6526 ( .A(n35620), .B(n5823), .Z(n5652) );
  NANDN U6527 ( .A(n5650), .B(n35621), .Z(n5651) );
  AND U6528 ( .A(n5652), .B(n5651), .Z(n5877) );
  XNOR U6529 ( .A(n5876), .B(n5877), .Z(n5878) );
  XNOR U6530 ( .A(n5879), .B(n5878), .Z(n5780) );
  NANDN U6531 ( .A(n5653), .B(n35188), .Z(n5655) );
  XNOR U6532 ( .A(n35540), .B(a[17]), .Z(n5795) );
  NANDN U6533 ( .A(n34968), .B(n5795), .Z(n5654) );
  NAND U6534 ( .A(n5655), .B(n5654), .Z(n5778) );
  NANDN U6535 ( .A(n5656), .B(n33283), .Z(n5658) );
  XNOR U6536 ( .A(n33020), .B(a[27]), .Z(n5808) );
  NANDN U6537 ( .A(n33021), .B(n5808), .Z(n5657) );
  AND U6538 ( .A(n5658), .B(n5657), .Z(n5777) );
  XNOR U6539 ( .A(n5778), .B(n5777), .Z(n5779) );
  XOR U6540 ( .A(n5780), .B(n5779), .Z(n5835) );
  XOR U6541 ( .A(n5836), .B(n5835), .Z(n5837) );
  NANDN U6542 ( .A(n977), .B(b[44]), .Z(n37331) );
  NAND U6543 ( .A(n37331), .B(b[45]), .Z(n37570) );
  NOR U6544 ( .A(b[43]), .B(b[44]), .Z(n5659) );
  OR U6545 ( .A(n5659), .B(n986), .Z(n5660) );
  NANDN U6546 ( .A(n37570), .B(n5660), .Z(n5804) );
  NAND U6547 ( .A(n36807), .B(n5661), .Z(n5663) );
  XNOR U6548 ( .A(b[41]), .B(n11202), .Z(n5915) );
  NANDN U6549 ( .A(n36905), .B(n5915), .Z(n5662) );
  NAND U6550 ( .A(n5663), .B(n5662), .Z(n5805) );
  XNOR U6551 ( .A(n5804), .B(n5805), .Z(n5806) );
  XNOR U6552 ( .A(b[25]), .B(a[21]), .Z(n5873) );
  OR U6553 ( .A(n5873), .B(n34219), .Z(n5666) );
  NANDN U6554 ( .A(n5664), .B(n34217), .Z(n5665) );
  AND U6555 ( .A(n5666), .B(n5665), .Z(n5807) );
  XNOR U6556 ( .A(n5806), .B(n5807), .Z(n5838) );
  XNOR U6557 ( .A(n5837), .B(n5838), .Z(n5850) );
  XNOR U6558 ( .A(n5849), .B(n5850), .Z(n5924) );
  NANDN U6559 ( .A(n5668), .B(n5667), .Z(n5672) );
  NAND U6560 ( .A(n5670), .B(n5669), .Z(n5671) );
  NAND U6561 ( .A(n5672), .B(n5671), .Z(n5843) );
  NAND U6562 ( .A(n34848), .B(n5673), .Z(n5675) );
  XOR U6563 ( .A(n35375), .B(n15113), .Z(n5865) );
  NAND U6564 ( .A(n34618), .B(n5865), .Z(n5674) );
  NAND U6565 ( .A(n5675), .B(n5674), .Z(n5832) );
  XOR U6566 ( .A(n967), .B(n21996), .Z(n5912) );
  NAND U6567 ( .A(n5912), .B(n28939), .Z(n5678) );
  NAND U6568 ( .A(n5676), .B(n28938), .Z(n5677) );
  NAND U6569 ( .A(n5678), .B(n5677), .Z(n5829) );
  XOR U6570 ( .A(b[39]), .B(n11694), .Z(n5859) );
  NANDN U6571 ( .A(n5859), .B(n36553), .Z(n5681) );
  NANDN U6572 ( .A(n5679), .B(n36643), .Z(n5680) );
  AND U6573 ( .A(n5681), .B(n5680), .Z(n5830) );
  XNOR U6574 ( .A(n5829), .B(n5830), .Z(n5831) );
  XNOR U6575 ( .A(n5832), .B(n5831), .Z(n5841) );
  XNOR U6576 ( .A(b[21]), .B(a[25]), .Z(n5826) );
  OR U6577 ( .A(n5826), .B(n33634), .Z(n5684) );
  NANDN U6578 ( .A(n5682), .B(n33464), .Z(n5683) );
  NAND U6579 ( .A(n5684), .B(n5683), .Z(n5891) );
  XOR U6580 ( .A(n31123), .B(n20867), .Z(n5801) );
  NAND U6581 ( .A(n5801), .B(n29949), .Z(n5687) );
  NAND U6582 ( .A(n29948), .B(n5685), .Z(n5686) );
  NAND U6583 ( .A(n5687), .B(n5686), .Z(n5888) );
  XOR U6584 ( .A(b[5]), .B(n21441), .Z(n5862) );
  OR U6585 ( .A(n5862), .B(n29363), .Z(n5690) );
  NANDN U6586 ( .A(n5688), .B(n29864), .Z(n5689) );
  AND U6587 ( .A(n5690), .B(n5689), .Z(n5889) );
  XNOR U6588 ( .A(n5888), .B(n5889), .Z(n5890) );
  XOR U6589 ( .A(n5891), .B(n5890), .Z(n5842) );
  XOR U6590 ( .A(n5841), .B(n5842), .Z(n5844) );
  XNOR U6591 ( .A(n5843), .B(n5844), .Z(n5856) );
  NANDN U6592 ( .A(n5692), .B(n5691), .Z(n5696) );
  NAND U6593 ( .A(n5694), .B(n5693), .Z(n5695) );
  NAND U6594 ( .A(n5696), .B(n5695), .Z(n5853) );
  NANDN U6595 ( .A(n5698), .B(n5697), .Z(n5702) );
  NAND U6596 ( .A(n5700), .B(n5699), .Z(n5701) );
  AND U6597 ( .A(n5702), .B(n5701), .Z(n5854) );
  XNOR U6598 ( .A(n5853), .B(n5854), .Z(n5855) );
  XNOR U6599 ( .A(n5856), .B(n5855), .Z(n5925) );
  XNOR U6600 ( .A(n5924), .B(n5925), .Z(n5926) );
  XOR U6601 ( .A(n5927), .B(n5926), .Z(n5931) );
  NANDN U6602 ( .A(n5704), .B(n5703), .Z(n5708) );
  NAND U6603 ( .A(n5706), .B(n5705), .Z(n5707) );
  NAND U6604 ( .A(n5708), .B(n5707), .Z(n5929) );
  NANDN U6605 ( .A(n5710), .B(n5709), .Z(n5714) );
  NANDN U6606 ( .A(n5712), .B(n5711), .Z(n5713) );
  AND U6607 ( .A(n5714), .B(n5713), .Z(n5928) );
  XNOR U6608 ( .A(n5929), .B(n5928), .Z(n5930) );
  XNOR U6609 ( .A(n5931), .B(n5930), .Z(n5759) );
  XNOR U6610 ( .A(n5760), .B(n5759), .Z(n5761) );
  XNOR U6611 ( .A(n5762), .B(n5761), .Z(n5756) );
  XOR U6612 ( .A(n5755), .B(n5756), .Z(n5750) );
  NANDN U6613 ( .A(n5716), .B(n5715), .Z(n5720) );
  NANDN U6614 ( .A(n5718), .B(n5717), .Z(n5719) );
  NAND U6615 ( .A(n5720), .B(n5719), .Z(n5748) );
  NANDN U6616 ( .A(n5722), .B(n5721), .Z(n5726) );
  NANDN U6617 ( .A(n5724), .B(n5723), .Z(n5725) );
  AND U6618 ( .A(n5726), .B(n5725), .Z(n5747) );
  XNOR U6619 ( .A(n5748), .B(n5747), .Z(n5749) );
  XNOR U6620 ( .A(n5750), .B(n5749), .Z(n5743) );
  OR U6621 ( .A(n5728), .B(n5727), .Z(n5732) );
  NAND U6622 ( .A(n5730), .B(n5729), .Z(n5731) );
  AND U6623 ( .A(n5732), .B(n5731), .Z(n5744) );
  XNOR U6624 ( .A(n5743), .B(n5744), .Z(n5745) );
  XNOR U6625 ( .A(n5746), .B(n5745), .Z(n5738) );
  XNOR U6626 ( .A(n5738), .B(sreg[109]), .Z(n5740) );
  NAND U6627 ( .A(n5733), .B(sreg[108]), .Z(n5737) );
  OR U6628 ( .A(n5735), .B(n5734), .Z(n5736) );
  AND U6629 ( .A(n5737), .B(n5736), .Z(n5739) );
  XOR U6630 ( .A(n5740), .B(n5739), .Z(c[109]) );
  NAND U6631 ( .A(n5738), .B(sreg[109]), .Z(n5742) );
  OR U6632 ( .A(n5740), .B(n5739), .Z(n5741) );
  NAND U6633 ( .A(n5742), .B(n5741), .Z(n6153) );
  XNOR U6634 ( .A(n6153), .B(sreg[110]), .Z(n6155) );
  NANDN U6635 ( .A(n5748), .B(n5747), .Z(n5752) );
  NAND U6636 ( .A(n5750), .B(n5749), .Z(n5751) );
  NAND U6637 ( .A(n5752), .B(n5751), .Z(n5941) );
  NANDN U6638 ( .A(n5754), .B(n5753), .Z(n5758) );
  NANDN U6639 ( .A(n5756), .B(n5755), .Z(n5757) );
  NAND U6640 ( .A(n5758), .B(n5757), .Z(n5946) );
  OR U6641 ( .A(n5760), .B(n5759), .Z(n5764) );
  OR U6642 ( .A(n5762), .B(n5761), .Z(n5763) );
  AND U6643 ( .A(n5764), .B(n5763), .Z(n5947) );
  XNOR U6644 ( .A(n5946), .B(n5947), .Z(n5948) );
  NANDN U6645 ( .A(n5766), .B(n5765), .Z(n5770) );
  NAND U6646 ( .A(n5768), .B(n5767), .Z(n5769) );
  NAND U6647 ( .A(n5770), .B(n5769), .Z(n5961) );
  NANDN U6648 ( .A(n5772), .B(n5771), .Z(n5776) );
  NANDN U6649 ( .A(n5774), .B(n5773), .Z(n5775) );
  NAND U6650 ( .A(n5776), .B(n5775), .Z(n6148) );
  NANDN U6651 ( .A(n5778), .B(n5777), .Z(n5782) );
  NAND U6652 ( .A(n5780), .B(n5779), .Z(n5781) );
  NAND U6653 ( .A(n5782), .B(n5781), .Z(n6089) );
  NANDN U6654 ( .A(n5784), .B(n5783), .Z(n5788) );
  NAND U6655 ( .A(n5786), .B(n5785), .Z(n5787) );
  NAND U6656 ( .A(n5788), .B(n5787), .Z(n5979) );
  XOR U6657 ( .A(b[45]), .B(b[46]), .Z(n37471) );
  AND U6658 ( .A(n37471), .B(a[0]), .Z(n6032) );
  NANDN U6659 ( .A(n966), .B(a[46]), .Z(n5789) );
  XOR U6660 ( .A(n29232), .B(n5789), .Z(n5791) );
  IV U6661 ( .A(a[45]), .Z(n22579) );
  NANDN U6662 ( .A(n22579), .B(n966), .Z(n5790) );
  AND U6663 ( .A(n5791), .B(n5790), .Z(n6030) );
  NANDN U6664 ( .A(n5792), .B(n37069), .Z(n5794) );
  XNOR U6665 ( .A(n977), .B(a[4]), .Z(n6102) );
  NAND U6666 ( .A(n6102), .B(n37068), .Z(n5793) );
  AND U6667 ( .A(n5794), .B(n5793), .Z(n6029) );
  XNOR U6668 ( .A(n6030), .B(n6029), .Z(n6031) );
  XOR U6669 ( .A(n6032), .B(n6031), .Z(n5976) );
  NAND U6670 ( .A(n5795), .B(n35188), .Z(n5797) );
  XOR U6671 ( .A(n35540), .B(n14905), .Z(n6059) );
  NANDN U6672 ( .A(n34968), .B(n6059), .Z(n5796) );
  NAND U6673 ( .A(n5797), .B(n5796), .Z(n6056) );
  XOR U6674 ( .A(b[9]), .B(n20686), .Z(n6105) );
  NANDN U6675 ( .A(n6105), .B(n30509), .Z(n5800) );
  NANDN U6676 ( .A(n5798), .B(n30846), .Z(n5799) );
  NAND U6677 ( .A(n5800), .B(n5799), .Z(n6053) );
  XOR U6678 ( .A(n31123), .B(n21149), .Z(n6068) );
  NAND U6679 ( .A(n6068), .B(n29949), .Z(n5803) );
  NAND U6680 ( .A(n29948), .B(n5801), .Z(n5802) );
  AND U6681 ( .A(n5803), .B(n5802), .Z(n6054) );
  XNOR U6682 ( .A(n6053), .B(n6054), .Z(n6055) );
  XNOR U6683 ( .A(n6056), .B(n6055), .Z(n5977) );
  XNOR U6684 ( .A(n5976), .B(n5977), .Z(n5978) );
  XOR U6685 ( .A(n5979), .B(n5978), .Z(n6090) );
  XNOR U6686 ( .A(n6089), .B(n6090), .Z(n6091) );
  NAND U6687 ( .A(n5808), .B(n33283), .Z(n5810) );
  XOR U6688 ( .A(n33020), .B(n17702), .Z(n6020) );
  NANDN U6689 ( .A(n33021), .B(n6020), .Z(n5809) );
  NAND U6690 ( .A(n5810), .B(n5809), .Z(n6082) );
  XNOR U6691 ( .A(b[17]), .B(a[30]), .Z(n6014) );
  NANDN U6692 ( .A(n6014), .B(n32543), .Z(n5813) );
  NAND U6693 ( .A(n5811), .B(n32541), .Z(n5812) );
  NAND U6694 ( .A(n5813), .B(n5812), .Z(n6079) );
  XOR U6695 ( .A(b[15]), .B(n18841), .Z(n6108) );
  OR U6696 ( .A(n6108), .B(n32010), .Z(n5816) );
  NAND U6697 ( .A(n5814), .B(n32011), .Z(n5815) );
  AND U6698 ( .A(n5816), .B(n5815), .Z(n6080) );
  XNOR U6699 ( .A(n6079), .B(n6080), .Z(n6081) );
  XNOR U6700 ( .A(n6082), .B(n6081), .Z(n6098) );
  XOR U6701 ( .A(b[13]), .B(n19513), .Z(n6035) );
  OR U6702 ( .A(n6035), .B(n31550), .Z(n5819) );
  NAND U6703 ( .A(n5817), .B(n31874), .Z(n5818) );
  NAND U6704 ( .A(n5819), .B(n5818), .Z(n5997) );
  XOR U6705 ( .A(b[31]), .B(n14259), .Z(n6076) );
  NANDN U6706 ( .A(n6076), .B(n35313), .Z(n5822) );
  NANDN U6707 ( .A(n5820), .B(n35311), .Z(n5821) );
  NAND U6708 ( .A(n5822), .B(n5821), .Z(n5994) );
  XOR U6709 ( .A(b[33]), .B(n14210), .Z(n6099) );
  NANDN U6710 ( .A(n6099), .B(n35620), .Z(n5825) );
  NAND U6711 ( .A(n5823), .B(n35621), .Z(n5824) );
  AND U6712 ( .A(n5825), .B(n5824), .Z(n5995) );
  XNOR U6713 ( .A(n5994), .B(n5995), .Z(n5996) );
  XNOR U6714 ( .A(n5997), .B(n5996), .Z(n6095) );
  XNOR U6715 ( .A(b[21]), .B(n17133), .Z(n6017) );
  NANDN U6716 ( .A(n33634), .B(n6017), .Z(n5828) );
  NANDN U6717 ( .A(n5826), .B(n33464), .Z(n5827) );
  NAND U6718 ( .A(n5828), .B(n5827), .Z(n6096) );
  XNOR U6719 ( .A(n6095), .B(n6096), .Z(n6097) );
  XOR U6720 ( .A(n6098), .B(n6097), .Z(n6135) );
  NANDN U6721 ( .A(n5830), .B(n5829), .Z(n5834) );
  NAND U6722 ( .A(n5832), .B(n5831), .Z(n5833) );
  AND U6723 ( .A(n5834), .B(n5833), .Z(n6136) );
  XNOR U6724 ( .A(n6135), .B(n6136), .Z(n6138) );
  XNOR U6725 ( .A(n6137), .B(n6138), .Z(n6092) );
  XOR U6726 ( .A(n6091), .B(n6092), .Z(n5966) );
  NAND U6727 ( .A(n5836), .B(n5835), .Z(n5840) );
  NANDN U6728 ( .A(n5838), .B(n5837), .Z(n5839) );
  NAND U6729 ( .A(n5840), .B(n5839), .Z(n5964) );
  NANDN U6730 ( .A(n5842), .B(n5841), .Z(n5846) );
  OR U6731 ( .A(n5844), .B(n5843), .Z(n5845) );
  AND U6732 ( .A(n5846), .B(n5845), .Z(n5965) );
  XNOR U6733 ( .A(n5964), .B(n5965), .Z(n5967) );
  XOR U6734 ( .A(n5966), .B(n5967), .Z(n6147) );
  XNOR U6735 ( .A(n6148), .B(n6147), .Z(n6150) );
  NANDN U6736 ( .A(n5848), .B(n5847), .Z(n5852) );
  NAND U6737 ( .A(n5850), .B(n5849), .Z(n5851) );
  NAND U6738 ( .A(n5852), .B(n5851), .Z(n6141) );
  NANDN U6739 ( .A(n5854), .B(n5853), .Z(n5858) );
  NAND U6740 ( .A(n5856), .B(n5855), .Z(n5857) );
  NAND U6741 ( .A(n5858), .B(n5857), .Z(n6142) );
  XNOR U6742 ( .A(n6141), .B(n6142), .Z(n6143) );
  XOR U6743 ( .A(b[39]), .B(n11986), .Z(n6041) );
  NANDN U6744 ( .A(n6041), .B(n36553), .Z(n5861) );
  NANDN U6745 ( .A(n5859), .B(n36643), .Z(n5860) );
  NAND U6746 ( .A(n5861), .B(n5860), .Z(n6025) );
  XOR U6747 ( .A(b[5]), .B(n22246), .Z(n6047) );
  OR U6748 ( .A(n6047), .B(n29363), .Z(n5864) );
  NANDN U6749 ( .A(n5862), .B(n29864), .Z(n5863) );
  AND U6750 ( .A(n5864), .B(n5863), .Z(n6023) );
  NAND U6751 ( .A(n34848), .B(n5865), .Z(n5867) );
  XOR U6752 ( .A(n35375), .B(n15484), .Z(n6044) );
  NAND U6753 ( .A(n34618), .B(n6044), .Z(n5866) );
  AND U6754 ( .A(n5867), .B(n5866), .Z(n6024) );
  XOR U6755 ( .A(n6025), .B(n6026), .Z(n5982) );
  AND U6756 ( .A(n5869), .B(n5868), .Z(n6132) );
  NANDN U6757 ( .A(n5870), .B(n37262), .Z(n5872) );
  XNOR U6758 ( .A(b[45]), .B(a[2]), .Z(n6011) );
  NANDN U6759 ( .A(n6011), .B(n37261), .Z(n5871) );
  NAND U6760 ( .A(n5872), .B(n5871), .Z(n6130) );
  XNOR U6761 ( .A(b[25]), .B(n15963), .Z(n6003) );
  NANDN U6762 ( .A(n34219), .B(n6003), .Z(n5875) );
  NANDN U6763 ( .A(n5873), .B(n34217), .Z(n5874) );
  NAND U6764 ( .A(n5875), .B(n5874), .Z(n6129) );
  XOR U6765 ( .A(n6132), .B(n6131), .Z(n5983) );
  XNOR U6766 ( .A(n5982), .B(n5983), .Z(n5984) );
  NANDN U6767 ( .A(n5877), .B(n5876), .Z(n5881) );
  NAND U6768 ( .A(n5879), .B(n5878), .Z(n5880) );
  AND U6769 ( .A(n5881), .B(n5880), .Z(n5985) );
  XNOR U6770 ( .A(n5984), .B(n5985), .Z(n5973) );
  NANDN U6771 ( .A(n5883), .B(n5882), .Z(n5887) );
  NAND U6772 ( .A(n5885), .B(n5884), .Z(n5886) );
  NAND U6773 ( .A(n5887), .B(n5886), .Z(n5970) );
  NANDN U6774 ( .A(n5889), .B(n5888), .Z(n5893) );
  NAND U6775 ( .A(n5891), .B(n5890), .Z(n5892) );
  NAND U6776 ( .A(n5893), .B(n5892), .Z(n5971) );
  XNOR U6777 ( .A(n5970), .B(n5971), .Z(n5972) );
  XNOR U6778 ( .A(n5973), .B(n5972), .Z(n6087) );
  NAND U6779 ( .A(n5895), .B(n5894), .Z(n5899) );
  NANDN U6780 ( .A(n5897), .B(n5896), .Z(n5898) );
  NAND U6781 ( .A(n5899), .B(n5898), .Z(n6085) );
  XOR U6782 ( .A(b[11]), .B(n19980), .Z(n6062) );
  OR U6783 ( .A(n6062), .B(n31369), .Z(n5902) );
  NANDN U6784 ( .A(n5900), .B(n31119), .Z(n5901) );
  NAND U6785 ( .A(n5902), .B(n5901), .Z(n6119) );
  XNOR U6786 ( .A(b[35]), .B(a[12]), .Z(n6114) );
  NANDN U6787 ( .A(n6114), .B(n35985), .Z(n5905) );
  NANDN U6788 ( .A(n5903), .B(n35986), .Z(n5904) );
  AND U6789 ( .A(n5905), .B(n5904), .Z(n6117) );
  XOR U6790 ( .A(b[37]), .B(n12555), .Z(n6038) );
  NANDN U6791 ( .A(n6038), .B(n36311), .Z(n5908) );
  NANDN U6792 ( .A(n5906), .B(n36309), .Z(n5907) );
  AND U6793 ( .A(n5908), .B(n5907), .Z(n6118) );
  XOR U6794 ( .A(n6119), .B(n6120), .Z(n5988) );
  NAND U6795 ( .A(n5909), .B(n34044), .Z(n5911) );
  XOR U6796 ( .A(n34510), .B(n16508), .Z(n6111) );
  NANDN U6797 ( .A(n33867), .B(n6111), .Z(n5910) );
  NAND U6798 ( .A(n5911), .B(n5910), .Z(n6126) );
  XOR U6799 ( .A(n967), .B(n22289), .Z(n6050) );
  NAND U6800 ( .A(n6050), .B(n28939), .Z(n5914) );
  NAND U6801 ( .A(n28938), .B(n5912), .Z(n5913) );
  AND U6802 ( .A(n5914), .B(n5913), .Z(n6123) );
  XNOR U6803 ( .A(b[41]), .B(a[6]), .Z(n6065) );
  OR U6804 ( .A(n6065), .B(n36905), .Z(n5917) );
  NAND U6805 ( .A(n5915), .B(n36807), .Z(n5916) );
  AND U6806 ( .A(n5917), .B(n5916), .Z(n6124) );
  XOR U6807 ( .A(n6126), .B(n6125), .Z(n5989) );
  XNOR U6808 ( .A(n5988), .B(n5989), .Z(n5990) );
  NANDN U6809 ( .A(n5919), .B(n5918), .Z(n5923) );
  NAND U6810 ( .A(n5921), .B(n5920), .Z(n5922) );
  AND U6811 ( .A(n5923), .B(n5922), .Z(n5991) );
  XNOR U6812 ( .A(n5990), .B(n5991), .Z(n6086) );
  XNOR U6813 ( .A(n6085), .B(n6086), .Z(n6088) );
  XOR U6814 ( .A(n6087), .B(n6088), .Z(n6144) );
  XOR U6815 ( .A(n6143), .B(n6144), .Z(n6149) );
  XOR U6816 ( .A(n6150), .B(n6149), .Z(n5958) );
  XNOR U6817 ( .A(n5958), .B(n5959), .Z(n5960) );
  XNOR U6818 ( .A(n5961), .B(n5960), .Z(n5955) );
  NANDN U6819 ( .A(n5929), .B(n5928), .Z(n5933) );
  NAND U6820 ( .A(n5931), .B(n5930), .Z(n5932) );
  NAND U6821 ( .A(n5933), .B(n5932), .Z(n5952) );
  NANDN U6822 ( .A(n5935), .B(n5934), .Z(n5939) );
  NAND U6823 ( .A(n5937), .B(n5936), .Z(n5938) );
  AND U6824 ( .A(n5939), .B(n5938), .Z(n5953) );
  XNOR U6825 ( .A(n5952), .B(n5953), .Z(n5954) );
  XOR U6826 ( .A(n5955), .B(n5954), .Z(n5949) );
  XOR U6827 ( .A(n5948), .B(n5949), .Z(n5940) );
  XNOR U6828 ( .A(n5941), .B(n5940), .Z(n5942) );
  XOR U6829 ( .A(n5943), .B(n5942), .Z(n6154) );
  XOR U6830 ( .A(n6155), .B(n6154), .Z(c[110]) );
  NANDN U6831 ( .A(n5941), .B(n5940), .Z(n5945) );
  NAND U6832 ( .A(n5943), .B(n5942), .Z(n5944) );
  NAND U6833 ( .A(n5945), .B(n5944), .Z(n6166) );
  NANDN U6834 ( .A(n5947), .B(n5946), .Z(n5951) );
  NAND U6835 ( .A(n5949), .B(n5948), .Z(n5950) );
  NAND U6836 ( .A(n5951), .B(n5950), .Z(n6163) );
  NANDN U6837 ( .A(n5953), .B(n5952), .Z(n5957) );
  NAND U6838 ( .A(n5955), .B(n5954), .Z(n5956) );
  NAND U6839 ( .A(n5957), .B(n5956), .Z(n6366) );
  NANDN U6840 ( .A(n5959), .B(n5958), .Z(n5963) );
  NAND U6841 ( .A(n5961), .B(n5960), .Z(n5962) );
  NAND U6842 ( .A(n5963), .B(n5962), .Z(n6364) );
  NANDN U6843 ( .A(n5965), .B(n5964), .Z(n5969) );
  NAND U6844 ( .A(n5967), .B(n5966), .Z(n5968) );
  NAND U6845 ( .A(n5969), .B(n5968), .Z(n6170) );
  NANDN U6846 ( .A(n5971), .B(n5970), .Z(n5975) );
  NANDN U6847 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U6848 ( .A(n5975), .B(n5974), .Z(n6175) );
  NANDN U6849 ( .A(n5977), .B(n5976), .Z(n5981) );
  NAND U6850 ( .A(n5979), .B(n5978), .Z(n5980) );
  NAND U6851 ( .A(n5981), .B(n5980), .Z(n6176) );
  XNOR U6852 ( .A(n6175), .B(n6176), .Z(n6177) );
  NANDN U6853 ( .A(n5983), .B(n5982), .Z(n5987) );
  NAND U6854 ( .A(n5985), .B(n5984), .Z(n5986) );
  NAND U6855 ( .A(n5987), .B(n5986), .Z(n6280) );
  NANDN U6856 ( .A(n5989), .B(n5988), .Z(n5993) );
  NAND U6857 ( .A(n5991), .B(n5990), .Z(n5992) );
  AND U6858 ( .A(n5993), .B(n5992), .Z(n6281) );
  XNOR U6859 ( .A(n6280), .B(n6281), .Z(n6282) );
  NANDN U6860 ( .A(n5995), .B(n5994), .Z(n5999) );
  NAND U6861 ( .A(n5997), .B(n5996), .Z(n5998) );
  NAND U6862 ( .A(n5999), .B(n5998), .Z(n6299) );
  NANDN U6863 ( .A(n966), .B(a[47]), .Z(n6000) );
  XOR U6864 ( .A(n29232), .B(n6000), .Z(n6002) );
  IV U6865 ( .A(a[46]), .Z(n22964) );
  NANDN U6866 ( .A(n22964), .B(n966), .Z(n6001) );
  AND U6867 ( .A(n6002), .B(n6001), .Z(n6255) );
  XNOR U6868 ( .A(b[25]), .B(n16269), .Z(n6193) );
  NANDN U6869 ( .A(n34219), .B(n6193), .Z(n6005) );
  NAND U6870 ( .A(n6003), .B(n34217), .Z(n6004) );
  AND U6871 ( .A(n6005), .B(n6004), .Z(n6256) );
  XNOR U6872 ( .A(n6255), .B(n6256), .Z(n6257) );
  XNOR U6873 ( .A(n978), .B(a[0]), .Z(n6008) );
  XNOR U6874 ( .A(n978), .B(b[45]), .Z(n6007) );
  XNOR U6875 ( .A(b[47]), .B(b[46]), .Z(n6006) );
  ANDN U6876 ( .B(n6007), .A(n6006), .Z(n37469) );
  NAND U6877 ( .A(n6008), .B(n37469), .Z(n6010) );
  XOR U6878 ( .A(b[47]), .B(n10457), .Z(n6190) );
  NANDN U6879 ( .A(n6190), .B(n37471), .Z(n6009) );
  AND U6880 ( .A(n6010), .B(n6009), .Z(n6196) );
  XNOR U6881 ( .A(b[45]), .B(n10524), .Z(n6322) );
  NAND U6882 ( .A(n6322), .B(n37261), .Z(n6013) );
  NANDN U6883 ( .A(n6011), .B(n37262), .Z(n6012) );
  AND U6884 ( .A(n6013), .B(n6012), .Z(n6197) );
  XNOR U6885 ( .A(n6196), .B(n6197), .Z(n6258) );
  XNOR U6886 ( .A(n6257), .B(n6258), .Z(n6298) );
  XNOR U6887 ( .A(n6299), .B(n6298), .Z(n6301) );
  XNOR U6888 ( .A(b[17]), .B(a[31]), .Z(n6259) );
  NANDN U6889 ( .A(n6259), .B(n32543), .Z(n6016) );
  NANDN U6890 ( .A(n6014), .B(n32541), .Z(n6015) );
  NAND U6891 ( .A(n6016), .B(n6015), .Z(n6237) );
  XNOR U6892 ( .A(b[21]), .B(a[27]), .Z(n6271) );
  OR U6893 ( .A(n6271), .B(n33634), .Z(n6019) );
  NAND U6894 ( .A(n6017), .B(n33464), .Z(n6018) );
  NAND U6895 ( .A(n6019), .B(n6018), .Z(n6234) );
  NAND U6896 ( .A(n33283), .B(n6020), .Z(n6022) );
  XOR U6897 ( .A(b[19]), .B(n18003), .Z(n6268) );
  OR U6898 ( .A(n6268), .B(n33021), .Z(n6021) );
  AND U6899 ( .A(n6022), .B(n6021), .Z(n6235) );
  XNOR U6900 ( .A(n6234), .B(n6235), .Z(n6236) );
  XOR U6901 ( .A(n6237), .B(n6236), .Z(n6300) );
  XOR U6902 ( .A(n6301), .B(n6300), .Z(n6356) );
  OR U6903 ( .A(n6024), .B(n6023), .Z(n6028) );
  NANDN U6904 ( .A(n6026), .B(n6025), .Z(n6027) );
  AND U6905 ( .A(n6028), .B(n6027), .Z(n6353) );
  NANDN U6906 ( .A(n6030), .B(n6029), .Z(n6034) );
  NANDN U6907 ( .A(n6032), .B(n6031), .Z(n6033) );
  NAND U6908 ( .A(n6034), .B(n6033), .Z(n6354) );
  XNOR U6909 ( .A(n6356), .B(n6355), .Z(n6277) );
  XOR U6910 ( .A(b[13]), .B(n20315), .Z(n6210) );
  OR U6911 ( .A(n6210), .B(n31550), .Z(n6037) );
  NANDN U6912 ( .A(n6035), .B(n31874), .Z(n6036) );
  NAND U6913 ( .A(n6037), .B(n6036), .Z(n6316) );
  XOR U6914 ( .A(b[37]), .B(n12830), .Z(n6310) );
  NANDN U6915 ( .A(n6310), .B(n36311), .Z(n6040) );
  NANDN U6916 ( .A(n6038), .B(n36309), .Z(n6039) );
  NAND U6917 ( .A(n6040), .B(n6039), .Z(n6313) );
  XOR U6918 ( .A(b[39]), .B(n12258), .Z(n6213) );
  NANDN U6919 ( .A(n6213), .B(n36553), .Z(n6043) );
  NANDN U6920 ( .A(n6041), .B(n36643), .Z(n6042) );
  AND U6921 ( .A(n6043), .B(n6042), .Z(n6314) );
  XNOR U6922 ( .A(n6313), .B(n6314), .Z(n6315) );
  XNOR U6923 ( .A(n6316), .B(n6315), .Z(n6337) );
  NAND U6924 ( .A(n34848), .B(n6044), .Z(n6046) );
  XOR U6925 ( .A(b[27]), .B(n16220), .Z(n6198) );
  NANDN U6926 ( .A(n6198), .B(n34618), .Z(n6045) );
  NAND U6927 ( .A(n6046), .B(n6045), .Z(n6243) );
  XOR U6928 ( .A(b[5]), .B(n21996), .Z(n6187) );
  OR U6929 ( .A(n6187), .B(n29363), .Z(n6049) );
  NANDN U6930 ( .A(n6047), .B(n29864), .Z(n6048) );
  NAND U6931 ( .A(n6049), .B(n6048), .Z(n6240) );
  XOR U6932 ( .A(b[3]), .B(n22579), .Z(n6201) );
  NANDN U6933 ( .A(n6201), .B(n28939), .Z(n6052) );
  NAND U6934 ( .A(n28938), .B(n6050), .Z(n6051) );
  AND U6935 ( .A(n6052), .B(n6051), .Z(n6241) );
  XNOR U6936 ( .A(n6240), .B(n6241), .Z(n6242) );
  XNOR U6937 ( .A(n6243), .B(n6242), .Z(n6335) );
  NANDN U6938 ( .A(n6054), .B(n6053), .Z(n6058) );
  NAND U6939 ( .A(n6056), .B(n6055), .Z(n6057) );
  NAND U6940 ( .A(n6058), .B(n6057), .Z(n6336) );
  XOR U6941 ( .A(n6335), .B(n6336), .Z(n6338) );
  XOR U6942 ( .A(n6337), .B(n6338), .Z(n6275) );
  NAND U6943 ( .A(n35188), .B(n6059), .Z(n6061) );
  XOR U6944 ( .A(n35540), .B(n15113), .Z(n6265) );
  NANDN U6945 ( .A(n34968), .B(n6265), .Z(n6060) );
  NAND U6946 ( .A(n6061), .B(n6060), .Z(n6207) );
  XOR U6947 ( .A(b[11]), .B(n20352), .Z(n6222) );
  OR U6948 ( .A(n6222), .B(n31369), .Z(n6064) );
  NANDN U6949 ( .A(n6062), .B(n31119), .Z(n6063) );
  NAND U6950 ( .A(n6064), .B(n6063), .Z(n6204) );
  XNOR U6951 ( .A(b[41]), .B(a[7]), .Z(n6216) );
  OR U6952 ( .A(n6216), .B(n36905), .Z(n6067) );
  NANDN U6953 ( .A(n6065), .B(n36807), .Z(n6066) );
  AND U6954 ( .A(n6067), .B(n6066), .Z(n6205) );
  XNOR U6955 ( .A(n6204), .B(n6205), .Z(n6206) );
  XNOR U6956 ( .A(n6207), .B(n6206), .Z(n6349) );
  XOR U6957 ( .A(n31123), .B(n21441), .Z(n6252) );
  NAND U6958 ( .A(n6252), .B(n29949), .Z(n6070) );
  NAND U6959 ( .A(n29948), .B(n6068), .Z(n6069) );
  NAND U6960 ( .A(n6070), .B(n6069), .Z(n6328) );
  NOR U6961 ( .A(n978), .B(b[45]), .Z(n6071) );
  NANDN U6962 ( .A(a[0]), .B(n6071), .Z(n6075) );
  ANDN U6963 ( .B(b[45]), .A(n986), .Z(n6073) );
  OR U6964 ( .A(b[46]), .B(n978), .Z(n6072) );
  OR U6965 ( .A(n6073), .B(n6072), .Z(n6074) );
  NAND U6966 ( .A(n6075), .B(n6074), .Z(n6325) );
  XOR U6967 ( .A(b[31]), .B(n14514), .Z(n6246) );
  NANDN U6968 ( .A(n6246), .B(n35313), .Z(n6078) );
  NANDN U6969 ( .A(n6076), .B(n35311), .Z(n6077) );
  AND U6970 ( .A(n6078), .B(n6077), .Z(n6326) );
  XNOR U6971 ( .A(n6325), .B(n6326), .Z(n6327) );
  XNOR U6972 ( .A(n6328), .B(n6327), .Z(n6347) );
  NANDN U6973 ( .A(n6080), .B(n6079), .Z(n6084) );
  NAND U6974 ( .A(n6082), .B(n6081), .Z(n6083) );
  NAND U6975 ( .A(n6084), .B(n6083), .Z(n6348) );
  XOR U6976 ( .A(n6347), .B(n6348), .Z(n6350) );
  XNOR U6977 ( .A(n6349), .B(n6350), .Z(n6274) );
  XOR U6978 ( .A(n6277), .B(n6276), .Z(n6283) );
  XNOR U6979 ( .A(n6282), .B(n6283), .Z(n6178) );
  XOR U6980 ( .A(n6177), .B(n6178), .Z(n6169) );
  XNOR U6981 ( .A(n6170), .B(n6169), .Z(n6172) );
  NANDN U6982 ( .A(n6090), .B(n6089), .Z(n6094) );
  NAND U6983 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U6984 ( .A(n6094), .B(n6093), .Z(n6181) );
  XOR U6985 ( .A(b[33]), .B(n13976), .Z(n6219) );
  NANDN U6986 ( .A(n6219), .B(n35620), .Z(n6101) );
  NANDN U6987 ( .A(n6099), .B(n35621), .Z(n6100) );
  NAND U6988 ( .A(n6101), .B(n6100), .Z(n6332) );
  XOR U6989 ( .A(b[43]), .B(n11202), .Z(n6225) );
  NANDN U6990 ( .A(n6225), .B(n37068), .Z(n6104) );
  NAND U6991 ( .A(n6102), .B(n37069), .Z(n6103) );
  NAND U6992 ( .A(n6104), .B(n6103), .Z(n6329) );
  XOR U6993 ( .A(b[9]), .B(n20867), .Z(n6249) );
  NANDN U6994 ( .A(n6249), .B(n30509), .Z(n6107) );
  NANDN U6995 ( .A(n6105), .B(n30846), .Z(n6106) );
  AND U6996 ( .A(n6107), .B(n6106), .Z(n6330) );
  XNOR U6997 ( .A(n6329), .B(n6330), .Z(n6331) );
  XOR U6998 ( .A(n6332), .B(n6331), .Z(n6344) );
  XOR U6999 ( .A(b[15]), .B(n19656), .Z(n6304) );
  OR U7000 ( .A(n6304), .B(n32010), .Z(n6110) );
  NANDN U7001 ( .A(n6108), .B(n32011), .Z(n6109) );
  NAND U7002 ( .A(n6110), .B(n6109), .Z(n6231) );
  NAND U7003 ( .A(n34044), .B(n6111), .Z(n6113) );
  XOR U7004 ( .A(n34510), .B(n16916), .Z(n6262) );
  NANDN U7005 ( .A(n33867), .B(n6262), .Z(n6112) );
  NAND U7006 ( .A(n6113), .B(n6112), .Z(n6228) );
  XNOR U7007 ( .A(b[35]), .B(a[13]), .Z(n6307) );
  NANDN U7008 ( .A(n6307), .B(n35985), .Z(n6116) );
  NANDN U7009 ( .A(n6114), .B(n35986), .Z(n6115) );
  AND U7010 ( .A(n6116), .B(n6115), .Z(n6229) );
  XNOR U7011 ( .A(n6228), .B(n6229), .Z(n6230) );
  XOR U7012 ( .A(n6231), .B(n6230), .Z(n6342) );
  OR U7013 ( .A(n6118), .B(n6117), .Z(n6122) );
  NANDN U7014 ( .A(n6120), .B(n6119), .Z(n6121) );
  NAND U7015 ( .A(n6122), .B(n6121), .Z(n6341) );
  XNOR U7016 ( .A(n6342), .B(n6341), .Z(n6343) );
  XOR U7017 ( .A(n6344), .B(n6343), .Z(n6295) );
  OR U7018 ( .A(n6124), .B(n6123), .Z(n6128) );
  NAND U7019 ( .A(n6126), .B(n6125), .Z(n6127) );
  NAND U7020 ( .A(n6128), .B(n6127), .Z(n6292) );
  OR U7021 ( .A(n6130), .B(n6129), .Z(n6134) );
  NANDN U7022 ( .A(n6132), .B(n6131), .Z(n6133) );
  NAND U7023 ( .A(n6134), .B(n6133), .Z(n6293) );
  XNOR U7024 ( .A(n6292), .B(n6293), .Z(n6294) );
  XOR U7025 ( .A(n6295), .B(n6294), .Z(n6287) );
  XOR U7026 ( .A(n6286), .B(n6287), .Z(n6288) );
  NAND U7027 ( .A(n6136), .B(n6135), .Z(n6140) );
  NANDN U7028 ( .A(n6138), .B(n6137), .Z(n6139) );
  NAND U7029 ( .A(n6140), .B(n6139), .Z(n6289) );
  XNOR U7030 ( .A(n6288), .B(n6289), .Z(n6182) );
  XNOR U7031 ( .A(n6181), .B(n6182), .Z(n6183) );
  XOR U7032 ( .A(n6184), .B(n6183), .Z(n6171) );
  XNOR U7033 ( .A(n6172), .B(n6171), .Z(n6361) );
  NANDN U7034 ( .A(n6142), .B(n6141), .Z(n6146) );
  NAND U7035 ( .A(n6144), .B(n6143), .Z(n6145) );
  NAND U7036 ( .A(n6146), .B(n6145), .Z(n6359) );
  NAND U7037 ( .A(n6148), .B(n6147), .Z(n6152) );
  NANDN U7038 ( .A(n6150), .B(n6149), .Z(n6151) );
  AND U7039 ( .A(n6152), .B(n6151), .Z(n6360) );
  XNOR U7040 ( .A(n6359), .B(n6360), .Z(n6362) );
  XOR U7041 ( .A(n6361), .B(n6362), .Z(n6363) );
  XNOR U7042 ( .A(n6364), .B(n6363), .Z(n6365) );
  XNOR U7043 ( .A(n6366), .B(n6365), .Z(n6164) );
  XNOR U7044 ( .A(n6163), .B(n6164), .Z(n6165) );
  XNOR U7045 ( .A(n6166), .B(n6165), .Z(n6158) );
  XNOR U7046 ( .A(n6158), .B(sreg[111]), .Z(n6160) );
  NAND U7047 ( .A(n6153), .B(sreg[110]), .Z(n6157) );
  OR U7048 ( .A(n6155), .B(n6154), .Z(n6156) );
  AND U7049 ( .A(n6157), .B(n6156), .Z(n6159) );
  XOR U7050 ( .A(n6160), .B(n6159), .Z(c[111]) );
  NAND U7051 ( .A(n6158), .B(sreg[111]), .Z(n6162) );
  OR U7052 ( .A(n6160), .B(n6159), .Z(n6161) );
  NAND U7053 ( .A(n6162), .B(n6161), .Z(n6584) );
  XNOR U7054 ( .A(n6584), .B(sreg[112]), .Z(n6586) );
  NANDN U7055 ( .A(n6164), .B(n6163), .Z(n6168) );
  NAND U7056 ( .A(n6166), .B(n6165), .Z(n6167) );
  NAND U7057 ( .A(n6168), .B(n6167), .Z(n6372) );
  NAND U7058 ( .A(n6170), .B(n6169), .Z(n6174) );
  NANDN U7059 ( .A(n6172), .B(n6171), .Z(n6173) );
  NAND U7060 ( .A(n6174), .B(n6173), .Z(n6378) );
  NANDN U7061 ( .A(n6176), .B(n6175), .Z(n6180) );
  NAND U7062 ( .A(n6178), .B(n6177), .Z(n6179) );
  NAND U7063 ( .A(n6180), .B(n6179), .Z(n6375) );
  NANDN U7064 ( .A(n6182), .B(n6181), .Z(n6186) );
  NAND U7065 ( .A(n6184), .B(n6183), .Z(n6185) );
  AND U7066 ( .A(n6186), .B(n6185), .Z(n6376) );
  XNOR U7067 ( .A(n6375), .B(n6376), .Z(n6377) );
  XNOR U7068 ( .A(n6378), .B(n6377), .Z(n6578) );
  XOR U7069 ( .A(b[5]), .B(n22289), .Z(n6419) );
  OR U7070 ( .A(n6419), .B(n29363), .Z(n6189) );
  NANDN U7071 ( .A(n6187), .B(n29864), .Z(n6188) );
  NAND U7072 ( .A(n6189), .B(n6188), .Z(n6498) );
  NANDN U7073 ( .A(n6190), .B(n37469), .Z(n6192) );
  XOR U7074 ( .A(n978), .B(n10363), .Z(n6466) );
  NAND U7075 ( .A(n6466), .B(n37471), .Z(n6191) );
  NAND U7076 ( .A(n6192), .B(n6191), .Z(n6495) );
  XNOR U7077 ( .A(b[25]), .B(a[24]), .Z(n6474) );
  OR U7078 ( .A(n6474), .B(n34219), .Z(n6195) );
  NAND U7079 ( .A(n34217), .B(n6193), .Z(n6194) );
  AND U7080 ( .A(n6195), .B(n6194), .Z(n6496) );
  XNOR U7081 ( .A(n6495), .B(n6496), .Z(n6497) );
  XNOR U7082 ( .A(n6498), .B(n6497), .Z(n6442) );
  NANDN U7083 ( .A(n6198), .B(n34848), .Z(n6200) );
  XOR U7084 ( .A(b[27]), .B(n15963), .Z(n6439) );
  NANDN U7085 ( .A(n6439), .B(n34618), .Z(n6199) );
  NAND U7086 ( .A(n6200), .B(n6199), .Z(n6449) );
  XNOR U7087 ( .A(n967), .B(a[46]), .Z(n6422) );
  NAND U7088 ( .A(n6422), .B(n28939), .Z(n6203) );
  NANDN U7089 ( .A(n6201), .B(n28938), .Z(n6202) );
  AND U7090 ( .A(n6203), .B(n6202), .Z(n6448) );
  XNOR U7091 ( .A(n6449), .B(n6448), .Z(n6450) );
  XNOR U7092 ( .A(n6451), .B(n6450), .Z(n6443) );
  XNOR U7093 ( .A(n6442), .B(n6443), .Z(n6444) );
  NANDN U7094 ( .A(n6205), .B(n6204), .Z(n6209) );
  NAND U7095 ( .A(n6207), .B(n6206), .Z(n6208) );
  AND U7096 ( .A(n6209), .B(n6208), .Z(n6445) );
  XNOR U7097 ( .A(n6444), .B(n6445), .Z(n6532) );
  XOR U7098 ( .A(n971), .B(n19980), .Z(n6507) );
  NANDN U7099 ( .A(n31550), .B(n6507), .Z(n6212) );
  NANDN U7100 ( .A(n6210), .B(n31874), .Z(n6211) );
  NAND U7101 ( .A(n6212), .B(n6211), .Z(n6431) );
  XOR U7102 ( .A(n976), .B(n12555), .Z(n6510) );
  NAND U7103 ( .A(n6510), .B(n36553), .Z(n6215) );
  NANDN U7104 ( .A(n6213), .B(n36643), .Z(n6214) );
  NAND U7105 ( .A(n6215), .B(n6214), .Z(n6428) );
  XNOR U7106 ( .A(b[41]), .B(n11986), .Z(n6513) );
  NANDN U7107 ( .A(n36905), .B(n6513), .Z(n6218) );
  NANDN U7108 ( .A(n6216), .B(n36807), .Z(n6217) );
  AND U7109 ( .A(n6218), .B(n6217), .Z(n6429) );
  XNOR U7110 ( .A(n6428), .B(n6429), .Z(n6430) );
  XNOR U7111 ( .A(n6431), .B(n6430), .Z(n6411) );
  XOR U7112 ( .A(b[33]), .B(n14259), .Z(n6480) );
  NANDN U7113 ( .A(n6480), .B(n35620), .Z(n6221) );
  NANDN U7114 ( .A(n6219), .B(n35621), .Z(n6220) );
  NAND U7115 ( .A(n6221), .B(n6220), .Z(n6548) );
  XOR U7116 ( .A(b[11]), .B(n20686), .Z(n6483) );
  OR U7117 ( .A(n6483), .B(n31369), .Z(n6224) );
  NANDN U7118 ( .A(n6222), .B(n31119), .Z(n6223) );
  NAND U7119 ( .A(n6224), .B(n6223), .Z(n6545) );
  XOR U7120 ( .A(n977), .B(n11406), .Z(n6519) );
  NAND U7121 ( .A(n6519), .B(n37068), .Z(n6227) );
  NANDN U7122 ( .A(n6225), .B(n37069), .Z(n6226) );
  AND U7123 ( .A(n6227), .B(n6226), .Z(n6546) );
  XNOR U7124 ( .A(n6545), .B(n6546), .Z(n6547) );
  XOR U7125 ( .A(n6548), .B(n6547), .Z(n6412) );
  XNOR U7126 ( .A(n6411), .B(n6412), .Z(n6413) );
  NANDN U7127 ( .A(n6229), .B(n6228), .Z(n6233) );
  NAND U7128 ( .A(n6231), .B(n6230), .Z(n6232) );
  AND U7129 ( .A(n6233), .B(n6232), .Z(n6414) );
  XNOR U7130 ( .A(n6413), .B(n6414), .Z(n6527) );
  NANDN U7131 ( .A(n6235), .B(n6234), .Z(n6239) );
  NAND U7132 ( .A(n6237), .B(n6236), .Z(n6238) );
  NAND U7133 ( .A(n6239), .B(n6238), .Z(n6525) );
  NANDN U7134 ( .A(n6241), .B(n6240), .Z(n6245) );
  NAND U7135 ( .A(n6243), .B(n6242), .Z(n6244) );
  NAND U7136 ( .A(n6245), .B(n6244), .Z(n6526) );
  XNOR U7137 ( .A(n6525), .B(n6526), .Z(n6528) );
  XNOR U7138 ( .A(n6527), .B(n6528), .Z(n6530) );
  XOR U7139 ( .A(b[31]), .B(n14905), .Z(n6516) );
  NANDN U7140 ( .A(n6516), .B(n35313), .Z(n6248) );
  NANDN U7141 ( .A(n6246), .B(n35311), .Z(n6247) );
  NAND U7142 ( .A(n6248), .B(n6247), .Z(n6575) );
  XOR U7143 ( .A(b[9]), .B(n21149), .Z(n6486) );
  NANDN U7144 ( .A(n6486), .B(n30509), .Z(n6251) );
  NANDN U7145 ( .A(n6249), .B(n30846), .Z(n6250) );
  NAND U7146 ( .A(n6251), .B(n6250), .Z(n6572) );
  XOR U7147 ( .A(b[7]), .B(n22246), .Z(n6522) );
  NANDN U7148 ( .A(n6522), .B(n29949), .Z(n6254) );
  NAND U7149 ( .A(n29948), .B(n6252), .Z(n6253) );
  AND U7150 ( .A(n6254), .B(n6253), .Z(n6573) );
  XNOR U7151 ( .A(n6572), .B(n6573), .Z(n6574) );
  XNOR U7152 ( .A(n6575), .B(n6574), .Z(n6544) );
  XNOR U7153 ( .A(b[17]), .B(a[32]), .Z(n6569) );
  NANDN U7154 ( .A(n6569), .B(n32543), .Z(n6261) );
  NANDN U7155 ( .A(n6259), .B(n32541), .Z(n6260) );
  NAND U7156 ( .A(n6261), .B(n6260), .Z(n6462) );
  NAND U7157 ( .A(n34044), .B(n6262), .Z(n6264) );
  XOR U7158 ( .A(n34510), .B(n17133), .Z(n6425) );
  NANDN U7159 ( .A(n33867), .B(n6425), .Z(n6263) );
  AND U7160 ( .A(n6264), .B(n6263), .Z(n6460) );
  NAND U7161 ( .A(n35188), .B(n6265), .Z(n6267) );
  XOR U7162 ( .A(n35540), .B(n15484), .Z(n6566) );
  NANDN U7163 ( .A(n34968), .B(n6566), .Z(n6266) );
  AND U7164 ( .A(n6267), .B(n6266), .Z(n6461) );
  XOR U7165 ( .A(n6462), .B(n6463), .Z(n6457) );
  NANDN U7166 ( .A(n6268), .B(n33283), .Z(n6270) );
  XNOR U7167 ( .A(n33020), .B(a[30]), .Z(n6563) );
  NANDN U7168 ( .A(n33021), .B(n6563), .Z(n6269) );
  NAND U7169 ( .A(n6270), .B(n6269), .Z(n6455) );
  XNOR U7170 ( .A(b[21]), .B(n17702), .Z(n6560) );
  NANDN U7171 ( .A(n33634), .B(n6560), .Z(n6273) );
  NANDN U7172 ( .A(n6271), .B(n33464), .Z(n6272) );
  AND U7173 ( .A(n6273), .B(n6272), .Z(n6454) );
  XNOR U7174 ( .A(n6455), .B(n6454), .Z(n6456) );
  XOR U7175 ( .A(n6457), .B(n6456), .Z(n6541) );
  XNOR U7176 ( .A(n6542), .B(n6541), .Z(n6543) );
  XOR U7177 ( .A(n6544), .B(n6543), .Z(n6529) );
  XNOR U7178 ( .A(n6530), .B(n6529), .Z(n6531) );
  XOR U7179 ( .A(n6532), .B(n6531), .Z(n6408) );
  NANDN U7180 ( .A(n6275), .B(n6274), .Z(n6279) );
  NANDN U7181 ( .A(n6277), .B(n6276), .Z(n6278) );
  NAND U7182 ( .A(n6279), .B(n6278), .Z(n6406) );
  NANDN U7183 ( .A(n6281), .B(n6280), .Z(n6285) );
  NANDN U7184 ( .A(n6283), .B(n6282), .Z(n6284) );
  AND U7185 ( .A(n6285), .B(n6284), .Z(n6405) );
  XNOR U7186 ( .A(n6406), .B(n6405), .Z(n6407) );
  XNOR U7187 ( .A(n6408), .B(n6407), .Z(n6381) );
  OR U7188 ( .A(n6287), .B(n6286), .Z(n6291) );
  NANDN U7189 ( .A(n6289), .B(n6288), .Z(n6290) );
  NAND U7190 ( .A(n6291), .B(n6290), .Z(n6382) );
  XNOR U7191 ( .A(n6381), .B(n6382), .Z(n6383) );
  NANDN U7192 ( .A(n6293), .B(n6292), .Z(n6297) );
  NANDN U7193 ( .A(n6295), .B(n6294), .Z(n6296) );
  NAND U7194 ( .A(n6297), .B(n6296), .Z(n6389) );
  NAND U7195 ( .A(n6299), .B(n6298), .Z(n6303) );
  NANDN U7196 ( .A(n6301), .B(n6300), .Z(n6302) );
  NAND U7197 ( .A(n6303), .B(n6302), .Z(n6388) );
  XOR U7198 ( .A(b[15]), .B(n19513), .Z(n6551) );
  OR U7199 ( .A(n6551), .B(n32010), .Z(n6306) );
  NANDN U7200 ( .A(n6304), .B(n32011), .Z(n6305) );
  NAND U7201 ( .A(n6306), .B(n6305), .Z(n6504) );
  XNOR U7202 ( .A(b[35]), .B(a[14]), .Z(n6554) );
  NANDN U7203 ( .A(n6554), .B(n35985), .Z(n6309) );
  NANDN U7204 ( .A(n6307), .B(n35986), .Z(n6308) );
  NAND U7205 ( .A(n6309), .B(n6308), .Z(n6501) );
  XOR U7206 ( .A(b[37]), .B(n13106), .Z(n6557) );
  NANDN U7207 ( .A(n6557), .B(n36311), .Z(n6312) );
  NANDN U7208 ( .A(n6310), .B(n36309), .Z(n6311) );
  AND U7209 ( .A(n6312), .B(n6311), .Z(n6502) );
  XNOR U7210 ( .A(n6501), .B(n6502), .Z(n6503) );
  XNOR U7211 ( .A(n6504), .B(n6503), .Z(n6415) );
  NANDN U7212 ( .A(n6314), .B(n6313), .Z(n6318) );
  NAND U7213 ( .A(n6316), .B(n6315), .Z(n6317) );
  NAND U7214 ( .A(n6318), .B(n6317), .Z(n6416) );
  XNOR U7215 ( .A(n6415), .B(n6416), .Z(n6417) );
  XOR U7216 ( .A(n978), .B(b[48]), .Z(n37756) );
  NOR U7217 ( .A(n986), .B(n37756), .Z(n6492) );
  NANDN U7218 ( .A(n966), .B(a[48]), .Z(n6319) );
  XOR U7219 ( .A(n29232), .B(n6319), .Z(n6321) );
  IV U7220 ( .A(a[47]), .Z(n23149) );
  NANDN U7221 ( .A(n23149), .B(n966), .Z(n6320) );
  AND U7222 ( .A(n6321), .B(n6320), .Z(n6490) );
  NAND U7223 ( .A(n37262), .B(n6322), .Z(n6324) );
  XOR U7224 ( .A(b[45]), .B(n10854), .Z(n6436) );
  NANDN U7225 ( .A(n6436), .B(n37261), .Z(n6323) );
  AND U7226 ( .A(n6324), .B(n6323), .Z(n6489) );
  XNOR U7227 ( .A(n6490), .B(n6489), .Z(n6491) );
  XOR U7228 ( .A(n6492), .B(n6491), .Z(n6418) );
  XNOR U7229 ( .A(n6417), .B(n6418), .Z(n6537) );
  NANDN U7230 ( .A(n6330), .B(n6329), .Z(n6334) );
  NAND U7231 ( .A(n6332), .B(n6331), .Z(n6333) );
  AND U7232 ( .A(n6334), .B(n6333), .Z(n6535) );
  XNOR U7233 ( .A(n6536), .B(n6535), .Z(n6538) );
  XOR U7234 ( .A(n6537), .B(n6538), .Z(n6387) );
  XOR U7235 ( .A(n6388), .B(n6387), .Z(n6390) );
  XOR U7236 ( .A(n6389), .B(n6390), .Z(n6401) );
  NANDN U7237 ( .A(n6336), .B(n6335), .Z(n6340) );
  NANDN U7238 ( .A(n6338), .B(n6337), .Z(n6339) );
  NAND U7239 ( .A(n6340), .B(n6339), .Z(n6399) );
  OR U7240 ( .A(n6342), .B(n6341), .Z(n6346) );
  OR U7241 ( .A(n6344), .B(n6343), .Z(n6345) );
  NAND U7242 ( .A(n6346), .B(n6345), .Z(n6396) );
  NANDN U7243 ( .A(n6348), .B(n6347), .Z(n6352) );
  NANDN U7244 ( .A(n6350), .B(n6349), .Z(n6351) );
  NAND U7245 ( .A(n6352), .B(n6351), .Z(n6393) );
  OR U7246 ( .A(n6354), .B(n6353), .Z(n6358) );
  NANDN U7247 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U7248 ( .A(n6358), .B(n6357), .Z(n6394) );
  XNOR U7249 ( .A(n6393), .B(n6394), .Z(n6395) );
  XNOR U7250 ( .A(n6396), .B(n6395), .Z(n6400) );
  XNOR U7251 ( .A(n6399), .B(n6400), .Z(n6402) );
  XOR U7252 ( .A(n6401), .B(n6402), .Z(n6384) );
  XOR U7253 ( .A(n6383), .B(n6384), .Z(n6579) );
  XOR U7254 ( .A(n6578), .B(n6579), .Z(n6581) );
  XNOR U7255 ( .A(n6581), .B(n6580), .Z(n6369) );
  NANDN U7256 ( .A(n6364), .B(n6363), .Z(n6368) );
  NAND U7257 ( .A(n6366), .B(n6365), .Z(n6367) );
  AND U7258 ( .A(n6368), .B(n6367), .Z(n6370) );
  XNOR U7259 ( .A(n6369), .B(n6370), .Z(n6371) );
  XOR U7260 ( .A(n6372), .B(n6371), .Z(n6585) );
  XOR U7261 ( .A(n6586), .B(n6585), .Z(c[112]) );
  NANDN U7262 ( .A(n6370), .B(n6369), .Z(n6374) );
  NAND U7263 ( .A(n6372), .B(n6371), .Z(n6373) );
  NAND U7264 ( .A(n6374), .B(n6373), .Z(n6597) );
  NANDN U7265 ( .A(n6376), .B(n6375), .Z(n6380) );
  NAND U7266 ( .A(n6378), .B(n6377), .Z(n6379) );
  NAND U7267 ( .A(n6380), .B(n6379), .Z(n6602) );
  NANDN U7268 ( .A(n6382), .B(n6381), .Z(n6386) );
  NAND U7269 ( .A(n6384), .B(n6383), .Z(n6385) );
  NAND U7270 ( .A(n6386), .B(n6385), .Z(n6601) );
  NANDN U7271 ( .A(n6388), .B(n6387), .Z(n6392) );
  OR U7272 ( .A(n6390), .B(n6389), .Z(n6391) );
  AND U7273 ( .A(n6392), .B(n6391), .Z(n6606) );
  NANDN U7274 ( .A(n6394), .B(n6393), .Z(n6398) );
  NAND U7275 ( .A(n6396), .B(n6395), .Z(n6397) );
  AND U7276 ( .A(n6398), .B(n6397), .Z(n6607) );
  XNOR U7277 ( .A(n6606), .B(n6607), .Z(n6608) );
  NANDN U7278 ( .A(n6400), .B(n6399), .Z(n6404) );
  NAND U7279 ( .A(n6402), .B(n6401), .Z(n6403) );
  AND U7280 ( .A(n6404), .B(n6403), .Z(n6609) );
  XOR U7281 ( .A(n6608), .B(n6609), .Z(n6612) );
  NANDN U7282 ( .A(n6406), .B(n6405), .Z(n6410) );
  NAND U7283 ( .A(n6408), .B(n6407), .Z(n6409) );
  AND U7284 ( .A(n6410), .B(n6409), .Z(n6613) );
  XNOR U7285 ( .A(n6612), .B(n6613), .Z(n6615) );
  XOR U7286 ( .A(b[5]), .B(n22579), .Z(n6652) );
  OR U7287 ( .A(n6652), .B(n29363), .Z(n6421) );
  NANDN U7288 ( .A(n6419), .B(n29864), .Z(n6420) );
  NAND U7289 ( .A(n6421), .B(n6420), .Z(n6735) );
  XOR U7290 ( .A(b[3]), .B(n23149), .Z(n6776) );
  NANDN U7291 ( .A(n6776), .B(n28939), .Z(n6424) );
  NAND U7292 ( .A(n6422), .B(n28938), .Z(n6423) );
  NAND U7293 ( .A(n6424), .B(n6423), .Z(n6732) );
  NAND U7294 ( .A(n34044), .B(n6425), .Z(n6427) );
  XOR U7295 ( .A(n34510), .B(n17960), .Z(n6765) );
  NANDN U7296 ( .A(n33867), .B(n6765), .Z(n6426) );
  AND U7297 ( .A(n6427), .B(n6426), .Z(n6733) );
  XNOR U7298 ( .A(n6732), .B(n6733), .Z(n6734) );
  XNOR U7299 ( .A(n6735), .B(n6734), .Z(n6704) );
  NANDN U7300 ( .A(n6429), .B(n6428), .Z(n6433) );
  NAND U7301 ( .A(n6431), .B(n6430), .Z(n6432) );
  NAND U7302 ( .A(n6433), .B(n6432), .Z(n6702) );
  NOR U7303 ( .A(b[47]), .B(b[48]), .Z(n6434) );
  OR U7304 ( .A(n6434), .B(n986), .Z(n6435) );
  NANDN U7305 ( .A(n978), .B(b[48]), .Z(n37754) );
  AND U7306 ( .A(n37754), .B(b[49]), .Z(n37862) );
  AND U7307 ( .A(n6435), .B(n37862), .Z(n6727) );
  NANDN U7308 ( .A(n6436), .B(n37262), .Z(n6438) );
  XNOR U7309 ( .A(b[45]), .B(a[5]), .Z(n6747) );
  NANDN U7310 ( .A(n6747), .B(n37261), .Z(n6437) );
  NAND U7311 ( .A(n6438), .B(n6437), .Z(n6726) );
  XOR U7312 ( .A(n6727), .B(n6726), .Z(n6728) );
  NANDN U7313 ( .A(n6439), .B(n34848), .Z(n6441) );
  XOR U7314 ( .A(b[27]), .B(n16269), .Z(n6773) );
  NANDN U7315 ( .A(n6773), .B(n34618), .Z(n6440) );
  AND U7316 ( .A(n6441), .B(n6440), .Z(n6729) );
  XOR U7317 ( .A(n6728), .B(n6729), .Z(n6701) );
  XNOR U7318 ( .A(n6702), .B(n6701), .Z(n6703) );
  XOR U7319 ( .A(n6704), .B(n6703), .Z(n6667) );
  XNOR U7320 ( .A(n6668), .B(n6667), .Z(n6670) );
  XNOR U7321 ( .A(n6669), .B(n6670), .Z(n6800) );
  NANDN U7322 ( .A(n6443), .B(n6442), .Z(n6447) );
  NAND U7323 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U7324 ( .A(n6447), .B(n6446), .Z(n6673) );
  NANDN U7325 ( .A(n6449), .B(n6448), .Z(n6453) );
  NAND U7326 ( .A(n6451), .B(n6450), .Z(n6452) );
  NAND U7327 ( .A(n6453), .B(n6452), .Z(n6692) );
  NANDN U7328 ( .A(n6455), .B(n6454), .Z(n6459) );
  NAND U7329 ( .A(n6457), .B(n6456), .Z(n6458) );
  NAND U7330 ( .A(n6459), .B(n6458), .Z(n6689) );
  OR U7331 ( .A(n6461), .B(n6460), .Z(n6465) );
  NANDN U7332 ( .A(n6463), .B(n6462), .Z(n6464) );
  NAND U7333 ( .A(n6465), .B(n6464), .Z(n6690) );
  XNOR U7334 ( .A(n6689), .B(n6690), .Z(n6691) );
  XNOR U7335 ( .A(n6692), .B(n6691), .Z(n6674) );
  XNOR U7336 ( .A(n6673), .B(n6674), .Z(n6675) );
  NAND U7337 ( .A(n37469), .B(n6466), .Z(n6468) );
  XOR U7338 ( .A(n978), .B(n10524), .Z(n6717) );
  NAND U7339 ( .A(n37471), .B(n6717), .Z(n6467) );
  NAND U7340 ( .A(n6468), .B(n6467), .Z(n6771) );
  XNOR U7341 ( .A(n979), .B(a[0]), .Z(n6471) );
  XNOR U7342 ( .A(n979), .B(b[47]), .Z(n6470) );
  XNOR U7343 ( .A(n979), .B(b[48]), .Z(n6469) );
  AND U7344 ( .A(n6470), .B(n6469), .Z(n37652) );
  NAND U7345 ( .A(n6471), .B(n37652), .Z(n6473) );
  XOR U7346 ( .A(n979), .B(n10457), .Z(n6640) );
  ANDN U7347 ( .B(n6640), .A(n37756), .Z(n6472) );
  ANDN U7348 ( .B(n6473), .A(n6472), .Z(n6772) );
  XNOR U7349 ( .A(n6771), .B(n6772), .Z(n6658) );
  XNOR U7350 ( .A(b[25]), .B(n16916), .Z(n6768) );
  NANDN U7351 ( .A(n34219), .B(n6768), .Z(n6476) );
  NANDN U7352 ( .A(n6474), .B(n34217), .Z(n6475) );
  NAND U7353 ( .A(n6476), .B(n6475), .Z(n6656) );
  NANDN U7354 ( .A(n966), .B(a[49]), .Z(n6477) );
  XOR U7355 ( .A(n29232), .B(n6477), .Z(n6479) );
  IV U7356 ( .A(a[48]), .Z(n23447) );
  NANDN U7357 ( .A(n23447), .B(n966), .Z(n6478) );
  AND U7358 ( .A(n6479), .B(n6478), .Z(n6655) );
  XNOR U7359 ( .A(n6656), .B(n6655), .Z(n6657) );
  XOR U7360 ( .A(n6658), .B(n6657), .Z(n6791) );
  XNOR U7361 ( .A(n974), .B(a[17]), .Z(n6637) );
  NAND U7362 ( .A(n35620), .B(n6637), .Z(n6482) );
  NANDN U7363 ( .A(n6480), .B(n35621), .Z(n6481) );
  AND U7364 ( .A(n6482), .B(n6481), .Z(n6741) );
  XNOR U7365 ( .A(n970), .B(a[39]), .Z(n6750) );
  NANDN U7366 ( .A(n31369), .B(n6750), .Z(n6485) );
  NANDN U7367 ( .A(n6483), .B(n31119), .Z(n6484) );
  AND U7368 ( .A(n6485), .B(n6484), .Z(n6738) );
  XOR U7369 ( .A(b[9]), .B(n21441), .Z(n6643) );
  NANDN U7370 ( .A(n6643), .B(n30509), .Z(n6488) );
  NANDN U7371 ( .A(n6486), .B(n30846), .Z(n6487) );
  AND U7372 ( .A(n6488), .B(n6487), .Z(n6739) );
  XNOR U7373 ( .A(n6738), .B(n6739), .Z(n6740) );
  XOR U7374 ( .A(n6791), .B(n6792), .Z(n6793) );
  NANDN U7375 ( .A(n6490), .B(n6489), .Z(n6494) );
  NANDN U7376 ( .A(n6492), .B(n6491), .Z(n6493) );
  NAND U7377 ( .A(n6494), .B(n6493), .Z(n6794) );
  XOR U7378 ( .A(n6793), .B(n6794), .Z(n6686) );
  NANDN U7379 ( .A(n6496), .B(n6495), .Z(n6500) );
  NAND U7380 ( .A(n6498), .B(n6497), .Z(n6499) );
  NAND U7381 ( .A(n6500), .B(n6499), .Z(n6683) );
  NANDN U7382 ( .A(n6502), .B(n6501), .Z(n6506) );
  NAND U7383 ( .A(n6504), .B(n6503), .Z(n6505) );
  NAND U7384 ( .A(n6506), .B(n6505), .Z(n6788) );
  NAND U7385 ( .A(n31874), .B(n6507), .Z(n6509) );
  XNOR U7386 ( .A(n971), .B(a[37]), .Z(n6628) );
  NANDN U7387 ( .A(n31550), .B(n6628), .Z(n6508) );
  NAND U7388 ( .A(n6509), .B(n6508), .Z(n6626) );
  NAND U7389 ( .A(n36643), .B(n6510), .Z(n6512) );
  XNOR U7390 ( .A(n976), .B(a[11]), .Z(n6756) );
  NAND U7391 ( .A(n6756), .B(n36553), .Z(n6511) );
  NAND U7392 ( .A(n6512), .B(n6511), .Z(n6624) );
  NAND U7393 ( .A(n36807), .B(n6513), .Z(n6515) );
  XNOR U7394 ( .A(b[41]), .B(n12258), .Z(n6759) );
  NANDN U7395 ( .A(n36905), .B(n6759), .Z(n6514) );
  NAND U7396 ( .A(n6515), .B(n6514), .Z(n6625) );
  XNOR U7397 ( .A(n6624), .B(n6625), .Z(n6627) );
  XOR U7398 ( .A(n6626), .B(n6627), .Z(n6785) );
  NANDN U7399 ( .A(n6516), .B(n35311), .Z(n6518) );
  XNOR U7400 ( .A(n973), .B(a[19]), .Z(n6631) );
  NAND U7401 ( .A(n6631), .B(n35313), .Z(n6517) );
  NAND U7402 ( .A(n6518), .B(n6517), .Z(n6663) );
  NAND U7403 ( .A(n37069), .B(n6519), .Z(n6521) );
  XNOR U7404 ( .A(n977), .B(a[7]), .Z(n6753) );
  NAND U7405 ( .A(n6753), .B(n37068), .Z(n6520) );
  AND U7406 ( .A(n6521), .B(n6520), .Z(n6662) );
  XNOR U7407 ( .A(n31123), .B(a[43]), .Z(n6649) );
  NAND U7408 ( .A(n6649), .B(n29949), .Z(n6524) );
  NANDN U7409 ( .A(n6522), .B(n29948), .Z(n6523) );
  NAND U7410 ( .A(n6524), .B(n6523), .Z(n6661) );
  XNOR U7411 ( .A(n6662), .B(n6661), .Z(n6664) );
  XOR U7412 ( .A(n6663), .B(n6664), .Z(n6786) );
  XNOR U7413 ( .A(n6785), .B(n6786), .Z(n6787) );
  XOR U7414 ( .A(n6788), .B(n6787), .Z(n6684) );
  XOR U7415 ( .A(n6683), .B(n6684), .Z(n6685) );
  XOR U7416 ( .A(n6686), .B(n6685), .Z(n6676) );
  XOR U7417 ( .A(n6675), .B(n6676), .Z(n6798) );
  XOR U7418 ( .A(n6798), .B(n6797), .Z(n6799) );
  XOR U7419 ( .A(n6800), .B(n6799), .Z(n6805) );
  NANDN U7420 ( .A(n6530), .B(n6529), .Z(n6534) );
  NANDN U7421 ( .A(n6532), .B(n6531), .Z(n6533) );
  NAND U7422 ( .A(n6534), .B(n6533), .Z(n6804) );
  NANDN U7423 ( .A(n6536), .B(n6535), .Z(n6540) );
  NAND U7424 ( .A(n6538), .B(n6537), .Z(n6539) );
  AND U7425 ( .A(n6540), .B(n6539), .Z(n6682) );
  NANDN U7426 ( .A(n6546), .B(n6545), .Z(n6550) );
  NAND U7427 ( .A(n6548), .B(n6547), .Z(n6549) );
  NAND U7428 ( .A(n6550), .B(n6549), .Z(n6698) );
  XOR U7429 ( .A(b[15]), .B(n20315), .Z(n6762) );
  OR U7430 ( .A(n6762), .B(n32010), .Z(n6553) );
  NANDN U7431 ( .A(n6551), .B(n32011), .Z(n6552) );
  NAND U7432 ( .A(n6553), .B(n6552), .Z(n6723) );
  XNOR U7433 ( .A(b[35]), .B(a[15]), .Z(n6744) );
  NANDN U7434 ( .A(n6744), .B(n35985), .Z(n6556) );
  NANDN U7435 ( .A(n6554), .B(n35986), .Z(n6555) );
  NAND U7436 ( .A(n6556), .B(n6555), .Z(n6720) );
  XOR U7437 ( .A(b[37]), .B(n13509), .Z(n6634) );
  NANDN U7438 ( .A(n6634), .B(n36311), .Z(n6559) );
  NANDN U7439 ( .A(n6557), .B(n36309), .Z(n6558) );
  AND U7440 ( .A(n6559), .B(n6558), .Z(n6721) );
  XNOR U7441 ( .A(n6720), .B(n6721), .Z(n6722) );
  XNOR U7442 ( .A(n6723), .B(n6722), .Z(n6621) );
  XNOR U7443 ( .A(b[21]), .B(a[29]), .Z(n6705) );
  OR U7444 ( .A(n6705), .B(n33634), .Z(n6562) );
  NAND U7445 ( .A(n6560), .B(n33464), .Z(n6561) );
  NAND U7446 ( .A(n6562), .B(n6561), .Z(n6782) );
  NAND U7447 ( .A(n6563), .B(n33283), .Z(n6565) );
  XOR U7448 ( .A(n33020), .B(n18639), .Z(n6711) );
  NANDN U7449 ( .A(n33021), .B(n6711), .Z(n6564) );
  NAND U7450 ( .A(n6565), .B(n6564), .Z(n6779) );
  NAND U7451 ( .A(n35188), .B(n6566), .Z(n6568) );
  XOR U7452 ( .A(n35540), .B(n16220), .Z(n6646) );
  NANDN U7453 ( .A(n34968), .B(n6646), .Z(n6567) );
  AND U7454 ( .A(n6568), .B(n6567), .Z(n6780) );
  XNOR U7455 ( .A(n6779), .B(n6780), .Z(n6781) );
  XNOR U7456 ( .A(n6782), .B(n6781), .Z(n6618) );
  XNOR U7457 ( .A(b[17]), .B(n19656), .Z(n6708) );
  NAND U7458 ( .A(n6708), .B(n32543), .Z(n6571) );
  NANDN U7459 ( .A(n6569), .B(n32541), .Z(n6570) );
  NAND U7460 ( .A(n6571), .B(n6570), .Z(n6619) );
  XNOR U7461 ( .A(n6618), .B(n6619), .Z(n6620) );
  XOR U7462 ( .A(n6621), .B(n6620), .Z(n6696) );
  NANDN U7463 ( .A(n6573), .B(n6572), .Z(n6577) );
  NAND U7464 ( .A(n6575), .B(n6574), .Z(n6576) );
  AND U7465 ( .A(n6577), .B(n6576), .Z(n6695) );
  XOR U7466 ( .A(n6696), .B(n6695), .Z(n6697) );
  XOR U7467 ( .A(n6698), .B(n6697), .Z(n6680) );
  XNOR U7468 ( .A(n6679), .B(n6680), .Z(n6681) );
  XNOR U7469 ( .A(n6682), .B(n6681), .Z(n6803) );
  XNOR U7470 ( .A(n6804), .B(n6803), .Z(n6806) );
  XOR U7471 ( .A(n6805), .B(n6806), .Z(n6614) );
  XNOR U7472 ( .A(n6615), .B(n6614), .Z(n6600) );
  XNOR U7473 ( .A(n6601), .B(n6600), .Z(n6603) );
  XNOR U7474 ( .A(n6602), .B(n6603), .Z(n6594) );
  NANDN U7475 ( .A(n6579), .B(n6578), .Z(n6583) );
  OR U7476 ( .A(n6581), .B(n6580), .Z(n6582) );
  AND U7477 ( .A(n6583), .B(n6582), .Z(n6595) );
  XOR U7478 ( .A(n6594), .B(n6595), .Z(n6596) );
  XNOR U7479 ( .A(n6597), .B(n6596), .Z(n6589) );
  XNOR U7480 ( .A(n6589), .B(sreg[113]), .Z(n6591) );
  NAND U7481 ( .A(n6584), .B(sreg[112]), .Z(n6588) );
  OR U7482 ( .A(n6586), .B(n6585), .Z(n6587) );
  AND U7483 ( .A(n6588), .B(n6587), .Z(n6590) );
  XOR U7484 ( .A(n6591), .B(n6590), .Z(c[113]) );
  NAND U7485 ( .A(n6589), .B(sreg[113]), .Z(n6593) );
  OR U7486 ( .A(n6591), .B(n6590), .Z(n6592) );
  NAND U7487 ( .A(n6593), .B(n6592), .Z(n7037) );
  XNOR U7488 ( .A(n7037), .B(sreg[114]), .Z(n7039) );
  NAND U7489 ( .A(n6595), .B(n6594), .Z(n6599) );
  NAND U7490 ( .A(n6597), .B(n6596), .Z(n6598) );
  NAND U7491 ( .A(n6599), .B(n6598), .Z(n6812) );
  NAND U7492 ( .A(n6601), .B(n6600), .Z(n6605) );
  NANDN U7493 ( .A(n6603), .B(n6602), .Z(n6604) );
  NAND U7494 ( .A(n6605), .B(n6604), .Z(n6809) );
  OR U7495 ( .A(n6607), .B(n6606), .Z(n6611) );
  OR U7496 ( .A(n6609), .B(n6608), .Z(n6610) );
  NAND U7497 ( .A(n6611), .B(n6610), .Z(n6818) );
  NAND U7498 ( .A(n6613), .B(n6612), .Z(n6617) );
  NANDN U7499 ( .A(n6615), .B(n6614), .Z(n6616) );
  NAND U7500 ( .A(n6617), .B(n6616), .Z(n6815) );
  NANDN U7501 ( .A(n6619), .B(n6618), .Z(n6623) );
  NAND U7502 ( .A(n6621), .B(n6620), .Z(n6622) );
  NAND U7503 ( .A(n6623), .B(n6622), .Z(n6838) );
  XOR U7504 ( .A(b[13]), .B(n20686), .Z(n6971) );
  OR U7505 ( .A(n6971), .B(n31550), .Z(n6630) );
  NAND U7506 ( .A(n6628), .B(n31874), .Z(n6629) );
  NAND U7507 ( .A(n6630), .B(n6629), .Z(n6886) );
  XOR U7508 ( .A(b[31]), .B(n15484), .Z(n6865) );
  NANDN U7509 ( .A(n6865), .B(n35313), .Z(n6633) );
  NAND U7510 ( .A(n6631), .B(n35311), .Z(n6632) );
  NAND U7511 ( .A(n6633), .B(n6632), .Z(n6883) );
  XOR U7512 ( .A(b[37]), .B(n14210), .Z(n6928) );
  NANDN U7513 ( .A(n6928), .B(n36311), .Z(n6636) );
  NANDN U7514 ( .A(n6634), .B(n36309), .Z(n6635) );
  AND U7515 ( .A(n6636), .B(n6635), .Z(n6884) );
  XNOR U7516 ( .A(n6883), .B(n6884), .Z(n6885) );
  XNOR U7517 ( .A(n6886), .B(n6885), .Z(n7019) );
  XOR U7518 ( .A(b[33]), .B(n14905), .Z(n6934) );
  NANDN U7519 ( .A(n6934), .B(n35620), .Z(n6639) );
  NAND U7520 ( .A(n6637), .B(n35621), .Z(n6638) );
  NAND U7521 ( .A(n6639), .B(n6638), .Z(n6910) );
  XOR U7522 ( .A(b[49]), .B(n10363), .Z(n6849) );
  OR U7523 ( .A(n6849), .B(n37756), .Z(n6642) );
  NAND U7524 ( .A(n6640), .B(n37652), .Z(n6641) );
  NAND U7525 ( .A(n6642), .B(n6641), .Z(n6907) );
  XOR U7526 ( .A(b[9]), .B(n22246), .Z(n6862) );
  NANDN U7527 ( .A(n6862), .B(n30509), .Z(n6645) );
  NANDN U7528 ( .A(n6643), .B(n30846), .Z(n6644) );
  AND U7529 ( .A(n6645), .B(n6644), .Z(n6908) );
  XNOR U7530 ( .A(n6907), .B(n6908), .Z(n6909) );
  XOR U7531 ( .A(n6910), .B(n6909), .Z(n7020) );
  XNOR U7532 ( .A(n7019), .B(n7020), .Z(n7021) );
  XNOR U7533 ( .A(n7022), .B(n7021), .Z(n6837) );
  XNOR U7534 ( .A(n6838), .B(n6837), .Z(n6840) );
  NAND U7535 ( .A(n35188), .B(n6646), .Z(n6648) );
  XOR U7536 ( .A(b[29]), .B(n15963), .Z(n6895) );
  OR U7537 ( .A(n6895), .B(n34968), .Z(n6647) );
  NAND U7538 ( .A(n6648), .B(n6647), .Z(n6916) );
  XOR U7539 ( .A(n31123), .B(n22289), .Z(n6937) );
  NAND U7540 ( .A(n6937), .B(n29949), .Z(n6651) );
  NAND U7541 ( .A(n6649), .B(n29948), .Z(n6650) );
  NAND U7542 ( .A(n6651), .B(n6650), .Z(n6913) );
  XOR U7543 ( .A(b[5]), .B(n22964), .Z(n6901) );
  OR U7544 ( .A(n6901), .B(n29363), .Z(n6654) );
  NANDN U7545 ( .A(n6652), .B(n29864), .Z(n6653) );
  AND U7546 ( .A(n6654), .B(n6653), .Z(n6914) );
  XNOR U7547 ( .A(n6913), .B(n6914), .Z(n6915) );
  XNOR U7548 ( .A(n6916), .B(n6915), .Z(n7009) );
  OR U7549 ( .A(n6656), .B(n6655), .Z(n6660) );
  OR U7550 ( .A(n6658), .B(n6657), .Z(n6659) );
  AND U7551 ( .A(n6660), .B(n6659), .Z(n7007) );
  NANDN U7552 ( .A(n6662), .B(n6661), .Z(n6666) );
  NAND U7553 ( .A(n6664), .B(n6663), .Z(n6665) );
  NAND U7554 ( .A(n6666), .B(n6665), .Z(n7008) );
  XOR U7555 ( .A(n6840), .B(n6839), .Z(n7031) );
  NAND U7556 ( .A(n6668), .B(n6667), .Z(n6672) );
  NANDN U7557 ( .A(n6670), .B(n6669), .Z(n6671) );
  NAND U7558 ( .A(n6672), .B(n6671), .Z(n7032) );
  XNOR U7559 ( .A(n7031), .B(n7032), .Z(n7033) );
  NANDN U7560 ( .A(n6674), .B(n6673), .Z(n6678) );
  NAND U7561 ( .A(n6676), .B(n6675), .Z(n6677) );
  AND U7562 ( .A(n6678), .B(n6677), .Z(n7034) );
  XOR U7563 ( .A(n7033), .B(n7034), .Z(n6824) );
  OR U7564 ( .A(n6684), .B(n6683), .Z(n6688) );
  NAND U7565 ( .A(n6686), .B(n6685), .Z(n6687) );
  NAND U7566 ( .A(n6688), .B(n6687), .Z(n6832) );
  NANDN U7567 ( .A(n6690), .B(n6689), .Z(n6694) );
  NAND U7568 ( .A(n6692), .B(n6691), .Z(n6693) );
  AND U7569 ( .A(n6694), .B(n6693), .Z(n7025) );
  OR U7570 ( .A(n6696), .B(n6695), .Z(n6700) );
  NAND U7571 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U7572 ( .A(n6700), .B(n6699), .Z(n7026) );
  XNOR U7573 ( .A(n7025), .B(n7026), .Z(n7027) );
  XOR U7574 ( .A(n7027), .B(n7028), .Z(n6831) );
  XNOR U7575 ( .A(n6832), .B(n6831), .Z(n6833) );
  XNOR U7576 ( .A(b[21]), .B(a[30]), .Z(n6974) );
  OR U7577 ( .A(n6974), .B(n33634), .Z(n6707) );
  NANDN U7578 ( .A(n6705), .B(n33464), .Z(n6706) );
  NAND U7579 ( .A(n6707), .B(n6706), .Z(n6880) );
  XNOR U7580 ( .A(b[17]), .B(n19513), .Z(n6980) );
  NAND U7581 ( .A(n6980), .B(n32543), .Z(n6710) );
  NAND U7582 ( .A(n6708), .B(n32541), .Z(n6709) );
  NAND U7583 ( .A(n6710), .B(n6709), .Z(n6877) );
  NAND U7584 ( .A(n33283), .B(n6711), .Z(n6713) );
  XOR U7585 ( .A(n33020), .B(n18841), .Z(n6925) );
  NANDN U7586 ( .A(n33021), .B(n6925), .Z(n6712) );
  AND U7587 ( .A(n6713), .B(n6712), .Z(n6878) );
  XNOR U7588 ( .A(n6877), .B(n6878), .Z(n6879) );
  XNOR U7589 ( .A(n6880), .B(n6879), .Z(n6983) );
  NANDN U7590 ( .A(n966), .B(a[50]), .Z(n6714) );
  XOR U7591 ( .A(n29232), .B(n6714), .Z(n6716) );
  IV U7592 ( .A(a[49]), .Z(n23852) );
  NANDN U7593 ( .A(n23852), .B(n966), .Z(n6715) );
  AND U7594 ( .A(n6716), .B(n6715), .Z(n6964) );
  NAND U7595 ( .A(n6717), .B(n37469), .Z(n6719) );
  XOR U7596 ( .A(n978), .B(n10854), .Z(n6959) );
  NAND U7597 ( .A(n6959), .B(n37471), .Z(n6718) );
  NAND U7598 ( .A(n6719), .B(n6718), .Z(n6962) );
  XNOR U7599 ( .A(n979), .B(b[50]), .Z(n37803) );
  NANDN U7600 ( .A(n986), .B(n37803), .Z(n6963) );
  XNOR U7601 ( .A(n6962), .B(n6963), .Z(n6965) );
  XOR U7602 ( .A(n6964), .B(n6965), .Z(n6984) );
  XNOR U7603 ( .A(n6983), .B(n6984), .Z(n6985) );
  NANDN U7604 ( .A(n6721), .B(n6720), .Z(n6725) );
  NAND U7605 ( .A(n6723), .B(n6722), .Z(n6724) );
  AND U7606 ( .A(n6725), .B(n6724), .Z(n6986) );
  XNOR U7607 ( .A(n6985), .B(n6986), .Z(n6992) );
  OR U7608 ( .A(n6727), .B(n6726), .Z(n6731) );
  NAND U7609 ( .A(n6729), .B(n6728), .Z(n6730) );
  NAND U7610 ( .A(n6731), .B(n6730), .Z(n6989) );
  NANDN U7611 ( .A(n6733), .B(n6732), .Z(n6737) );
  NAND U7612 ( .A(n6735), .B(n6734), .Z(n6736) );
  NAND U7613 ( .A(n6737), .B(n6736), .Z(n6990) );
  XNOR U7614 ( .A(n6989), .B(n6990), .Z(n6991) );
  XOR U7615 ( .A(n6992), .B(n6991), .Z(n7004) );
  OR U7616 ( .A(n6739), .B(n6738), .Z(n6743) );
  OR U7617 ( .A(n6741), .B(n6740), .Z(n6742) );
  NAND U7618 ( .A(n6743), .B(n6742), .Z(n7016) );
  XNOR U7619 ( .A(b[35]), .B(a[16]), .Z(n6868) );
  NANDN U7620 ( .A(n6868), .B(n35985), .Z(n6746) );
  NANDN U7621 ( .A(n6744), .B(n35986), .Z(n6745) );
  NAND U7622 ( .A(n6746), .B(n6745), .Z(n6946) );
  XNOR U7623 ( .A(b[45]), .B(n11406), .Z(n6892) );
  NAND U7624 ( .A(n6892), .B(n37261), .Z(n6749) );
  NANDN U7625 ( .A(n6747), .B(n37262), .Z(n6748) );
  NAND U7626 ( .A(n6749), .B(n6748), .Z(n6943) );
  XOR U7627 ( .A(b[11]), .B(n21149), .Z(n6968) );
  OR U7628 ( .A(n6968), .B(n31369), .Z(n6752) );
  NAND U7629 ( .A(n6750), .B(n31119), .Z(n6751) );
  AND U7630 ( .A(n6752), .B(n6751), .Z(n6944) );
  XNOR U7631 ( .A(n6943), .B(n6944), .Z(n6945) );
  XOR U7632 ( .A(n6946), .B(n6945), .Z(n7014) );
  XOR U7633 ( .A(n977), .B(n11986), .Z(n6889) );
  NAND U7634 ( .A(n6889), .B(n37068), .Z(n6755) );
  NAND U7635 ( .A(n6753), .B(n37069), .Z(n6754) );
  NAND U7636 ( .A(n6755), .B(n6754), .Z(n6846) );
  XOR U7637 ( .A(b[39]), .B(n13106), .Z(n6931) );
  NANDN U7638 ( .A(n6931), .B(n36553), .Z(n6758) );
  NAND U7639 ( .A(n6756), .B(n36643), .Z(n6757) );
  NAND U7640 ( .A(n6758), .B(n6757), .Z(n6843) );
  XNOR U7641 ( .A(b[41]), .B(a[10]), .Z(n6940) );
  OR U7642 ( .A(n6940), .B(n36905), .Z(n6761) );
  NAND U7643 ( .A(n6759), .B(n36807), .Z(n6760) );
  AND U7644 ( .A(n6761), .B(n6760), .Z(n6844) );
  XNOR U7645 ( .A(n6843), .B(n6844), .Z(n6845) );
  XNOR U7646 ( .A(n6846), .B(n6845), .Z(n7013) );
  XOR U7647 ( .A(n7014), .B(n7013), .Z(n7015) );
  XNOR U7648 ( .A(n7016), .B(n7015), .Z(n7002) );
  XNOR U7649 ( .A(n972), .B(a[36]), .Z(n6977) );
  NANDN U7650 ( .A(n32010), .B(n6977), .Z(n6764) );
  NANDN U7651 ( .A(n6762), .B(n32011), .Z(n6763) );
  NAND U7652 ( .A(n6764), .B(n6763), .Z(n6922) );
  NAND U7653 ( .A(n34044), .B(n6765), .Z(n6767) );
  XOR U7654 ( .A(n34510), .B(n17702), .Z(n6898) );
  NANDN U7655 ( .A(n33867), .B(n6898), .Z(n6766) );
  NAND U7656 ( .A(n6767), .B(n6766), .Z(n6919) );
  XNOR U7657 ( .A(b[25]), .B(n17133), .Z(n6953) );
  NANDN U7658 ( .A(n34219), .B(n6953), .Z(n6770) );
  NAND U7659 ( .A(n6768), .B(n34217), .Z(n6769) );
  AND U7660 ( .A(n6770), .B(n6769), .Z(n6920) );
  XNOR U7661 ( .A(n6919), .B(n6920), .Z(n6921) );
  XOR U7662 ( .A(n6922), .B(n6921), .Z(n6949) );
  NANDN U7663 ( .A(n6772), .B(n6771), .Z(n6874) );
  NANDN U7664 ( .A(n6773), .B(n34848), .Z(n6775) );
  XOR U7665 ( .A(b[27]), .B(n16508), .Z(n6859) );
  NANDN U7666 ( .A(n6859), .B(n34618), .Z(n6774) );
  NAND U7667 ( .A(n6775), .B(n6774), .Z(n6872) );
  XNOR U7668 ( .A(n967), .B(a[48]), .Z(n6904) );
  NAND U7669 ( .A(n6904), .B(n28939), .Z(n6778) );
  NANDN U7670 ( .A(n6776), .B(n28938), .Z(n6777) );
  AND U7671 ( .A(n6778), .B(n6777), .Z(n6871) );
  XNOR U7672 ( .A(n6872), .B(n6871), .Z(n6873) );
  XNOR U7673 ( .A(n6874), .B(n6873), .Z(n6950) );
  XNOR U7674 ( .A(n6949), .B(n6950), .Z(n6952) );
  NANDN U7675 ( .A(n6780), .B(n6779), .Z(n6784) );
  NAND U7676 ( .A(n6782), .B(n6781), .Z(n6783) );
  AND U7677 ( .A(n6784), .B(n6783), .Z(n6951) );
  XOR U7678 ( .A(n6952), .B(n6951), .Z(n7001) );
  XOR U7679 ( .A(n7004), .B(n7003), .Z(n6998) );
  NANDN U7680 ( .A(n6786), .B(n6785), .Z(n6790) );
  NANDN U7681 ( .A(n6788), .B(n6787), .Z(n6789) );
  NAND U7682 ( .A(n6790), .B(n6789), .Z(n6995) );
  OR U7683 ( .A(n6792), .B(n6791), .Z(n6796) );
  NANDN U7684 ( .A(n6794), .B(n6793), .Z(n6795) );
  NAND U7685 ( .A(n6796), .B(n6795), .Z(n6996) );
  XNOR U7686 ( .A(n6995), .B(n6996), .Z(n6997) );
  XOR U7687 ( .A(n6998), .B(n6997), .Z(n6834) );
  XOR U7688 ( .A(n6833), .B(n6834), .Z(n6821) );
  XNOR U7689 ( .A(n6822), .B(n6821), .Z(n6823) );
  XOR U7690 ( .A(n6824), .B(n6823), .Z(n6828) );
  NANDN U7691 ( .A(n6798), .B(n6797), .Z(n6802) );
  OR U7692 ( .A(n6800), .B(n6799), .Z(n6801) );
  NAND U7693 ( .A(n6802), .B(n6801), .Z(n6825) );
  NAND U7694 ( .A(n6804), .B(n6803), .Z(n6808) );
  OR U7695 ( .A(n6806), .B(n6805), .Z(n6807) );
  NAND U7696 ( .A(n6808), .B(n6807), .Z(n6826) );
  XNOR U7697 ( .A(n6825), .B(n6826), .Z(n6827) );
  XNOR U7698 ( .A(n6828), .B(n6827), .Z(n6816) );
  XNOR U7699 ( .A(n6815), .B(n6816), .Z(n6817) );
  XNOR U7700 ( .A(n6818), .B(n6817), .Z(n6810) );
  XNOR U7701 ( .A(n6809), .B(n6810), .Z(n6811) );
  XOR U7702 ( .A(n6812), .B(n6811), .Z(n7038) );
  XOR U7703 ( .A(n7039), .B(n7038), .Z(c[114]) );
  NANDN U7704 ( .A(n6810), .B(n6809), .Z(n6814) );
  NAND U7705 ( .A(n6812), .B(n6811), .Z(n6813) );
  NAND U7706 ( .A(n6814), .B(n6813), .Z(n7050) );
  NANDN U7707 ( .A(n6816), .B(n6815), .Z(n6820) );
  NAND U7708 ( .A(n6818), .B(n6817), .Z(n6819) );
  NAND U7709 ( .A(n6820), .B(n6819), .Z(n7048) );
  NANDN U7710 ( .A(n6826), .B(n6825), .Z(n6830) );
  NANDN U7711 ( .A(n6828), .B(n6827), .Z(n6829) );
  NAND U7712 ( .A(n6830), .B(n6829), .Z(n7054) );
  XNOR U7713 ( .A(n7053), .B(n7054), .Z(n7055) );
  NAND U7714 ( .A(n6832), .B(n6831), .Z(n6836) );
  OR U7715 ( .A(n6834), .B(n6833), .Z(n6835) );
  NAND U7716 ( .A(n6836), .B(n6835), .Z(n7259) );
  NAND U7717 ( .A(n6838), .B(n6837), .Z(n6842) );
  NANDN U7718 ( .A(n6840), .B(n6839), .Z(n6841) );
  NAND U7719 ( .A(n6842), .B(n6841), .Z(n7254) );
  NANDN U7720 ( .A(n6844), .B(n6843), .Z(n6848) );
  NAND U7721 ( .A(n6846), .B(n6845), .Z(n6847) );
  NAND U7722 ( .A(n6848), .B(n6847), .Z(n7091) );
  XOR U7723 ( .A(n979), .B(n10524), .Z(n7105) );
  NANDN U7724 ( .A(n37756), .B(n7105), .Z(n6851) );
  NANDN U7725 ( .A(n6849), .B(n37652), .Z(n6850) );
  NAND U7726 ( .A(n6851), .B(n6850), .Z(n7228) );
  XNOR U7727 ( .A(n980), .B(a[0]), .Z(n6854) );
  XNOR U7728 ( .A(n980), .B(b[49]), .Z(n6853) );
  XNOR U7729 ( .A(n980), .B(b[50]), .Z(n6852) );
  AND U7730 ( .A(n6853), .B(n6852), .Z(n37802) );
  NAND U7731 ( .A(n6854), .B(n37802), .Z(n6856) );
  XOR U7732 ( .A(n980), .B(n10457), .Z(n7096) );
  NAND U7733 ( .A(n37803), .B(n7096), .Z(n6855) );
  NAND U7734 ( .A(n6856), .B(n6855), .Z(n7227) );
  XNOR U7735 ( .A(n7228), .B(n7227), .Z(n7185) );
  NOR U7736 ( .A(b[49]), .B(b[50]), .Z(n6857) );
  OR U7737 ( .A(n6857), .B(n986), .Z(n6858) );
  NANDN U7738 ( .A(n979), .B(b[50]), .Z(n37868) );
  AND U7739 ( .A(n37868), .B(b[51]), .Z(n38024) );
  AND U7740 ( .A(n6858), .B(n38024), .Z(n7183) );
  NANDN U7741 ( .A(n6859), .B(n34848), .Z(n6861) );
  XNOR U7742 ( .A(n35375), .B(a[25]), .Z(n7218) );
  NAND U7743 ( .A(n34618), .B(n7218), .Z(n6860) );
  NAND U7744 ( .A(n6861), .B(n6860), .Z(n7182) );
  XOR U7745 ( .A(n7183), .B(n7182), .Z(n7184) );
  XOR U7746 ( .A(n7185), .B(n7184), .Z(n7090) );
  XOR U7747 ( .A(b[9]), .B(n21996), .Z(n7200) );
  NANDN U7748 ( .A(n7200), .B(n30509), .Z(n6864) );
  NANDN U7749 ( .A(n6862), .B(n30846), .Z(n6863) );
  NAND U7750 ( .A(n6864), .B(n6863), .Z(n7191) );
  XOR U7751 ( .A(b[31]), .B(n16220), .Z(n7093) );
  NANDN U7752 ( .A(n7093), .B(n35313), .Z(n6867) );
  NANDN U7753 ( .A(n6865), .B(n35311), .Z(n6866) );
  NAND U7754 ( .A(n6867), .B(n6866), .Z(n7188) );
  XNOR U7755 ( .A(b[35]), .B(a[17]), .Z(n7140) );
  NANDN U7756 ( .A(n7140), .B(n35985), .Z(n6870) );
  NANDN U7757 ( .A(n6868), .B(n35986), .Z(n6869) );
  AND U7758 ( .A(n6870), .B(n6869), .Z(n7189) );
  XNOR U7759 ( .A(n7188), .B(n7189), .Z(n7190) );
  XNOR U7760 ( .A(n7191), .B(n7190), .Z(n7089) );
  XOR U7761 ( .A(n7090), .B(n7089), .Z(n7092) );
  XNOR U7762 ( .A(n7091), .B(n7092), .Z(n7164) );
  NANDN U7763 ( .A(n6872), .B(n6871), .Z(n6876) );
  NAND U7764 ( .A(n6874), .B(n6873), .Z(n6875) );
  NAND U7765 ( .A(n6876), .B(n6875), .Z(n7161) );
  NANDN U7766 ( .A(n6878), .B(n6877), .Z(n6882) );
  NAND U7767 ( .A(n6880), .B(n6879), .Z(n6881) );
  NAND U7768 ( .A(n6882), .B(n6881), .Z(n7162) );
  XNOR U7769 ( .A(n7161), .B(n7162), .Z(n7163) );
  XOR U7770 ( .A(n7164), .B(n7163), .Z(n7170) );
  NANDN U7771 ( .A(n6884), .B(n6883), .Z(n6888) );
  NAND U7772 ( .A(n6886), .B(n6885), .Z(n6887) );
  NAND U7773 ( .A(n6888), .B(n6887), .Z(n7158) );
  NAND U7774 ( .A(n37069), .B(n6889), .Z(n6891) );
  XNOR U7775 ( .A(n977), .B(a[9]), .Z(n7176) );
  NAND U7776 ( .A(n7176), .B(n37068), .Z(n6890) );
  NAND U7777 ( .A(n6891), .B(n6890), .Z(n7122) );
  NAND U7778 ( .A(n37262), .B(n6892), .Z(n6894) );
  XNOR U7779 ( .A(b[45]), .B(a[7]), .Z(n7221) );
  NANDN U7780 ( .A(n7221), .B(n37261), .Z(n6893) );
  NAND U7781 ( .A(n6894), .B(n6893), .Z(n7120) );
  NANDN U7782 ( .A(n6895), .B(n35188), .Z(n6897) );
  XOR U7783 ( .A(b[29]), .B(n16269), .Z(n7229) );
  OR U7784 ( .A(n7229), .B(n34968), .Z(n6896) );
  NAND U7785 ( .A(n6897), .B(n6896), .Z(n7121) );
  XNOR U7786 ( .A(n7120), .B(n7121), .Z(n7123) );
  XOR U7787 ( .A(n7122), .B(n7123), .Z(n7155) );
  NAND U7788 ( .A(n34044), .B(n6898), .Z(n6900) );
  XOR U7789 ( .A(n34510), .B(n18003), .Z(n7131) );
  NANDN U7790 ( .A(n33867), .B(n7131), .Z(n6899) );
  NAND U7791 ( .A(n6900), .B(n6899), .Z(n7152) );
  XOR U7792 ( .A(b[5]), .B(n23149), .Z(n7099) );
  OR U7793 ( .A(n7099), .B(n29363), .Z(n6903) );
  NANDN U7794 ( .A(n6901), .B(n29864), .Z(n6902) );
  NAND U7795 ( .A(n6903), .B(n6902), .Z(n7149) );
  XOR U7796 ( .A(b[3]), .B(n23852), .Z(n7232) );
  NANDN U7797 ( .A(n7232), .B(n28939), .Z(n6906) );
  NAND U7798 ( .A(n6904), .B(n28938), .Z(n6905) );
  AND U7799 ( .A(n6906), .B(n6905), .Z(n7150) );
  XNOR U7800 ( .A(n7149), .B(n7150), .Z(n7151) );
  XOR U7801 ( .A(n7152), .B(n7151), .Z(n7156) );
  XNOR U7802 ( .A(n7155), .B(n7156), .Z(n7157) );
  XOR U7803 ( .A(n7158), .B(n7157), .Z(n7167) );
  NANDN U7804 ( .A(n6908), .B(n6907), .Z(n6912) );
  NAND U7805 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7806 ( .A(n6912), .B(n6911), .Z(n7168) );
  XNOR U7807 ( .A(n7167), .B(n7168), .Z(n7169) );
  XNOR U7808 ( .A(n7170), .B(n7169), .Z(n7073) );
  NANDN U7809 ( .A(n6914), .B(n6913), .Z(n6918) );
  NAND U7810 ( .A(n6916), .B(n6915), .Z(n6917) );
  NAND U7811 ( .A(n6918), .B(n6917), .Z(n7080) );
  NANDN U7812 ( .A(n6920), .B(n6919), .Z(n6924) );
  NAND U7813 ( .A(n6922), .B(n6921), .Z(n6923) );
  NAND U7814 ( .A(n6924), .B(n6923), .Z(n7085) );
  NAND U7815 ( .A(n33283), .B(n6925), .Z(n6927) );
  XNOR U7816 ( .A(n33020), .B(a[33]), .Z(n7146) );
  NANDN U7817 ( .A(n33021), .B(n7146), .Z(n6926) );
  NAND U7818 ( .A(n6927), .B(n6926), .Z(n7215) );
  XOR U7819 ( .A(b[37]), .B(n13976), .Z(n7206) );
  NANDN U7820 ( .A(n7206), .B(n36311), .Z(n6930) );
  NANDN U7821 ( .A(n6928), .B(n36309), .Z(n6929) );
  NAND U7822 ( .A(n6930), .B(n6929), .Z(n7212) );
  XOR U7823 ( .A(b[39]), .B(n13509), .Z(n7194) );
  NANDN U7824 ( .A(n7194), .B(n36553), .Z(n6933) );
  NANDN U7825 ( .A(n6931), .B(n36643), .Z(n6932) );
  AND U7826 ( .A(n6933), .B(n6932), .Z(n7213) );
  XNOR U7827 ( .A(n7212), .B(n7213), .Z(n7214) );
  XNOR U7828 ( .A(n7215), .B(n7214), .Z(n7083) );
  XOR U7829 ( .A(b[33]), .B(n15113), .Z(n7137) );
  NANDN U7830 ( .A(n7137), .B(n35620), .Z(n6936) );
  NANDN U7831 ( .A(n6934), .B(n35621), .Z(n6935) );
  NAND U7832 ( .A(n6936), .B(n6935), .Z(n7238) );
  XOR U7833 ( .A(n31123), .B(n22579), .Z(n7179) );
  NAND U7834 ( .A(n7179), .B(n29949), .Z(n6939) );
  NAND U7835 ( .A(n29948), .B(n6937), .Z(n6938) );
  NAND U7836 ( .A(n6939), .B(n6938), .Z(n7235) );
  XNOR U7837 ( .A(b[41]), .B(a[11]), .Z(n7209) );
  OR U7838 ( .A(n7209), .B(n36905), .Z(n6942) );
  NANDN U7839 ( .A(n6940), .B(n36807), .Z(n6941) );
  AND U7840 ( .A(n6942), .B(n6941), .Z(n7236) );
  XNOR U7841 ( .A(n7235), .B(n7236), .Z(n7237) );
  XOR U7842 ( .A(n7238), .B(n7237), .Z(n7084) );
  XOR U7843 ( .A(n7083), .B(n7084), .Z(n7086) );
  XNOR U7844 ( .A(n7085), .B(n7086), .Z(n7077) );
  NANDN U7845 ( .A(n6944), .B(n6943), .Z(n6948) );
  NAND U7846 ( .A(n6946), .B(n6945), .Z(n6947) );
  AND U7847 ( .A(n6948), .B(n6947), .Z(n7078) );
  XNOR U7848 ( .A(n7077), .B(n7078), .Z(n7079) );
  XNOR U7849 ( .A(n7080), .B(n7079), .Z(n7071) );
  XOR U7850 ( .A(n7071), .B(n7072), .Z(n7074) );
  XOR U7851 ( .A(n7073), .B(n7074), .Z(n7251) );
  XNOR U7852 ( .A(b[25]), .B(n17960), .Z(n7173) );
  NANDN U7853 ( .A(n34219), .B(n7173), .Z(n6955) );
  NAND U7854 ( .A(n34217), .B(n6953), .Z(n6954) );
  NAND U7855 ( .A(n6955), .B(n6954), .Z(n7127) );
  NANDN U7856 ( .A(n966), .B(a[51]), .Z(n6956) );
  XOR U7857 ( .A(n29232), .B(n6956), .Z(n6958) );
  IV U7858 ( .A(a[50]), .Z(n24671) );
  NANDN U7859 ( .A(n24671), .B(n966), .Z(n6957) );
  AND U7860 ( .A(n6958), .B(n6957), .Z(n7124) );
  NAND U7861 ( .A(n37469), .B(n6959), .Z(n6961) );
  XOR U7862 ( .A(n978), .B(n11202), .Z(n7224) );
  NAND U7863 ( .A(n7224), .B(n37471), .Z(n6960) );
  AND U7864 ( .A(n6961), .B(n6960), .Z(n7125) );
  XNOR U7865 ( .A(n7124), .B(n7125), .Z(n7126) );
  XNOR U7866 ( .A(n7127), .B(n7126), .Z(n7241) );
  NANDN U7867 ( .A(n6963), .B(n6962), .Z(n6967) );
  NAND U7868 ( .A(n6965), .B(n6964), .Z(n6966) );
  NAND U7869 ( .A(n6967), .B(n6966), .Z(n7242) );
  XNOR U7870 ( .A(n7241), .B(n7242), .Z(n7243) );
  XOR U7871 ( .A(b[11]), .B(n21441), .Z(n7197) );
  OR U7872 ( .A(n7197), .B(n31369), .Z(n6970) );
  NANDN U7873 ( .A(n6968), .B(n31119), .Z(n6969) );
  NAND U7874 ( .A(n6970), .B(n6969), .Z(n7111) );
  XOR U7875 ( .A(b[13]), .B(n20867), .Z(n7203) );
  OR U7876 ( .A(n7203), .B(n31550), .Z(n6973) );
  NANDN U7877 ( .A(n6971), .B(n31874), .Z(n6972) );
  NAND U7878 ( .A(n6973), .B(n6972), .Z(n7108) );
  XNOR U7879 ( .A(b[21]), .B(a[31]), .Z(n7128) );
  OR U7880 ( .A(n7128), .B(n33634), .Z(n6976) );
  NANDN U7881 ( .A(n6974), .B(n33464), .Z(n6975) );
  AND U7882 ( .A(n6976), .B(n6975), .Z(n7109) );
  XNOR U7883 ( .A(n7108), .B(n7109), .Z(n7110) );
  XNOR U7884 ( .A(n7111), .B(n7110), .Z(n7117) );
  NAND U7885 ( .A(n6977), .B(n32011), .Z(n6979) );
  XNOR U7886 ( .A(n972), .B(a[37]), .Z(n7143) );
  NANDN U7887 ( .A(n32010), .B(n7143), .Z(n6978) );
  NAND U7888 ( .A(n6979), .B(n6978), .Z(n7115) );
  XNOR U7889 ( .A(b[17]), .B(n20315), .Z(n7134) );
  NAND U7890 ( .A(n7134), .B(n32543), .Z(n6982) );
  NAND U7891 ( .A(n6980), .B(n32541), .Z(n6981) );
  AND U7892 ( .A(n6982), .B(n6981), .Z(n7114) );
  XNOR U7893 ( .A(n7115), .B(n7114), .Z(n7116) );
  XOR U7894 ( .A(n7117), .B(n7116), .Z(n7244) );
  XOR U7895 ( .A(n7243), .B(n7244), .Z(n7245) );
  NANDN U7896 ( .A(n6984), .B(n6983), .Z(n6988) );
  NAND U7897 ( .A(n6986), .B(n6985), .Z(n6987) );
  NAND U7898 ( .A(n6988), .B(n6987), .Z(n7246) );
  XOR U7899 ( .A(n7245), .B(n7246), .Z(n7247) );
  NANDN U7900 ( .A(n6990), .B(n6989), .Z(n6994) );
  NANDN U7901 ( .A(n6992), .B(n6991), .Z(n6993) );
  AND U7902 ( .A(n6994), .B(n6993), .Z(n7248) );
  XNOR U7903 ( .A(n7247), .B(n7248), .Z(n7252) );
  XOR U7904 ( .A(n7251), .B(n7252), .Z(n7253) );
  XOR U7905 ( .A(n7254), .B(n7253), .Z(n7258) );
  NANDN U7906 ( .A(n6996), .B(n6995), .Z(n7000) );
  NANDN U7907 ( .A(n6998), .B(n6997), .Z(n6999) );
  NAND U7908 ( .A(n7000), .B(n6999), .Z(n7059) );
  OR U7909 ( .A(n7002), .B(n7001), .Z(n7006) );
  NANDN U7910 ( .A(n7004), .B(n7003), .Z(n7005) );
  AND U7911 ( .A(n7006), .B(n7005), .Z(n7060) );
  XNOR U7912 ( .A(n7059), .B(n7060), .Z(n7061) );
  OR U7913 ( .A(n7008), .B(n7007), .Z(n7012) );
  NANDN U7914 ( .A(n7010), .B(n7009), .Z(n7011) );
  AND U7915 ( .A(n7012), .B(n7011), .Z(n7068) );
  NANDN U7916 ( .A(n7014), .B(n7013), .Z(n7018) );
  OR U7917 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U7918 ( .A(n7018), .B(n7017), .Z(n7065) );
  NANDN U7919 ( .A(n7020), .B(n7019), .Z(n7024) );
  NANDN U7920 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U7921 ( .A(n7024), .B(n7023), .Z(n7066) );
  XNOR U7922 ( .A(n7065), .B(n7066), .Z(n7067) );
  XNOR U7923 ( .A(n7061), .B(n7062), .Z(n7257) );
  XNOR U7924 ( .A(n7258), .B(n7257), .Z(n7260) );
  XNOR U7925 ( .A(n7259), .B(n7260), .Z(n7265) );
  OR U7926 ( .A(n7026), .B(n7025), .Z(n7030) );
  OR U7927 ( .A(n7028), .B(n7027), .Z(n7029) );
  NAND U7928 ( .A(n7030), .B(n7029), .Z(n7263) );
  NANDN U7929 ( .A(n7032), .B(n7031), .Z(n7036) );
  NAND U7930 ( .A(n7034), .B(n7033), .Z(n7035) );
  NAND U7931 ( .A(n7036), .B(n7035), .Z(n7264) );
  XNOR U7932 ( .A(n7263), .B(n7264), .Z(n7266) );
  XOR U7933 ( .A(n7265), .B(n7266), .Z(n7056) );
  XOR U7934 ( .A(n7055), .B(n7056), .Z(n7047) );
  XOR U7935 ( .A(n7048), .B(n7047), .Z(n7049) );
  XNOR U7936 ( .A(n7050), .B(n7049), .Z(n7042) );
  XNOR U7937 ( .A(n7042), .B(sreg[115]), .Z(n7044) );
  NAND U7938 ( .A(n7037), .B(sreg[114]), .Z(n7041) );
  OR U7939 ( .A(n7039), .B(n7038), .Z(n7040) );
  AND U7940 ( .A(n7041), .B(n7040), .Z(n7043) );
  XOR U7941 ( .A(n7044), .B(n7043), .Z(c[115]) );
  NAND U7942 ( .A(n7042), .B(sreg[115]), .Z(n7046) );
  OR U7943 ( .A(n7044), .B(n7043), .Z(n7045) );
  NAND U7944 ( .A(n7046), .B(n7045), .Z(n7506) );
  XNOR U7945 ( .A(n7506), .B(sreg[116]), .Z(n7508) );
  NAND U7946 ( .A(n7048), .B(n7047), .Z(n7052) );
  NAND U7947 ( .A(n7050), .B(n7049), .Z(n7051) );
  NAND U7948 ( .A(n7052), .B(n7051), .Z(n7272) );
  NANDN U7949 ( .A(n7054), .B(n7053), .Z(n7058) );
  NAND U7950 ( .A(n7056), .B(n7055), .Z(n7057) );
  NAND U7951 ( .A(n7058), .B(n7057), .Z(n7269) );
  NANDN U7952 ( .A(n7060), .B(n7059), .Z(n7064) );
  NANDN U7953 ( .A(n7062), .B(n7061), .Z(n7063) );
  NAND U7954 ( .A(n7064), .B(n7063), .Z(n7501) );
  OR U7955 ( .A(n7066), .B(n7065), .Z(n7070) );
  OR U7956 ( .A(n7068), .B(n7067), .Z(n7069) );
  NAND U7957 ( .A(n7070), .B(n7069), .Z(n7500) );
  NANDN U7958 ( .A(n7072), .B(n7071), .Z(n7076) );
  OR U7959 ( .A(n7074), .B(n7073), .Z(n7075) );
  NAND U7960 ( .A(n7076), .B(n7075), .Z(n7503) );
  XOR U7961 ( .A(n7502), .B(n7503), .Z(n7497) );
  NANDN U7962 ( .A(n7078), .B(n7077), .Z(n7082) );
  NAND U7963 ( .A(n7080), .B(n7079), .Z(n7081) );
  NAND U7964 ( .A(n7082), .B(n7081), .Z(n7284) );
  NANDN U7965 ( .A(n7084), .B(n7083), .Z(n7088) );
  OR U7966 ( .A(n7086), .B(n7085), .Z(n7087) );
  NAND U7967 ( .A(n7088), .B(n7087), .Z(n7281) );
  XNOR U7968 ( .A(n7281), .B(n7282), .Z(n7283) );
  XOR U7969 ( .A(n7284), .B(n7283), .Z(n7484) );
  NANDN U7970 ( .A(n7093), .B(n35311), .Z(n7095) );
  XNOR U7971 ( .A(n973), .B(a[22]), .Z(n7436) );
  NAND U7972 ( .A(n7436), .B(n35313), .Z(n7094) );
  AND U7973 ( .A(n7095), .B(n7094), .Z(n7448) );
  XOR U7974 ( .A(b[51]), .B(n10363), .Z(n7469) );
  NANDN U7975 ( .A(n7469), .B(n37803), .Z(n7098) );
  NAND U7976 ( .A(n7096), .B(n37802), .Z(n7097) );
  AND U7977 ( .A(n7098), .B(n7097), .Z(n7449) );
  XOR U7978 ( .A(n7448), .B(n7449), .Z(n7450) );
  XOR U7979 ( .A(b[5]), .B(n23447), .Z(n7311) );
  OR U7980 ( .A(n7311), .B(n29363), .Z(n7101) );
  NANDN U7981 ( .A(n7099), .B(n29864), .Z(n7100) );
  AND U7982 ( .A(n7101), .B(n7100), .Z(n7451) );
  XNOR U7983 ( .A(n7450), .B(n7451), .Z(n7383) );
  NANDN U7984 ( .A(n966), .B(a[52]), .Z(n7102) );
  XOR U7985 ( .A(n29232), .B(n7102), .Z(n7104) );
  IV U7986 ( .A(a[51]), .Z(n24288) );
  NANDN U7987 ( .A(n24288), .B(n966), .Z(n7103) );
  AND U7988 ( .A(n7104), .B(n7103), .Z(n7316) );
  XOR U7989 ( .A(b[49]), .B(n10854), .Z(n7400) );
  OR U7990 ( .A(n7400), .B(n37756), .Z(n7107) );
  NAND U7991 ( .A(n7105), .B(n37652), .Z(n7106) );
  NAND U7992 ( .A(n7107), .B(n7106), .Z(n7314) );
  XNOR U7993 ( .A(n980), .B(b[52]), .Z(n37940) );
  NANDN U7994 ( .A(n986), .B(n37940), .Z(n7315) );
  XNOR U7995 ( .A(n7314), .B(n7315), .Z(n7317) );
  XOR U7996 ( .A(n7316), .B(n7317), .Z(n7382) );
  XOR U7997 ( .A(n7383), .B(n7382), .Z(n7384) );
  NANDN U7998 ( .A(n7109), .B(n7108), .Z(n7113) );
  NAND U7999 ( .A(n7111), .B(n7110), .Z(n7112) );
  AND U8000 ( .A(n7113), .B(n7112), .Z(n7385) );
  XNOR U8001 ( .A(n7384), .B(n7385), .Z(n7290) );
  NANDN U8002 ( .A(n7115), .B(n7114), .Z(n7119) );
  NAND U8003 ( .A(n7117), .B(n7116), .Z(n7118) );
  NAND U8004 ( .A(n7119), .B(n7118), .Z(n7287) );
  XNOR U8005 ( .A(n7287), .B(n7288), .Z(n7289) );
  XOR U8006 ( .A(n7290), .B(n7289), .Z(n7483) );
  XNOR U8007 ( .A(b[21]), .B(a[32]), .Z(n7338) );
  OR U8008 ( .A(n7338), .B(n33634), .Z(n7130) );
  NANDN U8009 ( .A(n7128), .B(n33464), .Z(n7129) );
  NAND U8010 ( .A(n7130), .B(n7129), .Z(n7415) );
  NAND U8011 ( .A(n34044), .B(n7131), .Z(n7133) );
  XOR U8012 ( .A(n34510), .B(n18804), .Z(n7439) );
  NANDN U8013 ( .A(n33867), .B(n7439), .Z(n7132) );
  NAND U8014 ( .A(n7133), .B(n7132), .Z(n7412) );
  XNOR U8015 ( .A(b[17]), .B(a[36]), .Z(n7329) );
  NANDN U8016 ( .A(n7329), .B(n32543), .Z(n7136) );
  NAND U8017 ( .A(n7134), .B(n32541), .Z(n7135) );
  AND U8018 ( .A(n7136), .B(n7135), .Z(n7413) );
  XNOR U8019 ( .A(n7412), .B(n7413), .Z(n7414) );
  XOR U8020 ( .A(n7415), .B(n7414), .Z(n7295) );
  XOR U8021 ( .A(b[33]), .B(n15484), .Z(n7341) );
  NANDN U8022 ( .A(n7341), .B(n35620), .Z(n7139) );
  NANDN U8023 ( .A(n7137), .B(n35621), .Z(n7138) );
  NAND U8024 ( .A(n7139), .B(n7138), .Z(n7457) );
  XNOR U8025 ( .A(b[35]), .B(a[18]), .Z(n7308) );
  NANDN U8026 ( .A(n7308), .B(n35985), .Z(n7142) );
  NANDN U8027 ( .A(n7140), .B(n35986), .Z(n7141) );
  NAND U8028 ( .A(n7142), .B(n7141), .Z(n7454) );
  XOR U8029 ( .A(b[15]), .B(n20686), .Z(n7460) );
  OR U8030 ( .A(n7460), .B(n32010), .Z(n7145) );
  NAND U8031 ( .A(n7143), .B(n32011), .Z(n7144) );
  AND U8032 ( .A(n7145), .B(n7144), .Z(n7455) );
  XNOR U8033 ( .A(n7454), .B(n7455), .Z(n7456) );
  XOR U8034 ( .A(n7457), .B(n7456), .Z(n7293) );
  NAND U8035 ( .A(n7146), .B(n33283), .Z(n7148) );
  XNOR U8036 ( .A(n33020), .B(a[34]), .Z(n7332) );
  NANDN U8037 ( .A(n33021), .B(n7332), .Z(n7147) );
  NAND U8038 ( .A(n7148), .B(n7147), .Z(n7294) );
  XNOR U8039 ( .A(n7293), .B(n7294), .Z(n7296) );
  XNOR U8040 ( .A(n7295), .B(n7296), .Z(n7363) );
  NANDN U8041 ( .A(n7150), .B(n7149), .Z(n7154) );
  NAND U8042 ( .A(n7152), .B(n7151), .Z(n7153) );
  AND U8043 ( .A(n7154), .B(n7153), .Z(n7362) );
  XNOR U8044 ( .A(n7363), .B(n7362), .Z(n7364) );
  XOR U8045 ( .A(n7365), .B(n7364), .Z(n7344) );
  NANDN U8046 ( .A(n7156), .B(n7155), .Z(n7160) );
  NANDN U8047 ( .A(n7158), .B(n7157), .Z(n7159) );
  NAND U8048 ( .A(n7160), .B(n7159), .Z(n7345) );
  XNOR U8049 ( .A(n7344), .B(n7345), .Z(n7346) );
  NANDN U8050 ( .A(n7162), .B(n7161), .Z(n7166) );
  NAND U8051 ( .A(n7164), .B(n7163), .Z(n7165) );
  NAND U8052 ( .A(n7166), .B(n7165), .Z(n7347) );
  XNOR U8053 ( .A(n7346), .B(n7347), .Z(n7482) );
  XNOR U8054 ( .A(n7483), .B(n7482), .Z(n7485) );
  XNOR U8055 ( .A(n7484), .B(n7485), .Z(n7490) );
  NANDN U8056 ( .A(n7168), .B(n7167), .Z(n7172) );
  NANDN U8057 ( .A(n7170), .B(n7169), .Z(n7171) );
  NAND U8058 ( .A(n7172), .B(n7171), .Z(n7359) );
  XNOR U8059 ( .A(b[25]), .B(n17702), .Z(n7394) );
  NANDN U8060 ( .A(n34219), .B(n7394), .Z(n7175) );
  NAND U8061 ( .A(n34217), .B(n7173), .Z(n7174) );
  NAND U8062 ( .A(n7175), .B(n7174), .Z(n7427) );
  XOR U8063 ( .A(b[43]), .B(n12555), .Z(n7406) );
  NANDN U8064 ( .A(n7406), .B(n37068), .Z(n7178) );
  NAND U8065 ( .A(n7176), .B(n37069), .Z(n7177) );
  NAND U8066 ( .A(n7178), .B(n7177), .Z(n7424) );
  XOR U8067 ( .A(n31123), .B(n22964), .Z(n7335) );
  NAND U8068 ( .A(n7335), .B(n29949), .Z(n7181) );
  NAND U8069 ( .A(n29948), .B(n7179), .Z(n7180) );
  AND U8070 ( .A(n7181), .B(n7180), .Z(n7425) );
  XNOR U8071 ( .A(n7424), .B(n7425), .Z(n7426) );
  XOR U8072 ( .A(n7427), .B(n7426), .Z(n7381) );
  OR U8073 ( .A(n7183), .B(n7182), .Z(n7187) );
  NAND U8074 ( .A(n7185), .B(n7184), .Z(n7186) );
  NAND U8075 ( .A(n7187), .B(n7186), .Z(n7378) );
  NANDN U8076 ( .A(n7189), .B(n7188), .Z(n7193) );
  NAND U8077 ( .A(n7191), .B(n7190), .Z(n7192) );
  NAND U8078 ( .A(n7193), .B(n7192), .Z(n7379) );
  XNOR U8079 ( .A(n7378), .B(n7379), .Z(n7380) );
  XOR U8080 ( .A(n7381), .B(n7380), .Z(n7353) );
  XOR U8081 ( .A(b[39]), .B(n14210), .Z(n7430) );
  NANDN U8082 ( .A(n7430), .B(n36553), .Z(n7196) );
  NANDN U8083 ( .A(n7194), .B(n36643), .Z(n7195) );
  NAND U8084 ( .A(n7196), .B(n7195), .Z(n7323) );
  XOR U8085 ( .A(b[11]), .B(n22246), .Z(n7463) );
  OR U8086 ( .A(n7463), .B(n31369), .Z(n7199) );
  NANDN U8087 ( .A(n7197), .B(n31119), .Z(n7198) );
  NAND U8088 ( .A(n7199), .B(n7198), .Z(n7320) );
  XOR U8089 ( .A(b[9]), .B(n22289), .Z(n7326) );
  NANDN U8090 ( .A(n7326), .B(n30509), .Z(n7202) );
  NANDN U8091 ( .A(n7200), .B(n30846), .Z(n7201) );
  AND U8092 ( .A(n7202), .B(n7201), .Z(n7321) );
  XNOR U8093 ( .A(n7320), .B(n7321), .Z(n7322) );
  XNOR U8094 ( .A(n7323), .B(n7322), .Z(n7368) );
  XOR U8095 ( .A(b[13]), .B(n21149), .Z(n7466) );
  OR U8096 ( .A(n7466), .B(n31550), .Z(n7205) );
  NANDN U8097 ( .A(n7203), .B(n31874), .Z(n7204) );
  NAND U8098 ( .A(n7205), .B(n7204), .Z(n7302) );
  XOR U8099 ( .A(b[37]), .B(n14259), .Z(n7305) );
  NANDN U8100 ( .A(n7305), .B(n36311), .Z(n7208) );
  NANDN U8101 ( .A(n7206), .B(n36309), .Z(n7207) );
  NAND U8102 ( .A(n7208), .B(n7207), .Z(n7299) );
  XNOR U8103 ( .A(b[41]), .B(a[12]), .Z(n7433) );
  OR U8104 ( .A(n7433), .B(n36905), .Z(n7211) );
  NANDN U8105 ( .A(n7209), .B(n36807), .Z(n7210) );
  AND U8106 ( .A(n7211), .B(n7210), .Z(n7300) );
  XNOR U8107 ( .A(n7299), .B(n7300), .Z(n7301) );
  XOR U8108 ( .A(n7302), .B(n7301), .Z(n7369) );
  XNOR U8109 ( .A(n7368), .B(n7369), .Z(n7370) );
  NANDN U8110 ( .A(n7213), .B(n7212), .Z(n7217) );
  NAND U8111 ( .A(n7215), .B(n7214), .Z(n7216) );
  AND U8112 ( .A(n7217), .B(n7216), .Z(n7371) );
  XNOR U8113 ( .A(n7370), .B(n7371), .Z(n7350) );
  NAND U8114 ( .A(n7218), .B(n34848), .Z(n7220) );
  XOR U8115 ( .A(b[27]), .B(n17133), .Z(n7479) );
  NANDN U8116 ( .A(n7479), .B(n34618), .Z(n7219) );
  NAND U8117 ( .A(n7220), .B(n7219), .Z(n7421) );
  XNOR U8118 ( .A(b[45]), .B(a[8]), .Z(n7445) );
  NANDN U8119 ( .A(n7445), .B(n37261), .Z(n7223) );
  NANDN U8120 ( .A(n7221), .B(n37262), .Z(n7222) );
  NAND U8121 ( .A(n7223), .B(n7222), .Z(n7418) );
  NAND U8122 ( .A(n37469), .B(n7224), .Z(n7226) );
  XOR U8123 ( .A(n978), .B(n11406), .Z(n7397) );
  NAND U8124 ( .A(n7397), .B(n37471), .Z(n7225) );
  AND U8125 ( .A(n7226), .B(n7225), .Z(n7419) );
  XNOR U8126 ( .A(n7418), .B(n7419), .Z(n7420) );
  XNOR U8127 ( .A(n7421), .B(n7420), .Z(n7374) );
  NAND U8128 ( .A(n7228), .B(n7227), .Z(n7391) );
  NANDN U8129 ( .A(n7229), .B(n35188), .Z(n7231) );
  XNOR U8130 ( .A(n35540), .B(a[24]), .Z(n7409) );
  NANDN U8131 ( .A(n34968), .B(n7409), .Z(n7230) );
  NAND U8132 ( .A(n7231), .B(n7230), .Z(n7389) );
  XNOR U8133 ( .A(n967), .B(a[50]), .Z(n7403) );
  NAND U8134 ( .A(n7403), .B(n28939), .Z(n7234) );
  NANDN U8135 ( .A(n7232), .B(n28938), .Z(n7233) );
  AND U8136 ( .A(n7234), .B(n7233), .Z(n7388) );
  XNOR U8137 ( .A(n7389), .B(n7388), .Z(n7390) );
  XNOR U8138 ( .A(n7391), .B(n7390), .Z(n7375) );
  XNOR U8139 ( .A(n7374), .B(n7375), .Z(n7376) );
  NANDN U8140 ( .A(n7236), .B(n7235), .Z(n7240) );
  NAND U8141 ( .A(n7238), .B(n7237), .Z(n7239) );
  AND U8142 ( .A(n7240), .B(n7239), .Z(n7377) );
  XNOR U8143 ( .A(n7376), .B(n7377), .Z(n7351) );
  XOR U8144 ( .A(n7350), .B(n7351), .Z(n7352) );
  XOR U8145 ( .A(n7353), .B(n7352), .Z(n7356) );
  XNOR U8146 ( .A(n7356), .B(n7357), .Z(n7358) );
  XNOR U8147 ( .A(n7359), .B(n7358), .Z(n7488) );
  OR U8148 ( .A(n7246), .B(n7245), .Z(n7250) );
  NAND U8149 ( .A(n7248), .B(n7247), .Z(n7249) );
  NAND U8150 ( .A(n7250), .B(n7249), .Z(n7489) );
  XOR U8151 ( .A(n7488), .B(n7489), .Z(n7491) );
  XOR U8152 ( .A(n7490), .B(n7491), .Z(n7494) );
  OR U8153 ( .A(n7252), .B(n7251), .Z(n7256) );
  NANDN U8154 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U8155 ( .A(n7256), .B(n7255), .Z(n7495) );
  XOR U8156 ( .A(n7494), .B(n7495), .Z(n7496) );
  XNOR U8157 ( .A(n7497), .B(n7496), .Z(n7275) );
  NAND U8158 ( .A(n7258), .B(n7257), .Z(n7262) );
  NANDN U8159 ( .A(n7260), .B(n7259), .Z(n7261) );
  NAND U8160 ( .A(n7262), .B(n7261), .Z(n7276) );
  XOR U8161 ( .A(n7275), .B(n7276), .Z(n7278) );
  NANDN U8162 ( .A(n7264), .B(n7263), .Z(n7268) );
  NAND U8163 ( .A(n7266), .B(n7265), .Z(n7267) );
  NAND U8164 ( .A(n7268), .B(n7267), .Z(n7277) );
  XOR U8165 ( .A(n7278), .B(n7277), .Z(n7270) );
  XNOR U8166 ( .A(n7269), .B(n7270), .Z(n7271) );
  XOR U8167 ( .A(n7272), .B(n7271), .Z(n7507) );
  XOR U8168 ( .A(n7508), .B(n7507), .Z(c[116]) );
  NANDN U8169 ( .A(n7270), .B(n7269), .Z(n7274) );
  NAND U8170 ( .A(n7272), .B(n7271), .Z(n7273) );
  NAND U8171 ( .A(n7274), .B(n7273), .Z(n7519) );
  NANDN U8172 ( .A(n7276), .B(n7275), .Z(n7280) );
  OR U8173 ( .A(n7278), .B(n7277), .Z(n7279) );
  NAND U8174 ( .A(n7280), .B(n7279), .Z(n7516) );
  NANDN U8175 ( .A(n7282), .B(n7281), .Z(n7286) );
  NANDN U8176 ( .A(n7284), .B(n7283), .Z(n7285) );
  NAND U8177 ( .A(n7286), .B(n7285), .Z(n7735) );
  NANDN U8178 ( .A(n7288), .B(n7287), .Z(n7292) );
  NANDN U8179 ( .A(n7290), .B(n7289), .Z(n7291) );
  NAND U8180 ( .A(n7292), .B(n7291), .Z(n7734) );
  OR U8181 ( .A(n7294), .B(n7293), .Z(n7298) );
  OR U8182 ( .A(n7296), .B(n7295), .Z(n7297) );
  NAND U8183 ( .A(n7298), .B(n7297), .Z(n7529) );
  NANDN U8184 ( .A(n7300), .B(n7299), .Z(n7304) );
  NAND U8185 ( .A(n7302), .B(n7301), .Z(n7303) );
  NAND U8186 ( .A(n7304), .B(n7303), .Z(n7664) );
  XOR U8187 ( .A(b[37]), .B(n14514), .Z(n7677) );
  NANDN U8188 ( .A(n7677), .B(n36311), .Z(n7307) );
  NANDN U8189 ( .A(n7305), .B(n36309), .Z(n7306) );
  NAND U8190 ( .A(n7307), .B(n7306), .Z(n7561) );
  XNOR U8191 ( .A(b[35]), .B(a[19]), .Z(n7609) );
  NANDN U8192 ( .A(n7609), .B(n35985), .Z(n7310) );
  NANDN U8193 ( .A(n7308), .B(n35986), .Z(n7309) );
  NAND U8194 ( .A(n7310), .B(n7309), .Z(n7558) );
  XOR U8195 ( .A(b[5]), .B(n23852), .Z(n7585) );
  OR U8196 ( .A(n7585), .B(n29363), .Z(n7313) );
  NANDN U8197 ( .A(n7311), .B(n29864), .Z(n7312) );
  AND U8198 ( .A(n7313), .B(n7312), .Z(n7559) );
  XNOR U8199 ( .A(n7558), .B(n7559), .Z(n7560) );
  XNOR U8200 ( .A(n7561), .B(n7560), .Z(n7662) );
  NANDN U8201 ( .A(n7315), .B(n7314), .Z(n7319) );
  NAND U8202 ( .A(n7317), .B(n7316), .Z(n7318) );
  NAND U8203 ( .A(n7319), .B(n7318), .Z(n7663) );
  XOR U8204 ( .A(n7662), .B(n7663), .Z(n7665) );
  XOR U8205 ( .A(n7664), .B(n7665), .Z(n7528) );
  XNOR U8206 ( .A(n7529), .B(n7528), .Z(n7531) );
  NANDN U8207 ( .A(n7321), .B(n7320), .Z(n7325) );
  NAND U8208 ( .A(n7323), .B(n7322), .Z(n7324) );
  NAND U8209 ( .A(n7325), .B(n7324), .Z(n7670) );
  XOR U8210 ( .A(b[9]), .B(n22579), .Z(n7615) );
  NANDN U8211 ( .A(n7615), .B(n30509), .Z(n7328) );
  NANDN U8212 ( .A(n7326), .B(n30846), .Z(n7327) );
  NAND U8213 ( .A(n7328), .B(n7327), .Z(n7606) );
  XNOR U8214 ( .A(b[17]), .B(a[37]), .Z(n7540) );
  NANDN U8215 ( .A(n7540), .B(n32543), .Z(n7331) );
  NANDN U8216 ( .A(n7329), .B(n32541), .Z(n7330) );
  NAND U8217 ( .A(n7331), .B(n7330), .Z(n7603) );
  NAND U8218 ( .A(n7332), .B(n33283), .Z(n7334) );
  XOR U8219 ( .A(n33020), .B(n20315), .Z(n7674) );
  NANDN U8220 ( .A(n33021), .B(n7674), .Z(n7333) );
  AND U8221 ( .A(n7334), .B(n7333), .Z(n7604) );
  XNOR U8222 ( .A(n7603), .B(n7604), .Z(n7605) );
  XNOR U8223 ( .A(n7606), .B(n7605), .Z(n7668) );
  XOR U8224 ( .A(n31123), .B(n23149), .Z(n7582) );
  NAND U8225 ( .A(n7582), .B(n29949), .Z(n7337) );
  NAND U8226 ( .A(n29948), .B(n7335), .Z(n7336) );
  NAND U8227 ( .A(n7337), .B(n7336), .Z(n7692) );
  XNOR U8228 ( .A(b[21]), .B(a[33]), .Z(n7594) );
  OR U8229 ( .A(n7594), .B(n33634), .Z(n7340) );
  NANDN U8230 ( .A(n7338), .B(n33464), .Z(n7339) );
  NAND U8231 ( .A(n7340), .B(n7339), .Z(n7689) );
  XOR U8232 ( .A(b[33]), .B(n16220), .Z(n7591) );
  NANDN U8233 ( .A(n7591), .B(n35620), .Z(n7343) );
  NANDN U8234 ( .A(n7341), .B(n35621), .Z(n7342) );
  AND U8235 ( .A(n7343), .B(n7342), .Z(n7690) );
  XNOR U8236 ( .A(n7689), .B(n7690), .Z(n7691) );
  XOR U8237 ( .A(n7692), .B(n7691), .Z(n7669) );
  XOR U8238 ( .A(n7668), .B(n7669), .Z(n7671) );
  XOR U8239 ( .A(n7670), .B(n7671), .Z(n7530) );
  XNOR U8240 ( .A(n7531), .B(n7530), .Z(n7733) );
  XNOR U8241 ( .A(n7734), .B(n7733), .Z(n7736) );
  XOR U8242 ( .A(n7735), .B(n7736), .Z(n7740) );
  NANDN U8243 ( .A(n7345), .B(n7344), .Z(n7349) );
  NANDN U8244 ( .A(n7347), .B(n7346), .Z(n7348) );
  NAND U8245 ( .A(n7349), .B(n7348), .Z(n7737) );
  OR U8246 ( .A(n7351), .B(n7350), .Z(n7355) );
  NANDN U8247 ( .A(n7353), .B(n7352), .Z(n7354) );
  NAND U8248 ( .A(n7355), .B(n7354), .Z(n7738) );
  XNOR U8249 ( .A(n7737), .B(n7738), .Z(n7739) );
  XNOR U8250 ( .A(n7740), .B(n7739), .Z(n7730) );
  NANDN U8251 ( .A(n7357), .B(n7356), .Z(n7361) );
  NAND U8252 ( .A(n7359), .B(n7358), .Z(n7360) );
  NAND U8253 ( .A(n7361), .B(n7360), .Z(n7728) );
  NANDN U8254 ( .A(n7363), .B(n7362), .Z(n7367) );
  NANDN U8255 ( .A(n7365), .B(n7364), .Z(n7366) );
  NAND U8256 ( .A(n7367), .B(n7366), .Z(n7653) );
  NANDN U8257 ( .A(n7369), .B(n7368), .Z(n7373) );
  NAND U8258 ( .A(n7371), .B(n7370), .Z(n7372) );
  NAND U8259 ( .A(n7373), .B(n7372), .Z(n7650) );
  XNOR U8260 ( .A(n7650), .B(n7651), .Z(n7652) );
  XNOR U8261 ( .A(n7653), .B(n7652), .Z(n7726) );
  OR U8262 ( .A(n7383), .B(n7382), .Z(n7387) );
  NAND U8263 ( .A(n7385), .B(n7384), .Z(n7386) );
  NAND U8264 ( .A(n7387), .B(n7386), .Z(n7644) );
  NANDN U8265 ( .A(n7389), .B(n7388), .Z(n7393) );
  NAND U8266 ( .A(n7391), .B(n7390), .Z(n7392) );
  NAND U8267 ( .A(n7393), .B(n7392), .Z(n7714) );
  XNOR U8268 ( .A(b[25]), .B(n18003), .Z(n7600) );
  NANDN U8269 ( .A(n34219), .B(n7600), .Z(n7396) );
  NAND U8270 ( .A(n34217), .B(n7394), .Z(n7395) );
  NAND U8271 ( .A(n7396), .B(n7395), .Z(n7641) );
  NAND U8272 ( .A(n37469), .B(n7397), .Z(n7399) );
  XOR U8273 ( .A(n978), .B(n11694), .Z(n7546) );
  NAND U8274 ( .A(n7546), .B(n37471), .Z(n7398) );
  NAND U8275 ( .A(n7399), .B(n7398), .Z(n7638) );
  XOR U8276 ( .A(b[49]), .B(n11202), .Z(n7555) );
  OR U8277 ( .A(n7555), .B(n37756), .Z(n7402) );
  NANDN U8278 ( .A(n7400), .B(n37652), .Z(n7401) );
  AND U8279 ( .A(n7402), .B(n7401), .Z(n7639) );
  XNOR U8280 ( .A(n7638), .B(n7639), .Z(n7640) );
  XOR U8281 ( .A(n7641), .B(n7640), .Z(n7707) );
  XOR U8282 ( .A(b[3]), .B(n24288), .Z(n7623) );
  NANDN U8283 ( .A(n7623), .B(n28939), .Z(n7405) );
  NAND U8284 ( .A(n7403), .B(n28938), .Z(n7404) );
  NAND U8285 ( .A(n7405), .B(n7404), .Z(n7698) );
  XOR U8286 ( .A(b[43]), .B(n12830), .Z(n7680) );
  NANDN U8287 ( .A(n7680), .B(n37068), .Z(n7408) );
  NANDN U8288 ( .A(n7406), .B(n37069), .Z(n7407) );
  NAND U8289 ( .A(n7408), .B(n7407), .Z(n7695) );
  NAND U8290 ( .A(n7409), .B(n35188), .Z(n7411) );
  XNOR U8291 ( .A(n35540), .B(a[25]), .Z(n7620) );
  NANDN U8292 ( .A(n34968), .B(n7620), .Z(n7410) );
  AND U8293 ( .A(n7411), .B(n7410), .Z(n7696) );
  XNOR U8294 ( .A(n7695), .B(n7696), .Z(n7697) );
  XOR U8295 ( .A(n7698), .B(n7697), .Z(n7705) );
  NANDN U8296 ( .A(n7413), .B(n7412), .Z(n7417) );
  NAND U8297 ( .A(n7415), .B(n7414), .Z(n7416) );
  NAND U8298 ( .A(n7417), .B(n7416), .Z(n7706) );
  XNOR U8299 ( .A(n7705), .B(n7706), .Z(n7708) );
  XNOR U8300 ( .A(n7707), .B(n7708), .Z(n7712) );
  NANDN U8301 ( .A(n7419), .B(n7418), .Z(n7423) );
  NAND U8302 ( .A(n7421), .B(n7420), .Z(n7422) );
  AND U8303 ( .A(n7423), .B(n7422), .Z(n7711) );
  XNOR U8304 ( .A(n7712), .B(n7711), .Z(n7713) );
  XNOR U8305 ( .A(n7714), .B(n7713), .Z(n7645) );
  XNOR U8306 ( .A(n7644), .B(n7645), .Z(n7646) );
  NANDN U8307 ( .A(n7425), .B(n7424), .Z(n7429) );
  NAND U8308 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U8309 ( .A(n7429), .B(n7428), .Z(n7659) );
  XOR U8310 ( .A(n976), .B(n13976), .Z(n7570) );
  NAND U8311 ( .A(n7570), .B(n36553), .Z(n7432) );
  NANDN U8312 ( .A(n7430), .B(n36643), .Z(n7431) );
  NAND U8313 ( .A(n7432), .B(n7431), .Z(n7635) );
  XNOR U8314 ( .A(b[41]), .B(a[13]), .Z(n7549) );
  OR U8315 ( .A(n7549), .B(n36905), .Z(n7435) );
  NANDN U8316 ( .A(n7433), .B(n36807), .Z(n7434) );
  NAND U8317 ( .A(n7435), .B(n7434), .Z(n7632) );
  XOR U8318 ( .A(b[31]), .B(n16269), .Z(n7579) );
  NANDN U8319 ( .A(n7579), .B(n35313), .Z(n7438) );
  NAND U8320 ( .A(n7436), .B(n35311), .Z(n7437) );
  AND U8321 ( .A(n7438), .B(n7437), .Z(n7633) );
  XNOR U8322 ( .A(n7632), .B(n7633), .Z(n7634) );
  XOR U8323 ( .A(n7635), .B(n7634), .Z(n7657) );
  NAND U8324 ( .A(n34044), .B(n7439), .Z(n7441) );
  XOR U8325 ( .A(n34510), .B(n18639), .Z(n7588) );
  NANDN U8326 ( .A(n33867), .B(n7588), .Z(n7440) );
  NAND U8327 ( .A(n7441), .B(n7440), .Z(n7704) );
  NANDN U8328 ( .A(n966), .B(a[53]), .Z(n7442) );
  XOR U8329 ( .A(n29232), .B(n7442), .Z(n7444) );
  IV U8330 ( .A(a[52]), .Z(n25134) );
  NANDN U8331 ( .A(n25134), .B(n966), .Z(n7443) );
  AND U8332 ( .A(n7444), .B(n7443), .Z(n7701) );
  XNOR U8333 ( .A(b[45]), .B(a[9]), .Z(n7543) );
  NANDN U8334 ( .A(n7543), .B(n37261), .Z(n7447) );
  NANDN U8335 ( .A(n7445), .B(n37262), .Z(n7446) );
  AND U8336 ( .A(n7447), .B(n7446), .Z(n7702) );
  XNOR U8337 ( .A(n7701), .B(n7702), .Z(n7703) );
  XNOR U8338 ( .A(n7704), .B(n7703), .Z(n7656) );
  XOR U8339 ( .A(n7657), .B(n7656), .Z(n7658) );
  XNOR U8340 ( .A(n7659), .B(n7658), .Z(n7535) );
  OR U8341 ( .A(n7449), .B(n7448), .Z(n7453) );
  NANDN U8342 ( .A(n7451), .B(n7450), .Z(n7452) );
  NAND U8343 ( .A(n7453), .B(n7452), .Z(n7534) );
  XNOR U8344 ( .A(n7535), .B(n7534), .Z(n7536) );
  NANDN U8345 ( .A(n7455), .B(n7454), .Z(n7459) );
  NAND U8346 ( .A(n7457), .B(n7456), .Z(n7458) );
  NAND U8347 ( .A(n7459), .B(n7458), .Z(n7720) );
  XOR U8348 ( .A(b[15]), .B(n20867), .Z(n7552) );
  OR U8349 ( .A(n7552), .B(n32010), .Z(n7462) );
  NANDN U8350 ( .A(n7460), .B(n32011), .Z(n7461) );
  NAND U8351 ( .A(n7462), .B(n7461), .Z(n7629) );
  XOR U8352 ( .A(b[11]), .B(n21996), .Z(n7612) );
  OR U8353 ( .A(n7612), .B(n31369), .Z(n7465) );
  NANDN U8354 ( .A(n7463), .B(n31119), .Z(n7464) );
  NAND U8355 ( .A(n7465), .B(n7464), .Z(n7626) );
  XOR U8356 ( .A(b[13]), .B(n21441), .Z(n7573) );
  OR U8357 ( .A(n7573), .B(n31550), .Z(n7468) );
  NANDN U8358 ( .A(n7466), .B(n31874), .Z(n7467) );
  AND U8359 ( .A(n7468), .B(n7467), .Z(n7627) );
  XNOR U8360 ( .A(n7626), .B(n7627), .Z(n7628) );
  XNOR U8361 ( .A(n7629), .B(n7628), .Z(n7718) );
  XOR U8362 ( .A(n980), .B(n10524), .Z(n7686) );
  NAND U8363 ( .A(n7686), .B(n37803), .Z(n7471) );
  NANDN U8364 ( .A(n7469), .B(n37802), .Z(n7470) );
  NAND U8365 ( .A(n7471), .B(n7470), .Z(n7619) );
  XOR U8366 ( .A(b[53]), .B(n10457), .Z(n7576) );
  ANDN U8367 ( .B(n37940), .A(n7576), .Z(n7476) );
  XNOR U8368 ( .A(n981), .B(a[0]), .Z(n7474) );
  XNOR U8369 ( .A(n981), .B(b[51]), .Z(n7473) );
  XNOR U8370 ( .A(n981), .B(b[52]), .Z(n7472) );
  AND U8371 ( .A(n7473), .B(n7472), .Z(n37941) );
  NAND U8372 ( .A(n7474), .B(n37941), .Z(n7475) );
  NANDN U8373 ( .A(n7476), .B(n7475), .Z(n7618) );
  XNOR U8374 ( .A(n7619), .B(n7618), .Z(n7567) );
  NOR U8375 ( .A(b[51]), .B(b[52]), .Z(n7477) );
  OR U8376 ( .A(n7477), .B(n986), .Z(n7478) );
  NANDN U8377 ( .A(n980), .B(b[52]), .Z(n38041) );
  AND U8378 ( .A(n38041), .B(b[53]), .Z(n38117) );
  IV U8379 ( .A(n38117), .Z(n38081) );
  ANDN U8380 ( .B(n7478), .A(n38081), .Z(n7565) );
  NANDN U8381 ( .A(n7479), .B(n34848), .Z(n7481) );
  XOR U8382 ( .A(b[27]), .B(n17960), .Z(n7597) );
  NANDN U8383 ( .A(n7597), .B(n34618), .Z(n7480) );
  NAND U8384 ( .A(n7481), .B(n7480), .Z(n7564) );
  XOR U8385 ( .A(n7565), .B(n7564), .Z(n7566) );
  XOR U8386 ( .A(n7567), .B(n7566), .Z(n7717) );
  XOR U8387 ( .A(n7718), .B(n7717), .Z(n7719) );
  XOR U8388 ( .A(n7720), .B(n7719), .Z(n7537) );
  XNOR U8389 ( .A(n7646), .B(n7647), .Z(n7723) );
  XNOR U8390 ( .A(n7724), .B(n7723), .Z(n7725) );
  XOR U8391 ( .A(n7726), .B(n7725), .Z(n7727) );
  XNOR U8392 ( .A(n7728), .B(n7727), .Z(n7729) );
  XOR U8393 ( .A(n7730), .B(n7729), .Z(n7746) );
  NAND U8394 ( .A(n7483), .B(n7482), .Z(n7487) );
  NANDN U8395 ( .A(n7485), .B(n7484), .Z(n7486) );
  NAND U8396 ( .A(n7487), .B(n7486), .Z(n7743) );
  NANDN U8397 ( .A(n7489), .B(n7488), .Z(n7493) );
  OR U8398 ( .A(n7491), .B(n7490), .Z(n7492) );
  NAND U8399 ( .A(n7493), .B(n7492), .Z(n7744) );
  XNOR U8400 ( .A(n7743), .B(n7744), .Z(n7745) );
  XNOR U8401 ( .A(n7746), .B(n7745), .Z(n7525) );
  NAND U8402 ( .A(n7495), .B(n7494), .Z(n7499) );
  NAND U8403 ( .A(n7497), .B(n7496), .Z(n7498) );
  NAND U8404 ( .A(n7499), .B(n7498), .Z(n7522) );
  OR U8405 ( .A(n7501), .B(n7500), .Z(n7505) );
  NANDN U8406 ( .A(n7503), .B(n7502), .Z(n7504) );
  NAND U8407 ( .A(n7505), .B(n7504), .Z(n7523) );
  XNOR U8408 ( .A(n7522), .B(n7523), .Z(n7524) );
  XOR U8409 ( .A(n7525), .B(n7524), .Z(n7517) );
  XOR U8410 ( .A(n7516), .B(n7517), .Z(n7518) );
  XNOR U8411 ( .A(n7519), .B(n7518), .Z(n7511) );
  XNOR U8412 ( .A(n7511), .B(sreg[117]), .Z(n7513) );
  NAND U8413 ( .A(n7506), .B(sreg[116]), .Z(n7510) );
  OR U8414 ( .A(n7508), .B(n7507), .Z(n7509) );
  AND U8415 ( .A(n7510), .B(n7509), .Z(n7512) );
  XOR U8416 ( .A(n7513), .B(n7512), .Z(c[117]) );
  NAND U8417 ( .A(n7511), .B(sreg[117]), .Z(n7515) );
  OR U8418 ( .A(n7513), .B(n7512), .Z(n7514) );
  NAND U8419 ( .A(n7515), .B(n7514), .Z(n7993) );
  XNOR U8420 ( .A(n7993), .B(sreg[118]), .Z(n7995) );
  OR U8421 ( .A(n7517), .B(n7516), .Z(n7521) );
  NAND U8422 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U8423 ( .A(n7521), .B(n7520), .Z(n7752) );
  NANDN U8424 ( .A(n7523), .B(n7522), .Z(n7527) );
  NANDN U8425 ( .A(n7525), .B(n7524), .Z(n7526) );
  NAND U8426 ( .A(n7527), .B(n7526), .Z(n7749) );
  NAND U8427 ( .A(n7529), .B(n7528), .Z(n7533) );
  NANDN U8428 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U8429 ( .A(n7533), .B(n7532), .Z(n7972) );
  OR U8430 ( .A(n7535), .B(n7534), .Z(n7539) );
  OR U8431 ( .A(n7537), .B(n7536), .Z(n7538) );
  NAND U8432 ( .A(n7539), .B(n7538), .Z(n7970) );
  XNOR U8433 ( .A(b[17]), .B(a[38]), .Z(n7801) );
  NANDN U8434 ( .A(n7801), .B(n32543), .Z(n7542) );
  NANDN U8435 ( .A(n7540), .B(n32541), .Z(n7541) );
  NAND U8436 ( .A(n7542), .B(n7541), .Z(n7859) );
  XNOR U8437 ( .A(b[45]), .B(n12555), .Z(n7874) );
  NAND U8438 ( .A(n7874), .B(n37261), .Z(n7545) );
  NANDN U8439 ( .A(n7543), .B(n37262), .Z(n7544) );
  NAND U8440 ( .A(n7545), .B(n7544), .Z(n7856) );
  NAND U8441 ( .A(n37469), .B(n7546), .Z(n7548) );
  XOR U8442 ( .A(b[47]), .B(n11986), .Z(n7877) );
  NANDN U8443 ( .A(n7877), .B(n37471), .Z(n7547) );
  AND U8444 ( .A(n7548), .B(n7547), .Z(n7857) );
  XNOR U8445 ( .A(n7856), .B(n7857), .Z(n7858) );
  XNOR U8446 ( .A(n7859), .B(n7858), .Z(n7761) );
  XNOR U8447 ( .A(b[41]), .B(a[14]), .Z(n7810) );
  OR U8448 ( .A(n7810), .B(n36905), .Z(n7551) );
  NANDN U8449 ( .A(n7549), .B(n36807), .Z(n7550) );
  NAND U8450 ( .A(n7551), .B(n7550), .Z(n7786) );
  XOR U8451 ( .A(b[15]), .B(n21149), .Z(n7804) );
  OR U8452 ( .A(n7804), .B(n32010), .Z(n7554) );
  NANDN U8453 ( .A(n7552), .B(n32011), .Z(n7553) );
  NAND U8454 ( .A(n7554), .B(n7553), .Z(n7783) );
  XOR U8455 ( .A(b[49]), .B(n11406), .Z(n7798) );
  OR U8456 ( .A(n7798), .B(n37756), .Z(n7557) );
  NANDN U8457 ( .A(n7555), .B(n37652), .Z(n7556) );
  AND U8458 ( .A(n7557), .B(n7556), .Z(n7784) );
  XNOR U8459 ( .A(n7783), .B(n7784), .Z(n7785) );
  XOR U8460 ( .A(n7786), .B(n7785), .Z(n7762) );
  XNOR U8461 ( .A(n7761), .B(n7762), .Z(n7763) );
  NANDN U8462 ( .A(n7559), .B(n7558), .Z(n7563) );
  NAND U8463 ( .A(n7561), .B(n7560), .Z(n7562) );
  AND U8464 ( .A(n7563), .B(n7562), .Z(n7764) );
  XNOR U8465 ( .A(n7763), .B(n7764), .Z(n7881) );
  OR U8466 ( .A(n7565), .B(n7564), .Z(n7569) );
  NAND U8467 ( .A(n7567), .B(n7566), .Z(n7568) );
  NAND U8468 ( .A(n7569), .B(n7568), .Z(n7960) );
  NAND U8469 ( .A(n36643), .B(n7570), .Z(n7572) );
  XNOR U8470 ( .A(n976), .B(a[16]), .Z(n7927) );
  NAND U8471 ( .A(n7927), .B(n36553), .Z(n7571) );
  NAND U8472 ( .A(n7572), .B(n7571), .Z(n7854) );
  NANDN U8473 ( .A(n7573), .B(n31874), .Z(n7575) );
  XNOR U8474 ( .A(n971), .B(a[42]), .Z(n7930) );
  NANDN U8475 ( .A(n31550), .B(n7930), .Z(n7574) );
  NAND U8476 ( .A(n7575), .B(n7574), .Z(n7852) );
  NANDN U8477 ( .A(n7576), .B(n37941), .Z(n7578) );
  XOR U8478 ( .A(b[53]), .B(n10363), .Z(n7908) );
  NANDN U8479 ( .A(n7908), .B(n37940), .Z(n7577) );
  NAND U8480 ( .A(n7578), .B(n7577), .Z(n7853) );
  XNOR U8481 ( .A(n7852), .B(n7853), .Z(n7855) );
  XOR U8482 ( .A(n7854), .B(n7855), .Z(n7776) );
  XOR U8483 ( .A(b[31]), .B(n16508), .Z(n7816) );
  NANDN U8484 ( .A(n7816), .B(n35313), .Z(n7581) );
  NANDN U8485 ( .A(n7579), .B(n35311), .Z(n7580) );
  NAND U8486 ( .A(n7581), .B(n7580), .Z(n7837) );
  XOR U8487 ( .A(n31123), .B(n23447), .Z(n7792) );
  NAND U8488 ( .A(n7792), .B(n29949), .Z(n7584) );
  NAND U8489 ( .A(n29948), .B(n7582), .Z(n7583) );
  NAND U8490 ( .A(n7584), .B(n7583), .Z(n7834) );
  XOR U8491 ( .A(b[5]), .B(n24671), .Z(n7868) );
  OR U8492 ( .A(n7868), .B(n29363), .Z(n7587) );
  NANDN U8493 ( .A(n7585), .B(n29864), .Z(n7586) );
  AND U8494 ( .A(n7587), .B(n7586), .Z(n7835) );
  XNOR U8495 ( .A(n7834), .B(n7835), .Z(n7836) );
  XNOR U8496 ( .A(n7837), .B(n7836), .Z(n7773) );
  NAND U8497 ( .A(n34044), .B(n7588), .Z(n7590) );
  XOR U8498 ( .A(n34510), .B(n18841), .Z(n7822) );
  NANDN U8499 ( .A(n33867), .B(n7822), .Z(n7589) );
  NAND U8500 ( .A(n7590), .B(n7589), .Z(n7905) );
  XOR U8501 ( .A(b[33]), .B(n15963), .Z(n7862) );
  NANDN U8502 ( .A(n7862), .B(n35620), .Z(n7593) );
  NANDN U8503 ( .A(n7591), .B(n35621), .Z(n7592) );
  NAND U8504 ( .A(n7593), .B(n7592), .Z(n7902) );
  XNOR U8505 ( .A(b[21]), .B(a[34]), .Z(n7807) );
  OR U8506 ( .A(n7807), .B(n33634), .Z(n7596) );
  NANDN U8507 ( .A(n7594), .B(n33464), .Z(n7595) );
  AND U8508 ( .A(n7596), .B(n7595), .Z(n7903) );
  XNOR U8509 ( .A(n7902), .B(n7903), .Z(n7904) );
  XOR U8510 ( .A(n7905), .B(n7904), .Z(n7782) );
  NANDN U8511 ( .A(n7597), .B(n34848), .Z(n7599) );
  XNOR U8512 ( .A(n35375), .B(a[28]), .Z(n7942) );
  NAND U8513 ( .A(n34618), .B(n7942), .Z(n7598) );
  NAND U8514 ( .A(n7599), .B(n7598), .Z(n7780) );
  XNOR U8515 ( .A(b[25]), .B(a[30]), .Z(n7825) );
  OR U8516 ( .A(n7825), .B(n34219), .Z(n7602) );
  NAND U8517 ( .A(n34217), .B(n7600), .Z(n7601) );
  AND U8518 ( .A(n7602), .B(n7601), .Z(n7779) );
  XNOR U8519 ( .A(n7780), .B(n7779), .Z(n7781) );
  XOR U8520 ( .A(n7782), .B(n7781), .Z(n7774) );
  XNOR U8521 ( .A(n7773), .B(n7774), .Z(n7775) );
  XNOR U8522 ( .A(n7776), .B(n7775), .Z(n7958) );
  NANDN U8523 ( .A(n7604), .B(n7603), .Z(n7608) );
  NAND U8524 ( .A(n7606), .B(n7605), .Z(n7607) );
  AND U8525 ( .A(n7608), .B(n7607), .Z(n7957) );
  XNOR U8526 ( .A(n7958), .B(n7957), .Z(n7959) );
  XOR U8527 ( .A(n7960), .B(n7959), .Z(n7880) );
  XNOR U8528 ( .A(n7881), .B(n7880), .Z(n7882) );
  XNOR U8529 ( .A(b[35]), .B(a[20]), .Z(n7795) );
  NANDN U8530 ( .A(n7795), .B(n35985), .Z(n7611) );
  NANDN U8531 ( .A(n7609), .B(n35986), .Z(n7610) );
  NAND U8532 ( .A(n7611), .B(n7610), .Z(n7831) );
  XOR U8533 ( .A(b[11]), .B(n22289), .Z(n7933) );
  OR U8534 ( .A(n7933), .B(n31369), .Z(n7614) );
  NANDN U8535 ( .A(n7612), .B(n31119), .Z(n7613) );
  NAND U8536 ( .A(n7614), .B(n7613), .Z(n7828) );
  XOR U8537 ( .A(b[9]), .B(n22964), .Z(n7789) );
  NANDN U8538 ( .A(n7789), .B(n30509), .Z(n7617) );
  NANDN U8539 ( .A(n7615), .B(n30846), .Z(n7616) );
  AND U8540 ( .A(n7617), .B(n7616), .Z(n7829) );
  XNOR U8541 ( .A(n7828), .B(n7829), .Z(n7830) );
  XNOR U8542 ( .A(n7831), .B(n7830), .Z(n7840) );
  AND U8543 ( .A(n7619), .B(n7618), .Z(n7849) );
  NAND U8544 ( .A(n7620), .B(n35188), .Z(n7622) );
  XOR U8545 ( .A(b[29]), .B(n17133), .Z(n7918) );
  OR U8546 ( .A(n7918), .B(n34968), .Z(n7621) );
  NAND U8547 ( .A(n7622), .B(n7621), .Z(n7847) );
  XOR U8548 ( .A(n967), .B(n25134), .Z(n7936) );
  NAND U8549 ( .A(n7936), .B(n28939), .Z(n7625) );
  NANDN U8550 ( .A(n7623), .B(n28938), .Z(n7624) );
  NAND U8551 ( .A(n7625), .B(n7624), .Z(n7846) );
  XNOR U8552 ( .A(n7847), .B(n7846), .Z(n7848) );
  XNOR U8553 ( .A(n7840), .B(n7841), .Z(n7842) );
  NANDN U8554 ( .A(n7627), .B(n7626), .Z(n7631) );
  NAND U8555 ( .A(n7629), .B(n7628), .Z(n7630) );
  AND U8556 ( .A(n7631), .B(n7630), .Z(n7843) );
  XNOR U8557 ( .A(n7842), .B(n7843), .Z(n7954) );
  NANDN U8558 ( .A(n7633), .B(n7632), .Z(n7637) );
  NAND U8559 ( .A(n7635), .B(n7634), .Z(n7636) );
  NAND U8560 ( .A(n7637), .B(n7636), .Z(n7952) );
  NANDN U8561 ( .A(n7639), .B(n7638), .Z(n7643) );
  NAND U8562 ( .A(n7641), .B(n7640), .Z(n7642) );
  AND U8563 ( .A(n7643), .B(n7642), .Z(n7951) );
  XNOR U8564 ( .A(n7952), .B(n7951), .Z(n7953) );
  XOR U8565 ( .A(n7954), .B(n7953), .Z(n7883) );
  XNOR U8566 ( .A(n7882), .B(n7883), .Z(n7969) );
  XOR U8567 ( .A(n7970), .B(n7969), .Z(n7971) );
  XNOR U8568 ( .A(n7972), .B(n7971), .Z(n7978) );
  NANDN U8569 ( .A(n7645), .B(n7644), .Z(n7649) );
  NANDN U8570 ( .A(n7647), .B(n7646), .Z(n7648) );
  NAND U8571 ( .A(n7649), .B(n7648), .Z(n7755) );
  NANDN U8572 ( .A(n7651), .B(n7650), .Z(n7655) );
  NAND U8573 ( .A(n7653), .B(n7652), .Z(n7654) );
  AND U8574 ( .A(n7655), .B(n7654), .Z(n7756) );
  XNOR U8575 ( .A(n7755), .B(n7756), .Z(n7757) );
  NANDN U8576 ( .A(n7657), .B(n7656), .Z(n7661) );
  OR U8577 ( .A(n7659), .B(n7658), .Z(n7660) );
  AND U8578 ( .A(n7661), .B(n7660), .Z(n7964) );
  NANDN U8579 ( .A(n7663), .B(n7662), .Z(n7667) );
  OR U8580 ( .A(n7665), .B(n7664), .Z(n7666) );
  NAND U8581 ( .A(n7667), .B(n7666), .Z(n7892) );
  NANDN U8582 ( .A(n7669), .B(n7668), .Z(n7673) );
  OR U8583 ( .A(n7671), .B(n7670), .Z(n7672) );
  NAND U8584 ( .A(n7673), .B(n7672), .Z(n7891) );
  NAND U8585 ( .A(n33283), .B(n7674), .Z(n7676) );
  XOR U8586 ( .A(b[19]), .B(n19980), .Z(n7871) );
  OR U8587 ( .A(n7871), .B(n33021), .Z(n7675) );
  NAND U8588 ( .A(n7676), .B(n7675), .Z(n7948) );
  XOR U8589 ( .A(b[37]), .B(n14905), .Z(n7819) );
  NANDN U8590 ( .A(n7819), .B(n36311), .Z(n7679) );
  NANDN U8591 ( .A(n7677), .B(n36309), .Z(n7678) );
  NAND U8592 ( .A(n7679), .B(n7678), .Z(n7945) );
  XOR U8593 ( .A(b[43]), .B(n13106), .Z(n7813) );
  NANDN U8594 ( .A(n7813), .B(n37068), .Z(n7682) );
  NANDN U8595 ( .A(n7680), .B(n37069), .Z(n7681) );
  AND U8596 ( .A(n7682), .B(n7681), .Z(n7946) );
  XNOR U8597 ( .A(n7945), .B(n7946), .Z(n7947) );
  XNOR U8598 ( .A(n7948), .B(n7947), .Z(n7922) );
  XNOR U8599 ( .A(n981), .B(b[54]), .Z(n38075) );
  NAND U8600 ( .A(a[0]), .B(n38075), .Z(n7899) );
  NANDN U8601 ( .A(n966), .B(a[54]), .Z(n7683) );
  XOR U8602 ( .A(n29232), .B(n7683), .Z(n7685) );
  IV U8603 ( .A(a[53]), .Z(n25001) );
  NANDN U8604 ( .A(n25001), .B(n966), .Z(n7684) );
  AND U8605 ( .A(n7685), .B(n7684), .Z(n7897) );
  NAND U8606 ( .A(n37802), .B(n7686), .Z(n7688) );
  XOR U8607 ( .A(b[51]), .B(n10854), .Z(n7865) );
  NANDN U8608 ( .A(n7865), .B(n37803), .Z(n7687) );
  AND U8609 ( .A(n7688), .B(n7687), .Z(n7896) );
  XNOR U8610 ( .A(n7897), .B(n7896), .Z(n7898) );
  XOR U8611 ( .A(n7899), .B(n7898), .Z(n7921) );
  XNOR U8612 ( .A(n7922), .B(n7921), .Z(n7924) );
  NANDN U8613 ( .A(n7690), .B(n7689), .Z(n7694) );
  NAND U8614 ( .A(n7692), .B(n7691), .Z(n7693) );
  AND U8615 ( .A(n7694), .B(n7693), .Z(n7923) );
  XNOR U8616 ( .A(n7924), .B(n7923), .Z(n7770) );
  NANDN U8617 ( .A(n7696), .B(n7695), .Z(n7700) );
  NAND U8618 ( .A(n7698), .B(n7697), .Z(n7699) );
  NAND U8619 ( .A(n7700), .B(n7699), .Z(n7768) );
  XNOR U8620 ( .A(n7768), .B(n7767), .Z(n7769) );
  XOR U8621 ( .A(n7770), .B(n7769), .Z(n7890) );
  XNOR U8622 ( .A(n7891), .B(n7890), .Z(n7893) );
  XOR U8623 ( .A(n7892), .B(n7893), .Z(n7963) );
  OR U8624 ( .A(n7706), .B(n7705), .Z(n7710) );
  OR U8625 ( .A(n7708), .B(n7707), .Z(n7709) );
  NAND U8626 ( .A(n7710), .B(n7709), .Z(n7887) );
  NANDN U8627 ( .A(n7712), .B(n7711), .Z(n7716) );
  NAND U8628 ( .A(n7714), .B(n7713), .Z(n7715) );
  NAND U8629 ( .A(n7716), .B(n7715), .Z(n7884) );
  NAND U8630 ( .A(n7718), .B(n7717), .Z(n7722) );
  NANDN U8631 ( .A(n7720), .B(n7719), .Z(n7721) );
  AND U8632 ( .A(n7722), .B(n7721), .Z(n7885) );
  XNOR U8633 ( .A(n7884), .B(n7885), .Z(n7886) );
  XNOR U8634 ( .A(n7887), .B(n7886), .Z(n7965) );
  XNOR U8635 ( .A(n7966), .B(n7965), .Z(n7758) );
  XOR U8636 ( .A(n7757), .B(n7758), .Z(n7975) );
  XNOR U8637 ( .A(n7975), .B(n7976), .Z(n7977) );
  XOR U8638 ( .A(n7978), .B(n7977), .Z(n7987) );
  NANDN U8639 ( .A(n7728), .B(n7727), .Z(n7732) );
  NAND U8640 ( .A(n7730), .B(n7729), .Z(n7731) );
  NAND U8641 ( .A(n7732), .B(n7731), .Z(n7984) );
  NANDN U8642 ( .A(n7738), .B(n7737), .Z(n7742) );
  NAND U8643 ( .A(n7740), .B(n7739), .Z(n7741) );
  NAND U8644 ( .A(n7742), .B(n7741), .Z(n7982) );
  XNOR U8645 ( .A(n7981), .B(n7982), .Z(n7983) );
  XNOR U8646 ( .A(n7984), .B(n7983), .Z(n7988) );
  XOR U8647 ( .A(n7987), .B(n7988), .Z(n7989) );
  NANDN U8648 ( .A(n7744), .B(n7743), .Z(n7748) );
  NANDN U8649 ( .A(n7746), .B(n7745), .Z(n7747) );
  AND U8650 ( .A(n7748), .B(n7747), .Z(n7990) );
  XNOR U8651 ( .A(n7989), .B(n7990), .Z(n7750) );
  XNOR U8652 ( .A(n7749), .B(n7750), .Z(n7751) );
  XOR U8653 ( .A(n7752), .B(n7751), .Z(n7994) );
  XOR U8654 ( .A(n7995), .B(n7994), .Z(c[118]) );
  NANDN U8655 ( .A(n7750), .B(n7749), .Z(n7754) );
  NAND U8656 ( .A(n7752), .B(n7751), .Z(n7753) );
  NAND U8657 ( .A(n7754), .B(n7753), .Z(n8006) );
  NANDN U8658 ( .A(n7756), .B(n7755), .Z(n7760) );
  NANDN U8659 ( .A(n7758), .B(n7757), .Z(n7759) );
  NAND U8660 ( .A(n7760), .B(n7759), .Z(n8234) );
  NANDN U8661 ( .A(n7762), .B(n7761), .Z(n7766) );
  NAND U8662 ( .A(n7764), .B(n7763), .Z(n7765) );
  NAND U8663 ( .A(n7766), .B(n7765), .Z(n8109) );
  NANDN U8664 ( .A(n7768), .B(n7767), .Z(n7772) );
  NAND U8665 ( .A(n7770), .B(n7769), .Z(n7771) );
  NAND U8666 ( .A(n7772), .B(n7771), .Z(n8106) );
  NANDN U8667 ( .A(n7774), .B(n7773), .Z(n7778) );
  NAND U8668 ( .A(n7776), .B(n7775), .Z(n7777) );
  AND U8669 ( .A(n7778), .B(n7777), .Z(n8107) );
  XNOR U8670 ( .A(n8106), .B(n8107), .Z(n8108) );
  XOR U8671 ( .A(n8109), .B(n8108), .Z(n8222) );
  NANDN U8672 ( .A(n7784), .B(n7783), .Z(n7788) );
  NAND U8673 ( .A(n7786), .B(n7785), .Z(n7787) );
  NAND U8674 ( .A(n7788), .B(n7787), .Z(n8096) );
  XOR U8675 ( .A(b[9]), .B(n23149), .Z(n8028) );
  NANDN U8676 ( .A(n8028), .B(n30509), .Z(n7791) );
  NANDN U8677 ( .A(n7789), .B(n30846), .Z(n7790) );
  NAND U8678 ( .A(n7791), .B(n7790), .Z(n8058) );
  XOR U8679 ( .A(n31123), .B(n23852), .Z(n8158) );
  NAND U8680 ( .A(n8158), .B(n29949), .Z(n7794) );
  NAND U8681 ( .A(n29948), .B(n7792), .Z(n7793) );
  NAND U8682 ( .A(n7794), .B(n7793), .Z(n8055) );
  XNOR U8683 ( .A(b[35]), .B(a[21]), .Z(n8025) );
  NANDN U8684 ( .A(n8025), .B(n35985), .Z(n7797) );
  NANDN U8685 ( .A(n7795), .B(n35986), .Z(n7796) );
  AND U8686 ( .A(n7797), .B(n7796), .Z(n8056) );
  XNOR U8687 ( .A(n8055), .B(n8056), .Z(n8057) );
  XNOR U8688 ( .A(n8058), .B(n8057), .Z(n8094) );
  XOR U8689 ( .A(b[49]), .B(n11694), .Z(n8143) );
  OR U8690 ( .A(n8143), .B(n37756), .Z(n7800) );
  NANDN U8691 ( .A(n7798), .B(n37652), .Z(n7799) );
  NAND U8692 ( .A(n7800), .B(n7799), .Z(n8149) );
  XNOR U8693 ( .A(b[17]), .B(a[39]), .Z(n8067) );
  NANDN U8694 ( .A(n8067), .B(n32543), .Z(n7803) );
  NANDN U8695 ( .A(n7801), .B(n32541), .Z(n7802) );
  NAND U8696 ( .A(n7803), .B(n7802), .Z(n8146) );
  XOR U8697 ( .A(b[15]), .B(n21441), .Z(n8182) );
  OR U8698 ( .A(n8182), .B(n32010), .Z(n7806) );
  NANDN U8699 ( .A(n7804), .B(n32011), .Z(n7805) );
  AND U8700 ( .A(n7806), .B(n7805), .Z(n8147) );
  XNOR U8701 ( .A(n8146), .B(n8147), .Z(n8148) );
  XOR U8702 ( .A(n8149), .B(n8148), .Z(n8095) );
  XOR U8703 ( .A(n8094), .B(n8095), .Z(n8097) );
  XNOR U8704 ( .A(n8096), .B(n8097), .Z(n8215) );
  XNOR U8705 ( .A(b[21]), .B(a[35]), .Z(n8061) );
  OR U8706 ( .A(n8061), .B(n33634), .Z(n7809) );
  NANDN U8707 ( .A(n7807), .B(n33464), .Z(n7808) );
  NAND U8708 ( .A(n7809), .B(n7808), .Z(n8073) );
  XNOR U8709 ( .A(b[41]), .B(a[15]), .Z(n8161) );
  OR U8710 ( .A(n8161), .B(n36905), .Z(n7812) );
  NANDN U8711 ( .A(n7810), .B(n36807), .Z(n7811) );
  NAND U8712 ( .A(n7812), .B(n7811), .Z(n8070) );
  XOR U8713 ( .A(b[43]), .B(n13509), .Z(n8164) );
  NANDN U8714 ( .A(n8164), .B(n37068), .Z(n7815) );
  NANDN U8715 ( .A(n7813), .B(n37069), .Z(n7814) );
  AND U8716 ( .A(n7815), .B(n7814), .Z(n8071) );
  XNOR U8717 ( .A(n8070), .B(n8071), .Z(n8072) );
  XNOR U8718 ( .A(n8073), .B(n8072), .Z(n8022) );
  XOR U8719 ( .A(n973), .B(n16916), .Z(n8196) );
  NAND U8720 ( .A(n8196), .B(n35313), .Z(n7818) );
  NANDN U8721 ( .A(n7816), .B(n35311), .Z(n7817) );
  NAND U8722 ( .A(n7818), .B(n7817), .Z(n8179) );
  XOR U8723 ( .A(b[37]), .B(n15113), .Z(n8037) );
  NANDN U8724 ( .A(n8037), .B(n36311), .Z(n7821) );
  NANDN U8725 ( .A(n7819), .B(n36309), .Z(n7820) );
  NAND U8726 ( .A(n7821), .B(n7820), .Z(n8176) );
  NAND U8727 ( .A(n34044), .B(n7822), .Z(n7824) );
  XOR U8728 ( .A(n34510), .B(n19656), .Z(n8185) );
  NANDN U8729 ( .A(n33867), .B(n8185), .Z(n7823) );
  AND U8730 ( .A(n7824), .B(n7823), .Z(n8177) );
  XNOR U8731 ( .A(n8176), .B(n8177), .Z(n8178) );
  XNOR U8732 ( .A(n8179), .B(n8178), .Z(n8019) );
  XNOR U8733 ( .A(b[25]), .B(n18639), .Z(n8188) );
  NANDN U8734 ( .A(n34219), .B(n8188), .Z(n7827) );
  NANDN U8735 ( .A(n7825), .B(n34217), .Z(n7826) );
  NAND U8736 ( .A(n7827), .B(n7826), .Z(n8020) );
  XNOR U8737 ( .A(n8019), .B(n8020), .Z(n8021) );
  XOR U8738 ( .A(n8022), .B(n8021), .Z(n8085) );
  NANDN U8739 ( .A(n7829), .B(n7828), .Z(n7833) );
  NAND U8740 ( .A(n7831), .B(n7830), .Z(n7832) );
  NAND U8741 ( .A(n7833), .B(n7832), .Z(n8082) );
  NANDN U8742 ( .A(n7835), .B(n7834), .Z(n7839) );
  NAND U8743 ( .A(n7837), .B(n7836), .Z(n7838) );
  AND U8744 ( .A(n7839), .B(n7838), .Z(n8083) );
  XNOR U8745 ( .A(n8082), .B(n8083), .Z(n8084) );
  XNOR U8746 ( .A(n8085), .B(n8084), .Z(n8217) );
  XOR U8747 ( .A(n8218), .B(n8217), .Z(n8100) );
  NANDN U8748 ( .A(n7841), .B(n7840), .Z(n7845) );
  NAND U8749 ( .A(n7843), .B(n7842), .Z(n7844) );
  NAND U8750 ( .A(n7845), .B(n7844), .Z(n8101) );
  XOR U8751 ( .A(n8100), .B(n8101), .Z(n8102) );
  OR U8752 ( .A(n7847), .B(n7846), .Z(n7851) );
  OR U8753 ( .A(n7849), .B(n7848), .Z(n7850) );
  NAND U8754 ( .A(n7851), .B(n7850), .Z(n8210) );
  XOR U8755 ( .A(n8210), .B(n8209), .Z(n8211) );
  NANDN U8756 ( .A(n7857), .B(n7856), .Z(n7861) );
  NAND U8757 ( .A(n7859), .B(n7858), .Z(n7860) );
  NAND U8758 ( .A(n7861), .B(n7860), .Z(n8120) );
  XOR U8759 ( .A(n974), .B(n16269), .Z(n8137) );
  NAND U8760 ( .A(n35620), .B(n8137), .Z(n7864) );
  NANDN U8761 ( .A(n7862), .B(n35621), .Z(n7863) );
  NAND U8762 ( .A(n7864), .B(n7863), .Z(n8202) );
  XOR U8763 ( .A(b[51]), .B(n11202), .Z(n8134) );
  NANDN U8764 ( .A(n8134), .B(n37803), .Z(n7867) );
  NANDN U8765 ( .A(n7865), .B(n37802), .Z(n7866) );
  NAND U8766 ( .A(n7867), .B(n7866), .Z(n8199) );
  XOR U8767 ( .A(n968), .B(n24288), .Z(n8140) );
  NANDN U8768 ( .A(n29363), .B(n8140), .Z(n7870) );
  NANDN U8769 ( .A(n7868), .B(n29864), .Z(n7869) );
  AND U8770 ( .A(n7870), .B(n7869), .Z(n8200) );
  XNOR U8771 ( .A(n8199), .B(n8200), .Z(n8201) );
  XNOR U8772 ( .A(n8202), .B(n8201), .Z(n8118) );
  NANDN U8773 ( .A(n7871), .B(n33283), .Z(n7873) );
  XNOR U8774 ( .A(n33020), .B(a[37]), .Z(n8064) );
  NANDN U8775 ( .A(n33021), .B(n8064), .Z(n7872) );
  NAND U8776 ( .A(n7873), .B(n7872), .Z(n8045) );
  NAND U8777 ( .A(n37262), .B(n7874), .Z(n7876) );
  XNOR U8778 ( .A(b[45]), .B(a[11]), .Z(n8031) );
  NANDN U8779 ( .A(n8031), .B(n37261), .Z(n7875) );
  AND U8780 ( .A(n7876), .B(n7875), .Z(n8044) );
  NANDN U8781 ( .A(n7877), .B(n37469), .Z(n7879) );
  XNOR U8782 ( .A(n978), .B(a[9]), .Z(n8155) );
  NAND U8783 ( .A(n8155), .B(n37471), .Z(n7878) );
  NAND U8784 ( .A(n7879), .B(n7878), .Z(n8043) );
  XNOR U8785 ( .A(n8044), .B(n8043), .Z(n8046) );
  XOR U8786 ( .A(n8045), .B(n8046), .Z(n8119) );
  XOR U8787 ( .A(n8118), .B(n8119), .Z(n8121) );
  XOR U8788 ( .A(n8120), .B(n8121), .Z(n8212) );
  XOR U8789 ( .A(n8211), .B(n8212), .Z(n8103) );
  XNOR U8790 ( .A(n8102), .B(n8103), .Z(n8221) );
  XOR U8791 ( .A(n8222), .B(n8221), .Z(n8224) );
  XNOR U8792 ( .A(n8224), .B(n8223), .Z(n8230) );
  NANDN U8793 ( .A(n7885), .B(n7884), .Z(n7889) );
  NAND U8794 ( .A(n7887), .B(n7886), .Z(n7888) );
  NAND U8795 ( .A(n7889), .B(n7888), .Z(n8227) );
  NAND U8796 ( .A(n7891), .B(n7890), .Z(n7895) );
  NANDN U8797 ( .A(n7893), .B(n7892), .Z(n7894) );
  AND U8798 ( .A(n7895), .B(n7894), .Z(n8228) );
  XNOR U8799 ( .A(n8227), .B(n8228), .Z(n8229) );
  XOR U8800 ( .A(n8230), .B(n8229), .Z(n8233) );
  XNOR U8801 ( .A(n8234), .B(n8233), .Z(n8235) );
  NANDN U8802 ( .A(n7897), .B(n7896), .Z(n7901) );
  NAND U8803 ( .A(n7899), .B(n7898), .Z(n7900) );
  NAND U8804 ( .A(n7901), .B(n7900), .Z(n8088) );
  NANDN U8805 ( .A(n7903), .B(n7902), .Z(n7907) );
  NAND U8806 ( .A(n7905), .B(n7904), .Z(n7906) );
  NAND U8807 ( .A(n7907), .B(n7906), .Z(n8089) );
  XNOR U8808 ( .A(n8088), .B(n8089), .Z(n8090) );
  XOR U8809 ( .A(n981), .B(n10524), .Z(n8079) );
  NAND U8810 ( .A(n8079), .B(n37940), .Z(n7910) );
  NANDN U8811 ( .A(n7908), .B(n37941), .Z(n7909) );
  NAND U8812 ( .A(n7910), .B(n7909), .Z(n8192) );
  XNOR U8813 ( .A(n982), .B(a[0]), .Z(n7913) );
  XNOR U8814 ( .A(n982), .B(b[53]), .Z(n7912) );
  XNOR U8815 ( .A(n982), .B(b[54]), .Z(n7911) );
  AND U8816 ( .A(n7912), .B(n7911), .Z(n38073) );
  NAND U8817 ( .A(n7913), .B(n38073), .Z(n7915) );
  XOR U8818 ( .A(n982), .B(n10457), .Z(n8193) );
  NAND U8819 ( .A(n38075), .B(n8193), .Z(n7914) );
  NAND U8820 ( .A(n7915), .B(n7914), .Z(n8191) );
  XNOR U8821 ( .A(n8192), .B(n8191), .Z(n8052) );
  NOR U8822 ( .A(b[53]), .B(b[54]), .Z(n7916) );
  OR U8823 ( .A(n7916), .B(n986), .Z(n7917) );
  NANDN U8824 ( .A(n981), .B(b[54]), .Z(n38138) );
  AND U8825 ( .A(n38138), .B(b[55]), .Z(n38236) );
  IV U8826 ( .A(n38236), .Z(n38192) );
  ANDN U8827 ( .B(n7917), .A(n38192), .Z(n8050) );
  NANDN U8828 ( .A(n7918), .B(n35188), .Z(n7920) );
  XNOR U8829 ( .A(n35540), .B(a[27]), .Z(n8128) );
  NANDN U8830 ( .A(n34968), .B(n8128), .Z(n7919) );
  NAND U8831 ( .A(n7920), .B(n7919), .Z(n8049) );
  XOR U8832 ( .A(n8050), .B(n8049), .Z(n8051) );
  XOR U8833 ( .A(n8052), .B(n8051), .Z(n8091) );
  XOR U8834 ( .A(n8090), .B(n8091), .Z(n8016) );
  OR U8835 ( .A(n7922), .B(n7921), .Z(n7926) );
  OR U8836 ( .A(n7924), .B(n7923), .Z(n7925) );
  AND U8837 ( .A(n7926), .B(n7925), .Z(n8013) );
  XOR U8838 ( .A(b[39]), .B(n14514), .Z(n8040) );
  NANDN U8839 ( .A(n8040), .B(n36553), .Z(n7929) );
  NAND U8840 ( .A(n7927), .B(n36643), .Z(n7928) );
  NAND U8841 ( .A(n7929), .B(n7928), .Z(n8173) );
  XOR U8842 ( .A(b[13]), .B(n21996), .Z(n8034) );
  OR U8843 ( .A(n8034), .B(n31550), .Z(n7932) );
  NAND U8844 ( .A(n7930), .B(n31874), .Z(n7931) );
  NAND U8845 ( .A(n7932), .B(n7931), .Z(n8170) );
  XOR U8846 ( .A(b[11]), .B(n22579), .Z(n8167) );
  OR U8847 ( .A(n8167), .B(n31369), .Z(n7935) );
  NANDN U8848 ( .A(n7933), .B(n31119), .Z(n7934) );
  AND U8849 ( .A(n7935), .B(n7934), .Z(n8171) );
  XNOR U8850 ( .A(n8170), .B(n8171), .Z(n8172) );
  XNOR U8851 ( .A(n8173), .B(n8172), .Z(n8127) );
  XOR U8852 ( .A(n967), .B(n25001), .Z(n8131) );
  NAND U8853 ( .A(n8131), .B(n28939), .Z(n7938) );
  NAND U8854 ( .A(n28938), .B(n7936), .Z(n7937) );
  NAND U8855 ( .A(n7938), .B(n7937), .Z(n8208) );
  NANDN U8856 ( .A(n966), .B(a[55]), .Z(n7939) );
  XOR U8857 ( .A(n29232), .B(n7939), .Z(n7941) );
  IV U8858 ( .A(a[54]), .Z(n25177) );
  NANDN U8859 ( .A(n25177), .B(n966), .Z(n7940) );
  AND U8860 ( .A(n7941), .B(n7940), .Z(n8205) );
  NAND U8861 ( .A(n7942), .B(n34848), .Z(n7944) );
  XOR U8862 ( .A(n35375), .B(n18003), .Z(n8152) );
  NAND U8863 ( .A(n34618), .B(n8152), .Z(n7943) );
  AND U8864 ( .A(n7944), .B(n7943), .Z(n8206) );
  XNOR U8865 ( .A(n8205), .B(n8206), .Z(n8207) );
  XNOR U8866 ( .A(n8208), .B(n8207), .Z(n8124) );
  NANDN U8867 ( .A(n7946), .B(n7945), .Z(n7950) );
  NAND U8868 ( .A(n7948), .B(n7947), .Z(n7949) );
  NAND U8869 ( .A(n7950), .B(n7949), .Z(n8125) );
  XNOR U8870 ( .A(n8124), .B(n8125), .Z(n8126) );
  XOR U8871 ( .A(n8127), .B(n8126), .Z(n8014) );
  XNOR U8872 ( .A(n8013), .B(n8014), .Z(n8015) );
  XOR U8873 ( .A(n8016), .B(n8015), .Z(n8115) );
  NANDN U8874 ( .A(n7952), .B(n7951), .Z(n7956) );
  NANDN U8875 ( .A(n7954), .B(n7953), .Z(n7955) );
  NAND U8876 ( .A(n7956), .B(n7955), .Z(n8112) );
  NANDN U8877 ( .A(n7958), .B(n7957), .Z(n7962) );
  NAND U8878 ( .A(n7960), .B(n7959), .Z(n7961) );
  AND U8879 ( .A(n7962), .B(n7961), .Z(n8113) );
  XNOR U8880 ( .A(n8112), .B(n8113), .Z(n8114) );
  XOR U8881 ( .A(n8115), .B(n8114), .Z(n8242) );
  OR U8882 ( .A(n7964), .B(n7963), .Z(n7968) );
  OR U8883 ( .A(n7966), .B(n7965), .Z(n7967) );
  AND U8884 ( .A(n7968), .B(n7967), .Z(n8240) );
  NAND U8885 ( .A(n7970), .B(n7969), .Z(n7974) );
  NAND U8886 ( .A(n7972), .B(n7971), .Z(n7973) );
  AND U8887 ( .A(n7974), .B(n7973), .Z(n8239) );
  XNOR U8888 ( .A(n8240), .B(n8239), .Z(n8241) );
  XNOR U8889 ( .A(n8242), .B(n8241), .Z(n8236) );
  XNOR U8890 ( .A(n8235), .B(n8236), .Z(n8010) );
  NANDN U8891 ( .A(n7976), .B(n7975), .Z(n7980) );
  NAND U8892 ( .A(n7978), .B(n7977), .Z(n7979) );
  NAND U8893 ( .A(n7980), .B(n7979), .Z(n8007) );
  NANDN U8894 ( .A(n7982), .B(n7981), .Z(n7986) );
  NAND U8895 ( .A(n7984), .B(n7983), .Z(n7985) );
  NAND U8896 ( .A(n7986), .B(n7985), .Z(n8008) );
  XNOR U8897 ( .A(n8007), .B(n8008), .Z(n8009) );
  XNOR U8898 ( .A(n8010), .B(n8009), .Z(n8003) );
  OR U8899 ( .A(n7988), .B(n7987), .Z(n7992) );
  NAND U8900 ( .A(n7990), .B(n7989), .Z(n7991) );
  AND U8901 ( .A(n7992), .B(n7991), .Z(n8004) );
  XNOR U8902 ( .A(n8003), .B(n8004), .Z(n8005) );
  XNOR U8903 ( .A(n8006), .B(n8005), .Z(n7998) );
  XNOR U8904 ( .A(n7998), .B(sreg[119]), .Z(n8000) );
  NAND U8905 ( .A(n7993), .B(sreg[118]), .Z(n7997) );
  OR U8906 ( .A(n7995), .B(n7994), .Z(n7996) );
  AND U8907 ( .A(n7997), .B(n7996), .Z(n7999) );
  XOR U8908 ( .A(n8000), .B(n7999), .Z(c[119]) );
  NAND U8909 ( .A(n7998), .B(sreg[119]), .Z(n8002) );
  OR U8910 ( .A(n8000), .B(n7999), .Z(n8001) );
  NAND U8911 ( .A(n8002), .B(n8001), .Z(n8497) );
  XNOR U8912 ( .A(n8497), .B(sreg[120]), .Z(n8499) );
  NANDN U8913 ( .A(n8008), .B(n8007), .Z(n8012) );
  NAND U8914 ( .A(n8010), .B(n8009), .Z(n8011) );
  NAND U8915 ( .A(n8012), .B(n8011), .Z(n8245) );
  OR U8916 ( .A(n8014), .B(n8013), .Z(n8018) );
  OR U8917 ( .A(n8016), .B(n8015), .Z(n8017) );
  NAND U8918 ( .A(n8018), .B(n8017), .Z(n8270) );
  NANDN U8919 ( .A(n8020), .B(n8019), .Z(n8024) );
  NAND U8920 ( .A(n8022), .B(n8021), .Z(n8023) );
  NAND U8921 ( .A(n8024), .B(n8023), .Z(n8410) );
  XNOR U8922 ( .A(b[35]), .B(a[22]), .Z(n8374) );
  NANDN U8923 ( .A(n8374), .B(n35985), .Z(n8027) );
  NANDN U8924 ( .A(n8025), .B(n35986), .Z(n8026) );
  NAND U8925 ( .A(n8027), .B(n8026), .Z(n8329) );
  XOR U8926 ( .A(b[9]), .B(n23447), .Z(n8377) );
  NANDN U8927 ( .A(n8377), .B(n30509), .Z(n8030) );
  NANDN U8928 ( .A(n8028), .B(n30846), .Z(n8029) );
  NAND U8929 ( .A(n8030), .B(n8029), .Z(n8326) );
  XNOR U8930 ( .A(b[45]), .B(a[12]), .Z(n8341) );
  NANDN U8931 ( .A(n8341), .B(n37261), .Z(n8033) );
  NANDN U8932 ( .A(n8031), .B(n37262), .Z(n8032) );
  AND U8933 ( .A(n8033), .B(n8032), .Z(n8327) );
  XNOR U8934 ( .A(n8326), .B(n8327), .Z(n8328) );
  XOR U8935 ( .A(n8329), .B(n8328), .Z(n8394) );
  XOR U8936 ( .A(b[13]), .B(n22289), .Z(n8452) );
  OR U8937 ( .A(n8452), .B(n31550), .Z(n8036) );
  NANDN U8938 ( .A(n8034), .B(n31874), .Z(n8035) );
  NAND U8939 ( .A(n8036), .B(n8035), .Z(n8371) );
  XOR U8940 ( .A(b[37]), .B(n15484), .Z(n8302) );
  NANDN U8941 ( .A(n8302), .B(n36311), .Z(n8039) );
  NANDN U8942 ( .A(n8037), .B(n36309), .Z(n8038) );
  NAND U8943 ( .A(n8039), .B(n8038), .Z(n8368) );
  XOR U8944 ( .A(b[39]), .B(n14905), .Z(n8449) );
  NANDN U8945 ( .A(n8449), .B(n36553), .Z(n8042) );
  NANDN U8946 ( .A(n8040), .B(n36643), .Z(n8041) );
  AND U8947 ( .A(n8042), .B(n8041), .Z(n8369) );
  XNOR U8948 ( .A(n8368), .B(n8369), .Z(n8370) );
  XOR U8949 ( .A(n8371), .B(n8370), .Z(n8392) );
  NANDN U8950 ( .A(n8044), .B(n8043), .Z(n8048) );
  NAND U8951 ( .A(n8046), .B(n8045), .Z(n8047) );
  NAND U8952 ( .A(n8048), .B(n8047), .Z(n8393) );
  XNOR U8953 ( .A(n8392), .B(n8393), .Z(n8395) );
  XNOR U8954 ( .A(n8394), .B(n8395), .Z(n8411) );
  XNOR U8955 ( .A(n8410), .B(n8411), .Z(n8412) );
  OR U8956 ( .A(n8050), .B(n8049), .Z(n8054) );
  NAND U8957 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U8958 ( .A(n8054), .B(n8053), .Z(n8422) );
  NANDN U8959 ( .A(n8056), .B(n8055), .Z(n8060) );
  NAND U8960 ( .A(n8058), .B(n8057), .Z(n8059) );
  NAND U8961 ( .A(n8060), .B(n8059), .Z(n8423) );
  XNOR U8962 ( .A(n8422), .B(n8423), .Z(n8424) );
  XNOR U8963 ( .A(b[21]), .B(a[36]), .Z(n8467) );
  OR U8964 ( .A(n8467), .B(n33634), .Z(n8063) );
  NANDN U8965 ( .A(n8061), .B(n33464), .Z(n8062) );
  NAND U8966 ( .A(n8063), .B(n8062), .Z(n8476) );
  NAND U8967 ( .A(n8064), .B(n33283), .Z(n8066) );
  XOR U8968 ( .A(n33020), .B(n20686), .Z(n8461) );
  NANDN U8969 ( .A(n33021), .B(n8461), .Z(n8065) );
  NAND U8970 ( .A(n8066), .B(n8065), .Z(n8473) );
  XNOR U8971 ( .A(b[17]), .B(a[40]), .Z(n8299) );
  NANDN U8972 ( .A(n8299), .B(n32543), .Z(n8069) );
  NANDN U8973 ( .A(n8067), .B(n32541), .Z(n8068) );
  AND U8974 ( .A(n8069), .B(n8068), .Z(n8474) );
  XNOR U8975 ( .A(n8473), .B(n8474), .Z(n8475) );
  XOR U8976 ( .A(n8476), .B(n8475), .Z(n8428) );
  NANDN U8977 ( .A(n8071), .B(n8070), .Z(n8075) );
  NAND U8978 ( .A(n8073), .B(n8072), .Z(n8074) );
  NAND U8979 ( .A(n8075), .B(n8074), .Z(n8429) );
  XNOR U8980 ( .A(n8428), .B(n8429), .Z(n8431) );
  NAND U8981 ( .A(a[0]), .B(n964), .Z(n8437) );
  NANDN U8982 ( .A(n966), .B(a[56]), .Z(n8076) );
  XOR U8983 ( .A(n29232), .B(n8076), .Z(n8078) );
  IV U8984 ( .A(a[55]), .Z(n25466) );
  NANDN U8985 ( .A(n25466), .B(n966), .Z(n8077) );
  AND U8986 ( .A(n8078), .B(n8077), .Z(n8435) );
  NAND U8987 ( .A(n37941), .B(n8079), .Z(n8081) );
  XOR U8988 ( .A(b[53]), .B(n10854), .Z(n8350) );
  NANDN U8989 ( .A(n8350), .B(n37940), .Z(n8080) );
  AND U8990 ( .A(n8081), .B(n8080), .Z(n8434) );
  XNOR U8991 ( .A(n8435), .B(n8434), .Z(n8436) );
  XNOR U8992 ( .A(n8437), .B(n8436), .Z(n8430) );
  XNOR U8993 ( .A(n8431), .B(n8430), .Z(n8425) );
  XOR U8994 ( .A(n8424), .B(n8425), .Z(n8413) );
  XNOR U8995 ( .A(n8412), .B(n8413), .Z(n8269) );
  XNOR U8996 ( .A(n8270), .B(n8269), .Z(n8271) );
  NANDN U8997 ( .A(n8083), .B(n8082), .Z(n8087) );
  NANDN U8998 ( .A(n8085), .B(n8084), .Z(n8086) );
  NAND U8999 ( .A(n8087), .B(n8086), .Z(n8488) );
  NANDN U9000 ( .A(n8089), .B(n8088), .Z(n8093) );
  NAND U9001 ( .A(n8091), .B(n8090), .Z(n8092) );
  NAND U9002 ( .A(n8093), .B(n8092), .Z(n8485) );
  NANDN U9003 ( .A(n8095), .B(n8094), .Z(n8099) );
  OR U9004 ( .A(n8097), .B(n8096), .Z(n8098) );
  AND U9005 ( .A(n8099), .B(n8098), .Z(n8486) );
  XNOR U9006 ( .A(n8485), .B(n8486), .Z(n8487) );
  XOR U9007 ( .A(n8488), .B(n8487), .Z(n8272) );
  XNOR U9008 ( .A(n8271), .B(n8272), .Z(n8259) );
  OR U9009 ( .A(n8101), .B(n8100), .Z(n8105) );
  NANDN U9010 ( .A(n8103), .B(n8102), .Z(n8104) );
  NAND U9011 ( .A(n8105), .B(n8104), .Z(n8491) );
  NANDN U9012 ( .A(n8107), .B(n8106), .Z(n8111) );
  NAND U9013 ( .A(n8109), .B(n8108), .Z(n8110) );
  NAND U9014 ( .A(n8111), .B(n8110), .Z(n8492) );
  XNOR U9015 ( .A(n8491), .B(n8492), .Z(n8493) );
  NANDN U9016 ( .A(n8113), .B(n8112), .Z(n8117) );
  NANDN U9017 ( .A(n8115), .B(n8114), .Z(n8116) );
  AND U9018 ( .A(n8117), .B(n8116), .Z(n8494) );
  XOR U9019 ( .A(n8493), .B(n8494), .Z(n8257) );
  NANDN U9020 ( .A(n8119), .B(n8118), .Z(n8123) );
  OR U9021 ( .A(n8121), .B(n8120), .Z(n8122) );
  NAND U9022 ( .A(n8123), .B(n8122), .Z(n8479) );
  XNOR U9023 ( .A(n8479), .B(n8480), .Z(n8481) );
  NAND U9024 ( .A(n8128), .B(n35188), .Z(n8130) );
  XOR U9025 ( .A(n35540), .B(n17702), .Z(n8347) );
  NANDN U9026 ( .A(n34968), .B(n8347), .Z(n8129) );
  NAND U9027 ( .A(n8130), .B(n8129), .Z(n8317) );
  XOR U9028 ( .A(b[3]), .B(n25177), .Z(n8386) );
  NANDN U9029 ( .A(n8386), .B(n28939), .Z(n8133) );
  NAND U9030 ( .A(n28938), .B(n8131), .Z(n8132) );
  NAND U9031 ( .A(n8133), .B(n8132), .Z(n8314) );
  XOR U9032 ( .A(b[51]), .B(n11406), .Z(n8446) );
  NANDN U9033 ( .A(n8446), .B(n37803), .Z(n8136) );
  NANDN U9034 ( .A(n8134), .B(n37802), .Z(n8135) );
  AND U9035 ( .A(n8136), .B(n8135), .Z(n8315) );
  XNOR U9036 ( .A(n8314), .B(n8315), .Z(n8316) );
  XNOR U9037 ( .A(n8317), .B(n8316), .Z(n8401) );
  XOR U9038 ( .A(b[33]), .B(n16508), .Z(n8389) );
  NANDN U9039 ( .A(n8389), .B(n35620), .Z(n8139) );
  NAND U9040 ( .A(n8137), .B(n35621), .Z(n8138) );
  NAND U9041 ( .A(n8139), .B(n8138), .Z(n8364) );
  XOR U9042 ( .A(b[5]), .B(n25134), .Z(n8353) );
  OR U9043 ( .A(n8353), .B(n29363), .Z(n8142) );
  NAND U9044 ( .A(n8140), .B(n29864), .Z(n8141) );
  AND U9045 ( .A(n8142), .B(n8141), .Z(n8362) );
  XOR U9046 ( .A(b[49]), .B(n11986), .Z(n8443) );
  OR U9047 ( .A(n8443), .B(n37756), .Z(n8145) );
  NANDN U9048 ( .A(n8143), .B(n37652), .Z(n8144) );
  AND U9049 ( .A(n8145), .B(n8144), .Z(n8363) );
  XOR U9050 ( .A(n8364), .B(n8365), .Z(n8398) );
  NANDN U9051 ( .A(n8147), .B(n8146), .Z(n8151) );
  NAND U9052 ( .A(n8149), .B(n8148), .Z(n8150) );
  NAND U9053 ( .A(n8151), .B(n8150), .Z(n8399) );
  XNOR U9054 ( .A(n8398), .B(n8399), .Z(n8400) );
  XOR U9055 ( .A(n8401), .B(n8400), .Z(n8417) );
  NAND U9056 ( .A(n34848), .B(n8152), .Z(n8154) );
  XOR U9057 ( .A(n35375), .B(n18804), .Z(n8464) );
  NAND U9058 ( .A(n34618), .B(n8464), .Z(n8153) );
  NAND U9059 ( .A(n8154), .B(n8153), .Z(n8311) );
  NAND U9060 ( .A(n8155), .B(n37469), .Z(n8157) );
  XOR U9061 ( .A(n978), .B(n12555), .Z(n8344) );
  NAND U9062 ( .A(n8344), .B(n37471), .Z(n8156) );
  NAND U9063 ( .A(n8157), .B(n8156), .Z(n8308) );
  XOR U9064 ( .A(n31123), .B(n24671), .Z(n8380) );
  NAND U9065 ( .A(n8380), .B(n29949), .Z(n8160) );
  NAND U9066 ( .A(n29948), .B(n8158), .Z(n8159) );
  AND U9067 ( .A(n8160), .B(n8159), .Z(n8309) );
  XNOR U9068 ( .A(n8308), .B(n8309), .Z(n8310) );
  XNOR U9069 ( .A(n8311), .B(n8310), .Z(n8409) );
  XNOR U9070 ( .A(b[41]), .B(a[16]), .Z(n8305) );
  OR U9071 ( .A(n8305), .B(n36905), .Z(n8163) );
  NANDN U9072 ( .A(n8161), .B(n36807), .Z(n8162) );
  NAND U9073 ( .A(n8163), .B(n8162), .Z(n8282) );
  XOR U9074 ( .A(b[43]), .B(n14210), .Z(n8440) );
  NANDN U9075 ( .A(n8440), .B(n37068), .Z(n8166) );
  NANDN U9076 ( .A(n8164), .B(n37069), .Z(n8165) );
  NAND U9077 ( .A(n8166), .B(n8165), .Z(n8279) );
  XOR U9078 ( .A(b[11]), .B(n22964), .Z(n8455) );
  OR U9079 ( .A(n8455), .B(n31369), .Z(n8169) );
  NANDN U9080 ( .A(n8167), .B(n31119), .Z(n8168) );
  AND U9081 ( .A(n8169), .B(n8168), .Z(n8280) );
  XNOR U9082 ( .A(n8279), .B(n8280), .Z(n8281) );
  XNOR U9083 ( .A(n8282), .B(n8281), .Z(n8406) );
  NANDN U9084 ( .A(n8171), .B(n8170), .Z(n8175) );
  NAND U9085 ( .A(n8173), .B(n8172), .Z(n8174) );
  NAND U9086 ( .A(n8175), .B(n8174), .Z(n8407) );
  XNOR U9087 ( .A(n8406), .B(n8407), .Z(n8408) );
  XOR U9088 ( .A(n8409), .B(n8408), .Z(n8416) );
  XNOR U9089 ( .A(n8417), .B(n8416), .Z(n8419) );
  NANDN U9090 ( .A(n8177), .B(n8176), .Z(n8181) );
  NAND U9091 ( .A(n8179), .B(n8178), .Z(n8180) );
  NAND U9092 ( .A(n8181), .B(n8180), .Z(n8323) );
  XOR U9093 ( .A(b[15]), .B(n22246), .Z(n8338) );
  OR U9094 ( .A(n8338), .B(n32010), .Z(n8184) );
  NANDN U9095 ( .A(n8182), .B(n32011), .Z(n8183) );
  NAND U9096 ( .A(n8184), .B(n8183), .Z(n8359) );
  NAND U9097 ( .A(n34044), .B(n8185), .Z(n8187) );
  XOR U9098 ( .A(n34510), .B(n19513), .Z(n8458) );
  NANDN U9099 ( .A(n33867), .B(n8458), .Z(n8186) );
  NAND U9100 ( .A(n8187), .B(n8186), .Z(n8356) );
  XNOR U9101 ( .A(b[25]), .B(a[32]), .Z(n8470) );
  OR U9102 ( .A(n8470), .B(n34219), .Z(n8190) );
  NAND U9103 ( .A(n8188), .B(n34217), .Z(n8189) );
  AND U9104 ( .A(n8190), .B(n8189), .Z(n8357) );
  XNOR U9105 ( .A(n8356), .B(n8357), .Z(n8358) );
  XNOR U9106 ( .A(n8359), .B(n8358), .Z(n8320) );
  AND U9107 ( .A(n8192), .B(n8191), .Z(n8335) );
  XNOR U9108 ( .A(n982), .B(a[2]), .Z(n8285) );
  NAND U9109 ( .A(n38075), .B(n8285), .Z(n8195) );
  NAND U9110 ( .A(n8193), .B(n38073), .Z(n8194) );
  NAND U9111 ( .A(n8195), .B(n8194), .Z(n8333) );
  NAND U9112 ( .A(n8196), .B(n35311), .Z(n8198) );
  XOR U9113 ( .A(b[31]), .B(n17133), .Z(n8296) );
  NANDN U9114 ( .A(n8296), .B(n35313), .Z(n8197) );
  NAND U9115 ( .A(n8198), .B(n8197), .Z(n8332) );
  XOR U9116 ( .A(n8335), .B(n8334), .Z(n8321) );
  XNOR U9117 ( .A(n8320), .B(n8321), .Z(n8322) );
  XNOR U9118 ( .A(n8323), .B(n8322), .Z(n8404) );
  NANDN U9119 ( .A(n8200), .B(n8199), .Z(n8204) );
  NAND U9120 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U9121 ( .A(n8204), .B(n8203), .Z(n8403) );
  XNOR U9122 ( .A(n8403), .B(n8402), .Z(n8405) );
  XOR U9123 ( .A(n8404), .B(n8405), .Z(n8418) );
  XNOR U9124 ( .A(n8419), .B(n8418), .Z(n8482) );
  XNOR U9125 ( .A(n8481), .B(n8482), .Z(n8276) );
  OR U9126 ( .A(n8210), .B(n8209), .Z(n8214) );
  NANDN U9127 ( .A(n8212), .B(n8211), .Z(n8213) );
  NAND U9128 ( .A(n8214), .B(n8213), .Z(n8273) );
  OR U9129 ( .A(n8216), .B(n8215), .Z(n8220) );
  OR U9130 ( .A(n8218), .B(n8217), .Z(n8219) );
  NAND U9131 ( .A(n8220), .B(n8219), .Z(n8274) );
  XNOR U9132 ( .A(n8273), .B(n8274), .Z(n8275) );
  XOR U9133 ( .A(n8276), .B(n8275), .Z(n8258) );
  XNOR U9134 ( .A(n8257), .B(n8258), .Z(n8260) );
  XNOR U9135 ( .A(n8259), .B(n8260), .Z(n8266) );
  NANDN U9136 ( .A(n8222), .B(n8221), .Z(n8226) );
  OR U9137 ( .A(n8224), .B(n8223), .Z(n8225) );
  NAND U9138 ( .A(n8226), .B(n8225), .Z(n8263) );
  NANDN U9139 ( .A(n8228), .B(n8227), .Z(n8232) );
  NAND U9140 ( .A(n8230), .B(n8229), .Z(n8231) );
  NAND U9141 ( .A(n8232), .B(n8231), .Z(n8264) );
  XNOR U9142 ( .A(n8263), .B(n8264), .Z(n8265) );
  XNOR U9143 ( .A(n8266), .B(n8265), .Z(n8254) );
  NAND U9144 ( .A(n8234), .B(n8233), .Z(n8238) );
  OR U9145 ( .A(n8236), .B(n8235), .Z(n8237) );
  NAND U9146 ( .A(n8238), .B(n8237), .Z(n8251) );
  OR U9147 ( .A(n8240), .B(n8239), .Z(n8244) );
  OR U9148 ( .A(n8242), .B(n8241), .Z(n8243) );
  AND U9149 ( .A(n8244), .B(n8243), .Z(n8252) );
  XNOR U9150 ( .A(n8251), .B(n8252), .Z(n8253) );
  XOR U9151 ( .A(n8254), .B(n8253), .Z(n8246) );
  XOR U9152 ( .A(n8245), .B(n8246), .Z(n8247) );
  XOR U9153 ( .A(n8248), .B(n8247), .Z(n8498) );
  XOR U9154 ( .A(n8499), .B(n8498), .Z(c[120]) );
  OR U9155 ( .A(n8246), .B(n8245), .Z(n8250) );
  NAND U9156 ( .A(n8248), .B(n8247), .Z(n8249) );
  NAND U9157 ( .A(n8250), .B(n8249), .Z(n8510) );
  NANDN U9158 ( .A(n8252), .B(n8251), .Z(n8256) );
  NANDN U9159 ( .A(n8254), .B(n8253), .Z(n8255) );
  NAND U9160 ( .A(n8256), .B(n8255), .Z(n8508) );
  OR U9161 ( .A(n8258), .B(n8257), .Z(n8262) );
  NANDN U9162 ( .A(n8260), .B(n8259), .Z(n8261) );
  NAND U9163 ( .A(n8262), .B(n8261), .Z(n8513) );
  NANDN U9164 ( .A(n8264), .B(n8263), .Z(n8268) );
  NANDN U9165 ( .A(n8266), .B(n8265), .Z(n8267) );
  NAND U9166 ( .A(n8268), .B(n8267), .Z(n8514) );
  XNOR U9167 ( .A(n8513), .B(n8514), .Z(n8515) );
  NANDN U9168 ( .A(n8274), .B(n8273), .Z(n8278) );
  NAND U9169 ( .A(n8276), .B(n8275), .Z(n8277) );
  AND U9170 ( .A(n8278), .B(n8277), .Z(n8758) );
  XOR U9171 ( .A(n8759), .B(n8758), .Z(n8760) );
  NANDN U9172 ( .A(n8280), .B(n8279), .Z(n8284) );
  NAND U9173 ( .A(n8282), .B(n8281), .Z(n8283) );
  NAND U9174 ( .A(n8284), .B(n8283), .Z(n8698) );
  XOR U9175 ( .A(n982), .B(n10524), .Z(n8624) );
  NAND U9176 ( .A(n38075), .B(n8624), .Z(n8287) );
  NAND U9177 ( .A(n8285), .B(n38073), .Z(n8286) );
  NAND U9178 ( .A(n8287), .B(n8286), .Z(n8628) );
  XNOR U9179 ( .A(n983), .B(a[0]), .Z(n8290) );
  XNOR U9180 ( .A(n983), .B(b[55]), .Z(n8559) );
  IV U9181 ( .A(b[56]), .Z(n8383) );
  XOR U9182 ( .A(n983), .B(n8383), .Z(n8288) );
  AND U9183 ( .A(n8559), .B(n8288), .Z(n8289) );
  NAND U9184 ( .A(n8290), .B(n8289), .Z(n8292) );
  XOR U9185 ( .A(n983), .B(n10457), .Z(n8560) );
  NANDN U9186 ( .A(n965), .B(n8560), .Z(n8291) );
  NAND U9187 ( .A(n8292), .B(n8291), .Z(n8627) );
  XNOR U9188 ( .A(n8628), .B(n8627), .Z(n8644) );
  NANDN U9189 ( .A(n966), .B(a[57]), .Z(n8293) );
  XOR U9190 ( .A(n29232), .B(n8293), .Z(n8295) );
  IV U9191 ( .A(a[56]), .Z(n25860) );
  NANDN U9192 ( .A(n25860), .B(n966), .Z(n8294) );
  AND U9193 ( .A(n8295), .B(n8294), .Z(n8642) );
  NANDN U9194 ( .A(n8296), .B(n35311), .Z(n8298) );
  XOR U9195 ( .A(b[31]), .B(n17960), .Z(n8629) );
  NANDN U9196 ( .A(n8629), .B(n35313), .Z(n8297) );
  AND U9197 ( .A(n8298), .B(n8297), .Z(n8641) );
  XNOR U9198 ( .A(n8642), .B(n8641), .Z(n8643) );
  XOR U9199 ( .A(n8644), .B(n8643), .Z(n8695) );
  XNOR U9200 ( .A(b[17]), .B(a[41]), .Z(n8677) );
  NANDN U9201 ( .A(n8677), .B(n32543), .Z(n8301) );
  NANDN U9202 ( .A(n8299), .B(n32541), .Z(n8300) );
  NAND U9203 ( .A(n8301), .B(n8300), .Z(n8618) );
  XOR U9204 ( .A(b[37]), .B(n16220), .Z(n8552) );
  NANDN U9205 ( .A(n8552), .B(n36311), .Z(n8304) );
  NANDN U9206 ( .A(n8302), .B(n36309), .Z(n8303) );
  NAND U9207 ( .A(n8304), .B(n8303), .Z(n8615) );
  XNOR U9208 ( .A(b[41]), .B(a[17]), .Z(n8653) );
  OR U9209 ( .A(n8653), .B(n36905), .Z(n8307) );
  NANDN U9210 ( .A(n8305), .B(n36807), .Z(n8306) );
  AND U9211 ( .A(n8307), .B(n8306), .Z(n8616) );
  XNOR U9212 ( .A(n8615), .B(n8616), .Z(n8617) );
  XNOR U9213 ( .A(n8618), .B(n8617), .Z(n8696) );
  XOR U9214 ( .A(n8695), .B(n8696), .Z(n8697) );
  XNOR U9215 ( .A(n8698), .B(n8697), .Z(n8704) );
  NANDN U9216 ( .A(n8309), .B(n8308), .Z(n8313) );
  NAND U9217 ( .A(n8311), .B(n8310), .Z(n8312) );
  NAND U9218 ( .A(n8313), .B(n8312), .Z(n8701) );
  NANDN U9219 ( .A(n8315), .B(n8314), .Z(n8319) );
  NAND U9220 ( .A(n8317), .B(n8316), .Z(n8318) );
  AND U9221 ( .A(n8319), .B(n8318), .Z(n8702) );
  XNOR U9222 ( .A(n8701), .B(n8702), .Z(n8703) );
  XOR U9223 ( .A(n8704), .B(n8703), .Z(n8593) );
  NANDN U9224 ( .A(n8321), .B(n8320), .Z(n8325) );
  NANDN U9225 ( .A(n8323), .B(n8322), .Z(n8324) );
  NAND U9226 ( .A(n8325), .B(n8324), .Z(n8592) );
  NANDN U9227 ( .A(n8327), .B(n8326), .Z(n8331) );
  NAND U9228 ( .A(n8329), .B(n8328), .Z(n8330) );
  AND U9229 ( .A(n8331), .B(n8330), .Z(n8579) );
  OR U9230 ( .A(n8333), .B(n8332), .Z(n8337) );
  NANDN U9231 ( .A(n8335), .B(n8334), .Z(n8336) );
  NAND U9232 ( .A(n8337), .B(n8336), .Z(n8580) );
  XNOR U9233 ( .A(n8579), .B(n8580), .Z(n8581) );
  XOR U9234 ( .A(b[15]), .B(n21996), .Z(n8662) );
  OR U9235 ( .A(n8662), .B(n32010), .Z(n8340) );
  NANDN U9236 ( .A(n8338), .B(n32011), .Z(n8339) );
  NAND U9237 ( .A(n8340), .B(n8339), .Z(n8566) );
  XNOR U9238 ( .A(b[45]), .B(a[13]), .Z(n8683) );
  NANDN U9239 ( .A(n8683), .B(n37261), .Z(n8343) );
  NANDN U9240 ( .A(n8341), .B(n37262), .Z(n8342) );
  NAND U9241 ( .A(n8343), .B(n8342), .Z(n8563) );
  NAND U9242 ( .A(n37469), .B(n8344), .Z(n8346) );
  XOR U9243 ( .A(n978), .B(n12830), .Z(n8665) );
  NAND U9244 ( .A(n8665), .B(n37471), .Z(n8345) );
  AND U9245 ( .A(n8346), .B(n8345), .Z(n8564) );
  XNOR U9246 ( .A(n8563), .B(n8564), .Z(n8565) );
  XNOR U9247 ( .A(n8566), .B(n8565), .Z(n8534) );
  NAND U9248 ( .A(n35188), .B(n8347), .Z(n8349) );
  XOR U9249 ( .A(n35540), .B(n18003), .Z(n8716) );
  NANDN U9250 ( .A(n34968), .B(n8716), .Z(n8348) );
  NAND U9251 ( .A(n8349), .B(n8348), .Z(n8572) );
  XOR U9252 ( .A(b[53]), .B(n11202), .Z(n8555) );
  NANDN U9253 ( .A(n8555), .B(n37940), .Z(n8352) );
  NANDN U9254 ( .A(n8350), .B(n37941), .Z(n8351) );
  NAND U9255 ( .A(n8352), .B(n8351), .Z(n8569) );
  XOR U9256 ( .A(b[5]), .B(n25001), .Z(n8692) );
  OR U9257 ( .A(n8692), .B(n29363), .Z(n8355) );
  NANDN U9258 ( .A(n8353), .B(n29864), .Z(n8354) );
  AND U9259 ( .A(n8355), .B(n8354), .Z(n8570) );
  XNOR U9260 ( .A(n8569), .B(n8570), .Z(n8571) );
  XNOR U9261 ( .A(n8572), .B(n8571), .Z(n8531) );
  NANDN U9262 ( .A(n8357), .B(n8356), .Z(n8361) );
  NAND U9263 ( .A(n8359), .B(n8358), .Z(n8360) );
  NAND U9264 ( .A(n8361), .B(n8360), .Z(n8532) );
  XNOR U9265 ( .A(n8531), .B(n8532), .Z(n8533) );
  XOR U9266 ( .A(n8534), .B(n8533), .Z(n8582) );
  OR U9267 ( .A(n8363), .B(n8362), .Z(n8367) );
  NANDN U9268 ( .A(n8365), .B(n8364), .Z(n8366) );
  NAND U9269 ( .A(n8367), .B(n8366), .Z(n8586) );
  XNOR U9270 ( .A(n8585), .B(n8586), .Z(n8588) );
  NANDN U9271 ( .A(n8369), .B(n8368), .Z(n8373) );
  NAND U9272 ( .A(n8371), .B(n8370), .Z(n8372) );
  NAND U9273 ( .A(n8373), .B(n8372), .Z(n8605) );
  XNOR U9274 ( .A(b[35]), .B(a[23]), .Z(n8543) );
  NANDN U9275 ( .A(n8543), .B(n35985), .Z(n8376) );
  NANDN U9276 ( .A(n8374), .B(n35986), .Z(n8375) );
  NAND U9277 ( .A(n8376), .B(n8375), .Z(n8737) );
  XOR U9278 ( .A(b[9]), .B(n23852), .Z(n8549) );
  NANDN U9279 ( .A(n8549), .B(n30509), .Z(n8379) );
  NANDN U9280 ( .A(n8377), .B(n30846), .Z(n8378) );
  NAND U9281 ( .A(n8379), .B(n8378), .Z(n8734) );
  XOR U9282 ( .A(n31123), .B(n24288), .Z(n8689) );
  NAND U9283 ( .A(n8689), .B(n29949), .Z(n8382) );
  NAND U9284 ( .A(n29948), .B(n8380), .Z(n8381) );
  AND U9285 ( .A(n8382), .B(n8381), .Z(n8735) );
  XNOR U9286 ( .A(n8734), .B(n8735), .Z(n8736) );
  XNOR U9287 ( .A(n8737), .B(n8736), .Z(n8603) );
  ANDN U9288 ( .B(n8383), .A(b[55]), .Z(n8384) );
  OR U9289 ( .A(n8384), .B(n986), .Z(n8385) );
  AND U9290 ( .A(b[56]), .B(b[55]), .Z(n38247) );
  NOR U9291 ( .A(n983), .B(n38247), .Z(n38329) );
  AND U9292 ( .A(n8385), .B(n38329), .Z(n8708) );
  XOR U9293 ( .A(b[3]), .B(n25466), .Z(n8632) );
  NANDN U9294 ( .A(n8632), .B(n28939), .Z(n8388) );
  NANDN U9295 ( .A(n8386), .B(n28938), .Z(n8387) );
  NAND U9296 ( .A(n8388), .B(n8387), .Z(n8707) );
  XOR U9297 ( .A(n8708), .B(n8707), .Z(n8709) );
  XNOR U9298 ( .A(n974), .B(a[25]), .Z(n8686) );
  NAND U9299 ( .A(n35620), .B(n8686), .Z(n8391) );
  NANDN U9300 ( .A(n8389), .B(n35621), .Z(n8390) );
  AND U9301 ( .A(n8391), .B(n8390), .Z(n8710) );
  XNOR U9302 ( .A(n8709), .B(n8710), .Z(n8604) );
  XOR U9303 ( .A(n8603), .B(n8604), .Z(n8606) );
  XNOR U9304 ( .A(n8605), .B(n8606), .Z(n8587) );
  XOR U9305 ( .A(n8588), .B(n8587), .Z(n8591) );
  XNOR U9306 ( .A(n8592), .B(n8591), .Z(n8594) );
  XNOR U9307 ( .A(n8593), .B(n8594), .Z(n8748) );
  OR U9308 ( .A(n8393), .B(n8392), .Z(n8397) );
  OR U9309 ( .A(n8395), .B(n8394), .Z(n8396) );
  NAND U9310 ( .A(n8397), .B(n8396), .Z(n8746) );
  XNOR U9311 ( .A(n8597), .B(n8598), .Z(n8599) );
  XNOR U9312 ( .A(n8600), .B(n8599), .Z(n8747) );
  XNOR U9313 ( .A(n8746), .B(n8747), .Z(n8749) );
  XOR U9314 ( .A(n8748), .B(n8749), .Z(n8761) );
  XNOR U9315 ( .A(n8760), .B(n8761), .Z(n8522) );
  NANDN U9316 ( .A(n8411), .B(n8410), .Z(n8415) );
  NANDN U9317 ( .A(n8413), .B(n8412), .Z(n8414) );
  NAND U9318 ( .A(n8415), .B(n8414), .Z(n8527) );
  NAND U9319 ( .A(n8417), .B(n8416), .Z(n8421) );
  NANDN U9320 ( .A(n8419), .B(n8418), .Z(n8420) );
  NAND U9321 ( .A(n8421), .B(n8420), .Z(n8526) );
  NANDN U9322 ( .A(n8423), .B(n8422), .Z(n8427) );
  NANDN U9323 ( .A(n8425), .B(n8424), .Z(n8426) );
  NAND U9324 ( .A(n8427), .B(n8426), .Z(n8740) );
  OR U9325 ( .A(n8429), .B(n8428), .Z(n8433) );
  OR U9326 ( .A(n8431), .B(n8430), .Z(n8432) );
  AND U9327 ( .A(n8433), .B(n8432), .Z(n8741) );
  XNOR U9328 ( .A(n8740), .B(n8741), .Z(n8742) );
  NANDN U9329 ( .A(n8435), .B(n8434), .Z(n8439) );
  NAND U9330 ( .A(n8437), .B(n8436), .Z(n8438) );
  NAND U9331 ( .A(n8439), .B(n8438), .Z(n8611) );
  XOR U9332 ( .A(b[43]), .B(n13976), .Z(n8680) );
  NANDN U9333 ( .A(n8680), .B(n37068), .Z(n8442) );
  NANDN U9334 ( .A(n8440), .B(n37069), .Z(n8441) );
  NAND U9335 ( .A(n8442), .B(n8441), .Z(n8650) );
  XOR U9336 ( .A(b[49]), .B(n12258), .Z(n8668) );
  OR U9337 ( .A(n8668), .B(n37756), .Z(n8445) );
  NANDN U9338 ( .A(n8443), .B(n37652), .Z(n8444) );
  NAND U9339 ( .A(n8445), .B(n8444), .Z(n8647) );
  XOR U9340 ( .A(b[51]), .B(n11694), .Z(n8656) );
  NANDN U9341 ( .A(n8656), .B(n37803), .Z(n8448) );
  NANDN U9342 ( .A(n8446), .B(n37802), .Z(n8447) );
  AND U9343 ( .A(n8448), .B(n8447), .Z(n8648) );
  XNOR U9344 ( .A(n8647), .B(n8648), .Z(n8649) );
  XNOR U9345 ( .A(n8650), .B(n8649), .Z(n8575) );
  XOR U9346 ( .A(b[39]), .B(n15113), .Z(n8719) );
  NANDN U9347 ( .A(n8719), .B(n36553), .Z(n8451) );
  NANDN U9348 ( .A(n8449), .B(n36643), .Z(n8450) );
  NAND U9349 ( .A(n8451), .B(n8450), .Z(n8638) );
  XOR U9350 ( .A(b[13]), .B(n22579), .Z(n8659) );
  OR U9351 ( .A(n8659), .B(n31550), .Z(n8454) );
  NANDN U9352 ( .A(n8452), .B(n31874), .Z(n8453) );
  NAND U9353 ( .A(n8454), .B(n8453), .Z(n8635) );
  XOR U9354 ( .A(b[11]), .B(n23149), .Z(n8546) );
  OR U9355 ( .A(n8546), .B(n31369), .Z(n8457) );
  NANDN U9356 ( .A(n8455), .B(n31119), .Z(n8456) );
  AND U9357 ( .A(n8457), .B(n8456), .Z(n8636) );
  XNOR U9358 ( .A(n8635), .B(n8636), .Z(n8637) );
  XOR U9359 ( .A(n8638), .B(n8637), .Z(n8576) );
  XNOR U9360 ( .A(n8575), .B(n8576), .Z(n8577) );
  NAND U9361 ( .A(n34044), .B(n8458), .Z(n8460) );
  XOR U9362 ( .A(n34510), .B(n20315), .Z(n8728) );
  NANDN U9363 ( .A(n33867), .B(n8728), .Z(n8459) );
  NAND U9364 ( .A(n8460), .B(n8459), .Z(n8674) );
  NAND U9365 ( .A(n33283), .B(n8461), .Z(n8463) );
  XOR U9366 ( .A(n33020), .B(n20867), .Z(n8713) );
  NANDN U9367 ( .A(n33021), .B(n8713), .Z(n8462) );
  NAND U9368 ( .A(n8463), .B(n8462), .Z(n8671) );
  NAND U9369 ( .A(n34848), .B(n8464), .Z(n8466) );
  XOR U9370 ( .A(b[27]), .B(n18639), .Z(n8731) );
  NANDN U9371 ( .A(n8731), .B(n34618), .Z(n8465) );
  AND U9372 ( .A(n8466), .B(n8465), .Z(n8672) );
  XNOR U9373 ( .A(n8671), .B(n8672), .Z(n8673) );
  XNOR U9374 ( .A(n8674), .B(n8673), .Z(n8540) );
  XNOR U9375 ( .A(b[21]), .B(n20352), .Z(n8722) );
  NANDN U9376 ( .A(n33634), .B(n8722), .Z(n8469) );
  NANDN U9377 ( .A(n8467), .B(n33464), .Z(n8468) );
  NAND U9378 ( .A(n8469), .B(n8468), .Z(n8538) );
  XNOR U9379 ( .A(b[25]), .B(n19656), .Z(n8725) );
  NANDN U9380 ( .A(n34219), .B(n8725), .Z(n8472) );
  NANDN U9381 ( .A(n8470), .B(n34217), .Z(n8471) );
  AND U9382 ( .A(n8472), .B(n8471), .Z(n8537) );
  XNOR U9383 ( .A(n8538), .B(n8537), .Z(n8539) );
  XOR U9384 ( .A(n8540), .B(n8539), .Z(n8578) );
  XOR U9385 ( .A(n8577), .B(n8578), .Z(n8609) );
  NANDN U9386 ( .A(n8474), .B(n8473), .Z(n8478) );
  NAND U9387 ( .A(n8476), .B(n8475), .Z(n8477) );
  AND U9388 ( .A(n8478), .B(n8477), .Z(n8610) );
  XNOR U9389 ( .A(n8609), .B(n8610), .Z(n8612) );
  XNOR U9390 ( .A(n8611), .B(n8612), .Z(n8743) );
  XOR U9391 ( .A(n8742), .B(n8743), .Z(n8525) );
  XNOR U9392 ( .A(n8526), .B(n8525), .Z(n8528) );
  XOR U9393 ( .A(n8527), .B(n8528), .Z(n8752) );
  NANDN U9394 ( .A(n8480), .B(n8479), .Z(n8484) );
  NAND U9395 ( .A(n8482), .B(n8481), .Z(n8483) );
  NAND U9396 ( .A(n8484), .B(n8483), .Z(n8753) );
  XNOR U9397 ( .A(n8752), .B(n8753), .Z(n8754) );
  NANDN U9398 ( .A(n8486), .B(n8485), .Z(n8490) );
  NANDN U9399 ( .A(n8488), .B(n8487), .Z(n8489) );
  NAND U9400 ( .A(n8490), .B(n8489), .Z(n8755) );
  XOR U9401 ( .A(n8754), .B(n8755), .Z(n8519) );
  NANDN U9402 ( .A(n8492), .B(n8491), .Z(n8496) );
  NAND U9403 ( .A(n8494), .B(n8493), .Z(n8495) );
  NAND U9404 ( .A(n8496), .B(n8495), .Z(n8520) );
  XNOR U9405 ( .A(n8519), .B(n8520), .Z(n8521) );
  XOR U9406 ( .A(n8522), .B(n8521), .Z(n8516) );
  XNOR U9407 ( .A(n8515), .B(n8516), .Z(n8507) );
  XOR U9408 ( .A(n8508), .B(n8507), .Z(n8509) );
  XNOR U9409 ( .A(n8510), .B(n8509), .Z(n8502) );
  XNOR U9410 ( .A(n8502), .B(sreg[121]), .Z(n8504) );
  NAND U9411 ( .A(n8497), .B(sreg[120]), .Z(n8501) );
  OR U9412 ( .A(n8499), .B(n8498), .Z(n8500) );
  AND U9413 ( .A(n8501), .B(n8500), .Z(n8503) );
  XOR U9414 ( .A(n8504), .B(n8503), .Z(c[121]) );
  NAND U9415 ( .A(n8502), .B(sreg[121]), .Z(n8506) );
  OR U9416 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U9417 ( .A(n8506), .B(n8505), .Z(n9033) );
  XNOR U9418 ( .A(n9033), .B(sreg[122]), .Z(n9035) );
  NAND U9419 ( .A(n8508), .B(n8507), .Z(n8512) );
  NAND U9420 ( .A(n8510), .B(n8509), .Z(n8511) );
  NAND U9421 ( .A(n8512), .B(n8511), .Z(n8767) );
  NANDN U9422 ( .A(n8514), .B(n8513), .Z(n8518) );
  NANDN U9423 ( .A(n8516), .B(n8515), .Z(n8517) );
  NAND U9424 ( .A(n8518), .B(n8517), .Z(n8765) );
  NANDN U9425 ( .A(n8520), .B(n8519), .Z(n8524) );
  NANDN U9426 ( .A(n8522), .B(n8521), .Z(n8523) );
  NAND U9427 ( .A(n8524), .B(n8523), .Z(n9028) );
  NAND U9428 ( .A(n8526), .B(n8525), .Z(n8530) );
  NANDN U9429 ( .A(n8528), .B(n8527), .Z(n8529) );
  NAND U9430 ( .A(n8530), .B(n8529), .Z(n9018) );
  NANDN U9431 ( .A(n8532), .B(n8531), .Z(n8536) );
  NAND U9432 ( .A(n8534), .B(n8533), .Z(n8535) );
  NAND U9433 ( .A(n8536), .B(n8535), .Z(n8910) );
  NANDN U9434 ( .A(n8538), .B(n8537), .Z(n8542) );
  NAND U9435 ( .A(n8540), .B(n8539), .Z(n8541) );
  NAND U9436 ( .A(n8542), .B(n8541), .Z(n9000) );
  XNOR U9437 ( .A(b[35]), .B(a[24]), .Z(n8868) );
  NANDN U9438 ( .A(n8868), .B(n35985), .Z(n8545) );
  NANDN U9439 ( .A(n8543), .B(n35986), .Z(n8544) );
  NAND U9440 ( .A(n8545), .B(n8544), .Z(n8779) );
  XOR U9441 ( .A(b[11]), .B(n23447), .Z(n8952) );
  OR U9442 ( .A(n8952), .B(n31369), .Z(n8548) );
  NANDN U9443 ( .A(n8546), .B(n31119), .Z(n8547) );
  NAND U9444 ( .A(n8548), .B(n8547), .Z(n8776) );
  XOR U9445 ( .A(b[9]), .B(n24671), .Z(n8832) );
  NANDN U9446 ( .A(n8832), .B(n30509), .Z(n8551) );
  NANDN U9447 ( .A(n8549), .B(n30846), .Z(n8550) );
  AND U9448 ( .A(n8551), .B(n8550), .Z(n8777) );
  XNOR U9449 ( .A(n8776), .B(n8777), .Z(n8778) );
  XNOR U9450 ( .A(n8779), .B(n8778), .Z(n8841) );
  XOR U9451 ( .A(b[37]), .B(n15963), .Z(n8838) );
  NANDN U9452 ( .A(n8838), .B(n36311), .Z(n8554) );
  NANDN U9453 ( .A(n8552), .B(n36309), .Z(n8553) );
  NAND U9454 ( .A(n8554), .B(n8553), .Z(n8970) );
  XOR U9455 ( .A(b[53]), .B(n11406), .Z(n8880) );
  NANDN U9456 ( .A(n8880), .B(n37940), .Z(n8557) );
  NANDN U9457 ( .A(n8555), .B(n37941), .Z(n8556) );
  NAND U9458 ( .A(n8557), .B(n8556), .Z(n8967) );
  XOR U9459 ( .A(b[57]), .B(n10363), .Z(n8797) );
  OR U9460 ( .A(n8797), .B(n965), .Z(n8562) );
  XNOR U9461 ( .A(n983), .B(b[56]), .Z(n8558) );
  AND U9462 ( .A(n8559), .B(n8558), .Z(n38194) );
  NAND U9463 ( .A(n8560), .B(n38194), .Z(n8561) );
  AND U9464 ( .A(n8562), .B(n8561), .Z(n8968) );
  XNOR U9465 ( .A(n8967), .B(n8968), .Z(n8969) );
  XOR U9466 ( .A(n8970), .B(n8969), .Z(n8842) );
  XNOR U9467 ( .A(n8841), .B(n8842), .Z(n8843) );
  NANDN U9468 ( .A(n8564), .B(n8563), .Z(n8568) );
  NAND U9469 ( .A(n8566), .B(n8565), .Z(n8567) );
  AND U9470 ( .A(n8568), .B(n8567), .Z(n8844) );
  XOR U9471 ( .A(n8843), .B(n8844), .Z(n8997) );
  NANDN U9472 ( .A(n8570), .B(n8569), .Z(n8574) );
  NAND U9473 ( .A(n8572), .B(n8571), .Z(n8573) );
  AND U9474 ( .A(n8574), .B(n8573), .Z(n8998) );
  XNOR U9475 ( .A(n8997), .B(n8998), .Z(n8999) );
  XNOR U9476 ( .A(n9000), .B(n8999), .Z(n8907) );
  XNOR U9477 ( .A(n8907), .B(n8908), .Z(n8909) );
  XNOR U9478 ( .A(n8910), .B(n8909), .Z(n8916) );
  OR U9479 ( .A(n8580), .B(n8579), .Z(n8584) );
  OR U9480 ( .A(n8582), .B(n8581), .Z(n8583) );
  NAND U9481 ( .A(n8584), .B(n8583), .Z(n8914) );
  OR U9482 ( .A(n8586), .B(n8585), .Z(n8590) );
  OR U9483 ( .A(n8588), .B(n8587), .Z(n8589) );
  AND U9484 ( .A(n8590), .B(n8589), .Z(n8913) );
  XOR U9485 ( .A(n8914), .B(n8913), .Z(n8915) );
  XNOR U9486 ( .A(n8916), .B(n8915), .Z(n8928) );
  NAND U9487 ( .A(n8592), .B(n8591), .Z(n8596) );
  NANDN U9488 ( .A(n8594), .B(n8593), .Z(n8595) );
  NAND U9489 ( .A(n8596), .B(n8595), .Z(n8926) );
  NANDN U9490 ( .A(n8598), .B(n8597), .Z(n8602) );
  NAND U9491 ( .A(n8600), .B(n8599), .Z(n8601) );
  AND U9492 ( .A(n8602), .B(n8601), .Z(n8925) );
  XNOR U9493 ( .A(n8926), .B(n8925), .Z(n8927) );
  XOR U9494 ( .A(n8928), .B(n8927), .Z(n9016) );
  NANDN U9495 ( .A(n8604), .B(n8603), .Z(n8608) );
  OR U9496 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U9497 ( .A(n8608), .B(n8607), .Z(n8932) );
  NAND U9498 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U9499 ( .A(n8612), .B(n8611), .Z(n8613) );
  AND U9500 ( .A(n8614), .B(n8613), .Z(n8931) );
  XNOR U9501 ( .A(n8932), .B(n8931), .Z(n8933) );
  NANDN U9502 ( .A(n8616), .B(n8615), .Z(n8620) );
  NAND U9503 ( .A(n8618), .B(n8617), .Z(n8619) );
  NAND U9504 ( .A(n8620), .B(n8619), .Z(n8848) );
  XNOR U9505 ( .A(b[57]), .B(b[58]), .Z(n38273) );
  NANDN U9506 ( .A(n38273), .B(a[0]), .Z(n8773) );
  NANDN U9507 ( .A(n966), .B(a[58]), .Z(n8621) );
  XOR U9508 ( .A(n29232), .B(n8621), .Z(n8623) );
  IV U9509 ( .A(a[57]), .Z(n26122) );
  NANDN U9510 ( .A(n26122), .B(n966), .Z(n8622) );
  AND U9511 ( .A(n8623), .B(n8622), .Z(n8771) );
  XNOR U9512 ( .A(n982), .B(a[4]), .Z(n8883) );
  NAND U9513 ( .A(n38075), .B(n8883), .Z(n8626) );
  NAND U9514 ( .A(n8624), .B(n38073), .Z(n8625) );
  AND U9515 ( .A(n8626), .B(n8625), .Z(n8770) );
  XNOR U9516 ( .A(n8771), .B(n8770), .Z(n8772) );
  XNOR U9517 ( .A(n8773), .B(n8772), .Z(n8847) );
  XNOR U9518 ( .A(n8848), .B(n8847), .Z(n8850) );
  NAND U9519 ( .A(n8628), .B(n8627), .Z(n8976) );
  NANDN U9520 ( .A(n8629), .B(n35311), .Z(n8631) );
  XOR U9521 ( .A(b[31]), .B(n17702), .Z(n8808) );
  NANDN U9522 ( .A(n8808), .B(n35313), .Z(n8630) );
  NAND U9523 ( .A(n8631), .B(n8630), .Z(n8974) );
  XNOR U9524 ( .A(n967), .B(a[56]), .Z(n8946) );
  NAND U9525 ( .A(n8946), .B(n28939), .Z(n8634) );
  NANDN U9526 ( .A(n8632), .B(n28938), .Z(n8633) );
  AND U9527 ( .A(n8634), .B(n8633), .Z(n8973) );
  XNOR U9528 ( .A(n8974), .B(n8973), .Z(n8975) );
  XNOR U9529 ( .A(n8976), .B(n8975), .Z(n8849) );
  XNOR U9530 ( .A(n8850), .B(n8849), .Z(n8991) );
  NANDN U9531 ( .A(n8636), .B(n8635), .Z(n8640) );
  NAND U9532 ( .A(n8638), .B(n8637), .Z(n8639) );
  AND U9533 ( .A(n8640), .B(n8639), .Z(n8992) );
  XNOR U9534 ( .A(n8991), .B(n8992), .Z(n8993) );
  NANDN U9535 ( .A(n8642), .B(n8641), .Z(n8646) );
  NAND U9536 ( .A(n8644), .B(n8643), .Z(n8645) );
  AND U9537 ( .A(n8646), .B(n8645), .Z(n8994) );
  XNOR U9538 ( .A(n8993), .B(n8994), .Z(n9012) );
  NANDN U9539 ( .A(n8648), .B(n8647), .Z(n8652) );
  NAND U9540 ( .A(n8650), .B(n8649), .Z(n8651) );
  NAND U9541 ( .A(n8652), .B(n8651), .Z(n8939) );
  XNOR U9542 ( .A(b[41]), .B(a[18]), .Z(n8829) );
  OR U9543 ( .A(n8829), .B(n36905), .Z(n8655) );
  NANDN U9544 ( .A(n8653), .B(n36807), .Z(n8654) );
  NAND U9545 ( .A(n8655), .B(n8654), .Z(n8820) );
  XOR U9546 ( .A(n980), .B(n11986), .Z(n8895) );
  NAND U9547 ( .A(n8895), .B(n37803), .Z(n8658) );
  NANDN U9548 ( .A(n8656), .B(n37802), .Z(n8657) );
  NAND U9549 ( .A(n8658), .B(n8657), .Z(n8817) );
  XOR U9550 ( .A(b[13]), .B(n22964), .Z(n8958) );
  OR U9551 ( .A(n8958), .B(n31550), .Z(n8661) );
  NANDN U9552 ( .A(n8659), .B(n31874), .Z(n8660) );
  AND U9553 ( .A(n8661), .B(n8660), .Z(n8818) );
  XNOR U9554 ( .A(n8817), .B(n8818), .Z(n8819) );
  XNOR U9555 ( .A(n8820), .B(n8819), .Z(n8937) );
  XOR U9556 ( .A(b[15]), .B(n22289), .Z(n8782) );
  OR U9557 ( .A(n8782), .B(n32010), .Z(n8664) );
  NANDN U9558 ( .A(n8662), .B(n32011), .Z(n8663) );
  NAND U9559 ( .A(n8664), .B(n8663), .Z(n8856) );
  NAND U9560 ( .A(n37469), .B(n8665), .Z(n8667) );
  XOR U9561 ( .A(n978), .B(n13106), .Z(n8862) );
  NAND U9562 ( .A(n8862), .B(n37471), .Z(n8666) );
  NAND U9563 ( .A(n8667), .B(n8666), .Z(n8853) );
  XOR U9564 ( .A(b[49]), .B(n12555), .Z(n8949) );
  OR U9565 ( .A(n8949), .B(n37756), .Z(n8670) );
  NANDN U9566 ( .A(n8668), .B(n37652), .Z(n8669) );
  AND U9567 ( .A(n8670), .B(n8669), .Z(n8854) );
  XNOR U9568 ( .A(n8853), .B(n8854), .Z(n8855) );
  XOR U9569 ( .A(n8856), .B(n8855), .Z(n8938) );
  XOR U9570 ( .A(n8937), .B(n8938), .Z(n8940) );
  XNOR U9571 ( .A(n8939), .B(n8940), .Z(n9009) );
  NANDN U9572 ( .A(n8672), .B(n8671), .Z(n8676) );
  NAND U9573 ( .A(n8674), .B(n8673), .Z(n8675) );
  NAND U9574 ( .A(n8676), .B(n8675), .Z(n8987) );
  XNOR U9575 ( .A(b[17]), .B(a[42]), .Z(n8788) );
  NANDN U9576 ( .A(n8788), .B(n32543), .Z(n8679) );
  NANDN U9577 ( .A(n8677), .B(n32541), .Z(n8678) );
  NAND U9578 ( .A(n8679), .B(n8678), .Z(n8889) );
  XOR U9579 ( .A(b[43]), .B(n14259), .Z(n8874) );
  NANDN U9580 ( .A(n8874), .B(n37068), .Z(n8682) );
  NANDN U9581 ( .A(n8680), .B(n37069), .Z(n8681) );
  NAND U9582 ( .A(n8682), .B(n8681), .Z(n8886) );
  XNOR U9583 ( .A(b[45]), .B(a[14]), .Z(n8859) );
  NANDN U9584 ( .A(n8859), .B(n37261), .Z(n8685) );
  NANDN U9585 ( .A(n8683), .B(n37262), .Z(n8684) );
  AND U9586 ( .A(n8685), .B(n8684), .Z(n8887) );
  XNOR U9587 ( .A(n8886), .B(n8887), .Z(n8888) );
  XNOR U9588 ( .A(n8889), .B(n8888), .Z(n8985) );
  XOR U9589 ( .A(b[33]), .B(n17133), .Z(n8943) );
  NANDN U9590 ( .A(n8943), .B(n35620), .Z(n8688) );
  NAND U9591 ( .A(n8686), .B(n35621), .Z(n8687) );
  NAND U9592 ( .A(n8688), .B(n8687), .Z(n8904) );
  XOR U9593 ( .A(n31123), .B(n25134), .Z(n8823) );
  NAND U9594 ( .A(n8823), .B(n29949), .Z(n8691) );
  NAND U9595 ( .A(n29948), .B(n8689), .Z(n8690) );
  NAND U9596 ( .A(n8691), .B(n8690), .Z(n8901) );
  XOR U9597 ( .A(b[5]), .B(n25177), .Z(n8871) );
  OR U9598 ( .A(n8871), .B(n29363), .Z(n8694) );
  NANDN U9599 ( .A(n8692), .B(n29864), .Z(n8693) );
  AND U9600 ( .A(n8694), .B(n8693), .Z(n8902) );
  XNOR U9601 ( .A(n8901), .B(n8902), .Z(n8903) );
  XOR U9602 ( .A(n8904), .B(n8903), .Z(n8986) );
  XOR U9603 ( .A(n8985), .B(n8986), .Z(n8988) );
  XOR U9604 ( .A(n8987), .B(n8988), .Z(n9010) );
  XNOR U9605 ( .A(n9009), .B(n9010), .Z(n9011) );
  XOR U9606 ( .A(n9012), .B(n9011), .Z(n8934) );
  XNOR U9607 ( .A(n8933), .B(n8934), .Z(n8921) );
  OR U9608 ( .A(n8696), .B(n8695), .Z(n8700) );
  NAND U9609 ( .A(n8698), .B(n8697), .Z(n8699) );
  NAND U9610 ( .A(n8700), .B(n8699), .Z(n9004) );
  NANDN U9611 ( .A(n8702), .B(n8701), .Z(n8706) );
  NANDN U9612 ( .A(n8704), .B(n8703), .Z(n8705) );
  AND U9613 ( .A(n8706), .B(n8705), .Z(n9003) );
  XNOR U9614 ( .A(n9004), .B(n9003), .Z(n9005) );
  OR U9615 ( .A(n8708), .B(n8707), .Z(n8712) );
  NAND U9616 ( .A(n8710), .B(n8709), .Z(n8711) );
  NAND U9617 ( .A(n8712), .B(n8711), .Z(n8982) );
  NAND U9618 ( .A(n33283), .B(n8713), .Z(n8715) );
  XOR U9619 ( .A(n33020), .B(n21149), .Z(n8785) );
  NANDN U9620 ( .A(n33021), .B(n8785), .Z(n8714) );
  NAND U9621 ( .A(n8715), .B(n8714), .Z(n8794) );
  NAND U9622 ( .A(n35188), .B(n8716), .Z(n8718) );
  XOR U9623 ( .A(n35540), .B(n18804), .Z(n8877) );
  NANDN U9624 ( .A(n34968), .B(n8877), .Z(n8717) );
  NAND U9625 ( .A(n8718), .B(n8717), .Z(n8791) );
  XOR U9626 ( .A(b[39]), .B(n15484), .Z(n8826) );
  NANDN U9627 ( .A(n8826), .B(n36553), .Z(n8721) );
  NANDN U9628 ( .A(n8719), .B(n36643), .Z(n8720) );
  AND U9629 ( .A(n8721), .B(n8720), .Z(n8792) );
  XNOR U9630 ( .A(n8791), .B(n8792), .Z(n8793) );
  XOR U9631 ( .A(n8794), .B(n8793), .Z(n8813) );
  XNOR U9632 ( .A(b[21]), .B(a[38]), .Z(n8955) );
  OR U9633 ( .A(n8955), .B(n33634), .Z(n8724) );
  NAND U9634 ( .A(n8722), .B(n33464), .Z(n8723) );
  NAND U9635 ( .A(n8724), .B(n8723), .Z(n8964) );
  XNOR U9636 ( .A(b[25]), .B(n19513), .Z(n8865) );
  NANDN U9637 ( .A(n34219), .B(n8865), .Z(n8727) );
  NAND U9638 ( .A(n8725), .B(n34217), .Z(n8726) );
  NAND U9639 ( .A(n8727), .B(n8726), .Z(n8961) );
  NAND U9640 ( .A(n34044), .B(n8728), .Z(n8730) );
  XOR U9641 ( .A(n34510), .B(n19980), .Z(n8835) );
  NANDN U9642 ( .A(n33867), .B(n8835), .Z(n8729) );
  AND U9643 ( .A(n8730), .B(n8729), .Z(n8962) );
  XNOR U9644 ( .A(n8961), .B(n8962), .Z(n8963) );
  XOR U9645 ( .A(n8964), .B(n8963), .Z(n8811) );
  NANDN U9646 ( .A(n8731), .B(n34848), .Z(n8733) );
  XOR U9647 ( .A(b[27]), .B(n18841), .Z(n8898) );
  NANDN U9648 ( .A(n8898), .B(n34618), .Z(n8732) );
  NAND U9649 ( .A(n8733), .B(n8732), .Z(n8812) );
  XNOR U9650 ( .A(n8811), .B(n8812), .Z(n8814) );
  XNOR U9651 ( .A(n8813), .B(n8814), .Z(n8980) );
  NANDN U9652 ( .A(n8735), .B(n8734), .Z(n8739) );
  NAND U9653 ( .A(n8737), .B(n8736), .Z(n8738) );
  AND U9654 ( .A(n8739), .B(n8738), .Z(n8979) );
  XNOR U9655 ( .A(n8980), .B(n8979), .Z(n8981) );
  XNOR U9656 ( .A(n8982), .B(n8981), .Z(n9006) );
  XOR U9657 ( .A(n9005), .B(n9006), .Z(n8919) );
  NANDN U9658 ( .A(n8741), .B(n8740), .Z(n8745) );
  NAND U9659 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U9660 ( .A(n8745), .B(n8744), .Z(n8920) );
  XNOR U9661 ( .A(n8919), .B(n8920), .Z(n8922) );
  XOR U9662 ( .A(n8921), .B(n8922), .Z(n9015) );
  XNOR U9663 ( .A(n9016), .B(n9015), .Z(n9017) );
  XNOR U9664 ( .A(n9018), .B(n9017), .Z(n9024) );
  NANDN U9665 ( .A(n8747), .B(n8746), .Z(n8751) );
  NAND U9666 ( .A(n8749), .B(n8748), .Z(n8750) );
  NAND U9667 ( .A(n8751), .B(n8750), .Z(n9021) );
  NANDN U9668 ( .A(n8753), .B(n8752), .Z(n8757) );
  NANDN U9669 ( .A(n8755), .B(n8754), .Z(n8756) );
  NAND U9670 ( .A(n8757), .B(n8756), .Z(n9022) );
  XNOR U9671 ( .A(n9021), .B(n9022), .Z(n9023) );
  XNOR U9672 ( .A(n9024), .B(n9023), .Z(n9027) );
  XNOR U9673 ( .A(n9028), .B(n9027), .Z(n9030) );
  OR U9674 ( .A(n8759), .B(n8758), .Z(n8763) );
  NANDN U9675 ( .A(n8761), .B(n8760), .Z(n8762) );
  AND U9676 ( .A(n8763), .B(n8762), .Z(n9029) );
  XNOR U9677 ( .A(n9030), .B(n9029), .Z(n8764) );
  XOR U9678 ( .A(n8765), .B(n8764), .Z(n8766) );
  XOR U9679 ( .A(n8767), .B(n8766), .Z(n9034) );
  XOR U9680 ( .A(n9035), .B(n9034), .Z(c[122]) );
  NAND U9681 ( .A(n8765), .B(n8764), .Z(n8769) );
  NAND U9682 ( .A(n8767), .B(n8766), .Z(n8768) );
  NAND U9683 ( .A(n8769), .B(n8768), .Z(n9046) );
  NANDN U9684 ( .A(n8771), .B(n8770), .Z(n8775) );
  NAND U9685 ( .A(n8773), .B(n8772), .Z(n8774) );
  NAND U9686 ( .A(n8775), .B(n8774), .Z(n9061) );
  NANDN U9687 ( .A(n8777), .B(n8776), .Z(n8781) );
  NAND U9688 ( .A(n8779), .B(n8778), .Z(n8780) );
  NAND U9689 ( .A(n8781), .B(n8780), .Z(n9062) );
  XNOR U9690 ( .A(n9061), .B(n9062), .Z(n9063) );
  XOR U9691 ( .A(b[15]), .B(n22579), .Z(n9179) );
  OR U9692 ( .A(n9179), .B(n32010), .Z(n8784) );
  NANDN U9693 ( .A(n8782), .B(n32011), .Z(n8783) );
  NAND U9694 ( .A(n8784), .B(n8783), .Z(n9200) );
  NAND U9695 ( .A(n33283), .B(n8785), .Z(n8787) );
  XOR U9696 ( .A(b[19]), .B(n21441), .Z(n9275) );
  OR U9697 ( .A(n9275), .B(n33021), .Z(n8786) );
  NAND U9698 ( .A(n8787), .B(n8786), .Z(n9197) );
  XNOR U9699 ( .A(b[17]), .B(a[43]), .Z(n9170) );
  NANDN U9700 ( .A(n9170), .B(n32543), .Z(n8790) );
  NANDN U9701 ( .A(n8788), .B(n32541), .Z(n8789) );
  AND U9702 ( .A(n8790), .B(n8789), .Z(n9198) );
  XNOR U9703 ( .A(n9197), .B(n9198), .Z(n9199) );
  XOR U9704 ( .A(n9200), .B(n9199), .Z(n9239) );
  NANDN U9705 ( .A(n8792), .B(n8791), .Z(n8796) );
  NAND U9706 ( .A(n8794), .B(n8793), .Z(n8795) );
  NAND U9707 ( .A(n8796), .B(n8795), .Z(n9240) );
  XNOR U9708 ( .A(n9239), .B(n9240), .Z(n9242) );
  XOR U9709 ( .A(n983), .B(n10524), .Z(n9167) );
  NANDN U9710 ( .A(n965), .B(n9167), .Z(n8799) );
  NANDN U9711 ( .A(n8797), .B(n38194), .Z(n8798) );
  NAND U9712 ( .A(n8799), .B(n8798), .Z(n9089) );
  IV U9713 ( .A(b[59]), .Z(n38400) );
  XNOR U9714 ( .A(n38400), .B(a[0]), .Z(n8802) );
  XNOR U9715 ( .A(n38400), .B(b[57]), .Z(n9091) );
  XOR U9716 ( .A(b[59]), .B(b[58]), .Z(n8800) );
  AND U9717 ( .A(n9091), .B(n8800), .Z(n8801) );
  NAND U9718 ( .A(n8802), .B(n8801), .Z(n8804) );
  XOR U9719 ( .A(b[59]), .B(n10457), .Z(n9092) );
  OR U9720 ( .A(n9092), .B(n38273), .Z(n8803) );
  NAND U9721 ( .A(n8804), .B(n8803), .Z(n9088) );
  XNOR U9722 ( .A(n9089), .B(n9088), .Z(n9254) );
  NANDN U9723 ( .A(n38400), .B(n983), .Z(n8805) );
  OR U9724 ( .A(n8805), .B(b[58]), .Z(n8807) );
  ANDN U9725 ( .B(b[59]), .A(n38273), .Z(n38327) );
  NANDN U9726 ( .A(a[0]), .B(n38327), .Z(n8806) );
  NAND U9727 ( .A(n8807), .B(n8806), .Z(n9252) );
  NANDN U9728 ( .A(n8808), .B(n35311), .Z(n8810) );
  XNOR U9729 ( .A(n973), .B(a[29]), .Z(n9257) );
  NAND U9730 ( .A(n9257), .B(n35313), .Z(n8809) );
  AND U9731 ( .A(n8810), .B(n8809), .Z(n9251) );
  XNOR U9732 ( .A(n9252), .B(n9251), .Z(n9253) );
  XOR U9733 ( .A(n9254), .B(n9253), .Z(n9241) );
  XNOR U9734 ( .A(n9242), .B(n9241), .Z(n9064) );
  XOR U9735 ( .A(n9063), .B(n9064), .Z(n9229) );
  OR U9736 ( .A(n8812), .B(n8811), .Z(n8816) );
  OR U9737 ( .A(n8814), .B(n8813), .Z(n8815) );
  NAND U9738 ( .A(n8816), .B(n8815), .Z(n9228) );
  NANDN U9739 ( .A(n8818), .B(n8817), .Z(n8822) );
  NAND U9740 ( .A(n8820), .B(n8819), .Z(n8821) );
  NAND U9741 ( .A(n8822), .B(n8821), .Z(n9211) );
  XOR U9742 ( .A(n31123), .B(n25001), .Z(n9137) );
  NAND U9743 ( .A(n9137), .B(n29949), .Z(n8825) );
  NAND U9744 ( .A(n29948), .B(n8823), .Z(n8824) );
  NAND U9745 ( .A(n8825), .B(n8824), .Z(n9143) );
  XOR U9746 ( .A(b[39]), .B(n16220), .Z(n9122) );
  NANDN U9747 ( .A(n9122), .B(n36553), .Z(n8828) );
  NANDN U9748 ( .A(n8826), .B(n36643), .Z(n8827) );
  NAND U9749 ( .A(n8828), .B(n8827), .Z(n9140) );
  XNOR U9750 ( .A(b[41]), .B(a[19]), .Z(n9176) );
  OR U9751 ( .A(n9176), .B(n36905), .Z(n8831) );
  NANDN U9752 ( .A(n8829), .B(n36807), .Z(n8830) );
  AND U9753 ( .A(n8831), .B(n8830), .Z(n9141) );
  XNOR U9754 ( .A(n9140), .B(n9141), .Z(n9142) );
  XNOR U9755 ( .A(n9143), .B(n9142), .Z(n9209) );
  XOR U9756 ( .A(b[9]), .B(n24288), .Z(n9134) );
  NANDN U9757 ( .A(n9134), .B(n30509), .Z(n8834) );
  NANDN U9758 ( .A(n8832), .B(n30846), .Z(n8833) );
  NAND U9759 ( .A(n8834), .B(n8833), .Z(n9161) );
  NAND U9760 ( .A(n34044), .B(n8835), .Z(n8837) );
  XOR U9761 ( .A(n34510), .B(n20352), .Z(n9266) );
  NANDN U9762 ( .A(n33867), .B(n9266), .Z(n8836) );
  NAND U9763 ( .A(n8837), .B(n8836), .Z(n9158) );
  XOR U9764 ( .A(b[37]), .B(n16269), .Z(n9131) );
  NANDN U9765 ( .A(n9131), .B(n36311), .Z(n8840) );
  NANDN U9766 ( .A(n8838), .B(n36309), .Z(n8839) );
  AND U9767 ( .A(n8840), .B(n8839), .Z(n9159) );
  XNOR U9768 ( .A(n9158), .B(n9159), .Z(n9160) );
  XOR U9769 ( .A(n9161), .B(n9160), .Z(n9210) );
  XOR U9770 ( .A(n9209), .B(n9210), .Z(n9212) );
  XOR U9771 ( .A(n9211), .B(n9212), .Z(n9227) );
  XNOR U9772 ( .A(n9228), .B(n9227), .Z(n9230) );
  XOR U9773 ( .A(n9229), .B(n9230), .Z(n9281) );
  NANDN U9774 ( .A(n8842), .B(n8841), .Z(n8846) );
  NAND U9775 ( .A(n8844), .B(n8843), .Z(n8845) );
  NAND U9776 ( .A(n8846), .B(n8845), .Z(n9236) );
  OR U9777 ( .A(n8848), .B(n8847), .Z(n8852) );
  OR U9778 ( .A(n8850), .B(n8849), .Z(n8851) );
  NAND U9779 ( .A(n8852), .B(n8851), .Z(n9233) );
  NANDN U9780 ( .A(n8854), .B(n8853), .Z(n8858) );
  NAND U9781 ( .A(n8856), .B(n8855), .Z(n8857) );
  NAND U9782 ( .A(n8858), .B(n8857), .Z(n9118) );
  XNOR U9783 ( .A(b[45]), .B(a[15]), .Z(n9185) );
  NANDN U9784 ( .A(n9185), .B(n37261), .Z(n8861) );
  NANDN U9785 ( .A(n8859), .B(n37262), .Z(n8860) );
  NAND U9786 ( .A(n8861), .B(n8860), .Z(n9107) );
  NAND U9787 ( .A(n37469), .B(n8862), .Z(n8864) );
  XOR U9788 ( .A(n978), .B(n13509), .Z(n9076) );
  NAND U9789 ( .A(n9076), .B(n37471), .Z(n8863) );
  NAND U9790 ( .A(n8864), .B(n8863), .Z(n9104) );
  XNOR U9791 ( .A(b[25]), .B(n20315), .Z(n9269) );
  NANDN U9792 ( .A(n34219), .B(n9269), .Z(n8867) );
  NAND U9793 ( .A(n34217), .B(n8865), .Z(n8866) );
  AND U9794 ( .A(n8867), .B(n8866), .Z(n9105) );
  XNOR U9795 ( .A(n9104), .B(n9105), .Z(n9106) );
  XNOR U9796 ( .A(n9107), .B(n9106), .Z(n9116) );
  XNOR U9797 ( .A(b[35]), .B(a[25]), .Z(n9188) );
  NANDN U9798 ( .A(n9188), .B(n35985), .Z(n8870) );
  NANDN U9799 ( .A(n8868), .B(n35986), .Z(n8869) );
  NAND U9800 ( .A(n8870), .B(n8869), .Z(n9085) );
  XOR U9801 ( .A(b[5]), .B(n25466), .Z(n9194) );
  OR U9802 ( .A(n9194), .B(n29363), .Z(n8873) );
  NANDN U9803 ( .A(n8871), .B(n29864), .Z(n8872) );
  NAND U9804 ( .A(n8873), .B(n8872), .Z(n9082) );
  XOR U9805 ( .A(b[43]), .B(n14514), .Z(n9182) );
  NANDN U9806 ( .A(n9182), .B(n37068), .Z(n8876) );
  NANDN U9807 ( .A(n8874), .B(n37069), .Z(n8875) );
  AND U9808 ( .A(n8876), .B(n8875), .Z(n9083) );
  XNOR U9809 ( .A(n9082), .B(n9083), .Z(n9084) );
  XOR U9810 ( .A(n9085), .B(n9084), .Z(n9117) );
  XOR U9811 ( .A(n9116), .B(n9117), .Z(n9119) );
  XNOR U9812 ( .A(n9118), .B(n9119), .Z(n9113) );
  NAND U9813 ( .A(n35188), .B(n8877), .Z(n8879) );
  XOR U9814 ( .A(n35540), .B(n18639), .Z(n9173) );
  NANDN U9815 ( .A(n34968), .B(n9173), .Z(n8878) );
  NAND U9816 ( .A(n8879), .B(n8878), .Z(n9155) );
  XOR U9817 ( .A(b[53]), .B(n11694), .Z(n9191) );
  NANDN U9818 ( .A(n9191), .B(n37940), .Z(n8882) );
  NANDN U9819 ( .A(n8880), .B(n37941), .Z(n8881) );
  NAND U9820 ( .A(n8882), .B(n8881), .Z(n9152) );
  XOR U9821 ( .A(b[55]), .B(n11202), .Z(n9263) );
  NANDN U9822 ( .A(n9263), .B(n38075), .Z(n8885) );
  NAND U9823 ( .A(n8883), .B(n38073), .Z(n8884) );
  AND U9824 ( .A(n8885), .B(n8884), .Z(n9153) );
  XNOR U9825 ( .A(n9152), .B(n9153), .Z(n9154) );
  XNOR U9826 ( .A(n9155), .B(n9154), .Z(n9215) );
  NANDN U9827 ( .A(n8887), .B(n8886), .Z(n8891) );
  NAND U9828 ( .A(n8889), .B(n8888), .Z(n8890) );
  NAND U9829 ( .A(n8891), .B(n8890), .Z(n9216) );
  XOR U9830 ( .A(n9215), .B(n9216), .Z(n9218) );
  NANDN U9831 ( .A(n966), .B(a[59]), .Z(n8892) );
  XOR U9832 ( .A(n29232), .B(n8892), .Z(n8894) );
  IV U9833 ( .A(a[58]), .Z(n26347) );
  NANDN U9834 ( .A(n26347), .B(n966), .Z(n8893) );
  AND U9835 ( .A(n8894), .B(n8893), .Z(n9099) );
  NAND U9836 ( .A(n37802), .B(n8895), .Z(n8897) );
  XOR U9837 ( .A(b[51]), .B(n12258), .Z(n9073) );
  NANDN U9838 ( .A(n9073), .B(n37803), .Z(n8896) );
  AND U9839 ( .A(n8897), .B(n8896), .Z(n9098) );
  XNOR U9840 ( .A(n9099), .B(n9098), .Z(n9100) );
  NANDN U9841 ( .A(n8898), .B(n34848), .Z(n8900) );
  XNOR U9842 ( .A(n35375), .B(a[33]), .Z(n9272) );
  NAND U9843 ( .A(n34618), .B(n9272), .Z(n8899) );
  AND U9844 ( .A(n8900), .B(n8899), .Z(n9101) );
  XNOR U9845 ( .A(n9100), .B(n9101), .Z(n9217) );
  XNOR U9846 ( .A(n9218), .B(n9217), .Z(n9110) );
  NANDN U9847 ( .A(n8902), .B(n8901), .Z(n8906) );
  NAND U9848 ( .A(n8904), .B(n8903), .Z(n8905) );
  AND U9849 ( .A(n8906), .B(n8905), .Z(n9111) );
  XNOR U9850 ( .A(n9110), .B(n9111), .Z(n9112) );
  XOR U9851 ( .A(n9113), .B(n9112), .Z(n9234) );
  XNOR U9852 ( .A(n9233), .B(n9234), .Z(n9235) );
  XOR U9853 ( .A(n9236), .B(n9235), .Z(n9282) );
  XNOR U9854 ( .A(n9281), .B(n9282), .Z(n9283) );
  NANDN U9855 ( .A(n8908), .B(n8907), .Z(n8912) );
  NAND U9856 ( .A(n8910), .B(n8909), .Z(n8911) );
  AND U9857 ( .A(n8912), .B(n8911), .Z(n9284) );
  XNOR U9858 ( .A(n9283), .B(n9284), .Z(n9052) );
  OR U9859 ( .A(n8914), .B(n8913), .Z(n8918) );
  NANDN U9860 ( .A(n8916), .B(n8915), .Z(n8917) );
  NAND U9861 ( .A(n8918), .B(n8917), .Z(n9050) );
  NANDN U9862 ( .A(n8920), .B(n8919), .Z(n8924) );
  NAND U9863 ( .A(n8922), .B(n8921), .Z(n8923) );
  AND U9864 ( .A(n8924), .B(n8923), .Z(n9049) );
  XOR U9865 ( .A(n9050), .B(n9049), .Z(n9051) );
  XNOR U9866 ( .A(n9052), .B(n9051), .Z(n9300) );
  NANDN U9867 ( .A(n8926), .B(n8925), .Z(n8930) );
  NANDN U9868 ( .A(n8928), .B(n8927), .Z(n8929) );
  NAND U9869 ( .A(n8930), .B(n8929), .Z(n9297) );
  NANDN U9870 ( .A(n8932), .B(n8931), .Z(n8936) );
  NANDN U9871 ( .A(n8934), .B(n8933), .Z(n8935) );
  NAND U9872 ( .A(n8936), .B(n8935), .Z(n9290) );
  NANDN U9873 ( .A(n8938), .B(n8937), .Z(n8942) );
  OR U9874 ( .A(n8940), .B(n8939), .Z(n8941) );
  NAND U9875 ( .A(n8942), .B(n8941), .Z(n9058) );
  XOR U9876 ( .A(b[33]), .B(n17960), .Z(n9095) );
  NANDN U9877 ( .A(n9095), .B(n35620), .Z(n8945) );
  NANDN U9878 ( .A(n8943), .B(n35621), .Z(n8944) );
  NAND U9879 ( .A(n8945), .B(n8944), .Z(n9206) );
  XOR U9880 ( .A(n967), .B(n26122), .Z(n9260) );
  NAND U9881 ( .A(n9260), .B(n28939), .Z(n8948) );
  NAND U9882 ( .A(n8946), .B(n28938), .Z(n8947) );
  NAND U9883 ( .A(n8948), .B(n8947), .Z(n9203) );
  XOR U9884 ( .A(b[49]), .B(n12830), .Z(n9079) );
  OR U9885 ( .A(n9079), .B(n37756), .Z(n8951) );
  NANDN U9886 ( .A(n8949), .B(n37652), .Z(n8950) );
  AND U9887 ( .A(n8951), .B(n8950), .Z(n9204) );
  XNOR U9888 ( .A(n9203), .B(n9204), .Z(n9205) );
  XNOR U9889 ( .A(n9206), .B(n9205), .Z(n9069) );
  XOR U9890 ( .A(b[11]), .B(n23852), .Z(n9128) );
  OR U9891 ( .A(n9128), .B(n31369), .Z(n8954) );
  NANDN U9892 ( .A(n8952), .B(n31119), .Z(n8953) );
  NAND U9893 ( .A(n8954), .B(n8953), .Z(n9149) );
  XNOR U9894 ( .A(b[21]), .B(a[39]), .Z(n9278) );
  OR U9895 ( .A(n9278), .B(n33634), .Z(n8957) );
  NANDN U9896 ( .A(n8955), .B(n33464), .Z(n8956) );
  NAND U9897 ( .A(n8957), .B(n8956), .Z(n9146) );
  XOR U9898 ( .A(b[13]), .B(n23149), .Z(n9125) );
  OR U9899 ( .A(n9125), .B(n31550), .Z(n8960) );
  NANDN U9900 ( .A(n8958), .B(n31874), .Z(n8959) );
  AND U9901 ( .A(n8960), .B(n8959), .Z(n9147) );
  XNOR U9902 ( .A(n9146), .B(n9147), .Z(n9148) );
  XNOR U9903 ( .A(n9149), .B(n9148), .Z(n9067) );
  NANDN U9904 ( .A(n8962), .B(n8961), .Z(n8966) );
  NAND U9905 ( .A(n8964), .B(n8963), .Z(n8965) );
  NAND U9906 ( .A(n8966), .B(n8965), .Z(n9068) );
  XOR U9907 ( .A(n9067), .B(n9068), .Z(n9070) );
  XNOR U9908 ( .A(n9069), .B(n9070), .Z(n9248) );
  NANDN U9909 ( .A(n8968), .B(n8967), .Z(n8972) );
  NAND U9910 ( .A(n8970), .B(n8969), .Z(n8971) );
  NAND U9911 ( .A(n8972), .B(n8971), .Z(n9245) );
  NANDN U9912 ( .A(n8974), .B(n8973), .Z(n8978) );
  NAND U9913 ( .A(n8976), .B(n8975), .Z(n8977) );
  NAND U9914 ( .A(n8978), .B(n8977), .Z(n9246) );
  XNOR U9915 ( .A(n9245), .B(n9246), .Z(n9247) );
  XNOR U9916 ( .A(n9248), .B(n9247), .Z(n9224) );
  NANDN U9917 ( .A(n8980), .B(n8979), .Z(n8984) );
  NAND U9918 ( .A(n8982), .B(n8981), .Z(n8983) );
  NAND U9919 ( .A(n8984), .B(n8983), .Z(n9221) );
  NANDN U9920 ( .A(n8986), .B(n8985), .Z(n8990) );
  OR U9921 ( .A(n8988), .B(n8987), .Z(n8989) );
  AND U9922 ( .A(n8990), .B(n8989), .Z(n9222) );
  XNOR U9923 ( .A(n9221), .B(n9222), .Z(n9223) );
  XNOR U9924 ( .A(n9224), .B(n9223), .Z(n9056) );
  NANDN U9925 ( .A(n8992), .B(n8991), .Z(n8996) );
  NAND U9926 ( .A(n8994), .B(n8993), .Z(n8995) );
  AND U9927 ( .A(n8996), .B(n8995), .Z(n9055) );
  XOR U9928 ( .A(n9056), .B(n9055), .Z(n9057) );
  XOR U9929 ( .A(n9058), .B(n9057), .Z(n9288) );
  OR U9930 ( .A(n8998), .B(n8997), .Z(n9002) );
  OR U9931 ( .A(n9000), .B(n8999), .Z(n9001) );
  NAND U9932 ( .A(n9002), .B(n9001), .Z(n9296) );
  NANDN U9933 ( .A(n9004), .B(n9003), .Z(n9008) );
  NANDN U9934 ( .A(n9006), .B(n9005), .Z(n9007) );
  NAND U9935 ( .A(n9008), .B(n9007), .Z(n9294) );
  NANDN U9936 ( .A(n9010), .B(n9009), .Z(n9014) );
  NANDN U9937 ( .A(n9012), .B(n9011), .Z(n9013) );
  AND U9938 ( .A(n9014), .B(n9013), .Z(n9293) );
  XNOR U9939 ( .A(n9294), .B(n9293), .Z(n9295) );
  XOR U9940 ( .A(n9296), .B(n9295), .Z(n9287) );
  XOR U9941 ( .A(n9288), .B(n9287), .Z(n9289) );
  XOR U9942 ( .A(n9290), .B(n9289), .Z(n9298) );
  XOR U9943 ( .A(n9297), .B(n9298), .Z(n9299) );
  XNOR U9944 ( .A(n9300), .B(n9299), .Z(n9306) );
  NANDN U9945 ( .A(n9016), .B(n9015), .Z(n9020) );
  NANDN U9946 ( .A(n9018), .B(n9017), .Z(n9019) );
  NAND U9947 ( .A(n9020), .B(n9019), .Z(n9303) );
  NANDN U9948 ( .A(n9022), .B(n9021), .Z(n9026) );
  NANDN U9949 ( .A(n9024), .B(n9023), .Z(n9025) );
  NAND U9950 ( .A(n9026), .B(n9025), .Z(n9304) );
  XNOR U9951 ( .A(n9303), .B(n9304), .Z(n9305) );
  XNOR U9952 ( .A(n9306), .B(n9305), .Z(n9044) );
  NAND U9953 ( .A(n9028), .B(n9027), .Z(n9032) );
  NANDN U9954 ( .A(n9030), .B(n9029), .Z(n9031) );
  AND U9955 ( .A(n9032), .B(n9031), .Z(n9043) );
  XOR U9956 ( .A(n9044), .B(n9043), .Z(n9045) );
  XNOR U9957 ( .A(n9046), .B(n9045), .Z(n9038) );
  XNOR U9958 ( .A(n9038), .B(sreg[123]), .Z(n9040) );
  NAND U9959 ( .A(n9033), .B(sreg[122]), .Z(n9037) );
  OR U9960 ( .A(n9035), .B(n9034), .Z(n9036) );
  AND U9961 ( .A(n9037), .B(n9036), .Z(n9039) );
  XOR U9962 ( .A(n9040), .B(n9039), .Z(c[123]) );
  NAND U9963 ( .A(n9038), .B(sreg[123]), .Z(n9042) );
  OR U9964 ( .A(n9040), .B(n9039), .Z(n9041) );
  NAND U9965 ( .A(n9042), .B(n9041), .Z(n9573) );
  XNOR U9966 ( .A(n9573), .B(sreg[124]), .Z(n9575) );
  OR U9967 ( .A(n9044), .B(n9043), .Z(n9048) );
  NAND U9968 ( .A(n9046), .B(n9045), .Z(n9047) );
  NAND U9969 ( .A(n9048), .B(n9047), .Z(n9312) );
  OR U9970 ( .A(n9050), .B(n9049), .Z(n9054) );
  NANDN U9971 ( .A(n9052), .B(n9051), .Z(n9053) );
  NAND U9972 ( .A(n9054), .B(n9053), .Z(n9318) );
  OR U9973 ( .A(n9056), .B(n9055), .Z(n9060) );
  NANDN U9974 ( .A(n9058), .B(n9057), .Z(n9059) );
  NAND U9975 ( .A(n9060), .B(n9059), .Z(n9340) );
  NANDN U9976 ( .A(n9062), .B(n9061), .Z(n9066) );
  NAND U9977 ( .A(n9064), .B(n9063), .Z(n9065) );
  NAND U9978 ( .A(n9066), .B(n9065), .Z(n9510) );
  NANDN U9979 ( .A(n9068), .B(n9067), .Z(n9072) );
  NANDN U9980 ( .A(n9070), .B(n9069), .Z(n9071) );
  AND U9981 ( .A(n9072), .B(n9071), .Z(n9511) );
  XNOR U9982 ( .A(n9510), .B(n9511), .Z(n9512) );
  XOR U9983 ( .A(b[51]), .B(n12555), .Z(n9450) );
  NANDN U9984 ( .A(n9450), .B(n37803), .Z(n9075) );
  NANDN U9985 ( .A(n9073), .B(n37802), .Z(n9074) );
  NAND U9986 ( .A(n9075), .B(n9074), .Z(n9495) );
  NAND U9987 ( .A(n37469), .B(n9076), .Z(n9078) );
  XOR U9988 ( .A(n978), .B(n14210), .Z(n9486) );
  NAND U9989 ( .A(n9486), .B(n37471), .Z(n9077) );
  NAND U9990 ( .A(n9078), .B(n9077), .Z(n9492) );
  XOR U9991 ( .A(b[49]), .B(n13106), .Z(n9489) );
  OR U9992 ( .A(n9489), .B(n37756), .Z(n9081) );
  NANDN U9993 ( .A(n9079), .B(n37652), .Z(n9080) );
  AND U9994 ( .A(n9081), .B(n9080), .Z(n9493) );
  XNOR U9995 ( .A(n9492), .B(n9493), .Z(n9494) );
  XNOR U9996 ( .A(n9495), .B(n9494), .Z(n9416) );
  NANDN U9997 ( .A(n9083), .B(n9082), .Z(n9087) );
  NAND U9998 ( .A(n9085), .B(n9084), .Z(n9086) );
  NAND U9999 ( .A(n9087), .B(n9086), .Z(n9417) );
  XNOR U10000 ( .A(n9416), .B(n9417), .Z(n9418) );
  NAND U10001 ( .A(n9089), .B(n9088), .Z(n9534) );
  XOR U10002 ( .A(n38400), .B(b[58]), .Z(n9090) );
  ANDN U10003 ( .B(n9091), .A(n9090), .Z(n38326) );
  NANDN U10004 ( .A(n9092), .B(n38326), .Z(n9094) );
  XNOR U10005 ( .A(n38400), .B(a[2]), .Z(n9372) );
  NANDN U10006 ( .A(n38273), .B(n9372), .Z(n9093) );
  NAND U10007 ( .A(n9094), .B(n9093), .Z(n9533) );
  XNOR U10008 ( .A(n974), .B(a[28]), .Z(n9474) );
  NAND U10009 ( .A(n35620), .B(n9474), .Z(n9097) );
  NANDN U10010 ( .A(n9095), .B(n35621), .Z(n9096) );
  AND U10011 ( .A(n9097), .B(n9096), .Z(n9532) );
  XNOR U10012 ( .A(n9533), .B(n9532), .Z(n9535) );
  XNOR U10013 ( .A(n9534), .B(n9535), .Z(n9419) );
  XNOR U10014 ( .A(n9418), .B(n9419), .Z(n9522) );
  NANDN U10015 ( .A(n9099), .B(n9098), .Z(n9103) );
  NAND U10016 ( .A(n9101), .B(n9100), .Z(n9102) );
  NAND U10017 ( .A(n9103), .B(n9102), .Z(n9520) );
  NANDN U10018 ( .A(n9105), .B(n9104), .Z(n9109) );
  NAND U10019 ( .A(n9107), .B(n9106), .Z(n9108) );
  NAND U10020 ( .A(n9109), .B(n9108), .Z(n9521) );
  XNOR U10021 ( .A(n9520), .B(n9521), .Z(n9523) );
  XOR U10022 ( .A(n9522), .B(n9523), .Z(n9513) );
  XNOR U10023 ( .A(n9512), .B(n9513), .Z(n9518) );
  NANDN U10024 ( .A(n9111), .B(n9110), .Z(n9115) );
  NAND U10025 ( .A(n9113), .B(n9112), .Z(n9114) );
  NAND U10026 ( .A(n9115), .B(n9114), .Z(n9517) );
  NANDN U10027 ( .A(n9117), .B(n9116), .Z(n9121) );
  OR U10028 ( .A(n9119), .B(n9118), .Z(n9120) );
  NAND U10029 ( .A(n9121), .B(n9120), .Z(n9569) );
  XOR U10030 ( .A(b[39]), .B(n15963), .Z(n9426) );
  NANDN U10031 ( .A(n9426), .B(n36553), .Z(n9124) );
  NANDN U10032 ( .A(n9122), .B(n36643), .Z(n9123) );
  NAND U10033 ( .A(n9124), .B(n9123), .Z(n9352) );
  XOR U10034 ( .A(b[13]), .B(n23447), .Z(n9459) );
  OR U10035 ( .A(n9459), .B(n31550), .Z(n9127) );
  NANDN U10036 ( .A(n9125), .B(n31874), .Z(n9126) );
  NAND U10037 ( .A(n9127), .B(n9126), .Z(n9349) );
  XOR U10038 ( .A(b[11]), .B(n24671), .Z(n9429) );
  OR U10039 ( .A(n9429), .B(n31369), .Z(n9130) );
  NANDN U10040 ( .A(n9128), .B(n31119), .Z(n9129) );
  AND U10041 ( .A(n9130), .B(n9129), .Z(n9350) );
  XNOR U10042 ( .A(n9349), .B(n9350), .Z(n9351) );
  XNOR U10043 ( .A(n9352), .B(n9351), .Z(n9423) );
  XOR U10044 ( .A(b[37]), .B(n16508), .Z(n9551) );
  NANDN U10045 ( .A(n9551), .B(n36311), .Z(n9133) );
  NANDN U10046 ( .A(n9131), .B(n36309), .Z(n9132) );
  NAND U10047 ( .A(n9133), .B(n9132), .Z(n9560) );
  XOR U10048 ( .A(b[9]), .B(n25134), .Z(n9432) );
  NANDN U10049 ( .A(n9432), .B(n30509), .Z(n9136) );
  NANDN U10050 ( .A(n9134), .B(n30846), .Z(n9135) );
  NAND U10051 ( .A(n9136), .B(n9135), .Z(n9557) );
  XOR U10052 ( .A(n31123), .B(n25177), .Z(n9438) );
  NAND U10053 ( .A(n9438), .B(n29949), .Z(n9139) );
  NAND U10054 ( .A(n29948), .B(n9137), .Z(n9138) );
  AND U10055 ( .A(n9139), .B(n9138), .Z(n9558) );
  XNOR U10056 ( .A(n9557), .B(n9558), .Z(n9559) );
  XNOR U10057 ( .A(n9560), .B(n9559), .Z(n9420) );
  NANDN U10058 ( .A(n9141), .B(n9140), .Z(n9145) );
  NAND U10059 ( .A(n9143), .B(n9142), .Z(n9144) );
  NAND U10060 ( .A(n9145), .B(n9144), .Z(n9421) );
  XNOR U10061 ( .A(n9420), .B(n9421), .Z(n9422) );
  XOR U10062 ( .A(n9423), .B(n9422), .Z(n9407) );
  NANDN U10063 ( .A(n9147), .B(n9146), .Z(n9151) );
  NAND U10064 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U10065 ( .A(n9151), .B(n9150), .Z(n9404) );
  NANDN U10066 ( .A(n9153), .B(n9152), .Z(n9157) );
  NAND U10067 ( .A(n9155), .B(n9154), .Z(n9156) );
  AND U10068 ( .A(n9157), .B(n9156), .Z(n9405) );
  XNOR U10069 ( .A(n9404), .B(n9405), .Z(n9406) );
  XNOR U10070 ( .A(n9407), .B(n9406), .Z(n9570) );
  XNOR U10071 ( .A(n9569), .B(n9570), .Z(n9572) );
  NANDN U10072 ( .A(n9159), .B(n9158), .Z(n9163) );
  NAND U10073 ( .A(n9161), .B(n9160), .Z(n9162) );
  NAND U10074 ( .A(n9163), .B(n9162), .Z(n9397) );
  XOR U10075 ( .A(b[59]), .B(b[60]), .Z(n9375) );
  AND U10076 ( .A(a[0]), .B(n9375), .Z(n9381) );
  NANDN U10077 ( .A(n966), .B(a[60]), .Z(n9164) );
  XOR U10078 ( .A(n29232), .B(n9164), .Z(n9166) );
  NANDN U10079 ( .A(b[0]), .B(a[59]), .Z(n9165) );
  AND U10080 ( .A(n9166), .B(n9165), .Z(n9355) );
  XOR U10081 ( .A(b[57]), .B(n10854), .Z(n9480) );
  OR U10082 ( .A(n9480), .B(n965), .Z(n9169) );
  NAND U10083 ( .A(n9167), .B(n38194), .Z(n9168) );
  AND U10084 ( .A(n9169), .B(n9168), .Z(n9356) );
  XOR U10085 ( .A(n9355), .B(n9356), .Z(n9357) );
  XOR U10086 ( .A(n9381), .B(n9357), .Z(n9395) );
  XNOR U10087 ( .A(b[17]), .B(a[44]), .Z(n9539) );
  NANDN U10088 ( .A(n9539), .B(n32543), .Z(n9172) );
  NANDN U10089 ( .A(n9170), .B(n32541), .Z(n9171) );
  NAND U10090 ( .A(n9172), .B(n9171), .Z(n9471) );
  NAND U10091 ( .A(n35188), .B(n9173), .Z(n9175) );
  XOR U10092 ( .A(n35540), .B(n18841), .Z(n9385) );
  NANDN U10093 ( .A(n34968), .B(n9385), .Z(n9174) );
  NAND U10094 ( .A(n9175), .B(n9174), .Z(n9468) );
  XNOR U10095 ( .A(b[41]), .B(a[20]), .Z(n9542) );
  OR U10096 ( .A(n9542), .B(n36905), .Z(n9178) );
  NANDN U10097 ( .A(n9176), .B(n36807), .Z(n9177) );
  AND U10098 ( .A(n9178), .B(n9177), .Z(n9469) );
  XNOR U10099 ( .A(n9468), .B(n9469), .Z(n9470) );
  XOR U10100 ( .A(n9471), .B(n9470), .Z(n9394) );
  XNOR U10101 ( .A(n9395), .B(n9394), .Z(n9396) );
  XNOR U10102 ( .A(n9397), .B(n9396), .Z(n9413) );
  XOR U10103 ( .A(b[15]), .B(n22964), .Z(n9536) );
  OR U10104 ( .A(n9536), .B(n32010), .Z(n9181) );
  NANDN U10105 ( .A(n9179), .B(n32011), .Z(n9180) );
  NAND U10106 ( .A(n9181), .B(n9180), .Z(n9369) );
  XOR U10107 ( .A(b[43]), .B(n14905), .Z(n9462) );
  NANDN U10108 ( .A(n9462), .B(n37068), .Z(n9184) );
  NANDN U10109 ( .A(n9182), .B(n37069), .Z(n9183) );
  NAND U10110 ( .A(n9184), .B(n9183), .Z(n9366) );
  XNOR U10111 ( .A(b[45]), .B(a[16]), .Z(n9465) );
  NANDN U10112 ( .A(n9465), .B(n37261), .Z(n9187) );
  NANDN U10113 ( .A(n9185), .B(n37262), .Z(n9186) );
  AND U10114 ( .A(n9187), .B(n9186), .Z(n9367) );
  XNOR U10115 ( .A(n9366), .B(n9367), .Z(n9368) );
  XNOR U10116 ( .A(n9369), .B(n9368), .Z(n9526) );
  XNOR U10117 ( .A(b[35]), .B(a[26]), .Z(n9456) );
  NANDN U10118 ( .A(n9456), .B(n35985), .Z(n9190) );
  NANDN U10119 ( .A(n9188), .B(n35986), .Z(n9189) );
  NAND U10120 ( .A(n9190), .B(n9189), .Z(n9501) );
  XOR U10121 ( .A(b[53]), .B(n11986), .Z(n9453) );
  NANDN U10122 ( .A(n9453), .B(n37940), .Z(n9193) );
  NANDN U10123 ( .A(n9191), .B(n37941), .Z(n9192) );
  NAND U10124 ( .A(n9193), .B(n9192), .Z(n9498) );
  XOR U10125 ( .A(b[5]), .B(n25860), .Z(n9441) );
  OR U10126 ( .A(n9441), .B(n29363), .Z(n9196) );
  NANDN U10127 ( .A(n9194), .B(n29864), .Z(n9195) );
  AND U10128 ( .A(n9196), .B(n9195), .Z(n9499) );
  XNOR U10129 ( .A(n9498), .B(n9499), .Z(n9500) );
  XOR U10130 ( .A(n9501), .B(n9500), .Z(n9527) );
  XNOR U10131 ( .A(n9526), .B(n9527), .Z(n9528) );
  NANDN U10132 ( .A(n9198), .B(n9197), .Z(n9202) );
  NAND U10133 ( .A(n9200), .B(n9199), .Z(n9201) );
  AND U10134 ( .A(n9202), .B(n9201), .Z(n9529) );
  XNOR U10135 ( .A(n9528), .B(n9529), .Z(n9411) );
  NANDN U10136 ( .A(n9204), .B(n9203), .Z(n9208) );
  NAND U10137 ( .A(n9206), .B(n9205), .Z(n9207) );
  AND U10138 ( .A(n9208), .B(n9207), .Z(n9410) );
  XNOR U10139 ( .A(n9411), .B(n9410), .Z(n9412) );
  XOR U10140 ( .A(n9413), .B(n9412), .Z(n9571) );
  XOR U10141 ( .A(n9572), .B(n9571), .Z(n9346) );
  NANDN U10142 ( .A(n9210), .B(n9209), .Z(n9214) );
  OR U10143 ( .A(n9212), .B(n9211), .Z(n9213) );
  NAND U10144 ( .A(n9214), .B(n9213), .Z(n9344) );
  NANDN U10145 ( .A(n9216), .B(n9215), .Z(n9220) );
  OR U10146 ( .A(n9218), .B(n9217), .Z(n9219) );
  AND U10147 ( .A(n9220), .B(n9219), .Z(n9343) );
  XNOR U10148 ( .A(n9344), .B(n9343), .Z(n9345) );
  XNOR U10149 ( .A(n9346), .B(n9345), .Z(n9516) );
  XNOR U10150 ( .A(n9517), .B(n9516), .Z(n9519) );
  XNOR U10151 ( .A(n9518), .B(n9519), .Z(n9337) );
  NANDN U10152 ( .A(n9222), .B(n9221), .Z(n9226) );
  NANDN U10153 ( .A(n9224), .B(n9223), .Z(n9225) );
  AND U10154 ( .A(n9226), .B(n9225), .Z(n9338) );
  XOR U10155 ( .A(n9337), .B(n9338), .Z(n9339) );
  XNOR U10156 ( .A(n9340), .B(n9339), .Z(n9328) );
  NAND U10157 ( .A(n9228), .B(n9227), .Z(n9232) );
  NANDN U10158 ( .A(n9230), .B(n9229), .Z(n9231) );
  NAND U10159 ( .A(n9232), .B(n9231), .Z(n9333) );
  NANDN U10160 ( .A(n9234), .B(n9233), .Z(n9238) );
  NAND U10161 ( .A(n9236), .B(n9235), .Z(n9237) );
  NAND U10162 ( .A(n9238), .B(n9237), .Z(n9332) );
  OR U10163 ( .A(n9240), .B(n9239), .Z(n9244) );
  NANDN U10164 ( .A(n9242), .B(n9241), .Z(n9243) );
  NAND U10165 ( .A(n9244), .B(n9243), .Z(n9563) );
  NANDN U10166 ( .A(n9246), .B(n9245), .Z(n9250) );
  NANDN U10167 ( .A(n9248), .B(n9247), .Z(n9249) );
  NAND U10168 ( .A(n9250), .B(n9249), .Z(n9564) );
  XNOR U10169 ( .A(n9563), .B(n9564), .Z(n9565) );
  NANDN U10170 ( .A(n9252), .B(n9251), .Z(n9256) );
  NAND U10171 ( .A(n9254), .B(n9253), .Z(n9255) );
  NAND U10172 ( .A(n9256), .B(n9255), .Z(n9398) );
  XOR U10173 ( .A(b[31]), .B(n18804), .Z(n9382) );
  NANDN U10174 ( .A(n9382), .B(n35313), .Z(n9259) );
  NAND U10175 ( .A(n9257), .B(n35311), .Z(n9258) );
  NAND U10176 ( .A(n9259), .B(n9258), .Z(n9507) );
  XOR U10177 ( .A(n967), .B(n26347), .Z(n9391) );
  NAND U10178 ( .A(n9391), .B(n28939), .Z(n9262) );
  NAND U10179 ( .A(n28938), .B(n9260), .Z(n9261) );
  NAND U10180 ( .A(n9262), .B(n9261), .Z(n9504) );
  XOR U10181 ( .A(b[55]), .B(n11406), .Z(n9477) );
  NANDN U10182 ( .A(n9477), .B(n38075), .Z(n9265) );
  NANDN U10183 ( .A(n9263), .B(n38073), .Z(n9264) );
  AND U10184 ( .A(n9265), .B(n9264), .Z(n9505) );
  XNOR U10185 ( .A(n9504), .B(n9505), .Z(n9506) );
  XOR U10186 ( .A(n9507), .B(n9506), .Z(n9399) );
  XNOR U10187 ( .A(n9398), .B(n9399), .Z(n9400) );
  NAND U10188 ( .A(n34044), .B(n9266), .Z(n9268) );
  XOR U10189 ( .A(n34510), .B(n20686), .Z(n9483) );
  NANDN U10190 ( .A(n33867), .B(n9483), .Z(n9267) );
  NAND U10191 ( .A(n9268), .B(n9267), .Z(n9447) );
  XNOR U10192 ( .A(b[25]), .B(n19980), .Z(n9548) );
  NANDN U10193 ( .A(n34219), .B(n9548), .Z(n9271) );
  NAND U10194 ( .A(n34217), .B(n9269), .Z(n9270) );
  NAND U10195 ( .A(n9271), .B(n9270), .Z(n9444) );
  NAND U10196 ( .A(n9272), .B(n34848), .Z(n9274) );
  XOR U10197 ( .A(n35375), .B(n19513), .Z(n9435) );
  NAND U10198 ( .A(n34618), .B(n9435), .Z(n9273) );
  AND U10199 ( .A(n9274), .B(n9273), .Z(n9445) );
  XNOR U10200 ( .A(n9444), .B(n9445), .Z(n9446) );
  XNOR U10201 ( .A(n9447), .B(n9446), .Z(n9363) );
  NANDN U10202 ( .A(n9275), .B(n33283), .Z(n9277) );
  XNOR U10203 ( .A(n33020), .B(a[42]), .Z(n9545) );
  NANDN U10204 ( .A(n33021), .B(n9545), .Z(n9276) );
  NAND U10205 ( .A(n9277), .B(n9276), .Z(n9361) );
  XNOR U10206 ( .A(b[21]), .B(a[40]), .Z(n9554) );
  OR U10207 ( .A(n9554), .B(n33634), .Z(n9280) );
  NANDN U10208 ( .A(n9278), .B(n33464), .Z(n9279) );
  AND U10209 ( .A(n9280), .B(n9279), .Z(n9360) );
  XNOR U10210 ( .A(n9361), .B(n9360), .Z(n9362) );
  XOR U10211 ( .A(n9363), .B(n9362), .Z(n9401) );
  XOR U10212 ( .A(n9400), .B(n9401), .Z(n9566) );
  XOR U10213 ( .A(n9565), .B(n9566), .Z(n9331) );
  XNOR U10214 ( .A(n9332), .B(n9331), .Z(n9334) );
  XNOR U10215 ( .A(n9333), .B(n9334), .Z(n9325) );
  NANDN U10216 ( .A(n9282), .B(n9281), .Z(n9286) );
  NAND U10217 ( .A(n9284), .B(n9283), .Z(n9285) );
  AND U10218 ( .A(n9286), .B(n9285), .Z(n9326) );
  XOR U10219 ( .A(n9325), .B(n9326), .Z(n9327) );
  XOR U10220 ( .A(n9328), .B(n9327), .Z(n9322) );
  NAND U10221 ( .A(n9288), .B(n9287), .Z(n9292) );
  NANDN U10222 ( .A(n9290), .B(n9289), .Z(n9291) );
  NAND U10223 ( .A(n9292), .B(n9291), .Z(n9320) );
  XNOR U10224 ( .A(n9320), .B(n9319), .Z(n9321) );
  XNOR U10225 ( .A(n9322), .B(n9321), .Z(n9315) );
  OR U10226 ( .A(n9298), .B(n9297), .Z(n9302) );
  NANDN U10227 ( .A(n9300), .B(n9299), .Z(n9301) );
  AND U10228 ( .A(n9302), .B(n9301), .Z(n9316) );
  XOR U10229 ( .A(n9315), .B(n9316), .Z(n9317) );
  XNOR U10230 ( .A(n9318), .B(n9317), .Z(n9309) );
  NANDN U10231 ( .A(n9304), .B(n9303), .Z(n9308) );
  NANDN U10232 ( .A(n9306), .B(n9305), .Z(n9307) );
  NAND U10233 ( .A(n9308), .B(n9307), .Z(n9310) );
  XNOR U10234 ( .A(n9309), .B(n9310), .Z(n9311) );
  XOR U10235 ( .A(n9312), .B(n9311), .Z(n9574) );
  XOR U10236 ( .A(n9575), .B(n9574), .Z(c[124]) );
  NANDN U10237 ( .A(n9310), .B(n9309), .Z(n9314) );
  NAND U10238 ( .A(n9312), .B(n9311), .Z(n9313) );
  NAND U10239 ( .A(n9314), .B(n9313), .Z(n9586) );
  NANDN U10240 ( .A(n9320), .B(n9319), .Z(n9324) );
  NANDN U10241 ( .A(n9322), .B(n9321), .Z(n9323) );
  NAND U10242 ( .A(n9324), .B(n9323), .Z(n9592) );
  NAND U10243 ( .A(n9326), .B(n9325), .Z(n9330) );
  NAND U10244 ( .A(n9328), .B(n9327), .Z(n9329) );
  NAND U10245 ( .A(n9330), .B(n9329), .Z(n9590) );
  NAND U10246 ( .A(n9332), .B(n9331), .Z(n9336) );
  NANDN U10247 ( .A(n9334), .B(n9333), .Z(n9335) );
  NAND U10248 ( .A(n9336), .B(n9335), .Z(n9595) );
  NAND U10249 ( .A(n9338), .B(n9337), .Z(n9342) );
  NAND U10250 ( .A(n9340), .B(n9339), .Z(n9341) );
  NAND U10251 ( .A(n9342), .B(n9341), .Z(n9596) );
  XNOR U10252 ( .A(n9595), .B(n9596), .Z(n9597) );
  NANDN U10253 ( .A(n9344), .B(n9343), .Z(n9348) );
  NANDN U10254 ( .A(n9346), .B(n9345), .Z(n9347) );
  NAND U10255 ( .A(n9348), .B(n9347), .Z(n9614) );
  NANDN U10256 ( .A(n9350), .B(n9349), .Z(n9354) );
  NAND U10257 ( .A(n9352), .B(n9351), .Z(n9353) );
  NAND U10258 ( .A(n9354), .B(n9353), .Z(n9641) );
  NANDN U10259 ( .A(n9356), .B(n9355), .Z(n9359) );
  NANDN U10260 ( .A(n9357), .B(n9381), .Z(n9358) );
  AND U10261 ( .A(n9359), .B(n9358), .Z(n9642) );
  XNOR U10262 ( .A(n9641), .B(n9642), .Z(n9643) );
  NANDN U10263 ( .A(n9361), .B(n9360), .Z(n9365) );
  NAND U10264 ( .A(n9363), .B(n9362), .Z(n9364) );
  NAND U10265 ( .A(n9365), .B(n9364), .Z(n9644) );
  XOR U10266 ( .A(n9643), .B(n9644), .Z(n9782) );
  NANDN U10267 ( .A(n9367), .B(n9366), .Z(n9371) );
  NAND U10268 ( .A(n9369), .B(n9368), .Z(n9370) );
  NAND U10269 ( .A(n9371), .B(n9370), .Z(n9772) );
  NAND U10270 ( .A(n9372), .B(n38326), .Z(n9374) );
  XOR U10271 ( .A(b[59]), .B(n10524), .Z(n9666) );
  OR U10272 ( .A(n9666), .B(n38273), .Z(n9373) );
  NAND U10273 ( .A(n9374), .B(n9373), .Z(n9841) );
  IV U10274 ( .A(n9375), .Z(n38371) );
  XOR U10275 ( .A(b[61]), .B(n10457), .Z(n9705) );
  NOR U10276 ( .A(n38371), .B(n9705), .Z(n9380) );
  XNOR U10277 ( .A(n984), .B(a[0]), .Z(n9378) );
  XNOR U10278 ( .A(n984), .B(b[59]), .Z(n9377) );
  XNOR U10279 ( .A(n984), .B(b[60]), .Z(n9376) );
  AND U10280 ( .A(n9377), .B(n9376), .Z(n38369) );
  NAND U10281 ( .A(n9378), .B(n38369), .Z(n9379) );
  NANDN U10282 ( .A(n9380), .B(n9379), .Z(n9840) );
  XNOR U10283 ( .A(n9841), .B(n9840), .Z(n9714) );
  NANDN U10284 ( .A(n38400), .B(b[60]), .Z(n38399) );
  AND U10285 ( .A(n38399), .B(b[61]), .Z(n38440) );
  NANDN U10286 ( .A(n9381), .B(n38440), .Z(n9711) );
  NANDN U10287 ( .A(n9382), .B(n35311), .Z(n9384) );
  XNOR U10288 ( .A(n973), .B(a[31]), .Z(n9828) );
  NAND U10289 ( .A(n9828), .B(n35313), .Z(n9383) );
  NAND U10290 ( .A(n9384), .B(n9383), .Z(n9712) );
  XNOR U10291 ( .A(n9711), .B(n9712), .Z(n9713) );
  XOR U10292 ( .A(n9714), .B(n9713), .Z(n9770) );
  NAND U10293 ( .A(n9385), .B(n35188), .Z(n9387) );
  XNOR U10294 ( .A(n35540), .B(a[33]), .Z(n9672) );
  NANDN U10295 ( .A(n34968), .B(n9672), .Z(n9386) );
  NAND U10296 ( .A(n9387), .B(n9386), .Z(n9823) );
  NANDN U10297 ( .A(n966), .B(a[61]), .Z(n9388) );
  XOR U10298 ( .A(n29232), .B(n9388), .Z(n9390) );
  IV U10299 ( .A(a[60]), .Z(n27436) );
  NANDN U10300 ( .A(n27436), .B(n966), .Z(n9389) );
  AND U10301 ( .A(n9390), .B(n9389), .Z(n9821) );
  XNOR U10302 ( .A(b[3]), .B(a[59]), .Z(n9845) );
  NANDN U10303 ( .A(n9845), .B(n28939), .Z(n9393) );
  NAND U10304 ( .A(n28938), .B(n9391), .Z(n9392) );
  AND U10305 ( .A(n9393), .B(n9392), .Z(n9822) );
  XOR U10306 ( .A(n9821), .B(n9822), .Z(n9824) );
  XNOR U10307 ( .A(n9823), .B(n9824), .Z(n9769) );
  XNOR U10308 ( .A(n9770), .B(n9769), .Z(n9771) );
  XNOR U10309 ( .A(n9772), .B(n9771), .Z(n9779) );
  XNOR U10310 ( .A(n9779), .B(n9780), .Z(n9781) );
  XNOR U10311 ( .A(n9782), .B(n9781), .Z(n9626) );
  NANDN U10312 ( .A(n9399), .B(n9398), .Z(n9403) );
  NAND U10313 ( .A(n9401), .B(n9400), .Z(n9402) );
  NAND U10314 ( .A(n9403), .B(n9402), .Z(n9623) );
  NANDN U10315 ( .A(n9405), .B(n9404), .Z(n9409) );
  NANDN U10316 ( .A(n9407), .B(n9406), .Z(n9408) );
  NAND U10317 ( .A(n9409), .B(n9408), .Z(n9624) );
  XNOR U10318 ( .A(n9623), .B(n9624), .Z(n9625) );
  XOR U10319 ( .A(n9626), .B(n9625), .Z(n9620) );
  NANDN U10320 ( .A(n9411), .B(n9410), .Z(n9415) );
  NAND U10321 ( .A(n9413), .B(n9412), .Z(n9414) );
  NAND U10322 ( .A(n9415), .B(n9414), .Z(n9618) );
  NANDN U10323 ( .A(n9421), .B(n9420), .Z(n9425) );
  NAND U10324 ( .A(n9423), .B(n9422), .Z(n9424) );
  AND U10325 ( .A(n9425), .B(n9424), .Z(n9774) );
  XNOR U10326 ( .A(n9773), .B(n9774), .Z(n9775) );
  XOR U10327 ( .A(b[39]), .B(n16269), .Z(n9721) );
  NANDN U10328 ( .A(n9721), .B(n36553), .Z(n9428) );
  NANDN U10329 ( .A(n9426), .B(n36643), .Z(n9427) );
  NAND U10330 ( .A(n9428), .B(n9427), .Z(n9742) );
  XOR U10331 ( .A(b[11]), .B(n24288), .Z(n9724) );
  OR U10332 ( .A(n9724), .B(n31369), .Z(n9431) );
  NANDN U10333 ( .A(n9429), .B(n31119), .Z(n9430) );
  NAND U10334 ( .A(n9431), .B(n9430), .Z(n9739) );
  XOR U10335 ( .A(b[9]), .B(n25001), .Z(n9727) );
  NANDN U10336 ( .A(n9727), .B(n30509), .Z(n9434) );
  NANDN U10337 ( .A(n9432), .B(n30846), .Z(n9433) );
  AND U10338 ( .A(n9434), .B(n9433), .Z(n9740) );
  XNOR U10339 ( .A(n9739), .B(n9740), .Z(n9741) );
  XNOR U10340 ( .A(n9742), .B(n9741), .Z(n9791) );
  NAND U10341 ( .A(n34848), .B(n9435), .Z(n9437) );
  XOR U10342 ( .A(n35375), .B(n20315), .Z(n9669) );
  NAND U10343 ( .A(n34618), .B(n9669), .Z(n9436) );
  NAND U10344 ( .A(n9437), .B(n9436), .Z(n9718) );
  XOR U10345 ( .A(n31123), .B(n25466), .Z(n9812) );
  NAND U10346 ( .A(n9812), .B(n29949), .Z(n9440) );
  NAND U10347 ( .A(n29948), .B(n9438), .Z(n9439) );
  NAND U10348 ( .A(n9440), .B(n9439), .Z(n9715) );
  XOR U10349 ( .A(b[5]), .B(n26122), .Z(n9708) );
  OR U10350 ( .A(n9708), .B(n29363), .Z(n9443) );
  NANDN U10351 ( .A(n9441), .B(n29864), .Z(n9442) );
  AND U10352 ( .A(n9443), .B(n9442), .Z(n9716) );
  XNOR U10353 ( .A(n9715), .B(n9716), .Z(n9717) );
  XOR U10354 ( .A(n9718), .B(n9717), .Z(n9792) );
  XNOR U10355 ( .A(n9791), .B(n9792), .Z(n9793) );
  NANDN U10356 ( .A(n9445), .B(n9444), .Z(n9449) );
  NAND U10357 ( .A(n9447), .B(n9446), .Z(n9448) );
  AND U10358 ( .A(n9449), .B(n9448), .Z(n9794) );
  XNOR U10359 ( .A(n9793), .B(n9794), .Z(n9691) );
  XOR U10360 ( .A(b[51]), .B(n12830), .Z(n9730) );
  NANDN U10361 ( .A(n9730), .B(n37803), .Z(n9452) );
  NANDN U10362 ( .A(n9450), .B(n37802), .Z(n9451) );
  NAND U10363 ( .A(n9452), .B(n9451), .Z(n9687) );
  XOR U10364 ( .A(b[53]), .B(n12258), .Z(n9757) );
  NANDN U10365 ( .A(n9757), .B(n37940), .Z(n9455) );
  NANDN U10366 ( .A(n9453), .B(n37941), .Z(n9454) );
  NAND U10367 ( .A(n9455), .B(n9454), .Z(n9684) );
  XNOR U10368 ( .A(b[35]), .B(a[27]), .Z(n9702) );
  NANDN U10369 ( .A(n9702), .B(n35985), .Z(n9458) );
  NANDN U10370 ( .A(n9456), .B(n35986), .Z(n9457) );
  AND U10371 ( .A(n9458), .B(n9457), .Z(n9685) );
  XNOR U10372 ( .A(n9684), .B(n9685), .Z(n9686) );
  XNOR U10373 ( .A(n9687), .B(n9686), .Z(n9785) );
  XOR U10374 ( .A(b[13]), .B(n23852), .Z(n9736) );
  OR U10375 ( .A(n9736), .B(n31550), .Z(n9461) );
  NANDN U10376 ( .A(n9459), .B(n31874), .Z(n9460) );
  NAND U10377 ( .A(n9461), .B(n9460), .Z(n9766) );
  XOR U10378 ( .A(b[43]), .B(n15113), .Z(n9754) );
  NANDN U10379 ( .A(n9754), .B(n37068), .Z(n9464) );
  NANDN U10380 ( .A(n9462), .B(n37069), .Z(n9463) );
  NAND U10381 ( .A(n9464), .B(n9463), .Z(n9763) );
  XNOR U10382 ( .A(b[45]), .B(a[17]), .Z(n9751) );
  NANDN U10383 ( .A(n9751), .B(n37261), .Z(n9467) );
  NANDN U10384 ( .A(n9465), .B(n37262), .Z(n9466) );
  AND U10385 ( .A(n9467), .B(n9466), .Z(n9764) );
  XNOR U10386 ( .A(n9763), .B(n9764), .Z(n9765) );
  XOR U10387 ( .A(n9766), .B(n9765), .Z(n9786) );
  XOR U10388 ( .A(n9785), .B(n9786), .Z(n9788) );
  NANDN U10389 ( .A(n9469), .B(n9468), .Z(n9473) );
  NAND U10390 ( .A(n9471), .B(n9470), .Z(n9472) );
  NAND U10391 ( .A(n9473), .B(n9472), .Z(n9787) );
  XNOR U10392 ( .A(n9788), .B(n9787), .Z(n9690) );
  XOR U10393 ( .A(n9691), .B(n9690), .Z(n9692) );
  XOR U10394 ( .A(b[33]), .B(n18003), .Z(n9842) );
  NANDN U10395 ( .A(n9842), .B(n35620), .Z(n9476) );
  NAND U10396 ( .A(n9474), .B(n35621), .Z(n9475) );
  NAND U10397 ( .A(n9476), .B(n9475), .Z(n9681) );
  XOR U10398 ( .A(b[55]), .B(n11694), .Z(n9760) );
  NANDN U10399 ( .A(n9760), .B(n38075), .Z(n9479) );
  NANDN U10400 ( .A(n9477), .B(n38073), .Z(n9478) );
  NAND U10401 ( .A(n9479), .B(n9478), .Z(n9678) );
  XOR U10402 ( .A(b[57]), .B(n11202), .Z(n9809) );
  OR U10403 ( .A(n9809), .B(n965), .Z(n9482) );
  NANDN U10404 ( .A(n9480), .B(n38194), .Z(n9481) );
  AND U10405 ( .A(n9482), .B(n9481), .Z(n9679) );
  XNOR U10406 ( .A(n9678), .B(n9679), .Z(n9680) );
  XNOR U10407 ( .A(n9681), .B(n9680), .Z(n9696) );
  NAND U10408 ( .A(n34044), .B(n9483), .Z(n9485) );
  XOR U10409 ( .A(n34510), .B(n20867), .Z(n9831) );
  NANDN U10410 ( .A(n33867), .B(n9831), .Z(n9484) );
  NAND U10411 ( .A(n9485), .B(n9484), .Z(n9818) );
  NAND U10412 ( .A(n37469), .B(n9486), .Z(n9488) );
  XOR U10413 ( .A(n978), .B(n13976), .Z(n9800) );
  NAND U10414 ( .A(n9800), .B(n37471), .Z(n9487) );
  NAND U10415 ( .A(n9488), .B(n9487), .Z(n9815) );
  XOR U10416 ( .A(b[49]), .B(n13509), .Z(n9803) );
  OR U10417 ( .A(n9803), .B(n37756), .Z(n9491) );
  NANDN U10418 ( .A(n9489), .B(n37652), .Z(n9490) );
  AND U10419 ( .A(n9491), .B(n9490), .Z(n9816) );
  XNOR U10420 ( .A(n9815), .B(n9816), .Z(n9817) );
  XOR U10421 ( .A(n9818), .B(n9817), .Z(n9697) );
  XOR U10422 ( .A(n9696), .B(n9697), .Z(n9699) );
  NANDN U10423 ( .A(n9493), .B(n9492), .Z(n9497) );
  NAND U10424 ( .A(n9495), .B(n9494), .Z(n9496) );
  NAND U10425 ( .A(n9497), .B(n9496), .Z(n9698) );
  XNOR U10426 ( .A(n9699), .B(n9698), .Z(n9654) );
  NANDN U10427 ( .A(n9499), .B(n9498), .Z(n9503) );
  NAND U10428 ( .A(n9501), .B(n9500), .Z(n9502) );
  NAND U10429 ( .A(n9503), .B(n9502), .Z(n9651) );
  NANDN U10430 ( .A(n9505), .B(n9504), .Z(n9509) );
  NAND U10431 ( .A(n9507), .B(n9506), .Z(n9508) );
  AND U10432 ( .A(n9509), .B(n9508), .Z(n9652) );
  XNOR U10433 ( .A(n9651), .B(n9652), .Z(n9653) );
  XOR U10434 ( .A(n9654), .B(n9653), .Z(n9693) );
  XOR U10435 ( .A(n9692), .B(n9693), .Z(n9776) );
  XNOR U10436 ( .A(n9775), .B(n9776), .Z(n9617) );
  XNOR U10437 ( .A(n9618), .B(n9617), .Z(n9619) );
  XNOR U10438 ( .A(n9620), .B(n9619), .Z(n9611) );
  NANDN U10439 ( .A(n9511), .B(n9510), .Z(n9515) );
  NAND U10440 ( .A(n9513), .B(n9512), .Z(n9514) );
  NAND U10441 ( .A(n9515), .B(n9514), .Z(n9612) );
  XNOR U10442 ( .A(n9611), .B(n9612), .Z(n9613) );
  XNOR U10443 ( .A(n9614), .B(n9613), .Z(n9604) );
  NANDN U10444 ( .A(n9521), .B(n9520), .Z(n9525) );
  NAND U10445 ( .A(n9523), .B(n9522), .Z(n9524) );
  NAND U10446 ( .A(n9525), .B(n9524), .Z(n9631) );
  NANDN U10447 ( .A(n9527), .B(n9526), .Z(n9531) );
  NAND U10448 ( .A(n9529), .B(n9528), .Z(n9530) );
  NAND U10449 ( .A(n9531), .B(n9530), .Z(n9630) );
  XOR U10450 ( .A(b[15]), .B(n23149), .Z(n9733) );
  OR U10451 ( .A(n9733), .B(n32010), .Z(n9538) );
  NANDN U10452 ( .A(n9536), .B(n32011), .Z(n9537) );
  NAND U10453 ( .A(n9538), .B(n9537), .Z(n9660) );
  XNOR U10454 ( .A(b[17]), .B(a[45]), .Z(n9797) );
  NANDN U10455 ( .A(n9797), .B(n32543), .Z(n9541) );
  NANDN U10456 ( .A(n9539), .B(n32541), .Z(n9540) );
  NAND U10457 ( .A(n9541), .B(n9540), .Z(n9657) );
  XNOR U10458 ( .A(b[41]), .B(a[21]), .Z(n9748) );
  OR U10459 ( .A(n9748), .B(n36905), .Z(n9544) );
  NANDN U10460 ( .A(n9542), .B(n36807), .Z(n9543) );
  AND U10461 ( .A(n9544), .B(n9543), .Z(n9658) );
  XNOR U10462 ( .A(n9657), .B(n9658), .Z(n9659) );
  XNOR U10463 ( .A(n9660), .B(n9659), .Z(n9650) );
  NAND U10464 ( .A(n9545), .B(n33283), .Z(n9547) );
  XOR U10465 ( .A(n33020), .B(n21996), .Z(n9745) );
  NANDN U10466 ( .A(n33021), .B(n9745), .Z(n9546) );
  NAND U10467 ( .A(n9547), .B(n9546), .Z(n9837) );
  XNOR U10468 ( .A(b[25]), .B(n20352), .Z(n9675) );
  NANDN U10469 ( .A(n34219), .B(n9675), .Z(n9550) );
  NAND U10470 ( .A(n34217), .B(n9548), .Z(n9549) );
  NAND U10471 ( .A(n9550), .B(n9549), .Z(n9834) );
  XOR U10472 ( .A(b[37]), .B(n16916), .Z(n9806) );
  NANDN U10473 ( .A(n9806), .B(n36311), .Z(n9553) );
  NANDN U10474 ( .A(n9551), .B(n36309), .Z(n9552) );
  AND U10475 ( .A(n9553), .B(n9552), .Z(n9835) );
  XNOR U10476 ( .A(n9834), .B(n9835), .Z(n9836) );
  XNOR U10477 ( .A(n9837), .B(n9836), .Z(n9647) );
  XNOR U10478 ( .A(b[21]), .B(n21441), .Z(n9825) );
  NANDN U10479 ( .A(n33634), .B(n9825), .Z(n9556) );
  NANDN U10480 ( .A(n9554), .B(n33464), .Z(n9555) );
  NAND U10481 ( .A(n9556), .B(n9555), .Z(n9648) );
  XNOR U10482 ( .A(n9647), .B(n9648), .Z(n9649) );
  XOR U10483 ( .A(n9650), .B(n9649), .Z(n9635) );
  NANDN U10484 ( .A(n9558), .B(n9557), .Z(n9562) );
  NAND U10485 ( .A(n9560), .B(n9559), .Z(n9561) );
  AND U10486 ( .A(n9562), .B(n9561), .Z(n9636) );
  XNOR U10487 ( .A(n9635), .B(n9636), .Z(n9638) );
  XNOR U10488 ( .A(n9637), .B(n9638), .Z(n9629) );
  XNOR U10489 ( .A(n9630), .B(n9629), .Z(n9632) );
  XNOR U10490 ( .A(n9631), .B(n9632), .Z(n9607) );
  NANDN U10491 ( .A(n9564), .B(n9563), .Z(n9568) );
  NAND U10492 ( .A(n9566), .B(n9565), .Z(n9567) );
  NAND U10493 ( .A(n9568), .B(n9567), .Z(n9605) );
  XNOR U10494 ( .A(n9605), .B(n9606), .Z(n9608) );
  XOR U10495 ( .A(n9607), .B(n9608), .Z(n9601) );
  XNOR U10496 ( .A(n9602), .B(n9601), .Z(n9603) );
  XOR U10497 ( .A(n9604), .B(n9603), .Z(n9598) );
  XOR U10498 ( .A(n9597), .B(n9598), .Z(n9589) );
  XOR U10499 ( .A(n9590), .B(n9589), .Z(n9591) );
  XOR U10500 ( .A(n9592), .B(n9591), .Z(n9584) );
  XOR U10501 ( .A(n9583), .B(n9584), .Z(n9585) );
  XNOR U10502 ( .A(n9586), .B(n9585), .Z(n9578) );
  XNOR U10503 ( .A(n9578), .B(sreg[125]), .Z(n9580) );
  NAND U10504 ( .A(n9573), .B(sreg[124]), .Z(n9577) );
  OR U10505 ( .A(n9575), .B(n9574), .Z(n9576) );
  AND U10506 ( .A(n9577), .B(n9576), .Z(n9579) );
  XOR U10507 ( .A(n9580), .B(n9579), .Z(c[125]) );
  NAND U10508 ( .A(n9578), .B(sreg[125]), .Z(n9582) );
  OR U10509 ( .A(n9580), .B(n9579), .Z(n9581) );
  NAND U10510 ( .A(n9582), .B(n9581), .Z(n10130) );
  XNOR U10511 ( .A(n10130), .B(sreg[126]), .Z(n10132) );
  OR U10512 ( .A(n9584), .B(n9583), .Z(n9588) );
  NAND U10513 ( .A(n9586), .B(n9585), .Z(n9587) );
  NAND U10514 ( .A(n9588), .B(n9587), .Z(n9851) );
  NAND U10515 ( .A(n9590), .B(n9589), .Z(n9594) );
  NANDN U10516 ( .A(n9592), .B(n9591), .Z(n9593) );
  NAND U10517 ( .A(n9594), .B(n9593), .Z(n9849) );
  NANDN U10518 ( .A(n9596), .B(n9595), .Z(n9600) );
  NAND U10519 ( .A(n9598), .B(n9597), .Z(n9599) );
  NAND U10520 ( .A(n9600), .B(n9599), .Z(n9856) );
  NANDN U10521 ( .A(n9606), .B(n9605), .Z(n9610) );
  NAND U10522 ( .A(n9608), .B(n9607), .Z(n9609) );
  NAND U10523 ( .A(n9610), .B(n9609), .Z(n9866) );
  NANDN U10524 ( .A(n9612), .B(n9611), .Z(n9616) );
  NAND U10525 ( .A(n9614), .B(n9613), .Z(n9615) );
  NAND U10526 ( .A(n9616), .B(n9615), .Z(n9867) );
  XNOR U10527 ( .A(n9866), .B(n9867), .Z(n9868) );
  NAND U10528 ( .A(n9618), .B(n9617), .Z(n9622) );
  OR U10529 ( .A(n9620), .B(n9619), .Z(n9621) );
  NAND U10530 ( .A(n9622), .B(n9621), .Z(n9861) );
  NANDN U10531 ( .A(n9624), .B(n9623), .Z(n9628) );
  NANDN U10532 ( .A(n9626), .B(n9625), .Z(n9627) );
  NAND U10533 ( .A(n9628), .B(n9627), .Z(n10036) );
  NAND U10534 ( .A(n9630), .B(n9629), .Z(n9634) );
  NANDN U10535 ( .A(n9632), .B(n9631), .Z(n9633) );
  AND U10536 ( .A(n9634), .B(n9633), .Z(n10037) );
  XNOR U10537 ( .A(n10036), .B(n10037), .Z(n10038) );
  NAND U10538 ( .A(n9636), .B(n9635), .Z(n9640) );
  NANDN U10539 ( .A(n9638), .B(n9637), .Z(n9639) );
  NAND U10540 ( .A(n9640), .B(n9639), .Z(n10030) );
  NANDN U10541 ( .A(n9642), .B(n9641), .Z(n9646) );
  NANDN U10542 ( .A(n9644), .B(n9643), .Z(n9645) );
  NAND U10543 ( .A(n9646), .B(n9645), .Z(n10031) );
  XNOR U10544 ( .A(n10030), .B(n10031), .Z(n10032) );
  NANDN U10545 ( .A(n9652), .B(n9651), .Z(n9656) );
  NAND U10546 ( .A(n9654), .B(n9653), .Z(n9655) );
  NAND U10547 ( .A(n9656), .B(n9655), .Z(n10049) );
  XNOR U10548 ( .A(n10048), .B(n10049), .Z(n10050) );
  NANDN U10549 ( .A(n9658), .B(n9657), .Z(n9662) );
  NAND U10550 ( .A(n9660), .B(n9659), .Z(n9661) );
  NAND U10551 ( .A(n9662), .B(n9661), .Z(n10016) );
  NANDN U10552 ( .A(n966), .B(a[62]), .Z(n9663) );
  XOR U10553 ( .A(n29232), .B(n9663), .Z(n9665) );
  IV U10554 ( .A(a[61]), .Z(n27773) );
  NANDN U10555 ( .A(n27773), .B(n966), .Z(n9664) );
  AND U10556 ( .A(n9665), .B(n9664), .Z(n10097) );
  NANDN U10557 ( .A(n9666), .B(n38326), .Z(n9668) );
  XOR U10558 ( .A(n38400), .B(n10854), .Z(n10094) );
  NANDN U10559 ( .A(n38273), .B(n10094), .Z(n9667) );
  AND U10560 ( .A(n9668), .B(n9667), .Z(n10098) );
  XOR U10561 ( .A(n10097), .B(n10098), .Z(n10100) );
  IV U10562 ( .A(b[62]), .Z(n38433) );
  XOR U10563 ( .A(n38433), .B(n984), .Z(n38422) );
  NANDN U10564 ( .A(n986), .B(n38422), .Z(n10099) );
  XOR U10565 ( .A(n10100), .B(n10099), .Z(n10014) );
  NAND U10566 ( .A(n34848), .B(n9669), .Z(n9671) );
  XOR U10567 ( .A(n35375), .B(n19980), .Z(n9950) );
  NAND U10568 ( .A(n34618), .B(n9950), .Z(n9670) );
  NAND U10569 ( .A(n9671), .B(n9670), .Z(n9983) );
  NAND U10570 ( .A(n9672), .B(n35188), .Z(n9674) );
  XOR U10571 ( .A(n35540), .B(n19513), .Z(n9878) );
  NANDN U10572 ( .A(n34968), .B(n9878), .Z(n9673) );
  NAND U10573 ( .A(n9674), .B(n9673), .Z(n9980) );
  XNOR U10574 ( .A(b[25]), .B(n20686), .Z(n10109) );
  NANDN U10575 ( .A(n34219), .B(n10109), .Z(n9677) );
  NAND U10576 ( .A(n34217), .B(n9675), .Z(n9676) );
  AND U10577 ( .A(n9677), .B(n9676), .Z(n9981) );
  XNOR U10578 ( .A(n9980), .B(n9981), .Z(n9982) );
  XNOR U10579 ( .A(n9983), .B(n9982), .Z(n10015) );
  XNOR U10580 ( .A(n10014), .B(n10015), .Z(n10017) );
  XNOR U10581 ( .A(n10016), .B(n10017), .Z(n10021) );
  NANDN U10582 ( .A(n9679), .B(n9678), .Z(n9683) );
  NAND U10583 ( .A(n9681), .B(n9680), .Z(n9682) );
  NAND U10584 ( .A(n9683), .B(n9682), .Z(n10019) );
  NANDN U10585 ( .A(n9685), .B(n9684), .Z(n9689) );
  NAND U10586 ( .A(n9687), .B(n9686), .Z(n9688) );
  AND U10587 ( .A(n9689), .B(n9688), .Z(n10018) );
  XNOR U10588 ( .A(n10019), .B(n10018), .Z(n10020) );
  XOR U10589 ( .A(n10021), .B(n10020), .Z(n10051) );
  XOR U10590 ( .A(n10050), .B(n10051), .Z(n10033) );
  XOR U10591 ( .A(n10032), .B(n10033), .Z(n10126) );
  OR U10592 ( .A(n9691), .B(n9690), .Z(n9695) );
  NANDN U10593 ( .A(n9693), .B(n9692), .Z(n9694) );
  NAND U10594 ( .A(n9695), .B(n9694), .Z(n10124) );
  NANDN U10595 ( .A(n9697), .B(n9696), .Z(n9701) );
  OR U10596 ( .A(n9699), .B(n9698), .Z(n9700) );
  NAND U10597 ( .A(n9701), .B(n9700), .Z(n10027) );
  XNOR U10598 ( .A(b[35]), .B(a[28]), .Z(n9965) );
  NANDN U10599 ( .A(n9965), .B(n35985), .Z(n9704) );
  NANDN U10600 ( .A(n9702), .B(n35986), .Z(n9703) );
  NAND U10601 ( .A(n9704), .B(n9703), .Z(n9947) );
  XOR U10602 ( .A(b[61]), .B(n10363), .Z(n10006) );
  OR U10603 ( .A(n10006), .B(n38371), .Z(n9707) );
  NANDN U10604 ( .A(n9705), .B(n38369), .Z(n9706) );
  NAND U10605 ( .A(n9707), .B(n9706), .Z(n9944) );
  XOR U10606 ( .A(b[5]), .B(n26347), .Z(n9932) );
  OR U10607 ( .A(n9932), .B(n29363), .Z(n9710) );
  NANDN U10608 ( .A(n9708), .B(n29864), .Z(n9709) );
  AND U10609 ( .A(n9710), .B(n9709), .Z(n9945) );
  XNOR U10610 ( .A(n9944), .B(n9945), .Z(n9946) );
  XNOR U10611 ( .A(n9947), .B(n9946), .Z(n10079) );
  NANDN U10612 ( .A(n9716), .B(n9715), .Z(n9720) );
  NAND U10613 ( .A(n9718), .B(n9717), .Z(n9719) );
  NAND U10614 ( .A(n9720), .B(n9719), .Z(n10077) );
  XNOR U10615 ( .A(n10076), .B(n10077), .Z(n10078) );
  XOR U10616 ( .A(n10079), .B(n10078), .Z(n10056) );
  XOR U10617 ( .A(b[39]), .B(n16508), .Z(n9992) );
  NANDN U10618 ( .A(n9992), .B(n36553), .Z(n9723) );
  NANDN U10619 ( .A(n9721), .B(n36643), .Z(n9722) );
  NAND U10620 ( .A(n9723), .B(n9722), .Z(n9905) );
  XOR U10621 ( .A(b[11]), .B(n25134), .Z(n9986) );
  OR U10622 ( .A(n9986), .B(n31369), .Z(n9726) );
  NANDN U10623 ( .A(n9724), .B(n31119), .Z(n9725) );
  NAND U10624 ( .A(n9726), .B(n9725), .Z(n9902) );
  XOR U10625 ( .A(b[9]), .B(n25177), .Z(n9920) );
  NANDN U10626 ( .A(n9920), .B(n30509), .Z(n9729) );
  NANDN U10627 ( .A(n9727), .B(n30846), .Z(n9728) );
  AND U10628 ( .A(n9729), .B(n9728), .Z(n9903) );
  XNOR U10629 ( .A(n9902), .B(n9903), .Z(n9904) );
  XNOR U10630 ( .A(n9905), .B(n9904), .Z(n10070) );
  XOR U10631 ( .A(b[51]), .B(n13106), .Z(n9959) );
  NANDN U10632 ( .A(n9959), .B(n37803), .Z(n9732) );
  NANDN U10633 ( .A(n9730), .B(n37802), .Z(n9731) );
  NAND U10634 ( .A(n9732), .B(n9731), .Z(n9890) );
  XOR U10635 ( .A(b[15]), .B(n23447), .Z(n10115) );
  OR U10636 ( .A(n10115), .B(n32010), .Z(n9735) );
  NANDN U10637 ( .A(n9733), .B(n32011), .Z(n9734) );
  NAND U10638 ( .A(n9735), .B(n9734), .Z(n9887) );
  XOR U10639 ( .A(n971), .B(n24671), .Z(n10112) );
  NANDN U10640 ( .A(n31550), .B(n10112), .Z(n9738) );
  NANDN U10641 ( .A(n9736), .B(n31874), .Z(n9737) );
  AND U10642 ( .A(n9738), .B(n9737), .Z(n9888) );
  XNOR U10643 ( .A(n9887), .B(n9888), .Z(n9889) );
  XOR U10644 ( .A(n9890), .B(n9889), .Z(n10071) );
  XNOR U10645 ( .A(n10070), .B(n10071), .Z(n10072) );
  NANDN U10646 ( .A(n9740), .B(n9739), .Z(n9744) );
  NAND U10647 ( .A(n9742), .B(n9741), .Z(n9743) );
  AND U10648 ( .A(n9744), .B(n9743), .Z(n10073) );
  XNOR U10649 ( .A(n10072), .B(n10073), .Z(n10055) );
  NAND U10650 ( .A(n33283), .B(n9745), .Z(n9747) );
  XOR U10651 ( .A(n33020), .B(n22289), .Z(n9893) );
  NANDN U10652 ( .A(n33021), .B(n9893), .Z(n9746) );
  NAND U10653 ( .A(n9747), .B(n9746), .Z(n9971) );
  XNOR U10654 ( .A(b[41]), .B(a[22]), .Z(n9923) );
  OR U10655 ( .A(n9923), .B(n36905), .Z(n9750) );
  NANDN U10656 ( .A(n9748), .B(n36807), .Z(n9749) );
  NAND U10657 ( .A(n9750), .B(n9749), .Z(n9968) );
  XNOR U10658 ( .A(b[45]), .B(a[18]), .Z(n9896) );
  NANDN U10659 ( .A(n9896), .B(n37261), .Z(n9753) );
  NANDN U10660 ( .A(n9751), .B(n37262), .Z(n9752) );
  AND U10661 ( .A(n9753), .B(n9752), .Z(n9969) );
  XNOR U10662 ( .A(n9968), .B(n9969), .Z(n9970) );
  XNOR U10663 ( .A(n9971), .B(n9970), .Z(n10060) );
  XOR U10664 ( .A(b[43]), .B(n15484), .Z(n9926) );
  NANDN U10665 ( .A(n9926), .B(n37068), .Z(n9756) );
  NANDN U10666 ( .A(n9754), .B(n37069), .Z(n9755) );
  NAND U10667 ( .A(n9756), .B(n9755), .Z(n9941) );
  XOR U10668 ( .A(b[53]), .B(n12555), .Z(n9962) );
  NANDN U10669 ( .A(n9962), .B(n37940), .Z(n9759) );
  NANDN U10670 ( .A(n9757), .B(n37941), .Z(n9758) );
  NAND U10671 ( .A(n9759), .B(n9758), .Z(n9938) );
  XOR U10672 ( .A(b[55]), .B(n11986), .Z(n9881) );
  NANDN U10673 ( .A(n9881), .B(n38075), .Z(n9762) );
  NANDN U10674 ( .A(n9760), .B(n38073), .Z(n9761) );
  AND U10675 ( .A(n9762), .B(n9761), .Z(n9939) );
  XNOR U10676 ( .A(n9938), .B(n9939), .Z(n9940) );
  XOR U10677 ( .A(n9941), .B(n9940), .Z(n10061) );
  XNOR U10678 ( .A(n10060), .B(n10061), .Z(n10062) );
  NANDN U10679 ( .A(n9764), .B(n9763), .Z(n9768) );
  NAND U10680 ( .A(n9766), .B(n9765), .Z(n9767) );
  AND U10681 ( .A(n9768), .B(n9767), .Z(n10063) );
  XNOR U10682 ( .A(n10062), .B(n10063), .Z(n10054) );
  XNOR U10683 ( .A(n10055), .B(n10054), .Z(n10057) );
  XOR U10684 ( .A(n10056), .B(n10057), .Z(n10025) );
  XNOR U10685 ( .A(n10025), .B(n10024), .Z(n10026) );
  XNOR U10686 ( .A(n10027), .B(n10026), .Z(n10125) );
  XNOR U10687 ( .A(n10124), .B(n10125), .Z(n10127) );
  XOR U10688 ( .A(n10126), .B(n10127), .Z(n10039) );
  XOR U10689 ( .A(n10038), .B(n10039), .Z(n9860) );
  XNOR U10690 ( .A(n9861), .B(n9860), .Z(n9863) );
  NANDN U10691 ( .A(n9774), .B(n9773), .Z(n9778) );
  NANDN U10692 ( .A(n9776), .B(n9775), .Z(n9777) );
  NAND U10693 ( .A(n9778), .B(n9777), .Z(n9872) );
  NANDN U10694 ( .A(n9780), .B(n9779), .Z(n9784) );
  NAND U10695 ( .A(n9782), .B(n9781), .Z(n9783) );
  AND U10696 ( .A(n9784), .B(n9783), .Z(n9873) );
  XNOR U10697 ( .A(n9872), .B(n9873), .Z(n9874) );
  NANDN U10698 ( .A(n9786), .B(n9785), .Z(n9790) );
  OR U10699 ( .A(n9788), .B(n9787), .Z(n9789) );
  NAND U10700 ( .A(n9790), .B(n9789), .Z(n10118) );
  NANDN U10701 ( .A(n9792), .B(n9791), .Z(n9796) );
  NAND U10702 ( .A(n9794), .B(n9793), .Z(n9795) );
  AND U10703 ( .A(n9796), .B(n9795), .Z(n10119) );
  XNOR U10704 ( .A(n10118), .B(n10119), .Z(n10120) );
  XNOR U10705 ( .A(b[17]), .B(a[46]), .Z(n10103) );
  NANDN U10706 ( .A(n10103), .B(n32543), .Z(n9799) );
  NANDN U10707 ( .A(n9797), .B(n32541), .Z(n9798) );
  NAND U10708 ( .A(n9799), .B(n9798), .Z(n9998) );
  NAND U10709 ( .A(n37469), .B(n9800), .Z(n9802) );
  XOR U10710 ( .A(n978), .B(n14259), .Z(n9953) );
  NAND U10711 ( .A(n9953), .B(n37471), .Z(n9801) );
  NAND U10712 ( .A(n9802), .B(n9801), .Z(n9995) );
  XOR U10713 ( .A(b[49]), .B(n14210), .Z(n9956) );
  OR U10714 ( .A(n9956), .B(n37756), .Z(n9805) );
  NANDN U10715 ( .A(n9803), .B(n37652), .Z(n9804) );
  AND U10716 ( .A(n9805), .B(n9804), .Z(n9996) );
  XNOR U10717 ( .A(n9995), .B(n9996), .Z(n9997) );
  XNOR U10718 ( .A(n9998), .B(n9997), .Z(n10069) );
  XOR U10719 ( .A(b[37]), .B(n17133), .Z(n9989) );
  NANDN U10720 ( .A(n9989), .B(n36311), .Z(n9808) );
  NANDN U10721 ( .A(n9806), .B(n36309), .Z(n9807) );
  NAND U10722 ( .A(n9808), .B(n9807), .Z(n9911) );
  XOR U10723 ( .A(b[57]), .B(n11406), .Z(n10091) );
  OR U10724 ( .A(n10091), .B(n965), .Z(n9811) );
  NANDN U10725 ( .A(n9809), .B(n38194), .Z(n9810) );
  NAND U10726 ( .A(n9811), .B(n9810), .Z(n9908) );
  XOR U10727 ( .A(n31123), .B(n25860), .Z(n9899) );
  NAND U10728 ( .A(n9899), .B(n29949), .Z(n9814) );
  NAND U10729 ( .A(n29948), .B(n9812), .Z(n9813) );
  AND U10730 ( .A(n9814), .B(n9813), .Z(n9909) );
  XNOR U10731 ( .A(n9908), .B(n9909), .Z(n9910) );
  XNOR U10732 ( .A(n9911), .B(n9910), .Z(n10066) );
  NANDN U10733 ( .A(n9816), .B(n9815), .Z(n9820) );
  NAND U10734 ( .A(n9818), .B(n9817), .Z(n9819) );
  NAND U10735 ( .A(n9820), .B(n9819), .Z(n10067) );
  XNOR U10736 ( .A(n10066), .B(n10067), .Z(n10068) );
  XOR U10737 ( .A(n10069), .B(n10068), .Z(n10042) );
  XOR U10738 ( .A(n10042), .B(n10043), .Z(n10045) );
  XNOR U10739 ( .A(b[21]), .B(a[42]), .Z(n10106) );
  OR U10740 ( .A(n10106), .B(n33634), .Z(n9827) );
  NAND U10741 ( .A(n9825), .B(n33464), .Z(n9826) );
  NAND U10742 ( .A(n9827), .B(n9826), .Z(n9917) );
  XOR U10743 ( .A(b[31]), .B(n18841), .Z(n10088) );
  NANDN U10744 ( .A(n10088), .B(n35313), .Z(n9830) );
  NAND U10745 ( .A(n9828), .B(n35311), .Z(n9829) );
  NAND U10746 ( .A(n9830), .B(n9829), .Z(n9914) );
  NAND U10747 ( .A(n34044), .B(n9831), .Z(n9833) );
  XOR U10748 ( .A(n34510), .B(n21149), .Z(n9929) );
  NANDN U10749 ( .A(n33867), .B(n9929), .Z(n9832) );
  AND U10750 ( .A(n9833), .B(n9832), .Z(n9915) );
  XNOR U10751 ( .A(n9914), .B(n9915), .Z(n9916) );
  XNOR U10752 ( .A(n9917), .B(n9916), .Z(n10082) );
  NANDN U10753 ( .A(n9835), .B(n9834), .Z(n9839) );
  NAND U10754 ( .A(n9837), .B(n9836), .Z(n9838) );
  NAND U10755 ( .A(n9839), .B(n9838), .Z(n10083) );
  XOR U10756 ( .A(n10082), .B(n10083), .Z(n10085) );
  NAND U10757 ( .A(n9841), .B(n9840), .Z(n9977) );
  XOR U10758 ( .A(b[33]), .B(n18804), .Z(n10011) );
  NANDN U10759 ( .A(n10011), .B(n35620), .Z(n9844) );
  NANDN U10760 ( .A(n9842), .B(n35621), .Z(n9843) );
  NAND U10761 ( .A(n9844), .B(n9843), .Z(n9975) );
  XNOR U10762 ( .A(n967), .B(a[60]), .Z(n9935) );
  NAND U10763 ( .A(n9935), .B(n28939), .Z(n9847) );
  NANDN U10764 ( .A(n9845), .B(n28938), .Z(n9846) );
  AND U10765 ( .A(n9847), .B(n9846), .Z(n9974) );
  XNOR U10766 ( .A(n9975), .B(n9974), .Z(n9976) );
  XNOR U10767 ( .A(n9977), .B(n9976), .Z(n10084) );
  XNOR U10768 ( .A(n10085), .B(n10084), .Z(n10044) );
  XNOR U10769 ( .A(n10045), .B(n10044), .Z(n10121) );
  XNOR U10770 ( .A(n10120), .B(n10121), .Z(n9875) );
  XOR U10771 ( .A(n9874), .B(n9875), .Z(n9862) );
  XOR U10772 ( .A(n9863), .B(n9862), .Z(n9869) );
  XNOR U10773 ( .A(n9868), .B(n9869), .Z(n9854) );
  XNOR U10774 ( .A(n9855), .B(n9854), .Z(n9857) );
  XNOR U10775 ( .A(n9856), .B(n9857), .Z(n9848) );
  XOR U10776 ( .A(n9849), .B(n9848), .Z(n9850) );
  XOR U10777 ( .A(n9851), .B(n9850), .Z(n10131) );
  XOR U10778 ( .A(n10132), .B(n10131), .Z(c[126]) );
  NAND U10779 ( .A(n9849), .B(n9848), .Z(n9853) );
  NAND U10780 ( .A(n9851), .B(n9850), .Z(n9852) );
  NAND U10781 ( .A(n9853), .B(n9852), .Z(n10143) );
  NAND U10782 ( .A(n9855), .B(n9854), .Z(n9859) );
  NANDN U10783 ( .A(n9857), .B(n9856), .Z(n9858) );
  NAND U10784 ( .A(n9859), .B(n9858), .Z(n10141) );
  NAND U10785 ( .A(n9861), .B(n9860), .Z(n9865) );
  NANDN U10786 ( .A(n9863), .B(n9862), .Z(n9864) );
  NAND U10787 ( .A(n9865), .B(n9864), .Z(n10146) );
  NANDN U10788 ( .A(n9867), .B(n9866), .Z(n9871) );
  NANDN U10789 ( .A(n9869), .B(n9868), .Z(n9870) );
  AND U10790 ( .A(n9871), .B(n9870), .Z(n10147) );
  XNOR U10791 ( .A(n10146), .B(n10147), .Z(n10148) );
  NANDN U10792 ( .A(n9873), .B(n9872), .Z(n9877) );
  NAND U10793 ( .A(n9875), .B(n9874), .Z(n9876) );
  NAND U10794 ( .A(n9877), .B(n9876), .Z(n10406) );
  NAND U10795 ( .A(n35188), .B(n9878), .Z(n9880) );
  XOR U10796 ( .A(n35540), .B(n20315), .Z(n10254) );
  NANDN U10797 ( .A(n34968), .B(n10254), .Z(n9879) );
  NAND U10798 ( .A(n9880), .B(n9879), .Z(n10370) );
  XOR U10799 ( .A(b[55]), .B(n12258), .Z(n10300) );
  NANDN U10800 ( .A(n10300), .B(n38075), .Z(n9883) );
  NANDN U10801 ( .A(n9881), .B(n38073), .Z(n9882) );
  AND U10802 ( .A(n9883), .B(n9882), .Z(n10368) );
  NANDN U10803 ( .A(n966), .B(a[63]), .Z(n9884) );
  XOR U10804 ( .A(n29232), .B(n9884), .Z(n9886) );
  NANDN U10805 ( .A(b[0]), .B(a[62]), .Z(n9885) );
  AND U10806 ( .A(n9886), .B(n9885), .Z(n10367) );
  XNOR U10807 ( .A(n10368), .B(n10367), .Z(n10369) );
  XOR U10808 ( .A(n10370), .B(n10369), .Z(n10379) );
  NANDN U10809 ( .A(n9888), .B(n9887), .Z(n9892) );
  NAND U10810 ( .A(n9890), .B(n9889), .Z(n9891) );
  NAND U10811 ( .A(n9892), .B(n9891), .Z(n10380) );
  XNOR U10812 ( .A(n10379), .B(n10380), .Z(n10382) );
  NAND U10813 ( .A(n33283), .B(n9893), .Z(n9895) );
  XOR U10814 ( .A(n33020), .B(n22579), .Z(n10239) );
  NANDN U10815 ( .A(n33021), .B(n10239), .Z(n9894) );
  NAND U10816 ( .A(n9895), .B(n9894), .Z(n10230) );
  XNOR U10817 ( .A(b[45]), .B(a[19]), .Z(n10294) );
  NANDN U10818 ( .A(n10294), .B(n37261), .Z(n9898) );
  NANDN U10819 ( .A(n9896), .B(n37262), .Z(n9897) );
  NAND U10820 ( .A(n9898), .B(n9897), .Z(n10227) );
  XOR U10821 ( .A(n31123), .B(n26122), .Z(n10218) );
  NAND U10822 ( .A(n10218), .B(n29949), .Z(n9901) );
  NAND U10823 ( .A(n29948), .B(n9899), .Z(n9900) );
  AND U10824 ( .A(n9901), .B(n9900), .Z(n10228) );
  XNOR U10825 ( .A(n10227), .B(n10228), .Z(n10229) );
  XOR U10826 ( .A(n10230), .B(n10229), .Z(n10381) );
  XNOR U10827 ( .A(n10382), .B(n10381), .Z(n10394) );
  NANDN U10828 ( .A(n9903), .B(n9902), .Z(n9907) );
  NAND U10829 ( .A(n9905), .B(n9904), .Z(n9906) );
  NAND U10830 ( .A(n9907), .B(n9906), .Z(n10391) );
  NANDN U10831 ( .A(n9909), .B(n9908), .Z(n9913) );
  NAND U10832 ( .A(n9911), .B(n9910), .Z(n9912) );
  AND U10833 ( .A(n9913), .B(n9912), .Z(n10392) );
  XNOR U10834 ( .A(n10391), .B(n10392), .Z(n10393) );
  XOR U10835 ( .A(n10394), .B(n10393), .Z(n10285) );
  NANDN U10836 ( .A(n9915), .B(n9914), .Z(n9919) );
  NAND U10837 ( .A(n9917), .B(n9916), .Z(n9918) );
  NAND U10838 ( .A(n9919), .B(n9918), .Z(n10342) );
  XOR U10839 ( .A(b[9]), .B(n25466), .Z(n10191) );
  NANDN U10840 ( .A(n10191), .B(n30509), .Z(n9922) );
  NANDN U10841 ( .A(n9920), .B(n30846), .Z(n9921) );
  NAND U10842 ( .A(n9922), .B(n9921), .Z(n10209) );
  XNOR U10843 ( .A(b[41]), .B(n16269), .Z(n10297) );
  NANDN U10844 ( .A(n36905), .B(n10297), .Z(n9925) );
  NANDN U10845 ( .A(n9923), .B(n36807), .Z(n9924) );
  NAND U10846 ( .A(n9925), .B(n9924), .Z(n10206) );
  XOR U10847 ( .A(b[43]), .B(n16220), .Z(n10291) );
  NANDN U10848 ( .A(n10291), .B(n37068), .Z(n9928) );
  NANDN U10849 ( .A(n9926), .B(n37069), .Z(n9927) );
  AND U10850 ( .A(n9928), .B(n9927), .Z(n10207) );
  XNOR U10851 ( .A(n10206), .B(n10207), .Z(n10208) );
  XNOR U10852 ( .A(n10209), .B(n10208), .Z(n10339) );
  NAND U10853 ( .A(n34044), .B(n9929), .Z(n9931) );
  XOR U10854 ( .A(b[23]), .B(n21441), .Z(n10257) );
  OR U10855 ( .A(n10257), .B(n33867), .Z(n9930) );
  NAND U10856 ( .A(n9931), .B(n9930), .Z(n10324) );
  XNOR U10857 ( .A(b[5]), .B(a[59]), .Z(n10360) );
  OR U10858 ( .A(n10360), .B(n29363), .Z(n9934) );
  NANDN U10859 ( .A(n9932), .B(n29864), .Z(n9933) );
  NAND U10860 ( .A(n9934), .B(n9933), .Z(n10321) );
  XOR U10861 ( .A(b[3]), .B(n27773), .Z(n10332) );
  NANDN U10862 ( .A(n10332), .B(n28939), .Z(n9937) );
  NAND U10863 ( .A(n9935), .B(n28938), .Z(n9936) );
  AND U10864 ( .A(n9937), .B(n9936), .Z(n10322) );
  XNOR U10865 ( .A(n10321), .B(n10322), .Z(n10323) );
  XOR U10866 ( .A(n10324), .B(n10323), .Z(n10340) );
  XNOR U10867 ( .A(n10339), .B(n10340), .Z(n10341) );
  XOR U10868 ( .A(n10342), .B(n10341), .Z(n10275) );
  NANDN U10869 ( .A(n9939), .B(n9938), .Z(n9943) );
  NAND U10870 ( .A(n9941), .B(n9940), .Z(n9942) );
  NAND U10871 ( .A(n9943), .B(n9942), .Z(n10272) );
  NANDN U10872 ( .A(n9945), .B(n9944), .Z(n9949) );
  NAND U10873 ( .A(n9947), .B(n9946), .Z(n9948) );
  AND U10874 ( .A(n9949), .B(n9948), .Z(n10273) );
  XNOR U10875 ( .A(n10272), .B(n10273), .Z(n10274) );
  XNOR U10876 ( .A(n10275), .B(n10274), .Z(n10283) );
  NAND U10877 ( .A(n34848), .B(n9950), .Z(n9952) );
  XOR U10878 ( .A(n35375), .B(n20352), .Z(n10248) );
  NAND U10879 ( .A(n34618), .B(n10248), .Z(n9951) );
  NAND U10880 ( .A(n9952), .B(n9951), .Z(n10263) );
  NAND U10881 ( .A(n37469), .B(n9953), .Z(n9955) );
  XOR U10882 ( .A(n978), .B(n14514), .Z(n10315) );
  NAND U10883 ( .A(n10315), .B(n37471), .Z(n9954) );
  NAND U10884 ( .A(n9955), .B(n9954), .Z(n10260) );
  XOR U10885 ( .A(b[49]), .B(n13976), .Z(n10197) );
  OR U10886 ( .A(n10197), .B(n37756), .Z(n9958) );
  NANDN U10887 ( .A(n9956), .B(n37652), .Z(n9957) );
  AND U10888 ( .A(n9958), .B(n9957), .Z(n10261) );
  XNOR U10889 ( .A(n10260), .B(n10261), .Z(n10262) );
  XNOR U10890 ( .A(n10263), .B(n10262), .Z(n10338) );
  XOR U10891 ( .A(b[51]), .B(n13509), .Z(n10318) );
  NANDN U10892 ( .A(n10318), .B(n37803), .Z(n9961) );
  NANDN U10893 ( .A(n9959), .B(n37802), .Z(n9960) );
  NAND U10894 ( .A(n9961), .B(n9960), .Z(n10376) );
  XOR U10895 ( .A(b[53]), .B(n12830), .Z(n10194) );
  NANDN U10896 ( .A(n10194), .B(n37940), .Z(n9964) );
  NANDN U10897 ( .A(n9962), .B(n37941), .Z(n9963) );
  NAND U10898 ( .A(n9964), .B(n9963), .Z(n10373) );
  XNOR U10899 ( .A(b[35]), .B(n18003), .Z(n10329) );
  NAND U10900 ( .A(n35985), .B(n10329), .Z(n9967) );
  NANDN U10901 ( .A(n9965), .B(n35986), .Z(n9966) );
  AND U10902 ( .A(n9967), .B(n9966), .Z(n10374) );
  XNOR U10903 ( .A(n10373), .B(n10374), .Z(n10375) );
  XNOR U10904 ( .A(n10376), .B(n10375), .Z(n10335) );
  NANDN U10905 ( .A(n9969), .B(n9968), .Z(n9973) );
  NAND U10906 ( .A(n9971), .B(n9970), .Z(n9972) );
  NAND U10907 ( .A(n9973), .B(n9972), .Z(n10336) );
  XNOR U10908 ( .A(n10335), .B(n10336), .Z(n10337) );
  XOR U10909 ( .A(n10338), .B(n10337), .Z(n10282) );
  XOR U10910 ( .A(n10283), .B(n10282), .Z(n10284) );
  XNOR U10911 ( .A(n10285), .B(n10284), .Z(n10158) );
  NANDN U10912 ( .A(n9975), .B(n9974), .Z(n9979) );
  NAND U10913 ( .A(n9977), .B(n9976), .Z(n9978) );
  NAND U10914 ( .A(n9979), .B(n9978), .Z(n10385) );
  NANDN U10915 ( .A(n9981), .B(n9980), .Z(n9985) );
  NAND U10916 ( .A(n9983), .B(n9982), .Z(n9984) );
  NAND U10917 ( .A(n9985), .B(n9984), .Z(n10386) );
  XNOR U10918 ( .A(n10385), .B(n10386), .Z(n10387) );
  XOR U10919 ( .A(b[11]), .B(n25001), .Z(n10203) );
  OR U10920 ( .A(n10203), .B(n31369), .Z(n9988) );
  NANDN U10921 ( .A(n9986), .B(n31119), .Z(n9987) );
  NAND U10922 ( .A(n9988), .B(n9987), .Z(n10309) );
  XOR U10923 ( .A(b[37]), .B(n17960), .Z(n10357) );
  NANDN U10924 ( .A(n10357), .B(n36311), .Z(n9991) );
  NANDN U10925 ( .A(n9989), .B(n36309), .Z(n9990) );
  NAND U10926 ( .A(n9991), .B(n9990), .Z(n10306) );
  XOR U10927 ( .A(b[39]), .B(n16916), .Z(n10212) );
  NANDN U10928 ( .A(n10212), .B(n36553), .Z(n9994) );
  NANDN U10929 ( .A(n9992), .B(n36643), .Z(n9993) );
  AND U10930 ( .A(n9994), .B(n9993), .Z(n10307) );
  XNOR U10931 ( .A(n10306), .B(n10307), .Z(n10308) );
  XNOR U10932 ( .A(n10309), .B(n10308), .Z(n10233) );
  NANDN U10933 ( .A(n9996), .B(n9995), .Z(n10000) );
  NAND U10934 ( .A(n9998), .B(n9997), .Z(n9999) );
  NAND U10935 ( .A(n10000), .B(n9999), .Z(n10234) );
  XOR U10936 ( .A(n10233), .B(n10234), .Z(n10236) );
  XNOR U10937 ( .A(n985), .B(a[0]), .Z(n10003) );
  XNOR U10938 ( .A(n985), .B(b[62]), .Z(n10002) );
  XNOR U10939 ( .A(n985), .B(b[61]), .Z(n10001) );
  AND U10940 ( .A(n10002), .B(n10001), .Z(n38423) );
  NAND U10941 ( .A(n10003), .B(n38423), .Z(n10005) );
  XNOR U10942 ( .A(n985), .B(a[1]), .Z(n10364) );
  NAND U10943 ( .A(n10364), .B(n38422), .Z(n10004) );
  AND U10944 ( .A(n10005), .B(n10004), .Z(n10328) );
  XOR U10945 ( .A(b[61]), .B(n10524), .Z(n10354) );
  OR U10946 ( .A(n10354), .B(n38371), .Z(n10008) );
  NANDN U10947 ( .A(n10006), .B(n38369), .Z(n10007) );
  AND U10948 ( .A(n10008), .B(n10007), .Z(n10327) );
  XOR U10949 ( .A(n10328), .B(n10327), .Z(n10223) );
  AND U10950 ( .A(b[61]), .B(b[62]), .Z(n38462) );
  NOR U10951 ( .A(n985), .B(n38462), .Z(n10010) );
  ANDN U10952 ( .B(n38433), .A(b[61]), .Z(n38461) );
  OR U10953 ( .A(n38461), .B(n986), .Z(n10009) );
  NAND U10954 ( .A(n10010), .B(n10009), .Z(n10221) );
  XNOR U10955 ( .A(n974), .B(a[31]), .Z(n10245) );
  NAND U10956 ( .A(n35620), .B(n10245), .Z(n10013) );
  NANDN U10957 ( .A(n10011), .B(n35621), .Z(n10012) );
  NAND U10958 ( .A(n10013), .B(n10012), .Z(n10222) );
  XOR U10959 ( .A(n10221), .B(n10222), .Z(n10224) );
  XNOR U10960 ( .A(n10223), .B(n10224), .Z(n10235) );
  XOR U10961 ( .A(n10236), .B(n10235), .Z(n10388) );
  XNOR U10962 ( .A(n10387), .B(n10388), .Z(n10179) );
  NANDN U10963 ( .A(n10019), .B(n10018), .Z(n10023) );
  NAND U10964 ( .A(n10021), .B(n10020), .Z(n10022) );
  NAND U10965 ( .A(n10023), .B(n10022), .Z(n10177) );
  XNOR U10966 ( .A(n10176), .B(n10177), .Z(n10178) );
  XNOR U10967 ( .A(n10179), .B(n10178), .Z(n10159) );
  XOR U10968 ( .A(n10158), .B(n10159), .Z(n10160) );
  NANDN U10969 ( .A(n10025), .B(n10024), .Z(n10029) );
  NAND U10970 ( .A(n10027), .B(n10026), .Z(n10028) );
  NAND U10971 ( .A(n10029), .B(n10028), .Z(n10161) );
  XOR U10972 ( .A(n10160), .B(n10161), .Z(n10403) );
  NANDN U10973 ( .A(n10031), .B(n10030), .Z(n10035) );
  NAND U10974 ( .A(n10033), .B(n10032), .Z(n10034) );
  AND U10975 ( .A(n10035), .B(n10034), .Z(n10404) );
  XNOR U10976 ( .A(n10403), .B(n10404), .Z(n10405) );
  XNOR U10977 ( .A(n10406), .B(n10405), .Z(n10418) );
  NANDN U10978 ( .A(n10037), .B(n10036), .Z(n10041) );
  NAND U10979 ( .A(n10039), .B(n10038), .Z(n10040) );
  NAND U10980 ( .A(n10041), .B(n10040), .Z(n10415) );
  NANDN U10981 ( .A(n10043), .B(n10042), .Z(n10047) );
  OR U10982 ( .A(n10045), .B(n10044), .Z(n10046) );
  NAND U10983 ( .A(n10047), .B(n10046), .Z(n10155) );
  NANDN U10984 ( .A(n10049), .B(n10048), .Z(n10053) );
  NAND U10985 ( .A(n10051), .B(n10050), .Z(n10052) );
  NAND U10986 ( .A(n10053), .B(n10052), .Z(n10152) );
  OR U10987 ( .A(n10055), .B(n10054), .Z(n10059) );
  NANDN U10988 ( .A(n10057), .B(n10056), .Z(n10058) );
  AND U10989 ( .A(n10059), .B(n10058), .Z(n10153) );
  XNOR U10990 ( .A(n10152), .B(n10153), .Z(n10154) );
  XNOR U10991 ( .A(n10155), .B(n10154), .Z(n10409) );
  NANDN U10992 ( .A(n10061), .B(n10060), .Z(n10065) );
  NAND U10993 ( .A(n10063), .B(n10062), .Z(n10064) );
  NAND U10994 ( .A(n10065), .B(n10064), .Z(n10400) );
  NANDN U10995 ( .A(n10071), .B(n10070), .Z(n10075) );
  NAND U10996 ( .A(n10073), .B(n10072), .Z(n10074) );
  AND U10997 ( .A(n10075), .B(n10074), .Z(n10398) );
  XNOR U10998 ( .A(n10397), .B(n10398), .Z(n10399) );
  XNOR U10999 ( .A(n10400), .B(n10399), .Z(n10164) );
  NANDN U11000 ( .A(n10077), .B(n10076), .Z(n10081) );
  NAND U11001 ( .A(n10079), .B(n10078), .Z(n10080) );
  NAND U11002 ( .A(n10081), .B(n10080), .Z(n10173) );
  NANDN U11003 ( .A(n10083), .B(n10082), .Z(n10087) );
  OR U11004 ( .A(n10085), .B(n10084), .Z(n10086) );
  NAND U11005 ( .A(n10087), .B(n10086), .Z(n10171) );
  XOR U11006 ( .A(b[31]), .B(n19656), .Z(n10188) );
  NANDN U11007 ( .A(n10188), .B(n35313), .Z(n10090) );
  NANDN U11008 ( .A(n10088), .B(n35311), .Z(n10089) );
  NAND U11009 ( .A(n10090), .B(n10089), .Z(n10269) );
  XOR U11010 ( .A(b[57]), .B(n11694), .Z(n10303) );
  OR U11011 ( .A(n10303), .B(n965), .Z(n10093) );
  NANDN U11012 ( .A(n10091), .B(n38194), .Z(n10092) );
  NAND U11013 ( .A(n10093), .B(n10092), .Z(n10266) );
  NAND U11014 ( .A(n38326), .B(n10094), .Z(n10096) );
  XOR U11015 ( .A(n38400), .B(n11202), .Z(n10215) );
  NANDN U11016 ( .A(n38273), .B(n10215), .Z(n10095) );
  AND U11017 ( .A(n10096), .B(n10095), .Z(n10267) );
  XNOR U11018 ( .A(n10266), .B(n10267), .Z(n10268) );
  XNOR U11019 ( .A(n10269), .B(n10268), .Z(n10281) );
  NANDN U11020 ( .A(n10098), .B(n10097), .Z(n10102) );
  OR U11021 ( .A(n10100), .B(n10099), .Z(n10101) );
  NAND U11022 ( .A(n10102), .B(n10101), .Z(n10279) );
  XNOR U11023 ( .A(b[17]), .B(a[47]), .Z(n10288) );
  NANDN U11024 ( .A(n10288), .B(n32543), .Z(n10105) );
  NANDN U11025 ( .A(n10103), .B(n32541), .Z(n10104) );
  NAND U11026 ( .A(n10105), .B(n10104), .Z(n10348) );
  XNOR U11027 ( .A(b[21]), .B(a[43]), .Z(n10242) );
  OR U11028 ( .A(n10242), .B(n33634), .Z(n10108) );
  NANDN U11029 ( .A(n10106), .B(n33464), .Z(n10107) );
  NAND U11030 ( .A(n10108), .B(n10107), .Z(n10345) );
  XNOR U11031 ( .A(b[25]), .B(n20867), .Z(n10251) );
  NANDN U11032 ( .A(n34219), .B(n10251), .Z(n10111) );
  NAND U11033 ( .A(n34217), .B(n10109), .Z(n10110) );
  AND U11034 ( .A(n10111), .B(n10110), .Z(n10346) );
  XNOR U11035 ( .A(n10345), .B(n10346), .Z(n10347) );
  XNOR U11036 ( .A(n10348), .B(n10347), .Z(n10185) );
  NAND U11037 ( .A(n31874), .B(n10112), .Z(n10114) );
  XNOR U11038 ( .A(n971), .B(a[51]), .Z(n10200) );
  NANDN U11039 ( .A(n31550), .B(n10200), .Z(n10113) );
  NAND U11040 ( .A(n10114), .B(n10113), .Z(n10183) );
  NANDN U11041 ( .A(n10115), .B(n32011), .Z(n10117) );
  XNOR U11042 ( .A(n972), .B(a[49]), .Z(n10312) );
  NANDN U11043 ( .A(n32010), .B(n10312), .Z(n10116) );
  AND U11044 ( .A(n10117), .B(n10116), .Z(n10182) );
  XNOR U11045 ( .A(n10183), .B(n10182), .Z(n10184) );
  XOR U11046 ( .A(n10185), .B(n10184), .Z(n10278) );
  XNOR U11047 ( .A(n10279), .B(n10278), .Z(n10280) );
  XOR U11048 ( .A(n10281), .B(n10280), .Z(n10170) );
  XOR U11049 ( .A(n10171), .B(n10170), .Z(n10172) );
  XOR U11050 ( .A(n10173), .B(n10172), .Z(n10165) );
  XNOR U11051 ( .A(n10164), .B(n10165), .Z(n10166) );
  NANDN U11052 ( .A(n10119), .B(n10118), .Z(n10123) );
  NANDN U11053 ( .A(n10121), .B(n10120), .Z(n10122) );
  AND U11054 ( .A(n10123), .B(n10122), .Z(n10167) );
  XNOR U11055 ( .A(n10166), .B(n10167), .Z(n10410) );
  XOR U11056 ( .A(n10409), .B(n10410), .Z(n10412) );
  NANDN U11057 ( .A(n10125), .B(n10124), .Z(n10129) );
  NAND U11058 ( .A(n10127), .B(n10126), .Z(n10128) );
  NAND U11059 ( .A(n10129), .B(n10128), .Z(n10411) );
  XOR U11060 ( .A(n10412), .B(n10411), .Z(n10416) );
  XNOR U11061 ( .A(n10415), .B(n10416), .Z(n10417) );
  XOR U11062 ( .A(n10418), .B(n10417), .Z(n10149) );
  XNOR U11063 ( .A(n10148), .B(n10149), .Z(n10140) );
  XOR U11064 ( .A(n10141), .B(n10140), .Z(n10142) );
  XNOR U11065 ( .A(n10143), .B(n10142), .Z(n10135) );
  XNOR U11066 ( .A(n10135), .B(sreg[127]), .Z(n10137) );
  NAND U11067 ( .A(n10130), .B(sreg[126]), .Z(n10134) );
  OR U11068 ( .A(n10132), .B(n10131), .Z(n10133) );
  AND U11069 ( .A(n10134), .B(n10133), .Z(n10136) );
  XOR U11070 ( .A(n10137), .B(n10136), .Z(c[127]) );
  NAND U11071 ( .A(n10135), .B(sreg[127]), .Z(n10139) );
  OR U11072 ( .A(n10137), .B(n10136), .Z(n10138) );
  NAND U11073 ( .A(n10139), .B(n10138), .Z(n10709) );
  XNOR U11074 ( .A(n10709), .B(sreg[128]), .Z(n10711) );
  NAND U11075 ( .A(n10141), .B(n10140), .Z(n10145) );
  NAND U11076 ( .A(n10143), .B(n10142), .Z(n10144) );
  NAND U11077 ( .A(n10145), .B(n10144), .Z(n10424) );
  NANDN U11078 ( .A(n10147), .B(n10146), .Z(n10151) );
  NANDN U11079 ( .A(n10149), .B(n10148), .Z(n10150) );
  NAND U11080 ( .A(n10151), .B(n10150), .Z(n10421) );
  NANDN U11081 ( .A(n10153), .B(n10152), .Z(n10157) );
  NAND U11082 ( .A(n10155), .B(n10154), .Z(n10156) );
  NAND U11083 ( .A(n10157), .B(n10156), .Z(n10672) );
  OR U11084 ( .A(n10159), .B(n10158), .Z(n10163) );
  NANDN U11085 ( .A(n10161), .B(n10160), .Z(n10162) );
  NAND U11086 ( .A(n10163), .B(n10162), .Z(n10670) );
  NANDN U11087 ( .A(n10165), .B(n10164), .Z(n10169) );
  NAND U11088 ( .A(n10167), .B(n10166), .Z(n10168) );
  AND U11089 ( .A(n10169), .B(n10168), .Z(n10669) );
  XNOR U11090 ( .A(n10670), .B(n10669), .Z(n10671) );
  XNOR U11091 ( .A(n10672), .B(n10671), .Z(n10678) );
  NAND U11092 ( .A(n10171), .B(n10170), .Z(n10175) );
  NAND U11093 ( .A(n10173), .B(n10172), .Z(n10174) );
  NAND U11094 ( .A(n10175), .B(n10174), .Z(n10684) );
  NANDN U11095 ( .A(n10177), .B(n10176), .Z(n10181) );
  NAND U11096 ( .A(n10179), .B(n10178), .Z(n10180) );
  NAND U11097 ( .A(n10181), .B(n10180), .Z(n10681) );
  NANDN U11098 ( .A(n10183), .B(n10182), .Z(n10187) );
  NAND U11099 ( .A(n10185), .B(n10184), .Z(n10186) );
  AND U11100 ( .A(n10187), .B(n10186), .Z(n10703) );
  XOR U11101 ( .A(b[31]), .B(n19513), .Z(n10461) );
  NANDN U11102 ( .A(n10461), .B(n35313), .Z(n10190) );
  NANDN U11103 ( .A(n10188), .B(n35311), .Z(n10189) );
  NAND U11104 ( .A(n10190), .B(n10189), .Z(n10494) );
  XOR U11105 ( .A(n969), .B(n25860), .Z(n10609) );
  NAND U11106 ( .A(n30509), .B(n10609), .Z(n10193) );
  NANDN U11107 ( .A(n10191), .B(n30846), .Z(n10192) );
  NAND U11108 ( .A(n10193), .B(n10192), .Z(n10491) );
  XOR U11109 ( .A(b[53]), .B(n13106), .Z(n10579) );
  NANDN U11110 ( .A(n10579), .B(n37940), .Z(n10196) );
  NANDN U11111 ( .A(n10194), .B(n37941), .Z(n10195) );
  AND U11112 ( .A(n10196), .B(n10195), .Z(n10492) );
  XNOR U11113 ( .A(n10491), .B(n10492), .Z(n10493) );
  XNOR U11114 ( .A(n10494), .B(n10493), .Z(n10445) );
  XOR U11115 ( .A(n979), .B(n14259), .Z(n10603) );
  NANDN U11116 ( .A(n37756), .B(n10603), .Z(n10199) );
  NANDN U11117 ( .A(n10197), .B(n37652), .Z(n10198) );
  NAND U11118 ( .A(n10199), .B(n10198), .Z(n10636) );
  XOR U11119 ( .A(b[13]), .B(n25134), .Z(n10482) );
  OR U11120 ( .A(n10482), .B(n31550), .Z(n10202) );
  NAND U11121 ( .A(n10200), .B(n31874), .Z(n10201) );
  NAND U11122 ( .A(n10202), .B(n10201), .Z(n10633) );
  XOR U11123 ( .A(b[11]), .B(n25177), .Z(n10594) );
  OR U11124 ( .A(n10594), .B(n31369), .Z(n10205) );
  NANDN U11125 ( .A(n10203), .B(n31119), .Z(n10204) );
  AND U11126 ( .A(n10205), .B(n10204), .Z(n10634) );
  XNOR U11127 ( .A(n10633), .B(n10634), .Z(n10635) );
  XOR U11128 ( .A(n10636), .B(n10635), .Z(n10446) );
  XNOR U11129 ( .A(n10445), .B(n10446), .Z(n10447) );
  NANDN U11130 ( .A(n10207), .B(n10206), .Z(n10211) );
  NAND U11131 ( .A(n10209), .B(n10208), .Z(n10210) );
  AND U11132 ( .A(n10211), .B(n10210), .Z(n10448) );
  XNOR U11133 ( .A(n10447), .B(n10448), .Z(n10704) );
  XOR U11134 ( .A(n10703), .B(n10704), .Z(n10705) );
  XOR U11135 ( .A(b[39]), .B(n17133), .Z(n10573) );
  NANDN U11136 ( .A(n10573), .B(n36553), .Z(n10214) );
  NANDN U11137 ( .A(n10212), .B(n36643), .Z(n10213) );
  NAND U11138 ( .A(n10214), .B(n10213), .Z(n10537) );
  NAND U11139 ( .A(n38326), .B(n10215), .Z(n10217) );
  XOR U11140 ( .A(n38400), .B(n11406), .Z(n10515) );
  NANDN U11141 ( .A(n38273), .B(n10515), .Z(n10216) );
  NAND U11142 ( .A(n10217), .B(n10216), .Z(n10534) );
  XOR U11143 ( .A(n31123), .B(n26347), .Z(n10621) );
  NAND U11144 ( .A(n10621), .B(n29949), .Z(n10220) );
  NAND U11145 ( .A(n29948), .B(n10218), .Z(n10219) );
  AND U11146 ( .A(n10220), .B(n10219), .Z(n10535) );
  XNOR U11147 ( .A(n10534), .B(n10535), .Z(n10536) );
  XOR U11148 ( .A(n10537), .B(n10536), .Z(n10648) );
  NANDN U11149 ( .A(n10222), .B(n10221), .Z(n10226) );
  OR U11150 ( .A(n10224), .B(n10223), .Z(n10225) );
  NAND U11151 ( .A(n10226), .B(n10225), .Z(n10645) );
  NANDN U11152 ( .A(n10228), .B(n10227), .Z(n10232) );
  NAND U11153 ( .A(n10230), .B(n10229), .Z(n10231) );
  NAND U11154 ( .A(n10232), .B(n10231), .Z(n10646) );
  XNOR U11155 ( .A(n10645), .B(n10646), .Z(n10647) );
  XOR U11156 ( .A(n10648), .B(n10647), .Z(n10706) );
  XOR U11157 ( .A(n10705), .B(n10706), .Z(n10442) );
  NANDN U11158 ( .A(n10234), .B(n10233), .Z(n10238) );
  OR U11159 ( .A(n10236), .B(n10235), .Z(n10237) );
  NAND U11160 ( .A(n10238), .B(n10237), .Z(n10439) );
  NAND U11161 ( .A(n33283), .B(n10239), .Z(n10241) );
  XOR U11162 ( .A(n33020), .B(n22964), .Z(n10464) );
  NANDN U11163 ( .A(n33021), .B(n10464), .Z(n10240) );
  NAND U11164 ( .A(n10241), .B(n10240), .Z(n10454) );
  XNOR U11165 ( .A(b[21]), .B(a[44]), .Z(n10467) );
  OR U11166 ( .A(n10467), .B(n33634), .Z(n10244) );
  NANDN U11167 ( .A(n10242), .B(n33464), .Z(n10243) );
  NAND U11168 ( .A(n10244), .B(n10243), .Z(n10451) );
  XOR U11169 ( .A(b[33]), .B(n18841), .Z(n10518) );
  NANDN U11170 ( .A(n10518), .B(n35620), .Z(n10247) );
  NAND U11171 ( .A(n10245), .B(n35621), .Z(n10246) );
  AND U11172 ( .A(n10247), .B(n10246), .Z(n10452) );
  XNOR U11173 ( .A(n10451), .B(n10452), .Z(n10453) );
  XOR U11174 ( .A(n10454), .B(n10453), .Z(n10591) );
  NAND U11175 ( .A(n34848), .B(n10248), .Z(n10250) );
  XOR U11176 ( .A(n35375), .B(n20686), .Z(n10485) );
  NAND U11177 ( .A(n34618), .B(n10485), .Z(n10249) );
  NAND U11178 ( .A(n10250), .B(n10249), .Z(n10531) );
  XNOR U11179 ( .A(b[25]), .B(n21149), .Z(n10567) );
  NANDN U11180 ( .A(n34219), .B(n10567), .Z(n10253) );
  NAND U11181 ( .A(n34217), .B(n10251), .Z(n10252) );
  NAND U11182 ( .A(n10253), .B(n10252), .Z(n10528) );
  NAND U11183 ( .A(n35188), .B(n10254), .Z(n10256) );
  XOR U11184 ( .A(n35540), .B(n19980), .Z(n10488) );
  NANDN U11185 ( .A(n34968), .B(n10488), .Z(n10255) );
  AND U11186 ( .A(n10256), .B(n10255), .Z(n10529) );
  XNOR U11187 ( .A(n10528), .B(n10529), .Z(n10530) );
  XOR U11188 ( .A(n10531), .B(n10530), .Z(n10589) );
  NANDN U11189 ( .A(n10257), .B(n34044), .Z(n10259) );
  XOR U11190 ( .A(n34510), .B(n22246), .Z(n10470) );
  NANDN U11191 ( .A(n33867), .B(n10470), .Z(n10258) );
  NAND U11192 ( .A(n10259), .B(n10258), .Z(n10588) );
  XNOR U11193 ( .A(n10589), .B(n10588), .Z(n10590) );
  XOR U11194 ( .A(n10591), .B(n10590), .Z(n10549) );
  NANDN U11195 ( .A(n10261), .B(n10260), .Z(n10265) );
  NAND U11196 ( .A(n10263), .B(n10262), .Z(n10264) );
  NAND U11197 ( .A(n10265), .B(n10264), .Z(n10546) );
  NANDN U11198 ( .A(n10267), .B(n10266), .Z(n10271) );
  NAND U11199 ( .A(n10269), .B(n10268), .Z(n10270) );
  AND U11200 ( .A(n10271), .B(n10270), .Z(n10547) );
  XNOR U11201 ( .A(n10546), .B(n10547), .Z(n10548) );
  XNOR U11202 ( .A(n10549), .B(n10548), .Z(n10440) );
  XNOR U11203 ( .A(n10439), .B(n10440), .Z(n10441) );
  XOR U11204 ( .A(n10442), .B(n10441), .Z(n10660) );
  NANDN U11205 ( .A(n10273), .B(n10272), .Z(n10277) );
  NAND U11206 ( .A(n10275), .B(n10274), .Z(n10276) );
  NAND U11207 ( .A(n10277), .B(n10276), .Z(n10657) );
  XNOR U11208 ( .A(n10657), .B(n10658), .Z(n10659) );
  XNOR U11209 ( .A(n10660), .B(n10659), .Z(n10682) );
  XNOR U11210 ( .A(n10681), .B(n10682), .Z(n10683) );
  XOR U11211 ( .A(n10684), .B(n10683), .Z(n10436) );
  NAND U11212 ( .A(n10283), .B(n10282), .Z(n10287) );
  NANDN U11213 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U11214 ( .A(n10287), .B(n10286), .Z(n10690) );
  XNOR U11215 ( .A(b[17]), .B(a[48]), .Z(n10570) );
  NANDN U11216 ( .A(n10570), .B(n32543), .Z(n10290) );
  NANDN U11217 ( .A(n10288), .B(n32541), .Z(n10289) );
  NAND U11218 ( .A(n10290), .B(n10289), .Z(n10561) );
  XOR U11219 ( .A(b[43]), .B(n15963), .Z(n10597) );
  NANDN U11220 ( .A(n10597), .B(n37068), .Z(n10293) );
  NANDN U11221 ( .A(n10291), .B(n37069), .Z(n10292) );
  NAND U11222 ( .A(n10293), .B(n10292), .Z(n10558) );
  XNOR U11223 ( .A(b[45]), .B(a[20]), .Z(n10600) );
  NANDN U11224 ( .A(n10600), .B(n37261), .Z(n10296) );
  NANDN U11225 ( .A(n10294), .B(n37262), .Z(n10295) );
  AND U11226 ( .A(n10296), .B(n10295), .Z(n10559) );
  XNOR U11227 ( .A(n10558), .B(n10559), .Z(n10560) );
  XNOR U11228 ( .A(n10561), .B(n10560), .Z(n10497) );
  XNOR U11229 ( .A(b[41]), .B(a[24]), .Z(n10509) );
  OR U11230 ( .A(n10509), .B(n36905), .Z(n10299) );
  NAND U11231 ( .A(n10297), .B(n36807), .Z(n10298) );
  NAND U11232 ( .A(n10299), .B(n10298), .Z(n10585) );
  XOR U11233 ( .A(b[55]), .B(n12555), .Z(n10624) );
  NANDN U11234 ( .A(n10624), .B(n38075), .Z(n10302) );
  NANDN U11235 ( .A(n10300), .B(n38073), .Z(n10301) );
  NAND U11236 ( .A(n10302), .B(n10301), .Z(n10582) );
  XOR U11237 ( .A(b[57]), .B(n11986), .Z(n10512) );
  OR U11238 ( .A(n10512), .B(n965), .Z(n10305) );
  NANDN U11239 ( .A(n10303), .B(n38194), .Z(n10304) );
  AND U11240 ( .A(n10305), .B(n10304), .Z(n10583) );
  XNOR U11241 ( .A(n10582), .B(n10583), .Z(n10584) );
  XOR U11242 ( .A(n10585), .B(n10584), .Z(n10498) );
  XNOR U11243 ( .A(n10497), .B(n10498), .Z(n10499) );
  NANDN U11244 ( .A(n10307), .B(n10306), .Z(n10311) );
  NAND U11245 ( .A(n10309), .B(n10308), .Z(n10310) );
  AND U11246 ( .A(n10311), .B(n10310), .Z(n10500) );
  XOR U11247 ( .A(n10499), .B(n10500), .Z(n10693) );
  XOR U11248 ( .A(b[15]), .B(n24671), .Z(n10564) );
  OR U11249 ( .A(n10564), .B(n32010), .Z(n10314) );
  NAND U11250 ( .A(n10312), .B(n32011), .Z(n10313) );
  NAND U11251 ( .A(n10314), .B(n10313), .Z(n10615) );
  NAND U11252 ( .A(n37469), .B(n10315), .Z(n10317) );
  XOR U11253 ( .A(b[47]), .B(n14905), .Z(n10606) );
  NANDN U11254 ( .A(n10606), .B(n37471), .Z(n10316) );
  NAND U11255 ( .A(n10317), .B(n10316), .Z(n10612) );
  XOR U11256 ( .A(b[51]), .B(n14210), .Z(n10576) );
  NANDN U11257 ( .A(n10576), .B(n37803), .Z(n10320) );
  NANDN U11258 ( .A(n10318), .B(n37802), .Z(n10319) );
  AND U11259 ( .A(n10320), .B(n10319), .Z(n10613) );
  XNOR U11260 ( .A(n10612), .B(n10613), .Z(n10614) );
  XNOR U11261 ( .A(n10615), .B(n10614), .Z(n10639) );
  NANDN U11262 ( .A(n10322), .B(n10321), .Z(n10326) );
  NAND U11263 ( .A(n10324), .B(n10323), .Z(n10325) );
  NAND U11264 ( .A(n10326), .B(n10325), .Z(n10640) );
  XOR U11265 ( .A(n10639), .B(n10640), .Z(n10642) );
  OR U11266 ( .A(n10328), .B(n10327), .Z(n10555) );
  NAND U11267 ( .A(n35986), .B(n10329), .Z(n10331) );
  XNOR U11268 ( .A(b[35]), .B(a[30]), .Z(n10618) );
  NANDN U11269 ( .A(n10618), .B(n35985), .Z(n10330) );
  NAND U11270 ( .A(n10331), .B(n10330), .Z(n10553) );
  XNOR U11271 ( .A(n967), .B(a[62]), .Z(n10479) );
  NAND U11272 ( .A(n10479), .B(n28939), .Z(n10334) );
  NANDN U11273 ( .A(n10332), .B(n28938), .Z(n10333) );
  AND U11274 ( .A(n10334), .B(n10333), .Z(n10552) );
  XNOR U11275 ( .A(n10553), .B(n10552), .Z(n10554) );
  XNOR U11276 ( .A(n10555), .B(n10554), .Z(n10641) );
  XOR U11277 ( .A(n10642), .B(n10641), .Z(n10694) );
  XNOR U11278 ( .A(n10693), .B(n10694), .Z(n10696) );
  XNOR U11279 ( .A(n10696), .B(n10695), .Z(n10699) );
  NANDN U11280 ( .A(n10340), .B(n10339), .Z(n10344) );
  NANDN U11281 ( .A(n10342), .B(n10341), .Z(n10343) );
  AND U11282 ( .A(n10344), .B(n10343), .Z(n10700) );
  XNOR U11283 ( .A(n10699), .B(n10700), .Z(n10701) );
  NANDN U11284 ( .A(n10346), .B(n10345), .Z(n10350) );
  NAND U11285 ( .A(n10348), .B(n10347), .Z(n10349) );
  AND U11286 ( .A(n10350), .B(n10349), .Z(n10543) );
  NANDN U11287 ( .A(n966), .B(a[64]), .Z(n10351) );
  XOR U11288 ( .A(n29232), .B(n10351), .Z(n10353) );
  NANDN U11289 ( .A(b[0]), .B(a[63]), .Z(n10352) );
  AND U11290 ( .A(n10353), .B(n10352), .Z(n10627) );
  XOR U11291 ( .A(b[61]), .B(n10854), .Z(n10458) );
  OR U11292 ( .A(n10458), .B(n38371), .Z(n10356) );
  NANDN U11293 ( .A(n10354), .B(n38369), .Z(n10355) );
  AND U11294 ( .A(n10356), .B(n10355), .Z(n10628) );
  XOR U11295 ( .A(n10627), .B(n10628), .Z(n10630) );
  NANDN U11296 ( .A(n986), .B(b[63]), .Z(n10629) );
  XNOR U11297 ( .A(n10630), .B(n10629), .Z(n10541) );
  XOR U11298 ( .A(b[37]), .B(n17702), .Z(n10473) );
  NANDN U11299 ( .A(n10473), .B(n36311), .Z(n10359) );
  NANDN U11300 ( .A(n10357), .B(n36309), .Z(n10358) );
  NAND U11301 ( .A(n10359), .B(n10358), .Z(n10506) );
  XOR U11302 ( .A(b[5]), .B(n27436), .Z(n10476) );
  OR U11303 ( .A(n10476), .B(n29363), .Z(n10362) );
  NANDN U11304 ( .A(n10360), .B(n29864), .Z(n10361) );
  NAND U11305 ( .A(n10362), .B(n10361), .Z(n10503) );
  XOR U11306 ( .A(b[63]), .B(n10363), .Z(n10525) );
  NANDN U11307 ( .A(n10525), .B(n38422), .Z(n10366) );
  NAND U11308 ( .A(n10364), .B(n38423), .Z(n10365) );
  AND U11309 ( .A(n10366), .B(n10365), .Z(n10504) );
  XNOR U11310 ( .A(n10503), .B(n10504), .Z(n10505) );
  XOR U11311 ( .A(n10506), .B(n10505), .Z(n10540) );
  XOR U11312 ( .A(n10543), .B(n10542), .Z(n10654) );
  NANDN U11313 ( .A(n10368), .B(n10367), .Z(n10372) );
  NAND U11314 ( .A(n10370), .B(n10369), .Z(n10371) );
  NAND U11315 ( .A(n10372), .B(n10371), .Z(n10652) );
  NANDN U11316 ( .A(n10374), .B(n10373), .Z(n10378) );
  NAND U11317 ( .A(n10376), .B(n10375), .Z(n10377) );
  AND U11318 ( .A(n10378), .B(n10377), .Z(n10651) );
  XNOR U11319 ( .A(n10652), .B(n10651), .Z(n10653) );
  XOR U11320 ( .A(n10654), .B(n10653), .Z(n10702) );
  XOR U11321 ( .A(n10701), .B(n10702), .Z(n10687) );
  OR U11322 ( .A(n10380), .B(n10379), .Z(n10384) );
  OR U11323 ( .A(n10382), .B(n10381), .Z(n10383) );
  NAND U11324 ( .A(n10384), .B(n10383), .Z(n10666) );
  NANDN U11325 ( .A(n10386), .B(n10385), .Z(n10390) );
  NAND U11326 ( .A(n10388), .B(n10387), .Z(n10389) );
  NAND U11327 ( .A(n10390), .B(n10389), .Z(n10663) );
  NANDN U11328 ( .A(n10392), .B(n10391), .Z(n10396) );
  NAND U11329 ( .A(n10394), .B(n10393), .Z(n10395) );
  NAND U11330 ( .A(n10396), .B(n10395), .Z(n10664) );
  XNOR U11331 ( .A(n10663), .B(n10664), .Z(n10665) );
  XOR U11332 ( .A(n10666), .B(n10665), .Z(n10688) );
  XOR U11333 ( .A(n10687), .B(n10688), .Z(n10689) );
  XNOR U11334 ( .A(n10690), .B(n10689), .Z(n10433) );
  NANDN U11335 ( .A(n10398), .B(n10397), .Z(n10402) );
  NAND U11336 ( .A(n10400), .B(n10399), .Z(n10401) );
  AND U11337 ( .A(n10402), .B(n10401), .Z(n10434) );
  XNOR U11338 ( .A(n10433), .B(n10434), .Z(n10435) );
  XNOR U11339 ( .A(n10436), .B(n10435), .Z(n10675) );
  NANDN U11340 ( .A(n10404), .B(n10403), .Z(n10408) );
  NAND U11341 ( .A(n10406), .B(n10405), .Z(n10407) );
  AND U11342 ( .A(n10408), .B(n10407), .Z(n10676) );
  XNOR U11343 ( .A(n10675), .B(n10676), .Z(n10677) );
  XOR U11344 ( .A(n10678), .B(n10677), .Z(n10427) );
  NANDN U11345 ( .A(n10410), .B(n10409), .Z(n10414) );
  OR U11346 ( .A(n10412), .B(n10411), .Z(n10413) );
  AND U11347 ( .A(n10414), .B(n10413), .Z(n10428) );
  XNOR U11348 ( .A(n10427), .B(n10428), .Z(n10429) );
  NANDN U11349 ( .A(n10416), .B(n10415), .Z(n10420) );
  NANDN U11350 ( .A(n10418), .B(n10417), .Z(n10419) );
  NAND U11351 ( .A(n10420), .B(n10419), .Z(n10430) );
  XNOR U11352 ( .A(n10429), .B(n10430), .Z(n10422) );
  XNOR U11353 ( .A(n10421), .B(n10422), .Z(n10423) );
  XOR U11354 ( .A(n10424), .B(n10423), .Z(n10710) );
  XOR U11355 ( .A(n10711), .B(n10710), .Z(c[128]) );
  NANDN U11356 ( .A(n10422), .B(n10421), .Z(n10426) );
  NAND U11357 ( .A(n10424), .B(n10423), .Z(n10425) );
  NAND U11358 ( .A(n10426), .B(n10425), .Z(n10717) );
  NANDN U11359 ( .A(n10428), .B(n10427), .Z(n10432) );
  NANDN U11360 ( .A(n10430), .B(n10429), .Z(n10431) );
  NAND U11361 ( .A(n10432), .B(n10431), .Z(n10715) );
  NAND U11362 ( .A(n10434), .B(n10433), .Z(n10438) );
  OR U11363 ( .A(n10436), .B(n10435), .Z(n10437) );
  NAND U11364 ( .A(n10438), .B(n10437), .Z(n10725) );
  NANDN U11365 ( .A(n10440), .B(n10439), .Z(n10444) );
  NANDN U11366 ( .A(n10442), .B(n10441), .Z(n10443) );
  NAND U11367 ( .A(n10444), .B(n10443), .Z(n10745) );
  NANDN U11368 ( .A(n10446), .B(n10445), .Z(n10450) );
  NAND U11369 ( .A(n10448), .B(n10447), .Z(n10449) );
  NAND U11370 ( .A(n10450), .B(n10449), .Z(n10751) );
  NANDN U11371 ( .A(n10452), .B(n10451), .Z(n10456) );
  NAND U11372 ( .A(n10454), .B(n10453), .Z(n10455) );
  NAND U11373 ( .A(n10456), .B(n10455), .Z(n10896) );
  ANDN U11374 ( .B(b[63]), .A(n10457), .Z(n10910) );
  NANDN U11375 ( .A(n10458), .B(n38369), .Z(n10460) );
  XOR U11376 ( .A(b[61]), .B(n11202), .Z(n10806) );
  OR U11377 ( .A(n10806), .B(n38371), .Z(n10459) );
  NAND U11378 ( .A(n10460), .B(n10459), .Z(n10908) );
  NANDN U11379 ( .A(n10461), .B(n35311), .Z(n10463) );
  XOR U11380 ( .A(b[31]), .B(n20315), .Z(n10809) );
  NANDN U11381 ( .A(n10809), .B(n35313), .Z(n10462) );
  AND U11382 ( .A(n10463), .B(n10462), .Z(n10907) );
  XNOR U11383 ( .A(n10908), .B(n10907), .Z(n10909) );
  XOR U11384 ( .A(n10910), .B(n10909), .Z(n10894) );
  NAND U11385 ( .A(n33283), .B(n10464), .Z(n10466) );
  XOR U11386 ( .A(n33020), .B(n23149), .Z(n10812) );
  NANDN U11387 ( .A(n33021), .B(n10812), .Z(n10465) );
  NAND U11388 ( .A(n10466), .B(n10465), .Z(n10836) );
  XNOR U11389 ( .A(b[21]), .B(a[45]), .Z(n10815) );
  OR U11390 ( .A(n10815), .B(n33634), .Z(n10469) );
  NANDN U11391 ( .A(n10467), .B(n33464), .Z(n10468) );
  NAND U11392 ( .A(n10469), .B(n10468), .Z(n10833) );
  NAND U11393 ( .A(n34044), .B(n10470), .Z(n10472) );
  XOR U11394 ( .A(n34510), .B(n21996), .Z(n10818) );
  NANDN U11395 ( .A(n33867), .B(n10818), .Z(n10471) );
  AND U11396 ( .A(n10472), .B(n10471), .Z(n10834) );
  XNOR U11397 ( .A(n10833), .B(n10834), .Z(n10835) );
  XNOR U11398 ( .A(n10836), .B(n10835), .Z(n10895) );
  XNOR U11399 ( .A(n10894), .B(n10895), .Z(n10897) );
  XNOR U11400 ( .A(n10896), .B(n10897), .Z(n10749) );
  XOR U11401 ( .A(b[37]), .B(n18003), .Z(n10776) );
  NANDN U11402 ( .A(n10776), .B(n36311), .Z(n10475) );
  NANDN U11403 ( .A(n10473), .B(n36309), .Z(n10474) );
  NAND U11404 ( .A(n10475), .B(n10474), .Z(n10830) );
  XOR U11405 ( .A(b[5]), .B(n27773), .Z(n10779) );
  OR U11406 ( .A(n10779), .B(n29363), .Z(n10478) );
  NANDN U11407 ( .A(n10476), .B(n29864), .Z(n10477) );
  NAND U11408 ( .A(n10478), .B(n10477), .Z(n10827) );
  XNOR U11409 ( .A(n967), .B(a[63]), .Z(n10782) );
  NAND U11410 ( .A(n10782), .B(n28939), .Z(n10481) );
  NAND U11411 ( .A(n10479), .B(n28938), .Z(n10480) );
  AND U11412 ( .A(n10481), .B(n10480), .Z(n10828) );
  XNOR U11413 ( .A(n10827), .B(n10828), .Z(n10829) );
  XNOR U11414 ( .A(n10830), .B(n10829), .Z(n10757) );
  XOR U11415 ( .A(b[13]), .B(n25001), .Z(n10785) );
  OR U11416 ( .A(n10785), .B(n31550), .Z(n10484) );
  NANDN U11417 ( .A(n10482), .B(n31874), .Z(n10483) );
  NAND U11418 ( .A(n10484), .B(n10483), .Z(n10958) );
  NAND U11419 ( .A(n34848), .B(n10485), .Z(n10487) );
  XOR U11420 ( .A(n35375), .B(n20867), .Z(n10788) );
  NAND U11421 ( .A(n34618), .B(n10788), .Z(n10486) );
  NAND U11422 ( .A(n10487), .B(n10486), .Z(n10955) );
  NAND U11423 ( .A(n35188), .B(n10488), .Z(n10490) );
  XOR U11424 ( .A(n35540), .B(n20352), .Z(n10791) );
  NANDN U11425 ( .A(n34968), .B(n10791), .Z(n10489) );
  AND U11426 ( .A(n10490), .B(n10489), .Z(n10956) );
  XNOR U11427 ( .A(n10955), .B(n10956), .Z(n10957) );
  XNOR U11428 ( .A(n10958), .B(n10957), .Z(n10754) );
  NANDN U11429 ( .A(n10492), .B(n10491), .Z(n10496) );
  NAND U11430 ( .A(n10494), .B(n10493), .Z(n10495) );
  NAND U11431 ( .A(n10496), .B(n10495), .Z(n10755) );
  XNOR U11432 ( .A(n10754), .B(n10755), .Z(n10756) );
  XOR U11433 ( .A(n10757), .B(n10756), .Z(n10748) );
  XOR U11434 ( .A(n10749), .B(n10748), .Z(n10750) );
  XNOR U11435 ( .A(n10751), .B(n10750), .Z(n10867) );
  NANDN U11436 ( .A(n10498), .B(n10497), .Z(n10502) );
  NAND U11437 ( .A(n10500), .B(n10499), .Z(n10501) );
  NAND U11438 ( .A(n10502), .B(n10501), .Z(n10865) );
  NANDN U11439 ( .A(n10504), .B(n10503), .Z(n10508) );
  NAND U11440 ( .A(n10506), .B(n10505), .Z(n10507) );
  NAND U11441 ( .A(n10508), .B(n10507), .Z(n10761) );
  XNOR U11442 ( .A(b[41]), .B(a[25]), .Z(n10839) );
  OR U11443 ( .A(n10839), .B(n36905), .Z(n10511) );
  NANDN U11444 ( .A(n10509), .B(n36807), .Z(n10510) );
  NAND U11445 ( .A(n10511), .B(n10510), .Z(n10861) );
  XOR U11446 ( .A(b[57]), .B(n12258), .Z(n10842) );
  OR U11447 ( .A(n10842), .B(n965), .Z(n10514) );
  NANDN U11448 ( .A(n10512), .B(n38194), .Z(n10513) );
  NAND U11449 ( .A(n10514), .B(n10513), .Z(n10858) );
  NAND U11450 ( .A(n38326), .B(n10515), .Z(n10517) );
  XOR U11451 ( .A(n38400), .B(n11694), .Z(n10845) );
  NANDN U11452 ( .A(n38273), .B(n10845), .Z(n10516) );
  AND U11453 ( .A(n10517), .B(n10516), .Z(n10859) );
  XNOR U11454 ( .A(n10858), .B(n10859), .Z(n10860) );
  XOR U11455 ( .A(n10861), .B(n10860), .Z(n10925) );
  XOR U11456 ( .A(b[33]), .B(n19656), .Z(n10848) );
  NANDN U11457 ( .A(n10848), .B(n35620), .Z(n10520) );
  NANDN U11458 ( .A(n10518), .B(n35621), .Z(n10519) );
  NAND U11459 ( .A(n10520), .B(n10519), .Z(n10934) );
  NANDN U11460 ( .A(n966), .B(a[65]), .Z(n10521) );
  XOR U11461 ( .A(n29232), .B(n10521), .Z(n10523) );
  NANDN U11462 ( .A(b[0]), .B(a[64]), .Z(n10522) );
  AND U11463 ( .A(n10523), .B(n10522), .Z(n10931) );
  XOR U11464 ( .A(b[63]), .B(n10524), .Z(n10855) );
  NANDN U11465 ( .A(n10855), .B(n38422), .Z(n10527) );
  NANDN U11466 ( .A(n10525), .B(n38423), .Z(n10526) );
  AND U11467 ( .A(n10527), .B(n10526), .Z(n10932) );
  XNOR U11468 ( .A(n10931), .B(n10932), .Z(n10933) );
  XOR U11469 ( .A(n10934), .B(n10933), .Z(n10926) );
  XNOR U11470 ( .A(n10925), .B(n10926), .Z(n10928) );
  NANDN U11471 ( .A(n10529), .B(n10528), .Z(n10533) );
  NAND U11472 ( .A(n10531), .B(n10530), .Z(n10532) );
  NAND U11473 ( .A(n10533), .B(n10532), .Z(n10927) );
  XOR U11474 ( .A(n10928), .B(n10927), .Z(n10758) );
  NANDN U11475 ( .A(n10535), .B(n10534), .Z(n10539) );
  NAND U11476 ( .A(n10537), .B(n10536), .Z(n10538) );
  AND U11477 ( .A(n10539), .B(n10538), .Z(n10759) );
  XOR U11478 ( .A(n10758), .B(n10759), .Z(n10760) );
  XNOR U11479 ( .A(n10761), .B(n10760), .Z(n10864) );
  XNOR U11480 ( .A(n10865), .B(n10864), .Z(n10866) );
  XNOR U11481 ( .A(n10867), .B(n10866), .Z(n10742) );
  NANDN U11482 ( .A(n10541), .B(n10540), .Z(n10545) );
  NANDN U11483 ( .A(n10543), .B(n10542), .Z(n10544) );
  NAND U11484 ( .A(n10545), .B(n10544), .Z(n10986) );
  NANDN U11485 ( .A(n10547), .B(n10546), .Z(n10551) );
  NANDN U11486 ( .A(n10549), .B(n10548), .Z(n10550) );
  AND U11487 ( .A(n10551), .B(n10550), .Z(n10985) );
  XNOR U11488 ( .A(n10986), .B(n10985), .Z(n10988) );
  NANDN U11489 ( .A(n10553), .B(n10552), .Z(n10557) );
  NAND U11490 ( .A(n10555), .B(n10554), .Z(n10556) );
  NAND U11491 ( .A(n10557), .B(n10556), .Z(n10921) );
  NANDN U11492 ( .A(n10559), .B(n10558), .Z(n10563) );
  NAND U11493 ( .A(n10561), .B(n10560), .Z(n10562) );
  NAND U11494 ( .A(n10563), .B(n10562), .Z(n10824) );
  XOR U11495 ( .A(b[15]), .B(n24288), .Z(n10937) );
  OR U11496 ( .A(n10937), .B(n32010), .Z(n10566) );
  NANDN U11497 ( .A(n10564), .B(n32011), .Z(n10565) );
  NAND U11498 ( .A(n10566), .B(n10565), .Z(n10803) );
  XNOR U11499 ( .A(b[25]), .B(n21441), .Z(n10940) );
  NANDN U11500 ( .A(n34219), .B(n10940), .Z(n10569) );
  NAND U11501 ( .A(n34217), .B(n10567), .Z(n10568) );
  NAND U11502 ( .A(n10569), .B(n10568), .Z(n10800) );
  XNOR U11503 ( .A(b[17]), .B(a[49]), .Z(n10943) );
  NANDN U11504 ( .A(n10943), .B(n32543), .Z(n10572) );
  NANDN U11505 ( .A(n10570), .B(n32541), .Z(n10571) );
  AND U11506 ( .A(n10572), .B(n10571), .Z(n10801) );
  XNOR U11507 ( .A(n10800), .B(n10801), .Z(n10802) );
  XNOR U11508 ( .A(n10803), .B(n10802), .Z(n10821) );
  XOR U11509 ( .A(b[39]), .B(n17960), .Z(n10946) );
  NANDN U11510 ( .A(n10946), .B(n36553), .Z(n10575) );
  NANDN U11511 ( .A(n10573), .B(n36643), .Z(n10574) );
  NAND U11512 ( .A(n10575), .B(n10574), .Z(n10797) );
  XOR U11513 ( .A(b[51]), .B(n13976), .Z(n10949) );
  NANDN U11514 ( .A(n10949), .B(n37803), .Z(n10578) );
  NANDN U11515 ( .A(n10576), .B(n37802), .Z(n10577) );
  NAND U11516 ( .A(n10578), .B(n10577), .Z(n10794) );
  XOR U11517 ( .A(b[53]), .B(n13509), .Z(n10952) );
  NANDN U11518 ( .A(n10952), .B(n37940), .Z(n10581) );
  NANDN U11519 ( .A(n10579), .B(n37941), .Z(n10580) );
  AND U11520 ( .A(n10581), .B(n10580), .Z(n10795) );
  XNOR U11521 ( .A(n10794), .B(n10795), .Z(n10796) );
  XOR U11522 ( .A(n10797), .B(n10796), .Z(n10822) );
  XNOR U11523 ( .A(n10821), .B(n10822), .Z(n10823) );
  XNOR U11524 ( .A(n10824), .B(n10823), .Z(n10919) );
  NANDN U11525 ( .A(n10583), .B(n10582), .Z(n10587) );
  NAND U11526 ( .A(n10585), .B(n10584), .Z(n10586) );
  AND U11527 ( .A(n10587), .B(n10586), .Z(n10920) );
  XNOR U11528 ( .A(n10919), .B(n10920), .Z(n10922) );
  XNOR U11529 ( .A(n10921), .B(n10922), .Z(n10987) );
  XOR U11530 ( .A(n10988), .B(n10987), .Z(n10743) );
  XNOR U11531 ( .A(n10742), .B(n10743), .Z(n10744) );
  XOR U11532 ( .A(n10745), .B(n10744), .Z(n10733) );
  OR U11533 ( .A(n10589), .B(n10588), .Z(n10593) );
  OR U11534 ( .A(n10591), .B(n10590), .Z(n10592) );
  NAND U11535 ( .A(n10593), .B(n10592), .Z(n10973) );
  XOR U11536 ( .A(b[11]), .B(n25466), .Z(n10870) );
  OR U11537 ( .A(n10870), .B(n31369), .Z(n10596) );
  NANDN U11538 ( .A(n10594), .B(n31119), .Z(n10595) );
  NAND U11539 ( .A(n10596), .B(n10595), .Z(n10891) );
  XOR U11540 ( .A(b[43]), .B(n16269), .Z(n10873) );
  NANDN U11541 ( .A(n10873), .B(n37068), .Z(n10599) );
  NANDN U11542 ( .A(n10597), .B(n37069), .Z(n10598) );
  NAND U11543 ( .A(n10599), .B(n10598), .Z(n10888) );
  XNOR U11544 ( .A(b[45]), .B(a[21]), .Z(n10876) );
  NANDN U11545 ( .A(n10876), .B(n37261), .Z(n10602) );
  NANDN U11546 ( .A(n10600), .B(n37262), .Z(n10601) );
  AND U11547 ( .A(n10602), .B(n10601), .Z(n10889) );
  XNOR U11548 ( .A(n10888), .B(n10889), .Z(n10890) );
  XNOR U11549 ( .A(n10891), .B(n10890), .Z(n10770) );
  NAND U11550 ( .A(n37652), .B(n10603), .Z(n10605) );
  XOR U11551 ( .A(n979), .B(a[17]), .Z(n10879) );
  OR U11552 ( .A(n10879), .B(n37756), .Z(n10604) );
  NAND U11553 ( .A(n10605), .B(n10604), .Z(n10915) );
  NANDN U11554 ( .A(n10606), .B(n37469), .Z(n10608) );
  XOR U11555 ( .A(b[47]), .B(n15113), .Z(n10882) );
  NANDN U11556 ( .A(n10882), .B(n37471), .Z(n10607) );
  AND U11557 ( .A(n10608), .B(n10607), .Z(n10914) );
  NAND U11558 ( .A(n30846), .B(n10609), .Z(n10611) );
  XOR U11559 ( .A(n969), .B(n26122), .Z(n10885) );
  NAND U11560 ( .A(n30509), .B(n10885), .Z(n10610) );
  NAND U11561 ( .A(n10611), .B(n10610), .Z(n10913) );
  XNOR U11562 ( .A(n10914), .B(n10913), .Z(n10916) );
  XOR U11563 ( .A(n10915), .B(n10916), .Z(n10771) );
  XNOR U11564 ( .A(n10770), .B(n10771), .Z(n10772) );
  NANDN U11565 ( .A(n10613), .B(n10612), .Z(n10617) );
  NAND U11566 ( .A(n10615), .B(n10614), .Z(n10616) );
  AND U11567 ( .A(n10617), .B(n10616), .Z(n10773) );
  XNOR U11568 ( .A(n10772), .B(n10773), .Z(n10974) );
  XNOR U11569 ( .A(n10973), .B(n10974), .Z(n10975) );
  XNOR U11570 ( .A(b[35]), .B(a[31]), .Z(n10898) );
  NANDN U11571 ( .A(n10898), .B(n35985), .Z(n10620) );
  NANDN U11572 ( .A(n10618), .B(n35986), .Z(n10619) );
  NAND U11573 ( .A(n10620), .B(n10619), .Z(n10964) );
  XNOR U11574 ( .A(n31123), .B(a[59]), .Z(n10901) );
  NAND U11575 ( .A(n10901), .B(n29949), .Z(n10623) );
  NAND U11576 ( .A(n29948), .B(n10621), .Z(n10622) );
  NAND U11577 ( .A(n10623), .B(n10622), .Z(n10961) );
  XOR U11578 ( .A(b[55]), .B(n12830), .Z(n10904) );
  NANDN U11579 ( .A(n10904), .B(n38075), .Z(n10626) );
  NANDN U11580 ( .A(n10624), .B(n38073), .Z(n10625) );
  AND U11581 ( .A(n10626), .B(n10625), .Z(n10962) );
  XNOR U11582 ( .A(n10961), .B(n10962), .Z(n10963) );
  XNOR U11583 ( .A(n10964), .B(n10963), .Z(n10767) );
  NANDN U11584 ( .A(n10628), .B(n10627), .Z(n10632) );
  OR U11585 ( .A(n10630), .B(n10629), .Z(n10631) );
  NAND U11586 ( .A(n10632), .B(n10631), .Z(n10765) );
  NANDN U11587 ( .A(n10634), .B(n10633), .Z(n10638) );
  NAND U11588 ( .A(n10636), .B(n10635), .Z(n10637) );
  AND U11589 ( .A(n10638), .B(n10637), .Z(n10764) );
  XNOR U11590 ( .A(n10765), .B(n10764), .Z(n10766) );
  XOR U11591 ( .A(n10767), .B(n10766), .Z(n10976) );
  XOR U11592 ( .A(n10975), .B(n10976), .Z(n10730) );
  NANDN U11593 ( .A(n10640), .B(n10639), .Z(n10644) );
  OR U11594 ( .A(n10642), .B(n10641), .Z(n10643) );
  NAND U11595 ( .A(n10644), .B(n10643), .Z(n10982) );
  NANDN U11596 ( .A(n10646), .B(n10645), .Z(n10650) );
  NANDN U11597 ( .A(n10648), .B(n10647), .Z(n10649) );
  NAND U11598 ( .A(n10650), .B(n10649), .Z(n10979) );
  NANDN U11599 ( .A(n10652), .B(n10651), .Z(n10656) );
  NAND U11600 ( .A(n10654), .B(n10653), .Z(n10655) );
  AND U11601 ( .A(n10656), .B(n10655), .Z(n10980) );
  XNOR U11602 ( .A(n10979), .B(n10980), .Z(n10981) );
  XNOR U11603 ( .A(n10982), .B(n10981), .Z(n10731) );
  XNOR U11604 ( .A(n10730), .B(n10731), .Z(n10732) );
  XOR U11605 ( .A(n10733), .B(n10732), .Z(n10739) );
  NANDN U11606 ( .A(n10658), .B(n10657), .Z(n10662) );
  NAND U11607 ( .A(n10660), .B(n10659), .Z(n10661) );
  NAND U11608 ( .A(n10662), .B(n10661), .Z(n10736) );
  NANDN U11609 ( .A(n10664), .B(n10663), .Z(n10668) );
  NAND U11610 ( .A(n10666), .B(n10665), .Z(n10667) );
  NAND U11611 ( .A(n10668), .B(n10667), .Z(n10737) );
  XNOR U11612 ( .A(n10736), .B(n10737), .Z(n10738) );
  XNOR U11613 ( .A(n10739), .B(n10738), .Z(n10724) );
  XNOR U11614 ( .A(n10725), .B(n10724), .Z(n10727) );
  NANDN U11615 ( .A(n10670), .B(n10669), .Z(n10674) );
  NAND U11616 ( .A(n10672), .B(n10671), .Z(n10673) );
  NAND U11617 ( .A(n10674), .B(n10673), .Z(n10726) );
  XNOR U11618 ( .A(n10727), .B(n10726), .Z(n10720) );
  NANDN U11619 ( .A(n10676), .B(n10675), .Z(n10680) );
  NANDN U11620 ( .A(n10678), .B(n10677), .Z(n10679) );
  NAND U11621 ( .A(n10680), .B(n10679), .Z(n10719) );
  NANDN U11622 ( .A(n10682), .B(n10681), .Z(n10686) );
  NANDN U11623 ( .A(n10684), .B(n10683), .Z(n10685) );
  NAND U11624 ( .A(n10686), .B(n10685), .Z(n10992) );
  OR U11625 ( .A(n10688), .B(n10687), .Z(n10692) );
  NANDN U11626 ( .A(n10690), .B(n10689), .Z(n10691) );
  NAND U11627 ( .A(n10692), .B(n10691), .Z(n10989) );
  OR U11628 ( .A(n10694), .B(n10693), .Z(n10698) );
  OR U11629 ( .A(n10696), .B(n10695), .Z(n10697) );
  NAND U11630 ( .A(n10698), .B(n10697), .Z(n10970) );
  OR U11631 ( .A(n10704), .B(n10703), .Z(n10708) );
  NANDN U11632 ( .A(n10706), .B(n10705), .Z(n10707) );
  AND U11633 ( .A(n10708), .B(n10707), .Z(n10968) );
  XNOR U11634 ( .A(n10967), .B(n10968), .Z(n10969) );
  XOR U11635 ( .A(n10970), .B(n10969), .Z(n10990) );
  XOR U11636 ( .A(n10989), .B(n10990), .Z(n10991) );
  XNOR U11637 ( .A(n10992), .B(n10991), .Z(n10718) );
  XNOR U11638 ( .A(n10719), .B(n10718), .Z(n10721) );
  XNOR U11639 ( .A(n10720), .B(n10721), .Z(n10714) );
  XNOR U11640 ( .A(n10715), .B(n10714), .Z(n10716) );
  XNOR U11641 ( .A(n10717), .B(n10716), .Z(n10995) );
  XNOR U11642 ( .A(n10995), .B(sreg[129]), .Z(n10997) );
  NAND U11643 ( .A(n10709), .B(sreg[128]), .Z(n10713) );
  OR U11644 ( .A(n10711), .B(n10710), .Z(n10712) );
  AND U11645 ( .A(n10713), .B(n10712), .Z(n10996) );
  XOR U11646 ( .A(n10997), .B(n10996), .Z(c[129]) );
  NAND U11647 ( .A(n10719), .B(n10718), .Z(n10723) );
  NANDN U11648 ( .A(n10721), .B(n10720), .Z(n10722) );
  NAND U11649 ( .A(n10723), .B(n10722), .Z(n11000) );
  NAND U11650 ( .A(n10725), .B(n10724), .Z(n10729) );
  OR U11651 ( .A(n10727), .B(n10726), .Z(n10728) );
  NAND U11652 ( .A(n10729), .B(n10728), .Z(n11278) );
  NANDN U11653 ( .A(n10731), .B(n10730), .Z(n10735) );
  NAND U11654 ( .A(n10733), .B(n10732), .Z(n10734) );
  NAND U11655 ( .A(n10735), .B(n10734), .Z(n11269) );
  NANDN U11656 ( .A(n10737), .B(n10736), .Z(n10741) );
  NANDN U11657 ( .A(n10739), .B(n10738), .Z(n10740) );
  NAND U11658 ( .A(n10741), .B(n10740), .Z(n11270) );
  XNOR U11659 ( .A(n11269), .B(n11270), .Z(n11271) );
  NANDN U11660 ( .A(n10743), .B(n10742), .Z(n10747) );
  NANDN U11661 ( .A(n10745), .B(n10744), .Z(n10746) );
  NAND U11662 ( .A(n10747), .B(n10746), .Z(n11260) );
  NAND U11663 ( .A(n10749), .B(n10748), .Z(n10753) );
  NAND U11664 ( .A(n10751), .B(n10750), .Z(n10752) );
  NAND U11665 ( .A(n10753), .B(n10752), .Z(n11246) );
  NAND U11666 ( .A(n10759), .B(n10758), .Z(n10763) );
  NANDN U11667 ( .A(n10761), .B(n10760), .Z(n10762) );
  NAND U11668 ( .A(n10763), .B(n10762), .Z(n11012) );
  NANDN U11669 ( .A(n10765), .B(n10764), .Z(n10769) );
  NAND U11670 ( .A(n10767), .B(n10766), .Z(n10768) );
  AND U11671 ( .A(n10769), .B(n10768), .Z(n11013) );
  XNOR U11672 ( .A(n11012), .B(n11013), .Z(n11014) );
  XNOR U11673 ( .A(n11015), .B(n11014), .Z(n11245) );
  XNOR U11674 ( .A(n11246), .B(n11245), .Z(n11248) );
  NANDN U11675 ( .A(n10771), .B(n10770), .Z(n10775) );
  NAND U11676 ( .A(n10773), .B(n10772), .Z(n10774) );
  NAND U11677 ( .A(n10775), .B(n10774), .Z(n11241) );
  XOR U11678 ( .A(b[37]), .B(n18804), .Z(n11151) );
  NANDN U11679 ( .A(n11151), .B(n36311), .Z(n10778) );
  NANDN U11680 ( .A(n10776), .B(n36309), .Z(n10777) );
  NAND U11681 ( .A(n10778), .B(n10777), .Z(n11230) );
  XNOR U11682 ( .A(b[5]), .B(a[62]), .Z(n11154) );
  OR U11683 ( .A(n11154), .B(n29363), .Z(n10781) );
  NANDN U11684 ( .A(n10779), .B(n29864), .Z(n10780) );
  NAND U11685 ( .A(n10781), .B(n10780), .Z(n11227) );
  XNOR U11686 ( .A(n967), .B(a[64]), .Z(n11157) );
  NAND U11687 ( .A(n11157), .B(n28939), .Z(n10784) );
  NAND U11688 ( .A(n28938), .B(n10782), .Z(n10783) );
  AND U11689 ( .A(n10784), .B(n10783), .Z(n11228) );
  XNOR U11690 ( .A(n11227), .B(n11228), .Z(n11229) );
  XOR U11691 ( .A(n11230), .B(n11229), .Z(n11142) );
  XOR U11692 ( .A(b[13]), .B(n25177), .Z(n11160) );
  OR U11693 ( .A(n11160), .B(n31550), .Z(n10787) );
  NANDN U11694 ( .A(n10785), .B(n31874), .Z(n10786) );
  NAND U11695 ( .A(n10787), .B(n10786), .Z(n11102) );
  NAND U11696 ( .A(n34848), .B(n10788), .Z(n10790) );
  XOR U11697 ( .A(n35375), .B(n21149), .Z(n11163) );
  NAND U11698 ( .A(n34618), .B(n11163), .Z(n10789) );
  NAND U11699 ( .A(n10790), .B(n10789), .Z(n11099) );
  NAND U11700 ( .A(n35188), .B(n10791), .Z(n10793) );
  XOR U11701 ( .A(n35540), .B(n20686), .Z(n11166) );
  NANDN U11702 ( .A(n34968), .B(n11166), .Z(n10792) );
  AND U11703 ( .A(n10793), .B(n10792), .Z(n11100) );
  XNOR U11704 ( .A(n11099), .B(n11100), .Z(n11101) );
  XOR U11705 ( .A(n11102), .B(n11101), .Z(n11140) );
  NANDN U11706 ( .A(n10795), .B(n10794), .Z(n10799) );
  NAND U11707 ( .A(n10797), .B(n10796), .Z(n10798) );
  AND U11708 ( .A(n10799), .B(n10798), .Z(n11139) );
  XOR U11709 ( .A(n11140), .B(n11139), .Z(n11141) );
  XOR U11710 ( .A(n11142), .B(n11141), .Z(n11240) );
  NANDN U11711 ( .A(n10801), .B(n10800), .Z(n10805) );
  NAND U11712 ( .A(n10803), .B(n10802), .Z(n10804) );
  NAND U11713 ( .A(n10805), .B(n10804), .Z(n11054) );
  NAND U11714 ( .A(a[2]), .B(b[63]), .Z(n11068) );
  NANDN U11715 ( .A(n10806), .B(n38369), .Z(n10808) );
  XOR U11716 ( .A(b[61]), .B(n11406), .Z(n11181) );
  OR U11717 ( .A(n11181), .B(n38371), .Z(n10807) );
  NAND U11718 ( .A(n10808), .B(n10807), .Z(n11066) );
  NANDN U11719 ( .A(n10809), .B(n35311), .Z(n10811) );
  XOR U11720 ( .A(b[31]), .B(n19980), .Z(n11184) );
  NANDN U11721 ( .A(n11184), .B(n35313), .Z(n10810) );
  AND U11722 ( .A(n10811), .B(n10810), .Z(n11065) );
  XNOR U11723 ( .A(n11066), .B(n11065), .Z(n11067) );
  XOR U11724 ( .A(n11068), .B(n11067), .Z(n11052) );
  NAND U11725 ( .A(n33283), .B(n10812), .Z(n10814) );
  XOR U11726 ( .A(n33020), .B(n23447), .Z(n11187) );
  NANDN U11727 ( .A(n33021), .B(n11187), .Z(n10813) );
  NAND U11728 ( .A(n10814), .B(n10813), .Z(n11218) );
  XNOR U11729 ( .A(b[21]), .B(a[46]), .Z(n11190) );
  OR U11730 ( .A(n11190), .B(n33634), .Z(n10817) );
  NANDN U11731 ( .A(n10815), .B(n33464), .Z(n10816) );
  NAND U11732 ( .A(n10817), .B(n10816), .Z(n11215) );
  NAND U11733 ( .A(n34044), .B(n10818), .Z(n10820) );
  XOR U11734 ( .A(n34510), .B(n22289), .Z(n11193) );
  NANDN U11735 ( .A(n33867), .B(n11193), .Z(n10819) );
  AND U11736 ( .A(n10820), .B(n10819), .Z(n11216) );
  XNOR U11737 ( .A(n11215), .B(n11216), .Z(n11217) );
  XNOR U11738 ( .A(n11218), .B(n11217), .Z(n11053) );
  XNOR U11739 ( .A(n11052), .B(n11053), .Z(n11055) );
  XNOR U11740 ( .A(n11054), .B(n11055), .Z(n11239) );
  XOR U11741 ( .A(n11240), .B(n11239), .Z(n11242) );
  XNOR U11742 ( .A(n11241), .B(n11242), .Z(n11123) );
  NANDN U11743 ( .A(n10822), .B(n10821), .Z(n10826) );
  NANDN U11744 ( .A(n10824), .B(n10823), .Z(n10825) );
  NAND U11745 ( .A(n10826), .B(n10825), .Z(n11122) );
  NANDN U11746 ( .A(n10828), .B(n10827), .Z(n10832) );
  NAND U11747 ( .A(n10830), .B(n10829), .Z(n10831) );
  NAND U11748 ( .A(n10832), .B(n10831), .Z(n11136) );
  NANDN U11749 ( .A(n10834), .B(n10833), .Z(n10838) );
  NAND U11750 ( .A(n10836), .B(n10835), .Z(n10837) );
  NAND U11751 ( .A(n10838), .B(n10837), .Z(n11118) );
  XNOR U11752 ( .A(b[41]), .B(a[26]), .Z(n11206) );
  OR U11753 ( .A(n11206), .B(n36905), .Z(n10841) );
  NANDN U11754 ( .A(n10839), .B(n36807), .Z(n10840) );
  NAND U11755 ( .A(n10841), .B(n10840), .Z(n11224) );
  XOR U11756 ( .A(b[57]), .B(n12555), .Z(n11209) );
  OR U11757 ( .A(n11209), .B(n965), .Z(n10844) );
  NANDN U11758 ( .A(n10842), .B(n38194), .Z(n10843) );
  NAND U11759 ( .A(n10844), .B(n10843), .Z(n11221) );
  NAND U11760 ( .A(n38326), .B(n10845), .Z(n10847) );
  XOR U11761 ( .A(n38400), .B(n11986), .Z(n11212) );
  NANDN U11762 ( .A(n38273), .B(n11212), .Z(n10846) );
  AND U11763 ( .A(n10847), .B(n10846), .Z(n11222) );
  XNOR U11764 ( .A(n11221), .B(n11222), .Z(n11223) );
  XOR U11765 ( .A(n11224), .B(n11223), .Z(n11116) );
  XOR U11766 ( .A(b[33]), .B(n19513), .Z(n11196) );
  NANDN U11767 ( .A(n11196), .B(n35620), .Z(n10850) );
  NANDN U11768 ( .A(n10848), .B(n35621), .Z(n10849) );
  NAND U11769 ( .A(n10850), .B(n10849), .Z(n11114) );
  NANDN U11770 ( .A(n966), .B(a[66]), .Z(n10851) );
  XOR U11771 ( .A(n29232), .B(n10851), .Z(n10853) );
  IV U11772 ( .A(a[65]), .Z(n28403) );
  NANDN U11773 ( .A(n28403), .B(n966), .Z(n10852) );
  AND U11774 ( .A(n10853), .B(n10852), .Z(n11111) );
  XOR U11775 ( .A(b[63]), .B(n10854), .Z(n11203) );
  NANDN U11776 ( .A(n11203), .B(n38422), .Z(n10857) );
  NANDN U11777 ( .A(n10855), .B(n38423), .Z(n10856) );
  AND U11778 ( .A(n10857), .B(n10856), .Z(n11112) );
  XNOR U11779 ( .A(n11111), .B(n11112), .Z(n11113) );
  XNOR U11780 ( .A(n11114), .B(n11113), .Z(n11115) );
  XOR U11781 ( .A(n11116), .B(n11115), .Z(n11117) );
  XNOR U11782 ( .A(n11118), .B(n11117), .Z(n11134) );
  NANDN U11783 ( .A(n10859), .B(n10858), .Z(n10863) );
  NAND U11784 ( .A(n10861), .B(n10860), .Z(n10862) );
  AND U11785 ( .A(n10863), .B(n10862), .Z(n11133) );
  XNOR U11786 ( .A(n11134), .B(n11133), .Z(n11135) );
  XNOR U11787 ( .A(n11136), .B(n11135), .Z(n11121) );
  XNOR U11788 ( .A(n11122), .B(n11121), .Z(n11124) );
  XNOR U11789 ( .A(n11123), .B(n11124), .Z(n11247) );
  XOR U11790 ( .A(n11248), .B(n11247), .Z(n11257) );
  NAND U11791 ( .A(n10865), .B(n10864), .Z(n10869) );
  OR U11792 ( .A(n10867), .B(n10866), .Z(n10868) );
  NAND U11793 ( .A(n10869), .B(n10868), .Z(n11025) );
  XOR U11794 ( .A(b[11]), .B(n25860), .Z(n11028) );
  OR U11795 ( .A(n11028), .B(n31369), .Z(n10872) );
  NANDN U11796 ( .A(n10870), .B(n31119), .Z(n10871) );
  NAND U11797 ( .A(n10872), .B(n10871), .Z(n11049) );
  XOR U11798 ( .A(b[43]), .B(n16508), .Z(n11031) );
  NANDN U11799 ( .A(n11031), .B(n37068), .Z(n10875) );
  NANDN U11800 ( .A(n10873), .B(n37069), .Z(n10874) );
  NAND U11801 ( .A(n10875), .B(n10874), .Z(n11046) );
  XNOR U11802 ( .A(b[45]), .B(a[22]), .Z(n11034) );
  NANDN U11803 ( .A(n11034), .B(n37261), .Z(n10878) );
  NANDN U11804 ( .A(n10876), .B(n37262), .Z(n10877) );
  AND U11805 ( .A(n10878), .B(n10877), .Z(n11047) );
  XNOR U11806 ( .A(n11046), .B(n11047), .Z(n11048) );
  XNOR U11807 ( .A(n11049), .B(n11048), .Z(n11148) );
  NANDN U11808 ( .A(n10879), .B(n37652), .Z(n10881) );
  XOR U11809 ( .A(b[49]), .B(n14905), .Z(n11037) );
  OR U11810 ( .A(n11037), .B(n37756), .Z(n10880) );
  NAND U11811 ( .A(n10881), .B(n10880), .Z(n11073) );
  NANDN U11812 ( .A(n10882), .B(n37469), .Z(n10884) );
  XNOR U11813 ( .A(n978), .B(a[20]), .Z(n11040) );
  NAND U11814 ( .A(n11040), .B(n37471), .Z(n10883) );
  NAND U11815 ( .A(n10884), .B(n10883), .Z(n11071) );
  NAND U11816 ( .A(n30846), .B(n10885), .Z(n10887) );
  XNOR U11817 ( .A(n969), .B(a[58]), .Z(n11043) );
  NAND U11818 ( .A(n30509), .B(n11043), .Z(n10886) );
  NAND U11819 ( .A(n10887), .B(n10886), .Z(n11072) );
  XNOR U11820 ( .A(n11071), .B(n11072), .Z(n11074) );
  XOR U11821 ( .A(n11073), .B(n11074), .Z(n11145) );
  NANDN U11822 ( .A(n10889), .B(n10888), .Z(n10893) );
  NAND U11823 ( .A(n10891), .B(n10890), .Z(n10892) );
  NAND U11824 ( .A(n10893), .B(n10892), .Z(n11146) );
  XNOR U11825 ( .A(n11145), .B(n11146), .Z(n11147) );
  XOR U11826 ( .A(n11148), .B(n11147), .Z(n11006) );
  XNOR U11827 ( .A(n11006), .B(n11007), .Z(n11009) );
  XNOR U11828 ( .A(b[35]), .B(a[32]), .Z(n11056) );
  NANDN U11829 ( .A(n11056), .B(n35985), .Z(n10900) );
  NANDN U11830 ( .A(n10898), .B(n35986), .Z(n10899) );
  NAND U11831 ( .A(n10900), .B(n10899), .Z(n11108) );
  XOR U11832 ( .A(n31123), .B(n27436), .Z(n11059) );
  NAND U11833 ( .A(n11059), .B(n29949), .Z(n10903) );
  NAND U11834 ( .A(n29948), .B(n10901), .Z(n10902) );
  NAND U11835 ( .A(n10903), .B(n10902), .Z(n11105) );
  XOR U11836 ( .A(b[55]), .B(n13106), .Z(n11062) );
  NANDN U11837 ( .A(n11062), .B(n38075), .Z(n10906) );
  NANDN U11838 ( .A(n10904), .B(n38073), .Z(n10905) );
  AND U11839 ( .A(n10906), .B(n10905), .Z(n11106) );
  XNOR U11840 ( .A(n11105), .B(n11106), .Z(n11107) );
  XNOR U11841 ( .A(n11108), .B(n11107), .Z(n11130) );
  NANDN U11842 ( .A(n10908), .B(n10907), .Z(n10912) );
  NANDN U11843 ( .A(n10910), .B(n10909), .Z(n10911) );
  NAND U11844 ( .A(n10912), .B(n10911), .Z(n11127) );
  NANDN U11845 ( .A(n10914), .B(n10913), .Z(n10918) );
  NAND U11846 ( .A(n10916), .B(n10915), .Z(n10917) );
  NAND U11847 ( .A(n10918), .B(n10917), .Z(n11128) );
  XNOR U11848 ( .A(n11127), .B(n11128), .Z(n11129) );
  XOR U11849 ( .A(n11130), .B(n11129), .Z(n11008) );
  XOR U11850 ( .A(n11009), .B(n11008), .Z(n11023) );
  NAND U11851 ( .A(n10920), .B(n10919), .Z(n10924) );
  NANDN U11852 ( .A(n10922), .B(n10921), .Z(n10923) );
  NAND U11853 ( .A(n10924), .B(n10923), .Z(n11016) );
  OR U11854 ( .A(n10926), .B(n10925), .Z(n10930) );
  OR U11855 ( .A(n10928), .B(n10927), .Z(n10929) );
  AND U11856 ( .A(n10930), .B(n10929), .Z(n11017) );
  XNOR U11857 ( .A(n11016), .B(n11017), .Z(n11018) );
  NANDN U11858 ( .A(n10932), .B(n10931), .Z(n10936) );
  NAND U11859 ( .A(n10934), .B(n10933), .Z(n10935) );
  NAND U11860 ( .A(n10936), .B(n10935), .Z(n11078) );
  XOR U11861 ( .A(b[15]), .B(n25134), .Z(n11081) );
  OR U11862 ( .A(n11081), .B(n32010), .Z(n10939) );
  NANDN U11863 ( .A(n10937), .B(n32011), .Z(n10938) );
  NAND U11864 ( .A(n10939), .B(n10938), .Z(n11178) );
  XNOR U11865 ( .A(b[25]), .B(n22246), .Z(n11084) );
  NANDN U11866 ( .A(n34219), .B(n11084), .Z(n10942) );
  NAND U11867 ( .A(n34217), .B(n10940), .Z(n10941) );
  NAND U11868 ( .A(n10942), .B(n10941), .Z(n11175) );
  XNOR U11869 ( .A(b[17]), .B(a[50]), .Z(n11087) );
  NANDN U11870 ( .A(n11087), .B(n32543), .Z(n10945) );
  NANDN U11871 ( .A(n10943), .B(n32541), .Z(n10944) );
  AND U11872 ( .A(n10945), .B(n10944), .Z(n11176) );
  XNOR U11873 ( .A(n11175), .B(n11176), .Z(n11177) );
  XNOR U11874 ( .A(n11178), .B(n11177), .Z(n11233) );
  XOR U11875 ( .A(b[39]), .B(n17702), .Z(n11090) );
  NANDN U11876 ( .A(n11090), .B(n36553), .Z(n10948) );
  NANDN U11877 ( .A(n10946), .B(n36643), .Z(n10947) );
  NAND U11878 ( .A(n10948), .B(n10947), .Z(n11172) );
  XOR U11879 ( .A(b[51]), .B(n14259), .Z(n11093) );
  NANDN U11880 ( .A(n11093), .B(n37803), .Z(n10951) );
  NANDN U11881 ( .A(n10949), .B(n37802), .Z(n10950) );
  NAND U11882 ( .A(n10951), .B(n10950), .Z(n11169) );
  XOR U11883 ( .A(b[53]), .B(n14210), .Z(n11096) );
  NANDN U11884 ( .A(n11096), .B(n37940), .Z(n10954) );
  NANDN U11885 ( .A(n10952), .B(n37941), .Z(n10953) );
  AND U11886 ( .A(n10954), .B(n10953), .Z(n11170) );
  XNOR U11887 ( .A(n11169), .B(n11170), .Z(n11171) );
  XOR U11888 ( .A(n11172), .B(n11171), .Z(n11234) );
  XOR U11889 ( .A(n11233), .B(n11234), .Z(n11236) );
  NANDN U11890 ( .A(n10956), .B(n10955), .Z(n10960) );
  NAND U11891 ( .A(n10958), .B(n10957), .Z(n10959) );
  AND U11892 ( .A(n10960), .B(n10959), .Z(n11235) );
  XOR U11893 ( .A(n11236), .B(n11235), .Z(n11076) );
  NANDN U11894 ( .A(n10962), .B(n10961), .Z(n10966) );
  NAND U11895 ( .A(n10964), .B(n10963), .Z(n10965) );
  AND U11896 ( .A(n10966), .B(n10965), .Z(n11075) );
  XNOR U11897 ( .A(n11076), .B(n11075), .Z(n11077) );
  XOR U11898 ( .A(n11078), .B(n11077), .Z(n11019) );
  XNOR U11899 ( .A(n11018), .B(n11019), .Z(n11022) );
  XNOR U11900 ( .A(n11023), .B(n11022), .Z(n11024) );
  XOR U11901 ( .A(n11025), .B(n11024), .Z(n11258) );
  XNOR U11902 ( .A(n11257), .B(n11258), .Z(n11259) );
  XNOR U11903 ( .A(n11260), .B(n11259), .Z(n11265) );
  NANDN U11904 ( .A(n10968), .B(n10967), .Z(n10972) );
  NANDN U11905 ( .A(n10970), .B(n10969), .Z(n10971) );
  AND U11906 ( .A(n10972), .B(n10971), .Z(n11263) );
  NANDN U11907 ( .A(n10974), .B(n10973), .Z(n10978) );
  NAND U11908 ( .A(n10976), .B(n10975), .Z(n10977) );
  NAND U11909 ( .A(n10978), .B(n10977), .Z(n11254) );
  NANDN U11910 ( .A(n10980), .B(n10979), .Z(n10984) );
  NAND U11911 ( .A(n10982), .B(n10981), .Z(n10983) );
  NAND U11912 ( .A(n10984), .B(n10983), .Z(n11251) );
  XNOR U11913 ( .A(n11251), .B(n11252), .Z(n11253) );
  XNOR U11914 ( .A(n11254), .B(n11253), .Z(n11264) );
  XNOR U11915 ( .A(n11271), .B(n11272), .Z(n11275) );
  OR U11916 ( .A(n10990), .B(n10989), .Z(n10994) );
  NANDN U11917 ( .A(n10992), .B(n10991), .Z(n10993) );
  NAND U11918 ( .A(n10994), .B(n10993), .Z(n11276) );
  XNOR U11919 ( .A(n11275), .B(n11276), .Z(n11277) );
  XOR U11920 ( .A(n11278), .B(n11277), .Z(n11001) );
  XNOR U11921 ( .A(n11000), .B(n11001), .Z(n11002) );
  XNOR U11922 ( .A(n11003), .B(n11002), .Z(n11279) );
  XNOR U11923 ( .A(n11279), .B(sreg[130]), .Z(n11281) );
  NAND U11924 ( .A(n10995), .B(sreg[129]), .Z(n10999) );
  OR U11925 ( .A(n10997), .B(n10996), .Z(n10998) );
  AND U11926 ( .A(n10999), .B(n10998), .Z(n11280) );
  XOR U11927 ( .A(n11281), .B(n11280), .Z(c[130]) );
  NANDN U11928 ( .A(n11001), .B(n11000), .Z(n11005) );
  NAND U11929 ( .A(n11003), .B(n11002), .Z(n11004) );
  NAND U11930 ( .A(n11005), .B(n11004), .Z(n11287) );
  NAND U11931 ( .A(n11007), .B(n11006), .Z(n11011) );
  NANDN U11932 ( .A(n11009), .B(n11008), .Z(n11010) );
  NAND U11933 ( .A(n11011), .B(n11010), .Z(n11305) );
  NANDN U11934 ( .A(n11017), .B(n11016), .Z(n11021) );
  NANDN U11935 ( .A(n11019), .B(n11018), .Z(n11020) );
  AND U11936 ( .A(n11021), .B(n11020), .Z(n11303) );
  XNOR U11937 ( .A(n11302), .B(n11303), .Z(n11304) );
  XNOR U11938 ( .A(n11305), .B(n11304), .Z(n11296) );
  NANDN U11939 ( .A(n11023), .B(n11022), .Z(n11027) );
  NAND U11940 ( .A(n11025), .B(n11024), .Z(n11026) );
  NAND U11941 ( .A(n11027), .B(n11026), .Z(n11297) );
  XNOR U11942 ( .A(n11296), .B(n11297), .Z(n11298) );
  XOR U11943 ( .A(b[11]), .B(n26122), .Z(n11486) );
  OR U11944 ( .A(n11486), .B(n31369), .Z(n11030) );
  NANDN U11945 ( .A(n11028), .B(n31119), .Z(n11029) );
  NAND U11946 ( .A(n11030), .B(n11029), .Z(n11507) );
  XOR U11947 ( .A(b[43]), .B(n16916), .Z(n11489) );
  NANDN U11948 ( .A(n11489), .B(n37068), .Z(n11033) );
  NANDN U11949 ( .A(n11031), .B(n37069), .Z(n11032) );
  NAND U11950 ( .A(n11033), .B(n11032), .Z(n11504) );
  XNOR U11951 ( .A(b[45]), .B(a[23]), .Z(n11492) );
  NANDN U11952 ( .A(n11492), .B(n37261), .Z(n11036) );
  NANDN U11953 ( .A(n11034), .B(n37262), .Z(n11035) );
  AND U11954 ( .A(n11036), .B(n11035), .Z(n11505) );
  XNOR U11955 ( .A(n11504), .B(n11505), .Z(n11506) );
  XNOR U11956 ( .A(n11507), .B(n11506), .Z(n11345) );
  XOR U11957 ( .A(b[49]), .B(n15113), .Z(n11495) );
  OR U11958 ( .A(n11495), .B(n37756), .Z(n11039) );
  NANDN U11959 ( .A(n11037), .B(n37652), .Z(n11038) );
  NAND U11960 ( .A(n11039), .B(n11038), .Z(n11532) );
  NAND U11961 ( .A(n11040), .B(n37469), .Z(n11042) );
  XOR U11962 ( .A(n978), .B(n16220), .Z(n11498) );
  NAND U11963 ( .A(n11498), .B(n37471), .Z(n11041) );
  NAND U11964 ( .A(n11042), .B(n11041), .Z(n11529) );
  XNOR U11965 ( .A(b[9]), .B(a[59]), .Z(n11501) );
  NANDN U11966 ( .A(n11501), .B(n30509), .Z(n11045) );
  NAND U11967 ( .A(n11043), .B(n30846), .Z(n11044) );
  AND U11968 ( .A(n11045), .B(n11044), .Z(n11530) );
  XNOR U11969 ( .A(n11529), .B(n11530), .Z(n11531) );
  XNOR U11970 ( .A(n11532), .B(n11531), .Z(n11342) );
  NANDN U11971 ( .A(n11047), .B(n11046), .Z(n11051) );
  NAND U11972 ( .A(n11049), .B(n11048), .Z(n11050) );
  NAND U11973 ( .A(n11051), .B(n11050), .Z(n11343) );
  XNOR U11974 ( .A(n11342), .B(n11343), .Z(n11344) );
  XOR U11975 ( .A(n11345), .B(n11344), .Z(n11541) );
  XNOR U11976 ( .A(n11541), .B(n11542), .Z(n11544) );
  XNOR U11977 ( .A(b[35]), .B(a[33]), .Z(n11514) );
  NANDN U11978 ( .A(n11514), .B(n35985), .Z(n11058) );
  NANDN U11979 ( .A(n11056), .B(n35986), .Z(n11057) );
  NAND U11980 ( .A(n11058), .B(n11057), .Z(n11473) );
  XOR U11981 ( .A(n31123), .B(n27773), .Z(n11517) );
  NAND U11982 ( .A(n11517), .B(n29949), .Z(n11061) );
  NAND U11983 ( .A(n29948), .B(n11059), .Z(n11060) );
  NAND U11984 ( .A(n11061), .B(n11060), .Z(n11470) );
  XOR U11985 ( .A(b[55]), .B(n13509), .Z(n11520) );
  NANDN U11986 ( .A(n11520), .B(n38075), .Z(n11064) );
  NANDN U11987 ( .A(n11062), .B(n38073), .Z(n11063) );
  AND U11988 ( .A(n11064), .B(n11063), .Z(n11471) );
  XNOR U11989 ( .A(n11470), .B(n11471), .Z(n11472) );
  XNOR U11990 ( .A(n11473), .B(n11472), .Z(n11333) );
  NANDN U11991 ( .A(n11066), .B(n11065), .Z(n11070) );
  NAND U11992 ( .A(n11068), .B(n11067), .Z(n11069) );
  NAND U11993 ( .A(n11070), .B(n11069), .Z(n11330) );
  XNOR U11994 ( .A(n11330), .B(n11331), .Z(n11332) );
  XOR U11995 ( .A(n11333), .B(n11332), .Z(n11543) );
  XNOR U11996 ( .A(n11544), .B(n11543), .Z(n11535) );
  NANDN U11997 ( .A(n11076), .B(n11075), .Z(n11080) );
  NANDN U11998 ( .A(n11078), .B(n11077), .Z(n11079) );
  NAND U11999 ( .A(n11080), .B(n11079), .Z(n11554) );
  XOR U12000 ( .A(b[15]), .B(n25001), .Z(n11446) );
  OR U12001 ( .A(n11446), .B(n32010), .Z(n11083) );
  NANDN U12002 ( .A(n11081), .B(n32011), .Z(n11082) );
  NAND U12003 ( .A(n11083), .B(n11082), .Z(n11358) );
  XNOR U12004 ( .A(b[25]), .B(n21996), .Z(n11449) );
  NANDN U12005 ( .A(n34219), .B(n11449), .Z(n11086) );
  NAND U12006 ( .A(n34217), .B(n11084), .Z(n11085) );
  NAND U12007 ( .A(n11086), .B(n11085), .Z(n11355) );
  XNOR U12008 ( .A(b[17]), .B(a[51]), .Z(n11452) );
  NANDN U12009 ( .A(n11452), .B(n32543), .Z(n11089) );
  NANDN U12010 ( .A(n11087), .B(n32541), .Z(n11088) );
  AND U12011 ( .A(n11089), .B(n11088), .Z(n11356) );
  XNOR U12012 ( .A(n11355), .B(n11356), .Z(n11357) );
  XNOR U12013 ( .A(n11358), .B(n11357), .Z(n11428) );
  XOR U12014 ( .A(b[39]), .B(n18003), .Z(n11455) );
  NANDN U12015 ( .A(n11455), .B(n36553), .Z(n11092) );
  NANDN U12016 ( .A(n11090), .B(n36643), .Z(n11091) );
  NAND U12017 ( .A(n11092), .B(n11091), .Z(n11388) );
  XOR U12018 ( .A(b[51]), .B(n14514), .Z(n11458) );
  NANDN U12019 ( .A(n11458), .B(n37803), .Z(n11095) );
  NANDN U12020 ( .A(n11093), .B(n37802), .Z(n11094) );
  NAND U12021 ( .A(n11095), .B(n11094), .Z(n11385) );
  XOR U12022 ( .A(b[53]), .B(n13976), .Z(n11461) );
  NANDN U12023 ( .A(n11461), .B(n37940), .Z(n11098) );
  NANDN U12024 ( .A(n11096), .B(n37941), .Z(n11097) );
  AND U12025 ( .A(n11098), .B(n11097), .Z(n11386) );
  XNOR U12026 ( .A(n11385), .B(n11386), .Z(n11387) );
  XOR U12027 ( .A(n11388), .B(n11387), .Z(n11429) );
  XOR U12028 ( .A(n11428), .B(n11429), .Z(n11431) );
  NANDN U12029 ( .A(n11100), .B(n11099), .Z(n11104) );
  NAND U12030 ( .A(n11102), .B(n11101), .Z(n11103) );
  NAND U12031 ( .A(n11104), .B(n11103), .Z(n11430) );
  XNOR U12032 ( .A(n11431), .B(n11430), .Z(n11483) );
  NANDN U12033 ( .A(n11106), .B(n11105), .Z(n11110) );
  NAND U12034 ( .A(n11108), .B(n11107), .Z(n11109) );
  NAND U12035 ( .A(n11110), .B(n11109), .Z(n11480) );
  XNOR U12036 ( .A(n11480), .B(n11481), .Z(n11482) );
  XNOR U12037 ( .A(n11483), .B(n11482), .Z(n11551) );
  NANDN U12038 ( .A(n11116), .B(n11115), .Z(n11120) );
  OR U12039 ( .A(n11118), .B(n11117), .Z(n11119) );
  AND U12040 ( .A(n11120), .B(n11119), .Z(n11552) );
  XNOR U12041 ( .A(n11551), .B(n11552), .Z(n11553) );
  XOR U12042 ( .A(n11554), .B(n11553), .Z(n11536) );
  NAND U12043 ( .A(n11122), .B(n11121), .Z(n11126) );
  NANDN U12044 ( .A(n11124), .B(n11123), .Z(n11125) );
  AND U12045 ( .A(n11126), .B(n11125), .Z(n11538) );
  XNOR U12046 ( .A(n11537), .B(n11538), .Z(n11308) );
  NANDN U12047 ( .A(n11128), .B(n11127), .Z(n11132) );
  NAND U12048 ( .A(n11130), .B(n11129), .Z(n11131) );
  NAND U12049 ( .A(n11132), .B(n11131), .Z(n11549) );
  NANDN U12050 ( .A(n11134), .B(n11133), .Z(n11138) );
  NANDN U12051 ( .A(n11136), .B(n11135), .Z(n11137) );
  NAND U12052 ( .A(n11138), .B(n11137), .Z(n11547) );
  NANDN U12053 ( .A(n11140), .B(n11139), .Z(n11144) );
  OR U12054 ( .A(n11142), .B(n11141), .Z(n11143) );
  NAND U12055 ( .A(n11144), .B(n11143), .Z(n11548) );
  XNOR U12056 ( .A(n11547), .B(n11548), .Z(n11550) );
  XOR U12057 ( .A(n11549), .B(n11550), .Z(n11317) );
  NANDN U12058 ( .A(n11146), .B(n11145), .Z(n11150) );
  NAND U12059 ( .A(n11148), .B(n11147), .Z(n11149) );
  NAND U12060 ( .A(n11150), .B(n11149), .Z(n11321) );
  XOR U12061 ( .A(b[37]), .B(n18639), .Z(n11367) );
  NANDN U12062 ( .A(n11367), .B(n36311), .Z(n11153) );
  NANDN U12063 ( .A(n11151), .B(n36309), .Z(n11152) );
  NAND U12064 ( .A(n11153), .B(n11152), .Z(n11425) );
  XNOR U12065 ( .A(b[5]), .B(a[63]), .Z(n11370) );
  OR U12066 ( .A(n11370), .B(n29363), .Z(n11156) );
  NANDN U12067 ( .A(n11154), .B(n29864), .Z(n11155) );
  NAND U12068 ( .A(n11156), .B(n11155), .Z(n11422) );
  XOR U12069 ( .A(n967), .B(n28403), .Z(n11373) );
  NAND U12070 ( .A(n11373), .B(n28939), .Z(n11159) );
  NAND U12071 ( .A(n28938), .B(n11157), .Z(n11158) );
  AND U12072 ( .A(n11159), .B(n11158), .Z(n11423) );
  XNOR U12073 ( .A(n11422), .B(n11423), .Z(n11424) );
  XOR U12074 ( .A(n11425), .B(n11424), .Z(n11324) );
  XOR U12075 ( .A(b[13]), .B(n25466), .Z(n11376) );
  OR U12076 ( .A(n11376), .B(n31550), .Z(n11162) );
  NANDN U12077 ( .A(n11160), .B(n31874), .Z(n11161) );
  NAND U12078 ( .A(n11162), .B(n11161), .Z(n11467) );
  NAND U12079 ( .A(n34848), .B(n11163), .Z(n11165) );
  XOR U12080 ( .A(n35375), .B(n21441), .Z(n11379) );
  NAND U12081 ( .A(n34618), .B(n11379), .Z(n11164) );
  NAND U12082 ( .A(n11165), .B(n11164), .Z(n11464) );
  NAND U12083 ( .A(n35188), .B(n11166), .Z(n11168) );
  XOR U12084 ( .A(n35540), .B(n20867), .Z(n11382) );
  NANDN U12085 ( .A(n34968), .B(n11382), .Z(n11167) );
  AND U12086 ( .A(n11168), .B(n11167), .Z(n11465) );
  XNOR U12087 ( .A(n11464), .B(n11465), .Z(n11466) );
  XOR U12088 ( .A(n11467), .B(n11466), .Z(n11325) );
  XNOR U12089 ( .A(n11324), .B(n11325), .Z(n11327) );
  NANDN U12090 ( .A(n11170), .B(n11169), .Z(n11174) );
  NAND U12091 ( .A(n11172), .B(n11171), .Z(n11173) );
  NAND U12092 ( .A(n11174), .B(n11173), .Z(n11326) );
  XNOR U12093 ( .A(n11327), .B(n11326), .Z(n11319) );
  NANDN U12094 ( .A(n11176), .B(n11175), .Z(n11180) );
  NAND U12095 ( .A(n11178), .B(n11177), .Z(n11179) );
  NAND U12096 ( .A(n11180), .B(n11179), .Z(n11512) );
  NAND U12097 ( .A(a[3]), .B(b[63]), .Z(n11526) );
  NANDN U12098 ( .A(n11181), .B(n38369), .Z(n11183) );
  XOR U12099 ( .A(b[61]), .B(n11694), .Z(n11361) );
  OR U12100 ( .A(n11361), .B(n38371), .Z(n11182) );
  NAND U12101 ( .A(n11183), .B(n11182), .Z(n11524) );
  NANDN U12102 ( .A(n11184), .B(n35311), .Z(n11186) );
  XOR U12103 ( .A(b[31]), .B(n20352), .Z(n11364) );
  NANDN U12104 ( .A(n11364), .B(n35313), .Z(n11185) );
  AND U12105 ( .A(n11186), .B(n11185), .Z(n11523) );
  XNOR U12106 ( .A(n11524), .B(n11523), .Z(n11525) );
  XOR U12107 ( .A(n11526), .B(n11525), .Z(n11510) );
  NAND U12108 ( .A(n33283), .B(n11187), .Z(n11189) );
  XOR U12109 ( .A(n33020), .B(n23852), .Z(n11346) );
  NANDN U12110 ( .A(n33021), .B(n11346), .Z(n11188) );
  NAND U12111 ( .A(n11189), .B(n11188), .Z(n11413) );
  XNOR U12112 ( .A(b[21]), .B(a[47]), .Z(n11349) );
  OR U12113 ( .A(n11349), .B(n33634), .Z(n11192) );
  NANDN U12114 ( .A(n11190), .B(n33464), .Z(n11191) );
  NAND U12115 ( .A(n11192), .B(n11191), .Z(n11410) );
  NAND U12116 ( .A(n34044), .B(n11193), .Z(n11195) );
  XOR U12117 ( .A(n34510), .B(n22579), .Z(n11352) );
  NANDN U12118 ( .A(n33867), .B(n11352), .Z(n11194) );
  AND U12119 ( .A(n11195), .B(n11194), .Z(n11411) );
  XNOR U12120 ( .A(n11410), .B(n11411), .Z(n11412) );
  XNOR U12121 ( .A(n11413), .B(n11412), .Z(n11511) );
  XNOR U12122 ( .A(n11510), .B(n11511), .Z(n11513) );
  XNOR U12123 ( .A(n11512), .B(n11513), .Z(n11318) );
  XOR U12124 ( .A(n11319), .B(n11318), .Z(n11320) );
  XOR U12125 ( .A(n11321), .B(n11320), .Z(n11437) );
  XOR U12126 ( .A(b[33]), .B(n20315), .Z(n11400) );
  NANDN U12127 ( .A(n11400), .B(n35620), .Z(n11198) );
  NANDN U12128 ( .A(n11196), .B(n35621), .Z(n11197) );
  NAND U12129 ( .A(n11198), .B(n11197), .Z(n11479) );
  NANDN U12130 ( .A(n966), .B(a[67]), .Z(n11199) );
  XOR U12131 ( .A(n29232), .B(n11199), .Z(n11201) );
  IV U12132 ( .A(a[66]), .Z(n28701) );
  NANDN U12133 ( .A(n28701), .B(n966), .Z(n11200) );
  AND U12134 ( .A(n11201), .B(n11200), .Z(n11476) );
  XOR U12135 ( .A(b[63]), .B(n11202), .Z(n11407) );
  NANDN U12136 ( .A(n11407), .B(n38422), .Z(n11205) );
  NANDN U12137 ( .A(n11203), .B(n38423), .Z(n11204) );
  AND U12138 ( .A(n11205), .B(n11204), .Z(n11477) );
  XNOR U12139 ( .A(n11476), .B(n11477), .Z(n11478) );
  XNOR U12140 ( .A(n11479), .B(n11478), .Z(n11442) );
  XNOR U12141 ( .A(b[41]), .B(a[27]), .Z(n11391) );
  OR U12142 ( .A(n11391), .B(n36905), .Z(n11208) );
  NANDN U12143 ( .A(n11206), .B(n36807), .Z(n11207) );
  NAND U12144 ( .A(n11208), .B(n11207), .Z(n11419) );
  XOR U12145 ( .A(b[57]), .B(n12830), .Z(n11394) );
  OR U12146 ( .A(n11394), .B(n965), .Z(n11211) );
  NANDN U12147 ( .A(n11209), .B(n38194), .Z(n11210) );
  NAND U12148 ( .A(n11211), .B(n11210), .Z(n11416) );
  NAND U12149 ( .A(n38326), .B(n11212), .Z(n11214) );
  XOR U12150 ( .A(n38400), .B(n12258), .Z(n11397) );
  NANDN U12151 ( .A(n38273), .B(n11397), .Z(n11213) );
  AND U12152 ( .A(n11214), .B(n11213), .Z(n11417) );
  XNOR U12153 ( .A(n11416), .B(n11417), .Z(n11418) );
  XOR U12154 ( .A(n11419), .B(n11418), .Z(n11441) );
  NANDN U12155 ( .A(n11216), .B(n11215), .Z(n11220) );
  NAND U12156 ( .A(n11218), .B(n11217), .Z(n11219) );
  NAND U12157 ( .A(n11220), .B(n11219), .Z(n11440) );
  XNOR U12158 ( .A(n11441), .B(n11440), .Z(n11443) );
  XNOR U12159 ( .A(n11442), .B(n11443), .Z(n11339) );
  NANDN U12160 ( .A(n11222), .B(n11221), .Z(n11226) );
  NAND U12161 ( .A(n11224), .B(n11223), .Z(n11225) );
  NAND U12162 ( .A(n11226), .B(n11225), .Z(n11336) );
  NANDN U12163 ( .A(n11228), .B(n11227), .Z(n11232) );
  NAND U12164 ( .A(n11230), .B(n11229), .Z(n11231) );
  AND U12165 ( .A(n11232), .B(n11231), .Z(n11337) );
  XNOR U12166 ( .A(n11336), .B(n11337), .Z(n11338) );
  XNOR U12167 ( .A(n11339), .B(n11338), .Z(n11435) );
  NANDN U12168 ( .A(n11234), .B(n11233), .Z(n11238) );
  NANDN U12169 ( .A(n11236), .B(n11235), .Z(n11237) );
  AND U12170 ( .A(n11238), .B(n11237), .Z(n11434) );
  XOR U12171 ( .A(n11435), .B(n11434), .Z(n11436) );
  XNOR U12172 ( .A(n11437), .B(n11436), .Z(n11314) );
  NANDN U12173 ( .A(n11240), .B(n11239), .Z(n11244) );
  OR U12174 ( .A(n11242), .B(n11241), .Z(n11243) );
  AND U12175 ( .A(n11244), .B(n11243), .Z(n11315) );
  XNOR U12176 ( .A(n11314), .B(n11315), .Z(n11316) );
  XNOR U12177 ( .A(n11317), .B(n11316), .Z(n11309) );
  XOR U12178 ( .A(n11308), .B(n11309), .Z(n11310) );
  NAND U12179 ( .A(n11246), .B(n11245), .Z(n11250) );
  NANDN U12180 ( .A(n11248), .B(n11247), .Z(n11249) );
  AND U12181 ( .A(n11250), .B(n11249), .Z(n11311) );
  XNOR U12182 ( .A(n11310), .B(n11311), .Z(n11299) );
  XOR U12183 ( .A(n11298), .B(n11299), .Z(n11293) );
  NANDN U12184 ( .A(n11252), .B(n11251), .Z(n11256) );
  NAND U12185 ( .A(n11254), .B(n11253), .Z(n11255) );
  NAND U12186 ( .A(n11256), .B(n11255), .Z(n11290) );
  NANDN U12187 ( .A(n11258), .B(n11257), .Z(n11262) );
  NAND U12188 ( .A(n11260), .B(n11259), .Z(n11261) );
  NAND U12189 ( .A(n11262), .B(n11261), .Z(n11291) );
  XNOR U12190 ( .A(n11290), .B(n11291), .Z(n11292) );
  XNOR U12191 ( .A(n11293), .B(n11292), .Z(n11560) );
  OR U12192 ( .A(n11264), .B(n11263), .Z(n11268) );
  NANDN U12193 ( .A(n11266), .B(n11265), .Z(n11267) );
  NAND U12194 ( .A(n11268), .B(n11267), .Z(n11558) );
  NANDN U12195 ( .A(n11270), .B(n11269), .Z(n11274) );
  NAND U12196 ( .A(n11272), .B(n11271), .Z(n11273) );
  AND U12197 ( .A(n11274), .B(n11273), .Z(n11557) );
  XNOR U12198 ( .A(n11558), .B(n11557), .Z(n11559) );
  XOR U12199 ( .A(n11560), .B(n11559), .Z(n11284) );
  XOR U12200 ( .A(n11284), .B(n11285), .Z(n11286) );
  XNOR U12201 ( .A(n11287), .B(n11286), .Z(n11563) );
  XNOR U12202 ( .A(n11563), .B(sreg[131]), .Z(n11565) );
  NAND U12203 ( .A(n11279), .B(sreg[130]), .Z(n11283) );
  OR U12204 ( .A(n11281), .B(n11280), .Z(n11282) );
  AND U12205 ( .A(n11283), .B(n11282), .Z(n11564) );
  XOR U12206 ( .A(n11565), .B(n11564), .Z(c[131]) );
  OR U12207 ( .A(n11285), .B(n11284), .Z(n11289) );
  NAND U12208 ( .A(n11287), .B(n11286), .Z(n11288) );
  NAND U12209 ( .A(n11289), .B(n11288), .Z(n11571) );
  NANDN U12210 ( .A(n11291), .B(n11290), .Z(n11295) );
  NAND U12211 ( .A(n11293), .B(n11292), .Z(n11294) );
  NAND U12212 ( .A(n11295), .B(n11294), .Z(n11849) );
  NANDN U12213 ( .A(n11297), .B(n11296), .Z(n11301) );
  NANDN U12214 ( .A(n11299), .B(n11298), .Z(n11300) );
  NAND U12215 ( .A(n11301), .B(n11300), .Z(n11850) );
  XNOR U12216 ( .A(n11849), .B(n11850), .Z(n11851) );
  NANDN U12217 ( .A(n11303), .B(n11302), .Z(n11307) );
  NAND U12218 ( .A(n11305), .B(n11304), .Z(n11306) );
  NAND U12219 ( .A(n11307), .B(n11306), .Z(n11843) );
  OR U12220 ( .A(n11309), .B(n11308), .Z(n11313) );
  NAND U12221 ( .A(n11311), .B(n11310), .Z(n11312) );
  NAND U12222 ( .A(n11313), .B(n11312), .Z(n11844) );
  XNOR U12223 ( .A(n11843), .B(n11844), .Z(n11845) );
  NAND U12224 ( .A(n11319), .B(n11318), .Z(n11323) );
  NANDN U12225 ( .A(n11321), .B(n11320), .Z(n11322) );
  NAND U12226 ( .A(n11323), .B(n11322), .Z(n11809) );
  OR U12227 ( .A(n11325), .B(n11324), .Z(n11329) );
  OR U12228 ( .A(n11327), .B(n11326), .Z(n11328) );
  NAND U12229 ( .A(n11329), .B(n11328), .Z(n11829) );
  NANDN U12230 ( .A(n11331), .B(n11330), .Z(n11335) );
  NAND U12231 ( .A(n11333), .B(n11332), .Z(n11334) );
  NAND U12232 ( .A(n11335), .B(n11334), .Z(n11827) );
  NANDN U12233 ( .A(n11337), .B(n11336), .Z(n11341) );
  NANDN U12234 ( .A(n11339), .B(n11338), .Z(n11340) );
  NAND U12235 ( .A(n11341), .B(n11340), .Z(n11828) );
  XNOR U12236 ( .A(n11827), .B(n11828), .Z(n11830) );
  XNOR U12237 ( .A(n11829), .B(n11830), .Z(n11810) );
  XOR U12238 ( .A(n11809), .B(n11810), .Z(n11811) );
  NAND U12239 ( .A(n33283), .B(n11346), .Z(n11348) );
  XOR U12240 ( .A(n33020), .B(n24671), .Z(n11616) );
  NANDN U12241 ( .A(n33021), .B(n11616), .Z(n11347) );
  NAND U12242 ( .A(n11348), .B(n11347), .Z(n11676) );
  XNOR U12243 ( .A(b[21]), .B(a[48]), .Z(n11619) );
  OR U12244 ( .A(n11619), .B(n33634), .Z(n11351) );
  NANDN U12245 ( .A(n11349), .B(n33464), .Z(n11350) );
  NAND U12246 ( .A(n11351), .B(n11350), .Z(n11673) );
  NAND U12247 ( .A(n34044), .B(n11352), .Z(n11354) );
  XOR U12248 ( .A(n34510), .B(n22964), .Z(n11622) );
  NANDN U12249 ( .A(n33867), .B(n11622), .Z(n11353) );
  AND U12250 ( .A(n11354), .B(n11353), .Z(n11674) );
  XNOR U12251 ( .A(n11673), .B(n11674), .Z(n11675) );
  XOR U12252 ( .A(n11676), .B(n11675), .Z(n11731) );
  NANDN U12253 ( .A(n11356), .B(n11355), .Z(n11360) );
  NAND U12254 ( .A(n11358), .B(n11357), .Z(n11359) );
  NAND U12255 ( .A(n11360), .B(n11359), .Z(n11732) );
  XNOR U12256 ( .A(n11731), .B(n11732), .Z(n11734) );
  NAND U12257 ( .A(a[4]), .B(b[63]), .Z(n11722) );
  NANDN U12258 ( .A(n11361), .B(n38369), .Z(n11363) );
  XOR U12259 ( .A(b[61]), .B(n11986), .Z(n11631) );
  OR U12260 ( .A(n11631), .B(n38371), .Z(n11362) );
  NAND U12261 ( .A(n11363), .B(n11362), .Z(n11720) );
  NANDN U12262 ( .A(n11364), .B(n35311), .Z(n11366) );
  XOR U12263 ( .A(b[31]), .B(n20686), .Z(n11634) );
  NANDN U12264 ( .A(n11634), .B(n35313), .Z(n11365) );
  AND U12265 ( .A(n11366), .B(n11365), .Z(n11719) );
  XNOR U12266 ( .A(n11720), .B(n11719), .Z(n11721) );
  XNOR U12267 ( .A(n11722), .B(n11721), .Z(n11733) );
  XNOR U12268 ( .A(n11734), .B(n11733), .Z(n11604) );
  XOR U12269 ( .A(b[37]), .B(n18841), .Z(n11646) );
  NANDN U12270 ( .A(n11646), .B(n36311), .Z(n11369) );
  NANDN U12271 ( .A(n11367), .B(n36309), .Z(n11368) );
  NAND U12272 ( .A(n11369), .B(n11368), .Z(n11670) );
  XNOR U12273 ( .A(b[5]), .B(a[64]), .Z(n11649) );
  OR U12274 ( .A(n11649), .B(n29363), .Z(n11372) );
  NANDN U12275 ( .A(n11370), .B(n29864), .Z(n11371) );
  NAND U12276 ( .A(n11372), .B(n11371), .Z(n11667) );
  XOR U12277 ( .A(n967), .B(n28701), .Z(n11652) );
  NAND U12278 ( .A(n11652), .B(n28939), .Z(n11375) );
  NAND U12279 ( .A(n28938), .B(n11373), .Z(n11374) );
  AND U12280 ( .A(n11375), .B(n11374), .Z(n11668) );
  XNOR U12281 ( .A(n11667), .B(n11668), .Z(n11669) );
  XNOR U12282 ( .A(n11670), .B(n11669), .Z(n11586) );
  XOR U12283 ( .A(b[13]), .B(n25860), .Z(n11637) );
  OR U12284 ( .A(n11637), .B(n31550), .Z(n11378) );
  NANDN U12285 ( .A(n11376), .B(n31874), .Z(n11377) );
  NAND U12286 ( .A(n11378), .B(n11377), .Z(n11782) );
  NAND U12287 ( .A(n34848), .B(n11379), .Z(n11381) );
  XOR U12288 ( .A(n35375), .B(n22246), .Z(n11640) );
  NAND U12289 ( .A(n34618), .B(n11640), .Z(n11380) );
  NAND U12290 ( .A(n11381), .B(n11380), .Z(n11779) );
  NAND U12291 ( .A(n35188), .B(n11382), .Z(n11384) );
  XOR U12292 ( .A(n35540), .B(n21149), .Z(n11643) );
  NANDN U12293 ( .A(n34968), .B(n11643), .Z(n11383) );
  AND U12294 ( .A(n11384), .B(n11383), .Z(n11780) );
  XNOR U12295 ( .A(n11779), .B(n11780), .Z(n11781) );
  XOR U12296 ( .A(n11782), .B(n11781), .Z(n11587) );
  XOR U12297 ( .A(n11586), .B(n11587), .Z(n11589) );
  NANDN U12298 ( .A(n11386), .B(n11385), .Z(n11390) );
  NAND U12299 ( .A(n11388), .B(n11387), .Z(n11389) );
  NAND U12300 ( .A(n11390), .B(n11389), .Z(n11588) );
  XOR U12301 ( .A(n11589), .B(n11588), .Z(n11605) );
  XOR U12302 ( .A(n11604), .B(n11605), .Z(n11607) );
  XNOR U12303 ( .A(n11606), .B(n11607), .Z(n11707) );
  XNOR U12304 ( .A(b[41]), .B(a[28]), .Z(n11679) );
  OR U12305 ( .A(n11679), .B(n36905), .Z(n11393) );
  NANDN U12306 ( .A(n11391), .B(n36807), .Z(n11392) );
  NAND U12307 ( .A(n11393), .B(n11392), .Z(n11701) );
  XOR U12308 ( .A(b[57]), .B(n13106), .Z(n11682) );
  OR U12309 ( .A(n11682), .B(n965), .Z(n11396) );
  NANDN U12310 ( .A(n11394), .B(n38194), .Z(n11395) );
  NAND U12311 ( .A(n11396), .B(n11395), .Z(n11698) );
  NAND U12312 ( .A(n38326), .B(n11397), .Z(n11399) );
  XOR U12313 ( .A(n38400), .B(n12555), .Z(n11685) );
  NANDN U12314 ( .A(n38273), .B(n11685), .Z(n11398) );
  AND U12315 ( .A(n11399), .B(n11398), .Z(n11699) );
  XNOR U12316 ( .A(n11698), .B(n11699), .Z(n11700) );
  XOR U12317 ( .A(n11701), .B(n11700), .Z(n11797) );
  XOR U12318 ( .A(b[33]), .B(n19980), .Z(n11688) );
  NANDN U12319 ( .A(n11688), .B(n35620), .Z(n11402) );
  NANDN U12320 ( .A(n11400), .B(n35621), .Z(n11401) );
  NAND U12321 ( .A(n11402), .B(n11401), .Z(n11794) );
  NANDN U12322 ( .A(n966), .B(a[68]), .Z(n11403) );
  XOR U12323 ( .A(n29232), .B(n11403), .Z(n11405) );
  IV U12324 ( .A(a[67]), .Z(n29372) );
  NANDN U12325 ( .A(n29372), .B(n966), .Z(n11404) );
  AND U12326 ( .A(n11405), .B(n11404), .Z(n11791) );
  XOR U12327 ( .A(b[63]), .B(n11406), .Z(n11695) );
  NANDN U12328 ( .A(n11695), .B(n38422), .Z(n11409) );
  NANDN U12329 ( .A(n11407), .B(n38423), .Z(n11408) );
  AND U12330 ( .A(n11409), .B(n11408), .Z(n11792) );
  XNOR U12331 ( .A(n11791), .B(n11792), .Z(n11793) );
  XOR U12332 ( .A(n11794), .B(n11793), .Z(n11798) );
  XNOR U12333 ( .A(n11797), .B(n11798), .Z(n11800) );
  NANDN U12334 ( .A(n11411), .B(n11410), .Z(n11415) );
  NAND U12335 ( .A(n11413), .B(n11412), .Z(n11414) );
  NAND U12336 ( .A(n11415), .B(n11414), .Z(n11799) );
  XNOR U12337 ( .A(n11800), .B(n11799), .Z(n11601) );
  NANDN U12338 ( .A(n11417), .B(n11416), .Z(n11421) );
  NAND U12339 ( .A(n11419), .B(n11418), .Z(n11420) );
  NAND U12340 ( .A(n11421), .B(n11420), .Z(n11598) );
  NANDN U12341 ( .A(n11423), .B(n11422), .Z(n11427) );
  NAND U12342 ( .A(n11425), .B(n11424), .Z(n11426) );
  AND U12343 ( .A(n11427), .B(n11426), .Z(n11599) );
  XNOR U12344 ( .A(n11598), .B(n11599), .Z(n11600) );
  XOR U12345 ( .A(n11601), .B(n11600), .Z(n11705) );
  NANDN U12346 ( .A(n11429), .B(n11428), .Z(n11433) );
  OR U12347 ( .A(n11431), .B(n11430), .Z(n11432) );
  AND U12348 ( .A(n11433), .B(n11432), .Z(n11704) );
  XOR U12349 ( .A(n11705), .B(n11704), .Z(n11706) );
  XNOR U12350 ( .A(n11707), .B(n11706), .Z(n11812) );
  XOR U12351 ( .A(n11811), .B(n11812), .Z(n11580) );
  OR U12352 ( .A(n11435), .B(n11434), .Z(n11439) );
  NAND U12353 ( .A(n11437), .B(n11436), .Z(n11438) );
  NAND U12354 ( .A(n11439), .B(n11438), .Z(n11833) );
  OR U12355 ( .A(n11441), .B(n11440), .Z(n11445) );
  NANDN U12356 ( .A(n11443), .B(n11442), .Z(n11444) );
  NAND U12357 ( .A(n11445), .B(n11444), .Z(n11821) );
  XOR U12358 ( .A(b[15]), .B(n25177), .Z(n11761) );
  OR U12359 ( .A(n11761), .B(n32010), .Z(n11448) );
  NANDN U12360 ( .A(n11446), .B(n32011), .Z(n11447) );
  NAND U12361 ( .A(n11448), .B(n11447), .Z(n11628) );
  XNOR U12362 ( .A(b[25]), .B(n22289), .Z(n11764) );
  NANDN U12363 ( .A(n34219), .B(n11764), .Z(n11451) );
  NAND U12364 ( .A(n34217), .B(n11449), .Z(n11450) );
  NAND U12365 ( .A(n11451), .B(n11450), .Z(n11625) );
  XNOR U12366 ( .A(b[17]), .B(a[52]), .Z(n11767) );
  NANDN U12367 ( .A(n11767), .B(n32543), .Z(n11454) );
  NANDN U12368 ( .A(n11452), .B(n32541), .Z(n11453) );
  AND U12369 ( .A(n11454), .B(n11453), .Z(n11626) );
  XNOR U12370 ( .A(n11625), .B(n11626), .Z(n11627) );
  XNOR U12371 ( .A(n11628), .B(n11627), .Z(n11661) );
  XOR U12372 ( .A(b[39]), .B(n18804), .Z(n11770) );
  NANDN U12373 ( .A(n11770), .B(n36553), .Z(n11457) );
  NANDN U12374 ( .A(n11455), .B(n36643), .Z(n11456) );
  NAND U12375 ( .A(n11457), .B(n11456), .Z(n11658) );
  XOR U12376 ( .A(b[51]), .B(n14905), .Z(n11773) );
  NANDN U12377 ( .A(n11773), .B(n37803), .Z(n11460) );
  NANDN U12378 ( .A(n11458), .B(n37802), .Z(n11459) );
  NAND U12379 ( .A(n11460), .B(n11459), .Z(n11655) );
  XOR U12380 ( .A(b[53]), .B(n14259), .Z(n11776) );
  NANDN U12381 ( .A(n11776), .B(n37940), .Z(n11463) );
  NANDN U12382 ( .A(n11461), .B(n37941), .Z(n11462) );
  AND U12383 ( .A(n11463), .B(n11462), .Z(n11656) );
  XNOR U12384 ( .A(n11655), .B(n11656), .Z(n11657) );
  XOR U12385 ( .A(n11658), .B(n11657), .Z(n11662) );
  XOR U12386 ( .A(n11661), .B(n11662), .Z(n11664) );
  NANDN U12387 ( .A(n11465), .B(n11464), .Z(n11469) );
  NAND U12388 ( .A(n11467), .B(n11466), .Z(n11468) );
  NAND U12389 ( .A(n11469), .B(n11468), .Z(n11663) );
  XNOR U12390 ( .A(n11664), .B(n11663), .Z(n11806) );
  NANDN U12391 ( .A(n11471), .B(n11470), .Z(n11475) );
  NAND U12392 ( .A(n11473), .B(n11472), .Z(n11474) );
  NAND U12393 ( .A(n11475), .B(n11474), .Z(n11803) );
  XNOR U12394 ( .A(n11803), .B(n11804), .Z(n11805) );
  XOR U12395 ( .A(n11806), .B(n11805), .Z(n11822) );
  XNOR U12396 ( .A(n11821), .B(n11822), .Z(n11823) );
  NANDN U12397 ( .A(n11481), .B(n11480), .Z(n11485) );
  NAND U12398 ( .A(n11483), .B(n11482), .Z(n11484) );
  AND U12399 ( .A(n11485), .B(n11484), .Z(n11824) );
  XNOR U12400 ( .A(n11823), .B(n11824), .Z(n11832) );
  XOR U12401 ( .A(b[11]), .B(n26347), .Z(n11746) );
  OR U12402 ( .A(n11746), .B(n31369), .Z(n11488) );
  NANDN U12403 ( .A(n11486), .B(n31119), .Z(n11487) );
  NAND U12404 ( .A(n11488), .B(n11487), .Z(n11758) );
  XOR U12405 ( .A(b[43]), .B(n17133), .Z(n11749) );
  NANDN U12406 ( .A(n11749), .B(n37068), .Z(n11491) );
  NANDN U12407 ( .A(n11489), .B(n37069), .Z(n11490) );
  NAND U12408 ( .A(n11491), .B(n11490), .Z(n11755) );
  XNOR U12409 ( .A(b[45]), .B(a[24]), .Z(n11752) );
  NANDN U12410 ( .A(n11752), .B(n37261), .Z(n11494) );
  NANDN U12411 ( .A(n11492), .B(n37262), .Z(n11493) );
  AND U12412 ( .A(n11494), .B(n11493), .Z(n11756) );
  XNOR U12413 ( .A(n11755), .B(n11756), .Z(n11757) );
  XNOR U12414 ( .A(n11758), .B(n11757), .Z(n11610) );
  XOR U12415 ( .A(n979), .B(n15484), .Z(n11737) );
  NANDN U12416 ( .A(n37756), .B(n11737), .Z(n11497) );
  NANDN U12417 ( .A(n11495), .B(n37652), .Z(n11496) );
  NAND U12418 ( .A(n11497), .B(n11496), .Z(n11728) );
  NAND U12419 ( .A(n37469), .B(n11498), .Z(n11500) );
  XOR U12420 ( .A(b[47]), .B(n15963), .Z(n11740) );
  NANDN U12421 ( .A(n11740), .B(n37471), .Z(n11499) );
  NAND U12422 ( .A(n11500), .B(n11499), .Z(n11725) );
  XOR U12423 ( .A(n969), .B(n27436), .Z(n11743) );
  NAND U12424 ( .A(n30509), .B(n11743), .Z(n11503) );
  NANDN U12425 ( .A(n11501), .B(n30846), .Z(n11502) );
  AND U12426 ( .A(n11503), .B(n11502), .Z(n11726) );
  XNOR U12427 ( .A(n11725), .B(n11726), .Z(n11727) );
  XOR U12428 ( .A(n11728), .B(n11727), .Z(n11611) );
  XNOR U12429 ( .A(n11610), .B(n11611), .Z(n11612) );
  NANDN U12430 ( .A(n11505), .B(n11504), .Z(n11509) );
  NAND U12431 ( .A(n11507), .B(n11506), .Z(n11508) );
  AND U12432 ( .A(n11509), .B(n11508), .Z(n11613) );
  XNOR U12433 ( .A(n11612), .B(n11613), .Z(n11816) );
  XNOR U12434 ( .A(n11816), .B(n11815), .Z(n11817) );
  XNOR U12435 ( .A(b[35]), .B(a[34]), .Z(n11710) );
  NANDN U12436 ( .A(n11710), .B(n35985), .Z(n11516) );
  NANDN U12437 ( .A(n11514), .B(n35986), .Z(n11515) );
  NAND U12438 ( .A(n11516), .B(n11515), .Z(n11788) );
  XNOR U12439 ( .A(n31123), .B(a[62]), .Z(n11713) );
  NAND U12440 ( .A(n11713), .B(n29949), .Z(n11519) );
  NAND U12441 ( .A(n29948), .B(n11517), .Z(n11518) );
  NAND U12442 ( .A(n11519), .B(n11518), .Z(n11785) );
  XOR U12443 ( .A(b[55]), .B(n14210), .Z(n11716) );
  NANDN U12444 ( .A(n11716), .B(n38075), .Z(n11522) );
  NANDN U12445 ( .A(n11520), .B(n38073), .Z(n11521) );
  AND U12446 ( .A(n11522), .B(n11521), .Z(n11786) );
  XNOR U12447 ( .A(n11785), .B(n11786), .Z(n11787) );
  XNOR U12448 ( .A(n11788), .B(n11787), .Z(n11595) );
  NANDN U12449 ( .A(n11524), .B(n11523), .Z(n11528) );
  NAND U12450 ( .A(n11526), .B(n11525), .Z(n11527) );
  NAND U12451 ( .A(n11528), .B(n11527), .Z(n11592) );
  NANDN U12452 ( .A(n11530), .B(n11529), .Z(n11534) );
  NAND U12453 ( .A(n11532), .B(n11531), .Z(n11533) );
  NAND U12454 ( .A(n11534), .B(n11533), .Z(n11593) );
  XNOR U12455 ( .A(n11592), .B(n11593), .Z(n11594) );
  XOR U12456 ( .A(n11595), .B(n11594), .Z(n11818) );
  XOR U12457 ( .A(n11817), .B(n11818), .Z(n11831) );
  XOR U12458 ( .A(n11832), .B(n11831), .Z(n11834) );
  XNOR U12459 ( .A(n11833), .B(n11834), .Z(n11581) );
  XNOR U12460 ( .A(n11580), .B(n11581), .Z(n11582) );
  XNOR U12461 ( .A(n11583), .B(n11582), .Z(n11839) );
  OR U12462 ( .A(n11536), .B(n11535), .Z(n11540) );
  NAND U12463 ( .A(n11538), .B(n11537), .Z(n11539) );
  NAND U12464 ( .A(n11540), .B(n11539), .Z(n11838) );
  NAND U12465 ( .A(n11542), .B(n11541), .Z(n11546) );
  NANDN U12466 ( .A(n11544), .B(n11543), .Z(n11545) );
  NAND U12467 ( .A(n11546), .B(n11545), .Z(n11577) );
  NANDN U12468 ( .A(n11552), .B(n11551), .Z(n11556) );
  NAND U12469 ( .A(n11554), .B(n11553), .Z(n11555) );
  AND U12470 ( .A(n11556), .B(n11555), .Z(n11575) );
  XNOR U12471 ( .A(n11574), .B(n11575), .Z(n11576) );
  XOR U12472 ( .A(n11577), .B(n11576), .Z(n11837) );
  XOR U12473 ( .A(n11838), .B(n11837), .Z(n11840) );
  XNOR U12474 ( .A(n11839), .B(n11840), .Z(n11846) );
  XOR U12475 ( .A(n11845), .B(n11846), .Z(n11852) );
  XOR U12476 ( .A(n11851), .B(n11852), .Z(n11568) );
  NANDN U12477 ( .A(n11558), .B(n11557), .Z(n11562) );
  NAND U12478 ( .A(n11560), .B(n11559), .Z(n11561) );
  AND U12479 ( .A(n11562), .B(n11561), .Z(n11569) );
  XOR U12480 ( .A(n11568), .B(n11569), .Z(n11570) );
  XNOR U12481 ( .A(n11571), .B(n11570), .Z(n11855) );
  XNOR U12482 ( .A(n11855), .B(sreg[132]), .Z(n11857) );
  NAND U12483 ( .A(n11563), .B(sreg[131]), .Z(n11567) );
  OR U12484 ( .A(n11565), .B(n11564), .Z(n11566) );
  AND U12485 ( .A(n11567), .B(n11566), .Z(n11856) );
  XOR U12486 ( .A(n11857), .B(n11856), .Z(c[132]) );
  NAND U12487 ( .A(n11569), .B(n11568), .Z(n11573) );
  NAND U12488 ( .A(n11571), .B(n11570), .Z(n11572) );
  NAND U12489 ( .A(n11573), .B(n11572), .Z(n11863) );
  NANDN U12490 ( .A(n11575), .B(n11574), .Z(n11579) );
  NAND U12491 ( .A(n11577), .B(n11576), .Z(n11578) );
  NAND U12492 ( .A(n11579), .B(n11578), .Z(n12127) );
  NANDN U12493 ( .A(n11581), .B(n11580), .Z(n11585) );
  NAND U12494 ( .A(n11583), .B(n11582), .Z(n11584) );
  NAND U12495 ( .A(n11585), .B(n11584), .Z(n12128) );
  XNOR U12496 ( .A(n12127), .B(n12128), .Z(n12129) );
  NANDN U12497 ( .A(n11587), .B(n11586), .Z(n11591) );
  OR U12498 ( .A(n11589), .B(n11588), .Z(n11590) );
  AND U12499 ( .A(n11591), .B(n11590), .Z(n11883) );
  NANDN U12500 ( .A(n11593), .B(n11592), .Z(n11597) );
  NAND U12501 ( .A(n11595), .B(n11594), .Z(n11596) );
  NAND U12502 ( .A(n11597), .B(n11596), .Z(n11880) );
  NANDN U12503 ( .A(n11599), .B(n11598), .Z(n11603) );
  NAND U12504 ( .A(n11601), .B(n11600), .Z(n11602) );
  NAND U12505 ( .A(n11603), .B(n11602), .Z(n11881) );
  XNOR U12506 ( .A(n11880), .B(n11881), .Z(n11882) );
  XNOR U12507 ( .A(n11883), .B(n11882), .Z(n12103) );
  NANDN U12508 ( .A(n11605), .B(n11604), .Z(n11609) );
  OR U12509 ( .A(n11607), .B(n11606), .Z(n11608) );
  AND U12510 ( .A(n11609), .B(n11608), .Z(n12104) );
  XNOR U12511 ( .A(n12103), .B(n12104), .Z(n12106) );
  NANDN U12512 ( .A(n11611), .B(n11610), .Z(n11615) );
  NAND U12513 ( .A(n11613), .B(n11612), .Z(n11614) );
  NAND U12514 ( .A(n11615), .B(n11614), .Z(n11904) );
  NAND U12515 ( .A(n33283), .B(n11616), .Z(n11618) );
  XOR U12516 ( .A(n33020), .B(n24288), .Z(n11908) );
  NANDN U12517 ( .A(n33021), .B(n11908), .Z(n11617) );
  NAND U12518 ( .A(n11618), .B(n11617), .Z(n11993) );
  XNOR U12519 ( .A(b[21]), .B(a[49]), .Z(n11911) );
  OR U12520 ( .A(n11911), .B(n33634), .Z(n11621) );
  NANDN U12521 ( .A(n11619), .B(n33464), .Z(n11620) );
  NAND U12522 ( .A(n11621), .B(n11620), .Z(n11990) );
  NAND U12523 ( .A(n34044), .B(n11622), .Z(n11624) );
  XOR U12524 ( .A(n34510), .B(n23149), .Z(n11914) );
  NANDN U12525 ( .A(n33867), .B(n11914), .Z(n11623) );
  AND U12526 ( .A(n11624), .B(n11623), .Z(n11991) );
  XNOR U12527 ( .A(n11990), .B(n11991), .Z(n11992) );
  XOR U12528 ( .A(n11993), .B(n11992), .Z(n12027) );
  NANDN U12529 ( .A(n11626), .B(n11625), .Z(n11630) );
  NAND U12530 ( .A(n11628), .B(n11627), .Z(n11629) );
  NAND U12531 ( .A(n11630), .B(n11629), .Z(n12028) );
  XNOR U12532 ( .A(n12027), .B(n12028), .Z(n12030) );
  NAND U12533 ( .A(a[5]), .B(b[63]), .Z(n12020) );
  NANDN U12534 ( .A(n11631), .B(n38369), .Z(n11633) );
  XOR U12535 ( .A(b[61]), .B(n12258), .Z(n11923) );
  OR U12536 ( .A(n11923), .B(n38371), .Z(n11632) );
  NAND U12537 ( .A(n11633), .B(n11632), .Z(n12018) );
  NANDN U12538 ( .A(n11634), .B(n35311), .Z(n11636) );
  XOR U12539 ( .A(b[31]), .B(n20867), .Z(n11926) );
  NANDN U12540 ( .A(n11926), .B(n35313), .Z(n11635) );
  AND U12541 ( .A(n11636), .B(n11635), .Z(n12017) );
  XNOR U12542 ( .A(n12018), .B(n12017), .Z(n12019) );
  XNOR U12543 ( .A(n12020), .B(n12019), .Z(n12029) );
  XNOR U12544 ( .A(n12030), .B(n12029), .Z(n11902) );
  XOR U12545 ( .A(b[13]), .B(n26122), .Z(n11938) );
  OR U12546 ( .A(n11938), .B(n31550), .Z(n11639) );
  NANDN U12547 ( .A(n11637), .B(n31874), .Z(n11638) );
  NAND U12548 ( .A(n11639), .B(n11638), .Z(n12094) );
  NAND U12549 ( .A(n34848), .B(n11640), .Z(n11642) );
  XOR U12550 ( .A(n35375), .B(n21996), .Z(n11941) );
  NAND U12551 ( .A(n34618), .B(n11941), .Z(n11641) );
  NAND U12552 ( .A(n11642), .B(n11641), .Z(n12091) );
  NAND U12553 ( .A(n35188), .B(n11643), .Z(n11645) );
  XOR U12554 ( .A(n35540), .B(n21441), .Z(n11944) );
  NANDN U12555 ( .A(n34968), .B(n11944), .Z(n11644) );
  AND U12556 ( .A(n11645), .B(n11644), .Z(n12092) );
  XNOR U12557 ( .A(n12091), .B(n12092), .Z(n12093) );
  XNOR U12558 ( .A(n12094), .B(n12093), .Z(n11896) );
  XOR U12559 ( .A(b[37]), .B(n19656), .Z(n11929) );
  NANDN U12560 ( .A(n11929), .B(n36311), .Z(n11648) );
  NANDN U12561 ( .A(n11646), .B(n36309), .Z(n11647) );
  NAND U12562 ( .A(n11648), .B(n11647), .Z(n11968) );
  XOR U12563 ( .A(b[5]), .B(n28403), .Z(n11932) );
  OR U12564 ( .A(n11932), .B(n29363), .Z(n11651) );
  NANDN U12565 ( .A(n11649), .B(n29864), .Z(n11650) );
  NAND U12566 ( .A(n11651), .B(n11650), .Z(n11965) );
  XOR U12567 ( .A(n967), .B(n29372), .Z(n11935) );
  NAND U12568 ( .A(n11935), .B(n28939), .Z(n11654) );
  NAND U12569 ( .A(n28938), .B(n11652), .Z(n11653) );
  AND U12570 ( .A(n11654), .B(n11653), .Z(n11966) );
  XNOR U12571 ( .A(n11965), .B(n11966), .Z(n11967) );
  XOR U12572 ( .A(n11968), .B(n11967), .Z(n11897) );
  XOR U12573 ( .A(n11896), .B(n11897), .Z(n11899) );
  NANDN U12574 ( .A(n11656), .B(n11655), .Z(n11660) );
  NAND U12575 ( .A(n11658), .B(n11657), .Z(n11659) );
  NAND U12576 ( .A(n11660), .B(n11659), .Z(n11898) );
  XOR U12577 ( .A(n11899), .B(n11898), .Z(n11903) );
  XOR U12578 ( .A(n11902), .B(n11903), .Z(n11905) );
  XNOR U12579 ( .A(n11904), .B(n11905), .Z(n12004) );
  NANDN U12580 ( .A(n11662), .B(n11661), .Z(n11666) );
  OR U12581 ( .A(n11664), .B(n11663), .Z(n11665) );
  NAND U12582 ( .A(n11666), .B(n11665), .Z(n12003) );
  NANDN U12583 ( .A(n11668), .B(n11667), .Z(n11672) );
  NAND U12584 ( .A(n11670), .B(n11669), .Z(n11671) );
  NAND U12585 ( .A(n11672), .B(n11671), .Z(n11893) );
  NANDN U12586 ( .A(n11674), .B(n11673), .Z(n11678) );
  NAND U12587 ( .A(n11676), .B(n11675), .Z(n11677) );
  NAND U12588 ( .A(n11678), .B(n11677), .Z(n12060) );
  XNOR U12589 ( .A(b[41]), .B(a[29]), .Z(n11971) );
  OR U12590 ( .A(n11971), .B(n36905), .Z(n11681) );
  NANDN U12591 ( .A(n11679), .B(n36807), .Z(n11680) );
  NAND U12592 ( .A(n11681), .B(n11680), .Z(n11999) );
  XOR U12593 ( .A(b[57]), .B(n13509), .Z(n11974) );
  OR U12594 ( .A(n11974), .B(n965), .Z(n11684) );
  NANDN U12595 ( .A(n11682), .B(n38194), .Z(n11683) );
  NAND U12596 ( .A(n11684), .B(n11683), .Z(n11996) );
  NAND U12597 ( .A(n38326), .B(n11685), .Z(n11687) );
  XOR U12598 ( .A(n38400), .B(n12830), .Z(n11977) );
  NANDN U12599 ( .A(n38273), .B(n11977), .Z(n11686) );
  AND U12600 ( .A(n11687), .B(n11686), .Z(n11997) );
  XNOR U12601 ( .A(n11996), .B(n11997), .Z(n11998) );
  XOR U12602 ( .A(n11999), .B(n11998), .Z(n12058) );
  XOR U12603 ( .A(b[33]), .B(n20352), .Z(n11980) );
  NANDN U12604 ( .A(n11980), .B(n35620), .Z(n11690) );
  NANDN U12605 ( .A(n11688), .B(n35621), .Z(n11689) );
  NAND U12606 ( .A(n11690), .B(n11689), .Z(n12072) );
  NANDN U12607 ( .A(n966), .B(a[69]), .Z(n11691) );
  XOR U12608 ( .A(n29232), .B(n11691), .Z(n11693) );
  IV U12609 ( .A(a[68]), .Z(n29868) );
  NANDN U12610 ( .A(n29868), .B(n966), .Z(n11692) );
  AND U12611 ( .A(n11693), .B(n11692), .Z(n12069) );
  XOR U12612 ( .A(b[63]), .B(n11694), .Z(n11987) );
  NANDN U12613 ( .A(n11987), .B(n38422), .Z(n11697) );
  NANDN U12614 ( .A(n11695), .B(n38423), .Z(n11696) );
  AND U12615 ( .A(n11697), .B(n11696), .Z(n12070) );
  XNOR U12616 ( .A(n12069), .B(n12070), .Z(n12071) );
  XNOR U12617 ( .A(n12072), .B(n12071), .Z(n12057) );
  XNOR U12618 ( .A(n12058), .B(n12057), .Z(n12059) );
  XOR U12619 ( .A(n12060), .B(n12059), .Z(n11891) );
  NANDN U12620 ( .A(n11699), .B(n11698), .Z(n11703) );
  NAND U12621 ( .A(n11701), .B(n11700), .Z(n11702) );
  AND U12622 ( .A(n11703), .B(n11702), .Z(n11890) );
  XNOR U12623 ( .A(n11891), .B(n11890), .Z(n11892) );
  XNOR U12624 ( .A(n11893), .B(n11892), .Z(n12002) );
  XNOR U12625 ( .A(n12003), .B(n12002), .Z(n12005) );
  XNOR U12626 ( .A(n12004), .B(n12005), .Z(n12105) );
  XOR U12627 ( .A(n12106), .B(n12105), .Z(n12110) );
  OR U12628 ( .A(n11705), .B(n11704), .Z(n11709) );
  NAND U12629 ( .A(n11707), .B(n11706), .Z(n11708) );
  NAND U12630 ( .A(n11709), .B(n11708), .Z(n11866) );
  XNOR U12631 ( .A(b[35]), .B(a[35]), .Z(n12008) );
  NANDN U12632 ( .A(n12008), .B(n35985), .Z(n11712) );
  NANDN U12633 ( .A(n11710), .B(n35986), .Z(n11711) );
  NAND U12634 ( .A(n11712), .B(n11711), .Z(n12100) );
  XNOR U12635 ( .A(n31123), .B(a[63]), .Z(n12011) );
  NAND U12636 ( .A(n12011), .B(n29949), .Z(n11715) );
  NAND U12637 ( .A(n29948), .B(n11713), .Z(n11714) );
  NAND U12638 ( .A(n11715), .B(n11714), .Z(n12097) );
  XOR U12639 ( .A(b[55]), .B(n13976), .Z(n12014) );
  NANDN U12640 ( .A(n12014), .B(n38075), .Z(n11718) );
  NANDN U12641 ( .A(n11716), .B(n38073), .Z(n11717) );
  AND U12642 ( .A(n11718), .B(n11717), .Z(n12098) );
  XNOR U12643 ( .A(n12097), .B(n12098), .Z(n12099) );
  XNOR U12644 ( .A(n12100), .B(n12099), .Z(n11887) );
  NANDN U12645 ( .A(n11720), .B(n11719), .Z(n11724) );
  NAND U12646 ( .A(n11722), .B(n11721), .Z(n11723) );
  NAND U12647 ( .A(n11724), .B(n11723), .Z(n11884) );
  NANDN U12648 ( .A(n11726), .B(n11725), .Z(n11730) );
  NAND U12649 ( .A(n11728), .B(n11727), .Z(n11729) );
  NAND U12650 ( .A(n11730), .B(n11729), .Z(n11885) );
  XNOR U12651 ( .A(n11884), .B(n11885), .Z(n11886) );
  XOR U12652 ( .A(n11887), .B(n11886), .Z(n11870) );
  OR U12653 ( .A(n11732), .B(n11731), .Z(n11736) );
  OR U12654 ( .A(n11734), .B(n11733), .Z(n11735) );
  NAND U12655 ( .A(n11736), .B(n11735), .Z(n11868) );
  NAND U12656 ( .A(n37652), .B(n11737), .Z(n11739) );
  XOR U12657 ( .A(b[49]), .B(n16220), .Z(n12042) );
  OR U12658 ( .A(n12042), .B(n37756), .Z(n11738) );
  NAND U12659 ( .A(n11739), .B(n11738), .Z(n12025) );
  NANDN U12660 ( .A(n11740), .B(n37469), .Z(n11742) );
  XNOR U12661 ( .A(n978), .B(a[23]), .Z(n12045) );
  NAND U12662 ( .A(n12045), .B(n37471), .Z(n11741) );
  NAND U12663 ( .A(n11742), .B(n11741), .Z(n12023) );
  NAND U12664 ( .A(n30846), .B(n11743), .Z(n11745) );
  XNOR U12665 ( .A(n969), .B(a[61]), .Z(n12048) );
  NAND U12666 ( .A(n30509), .B(n12048), .Z(n11744) );
  NAND U12667 ( .A(n11745), .B(n11744), .Z(n12024) );
  XNOR U12668 ( .A(n12023), .B(n12024), .Z(n12026) );
  XOR U12669 ( .A(n12025), .B(n12026), .Z(n11953) );
  XNOR U12670 ( .A(b[11]), .B(a[59]), .Z(n12033) );
  OR U12671 ( .A(n12033), .B(n31369), .Z(n11748) );
  NANDN U12672 ( .A(n11746), .B(n31119), .Z(n11747) );
  NAND U12673 ( .A(n11748), .B(n11747), .Z(n12054) );
  XOR U12674 ( .A(b[43]), .B(n17960), .Z(n12036) );
  NANDN U12675 ( .A(n12036), .B(n37068), .Z(n11751) );
  NANDN U12676 ( .A(n11749), .B(n37069), .Z(n11750) );
  NAND U12677 ( .A(n11751), .B(n11750), .Z(n12051) );
  XNOR U12678 ( .A(b[45]), .B(a[25]), .Z(n12039) );
  NANDN U12679 ( .A(n12039), .B(n37261), .Z(n11754) );
  NANDN U12680 ( .A(n11752), .B(n37262), .Z(n11753) );
  AND U12681 ( .A(n11754), .B(n11753), .Z(n12052) );
  XNOR U12682 ( .A(n12051), .B(n12052), .Z(n12053) );
  XOR U12683 ( .A(n12054), .B(n12053), .Z(n11954) );
  XNOR U12684 ( .A(n11953), .B(n11954), .Z(n11955) );
  NANDN U12685 ( .A(n11756), .B(n11755), .Z(n11760) );
  NAND U12686 ( .A(n11758), .B(n11757), .Z(n11759) );
  AND U12687 ( .A(n11760), .B(n11759), .Z(n11956) );
  XNOR U12688 ( .A(n11955), .B(n11956), .Z(n11869) );
  XNOR U12689 ( .A(n11868), .B(n11869), .Z(n11871) );
  XOR U12690 ( .A(n11870), .B(n11871), .Z(n11864) );
  XOR U12691 ( .A(b[15]), .B(n25466), .Z(n12073) );
  OR U12692 ( .A(n12073), .B(n32010), .Z(n11763) );
  NANDN U12693 ( .A(n11761), .B(n32011), .Z(n11762) );
  NAND U12694 ( .A(n11763), .B(n11762), .Z(n11920) );
  XNOR U12695 ( .A(b[25]), .B(n22579), .Z(n12076) );
  NANDN U12696 ( .A(n34219), .B(n12076), .Z(n11766) );
  NAND U12697 ( .A(n34217), .B(n11764), .Z(n11765) );
  NAND U12698 ( .A(n11766), .B(n11765), .Z(n11917) );
  XNOR U12699 ( .A(b[17]), .B(a[53]), .Z(n12079) );
  NANDN U12700 ( .A(n12079), .B(n32543), .Z(n11769) );
  NANDN U12701 ( .A(n11767), .B(n32541), .Z(n11768) );
  AND U12702 ( .A(n11769), .B(n11768), .Z(n11918) );
  XNOR U12703 ( .A(n11917), .B(n11918), .Z(n11919) );
  XNOR U12704 ( .A(n11920), .B(n11919), .Z(n11959) );
  XOR U12705 ( .A(b[39]), .B(n18639), .Z(n12082) );
  NANDN U12706 ( .A(n12082), .B(n36553), .Z(n11772) );
  NANDN U12707 ( .A(n11770), .B(n36643), .Z(n11771) );
  NAND U12708 ( .A(n11772), .B(n11771), .Z(n11950) );
  XOR U12709 ( .A(b[51]), .B(n15113), .Z(n12085) );
  NANDN U12710 ( .A(n12085), .B(n37803), .Z(n11775) );
  NANDN U12711 ( .A(n11773), .B(n37802), .Z(n11774) );
  NAND U12712 ( .A(n11775), .B(n11774), .Z(n11947) );
  XOR U12713 ( .A(b[53]), .B(n14514), .Z(n12088) );
  NANDN U12714 ( .A(n12088), .B(n37940), .Z(n11778) );
  NANDN U12715 ( .A(n11776), .B(n37941), .Z(n11777) );
  AND U12716 ( .A(n11778), .B(n11777), .Z(n11948) );
  XNOR U12717 ( .A(n11947), .B(n11948), .Z(n11949) );
  XOR U12718 ( .A(n11950), .B(n11949), .Z(n11960) );
  XNOR U12719 ( .A(n11959), .B(n11960), .Z(n11961) );
  NANDN U12720 ( .A(n11780), .B(n11779), .Z(n11784) );
  NAND U12721 ( .A(n11782), .B(n11781), .Z(n11783) );
  NAND U12722 ( .A(n11784), .B(n11783), .Z(n11962) );
  XOR U12723 ( .A(n11961), .B(n11962), .Z(n12066) );
  NANDN U12724 ( .A(n11786), .B(n11785), .Z(n11790) );
  NAND U12725 ( .A(n11788), .B(n11787), .Z(n11789) );
  NAND U12726 ( .A(n11790), .B(n11789), .Z(n12063) );
  NANDN U12727 ( .A(n11792), .B(n11791), .Z(n11796) );
  NAND U12728 ( .A(n11794), .B(n11793), .Z(n11795) );
  AND U12729 ( .A(n11796), .B(n11795), .Z(n12064) );
  XNOR U12730 ( .A(n12063), .B(n12064), .Z(n12065) );
  XNOR U12731 ( .A(n12066), .B(n12065), .Z(n11874) );
  OR U12732 ( .A(n11798), .B(n11797), .Z(n11802) );
  OR U12733 ( .A(n11800), .B(n11799), .Z(n11801) );
  AND U12734 ( .A(n11802), .B(n11801), .Z(n11875) );
  XNOR U12735 ( .A(n11874), .B(n11875), .Z(n11876) );
  NANDN U12736 ( .A(n11804), .B(n11803), .Z(n11808) );
  NAND U12737 ( .A(n11806), .B(n11805), .Z(n11807) );
  AND U12738 ( .A(n11808), .B(n11807), .Z(n11877) );
  XNOR U12739 ( .A(n11876), .B(n11877), .Z(n11865) );
  XNOR U12740 ( .A(n11864), .B(n11865), .Z(n11867) );
  XNOR U12741 ( .A(n11866), .B(n11867), .Z(n12109) );
  XNOR U12742 ( .A(n12110), .B(n12109), .Z(n12112) );
  OR U12743 ( .A(n11810), .B(n11809), .Z(n11814) );
  NANDN U12744 ( .A(n11812), .B(n11811), .Z(n11813) );
  NAND U12745 ( .A(n11814), .B(n11813), .Z(n12111) );
  XNOR U12746 ( .A(n12112), .B(n12111), .Z(n12124) );
  NANDN U12747 ( .A(n11816), .B(n11815), .Z(n11820) );
  NAND U12748 ( .A(n11818), .B(n11817), .Z(n11819) );
  NAND U12749 ( .A(n11820), .B(n11819), .Z(n12118) );
  NANDN U12750 ( .A(n11822), .B(n11821), .Z(n11826) );
  NAND U12751 ( .A(n11824), .B(n11823), .Z(n11825) );
  NAND U12752 ( .A(n11826), .B(n11825), .Z(n12116) );
  XNOR U12753 ( .A(n12116), .B(n12115), .Z(n12117) );
  XNOR U12754 ( .A(n12118), .B(n12117), .Z(n12121) );
  NANDN U12755 ( .A(n11832), .B(n11831), .Z(n11836) );
  NANDN U12756 ( .A(n11834), .B(n11833), .Z(n11835) );
  AND U12757 ( .A(n11836), .B(n11835), .Z(n12122) );
  XNOR U12758 ( .A(n12124), .B(n12123), .Z(n12130) );
  XOR U12759 ( .A(n12129), .B(n12130), .Z(n12136) );
  NANDN U12760 ( .A(n11838), .B(n11837), .Z(n11842) );
  NANDN U12761 ( .A(n11840), .B(n11839), .Z(n11841) );
  NAND U12762 ( .A(n11842), .B(n11841), .Z(n12134) );
  NANDN U12763 ( .A(n11844), .B(n11843), .Z(n11848) );
  NAND U12764 ( .A(n11846), .B(n11845), .Z(n11847) );
  AND U12765 ( .A(n11848), .B(n11847), .Z(n12133) );
  XNOR U12766 ( .A(n12134), .B(n12133), .Z(n12135) );
  XNOR U12767 ( .A(n12136), .B(n12135), .Z(n11860) );
  NANDN U12768 ( .A(n11850), .B(n11849), .Z(n11854) );
  NAND U12769 ( .A(n11852), .B(n11851), .Z(n11853) );
  AND U12770 ( .A(n11854), .B(n11853), .Z(n11861) );
  XNOR U12771 ( .A(n11860), .B(n11861), .Z(n11862) );
  XNOR U12772 ( .A(n11863), .B(n11862), .Z(n12139) );
  XNOR U12773 ( .A(n12139), .B(sreg[133]), .Z(n12141) );
  NAND U12774 ( .A(n11855), .B(sreg[132]), .Z(n11859) );
  OR U12775 ( .A(n11857), .B(n11856), .Z(n11858) );
  AND U12776 ( .A(n11859), .B(n11858), .Z(n12140) );
  XOR U12777 ( .A(n12141), .B(n12140), .Z(c[133]) );
  NANDN U12778 ( .A(n11869), .B(n11868), .Z(n11873) );
  NAND U12779 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12780 ( .A(n11873), .B(n11872), .Z(n12409) );
  NANDN U12781 ( .A(n11875), .B(n11874), .Z(n11879) );
  NAND U12782 ( .A(n11877), .B(n11876), .Z(n11878) );
  NAND U12783 ( .A(n11879), .B(n11878), .Z(n12407) );
  XNOR U12784 ( .A(n12407), .B(n12406), .Z(n12408) );
  XNOR U12785 ( .A(n12409), .B(n12408), .Z(n12412) );
  XNOR U12786 ( .A(n12413), .B(n12412), .Z(n12414) );
  NANDN U12787 ( .A(n11885), .B(n11884), .Z(n11889) );
  NAND U12788 ( .A(n11887), .B(n11886), .Z(n11888) );
  AND U12789 ( .A(n11889), .B(n11888), .Z(n12380) );
  NANDN U12790 ( .A(n11891), .B(n11890), .Z(n11895) );
  NANDN U12791 ( .A(n11893), .B(n11892), .Z(n11894) );
  NAND U12792 ( .A(n11895), .B(n11894), .Z(n12377) );
  NANDN U12793 ( .A(n11897), .B(n11896), .Z(n11901) );
  OR U12794 ( .A(n11899), .B(n11898), .Z(n11900) );
  AND U12795 ( .A(n11901), .B(n11900), .Z(n12378) );
  XNOR U12796 ( .A(n12377), .B(n12378), .Z(n12379) );
  XNOR U12797 ( .A(n12380), .B(n12379), .Z(n12371) );
  NANDN U12798 ( .A(n11903), .B(n11902), .Z(n11907) );
  OR U12799 ( .A(n11905), .B(n11904), .Z(n11906) );
  AND U12800 ( .A(n11907), .B(n11906), .Z(n12372) );
  XNOR U12801 ( .A(n12371), .B(n12372), .Z(n12374) );
  NAND U12802 ( .A(n33283), .B(n11908), .Z(n11910) );
  XOR U12803 ( .A(n33020), .B(n25134), .Z(n12210) );
  NANDN U12804 ( .A(n33021), .B(n12210), .Z(n11909) );
  NAND U12805 ( .A(n11910), .B(n11909), .Z(n12240) );
  XNOR U12806 ( .A(b[21]), .B(a[50]), .Z(n12213) );
  OR U12807 ( .A(n12213), .B(n33634), .Z(n11913) );
  NANDN U12808 ( .A(n11911), .B(n33464), .Z(n11912) );
  NAND U12809 ( .A(n11913), .B(n11912), .Z(n12237) );
  NAND U12810 ( .A(n34044), .B(n11914), .Z(n11916) );
  XOR U12811 ( .A(n34510), .B(n23447), .Z(n12216) );
  NANDN U12812 ( .A(n33867), .B(n12216), .Z(n11915) );
  AND U12813 ( .A(n11916), .B(n11915), .Z(n12238) );
  XNOR U12814 ( .A(n12237), .B(n12238), .Z(n12239) );
  XOR U12815 ( .A(n12240), .B(n12239), .Z(n12295) );
  NANDN U12816 ( .A(n11918), .B(n11917), .Z(n11922) );
  NAND U12817 ( .A(n11920), .B(n11919), .Z(n11921) );
  NAND U12818 ( .A(n11922), .B(n11921), .Z(n12296) );
  XNOR U12819 ( .A(n12295), .B(n12296), .Z(n12298) );
  NAND U12820 ( .A(a[6]), .B(b[63]), .Z(n12286) );
  NANDN U12821 ( .A(n11923), .B(n38369), .Z(n11925) );
  XOR U12822 ( .A(b[61]), .B(n12555), .Z(n12204) );
  OR U12823 ( .A(n12204), .B(n38371), .Z(n11924) );
  NAND U12824 ( .A(n11925), .B(n11924), .Z(n12284) );
  NANDN U12825 ( .A(n11926), .B(n35311), .Z(n11928) );
  XOR U12826 ( .A(b[31]), .B(n21149), .Z(n12207) );
  NANDN U12827 ( .A(n12207), .B(n35313), .Z(n11927) );
  AND U12828 ( .A(n11928), .B(n11927), .Z(n12283) );
  XNOR U12829 ( .A(n12284), .B(n12283), .Z(n12285) );
  XNOR U12830 ( .A(n12286), .B(n12285), .Z(n12297) );
  XNOR U12831 ( .A(n12298), .B(n12297), .Z(n12150) );
  XOR U12832 ( .A(b[37]), .B(n19513), .Z(n12174) );
  NANDN U12833 ( .A(n12174), .B(n36311), .Z(n11931) );
  NANDN U12834 ( .A(n11929), .B(n36309), .Z(n11930) );
  NAND U12835 ( .A(n11931), .B(n11930), .Z(n12234) );
  XOR U12836 ( .A(b[5]), .B(n28701), .Z(n12177) );
  OR U12837 ( .A(n12177), .B(n29363), .Z(n11934) );
  NANDN U12838 ( .A(n11932), .B(n29864), .Z(n11933) );
  NAND U12839 ( .A(n11934), .B(n11933), .Z(n12231) );
  XOR U12840 ( .A(n967), .B(n29868), .Z(n12180) );
  NAND U12841 ( .A(n12180), .B(n28939), .Z(n11937) );
  NAND U12842 ( .A(n28938), .B(n11935), .Z(n11936) );
  AND U12843 ( .A(n11937), .B(n11936), .Z(n12232) );
  XNOR U12844 ( .A(n12231), .B(n12232), .Z(n12233) );
  XOR U12845 ( .A(n12234), .B(n12233), .Z(n12171) );
  XOR U12846 ( .A(b[13]), .B(n26347), .Z(n12183) );
  OR U12847 ( .A(n12183), .B(n31550), .Z(n11940) );
  NANDN U12848 ( .A(n11938), .B(n31874), .Z(n11939) );
  NAND U12849 ( .A(n11940), .B(n11939), .Z(n12362) );
  NAND U12850 ( .A(n34848), .B(n11941), .Z(n11943) );
  XOR U12851 ( .A(n35375), .B(n22289), .Z(n12186) );
  NAND U12852 ( .A(n34618), .B(n12186), .Z(n11942) );
  NAND U12853 ( .A(n11943), .B(n11942), .Z(n12359) );
  NAND U12854 ( .A(n35188), .B(n11944), .Z(n11946) );
  XOR U12855 ( .A(n35540), .B(n22246), .Z(n12189) );
  NANDN U12856 ( .A(n34968), .B(n12189), .Z(n11945) );
  AND U12857 ( .A(n11946), .B(n11945), .Z(n12360) );
  XNOR U12858 ( .A(n12359), .B(n12360), .Z(n12361) );
  XOR U12859 ( .A(n12362), .B(n12361), .Z(n12169) );
  NANDN U12860 ( .A(n11948), .B(n11947), .Z(n11952) );
  NAND U12861 ( .A(n11950), .B(n11949), .Z(n11951) );
  AND U12862 ( .A(n11952), .B(n11951), .Z(n12168) );
  XOR U12863 ( .A(n12169), .B(n12168), .Z(n12170) );
  XOR U12864 ( .A(n12171), .B(n12170), .Z(n12151) );
  XOR U12865 ( .A(n12150), .B(n12151), .Z(n12153) );
  NANDN U12866 ( .A(n11954), .B(n11953), .Z(n11958) );
  NAND U12867 ( .A(n11956), .B(n11955), .Z(n11957) );
  NAND U12868 ( .A(n11958), .B(n11957), .Z(n12152) );
  XNOR U12869 ( .A(n12153), .B(n12152), .Z(n12270) );
  NANDN U12870 ( .A(n11960), .B(n11959), .Z(n11964) );
  NANDN U12871 ( .A(n11962), .B(n11961), .Z(n11963) );
  NAND U12872 ( .A(n11964), .B(n11963), .Z(n12269) );
  NANDN U12873 ( .A(n11966), .B(n11965), .Z(n11970) );
  NAND U12874 ( .A(n11968), .B(n11967), .Z(n11969) );
  NAND U12875 ( .A(n11970), .B(n11969), .Z(n12165) );
  XNOR U12876 ( .A(b[41]), .B(a[30]), .Z(n12243) );
  OR U12877 ( .A(n12243), .B(n36905), .Z(n11973) );
  NANDN U12878 ( .A(n11971), .B(n36807), .Z(n11972) );
  NAND U12879 ( .A(n11973), .B(n11972), .Z(n12265) );
  XOR U12880 ( .A(b[57]), .B(n14210), .Z(n12246) );
  OR U12881 ( .A(n12246), .B(n965), .Z(n11976) );
  NANDN U12882 ( .A(n11974), .B(n38194), .Z(n11975) );
  NAND U12883 ( .A(n11976), .B(n11975), .Z(n12262) );
  NAND U12884 ( .A(n38326), .B(n11977), .Z(n11979) );
  XOR U12885 ( .A(n38400), .B(n13106), .Z(n12249) );
  NANDN U12886 ( .A(n38273), .B(n12249), .Z(n11978) );
  AND U12887 ( .A(n11979), .B(n11978), .Z(n12263) );
  XNOR U12888 ( .A(n12262), .B(n12263), .Z(n12264) );
  XOR U12889 ( .A(n12265), .B(n12264), .Z(n12331) );
  XOR U12890 ( .A(b[33]), .B(n20686), .Z(n12252) );
  NANDN U12891 ( .A(n12252), .B(n35620), .Z(n11982) );
  NANDN U12892 ( .A(n11980), .B(n35621), .Z(n11981) );
  NAND U12893 ( .A(n11982), .B(n11981), .Z(n12338) );
  NANDN U12894 ( .A(n966), .B(a[70]), .Z(n11983) );
  XOR U12895 ( .A(n29232), .B(n11983), .Z(n11985) );
  NANDN U12896 ( .A(b[0]), .B(a[69]), .Z(n11984) );
  AND U12897 ( .A(n11985), .B(n11984), .Z(n12335) );
  XOR U12898 ( .A(b[63]), .B(n11986), .Z(n12259) );
  NANDN U12899 ( .A(n12259), .B(n38422), .Z(n11989) );
  NANDN U12900 ( .A(n11987), .B(n38423), .Z(n11988) );
  AND U12901 ( .A(n11989), .B(n11988), .Z(n12336) );
  XNOR U12902 ( .A(n12335), .B(n12336), .Z(n12337) );
  XOR U12903 ( .A(n12338), .B(n12337), .Z(n12332) );
  XNOR U12904 ( .A(n12331), .B(n12332), .Z(n12334) );
  NANDN U12905 ( .A(n11991), .B(n11990), .Z(n11995) );
  NAND U12906 ( .A(n11993), .B(n11992), .Z(n11994) );
  AND U12907 ( .A(n11995), .B(n11994), .Z(n12333) );
  XNOR U12908 ( .A(n12334), .B(n12333), .Z(n12162) );
  NANDN U12909 ( .A(n11997), .B(n11996), .Z(n12001) );
  NAND U12910 ( .A(n11999), .B(n11998), .Z(n12000) );
  AND U12911 ( .A(n12001), .B(n12000), .Z(n12163) );
  XOR U12912 ( .A(n12162), .B(n12163), .Z(n12164) );
  XNOR U12913 ( .A(n12165), .B(n12164), .Z(n12268) );
  XNOR U12914 ( .A(n12269), .B(n12268), .Z(n12271) );
  XNOR U12915 ( .A(n12270), .B(n12271), .Z(n12373) );
  XOR U12916 ( .A(n12374), .B(n12373), .Z(n12400) );
  NAND U12917 ( .A(n12003), .B(n12002), .Z(n12007) );
  NANDN U12918 ( .A(n12005), .B(n12004), .Z(n12006) );
  NAND U12919 ( .A(n12007), .B(n12006), .Z(n12396) );
  XNOR U12920 ( .A(b[35]), .B(a[36]), .Z(n12274) );
  NANDN U12921 ( .A(n12274), .B(n35985), .Z(n12010) );
  NANDN U12922 ( .A(n12008), .B(n35986), .Z(n12009) );
  NAND U12923 ( .A(n12010), .B(n12009), .Z(n12368) );
  XNOR U12924 ( .A(n31123), .B(a[64]), .Z(n12277) );
  NAND U12925 ( .A(n12277), .B(n29949), .Z(n12013) );
  NAND U12926 ( .A(n29948), .B(n12011), .Z(n12012) );
  NAND U12927 ( .A(n12013), .B(n12012), .Z(n12365) );
  XOR U12928 ( .A(b[55]), .B(n14259), .Z(n12280) );
  NANDN U12929 ( .A(n12280), .B(n38075), .Z(n12016) );
  NANDN U12930 ( .A(n12014), .B(n38073), .Z(n12015) );
  AND U12931 ( .A(n12016), .B(n12015), .Z(n12366) );
  XNOR U12932 ( .A(n12365), .B(n12366), .Z(n12367) );
  XNOR U12933 ( .A(n12368), .B(n12367), .Z(n12159) );
  NANDN U12934 ( .A(n12018), .B(n12017), .Z(n12022) );
  NAND U12935 ( .A(n12020), .B(n12019), .Z(n12021) );
  NAND U12936 ( .A(n12022), .B(n12021), .Z(n12156) );
  XNOR U12937 ( .A(n12156), .B(n12157), .Z(n12158) );
  XOR U12938 ( .A(n12159), .B(n12158), .Z(n12389) );
  OR U12939 ( .A(n12028), .B(n12027), .Z(n12032) );
  OR U12940 ( .A(n12030), .B(n12029), .Z(n12031) );
  NAND U12941 ( .A(n12032), .B(n12031), .Z(n12387) );
  XOR U12942 ( .A(b[11]), .B(n27436), .Z(n12301) );
  OR U12943 ( .A(n12301), .B(n31369), .Z(n12035) );
  NANDN U12944 ( .A(n12033), .B(n31119), .Z(n12034) );
  NAND U12945 ( .A(n12035), .B(n12034), .Z(n12322) );
  XOR U12946 ( .A(b[43]), .B(n17702), .Z(n12304) );
  NANDN U12947 ( .A(n12304), .B(n37068), .Z(n12038) );
  NANDN U12948 ( .A(n12036), .B(n37069), .Z(n12037) );
  NAND U12949 ( .A(n12038), .B(n12037), .Z(n12319) );
  XNOR U12950 ( .A(b[45]), .B(a[26]), .Z(n12307) );
  NANDN U12951 ( .A(n12307), .B(n37261), .Z(n12041) );
  NANDN U12952 ( .A(n12039), .B(n37262), .Z(n12040) );
  AND U12953 ( .A(n12041), .B(n12040), .Z(n12320) );
  XNOR U12954 ( .A(n12319), .B(n12320), .Z(n12321) );
  XNOR U12955 ( .A(n12322), .B(n12321), .Z(n12219) );
  XOR U12956 ( .A(b[49]), .B(n15963), .Z(n12310) );
  OR U12957 ( .A(n12310), .B(n37756), .Z(n12044) );
  NANDN U12958 ( .A(n12042), .B(n37652), .Z(n12043) );
  NAND U12959 ( .A(n12044), .B(n12043), .Z(n12292) );
  NAND U12960 ( .A(n12045), .B(n37469), .Z(n12047) );
  XOR U12961 ( .A(n978), .B(n16508), .Z(n12313) );
  NAND U12962 ( .A(n12313), .B(n37471), .Z(n12046) );
  NAND U12963 ( .A(n12047), .B(n12046), .Z(n12289) );
  XNOR U12964 ( .A(b[9]), .B(a[62]), .Z(n12316) );
  NANDN U12965 ( .A(n12316), .B(n30509), .Z(n12050) );
  NAND U12966 ( .A(n12048), .B(n30846), .Z(n12049) );
  AND U12967 ( .A(n12050), .B(n12049), .Z(n12290) );
  XNOR U12968 ( .A(n12289), .B(n12290), .Z(n12291) );
  XOR U12969 ( .A(n12292), .B(n12291), .Z(n12220) );
  XNOR U12970 ( .A(n12219), .B(n12220), .Z(n12221) );
  NANDN U12971 ( .A(n12052), .B(n12051), .Z(n12056) );
  NAND U12972 ( .A(n12054), .B(n12053), .Z(n12055) );
  AND U12973 ( .A(n12056), .B(n12055), .Z(n12222) );
  XNOR U12974 ( .A(n12221), .B(n12222), .Z(n12388) );
  XNOR U12975 ( .A(n12387), .B(n12388), .Z(n12390) );
  XOR U12976 ( .A(n12389), .B(n12390), .Z(n12393) );
  NANDN U12977 ( .A(n12058), .B(n12057), .Z(n12062) );
  NANDN U12978 ( .A(n12060), .B(n12059), .Z(n12061) );
  NAND U12979 ( .A(n12062), .B(n12061), .Z(n12381) );
  NANDN U12980 ( .A(n12064), .B(n12063), .Z(n12068) );
  NAND U12981 ( .A(n12066), .B(n12065), .Z(n12067) );
  NAND U12982 ( .A(n12068), .B(n12067), .Z(n12382) );
  XNOR U12983 ( .A(n12381), .B(n12382), .Z(n12383) );
  XOR U12984 ( .A(b[15]), .B(n25860), .Z(n12350) );
  OR U12985 ( .A(n12350), .B(n32010), .Z(n12075) );
  NANDN U12986 ( .A(n12073), .B(n32011), .Z(n12074) );
  NAND U12987 ( .A(n12075), .B(n12074), .Z(n12201) );
  XNOR U12988 ( .A(b[25]), .B(n22964), .Z(n12353) );
  NANDN U12989 ( .A(n34219), .B(n12353), .Z(n12078) );
  NAND U12990 ( .A(n34217), .B(n12076), .Z(n12077) );
  NAND U12991 ( .A(n12078), .B(n12077), .Z(n12198) );
  XNOR U12992 ( .A(b[17]), .B(a[54]), .Z(n12356) );
  NANDN U12993 ( .A(n12356), .B(n32543), .Z(n12081) );
  NANDN U12994 ( .A(n12079), .B(n32541), .Z(n12080) );
  AND U12995 ( .A(n12081), .B(n12080), .Z(n12199) );
  XNOR U12996 ( .A(n12198), .B(n12199), .Z(n12200) );
  XNOR U12997 ( .A(n12201), .B(n12200), .Z(n12225) );
  XOR U12998 ( .A(b[39]), .B(n18841), .Z(n12341) );
  NANDN U12999 ( .A(n12341), .B(n36553), .Z(n12084) );
  NANDN U13000 ( .A(n12082), .B(n36643), .Z(n12083) );
  NAND U13001 ( .A(n12084), .B(n12083), .Z(n12195) );
  XOR U13002 ( .A(b[51]), .B(n15484), .Z(n12344) );
  NANDN U13003 ( .A(n12344), .B(n37803), .Z(n12087) );
  NANDN U13004 ( .A(n12085), .B(n37802), .Z(n12086) );
  NAND U13005 ( .A(n12087), .B(n12086), .Z(n12192) );
  XOR U13006 ( .A(b[53]), .B(n14905), .Z(n12347) );
  NANDN U13007 ( .A(n12347), .B(n37940), .Z(n12090) );
  NANDN U13008 ( .A(n12088), .B(n37941), .Z(n12089) );
  AND U13009 ( .A(n12090), .B(n12089), .Z(n12193) );
  XNOR U13010 ( .A(n12192), .B(n12193), .Z(n12194) );
  XOR U13011 ( .A(n12195), .B(n12194), .Z(n12226) );
  XOR U13012 ( .A(n12225), .B(n12226), .Z(n12228) );
  NANDN U13013 ( .A(n12092), .B(n12091), .Z(n12096) );
  NAND U13014 ( .A(n12094), .B(n12093), .Z(n12095) );
  AND U13015 ( .A(n12096), .B(n12095), .Z(n12227) );
  XOR U13016 ( .A(n12228), .B(n12227), .Z(n12326) );
  NANDN U13017 ( .A(n12098), .B(n12097), .Z(n12102) );
  NAND U13018 ( .A(n12100), .B(n12099), .Z(n12101) );
  AND U13019 ( .A(n12102), .B(n12101), .Z(n12325) );
  XNOR U13020 ( .A(n12326), .B(n12325), .Z(n12327) );
  XOR U13021 ( .A(n12328), .B(n12327), .Z(n12384) );
  XNOR U13022 ( .A(n12383), .B(n12384), .Z(n12394) );
  XOR U13023 ( .A(n12393), .B(n12394), .Z(n12395) );
  XOR U13024 ( .A(n12396), .B(n12395), .Z(n12401) );
  XNOR U13025 ( .A(n12400), .B(n12401), .Z(n12402) );
  NAND U13026 ( .A(n12104), .B(n12103), .Z(n12108) );
  NANDN U13027 ( .A(n12106), .B(n12105), .Z(n12107) );
  AND U13028 ( .A(n12108), .B(n12107), .Z(n12403) );
  XNOR U13029 ( .A(n12402), .B(n12403), .Z(n12415) );
  XNOR U13030 ( .A(n12414), .B(n12415), .Z(n12419) );
  NAND U13031 ( .A(n12110), .B(n12109), .Z(n12114) );
  OR U13032 ( .A(n12112), .B(n12111), .Z(n12113) );
  NAND U13033 ( .A(n12114), .B(n12113), .Z(n12417) );
  NANDN U13034 ( .A(n12116), .B(n12115), .Z(n12120) );
  NANDN U13035 ( .A(n12118), .B(n12117), .Z(n12119) );
  AND U13036 ( .A(n12120), .B(n12119), .Z(n12416) );
  XNOR U13037 ( .A(n12417), .B(n12416), .Z(n12418) );
  XNOR U13038 ( .A(n12419), .B(n12418), .Z(n12425) );
  OR U13039 ( .A(n12122), .B(n12121), .Z(n12126) );
  NAND U13040 ( .A(n12124), .B(n12123), .Z(n12125) );
  NAND U13041 ( .A(n12126), .B(n12125), .Z(n12423) );
  NANDN U13042 ( .A(n12128), .B(n12127), .Z(n12132) );
  NANDN U13043 ( .A(n12130), .B(n12129), .Z(n12131) );
  AND U13044 ( .A(n12132), .B(n12131), .Z(n12422) );
  XNOR U13045 ( .A(n12423), .B(n12422), .Z(n12424) );
  XNOR U13046 ( .A(n12425), .B(n12424), .Z(n12144) );
  NANDN U13047 ( .A(n12134), .B(n12133), .Z(n12138) );
  NAND U13048 ( .A(n12136), .B(n12135), .Z(n12137) );
  NAND U13049 ( .A(n12138), .B(n12137), .Z(n12145) );
  XOR U13050 ( .A(n12144), .B(n12145), .Z(n12146) );
  XNOR U13051 ( .A(n12147), .B(n12146), .Z(n12428) );
  XNOR U13052 ( .A(n12428), .B(sreg[134]), .Z(n12430) );
  NAND U13053 ( .A(n12139), .B(sreg[133]), .Z(n12143) );
  OR U13054 ( .A(n12141), .B(n12140), .Z(n12142) );
  AND U13055 ( .A(n12143), .B(n12142), .Z(n12429) );
  XOR U13056 ( .A(n12430), .B(n12429), .Z(c[134]) );
  OR U13057 ( .A(n12145), .B(n12144), .Z(n12149) );
  NAND U13058 ( .A(n12147), .B(n12146), .Z(n12148) );
  NAND U13059 ( .A(n12149), .B(n12148), .Z(n12436) );
  NANDN U13060 ( .A(n12151), .B(n12150), .Z(n12155) );
  OR U13061 ( .A(n12153), .B(n12152), .Z(n12154) );
  NAND U13062 ( .A(n12155), .B(n12154), .Z(n12666) );
  NANDN U13063 ( .A(n12157), .B(n12156), .Z(n12161) );
  NAND U13064 ( .A(n12159), .B(n12158), .Z(n12160) );
  NAND U13065 ( .A(n12161), .B(n12160), .Z(n12680) );
  NAND U13066 ( .A(n12163), .B(n12162), .Z(n12167) );
  NANDN U13067 ( .A(n12165), .B(n12164), .Z(n12166) );
  NAND U13068 ( .A(n12167), .B(n12166), .Z(n12678) );
  NANDN U13069 ( .A(n12169), .B(n12168), .Z(n12173) );
  OR U13070 ( .A(n12171), .B(n12170), .Z(n12172) );
  AND U13071 ( .A(n12173), .B(n12172), .Z(n12679) );
  XNOR U13072 ( .A(n12678), .B(n12679), .Z(n12681) );
  XNOR U13073 ( .A(n12680), .B(n12681), .Z(n12667) );
  XOR U13074 ( .A(n12666), .B(n12667), .Z(n12668) );
  XOR U13075 ( .A(b[37]), .B(n20315), .Z(n12477) );
  NANDN U13076 ( .A(n12477), .B(n36311), .Z(n12176) );
  NANDN U13077 ( .A(n12174), .B(n36309), .Z(n12175) );
  NAND U13078 ( .A(n12176), .B(n12175), .Z(n12531) );
  XOR U13079 ( .A(b[5]), .B(n29372), .Z(n12480) );
  OR U13080 ( .A(n12480), .B(n29363), .Z(n12179) );
  NANDN U13081 ( .A(n12177), .B(n29864), .Z(n12178) );
  NAND U13082 ( .A(n12179), .B(n12178), .Z(n12528) );
  XNOR U13083 ( .A(n967), .B(a[69]), .Z(n12483) );
  NAND U13084 ( .A(n12483), .B(n28939), .Z(n12182) );
  NAND U13085 ( .A(n28938), .B(n12180), .Z(n12181) );
  AND U13086 ( .A(n12182), .B(n12181), .Z(n12529) );
  XNOR U13087 ( .A(n12528), .B(n12529), .Z(n12530) );
  XNOR U13088 ( .A(n12531), .B(n12530), .Z(n12464) );
  XNOR U13089 ( .A(b[13]), .B(a[59]), .Z(n12486) );
  OR U13090 ( .A(n12486), .B(n31550), .Z(n12185) );
  NANDN U13091 ( .A(n12183), .B(n31874), .Z(n12184) );
  NAND U13092 ( .A(n12185), .B(n12184), .Z(n12592) );
  NAND U13093 ( .A(n34848), .B(n12186), .Z(n12188) );
  XOR U13094 ( .A(n35375), .B(n22579), .Z(n12489) );
  NAND U13095 ( .A(n34618), .B(n12489), .Z(n12187) );
  NAND U13096 ( .A(n12188), .B(n12187), .Z(n12589) );
  NAND U13097 ( .A(n35188), .B(n12189), .Z(n12191) );
  XOR U13098 ( .A(n35540), .B(n21996), .Z(n12492) );
  NANDN U13099 ( .A(n34968), .B(n12492), .Z(n12190) );
  AND U13100 ( .A(n12191), .B(n12190), .Z(n12590) );
  XNOR U13101 ( .A(n12589), .B(n12590), .Z(n12591) );
  XNOR U13102 ( .A(n12592), .B(n12591), .Z(n12461) );
  NANDN U13103 ( .A(n12193), .B(n12192), .Z(n12197) );
  NAND U13104 ( .A(n12195), .B(n12194), .Z(n12196) );
  NAND U13105 ( .A(n12197), .B(n12196), .Z(n12462) );
  XNOR U13106 ( .A(n12461), .B(n12462), .Z(n12463) );
  XOR U13107 ( .A(n12464), .B(n12463), .Z(n12468) );
  NANDN U13108 ( .A(n12199), .B(n12198), .Z(n12203) );
  NAND U13109 ( .A(n12201), .B(n12200), .Z(n12202) );
  NAND U13110 ( .A(n12203), .B(n12202), .Z(n12637) );
  NAND U13111 ( .A(a[7]), .B(b[63]), .Z(n12651) );
  NANDN U13112 ( .A(n12204), .B(n38369), .Z(n12206) );
  XOR U13113 ( .A(b[61]), .B(n12830), .Z(n12507) );
  OR U13114 ( .A(n12507), .B(n38371), .Z(n12205) );
  NAND U13115 ( .A(n12206), .B(n12205), .Z(n12649) );
  NANDN U13116 ( .A(n12207), .B(n35311), .Z(n12209) );
  XOR U13117 ( .A(b[31]), .B(n21441), .Z(n12510) );
  NANDN U13118 ( .A(n12510), .B(n35313), .Z(n12208) );
  AND U13119 ( .A(n12209), .B(n12208), .Z(n12648) );
  XNOR U13120 ( .A(n12649), .B(n12648), .Z(n12650) );
  XOR U13121 ( .A(n12651), .B(n12650), .Z(n12635) );
  NAND U13122 ( .A(n33283), .B(n12210), .Z(n12212) );
  XOR U13123 ( .A(n33020), .B(n25001), .Z(n12513) );
  NANDN U13124 ( .A(n33021), .B(n12513), .Z(n12211) );
  NAND U13125 ( .A(n12212), .B(n12211), .Z(n12537) );
  XNOR U13126 ( .A(b[21]), .B(a[51]), .Z(n12516) );
  OR U13127 ( .A(n12516), .B(n33634), .Z(n12215) );
  NANDN U13128 ( .A(n12213), .B(n33464), .Z(n12214) );
  NAND U13129 ( .A(n12215), .B(n12214), .Z(n12534) );
  NAND U13130 ( .A(n34044), .B(n12216), .Z(n12218) );
  XOR U13131 ( .A(n34510), .B(n23852), .Z(n12519) );
  NANDN U13132 ( .A(n33867), .B(n12519), .Z(n12217) );
  AND U13133 ( .A(n12218), .B(n12217), .Z(n12535) );
  XNOR U13134 ( .A(n12534), .B(n12535), .Z(n12536) );
  XNOR U13135 ( .A(n12537), .B(n12536), .Z(n12636) );
  XNOR U13136 ( .A(n12635), .B(n12636), .Z(n12638) );
  XNOR U13137 ( .A(n12637), .B(n12638), .Z(n12467) );
  XOR U13138 ( .A(n12468), .B(n12467), .Z(n12470) );
  NANDN U13139 ( .A(n12220), .B(n12219), .Z(n12224) );
  NAND U13140 ( .A(n12222), .B(n12221), .Z(n12223) );
  NAND U13141 ( .A(n12224), .B(n12223), .Z(n12469) );
  XNOR U13142 ( .A(n12470), .B(n12469), .Z(n12662) );
  NANDN U13143 ( .A(n12226), .B(n12225), .Z(n12230) );
  NANDN U13144 ( .A(n12228), .B(n12227), .Z(n12229) );
  NAND U13145 ( .A(n12230), .B(n12229), .Z(n12661) );
  NANDN U13146 ( .A(n12232), .B(n12231), .Z(n12236) );
  NAND U13147 ( .A(n12234), .B(n12233), .Z(n12235) );
  NAND U13148 ( .A(n12236), .B(n12235), .Z(n12458) );
  NANDN U13149 ( .A(n12238), .B(n12237), .Z(n12242) );
  NAND U13150 ( .A(n12240), .B(n12239), .Z(n12241) );
  NAND U13151 ( .A(n12242), .B(n12241), .Z(n12608) );
  XNOR U13152 ( .A(b[41]), .B(a[31]), .Z(n12540) );
  OR U13153 ( .A(n12540), .B(n36905), .Z(n12245) );
  NANDN U13154 ( .A(n12243), .B(n36807), .Z(n12244) );
  NAND U13155 ( .A(n12245), .B(n12244), .Z(n12562) );
  XOR U13156 ( .A(b[57]), .B(n13976), .Z(n12543) );
  OR U13157 ( .A(n12543), .B(n965), .Z(n12248) );
  NANDN U13158 ( .A(n12246), .B(n38194), .Z(n12247) );
  NAND U13159 ( .A(n12248), .B(n12247), .Z(n12559) );
  NAND U13160 ( .A(n38326), .B(n12249), .Z(n12251) );
  XOR U13161 ( .A(n38400), .B(n13509), .Z(n12546) );
  NANDN U13162 ( .A(n38273), .B(n12546), .Z(n12250) );
  AND U13163 ( .A(n12251), .B(n12250), .Z(n12560) );
  XNOR U13164 ( .A(n12559), .B(n12560), .Z(n12561) );
  XOR U13165 ( .A(n12562), .B(n12561), .Z(n12606) );
  XOR U13166 ( .A(b[33]), .B(n20867), .Z(n12549) );
  NANDN U13167 ( .A(n12549), .B(n35620), .Z(n12254) );
  NANDN U13168 ( .A(n12252), .B(n35621), .Z(n12253) );
  NAND U13169 ( .A(n12254), .B(n12253), .Z(n12604) );
  NANDN U13170 ( .A(n966), .B(a[71]), .Z(n12255) );
  XOR U13171 ( .A(n29232), .B(n12255), .Z(n12257) );
  IV U13172 ( .A(a[70]), .Z(n30379) );
  NANDN U13173 ( .A(n30379), .B(n966), .Z(n12256) );
  AND U13174 ( .A(n12257), .B(n12256), .Z(n12601) );
  XOR U13175 ( .A(b[63]), .B(n12258), .Z(n12556) );
  NANDN U13176 ( .A(n12556), .B(n38422), .Z(n12261) );
  NANDN U13177 ( .A(n12259), .B(n38423), .Z(n12260) );
  AND U13178 ( .A(n12261), .B(n12260), .Z(n12602) );
  XNOR U13179 ( .A(n12601), .B(n12602), .Z(n12603) );
  XNOR U13180 ( .A(n12604), .B(n12603), .Z(n12605) );
  XNOR U13181 ( .A(n12606), .B(n12605), .Z(n12607) );
  XOR U13182 ( .A(n12608), .B(n12607), .Z(n12456) );
  NANDN U13183 ( .A(n12263), .B(n12262), .Z(n12267) );
  NAND U13184 ( .A(n12265), .B(n12264), .Z(n12266) );
  AND U13185 ( .A(n12267), .B(n12266), .Z(n12455) );
  XNOR U13186 ( .A(n12456), .B(n12455), .Z(n12457) );
  XNOR U13187 ( .A(n12458), .B(n12457), .Z(n12660) );
  XNOR U13188 ( .A(n12661), .B(n12660), .Z(n12663) );
  XNOR U13189 ( .A(n12662), .B(n12663), .Z(n12669) );
  XNOR U13190 ( .A(n12668), .B(n12669), .Z(n12445) );
  NAND U13191 ( .A(n12269), .B(n12268), .Z(n12273) );
  NANDN U13192 ( .A(n12271), .B(n12270), .Z(n12272) );
  NAND U13193 ( .A(n12273), .B(n12272), .Z(n12691) );
  XNOR U13194 ( .A(b[35]), .B(a[37]), .Z(n12639) );
  NANDN U13195 ( .A(n12639), .B(n35985), .Z(n12276) );
  NANDN U13196 ( .A(n12274), .B(n35986), .Z(n12275) );
  NAND U13197 ( .A(n12276), .B(n12275), .Z(n12598) );
  XOR U13198 ( .A(n31123), .B(n28403), .Z(n12642) );
  NAND U13199 ( .A(n12642), .B(n29949), .Z(n12279) );
  NAND U13200 ( .A(n29948), .B(n12277), .Z(n12278) );
  NAND U13201 ( .A(n12279), .B(n12278), .Z(n12595) );
  XOR U13202 ( .A(b[55]), .B(n14514), .Z(n12645) );
  NANDN U13203 ( .A(n12645), .B(n38075), .Z(n12282) );
  NANDN U13204 ( .A(n12280), .B(n38073), .Z(n12281) );
  AND U13205 ( .A(n12282), .B(n12281), .Z(n12596) );
  XNOR U13206 ( .A(n12595), .B(n12596), .Z(n12597) );
  XNOR U13207 ( .A(n12598), .B(n12597), .Z(n12452) );
  NANDN U13208 ( .A(n12284), .B(n12283), .Z(n12288) );
  NAND U13209 ( .A(n12286), .B(n12285), .Z(n12287) );
  NAND U13210 ( .A(n12288), .B(n12287), .Z(n12449) );
  NANDN U13211 ( .A(n12290), .B(n12289), .Z(n12294) );
  NAND U13212 ( .A(n12292), .B(n12291), .Z(n12293) );
  NAND U13213 ( .A(n12294), .B(n12293), .Z(n12450) );
  XNOR U13214 ( .A(n12449), .B(n12450), .Z(n12451) );
  XOR U13215 ( .A(n12452), .B(n12451), .Z(n12674) );
  OR U13216 ( .A(n12296), .B(n12295), .Z(n12300) );
  OR U13217 ( .A(n12298), .B(n12297), .Z(n12299) );
  NAND U13218 ( .A(n12300), .B(n12299), .Z(n12673) );
  XOR U13219 ( .A(b[11]), .B(n27773), .Z(n12611) );
  OR U13220 ( .A(n12611), .B(n31369), .Z(n12303) );
  NANDN U13221 ( .A(n12301), .B(n31119), .Z(n12302) );
  NAND U13222 ( .A(n12303), .B(n12302), .Z(n12632) );
  XOR U13223 ( .A(b[43]), .B(n18003), .Z(n12614) );
  NANDN U13224 ( .A(n12614), .B(n37068), .Z(n12306) );
  NANDN U13225 ( .A(n12304), .B(n37069), .Z(n12305) );
  NAND U13226 ( .A(n12306), .B(n12305), .Z(n12629) );
  XNOR U13227 ( .A(b[45]), .B(a[27]), .Z(n12617) );
  NANDN U13228 ( .A(n12617), .B(n37261), .Z(n12309) );
  NANDN U13229 ( .A(n12307), .B(n37262), .Z(n12308) );
  AND U13230 ( .A(n12309), .B(n12308), .Z(n12630) );
  XNOR U13231 ( .A(n12629), .B(n12630), .Z(n12631) );
  XNOR U13232 ( .A(n12632), .B(n12631), .Z(n12476) );
  XOR U13233 ( .A(b[49]), .B(n16269), .Z(n12620) );
  OR U13234 ( .A(n12620), .B(n37756), .Z(n12312) );
  NANDN U13235 ( .A(n12310), .B(n37652), .Z(n12311) );
  NAND U13236 ( .A(n12312), .B(n12311), .Z(n12657) );
  NAND U13237 ( .A(n37469), .B(n12313), .Z(n12315) );
  XOR U13238 ( .A(n978), .B(n16916), .Z(n12623) );
  NAND U13239 ( .A(n12623), .B(n37471), .Z(n12314) );
  NAND U13240 ( .A(n12315), .B(n12314), .Z(n12654) );
  XNOR U13241 ( .A(b[9]), .B(a[63]), .Z(n12626) );
  NANDN U13242 ( .A(n12626), .B(n30509), .Z(n12318) );
  NANDN U13243 ( .A(n12316), .B(n30846), .Z(n12317) );
  AND U13244 ( .A(n12318), .B(n12317), .Z(n12655) );
  XNOR U13245 ( .A(n12654), .B(n12655), .Z(n12656) );
  XNOR U13246 ( .A(n12657), .B(n12656), .Z(n12473) );
  NANDN U13247 ( .A(n12320), .B(n12319), .Z(n12324) );
  NAND U13248 ( .A(n12322), .B(n12321), .Z(n12323) );
  NAND U13249 ( .A(n12324), .B(n12323), .Z(n12474) );
  XNOR U13250 ( .A(n12473), .B(n12474), .Z(n12475) );
  XOR U13251 ( .A(n12476), .B(n12475), .Z(n12672) );
  XOR U13252 ( .A(n12673), .B(n12672), .Z(n12675) );
  XNOR U13253 ( .A(n12674), .B(n12675), .Z(n12689) );
  NANDN U13254 ( .A(n12326), .B(n12325), .Z(n12330) );
  NANDN U13255 ( .A(n12328), .B(n12327), .Z(n12329) );
  NAND U13256 ( .A(n12330), .B(n12329), .Z(n12682) );
  XNOR U13257 ( .A(n12682), .B(n12683), .Z(n12684) );
  NANDN U13258 ( .A(n12336), .B(n12335), .Z(n12340) );
  NAND U13259 ( .A(n12338), .B(n12337), .Z(n12339) );
  NAND U13260 ( .A(n12340), .B(n12339), .Z(n12568) );
  XOR U13261 ( .A(b[39]), .B(n19656), .Z(n12580) );
  NANDN U13262 ( .A(n12580), .B(n36553), .Z(n12343) );
  NANDN U13263 ( .A(n12341), .B(n36643), .Z(n12342) );
  NAND U13264 ( .A(n12343), .B(n12342), .Z(n12498) );
  XOR U13265 ( .A(b[51]), .B(n16220), .Z(n12583) );
  NANDN U13266 ( .A(n12583), .B(n37803), .Z(n12346) );
  NANDN U13267 ( .A(n12344), .B(n37802), .Z(n12345) );
  NAND U13268 ( .A(n12346), .B(n12345), .Z(n12495) );
  XOR U13269 ( .A(b[53]), .B(n15113), .Z(n12586) );
  NANDN U13270 ( .A(n12586), .B(n37940), .Z(n12349) );
  NANDN U13271 ( .A(n12347), .B(n37941), .Z(n12348) );
  AND U13272 ( .A(n12349), .B(n12348), .Z(n12496) );
  XNOR U13273 ( .A(n12495), .B(n12496), .Z(n12497) );
  XNOR U13274 ( .A(n12498), .B(n12497), .Z(n12524) );
  XOR U13275 ( .A(b[15]), .B(n26122), .Z(n12571) );
  OR U13276 ( .A(n12571), .B(n32010), .Z(n12352) );
  NANDN U13277 ( .A(n12350), .B(n32011), .Z(n12351) );
  NAND U13278 ( .A(n12352), .B(n12351), .Z(n12504) );
  XNOR U13279 ( .A(b[25]), .B(n23149), .Z(n12574) );
  NANDN U13280 ( .A(n34219), .B(n12574), .Z(n12355) );
  NAND U13281 ( .A(n34217), .B(n12353), .Z(n12354) );
  NAND U13282 ( .A(n12355), .B(n12354), .Z(n12501) );
  XNOR U13283 ( .A(b[17]), .B(a[55]), .Z(n12577) );
  NANDN U13284 ( .A(n12577), .B(n32543), .Z(n12358) );
  NANDN U13285 ( .A(n12356), .B(n32541), .Z(n12357) );
  AND U13286 ( .A(n12358), .B(n12357), .Z(n12502) );
  XNOR U13287 ( .A(n12501), .B(n12502), .Z(n12503) );
  XNOR U13288 ( .A(n12504), .B(n12503), .Z(n12522) );
  NANDN U13289 ( .A(n12360), .B(n12359), .Z(n12364) );
  NAND U13290 ( .A(n12362), .B(n12361), .Z(n12363) );
  NAND U13291 ( .A(n12364), .B(n12363), .Z(n12523) );
  XOR U13292 ( .A(n12522), .B(n12523), .Z(n12525) );
  XNOR U13293 ( .A(n12524), .B(n12525), .Z(n12565) );
  NANDN U13294 ( .A(n12366), .B(n12365), .Z(n12370) );
  NAND U13295 ( .A(n12368), .B(n12367), .Z(n12369) );
  AND U13296 ( .A(n12370), .B(n12369), .Z(n12566) );
  XOR U13297 ( .A(n12565), .B(n12566), .Z(n12567) );
  XOR U13298 ( .A(n12568), .B(n12567), .Z(n12685) );
  XNOR U13299 ( .A(n12684), .B(n12685), .Z(n12688) );
  XOR U13300 ( .A(n12691), .B(n12690), .Z(n12446) );
  XNOR U13301 ( .A(n12445), .B(n12446), .Z(n12447) );
  NAND U13302 ( .A(n12372), .B(n12371), .Z(n12376) );
  NANDN U13303 ( .A(n12374), .B(n12373), .Z(n12375) );
  NAND U13304 ( .A(n12376), .B(n12375), .Z(n12448) );
  XOR U13305 ( .A(n12447), .B(n12448), .Z(n12696) );
  NANDN U13306 ( .A(n12382), .B(n12381), .Z(n12386) );
  NANDN U13307 ( .A(n12384), .B(n12383), .Z(n12385) );
  NAND U13308 ( .A(n12386), .B(n12385), .Z(n12439) );
  NANDN U13309 ( .A(n12388), .B(n12387), .Z(n12392) );
  NAND U13310 ( .A(n12390), .B(n12389), .Z(n12391) );
  AND U13311 ( .A(n12392), .B(n12391), .Z(n12440) );
  XNOR U13312 ( .A(n12439), .B(n12440), .Z(n12441) );
  XNOR U13313 ( .A(n12442), .B(n12441), .Z(n12694) );
  NAND U13314 ( .A(n12394), .B(n12393), .Z(n12398) );
  NAND U13315 ( .A(n12396), .B(n12395), .Z(n12397) );
  AND U13316 ( .A(n12398), .B(n12397), .Z(n12695) );
  XOR U13317 ( .A(n12694), .B(n12695), .Z(n12399) );
  XOR U13318 ( .A(n12696), .B(n12399), .Z(n12700) );
  NANDN U13319 ( .A(n12401), .B(n12400), .Z(n12405) );
  NAND U13320 ( .A(n12403), .B(n12402), .Z(n12404) );
  NAND U13321 ( .A(n12405), .B(n12404), .Z(n12698) );
  NANDN U13322 ( .A(n12407), .B(n12406), .Z(n12411) );
  NANDN U13323 ( .A(n12409), .B(n12408), .Z(n12410) );
  AND U13324 ( .A(n12411), .B(n12410), .Z(n12697) );
  XNOR U13325 ( .A(n12698), .B(n12697), .Z(n12699) );
  XOR U13326 ( .A(n12700), .B(n12699), .Z(n12706) );
  NANDN U13327 ( .A(n12417), .B(n12416), .Z(n12421) );
  NANDN U13328 ( .A(n12419), .B(n12418), .Z(n12420) );
  NAND U13329 ( .A(n12421), .B(n12420), .Z(n12704) );
  XNOR U13330 ( .A(n12703), .B(n12704), .Z(n12705) );
  XNOR U13331 ( .A(n12706), .B(n12705), .Z(n12433) );
  NANDN U13332 ( .A(n12423), .B(n12422), .Z(n12427) );
  NANDN U13333 ( .A(n12425), .B(n12424), .Z(n12426) );
  NAND U13334 ( .A(n12427), .B(n12426), .Z(n12434) );
  XOR U13335 ( .A(n12433), .B(n12434), .Z(n12435) );
  XNOR U13336 ( .A(n12436), .B(n12435), .Z(n12709) );
  XNOR U13337 ( .A(n12709), .B(sreg[135]), .Z(n12711) );
  NAND U13338 ( .A(n12428), .B(sreg[134]), .Z(n12432) );
  OR U13339 ( .A(n12430), .B(n12429), .Z(n12431) );
  AND U13340 ( .A(n12432), .B(n12431), .Z(n12710) );
  XOR U13341 ( .A(n12711), .B(n12710), .Z(c[135]) );
  OR U13342 ( .A(n12434), .B(n12433), .Z(n12438) );
  NAND U13343 ( .A(n12436), .B(n12435), .Z(n12437) );
  NAND U13344 ( .A(n12438), .B(n12437), .Z(n12717) );
  NANDN U13345 ( .A(n12440), .B(n12439), .Z(n12444) );
  NAND U13346 ( .A(n12442), .B(n12441), .Z(n12443) );
  NAND U13347 ( .A(n12444), .B(n12443), .Z(n12979) );
  XNOR U13348 ( .A(n12979), .B(n12980), .Z(n12981) );
  NANDN U13349 ( .A(n12450), .B(n12449), .Z(n12454) );
  NAND U13350 ( .A(n12452), .B(n12451), .Z(n12453) );
  AND U13351 ( .A(n12454), .B(n12453), .Z(n12962) );
  NANDN U13352 ( .A(n12456), .B(n12455), .Z(n12460) );
  NANDN U13353 ( .A(n12458), .B(n12457), .Z(n12459) );
  NAND U13354 ( .A(n12460), .B(n12459), .Z(n12959) );
  NANDN U13355 ( .A(n12462), .B(n12461), .Z(n12466) );
  NAND U13356 ( .A(n12464), .B(n12463), .Z(n12465) );
  AND U13357 ( .A(n12466), .B(n12465), .Z(n12960) );
  XNOR U13358 ( .A(n12959), .B(n12960), .Z(n12961) );
  XNOR U13359 ( .A(n12962), .B(n12961), .Z(n12947) );
  NANDN U13360 ( .A(n12468), .B(n12467), .Z(n12472) );
  OR U13361 ( .A(n12470), .B(n12469), .Z(n12471) );
  AND U13362 ( .A(n12472), .B(n12471), .Z(n12948) );
  XNOR U13363 ( .A(n12947), .B(n12948), .Z(n12950) );
  XOR U13364 ( .A(b[37]), .B(n19980), .Z(n12788) );
  NANDN U13365 ( .A(n12788), .B(n36311), .Z(n12479) );
  NANDN U13366 ( .A(n12477), .B(n36309), .Z(n12478) );
  NAND U13367 ( .A(n12479), .B(n12478), .Z(n12812) );
  XOR U13368 ( .A(b[5]), .B(n29868), .Z(n12791) );
  OR U13369 ( .A(n12791), .B(n29363), .Z(n12482) );
  NANDN U13370 ( .A(n12480), .B(n29864), .Z(n12481) );
  NAND U13371 ( .A(n12482), .B(n12481), .Z(n12809) );
  XOR U13372 ( .A(n30379), .B(n967), .Z(n12794) );
  NAND U13373 ( .A(n12794), .B(n28939), .Z(n12485) );
  NAND U13374 ( .A(n28938), .B(n12483), .Z(n12484) );
  AND U13375 ( .A(n12485), .B(n12484), .Z(n12810) );
  XNOR U13376 ( .A(n12809), .B(n12810), .Z(n12811) );
  XNOR U13377 ( .A(n12812), .B(n12811), .Z(n12745) );
  XOR U13378 ( .A(b[13]), .B(n27436), .Z(n12779) );
  OR U13379 ( .A(n12779), .B(n31550), .Z(n12488) );
  NANDN U13380 ( .A(n12486), .B(n31874), .Z(n12487) );
  NAND U13381 ( .A(n12488), .B(n12487), .Z(n12938) );
  NAND U13382 ( .A(n34848), .B(n12489), .Z(n12491) );
  XOR U13383 ( .A(n35375), .B(n22964), .Z(n12782) );
  NAND U13384 ( .A(n34618), .B(n12782), .Z(n12490) );
  NAND U13385 ( .A(n12491), .B(n12490), .Z(n12935) );
  NAND U13386 ( .A(n35188), .B(n12492), .Z(n12494) );
  XOR U13387 ( .A(n35540), .B(n22289), .Z(n12785) );
  NANDN U13388 ( .A(n34968), .B(n12785), .Z(n12493) );
  AND U13389 ( .A(n12494), .B(n12493), .Z(n12936) );
  XNOR U13390 ( .A(n12935), .B(n12936), .Z(n12937) );
  XNOR U13391 ( .A(n12938), .B(n12937), .Z(n12742) );
  NANDN U13392 ( .A(n12496), .B(n12495), .Z(n12500) );
  NAND U13393 ( .A(n12498), .B(n12497), .Z(n12499) );
  NAND U13394 ( .A(n12500), .B(n12499), .Z(n12743) );
  XNOR U13395 ( .A(n12742), .B(n12743), .Z(n12744) );
  XOR U13396 ( .A(n12745), .B(n12744), .Z(n12749) );
  NANDN U13397 ( .A(n12502), .B(n12501), .Z(n12506) );
  NAND U13398 ( .A(n12504), .B(n12503), .Z(n12505) );
  NAND U13399 ( .A(n12506), .B(n12505), .Z(n12878) );
  NAND U13400 ( .A(a[8]), .B(b[63]), .Z(n12892) );
  NANDN U13401 ( .A(n12507), .B(n38369), .Z(n12509) );
  XOR U13402 ( .A(b[61]), .B(n13106), .Z(n12773) );
  OR U13403 ( .A(n12773), .B(n38371), .Z(n12508) );
  NAND U13404 ( .A(n12509), .B(n12508), .Z(n12890) );
  NANDN U13405 ( .A(n12510), .B(n35311), .Z(n12512) );
  XOR U13406 ( .A(b[31]), .B(n22246), .Z(n12776) );
  NANDN U13407 ( .A(n12776), .B(n35313), .Z(n12511) );
  AND U13408 ( .A(n12512), .B(n12511), .Z(n12889) );
  XNOR U13409 ( .A(n12890), .B(n12889), .Z(n12891) );
  XOR U13410 ( .A(n12892), .B(n12891), .Z(n12876) );
  NAND U13411 ( .A(n33283), .B(n12513), .Z(n12515) );
  XOR U13412 ( .A(n33020), .B(n25177), .Z(n12758) );
  NANDN U13413 ( .A(n33021), .B(n12758), .Z(n12514) );
  NAND U13414 ( .A(n12515), .B(n12514), .Z(n12837) );
  XNOR U13415 ( .A(b[21]), .B(a[52]), .Z(n12761) );
  OR U13416 ( .A(n12761), .B(n33634), .Z(n12518) );
  NANDN U13417 ( .A(n12516), .B(n33464), .Z(n12517) );
  NAND U13418 ( .A(n12518), .B(n12517), .Z(n12834) );
  NAND U13419 ( .A(n34044), .B(n12519), .Z(n12521) );
  XOR U13420 ( .A(n34510), .B(n24671), .Z(n12764) );
  NANDN U13421 ( .A(n33867), .B(n12764), .Z(n12520) );
  AND U13422 ( .A(n12521), .B(n12520), .Z(n12835) );
  XNOR U13423 ( .A(n12834), .B(n12835), .Z(n12836) );
  XNOR U13424 ( .A(n12837), .B(n12836), .Z(n12877) );
  XNOR U13425 ( .A(n12876), .B(n12877), .Z(n12879) );
  XNOR U13426 ( .A(n12878), .B(n12879), .Z(n12748) );
  XOR U13427 ( .A(n12749), .B(n12748), .Z(n12751) );
  XNOR U13428 ( .A(n12750), .B(n12751), .Z(n12848) );
  NANDN U13429 ( .A(n12523), .B(n12522), .Z(n12527) );
  NANDN U13430 ( .A(n12525), .B(n12524), .Z(n12526) );
  NAND U13431 ( .A(n12527), .B(n12526), .Z(n12847) );
  NANDN U13432 ( .A(n12529), .B(n12528), .Z(n12533) );
  NAND U13433 ( .A(n12531), .B(n12530), .Z(n12532) );
  NAND U13434 ( .A(n12533), .B(n12532), .Z(n12739) );
  NANDN U13435 ( .A(n12535), .B(n12534), .Z(n12539) );
  NAND U13436 ( .A(n12537), .B(n12536), .Z(n12538) );
  NAND U13437 ( .A(n12539), .B(n12538), .Z(n12904) );
  XNOR U13438 ( .A(b[41]), .B(a[32]), .Z(n12815) );
  OR U13439 ( .A(n12815), .B(n36905), .Z(n12542) );
  NANDN U13440 ( .A(n12540), .B(n36807), .Z(n12541) );
  NAND U13441 ( .A(n12542), .B(n12541), .Z(n12843) );
  XOR U13442 ( .A(b[57]), .B(n14259), .Z(n12818) );
  OR U13443 ( .A(n12818), .B(n965), .Z(n12545) );
  NANDN U13444 ( .A(n12543), .B(n38194), .Z(n12544) );
  NAND U13445 ( .A(n12545), .B(n12544), .Z(n12840) );
  NAND U13446 ( .A(n38326), .B(n12546), .Z(n12548) );
  XOR U13447 ( .A(n38400), .B(n14210), .Z(n12821) );
  NANDN U13448 ( .A(n38273), .B(n12821), .Z(n12547) );
  AND U13449 ( .A(n12548), .B(n12547), .Z(n12841) );
  XNOR U13450 ( .A(n12840), .B(n12841), .Z(n12842) );
  XOR U13451 ( .A(n12843), .B(n12842), .Z(n12902) );
  XOR U13452 ( .A(b[33]), .B(n21149), .Z(n12824) );
  NANDN U13453 ( .A(n12824), .B(n35620), .Z(n12551) );
  NANDN U13454 ( .A(n12549), .B(n35621), .Z(n12550) );
  NAND U13455 ( .A(n12551), .B(n12550), .Z(n12916) );
  NANDN U13456 ( .A(n966), .B(a[72]), .Z(n12552) );
  XOR U13457 ( .A(n29232), .B(n12552), .Z(n12554) );
  IV U13458 ( .A(a[71]), .Z(n30543) );
  NANDN U13459 ( .A(n30543), .B(n966), .Z(n12553) );
  AND U13460 ( .A(n12554), .B(n12553), .Z(n12913) );
  XOR U13461 ( .A(b[63]), .B(n12555), .Z(n12831) );
  NANDN U13462 ( .A(n12831), .B(n38422), .Z(n12558) );
  NANDN U13463 ( .A(n12556), .B(n38423), .Z(n12557) );
  AND U13464 ( .A(n12558), .B(n12557), .Z(n12914) );
  XNOR U13465 ( .A(n12913), .B(n12914), .Z(n12915) );
  XNOR U13466 ( .A(n12916), .B(n12915), .Z(n12901) );
  XNOR U13467 ( .A(n12902), .B(n12901), .Z(n12903) );
  XOR U13468 ( .A(n12904), .B(n12903), .Z(n12737) );
  NANDN U13469 ( .A(n12560), .B(n12559), .Z(n12564) );
  NAND U13470 ( .A(n12562), .B(n12561), .Z(n12563) );
  AND U13471 ( .A(n12564), .B(n12563), .Z(n12736) );
  XNOR U13472 ( .A(n12737), .B(n12736), .Z(n12738) );
  XNOR U13473 ( .A(n12739), .B(n12738), .Z(n12846) );
  XNOR U13474 ( .A(n12847), .B(n12846), .Z(n12849) );
  XNOR U13475 ( .A(n12848), .B(n12849), .Z(n12949) );
  XOR U13476 ( .A(n12950), .B(n12949), .Z(n12718) );
  NAND U13477 ( .A(n12566), .B(n12565), .Z(n12570) );
  NANDN U13478 ( .A(n12568), .B(n12567), .Z(n12569) );
  NAND U13479 ( .A(n12570), .B(n12569), .Z(n12966) );
  XOR U13480 ( .A(b[15]), .B(n26347), .Z(n12917) );
  OR U13481 ( .A(n12917), .B(n32010), .Z(n12573) );
  NANDN U13482 ( .A(n12571), .B(n32011), .Z(n12572) );
  NAND U13483 ( .A(n12573), .B(n12572), .Z(n12770) );
  XNOR U13484 ( .A(b[25]), .B(n23447), .Z(n12920) );
  NANDN U13485 ( .A(n34219), .B(n12920), .Z(n12576) );
  NAND U13486 ( .A(n34217), .B(n12574), .Z(n12575) );
  NAND U13487 ( .A(n12576), .B(n12575), .Z(n12767) );
  XNOR U13488 ( .A(b[17]), .B(a[56]), .Z(n12923) );
  NANDN U13489 ( .A(n12923), .B(n32543), .Z(n12579) );
  NANDN U13490 ( .A(n12577), .B(n32541), .Z(n12578) );
  AND U13491 ( .A(n12579), .B(n12578), .Z(n12768) );
  XNOR U13492 ( .A(n12767), .B(n12768), .Z(n12769) );
  XNOR U13493 ( .A(n12770), .B(n12769), .Z(n12803) );
  XOR U13494 ( .A(b[39]), .B(n19513), .Z(n12926) );
  NANDN U13495 ( .A(n12926), .B(n36553), .Z(n12582) );
  NANDN U13496 ( .A(n12580), .B(n36643), .Z(n12581) );
  NAND U13497 ( .A(n12582), .B(n12581), .Z(n12800) );
  XOR U13498 ( .A(b[51]), .B(n15963), .Z(n12929) );
  NANDN U13499 ( .A(n12929), .B(n37803), .Z(n12585) );
  NANDN U13500 ( .A(n12583), .B(n37802), .Z(n12584) );
  NAND U13501 ( .A(n12585), .B(n12584), .Z(n12797) );
  XOR U13502 ( .A(b[53]), .B(n15484), .Z(n12932) );
  NANDN U13503 ( .A(n12932), .B(n37940), .Z(n12588) );
  NANDN U13504 ( .A(n12586), .B(n37941), .Z(n12587) );
  AND U13505 ( .A(n12588), .B(n12587), .Z(n12798) );
  XNOR U13506 ( .A(n12797), .B(n12798), .Z(n12799) );
  XOR U13507 ( .A(n12800), .B(n12799), .Z(n12804) );
  XNOR U13508 ( .A(n12803), .B(n12804), .Z(n12805) );
  NANDN U13509 ( .A(n12590), .B(n12589), .Z(n12594) );
  NAND U13510 ( .A(n12592), .B(n12591), .Z(n12593) );
  NAND U13511 ( .A(n12594), .B(n12593), .Z(n12806) );
  XOR U13512 ( .A(n12805), .B(n12806), .Z(n12910) );
  NANDN U13513 ( .A(n12596), .B(n12595), .Z(n12600) );
  NAND U13514 ( .A(n12598), .B(n12597), .Z(n12599) );
  NAND U13515 ( .A(n12600), .B(n12599), .Z(n12907) );
  XNOR U13516 ( .A(n12907), .B(n12908), .Z(n12909) );
  XNOR U13517 ( .A(n12910), .B(n12909), .Z(n12963) );
  NANDN U13518 ( .A(n12606), .B(n12605), .Z(n12610) );
  NANDN U13519 ( .A(n12608), .B(n12607), .Z(n12609) );
  AND U13520 ( .A(n12610), .B(n12609), .Z(n12964) );
  XNOR U13521 ( .A(n12963), .B(n12964), .Z(n12965) );
  XNOR U13522 ( .A(n12966), .B(n12965), .Z(n12967) );
  XNOR U13523 ( .A(b[11]), .B(a[62]), .Z(n12852) );
  OR U13524 ( .A(n12852), .B(n31369), .Z(n12613) );
  NANDN U13525 ( .A(n12611), .B(n31119), .Z(n12612) );
  NAND U13526 ( .A(n12613), .B(n12612), .Z(n12873) );
  XOR U13527 ( .A(b[43]), .B(n18804), .Z(n12855) );
  NANDN U13528 ( .A(n12855), .B(n37068), .Z(n12616) );
  NANDN U13529 ( .A(n12614), .B(n37069), .Z(n12615) );
  NAND U13530 ( .A(n12616), .B(n12615), .Z(n12870) );
  XNOR U13531 ( .A(b[45]), .B(a[28]), .Z(n12858) );
  NANDN U13532 ( .A(n12858), .B(n37261), .Z(n12619) );
  NANDN U13533 ( .A(n12617), .B(n37262), .Z(n12618) );
  AND U13534 ( .A(n12619), .B(n12618), .Z(n12871) );
  XNOR U13535 ( .A(n12870), .B(n12871), .Z(n12872) );
  XNOR U13536 ( .A(n12873), .B(n12872), .Z(n12757) );
  XOR U13537 ( .A(b[49]), .B(n16508), .Z(n12861) );
  OR U13538 ( .A(n12861), .B(n37756), .Z(n12622) );
  NANDN U13539 ( .A(n12620), .B(n37652), .Z(n12621) );
  NAND U13540 ( .A(n12622), .B(n12621), .Z(n12897) );
  NAND U13541 ( .A(n37469), .B(n12623), .Z(n12625) );
  XOR U13542 ( .A(n978), .B(n17133), .Z(n12864) );
  NAND U13543 ( .A(n12864), .B(n37471), .Z(n12624) );
  AND U13544 ( .A(n12625), .B(n12624), .Z(n12895) );
  XNOR U13545 ( .A(b[9]), .B(a[64]), .Z(n12867) );
  NANDN U13546 ( .A(n12867), .B(n30509), .Z(n12628) );
  NANDN U13547 ( .A(n12626), .B(n30846), .Z(n12627) );
  AND U13548 ( .A(n12628), .B(n12627), .Z(n12896) );
  XOR U13549 ( .A(n12897), .B(n12898), .Z(n12754) );
  NANDN U13550 ( .A(n12630), .B(n12629), .Z(n12634) );
  NAND U13551 ( .A(n12632), .B(n12631), .Z(n12633) );
  NAND U13552 ( .A(n12634), .B(n12633), .Z(n12755) );
  XNOR U13553 ( .A(n12754), .B(n12755), .Z(n12756) );
  XOR U13554 ( .A(n12757), .B(n12756), .Z(n12953) );
  XNOR U13555 ( .A(n12953), .B(n12954), .Z(n12956) );
  XNOR U13556 ( .A(b[35]), .B(a[38]), .Z(n12880) );
  NANDN U13557 ( .A(n12880), .B(n35985), .Z(n12641) );
  NANDN U13558 ( .A(n12639), .B(n35986), .Z(n12640) );
  NAND U13559 ( .A(n12641), .B(n12640), .Z(n12944) );
  XOR U13560 ( .A(n31123), .B(n28701), .Z(n12883) );
  NAND U13561 ( .A(n12883), .B(n29949), .Z(n12644) );
  NAND U13562 ( .A(n29948), .B(n12642), .Z(n12643) );
  NAND U13563 ( .A(n12644), .B(n12643), .Z(n12941) );
  XOR U13564 ( .A(b[55]), .B(n14905), .Z(n12886) );
  NANDN U13565 ( .A(n12886), .B(n38075), .Z(n12647) );
  NANDN U13566 ( .A(n12645), .B(n38073), .Z(n12646) );
  AND U13567 ( .A(n12647), .B(n12646), .Z(n12942) );
  XNOR U13568 ( .A(n12941), .B(n12942), .Z(n12943) );
  XNOR U13569 ( .A(n12944), .B(n12943), .Z(n12733) );
  NANDN U13570 ( .A(n12649), .B(n12648), .Z(n12653) );
  NAND U13571 ( .A(n12651), .B(n12650), .Z(n12652) );
  NAND U13572 ( .A(n12653), .B(n12652), .Z(n12730) );
  NANDN U13573 ( .A(n12655), .B(n12654), .Z(n12659) );
  NAND U13574 ( .A(n12657), .B(n12656), .Z(n12658) );
  NAND U13575 ( .A(n12659), .B(n12658), .Z(n12731) );
  XNOR U13576 ( .A(n12730), .B(n12731), .Z(n12732) );
  XOR U13577 ( .A(n12733), .B(n12732), .Z(n12955) );
  XNOR U13578 ( .A(n12956), .B(n12955), .Z(n12968) );
  XOR U13579 ( .A(n12967), .B(n12968), .Z(n12970) );
  NAND U13580 ( .A(n12661), .B(n12660), .Z(n12665) );
  NANDN U13581 ( .A(n12663), .B(n12662), .Z(n12664) );
  AND U13582 ( .A(n12665), .B(n12664), .Z(n12969) );
  XOR U13583 ( .A(n12970), .B(n12969), .Z(n12719) );
  XNOR U13584 ( .A(n12718), .B(n12719), .Z(n12720) );
  OR U13585 ( .A(n12667), .B(n12666), .Z(n12671) );
  NAND U13586 ( .A(n12669), .B(n12668), .Z(n12670) );
  NAND U13587 ( .A(n12671), .B(n12670), .Z(n12721) );
  XOR U13588 ( .A(n12720), .B(n12721), .Z(n12976) );
  NAND U13589 ( .A(n12673), .B(n12672), .Z(n12677) );
  NAND U13590 ( .A(n12675), .B(n12674), .Z(n12676) );
  NAND U13591 ( .A(n12677), .B(n12676), .Z(n12727) );
  NANDN U13592 ( .A(n12683), .B(n12682), .Z(n12687) );
  NANDN U13593 ( .A(n12685), .B(n12684), .Z(n12686) );
  AND U13594 ( .A(n12687), .B(n12686), .Z(n12724) );
  XNOR U13595 ( .A(n12725), .B(n12724), .Z(n12726) );
  XNOR U13596 ( .A(n12727), .B(n12726), .Z(n12973) );
  NANDN U13597 ( .A(n12689), .B(n12688), .Z(n12693) );
  NAND U13598 ( .A(n12691), .B(n12690), .Z(n12692) );
  AND U13599 ( .A(n12693), .B(n12692), .Z(n12974) );
  XNOR U13600 ( .A(n12976), .B(n12975), .Z(n12982) );
  XOR U13601 ( .A(n12981), .B(n12982), .Z(n12988) );
  NANDN U13602 ( .A(n12698), .B(n12697), .Z(n12702) );
  NAND U13603 ( .A(n12700), .B(n12699), .Z(n12701) );
  NAND U13604 ( .A(n12702), .B(n12701), .Z(n12986) );
  XNOR U13605 ( .A(n12985), .B(n12986), .Z(n12987) );
  XNOR U13606 ( .A(n12988), .B(n12987), .Z(n12714) );
  NANDN U13607 ( .A(n12704), .B(n12703), .Z(n12708) );
  NANDN U13608 ( .A(n12706), .B(n12705), .Z(n12707) );
  NAND U13609 ( .A(n12708), .B(n12707), .Z(n12715) );
  XNOR U13610 ( .A(n12714), .B(n12715), .Z(n12716) );
  XNOR U13611 ( .A(n12717), .B(n12716), .Z(n12989) );
  XNOR U13612 ( .A(n12989), .B(sreg[136]), .Z(n12991) );
  NAND U13613 ( .A(n12709), .B(sreg[135]), .Z(n12713) );
  OR U13614 ( .A(n12711), .B(n12710), .Z(n12712) );
  AND U13615 ( .A(n12713), .B(n12712), .Z(n12990) );
  XOR U13616 ( .A(n12991), .B(n12990), .Z(c[136]) );
  NANDN U13617 ( .A(n12719), .B(n12718), .Z(n12723) );
  NANDN U13618 ( .A(n12721), .B(n12720), .Z(n12722) );
  NAND U13619 ( .A(n12723), .B(n12722), .Z(n13268) );
  NANDN U13620 ( .A(n12725), .B(n12724), .Z(n12729) );
  NANDN U13621 ( .A(n12727), .B(n12726), .Z(n12728) );
  AND U13622 ( .A(n12729), .B(n12728), .Z(n13267) );
  XNOR U13623 ( .A(n13268), .B(n13267), .Z(n13269) );
  NANDN U13624 ( .A(n12731), .B(n12730), .Z(n12735) );
  NAND U13625 ( .A(n12733), .B(n12732), .Z(n12734) );
  AND U13626 ( .A(n12735), .B(n12734), .Z(n13236) );
  NANDN U13627 ( .A(n12737), .B(n12736), .Z(n12741) );
  NANDN U13628 ( .A(n12739), .B(n12738), .Z(n12740) );
  NAND U13629 ( .A(n12741), .B(n12740), .Z(n13233) );
  NANDN U13630 ( .A(n12743), .B(n12742), .Z(n12747) );
  NAND U13631 ( .A(n12745), .B(n12744), .Z(n12746) );
  AND U13632 ( .A(n12747), .B(n12746), .Z(n13234) );
  XNOR U13633 ( .A(n13233), .B(n13234), .Z(n13235) );
  XNOR U13634 ( .A(n13236), .B(n13235), .Z(n13221) );
  NANDN U13635 ( .A(n12749), .B(n12748), .Z(n12753) );
  OR U13636 ( .A(n12751), .B(n12750), .Z(n12752) );
  AND U13637 ( .A(n12753), .B(n12752), .Z(n13222) );
  XNOR U13638 ( .A(n13221), .B(n13222), .Z(n13224) );
  NAND U13639 ( .A(n33283), .B(n12758), .Z(n12760) );
  XOR U13640 ( .A(n33020), .B(n25466), .Z(n13064) );
  NANDN U13641 ( .A(n33021), .B(n13064), .Z(n12759) );
  NAND U13642 ( .A(n12760), .B(n12759), .Z(n13088) );
  XNOR U13643 ( .A(b[21]), .B(a[53]), .Z(n13067) );
  OR U13644 ( .A(n13067), .B(n33634), .Z(n12763) );
  NANDN U13645 ( .A(n12761), .B(n33464), .Z(n12762) );
  NAND U13646 ( .A(n12763), .B(n12762), .Z(n13085) );
  NAND U13647 ( .A(n34044), .B(n12764), .Z(n12766) );
  XOR U13648 ( .A(n34510), .B(n24288), .Z(n13070) );
  NANDN U13649 ( .A(n33867), .B(n13070), .Z(n12765) );
  AND U13650 ( .A(n12766), .B(n12765), .Z(n13086) );
  XNOR U13651 ( .A(n13085), .B(n13086), .Z(n13087) );
  XNOR U13652 ( .A(n13088), .B(n13087), .Z(n13185) );
  NANDN U13653 ( .A(n12768), .B(n12767), .Z(n12772) );
  NAND U13654 ( .A(n12770), .B(n12769), .Z(n12771) );
  NAND U13655 ( .A(n12772), .B(n12771), .Z(n13186) );
  XNOR U13656 ( .A(n13185), .B(n13186), .Z(n13187) );
  NAND U13657 ( .A(a[9]), .B(b[63]), .Z(n13176) );
  NANDN U13658 ( .A(n12773), .B(n38369), .Z(n12775) );
  XOR U13659 ( .A(b[61]), .B(n13509), .Z(n13058) );
  OR U13660 ( .A(n13058), .B(n38371), .Z(n12774) );
  NAND U13661 ( .A(n12775), .B(n12774), .Z(n13174) );
  NANDN U13662 ( .A(n12776), .B(n35311), .Z(n12778) );
  XOR U13663 ( .A(b[31]), .B(n21996), .Z(n13061) );
  NANDN U13664 ( .A(n13061), .B(n35313), .Z(n12777) );
  AND U13665 ( .A(n12778), .B(n12777), .Z(n13173) );
  XNOR U13666 ( .A(n13174), .B(n13173), .Z(n13175) );
  XNOR U13667 ( .A(n13176), .B(n13175), .Z(n13188) );
  XOR U13668 ( .A(n13187), .B(n13188), .Z(n13016) );
  XOR U13669 ( .A(b[13]), .B(n27773), .Z(n13037) );
  OR U13670 ( .A(n13037), .B(n31550), .Z(n12781) );
  NANDN U13671 ( .A(n12779), .B(n31874), .Z(n12780) );
  NAND U13672 ( .A(n12781), .B(n12780), .Z(n13155) );
  NAND U13673 ( .A(n34848), .B(n12782), .Z(n12784) );
  XOR U13674 ( .A(n35375), .B(n23149), .Z(n13040) );
  NAND U13675 ( .A(n34618), .B(n13040), .Z(n12783) );
  NAND U13676 ( .A(n12784), .B(n12783), .Z(n13152) );
  NAND U13677 ( .A(n35188), .B(n12785), .Z(n12787) );
  XOR U13678 ( .A(n35540), .B(n22579), .Z(n13043) );
  NANDN U13679 ( .A(n34968), .B(n13043), .Z(n12786) );
  AND U13680 ( .A(n12787), .B(n12786), .Z(n13153) );
  XNOR U13681 ( .A(n13152), .B(n13153), .Z(n13154) );
  XNOR U13682 ( .A(n13155), .B(n13154), .Z(n13010) );
  XOR U13683 ( .A(b[37]), .B(n20352), .Z(n13028) );
  NANDN U13684 ( .A(n13028), .B(n36311), .Z(n12790) );
  NANDN U13685 ( .A(n12788), .B(n36309), .Z(n12789) );
  NAND U13686 ( .A(n12790), .B(n12789), .Z(n13082) );
  XNOR U13687 ( .A(b[5]), .B(a[69]), .Z(n13031) );
  OR U13688 ( .A(n13031), .B(n29363), .Z(n12793) );
  NANDN U13689 ( .A(n12791), .B(n29864), .Z(n12792) );
  NAND U13690 ( .A(n12793), .B(n12792), .Z(n13079) );
  XOR U13691 ( .A(n30543), .B(n967), .Z(n13034) );
  NAND U13692 ( .A(n13034), .B(n28939), .Z(n12796) );
  NAND U13693 ( .A(n28938), .B(n12794), .Z(n12795) );
  AND U13694 ( .A(n12796), .B(n12795), .Z(n13080) );
  XNOR U13695 ( .A(n13079), .B(n13080), .Z(n13081) );
  XOR U13696 ( .A(n13082), .B(n13081), .Z(n13011) );
  XOR U13697 ( .A(n13010), .B(n13011), .Z(n13013) );
  NANDN U13698 ( .A(n12798), .B(n12797), .Z(n12802) );
  NAND U13699 ( .A(n12800), .B(n12799), .Z(n12801) );
  NAND U13700 ( .A(n12802), .B(n12801), .Z(n13012) );
  XOR U13701 ( .A(n13013), .B(n13012), .Z(n13017) );
  XNOR U13702 ( .A(n13016), .B(n13017), .Z(n13018) );
  XOR U13703 ( .A(n13019), .B(n13018), .Z(n13217) );
  NANDN U13704 ( .A(n12804), .B(n12803), .Z(n12808) );
  NANDN U13705 ( .A(n12806), .B(n12805), .Z(n12807) );
  NAND U13706 ( .A(n12808), .B(n12807), .Z(n13216) );
  NANDN U13707 ( .A(n12810), .B(n12809), .Z(n12814) );
  NAND U13708 ( .A(n12812), .B(n12811), .Z(n12813) );
  NAND U13709 ( .A(n12814), .B(n12813), .Z(n13007) );
  XNOR U13710 ( .A(b[41]), .B(a[33]), .Z(n13091) );
  OR U13711 ( .A(n13091), .B(n36905), .Z(n12817) );
  NANDN U13712 ( .A(n12815), .B(n36807), .Z(n12816) );
  NAND U13713 ( .A(n12817), .B(n12816), .Z(n13113) );
  XOR U13714 ( .A(b[57]), .B(n14514), .Z(n13094) );
  OR U13715 ( .A(n13094), .B(n965), .Z(n12820) );
  NANDN U13716 ( .A(n12818), .B(n38194), .Z(n12819) );
  NAND U13717 ( .A(n12820), .B(n12819), .Z(n13110) );
  NAND U13718 ( .A(n38326), .B(n12821), .Z(n12823) );
  XOR U13719 ( .A(n38400), .B(n13976), .Z(n13097) );
  NANDN U13720 ( .A(n38273), .B(n13097), .Z(n12822) );
  AND U13721 ( .A(n12823), .B(n12822), .Z(n13111) );
  XNOR U13722 ( .A(n13110), .B(n13111), .Z(n13112) );
  XOR U13723 ( .A(n13113), .B(n13112), .Z(n13122) );
  XOR U13724 ( .A(b[33]), .B(n21441), .Z(n13100) );
  NANDN U13725 ( .A(n13100), .B(n35620), .Z(n12826) );
  NANDN U13726 ( .A(n12824), .B(n35621), .Z(n12825) );
  NAND U13727 ( .A(n12826), .B(n12825), .Z(n13131) );
  NANDN U13728 ( .A(n966), .B(a[73]), .Z(n12827) );
  XOR U13729 ( .A(n29232), .B(n12827), .Z(n12829) );
  IV U13730 ( .A(a[72]), .Z(n30210) );
  NANDN U13731 ( .A(n30210), .B(n966), .Z(n12828) );
  AND U13732 ( .A(n12829), .B(n12828), .Z(n13128) );
  XOR U13733 ( .A(b[63]), .B(n12830), .Z(n13107) );
  NANDN U13734 ( .A(n13107), .B(n38422), .Z(n12833) );
  NANDN U13735 ( .A(n12831), .B(n38423), .Z(n12832) );
  AND U13736 ( .A(n12833), .B(n12832), .Z(n13129) );
  XNOR U13737 ( .A(n13128), .B(n13129), .Z(n13130) );
  XOR U13738 ( .A(n13131), .B(n13130), .Z(n13123) );
  XNOR U13739 ( .A(n13122), .B(n13123), .Z(n13125) );
  NANDN U13740 ( .A(n12835), .B(n12834), .Z(n12839) );
  NAND U13741 ( .A(n12837), .B(n12836), .Z(n12838) );
  NAND U13742 ( .A(n12839), .B(n12838), .Z(n13124) );
  XOR U13743 ( .A(n13125), .B(n13124), .Z(n13004) );
  NANDN U13744 ( .A(n12841), .B(n12840), .Z(n12845) );
  NAND U13745 ( .A(n12843), .B(n12842), .Z(n12844) );
  AND U13746 ( .A(n12845), .B(n12844), .Z(n13005) );
  XOR U13747 ( .A(n13004), .B(n13005), .Z(n13006) );
  XNOR U13748 ( .A(n13007), .B(n13006), .Z(n13215) );
  XNOR U13749 ( .A(n13216), .B(n13215), .Z(n13218) );
  XNOR U13750 ( .A(n13217), .B(n13218), .Z(n13223) );
  XOR U13751 ( .A(n13224), .B(n13223), .Z(n13249) );
  NAND U13752 ( .A(n12847), .B(n12846), .Z(n12851) );
  NANDN U13753 ( .A(n12849), .B(n12848), .Z(n12850) );
  NAND U13754 ( .A(n12851), .B(n12850), .Z(n13230) );
  XNOR U13755 ( .A(b[11]), .B(a[63]), .Z(n13191) );
  OR U13756 ( .A(n13191), .B(n31369), .Z(n12854) );
  NANDN U13757 ( .A(n12852), .B(n31119), .Z(n12853) );
  NAND U13758 ( .A(n12854), .B(n12853), .Z(n13212) );
  XOR U13759 ( .A(b[43]), .B(n18639), .Z(n13194) );
  NANDN U13760 ( .A(n13194), .B(n37068), .Z(n12857) );
  NANDN U13761 ( .A(n12855), .B(n37069), .Z(n12856) );
  NAND U13762 ( .A(n12857), .B(n12856), .Z(n13209) );
  XNOR U13763 ( .A(b[45]), .B(a[29]), .Z(n13197) );
  NANDN U13764 ( .A(n13197), .B(n37261), .Z(n12860) );
  NANDN U13765 ( .A(n12858), .B(n37262), .Z(n12859) );
  AND U13766 ( .A(n12860), .B(n12859), .Z(n13210) );
  XNOR U13767 ( .A(n13209), .B(n13210), .Z(n13211) );
  XNOR U13768 ( .A(n13212), .B(n13211), .Z(n13022) );
  XOR U13769 ( .A(n979), .B(n16916), .Z(n13200) );
  NANDN U13770 ( .A(n37756), .B(n13200), .Z(n12863) );
  NANDN U13771 ( .A(n12861), .B(n37652), .Z(n12862) );
  NAND U13772 ( .A(n12863), .B(n12862), .Z(n13182) );
  NAND U13773 ( .A(n37469), .B(n12864), .Z(n12866) );
  XOR U13774 ( .A(b[47]), .B(n17960), .Z(n13203) );
  NANDN U13775 ( .A(n13203), .B(n37471), .Z(n12865) );
  NAND U13776 ( .A(n12866), .B(n12865), .Z(n13179) );
  XOR U13777 ( .A(n969), .B(n28403), .Z(n13206) );
  NAND U13778 ( .A(n30509), .B(n13206), .Z(n12869) );
  NANDN U13779 ( .A(n12867), .B(n30846), .Z(n12868) );
  AND U13780 ( .A(n12869), .B(n12868), .Z(n13180) );
  XNOR U13781 ( .A(n13179), .B(n13180), .Z(n13181) );
  XOR U13782 ( .A(n13182), .B(n13181), .Z(n13023) );
  XNOR U13783 ( .A(n13022), .B(n13023), .Z(n13024) );
  NANDN U13784 ( .A(n12871), .B(n12870), .Z(n12875) );
  NAND U13785 ( .A(n12873), .B(n12872), .Z(n12874) );
  AND U13786 ( .A(n12875), .B(n12874), .Z(n13025) );
  XNOR U13787 ( .A(n13024), .B(n13025), .Z(n13244) );
  XNOR U13788 ( .A(n13244), .B(n13243), .Z(n13245) );
  XNOR U13789 ( .A(b[35]), .B(a[39]), .Z(n13164) );
  NANDN U13790 ( .A(n13164), .B(n35985), .Z(n12882) );
  NANDN U13791 ( .A(n12880), .B(n35986), .Z(n12881) );
  NAND U13792 ( .A(n12882), .B(n12881), .Z(n13161) );
  XOR U13793 ( .A(n31123), .B(n29372), .Z(n13167) );
  NAND U13794 ( .A(n13167), .B(n29949), .Z(n12885) );
  NAND U13795 ( .A(n29948), .B(n12883), .Z(n12884) );
  NAND U13796 ( .A(n12885), .B(n12884), .Z(n13158) );
  XOR U13797 ( .A(b[55]), .B(n15113), .Z(n13170) );
  NANDN U13798 ( .A(n13170), .B(n38075), .Z(n12888) );
  NANDN U13799 ( .A(n12886), .B(n38073), .Z(n12887) );
  AND U13800 ( .A(n12888), .B(n12887), .Z(n13159) );
  XNOR U13801 ( .A(n13158), .B(n13159), .Z(n13160) );
  XNOR U13802 ( .A(n13161), .B(n13160), .Z(n13001) );
  NANDN U13803 ( .A(n12890), .B(n12889), .Z(n12894) );
  NAND U13804 ( .A(n12892), .B(n12891), .Z(n12893) );
  NAND U13805 ( .A(n12894), .B(n12893), .Z(n12998) );
  OR U13806 ( .A(n12896), .B(n12895), .Z(n12900) );
  NANDN U13807 ( .A(n12898), .B(n12897), .Z(n12899) );
  NAND U13808 ( .A(n12900), .B(n12899), .Z(n12999) );
  XNOR U13809 ( .A(n12998), .B(n12999), .Z(n13000) );
  XOR U13810 ( .A(n13001), .B(n13000), .Z(n13246) );
  XNOR U13811 ( .A(n13245), .B(n13246), .Z(n13228) );
  NANDN U13812 ( .A(n12902), .B(n12901), .Z(n12906) );
  NANDN U13813 ( .A(n12904), .B(n12903), .Z(n12905) );
  NAND U13814 ( .A(n12906), .B(n12905), .Z(n13237) );
  NANDN U13815 ( .A(n12908), .B(n12907), .Z(n12912) );
  NAND U13816 ( .A(n12910), .B(n12909), .Z(n12911) );
  NAND U13817 ( .A(n12912), .B(n12911), .Z(n13238) );
  XNOR U13818 ( .A(n13237), .B(n13238), .Z(n13239) );
  XNOR U13819 ( .A(b[15]), .B(a[59]), .Z(n13134) );
  OR U13820 ( .A(n13134), .B(n32010), .Z(n12919) );
  NANDN U13821 ( .A(n12917), .B(n32011), .Z(n12918) );
  NAND U13822 ( .A(n12919), .B(n12918), .Z(n13055) );
  XNOR U13823 ( .A(b[25]), .B(n23852), .Z(n13137) );
  NANDN U13824 ( .A(n34219), .B(n13137), .Z(n12922) );
  NAND U13825 ( .A(n34217), .B(n12920), .Z(n12921) );
  NAND U13826 ( .A(n12922), .B(n12921), .Z(n13052) );
  XNOR U13827 ( .A(b[17]), .B(a[57]), .Z(n13140) );
  NANDN U13828 ( .A(n13140), .B(n32543), .Z(n12925) );
  NANDN U13829 ( .A(n12923), .B(n32541), .Z(n12924) );
  AND U13830 ( .A(n12925), .B(n12924), .Z(n13053) );
  XNOR U13831 ( .A(n13052), .B(n13053), .Z(n13054) );
  XNOR U13832 ( .A(n13055), .B(n13054), .Z(n13073) );
  XOR U13833 ( .A(b[39]), .B(n20315), .Z(n13143) );
  NANDN U13834 ( .A(n13143), .B(n36553), .Z(n12928) );
  NANDN U13835 ( .A(n12926), .B(n36643), .Z(n12927) );
  NAND U13836 ( .A(n12928), .B(n12927), .Z(n13049) );
  XOR U13837 ( .A(b[51]), .B(n16269), .Z(n13146) );
  NANDN U13838 ( .A(n13146), .B(n37803), .Z(n12931) );
  NANDN U13839 ( .A(n12929), .B(n37802), .Z(n12930) );
  NAND U13840 ( .A(n12931), .B(n12930), .Z(n13046) );
  XOR U13841 ( .A(b[53]), .B(n16220), .Z(n13149) );
  NANDN U13842 ( .A(n13149), .B(n37940), .Z(n12934) );
  NANDN U13843 ( .A(n12932), .B(n37941), .Z(n12933) );
  AND U13844 ( .A(n12934), .B(n12933), .Z(n13047) );
  XNOR U13845 ( .A(n13046), .B(n13047), .Z(n13048) );
  XOR U13846 ( .A(n13049), .B(n13048), .Z(n13074) );
  XNOR U13847 ( .A(n13073), .B(n13074), .Z(n13075) );
  NANDN U13848 ( .A(n12936), .B(n12935), .Z(n12940) );
  NAND U13849 ( .A(n12938), .B(n12937), .Z(n12939) );
  AND U13850 ( .A(n12940), .B(n12939), .Z(n13076) );
  XNOR U13851 ( .A(n13075), .B(n13076), .Z(n13117) );
  NANDN U13852 ( .A(n12942), .B(n12941), .Z(n12946) );
  NAND U13853 ( .A(n12944), .B(n12943), .Z(n12945) );
  AND U13854 ( .A(n12946), .B(n12945), .Z(n13116) );
  XNOR U13855 ( .A(n13117), .B(n13116), .Z(n13118) );
  XOR U13856 ( .A(n13119), .B(n13118), .Z(n13240) );
  XNOR U13857 ( .A(n13239), .B(n13240), .Z(n13227) );
  XOR U13858 ( .A(n13230), .B(n13229), .Z(n13250) );
  XNOR U13859 ( .A(n13249), .B(n13250), .Z(n13251) );
  NAND U13860 ( .A(n12948), .B(n12947), .Z(n12952) );
  NANDN U13861 ( .A(n12950), .B(n12949), .Z(n12951) );
  NAND U13862 ( .A(n12952), .B(n12951), .Z(n13252) );
  XOR U13863 ( .A(n13251), .B(n13252), .Z(n13264) );
  NAND U13864 ( .A(n12954), .B(n12953), .Z(n12958) );
  NANDN U13865 ( .A(n12956), .B(n12955), .Z(n12957) );
  NAND U13866 ( .A(n12958), .B(n12957), .Z(n13258) );
  XNOR U13867 ( .A(n13256), .B(n13255), .Z(n13257) );
  XNOR U13868 ( .A(n13258), .B(n13257), .Z(n13261) );
  NANDN U13869 ( .A(n12968), .B(n12967), .Z(n12972) );
  NANDN U13870 ( .A(n12970), .B(n12969), .Z(n12971) );
  NAND U13871 ( .A(n12972), .B(n12971), .Z(n13262) );
  XNOR U13872 ( .A(n13264), .B(n13263), .Z(n13270) );
  XOR U13873 ( .A(n13269), .B(n13270), .Z(n13276) );
  OR U13874 ( .A(n12974), .B(n12973), .Z(n12978) );
  NAND U13875 ( .A(n12976), .B(n12975), .Z(n12977) );
  NAND U13876 ( .A(n12978), .B(n12977), .Z(n13274) );
  NANDN U13877 ( .A(n12980), .B(n12979), .Z(n12984) );
  NANDN U13878 ( .A(n12982), .B(n12981), .Z(n12983) );
  AND U13879 ( .A(n12984), .B(n12983), .Z(n13273) );
  XNOR U13880 ( .A(n13274), .B(n13273), .Z(n13275) );
  XNOR U13881 ( .A(n13276), .B(n13275), .Z(n12994) );
  XNOR U13882 ( .A(n12994), .B(n12995), .Z(n12996) );
  XNOR U13883 ( .A(n12997), .B(n12996), .Z(n13279) );
  XNOR U13884 ( .A(n13279), .B(sreg[137]), .Z(n13281) );
  NAND U13885 ( .A(n12989), .B(sreg[136]), .Z(n12993) );
  OR U13886 ( .A(n12991), .B(n12990), .Z(n12992) );
  AND U13887 ( .A(n12993), .B(n12992), .Z(n13280) );
  XOR U13888 ( .A(n13281), .B(n13280), .Z(c[137]) );
  NANDN U13889 ( .A(n12999), .B(n12998), .Z(n13003) );
  NAND U13890 ( .A(n13001), .B(n13000), .Z(n13002) );
  NAND U13891 ( .A(n13003), .B(n13002), .Z(n13534) );
  NAND U13892 ( .A(n13005), .B(n13004), .Z(n13009) );
  NANDN U13893 ( .A(n13007), .B(n13006), .Z(n13008) );
  AND U13894 ( .A(n13009), .B(n13008), .Z(n13531) );
  NANDN U13895 ( .A(n13011), .B(n13010), .Z(n13015) );
  OR U13896 ( .A(n13013), .B(n13012), .Z(n13014) );
  AND U13897 ( .A(n13015), .B(n13014), .Z(n13532) );
  XNOR U13898 ( .A(n13534), .B(n13533), .Z(n13301) );
  NANDN U13899 ( .A(n13017), .B(n13016), .Z(n13021) );
  NANDN U13900 ( .A(n13019), .B(n13018), .Z(n13020) );
  AND U13901 ( .A(n13021), .B(n13020), .Z(n13300) );
  XNOR U13902 ( .A(n13301), .B(n13300), .Z(n13302) );
  NANDN U13903 ( .A(n13023), .B(n13022), .Z(n13027) );
  NAND U13904 ( .A(n13025), .B(n13024), .Z(n13026) );
  NAND U13905 ( .A(n13027), .B(n13026), .Z(n13427) );
  XOR U13906 ( .A(b[37]), .B(n20686), .Z(n13452) );
  NANDN U13907 ( .A(n13452), .B(n36311), .Z(n13030) );
  NANDN U13908 ( .A(n13028), .B(n36309), .Z(n13029) );
  NAND U13909 ( .A(n13030), .B(n13029), .Z(n13491) );
  XOR U13910 ( .A(a[70]), .B(n968), .Z(n13455) );
  OR U13911 ( .A(n13455), .B(n29363), .Z(n13033) );
  NANDN U13912 ( .A(n13031), .B(n29864), .Z(n13032) );
  NAND U13913 ( .A(n13033), .B(n13032), .Z(n13488) );
  XOR U13914 ( .A(n30210), .B(n967), .Z(n13458) );
  NAND U13915 ( .A(n13458), .B(n28939), .Z(n13036) );
  NAND U13916 ( .A(n28938), .B(n13034), .Z(n13035) );
  AND U13917 ( .A(n13036), .B(n13035), .Z(n13489) );
  XNOR U13918 ( .A(n13488), .B(n13489), .Z(n13490) );
  XNOR U13919 ( .A(n13491), .B(n13490), .Z(n13422) );
  XNOR U13920 ( .A(b[13]), .B(a[62]), .Z(n13461) );
  OR U13921 ( .A(n13461), .B(n31550), .Z(n13039) );
  NANDN U13922 ( .A(n13037), .B(n31874), .Z(n13038) );
  NAND U13923 ( .A(n13039), .B(n13038), .Z(n13333) );
  NAND U13924 ( .A(n34848), .B(n13040), .Z(n13042) );
  XOR U13925 ( .A(n35375), .B(n23447), .Z(n13464) );
  NAND U13926 ( .A(n34618), .B(n13464), .Z(n13041) );
  NAND U13927 ( .A(n13042), .B(n13041), .Z(n13330) );
  NAND U13928 ( .A(n35188), .B(n13043), .Z(n13045) );
  XOR U13929 ( .A(n35540), .B(n22964), .Z(n13467) );
  NANDN U13930 ( .A(n34968), .B(n13467), .Z(n13044) );
  AND U13931 ( .A(n13045), .B(n13044), .Z(n13331) );
  XNOR U13932 ( .A(n13330), .B(n13331), .Z(n13332) );
  XNOR U13933 ( .A(n13333), .B(n13332), .Z(n13419) );
  NANDN U13934 ( .A(n13047), .B(n13046), .Z(n13051) );
  NAND U13935 ( .A(n13049), .B(n13048), .Z(n13050) );
  NAND U13936 ( .A(n13051), .B(n13050), .Z(n13420) );
  XNOR U13937 ( .A(n13419), .B(n13420), .Z(n13421) );
  XOR U13938 ( .A(n13422), .B(n13421), .Z(n13426) );
  NANDN U13939 ( .A(n13053), .B(n13052), .Z(n13057) );
  NAND U13940 ( .A(n13055), .B(n13054), .Z(n13056) );
  NAND U13941 ( .A(n13057), .B(n13056), .Z(n13378) );
  NAND U13942 ( .A(a[10]), .B(b[63]), .Z(n13392) );
  NANDN U13943 ( .A(n13058), .B(n38369), .Z(n13060) );
  XOR U13944 ( .A(b[61]), .B(n14210), .Z(n13446) );
  OR U13945 ( .A(n13446), .B(n38371), .Z(n13059) );
  NAND U13946 ( .A(n13060), .B(n13059), .Z(n13390) );
  NANDN U13947 ( .A(n13061), .B(n35311), .Z(n13063) );
  XOR U13948 ( .A(b[31]), .B(n22289), .Z(n13449) );
  NANDN U13949 ( .A(n13449), .B(n35313), .Z(n13062) );
  AND U13950 ( .A(n13063), .B(n13062), .Z(n13389) );
  XNOR U13951 ( .A(n13390), .B(n13389), .Z(n13391) );
  XOR U13952 ( .A(n13392), .B(n13391), .Z(n13376) );
  NAND U13953 ( .A(n33283), .B(n13064), .Z(n13066) );
  XOR U13954 ( .A(n33020), .B(n25860), .Z(n13431) );
  NANDN U13955 ( .A(n33021), .B(n13431), .Z(n13065) );
  NAND U13956 ( .A(n13066), .B(n13065), .Z(n13516) );
  XNOR U13957 ( .A(b[21]), .B(a[54]), .Z(n13434) );
  OR U13958 ( .A(n13434), .B(n33634), .Z(n13069) );
  NANDN U13959 ( .A(n13067), .B(n33464), .Z(n13068) );
  NAND U13960 ( .A(n13069), .B(n13068), .Z(n13513) );
  NAND U13961 ( .A(n34044), .B(n13070), .Z(n13072) );
  XOR U13962 ( .A(n34510), .B(n25134), .Z(n13437) );
  NANDN U13963 ( .A(n33867), .B(n13437), .Z(n13071) );
  AND U13964 ( .A(n13072), .B(n13071), .Z(n13514) );
  XNOR U13965 ( .A(n13513), .B(n13514), .Z(n13515) );
  XNOR U13966 ( .A(n13516), .B(n13515), .Z(n13377) );
  XNOR U13967 ( .A(n13376), .B(n13377), .Z(n13379) );
  XNOR U13968 ( .A(n13378), .B(n13379), .Z(n13425) );
  XOR U13969 ( .A(n13426), .B(n13425), .Z(n13428) );
  XNOR U13970 ( .A(n13427), .B(n13428), .Z(n13403) );
  NANDN U13971 ( .A(n13074), .B(n13073), .Z(n13078) );
  NAND U13972 ( .A(n13076), .B(n13075), .Z(n13077) );
  NAND U13973 ( .A(n13078), .B(n13077), .Z(n13402) );
  NANDN U13974 ( .A(n13080), .B(n13079), .Z(n13084) );
  NAND U13975 ( .A(n13082), .B(n13081), .Z(n13083) );
  NAND U13976 ( .A(n13084), .B(n13083), .Z(n13416) );
  NANDN U13977 ( .A(n13086), .B(n13085), .Z(n13090) );
  NAND U13978 ( .A(n13088), .B(n13087), .Z(n13089) );
  NAND U13979 ( .A(n13090), .B(n13089), .Z(n13349) );
  XNOR U13980 ( .A(b[41]), .B(a[34]), .Z(n13494) );
  OR U13981 ( .A(n13494), .B(n36905), .Z(n13093) );
  NANDN U13982 ( .A(n13091), .B(n36807), .Z(n13092) );
  NAND U13983 ( .A(n13093), .B(n13092), .Z(n13522) );
  XOR U13984 ( .A(b[57]), .B(n14905), .Z(n13497) );
  OR U13985 ( .A(n13497), .B(n965), .Z(n13096) );
  NANDN U13986 ( .A(n13094), .B(n38194), .Z(n13095) );
  NAND U13987 ( .A(n13096), .B(n13095), .Z(n13519) );
  NAND U13988 ( .A(n38326), .B(n13097), .Z(n13099) );
  XOR U13989 ( .A(n38400), .B(n14259), .Z(n13500) );
  NANDN U13990 ( .A(n38273), .B(n13500), .Z(n13098) );
  AND U13991 ( .A(n13099), .B(n13098), .Z(n13520) );
  XNOR U13992 ( .A(n13519), .B(n13520), .Z(n13521) );
  XOR U13993 ( .A(n13522), .B(n13521), .Z(n13347) );
  XOR U13994 ( .A(b[33]), .B(n22246), .Z(n13503) );
  NANDN U13995 ( .A(n13503), .B(n35620), .Z(n13102) );
  NANDN U13996 ( .A(n13100), .B(n35621), .Z(n13101) );
  NAND U13997 ( .A(n13102), .B(n13101), .Z(n13345) );
  NANDN U13998 ( .A(n966), .B(a[74]), .Z(n13103) );
  XOR U13999 ( .A(n29232), .B(n13103), .Z(n13105) );
  NANDN U14000 ( .A(b[0]), .B(a[73]), .Z(n13104) );
  AND U14001 ( .A(n13105), .B(n13104), .Z(n13342) );
  XOR U14002 ( .A(b[63]), .B(n13106), .Z(n13510) );
  NANDN U14003 ( .A(n13510), .B(n38422), .Z(n13109) );
  NANDN U14004 ( .A(n13107), .B(n38423), .Z(n13108) );
  AND U14005 ( .A(n13109), .B(n13108), .Z(n13343) );
  XNOR U14006 ( .A(n13342), .B(n13343), .Z(n13344) );
  XNOR U14007 ( .A(n13345), .B(n13344), .Z(n13346) );
  XNOR U14008 ( .A(n13347), .B(n13346), .Z(n13348) );
  XOR U14009 ( .A(n13349), .B(n13348), .Z(n13414) );
  NANDN U14010 ( .A(n13111), .B(n13110), .Z(n13115) );
  NAND U14011 ( .A(n13113), .B(n13112), .Z(n13114) );
  AND U14012 ( .A(n13115), .B(n13114), .Z(n13413) );
  XNOR U14013 ( .A(n13414), .B(n13413), .Z(n13415) );
  XNOR U14014 ( .A(n13416), .B(n13415), .Z(n13401) );
  XNOR U14015 ( .A(n13402), .B(n13401), .Z(n13404) );
  XNOR U14016 ( .A(n13403), .B(n13404), .Z(n13303) );
  XNOR U14017 ( .A(n13302), .B(n13303), .Z(n13296) );
  NANDN U14018 ( .A(n13117), .B(n13116), .Z(n13121) );
  NANDN U14019 ( .A(n13119), .B(n13118), .Z(n13120) );
  NAND U14020 ( .A(n13121), .B(n13120), .Z(n13537) );
  OR U14021 ( .A(n13123), .B(n13122), .Z(n13127) );
  OR U14022 ( .A(n13125), .B(n13124), .Z(n13126) );
  AND U14023 ( .A(n13127), .B(n13126), .Z(n13538) );
  XNOR U14024 ( .A(n13537), .B(n13538), .Z(n13539) );
  NANDN U14025 ( .A(n13129), .B(n13128), .Z(n13133) );
  NAND U14026 ( .A(n13131), .B(n13130), .Z(n13132) );
  NAND U14027 ( .A(n13133), .B(n13132), .Z(n13309) );
  XOR U14028 ( .A(b[15]), .B(n27436), .Z(n13312) );
  OR U14029 ( .A(n13312), .B(n32010), .Z(n13136) );
  NANDN U14030 ( .A(n13134), .B(n32011), .Z(n13135) );
  NAND U14031 ( .A(n13136), .B(n13135), .Z(n13443) );
  XNOR U14032 ( .A(b[25]), .B(n24671), .Z(n13315) );
  NANDN U14033 ( .A(n34219), .B(n13315), .Z(n13139) );
  NAND U14034 ( .A(n34217), .B(n13137), .Z(n13138) );
  NAND U14035 ( .A(n13139), .B(n13138), .Z(n13440) );
  XNOR U14036 ( .A(b[17]), .B(a[58]), .Z(n13318) );
  NANDN U14037 ( .A(n13318), .B(n32543), .Z(n13142) );
  NANDN U14038 ( .A(n13140), .B(n32541), .Z(n13141) );
  AND U14039 ( .A(n13142), .B(n13141), .Z(n13441) );
  XNOR U14040 ( .A(n13440), .B(n13441), .Z(n13442) );
  XNOR U14041 ( .A(n13443), .B(n13442), .Z(n13482) );
  XOR U14042 ( .A(b[39]), .B(n19980), .Z(n13321) );
  NANDN U14043 ( .A(n13321), .B(n36553), .Z(n13145) );
  NANDN U14044 ( .A(n13143), .B(n36643), .Z(n13144) );
  NAND U14045 ( .A(n13145), .B(n13144), .Z(n13473) );
  XOR U14046 ( .A(b[51]), .B(n16508), .Z(n13324) );
  NANDN U14047 ( .A(n13324), .B(n37803), .Z(n13148) );
  NANDN U14048 ( .A(n13146), .B(n37802), .Z(n13147) );
  NAND U14049 ( .A(n13148), .B(n13147), .Z(n13470) );
  XOR U14050 ( .A(b[53]), .B(n15963), .Z(n13327) );
  NANDN U14051 ( .A(n13327), .B(n37940), .Z(n13151) );
  NANDN U14052 ( .A(n13149), .B(n37941), .Z(n13150) );
  AND U14053 ( .A(n13151), .B(n13150), .Z(n13471) );
  XNOR U14054 ( .A(n13470), .B(n13471), .Z(n13472) );
  XOR U14055 ( .A(n13473), .B(n13472), .Z(n13483) );
  XNOR U14056 ( .A(n13482), .B(n13483), .Z(n13484) );
  NANDN U14057 ( .A(n13153), .B(n13152), .Z(n13157) );
  NAND U14058 ( .A(n13155), .B(n13154), .Z(n13156) );
  AND U14059 ( .A(n13157), .B(n13156), .Z(n13485) );
  XNOR U14060 ( .A(n13484), .B(n13485), .Z(n13307) );
  NANDN U14061 ( .A(n13159), .B(n13158), .Z(n13163) );
  NAND U14062 ( .A(n13161), .B(n13160), .Z(n13162) );
  AND U14063 ( .A(n13163), .B(n13162), .Z(n13306) );
  XNOR U14064 ( .A(n13307), .B(n13306), .Z(n13308) );
  XOR U14065 ( .A(n13309), .B(n13308), .Z(n13540) );
  XNOR U14066 ( .A(n13539), .B(n13540), .Z(n13543) );
  XNOR U14067 ( .A(b[35]), .B(a[40]), .Z(n13380) );
  NANDN U14068 ( .A(n13380), .B(n35985), .Z(n13166) );
  NANDN U14069 ( .A(n13164), .B(n35986), .Z(n13165) );
  NAND U14070 ( .A(n13166), .B(n13165), .Z(n13339) );
  XOR U14071 ( .A(n31123), .B(n29868), .Z(n13383) );
  NAND U14072 ( .A(n13383), .B(n29949), .Z(n13169) );
  NAND U14073 ( .A(n29948), .B(n13167), .Z(n13168) );
  NAND U14074 ( .A(n13169), .B(n13168), .Z(n13336) );
  XOR U14075 ( .A(b[55]), .B(n15484), .Z(n13386) );
  NANDN U14076 ( .A(n13386), .B(n38075), .Z(n13172) );
  NANDN U14077 ( .A(n13170), .B(n38073), .Z(n13171) );
  AND U14078 ( .A(n13172), .B(n13171), .Z(n13337) );
  XNOR U14079 ( .A(n13336), .B(n13337), .Z(n13338) );
  XNOR U14080 ( .A(n13339), .B(n13338), .Z(n13410) );
  NANDN U14081 ( .A(n13174), .B(n13173), .Z(n13178) );
  NAND U14082 ( .A(n13176), .B(n13175), .Z(n13177) );
  NAND U14083 ( .A(n13178), .B(n13177), .Z(n13407) );
  NANDN U14084 ( .A(n13180), .B(n13179), .Z(n13184) );
  NAND U14085 ( .A(n13182), .B(n13181), .Z(n13183) );
  NAND U14086 ( .A(n13184), .B(n13183), .Z(n13408) );
  XNOR U14087 ( .A(n13407), .B(n13408), .Z(n13409) );
  XOR U14088 ( .A(n13410), .B(n13409), .Z(n13527) );
  NANDN U14089 ( .A(n13186), .B(n13185), .Z(n13190) );
  NANDN U14090 ( .A(n13188), .B(n13187), .Z(n13189) );
  NAND U14091 ( .A(n13190), .B(n13189), .Z(n13525) );
  XNOR U14092 ( .A(b[11]), .B(a[64]), .Z(n13352) );
  OR U14093 ( .A(n13352), .B(n31369), .Z(n13193) );
  NANDN U14094 ( .A(n13191), .B(n31119), .Z(n13192) );
  NAND U14095 ( .A(n13193), .B(n13192), .Z(n13373) );
  XOR U14096 ( .A(b[43]), .B(n18841), .Z(n13355) );
  NANDN U14097 ( .A(n13355), .B(n37068), .Z(n13196) );
  NANDN U14098 ( .A(n13194), .B(n37069), .Z(n13195) );
  NAND U14099 ( .A(n13196), .B(n13195), .Z(n13370) );
  XNOR U14100 ( .A(b[45]), .B(a[30]), .Z(n13358) );
  NANDN U14101 ( .A(n13358), .B(n37261), .Z(n13199) );
  NANDN U14102 ( .A(n13197), .B(n37262), .Z(n13198) );
  AND U14103 ( .A(n13199), .B(n13198), .Z(n13371) );
  XNOR U14104 ( .A(n13370), .B(n13371), .Z(n13372) );
  XNOR U14105 ( .A(n13373), .B(n13372), .Z(n13476) );
  NAND U14106 ( .A(n37652), .B(n13200), .Z(n13202) );
  XOR U14107 ( .A(n979), .B(a[26]), .Z(n13361) );
  OR U14108 ( .A(n13361), .B(n37756), .Z(n13201) );
  NAND U14109 ( .A(n13202), .B(n13201), .Z(n13397) );
  NANDN U14110 ( .A(n13203), .B(n37469), .Z(n13205) );
  XOR U14111 ( .A(b[47]), .B(n17702), .Z(n13364) );
  NANDN U14112 ( .A(n13364), .B(n37471), .Z(n13204) );
  AND U14113 ( .A(n13205), .B(n13204), .Z(n13396) );
  NAND U14114 ( .A(n30846), .B(n13206), .Z(n13208) );
  XOR U14115 ( .A(n969), .B(n28701), .Z(n13367) );
  NAND U14116 ( .A(n30509), .B(n13367), .Z(n13207) );
  NAND U14117 ( .A(n13208), .B(n13207), .Z(n13395) );
  XNOR U14118 ( .A(n13396), .B(n13395), .Z(n13398) );
  XOR U14119 ( .A(n13397), .B(n13398), .Z(n13477) );
  XNOR U14120 ( .A(n13476), .B(n13477), .Z(n13478) );
  NANDN U14121 ( .A(n13210), .B(n13209), .Z(n13214) );
  NAND U14122 ( .A(n13212), .B(n13211), .Z(n13213) );
  AND U14123 ( .A(n13214), .B(n13213), .Z(n13479) );
  XNOR U14124 ( .A(n13478), .B(n13479), .Z(n13526) );
  XNOR U14125 ( .A(n13525), .B(n13526), .Z(n13528) );
  XOR U14126 ( .A(n13527), .B(n13528), .Z(n13544) );
  NAND U14127 ( .A(n13216), .B(n13215), .Z(n13220) );
  NANDN U14128 ( .A(n13218), .B(n13217), .Z(n13219) );
  AND U14129 ( .A(n13220), .B(n13219), .Z(n13546) );
  XNOR U14130 ( .A(n13545), .B(n13546), .Z(n13297) );
  XNOR U14131 ( .A(n13296), .B(n13297), .Z(n13298) );
  NAND U14132 ( .A(n13222), .B(n13221), .Z(n13226) );
  NANDN U14133 ( .A(n13224), .B(n13223), .Z(n13225) );
  AND U14134 ( .A(n13226), .B(n13225), .Z(n13299) );
  XNOR U14135 ( .A(n13298), .B(n13299), .Z(n13551) );
  NANDN U14136 ( .A(n13228), .B(n13227), .Z(n13232) );
  NAND U14137 ( .A(n13230), .B(n13229), .Z(n13231) );
  AND U14138 ( .A(n13232), .B(n13231), .Z(n13550) );
  NANDN U14139 ( .A(n13238), .B(n13237), .Z(n13242) );
  NANDN U14140 ( .A(n13240), .B(n13239), .Z(n13241) );
  NAND U14141 ( .A(n13242), .B(n13241), .Z(n13290) );
  NANDN U14142 ( .A(n13244), .B(n13243), .Z(n13248) );
  NAND U14143 ( .A(n13246), .B(n13245), .Z(n13247) );
  AND U14144 ( .A(n13248), .B(n13247), .Z(n13291) );
  XNOR U14145 ( .A(n13290), .B(n13291), .Z(n13292) );
  XOR U14146 ( .A(n13293), .B(n13292), .Z(n13549) );
  NANDN U14147 ( .A(n13250), .B(n13249), .Z(n13254) );
  NANDN U14148 ( .A(n13252), .B(n13251), .Z(n13253) );
  NAND U14149 ( .A(n13254), .B(n13253), .Z(n13553) );
  NANDN U14150 ( .A(n13256), .B(n13255), .Z(n13260) );
  NANDN U14151 ( .A(n13258), .B(n13257), .Z(n13259) );
  AND U14152 ( .A(n13260), .B(n13259), .Z(n13552) );
  XNOR U14153 ( .A(n13553), .B(n13552), .Z(n13554) );
  XOR U14154 ( .A(n13555), .B(n13554), .Z(n13561) );
  OR U14155 ( .A(n13262), .B(n13261), .Z(n13266) );
  NAND U14156 ( .A(n13264), .B(n13263), .Z(n13265) );
  NAND U14157 ( .A(n13266), .B(n13265), .Z(n13559) );
  NANDN U14158 ( .A(n13268), .B(n13267), .Z(n13272) );
  NANDN U14159 ( .A(n13270), .B(n13269), .Z(n13271) );
  AND U14160 ( .A(n13272), .B(n13271), .Z(n13558) );
  XNOR U14161 ( .A(n13559), .B(n13558), .Z(n13560) );
  XNOR U14162 ( .A(n13561), .B(n13560), .Z(n13284) );
  NANDN U14163 ( .A(n13274), .B(n13273), .Z(n13278) );
  NAND U14164 ( .A(n13276), .B(n13275), .Z(n13277) );
  NAND U14165 ( .A(n13278), .B(n13277), .Z(n13285) );
  XOR U14166 ( .A(n13284), .B(n13285), .Z(n13286) );
  XNOR U14167 ( .A(n13287), .B(n13286), .Z(n13564) );
  XNOR U14168 ( .A(n13564), .B(sreg[138]), .Z(n13566) );
  NAND U14169 ( .A(n13279), .B(sreg[137]), .Z(n13283) );
  OR U14170 ( .A(n13281), .B(n13280), .Z(n13282) );
  AND U14171 ( .A(n13283), .B(n13282), .Z(n13565) );
  XOR U14172 ( .A(n13566), .B(n13565), .Z(c[138]) );
  OR U14173 ( .A(n13285), .B(n13284), .Z(n13289) );
  NAND U14174 ( .A(n13287), .B(n13286), .Z(n13288) );
  NAND U14175 ( .A(n13289), .B(n13288), .Z(n13572) );
  NANDN U14176 ( .A(n13291), .B(n13290), .Z(n13295) );
  NAND U14177 ( .A(n13293), .B(n13292), .Z(n13294) );
  NAND U14178 ( .A(n13295), .B(n13294), .Z(n13837) );
  XNOR U14179 ( .A(n13837), .B(n13838), .Z(n13839) );
  NANDN U14180 ( .A(n13301), .B(n13300), .Z(n13305) );
  NAND U14181 ( .A(n13303), .B(n13302), .Z(n13304) );
  NAND U14182 ( .A(n13305), .B(n13304), .Z(n13575) );
  NANDN U14183 ( .A(n13307), .B(n13306), .Z(n13311) );
  NANDN U14184 ( .A(n13309), .B(n13308), .Z(n13310) );
  NAND U14185 ( .A(n13311), .B(n13310), .Z(n13826) );
  XOR U14186 ( .A(b[15]), .B(n27773), .Z(n13600) );
  OR U14187 ( .A(n13600), .B(n32010), .Z(n13314) );
  NANDN U14188 ( .A(n13312), .B(n32011), .Z(n13313) );
  NAND U14189 ( .A(n13314), .B(n13313), .Z(n13739) );
  XNOR U14190 ( .A(b[25]), .B(n24288), .Z(n13603) );
  NANDN U14191 ( .A(n34219), .B(n13603), .Z(n13317) );
  NAND U14192 ( .A(n34217), .B(n13315), .Z(n13316) );
  NAND U14193 ( .A(n13317), .B(n13316), .Z(n13736) );
  XOR U14194 ( .A(b[17]), .B(a[59]), .Z(n13606) );
  NAND U14195 ( .A(n13606), .B(n32543), .Z(n13320) );
  NANDN U14196 ( .A(n13318), .B(n32541), .Z(n13319) );
  AND U14197 ( .A(n13320), .B(n13319), .Z(n13737) );
  XNOR U14198 ( .A(n13736), .B(n13737), .Z(n13738) );
  XNOR U14199 ( .A(n13739), .B(n13738), .Z(n13757) );
  XOR U14200 ( .A(b[39]), .B(n20352), .Z(n13591) );
  NANDN U14201 ( .A(n13591), .B(n36553), .Z(n13323) );
  NANDN U14202 ( .A(n13321), .B(n36643), .Z(n13322) );
  NAND U14203 ( .A(n13323), .B(n13322), .Z(n13733) );
  XOR U14204 ( .A(b[51]), .B(n16916), .Z(n13594) );
  NANDN U14205 ( .A(n13594), .B(n37803), .Z(n13326) );
  NANDN U14206 ( .A(n13324), .B(n37802), .Z(n13325) );
  NAND U14207 ( .A(n13326), .B(n13325), .Z(n13730) );
  XOR U14208 ( .A(b[53]), .B(n16269), .Z(n13597) );
  NANDN U14209 ( .A(n13597), .B(n37940), .Z(n13329) );
  NANDN U14210 ( .A(n13327), .B(n37941), .Z(n13328) );
  AND U14211 ( .A(n13329), .B(n13328), .Z(n13731) );
  XNOR U14212 ( .A(n13730), .B(n13731), .Z(n13732) );
  XOR U14213 ( .A(n13733), .B(n13732), .Z(n13758) );
  XNOR U14214 ( .A(n13757), .B(n13758), .Z(n13759) );
  NANDN U14215 ( .A(n13331), .B(n13330), .Z(n13335) );
  NAND U14216 ( .A(n13333), .B(n13332), .Z(n13334) );
  NAND U14217 ( .A(n13335), .B(n13334), .Z(n13760) );
  XOR U14218 ( .A(n13759), .B(n13760), .Z(n13636) );
  NANDN U14219 ( .A(n13337), .B(n13336), .Z(n13341) );
  NAND U14220 ( .A(n13339), .B(n13338), .Z(n13340) );
  NAND U14221 ( .A(n13341), .B(n13340), .Z(n13633) );
  XNOR U14222 ( .A(n13633), .B(n13634), .Z(n13635) );
  XNOR U14223 ( .A(n13636), .B(n13635), .Z(n13823) );
  NANDN U14224 ( .A(n13347), .B(n13346), .Z(n13351) );
  NANDN U14225 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U14226 ( .A(n13351), .B(n13350), .Z(n13824) );
  XNOR U14227 ( .A(n13823), .B(n13824), .Z(n13825) );
  XNOR U14228 ( .A(n13826), .B(n13825), .Z(n13811) );
  XOR U14229 ( .A(b[11]), .B(n28403), .Z(n13673) );
  OR U14230 ( .A(n13673), .B(n31369), .Z(n13354) );
  NANDN U14231 ( .A(n13352), .B(n31119), .Z(n13353) );
  NAND U14232 ( .A(n13354), .B(n13353), .Z(n13685) );
  XOR U14233 ( .A(b[43]), .B(n19656), .Z(n13676) );
  NANDN U14234 ( .A(n13676), .B(n37068), .Z(n13357) );
  NANDN U14235 ( .A(n13355), .B(n37069), .Z(n13356) );
  NAND U14236 ( .A(n13357), .B(n13356), .Z(n13682) );
  XNOR U14237 ( .A(b[45]), .B(a[31]), .Z(n13679) );
  NANDN U14238 ( .A(n13679), .B(n37261), .Z(n13360) );
  NANDN U14239 ( .A(n13358), .B(n37262), .Z(n13359) );
  AND U14240 ( .A(n13360), .B(n13359), .Z(n13683) );
  XNOR U14241 ( .A(n13682), .B(n13683), .Z(n13684) );
  XNOR U14242 ( .A(n13685), .B(n13684), .Z(n13709) );
  NANDN U14243 ( .A(n13361), .B(n37652), .Z(n13363) );
  XOR U14244 ( .A(b[49]), .B(n17960), .Z(n13664) );
  OR U14245 ( .A(n13664), .B(n37756), .Z(n13362) );
  NAND U14246 ( .A(n13363), .B(n13362), .Z(n13656) );
  NANDN U14247 ( .A(n13364), .B(n37469), .Z(n13366) );
  XNOR U14248 ( .A(n978), .B(a[29]), .Z(n13667) );
  NAND U14249 ( .A(n13667), .B(n37471), .Z(n13365) );
  NAND U14250 ( .A(n13366), .B(n13365), .Z(n13654) );
  NAND U14251 ( .A(n30846), .B(n13367), .Z(n13369) );
  XNOR U14252 ( .A(n969), .B(a[67]), .Z(n13670) );
  NAND U14253 ( .A(n30509), .B(n13670), .Z(n13368) );
  NAND U14254 ( .A(n13369), .B(n13368), .Z(n13655) );
  XNOR U14255 ( .A(n13654), .B(n13655), .Z(n13657) );
  XOR U14256 ( .A(n13656), .B(n13657), .Z(n13706) );
  NANDN U14257 ( .A(n13371), .B(n13370), .Z(n13375) );
  NAND U14258 ( .A(n13373), .B(n13372), .Z(n13374) );
  NAND U14259 ( .A(n13375), .B(n13374), .Z(n13707) );
  XNOR U14260 ( .A(n13706), .B(n13707), .Z(n13708) );
  XOR U14261 ( .A(n13709), .B(n13708), .Z(n13817) );
  XNOR U14262 ( .A(n13817), .B(n13818), .Z(n13820) );
  XNOR U14263 ( .A(b[35]), .B(a[41]), .Z(n13639) );
  NANDN U14264 ( .A(n13639), .B(n35985), .Z(n13382) );
  NANDN U14265 ( .A(n13380), .B(n35986), .Z(n13381) );
  NAND U14266 ( .A(n13382), .B(n13381), .Z(n13618) );
  XNOR U14267 ( .A(n31123), .B(a[69]), .Z(n13642) );
  NAND U14268 ( .A(n13642), .B(n29949), .Z(n13385) );
  NAND U14269 ( .A(n29948), .B(n13383), .Z(n13384) );
  NAND U14270 ( .A(n13385), .B(n13384), .Z(n13615) );
  XOR U14271 ( .A(b[55]), .B(n16220), .Z(n13645) );
  NANDN U14272 ( .A(n13645), .B(n38075), .Z(n13388) );
  NANDN U14273 ( .A(n13386), .B(n38073), .Z(n13387) );
  AND U14274 ( .A(n13388), .B(n13387), .Z(n13616) );
  XNOR U14275 ( .A(n13615), .B(n13616), .Z(n13617) );
  XNOR U14276 ( .A(n13618), .B(n13617), .Z(n13703) );
  NANDN U14277 ( .A(n13390), .B(n13389), .Z(n13394) );
  NAND U14278 ( .A(n13392), .B(n13391), .Z(n13393) );
  NAND U14279 ( .A(n13394), .B(n13393), .Z(n13700) );
  NANDN U14280 ( .A(n13396), .B(n13395), .Z(n13400) );
  NAND U14281 ( .A(n13398), .B(n13397), .Z(n13399) );
  NAND U14282 ( .A(n13400), .B(n13399), .Z(n13701) );
  XNOR U14283 ( .A(n13700), .B(n13701), .Z(n13702) );
  XOR U14284 ( .A(n13703), .B(n13702), .Z(n13819) );
  XNOR U14285 ( .A(n13820), .B(n13819), .Z(n13812) );
  XOR U14286 ( .A(n13811), .B(n13812), .Z(n13814) );
  NAND U14287 ( .A(n13402), .B(n13401), .Z(n13406) );
  NANDN U14288 ( .A(n13404), .B(n13403), .Z(n13405) );
  NAND U14289 ( .A(n13406), .B(n13405), .Z(n13813) );
  XNOR U14290 ( .A(n13814), .B(n13813), .Z(n13574) );
  NANDN U14291 ( .A(n13408), .B(n13407), .Z(n13412) );
  NAND U14292 ( .A(n13410), .B(n13409), .Z(n13411) );
  AND U14293 ( .A(n13412), .B(n13411), .Z(n13830) );
  NANDN U14294 ( .A(n13414), .B(n13413), .Z(n13418) );
  NANDN U14295 ( .A(n13416), .B(n13415), .Z(n13417) );
  NAND U14296 ( .A(n13418), .B(n13417), .Z(n13827) );
  NANDN U14297 ( .A(n13420), .B(n13419), .Z(n13424) );
  NAND U14298 ( .A(n13422), .B(n13421), .Z(n13423) );
  AND U14299 ( .A(n13424), .B(n13423), .Z(n13828) );
  XNOR U14300 ( .A(n13827), .B(n13828), .Z(n13829) );
  XNOR U14301 ( .A(n13830), .B(n13829), .Z(n13805) );
  NANDN U14302 ( .A(n13426), .B(n13425), .Z(n13430) );
  OR U14303 ( .A(n13428), .B(n13427), .Z(n13429) );
  AND U14304 ( .A(n13430), .B(n13429), .Z(n13806) );
  XNOR U14305 ( .A(n13805), .B(n13806), .Z(n13808) );
  NAND U14306 ( .A(n33283), .B(n13431), .Z(n13433) );
  XOR U14307 ( .A(n33020), .B(n26122), .Z(n13748) );
  NANDN U14308 ( .A(n33021), .B(n13748), .Z(n13432) );
  NAND U14309 ( .A(n13433), .B(n13432), .Z(n13772) );
  XNOR U14310 ( .A(b[21]), .B(a[55]), .Z(n13751) );
  OR U14311 ( .A(n13751), .B(n33634), .Z(n13436) );
  NANDN U14312 ( .A(n13434), .B(n33464), .Z(n13435) );
  NAND U14313 ( .A(n13436), .B(n13435), .Z(n13769) );
  NAND U14314 ( .A(n34044), .B(n13437), .Z(n13439) );
  XOR U14315 ( .A(n34510), .B(n25001), .Z(n13754) );
  NANDN U14316 ( .A(n33867), .B(n13754), .Z(n13438) );
  AND U14317 ( .A(n13439), .B(n13438), .Z(n13770) );
  XNOR U14318 ( .A(n13769), .B(n13770), .Z(n13771) );
  XOR U14319 ( .A(n13772), .B(n13771), .Z(n13658) );
  NANDN U14320 ( .A(n13441), .B(n13440), .Z(n13445) );
  NAND U14321 ( .A(n13443), .B(n13442), .Z(n13444) );
  NAND U14322 ( .A(n13445), .B(n13444), .Z(n13659) );
  XNOR U14323 ( .A(n13658), .B(n13659), .Z(n13661) );
  NAND U14324 ( .A(a[11]), .B(b[63]), .Z(n13651) );
  NANDN U14325 ( .A(n13446), .B(n38369), .Z(n13448) );
  XOR U14326 ( .A(b[61]), .B(n13976), .Z(n13742) );
  OR U14327 ( .A(n13742), .B(n38371), .Z(n13447) );
  NAND U14328 ( .A(n13448), .B(n13447), .Z(n13649) );
  NANDN U14329 ( .A(n13449), .B(n35311), .Z(n13451) );
  XOR U14330 ( .A(b[31]), .B(n22579), .Z(n13745) );
  NANDN U14331 ( .A(n13745), .B(n35313), .Z(n13450) );
  AND U14332 ( .A(n13451), .B(n13450), .Z(n13648) );
  XNOR U14333 ( .A(n13649), .B(n13648), .Z(n13650) );
  XNOR U14334 ( .A(n13651), .B(n13650), .Z(n13660) );
  XNOR U14335 ( .A(n13661), .B(n13660), .Z(n13799) );
  XOR U14336 ( .A(b[37]), .B(n20867), .Z(n13712) );
  NANDN U14337 ( .A(n13712), .B(n36311), .Z(n13454) );
  NANDN U14338 ( .A(n13452), .B(n36309), .Z(n13453) );
  NAND U14339 ( .A(n13454), .B(n13453), .Z(n13766) );
  XOR U14340 ( .A(a[71]), .B(n968), .Z(n13715) );
  OR U14341 ( .A(n13715), .B(n29363), .Z(n13457) );
  NANDN U14342 ( .A(n13455), .B(n29864), .Z(n13456) );
  NAND U14343 ( .A(n13457), .B(n13456), .Z(n13763) );
  XNOR U14344 ( .A(a[73]), .B(n967), .Z(n13718) );
  NAND U14345 ( .A(n13718), .B(n28939), .Z(n13460) );
  NAND U14346 ( .A(n28938), .B(n13458), .Z(n13459) );
  AND U14347 ( .A(n13460), .B(n13459), .Z(n13764) );
  XNOR U14348 ( .A(n13763), .B(n13764), .Z(n13765) );
  XOR U14349 ( .A(n13766), .B(n13765), .Z(n13691) );
  XNOR U14350 ( .A(b[13]), .B(a[63]), .Z(n13721) );
  OR U14351 ( .A(n13721), .B(n31550), .Z(n13463) );
  NANDN U14352 ( .A(n13461), .B(n31874), .Z(n13462) );
  NAND U14353 ( .A(n13463), .B(n13462), .Z(n13612) );
  NAND U14354 ( .A(n34848), .B(n13464), .Z(n13466) );
  XOR U14355 ( .A(n35375), .B(n23852), .Z(n13724) );
  NAND U14356 ( .A(n34618), .B(n13724), .Z(n13465) );
  NAND U14357 ( .A(n13466), .B(n13465), .Z(n13609) );
  NAND U14358 ( .A(n35188), .B(n13467), .Z(n13469) );
  XOR U14359 ( .A(n35540), .B(n23149), .Z(n13727) );
  NANDN U14360 ( .A(n34968), .B(n13727), .Z(n13468) );
  AND U14361 ( .A(n13469), .B(n13468), .Z(n13610) );
  XNOR U14362 ( .A(n13609), .B(n13610), .Z(n13611) );
  XOR U14363 ( .A(n13612), .B(n13611), .Z(n13689) );
  NANDN U14364 ( .A(n13471), .B(n13470), .Z(n13475) );
  NAND U14365 ( .A(n13473), .B(n13472), .Z(n13474) );
  AND U14366 ( .A(n13475), .B(n13474), .Z(n13688) );
  XOR U14367 ( .A(n13689), .B(n13688), .Z(n13690) );
  XOR U14368 ( .A(n13691), .B(n13690), .Z(n13800) );
  XOR U14369 ( .A(n13799), .B(n13800), .Z(n13802) );
  NANDN U14370 ( .A(n13477), .B(n13476), .Z(n13481) );
  NAND U14371 ( .A(n13479), .B(n13478), .Z(n13480) );
  NAND U14372 ( .A(n13481), .B(n13480), .Z(n13801) );
  XNOR U14373 ( .A(n13802), .B(n13801), .Z(n13587) );
  NANDN U14374 ( .A(n13483), .B(n13482), .Z(n13487) );
  NAND U14375 ( .A(n13485), .B(n13484), .Z(n13486) );
  NAND U14376 ( .A(n13487), .B(n13486), .Z(n13586) );
  NANDN U14377 ( .A(n13489), .B(n13488), .Z(n13493) );
  NAND U14378 ( .A(n13491), .B(n13490), .Z(n13492) );
  NAND U14379 ( .A(n13493), .B(n13492), .Z(n13697) );
  XNOR U14380 ( .A(b[41]), .B(a[35]), .Z(n13775) );
  OR U14381 ( .A(n13775), .B(n36905), .Z(n13496) );
  NANDN U14382 ( .A(n13494), .B(n36807), .Z(n13495) );
  NAND U14383 ( .A(n13496), .B(n13495), .Z(n13796) );
  XOR U14384 ( .A(b[57]), .B(n15113), .Z(n13778) );
  OR U14385 ( .A(n13778), .B(n965), .Z(n13499) );
  NANDN U14386 ( .A(n13497), .B(n38194), .Z(n13498) );
  NAND U14387 ( .A(n13499), .B(n13498), .Z(n13793) );
  NAND U14388 ( .A(n38326), .B(n13500), .Z(n13502) );
  XOR U14389 ( .A(n38400), .B(n14514), .Z(n13781) );
  NANDN U14390 ( .A(n38273), .B(n13781), .Z(n13501) );
  AND U14391 ( .A(n13502), .B(n13501), .Z(n13794) );
  XNOR U14392 ( .A(n13793), .B(n13794), .Z(n13795) );
  XOR U14393 ( .A(n13796), .B(n13795), .Z(n13627) );
  XOR U14394 ( .A(b[33]), .B(n21996), .Z(n13784) );
  NANDN U14395 ( .A(n13784), .B(n35620), .Z(n13505) );
  NANDN U14396 ( .A(n13503), .B(n35621), .Z(n13504) );
  NAND U14397 ( .A(n13505), .B(n13504), .Z(n13624) );
  NANDN U14398 ( .A(n966), .B(a[75]), .Z(n13506) );
  XOR U14399 ( .A(n29232), .B(n13506), .Z(n13508) );
  IV U14400 ( .A(a[74]), .Z(n31372) );
  NANDN U14401 ( .A(n31372), .B(n966), .Z(n13507) );
  AND U14402 ( .A(n13508), .B(n13507), .Z(n13621) );
  XOR U14403 ( .A(b[63]), .B(n13509), .Z(n13790) );
  NANDN U14404 ( .A(n13790), .B(n38422), .Z(n13512) );
  NANDN U14405 ( .A(n13510), .B(n38423), .Z(n13511) );
  AND U14406 ( .A(n13512), .B(n13511), .Z(n13622) );
  XNOR U14407 ( .A(n13621), .B(n13622), .Z(n13623) );
  XOR U14408 ( .A(n13624), .B(n13623), .Z(n13628) );
  XNOR U14409 ( .A(n13627), .B(n13628), .Z(n13630) );
  NANDN U14410 ( .A(n13514), .B(n13513), .Z(n13518) );
  NAND U14411 ( .A(n13516), .B(n13515), .Z(n13517) );
  NAND U14412 ( .A(n13518), .B(n13517), .Z(n13629) );
  XOR U14413 ( .A(n13630), .B(n13629), .Z(n13694) );
  NANDN U14414 ( .A(n13520), .B(n13519), .Z(n13524) );
  NAND U14415 ( .A(n13522), .B(n13521), .Z(n13523) );
  AND U14416 ( .A(n13524), .B(n13523), .Z(n13695) );
  XOR U14417 ( .A(n13694), .B(n13695), .Z(n13696) );
  XNOR U14418 ( .A(n13697), .B(n13696), .Z(n13585) );
  XNOR U14419 ( .A(n13586), .B(n13585), .Z(n13588) );
  XNOR U14420 ( .A(n13587), .B(n13588), .Z(n13807) );
  XNOR U14421 ( .A(n13808), .B(n13807), .Z(n13573) );
  XNOR U14422 ( .A(n13574), .B(n13573), .Z(n13576) );
  XOR U14423 ( .A(n13575), .B(n13576), .Z(n13834) );
  NANDN U14424 ( .A(n13526), .B(n13525), .Z(n13530) );
  NAND U14425 ( .A(n13528), .B(n13527), .Z(n13529) );
  NAND U14426 ( .A(n13530), .B(n13529), .Z(n13582) );
  OR U14427 ( .A(n13532), .B(n13531), .Z(n13536) );
  NAND U14428 ( .A(n13534), .B(n13533), .Z(n13535) );
  NAND U14429 ( .A(n13536), .B(n13535), .Z(n13580) );
  NANDN U14430 ( .A(n13538), .B(n13537), .Z(n13542) );
  NANDN U14431 ( .A(n13540), .B(n13539), .Z(n13541) );
  AND U14432 ( .A(n13542), .B(n13541), .Z(n13579) );
  XNOR U14433 ( .A(n13580), .B(n13579), .Z(n13581) );
  XNOR U14434 ( .A(n13582), .B(n13581), .Z(n13831) );
  OR U14435 ( .A(n13544), .B(n13543), .Z(n13548) );
  NAND U14436 ( .A(n13546), .B(n13545), .Z(n13547) );
  NAND U14437 ( .A(n13548), .B(n13547), .Z(n13832) );
  XNOR U14438 ( .A(n13839), .B(n13840), .Z(n13845) );
  NANDN U14439 ( .A(n13553), .B(n13552), .Z(n13557) );
  NAND U14440 ( .A(n13555), .B(n13554), .Z(n13556) );
  AND U14441 ( .A(n13557), .B(n13556), .Z(n13843) );
  XNOR U14442 ( .A(n13844), .B(n13843), .Z(n13846) );
  XNOR U14443 ( .A(n13845), .B(n13846), .Z(n13569) );
  NANDN U14444 ( .A(n13559), .B(n13558), .Z(n13563) );
  NANDN U14445 ( .A(n13561), .B(n13560), .Z(n13562) );
  NAND U14446 ( .A(n13563), .B(n13562), .Z(n13570) );
  XNOR U14447 ( .A(n13569), .B(n13570), .Z(n13571) );
  XNOR U14448 ( .A(n13572), .B(n13571), .Z(n13847) );
  XNOR U14449 ( .A(n13847), .B(sreg[139]), .Z(n13849) );
  NAND U14450 ( .A(n13564), .B(sreg[138]), .Z(n13568) );
  OR U14451 ( .A(n13566), .B(n13565), .Z(n13567) );
  AND U14452 ( .A(n13568), .B(n13567), .Z(n13848) );
  XOR U14453 ( .A(n13849), .B(n13848), .Z(c[139]) );
  NAND U14454 ( .A(n13574), .B(n13573), .Z(n13578) );
  NANDN U14455 ( .A(n13576), .B(n13575), .Z(n13577) );
  NAND U14456 ( .A(n13578), .B(n13577), .Z(n13856) );
  NANDN U14457 ( .A(n13580), .B(n13579), .Z(n13584) );
  NANDN U14458 ( .A(n13582), .B(n13581), .Z(n13583) );
  NAND U14459 ( .A(n13584), .B(n13583), .Z(n13857) );
  XNOR U14460 ( .A(n13856), .B(n13857), .Z(n13858) );
  NAND U14461 ( .A(n13586), .B(n13585), .Z(n13590) );
  NANDN U14462 ( .A(n13588), .B(n13587), .Z(n13589) );
  NAND U14463 ( .A(n13590), .B(n13589), .Z(n14109) );
  XOR U14464 ( .A(b[39]), .B(n20686), .Z(n14017) );
  NANDN U14465 ( .A(n14017), .B(n36553), .Z(n13593) );
  NANDN U14466 ( .A(n13591), .B(n36643), .Z(n13592) );
  NAND U14467 ( .A(n13593), .B(n13592), .Z(n13946) );
  XOR U14468 ( .A(b[51]), .B(n17133), .Z(n14020) );
  NANDN U14469 ( .A(n14020), .B(n37803), .Z(n13596) );
  NANDN U14470 ( .A(n13594), .B(n37802), .Z(n13595) );
  NAND U14471 ( .A(n13596), .B(n13595), .Z(n13943) );
  XOR U14472 ( .A(b[53]), .B(n16508), .Z(n14023) );
  NANDN U14473 ( .A(n14023), .B(n37940), .Z(n13599) );
  NANDN U14474 ( .A(n13597), .B(n37941), .Z(n13598) );
  AND U14475 ( .A(n13599), .B(n13598), .Z(n13944) );
  XNOR U14476 ( .A(n13943), .B(n13944), .Z(n13945) );
  XNOR U14477 ( .A(n13946), .B(n13945), .Z(n13949) );
  XNOR U14478 ( .A(b[15]), .B(a[62]), .Z(n14008) );
  OR U14479 ( .A(n14008), .B(n32010), .Z(n13602) );
  NANDN U14480 ( .A(n13600), .B(n32011), .Z(n13601) );
  NAND U14481 ( .A(n13602), .B(n13601), .Z(n13916) );
  XNOR U14482 ( .A(b[25]), .B(n25134), .Z(n14011) );
  NANDN U14483 ( .A(n34219), .B(n14011), .Z(n13605) );
  NAND U14484 ( .A(n34217), .B(n13603), .Z(n13604) );
  NAND U14485 ( .A(n13605), .B(n13604), .Z(n13913) );
  XNOR U14486 ( .A(b[17]), .B(a[60]), .Z(n14014) );
  NANDN U14487 ( .A(n14014), .B(n32543), .Z(n13608) );
  NAND U14488 ( .A(n13606), .B(n32541), .Z(n13607) );
  AND U14489 ( .A(n13608), .B(n13607), .Z(n13914) );
  XNOR U14490 ( .A(n13913), .B(n13914), .Z(n13915) );
  XOR U14491 ( .A(n13916), .B(n13915), .Z(n13950) );
  XOR U14492 ( .A(n13949), .B(n13950), .Z(n13952) );
  NANDN U14493 ( .A(n13610), .B(n13609), .Z(n13614) );
  NAND U14494 ( .A(n13612), .B(n13611), .Z(n13613) );
  NAND U14495 ( .A(n13614), .B(n13613), .Z(n13951) );
  XNOR U14496 ( .A(n13952), .B(n13951), .Z(n13999) );
  NANDN U14497 ( .A(n13616), .B(n13615), .Z(n13620) );
  NAND U14498 ( .A(n13618), .B(n13617), .Z(n13619) );
  NAND U14499 ( .A(n13620), .B(n13619), .Z(n13996) );
  NANDN U14500 ( .A(n13622), .B(n13621), .Z(n13626) );
  NAND U14501 ( .A(n13624), .B(n13623), .Z(n13625) );
  AND U14502 ( .A(n13626), .B(n13625), .Z(n13997) );
  XNOR U14503 ( .A(n13996), .B(n13997), .Z(n13998) );
  XNOR U14504 ( .A(n13999), .B(n13998), .Z(n14101) );
  OR U14505 ( .A(n13628), .B(n13627), .Z(n13632) );
  OR U14506 ( .A(n13630), .B(n13629), .Z(n13631) );
  AND U14507 ( .A(n13632), .B(n13631), .Z(n14102) );
  XNOR U14508 ( .A(n14101), .B(n14102), .Z(n14103) );
  NANDN U14509 ( .A(n13634), .B(n13633), .Z(n13638) );
  NAND U14510 ( .A(n13636), .B(n13635), .Z(n13637) );
  AND U14511 ( .A(n13638), .B(n13637), .Z(n14104) );
  XNOR U14512 ( .A(n14103), .B(n14104), .Z(n14108) );
  XNOR U14513 ( .A(b[35]), .B(a[42]), .Z(n14070) );
  NANDN U14514 ( .A(n14070), .B(n35985), .Z(n13641) );
  NANDN U14515 ( .A(n13639), .B(n35986), .Z(n13640) );
  NAND U14516 ( .A(n13641), .B(n13640), .Z(n14035) );
  XOR U14517 ( .A(n31123), .B(n30379), .Z(n14073) );
  NAND U14518 ( .A(n14073), .B(n29949), .Z(n13644) );
  NAND U14519 ( .A(n29948), .B(n13642), .Z(n13643) );
  NAND U14520 ( .A(n13644), .B(n13643), .Z(n14032) );
  XOR U14521 ( .A(b[55]), .B(n15963), .Z(n14076) );
  NANDN U14522 ( .A(n14076), .B(n38075), .Z(n13647) );
  NANDN U14523 ( .A(n13645), .B(n38073), .Z(n13646) );
  AND U14524 ( .A(n13647), .B(n13646), .Z(n14033) );
  XNOR U14525 ( .A(n14032), .B(n14033), .Z(n14034) );
  XNOR U14526 ( .A(n14035), .B(n14034), .Z(n13877) );
  NANDN U14527 ( .A(n13649), .B(n13648), .Z(n13653) );
  NAND U14528 ( .A(n13651), .B(n13650), .Z(n13652) );
  NAND U14529 ( .A(n13653), .B(n13652), .Z(n13874) );
  XNOR U14530 ( .A(n13874), .B(n13875), .Z(n13876) );
  XOR U14531 ( .A(n13877), .B(n13876), .Z(n14093) );
  OR U14532 ( .A(n13659), .B(n13658), .Z(n13663) );
  OR U14533 ( .A(n13661), .B(n13660), .Z(n13662) );
  NAND U14534 ( .A(n13663), .B(n13662), .Z(n14091) );
  XOR U14535 ( .A(b[49]), .B(n17702), .Z(n14042) );
  OR U14536 ( .A(n14042), .B(n37756), .Z(n13666) );
  NANDN U14537 ( .A(n13664), .B(n37652), .Z(n13665) );
  NAND U14538 ( .A(n13666), .B(n13665), .Z(n14088) );
  NAND U14539 ( .A(n13667), .B(n37469), .Z(n13669) );
  XOR U14540 ( .A(n978), .B(n18804), .Z(n14045) );
  NAND U14541 ( .A(n14045), .B(n37471), .Z(n13668) );
  NAND U14542 ( .A(n13669), .B(n13668), .Z(n14085) );
  XOR U14543 ( .A(b[9]), .B(n29868), .Z(n14048) );
  NANDN U14544 ( .A(n14048), .B(n30509), .Z(n13672) );
  NAND U14545 ( .A(n13670), .B(n30846), .Z(n13671) );
  AND U14546 ( .A(n13672), .B(n13671), .Z(n14086) );
  XNOR U14547 ( .A(n14085), .B(n14086), .Z(n14087) );
  XNOR U14548 ( .A(n14088), .B(n14087), .Z(n13898) );
  XOR U14549 ( .A(b[11]), .B(n28701), .Z(n14051) );
  OR U14550 ( .A(n14051), .B(n31369), .Z(n13675) );
  NANDN U14551 ( .A(n13673), .B(n31119), .Z(n13674) );
  NAND U14552 ( .A(n13675), .B(n13674), .Z(n14063) );
  XOR U14553 ( .A(b[43]), .B(n19513), .Z(n14054) );
  NANDN U14554 ( .A(n14054), .B(n37068), .Z(n13678) );
  NANDN U14555 ( .A(n13676), .B(n37069), .Z(n13677) );
  NAND U14556 ( .A(n13678), .B(n13677), .Z(n14060) );
  XNOR U14557 ( .A(b[45]), .B(a[32]), .Z(n14057) );
  NANDN U14558 ( .A(n14057), .B(n37261), .Z(n13681) );
  NANDN U14559 ( .A(n13679), .B(n37262), .Z(n13680) );
  AND U14560 ( .A(n13681), .B(n13680), .Z(n14061) );
  XNOR U14561 ( .A(n14060), .B(n14061), .Z(n14062) );
  XOR U14562 ( .A(n14063), .B(n14062), .Z(n13899) );
  XNOR U14563 ( .A(n13898), .B(n13899), .Z(n13900) );
  NANDN U14564 ( .A(n13683), .B(n13682), .Z(n13687) );
  NAND U14565 ( .A(n13685), .B(n13684), .Z(n13686) );
  AND U14566 ( .A(n13687), .B(n13686), .Z(n13901) );
  XNOR U14567 ( .A(n13900), .B(n13901), .Z(n14092) );
  XNOR U14568 ( .A(n14091), .B(n14092), .Z(n14094) );
  XOR U14569 ( .A(n14093), .B(n14094), .Z(n14107) );
  XNOR U14570 ( .A(n14108), .B(n14107), .Z(n14110) );
  XNOR U14571 ( .A(n14109), .B(n14110), .Z(n14117) );
  NANDN U14572 ( .A(n13689), .B(n13688), .Z(n13693) );
  OR U14573 ( .A(n13691), .B(n13690), .Z(n13692) );
  NAND U14574 ( .A(n13693), .B(n13692), .Z(n14099) );
  NAND U14575 ( .A(n13695), .B(n13694), .Z(n13699) );
  NANDN U14576 ( .A(n13697), .B(n13696), .Z(n13698) );
  NAND U14577 ( .A(n13699), .B(n13698), .Z(n14097) );
  NANDN U14578 ( .A(n13701), .B(n13700), .Z(n13705) );
  NAND U14579 ( .A(n13703), .B(n13702), .Z(n13704) );
  NAND U14580 ( .A(n13705), .B(n13704), .Z(n14098) );
  XNOR U14581 ( .A(n14097), .B(n14098), .Z(n14100) );
  XOR U14582 ( .A(n14099), .B(n14100), .Z(n13871) );
  NANDN U14583 ( .A(n13707), .B(n13706), .Z(n13711) );
  NAND U14584 ( .A(n13709), .B(n13708), .Z(n13710) );
  NAND U14585 ( .A(n13711), .B(n13710), .Z(n13894) );
  XOR U14586 ( .A(b[37]), .B(n21149), .Z(n13934) );
  NANDN U14587 ( .A(n13934), .B(n36311), .Z(n13714) );
  NANDN U14588 ( .A(n13712), .B(n36309), .Z(n13713) );
  NAND U14589 ( .A(n13714), .B(n13713), .Z(n13958) );
  XOR U14590 ( .A(a[72]), .B(n968), .Z(n13937) );
  OR U14591 ( .A(n13937), .B(n29363), .Z(n13717) );
  NANDN U14592 ( .A(n13715), .B(n29864), .Z(n13716) );
  NAND U14593 ( .A(n13717), .B(n13716), .Z(n13955) );
  XOR U14594 ( .A(n31372), .B(n967), .Z(n13940) );
  NAND U14595 ( .A(n13940), .B(n28939), .Z(n13720) );
  NAND U14596 ( .A(n28938), .B(n13718), .Z(n13719) );
  AND U14597 ( .A(n13720), .B(n13719), .Z(n13956) );
  XNOR U14598 ( .A(n13955), .B(n13956), .Z(n13957) );
  XOR U14599 ( .A(n13958), .B(n13957), .Z(n13883) );
  XNOR U14600 ( .A(b[13]), .B(a[64]), .Z(n13925) );
  OR U14601 ( .A(n13925), .B(n31550), .Z(n13723) );
  NANDN U14602 ( .A(n13721), .B(n31874), .Z(n13722) );
  NAND U14603 ( .A(n13723), .B(n13722), .Z(n14029) );
  NAND U14604 ( .A(n34848), .B(n13724), .Z(n13726) );
  XOR U14605 ( .A(n35375), .B(n24671), .Z(n13928) );
  NAND U14606 ( .A(n34618), .B(n13928), .Z(n13725) );
  NAND U14607 ( .A(n13726), .B(n13725), .Z(n14026) );
  NAND U14608 ( .A(n35188), .B(n13727), .Z(n13729) );
  XOR U14609 ( .A(n35540), .B(n23447), .Z(n13931) );
  NANDN U14610 ( .A(n34968), .B(n13931), .Z(n13728) );
  AND U14611 ( .A(n13729), .B(n13728), .Z(n14027) );
  XNOR U14612 ( .A(n14026), .B(n14027), .Z(n14028) );
  XOR U14613 ( .A(n14029), .B(n14028), .Z(n13881) );
  NANDN U14614 ( .A(n13731), .B(n13730), .Z(n13735) );
  NAND U14615 ( .A(n13733), .B(n13732), .Z(n13734) );
  AND U14616 ( .A(n13735), .B(n13734), .Z(n13880) );
  XOR U14617 ( .A(n13881), .B(n13880), .Z(n13882) );
  XOR U14618 ( .A(n13883), .B(n13882), .Z(n13893) );
  NANDN U14619 ( .A(n13737), .B(n13736), .Z(n13741) );
  NAND U14620 ( .A(n13739), .B(n13738), .Z(n13740) );
  NAND U14621 ( .A(n13741), .B(n13740), .Z(n14068) );
  NAND U14622 ( .A(a[12]), .B(b[63]), .Z(n14082) );
  NANDN U14623 ( .A(n13742), .B(n38369), .Z(n13744) );
  XOR U14624 ( .A(b[61]), .B(n14259), .Z(n13919) );
  OR U14625 ( .A(n13919), .B(n38371), .Z(n13743) );
  NAND U14626 ( .A(n13744), .B(n13743), .Z(n14080) );
  NANDN U14627 ( .A(n13745), .B(n35311), .Z(n13747) );
  XOR U14628 ( .A(b[31]), .B(n22964), .Z(n13922) );
  NANDN U14629 ( .A(n13922), .B(n35313), .Z(n13746) );
  AND U14630 ( .A(n13747), .B(n13746), .Z(n14079) );
  XNOR U14631 ( .A(n14080), .B(n14079), .Z(n14081) );
  XOR U14632 ( .A(n14082), .B(n14081), .Z(n14066) );
  NAND U14633 ( .A(n33283), .B(n13748), .Z(n13750) );
  XOR U14634 ( .A(n33020), .B(n26347), .Z(n13904) );
  NANDN U14635 ( .A(n33021), .B(n13904), .Z(n13749) );
  NAND U14636 ( .A(n13750), .B(n13749), .Z(n13983) );
  XNOR U14637 ( .A(b[21]), .B(a[56]), .Z(n13907) );
  OR U14638 ( .A(n13907), .B(n33634), .Z(n13753) );
  NANDN U14639 ( .A(n13751), .B(n33464), .Z(n13752) );
  NAND U14640 ( .A(n13753), .B(n13752), .Z(n13980) );
  NAND U14641 ( .A(n34044), .B(n13754), .Z(n13756) );
  XOR U14642 ( .A(n34510), .B(n25177), .Z(n13910) );
  NANDN U14643 ( .A(n33867), .B(n13910), .Z(n13755) );
  AND U14644 ( .A(n13756), .B(n13755), .Z(n13981) );
  XNOR U14645 ( .A(n13980), .B(n13981), .Z(n13982) );
  XNOR U14646 ( .A(n13983), .B(n13982), .Z(n14067) );
  XNOR U14647 ( .A(n14066), .B(n14067), .Z(n14069) );
  XNOR U14648 ( .A(n14068), .B(n14069), .Z(n13892) );
  XOR U14649 ( .A(n13893), .B(n13892), .Z(n13895) );
  XNOR U14650 ( .A(n13894), .B(n13895), .Z(n13995) );
  NANDN U14651 ( .A(n13758), .B(n13757), .Z(n13762) );
  NANDN U14652 ( .A(n13760), .B(n13759), .Z(n13761) );
  NAND U14653 ( .A(n13762), .B(n13761), .Z(n13993) );
  NANDN U14654 ( .A(n13764), .B(n13763), .Z(n13768) );
  NAND U14655 ( .A(n13766), .B(n13765), .Z(n13767) );
  NAND U14656 ( .A(n13768), .B(n13767), .Z(n13889) );
  NANDN U14657 ( .A(n13770), .B(n13769), .Z(n13774) );
  NAND U14658 ( .A(n13772), .B(n13771), .Z(n13773) );
  NAND U14659 ( .A(n13774), .B(n13773), .Z(n14005) );
  XNOR U14660 ( .A(b[41]), .B(a[36]), .Z(n13961) );
  OR U14661 ( .A(n13961), .B(n36905), .Z(n13777) );
  NANDN U14662 ( .A(n13775), .B(n36807), .Z(n13776) );
  NAND U14663 ( .A(n13777), .B(n13776), .Z(n13989) );
  XOR U14664 ( .A(b[57]), .B(n15484), .Z(n13964) );
  OR U14665 ( .A(n13964), .B(n965), .Z(n13780) );
  NANDN U14666 ( .A(n13778), .B(n38194), .Z(n13779) );
  NAND U14667 ( .A(n13780), .B(n13779), .Z(n13986) );
  NAND U14668 ( .A(n38326), .B(n13781), .Z(n13783) );
  XOR U14669 ( .A(n38400), .B(n14905), .Z(n13967) );
  NANDN U14670 ( .A(n38273), .B(n13967), .Z(n13782) );
  AND U14671 ( .A(n13783), .B(n13782), .Z(n13987) );
  XNOR U14672 ( .A(n13986), .B(n13987), .Z(n13988) );
  XOR U14673 ( .A(n13989), .B(n13988), .Z(n14003) );
  XOR U14674 ( .A(b[33]), .B(n22289), .Z(n13970) );
  NANDN U14675 ( .A(n13970), .B(n35620), .Z(n13786) );
  NANDN U14676 ( .A(n13784), .B(n35621), .Z(n13785) );
  NAND U14677 ( .A(n13786), .B(n13785), .Z(n14041) );
  NANDN U14678 ( .A(n966), .B(a[76]), .Z(n13787) );
  XOR U14679 ( .A(n29232), .B(n13787), .Z(n13789) );
  NANDN U14680 ( .A(b[0]), .B(a[75]), .Z(n13788) );
  AND U14681 ( .A(n13789), .B(n13788), .Z(n14038) );
  XOR U14682 ( .A(b[63]), .B(n14210), .Z(n13977) );
  NANDN U14683 ( .A(n13977), .B(n38422), .Z(n13792) );
  NANDN U14684 ( .A(n13790), .B(n38423), .Z(n13791) );
  AND U14685 ( .A(n13792), .B(n13791), .Z(n14039) );
  XNOR U14686 ( .A(n14038), .B(n14039), .Z(n14040) );
  XNOR U14687 ( .A(n14041), .B(n14040), .Z(n14002) );
  XOR U14688 ( .A(n14003), .B(n14002), .Z(n14004) );
  XNOR U14689 ( .A(n14005), .B(n14004), .Z(n13887) );
  NANDN U14690 ( .A(n13794), .B(n13793), .Z(n13798) );
  NAND U14691 ( .A(n13796), .B(n13795), .Z(n13797) );
  AND U14692 ( .A(n13798), .B(n13797), .Z(n13886) );
  XNOR U14693 ( .A(n13887), .B(n13886), .Z(n13888) );
  XNOR U14694 ( .A(n13889), .B(n13888), .Z(n13992) );
  XOR U14695 ( .A(n13993), .B(n13992), .Z(n13994) );
  XNOR U14696 ( .A(n13995), .B(n13994), .Z(n13868) );
  NANDN U14697 ( .A(n13800), .B(n13799), .Z(n13804) );
  OR U14698 ( .A(n13802), .B(n13801), .Z(n13803) );
  AND U14699 ( .A(n13804), .B(n13803), .Z(n13869) );
  XNOR U14700 ( .A(n13868), .B(n13869), .Z(n13870) );
  XNOR U14701 ( .A(n13871), .B(n13870), .Z(n14118) );
  XOR U14702 ( .A(n14117), .B(n14118), .Z(n14120) );
  NAND U14703 ( .A(n13806), .B(n13805), .Z(n13810) );
  NANDN U14704 ( .A(n13808), .B(n13807), .Z(n13809) );
  NAND U14705 ( .A(n13810), .B(n13809), .Z(n14119) );
  XNOR U14706 ( .A(n14120), .B(n14119), .Z(n13865) );
  NANDN U14707 ( .A(n13812), .B(n13811), .Z(n13816) );
  OR U14708 ( .A(n13814), .B(n13813), .Z(n13815) );
  NAND U14709 ( .A(n13816), .B(n13815), .Z(n13863) );
  NAND U14710 ( .A(n13818), .B(n13817), .Z(n13822) );
  NANDN U14711 ( .A(n13820), .B(n13819), .Z(n13821) );
  NAND U14712 ( .A(n13822), .B(n13821), .Z(n14114) );
  XNOR U14713 ( .A(n14111), .B(n14112), .Z(n14113) );
  XOR U14714 ( .A(n14114), .B(n14113), .Z(n13862) );
  XNOR U14715 ( .A(n13863), .B(n13862), .Z(n13864) );
  XNOR U14716 ( .A(n13865), .B(n13864), .Z(n13859) );
  XOR U14717 ( .A(n13858), .B(n13859), .Z(n14126) );
  OR U14718 ( .A(n13832), .B(n13831), .Z(n13836) );
  NANDN U14719 ( .A(n13834), .B(n13833), .Z(n13835) );
  NAND U14720 ( .A(n13836), .B(n13835), .Z(n14124) );
  NANDN U14721 ( .A(n13838), .B(n13837), .Z(n13842) );
  NAND U14722 ( .A(n13840), .B(n13839), .Z(n13841) );
  AND U14723 ( .A(n13842), .B(n13841), .Z(n14123) );
  XNOR U14724 ( .A(n14124), .B(n14123), .Z(n14125) );
  XNOR U14725 ( .A(n14126), .B(n14125), .Z(n13852) );
  XNOR U14726 ( .A(n13852), .B(n13853), .Z(n13854) );
  XNOR U14727 ( .A(n13855), .B(n13854), .Z(n14129) );
  XNOR U14728 ( .A(n14129), .B(sreg[140]), .Z(n14131) );
  NAND U14729 ( .A(n13847), .B(sreg[139]), .Z(n13851) );
  OR U14730 ( .A(n13849), .B(n13848), .Z(n13850) );
  AND U14731 ( .A(n13851), .B(n13850), .Z(n14130) );
  XOR U14732 ( .A(n14131), .B(n14130), .Z(c[140]) );
  NANDN U14733 ( .A(n13857), .B(n13856), .Z(n13861) );
  NANDN U14734 ( .A(n13859), .B(n13858), .Z(n13860) );
  NAND U14735 ( .A(n13861), .B(n13860), .Z(n14412) );
  NANDN U14736 ( .A(n13863), .B(n13862), .Z(n13867) );
  NAND U14737 ( .A(n13865), .B(n13864), .Z(n13866) );
  NAND U14738 ( .A(n13867), .B(n13866), .Z(n14411) );
  NANDN U14739 ( .A(n13869), .B(n13868), .Z(n13873) );
  NAND U14740 ( .A(n13871), .B(n13870), .Z(n13872) );
  NAND U14741 ( .A(n13873), .B(n13872), .Z(n14149) );
  NANDN U14742 ( .A(n13875), .B(n13874), .Z(n13879) );
  NAND U14743 ( .A(n13877), .B(n13876), .Z(n13878) );
  NAND U14744 ( .A(n13879), .B(n13878), .Z(n14397) );
  NANDN U14745 ( .A(n13881), .B(n13880), .Z(n13885) );
  OR U14746 ( .A(n13883), .B(n13882), .Z(n13884) );
  NAND U14747 ( .A(n13885), .B(n13884), .Z(n14395) );
  NANDN U14748 ( .A(n13887), .B(n13886), .Z(n13891) );
  NANDN U14749 ( .A(n13889), .B(n13888), .Z(n13890) );
  AND U14750 ( .A(n13891), .B(n13890), .Z(n14394) );
  XNOR U14751 ( .A(n14395), .B(n14394), .Z(n14396) );
  XNOR U14752 ( .A(n14397), .B(n14396), .Z(n14372) );
  NANDN U14753 ( .A(n13893), .B(n13892), .Z(n13897) );
  OR U14754 ( .A(n13895), .B(n13894), .Z(n13896) );
  NAND U14755 ( .A(n13897), .B(n13896), .Z(n14373) );
  XOR U14756 ( .A(n14372), .B(n14373), .Z(n14374) );
  NANDN U14757 ( .A(n13899), .B(n13898), .Z(n13903) );
  NAND U14758 ( .A(n13901), .B(n13900), .Z(n13902) );
  NAND U14759 ( .A(n13903), .B(n13902), .Z(n14170) );
  NAND U14760 ( .A(n33283), .B(n13904), .Z(n13906) );
  XNOR U14761 ( .A(n33020), .B(a[59]), .Z(n14217) );
  NANDN U14762 ( .A(n33021), .B(n14217), .Z(n13905) );
  NAND U14763 ( .A(n13906), .B(n13905), .Z(n14241) );
  XNOR U14764 ( .A(b[21]), .B(a[57]), .Z(n14220) );
  OR U14765 ( .A(n14220), .B(n33634), .Z(n13909) );
  NANDN U14766 ( .A(n13907), .B(n33464), .Z(n13908) );
  NAND U14767 ( .A(n13909), .B(n13908), .Z(n14238) );
  NAND U14768 ( .A(n34044), .B(n13910), .Z(n13912) );
  XOR U14769 ( .A(n34510), .B(n25466), .Z(n14223) );
  NANDN U14770 ( .A(n33867), .B(n14223), .Z(n13911) );
  AND U14771 ( .A(n13912), .B(n13911), .Z(n14239) );
  XNOR U14772 ( .A(n14238), .B(n14239), .Z(n14240) );
  XOR U14773 ( .A(n14241), .B(n14240), .Z(n14275) );
  NANDN U14774 ( .A(n13914), .B(n13913), .Z(n13918) );
  NAND U14775 ( .A(n13916), .B(n13915), .Z(n13917) );
  NAND U14776 ( .A(n13918), .B(n13917), .Z(n14276) );
  XNOR U14777 ( .A(n14275), .B(n14276), .Z(n14278) );
  NAND U14778 ( .A(a[13]), .B(b[63]), .Z(n14317) );
  NANDN U14779 ( .A(n13919), .B(n38369), .Z(n13921) );
  XOR U14780 ( .A(b[61]), .B(n14514), .Z(n14211) );
  OR U14781 ( .A(n14211), .B(n38371), .Z(n13920) );
  NAND U14782 ( .A(n13921), .B(n13920), .Z(n14315) );
  NANDN U14783 ( .A(n13922), .B(n35311), .Z(n13924) );
  XOR U14784 ( .A(b[31]), .B(n23149), .Z(n14214) );
  NANDN U14785 ( .A(n14214), .B(n35313), .Z(n13923) );
  AND U14786 ( .A(n13924), .B(n13923), .Z(n14314) );
  XNOR U14787 ( .A(n14315), .B(n14314), .Z(n14316) );
  XNOR U14788 ( .A(n14317), .B(n14316), .Z(n14277) );
  XNOR U14789 ( .A(n14278), .B(n14277), .Z(n14168) );
  XOR U14790 ( .A(b[13]), .B(n28403), .Z(n14189) );
  OR U14791 ( .A(n14189), .B(n31550), .Z(n13927) );
  NANDN U14792 ( .A(n13925), .B(n31874), .Z(n13926) );
  NAND U14793 ( .A(n13927), .B(n13926), .Z(n14363) );
  NAND U14794 ( .A(n34848), .B(n13928), .Z(n13930) );
  XOR U14795 ( .A(n35375), .B(n24288), .Z(n14192) );
  NAND U14796 ( .A(n34618), .B(n14192), .Z(n13929) );
  NAND U14797 ( .A(n13930), .B(n13929), .Z(n14360) );
  NAND U14798 ( .A(n35188), .B(n13931), .Z(n13933) );
  XOR U14799 ( .A(n35540), .B(n23852), .Z(n14195) );
  NANDN U14800 ( .A(n34968), .B(n14195), .Z(n13932) );
  AND U14801 ( .A(n13933), .B(n13932), .Z(n14361) );
  XNOR U14802 ( .A(n14360), .B(n14361), .Z(n14362) );
  XNOR U14803 ( .A(n14363), .B(n14362), .Z(n14162) );
  XOR U14804 ( .A(b[37]), .B(n21441), .Z(n14180) );
  NANDN U14805 ( .A(n14180), .B(n36311), .Z(n13936) );
  NANDN U14806 ( .A(n13934), .B(n36309), .Z(n13935) );
  NAND U14807 ( .A(n13936), .B(n13935), .Z(n14235) );
  XNOR U14808 ( .A(a[73]), .B(b[5]), .Z(n14183) );
  OR U14809 ( .A(n14183), .B(n29363), .Z(n13939) );
  NANDN U14810 ( .A(n13937), .B(n29864), .Z(n13938) );
  NAND U14811 ( .A(n13939), .B(n13938), .Z(n14232) );
  XNOR U14812 ( .A(a[75]), .B(n967), .Z(n14186) );
  NAND U14813 ( .A(n14186), .B(n28939), .Z(n13942) );
  NAND U14814 ( .A(n28938), .B(n13940), .Z(n13941) );
  AND U14815 ( .A(n13942), .B(n13941), .Z(n14233) );
  XNOR U14816 ( .A(n14232), .B(n14233), .Z(n14234) );
  XOR U14817 ( .A(n14235), .B(n14234), .Z(n14163) );
  XOR U14818 ( .A(n14162), .B(n14163), .Z(n14165) );
  NANDN U14819 ( .A(n13944), .B(n13943), .Z(n13948) );
  NAND U14820 ( .A(n13946), .B(n13945), .Z(n13947) );
  NAND U14821 ( .A(n13948), .B(n13947), .Z(n14164) );
  XOR U14822 ( .A(n14165), .B(n14164), .Z(n14169) );
  XOR U14823 ( .A(n14168), .B(n14169), .Z(n14171) );
  XNOR U14824 ( .A(n14170), .B(n14171), .Z(n14271) );
  NANDN U14825 ( .A(n13950), .B(n13949), .Z(n13954) );
  OR U14826 ( .A(n13952), .B(n13951), .Z(n13953) );
  NAND U14827 ( .A(n13954), .B(n13953), .Z(n14270) );
  NANDN U14828 ( .A(n13956), .B(n13955), .Z(n13960) );
  NAND U14829 ( .A(n13958), .B(n13957), .Z(n13959) );
  NAND U14830 ( .A(n13960), .B(n13959), .Z(n14159) );
  XNOR U14831 ( .A(b[41]), .B(a[37]), .Z(n14244) );
  OR U14832 ( .A(n14244), .B(n36905), .Z(n13963) );
  NANDN U14833 ( .A(n13961), .B(n36807), .Z(n13962) );
  NAND U14834 ( .A(n13963), .B(n13962), .Z(n14266) );
  XOR U14835 ( .A(b[57]), .B(n16220), .Z(n14247) );
  OR U14836 ( .A(n14247), .B(n965), .Z(n13966) );
  NANDN U14837 ( .A(n13964), .B(n38194), .Z(n13965) );
  NAND U14838 ( .A(n13966), .B(n13965), .Z(n14263) );
  NAND U14839 ( .A(n38326), .B(n13967), .Z(n13969) );
  XOR U14840 ( .A(n38400), .B(n15113), .Z(n14250) );
  NANDN U14841 ( .A(n38273), .B(n14250), .Z(n13968) );
  AND U14842 ( .A(n13969), .B(n13968), .Z(n14264) );
  XNOR U14843 ( .A(n14263), .B(n14264), .Z(n14265) );
  XOR U14844 ( .A(n14266), .B(n14265), .Z(n14326) );
  XOR U14845 ( .A(b[33]), .B(n22579), .Z(n14253) );
  NANDN U14846 ( .A(n14253), .B(n35620), .Z(n13972) );
  NANDN U14847 ( .A(n13970), .B(n35621), .Z(n13971) );
  NAND U14848 ( .A(n13972), .B(n13971), .Z(n14339) );
  NANDN U14849 ( .A(n966), .B(a[77]), .Z(n13973) );
  XOR U14850 ( .A(n29232), .B(n13973), .Z(n13975) );
  IV U14851 ( .A(a[76]), .Z(n31363) );
  NANDN U14852 ( .A(n31363), .B(n966), .Z(n13974) );
  AND U14853 ( .A(n13975), .B(n13974), .Z(n14336) );
  XOR U14854 ( .A(b[63]), .B(n13976), .Z(n14260) );
  NANDN U14855 ( .A(n14260), .B(n38422), .Z(n13979) );
  NANDN U14856 ( .A(n13977), .B(n38423), .Z(n13978) );
  AND U14857 ( .A(n13979), .B(n13978), .Z(n14337) );
  XNOR U14858 ( .A(n14336), .B(n14337), .Z(n14338) );
  XOR U14859 ( .A(n14339), .B(n14338), .Z(n14327) );
  XNOR U14860 ( .A(n14326), .B(n14327), .Z(n14329) );
  NANDN U14861 ( .A(n13981), .B(n13980), .Z(n13985) );
  NAND U14862 ( .A(n13983), .B(n13982), .Z(n13984) );
  AND U14863 ( .A(n13985), .B(n13984), .Z(n14328) );
  XNOR U14864 ( .A(n14329), .B(n14328), .Z(n14156) );
  NANDN U14865 ( .A(n13987), .B(n13986), .Z(n13991) );
  NAND U14866 ( .A(n13989), .B(n13988), .Z(n13990) );
  AND U14867 ( .A(n13991), .B(n13990), .Z(n14157) );
  XOR U14868 ( .A(n14156), .B(n14157), .Z(n14158) );
  XNOR U14869 ( .A(n14159), .B(n14158), .Z(n14269) );
  XNOR U14870 ( .A(n14270), .B(n14269), .Z(n14272) );
  XNOR U14871 ( .A(n14271), .B(n14272), .Z(n14375) );
  XNOR U14872 ( .A(n14374), .B(n14375), .Z(n14146) );
  NANDN U14873 ( .A(n13997), .B(n13996), .Z(n14001) );
  NAND U14874 ( .A(n13999), .B(n13998), .Z(n14000) );
  NAND U14875 ( .A(n14001), .B(n14000), .Z(n14393) );
  NANDN U14876 ( .A(n14003), .B(n14002), .Z(n14007) );
  OR U14877 ( .A(n14005), .B(n14004), .Z(n14006) );
  NAND U14878 ( .A(n14007), .B(n14006), .Z(n14391) );
  XNOR U14879 ( .A(b[15]), .B(a[63]), .Z(n14342) );
  OR U14880 ( .A(n14342), .B(n32010), .Z(n14010) );
  NANDN U14881 ( .A(n14008), .B(n32011), .Z(n14009) );
  NAND U14882 ( .A(n14010), .B(n14009), .Z(n14207) );
  XNOR U14883 ( .A(b[25]), .B(n25001), .Z(n14345) );
  NANDN U14884 ( .A(n34219), .B(n14345), .Z(n14013) );
  NAND U14885 ( .A(n34217), .B(n14011), .Z(n14012) );
  NAND U14886 ( .A(n14013), .B(n14012), .Z(n14204) );
  XNOR U14887 ( .A(b[17]), .B(a[61]), .Z(n14348) );
  NANDN U14888 ( .A(n14348), .B(n32543), .Z(n14016) );
  NANDN U14889 ( .A(n14014), .B(n32541), .Z(n14015) );
  AND U14890 ( .A(n14016), .B(n14015), .Z(n14205) );
  XNOR U14891 ( .A(n14204), .B(n14205), .Z(n14206) );
  XNOR U14892 ( .A(n14207), .B(n14206), .Z(n14226) );
  XOR U14893 ( .A(b[39]), .B(n20867), .Z(n14351) );
  NANDN U14894 ( .A(n14351), .B(n36553), .Z(n14019) );
  NANDN U14895 ( .A(n14017), .B(n36643), .Z(n14018) );
  NAND U14896 ( .A(n14019), .B(n14018), .Z(n14201) );
  XOR U14897 ( .A(b[51]), .B(n17960), .Z(n14354) );
  NANDN U14898 ( .A(n14354), .B(n37803), .Z(n14022) );
  NANDN U14899 ( .A(n14020), .B(n37802), .Z(n14021) );
  NAND U14900 ( .A(n14022), .B(n14021), .Z(n14198) );
  XOR U14901 ( .A(b[53]), .B(n16916), .Z(n14357) );
  NANDN U14902 ( .A(n14357), .B(n37940), .Z(n14025) );
  NANDN U14903 ( .A(n14023), .B(n37941), .Z(n14024) );
  AND U14904 ( .A(n14025), .B(n14024), .Z(n14199) );
  XNOR U14905 ( .A(n14198), .B(n14199), .Z(n14200) );
  XOR U14906 ( .A(n14201), .B(n14200), .Z(n14227) );
  XNOR U14907 ( .A(n14226), .B(n14227), .Z(n14228) );
  NANDN U14908 ( .A(n14027), .B(n14026), .Z(n14031) );
  NAND U14909 ( .A(n14029), .B(n14028), .Z(n14030) );
  NAND U14910 ( .A(n14031), .B(n14030), .Z(n14229) );
  XOR U14911 ( .A(n14228), .B(n14229), .Z(n14333) );
  NANDN U14912 ( .A(n14033), .B(n14032), .Z(n14037) );
  NAND U14913 ( .A(n14035), .B(n14034), .Z(n14036) );
  NAND U14914 ( .A(n14037), .B(n14036), .Z(n14330) );
  XNOR U14915 ( .A(n14330), .B(n14331), .Z(n14332) );
  XOR U14916 ( .A(n14333), .B(n14332), .Z(n14390) );
  XNOR U14917 ( .A(n14391), .B(n14390), .Z(n14392) );
  XNOR U14918 ( .A(n14393), .B(n14392), .Z(n14378) );
  XOR U14919 ( .A(b[49]), .B(n18003), .Z(n14290) );
  OR U14920 ( .A(n14290), .B(n37756), .Z(n14044) );
  NANDN U14921 ( .A(n14042), .B(n37652), .Z(n14043) );
  NAND U14922 ( .A(n14044), .B(n14043), .Z(n14322) );
  NAND U14923 ( .A(n37469), .B(n14045), .Z(n14047) );
  XOR U14924 ( .A(n978), .B(n18639), .Z(n14293) );
  NAND U14925 ( .A(n14293), .B(n37471), .Z(n14046) );
  AND U14926 ( .A(n14047), .B(n14046), .Z(n14320) );
  XNOR U14927 ( .A(b[9]), .B(a[69]), .Z(n14296) );
  NANDN U14928 ( .A(n14296), .B(n30509), .Z(n14050) );
  NANDN U14929 ( .A(n14048), .B(n30846), .Z(n14049) );
  AND U14930 ( .A(n14050), .B(n14049), .Z(n14321) );
  XOR U14931 ( .A(n14322), .B(n14323), .Z(n14174) );
  XOR U14932 ( .A(b[11]), .B(n29372), .Z(n14281) );
  OR U14933 ( .A(n14281), .B(n31369), .Z(n14053) );
  NANDN U14934 ( .A(n14051), .B(n31119), .Z(n14052) );
  NAND U14935 ( .A(n14053), .B(n14052), .Z(n14302) );
  XOR U14936 ( .A(b[43]), .B(n20315), .Z(n14284) );
  NANDN U14937 ( .A(n14284), .B(n37068), .Z(n14056) );
  NANDN U14938 ( .A(n14054), .B(n37069), .Z(n14055) );
  NAND U14939 ( .A(n14056), .B(n14055), .Z(n14299) );
  XNOR U14940 ( .A(b[45]), .B(a[33]), .Z(n14287) );
  NANDN U14941 ( .A(n14287), .B(n37261), .Z(n14059) );
  NANDN U14942 ( .A(n14057), .B(n37262), .Z(n14058) );
  AND U14943 ( .A(n14059), .B(n14058), .Z(n14300) );
  XNOR U14944 ( .A(n14299), .B(n14300), .Z(n14301) );
  XOR U14945 ( .A(n14302), .B(n14301), .Z(n14175) );
  XNOR U14946 ( .A(n14174), .B(n14175), .Z(n14176) );
  NANDN U14947 ( .A(n14061), .B(n14060), .Z(n14065) );
  NAND U14948 ( .A(n14063), .B(n14062), .Z(n14064) );
  AND U14949 ( .A(n14065), .B(n14064), .Z(n14177) );
  XNOR U14950 ( .A(n14176), .B(n14177), .Z(n14385) );
  XNOR U14951 ( .A(n14385), .B(n14384), .Z(n14386) );
  XNOR U14952 ( .A(b[35]), .B(a[43]), .Z(n14305) );
  NANDN U14953 ( .A(n14305), .B(n35985), .Z(n14072) );
  NANDN U14954 ( .A(n14070), .B(n35986), .Z(n14071) );
  NAND U14955 ( .A(n14072), .B(n14071), .Z(n14369) );
  XOR U14956 ( .A(n31123), .B(n30543), .Z(n14308) );
  NAND U14957 ( .A(n14308), .B(n29949), .Z(n14075) );
  NAND U14958 ( .A(n29948), .B(n14073), .Z(n14074) );
  NAND U14959 ( .A(n14075), .B(n14074), .Z(n14366) );
  XOR U14960 ( .A(b[55]), .B(n16269), .Z(n14311) );
  NANDN U14961 ( .A(n14311), .B(n38075), .Z(n14078) );
  NANDN U14962 ( .A(n14076), .B(n38073), .Z(n14077) );
  AND U14963 ( .A(n14078), .B(n14077), .Z(n14367) );
  XNOR U14964 ( .A(n14366), .B(n14367), .Z(n14368) );
  XNOR U14965 ( .A(n14369), .B(n14368), .Z(n14153) );
  NANDN U14966 ( .A(n14080), .B(n14079), .Z(n14084) );
  NAND U14967 ( .A(n14082), .B(n14081), .Z(n14083) );
  NAND U14968 ( .A(n14084), .B(n14083), .Z(n14150) );
  NANDN U14969 ( .A(n14086), .B(n14085), .Z(n14090) );
  NAND U14970 ( .A(n14088), .B(n14087), .Z(n14089) );
  NAND U14971 ( .A(n14090), .B(n14089), .Z(n14151) );
  XNOR U14972 ( .A(n14150), .B(n14151), .Z(n14152) );
  XOR U14973 ( .A(n14153), .B(n14152), .Z(n14387) );
  XNOR U14974 ( .A(n14386), .B(n14387), .Z(n14379) );
  XOR U14975 ( .A(n14381), .B(n14380), .Z(n14147) );
  XNOR U14976 ( .A(n14146), .B(n14147), .Z(n14148) );
  XNOR U14977 ( .A(n14149), .B(n14148), .Z(n14401) );
  NANDN U14978 ( .A(n14092), .B(n14091), .Z(n14096) );
  NAND U14979 ( .A(n14094), .B(n14093), .Z(n14095) );
  NAND U14980 ( .A(n14096), .B(n14095), .Z(n14143) );
  NANDN U14981 ( .A(n14102), .B(n14101), .Z(n14106) );
  NAND U14982 ( .A(n14104), .B(n14103), .Z(n14105) );
  AND U14983 ( .A(n14106), .B(n14105), .Z(n14141) );
  XNOR U14984 ( .A(n14140), .B(n14141), .Z(n14142) );
  XOR U14985 ( .A(n14143), .B(n14142), .Z(n14398) );
  XNOR U14986 ( .A(n14398), .B(n14399), .Z(n14400) );
  XNOR U14987 ( .A(n14401), .B(n14400), .Z(n14407) );
  NANDN U14988 ( .A(n14112), .B(n14111), .Z(n14116) );
  NAND U14989 ( .A(n14114), .B(n14113), .Z(n14115) );
  NAND U14990 ( .A(n14116), .B(n14115), .Z(n14404) );
  NANDN U14991 ( .A(n14118), .B(n14117), .Z(n14122) );
  OR U14992 ( .A(n14120), .B(n14119), .Z(n14121) );
  NAND U14993 ( .A(n14122), .B(n14121), .Z(n14405) );
  XNOR U14994 ( .A(n14404), .B(n14405), .Z(n14406) );
  XOR U14995 ( .A(n14407), .B(n14406), .Z(n14410) );
  XNOR U14996 ( .A(n14411), .B(n14410), .Z(n14413) );
  XNOR U14997 ( .A(n14412), .B(n14413), .Z(n14134) );
  NANDN U14998 ( .A(n14124), .B(n14123), .Z(n14128) );
  NAND U14999 ( .A(n14126), .B(n14125), .Z(n14127) );
  AND U15000 ( .A(n14128), .B(n14127), .Z(n14135) );
  XOR U15001 ( .A(n14134), .B(n14135), .Z(n14136) );
  XNOR U15002 ( .A(n14137), .B(n14136), .Z(n14416) );
  XNOR U15003 ( .A(n14416), .B(sreg[141]), .Z(n14418) );
  NAND U15004 ( .A(n14129), .B(sreg[140]), .Z(n14133) );
  OR U15005 ( .A(n14131), .B(n14130), .Z(n14132) );
  AND U15006 ( .A(n14133), .B(n14132), .Z(n14417) );
  XOR U15007 ( .A(n14418), .B(n14417), .Z(c[141]) );
  NAND U15008 ( .A(n14135), .B(n14134), .Z(n14139) );
  NAND U15009 ( .A(n14137), .B(n14136), .Z(n14138) );
  NAND U15010 ( .A(n14139), .B(n14138), .Z(n14424) );
  NANDN U15011 ( .A(n14141), .B(n14140), .Z(n14145) );
  NAND U15012 ( .A(n14143), .B(n14142), .Z(n14144) );
  NAND U15013 ( .A(n14145), .B(n14144), .Z(n14686) );
  XNOR U15014 ( .A(n14686), .B(n14687), .Z(n14688) );
  NANDN U15015 ( .A(n14151), .B(n14150), .Z(n14155) );
  NAND U15016 ( .A(n14153), .B(n14152), .Z(n14154) );
  AND U15017 ( .A(n14155), .B(n14154), .Z(n14679) );
  NAND U15018 ( .A(n14157), .B(n14156), .Z(n14161) );
  NANDN U15019 ( .A(n14159), .B(n14158), .Z(n14160) );
  NAND U15020 ( .A(n14161), .B(n14160), .Z(n14676) );
  NANDN U15021 ( .A(n14163), .B(n14162), .Z(n14167) );
  OR U15022 ( .A(n14165), .B(n14164), .Z(n14166) );
  AND U15023 ( .A(n14167), .B(n14166), .Z(n14677) );
  XNOR U15024 ( .A(n14676), .B(n14677), .Z(n14678) );
  XNOR U15025 ( .A(n14679), .B(n14678), .Z(n14654) );
  NANDN U15026 ( .A(n14169), .B(n14168), .Z(n14173) );
  OR U15027 ( .A(n14171), .B(n14170), .Z(n14172) );
  AND U15028 ( .A(n14173), .B(n14172), .Z(n14655) );
  XNOR U15029 ( .A(n14654), .B(n14655), .Z(n14657) );
  NANDN U15030 ( .A(n14175), .B(n14174), .Z(n14179) );
  NAND U15031 ( .A(n14177), .B(n14176), .Z(n14178) );
  NAND U15032 ( .A(n14179), .B(n14178), .Z(n14456) );
  XOR U15033 ( .A(b[37]), .B(n22246), .Z(n14463) );
  NANDN U15034 ( .A(n14463), .B(n36311), .Z(n14182) );
  NANDN U15035 ( .A(n14180), .B(n36309), .Z(n14181) );
  NAND U15036 ( .A(n14182), .B(n14181), .Z(n14542) );
  XOR U15037 ( .A(a[74]), .B(n968), .Z(n14466) );
  OR U15038 ( .A(n14466), .B(n29363), .Z(n14185) );
  NANDN U15039 ( .A(n14183), .B(n29864), .Z(n14184) );
  NAND U15040 ( .A(n14185), .B(n14184), .Z(n14539) );
  XOR U15041 ( .A(n31363), .B(n967), .Z(n14469) );
  NAND U15042 ( .A(n14469), .B(n28939), .Z(n14188) );
  NAND U15043 ( .A(n28938), .B(n14186), .Z(n14187) );
  AND U15044 ( .A(n14188), .B(n14187), .Z(n14540) );
  XNOR U15045 ( .A(n14539), .B(n14540), .Z(n14541) );
  XNOR U15046 ( .A(n14542), .B(n14541), .Z(n14447) );
  XOR U15047 ( .A(b[13]), .B(n28701), .Z(n14472) );
  OR U15048 ( .A(n14472), .B(n31550), .Z(n14191) );
  NANDN U15049 ( .A(n14189), .B(n31874), .Z(n14190) );
  NAND U15050 ( .A(n14191), .B(n14190), .Z(n14627) );
  NAND U15051 ( .A(n34848), .B(n14192), .Z(n14194) );
  XOR U15052 ( .A(n35375), .B(n25134), .Z(n14475) );
  NAND U15053 ( .A(n34618), .B(n14475), .Z(n14193) );
  NAND U15054 ( .A(n14194), .B(n14193), .Z(n14624) );
  NAND U15055 ( .A(n35188), .B(n14195), .Z(n14197) );
  XOR U15056 ( .A(n35540), .B(n24671), .Z(n14478) );
  NANDN U15057 ( .A(n34968), .B(n14478), .Z(n14196) );
  AND U15058 ( .A(n14197), .B(n14196), .Z(n14625) );
  XNOR U15059 ( .A(n14624), .B(n14625), .Z(n14626) );
  XOR U15060 ( .A(n14627), .B(n14626), .Z(n14448) );
  XNOR U15061 ( .A(n14447), .B(n14448), .Z(n14449) );
  NANDN U15062 ( .A(n14199), .B(n14198), .Z(n14203) );
  NAND U15063 ( .A(n14201), .B(n14200), .Z(n14202) );
  NAND U15064 ( .A(n14203), .B(n14202), .Z(n14450) );
  XOR U15065 ( .A(n14449), .B(n14450), .Z(n14453) );
  NANDN U15066 ( .A(n14205), .B(n14204), .Z(n14209) );
  NAND U15067 ( .A(n14207), .B(n14206), .Z(n14208) );
  NAND U15068 ( .A(n14209), .B(n14208), .Z(n14596) );
  ANDN U15069 ( .B(b[63]), .A(n14210), .Z(n14561) );
  NANDN U15070 ( .A(n14211), .B(n38369), .Z(n14213) );
  XOR U15071 ( .A(b[61]), .B(n14905), .Z(n14493) );
  OR U15072 ( .A(n14493), .B(n38371), .Z(n14212) );
  NAND U15073 ( .A(n14213), .B(n14212), .Z(n14559) );
  NANDN U15074 ( .A(n14214), .B(n35311), .Z(n14216) );
  XOR U15075 ( .A(b[31]), .B(n23447), .Z(n14496) );
  NANDN U15076 ( .A(n14496), .B(n35313), .Z(n14215) );
  AND U15077 ( .A(n14216), .B(n14215), .Z(n14558) );
  XNOR U15078 ( .A(n14559), .B(n14558), .Z(n14560) );
  XOR U15079 ( .A(n14561), .B(n14560), .Z(n14594) );
  NAND U15080 ( .A(n33283), .B(n14217), .Z(n14219) );
  XOR U15081 ( .A(n33020), .B(n27436), .Z(n14499) );
  NANDN U15082 ( .A(n33021), .B(n14499), .Z(n14218) );
  NAND U15083 ( .A(n14219), .B(n14218), .Z(n14530) );
  XNOR U15084 ( .A(b[21]), .B(a[58]), .Z(n14502) );
  OR U15085 ( .A(n14502), .B(n33634), .Z(n14222) );
  NANDN U15086 ( .A(n14220), .B(n33464), .Z(n14221) );
  NAND U15087 ( .A(n14222), .B(n14221), .Z(n14527) );
  NAND U15088 ( .A(n34044), .B(n14223), .Z(n14225) );
  XOR U15089 ( .A(n34510), .B(n25860), .Z(n14505) );
  NANDN U15090 ( .A(n33867), .B(n14505), .Z(n14224) );
  AND U15091 ( .A(n14225), .B(n14224), .Z(n14528) );
  XNOR U15092 ( .A(n14527), .B(n14528), .Z(n14529) );
  XNOR U15093 ( .A(n14530), .B(n14529), .Z(n14595) );
  XOR U15094 ( .A(n14594), .B(n14595), .Z(n14597) );
  XOR U15095 ( .A(n14596), .B(n14597), .Z(n14454) );
  XNOR U15096 ( .A(n14453), .B(n14454), .Z(n14455) );
  XOR U15097 ( .A(n14456), .B(n14455), .Z(n14650) );
  NANDN U15098 ( .A(n14227), .B(n14226), .Z(n14231) );
  NANDN U15099 ( .A(n14229), .B(n14228), .Z(n14230) );
  NAND U15100 ( .A(n14231), .B(n14230), .Z(n14649) );
  NANDN U15101 ( .A(n14233), .B(n14232), .Z(n14237) );
  NAND U15102 ( .A(n14235), .B(n14234), .Z(n14236) );
  NAND U15103 ( .A(n14237), .B(n14236), .Z(n14445) );
  NANDN U15104 ( .A(n14239), .B(n14238), .Z(n14243) );
  NAND U15105 ( .A(n14241), .B(n14240), .Z(n14242) );
  NAND U15106 ( .A(n14243), .B(n14242), .Z(n14645) );
  XNOR U15107 ( .A(b[41]), .B(a[38]), .Z(n14518) );
  OR U15108 ( .A(n14518), .B(n36905), .Z(n14246) );
  NANDN U15109 ( .A(n14244), .B(n36807), .Z(n14245) );
  NAND U15110 ( .A(n14246), .B(n14245), .Z(n14536) );
  XOR U15111 ( .A(b[57]), .B(n15963), .Z(n14521) );
  OR U15112 ( .A(n14521), .B(n965), .Z(n14249) );
  NANDN U15113 ( .A(n14247), .B(n38194), .Z(n14248) );
  NAND U15114 ( .A(n14249), .B(n14248), .Z(n14533) );
  NAND U15115 ( .A(n38326), .B(n14250), .Z(n14252) );
  XOR U15116 ( .A(n38400), .B(n15484), .Z(n14524) );
  NANDN U15117 ( .A(n38273), .B(n14524), .Z(n14251) );
  AND U15118 ( .A(n14252), .B(n14251), .Z(n14534) );
  XNOR U15119 ( .A(n14533), .B(n14534), .Z(n14535) );
  XNOR U15120 ( .A(n14536), .B(n14535), .Z(n14642) );
  XOR U15121 ( .A(b[33]), .B(n22964), .Z(n14508) );
  NANDN U15122 ( .A(n14508), .B(n35620), .Z(n14255) );
  NANDN U15123 ( .A(n14253), .B(n35621), .Z(n14254) );
  NAND U15124 ( .A(n14255), .B(n14254), .Z(n14639) );
  NANDN U15125 ( .A(n966), .B(a[78]), .Z(n14256) );
  XOR U15126 ( .A(n29232), .B(n14256), .Z(n14258) );
  NANDN U15127 ( .A(b[0]), .B(a[77]), .Z(n14257) );
  AND U15128 ( .A(n14258), .B(n14257), .Z(n14636) );
  XOR U15129 ( .A(b[63]), .B(n14259), .Z(n14515) );
  NANDN U15130 ( .A(n14515), .B(n38422), .Z(n14262) );
  NANDN U15131 ( .A(n14260), .B(n38423), .Z(n14261) );
  AND U15132 ( .A(n14262), .B(n14261), .Z(n14637) );
  XNOR U15133 ( .A(n14636), .B(n14637), .Z(n14638) );
  XOR U15134 ( .A(n14639), .B(n14638), .Z(n14643) );
  XNOR U15135 ( .A(n14642), .B(n14643), .Z(n14644) );
  XNOR U15136 ( .A(n14645), .B(n14644), .Z(n14443) );
  NANDN U15137 ( .A(n14264), .B(n14263), .Z(n14268) );
  NAND U15138 ( .A(n14266), .B(n14265), .Z(n14267) );
  AND U15139 ( .A(n14268), .B(n14267), .Z(n14444) );
  XNOR U15140 ( .A(n14443), .B(n14444), .Z(n14446) );
  XOR U15141 ( .A(n14445), .B(n14446), .Z(n14648) );
  XNOR U15142 ( .A(n14649), .B(n14648), .Z(n14651) );
  XNOR U15143 ( .A(n14650), .B(n14651), .Z(n14656) );
  XOR U15144 ( .A(n14657), .B(n14656), .Z(n14431) );
  NAND U15145 ( .A(n14270), .B(n14269), .Z(n14274) );
  NANDN U15146 ( .A(n14272), .B(n14271), .Z(n14273) );
  NAND U15147 ( .A(n14274), .B(n14273), .Z(n14663) );
  OR U15148 ( .A(n14276), .B(n14275), .Z(n14280) );
  OR U15149 ( .A(n14278), .B(n14277), .Z(n14279) );
  NAND U15150 ( .A(n14280), .B(n14279), .Z(n14665) );
  XOR U15151 ( .A(b[11]), .B(n29868), .Z(n14570) );
  OR U15152 ( .A(n14570), .B(n31369), .Z(n14283) );
  NANDN U15153 ( .A(n14281), .B(n31119), .Z(n14282) );
  NAND U15154 ( .A(n14283), .B(n14282), .Z(n14591) );
  XOR U15155 ( .A(b[43]), .B(n19980), .Z(n14573) );
  NANDN U15156 ( .A(n14573), .B(n37068), .Z(n14286) );
  NANDN U15157 ( .A(n14284), .B(n37069), .Z(n14285) );
  NAND U15158 ( .A(n14286), .B(n14285), .Z(n14588) );
  XNOR U15159 ( .A(b[45]), .B(a[34]), .Z(n14576) );
  NANDN U15160 ( .A(n14576), .B(n37261), .Z(n14289) );
  NANDN U15161 ( .A(n14287), .B(n37262), .Z(n14288) );
  AND U15162 ( .A(n14289), .B(n14288), .Z(n14589) );
  XNOR U15163 ( .A(n14588), .B(n14589), .Z(n14590) );
  XNOR U15164 ( .A(n14591), .B(n14590), .Z(n14462) );
  XOR U15165 ( .A(b[49]), .B(n18804), .Z(n14579) );
  OR U15166 ( .A(n14579), .B(n37756), .Z(n14292) );
  NANDN U15167 ( .A(n14290), .B(n37652), .Z(n14291) );
  NAND U15168 ( .A(n14292), .B(n14291), .Z(n14567) );
  NAND U15169 ( .A(n37469), .B(n14293), .Z(n14295) );
  XOR U15170 ( .A(n978), .B(n18841), .Z(n14582) );
  NAND U15171 ( .A(n14582), .B(n37471), .Z(n14294) );
  NAND U15172 ( .A(n14295), .B(n14294), .Z(n14564) );
  XOR U15173 ( .A(b[9]), .B(n30379), .Z(n14585) );
  NANDN U15174 ( .A(n14585), .B(n30509), .Z(n14298) );
  NANDN U15175 ( .A(n14296), .B(n30846), .Z(n14297) );
  AND U15176 ( .A(n14298), .B(n14297), .Z(n14565) );
  XNOR U15177 ( .A(n14564), .B(n14565), .Z(n14566) );
  XNOR U15178 ( .A(n14567), .B(n14566), .Z(n14459) );
  NANDN U15179 ( .A(n14300), .B(n14299), .Z(n14304) );
  NAND U15180 ( .A(n14302), .B(n14301), .Z(n14303) );
  NAND U15181 ( .A(n14304), .B(n14303), .Z(n14460) );
  XNOR U15182 ( .A(n14459), .B(n14460), .Z(n14461) );
  XOR U15183 ( .A(n14462), .B(n14461), .Z(n14664) );
  XNOR U15184 ( .A(n14665), .B(n14664), .Z(n14667) );
  XNOR U15185 ( .A(b[35]), .B(a[44]), .Z(n14549) );
  NANDN U15186 ( .A(n14549), .B(n35985), .Z(n14307) );
  NANDN U15187 ( .A(n14305), .B(n35986), .Z(n14306) );
  NAND U15188 ( .A(n14307), .B(n14306), .Z(n14633) );
  XOR U15189 ( .A(n31123), .B(n30210), .Z(n14552) );
  NAND U15190 ( .A(n14552), .B(n29949), .Z(n14310) );
  NAND U15191 ( .A(n29948), .B(n14308), .Z(n14309) );
  NAND U15192 ( .A(n14310), .B(n14309), .Z(n14630) );
  XOR U15193 ( .A(b[55]), .B(n16508), .Z(n14555) );
  NANDN U15194 ( .A(n14555), .B(n38075), .Z(n14313) );
  NANDN U15195 ( .A(n14311), .B(n38073), .Z(n14312) );
  AND U15196 ( .A(n14313), .B(n14312), .Z(n14631) );
  XNOR U15197 ( .A(n14630), .B(n14631), .Z(n14632) );
  XNOR U15198 ( .A(n14633), .B(n14632), .Z(n14440) );
  NANDN U15199 ( .A(n14315), .B(n14314), .Z(n14319) );
  NAND U15200 ( .A(n14317), .B(n14316), .Z(n14318) );
  NAND U15201 ( .A(n14319), .B(n14318), .Z(n14437) );
  OR U15202 ( .A(n14321), .B(n14320), .Z(n14325) );
  NANDN U15203 ( .A(n14323), .B(n14322), .Z(n14324) );
  NAND U15204 ( .A(n14325), .B(n14324), .Z(n14438) );
  XNOR U15205 ( .A(n14437), .B(n14438), .Z(n14439) );
  XOR U15206 ( .A(n14440), .B(n14439), .Z(n14666) );
  XNOR U15207 ( .A(n14667), .B(n14666), .Z(n14660) );
  NANDN U15208 ( .A(n14331), .B(n14330), .Z(n14335) );
  NAND U15209 ( .A(n14333), .B(n14332), .Z(n14334) );
  NAND U15210 ( .A(n14335), .B(n14334), .Z(n14671) );
  XNOR U15211 ( .A(n14670), .B(n14671), .Z(n14672) );
  NANDN U15212 ( .A(n14337), .B(n14336), .Z(n14341) );
  NAND U15213 ( .A(n14339), .B(n14338), .Z(n14340) );
  NAND U15214 ( .A(n14341), .B(n14340), .Z(n14603) );
  XNOR U15215 ( .A(b[15]), .B(a[64]), .Z(n14606) );
  OR U15216 ( .A(n14606), .B(n32010), .Z(n14344) );
  NANDN U15217 ( .A(n14342), .B(n32011), .Z(n14343) );
  NAND U15218 ( .A(n14344), .B(n14343), .Z(n14490) );
  XNOR U15219 ( .A(b[25]), .B(n25177), .Z(n14609) );
  NANDN U15220 ( .A(n34219), .B(n14609), .Z(n14347) );
  NAND U15221 ( .A(n34217), .B(n14345), .Z(n14346) );
  NAND U15222 ( .A(n14347), .B(n14346), .Z(n14487) );
  XOR U15223 ( .A(b[17]), .B(a[62]), .Z(n14612) );
  NAND U15224 ( .A(n14612), .B(n32543), .Z(n14350) );
  NANDN U15225 ( .A(n14348), .B(n32541), .Z(n14349) );
  AND U15226 ( .A(n14350), .B(n14349), .Z(n14488) );
  XNOR U15227 ( .A(n14487), .B(n14488), .Z(n14489) );
  XNOR U15228 ( .A(n14490), .B(n14489), .Z(n14548) );
  XOR U15229 ( .A(b[39]), .B(n21149), .Z(n14615) );
  NANDN U15230 ( .A(n14615), .B(n36553), .Z(n14353) );
  NANDN U15231 ( .A(n14351), .B(n36643), .Z(n14352) );
  NAND U15232 ( .A(n14353), .B(n14352), .Z(n14484) );
  XOR U15233 ( .A(b[51]), .B(n17702), .Z(n14618) );
  NANDN U15234 ( .A(n14618), .B(n37803), .Z(n14356) );
  NANDN U15235 ( .A(n14354), .B(n37802), .Z(n14355) );
  NAND U15236 ( .A(n14356), .B(n14355), .Z(n14481) );
  XOR U15237 ( .A(b[53]), .B(n17133), .Z(n14621) );
  NANDN U15238 ( .A(n14621), .B(n37940), .Z(n14359) );
  NANDN U15239 ( .A(n14357), .B(n37941), .Z(n14358) );
  AND U15240 ( .A(n14359), .B(n14358), .Z(n14482) );
  XNOR U15241 ( .A(n14481), .B(n14482), .Z(n14483) );
  XNOR U15242 ( .A(n14484), .B(n14483), .Z(n14545) );
  NANDN U15243 ( .A(n14361), .B(n14360), .Z(n14365) );
  NAND U15244 ( .A(n14363), .B(n14362), .Z(n14364) );
  NAND U15245 ( .A(n14365), .B(n14364), .Z(n14546) );
  XNOR U15246 ( .A(n14545), .B(n14546), .Z(n14547) );
  XOR U15247 ( .A(n14548), .B(n14547), .Z(n14600) );
  NANDN U15248 ( .A(n14367), .B(n14366), .Z(n14371) );
  NAND U15249 ( .A(n14369), .B(n14368), .Z(n14370) );
  AND U15250 ( .A(n14371), .B(n14370), .Z(n14601) );
  XOR U15251 ( .A(n14600), .B(n14601), .Z(n14602) );
  XOR U15252 ( .A(n14603), .B(n14602), .Z(n14673) );
  XNOR U15253 ( .A(n14672), .B(n14673), .Z(n14661) );
  XOR U15254 ( .A(n14660), .B(n14661), .Z(n14662) );
  XOR U15255 ( .A(n14663), .B(n14662), .Z(n14432) );
  XNOR U15256 ( .A(n14431), .B(n14432), .Z(n14433) );
  OR U15257 ( .A(n14373), .B(n14372), .Z(n14377) );
  NAND U15258 ( .A(n14375), .B(n14374), .Z(n14376) );
  NAND U15259 ( .A(n14377), .B(n14376), .Z(n14434) );
  XOR U15260 ( .A(n14433), .B(n14434), .Z(n14683) );
  NANDN U15261 ( .A(n14379), .B(n14378), .Z(n14383) );
  NAND U15262 ( .A(n14381), .B(n14380), .Z(n14382) );
  AND U15263 ( .A(n14383), .B(n14382), .Z(n14680) );
  NANDN U15264 ( .A(n14385), .B(n14384), .Z(n14389) );
  NAND U15265 ( .A(n14387), .B(n14386), .Z(n14388) );
  NAND U15266 ( .A(n14389), .B(n14388), .Z(n14428) );
  XNOR U15267 ( .A(n14426), .B(n14425), .Z(n14427) );
  XNOR U15268 ( .A(n14428), .B(n14427), .Z(n14681) );
  XNOR U15269 ( .A(n14683), .B(n14682), .Z(n14689) );
  XOR U15270 ( .A(n14688), .B(n14689), .Z(n14695) );
  OR U15271 ( .A(n14399), .B(n14398), .Z(n14403) );
  OR U15272 ( .A(n14401), .B(n14400), .Z(n14402) );
  NAND U15273 ( .A(n14403), .B(n14402), .Z(n14692) );
  NANDN U15274 ( .A(n14405), .B(n14404), .Z(n14409) );
  NAND U15275 ( .A(n14407), .B(n14406), .Z(n14408) );
  NAND U15276 ( .A(n14409), .B(n14408), .Z(n14693) );
  XNOR U15277 ( .A(n14692), .B(n14693), .Z(n14694) );
  XNOR U15278 ( .A(n14695), .B(n14694), .Z(n14421) );
  NAND U15279 ( .A(n14411), .B(n14410), .Z(n14415) );
  NANDN U15280 ( .A(n14413), .B(n14412), .Z(n14414) );
  AND U15281 ( .A(n14415), .B(n14414), .Z(n14422) );
  XNOR U15282 ( .A(n14421), .B(n14422), .Z(n14423) );
  XNOR U15283 ( .A(n14424), .B(n14423), .Z(n14698) );
  XNOR U15284 ( .A(n14698), .B(sreg[142]), .Z(n14700) );
  NAND U15285 ( .A(n14416), .B(sreg[141]), .Z(n14420) );
  OR U15286 ( .A(n14418), .B(n14417), .Z(n14419) );
  AND U15287 ( .A(n14420), .B(n14419), .Z(n14699) );
  XOR U15288 ( .A(n14700), .B(n14699), .Z(c[142]) );
  NANDN U15289 ( .A(n14426), .B(n14425), .Z(n14430) );
  NAND U15290 ( .A(n14428), .B(n14427), .Z(n14429) );
  NAND U15291 ( .A(n14430), .B(n14429), .Z(n14972) );
  NANDN U15292 ( .A(n14432), .B(n14431), .Z(n14436) );
  NANDN U15293 ( .A(n14434), .B(n14433), .Z(n14435) );
  NAND U15294 ( .A(n14436), .B(n14435), .Z(n14973) );
  XNOR U15295 ( .A(n14972), .B(n14973), .Z(n14974) );
  NANDN U15296 ( .A(n14438), .B(n14437), .Z(n14442) );
  NAND U15297 ( .A(n14440), .B(n14439), .Z(n14441) );
  NAND U15298 ( .A(n14442), .B(n14441), .Z(n14951) );
  NANDN U15299 ( .A(n14448), .B(n14447), .Z(n14452) );
  NANDN U15300 ( .A(n14450), .B(n14449), .Z(n14451) );
  AND U15301 ( .A(n14452), .B(n14451), .Z(n14949) );
  XNOR U15302 ( .A(n14951), .B(n14950), .Z(n14708) );
  NANDN U15303 ( .A(n14454), .B(n14453), .Z(n14458) );
  NANDN U15304 ( .A(n14456), .B(n14455), .Z(n14457) );
  AND U15305 ( .A(n14458), .B(n14457), .Z(n14707) );
  XNOR U15306 ( .A(n14708), .B(n14707), .Z(n14709) );
  XOR U15307 ( .A(b[37]), .B(n21996), .Z(n14872) );
  NANDN U15308 ( .A(n14872), .B(n36311), .Z(n14465) );
  NANDN U15309 ( .A(n14463), .B(n36309), .Z(n14464) );
  NAND U15310 ( .A(n14465), .B(n14464), .Z(n14896) );
  XNOR U15311 ( .A(a[75]), .B(b[5]), .Z(n14875) );
  OR U15312 ( .A(n14875), .B(n29363), .Z(n14468) );
  NANDN U15313 ( .A(n14466), .B(n29864), .Z(n14467) );
  NAND U15314 ( .A(n14468), .B(n14467), .Z(n14893) );
  XNOR U15315 ( .A(a[77]), .B(n967), .Z(n14878) );
  NAND U15316 ( .A(n14878), .B(n28939), .Z(n14471) );
  NAND U15317 ( .A(n28938), .B(n14469), .Z(n14470) );
  AND U15318 ( .A(n14471), .B(n14470), .Z(n14894) );
  XNOR U15319 ( .A(n14893), .B(n14894), .Z(n14895) );
  XNOR U15320 ( .A(n14896), .B(n14895), .Z(n14814) );
  XOR U15321 ( .A(b[13]), .B(n29372), .Z(n14863) );
  OR U15322 ( .A(n14863), .B(n31550), .Z(n14474) );
  NANDN U15323 ( .A(n14472), .B(n31874), .Z(n14473) );
  NAND U15324 ( .A(n14474), .B(n14473), .Z(n14746) );
  NAND U15325 ( .A(n34848), .B(n14475), .Z(n14477) );
  XOR U15326 ( .A(n35375), .B(n25001), .Z(n14866) );
  NAND U15327 ( .A(n34618), .B(n14866), .Z(n14476) );
  NAND U15328 ( .A(n14477), .B(n14476), .Z(n14743) );
  NAND U15329 ( .A(n35188), .B(n14478), .Z(n14480) );
  XOR U15330 ( .A(n35540), .B(n24288), .Z(n14869) );
  NANDN U15331 ( .A(n34968), .B(n14869), .Z(n14479) );
  AND U15332 ( .A(n14480), .B(n14479), .Z(n14744) );
  XNOR U15333 ( .A(n14743), .B(n14744), .Z(n14745) );
  XOR U15334 ( .A(n14746), .B(n14745), .Z(n14815) );
  XOR U15335 ( .A(n14814), .B(n14815), .Z(n14817) );
  NANDN U15336 ( .A(n14482), .B(n14481), .Z(n14486) );
  NAND U15337 ( .A(n14484), .B(n14483), .Z(n14485) );
  NAND U15338 ( .A(n14486), .B(n14485), .Z(n14816) );
  XNOR U15339 ( .A(n14817), .B(n14816), .Z(n14833) );
  NANDN U15340 ( .A(n14488), .B(n14487), .Z(n14492) );
  NAND U15341 ( .A(n14490), .B(n14489), .Z(n14491) );
  NAND U15342 ( .A(n14492), .B(n14491), .Z(n14791) );
  NAND U15343 ( .A(a[15]), .B(b[63]), .Z(n14805) );
  NANDN U15344 ( .A(n14493), .B(n38369), .Z(n14495) );
  XOR U15345 ( .A(b[61]), .B(n15113), .Z(n14857) );
  OR U15346 ( .A(n14857), .B(n38371), .Z(n14494) );
  NAND U15347 ( .A(n14495), .B(n14494), .Z(n14803) );
  NANDN U15348 ( .A(n14496), .B(n35311), .Z(n14498) );
  XOR U15349 ( .A(b[31]), .B(n23852), .Z(n14860) );
  NANDN U15350 ( .A(n14860), .B(n35313), .Z(n14497) );
  AND U15351 ( .A(n14498), .B(n14497), .Z(n14802) );
  XNOR U15352 ( .A(n14803), .B(n14802), .Z(n14804) );
  XOR U15353 ( .A(n14805), .B(n14804), .Z(n14789) );
  NAND U15354 ( .A(n33283), .B(n14499), .Z(n14501) );
  XOR U15355 ( .A(n33020), .B(n27773), .Z(n14842) );
  NANDN U15356 ( .A(n33021), .B(n14842), .Z(n14500) );
  NAND U15357 ( .A(n14501), .B(n14500), .Z(n14921) );
  XOR U15358 ( .A(b[21]), .B(a[59]), .Z(n14845) );
  NANDN U15359 ( .A(n33634), .B(n14845), .Z(n14504) );
  NANDN U15360 ( .A(n14502), .B(n33464), .Z(n14503) );
  NAND U15361 ( .A(n14504), .B(n14503), .Z(n14918) );
  NAND U15362 ( .A(n34044), .B(n14505), .Z(n14507) );
  XOR U15363 ( .A(n34510), .B(n26122), .Z(n14848) );
  NANDN U15364 ( .A(n33867), .B(n14848), .Z(n14506) );
  AND U15365 ( .A(n14507), .B(n14506), .Z(n14919) );
  XNOR U15366 ( .A(n14918), .B(n14919), .Z(n14920) );
  XNOR U15367 ( .A(n14921), .B(n14920), .Z(n14790) );
  XNOR U15368 ( .A(n14789), .B(n14790), .Z(n14792) );
  XNOR U15369 ( .A(n14791), .B(n14792), .Z(n14832) );
  XNOR U15370 ( .A(n14833), .B(n14832), .Z(n14834) );
  XNOR U15371 ( .A(n14835), .B(n14834), .Z(n14716) );
  XOR U15372 ( .A(b[33]), .B(n23149), .Z(n14899) );
  NANDN U15373 ( .A(n14899), .B(n35620), .Z(n14510) );
  NANDN U15374 ( .A(n14508), .B(n35621), .Z(n14509) );
  NAND U15375 ( .A(n14510), .B(n14509), .Z(n14758) );
  NANDN U15376 ( .A(n966), .B(a[79]), .Z(n14511) );
  XOR U15377 ( .A(n29232), .B(n14511), .Z(n14513) );
  IV U15378 ( .A(a[78]), .Z(n31870) );
  NANDN U15379 ( .A(n31870), .B(n966), .Z(n14512) );
  AND U15380 ( .A(n14513), .B(n14512), .Z(n14755) );
  XOR U15381 ( .A(b[63]), .B(n14514), .Z(n14906) );
  NANDN U15382 ( .A(n14906), .B(n38422), .Z(n14517) );
  NANDN U15383 ( .A(n14515), .B(n38423), .Z(n14516) );
  AND U15384 ( .A(n14517), .B(n14516), .Z(n14756) );
  XNOR U15385 ( .A(n14755), .B(n14756), .Z(n14757) );
  XNOR U15386 ( .A(n14758), .B(n14757), .Z(n14761) );
  XNOR U15387 ( .A(b[41]), .B(a[39]), .Z(n14909) );
  OR U15388 ( .A(n14909), .B(n36905), .Z(n14520) );
  NANDN U15389 ( .A(n14518), .B(n36807), .Z(n14519) );
  NAND U15390 ( .A(n14520), .B(n14519), .Z(n14927) );
  XOR U15391 ( .A(b[57]), .B(n16269), .Z(n14912) );
  OR U15392 ( .A(n14912), .B(n965), .Z(n14523) );
  NANDN U15393 ( .A(n14521), .B(n38194), .Z(n14522) );
  NAND U15394 ( .A(n14523), .B(n14522), .Z(n14924) );
  NAND U15395 ( .A(n38326), .B(n14524), .Z(n14526) );
  XOR U15396 ( .A(n38400), .B(n16220), .Z(n14915) );
  NANDN U15397 ( .A(n38273), .B(n14915), .Z(n14525) );
  AND U15398 ( .A(n14526), .B(n14525), .Z(n14925) );
  XNOR U15399 ( .A(n14924), .B(n14925), .Z(n14926) );
  XOR U15400 ( .A(n14927), .B(n14926), .Z(n14760) );
  NANDN U15401 ( .A(n14528), .B(n14527), .Z(n14532) );
  NAND U15402 ( .A(n14530), .B(n14529), .Z(n14531) );
  NAND U15403 ( .A(n14532), .B(n14531), .Z(n14759) );
  XNOR U15404 ( .A(n14760), .B(n14759), .Z(n14762) );
  XNOR U15405 ( .A(n14761), .B(n14762), .Z(n14829) );
  NANDN U15406 ( .A(n14534), .B(n14533), .Z(n14538) );
  NAND U15407 ( .A(n14536), .B(n14535), .Z(n14537) );
  NAND U15408 ( .A(n14538), .B(n14537), .Z(n14826) );
  NANDN U15409 ( .A(n14540), .B(n14539), .Z(n14544) );
  NAND U15410 ( .A(n14542), .B(n14541), .Z(n14543) );
  AND U15411 ( .A(n14544), .B(n14543), .Z(n14827) );
  XNOR U15412 ( .A(n14826), .B(n14827), .Z(n14828) );
  XNOR U15413 ( .A(n14829), .B(n14828), .Z(n14714) );
  XOR U15414 ( .A(n14714), .B(n14713), .Z(n14715) );
  XNOR U15415 ( .A(n14716), .B(n14715), .Z(n14710) );
  XOR U15416 ( .A(n14709), .B(n14710), .Z(n14960) );
  XNOR U15417 ( .A(b[35]), .B(a[45]), .Z(n14793) );
  NANDN U15418 ( .A(n14793), .B(n35985), .Z(n14551) );
  NANDN U15419 ( .A(n14549), .B(n35986), .Z(n14550) );
  NAND U15420 ( .A(n14551), .B(n14550), .Z(n14752) );
  XNOR U15421 ( .A(n31123), .B(a[73]), .Z(n14796) );
  NAND U15422 ( .A(n14796), .B(n29949), .Z(n14554) );
  NAND U15423 ( .A(n29948), .B(n14552), .Z(n14553) );
  NAND U15424 ( .A(n14554), .B(n14553), .Z(n14749) );
  XOR U15425 ( .A(b[55]), .B(n16916), .Z(n14799) );
  NANDN U15426 ( .A(n14799), .B(n38075), .Z(n14557) );
  NANDN U15427 ( .A(n14555), .B(n38073), .Z(n14556) );
  AND U15428 ( .A(n14557), .B(n14556), .Z(n14750) );
  XNOR U15429 ( .A(n14749), .B(n14750), .Z(n14751) );
  XNOR U15430 ( .A(n14752), .B(n14751), .Z(n14823) );
  NANDN U15431 ( .A(n14559), .B(n14558), .Z(n14563) );
  NANDN U15432 ( .A(n14561), .B(n14560), .Z(n14562) );
  NAND U15433 ( .A(n14563), .B(n14562), .Z(n14820) );
  NANDN U15434 ( .A(n14565), .B(n14564), .Z(n14569) );
  NAND U15435 ( .A(n14567), .B(n14566), .Z(n14568) );
  NAND U15436 ( .A(n14569), .B(n14568), .Z(n14821) );
  XNOR U15437 ( .A(n14820), .B(n14821), .Z(n14822) );
  XOR U15438 ( .A(n14823), .B(n14822), .Z(n14938) );
  XNOR U15439 ( .A(b[11]), .B(a[69]), .Z(n14765) );
  OR U15440 ( .A(n14765), .B(n31369), .Z(n14572) );
  NANDN U15441 ( .A(n14570), .B(n31119), .Z(n14571) );
  NAND U15442 ( .A(n14572), .B(n14571), .Z(n14786) );
  XOR U15443 ( .A(b[43]), .B(n20352), .Z(n14768) );
  NANDN U15444 ( .A(n14768), .B(n37068), .Z(n14575) );
  NANDN U15445 ( .A(n14573), .B(n37069), .Z(n14574) );
  NAND U15446 ( .A(n14575), .B(n14574), .Z(n14783) );
  XNOR U15447 ( .A(b[45]), .B(a[35]), .Z(n14771) );
  NANDN U15448 ( .A(n14771), .B(n37261), .Z(n14578) );
  NANDN U15449 ( .A(n14576), .B(n37262), .Z(n14577) );
  AND U15450 ( .A(n14578), .B(n14577), .Z(n14784) );
  XNOR U15451 ( .A(n14783), .B(n14784), .Z(n14785) );
  XNOR U15452 ( .A(n14786), .B(n14785), .Z(n14841) );
  XOR U15453 ( .A(b[49]), .B(n18639), .Z(n14774) );
  OR U15454 ( .A(n14774), .B(n37756), .Z(n14581) );
  NANDN U15455 ( .A(n14579), .B(n37652), .Z(n14580) );
  NAND U15456 ( .A(n14581), .B(n14580), .Z(n14811) );
  NAND U15457 ( .A(n37469), .B(n14582), .Z(n14584) );
  XOR U15458 ( .A(n978), .B(n19656), .Z(n14777) );
  NAND U15459 ( .A(n14777), .B(n37471), .Z(n14583) );
  NAND U15460 ( .A(n14584), .B(n14583), .Z(n14808) );
  XOR U15461 ( .A(b[9]), .B(n30543), .Z(n14780) );
  NANDN U15462 ( .A(n14780), .B(n30509), .Z(n14587) );
  NANDN U15463 ( .A(n14585), .B(n30846), .Z(n14586) );
  AND U15464 ( .A(n14587), .B(n14586), .Z(n14809) );
  XNOR U15465 ( .A(n14808), .B(n14809), .Z(n14810) );
  XNOR U15466 ( .A(n14811), .B(n14810), .Z(n14838) );
  NANDN U15467 ( .A(n14589), .B(n14588), .Z(n14593) );
  NAND U15468 ( .A(n14591), .B(n14590), .Z(n14592) );
  NAND U15469 ( .A(n14593), .B(n14592), .Z(n14839) );
  XNOR U15470 ( .A(n14838), .B(n14839), .Z(n14840) );
  XOR U15471 ( .A(n14841), .B(n14840), .Z(n14936) );
  NANDN U15472 ( .A(n14595), .B(n14594), .Z(n14599) );
  NANDN U15473 ( .A(n14597), .B(n14596), .Z(n14598) );
  AND U15474 ( .A(n14599), .B(n14598), .Z(n14937) );
  XNOR U15475 ( .A(n14936), .B(n14937), .Z(n14939) );
  XNOR U15476 ( .A(n14938), .B(n14939), .Z(n14930) );
  NAND U15477 ( .A(n14601), .B(n14600), .Z(n14605) );
  NANDN U15478 ( .A(n14603), .B(n14602), .Z(n14604) );
  NAND U15479 ( .A(n14605), .B(n14604), .Z(n14945) );
  XOR U15480 ( .A(b[15]), .B(n28403), .Z(n14734) );
  OR U15481 ( .A(n14734), .B(n32010), .Z(n14608) );
  NANDN U15482 ( .A(n14606), .B(n32011), .Z(n14607) );
  NAND U15483 ( .A(n14608), .B(n14607), .Z(n14854) );
  XNOR U15484 ( .A(b[25]), .B(n25466), .Z(n14737) );
  NANDN U15485 ( .A(n34219), .B(n14737), .Z(n14611) );
  NAND U15486 ( .A(n34217), .B(n14609), .Z(n14610) );
  NAND U15487 ( .A(n14611), .B(n14610), .Z(n14851) );
  XOR U15488 ( .A(b[17]), .B(a[63]), .Z(n14740) );
  NAND U15489 ( .A(n14740), .B(n32543), .Z(n14614) );
  NAND U15490 ( .A(n14612), .B(n32541), .Z(n14613) );
  AND U15491 ( .A(n14614), .B(n14613), .Z(n14852) );
  XNOR U15492 ( .A(n14851), .B(n14852), .Z(n14853) );
  XNOR U15493 ( .A(n14854), .B(n14853), .Z(n14887) );
  XOR U15494 ( .A(b[39]), .B(n21441), .Z(n14725) );
  NANDN U15495 ( .A(n14725), .B(n36553), .Z(n14617) );
  NANDN U15496 ( .A(n14615), .B(n36643), .Z(n14616) );
  NAND U15497 ( .A(n14617), .B(n14616), .Z(n14884) );
  XOR U15498 ( .A(b[51]), .B(n18003), .Z(n14728) );
  NANDN U15499 ( .A(n14728), .B(n37803), .Z(n14620) );
  NANDN U15500 ( .A(n14618), .B(n37802), .Z(n14619) );
  NAND U15501 ( .A(n14620), .B(n14619), .Z(n14881) );
  XOR U15502 ( .A(b[53]), .B(n17960), .Z(n14731) );
  NANDN U15503 ( .A(n14731), .B(n37940), .Z(n14623) );
  NANDN U15504 ( .A(n14621), .B(n37941), .Z(n14622) );
  AND U15505 ( .A(n14623), .B(n14622), .Z(n14882) );
  XNOR U15506 ( .A(n14881), .B(n14882), .Z(n14883) );
  XOR U15507 ( .A(n14884), .B(n14883), .Z(n14888) );
  XNOR U15508 ( .A(n14887), .B(n14888), .Z(n14889) );
  NANDN U15509 ( .A(n14625), .B(n14624), .Z(n14629) );
  NAND U15510 ( .A(n14627), .B(n14626), .Z(n14628) );
  NAND U15511 ( .A(n14629), .B(n14628), .Z(n14890) );
  XOR U15512 ( .A(n14889), .B(n14890), .Z(n14722) );
  NANDN U15513 ( .A(n14631), .B(n14630), .Z(n14635) );
  NAND U15514 ( .A(n14633), .B(n14632), .Z(n14634) );
  NAND U15515 ( .A(n14635), .B(n14634), .Z(n14719) );
  NANDN U15516 ( .A(n14637), .B(n14636), .Z(n14641) );
  NAND U15517 ( .A(n14639), .B(n14638), .Z(n14640) );
  AND U15518 ( .A(n14641), .B(n14640), .Z(n14720) );
  XNOR U15519 ( .A(n14719), .B(n14720), .Z(n14721) );
  XNOR U15520 ( .A(n14722), .B(n14721), .Z(n14942) );
  NANDN U15521 ( .A(n14643), .B(n14642), .Z(n14647) );
  NANDN U15522 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U15523 ( .A(n14647), .B(n14646), .Z(n14943) );
  XNOR U15524 ( .A(n14942), .B(n14943), .Z(n14944) );
  XOR U15525 ( .A(n14945), .B(n14944), .Z(n14931) );
  NAND U15526 ( .A(n14649), .B(n14648), .Z(n14653) );
  NANDN U15527 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U15528 ( .A(n14653), .B(n14652), .Z(n14933) );
  XNOR U15529 ( .A(n14932), .B(n14933), .Z(n14961) );
  XNOR U15530 ( .A(n14960), .B(n14961), .Z(n14962) );
  NAND U15531 ( .A(n14655), .B(n14654), .Z(n14659) );
  NANDN U15532 ( .A(n14657), .B(n14656), .Z(n14658) );
  NAND U15533 ( .A(n14659), .B(n14658), .Z(n14963) );
  XOR U15534 ( .A(n14962), .B(n14963), .Z(n14969) );
  NAND U15535 ( .A(n14665), .B(n14664), .Z(n14669) );
  NANDN U15536 ( .A(n14667), .B(n14666), .Z(n14668) );
  NAND U15537 ( .A(n14669), .B(n14668), .Z(n14957) );
  NANDN U15538 ( .A(n14671), .B(n14670), .Z(n14675) );
  NANDN U15539 ( .A(n14673), .B(n14672), .Z(n14674) );
  NAND U15540 ( .A(n14675), .B(n14674), .Z(n14954) );
  XNOR U15541 ( .A(n14954), .B(n14955), .Z(n14956) );
  XNOR U15542 ( .A(n14957), .B(n14956), .Z(n14967) );
  XNOR U15543 ( .A(n14966), .B(n14967), .Z(n14968) );
  XNOR U15544 ( .A(n14969), .B(n14968), .Z(n14975) );
  XOR U15545 ( .A(n14974), .B(n14975), .Z(n14981) );
  OR U15546 ( .A(n14681), .B(n14680), .Z(n14685) );
  NAND U15547 ( .A(n14683), .B(n14682), .Z(n14684) );
  NAND U15548 ( .A(n14685), .B(n14684), .Z(n14979) );
  NANDN U15549 ( .A(n14687), .B(n14686), .Z(n14691) );
  NANDN U15550 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15551 ( .A(n14691), .B(n14690), .Z(n14978) );
  XNOR U15552 ( .A(n14979), .B(n14978), .Z(n14980) );
  XNOR U15553 ( .A(n14981), .B(n14980), .Z(n14703) );
  NANDN U15554 ( .A(n14693), .B(n14692), .Z(n14697) );
  NAND U15555 ( .A(n14695), .B(n14694), .Z(n14696) );
  NAND U15556 ( .A(n14697), .B(n14696), .Z(n14704) );
  XNOR U15557 ( .A(n14703), .B(n14704), .Z(n14705) );
  XNOR U15558 ( .A(n14706), .B(n14705), .Z(n14984) );
  XNOR U15559 ( .A(n14984), .B(sreg[143]), .Z(n14986) );
  NAND U15560 ( .A(n14698), .B(sreg[142]), .Z(n14702) );
  OR U15561 ( .A(n14700), .B(n14699), .Z(n14701) );
  AND U15562 ( .A(n14702), .B(n14701), .Z(n14985) );
  XOR U15563 ( .A(n14986), .B(n14985), .Z(c[143]) );
  NANDN U15564 ( .A(n14708), .B(n14707), .Z(n14712) );
  NANDN U15565 ( .A(n14710), .B(n14709), .Z(n14711) );
  NAND U15566 ( .A(n14712), .B(n14711), .Z(n15010) );
  OR U15567 ( .A(n14714), .B(n14713), .Z(n14718) );
  NAND U15568 ( .A(n14716), .B(n14715), .Z(n14717) );
  NAND U15569 ( .A(n14718), .B(n14717), .Z(n15247) );
  NANDN U15570 ( .A(n14720), .B(n14719), .Z(n14724) );
  NAND U15571 ( .A(n14722), .B(n14721), .Z(n14723) );
  NAND U15572 ( .A(n14724), .B(n14723), .Z(n15261) );
  XOR U15573 ( .A(b[39]), .B(n22246), .Z(n15195) );
  NANDN U15574 ( .A(n15195), .B(n36553), .Z(n14727) );
  NANDN U15575 ( .A(n14725), .B(n36643), .Z(n14726) );
  NAND U15576 ( .A(n14727), .B(n14726), .Z(n15089) );
  XOR U15577 ( .A(b[51]), .B(n18804), .Z(n15198) );
  NANDN U15578 ( .A(n15198), .B(n37803), .Z(n14730) );
  NANDN U15579 ( .A(n14728), .B(n37802), .Z(n14729) );
  NAND U15580 ( .A(n14730), .B(n14729), .Z(n15086) );
  XOR U15581 ( .A(b[53]), .B(n17702), .Z(n15201) );
  NANDN U15582 ( .A(n15201), .B(n37940), .Z(n14733) );
  NANDN U15583 ( .A(n14731), .B(n37941), .Z(n14732) );
  AND U15584 ( .A(n14733), .B(n14732), .Z(n15087) );
  XNOR U15585 ( .A(n15086), .B(n15087), .Z(n15088) );
  XNOR U15586 ( .A(n15089), .B(n15088), .Z(n15132) );
  XOR U15587 ( .A(b[15]), .B(n28701), .Z(n15186) );
  OR U15588 ( .A(n15186), .B(n32010), .Z(n14736) );
  NANDN U15589 ( .A(n14734), .B(n32011), .Z(n14735) );
  NAND U15590 ( .A(n14736), .B(n14735), .Z(n15059) );
  XNOR U15591 ( .A(b[25]), .B(n25860), .Z(n15189) );
  NANDN U15592 ( .A(n34219), .B(n15189), .Z(n14739) );
  NAND U15593 ( .A(n34217), .B(n14737), .Z(n14738) );
  NAND U15594 ( .A(n14739), .B(n14738), .Z(n15056) );
  XOR U15595 ( .A(b[17]), .B(a[64]), .Z(n15192) );
  NAND U15596 ( .A(n15192), .B(n32543), .Z(n14742) );
  NAND U15597 ( .A(n14740), .B(n32541), .Z(n14741) );
  AND U15598 ( .A(n14742), .B(n14741), .Z(n15057) );
  XNOR U15599 ( .A(n15056), .B(n15057), .Z(n15058) );
  XNOR U15600 ( .A(n15059), .B(n15058), .Z(n15129) );
  NANDN U15601 ( .A(n14744), .B(n14743), .Z(n14748) );
  NAND U15602 ( .A(n14746), .B(n14745), .Z(n14747) );
  NAND U15603 ( .A(n14748), .B(n14747), .Z(n15130) );
  XNOR U15604 ( .A(n15129), .B(n15130), .Z(n15131) );
  XOR U15605 ( .A(n15132), .B(n15131), .Z(n15229) );
  NANDN U15606 ( .A(n14750), .B(n14749), .Z(n14754) );
  NAND U15607 ( .A(n14752), .B(n14751), .Z(n14753) );
  NAND U15608 ( .A(n14754), .B(n14753), .Z(n15226) );
  XNOR U15609 ( .A(n15226), .B(n15227), .Z(n15228) );
  XNOR U15610 ( .A(n15229), .B(n15228), .Z(n15258) );
  OR U15611 ( .A(n14760), .B(n14759), .Z(n14764) );
  NANDN U15612 ( .A(n14762), .B(n14761), .Z(n14763) );
  AND U15613 ( .A(n14764), .B(n14763), .Z(n15259) );
  XOR U15614 ( .A(n15258), .B(n15259), .Z(n15260) );
  XNOR U15615 ( .A(n15261), .B(n15260), .Z(n15245) );
  XOR U15616 ( .A(b[11]), .B(n30379), .Z(n15162) );
  OR U15617 ( .A(n15162), .B(n31369), .Z(n14767) );
  NANDN U15618 ( .A(n14765), .B(n31119), .Z(n14766) );
  NAND U15619 ( .A(n14767), .B(n14766), .Z(n15183) );
  XOR U15620 ( .A(b[43]), .B(n20686), .Z(n15165) );
  NANDN U15621 ( .A(n15165), .B(n37068), .Z(n14770) );
  NANDN U15622 ( .A(n14768), .B(n37069), .Z(n14769) );
  NAND U15623 ( .A(n14770), .B(n14769), .Z(n15180) );
  XNOR U15624 ( .A(b[45]), .B(a[36]), .Z(n15168) );
  NANDN U15625 ( .A(n15168), .B(n37261), .Z(n14773) );
  NANDN U15626 ( .A(n14771), .B(n37262), .Z(n14772) );
  AND U15627 ( .A(n14773), .B(n14772), .Z(n15181) );
  XNOR U15628 ( .A(n15180), .B(n15181), .Z(n15182) );
  XNOR U15629 ( .A(n15183), .B(n15182), .Z(n15046) );
  XOR U15630 ( .A(n979), .B(n18841), .Z(n15171) );
  NANDN U15631 ( .A(n37756), .B(n15171), .Z(n14776) );
  NANDN U15632 ( .A(n14774), .B(n37652), .Z(n14775) );
  NAND U15633 ( .A(n14776), .B(n14775), .Z(n15153) );
  NAND U15634 ( .A(n37469), .B(n14777), .Z(n14779) );
  XOR U15635 ( .A(b[47]), .B(n19513), .Z(n15174) );
  NANDN U15636 ( .A(n15174), .B(n37471), .Z(n14778) );
  NAND U15637 ( .A(n14779), .B(n14778), .Z(n15150) );
  XOR U15638 ( .A(n969), .B(n30210), .Z(n15177) );
  NAND U15639 ( .A(n30509), .B(n15177), .Z(n14782) );
  NANDN U15640 ( .A(n14780), .B(n30846), .Z(n14781) );
  AND U15641 ( .A(n14782), .B(n14781), .Z(n15151) );
  XNOR U15642 ( .A(n15150), .B(n15151), .Z(n15152) );
  XNOR U15643 ( .A(n15153), .B(n15152), .Z(n15043) );
  NANDN U15644 ( .A(n14784), .B(n14783), .Z(n14788) );
  NAND U15645 ( .A(n14786), .B(n14785), .Z(n14787) );
  NAND U15646 ( .A(n14788), .B(n14787), .Z(n15044) );
  XNOR U15647 ( .A(n15043), .B(n15044), .Z(n15045) );
  XOR U15648 ( .A(n15046), .B(n15045), .Z(n15248) );
  XNOR U15649 ( .A(n15248), .B(n15249), .Z(n15251) );
  XNOR U15650 ( .A(b[35]), .B(a[46]), .Z(n15135) );
  NANDN U15651 ( .A(n15135), .B(n35985), .Z(n14795) );
  NANDN U15652 ( .A(n14793), .B(n35986), .Z(n14794) );
  NAND U15653 ( .A(n14795), .B(n14794), .Z(n15213) );
  XOR U15654 ( .A(n31372), .B(n31123), .Z(n15138) );
  NAND U15655 ( .A(n15138), .B(n29949), .Z(n14798) );
  NAND U15656 ( .A(n29948), .B(n14796), .Z(n14797) );
  NAND U15657 ( .A(n14798), .B(n14797), .Z(n15210) );
  XOR U15658 ( .A(b[55]), .B(n17133), .Z(n15141) );
  NANDN U15659 ( .A(n15141), .B(n38075), .Z(n14801) );
  NANDN U15660 ( .A(n14799), .B(n38073), .Z(n14800) );
  AND U15661 ( .A(n14801), .B(n14800), .Z(n15211) );
  XNOR U15662 ( .A(n15210), .B(n15211), .Z(n15212) );
  XNOR U15663 ( .A(n15213), .B(n15212), .Z(n15034) );
  NANDN U15664 ( .A(n14803), .B(n14802), .Z(n14807) );
  NAND U15665 ( .A(n14805), .B(n14804), .Z(n14806) );
  NAND U15666 ( .A(n14807), .B(n14806), .Z(n15031) );
  NANDN U15667 ( .A(n14809), .B(n14808), .Z(n14813) );
  NAND U15668 ( .A(n14811), .B(n14810), .Z(n14812) );
  NAND U15669 ( .A(n14813), .B(n14812), .Z(n15032) );
  XNOR U15670 ( .A(n15031), .B(n15032), .Z(n15033) );
  XOR U15671 ( .A(n15034), .B(n15033), .Z(n15250) );
  XNOR U15672 ( .A(n15251), .B(n15250), .Z(n15244) );
  XOR U15673 ( .A(n15245), .B(n15244), .Z(n15246) );
  XNOR U15674 ( .A(n15247), .B(n15246), .Z(n15007) );
  NANDN U15675 ( .A(n14815), .B(n14814), .Z(n14819) );
  OR U15676 ( .A(n14817), .B(n14816), .Z(n14818) );
  AND U15677 ( .A(n14819), .B(n14818), .Z(n15257) );
  NANDN U15678 ( .A(n14821), .B(n14820), .Z(n14825) );
  NAND U15679 ( .A(n14823), .B(n14822), .Z(n14824) );
  NAND U15680 ( .A(n14825), .B(n14824), .Z(n15254) );
  NANDN U15681 ( .A(n14827), .B(n14826), .Z(n14831) );
  NANDN U15682 ( .A(n14829), .B(n14828), .Z(n14830) );
  NAND U15683 ( .A(n14831), .B(n14830), .Z(n15255) );
  XNOR U15684 ( .A(n15254), .B(n15255), .Z(n15256) );
  XNOR U15685 ( .A(n15257), .B(n15256), .Z(n15238) );
  NAND U15686 ( .A(n14833), .B(n14832), .Z(n14837) );
  OR U15687 ( .A(n14835), .B(n14834), .Z(n14836) );
  AND U15688 ( .A(n14837), .B(n14836), .Z(n15239) );
  XNOR U15689 ( .A(n15238), .B(n15239), .Z(n15241) );
  NAND U15690 ( .A(n33283), .B(n14842), .Z(n14844) );
  XNOR U15691 ( .A(n33020), .B(a[62]), .Z(n15047) );
  NANDN U15692 ( .A(n33021), .B(n15047), .Z(n14843) );
  NAND U15693 ( .A(n14844), .B(n14843), .Z(n15095) );
  XNOR U15694 ( .A(b[21]), .B(a[60]), .Z(n15050) );
  OR U15695 ( .A(n15050), .B(n33634), .Z(n14847) );
  NAND U15696 ( .A(n14845), .B(n33464), .Z(n14846) );
  NAND U15697 ( .A(n14847), .B(n14846), .Z(n15092) );
  NAND U15698 ( .A(n34044), .B(n14848), .Z(n14850) );
  XOR U15699 ( .A(n34510), .B(n26347), .Z(n15053) );
  NANDN U15700 ( .A(n33867), .B(n15053), .Z(n14849) );
  AND U15701 ( .A(n14850), .B(n14849), .Z(n15093) );
  XNOR U15702 ( .A(n15092), .B(n15093), .Z(n15094) );
  XNOR U15703 ( .A(n15095), .B(n15094), .Z(n15156) );
  NANDN U15704 ( .A(n14852), .B(n14851), .Z(n14856) );
  NAND U15705 ( .A(n14854), .B(n14853), .Z(n14855) );
  NAND U15706 ( .A(n14856), .B(n14855), .Z(n15157) );
  XNOR U15707 ( .A(n15156), .B(n15157), .Z(n15158) );
  NAND U15708 ( .A(a[16]), .B(b[63]), .Z(n15147) );
  NANDN U15709 ( .A(n14857), .B(n38369), .Z(n14859) );
  XOR U15710 ( .A(b[61]), .B(n15484), .Z(n15062) );
  OR U15711 ( .A(n15062), .B(n38371), .Z(n14858) );
  NAND U15712 ( .A(n14859), .B(n14858), .Z(n15145) );
  NANDN U15713 ( .A(n14860), .B(n35311), .Z(n14862) );
  XOR U15714 ( .A(b[31]), .B(n24671), .Z(n15065) );
  NANDN U15715 ( .A(n15065), .B(n35313), .Z(n14861) );
  AND U15716 ( .A(n14862), .B(n14861), .Z(n15144) );
  XNOR U15717 ( .A(n15145), .B(n15144), .Z(n15146) );
  XNOR U15718 ( .A(n15147), .B(n15146), .Z(n15159) );
  XOR U15719 ( .A(n15158), .B(n15159), .Z(n15019) );
  XOR U15720 ( .A(b[13]), .B(n29868), .Z(n15077) );
  OR U15721 ( .A(n15077), .B(n31550), .Z(n14865) );
  NANDN U15722 ( .A(n14863), .B(n31874), .Z(n14864) );
  NAND U15723 ( .A(n14865), .B(n14864), .Z(n15207) );
  NAND U15724 ( .A(n34848), .B(n14866), .Z(n14868) );
  XOR U15725 ( .A(n35375), .B(n25177), .Z(n15080) );
  NAND U15726 ( .A(n34618), .B(n15080), .Z(n14867) );
  NAND U15727 ( .A(n14868), .B(n14867), .Z(n15204) );
  NAND U15728 ( .A(n35188), .B(n14869), .Z(n14871) );
  XOR U15729 ( .A(n35540), .B(n25134), .Z(n15083) );
  NANDN U15730 ( .A(n34968), .B(n15083), .Z(n14870) );
  AND U15731 ( .A(n14871), .B(n14870), .Z(n15205) );
  XNOR U15732 ( .A(n15204), .B(n15205), .Z(n15206) );
  XNOR U15733 ( .A(n15207), .B(n15206), .Z(n15025) );
  XOR U15734 ( .A(b[37]), .B(n22289), .Z(n15068) );
  NANDN U15735 ( .A(n15068), .B(n36311), .Z(n14874) );
  NANDN U15736 ( .A(n14872), .B(n36309), .Z(n14873) );
  NAND U15737 ( .A(n14874), .B(n14873), .Z(n15126) );
  XOR U15738 ( .A(a[76]), .B(n968), .Z(n15071) );
  OR U15739 ( .A(n15071), .B(n29363), .Z(n14877) );
  NANDN U15740 ( .A(n14875), .B(n29864), .Z(n14876) );
  NAND U15741 ( .A(n14877), .B(n14876), .Z(n15123) );
  XOR U15742 ( .A(n31870), .B(n967), .Z(n15074) );
  NAND U15743 ( .A(n15074), .B(n28939), .Z(n14880) );
  NAND U15744 ( .A(n28938), .B(n14878), .Z(n14879) );
  AND U15745 ( .A(n14880), .B(n14879), .Z(n15124) );
  XNOR U15746 ( .A(n15123), .B(n15124), .Z(n15125) );
  XOR U15747 ( .A(n15126), .B(n15125), .Z(n15026) );
  XOR U15748 ( .A(n15025), .B(n15026), .Z(n15028) );
  NANDN U15749 ( .A(n14882), .B(n14881), .Z(n14886) );
  NAND U15750 ( .A(n14884), .B(n14883), .Z(n14885) );
  NAND U15751 ( .A(n14886), .B(n14885), .Z(n15027) );
  XOR U15752 ( .A(n15028), .B(n15027), .Z(n15020) );
  XNOR U15753 ( .A(n15019), .B(n15020), .Z(n15021) );
  XOR U15754 ( .A(n15022), .B(n15021), .Z(n15234) );
  NANDN U15755 ( .A(n14888), .B(n14887), .Z(n14892) );
  NANDN U15756 ( .A(n14890), .B(n14889), .Z(n14891) );
  NAND U15757 ( .A(n14892), .B(n14891), .Z(n15233) );
  NANDN U15758 ( .A(n14894), .B(n14893), .Z(n14898) );
  NAND U15759 ( .A(n14896), .B(n14895), .Z(n14897) );
  NAND U15760 ( .A(n14898), .B(n14897), .Z(n15040) );
  XOR U15761 ( .A(b[33]), .B(n23447), .Z(n15107) );
  NANDN U15762 ( .A(n15107), .B(n35620), .Z(n14901) );
  NANDN U15763 ( .A(n14899), .B(n35621), .Z(n14900) );
  NAND U15764 ( .A(n14901), .B(n14900), .Z(n15219) );
  NANDN U15765 ( .A(n966), .B(a[80]), .Z(n14902) );
  XOR U15766 ( .A(n29232), .B(n14902), .Z(n14904) );
  NANDN U15767 ( .A(b[0]), .B(a[79]), .Z(n14903) );
  AND U15768 ( .A(n14904), .B(n14903), .Z(n15216) );
  XOR U15769 ( .A(b[63]), .B(n14905), .Z(n15114) );
  NANDN U15770 ( .A(n15114), .B(n38422), .Z(n14908) );
  NANDN U15771 ( .A(n14906), .B(n38423), .Z(n14907) );
  AND U15772 ( .A(n14908), .B(n14907), .Z(n15217) );
  XNOR U15773 ( .A(n15216), .B(n15217), .Z(n15218) );
  XNOR U15774 ( .A(n15219), .B(n15218), .Z(n15222) );
  XNOR U15775 ( .A(b[41]), .B(a[40]), .Z(n15098) );
  OR U15776 ( .A(n15098), .B(n36905), .Z(n14911) );
  NANDN U15777 ( .A(n14909), .B(n36807), .Z(n14910) );
  NAND U15778 ( .A(n14911), .B(n14910), .Z(n15120) );
  XOR U15779 ( .A(b[57]), .B(n16508), .Z(n15101) );
  OR U15780 ( .A(n15101), .B(n965), .Z(n14914) );
  NANDN U15781 ( .A(n14912), .B(n38194), .Z(n14913) );
  NAND U15782 ( .A(n14914), .B(n14913), .Z(n15117) );
  NAND U15783 ( .A(n38326), .B(n14915), .Z(n14917) );
  XOR U15784 ( .A(n38400), .B(n15963), .Z(n15104) );
  NANDN U15785 ( .A(n38273), .B(n15104), .Z(n14916) );
  AND U15786 ( .A(n14917), .B(n14916), .Z(n15118) );
  XNOR U15787 ( .A(n15117), .B(n15118), .Z(n15119) );
  XNOR U15788 ( .A(n15120), .B(n15119), .Z(n15220) );
  NANDN U15789 ( .A(n14919), .B(n14918), .Z(n14923) );
  NAND U15790 ( .A(n14921), .B(n14920), .Z(n14922) );
  NAND U15791 ( .A(n14923), .B(n14922), .Z(n15221) );
  XOR U15792 ( .A(n15220), .B(n15221), .Z(n15223) );
  XNOR U15793 ( .A(n15222), .B(n15223), .Z(n15037) );
  NANDN U15794 ( .A(n14925), .B(n14924), .Z(n14929) );
  NAND U15795 ( .A(n14927), .B(n14926), .Z(n14928) );
  AND U15796 ( .A(n14929), .B(n14928), .Z(n15038) );
  XOR U15797 ( .A(n15037), .B(n15038), .Z(n15039) );
  XNOR U15798 ( .A(n15040), .B(n15039), .Z(n15232) );
  XNOR U15799 ( .A(n15233), .B(n15232), .Z(n15235) );
  XNOR U15800 ( .A(n15234), .B(n15235), .Z(n15240) );
  XOR U15801 ( .A(n15241), .B(n15240), .Z(n15008) );
  XOR U15802 ( .A(n15007), .B(n15008), .Z(n15009) );
  XNOR U15803 ( .A(n15010), .B(n15009), .Z(n15003) );
  OR U15804 ( .A(n14931), .B(n14930), .Z(n14935) );
  NAND U15805 ( .A(n14933), .B(n14932), .Z(n14934) );
  AND U15806 ( .A(n14935), .B(n14934), .Z(n15001) );
  NAND U15807 ( .A(n14937), .B(n14936), .Z(n14941) );
  NANDN U15808 ( .A(n14939), .B(n14938), .Z(n14940) );
  NAND U15809 ( .A(n14941), .B(n14940), .Z(n15016) );
  NANDN U15810 ( .A(n14943), .B(n14942), .Z(n14947) );
  NAND U15811 ( .A(n14945), .B(n14944), .Z(n14946) );
  NAND U15812 ( .A(n14947), .B(n14946), .Z(n15014) );
  OR U15813 ( .A(n14949), .B(n14948), .Z(n14953) );
  NAND U15814 ( .A(n14951), .B(n14950), .Z(n14952) );
  AND U15815 ( .A(n14953), .B(n14952), .Z(n15013) );
  XNOR U15816 ( .A(n15014), .B(n15013), .Z(n15015) );
  XOR U15817 ( .A(n15016), .B(n15015), .Z(n15002) );
  XNOR U15818 ( .A(n15003), .B(n15004), .Z(n14998) );
  NANDN U15819 ( .A(n14955), .B(n14954), .Z(n14959) );
  NAND U15820 ( .A(n14957), .B(n14956), .Z(n14958) );
  NAND U15821 ( .A(n14959), .B(n14958), .Z(n14995) );
  NANDN U15822 ( .A(n14961), .B(n14960), .Z(n14965) );
  NANDN U15823 ( .A(n14963), .B(n14962), .Z(n14964) );
  NAND U15824 ( .A(n14965), .B(n14964), .Z(n14996) );
  XNOR U15825 ( .A(n14995), .B(n14996), .Z(n14997) );
  XNOR U15826 ( .A(n14998), .B(n14997), .Z(n15262) );
  NANDN U15827 ( .A(n14967), .B(n14966), .Z(n14971) );
  NAND U15828 ( .A(n14969), .B(n14968), .Z(n14970) );
  NAND U15829 ( .A(n14971), .B(n14970), .Z(n15263) );
  XOR U15830 ( .A(n15262), .B(n15263), .Z(n15264) );
  NANDN U15831 ( .A(n14973), .B(n14972), .Z(n14977) );
  NANDN U15832 ( .A(n14975), .B(n14974), .Z(n14976) );
  NAND U15833 ( .A(n14977), .B(n14976), .Z(n15265) );
  XOR U15834 ( .A(n15264), .B(n15265), .Z(n14989) );
  NANDN U15835 ( .A(n14979), .B(n14978), .Z(n14983) );
  NAND U15836 ( .A(n14981), .B(n14980), .Z(n14982) );
  NAND U15837 ( .A(n14983), .B(n14982), .Z(n14990) );
  XNOR U15838 ( .A(n14989), .B(n14990), .Z(n14991) );
  XNOR U15839 ( .A(n14992), .B(n14991), .Z(n15268) );
  XNOR U15840 ( .A(n15268), .B(sreg[144]), .Z(n15270) );
  NAND U15841 ( .A(n14984), .B(sreg[143]), .Z(n14988) );
  OR U15842 ( .A(n14986), .B(n14985), .Z(n14987) );
  AND U15843 ( .A(n14988), .B(n14987), .Z(n15269) );
  XOR U15844 ( .A(n15270), .B(n15269), .Z(c[144]) );
  NANDN U15845 ( .A(n14990), .B(n14989), .Z(n14994) );
  NAND U15846 ( .A(n14992), .B(n14991), .Z(n14993) );
  NAND U15847 ( .A(n14994), .B(n14993), .Z(n15276) );
  NANDN U15848 ( .A(n14996), .B(n14995), .Z(n15000) );
  NANDN U15849 ( .A(n14998), .B(n14997), .Z(n14999) );
  NAND U15850 ( .A(n15000), .B(n14999), .Z(n15554) );
  OR U15851 ( .A(n15002), .B(n15001), .Z(n15006) );
  NANDN U15852 ( .A(n15004), .B(n15003), .Z(n15005) );
  NAND U15853 ( .A(n15006), .B(n15005), .Z(n15555) );
  XNOR U15854 ( .A(n15554), .B(n15555), .Z(n15556) );
  OR U15855 ( .A(n15008), .B(n15007), .Z(n15012) );
  NAND U15856 ( .A(n15010), .B(n15009), .Z(n15011) );
  NAND U15857 ( .A(n15012), .B(n15011), .Z(n15548) );
  NANDN U15858 ( .A(n15014), .B(n15013), .Z(n15018) );
  NANDN U15859 ( .A(n15016), .B(n15015), .Z(n15017) );
  NAND U15860 ( .A(n15018), .B(n15017), .Z(n15549) );
  XNOR U15861 ( .A(n15548), .B(n15549), .Z(n15550) );
  NANDN U15862 ( .A(n15020), .B(n15019), .Z(n15024) );
  NANDN U15863 ( .A(n15022), .B(n15021), .Z(n15023) );
  NAND U15864 ( .A(n15024), .B(n15023), .Z(n15279) );
  NANDN U15865 ( .A(n15026), .B(n15025), .Z(n15030) );
  OR U15866 ( .A(n15028), .B(n15027), .Z(n15029) );
  NAND U15867 ( .A(n15030), .B(n15029), .Z(n15526) );
  NANDN U15868 ( .A(n15032), .B(n15031), .Z(n15036) );
  NAND U15869 ( .A(n15034), .B(n15033), .Z(n15035) );
  AND U15870 ( .A(n15036), .B(n15035), .Z(n15524) );
  NAND U15871 ( .A(n15038), .B(n15037), .Z(n15042) );
  NANDN U15872 ( .A(n15040), .B(n15039), .Z(n15041) );
  AND U15873 ( .A(n15042), .B(n15041), .Z(n15525) );
  XOR U15874 ( .A(n15526), .B(n15527), .Z(n15280) );
  XOR U15875 ( .A(n15279), .B(n15280), .Z(n15281) );
  NAND U15876 ( .A(n33283), .B(n15047), .Z(n15049) );
  XNOR U15877 ( .A(n33020), .B(a[63]), .Z(n15454) );
  NANDN U15878 ( .A(n33021), .B(n15454), .Z(n15048) );
  NAND U15879 ( .A(n15049), .B(n15048), .Z(n15466) );
  XNOR U15880 ( .A(b[21]), .B(a[61]), .Z(n15457) );
  OR U15881 ( .A(n15457), .B(n33634), .Z(n15052) );
  NANDN U15882 ( .A(n15050), .B(n33464), .Z(n15051) );
  NAND U15883 ( .A(n15052), .B(n15051), .Z(n15463) );
  NAND U15884 ( .A(n34044), .B(n15053), .Z(n15055) );
  XNOR U15885 ( .A(n34510), .B(a[59]), .Z(n15460) );
  NANDN U15886 ( .A(n33867), .B(n15460), .Z(n15054) );
  AND U15887 ( .A(n15055), .B(n15054), .Z(n15464) );
  XNOR U15888 ( .A(n15463), .B(n15464), .Z(n15465) );
  XOR U15889 ( .A(n15466), .B(n15465), .Z(n15291) );
  NANDN U15890 ( .A(n15057), .B(n15056), .Z(n15061) );
  NAND U15891 ( .A(n15059), .B(n15058), .Z(n15060) );
  NAND U15892 ( .A(n15061), .B(n15060), .Z(n15292) );
  XNOR U15893 ( .A(n15291), .B(n15292), .Z(n15294) );
  NAND U15894 ( .A(a[17]), .B(b[63]), .Z(n15333) );
  NANDN U15895 ( .A(n15062), .B(n38369), .Z(n15064) );
  XOR U15896 ( .A(b[61]), .B(n16220), .Z(n15448) );
  OR U15897 ( .A(n15448), .B(n38371), .Z(n15063) );
  NAND U15898 ( .A(n15064), .B(n15063), .Z(n15331) );
  NANDN U15899 ( .A(n15065), .B(n35311), .Z(n15067) );
  XOR U15900 ( .A(b[31]), .B(n24288), .Z(n15451) );
  NANDN U15901 ( .A(n15451), .B(n35313), .Z(n15066) );
  AND U15902 ( .A(n15067), .B(n15066), .Z(n15330) );
  XNOR U15903 ( .A(n15331), .B(n15330), .Z(n15332) );
  XNOR U15904 ( .A(n15333), .B(n15332), .Z(n15293) );
  XNOR U15905 ( .A(n15294), .B(n15293), .Z(n15406) );
  XOR U15906 ( .A(b[37]), .B(n22579), .Z(n15418) );
  NANDN U15907 ( .A(n15418), .B(n36311), .Z(n15070) );
  NANDN U15908 ( .A(n15068), .B(n36309), .Z(n15069) );
  NAND U15909 ( .A(n15070), .B(n15069), .Z(n15497) );
  XNOR U15910 ( .A(a[77]), .B(b[5]), .Z(n15421) );
  OR U15911 ( .A(n15421), .B(n29363), .Z(n15073) );
  NANDN U15912 ( .A(n15071), .B(n29864), .Z(n15072) );
  NAND U15913 ( .A(n15073), .B(n15072), .Z(n15494) );
  XNOR U15914 ( .A(a[79]), .B(n967), .Z(n15424) );
  NAND U15915 ( .A(n15424), .B(n28939), .Z(n15076) );
  NAND U15916 ( .A(n28938), .B(n15074), .Z(n15075) );
  AND U15917 ( .A(n15076), .B(n15075), .Z(n15495) );
  XNOR U15918 ( .A(n15494), .B(n15495), .Z(n15496) );
  XNOR U15919 ( .A(n15497), .B(n15496), .Z(n15388) );
  XNOR U15920 ( .A(b[13]), .B(a[69]), .Z(n15427) );
  OR U15921 ( .A(n15427), .B(n31550), .Z(n15079) );
  NANDN U15922 ( .A(n15077), .B(n31874), .Z(n15078) );
  NAND U15923 ( .A(n15079), .B(n15078), .Z(n15361) );
  NAND U15924 ( .A(n34848), .B(n15080), .Z(n15082) );
  XOR U15925 ( .A(n35375), .B(n25466), .Z(n15430) );
  NAND U15926 ( .A(n34618), .B(n15430), .Z(n15081) );
  NAND U15927 ( .A(n15082), .B(n15081), .Z(n15358) );
  NAND U15928 ( .A(n35188), .B(n15083), .Z(n15085) );
  XOR U15929 ( .A(n35540), .B(n25001), .Z(n15433) );
  NANDN U15930 ( .A(n34968), .B(n15433), .Z(n15084) );
  AND U15931 ( .A(n15085), .B(n15084), .Z(n15359) );
  XNOR U15932 ( .A(n15358), .B(n15359), .Z(n15360) );
  XOR U15933 ( .A(n15361), .B(n15360), .Z(n15389) );
  XOR U15934 ( .A(n15388), .B(n15389), .Z(n15391) );
  NANDN U15935 ( .A(n15087), .B(n15086), .Z(n15091) );
  NAND U15936 ( .A(n15089), .B(n15088), .Z(n15090) );
  NAND U15937 ( .A(n15091), .B(n15090), .Z(n15390) );
  XOR U15938 ( .A(n15391), .B(n15390), .Z(n15407) );
  XOR U15939 ( .A(n15406), .B(n15407), .Z(n15409) );
  XNOR U15940 ( .A(n15408), .B(n15409), .Z(n15288) );
  NANDN U15941 ( .A(n15093), .B(n15092), .Z(n15097) );
  NAND U15942 ( .A(n15095), .B(n15094), .Z(n15096) );
  NAND U15943 ( .A(n15097), .B(n15096), .Z(n15379) );
  XNOR U15944 ( .A(b[41]), .B(a[41]), .Z(n15469) );
  OR U15945 ( .A(n15469), .B(n36905), .Z(n15100) );
  NANDN U15946 ( .A(n15098), .B(n36807), .Z(n15099) );
  NAND U15947 ( .A(n15100), .B(n15099), .Z(n15491) );
  XOR U15948 ( .A(b[57]), .B(n16916), .Z(n15472) );
  OR U15949 ( .A(n15472), .B(n965), .Z(n15103) );
  NANDN U15950 ( .A(n15101), .B(n38194), .Z(n15102) );
  NAND U15951 ( .A(n15103), .B(n15102), .Z(n15488) );
  NAND U15952 ( .A(n38326), .B(n15104), .Z(n15106) );
  XOR U15953 ( .A(n38400), .B(n16269), .Z(n15475) );
  NANDN U15954 ( .A(n38273), .B(n15475), .Z(n15105) );
  AND U15955 ( .A(n15106), .B(n15105), .Z(n15489) );
  XNOR U15956 ( .A(n15488), .B(n15489), .Z(n15490) );
  XOR U15957 ( .A(n15491), .B(n15490), .Z(n15376) );
  XOR U15958 ( .A(b[33]), .B(n23852), .Z(n15478) );
  NANDN U15959 ( .A(n15478), .B(n35620), .Z(n15109) );
  NANDN U15960 ( .A(n15107), .B(n35621), .Z(n15108) );
  NAND U15961 ( .A(n15109), .B(n15108), .Z(n15373) );
  NANDN U15962 ( .A(n966), .B(a[81]), .Z(n15110) );
  XOR U15963 ( .A(n29232), .B(n15110), .Z(n15112) );
  IV U15964 ( .A(a[80]), .Z(n32814) );
  NANDN U15965 ( .A(n32814), .B(n966), .Z(n15111) );
  AND U15966 ( .A(n15112), .B(n15111), .Z(n15370) );
  XOR U15967 ( .A(b[63]), .B(n15113), .Z(n15485) );
  NANDN U15968 ( .A(n15485), .B(n38422), .Z(n15116) );
  NANDN U15969 ( .A(n15114), .B(n38423), .Z(n15115) );
  AND U15970 ( .A(n15116), .B(n15115), .Z(n15371) );
  XNOR U15971 ( .A(n15370), .B(n15371), .Z(n15372) );
  XOR U15972 ( .A(n15373), .B(n15372), .Z(n15377) );
  XNOR U15973 ( .A(n15376), .B(n15377), .Z(n15378) );
  XNOR U15974 ( .A(n15379), .B(n15378), .Z(n15403) );
  NANDN U15975 ( .A(n15118), .B(n15117), .Z(n15122) );
  NAND U15976 ( .A(n15120), .B(n15119), .Z(n15121) );
  NAND U15977 ( .A(n15122), .B(n15121), .Z(n15400) );
  NANDN U15978 ( .A(n15124), .B(n15123), .Z(n15128) );
  NAND U15979 ( .A(n15126), .B(n15125), .Z(n15127) );
  AND U15980 ( .A(n15128), .B(n15127), .Z(n15401) );
  XNOR U15981 ( .A(n15400), .B(n15401), .Z(n15402) );
  XOR U15982 ( .A(n15403), .B(n15402), .Z(n15286) );
  NANDN U15983 ( .A(n15130), .B(n15129), .Z(n15134) );
  NAND U15984 ( .A(n15132), .B(n15131), .Z(n15133) );
  AND U15985 ( .A(n15134), .B(n15133), .Z(n15285) );
  XOR U15986 ( .A(n15286), .B(n15285), .Z(n15287) );
  XNOR U15987 ( .A(n15288), .B(n15287), .Z(n15282) );
  XOR U15988 ( .A(n15281), .B(n15282), .Z(n15536) );
  XNOR U15989 ( .A(b[35]), .B(a[47]), .Z(n15321) );
  NANDN U15990 ( .A(n15321), .B(n35985), .Z(n15137) );
  NANDN U15991 ( .A(n15135), .B(n35986), .Z(n15136) );
  NAND U15992 ( .A(n15137), .B(n15136), .Z(n15367) );
  XNOR U15993 ( .A(a[75]), .B(n31123), .Z(n15324) );
  NAND U15994 ( .A(n15324), .B(n29949), .Z(n15140) );
  NAND U15995 ( .A(n29948), .B(n15138), .Z(n15139) );
  NAND U15996 ( .A(n15140), .B(n15139), .Z(n15364) );
  XOR U15997 ( .A(b[55]), .B(n17960), .Z(n15327) );
  NANDN U15998 ( .A(n15327), .B(n38075), .Z(n15143) );
  NANDN U15999 ( .A(n15141), .B(n38073), .Z(n15142) );
  AND U16000 ( .A(n15143), .B(n15142), .Z(n15365) );
  XNOR U16001 ( .A(n15364), .B(n15365), .Z(n15366) );
  XNOR U16002 ( .A(n15367), .B(n15366), .Z(n15397) );
  NANDN U16003 ( .A(n15145), .B(n15144), .Z(n15149) );
  NAND U16004 ( .A(n15147), .B(n15146), .Z(n15148) );
  NAND U16005 ( .A(n15149), .B(n15148), .Z(n15394) );
  NANDN U16006 ( .A(n15151), .B(n15150), .Z(n15155) );
  NAND U16007 ( .A(n15153), .B(n15152), .Z(n15154) );
  NAND U16008 ( .A(n15155), .B(n15154), .Z(n15395) );
  XNOR U16009 ( .A(n15394), .B(n15395), .Z(n15396) );
  XOR U16010 ( .A(n15397), .B(n15396), .Z(n15514) );
  NANDN U16011 ( .A(n15157), .B(n15156), .Z(n15161) );
  NANDN U16012 ( .A(n15159), .B(n15158), .Z(n15160) );
  NAND U16013 ( .A(n15161), .B(n15160), .Z(n15513) );
  XOR U16014 ( .A(b[11]), .B(n30543), .Z(n15306) );
  OR U16015 ( .A(n15306), .B(n31369), .Z(n15164) );
  NANDN U16016 ( .A(n15162), .B(n31119), .Z(n15163) );
  NAND U16017 ( .A(n15164), .B(n15163), .Z(n15318) );
  XOR U16018 ( .A(b[43]), .B(n20867), .Z(n15309) );
  NANDN U16019 ( .A(n15309), .B(n37068), .Z(n15167) );
  NANDN U16020 ( .A(n15165), .B(n37069), .Z(n15166) );
  NAND U16021 ( .A(n15167), .B(n15166), .Z(n15315) );
  XNOR U16022 ( .A(b[45]), .B(a[37]), .Z(n15312) );
  NANDN U16023 ( .A(n15312), .B(n37261), .Z(n15170) );
  NANDN U16024 ( .A(n15168), .B(n37262), .Z(n15169) );
  AND U16025 ( .A(n15170), .B(n15169), .Z(n15316) );
  XNOR U16026 ( .A(n15315), .B(n15316), .Z(n15317) );
  XNOR U16027 ( .A(n15318), .B(n15317), .Z(n15415) );
  NAND U16028 ( .A(n37652), .B(n15171), .Z(n15173) );
  XOR U16029 ( .A(b[49]), .B(n19656), .Z(n15297) );
  OR U16030 ( .A(n15297), .B(n37756), .Z(n15172) );
  NAND U16031 ( .A(n15173), .B(n15172), .Z(n15338) );
  NANDN U16032 ( .A(n15174), .B(n37469), .Z(n15176) );
  XNOR U16033 ( .A(n978), .B(a[35]), .Z(n15300) );
  NAND U16034 ( .A(n15300), .B(n37471), .Z(n15175) );
  NAND U16035 ( .A(n15176), .B(n15175), .Z(n15336) );
  NAND U16036 ( .A(n30846), .B(n15177), .Z(n15179) );
  XNOR U16037 ( .A(n969), .B(a[73]), .Z(n15303) );
  NAND U16038 ( .A(n30509), .B(n15303), .Z(n15178) );
  NAND U16039 ( .A(n15179), .B(n15178), .Z(n15337) );
  XNOR U16040 ( .A(n15336), .B(n15337), .Z(n15339) );
  XOR U16041 ( .A(n15338), .B(n15339), .Z(n15412) );
  NANDN U16042 ( .A(n15181), .B(n15180), .Z(n15185) );
  NAND U16043 ( .A(n15183), .B(n15182), .Z(n15184) );
  NAND U16044 ( .A(n15185), .B(n15184), .Z(n15413) );
  XNOR U16045 ( .A(n15412), .B(n15413), .Z(n15414) );
  XOR U16046 ( .A(n15415), .B(n15414), .Z(n15512) );
  XNOR U16047 ( .A(n15513), .B(n15512), .Z(n15515) );
  XNOR U16048 ( .A(n15514), .B(n15515), .Z(n15506) );
  XOR U16049 ( .A(b[15]), .B(n29372), .Z(n15340) );
  OR U16050 ( .A(n15340), .B(n32010), .Z(n15188) );
  NANDN U16051 ( .A(n15186), .B(n32011), .Z(n15187) );
  NAND U16052 ( .A(n15188), .B(n15187), .Z(n15445) );
  XNOR U16053 ( .A(b[25]), .B(n26122), .Z(n15343) );
  NANDN U16054 ( .A(n34219), .B(n15343), .Z(n15191) );
  NAND U16055 ( .A(n34217), .B(n15189), .Z(n15190) );
  NAND U16056 ( .A(n15191), .B(n15190), .Z(n15442) );
  XNOR U16057 ( .A(b[17]), .B(a[65]), .Z(n15346) );
  NANDN U16058 ( .A(n15346), .B(n32543), .Z(n15194) );
  NAND U16059 ( .A(n15192), .B(n32541), .Z(n15193) );
  AND U16060 ( .A(n15194), .B(n15193), .Z(n15443) );
  XNOR U16061 ( .A(n15442), .B(n15443), .Z(n15444) );
  XNOR U16062 ( .A(n15445), .B(n15444), .Z(n15500) );
  XOR U16063 ( .A(b[39]), .B(n21996), .Z(n15349) );
  NANDN U16064 ( .A(n15349), .B(n36553), .Z(n15197) );
  NANDN U16065 ( .A(n15195), .B(n36643), .Z(n15196) );
  NAND U16066 ( .A(n15197), .B(n15196), .Z(n15439) );
  XOR U16067 ( .A(b[51]), .B(n18639), .Z(n15352) );
  NANDN U16068 ( .A(n15352), .B(n37803), .Z(n15200) );
  NANDN U16069 ( .A(n15198), .B(n37802), .Z(n15199) );
  NAND U16070 ( .A(n15200), .B(n15199), .Z(n15436) );
  XOR U16071 ( .A(b[53]), .B(n18003), .Z(n15355) );
  NANDN U16072 ( .A(n15355), .B(n37940), .Z(n15203) );
  NANDN U16073 ( .A(n15201), .B(n37941), .Z(n15202) );
  AND U16074 ( .A(n15203), .B(n15202), .Z(n15437) );
  XNOR U16075 ( .A(n15436), .B(n15437), .Z(n15438) );
  XOR U16076 ( .A(n15439), .B(n15438), .Z(n15501) );
  XOR U16077 ( .A(n15500), .B(n15501), .Z(n15503) );
  NANDN U16078 ( .A(n15205), .B(n15204), .Z(n15209) );
  NAND U16079 ( .A(n15207), .B(n15206), .Z(n15208) );
  NAND U16080 ( .A(n15209), .B(n15208), .Z(n15502) );
  XNOR U16081 ( .A(n15503), .B(n15502), .Z(n15385) );
  NANDN U16082 ( .A(n15211), .B(n15210), .Z(n15215) );
  NAND U16083 ( .A(n15213), .B(n15212), .Z(n15214) );
  NAND U16084 ( .A(n15215), .B(n15214), .Z(n15382) );
  XNOR U16085 ( .A(n15382), .B(n15383), .Z(n15384) );
  XNOR U16086 ( .A(n15385), .B(n15384), .Z(n15521) );
  NANDN U16087 ( .A(n15221), .B(n15220), .Z(n15225) );
  NANDN U16088 ( .A(n15223), .B(n15222), .Z(n15224) );
  NAND U16089 ( .A(n15225), .B(n15224), .Z(n15518) );
  NANDN U16090 ( .A(n15227), .B(n15226), .Z(n15231) );
  NANDN U16091 ( .A(n15229), .B(n15228), .Z(n15230) );
  NAND U16092 ( .A(n15231), .B(n15230), .Z(n15519) );
  XNOR U16093 ( .A(n15518), .B(n15519), .Z(n15520) );
  XOR U16094 ( .A(n15521), .B(n15520), .Z(n15507) );
  NAND U16095 ( .A(n15233), .B(n15232), .Z(n15237) );
  NANDN U16096 ( .A(n15235), .B(n15234), .Z(n15236) );
  AND U16097 ( .A(n15237), .B(n15236), .Z(n15509) );
  XNOR U16098 ( .A(n15508), .B(n15509), .Z(n15537) );
  XNOR U16099 ( .A(n15536), .B(n15537), .Z(n15538) );
  NAND U16100 ( .A(n15239), .B(n15238), .Z(n15243) );
  NANDN U16101 ( .A(n15241), .B(n15240), .Z(n15242) );
  NAND U16102 ( .A(n15243), .B(n15242), .Z(n15539) );
  XOR U16103 ( .A(n15538), .B(n15539), .Z(n15545) );
  NAND U16104 ( .A(n15249), .B(n15248), .Z(n15253) );
  NANDN U16105 ( .A(n15251), .B(n15250), .Z(n15252) );
  NAND U16106 ( .A(n15253), .B(n15252), .Z(n15533) );
  XNOR U16107 ( .A(n15530), .B(n15531), .Z(n15532) );
  XNOR U16108 ( .A(n15533), .B(n15532), .Z(n15543) );
  XNOR U16109 ( .A(n15542), .B(n15543), .Z(n15544) );
  XOR U16110 ( .A(n15545), .B(n15544), .Z(n15551) );
  XOR U16111 ( .A(n15550), .B(n15551), .Z(n15557) );
  XOR U16112 ( .A(n15556), .B(n15557), .Z(n15273) );
  OR U16113 ( .A(n15263), .B(n15262), .Z(n15267) );
  NANDN U16114 ( .A(n15265), .B(n15264), .Z(n15266) );
  AND U16115 ( .A(n15267), .B(n15266), .Z(n15274) );
  XOR U16116 ( .A(n15273), .B(n15274), .Z(n15275) );
  XNOR U16117 ( .A(n15276), .B(n15275), .Z(n15560) );
  XNOR U16118 ( .A(n15560), .B(sreg[145]), .Z(n15562) );
  NAND U16119 ( .A(n15268), .B(sreg[144]), .Z(n15272) );
  OR U16120 ( .A(n15270), .B(n15269), .Z(n15271) );
  AND U16121 ( .A(n15272), .B(n15271), .Z(n15561) );
  XOR U16122 ( .A(n15562), .B(n15561), .Z(c[145]) );
  NAND U16123 ( .A(n15274), .B(n15273), .Z(n15278) );
  NAND U16124 ( .A(n15276), .B(n15275), .Z(n15277) );
  NAND U16125 ( .A(n15278), .B(n15277), .Z(n15568) );
  OR U16126 ( .A(n15280), .B(n15279), .Z(n15284) );
  NANDN U16127 ( .A(n15282), .B(n15281), .Z(n15283) );
  NAND U16128 ( .A(n15284), .B(n15283), .Z(n15586) );
  OR U16129 ( .A(n15286), .B(n15285), .Z(n15290) );
  NAND U16130 ( .A(n15288), .B(n15287), .Z(n15289) );
  NAND U16131 ( .A(n15290), .B(n15289), .Z(n15837) );
  OR U16132 ( .A(n15292), .B(n15291), .Z(n15296) );
  OR U16133 ( .A(n15294), .B(n15293), .Z(n15295) );
  NAND U16134 ( .A(n15296), .B(n15295), .Z(n15821) );
  XOR U16135 ( .A(b[49]), .B(n19513), .Z(n15774) );
  OR U16136 ( .A(n15774), .B(n37756), .Z(n15299) );
  NANDN U16137 ( .A(n15297), .B(n37652), .Z(n15298) );
  NAND U16138 ( .A(n15299), .B(n15298), .Z(n15811) );
  NAND U16139 ( .A(n15300), .B(n37469), .Z(n15302) );
  XOR U16140 ( .A(n978), .B(n19980), .Z(n15777) );
  NAND U16141 ( .A(n15777), .B(n37471), .Z(n15301) );
  NAND U16142 ( .A(n15302), .B(n15301), .Z(n15808) );
  XOR U16143 ( .A(b[9]), .B(n31372), .Z(n15780) );
  NANDN U16144 ( .A(n15780), .B(n30509), .Z(n15305) );
  NAND U16145 ( .A(n15303), .B(n30846), .Z(n15304) );
  AND U16146 ( .A(n15305), .B(n15304), .Z(n15809) );
  XNOR U16147 ( .A(n15808), .B(n15809), .Z(n15810) );
  XNOR U16148 ( .A(n15811), .B(n15810), .Z(n15623) );
  XOR U16149 ( .A(b[11]), .B(n30210), .Z(n15765) );
  OR U16150 ( .A(n15765), .B(n31369), .Z(n15308) );
  NANDN U16151 ( .A(n15306), .B(n31119), .Z(n15307) );
  NAND U16152 ( .A(n15308), .B(n15307), .Z(n15786) );
  XOR U16153 ( .A(b[43]), .B(n21149), .Z(n15768) );
  NANDN U16154 ( .A(n15768), .B(n37068), .Z(n15311) );
  NANDN U16155 ( .A(n15309), .B(n37069), .Z(n15310) );
  NAND U16156 ( .A(n15311), .B(n15310), .Z(n15783) );
  XNOR U16157 ( .A(b[45]), .B(a[38]), .Z(n15771) );
  NANDN U16158 ( .A(n15771), .B(n37261), .Z(n15314) );
  NANDN U16159 ( .A(n15312), .B(n37262), .Z(n15313) );
  AND U16160 ( .A(n15314), .B(n15313), .Z(n15784) );
  XNOR U16161 ( .A(n15783), .B(n15784), .Z(n15785) );
  XNOR U16162 ( .A(n15786), .B(n15785), .Z(n15620) );
  NANDN U16163 ( .A(n15316), .B(n15315), .Z(n15320) );
  NAND U16164 ( .A(n15318), .B(n15317), .Z(n15319) );
  NAND U16165 ( .A(n15320), .B(n15319), .Z(n15621) );
  XNOR U16166 ( .A(n15620), .B(n15621), .Z(n15622) );
  XOR U16167 ( .A(n15623), .B(n15622), .Z(n15820) );
  XNOR U16168 ( .A(n15821), .B(n15820), .Z(n15823) );
  XNOR U16169 ( .A(b[35]), .B(a[48]), .Z(n15793) );
  NANDN U16170 ( .A(n15793), .B(n35985), .Z(n15323) );
  NANDN U16171 ( .A(n15321), .B(n35986), .Z(n15322) );
  NAND U16172 ( .A(n15323), .B(n15322), .Z(n15744) );
  XOR U16173 ( .A(n31363), .B(n31123), .Z(n15796) );
  NAND U16174 ( .A(n15796), .B(n29949), .Z(n15326) );
  NAND U16175 ( .A(n29948), .B(n15324), .Z(n15325) );
  NAND U16176 ( .A(n15326), .B(n15325), .Z(n15741) );
  XOR U16177 ( .A(b[55]), .B(n17702), .Z(n15799) );
  NANDN U16178 ( .A(n15799), .B(n38075), .Z(n15329) );
  NANDN U16179 ( .A(n15327), .B(n38073), .Z(n15328) );
  AND U16180 ( .A(n15329), .B(n15328), .Z(n15742) );
  XNOR U16181 ( .A(n15741), .B(n15742), .Z(n15743) );
  XNOR U16182 ( .A(n15744), .B(n15743), .Z(n15610) );
  NANDN U16183 ( .A(n15331), .B(n15330), .Z(n15335) );
  NAND U16184 ( .A(n15333), .B(n15332), .Z(n15334) );
  NAND U16185 ( .A(n15335), .B(n15334), .Z(n15607) );
  XNOR U16186 ( .A(n15607), .B(n15608), .Z(n15609) );
  XOR U16187 ( .A(n15610), .B(n15609), .Z(n15822) );
  XNOR U16188 ( .A(n15823), .B(n15822), .Z(n15834) );
  XOR U16189 ( .A(b[15]), .B(n29868), .Z(n15717) );
  OR U16190 ( .A(n15717), .B(n32010), .Z(n15342) );
  NANDN U16191 ( .A(n15340), .B(n32011), .Z(n15341) );
  NAND U16192 ( .A(n15342), .B(n15341), .Z(n15651) );
  XNOR U16193 ( .A(b[25]), .B(n26347), .Z(n15720) );
  NANDN U16194 ( .A(n34219), .B(n15720), .Z(n15345) );
  NAND U16195 ( .A(n34217), .B(n15343), .Z(n15344) );
  NAND U16196 ( .A(n15345), .B(n15344), .Z(n15648) );
  XNOR U16197 ( .A(b[17]), .B(a[66]), .Z(n15723) );
  NANDN U16198 ( .A(n15723), .B(n32543), .Z(n15348) );
  NANDN U16199 ( .A(n15346), .B(n32541), .Z(n15347) );
  AND U16200 ( .A(n15348), .B(n15347), .Z(n15649) );
  XNOR U16201 ( .A(n15648), .B(n15649), .Z(n15650) );
  XNOR U16202 ( .A(n15651), .B(n15650), .Z(n15705) );
  XOR U16203 ( .A(b[39]), .B(n22289), .Z(n15726) );
  NANDN U16204 ( .A(n15726), .B(n36553), .Z(n15351) );
  NANDN U16205 ( .A(n15349), .B(n36643), .Z(n15350) );
  NAND U16206 ( .A(n15351), .B(n15350), .Z(n15645) );
  XOR U16207 ( .A(b[51]), .B(n18841), .Z(n15729) );
  NANDN U16208 ( .A(n15729), .B(n37803), .Z(n15354) );
  NANDN U16209 ( .A(n15352), .B(n37802), .Z(n15353) );
  NAND U16210 ( .A(n15354), .B(n15353), .Z(n15642) );
  XOR U16211 ( .A(b[53]), .B(n18804), .Z(n15732) );
  NANDN U16212 ( .A(n15732), .B(n37940), .Z(n15357) );
  NANDN U16213 ( .A(n15355), .B(n37941), .Z(n15356) );
  AND U16214 ( .A(n15357), .B(n15356), .Z(n15643) );
  XNOR U16215 ( .A(n15642), .B(n15643), .Z(n15644) );
  XOR U16216 ( .A(n15645), .B(n15644), .Z(n15706) );
  XOR U16217 ( .A(n15705), .B(n15706), .Z(n15708) );
  NANDN U16218 ( .A(n15359), .B(n15358), .Z(n15363) );
  NAND U16219 ( .A(n15361), .B(n15360), .Z(n15362) );
  NAND U16220 ( .A(n15363), .B(n15362), .Z(n15707) );
  XNOR U16221 ( .A(n15708), .B(n15707), .Z(n15762) );
  NANDN U16222 ( .A(n15365), .B(n15364), .Z(n15369) );
  NAND U16223 ( .A(n15367), .B(n15366), .Z(n15368) );
  NAND U16224 ( .A(n15369), .B(n15368), .Z(n15759) );
  NANDN U16225 ( .A(n15371), .B(n15370), .Z(n15375) );
  NAND U16226 ( .A(n15373), .B(n15372), .Z(n15374) );
  AND U16227 ( .A(n15375), .B(n15374), .Z(n15760) );
  XNOR U16228 ( .A(n15759), .B(n15760), .Z(n15761) );
  XNOR U16229 ( .A(n15762), .B(n15761), .Z(n15826) );
  OR U16230 ( .A(n15377), .B(n15376), .Z(n15381) );
  OR U16231 ( .A(n15379), .B(n15378), .Z(n15380) );
  AND U16232 ( .A(n15381), .B(n15380), .Z(n15827) );
  XNOR U16233 ( .A(n15826), .B(n15827), .Z(n15828) );
  NANDN U16234 ( .A(n15383), .B(n15382), .Z(n15387) );
  NAND U16235 ( .A(n15385), .B(n15384), .Z(n15386) );
  AND U16236 ( .A(n15387), .B(n15386), .Z(n15829) );
  XNOR U16237 ( .A(n15828), .B(n15829), .Z(n15835) );
  XNOR U16238 ( .A(n15834), .B(n15835), .Z(n15836) );
  XNOR U16239 ( .A(n15837), .B(n15836), .Z(n15583) );
  NANDN U16240 ( .A(n15389), .B(n15388), .Z(n15393) );
  OR U16241 ( .A(n15391), .B(n15390), .Z(n15392) );
  AND U16242 ( .A(n15393), .B(n15392), .Z(n15833) );
  NANDN U16243 ( .A(n15395), .B(n15394), .Z(n15399) );
  NAND U16244 ( .A(n15397), .B(n15396), .Z(n15398) );
  NAND U16245 ( .A(n15399), .B(n15398), .Z(n15830) );
  NANDN U16246 ( .A(n15401), .B(n15400), .Z(n15405) );
  NAND U16247 ( .A(n15403), .B(n15402), .Z(n15404) );
  NAND U16248 ( .A(n15405), .B(n15404), .Z(n15831) );
  XNOR U16249 ( .A(n15830), .B(n15831), .Z(n15832) );
  XNOR U16250 ( .A(n15833), .B(n15832), .Z(n15814) );
  NANDN U16251 ( .A(n15407), .B(n15406), .Z(n15411) );
  OR U16252 ( .A(n15409), .B(n15408), .Z(n15410) );
  AND U16253 ( .A(n15411), .B(n15410), .Z(n15815) );
  XNOR U16254 ( .A(n15814), .B(n15815), .Z(n15817) );
  NANDN U16255 ( .A(n15413), .B(n15412), .Z(n15417) );
  NAND U16256 ( .A(n15415), .B(n15414), .Z(n15416) );
  NAND U16257 ( .A(n15417), .B(n15416), .Z(n15616) );
  XOR U16258 ( .A(b[37]), .B(n22964), .Z(n15624) );
  NANDN U16259 ( .A(n15624), .B(n36311), .Z(n15420) );
  NANDN U16260 ( .A(n15418), .B(n36309), .Z(n15419) );
  NAND U16261 ( .A(n15420), .B(n15419), .Z(n15702) );
  XOR U16262 ( .A(a[78]), .B(n968), .Z(n15627) );
  OR U16263 ( .A(n15627), .B(n29363), .Z(n15423) );
  NANDN U16264 ( .A(n15421), .B(n29864), .Z(n15422) );
  NAND U16265 ( .A(n15423), .B(n15422), .Z(n15699) );
  XOR U16266 ( .A(n32814), .B(n967), .Z(n15630) );
  NAND U16267 ( .A(n15630), .B(n28939), .Z(n15426) );
  NAND U16268 ( .A(n28938), .B(n15424), .Z(n15425) );
  AND U16269 ( .A(n15426), .B(n15425), .Z(n15700) );
  XNOR U16270 ( .A(n15699), .B(n15700), .Z(n15701) );
  XOR U16271 ( .A(n15702), .B(n15701), .Z(n15604) );
  XOR U16272 ( .A(b[13]), .B(n30379), .Z(n15633) );
  OR U16273 ( .A(n15633), .B(n31550), .Z(n15429) );
  NANDN U16274 ( .A(n15427), .B(n31874), .Z(n15428) );
  NAND U16275 ( .A(n15429), .B(n15428), .Z(n15738) );
  NAND U16276 ( .A(n34848), .B(n15430), .Z(n15432) );
  XOR U16277 ( .A(n35375), .B(n25860), .Z(n15636) );
  NAND U16278 ( .A(n34618), .B(n15636), .Z(n15431) );
  NAND U16279 ( .A(n15432), .B(n15431), .Z(n15735) );
  NAND U16280 ( .A(n35188), .B(n15433), .Z(n15435) );
  XOR U16281 ( .A(n35540), .B(n25177), .Z(n15639) );
  NANDN U16282 ( .A(n34968), .B(n15639), .Z(n15434) );
  AND U16283 ( .A(n15435), .B(n15434), .Z(n15736) );
  XNOR U16284 ( .A(n15735), .B(n15736), .Z(n15737) );
  XOR U16285 ( .A(n15738), .B(n15737), .Z(n15602) );
  NANDN U16286 ( .A(n15437), .B(n15436), .Z(n15441) );
  NAND U16287 ( .A(n15439), .B(n15438), .Z(n15440) );
  AND U16288 ( .A(n15441), .B(n15440), .Z(n15601) );
  XOR U16289 ( .A(n15602), .B(n15601), .Z(n15603) );
  XOR U16290 ( .A(n15604), .B(n15603), .Z(n15615) );
  NANDN U16291 ( .A(n15443), .B(n15442), .Z(n15447) );
  NAND U16292 ( .A(n15445), .B(n15444), .Z(n15446) );
  NAND U16293 ( .A(n15447), .B(n15446), .Z(n15791) );
  NAND U16294 ( .A(a[18]), .B(b[63]), .Z(n15805) );
  NANDN U16295 ( .A(n15448), .B(n38369), .Z(n15450) );
  XOR U16296 ( .A(b[61]), .B(n15963), .Z(n15654) );
  OR U16297 ( .A(n15654), .B(n38371), .Z(n15449) );
  NAND U16298 ( .A(n15450), .B(n15449), .Z(n15803) );
  NANDN U16299 ( .A(n15451), .B(n35311), .Z(n15453) );
  XOR U16300 ( .A(b[31]), .B(n25134), .Z(n15657) );
  NANDN U16301 ( .A(n15657), .B(n35313), .Z(n15452) );
  AND U16302 ( .A(n15453), .B(n15452), .Z(n15802) );
  XNOR U16303 ( .A(n15803), .B(n15802), .Z(n15804) );
  XOR U16304 ( .A(n15805), .B(n15804), .Z(n15789) );
  NAND U16305 ( .A(n33283), .B(n15454), .Z(n15456) );
  XNOR U16306 ( .A(n33020), .B(a[64]), .Z(n15660) );
  NANDN U16307 ( .A(n33021), .B(n15660), .Z(n15455) );
  NAND U16308 ( .A(n15456), .B(n15455), .Z(n15672) );
  XOR U16309 ( .A(b[21]), .B(a[62]), .Z(n15663) );
  NANDN U16310 ( .A(n33634), .B(n15663), .Z(n15459) );
  NANDN U16311 ( .A(n15457), .B(n33464), .Z(n15458) );
  NAND U16312 ( .A(n15459), .B(n15458), .Z(n15669) );
  NAND U16313 ( .A(n34044), .B(n15460), .Z(n15462) );
  XOR U16314 ( .A(n34510), .B(n27436), .Z(n15666) );
  NANDN U16315 ( .A(n33867), .B(n15666), .Z(n15461) );
  AND U16316 ( .A(n15462), .B(n15461), .Z(n15670) );
  XNOR U16317 ( .A(n15669), .B(n15670), .Z(n15671) );
  XNOR U16318 ( .A(n15672), .B(n15671), .Z(n15790) );
  XNOR U16319 ( .A(n15789), .B(n15790), .Z(n15792) );
  XNOR U16320 ( .A(n15791), .B(n15792), .Z(n15614) );
  XOR U16321 ( .A(n15615), .B(n15614), .Z(n15617) );
  XNOR U16322 ( .A(n15616), .B(n15617), .Z(n15714) );
  NANDN U16323 ( .A(n15464), .B(n15463), .Z(n15468) );
  NAND U16324 ( .A(n15466), .B(n15465), .Z(n15467) );
  NAND U16325 ( .A(n15468), .B(n15467), .Z(n15756) );
  XNOR U16326 ( .A(b[41]), .B(a[42]), .Z(n15675) );
  OR U16327 ( .A(n15675), .B(n36905), .Z(n15471) );
  NANDN U16328 ( .A(n15469), .B(n36807), .Z(n15470) );
  NAND U16329 ( .A(n15471), .B(n15470), .Z(n15696) );
  XOR U16330 ( .A(b[57]), .B(n17133), .Z(n15678) );
  OR U16331 ( .A(n15678), .B(n965), .Z(n15474) );
  NANDN U16332 ( .A(n15472), .B(n38194), .Z(n15473) );
  NAND U16333 ( .A(n15474), .B(n15473), .Z(n15693) );
  NAND U16334 ( .A(n38326), .B(n15475), .Z(n15477) );
  XOR U16335 ( .A(n38400), .B(n16508), .Z(n15681) );
  NANDN U16336 ( .A(n38273), .B(n15681), .Z(n15476) );
  AND U16337 ( .A(n15477), .B(n15476), .Z(n15694) );
  XNOR U16338 ( .A(n15693), .B(n15694), .Z(n15695) );
  XOR U16339 ( .A(n15696), .B(n15695), .Z(n15753) );
  XOR U16340 ( .A(b[33]), .B(n24671), .Z(n15684) );
  NANDN U16341 ( .A(n15684), .B(n35620), .Z(n15480) );
  NANDN U16342 ( .A(n15478), .B(n35621), .Z(n15479) );
  NAND U16343 ( .A(n15480), .B(n15479), .Z(n15750) );
  NANDN U16344 ( .A(n966), .B(a[82]), .Z(n15481) );
  XOR U16345 ( .A(n29232), .B(n15481), .Z(n15483) );
  NANDN U16346 ( .A(b[0]), .B(a[81]), .Z(n15482) );
  AND U16347 ( .A(n15483), .B(n15482), .Z(n15747) );
  XOR U16348 ( .A(b[63]), .B(n15484), .Z(n15690) );
  NANDN U16349 ( .A(n15690), .B(n38422), .Z(n15487) );
  NANDN U16350 ( .A(n15485), .B(n38423), .Z(n15486) );
  AND U16351 ( .A(n15487), .B(n15486), .Z(n15748) );
  XNOR U16352 ( .A(n15747), .B(n15748), .Z(n15749) );
  XOR U16353 ( .A(n15750), .B(n15749), .Z(n15754) );
  XNOR U16354 ( .A(n15753), .B(n15754), .Z(n15755) );
  XNOR U16355 ( .A(n15756), .B(n15755), .Z(n15598) );
  NANDN U16356 ( .A(n15489), .B(n15488), .Z(n15493) );
  NAND U16357 ( .A(n15491), .B(n15490), .Z(n15492) );
  NAND U16358 ( .A(n15493), .B(n15492), .Z(n15595) );
  NANDN U16359 ( .A(n15495), .B(n15494), .Z(n15499) );
  NAND U16360 ( .A(n15497), .B(n15496), .Z(n15498) );
  AND U16361 ( .A(n15499), .B(n15498), .Z(n15596) );
  XNOR U16362 ( .A(n15595), .B(n15596), .Z(n15597) );
  XOR U16363 ( .A(n15598), .B(n15597), .Z(n15712) );
  NANDN U16364 ( .A(n15501), .B(n15500), .Z(n15505) );
  OR U16365 ( .A(n15503), .B(n15502), .Z(n15504) );
  AND U16366 ( .A(n15505), .B(n15504), .Z(n15711) );
  XOR U16367 ( .A(n15712), .B(n15711), .Z(n15713) );
  XOR U16368 ( .A(n15714), .B(n15713), .Z(n15816) );
  XOR U16369 ( .A(n15817), .B(n15816), .Z(n15584) );
  XOR U16370 ( .A(n15583), .B(n15584), .Z(n15585) );
  XNOR U16371 ( .A(n15586), .B(n15585), .Z(n15579) );
  OR U16372 ( .A(n15507), .B(n15506), .Z(n15511) );
  NAND U16373 ( .A(n15509), .B(n15508), .Z(n15510) );
  AND U16374 ( .A(n15511), .B(n15510), .Z(n15577) );
  NAND U16375 ( .A(n15513), .B(n15512), .Z(n15517) );
  NANDN U16376 ( .A(n15515), .B(n15514), .Z(n15516) );
  NAND U16377 ( .A(n15517), .B(n15516), .Z(n15592) );
  NANDN U16378 ( .A(n15519), .B(n15518), .Z(n15523) );
  NAND U16379 ( .A(n15521), .B(n15520), .Z(n15522) );
  NAND U16380 ( .A(n15523), .B(n15522), .Z(n15590) );
  OR U16381 ( .A(n15525), .B(n15524), .Z(n15529) );
  NANDN U16382 ( .A(n15527), .B(n15526), .Z(n15528) );
  AND U16383 ( .A(n15529), .B(n15528), .Z(n15589) );
  XNOR U16384 ( .A(n15590), .B(n15589), .Z(n15591) );
  XOR U16385 ( .A(n15592), .B(n15591), .Z(n15578) );
  XNOR U16386 ( .A(n15579), .B(n15580), .Z(n15574) );
  NANDN U16387 ( .A(n15531), .B(n15530), .Z(n15535) );
  NAND U16388 ( .A(n15533), .B(n15532), .Z(n15534) );
  NAND U16389 ( .A(n15535), .B(n15534), .Z(n15571) );
  NANDN U16390 ( .A(n15537), .B(n15536), .Z(n15541) );
  NANDN U16391 ( .A(n15539), .B(n15538), .Z(n15540) );
  NAND U16392 ( .A(n15541), .B(n15540), .Z(n15572) );
  XNOR U16393 ( .A(n15571), .B(n15572), .Z(n15573) );
  XNOR U16394 ( .A(n15574), .B(n15573), .Z(n15838) );
  NANDN U16395 ( .A(n15543), .B(n15542), .Z(n15547) );
  NAND U16396 ( .A(n15545), .B(n15544), .Z(n15546) );
  NAND U16397 ( .A(n15547), .B(n15546), .Z(n15839) );
  XOR U16398 ( .A(n15838), .B(n15839), .Z(n15840) );
  NANDN U16399 ( .A(n15549), .B(n15548), .Z(n15553) );
  NAND U16400 ( .A(n15551), .B(n15550), .Z(n15552) );
  NAND U16401 ( .A(n15553), .B(n15552), .Z(n15841) );
  XOR U16402 ( .A(n15840), .B(n15841), .Z(n15565) );
  NANDN U16403 ( .A(n15555), .B(n15554), .Z(n15559) );
  NAND U16404 ( .A(n15557), .B(n15556), .Z(n15558) );
  AND U16405 ( .A(n15559), .B(n15558), .Z(n15566) );
  XNOR U16406 ( .A(n15565), .B(n15566), .Z(n15567) );
  XNOR U16407 ( .A(n15568), .B(n15567), .Z(n15844) );
  XNOR U16408 ( .A(n15844), .B(sreg[146]), .Z(n15846) );
  NAND U16409 ( .A(n15560), .B(sreg[145]), .Z(n15564) );
  OR U16410 ( .A(n15562), .B(n15561), .Z(n15563) );
  AND U16411 ( .A(n15564), .B(n15563), .Z(n15845) );
  XOR U16412 ( .A(n15846), .B(n15845), .Z(c[146]) );
  NANDN U16413 ( .A(n15566), .B(n15565), .Z(n15570) );
  NAND U16414 ( .A(n15568), .B(n15567), .Z(n15569) );
  NAND U16415 ( .A(n15570), .B(n15569), .Z(n15852) );
  NANDN U16416 ( .A(n15572), .B(n15571), .Z(n15576) );
  NANDN U16417 ( .A(n15574), .B(n15573), .Z(n15575) );
  NAND U16418 ( .A(n15576), .B(n15575), .Z(n15855) );
  OR U16419 ( .A(n15578), .B(n15577), .Z(n15582) );
  NANDN U16420 ( .A(n15580), .B(n15579), .Z(n15581) );
  NAND U16421 ( .A(n15582), .B(n15581), .Z(n15856) );
  XNOR U16422 ( .A(n15855), .B(n15856), .Z(n15857) );
  OR U16423 ( .A(n15584), .B(n15583), .Z(n15588) );
  NAND U16424 ( .A(n15586), .B(n15585), .Z(n15587) );
  NAND U16425 ( .A(n15588), .B(n15587), .Z(n16127) );
  NANDN U16426 ( .A(n15590), .B(n15589), .Z(n15594) );
  NANDN U16427 ( .A(n15592), .B(n15591), .Z(n15593) );
  NAND U16428 ( .A(n15594), .B(n15593), .Z(n16128) );
  XNOR U16429 ( .A(n16127), .B(n16128), .Z(n16129) );
  NANDN U16430 ( .A(n15596), .B(n15595), .Z(n15600) );
  NAND U16431 ( .A(n15598), .B(n15597), .Z(n15599) );
  NAND U16432 ( .A(n15600), .B(n15599), .Z(n16106) );
  NANDN U16433 ( .A(n15602), .B(n15601), .Z(n15606) );
  OR U16434 ( .A(n15604), .B(n15603), .Z(n15605) );
  NAND U16435 ( .A(n15606), .B(n15605), .Z(n16108) );
  NANDN U16436 ( .A(n15608), .B(n15607), .Z(n15612) );
  NAND U16437 ( .A(n15610), .B(n15609), .Z(n15611) );
  AND U16438 ( .A(n15612), .B(n15611), .Z(n16107) );
  XOR U16439 ( .A(n16108), .B(n16107), .Z(n15613) );
  XOR U16440 ( .A(n16106), .B(n15613), .Z(n16094) );
  NANDN U16441 ( .A(n15615), .B(n15614), .Z(n15619) );
  OR U16442 ( .A(n15617), .B(n15616), .Z(n15618) );
  NAND U16443 ( .A(n15619), .B(n15618), .Z(n16095) );
  XOR U16444 ( .A(n16094), .B(n16095), .Z(n16097) );
  XOR U16445 ( .A(b[37]), .B(n23149), .Z(n15903) );
  NANDN U16446 ( .A(n15903), .B(n36311), .Z(n15626) );
  NANDN U16447 ( .A(n15624), .B(n36309), .Z(n15625) );
  NAND U16448 ( .A(n15626), .B(n15625), .Z(n15982) );
  XNOR U16449 ( .A(a[79]), .B(b[5]), .Z(n15906) );
  OR U16450 ( .A(n15906), .B(n29363), .Z(n15629) );
  NANDN U16451 ( .A(n15627), .B(n29864), .Z(n15628) );
  NAND U16452 ( .A(n15629), .B(n15628), .Z(n15979) );
  XNOR U16453 ( .A(a[81]), .B(n967), .Z(n15909) );
  NAND U16454 ( .A(n15909), .B(n28939), .Z(n15632) );
  NAND U16455 ( .A(n28938), .B(n15630), .Z(n15631) );
  AND U16456 ( .A(n15632), .B(n15631), .Z(n15980) );
  XNOR U16457 ( .A(n15979), .B(n15980), .Z(n15981) );
  XNOR U16458 ( .A(n15982), .B(n15981), .Z(n15882) );
  XOR U16459 ( .A(b[13]), .B(n30543), .Z(n15912) );
  OR U16460 ( .A(n15912), .B(n31550), .Z(n15635) );
  NANDN U16461 ( .A(n15633), .B(n31874), .Z(n15634) );
  NAND U16462 ( .A(n15635), .B(n15634), .Z(n16067) );
  NAND U16463 ( .A(n34848), .B(n15636), .Z(n15638) );
  XOR U16464 ( .A(n35375), .B(n26122), .Z(n15915) );
  NAND U16465 ( .A(n34618), .B(n15915), .Z(n15637) );
  NAND U16466 ( .A(n15638), .B(n15637), .Z(n16064) );
  NAND U16467 ( .A(n35188), .B(n15639), .Z(n15641) );
  XOR U16468 ( .A(n35540), .B(n25466), .Z(n15918) );
  NANDN U16469 ( .A(n34968), .B(n15918), .Z(n15640) );
  AND U16470 ( .A(n15641), .B(n15640), .Z(n16065) );
  XNOR U16471 ( .A(n16064), .B(n16065), .Z(n16066) );
  XNOR U16472 ( .A(n16067), .B(n16066), .Z(n15879) );
  NANDN U16473 ( .A(n15643), .B(n15642), .Z(n15647) );
  NAND U16474 ( .A(n15645), .B(n15644), .Z(n15646) );
  NAND U16475 ( .A(n15647), .B(n15646), .Z(n15880) );
  XNOR U16476 ( .A(n15879), .B(n15880), .Z(n15881) );
  XOR U16477 ( .A(n15882), .B(n15881), .Z(n15892) );
  NANDN U16478 ( .A(n15649), .B(n15648), .Z(n15653) );
  NAND U16479 ( .A(n15651), .B(n15650), .Z(n15652) );
  NAND U16480 ( .A(n15653), .B(n15652), .Z(n16023) );
  NAND U16481 ( .A(a[19]), .B(b[63]), .Z(n16037) );
  NANDN U16482 ( .A(n15654), .B(n38369), .Z(n15656) );
  XOR U16483 ( .A(b[61]), .B(n16269), .Z(n15933) );
  OR U16484 ( .A(n15933), .B(n38371), .Z(n15655) );
  NAND U16485 ( .A(n15656), .B(n15655), .Z(n16035) );
  NANDN U16486 ( .A(n15657), .B(n35311), .Z(n15659) );
  XOR U16487 ( .A(b[31]), .B(n25001), .Z(n15936) );
  NANDN U16488 ( .A(n15936), .B(n35313), .Z(n15658) );
  AND U16489 ( .A(n15659), .B(n15658), .Z(n16034) );
  XNOR U16490 ( .A(n16035), .B(n16034), .Z(n16036) );
  XOR U16491 ( .A(n16037), .B(n16036), .Z(n16021) );
  NAND U16492 ( .A(n33283), .B(n15660), .Z(n15662) );
  XOR U16493 ( .A(n33020), .B(n28403), .Z(n15939) );
  NANDN U16494 ( .A(n33021), .B(n15939), .Z(n15661) );
  NAND U16495 ( .A(n15662), .B(n15661), .Z(n15970) );
  XOR U16496 ( .A(b[21]), .B(a[63]), .Z(n15942) );
  NANDN U16497 ( .A(n33634), .B(n15942), .Z(n15665) );
  NAND U16498 ( .A(n15663), .B(n33464), .Z(n15664) );
  NAND U16499 ( .A(n15665), .B(n15664), .Z(n15967) );
  NAND U16500 ( .A(n34044), .B(n15666), .Z(n15668) );
  XOR U16501 ( .A(n34510), .B(n27773), .Z(n15945) );
  NANDN U16502 ( .A(n33867), .B(n15945), .Z(n15667) );
  AND U16503 ( .A(n15668), .B(n15667), .Z(n15968) );
  XNOR U16504 ( .A(n15967), .B(n15968), .Z(n15969) );
  XNOR U16505 ( .A(n15970), .B(n15969), .Z(n16022) );
  XNOR U16506 ( .A(n16021), .B(n16022), .Z(n16024) );
  XNOR U16507 ( .A(n16023), .B(n16024), .Z(n15891) );
  XOR U16508 ( .A(n15892), .B(n15891), .Z(n15894) );
  XNOR U16509 ( .A(n15893), .B(n15894), .Z(n15994) );
  NANDN U16510 ( .A(n15670), .B(n15669), .Z(n15674) );
  NAND U16511 ( .A(n15672), .B(n15671), .Z(n15673) );
  NAND U16512 ( .A(n15674), .B(n15673), .Z(n16085) );
  XNOR U16513 ( .A(b[41]), .B(a[43]), .Z(n15948) );
  OR U16514 ( .A(n15948), .B(n36905), .Z(n15677) );
  NANDN U16515 ( .A(n15675), .B(n36807), .Z(n15676) );
  NAND U16516 ( .A(n15677), .B(n15676), .Z(n15976) );
  XOR U16517 ( .A(b[57]), .B(n17960), .Z(n15951) );
  OR U16518 ( .A(n15951), .B(n965), .Z(n15680) );
  NANDN U16519 ( .A(n15678), .B(n38194), .Z(n15679) );
  NAND U16520 ( .A(n15680), .B(n15679), .Z(n15973) );
  NAND U16521 ( .A(n38326), .B(n15681), .Z(n15683) );
  XOR U16522 ( .A(n38400), .B(n16916), .Z(n15954) );
  NANDN U16523 ( .A(n38273), .B(n15954), .Z(n15682) );
  AND U16524 ( .A(n15683), .B(n15682), .Z(n15974) );
  XNOR U16525 ( .A(n15973), .B(n15974), .Z(n15975) );
  XOR U16526 ( .A(n15976), .B(n15975), .Z(n16082) );
  XOR U16527 ( .A(b[33]), .B(n24288), .Z(n15957) );
  NANDN U16528 ( .A(n15957), .B(n35620), .Z(n15686) );
  NANDN U16529 ( .A(n15684), .B(n35621), .Z(n15685) );
  NAND U16530 ( .A(n15686), .B(n15685), .Z(n16079) );
  NANDN U16531 ( .A(n966), .B(a[83]), .Z(n15687) );
  XOR U16532 ( .A(n29232), .B(n15687), .Z(n15689) );
  IV U16533 ( .A(a[82]), .Z(n32815) );
  NANDN U16534 ( .A(n32815), .B(n966), .Z(n15688) );
  AND U16535 ( .A(n15689), .B(n15688), .Z(n16076) );
  XOR U16536 ( .A(b[63]), .B(n16220), .Z(n15964) );
  NANDN U16537 ( .A(n15964), .B(n38422), .Z(n15692) );
  NANDN U16538 ( .A(n15690), .B(n38423), .Z(n15691) );
  AND U16539 ( .A(n15692), .B(n15691), .Z(n16077) );
  XNOR U16540 ( .A(n16076), .B(n16077), .Z(n16078) );
  XOR U16541 ( .A(n16079), .B(n16078), .Z(n16083) );
  XNOR U16542 ( .A(n16082), .B(n16083), .Z(n16084) );
  XNOR U16543 ( .A(n16085), .B(n16084), .Z(n15888) );
  NANDN U16544 ( .A(n15694), .B(n15693), .Z(n15698) );
  NAND U16545 ( .A(n15696), .B(n15695), .Z(n15697) );
  NAND U16546 ( .A(n15698), .B(n15697), .Z(n15885) );
  NANDN U16547 ( .A(n15700), .B(n15699), .Z(n15704) );
  NAND U16548 ( .A(n15702), .B(n15701), .Z(n15703) );
  AND U16549 ( .A(n15704), .B(n15703), .Z(n15886) );
  XNOR U16550 ( .A(n15885), .B(n15886), .Z(n15887) );
  XOR U16551 ( .A(n15888), .B(n15887), .Z(n15992) );
  NANDN U16552 ( .A(n15706), .B(n15705), .Z(n15710) );
  OR U16553 ( .A(n15708), .B(n15707), .Z(n15709) );
  AND U16554 ( .A(n15710), .B(n15709), .Z(n15991) );
  XOR U16555 ( .A(n15992), .B(n15991), .Z(n15993) );
  XNOR U16556 ( .A(n15994), .B(n15993), .Z(n16096) );
  XNOR U16557 ( .A(n16097), .B(n16096), .Z(n15861) );
  OR U16558 ( .A(n15712), .B(n15711), .Z(n15716) );
  NAND U16559 ( .A(n15714), .B(n15713), .Z(n15715) );
  NAND U16560 ( .A(n15716), .B(n15715), .Z(n16118) );
  XNOR U16561 ( .A(b[15]), .B(a[69]), .Z(n16046) );
  OR U16562 ( .A(n16046), .B(n32010), .Z(n15719) );
  NANDN U16563 ( .A(n15717), .B(n32011), .Z(n15718) );
  NAND U16564 ( .A(n15719), .B(n15718), .Z(n15930) );
  XOR U16565 ( .A(b[25]), .B(a[59]), .Z(n16049) );
  NANDN U16566 ( .A(n34219), .B(n16049), .Z(n15722) );
  NAND U16567 ( .A(n34217), .B(n15720), .Z(n15721) );
  NAND U16568 ( .A(n15722), .B(n15721), .Z(n15927) );
  XNOR U16569 ( .A(b[17]), .B(a[67]), .Z(n16052) );
  NANDN U16570 ( .A(n16052), .B(n32543), .Z(n15725) );
  NANDN U16571 ( .A(n15723), .B(n32541), .Z(n15724) );
  AND U16572 ( .A(n15725), .B(n15724), .Z(n15928) );
  XNOR U16573 ( .A(n15927), .B(n15928), .Z(n15929) );
  XNOR U16574 ( .A(n15930), .B(n15929), .Z(n15985) );
  XOR U16575 ( .A(b[39]), .B(n22579), .Z(n16055) );
  NANDN U16576 ( .A(n16055), .B(n36553), .Z(n15728) );
  NANDN U16577 ( .A(n15726), .B(n36643), .Z(n15727) );
  NAND U16578 ( .A(n15728), .B(n15727), .Z(n15924) );
  XOR U16579 ( .A(b[51]), .B(n19656), .Z(n16058) );
  NANDN U16580 ( .A(n16058), .B(n37803), .Z(n15731) );
  NANDN U16581 ( .A(n15729), .B(n37802), .Z(n15730) );
  NAND U16582 ( .A(n15731), .B(n15730), .Z(n15921) );
  XOR U16583 ( .A(b[53]), .B(n18639), .Z(n16061) );
  NANDN U16584 ( .A(n16061), .B(n37940), .Z(n15734) );
  NANDN U16585 ( .A(n15732), .B(n37941), .Z(n15733) );
  AND U16586 ( .A(n15734), .B(n15733), .Z(n15922) );
  XNOR U16587 ( .A(n15921), .B(n15922), .Z(n15923) );
  XOR U16588 ( .A(n15924), .B(n15923), .Z(n15986) );
  XOR U16589 ( .A(n15985), .B(n15986), .Z(n15988) );
  NANDN U16590 ( .A(n15736), .B(n15735), .Z(n15740) );
  NAND U16591 ( .A(n15738), .B(n15737), .Z(n15739) );
  NAND U16592 ( .A(n15740), .B(n15739), .Z(n15987) );
  XNOR U16593 ( .A(n15988), .B(n15987), .Z(n16091) );
  NANDN U16594 ( .A(n15742), .B(n15741), .Z(n15746) );
  NAND U16595 ( .A(n15744), .B(n15743), .Z(n15745) );
  NAND U16596 ( .A(n15746), .B(n15745), .Z(n16088) );
  NANDN U16597 ( .A(n15748), .B(n15747), .Z(n15752) );
  NAND U16598 ( .A(n15750), .B(n15749), .Z(n15751) );
  AND U16599 ( .A(n15752), .B(n15751), .Z(n16089) );
  XNOR U16600 ( .A(n16088), .B(n16089), .Z(n16090) );
  XNOR U16601 ( .A(n16091), .B(n16090), .Z(n16109) );
  OR U16602 ( .A(n15754), .B(n15753), .Z(n15758) );
  OR U16603 ( .A(n15756), .B(n15755), .Z(n15757) );
  AND U16604 ( .A(n15758), .B(n15757), .Z(n16110) );
  XNOR U16605 ( .A(n16109), .B(n16110), .Z(n16111) );
  NANDN U16606 ( .A(n15760), .B(n15759), .Z(n15764) );
  NAND U16607 ( .A(n15762), .B(n15761), .Z(n15763) );
  AND U16608 ( .A(n15764), .B(n15763), .Z(n16112) );
  XNOR U16609 ( .A(n16111), .B(n16112), .Z(n16116) );
  XNOR U16610 ( .A(b[11]), .B(a[73]), .Z(n15997) );
  OR U16611 ( .A(n15997), .B(n31369), .Z(n15767) );
  NANDN U16612 ( .A(n15765), .B(n31119), .Z(n15766) );
  NAND U16613 ( .A(n15767), .B(n15766), .Z(n16018) );
  XOR U16614 ( .A(b[43]), .B(n21441), .Z(n16000) );
  NANDN U16615 ( .A(n16000), .B(n37068), .Z(n15770) );
  NANDN U16616 ( .A(n15768), .B(n37069), .Z(n15769) );
  NAND U16617 ( .A(n15770), .B(n15769), .Z(n16015) );
  XNOR U16618 ( .A(b[45]), .B(a[39]), .Z(n16003) );
  NANDN U16619 ( .A(n16003), .B(n37261), .Z(n15773) );
  NANDN U16620 ( .A(n15771), .B(n37262), .Z(n15772) );
  AND U16621 ( .A(n15773), .B(n15772), .Z(n16016) );
  XNOR U16622 ( .A(n16015), .B(n16016), .Z(n16017) );
  XNOR U16623 ( .A(n16018), .B(n16017), .Z(n15897) );
  XOR U16624 ( .A(b[49]), .B(n20315), .Z(n16006) );
  OR U16625 ( .A(n16006), .B(n37756), .Z(n15776) );
  NANDN U16626 ( .A(n15774), .B(n37652), .Z(n15775) );
  NAND U16627 ( .A(n15776), .B(n15775), .Z(n16043) );
  NAND U16628 ( .A(n37469), .B(n15777), .Z(n15779) );
  XOR U16629 ( .A(n978), .B(n20352), .Z(n16009) );
  NAND U16630 ( .A(n16009), .B(n37471), .Z(n15778) );
  NAND U16631 ( .A(n15779), .B(n15778), .Z(n16040) );
  XNOR U16632 ( .A(b[9]), .B(a[75]), .Z(n16012) );
  NANDN U16633 ( .A(n16012), .B(n30509), .Z(n15782) );
  NANDN U16634 ( .A(n15780), .B(n30846), .Z(n15781) );
  AND U16635 ( .A(n15782), .B(n15781), .Z(n16041) );
  XNOR U16636 ( .A(n16040), .B(n16041), .Z(n16042) );
  XOR U16637 ( .A(n16043), .B(n16042), .Z(n15898) );
  XNOR U16638 ( .A(n15897), .B(n15898), .Z(n15899) );
  NANDN U16639 ( .A(n15784), .B(n15783), .Z(n15788) );
  NAND U16640 ( .A(n15786), .B(n15785), .Z(n15787) );
  AND U16641 ( .A(n15788), .B(n15787), .Z(n15900) );
  XNOR U16642 ( .A(n15899), .B(n15900), .Z(n16101) );
  XNOR U16643 ( .A(n16101), .B(n16100), .Z(n16102) );
  XNOR U16644 ( .A(b[35]), .B(a[49]), .Z(n16025) );
  NANDN U16645 ( .A(n16025), .B(n35985), .Z(n15795) );
  NANDN U16646 ( .A(n15793), .B(n35986), .Z(n15794) );
  NAND U16647 ( .A(n15795), .B(n15794), .Z(n16073) );
  XNOR U16648 ( .A(a[77]), .B(n31123), .Z(n16028) );
  NAND U16649 ( .A(n16028), .B(n29949), .Z(n15798) );
  NAND U16650 ( .A(n29948), .B(n15796), .Z(n15797) );
  NAND U16651 ( .A(n15798), .B(n15797), .Z(n16070) );
  XOR U16652 ( .A(b[55]), .B(n18003), .Z(n16031) );
  NANDN U16653 ( .A(n16031), .B(n38075), .Z(n15801) );
  NANDN U16654 ( .A(n15799), .B(n38073), .Z(n15800) );
  AND U16655 ( .A(n15801), .B(n15800), .Z(n16071) );
  XNOR U16656 ( .A(n16070), .B(n16071), .Z(n16072) );
  XNOR U16657 ( .A(n16073), .B(n16072), .Z(n15876) );
  NANDN U16658 ( .A(n15803), .B(n15802), .Z(n15807) );
  NAND U16659 ( .A(n15805), .B(n15804), .Z(n15806) );
  NAND U16660 ( .A(n15807), .B(n15806), .Z(n15873) );
  NANDN U16661 ( .A(n15809), .B(n15808), .Z(n15813) );
  NAND U16662 ( .A(n15811), .B(n15810), .Z(n15812) );
  NAND U16663 ( .A(n15813), .B(n15812), .Z(n15874) );
  XNOR U16664 ( .A(n15873), .B(n15874), .Z(n15875) );
  XOR U16665 ( .A(n15876), .B(n15875), .Z(n16103) );
  XOR U16666 ( .A(n16102), .B(n16103), .Z(n16115) );
  XNOR U16667 ( .A(n16116), .B(n16115), .Z(n16117) );
  XOR U16668 ( .A(n16118), .B(n16117), .Z(n15862) );
  XNOR U16669 ( .A(n15861), .B(n15862), .Z(n15863) );
  NAND U16670 ( .A(n15815), .B(n15814), .Z(n15819) );
  NANDN U16671 ( .A(n15817), .B(n15816), .Z(n15818) );
  NAND U16672 ( .A(n15819), .B(n15818), .Z(n15864) );
  XOR U16673 ( .A(n15863), .B(n15864), .Z(n16124) );
  NAND U16674 ( .A(n15821), .B(n15820), .Z(n15825) );
  NANDN U16675 ( .A(n15823), .B(n15822), .Z(n15824) );
  NAND U16676 ( .A(n15825), .B(n15824), .Z(n15870) );
  XNOR U16677 ( .A(n15868), .B(n15867), .Z(n15869) );
  XOR U16678 ( .A(n15870), .B(n15869), .Z(n16121) );
  XNOR U16679 ( .A(n16121), .B(n16122), .Z(n16123) );
  XOR U16680 ( .A(n16124), .B(n16123), .Z(n16130) );
  XOR U16681 ( .A(n16129), .B(n16130), .Z(n15858) );
  XOR U16682 ( .A(n15857), .B(n15858), .Z(n15849) );
  OR U16683 ( .A(n15839), .B(n15838), .Z(n15843) );
  NANDN U16684 ( .A(n15841), .B(n15840), .Z(n15842) );
  AND U16685 ( .A(n15843), .B(n15842), .Z(n15850) );
  XOR U16686 ( .A(n15849), .B(n15850), .Z(n15851) );
  XNOR U16687 ( .A(n15852), .B(n15851), .Z(n16133) );
  XNOR U16688 ( .A(n16133), .B(sreg[147]), .Z(n16135) );
  NAND U16689 ( .A(n15844), .B(sreg[146]), .Z(n15848) );
  OR U16690 ( .A(n15846), .B(n15845), .Z(n15847) );
  AND U16691 ( .A(n15848), .B(n15847), .Z(n16134) );
  XOR U16692 ( .A(n16135), .B(n16134), .Z(c[147]) );
  NAND U16693 ( .A(n15850), .B(n15849), .Z(n15854) );
  NAND U16694 ( .A(n15852), .B(n15851), .Z(n15853) );
  NAND U16695 ( .A(n15854), .B(n15853), .Z(n16141) );
  NANDN U16696 ( .A(n15856), .B(n15855), .Z(n15860) );
  NAND U16697 ( .A(n15858), .B(n15857), .Z(n15859) );
  NAND U16698 ( .A(n15860), .B(n15859), .Z(n16138) );
  NANDN U16699 ( .A(n15862), .B(n15861), .Z(n15866) );
  NANDN U16700 ( .A(n15864), .B(n15863), .Z(n15865) );
  NAND U16701 ( .A(n15866), .B(n15865), .Z(n16407) );
  NANDN U16702 ( .A(n15868), .B(n15867), .Z(n15872) );
  NANDN U16703 ( .A(n15870), .B(n15869), .Z(n15871) );
  AND U16704 ( .A(n15872), .B(n15871), .Z(n16406) );
  XNOR U16705 ( .A(n16407), .B(n16406), .Z(n16408) );
  NANDN U16706 ( .A(n15874), .B(n15873), .Z(n15878) );
  NAND U16707 ( .A(n15876), .B(n15875), .Z(n15877) );
  AND U16708 ( .A(n15878), .B(n15877), .Z(n16153) );
  NANDN U16709 ( .A(n15880), .B(n15879), .Z(n15884) );
  NAND U16710 ( .A(n15882), .B(n15881), .Z(n15883) );
  NAND U16711 ( .A(n15884), .B(n15883), .Z(n16150) );
  NANDN U16712 ( .A(n15886), .B(n15885), .Z(n15890) );
  NAND U16713 ( .A(n15888), .B(n15887), .Z(n15889) );
  NAND U16714 ( .A(n15890), .B(n15889), .Z(n16151) );
  XNOR U16715 ( .A(n16150), .B(n16151), .Z(n16152) );
  XNOR U16716 ( .A(n16153), .B(n16152), .Z(n16382) );
  NANDN U16717 ( .A(n15892), .B(n15891), .Z(n15896) );
  OR U16718 ( .A(n15894), .B(n15893), .Z(n15895) );
  AND U16719 ( .A(n15896), .B(n15895), .Z(n16383) );
  XNOR U16720 ( .A(n16382), .B(n16383), .Z(n16385) );
  NANDN U16721 ( .A(n15898), .B(n15897), .Z(n15902) );
  NAND U16722 ( .A(n15900), .B(n15899), .Z(n15901) );
  NAND U16723 ( .A(n15902), .B(n15901), .Z(n16183) );
  XOR U16724 ( .A(b[37]), .B(n23447), .Z(n16190) );
  NANDN U16725 ( .A(n16190), .B(n36311), .Z(n15905) );
  NANDN U16726 ( .A(n15903), .B(n36309), .Z(n15904) );
  NAND U16727 ( .A(n15905), .B(n15904), .Z(n16245) );
  XOR U16728 ( .A(a[80]), .B(n968), .Z(n16193) );
  OR U16729 ( .A(n16193), .B(n29363), .Z(n15908) );
  NANDN U16730 ( .A(n15906), .B(n29864), .Z(n15907) );
  NAND U16731 ( .A(n15908), .B(n15907), .Z(n16242) );
  XOR U16732 ( .A(n32815), .B(n967), .Z(n16196) );
  NAND U16733 ( .A(n16196), .B(n28939), .Z(n15911) );
  NAND U16734 ( .A(n28938), .B(n15909), .Z(n15910) );
  AND U16735 ( .A(n15911), .B(n15910), .Z(n16243) );
  XNOR U16736 ( .A(n16242), .B(n16243), .Z(n16244) );
  XNOR U16737 ( .A(n16245), .B(n16244), .Z(n16162) );
  XOR U16738 ( .A(b[13]), .B(n30210), .Z(n16199) );
  OR U16739 ( .A(n16199), .B(n31550), .Z(n15914) );
  NANDN U16740 ( .A(n15912), .B(n31874), .Z(n15913) );
  NAND U16741 ( .A(n15914), .B(n15913), .Z(n16373) );
  NAND U16742 ( .A(n34848), .B(n15915), .Z(n15917) );
  XOR U16743 ( .A(n35375), .B(n26347), .Z(n16202) );
  NAND U16744 ( .A(n34618), .B(n16202), .Z(n15916) );
  NAND U16745 ( .A(n15917), .B(n15916), .Z(n16370) );
  NAND U16746 ( .A(n35188), .B(n15918), .Z(n15920) );
  XOR U16747 ( .A(n35540), .B(n25860), .Z(n16205) );
  NANDN U16748 ( .A(n34968), .B(n16205), .Z(n15919) );
  AND U16749 ( .A(n15920), .B(n15919), .Z(n16371) );
  XNOR U16750 ( .A(n16370), .B(n16371), .Z(n16372) );
  XOR U16751 ( .A(n16373), .B(n16372), .Z(n16163) );
  XOR U16752 ( .A(n16162), .B(n16163), .Z(n16165) );
  NANDN U16753 ( .A(n15922), .B(n15921), .Z(n15926) );
  NAND U16754 ( .A(n15924), .B(n15923), .Z(n15925) );
  NAND U16755 ( .A(n15926), .B(n15925), .Z(n16164) );
  XNOR U16756 ( .A(n16165), .B(n16164), .Z(n16181) );
  NANDN U16757 ( .A(n15928), .B(n15927), .Z(n15932) );
  NAND U16758 ( .A(n15930), .B(n15929), .Z(n15931) );
  NAND U16759 ( .A(n15932), .B(n15931), .Z(n16311) );
  NAND U16760 ( .A(a[20]), .B(b[63]), .Z(n16325) );
  NANDN U16761 ( .A(n15933), .B(n38369), .Z(n15935) );
  XOR U16762 ( .A(b[61]), .B(n16508), .Z(n16221) );
  OR U16763 ( .A(n16221), .B(n38371), .Z(n15934) );
  NAND U16764 ( .A(n15935), .B(n15934), .Z(n16323) );
  NANDN U16765 ( .A(n15936), .B(n35311), .Z(n15938) );
  XOR U16766 ( .A(b[31]), .B(n25177), .Z(n16224) );
  NANDN U16767 ( .A(n16224), .B(n35313), .Z(n15937) );
  AND U16768 ( .A(n15938), .B(n15937), .Z(n16322) );
  XNOR U16769 ( .A(n16323), .B(n16322), .Z(n16324) );
  XOR U16770 ( .A(n16325), .B(n16324), .Z(n16309) );
  NAND U16771 ( .A(n33283), .B(n15939), .Z(n15941) );
  XOR U16772 ( .A(n33020), .B(n28701), .Z(n16227) );
  NANDN U16773 ( .A(n33021), .B(n16227), .Z(n15940) );
  NAND U16774 ( .A(n15941), .B(n15940), .Z(n16251) );
  XOR U16775 ( .A(b[21]), .B(a[64]), .Z(n16230) );
  NANDN U16776 ( .A(n33634), .B(n16230), .Z(n15944) );
  NAND U16777 ( .A(n15942), .B(n33464), .Z(n15943) );
  NAND U16778 ( .A(n15944), .B(n15943), .Z(n16248) );
  NAND U16779 ( .A(n34044), .B(n15945), .Z(n15947) );
  XNOR U16780 ( .A(n34510), .B(a[62]), .Z(n16233) );
  NANDN U16781 ( .A(n33867), .B(n16233), .Z(n15946) );
  AND U16782 ( .A(n15947), .B(n15946), .Z(n16249) );
  XNOR U16783 ( .A(n16248), .B(n16249), .Z(n16250) );
  XNOR U16784 ( .A(n16251), .B(n16250), .Z(n16310) );
  XNOR U16785 ( .A(n16309), .B(n16310), .Z(n16312) );
  XNOR U16786 ( .A(n16311), .B(n16312), .Z(n16180) );
  XNOR U16787 ( .A(n16181), .B(n16180), .Z(n16182) );
  XNOR U16788 ( .A(n16183), .B(n16182), .Z(n16282) );
  XNOR U16789 ( .A(b[41]), .B(a[44]), .Z(n16254) );
  OR U16790 ( .A(n16254), .B(n36905), .Z(n15950) );
  NANDN U16791 ( .A(n15948), .B(n36807), .Z(n15949) );
  NAND U16792 ( .A(n15950), .B(n15949), .Z(n16276) );
  XOR U16793 ( .A(b[57]), .B(n17702), .Z(n16257) );
  OR U16794 ( .A(n16257), .B(n965), .Z(n15953) );
  NANDN U16795 ( .A(n15951), .B(n38194), .Z(n15952) );
  NAND U16796 ( .A(n15953), .B(n15952), .Z(n16273) );
  NAND U16797 ( .A(n38326), .B(n15954), .Z(n15956) );
  XOR U16798 ( .A(n38400), .B(n17133), .Z(n16260) );
  NANDN U16799 ( .A(n38273), .B(n16260), .Z(n15955) );
  AND U16800 ( .A(n15956), .B(n15955), .Z(n16274) );
  XNOR U16801 ( .A(n16273), .B(n16274), .Z(n16275) );
  XOR U16802 ( .A(n16276), .B(n16275), .Z(n16334) );
  XOR U16803 ( .A(b[33]), .B(n25134), .Z(n16263) );
  NANDN U16804 ( .A(n16263), .B(n35620), .Z(n15959) );
  NANDN U16805 ( .A(n15957), .B(n35621), .Z(n15958) );
  NAND U16806 ( .A(n15959), .B(n15958), .Z(n16349) );
  NANDN U16807 ( .A(n966), .B(a[84]), .Z(n15960) );
  XOR U16808 ( .A(n29232), .B(n15960), .Z(n15962) );
  NANDN U16809 ( .A(b[0]), .B(a[83]), .Z(n15961) );
  AND U16810 ( .A(n15962), .B(n15961), .Z(n16346) );
  XOR U16811 ( .A(b[63]), .B(n15963), .Z(n16270) );
  NANDN U16812 ( .A(n16270), .B(n38422), .Z(n15966) );
  NANDN U16813 ( .A(n15964), .B(n38423), .Z(n15965) );
  AND U16814 ( .A(n15966), .B(n15965), .Z(n16347) );
  XNOR U16815 ( .A(n16346), .B(n16347), .Z(n16348) );
  XOR U16816 ( .A(n16349), .B(n16348), .Z(n16335) );
  XNOR U16817 ( .A(n16334), .B(n16335), .Z(n16337) );
  NANDN U16818 ( .A(n15968), .B(n15967), .Z(n15972) );
  NAND U16819 ( .A(n15970), .B(n15969), .Z(n15971) );
  NAND U16820 ( .A(n15972), .B(n15971), .Z(n16336) );
  XNOR U16821 ( .A(n16337), .B(n16336), .Z(n16177) );
  NANDN U16822 ( .A(n15974), .B(n15973), .Z(n15978) );
  NAND U16823 ( .A(n15976), .B(n15975), .Z(n15977) );
  NAND U16824 ( .A(n15978), .B(n15977), .Z(n16174) );
  NANDN U16825 ( .A(n15980), .B(n15979), .Z(n15984) );
  NAND U16826 ( .A(n15982), .B(n15981), .Z(n15983) );
  AND U16827 ( .A(n15984), .B(n15983), .Z(n16175) );
  XNOR U16828 ( .A(n16174), .B(n16175), .Z(n16176) );
  XOR U16829 ( .A(n16177), .B(n16176), .Z(n16280) );
  NANDN U16830 ( .A(n15986), .B(n15985), .Z(n15990) );
  OR U16831 ( .A(n15988), .B(n15987), .Z(n15989) );
  AND U16832 ( .A(n15990), .B(n15989), .Z(n16279) );
  XOR U16833 ( .A(n16280), .B(n16279), .Z(n16281) );
  XNOR U16834 ( .A(n16282), .B(n16281), .Z(n16384) );
  XNOR U16835 ( .A(n16385), .B(n16384), .Z(n16388) );
  OR U16836 ( .A(n15992), .B(n15991), .Z(n15996) );
  NAND U16837 ( .A(n15994), .B(n15993), .Z(n15995) );
  NAND U16838 ( .A(n15996), .B(n15995), .Z(n16161) );
  XOR U16839 ( .A(b[11]), .B(n31372), .Z(n16294) );
  OR U16840 ( .A(n16294), .B(n31369), .Z(n15999) );
  NANDN U16841 ( .A(n15997), .B(n31119), .Z(n15998) );
  NAND U16842 ( .A(n15999), .B(n15998), .Z(n16306) );
  XOR U16843 ( .A(b[43]), .B(n22246), .Z(n16297) );
  NANDN U16844 ( .A(n16297), .B(n37068), .Z(n16002) );
  NANDN U16845 ( .A(n16000), .B(n37069), .Z(n16001) );
  NAND U16846 ( .A(n16002), .B(n16001), .Z(n16303) );
  XNOR U16847 ( .A(b[45]), .B(a[40]), .Z(n16300) );
  NANDN U16848 ( .A(n16300), .B(n37261), .Z(n16005) );
  NANDN U16849 ( .A(n16003), .B(n37262), .Z(n16004) );
  AND U16850 ( .A(n16005), .B(n16004), .Z(n16304) );
  XNOR U16851 ( .A(n16303), .B(n16304), .Z(n16305) );
  XNOR U16852 ( .A(n16306), .B(n16305), .Z(n16189) );
  XOR U16853 ( .A(b[49]), .B(n19980), .Z(n16285) );
  OR U16854 ( .A(n16285), .B(n37756), .Z(n16008) );
  NANDN U16855 ( .A(n16006), .B(n37652), .Z(n16007) );
  NAND U16856 ( .A(n16008), .B(n16007), .Z(n16331) );
  NAND U16857 ( .A(n37469), .B(n16009), .Z(n16011) );
  XOR U16858 ( .A(n978), .B(n20686), .Z(n16288) );
  NAND U16859 ( .A(n16288), .B(n37471), .Z(n16010) );
  NAND U16860 ( .A(n16011), .B(n16010), .Z(n16328) );
  XOR U16861 ( .A(a[76]), .B(n969), .Z(n16291) );
  NANDN U16862 ( .A(n16291), .B(n30509), .Z(n16014) );
  NANDN U16863 ( .A(n16012), .B(n30846), .Z(n16013) );
  AND U16864 ( .A(n16014), .B(n16013), .Z(n16329) );
  XNOR U16865 ( .A(n16328), .B(n16329), .Z(n16330) );
  XNOR U16866 ( .A(n16331), .B(n16330), .Z(n16186) );
  NANDN U16867 ( .A(n16016), .B(n16015), .Z(n16020) );
  NAND U16868 ( .A(n16018), .B(n16017), .Z(n16019) );
  NAND U16869 ( .A(n16020), .B(n16019), .Z(n16187) );
  XNOR U16870 ( .A(n16186), .B(n16187), .Z(n16188) );
  XOR U16871 ( .A(n16189), .B(n16188), .Z(n16144) );
  XNOR U16872 ( .A(n16144), .B(n16145), .Z(n16147) );
  XNOR U16873 ( .A(b[35]), .B(a[50]), .Z(n16313) );
  NANDN U16874 ( .A(n16313), .B(n35985), .Z(n16027) );
  NANDN U16875 ( .A(n16025), .B(n35986), .Z(n16026) );
  NAND U16876 ( .A(n16027), .B(n16026), .Z(n16379) );
  XOR U16877 ( .A(n31870), .B(n31123), .Z(n16316) );
  NAND U16878 ( .A(n16316), .B(n29949), .Z(n16030) );
  NAND U16879 ( .A(n29948), .B(n16028), .Z(n16029) );
  NAND U16880 ( .A(n16030), .B(n16029), .Z(n16376) );
  XOR U16881 ( .A(b[55]), .B(n18804), .Z(n16319) );
  NANDN U16882 ( .A(n16319), .B(n38075), .Z(n16033) );
  NANDN U16883 ( .A(n16031), .B(n38073), .Z(n16032) );
  AND U16884 ( .A(n16033), .B(n16032), .Z(n16377) );
  XNOR U16885 ( .A(n16376), .B(n16377), .Z(n16378) );
  XNOR U16886 ( .A(n16379), .B(n16378), .Z(n16171) );
  NANDN U16887 ( .A(n16035), .B(n16034), .Z(n16039) );
  NAND U16888 ( .A(n16037), .B(n16036), .Z(n16038) );
  NAND U16889 ( .A(n16039), .B(n16038), .Z(n16168) );
  NANDN U16890 ( .A(n16041), .B(n16040), .Z(n16045) );
  NAND U16891 ( .A(n16043), .B(n16042), .Z(n16044) );
  NAND U16892 ( .A(n16045), .B(n16044), .Z(n16169) );
  XNOR U16893 ( .A(n16168), .B(n16169), .Z(n16170) );
  XOR U16894 ( .A(n16171), .B(n16170), .Z(n16146) );
  XNOR U16895 ( .A(n16147), .B(n16146), .Z(n16158) );
  XOR U16896 ( .A(b[15]), .B(n30379), .Z(n16352) );
  OR U16897 ( .A(n16352), .B(n32010), .Z(n16048) );
  NANDN U16898 ( .A(n16046), .B(n32011), .Z(n16047) );
  NAND U16899 ( .A(n16048), .B(n16047), .Z(n16217) );
  XNOR U16900 ( .A(b[25]), .B(n27436), .Z(n16355) );
  NANDN U16901 ( .A(n34219), .B(n16355), .Z(n16051) );
  NAND U16902 ( .A(n34217), .B(n16049), .Z(n16050) );
  NAND U16903 ( .A(n16051), .B(n16050), .Z(n16214) );
  XNOR U16904 ( .A(b[17]), .B(a[68]), .Z(n16358) );
  NANDN U16905 ( .A(n16358), .B(n32543), .Z(n16054) );
  NANDN U16906 ( .A(n16052), .B(n32541), .Z(n16053) );
  AND U16907 ( .A(n16054), .B(n16053), .Z(n16215) );
  XNOR U16908 ( .A(n16214), .B(n16215), .Z(n16216) );
  XNOR U16909 ( .A(n16217), .B(n16216), .Z(n16236) );
  XOR U16910 ( .A(b[39]), .B(n22964), .Z(n16361) );
  NANDN U16911 ( .A(n16361), .B(n36553), .Z(n16057) );
  NANDN U16912 ( .A(n16055), .B(n36643), .Z(n16056) );
  NAND U16913 ( .A(n16057), .B(n16056), .Z(n16211) );
  XOR U16914 ( .A(b[51]), .B(n19513), .Z(n16364) );
  NANDN U16915 ( .A(n16364), .B(n37803), .Z(n16060) );
  NANDN U16916 ( .A(n16058), .B(n37802), .Z(n16059) );
  NAND U16917 ( .A(n16060), .B(n16059), .Z(n16208) );
  XOR U16918 ( .A(b[53]), .B(n18841), .Z(n16367) );
  NANDN U16919 ( .A(n16367), .B(n37940), .Z(n16063) );
  NANDN U16920 ( .A(n16061), .B(n37941), .Z(n16062) );
  AND U16921 ( .A(n16063), .B(n16062), .Z(n16209) );
  XNOR U16922 ( .A(n16208), .B(n16209), .Z(n16210) );
  XOR U16923 ( .A(n16211), .B(n16210), .Z(n16237) );
  XNOR U16924 ( .A(n16236), .B(n16237), .Z(n16238) );
  NANDN U16925 ( .A(n16065), .B(n16064), .Z(n16069) );
  NAND U16926 ( .A(n16067), .B(n16066), .Z(n16068) );
  NAND U16927 ( .A(n16069), .B(n16068), .Z(n16239) );
  XOR U16928 ( .A(n16238), .B(n16239), .Z(n16343) );
  NANDN U16929 ( .A(n16071), .B(n16070), .Z(n16075) );
  NAND U16930 ( .A(n16073), .B(n16072), .Z(n16074) );
  NAND U16931 ( .A(n16075), .B(n16074), .Z(n16340) );
  NANDN U16932 ( .A(n16077), .B(n16076), .Z(n16081) );
  NAND U16933 ( .A(n16079), .B(n16078), .Z(n16080) );
  AND U16934 ( .A(n16081), .B(n16080), .Z(n16341) );
  XNOR U16935 ( .A(n16340), .B(n16341), .Z(n16342) );
  XNOR U16936 ( .A(n16343), .B(n16342), .Z(n16154) );
  OR U16937 ( .A(n16083), .B(n16082), .Z(n16087) );
  OR U16938 ( .A(n16085), .B(n16084), .Z(n16086) );
  AND U16939 ( .A(n16087), .B(n16086), .Z(n16155) );
  XNOR U16940 ( .A(n16154), .B(n16155), .Z(n16156) );
  NANDN U16941 ( .A(n16089), .B(n16088), .Z(n16093) );
  NAND U16942 ( .A(n16091), .B(n16090), .Z(n16092) );
  AND U16943 ( .A(n16093), .B(n16092), .Z(n16157) );
  XNOR U16944 ( .A(n16156), .B(n16157), .Z(n16159) );
  XNOR U16945 ( .A(n16158), .B(n16159), .Z(n16160) );
  XOR U16946 ( .A(n16161), .B(n16160), .Z(n16389) );
  XNOR U16947 ( .A(n16388), .B(n16389), .Z(n16390) );
  NANDN U16948 ( .A(n16095), .B(n16094), .Z(n16099) );
  OR U16949 ( .A(n16097), .B(n16096), .Z(n16098) );
  NAND U16950 ( .A(n16099), .B(n16098), .Z(n16391) );
  XOR U16951 ( .A(n16390), .B(n16391), .Z(n16403) );
  NANDN U16952 ( .A(n16101), .B(n16100), .Z(n16105) );
  NAND U16953 ( .A(n16103), .B(n16102), .Z(n16104) );
  NAND U16954 ( .A(n16105), .B(n16104), .Z(n16397) );
  NANDN U16955 ( .A(n16110), .B(n16109), .Z(n16114) );
  NAND U16956 ( .A(n16112), .B(n16111), .Z(n16113) );
  AND U16957 ( .A(n16114), .B(n16113), .Z(n16394) );
  XNOR U16958 ( .A(n16395), .B(n16394), .Z(n16396) );
  XOR U16959 ( .A(n16397), .B(n16396), .Z(n16400) );
  NANDN U16960 ( .A(n16116), .B(n16115), .Z(n16120) );
  NAND U16961 ( .A(n16118), .B(n16117), .Z(n16119) );
  AND U16962 ( .A(n16120), .B(n16119), .Z(n16401) );
  XNOR U16963 ( .A(n16400), .B(n16401), .Z(n16402) );
  XNOR U16964 ( .A(n16403), .B(n16402), .Z(n16409) );
  XOR U16965 ( .A(n16408), .B(n16409), .Z(n16412) );
  NANDN U16966 ( .A(n16122), .B(n16121), .Z(n16126) );
  NAND U16967 ( .A(n16124), .B(n16123), .Z(n16125) );
  NAND U16968 ( .A(n16126), .B(n16125), .Z(n16413) );
  XNOR U16969 ( .A(n16412), .B(n16413), .Z(n16414) );
  NANDN U16970 ( .A(n16128), .B(n16127), .Z(n16132) );
  NAND U16971 ( .A(n16130), .B(n16129), .Z(n16131) );
  NAND U16972 ( .A(n16132), .B(n16131), .Z(n16415) );
  XNOR U16973 ( .A(n16414), .B(n16415), .Z(n16139) );
  XNOR U16974 ( .A(n16138), .B(n16139), .Z(n16140) );
  XNOR U16975 ( .A(n16141), .B(n16140), .Z(n16418) );
  XNOR U16976 ( .A(n16418), .B(sreg[148]), .Z(n16420) );
  NAND U16977 ( .A(n16133), .B(sreg[147]), .Z(n16137) );
  OR U16978 ( .A(n16135), .B(n16134), .Z(n16136) );
  AND U16979 ( .A(n16137), .B(n16136), .Z(n16419) );
  XOR U16980 ( .A(n16420), .B(n16419), .Z(c[148]) );
  NANDN U16981 ( .A(n16139), .B(n16138), .Z(n16143) );
  NAND U16982 ( .A(n16141), .B(n16140), .Z(n16142) );
  NAND U16983 ( .A(n16143), .B(n16142), .Z(n16426) );
  NAND U16984 ( .A(n16145), .B(n16144), .Z(n16149) );
  NANDN U16985 ( .A(n16147), .B(n16146), .Z(n16148) );
  NAND U16986 ( .A(n16149), .B(n16148), .Z(n16679) );
  XNOR U16987 ( .A(n16676), .B(n16677), .Z(n16678) );
  XNOR U16988 ( .A(n16679), .B(n16678), .Z(n16688) );
  XNOR U16989 ( .A(n16688), .B(n16689), .Z(n16690) );
  NANDN U16990 ( .A(n16163), .B(n16162), .Z(n16167) );
  OR U16991 ( .A(n16165), .B(n16164), .Z(n16166) );
  AND U16992 ( .A(n16167), .B(n16166), .Z(n16675) );
  NANDN U16993 ( .A(n16169), .B(n16168), .Z(n16173) );
  NAND U16994 ( .A(n16171), .B(n16170), .Z(n16172) );
  NAND U16995 ( .A(n16173), .B(n16172), .Z(n16672) );
  NANDN U16996 ( .A(n16175), .B(n16174), .Z(n16179) );
  NAND U16997 ( .A(n16177), .B(n16176), .Z(n16178) );
  NAND U16998 ( .A(n16179), .B(n16178), .Z(n16673) );
  XNOR U16999 ( .A(n16672), .B(n16673), .Z(n16674) );
  XNOR U17000 ( .A(n16675), .B(n16674), .Z(n16650) );
  NAND U17001 ( .A(n16181), .B(n16180), .Z(n16185) );
  OR U17002 ( .A(n16183), .B(n16182), .Z(n16184) );
  AND U17003 ( .A(n16185), .B(n16184), .Z(n16651) );
  XNOR U17004 ( .A(n16650), .B(n16651), .Z(n16653) );
  XOR U17005 ( .A(b[37]), .B(n23852), .Z(n16457) );
  NANDN U17006 ( .A(n16457), .B(n36311), .Z(n16192) );
  NANDN U17007 ( .A(n16190), .B(n36309), .Z(n16191) );
  NAND U17008 ( .A(n16192), .B(n16191), .Z(n16536) );
  XNOR U17009 ( .A(a[81]), .B(b[5]), .Z(n16460) );
  OR U17010 ( .A(n16460), .B(n29363), .Z(n16195) );
  NANDN U17011 ( .A(n16193), .B(n29864), .Z(n16194) );
  NAND U17012 ( .A(n16195), .B(n16194), .Z(n16533) );
  XNOR U17013 ( .A(a[83]), .B(n967), .Z(n16463) );
  NAND U17014 ( .A(n16463), .B(n28939), .Z(n16198) );
  NAND U17015 ( .A(n28938), .B(n16196), .Z(n16197) );
  AND U17016 ( .A(n16198), .B(n16197), .Z(n16534) );
  XNOR U17017 ( .A(n16533), .B(n16534), .Z(n16535) );
  XNOR U17018 ( .A(n16536), .B(n16535), .Z(n16438) );
  XNOR U17019 ( .A(b[13]), .B(a[73]), .Z(n16466) );
  OR U17020 ( .A(n16466), .B(n31550), .Z(n16201) );
  NANDN U17021 ( .A(n16199), .B(n31874), .Z(n16200) );
  NAND U17022 ( .A(n16201), .B(n16200), .Z(n16623) );
  NAND U17023 ( .A(n34848), .B(n16202), .Z(n16204) );
  XNOR U17024 ( .A(n35375), .B(a[59]), .Z(n16469) );
  NAND U17025 ( .A(n34618), .B(n16469), .Z(n16203) );
  NAND U17026 ( .A(n16204), .B(n16203), .Z(n16620) );
  NAND U17027 ( .A(n35188), .B(n16205), .Z(n16207) );
  XOR U17028 ( .A(n35540), .B(n26122), .Z(n16472) );
  NANDN U17029 ( .A(n34968), .B(n16472), .Z(n16206) );
  AND U17030 ( .A(n16207), .B(n16206), .Z(n16621) );
  XNOR U17031 ( .A(n16620), .B(n16621), .Z(n16622) );
  XNOR U17032 ( .A(n16623), .B(n16622), .Z(n16435) );
  NANDN U17033 ( .A(n16209), .B(n16208), .Z(n16213) );
  NAND U17034 ( .A(n16211), .B(n16210), .Z(n16212) );
  NAND U17035 ( .A(n16213), .B(n16212), .Z(n16436) );
  XNOR U17036 ( .A(n16435), .B(n16436), .Z(n16437) );
  XOR U17037 ( .A(n16438), .B(n16437), .Z(n16429) );
  NANDN U17038 ( .A(n16215), .B(n16214), .Z(n16219) );
  NAND U17039 ( .A(n16217), .B(n16216), .Z(n16218) );
  NAND U17040 ( .A(n16219), .B(n16218), .Z(n16571) );
  ANDN U17041 ( .B(b[63]), .A(n16220), .Z(n16587) );
  NANDN U17042 ( .A(n16221), .B(n38369), .Z(n16223) );
  XOR U17043 ( .A(b[61]), .B(n16916), .Z(n16487) );
  OR U17044 ( .A(n16487), .B(n38371), .Z(n16222) );
  NAND U17045 ( .A(n16223), .B(n16222), .Z(n16585) );
  NANDN U17046 ( .A(n16224), .B(n35311), .Z(n16226) );
  XOR U17047 ( .A(b[31]), .B(n25466), .Z(n16490) );
  NANDN U17048 ( .A(n16490), .B(n35313), .Z(n16225) );
  AND U17049 ( .A(n16226), .B(n16225), .Z(n16584) );
  XNOR U17050 ( .A(n16585), .B(n16584), .Z(n16586) );
  XOR U17051 ( .A(n16587), .B(n16586), .Z(n16569) );
  NAND U17052 ( .A(n33283), .B(n16227), .Z(n16229) );
  XOR U17053 ( .A(n33020), .B(n29372), .Z(n16493) );
  NANDN U17054 ( .A(n33021), .B(n16493), .Z(n16228) );
  NAND U17055 ( .A(n16229), .B(n16228), .Z(n16524) );
  XNOR U17056 ( .A(b[21]), .B(a[65]), .Z(n16496) );
  OR U17057 ( .A(n16496), .B(n33634), .Z(n16232) );
  NAND U17058 ( .A(n16230), .B(n33464), .Z(n16231) );
  NAND U17059 ( .A(n16232), .B(n16231), .Z(n16521) );
  NAND U17060 ( .A(n34044), .B(n16233), .Z(n16235) );
  XNOR U17061 ( .A(n34510), .B(a[63]), .Z(n16499) );
  NANDN U17062 ( .A(n33867), .B(n16499), .Z(n16234) );
  AND U17063 ( .A(n16235), .B(n16234), .Z(n16522) );
  XNOR U17064 ( .A(n16521), .B(n16522), .Z(n16523) );
  XNOR U17065 ( .A(n16524), .B(n16523), .Z(n16570) );
  XOR U17066 ( .A(n16569), .B(n16570), .Z(n16572) );
  XOR U17067 ( .A(n16571), .B(n16572), .Z(n16430) );
  XOR U17068 ( .A(n16429), .B(n16430), .Z(n16431) );
  XOR U17069 ( .A(n16432), .B(n16431), .Z(n16646) );
  NANDN U17070 ( .A(n16237), .B(n16236), .Z(n16241) );
  NANDN U17071 ( .A(n16239), .B(n16238), .Z(n16240) );
  NAND U17072 ( .A(n16241), .B(n16240), .Z(n16645) );
  NANDN U17073 ( .A(n16243), .B(n16242), .Z(n16247) );
  NAND U17074 ( .A(n16245), .B(n16244), .Z(n16246) );
  NAND U17075 ( .A(n16247), .B(n16246), .Z(n16443) );
  NANDN U17076 ( .A(n16249), .B(n16248), .Z(n16253) );
  NAND U17077 ( .A(n16251), .B(n16250), .Z(n16252) );
  NAND U17078 ( .A(n16253), .B(n16252), .Z(n16641) );
  XNOR U17079 ( .A(b[41]), .B(a[45]), .Z(n16512) );
  OR U17080 ( .A(n16512), .B(n36905), .Z(n16256) );
  NANDN U17081 ( .A(n16254), .B(n36807), .Z(n16255) );
  NAND U17082 ( .A(n16256), .B(n16255), .Z(n16530) );
  XOR U17083 ( .A(b[57]), .B(n18003), .Z(n16515) );
  OR U17084 ( .A(n16515), .B(n965), .Z(n16259) );
  NANDN U17085 ( .A(n16257), .B(n38194), .Z(n16258) );
  NAND U17086 ( .A(n16259), .B(n16258), .Z(n16527) );
  NAND U17087 ( .A(n38326), .B(n16260), .Z(n16262) );
  XOR U17088 ( .A(n38400), .B(n17960), .Z(n16518) );
  NANDN U17089 ( .A(n38273), .B(n16518), .Z(n16261) );
  AND U17090 ( .A(n16262), .B(n16261), .Z(n16528) );
  XNOR U17091 ( .A(n16527), .B(n16528), .Z(n16529) );
  XNOR U17092 ( .A(n16530), .B(n16529), .Z(n16638) );
  XOR U17093 ( .A(b[33]), .B(n25001), .Z(n16502) );
  NANDN U17094 ( .A(n16502), .B(n35620), .Z(n16265) );
  NANDN U17095 ( .A(n16263), .B(n35621), .Z(n16264) );
  NAND U17096 ( .A(n16265), .B(n16264), .Z(n16635) );
  NANDN U17097 ( .A(n966), .B(a[85]), .Z(n16266) );
  XOR U17098 ( .A(n29232), .B(n16266), .Z(n16268) );
  IV U17099 ( .A(a[84]), .Z(n33185) );
  NANDN U17100 ( .A(n33185), .B(n966), .Z(n16267) );
  AND U17101 ( .A(n16268), .B(n16267), .Z(n16632) );
  XOR U17102 ( .A(b[63]), .B(n16269), .Z(n16509) );
  NANDN U17103 ( .A(n16509), .B(n38422), .Z(n16272) );
  NANDN U17104 ( .A(n16270), .B(n38423), .Z(n16271) );
  AND U17105 ( .A(n16272), .B(n16271), .Z(n16633) );
  XNOR U17106 ( .A(n16632), .B(n16633), .Z(n16634) );
  XOR U17107 ( .A(n16635), .B(n16634), .Z(n16639) );
  XNOR U17108 ( .A(n16638), .B(n16639), .Z(n16640) );
  XNOR U17109 ( .A(n16641), .B(n16640), .Z(n16441) );
  NANDN U17110 ( .A(n16274), .B(n16273), .Z(n16278) );
  NAND U17111 ( .A(n16276), .B(n16275), .Z(n16277) );
  AND U17112 ( .A(n16278), .B(n16277), .Z(n16442) );
  XNOR U17113 ( .A(n16441), .B(n16442), .Z(n16444) );
  XOR U17114 ( .A(n16443), .B(n16444), .Z(n16644) );
  XNOR U17115 ( .A(n16645), .B(n16644), .Z(n16647) );
  XNOR U17116 ( .A(n16646), .B(n16647), .Z(n16652) );
  XOR U17117 ( .A(n16653), .B(n16652), .Z(n16683) );
  OR U17118 ( .A(n16280), .B(n16279), .Z(n16284) );
  NAND U17119 ( .A(n16282), .B(n16281), .Z(n16283) );
  NAND U17120 ( .A(n16284), .B(n16283), .Z(n16658) );
  XOR U17121 ( .A(b[49]), .B(n20352), .Z(n16554) );
  OR U17122 ( .A(n16554), .B(n37756), .Z(n16287) );
  NANDN U17123 ( .A(n16285), .B(n37652), .Z(n16286) );
  NAND U17124 ( .A(n16287), .B(n16286), .Z(n16593) );
  NAND U17125 ( .A(n37469), .B(n16288), .Z(n16290) );
  XOR U17126 ( .A(n978), .B(n20867), .Z(n16557) );
  NAND U17127 ( .A(n16557), .B(n37471), .Z(n16289) );
  NAND U17128 ( .A(n16290), .B(n16289), .Z(n16590) );
  XNOR U17129 ( .A(a[77]), .B(b[9]), .Z(n16560) );
  NANDN U17130 ( .A(n16560), .B(n30509), .Z(n16293) );
  NANDN U17131 ( .A(n16291), .B(n30846), .Z(n16292) );
  AND U17132 ( .A(n16293), .B(n16292), .Z(n16591) );
  XNOR U17133 ( .A(n16590), .B(n16591), .Z(n16592) );
  XNOR U17134 ( .A(n16593), .B(n16592), .Z(n16451) );
  XNOR U17135 ( .A(b[11]), .B(a[75]), .Z(n16545) );
  OR U17136 ( .A(n16545), .B(n31369), .Z(n16296) );
  NANDN U17137 ( .A(n16294), .B(n31119), .Z(n16295) );
  NAND U17138 ( .A(n16296), .B(n16295), .Z(n16566) );
  XOR U17139 ( .A(b[43]), .B(n21996), .Z(n16548) );
  NANDN U17140 ( .A(n16548), .B(n37068), .Z(n16299) );
  NANDN U17141 ( .A(n16297), .B(n37069), .Z(n16298) );
  NAND U17142 ( .A(n16299), .B(n16298), .Z(n16563) );
  XNOR U17143 ( .A(b[45]), .B(a[41]), .Z(n16551) );
  NANDN U17144 ( .A(n16551), .B(n37261), .Z(n16302) );
  NANDN U17145 ( .A(n16300), .B(n37262), .Z(n16301) );
  AND U17146 ( .A(n16302), .B(n16301), .Z(n16564) );
  XNOR U17147 ( .A(n16563), .B(n16564), .Z(n16565) );
  XOR U17148 ( .A(n16566), .B(n16565), .Z(n16452) );
  XNOR U17149 ( .A(n16451), .B(n16452), .Z(n16453) );
  NANDN U17150 ( .A(n16304), .B(n16303), .Z(n16308) );
  NAND U17151 ( .A(n16306), .B(n16305), .Z(n16307) );
  AND U17152 ( .A(n16308), .B(n16307), .Z(n16454) );
  XNOR U17153 ( .A(n16453), .B(n16454), .Z(n16661) );
  XNOR U17154 ( .A(n16661), .B(n16660), .Z(n16662) );
  XNOR U17155 ( .A(b[35]), .B(a[51]), .Z(n16575) );
  NANDN U17156 ( .A(n16575), .B(n35985), .Z(n16315) );
  NANDN U17157 ( .A(n16313), .B(n35986), .Z(n16314) );
  NAND U17158 ( .A(n16315), .B(n16314), .Z(n16629) );
  XNOR U17159 ( .A(a[79]), .B(n31123), .Z(n16578) );
  NAND U17160 ( .A(n16578), .B(n29949), .Z(n16318) );
  NAND U17161 ( .A(n29948), .B(n16316), .Z(n16317) );
  NAND U17162 ( .A(n16318), .B(n16317), .Z(n16626) );
  XOR U17163 ( .A(b[55]), .B(n18639), .Z(n16581) );
  NANDN U17164 ( .A(n16581), .B(n38075), .Z(n16321) );
  NANDN U17165 ( .A(n16319), .B(n38073), .Z(n16320) );
  AND U17166 ( .A(n16321), .B(n16320), .Z(n16627) );
  XNOR U17167 ( .A(n16626), .B(n16627), .Z(n16628) );
  XNOR U17168 ( .A(n16629), .B(n16628), .Z(n16448) );
  NANDN U17169 ( .A(n16323), .B(n16322), .Z(n16327) );
  NAND U17170 ( .A(n16325), .B(n16324), .Z(n16326) );
  NAND U17171 ( .A(n16327), .B(n16326), .Z(n16445) );
  NANDN U17172 ( .A(n16329), .B(n16328), .Z(n16333) );
  NAND U17173 ( .A(n16331), .B(n16330), .Z(n16332) );
  NAND U17174 ( .A(n16333), .B(n16332), .Z(n16446) );
  XNOR U17175 ( .A(n16445), .B(n16446), .Z(n16447) );
  XOR U17176 ( .A(n16448), .B(n16447), .Z(n16663) );
  XOR U17177 ( .A(n16662), .B(n16663), .Z(n16657) );
  OR U17178 ( .A(n16335), .B(n16334), .Z(n16339) );
  OR U17179 ( .A(n16337), .B(n16336), .Z(n16338) );
  NAND U17180 ( .A(n16339), .B(n16338), .Z(n16666) );
  NANDN U17181 ( .A(n16341), .B(n16340), .Z(n16345) );
  NAND U17182 ( .A(n16343), .B(n16342), .Z(n16344) );
  NAND U17183 ( .A(n16345), .B(n16344), .Z(n16667) );
  XNOR U17184 ( .A(n16666), .B(n16667), .Z(n16668) );
  NANDN U17185 ( .A(n16347), .B(n16346), .Z(n16351) );
  NAND U17186 ( .A(n16349), .B(n16348), .Z(n16350) );
  NAND U17187 ( .A(n16351), .B(n16350), .Z(n16599) );
  XOR U17188 ( .A(b[15]), .B(n30543), .Z(n16602) );
  OR U17189 ( .A(n16602), .B(n32010), .Z(n16354) );
  NANDN U17190 ( .A(n16352), .B(n32011), .Z(n16353) );
  NAND U17191 ( .A(n16354), .B(n16353), .Z(n16484) );
  XNOR U17192 ( .A(b[25]), .B(n27773), .Z(n16605) );
  NANDN U17193 ( .A(n34219), .B(n16605), .Z(n16357) );
  NAND U17194 ( .A(n34217), .B(n16355), .Z(n16356) );
  NAND U17195 ( .A(n16357), .B(n16356), .Z(n16481) );
  XOR U17196 ( .A(b[17]), .B(a[69]), .Z(n16608) );
  NAND U17197 ( .A(n16608), .B(n32543), .Z(n16360) );
  NANDN U17198 ( .A(n16358), .B(n32541), .Z(n16359) );
  AND U17199 ( .A(n16360), .B(n16359), .Z(n16482) );
  XNOR U17200 ( .A(n16481), .B(n16482), .Z(n16483) );
  XNOR U17201 ( .A(n16484), .B(n16483), .Z(n16539) );
  XOR U17202 ( .A(b[39]), .B(n23149), .Z(n16611) );
  NANDN U17203 ( .A(n16611), .B(n36553), .Z(n16363) );
  NANDN U17204 ( .A(n16361), .B(n36643), .Z(n16362) );
  NAND U17205 ( .A(n16363), .B(n16362), .Z(n16478) );
  XOR U17206 ( .A(b[51]), .B(n20315), .Z(n16614) );
  NANDN U17207 ( .A(n16614), .B(n37803), .Z(n16366) );
  NANDN U17208 ( .A(n16364), .B(n37802), .Z(n16365) );
  NAND U17209 ( .A(n16366), .B(n16365), .Z(n16475) );
  XOR U17210 ( .A(b[53]), .B(n19656), .Z(n16617) );
  NANDN U17211 ( .A(n16617), .B(n37940), .Z(n16369) );
  NANDN U17212 ( .A(n16367), .B(n37941), .Z(n16368) );
  AND U17213 ( .A(n16369), .B(n16368), .Z(n16476) );
  XNOR U17214 ( .A(n16475), .B(n16476), .Z(n16477) );
  XOR U17215 ( .A(n16478), .B(n16477), .Z(n16540) );
  XNOR U17216 ( .A(n16539), .B(n16540), .Z(n16541) );
  NANDN U17217 ( .A(n16371), .B(n16370), .Z(n16375) );
  NAND U17218 ( .A(n16373), .B(n16372), .Z(n16374) );
  AND U17219 ( .A(n16375), .B(n16374), .Z(n16542) );
  XNOR U17220 ( .A(n16541), .B(n16542), .Z(n16597) );
  NANDN U17221 ( .A(n16377), .B(n16376), .Z(n16381) );
  NAND U17222 ( .A(n16379), .B(n16378), .Z(n16380) );
  AND U17223 ( .A(n16381), .B(n16380), .Z(n16596) );
  XNOR U17224 ( .A(n16597), .B(n16596), .Z(n16598) );
  XOR U17225 ( .A(n16599), .B(n16598), .Z(n16669) );
  XNOR U17226 ( .A(n16668), .B(n16669), .Z(n16656) );
  XOR U17227 ( .A(n16657), .B(n16656), .Z(n16659) );
  XNOR U17228 ( .A(n16658), .B(n16659), .Z(n16682) );
  XNOR U17229 ( .A(n16683), .B(n16682), .Z(n16685) );
  NAND U17230 ( .A(n16383), .B(n16382), .Z(n16387) );
  OR U17231 ( .A(n16385), .B(n16384), .Z(n16386) );
  AND U17232 ( .A(n16387), .B(n16386), .Z(n16684) );
  XNOR U17233 ( .A(n16685), .B(n16684), .Z(n16691) );
  XOR U17234 ( .A(n16690), .B(n16691), .Z(n16695) );
  NANDN U17235 ( .A(n16389), .B(n16388), .Z(n16393) );
  NANDN U17236 ( .A(n16391), .B(n16390), .Z(n16392) );
  NAND U17237 ( .A(n16393), .B(n16392), .Z(n16693) );
  NANDN U17238 ( .A(n16395), .B(n16394), .Z(n16399) );
  NANDN U17239 ( .A(n16397), .B(n16396), .Z(n16398) );
  AND U17240 ( .A(n16399), .B(n16398), .Z(n16692) );
  XNOR U17241 ( .A(n16693), .B(n16692), .Z(n16694) );
  XOR U17242 ( .A(n16695), .B(n16694), .Z(n16698) );
  NANDN U17243 ( .A(n16401), .B(n16400), .Z(n16405) );
  NAND U17244 ( .A(n16403), .B(n16402), .Z(n16404) );
  NAND U17245 ( .A(n16405), .B(n16404), .Z(n16699) );
  XOR U17246 ( .A(n16698), .B(n16699), .Z(n16701) );
  NANDN U17247 ( .A(n16407), .B(n16406), .Z(n16411) );
  NANDN U17248 ( .A(n16409), .B(n16408), .Z(n16410) );
  NAND U17249 ( .A(n16411), .B(n16410), .Z(n16700) );
  XNOR U17250 ( .A(n16701), .B(n16700), .Z(n16423) );
  NANDN U17251 ( .A(n16413), .B(n16412), .Z(n16417) );
  NANDN U17252 ( .A(n16415), .B(n16414), .Z(n16416) );
  NAND U17253 ( .A(n16417), .B(n16416), .Z(n16424) );
  XNOR U17254 ( .A(n16423), .B(n16424), .Z(n16425) );
  XNOR U17255 ( .A(n16426), .B(n16425), .Z(n16704) );
  XNOR U17256 ( .A(n16704), .B(sreg[149]), .Z(n16706) );
  NAND U17257 ( .A(n16418), .B(sreg[148]), .Z(n16422) );
  OR U17258 ( .A(n16420), .B(n16419), .Z(n16421) );
  AND U17259 ( .A(n16422), .B(n16421), .Z(n16705) );
  XOR U17260 ( .A(n16706), .B(n16705), .Z(c[149]) );
  NANDN U17261 ( .A(n16424), .B(n16423), .Z(n16428) );
  NAND U17262 ( .A(n16426), .B(n16425), .Z(n16427) );
  NAND U17263 ( .A(n16428), .B(n16427), .Z(n16712) );
  OR U17264 ( .A(n16430), .B(n16429), .Z(n16434) );
  NANDN U17265 ( .A(n16432), .B(n16431), .Z(n16433) );
  NAND U17266 ( .A(n16434), .B(n16433), .Z(n16715) );
  NANDN U17267 ( .A(n16436), .B(n16435), .Z(n16440) );
  NAND U17268 ( .A(n16438), .B(n16437), .Z(n16439) );
  NAND U17269 ( .A(n16440), .B(n16439), .Z(n16958) );
  NANDN U17270 ( .A(n16446), .B(n16445), .Z(n16450) );
  NAND U17271 ( .A(n16448), .B(n16447), .Z(n16449) );
  AND U17272 ( .A(n16450), .B(n16449), .Z(n16957) );
  XOR U17273 ( .A(n16958), .B(n16959), .Z(n16716) );
  XOR U17274 ( .A(n16715), .B(n16716), .Z(n16717) );
  NANDN U17275 ( .A(n16452), .B(n16451), .Z(n16456) );
  NAND U17276 ( .A(n16454), .B(n16453), .Z(n16455) );
  NAND U17277 ( .A(n16456), .B(n16455), .Z(n16843) );
  XOR U17278 ( .A(b[37]), .B(n24671), .Z(n16871) );
  NANDN U17279 ( .A(n16871), .B(n36311), .Z(n16459) );
  NANDN U17280 ( .A(n16457), .B(n36309), .Z(n16458) );
  NAND U17281 ( .A(n16459), .B(n16458), .Z(n16929) );
  XOR U17282 ( .A(a[82]), .B(n968), .Z(n16874) );
  OR U17283 ( .A(n16874), .B(n29363), .Z(n16462) );
  NANDN U17284 ( .A(n16460), .B(n29864), .Z(n16461) );
  NAND U17285 ( .A(n16462), .B(n16461), .Z(n16926) );
  XOR U17286 ( .A(n33185), .B(n967), .Z(n16877) );
  NAND U17287 ( .A(n16877), .B(n28939), .Z(n16465) );
  NAND U17288 ( .A(n28938), .B(n16463), .Z(n16464) );
  AND U17289 ( .A(n16465), .B(n16464), .Z(n16927) );
  XNOR U17290 ( .A(n16926), .B(n16927), .Z(n16928) );
  XNOR U17291 ( .A(n16929), .B(n16928), .Z(n16822) );
  XOR U17292 ( .A(b[13]), .B(n31372), .Z(n16880) );
  OR U17293 ( .A(n16880), .B(n31550), .Z(n16468) );
  NANDN U17294 ( .A(n16466), .B(n31874), .Z(n16467) );
  NAND U17295 ( .A(n16468), .B(n16467), .Z(n16754) );
  NAND U17296 ( .A(n34848), .B(n16469), .Z(n16471) );
  XOR U17297 ( .A(n35375), .B(n27436), .Z(n16883) );
  NAND U17298 ( .A(n34618), .B(n16883), .Z(n16470) );
  NAND U17299 ( .A(n16471), .B(n16470), .Z(n16751) );
  NAND U17300 ( .A(n35188), .B(n16472), .Z(n16474) );
  XOR U17301 ( .A(n35540), .B(n26347), .Z(n16886) );
  NANDN U17302 ( .A(n34968), .B(n16886), .Z(n16473) );
  AND U17303 ( .A(n16474), .B(n16473), .Z(n16752) );
  XNOR U17304 ( .A(n16751), .B(n16752), .Z(n16753) );
  XOR U17305 ( .A(n16754), .B(n16753), .Z(n16823) );
  XOR U17306 ( .A(n16822), .B(n16823), .Z(n16825) );
  NANDN U17307 ( .A(n16476), .B(n16475), .Z(n16480) );
  NAND U17308 ( .A(n16478), .B(n16477), .Z(n16479) );
  NAND U17309 ( .A(n16480), .B(n16479), .Z(n16824) );
  XNOR U17310 ( .A(n16825), .B(n16824), .Z(n16841) );
  NANDN U17311 ( .A(n16482), .B(n16481), .Z(n16486) );
  NAND U17312 ( .A(n16484), .B(n16483), .Z(n16485) );
  NAND U17313 ( .A(n16486), .B(n16485), .Z(n16799) );
  NAND U17314 ( .A(a[22]), .B(b[63]), .Z(n16813) );
  NANDN U17315 ( .A(n16487), .B(n38369), .Z(n16489) );
  XOR U17316 ( .A(b[61]), .B(n17133), .Z(n16865) );
  OR U17317 ( .A(n16865), .B(n38371), .Z(n16488) );
  NAND U17318 ( .A(n16489), .B(n16488), .Z(n16811) );
  NANDN U17319 ( .A(n16490), .B(n35311), .Z(n16492) );
  XOR U17320 ( .A(b[31]), .B(n25860), .Z(n16868) );
  NANDN U17321 ( .A(n16868), .B(n35313), .Z(n16491) );
  AND U17322 ( .A(n16492), .B(n16491), .Z(n16810) );
  XNOR U17323 ( .A(n16811), .B(n16810), .Z(n16812) );
  XOR U17324 ( .A(n16813), .B(n16812), .Z(n16797) );
  NAND U17325 ( .A(n33283), .B(n16493), .Z(n16495) );
  XOR U17326 ( .A(n33020), .B(n29868), .Z(n16850) );
  NANDN U17327 ( .A(n33021), .B(n16850), .Z(n16494) );
  NAND U17328 ( .A(n16495), .B(n16494), .Z(n16898) );
  XNOR U17329 ( .A(b[21]), .B(a[66]), .Z(n16853) );
  OR U17330 ( .A(n16853), .B(n33634), .Z(n16498) );
  NANDN U17331 ( .A(n16496), .B(n33464), .Z(n16497) );
  NAND U17332 ( .A(n16498), .B(n16497), .Z(n16895) );
  NAND U17333 ( .A(n34044), .B(n16499), .Z(n16501) );
  XNOR U17334 ( .A(n34510), .B(a[64]), .Z(n16856) );
  NANDN U17335 ( .A(n33867), .B(n16856), .Z(n16500) );
  AND U17336 ( .A(n16501), .B(n16500), .Z(n16896) );
  XNOR U17337 ( .A(n16895), .B(n16896), .Z(n16897) );
  XNOR U17338 ( .A(n16898), .B(n16897), .Z(n16798) );
  XNOR U17339 ( .A(n16797), .B(n16798), .Z(n16800) );
  XNOR U17340 ( .A(n16799), .B(n16800), .Z(n16840) );
  XNOR U17341 ( .A(n16841), .B(n16840), .Z(n16842) );
  XNOR U17342 ( .A(n16843), .B(n16842), .Z(n16724) );
  XOR U17343 ( .A(b[33]), .B(n25177), .Z(n16910) );
  NANDN U17344 ( .A(n16910), .B(n35620), .Z(n16504) );
  NANDN U17345 ( .A(n16502), .B(n35621), .Z(n16503) );
  NAND U17346 ( .A(n16504), .B(n16503), .Z(n16766) );
  NANDN U17347 ( .A(n966), .B(a[86]), .Z(n16505) );
  XOR U17348 ( .A(n29232), .B(n16505), .Z(n16507) );
  NANDN U17349 ( .A(b[0]), .B(a[85]), .Z(n16506) );
  AND U17350 ( .A(n16507), .B(n16506), .Z(n16763) );
  XOR U17351 ( .A(b[63]), .B(n16508), .Z(n16917) );
  NANDN U17352 ( .A(n16917), .B(n38422), .Z(n16511) );
  NANDN U17353 ( .A(n16509), .B(n38423), .Z(n16510) );
  AND U17354 ( .A(n16511), .B(n16510), .Z(n16764) );
  XNOR U17355 ( .A(n16763), .B(n16764), .Z(n16765) );
  XNOR U17356 ( .A(n16766), .B(n16765), .Z(n16729) );
  XNOR U17357 ( .A(b[41]), .B(a[46]), .Z(n16901) );
  OR U17358 ( .A(n16901), .B(n36905), .Z(n16514) );
  NANDN U17359 ( .A(n16512), .B(n36807), .Z(n16513) );
  NAND U17360 ( .A(n16514), .B(n16513), .Z(n16923) );
  XOR U17361 ( .A(b[57]), .B(n18804), .Z(n16904) );
  OR U17362 ( .A(n16904), .B(n965), .Z(n16517) );
  NANDN U17363 ( .A(n16515), .B(n38194), .Z(n16516) );
  NAND U17364 ( .A(n16517), .B(n16516), .Z(n16920) );
  NAND U17365 ( .A(n38326), .B(n16518), .Z(n16520) );
  XOR U17366 ( .A(n38400), .B(n17702), .Z(n16907) );
  NANDN U17367 ( .A(n38273), .B(n16907), .Z(n16519) );
  AND U17368 ( .A(n16520), .B(n16519), .Z(n16921) );
  XNOR U17369 ( .A(n16920), .B(n16921), .Z(n16922) );
  XOR U17370 ( .A(n16923), .B(n16922), .Z(n16728) );
  NANDN U17371 ( .A(n16522), .B(n16521), .Z(n16526) );
  NAND U17372 ( .A(n16524), .B(n16523), .Z(n16525) );
  NAND U17373 ( .A(n16526), .B(n16525), .Z(n16727) );
  XNOR U17374 ( .A(n16728), .B(n16727), .Z(n16730) );
  XNOR U17375 ( .A(n16729), .B(n16730), .Z(n16837) );
  NANDN U17376 ( .A(n16528), .B(n16527), .Z(n16532) );
  NAND U17377 ( .A(n16530), .B(n16529), .Z(n16531) );
  NAND U17378 ( .A(n16532), .B(n16531), .Z(n16834) );
  NANDN U17379 ( .A(n16534), .B(n16533), .Z(n16538) );
  NAND U17380 ( .A(n16536), .B(n16535), .Z(n16537) );
  AND U17381 ( .A(n16538), .B(n16537), .Z(n16835) );
  XNOR U17382 ( .A(n16834), .B(n16835), .Z(n16836) );
  XNOR U17383 ( .A(n16837), .B(n16836), .Z(n16722) );
  NANDN U17384 ( .A(n16540), .B(n16539), .Z(n16544) );
  NAND U17385 ( .A(n16542), .B(n16541), .Z(n16543) );
  AND U17386 ( .A(n16544), .B(n16543), .Z(n16721) );
  XOR U17387 ( .A(n16722), .B(n16721), .Z(n16723) );
  XNOR U17388 ( .A(n16724), .B(n16723), .Z(n16718) );
  XOR U17389 ( .A(n16717), .B(n16718), .Z(n16962) );
  XOR U17390 ( .A(a[76]), .B(n970), .Z(n16773) );
  OR U17391 ( .A(n16773), .B(n31369), .Z(n16547) );
  NANDN U17392 ( .A(n16545), .B(n31119), .Z(n16546) );
  NAND U17393 ( .A(n16547), .B(n16546), .Z(n16794) );
  XOR U17394 ( .A(b[43]), .B(n22289), .Z(n16776) );
  NANDN U17395 ( .A(n16776), .B(n37068), .Z(n16550) );
  NANDN U17396 ( .A(n16548), .B(n37069), .Z(n16549) );
  NAND U17397 ( .A(n16550), .B(n16549), .Z(n16791) );
  XNOR U17398 ( .A(b[45]), .B(a[42]), .Z(n16779) );
  NANDN U17399 ( .A(n16779), .B(n37261), .Z(n16553) );
  NANDN U17400 ( .A(n16551), .B(n37262), .Z(n16552) );
  AND U17401 ( .A(n16553), .B(n16552), .Z(n16792) );
  XNOR U17402 ( .A(n16791), .B(n16792), .Z(n16793) );
  XNOR U17403 ( .A(n16794), .B(n16793), .Z(n16849) );
  XOR U17404 ( .A(n979), .B(n20686), .Z(n16782) );
  NANDN U17405 ( .A(n37756), .B(n16782), .Z(n16556) );
  NANDN U17406 ( .A(n16554), .B(n37652), .Z(n16555) );
  NAND U17407 ( .A(n16556), .B(n16555), .Z(n16819) );
  NAND U17408 ( .A(n37469), .B(n16557), .Z(n16559) );
  XOR U17409 ( .A(b[47]), .B(n21149), .Z(n16785) );
  NANDN U17410 ( .A(n16785), .B(n37471), .Z(n16558) );
  NAND U17411 ( .A(n16559), .B(n16558), .Z(n16816) );
  XOR U17412 ( .A(n31870), .B(n969), .Z(n16788) );
  NAND U17413 ( .A(n30509), .B(n16788), .Z(n16562) );
  NANDN U17414 ( .A(n16560), .B(n30846), .Z(n16561) );
  AND U17415 ( .A(n16562), .B(n16561), .Z(n16817) );
  XNOR U17416 ( .A(n16816), .B(n16817), .Z(n16818) );
  XNOR U17417 ( .A(n16819), .B(n16818), .Z(n16846) );
  NANDN U17418 ( .A(n16564), .B(n16563), .Z(n16568) );
  NAND U17419 ( .A(n16566), .B(n16565), .Z(n16567) );
  NAND U17420 ( .A(n16568), .B(n16567), .Z(n16847) );
  XNOR U17421 ( .A(n16846), .B(n16847), .Z(n16848) );
  XOR U17422 ( .A(n16849), .B(n16848), .Z(n16944) );
  NANDN U17423 ( .A(n16570), .B(n16569), .Z(n16574) );
  NANDN U17424 ( .A(n16572), .B(n16571), .Z(n16573) );
  AND U17425 ( .A(n16574), .B(n16573), .Z(n16945) );
  XNOR U17426 ( .A(n16944), .B(n16945), .Z(n16947) );
  XNOR U17427 ( .A(b[35]), .B(a[52]), .Z(n16801) );
  NANDN U17428 ( .A(n16801), .B(n35985), .Z(n16577) );
  NANDN U17429 ( .A(n16575), .B(n35986), .Z(n16576) );
  NAND U17430 ( .A(n16577), .B(n16576), .Z(n16760) );
  XOR U17431 ( .A(n32814), .B(n31123), .Z(n16804) );
  NAND U17432 ( .A(n16804), .B(n29949), .Z(n16580) );
  NAND U17433 ( .A(n29948), .B(n16578), .Z(n16579) );
  NAND U17434 ( .A(n16580), .B(n16579), .Z(n16757) );
  XOR U17435 ( .A(b[55]), .B(n18841), .Z(n16807) );
  NANDN U17436 ( .A(n16807), .B(n38075), .Z(n16583) );
  NANDN U17437 ( .A(n16581), .B(n38073), .Z(n16582) );
  AND U17438 ( .A(n16583), .B(n16582), .Z(n16758) );
  XNOR U17439 ( .A(n16757), .B(n16758), .Z(n16759) );
  XNOR U17440 ( .A(n16760), .B(n16759), .Z(n16831) );
  NANDN U17441 ( .A(n16585), .B(n16584), .Z(n16589) );
  NANDN U17442 ( .A(n16587), .B(n16586), .Z(n16588) );
  NAND U17443 ( .A(n16589), .B(n16588), .Z(n16828) );
  NANDN U17444 ( .A(n16591), .B(n16590), .Z(n16595) );
  NAND U17445 ( .A(n16593), .B(n16592), .Z(n16594) );
  NAND U17446 ( .A(n16595), .B(n16594), .Z(n16829) );
  XNOR U17447 ( .A(n16828), .B(n16829), .Z(n16830) );
  XOR U17448 ( .A(n16831), .B(n16830), .Z(n16946) );
  XNOR U17449 ( .A(n16947), .B(n16946), .Z(n16938) );
  NANDN U17450 ( .A(n16597), .B(n16596), .Z(n16601) );
  NANDN U17451 ( .A(n16599), .B(n16598), .Z(n16600) );
  NAND U17452 ( .A(n16601), .B(n16600), .Z(n16953) );
  XOR U17453 ( .A(b[15]), .B(n30210), .Z(n16733) );
  OR U17454 ( .A(n16733), .B(n32010), .Z(n16604) );
  NANDN U17455 ( .A(n16602), .B(n32011), .Z(n16603) );
  NAND U17456 ( .A(n16604), .B(n16603), .Z(n16862) );
  XOR U17457 ( .A(b[25]), .B(a[62]), .Z(n16736) );
  NANDN U17458 ( .A(n34219), .B(n16736), .Z(n16607) );
  NAND U17459 ( .A(n34217), .B(n16605), .Z(n16606) );
  NAND U17460 ( .A(n16607), .B(n16606), .Z(n16859) );
  XNOR U17461 ( .A(b[17]), .B(a[70]), .Z(n16739) );
  NANDN U17462 ( .A(n16739), .B(n32543), .Z(n16610) );
  NAND U17463 ( .A(n16608), .B(n32541), .Z(n16609) );
  AND U17464 ( .A(n16610), .B(n16609), .Z(n16860) );
  XNOR U17465 ( .A(n16859), .B(n16860), .Z(n16861) );
  XNOR U17466 ( .A(n16862), .B(n16861), .Z(n16932) );
  XOR U17467 ( .A(b[39]), .B(n23447), .Z(n16742) );
  NANDN U17468 ( .A(n16742), .B(n36553), .Z(n16613) );
  NANDN U17469 ( .A(n16611), .B(n36643), .Z(n16612) );
  NAND U17470 ( .A(n16613), .B(n16612), .Z(n16892) );
  XOR U17471 ( .A(b[51]), .B(n19980), .Z(n16745) );
  NANDN U17472 ( .A(n16745), .B(n37803), .Z(n16616) );
  NANDN U17473 ( .A(n16614), .B(n37802), .Z(n16615) );
  NAND U17474 ( .A(n16616), .B(n16615), .Z(n16889) );
  XOR U17475 ( .A(b[53]), .B(n19513), .Z(n16748) );
  NANDN U17476 ( .A(n16748), .B(n37940), .Z(n16619) );
  NANDN U17477 ( .A(n16617), .B(n37941), .Z(n16618) );
  AND U17478 ( .A(n16619), .B(n16618), .Z(n16890) );
  XNOR U17479 ( .A(n16889), .B(n16890), .Z(n16891) );
  XOR U17480 ( .A(n16892), .B(n16891), .Z(n16933) );
  XOR U17481 ( .A(n16932), .B(n16933), .Z(n16935) );
  NANDN U17482 ( .A(n16621), .B(n16620), .Z(n16625) );
  NAND U17483 ( .A(n16623), .B(n16622), .Z(n16624) );
  NAND U17484 ( .A(n16625), .B(n16624), .Z(n16934) );
  XNOR U17485 ( .A(n16935), .B(n16934), .Z(n16770) );
  NANDN U17486 ( .A(n16627), .B(n16626), .Z(n16631) );
  NAND U17487 ( .A(n16629), .B(n16628), .Z(n16630) );
  NAND U17488 ( .A(n16631), .B(n16630), .Z(n16767) );
  NANDN U17489 ( .A(n16633), .B(n16632), .Z(n16637) );
  NAND U17490 ( .A(n16635), .B(n16634), .Z(n16636) );
  AND U17491 ( .A(n16637), .B(n16636), .Z(n16768) );
  XNOR U17492 ( .A(n16767), .B(n16768), .Z(n16769) );
  XNOR U17493 ( .A(n16770), .B(n16769), .Z(n16950) );
  NANDN U17494 ( .A(n16639), .B(n16638), .Z(n16643) );
  NANDN U17495 ( .A(n16641), .B(n16640), .Z(n16642) );
  AND U17496 ( .A(n16643), .B(n16642), .Z(n16951) );
  XNOR U17497 ( .A(n16950), .B(n16951), .Z(n16952) );
  XOR U17498 ( .A(n16953), .B(n16952), .Z(n16939) );
  NAND U17499 ( .A(n16645), .B(n16644), .Z(n16649) );
  NANDN U17500 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U17501 ( .A(n16649), .B(n16648), .Z(n16941) );
  XNOR U17502 ( .A(n16940), .B(n16941), .Z(n16963) );
  XNOR U17503 ( .A(n16962), .B(n16963), .Z(n16964) );
  NAND U17504 ( .A(n16651), .B(n16650), .Z(n16655) );
  NANDN U17505 ( .A(n16653), .B(n16652), .Z(n16654) );
  AND U17506 ( .A(n16655), .B(n16654), .Z(n16965) );
  XNOR U17507 ( .A(n16964), .B(n16965), .Z(n16977) );
  NANDN U17508 ( .A(n16661), .B(n16660), .Z(n16665) );
  NAND U17509 ( .A(n16663), .B(n16662), .Z(n16664) );
  NAND U17510 ( .A(n16665), .B(n16664), .Z(n16969) );
  NANDN U17511 ( .A(n16667), .B(n16666), .Z(n16671) );
  NANDN U17512 ( .A(n16669), .B(n16668), .Z(n16670) );
  AND U17513 ( .A(n16671), .B(n16670), .Z(n16968) );
  XNOR U17514 ( .A(n16969), .B(n16968), .Z(n16970) );
  XNOR U17515 ( .A(n16970), .B(n16971), .Z(n16974) );
  XNOR U17516 ( .A(n16975), .B(n16974), .Z(n16976) );
  XNOR U17517 ( .A(n16977), .B(n16976), .Z(n16981) );
  NANDN U17518 ( .A(n16677), .B(n16676), .Z(n16681) );
  NAND U17519 ( .A(n16679), .B(n16678), .Z(n16680) );
  NAND U17520 ( .A(n16681), .B(n16680), .Z(n16978) );
  NAND U17521 ( .A(n16683), .B(n16682), .Z(n16687) );
  NANDN U17522 ( .A(n16685), .B(n16684), .Z(n16686) );
  NAND U17523 ( .A(n16687), .B(n16686), .Z(n16979) );
  XNOR U17524 ( .A(n16978), .B(n16979), .Z(n16980) );
  XNOR U17525 ( .A(n16981), .B(n16980), .Z(n16985) );
  XOR U17526 ( .A(n16985), .B(n16984), .Z(n16986) );
  NANDN U17527 ( .A(n16693), .B(n16692), .Z(n16697) );
  NANDN U17528 ( .A(n16695), .B(n16694), .Z(n16696) );
  NAND U17529 ( .A(n16697), .B(n16696), .Z(n16987) );
  XOR U17530 ( .A(n16986), .B(n16987), .Z(n16709) );
  NANDN U17531 ( .A(n16699), .B(n16698), .Z(n16703) );
  OR U17532 ( .A(n16701), .B(n16700), .Z(n16702) );
  NAND U17533 ( .A(n16703), .B(n16702), .Z(n16710) );
  XNOR U17534 ( .A(n16709), .B(n16710), .Z(n16711) );
  XNOR U17535 ( .A(n16712), .B(n16711), .Z(n16990) );
  XNOR U17536 ( .A(n16990), .B(sreg[150]), .Z(n16992) );
  NAND U17537 ( .A(n16704), .B(sreg[149]), .Z(n16708) );
  OR U17538 ( .A(n16706), .B(n16705), .Z(n16707) );
  AND U17539 ( .A(n16708), .B(n16707), .Z(n16991) );
  XOR U17540 ( .A(n16992), .B(n16991), .Z(c[150]) );
  NANDN U17541 ( .A(n16710), .B(n16709), .Z(n16714) );
  NAND U17542 ( .A(n16712), .B(n16711), .Z(n16713) );
  NAND U17543 ( .A(n16714), .B(n16713), .Z(n16998) );
  OR U17544 ( .A(n16716), .B(n16715), .Z(n16720) );
  NANDN U17545 ( .A(n16718), .B(n16717), .Z(n16719) );
  NAND U17546 ( .A(n16720), .B(n16719), .Z(n17022) );
  OR U17547 ( .A(n16722), .B(n16721), .Z(n16726) );
  NAND U17548 ( .A(n16724), .B(n16723), .Z(n16725) );
  NAND U17549 ( .A(n16726), .B(n16725), .Z(n17278) );
  OR U17550 ( .A(n16728), .B(n16727), .Z(n16732) );
  NANDN U17551 ( .A(n16730), .B(n16729), .Z(n16731) );
  NAND U17552 ( .A(n16732), .B(n16731), .Z(n17266) );
  XNOR U17553 ( .A(b[15]), .B(a[73]), .Z(n17155) );
  OR U17554 ( .A(n17155), .B(n32010), .Z(n16735) );
  NANDN U17555 ( .A(n16733), .B(n32011), .Z(n16734) );
  NAND U17556 ( .A(n16735), .B(n16734), .Z(n17088) );
  XOR U17557 ( .A(b[25]), .B(a[63]), .Z(n17158) );
  NANDN U17558 ( .A(n34219), .B(n17158), .Z(n16738) );
  NAND U17559 ( .A(n34217), .B(n16736), .Z(n16737) );
  NAND U17560 ( .A(n16738), .B(n16737), .Z(n17085) );
  XNOR U17561 ( .A(b[17]), .B(a[71]), .Z(n17161) );
  NANDN U17562 ( .A(n17161), .B(n32543), .Z(n16741) );
  NANDN U17563 ( .A(n16739), .B(n32541), .Z(n16740) );
  AND U17564 ( .A(n16741), .B(n16740), .Z(n17086) );
  XNOR U17565 ( .A(n17085), .B(n17086), .Z(n17087) );
  XNOR U17566 ( .A(n17088), .B(n17087), .Z(n17106) );
  XOR U17567 ( .A(b[39]), .B(n23852), .Z(n17164) );
  NANDN U17568 ( .A(n17164), .B(n36553), .Z(n16744) );
  NANDN U17569 ( .A(n16742), .B(n36643), .Z(n16743) );
  NAND U17570 ( .A(n16744), .B(n16743), .Z(n17082) );
  XOR U17571 ( .A(b[51]), .B(n20352), .Z(n17167) );
  NANDN U17572 ( .A(n17167), .B(n37803), .Z(n16747) );
  NANDN U17573 ( .A(n16745), .B(n37802), .Z(n16746) );
  NAND U17574 ( .A(n16747), .B(n16746), .Z(n17079) );
  XOR U17575 ( .A(b[53]), .B(n20315), .Z(n17170) );
  NANDN U17576 ( .A(n17170), .B(n37940), .Z(n16750) );
  NANDN U17577 ( .A(n16748), .B(n37941), .Z(n16749) );
  AND U17578 ( .A(n16750), .B(n16749), .Z(n17080) );
  XNOR U17579 ( .A(n17079), .B(n17080), .Z(n17081) );
  XOR U17580 ( .A(n17082), .B(n17081), .Z(n17107) );
  XNOR U17581 ( .A(n17106), .B(n17107), .Z(n17108) );
  NANDN U17582 ( .A(n16752), .B(n16751), .Z(n16756) );
  NAND U17583 ( .A(n16754), .B(n16753), .Z(n16755) );
  NAND U17584 ( .A(n16756), .B(n16755), .Z(n17109) );
  XOR U17585 ( .A(n17108), .B(n17109), .Z(n17200) );
  NANDN U17586 ( .A(n16758), .B(n16757), .Z(n16762) );
  NAND U17587 ( .A(n16760), .B(n16759), .Z(n16761) );
  NAND U17588 ( .A(n16762), .B(n16761), .Z(n17197) );
  XNOR U17589 ( .A(n17197), .B(n17198), .Z(n17199) );
  XOR U17590 ( .A(n17200), .B(n17199), .Z(n17267) );
  XNOR U17591 ( .A(n17266), .B(n17267), .Z(n17268) );
  NANDN U17592 ( .A(n16768), .B(n16767), .Z(n16772) );
  NAND U17593 ( .A(n16770), .B(n16769), .Z(n16771) );
  AND U17594 ( .A(n16772), .B(n16771), .Z(n17269) );
  XNOR U17595 ( .A(n17268), .B(n17269), .Z(n17277) );
  XNOR U17596 ( .A(a[77]), .B(b[11]), .Z(n17209) );
  OR U17597 ( .A(n17209), .B(n31369), .Z(n16775) );
  NANDN U17598 ( .A(n16773), .B(n31119), .Z(n16774) );
  NAND U17599 ( .A(n16775), .B(n16774), .Z(n17230) );
  XOR U17600 ( .A(b[43]), .B(n22579), .Z(n17212) );
  NANDN U17601 ( .A(n17212), .B(n37068), .Z(n16778) );
  NANDN U17602 ( .A(n16776), .B(n37069), .Z(n16777) );
  NAND U17603 ( .A(n16778), .B(n16777), .Z(n17227) );
  XNOR U17604 ( .A(b[45]), .B(a[43]), .Z(n17215) );
  NANDN U17605 ( .A(n17215), .B(n37261), .Z(n16781) );
  NANDN U17606 ( .A(n16779), .B(n37262), .Z(n16780) );
  AND U17607 ( .A(n16781), .B(n16780), .Z(n17228) );
  XNOR U17608 ( .A(n17227), .B(n17228), .Z(n17229) );
  XNOR U17609 ( .A(n17230), .B(n17229), .Z(n17055) );
  NAND U17610 ( .A(n37652), .B(n16782), .Z(n16784) );
  XOR U17611 ( .A(n979), .B(a[39]), .Z(n17218) );
  OR U17612 ( .A(n17218), .B(n37756), .Z(n16783) );
  NAND U17613 ( .A(n16784), .B(n16783), .Z(n17250) );
  NANDN U17614 ( .A(n16785), .B(n37469), .Z(n16787) );
  XOR U17615 ( .A(b[47]), .B(n21441), .Z(n17221) );
  NANDN U17616 ( .A(n17221), .B(n37471), .Z(n16786) );
  AND U17617 ( .A(n16787), .B(n16786), .Z(n17249) );
  NAND U17618 ( .A(n30846), .B(n16788), .Z(n16790) );
  XNOR U17619 ( .A(a[79]), .B(n969), .Z(n17224) );
  NAND U17620 ( .A(n30509), .B(n17224), .Z(n16789) );
  NAND U17621 ( .A(n16790), .B(n16789), .Z(n17248) );
  XNOR U17622 ( .A(n17249), .B(n17248), .Z(n17251) );
  XOR U17623 ( .A(n17250), .B(n17251), .Z(n17056) );
  XNOR U17624 ( .A(n17055), .B(n17056), .Z(n17057) );
  NANDN U17625 ( .A(n16792), .B(n16791), .Z(n16796) );
  NAND U17626 ( .A(n16794), .B(n16793), .Z(n16795) );
  AND U17627 ( .A(n16796), .B(n16795), .Z(n17058) );
  XNOR U17628 ( .A(n17057), .B(n17058), .Z(n17261) );
  XNOR U17629 ( .A(n17261), .B(n17260), .Z(n17262) );
  XNOR U17630 ( .A(b[35]), .B(a[53]), .Z(n17233) );
  NANDN U17631 ( .A(n17233), .B(n35985), .Z(n16803) );
  NANDN U17632 ( .A(n16801), .B(n35986), .Z(n16802) );
  NAND U17633 ( .A(n16803), .B(n16802), .Z(n17182) );
  XNOR U17634 ( .A(a[81]), .B(n31123), .Z(n17236) );
  NAND U17635 ( .A(n17236), .B(n29949), .Z(n16806) );
  NAND U17636 ( .A(n29948), .B(n16804), .Z(n16805) );
  NAND U17637 ( .A(n16806), .B(n16805), .Z(n17179) );
  XOR U17638 ( .A(b[55]), .B(n19656), .Z(n17239) );
  NANDN U17639 ( .A(n17239), .B(n38075), .Z(n16809) );
  NANDN U17640 ( .A(n16807), .B(n38073), .Z(n16808) );
  AND U17641 ( .A(n16809), .B(n16808), .Z(n17180) );
  XNOR U17642 ( .A(n17179), .B(n17180), .Z(n17181) );
  XNOR U17643 ( .A(n17182), .B(n17181), .Z(n17034) );
  NANDN U17644 ( .A(n16811), .B(n16810), .Z(n16815) );
  NAND U17645 ( .A(n16813), .B(n16812), .Z(n16814) );
  NAND U17646 ( .A(n16815), .B(n16814), .Z(n17031) );
  NANDN U17647 ( .A(n16817), .B(n16816), .Z(n16821) );
  NAND U17648 ( .A(n16819), .B(n16818), .Z(n16820) );
  NAND U17649 ( .A(n16821), .B(n16820), .Z(n17032) );
  XNOR U17650 ( .A(n17031), .B(n17032), .Z(n17033) );
  XOR U17651 ( .A(n17034), .B(n17033), .Z(n17263) );
  XOR U17652 ( .A(n17262), .B(n17263), .Z(n17276) );
  XOR U17653 ( .A(n17277), .B(n17276), .Z(n17279) );
  XOR U17654 ( .A(n17278), .B(n17279), .Z(n17019) );
  NANDN U17655 ( .A(n16823), .B(n16822), .Z(n16827) );
  OR U17656 ( .A(n16825), .B(n16824), .Z(n16826) );
  AND U17657 ( .A(n16827), .B(n16826), .Z(n17275) );
  NANDN U17658 ( .A(n16829), .B(n16828), .Z(n16833) );
  NAND U17659 ( .A(n16831), .B(n16830), .Z(n16832) );
  NAND U17660 ( .A(n16833), .B(n16832), .Z(n17272) );
  NANDN U17661 ( .A(n16835), .B(n16834), .Z(n16839) );
  NANDN U17662 ( .A(n16837), .B(n16836), .Z(n16838) );
  NAND U17663 ( .A(n16839), .B(n16838), .Z(n17273) );
  XNOR U17664 ( .A(n17272), .B(n17273), .Z(n17274) );
  XNOR U17665 ( .A(n17275), .B(n17274), .Z(n17254) );
  NAND U17666 ( .A(n16841), .B(n16840), .Z(n16845) );
  OR U17667 ( .A(n16843), .B(n16842), .Z(n16844) );
  AND U17668 ( .A(n16845), .B(n16844), .Z(n17255) );
  XNOR U17669 ( .A(n17254), .B(n17255), .Z(n17257) );
  NAND U17670 ( .A(n33283), .B(n16850), .Z(n16852) );
  XNOR U17671 ( .A(n33020), .B(a[69]), .Z(n17097) );
  NANDN U17672 ( .A(n33021), .B(n17097), .Z(n16851) );
  NAND U17673 ( .A(n16852), .B(n16851), .Z(n17140) );
  XNOR U17674 ( .A(b[21]), .B(a[67]), .Z(n17100) );
  OR U17675 ( .A(n17100), .B(n33634), .Z(n16855) );
  NANDN U17676 ( .A(n16853), .B(n33464), .Z(n16854) );
  NAND U17677 ( .A(n16855), .B(n16854), .Z(n17137) );
  NAND U17678 ( .A(n34044), .B(n16856), .Z(n16858) );
  XOR U17679 ( .A(n34510), .B(n28403), .Z(n17103) );
  NANDN U17680 ( .A(n33867), .B(n17103), .Z(n16857) );
  AND U17681 ( .A(n16858), .B(n16857), .Z(n17138) );
  XNOR U17682 ( .A(n17137), .B(n17138), .Z(n17139) );
  XOR U17683 ( .A(n17140), .B(n17139), .Z(n17203) );
  NANDN U17684 ( .A(n16860), .B(n16859), .Z(n16864) );
  NAND U17685 ( .A(n16862), .B(n16861), .Z(n16863) );
  NAND U17686 ( .A(n16864), .B(n16863), .Z(n17204) );
  XNOR U17687 ( .A(n17203), .B(n17204), .Z(n17206) );
  NAND U17688 ( .A(a[23]), .B(b[63]), .Z(n17245) );
  NANDN U17689 ( .A(n16865), .B(n38369), .Z(n16867) );
  XOR U17690 ( .A(b[61]), .B(n17960), .Z(n17091) );
  OR U17691 ( .A(n17091), .B(n38371), .Z(n16866) );
  NAND U17692 ( .A(n16867), .B(n16866), .Z(n17243) );
  NANDN U17693 ( .A(n16868), .B(n35311), .Z(n16870) );
  XOR U17694 ( .A(b[31]), .B(n26122), .Z(n17094) );
  NANDN U17695 ( .A(n17094), .B(n35313), .Z(n16869) );
  AND U17696 ( .A(n16870), .B(n16869), .Z(n17242) );
  XNOR U17697 ( .A(n17243), .B(n17242), .Z(n17244) );
  XNOR U17698 ( .A(n17245), .B(n17244), .Z(n17205) );
  XNOR U17699 ( .A(n17206), .B(n17205), .Z(n17049) );
  XOR U17700 ( .A(b[37]), .B(n24288), .Z(n17061) );
  NANDN U17701 ( .A(n17061), .B(n36311), .Z(n16873) );
  NANDN U17702 ( .A(n16871), .B(n36309), .Z(n16872) );
  NAND U17703 ( .A(n16873), .B(n16872), .Z(n17115) );
  XNOR U17704 ( .A(a[83]), .B(b[5]), .Z(n17064) );
  OR U17705 ( .A(n17064), .B(n29363), .Z(n16876) );
  NANDN U17706 ( .A(n16874), .B(n29864), .Z(n16875) );
  NAND U17707 ( .A(n16876), .B(n16875), .Z(n17112) );
  XNOR U17708 ( .A(a[85]), .B(n967), .Z(n17067) );
  NAND U17709 ( .A(n17067), .B(n28939), .Z(n16879) );
  NAND U17710 ( .A(n28938), .B(n16877), .Z(n16878) );
  AND U17711 ( .A(n16879), .B(n16878), .Z(n17113) );
  XNOR U17712 ( .A(n17112), .B(n17113), .Z(n17114) );
  XNOR U17713 ( .A(n17115), .B(n17114), .Z(n17037) );
  XNOR U17714 ( .A(b[13]), .B(a[75]), .Z(n17070) );
  OR U17715 ( .A(n17070), .B(n31550), .Z(n16882) );
  NANDN U17716 ( .A(n16880), .B(n31874), .Z(n16881) );
  NAND U17717 ( .A(n16882), .B(n16881), .Z(n17176) );
  NAND U17718 ( .A(n34848), .B(n16883), .Z(n16885) );
  XOR U17719 ( .A(n35375), .B(n27773), .Z(n17073) );
  NAND U17720 ( .A(n34618), .B(n17073), .Z(n16884) );
  NAND U17721 ( .A(n16885), .B(n16884), .Z(n17173) );
  NAND U17722 ( .A(n35188), .B(n16886), .Z(n16888) );
  XNOR U17723 ( .A(n35540), .B(a[59]), .Z(n17076) );
  NANDN U17724 ( .A(n34968), .B(n17076), .Z(n16887) );
  AND U17725 ( .A(n16888), .B(n16887), .Z(n17174) );
  XNOR U17726 ( .A(n17173), .B(n17174), .Z(n17175) );
  XOR U17727 ( .A(n17176), .B(n17175), .Z(n17038) );
  XOR U17728 ( .A(n17037), .B(n17038), .Z(n17040) );
  NANDN U17729 ( .A(n16890), .B(n16889), .Z(n16894) );
  NAND U17730 ( .A(n16892), .B(n16891), .Z(n16893) );
  NAND U17731 ( .A(n16894), .B(n16893), .Z(n17039) );
  XOR U17732 ( .A(n17040), .B(n17039), .Z(n17050) );
  XOR U17733 ( .A(n17049), .B(n17050), .Z(n17052) );
  XNOR U17734 ( .A(n17051), .B(n17052), .Z(n17152) );
  NANDN U17735 ( .A(n16896), .B(n16895), .Z(n16900) );
  NAND U17736 ( .A(n16898), .B(n16897), .Z(n16899) );
  NAND U17737 ( .A(n16900), .B(n16899), .Z(n17194) );
  XNOR U17738 ( .A(b[41]), .B(a[47]), .Z(n17118) );
  OR U17739 ( .A(n17118), .B(n36905), .Z(n16903) );
  NANDN U17740 ( .A(n16901), .B(n36807), .Z(n16902) );
  NAND U17741 ( .A(n16903), .B(n16902), .Z(n17146) );
  XOR U17742 ( .A(b[57]), .B(n18639), .Z(n17121) );
  OR U17743 ( .A(n17121), .B(n965), .Z(n16906) );
  NANDN U17744 ( .A(n16904), .B(n38194), .Z(n16905) );
  NAND U17745 ( .A(n16906), .B(n16905), .Z(n17143) );
  NAND U17746 ( .A(n38326), .B(n16907), .Z(n16909) );
  XOR U17747 ( .A(n38400), .B(n18003), .Z(n17124) );
  NANDN U17748 ( .A(n38273), .B(n17124), .Z(n16908) );
  AND U17749 ( .A(n16909), .B(n16908), .Z(n17144) );
  XNOR U17750 ( .A(n17143), .B(n17144), .Z(n17145) );
  XOR U17751 ( .A(n17146), .B(n17145), .Z(n17191) );
  XOR U17752 ( .A(b[33]), .B(n25466), .Z(n17127) );
  NANDN U17753 ( .A(n17127), .B(n35620), .Z(n16912) );
  NANDN U17754 ( .A(n16910), .B(n35621), .Z(n16911) );
  NAND U17755 ( .A(n16912), .B(n16911), .Z(n17188) );
  NANDN U17756 ( .A(n966), .B(a[87]), .Z(n16913) );
  XOR U17757 ( .A(n29232), .B(n16913), .Z(n16915) );
  IV U17758 ( .A(a[86]), .Z(n33628) );
  NANDN U17759 ( .A(n33628), .B(n966), .Z(n16914) );
  AND U17760 ( .A(n16915), .B(n16914), .Z(n17185) );
  XOR U17761 ( .A(b[63]), .B(n16916), .Z(n17134) );
  NANDN U17762 ( .A(n17134), .B(n38422), .Z(n16919) );
  NANDN U17763 ( .A(n16917), .B(n38423), .Z(n16918) );
  AND U17764 ( .A(n16919), .B(n16918), .Z(n17186) );
  XNOR U17765 ( .A(n17185), .B(n17186), .Z(n17187) );
  XOR U17766 ( .A(n17188), .B(n17187), .Z(n17192) );
  XNOR U17767 ( .A(n17191), .B(n17192), .Z(n17193) );
  XNOR U17768 ( .A(n17194), .B(n17193), .Z(n17046) );
  NANDN U17769 ( .A(n16921), .B(n16920), .Z(n16925) );
  NAND U17770 ( .A(n16923), .B(n16922), .Z(n16924) );
  NAND U17771 ( .A(n16925), .B(n16924), .Z(n17043) );
  NANDN U17772 ( .A(n16927), .B(n16926), .Z(n16931) );
  NAND U17773 ( .A(n16929), .B(n16928), .Z(n16930) );
  AND U17774 ( .A(n16931), .B(n16930), .Z(n17044) );
  XNOR U17775 ( .A(n17043), .B(n17044), .Z(n17045) );
  XOR U17776 ( .A(n17046), .B(n17045), .Z(n17150) );
  NANDN U17777 ( .A(n16933), .B(n16932), .Z(n16937) );
  OR U17778 ( .A(n16935), .B(n16934), .Z(n16936) );
  AND U17779 ( .A(n16937), .B(n16936), .Z(n17149) );
  XOR U17780 ( .A(n17150), .B(n17149), .Z(n17151) );
  XOR U17781 ( .A(n17152), .B(n17151), .Z(n17256) );
  XOR U17782 ( .A(n17257), .B(n17256), .Z(n17020) );
  XOR U17783 ( .A(n17019), .B(n17020), .Z(n17021) );
  XNOR U17784 ( .A(n17022), .B(n17021), .Z(n17015) );
  OR U17785 ( .A(n16939), .B(n16938), .Z(n16943) );
  NAND U17786 ( .A(n16941), .B(n16940), .Z(n16942) );
  AND U17787 ( .A(n16943), .B(n16942), .Z(n17013) );
  NAND U17788 ( .A(n16945), .B(n16944), .Z(n16949) );
  NANDN U17789 ( .A(n16947), .B(n16946), .Z(n16948) );
  NAND U17790 ( .A(n16949), .B(n16948), .Z(n17028) );
  NANDN U17791 ( .A(n16951), .B(n16950), .Z(n16955) );
  NAND U17792 ( .A(n16953), .B(n16952), .Z(n16954) );
  NAND U17793 ( .A(n16955), .B(n16954), .Z(n17026) );
  OR U17794 ( .A(n16957), .B(n16956), .Z(n16961) );
  NANDN U17795 ( .A(n16959), .B(n16958), .Z(n16960) );
  AND U17796 ( .A(n16961), .B(n16960), .Z(n17025) );
  XNOR U17797 ( .A(n17026), .B(n17025), .Z(n17027) );
  XOR U17798 ( .A(n17028), .B(n17027), .Z(n17014) );
  XNOR U17799 ( .A(n17015), .B(n17016), .Z(n17010) );
  NANDN U17800 ( .A(n16963), .B(n16962), .Z(n16967) );
  NAND U17801 ( .A(n16965), .B(n16964), .Z(n16966) );
  NAND U17802 ( .A(n16967), .B(n16966), .Z(n17008) );
  NANDN U17803 ( .A(n16969), .B(n16968), .Z(n16973) );
  NANDN U17804 ( .A(n16971), .B(n16970), .Z(n16972) );
  AND U17805 ( .A(n16973), .B(n16972), .Z(n17007) );
  XNOR U17806 ( .A(n17008), .B(n17007), .Z(n17009) );
  XNOR U17807 ( .A(n17010), .B(n17009), .Z(n17004) );
  NANDN U17808 ( .A(n16979), .B(n16978), .Z(n16983) );
  NANDN U17809 ( .A(n16981), .B(n16980), .Z(n16982) );
  NAND U17810 ( .A(n16983), .B(n16982), .Z(n17002) );
  XNOR U17811 ( .A(n17001), .B(n17002), .Z(n17003) );
  XNOR U17812 ( .A(n17004), .B(n17003), .Z(n16995) );
  OR U17813 ( .A(n16985), .B(n16984), .Z(n16989) );
  NANDN U17814 ( .A(n16987), .B(n16986), .Z(n16988) );
  NAND U17815 ( .A(n16989), .B(n16988), .Z(n16996) );
  XOR U17816 ( .A(n16995), .B(n16996), .Z(n16997) );
  XNOR U17817 ( .A(n16998), .B(n16997), .Z(n17282) );
  XNOR U17818 ( .A(n17282), .B(sreg[151]), .Z(n17284) );
  NAND U17819 ( .A(n16990), .B(sreg[150]), .Z(n16994) );
  OR U17820 ( .A(n16992), .B(n16991), .Z(n16993) );
  AND U17821 ( .A(n16994), .B(n16993), .Z(n17283) );
  XOR U17822 ( .A(n17284), .B(n17283), .Z(c[151]) );
  OR U17823 ( .A(n16996), .B(n16995), .Z(n17000) );
  NAND U17824 ( .A(n16998), .B(n16997), .Z(n16999) );
  NAND U17825 ( .A(n17000), .B(n16999), .Z(n17290) );
  NANDN U17826 ( .A(n17002), .B(n17001), .Z(n17006) );
  NANDN U17827 ( .A(n17004), .B(n17003), .Z(n17005) );
  NAND U17828 ( .A(n17006), .B(n17005), .Z(n17288) );
  NANDN U17829 ( .A(n17008), .B(n17007), .Z(n17012) );
  NANDN U17830 ( .A(n17010), .B(n17009), .Z(n17011) );
  NAND U17831 ( .A(n17012), .B(n17011), .Z(n17561) );
  OR U17832 ( .A(n17014), .B(n17013), .Z(n17018) );
  NANDN U17833 ( .A(n17016), .B(n17015), .Z(n17017) );
  NAND U17834 ( .A(n17018), .B(n17017), .Z(n17562) );
  XNOR U17835 ( .A(n17561), .B(n17562), .Z(n17563) );
  OR U17836 ( .A(n17020), .B(n17019), .Z(n17024) );
  NAND U17837 ( .A(n17022), .B(n17021), .Z(n17023) );
  NAND U17838 ( .A(n17024), .B(n17023), .Z(n17555) );
  NANDN U17839 ( .A(n17026), .B(n17025), .Z(n17030) );
  NANDN U17840 ( .A(n17028), .B(n17027), .Z(n17029) );
  NAND U17841 ( .A(n17030), .B(n17029), .Z(n17556) );
  XNOR U17842 ( .A(n17555), .B(n17556), .Z(n17557) );
  NANDN U17843 ( .A(n17032), .B(n17031), .Z(n17036) );
  NAND U17844 ( .A(n17034), .B(n17033), .Z(n17035) );
  AND U17845 ( .A(n17036), .B(n17035), .Z(n17312) );
  NANDN U17846 ( .A(n17038), .B(n17037), .Z(n17042) );
  OR U17847 ( .A(n17040), .B(n17039), .Z(n17041) );
  NAND U17848 ( .A(n17042), .B(n17041), .Z(n17309) );
  NANDN U17849 ( .A(n17044), .B(n17043), .Z(n17048) );
  NAND U17850 ( .A(n17046), .B(n17045), .Z(n17047) );
  NAND U17851 ( .A(n17048), .B(n17047), .Z(n17310) );
  XNOR U17852 ( .A(n17309), .B(n17310), .Z(n17311) );
  XNOR U17853 ( .A(n17312), .B(n17311), .Z(n17531) );
  NANDN U17854 ( .A(n17050), .B(n17049), .Z(n17054) );
  OR U17855 ( .A(n17052), .B(n17051), .Z(n17053) );
  AND U17856 ( .A(n17054), .B(n17053), .Z(n17532) );
  XNOR U17857 ( .A(n17531), .B(n17532), .Z(n17534) );
  NANDN U17858 ( .A(n17056), .B(n17055), .Z(n17060) );
  NAND U17859 ( .A(n17058), .B(n17057), .Z(n17059) );
  NAND U17860 ( .A(n17060), .B(n17059), .Z(n17316) );
  XOR U17861 ( .A(b[37]), .B(n25134), .Z(n17364) );
  NANDN U17862 ( .A(n17364), .B(n36311), .Z(n17063) );
  NANDN U17863 ( .A(n17061), .B(n36309), .Z(n17062) );
  NAND U17864 ( .A(n17063), .B(n17062), .Z(n17397) );
  XOR U17865 ( .A(a[84]), .B(n968), .Z(n17367) );
  OR U17866 ( .A(n17367), .B(n29363), .Z(n17066) );
  NANDN U17867 ( .A(n17064), .B(n29864), .Z(n17065) );
  NAND U17868 ( .A(n17066), .B(n17065), .Z(n17394) );
  XOR U17869 ( .A(n33628), .B(n967), .Z(n17370) );
  NAND U17870 ( .A(n17370), .B(n28939), .Z(n17069) );
  NAND U17871 ( .A(n28938), .B(n17067), .Z(n17068) );
  AND U17872 ( .A(n17069), .B(n17068), .Z(n17395) );
  XNOR U17873 ( .A(n17394), .B(n17395), .Z(n17396) );
  XOR U17874 ( .A(n17397), .B(n17396), .Z(n17319) );
  XOR U17875 ( .A(b[13]), .B(n31363), .Z(n17373) );
  OR U17876 ( .A(n17373), .B(n31550), .Z(n17072) );
  NANDN U17877 ( .A(n17070), .B(n31874), .Z(n17071) );
  NAND U17878 ( .A(n17072), .B(n17071), .Z(n17457) );
  NAND U17879 ( .A(n34848), .B(n17073), .Z(n17075) );
  XNOR U17880 ( .A(n35375), .B(a[62]), .Z(n17376) );
  NAND U17881 ( .A(n34618), .B(n17376), .Z(n17074) );
  NAND U17882 ( .A(n17075), .B(n17074), .Z(n17454) );
  NAND U17883 ( .A(n35188), .B(n17076), .Z(n17078) );
  XOR U17884 ( .A(n35540), .B(n27436), .Z(n17379) );
  NANDN U17885 ( .A(n34968), .B(n17379), .Z(n17077) );
  AND U17886 ( .A(n17078), .B(n17077), .Z(n17455) );
  XNOR U17887 ( .A(n17454), .B(n17455), .Z(n17456) );
  XOR U17888 ( .A(n17457), .B(n17456), .Z(n17320) );
  XNOR U17889 ( .A(n17319), .B(n17320), .Z(n17322) );
  NANDN U17890 ( .A(n17080), .B(n17079), .Z(n17084) );
  NAND U17891 ( .A(n17082), .B(n17081), .Z(n17083) );
  NAND U17892 ( .A(n17084), .B(n17083), .Z(n17321) );
  XNOR U17893 ( .A(n17322), .B(n17321), .Z(n17314) );
  NANDN U17894 ( .A(n17086), .B(n17085), .Z(n17090) );
  NAND U17895 ( .A(n17088), .B(n17087), .Z(n17089) );
  NAND U17896 ( .A(n17090), .B(n17089), .Z(n17510) );
  NAND U17897 ( .A(a[24]), .B(b[63]), .Z(n17524) );
  NANDN U17898 ( .A(n17091), .B(n38369), .Z(n17093) );
  XOR U17899 ( .A(b[61]), .B(n17702), .Z(n17358) );
  OR U17900 ( .A(n17358), .B(n38371), .Z(n17092) );
  NAND U17901 ( .A(n17093), .B(n17092), .Z(n17522) );
  NANDN U17902 ( .A(n17094), .B(n35311), .Z(n17096) );
  XOR U17903 ( .A(b[31]), .B(n26347), .Z(n17361) );
  NANDN U17904 ( .A(n17361), .B(n35313), .Z(n17095) );
  AND U17905 ( .A(n17096), .B(n17095), .Z(n17521) );
  XNOR U17906 ( .A(n17522), .B(n17521), .Z(n17523) );
  XOR U17907 ( .A(n17524), .B(n17523), .Z(n17508) );
  NAND U17908 ( .A(n33283), .B(n17097), .Z(n17099) );
  XOR U17909 ( .A(n33020), .B(n30379), .Z(n17343) );
  NANDN U17910 ( .A(n33021), .B(n17343), .Z(n17098) );
  NAND U17911 ( .A(n17099), .B(n17098), .Z(n17421) );
  XNOR U17912 ( .A(b[21]), .B(a[68]), .Z(n17346) );
  OR U17913 ( .A(n17346), .B(n33634), .Z(n17102) );
  NANDN U17914 ( .A(n17100), .B(n33464), .Z(n17101) );
  NAND U17915 ( .A(n17102), .B(n17101), .Z(n17418) );
  NAND U17916 ( .A(n34044), .B(n17103), .Z(n17105) );
  XOR U17917 ( .A(n34510), .B(n28701), .Z(n17349) );
  NANDN U17918 ( .A(n33867), .B(n17349), .Z(n17104) );
  AND U17919 ( .A(n17105), .B(n17104), .Z(n17419) );
  XNOR U17920 ( .A(n17418), .B(n17419), .Z(n17420) );
  XNOR U17921 ( .A(n17421), .B(n17420), .Z(n17509) );
  XNOR U17922 ( .A(n17508), .B(n17509), .Z(n17511) );
  XNOR U17923 ( .A(n17510), .B(n17511), .Z(n17313) );
  XOR U17924 ( .A(n17314), .B(n17313), .Z(n17315) );
  XOR U17925 ( .A(n17316), .B(n17315), .Z(n17432) );
  NANDN U17926 ( .A(n17107), .B(n17106), .Z(n17111) );
  NANDN U17927 ( .A(n17109), .B(n17108), .Z(n17110) );
  NAND U17928 ( .A(n17111), .B(n17110), .Z(n17431) );
  NANDN U17929 ( .A(n17113), .B(n17112), .Z(n17117) );
  NAND U17930 ( .A(n17115), .B(n17114), .Z(n17116) );
  NAND U17931 ( .A(n17117), .B(n17116), .Z(n17328) );
  XNOR U17932 ( .A(b[41]), .B(a[48]), .Z(n17400) );
  OR U17933 ( .A(n17400), .B(n36905), .Z(n17120) );
  NANDN U17934 ( .A(n17118), .B(n36807), .Z(n17119) );
  NAND U17935 ( .A(n17120), .B(n17119), .Z(n17427) );
  XOR U17936 ( .A(b[57]), .B(n18841), .Z(n17403) );
  OR U17937 ( .A(n17403), .B(n965), .Z(n17123) );
  NANDN U17938 ( .A(n17121), .B(n38194), .Z(n17122) );
  NAND U17939 ( .A(n17123), .B(n17122), .Z(n17424) );
  NAND U17940 ( .A(n38326), .B(n17124), .Z(n17126) );
  XOR U17941 ( .A(n38400), .B(n18804), .Z(n17406) );
  NANDN U17942 ( .A(n38273), .B(n17406), .Z(n17125) );
  AND U17943 ( .A(n17126), .B(n17125), .Z(n17425) );
  XNOR U17944 ( .A(n17424), .B(n17425), .Z(n17426) );
  XOR U17945 ( .A(n17427), .B(n17426), .Z(n17472) );
  XOR U17946 ( .A(b[33]), .B(n25860), .Z(n17409) );
  NANDN U17947 ( .A(n17409), .B(n35620), .Z(n17129) );
  NANDN U17948 ( .A(n17127), .B(n35621), .Z(n17128) );
  NAND U17949 ( .A(n17129), .B(n17128), .Z(n17469) );
  NANDN U17950 ( .A(n966), .B(a[88]), .Z(n17130) );
  XOR U17951 ( .A(n29232), .B(n17130), .Z(n17132) );
  NANDN U17952 ( .A(b[0]), .B(a[87]), .Z(n17131) );
  AND U17953 ( .A(n17132), .B(n17131), .Z(n17466) );
  XOR U17954 ( .A(b[63]), .B(n17133), .Z(n17415) );
  NANDN U17955 ( .A(n17415), .B(n38422), .Z(n17136) );
  NANDN U17956 ( .A(n17134), .B(n38423), .Z(n17135) );
  AND U17957 ( .A(n17136), .B(n17135), .Z(n17467) );
  XNOR U17958 ( .A(n17466), .B(n17467), .Z(n17468) );
  XOR U17959 ( .A(n17469), .B(n17468), .Z(n17473) );
  XNOR U17960 ( .A(n17472), .B(n17473), .Z(n17475) );
  NANDN U17961 ( .A(n17138), .B(n17137), .Z(n17142) );
  NAND U17962 ( .A(n17140), .B(n17139), .Z(n17141) );
  NAND U17963 ( .A(n17142), .B(n17141), .Z(n17474) );
  XOR U17964 ( .A(n17475), .B(n17474), .Z(n17325) );
  NANDN U17965 ( .A(n17144), .B(n17143), .Z(n17148) );
  NAND U17966 ( .A(n17146), .B(n17145), .Z(n17147) );
  AND U17967 ( .A(n17148), .B(n17147), .Z(n17326) );
  XOR U17968 ( .A(n17325), .B(n17326), .Z(n17327) );
  XNOR U17969 ( .A(n17328), .B(n17327), .Z(n17430) );
  XNOR U17970 ( .A(n17431), .B(n17430), .Z(n17433) );
  XNOR U17971 ( .A(n17432), .B(n17433), .Z(n17533) );
  XOR U17972 ( .A(n17534), .B(n17533), .Z(n17537) );
  OR U17973 ( .A(n17150), .B(n17149), .Z(n17154) );
  NAND U17974 ( .A(n17152), .B(n17151), .Z(n17153) );
  NAND U17975 ( .A(n17154), .B(n17153), .Z(n17294) );
  XOR U17976 ( .A(b[15]), .B(n31372), .Z(n17436) );
  OR U17977 ( .A(n17436), .B(n32010), .Z(n17157) );
  NANDN U17978 ( .A(n17155), .B(n32011), .Z(n17156) );
  NAND U17979 ( .A(n17157), .B(n17156), .Z(n17355) );
  XOR U17980 ( .A(b[25]), .B(a[64]), .Z(n17439) );
  NANDN U17981 ( .A(n34219), .B(n17439), .Z(n17160) );
  NAND U17982 ( .A(n34217), .B(n17158), .Z(n17159) );
  NAND U17983 ( .A(n17160), .B(n17159), .Z(n17352) );
  XNOR U17984 ( .A(b[17]), .B(a[72]), .Z(n17442) );
  NANDN U17985 ( .A(n17442), .B(n32543), .Z(n17163) );
  NANDN U17986 ( .A(n17161), .B(n32541), .Z(n17162) );
  AND U17987 ( .A(n17163), .B(n17162), .Z(n17353) );
  XNOR U17988 ( .A(n17352), .B(n17353), .Z(n17354) );
  XNOR U17989 ( .A(n17355), .B(n17354), .Z(n17388) );
  XOR U17990 ( .A(b[39]), .B(n24671), .Z(n17445) );
  NANDN U17991 ( .A(n17445), .B(n36553), .Z(n17166) );
  NANDN U17992 ( .A(n17164), .B(n36643), .Z(n17165) );
  NAND U17993 ( .A(n17166), .B(n17165), .Z(n17385) );
  XOR U17994 ( .A(b[51]), .B(n20686), .Z(n17448) );
  NANDN U17995 ( .A(n17448), .B(n37803), .Z(n17169) );
  NANDN U17996 ( .A(n17167), .B(n37802), .Z(n17168) );
  NAND U17997 ( .A(n17169), .B(n17168), .Z(n17382) );
  XOR U17998 ( .A(b[53]), .B(n19980), .Z(n17451) );
  NANDN U17999 ( .A(n17451), .B(n37940), .Z(n17172) );
  NANDN U18000 ( .A(n17170), .B(n37941), .Z(n17171) );
  AND U18001 ( .A(n17172), .B(n17171), .Z(n17383) );
  XNOR U18002 ( .A(n17382), .B(n17383), .Z(n17384) );
  XOR U18003 ( .A(n17385), .B(n17384), .Z(n17389) );
  XOR U18004 ( .A(n17388), .B(n17389), .Z(n17391) );
  NANDN U18005 ( .A(n17174), .B(n17173), .Z(n17178) );
  NAND U18006 ( .A(n17176), .B(n17175), .Z(n17177) );
  NAND U18007 ( .A(n17178), .B(n17177), .Z(n17390) );
  XNOR U18008 ( .A(n17391), .B(n17390), .Z(n17481) );
  NANDN U18009 ( .A(n17180), .B(n17179), .Z(n17184) );
  NAND U18010 ( .A(n17182), .B(n17181), .Z(n17183) );
  NAND U18011 ( .A(n17184), .B(n17183), .Z(n17478) );
  NANDN U18012 ( .A(n17186), .B(n17185), .Z(n17190) );
  NAND U18013 ( .A(n17188), .B(n17187), .Z(n17189) );
  AND U18014 ( .A(n17190), .B(n17189), .Z(n17479) );
  XNOR U18015 ( .A(n17478), .B(n17479), .Z(n17480) );
  XNOR U18016 ( .A(n17481), .B(n17480), .Z(n17303) );
  OR U18017 ( .A(n17192), .B(n17191), .Z(n17196) );
  OR U18018 ( .A(n17194), .B(n17193), .Z(n17195) );
  AND U18019 ( .A(n17196), .B(n17195), .Z(n17304) );
  XNOR U18020 ( .A(n17303), .B(n17304), .Z(n17305) );
  NANDN U18021 ( .A(n17198), .B(n17197), .Z(n17202) );
  NAND U18022 ( .A(n17200), .B(n17199), .Z(n17201) );
  AND U18023 ( .A(n17202), .B(n17201), .Z(n17306) );
  XNOR U18024 ( .A(n17305), .B(n17306), .Z(n17291) );
  OR U18025 ( .A(n17204), .B(n17203), .Z(n17208) );
  OR U18026 ( .A(n17206), .B(n17205), .Z(n17207) );
  NAND U18027 ( .A(n17208), .B(n17207), .Z(n17298) );
  XOR U18028 ( .A(a[78]), .B(n970), .Z(n17484) );
  OR U18029 ( .A(n17484), .B(n31369), .Z(n17211) );
  NANDN U18030 ( .A(n17209), .B(n31119), .Z(n17210) );
  NAND U18031 ( .A(n17211), .B(n17210), .Z(n17505) );
  XOR U18032 ( .A(b[43]), .B(n22964), .Z(n17487) );
  NANDN U18033 ( .A(n17487), .B(n37068), .Z(n17214) );
  NANDN U18034 ( .A(n17212), .B(n37069), .Z(n17213) );
  NAND U18035 ( .A(n17214), .B(n17213), .Z(n17502) );
  XNOR U18036 ( .A(b[45]), .B(a[44]), .Z(n17490) );
  NANDN U18037 ( .A(n17490), .B(n37261), .Z(n17217) );
  NANDN U18038 ( .A(n17215), .B(n37262), .Z(n17216) );
  AND U18039 ( .A(n17217), .B(n17216), .Z(n17503) );
  XNOR U18040 ( .A(n17502), .B(n17503), .Z(n17504) );
  XNOR U18041 ( .A(n17505), .B(n17504), .Z(n17340) );
  NANDN U18042 ( .A(n17218), .B(n37652), .Z(n17220) );
  XOR U18043 ( .A(b[49]), .B(n21149), .Z(n17493) );
  OR U18044 ( .A(n17493), .B(n37756), .Z(n17219) );
  NAND U18045 ( .A(n17220), .B(n17219), .Z(n17529) );
  NANDN U18046 ( .A(n17221), .B(n37469), .Z(n17223) );
  XNOR U18047 ( .A(n978), .B(a[42]), .Z(n17496) );
  NAND U18048 ( .A(n17496), .B(n37471), .Z(n17222) );
  NAND U18049 ( .A(n17223), .B(n17222), .Z(n17527) );
  NAND U18050 ( .A(n30846), .B(n17224), .Z(n17226) );
  XNOR U18051 ( .A(n32814), .B(b[9]), .Z(n17499) );
  NAND U18052 ( .A(n30509), .B(n17499), .Z(n17225) );
  NAND U18053 ( .A(n17226), .B(n17225), .Z(n17528) );
  XNOR U18054 ( .A(n17527), .B(n17528), .Z(n17530) );
  XOR U18055 ( .A(n17529), .B(n17530), .Z(n17337) );
  NANDN U18056 ( .A(n17228), .B(n17227), .Z(n17232) );
  NAND U18057 ( .A(n17230), .B(n17229), .Z(n17231) );
  NAND U18058 ( .A(n17232), .B(n17231), .Z(n17338) );
  XNOR U18059 ( .A(n17337), .B(n17338), .Z(n17339) );
  XOR U18060 ( .A(n17340), .B(n17339), .Z(n17297) );
  XNOR U18061 ( .A(n17298), .B(n17297), .Z(n17300) );
  XNOR U18062 ( .A(b[35]), .B(a[54]), .Z(n17512) );
  NANDN U18063 ( .A(n17512), .B(n35985), .Z(n17235) );
  NANDN U18064 ( .A(n17233), .B(n35986), .Z(n17234) );
  NAND U18065 ( .A(n17235), .B(n17234), .Z(n17463) );
  XOR U18066 ( .A(n32815), .B(n31123), .Z(n17515) );
  NAND U18067 ( .A(n17515), .B(n29949), .Z(n17238) );
  NAND U18068 ( .A(n29948), .B(n17236), .Z(n17237) );
  NAND U18069 ( .A(n17238), .B(n17237), .Z(n17460) );
  XOR U18070 ( .A(b[55]), .B(n19513), .Z(n17518) );
  NANDN U18071 ( .A(n17518), .B(n38075), .Z(n17241) );
  NANDN U18072 ( .A(n17239), .B(n38073), .Z(n17240) );
  AND U18073 ( .A(n17241), .B(n17240), .Z(n17461) );
  XNOR U18074 ( .A(n17460), .B(n17461), .Z(n17462) );
  XNOR U18075 ( .A(n17463), .B(n17462), .Z(n17334) );
  NANDN U18076 ( .A(n17243), .B(n17242), .Z(n17247) );
  NAND U18077 ( .A(n17245), .B(n17244), .Z(n17246) );
  NAND U18078 ( .A(n17247), .B(n17246), .Z(n17331) );
  NANDN U18079 ( .A(n17249), .B(n17248), .Z(n17253) );
  NAND U18080 ( .A(n17251), .B(n17250), .Z(n17252) );
  NAND U18081 ( .A(n17253), .B(n17252), .Z(n17332) );
  XNOR U18082 ( .A(n17331), .B(n17332), .Z(n17333) );
  XOR U18083 ( .A(n17334), .B(n17333), .Z(n17299) );
  XOR U18084 ( .A(n17300), .B(n17299), .Z(n17292) );
  XOR U18085 ( .A(n17291), .B(n17292), .Z(n17293) );
  XOR U18086 ( .A(n17294), .B(n17293), .Z(n17538) );
  XNOR U18087 ( .A(n17537), .B(n17538), .Z(n17539) );
  NAND U18088 ( .A(n17255), .B(n17254), .Z(n17259) );
  NANDN U18089 ( .A(n17257), .B(n17256), .Z(n17258) );
  NAND U18090 ( .A(n17259), .B(n17258), .Z(n17540) );
  XOR U18091 ( .A(n17539), .B(n17540), .Z(n17551) );
  NANDN U18092 ( .A(n17261), .B(n17260), .Z(n17265) );
  NAND U18093 ( .A(n17263), .B(n17262), .Z(n17264) );
  NAND U18094 ( .A(n17265), .B(n17264), .Z(n17546) );
  NANDN U18095 ( .A(n17267), .B(n17266), .Z(n17271) );
  NAND U18096 ( .A(n17269), .B(n17268), .Z(n17270) );
  NAND U18097 ( .A(n17271), .B(n17270), .Z(n17544) );
  XNOR U18098 ( .A(n17544), .B(n17543), .Z(n17545) );
  XNOR U18099 ( .A(n17546), .B(n17545), .Z(n17549) );
  NANDN U18100 ( .A(n17277), .B(n17276), .Z(n17281) );
  NANDN U18101 ( .A(n17279), .B(n17278), .Z(n17280) );
  AND U18102 ( .A(n17281), .B(n17280), .Z(n17550) );
  XOR U18103 ( .A(n17551), .B(n17552), .Z(n17558) );
  XNOR U18104 ( .A(n17557), .B(n17558), .Z(n17564) );
  XOR U18105 ( .A(n17563), .B(n17564), .Z(n17287) );
  XNOR U18106 ( .A(n17288), .B(n17287), .Z(n17289) );
  XNOR U18107 ( .A(n17290), .B(n17289), .Z(n17567) );
  XNOR U18108 ( .A(n17567), .B(sreg[152]), .Z(n17569) );
  NAND U18109 ( .A(n17282), .B(sreg[151]), .Z(n17286) );
  OR U18110 ( .A(n17284), .B(n17283), .Z(n17285) );
  AND U18111 ( .A(n17286), .B(n17285), .Z(n17568) );
  XOR U18112 ( .A(n17569), .B(n17568), .Z(c[152]) );
  OR U18113 ( .A(n17292), .B(n17291), .Z(n17296) );
  NAND U18114 ( .A(n17294), .B(n17293), .Z(n17295) );
  NAND U18115 ( .A(n17296), .B(n17295), .Z(n17837) );
  NAND U18116 ( .A(n17298), .B(n17297), .Z(n17302) );
  NANDN U18117 ( .A(n17300), .B(n17299), .Z(n17301) );
  NAND U18118 ( .A(n17302), .B(n17301), .Z(n17834) );
  NANDN U18119 ( .A(n17304), .B(n17303), .Z(n17308) );
  NAND U18120 ( .A(n17306), .B(n17305), .Z(n17307) );
  NAND U18121 ( .A(n17308), .B(n17307), .Z(n17832) );
  XNOR U18122 ( .A(n17832), .B(n17831), .Z(n17833) );
  XOR U18123 ( .A(n17834), .B(n17833), .Z(n17838) );
  XOR U18124 ( .A(n17837), .B(n17838), .Z(n17839) );
  NAND U18125 ( .A(n17314), .B(n17313), .Z(n17318) );
  NANDN U18126 ( .A(n17316), .B(n17315), .Z(n17317) );
  NAND U18127 ( .A(n17318), .B(n17317), .Z(n17821) );
  OR U18128 ( .A(n17320), .B(n17319), .Z(n17324) );
  OR U18129 ( .A(n17322), .B(n17321), .Z(n17323) );
  NAND U18130 ( .A(n17324), .B(n17323), .Z(n17586) );
  NAND U18131 ( .A(n17326), .B(n17325), .Z(n17330) );
  NANDN U18132 ( .A(n17328), .B(n17327), .Z(n17329) );
  NAND U18133 ( .A(n17330), .B(n17329), .Z(n17584) );
  NANDN U18134 ( .A(n17332), .B(n17331), .Z(n17336) );
  NAND U18135 ( .A(n17334), .B(n17333), .Z(n17335) );
  AND U18136 ( .A(n17336), .B(n17335), .Z(n17585) );
  XNOR U18137 ( .A(n17584), .B(n17585), .Z(n17587) );
  XNOR U18138 ( .A(n17586), .B(n17587), .Z(n17822) );
  XOR U18139 ( .A(n17821), .B(n17822), .Z(n17823) );
  NANDN U18140 ( .A(n17338), .B(n17337), .Z(n17342) );
  NAND U18141 ( .A(n17340), .B(n17339), .Z(n17341) );
  NAND U18142 ( .A(n17342), .B(n17341), .Z(n17602) );
  NAND U18143 ( .A(n33283), .B(n17343), .Z(n17345) );
  XOR U18144 ( .A(n33020), .B(n30543), .Z(n17630) );
  NANDN U18145 ( .A(n33021), .B(n17630), .Z(n17344) );
  NAND U18146 ( .A(n17345), .B(n17344), .Z(n17709) );
  XOR U18147 ( .A(b[21]), .B(a[69]), .Z(n17633) );
  NANDN U18148 ( .A(n33634), .B(n17633), .Z(n17348) );
  NANDN U18149 ( .A(n17346), .B(n33464), .Z(n17347) );
  NAND U18150 ( .A(n17348), .B(n17347), .Z(n17706) );
  NAND U18151 ( .A(n34044), .B(n17349), .Z(n17351) );
  XOR U18152 ( .A(n34510), .B(n29372), .Z(n17636) );
  NANDN U18153 ( .A(n33867), .B(n17636), .Z(n17350) );
  AND U18154 ( .A(n17351), .B(n17350), .Z(n17707) );
  XNOR U18155 ( .A(n17706), .B(n17707), .Z(n17708) );
  XOR U18156 ( .A(n17709), .B(n17708), .Z(n17724) );
  NANDN U18157 ( .A(n17353), .B(n17352), .Z(n17357) );
  NAND U18158 ( .A(n17355), .B(n17354), .Z(n17356) );
  NAND U18159 ( .A(n17357), .B(n17356), .Z(n17725) );
  XNOR U18160 ( .A(n17724), .B(n17725), .Z(n17727) );
  NAND U18161 ( .A(a[25]), .B(b[63]), .Z(n17766) );
  NANDN U18162 ( .A(n17358), .B(n38369), .Z(n17360) );
  XOR U18163 ( .A(b[61]), .B(n18003), .Z(n17645) );
  OR U18164 ( .A(n17645), .B(n38371), .Z(n17359) );
  NAND U18165 ( .A(n17360), .B(n17359), .Z(n17764) );
  NANDN U18166 ( .A(n17361), .B(n35311), .Z(n17363) );
  XNOR U18167 ( .A(b[31]), .B(a[59]), .Z(n17648) );
  NANDN U18168 ( .A(n17648), .B(n35313), .Z(n17362) );
  AND U18169 ( .A(n17363), .B(n17362), .Z(n17763) );
  XNOR U18170 ( .A(n17764), .B(n17763), .Z(n17765) );
  XNOR U18171 ( .A(n17766), .B(n17765), .Z(n17726) );
  XNOR U18172 ( .A(n17727), .B(n17726), .Z(n17600) );
  XOR U18173 ( .A(b[37]), .B(n25001), .Z(n17651) );
  NANDN U18174 ( .A(n17651), .B(n36311), .Z(n17366) );
  NANDN U18175 ( .A(n17364), .B(n36309), .Z(n17365) );
  NAND U18176 ( .A(n17366), .B(n17365), .Z(n17684) );
  XNOR U18177 ( .A(a[85]), .B(b[5]), .Z(n17654) );
  OR U18178 ( .A(n17654), .B(n29363), .Z(n17369) );
  NANDN U18179 ( .A(n17367), .B(n29864), .Z(n17368) );
  NAND U18180 ( .A(n17369), .B(n17368), .Z(n17681) );
  XNOR U18181 ( .A(a[87]), .B(n967), .Z(n17657) );
  NAND U18182 ( .A(n17657), .B(n28939), .Z(n17372) );
  NAND U18183 ( .A(n28938), .B(n17370), .Z(n17371) );
  AND U18184 ( .A(n17372), .B(n17371), .Z(n17682) );
  XNOR U18185 ( .A(n17681), .B(n17682), .Z(n17683) );
  XOR U18186 ( .A(n17684), .B(n17683), .Z(n17621) );
  XNOR U18187 ( .A(b[13]), .B(a[77]), .Z(n17660) );
  OR U18188 ( .A(n17660), .B(n31550), .Z(n17375) );
  NANDN U18189 ( .A(n17373), .B(n31874), .Z(n17374) );
  NAND U18190 ( .A(n17375), .B(n17374), .Z(n17812) );
  NAND U18191 ( .A(n34848), .B(n17376), .Z(n17378) );
  XNOR U18192 ( .A(n35375), .B(a[63]), .Z(n17663) );
  NAND U18193 ( .A(n34618), .B(n17663), .Z(n17377) );
  NAND U18194 ( .A(n17378), .B(n17377), .Z(n17809) );
  NAND U18195 ( .A(n35188), .B(n17379), .Z(n17381) );
  XOR U18196 ( .A(n35540), .B(n27773), .Z(n17666) );
  NANDN U18197 ( .A(n34968), .B(n17666), .Z(n17380) );
  AND U18198 ( .A(n17381), .B(n17380), .Z(n17810) );
  XNOR U18199 ( .A(n17809), .B(n17810), .Z(n17811) );
  XOR U18200 ( .A(n17812), .B(n17811), .Z(n17619) );
  NANDN U18201 ( .A(n17383), .B(n17382), .Z(n17387) );
  NAND U18202 ( .A(n17385), .B(n17384), .Z(n17386) );
  AND U18203 ( .A(n17387), .B(n17386), .Z(n17618) );
  XOR U18204 ( .A(n17619), .B(n17618), .Z(n17620) );
  XOR U18205 ( .A(n17621), .B(n17620), .Z(n17601) );
  XOR U18206 ( .A(n17600), .B(n17601), .Z(n17603) );
  XNOR U18207 ( .A(n17602), .B(n17603), .Z(n17720) );
  NANDN U18208 ( .A(n17389), .B(n17388), .Z(n17393) );
  OR U18209 ( .A(n17391), .B(n17390), .Z(n17392) );
  NAND U18210 ( .A(n17393), .B(n17392), .Z(n17719) );
  NANDN U18211 ( .A(n17395), .B(n17394), .Z(n17399) );
  NAND U18212 ( .A(n17397), .B(n17396), .Z(n17398) );
  NAND U18213 ( .A(n17399), .B(n17398), .Z(n17615) );
  XNOR U18214 ( .A(b[41]), .B(a[49]), .Z(n17687) );
  OR U18215 ( .A(n17687), .B(n36905), .Z(n17402) );
  NANDN U18216 ( .A(n17400), .B(n36807), .Z(n17401) );
  NAND U18217 ( .A(n17402), .B(n17401), .Z(n17715) );
  XOR U18218 ( .A(b[57]), .B(n19656), .Z(n17690) );
  OR U18219 ( .A(n17690), .B(n965), .Z(n17405) );
  NANDN U18220 ( .A(n17403), .B(n38194), .Z(n17404) );
  NAND U18221 ( .A(n17405), .B(n17404), .Z(n17712) );
  NAND U18222 ( .A(n38326), .B(n17406), .Z(n17408) );
  XOR U18223 ( .A(n38400), .B(n18639), .Z(n17693) );
  NANDN U18224 ( .A(n38273), .B(n17693), .Z(n17407) );
  AND U18225 ( .A(n17408), .B(n17407), .Z(n17713) );
  XNOR U18226 ( .A(n17712), .B(n17713), .Z(n17714) );
  XOR U18227 ( .A(n17715), .B(n17714), .Z(n17775) );
  XOR U18228 ( .A(b[33]), .B(n26122), .Z(n17696) );
  NANDN U18229 ( .A(n17696), .B(n35620), .Z(n17411) );
  NANDN U18230 ( .A(n17409), .B(n35621), .Z(n17410) );
  NAND U18231 ( .A(n17411), .B(n17410), .Z(n17788) );
  NANDN U18232 ( .A(n966), .B(a[89]), .Z(n17412) );
  XOR U18233 ( .A(n29232), .B(n17412), .Z(n17414) );
  IV U18234 ( .A(a[88]), .Z(n34048) );
  NANDN U18235 ( .A(n34048), .B(n966), .Z(n17413) );
  AND U18236 ( .A(n17414), .B(n17413), .Z(n17785) );
  XOR U18237 ( .A(b[63]), .B(n17960), .Z(n17703) );
  NANDN U18238 ( .A(n17703), .B(n38422), .Z(n17417) );
  NANDN U18239 ( .A(n17415), .B(n38423), .Z(n17416) );
  AND U18240 ( .A(n17417), .B(n17416), .Z(n17786) );
  XNOR U18241 ( .A(n17785), .B(n17786), .Z(n17787) );
  XOR U18242 ( .A(n17788), .B(n17787), .Z(n17776) );
  XNOR U18243 ( .A(n17775), .B(n17776), .Z(n17778) );
  NANDN U18244 ( .A(n17419), .B(n17418), .Z(n17423) );
  NAND U18245 ( .A(n17421), .B(n17420), .Z(n17422) );
  AND U18246 ( .A(n17423), .B(n17422), .Z(n17777) );
  XNOR U18247 ( .A(n17778), .B(n17777), .Z(n17612) );
  NANDN U18248 ( .A(n17425), .B(n17424), .Z(n17429) );
  NAND U18249 ( .A(n17427), .B(n17426), .Z(n17428) );
  AND U18250 ( .A(n17429), .B(n17428), .Z(n17613) );
  XOR U18251 ( .A(n17612), .B(n17613), .Z(n17614) );
  XNOR U18252 ( .A(n17615), .B(n17614), .Z(n17718) );
  XNOR U18253 ( .A(n17719), .B(n17718), .Z(n17721) );
  XNOR U18254 ( .A(n17720), .B(n17721), .Z(n17824) );
  XNOR U18255 ( .A(n17823), .B(n17824), .Z(n17827) );
  NAND U18256 ( .A(n17431), .B(n17430), .Z(n17435) );
  NANDN U18257 ( .A(n17433), .B(n17432), .Z(n17434) );
  NAND U18258 ( .A(n17435), .B(n17434), .Z(n17596) );
  XNOR U18259 ( .A(b[15]), .B(a[75]), .Z(n17791) );
  OR U18260 ( .A(n17791), .B(n32010), .Z(n17438) );
  NANDN U18261 ( .A(n17436), .B(n32011), .Z(n17437) );
  NAND U18262 ( .A(n17438), .B(n17437), .Z(n17642) );
  XNOR U18263 ( .A(b[25]), .B(n28403), .Z(n17794) );
  NANDN U18264 ( .A(n34219), .B(n17794), .Z(n17441) );
  NAND U18265 ( .A(n34217), .B(n17439), .Z(n17440) );
  NAND U18266 ( .A(n17441), .B(n17440), .Z(n17639) );
  XOR U18267 ( .A(b[17]), .B(a[73]), .Z(n17797) );
  NAND U18268 ( .A(n17797), .B(n32543), .Z(n17444) );
  NANDN U18269 ( .A(n17442), .B(n32541), .Z(n17443) );
  AND U18270 ( .A(n17444), .B(n17443), .Z(n17640) );
  XNOR U18271 ( .A(n17639), .B(n17640), .Z(n17641) );
  XNOR U18272 ( .A(n17642), .B(n17641), .Z(n17675) );
  XOR U18273 ( .A(b[39]), .B(n24288), .Z(n17800) );
  NANDN U18274 ( .A(n17800), .B(n36553), .Z(n17447) );
  NANDN U18275 ( .A(n17445), .B(n36643), .Z(n17446) );
  NAND U18276 ( .A(n17447), .B(n17446), .Z(n17672) );
  XOR U18277 ( .A(b[51]), .B(n20867), .Z(n17803) );
  NANDN U18278 ( .A(n17803), .B(n37803), .Z(n17450) );
  NANDN U18279 ( .A(n17448), .B(n37802), .Z(n17449) );
  NAND U18280 ( .A(n17450), .B(n17449), .Z(n17669) );
  XOR U18281 ( .A(b[53]), .B(n20352), .Z(n17806) );
  NANDN U18282 ( .A(n17806), .B(n37940), .Z(n17453) );
  NANDN U18283 ( .A(n17451), .B(n37941), .Z(n17452) );
  AND U18284 ( .A(n17453), .B(n17452), .Z(n17670) );
  XNOR U18285 ( .A(n17669), .B(n17670), .Z(n17671) );
  XOR U18286 ( .A(n17672), .B(n17671), .Z(n17676) );
  XNOR U18287 ( .A(n17675), .B(n17676), .Z(n17677) );
  NANDN U18288 ( .A(n17455), .B(n17454), .Z(n17459) );
  NAND U18289 ( .A(n17457), .B(n17456), .Z(n17458) );
  NAND U18290 ( .A(n17459), .B(n17458), .Z(n17678) );
  XOR U18291 ( .A(n17677), .B(n17678), .Z(n17782) );
  NANDN U18292 ( .A(n17461), .B(n17460), .Z(n17465) );
  NAND U18293 ( .A(n17463), .B(n17462), .Z(n17464) );
  NAND U18294 ( .A(n17465), .B(n17464), .Z(n17779) );
  NANDN U18295 ( .A(n17467), .B(n17466), .Z(n17471) );
  NAND U18296 ( .A(n17469), .B(n17468), .Z(n17470) );
  AND U18297 ( .A(n17471), .B(n17470), .Z(n17780) );
  XNOR U18298 ( .A(n17779), .B(n17780), .Z(n17781) );
  XNOR U18299 ( .A(n17782), .B(n17781), .Z(n17588) );
  OR U18300 ( .A(n17473), .B(n17472), .Z(n17477) );
  OR U18301 ( .A(n17475), .B(n17474), .Z(n17476) );
  AND U18302 ( .A(n17477), .B(n17476), .Z(n17589) );
  XNOR U18303 ( .A(n17588), .B(n17589), .Z(n17590) );
  NANDN U18304 ( .A(n17479), .B(n17478), .Z(n17483) );
  NAND U18305 ( .A(n17481), .B(n17480), .Z(n17482) );
  AND U18306 ( .A(n17483), .B(n17482), .Z(n17591) );
  XNOR U18307 ( .A(n17590), .B(n17591), .Z(n17595) );
  XNOR U18308 ( .A(a[79]), .B(b[11]), .Z(n17730) );
  OR U18309 ( .A(n17730), .B(n31369), .Z(n17486) );
  NANDN U18310 ( .A(n17484), .B(n31119), .Z(n17485) );
  NAND U18311 ( .A(n17486), .B(n17485), .Z(n17751) );
  XOR U18312 ( .A(b[43]), .B(n23149), .Z(n17733) );
  NANDN U18313 ( .A(n17733), .B(n37068), .Z(n17489) );
  NANDN U18314 ( .A(n17487), .B(n37069), .Z(n17488) );
  NAND U18315 ( .A(n17489), .B(n17488), .Z(n17748) );
  XNOR U18316 ( .A(b[45]), .B(a[45]), .Z(n17736) );
  NANDN U18317 ( .A(n17736), .B(n37261), .Z(n17492) );
  NANDN U18318 ( .A(n17490), .B(n37262), .Z(n17491) );
  AND U18319 ( .A(n17492), .B(n17491), .Z(n17749) );
  XNOR U18320 ( .A(n17748), .B(n17749), .Z(n17750) );
  XNOR U18321 ( .A(n17751), .B(n17750), .Z(n17624) );
  XOR U18322 ( .A(b[49]), .B(n21441), .Z(n17739) );
  OR U18323 ( .A(n17739), .B(n37756), .Z(n17495) );
  NANDN U18324 ( .A(n17493), .B(n37652), .Z(n17494) );
  NAND U18325 ( .A(n17495), .B(n17494), .Z(n17772) );
  NAND U18326 ( .A(n17496), .B(n37469), .Z(n17498) );
  XOR U18327 ( .A(n978), .B(n21996), .Z(n17742) );
  NAND U18328 ( .A(n17742), .B(n37471), .Z(n17497) );
  NAND U18329 ( .A(n17498), .B(n17497), .Z(n17769) );
  XNOR U18330 ( .A(a[81]), .B(b[9]), .Z(n17745) );
  NANDN U18331 ( .A(n17745), .B(n30509), .Z(n17501) );
  NAND U18332 ( .A(n17499), .B(n30846), .Z(n17500) );
  AND U18333 ( .A(n17501), .B(n17500), .Z(n17770) );
  XNOR U18334 ( .A(n17769), .B(n17770), .Z(n17771) );
  XOR U18335 ( .A(n17772), .B(n17771), .Z(n17625) );
  XNOR U18336 ( .A(n17624), .B(n17625), .Z(n17626) );
  NANDN U18337 ( .A(n17503), .B(n17502), .Z(n17507) );
  NAND U18338 ( .A(n17505), .B(n17504), .Z(n17506) );
  AND U18339 ( .A(n17507), .B(n17506), .Z(n17627) );
  XNOR U18340 ( .A(n17626), .B(n17627), .Z(n17579) );
  XNOR U18341 ( .A(n17579), .B(n17578), .Z(n17580) );
  XNOR U18342 ( .A(b[35]), .B(a[55]), .Z(n17754) );
  NANDN U18343 ( .A(n17754), .B(n35985), .Z(n17514) );
  NANDN U18344 ( .A(n17512), .B(n35986), .Z(n17513) );
  NAND U18345 ( .A(n17514), .B(n17513), .Z(n17818) );
  XNOR U18346 ( .A(a[83]), .B(n31123), .Z(n17757) );
  NAND U18347 ( .A(n17757), .B(n29949), .Z(n17517) );
  NAND U18348 ( .A(n29948), .B(n17515), .Z(n17516) );
  NAND U18349 ( .A(n17517), .B(n17516), .Z(n17815) );
  XOR U18350 ( .A(b[55]), .B(n20315), .Z(n17760) );
  NANDN U18351 ( .A(n17760), .B(n38075), .Z(n17520) );
  NANDN U18352 ( .A(n17518), .B(n38073), .Z(n17519) );
  AND U18353 ( .A(n17520), .B(n17519), .Z(n17816) );
  XNOR U18354 ( .A(n17815), .B(n17816), .Z(n17817) );
  XNOR U18355 ( .A(n17818), .B(n17817), .Z(n17609) );
  NANDN U18356 ( .A(n17522), .B(n17521), .Z(n17526) );
  NAND U18357 ( .A(n17524), .B(n17523), .Z(n17525) );
  NAND U18358 ( .A(n17526), .B(n17525), .Z(n17606) );
  XNOR U18359 ( .A(n17606), .B(n17607), .Z(n17608) );
  XOR U18360 ( .A(n17609), .B(n17608), .Z(n17581) );
  XOR U18361 ( .A(n17580), .B(n17581), .Z(n17594) );
  XOR U18362 ( .A(n17595), .B(n17594), .Z(n17597) );
  XNOR U18363 ( .A(n17596), .B(n17597), .Z(n17828) );
  XNOR U18364 ( .A(n17827), .B(n17828), .Z(n17829) );
  NAND U18365 ( .A(n17532), .B(n17531), .Z(n17536) );
  NANDN U18366 ( .A(n17534), .B(n17533), .Z(n17535) );
  AND U18367 ( .A(n17536), .B(n17535), .Z(n17830) );
  XNOR U18368 ( .A(n17829), .B(n17830), .Z(n17840) );
  XOR U18369 ( .A(n17839), .B(n17840), .Z(n17846) );
  NANDN U18370 ( .A(n17538), .B(n17537), .Z(n17542) );
  NANDN U18371 ( .A(n17540), .B(n17539), .Z(n17541) );
  NAND U18372 ( .A(n17542), .B(n17541), .Z(n17844) );
  NANDN U18373 ( .A(n17544), .B(n17543), .Z(n17548) );
  NANDN U18374 ( .A(n17546), .B(n17545), .Z(n17547) );
  AND U18375 ( .A(n17548), .B(n17547), .Z(n17843) );
  XNOR U18376 ( .A(n17844), .B(n17843), .Z(n17845) );
  XNOR U18377 ( .A(n17846), .B(n17845), .Z(n17852) );
  OR U18378 ( .A(n17550), .B(n17549), .Z(n17554) );
  NANDN U18379 ( .A(n17552), .B(n17551), .Z(n17553) );
  NAND U18380 ( .A(n17554), .B(n17553), .Z(n17850) );
  NANDN U18381 ( .A(n17556), .B(n17555), .Z(n17560) );
  NANDN U18382 ( .A(n17558), .B(n17557), .Z(n17559) );
  AND U18383 ( .A(n17560), .B(n17559), .Z(n17849) );
  XNOR U18384 ( .A(n17850), .B(n17849), .Z(n17851) );
  XOR U18385 ( .A(n17852), .B(n17851), .Z(n17573) );
  NANDN U18386 ( .A(n17562), .B(n17561), .Z(n17566) );
  NAND U18387 ( .A(n17564), .B(n17563), .Z(n17565) );
  AND U18388 ( .A(n17566), .B(n17565), .Z(n17572) );
  XOR U18389 ( .A(n17573), .B(n17572), .Z(n17574) );
  XNOR U18390 ( .A(n17575), .B(n17574), .Z(n17855) );
  XNOR U18391 ( .A(n17855), .B(sreg[153]), .Z(n17857) );
  NAND U18392 ( .A(n17567), .B(sreg[152]), .Z(n17571) );
  OR U18393 ( .A(n17569), .B(n17568), .Z(n17570) );
  AND U18394 ( .A(n17571), .B(n17570), .Z(n17856) );
  XOR U18395 ( .A(n17857), .B(n17856), .Z(c[153]) );
  OR U18396 ( .A(n17573), .B(n17572), .Z(n17577) );
  NAND U18397 ( .A(n17575), .B(n17574), .Z(n17576) );
  NAND U18398 ( .A(n17577), .B(n17576), .Z(n17863) );
  NANDN U18399 ( .A(n17579), .B(n17578), .Z(n17583) );
  NAND U18400 ( .A(n17581), .B(n17580), .Z(n17582) );
  NAND U18401 ( .A(n17583), .B(n17582), .Z(n18131) );
  NANDN U18402 ( .A(n17589), .B(n17588), .Z(n17593) );
  NAND U18403 ( .A(n17591), .B(n17590), .Z(n17592) );
  AND U18404 ( .A(n17593), .B(n17592), .Z(n18129) );
  XNOR U18405 ( .A(n18128), .B(n18129), .Z(n18130) );
  XNOR U18406 ( .A(n18131), .B(n18130), .Z(n17876) );
  NANDN U18407 ( .A(n17595), .B(n17594), .Z(n17599) );
  NANDN U18408 ( .A(n17597), .B(n17596), .Z(n17598) );
  NAND U18409 ( .A(n17599), .B(n17598), .Z(n17877) );
  XOR U18410 ( .A(n17876), .B(n17877), .Z(n17879) );
  NANDN U18411 ( .A(n17601), .B(n17600), .Z(n17605) );
  OR U18412 ( .A(n17603), .B(n17602), .Z(n17604) );
  NAND U18413 ( .A(n17605), .B(n17604), .Z(n18122) );
  NANDN U18414 ( .A(n17607), .B(n17606), .Z(n17611) );
  NAND U18415 ( .A(n17609), .B(n17608), .Z(n17610) );
  NAND U18416 ( .A(n17611), .B(n17610), .Z(n17896) );
  NAND U18417 ( .A(n17613), .B(n17612), .Z(n17617) );
  NANDN U18418 ( .A(n17615), .B(n17614), .Z(n17616) );
  NAND U18419 ( .A(n17617), .B(n17616), .Z(n17894) );
  NANDN U18420 ( .A(n17619), .B(n17618), .Z(n17623) );
  OR U18421 ( .A(n17621), .B(n17620), .Z(n17622) );
  AND U18422 ( .A(n17623), .B(n17622), .Z(n17895) );
  XNOR U18423 ( .A(n17894), .B(n17895), .Z(n17897) );
  XNOR U18424 ( .A(n17896), .B(n17897), .Z(n18123) );
  XOR U18425 ( .A(n18122), .B(n18123), .Z(n18124) );
  NANDN U18426 ( .A(n17625), .B(n17624), .Z(n17629) );
  NAND U18427 ( .A(n17627), .B(n17626), .Z(n17628) );
  NAND U18428 ( .A(n17629), .B(n17628), .Z(n17922) );
  NAND U18429 ( .A(n33283), .B(n17630), .Z(n17632) );
  XOR U18430 ( .A(n33020), .B(n30210), .Z(n17967) );
  NANDN U18431 ( .A(n33021), .B(n17967), .Z(n17631) );
  NAND U18432 ( .A(n17632), .B(n17631), .Z(n18010) );
  XNOR U18433 ( .A(b[21]), .B(a[70]), .Z(n17970) );
  OR U18434 ( .A(n17970), .B(n33634), .Z(n17635) );
  NAND U18435 ( .A(n17633), .B(n33464), .Z(n17634) );
  NAND U18436 ( .A(n17635), .B(n17634), .Z(n18007) );
  NAND U18437 ( .A(n34044), .B(n17636), .Z(n17638) );
  XOR U18438 ( .A(n34510), .B(n29868), .Z(n17973) );
  NANDN U18439 ( .A(n33867), .B(n17973), .Z(n17637) );
  AND U18440 ( .A(n17638), .B(n17637), .Z(n18008) );
  XNOR U18441 ( .A(n18007), .B(n18008), .Z(n18009) );
  XOR U18442 ( .A(n18010), .B(n18009), .Z(n18086) );
  NANDN U18443 ( .A(n17640), .B(n17639), .Z(n17644) );
  NAND U18444 ( .A(n17642), .B(n17641), .Z(n17643) );
  NAND U18445 ( .A(n17644), .B(n17643), .Z(n18087) );
  XNOR U18446 ( .A(n18086), .B(n18087), .Z(n18089) );
  NAND U18447 ( .A(a[26]), .B(b[63]), .Z(n18077) );
  NANDN U18448 ( .A(n17645), .B(n38369), .Z(n17647) );
  XOR U18449 ( .A(b[61]), .B(n18804), .Z(n17961) );
  OR U18450 ( .A(n17961), .B(n38371), .Z(n17646) );
  NAND U18451 ( .A(n17647), .B(n17646), .Z(n18075) );
  NANDN U18452 ( .A(n17648), .B(n35311), .Z(n17650) );
  XOR U18453 ( .A(b[31]), .B(n27436), .Z(n17964) );
  NANDN U18454 ( .A(n17964), .B(n35313), .Z(n17649) );
  AND U18455 ( .A(n17650), .B(n17649), .Z(n18074) );
  XNOR U18456 ( .A(n18075), .B(n18074), .Z(n18076) );
  XNOR U18457 ( .A(n18077), .B(n18076), .Z(n18088) );
  XNOR U18458 ( .A(n18089), .B(n18088), .Z(n17920) );
  XOR U18459 ( .A(b[37]), .B(n25177), .Z(n17930) );
  NANDN U18460 ( .A(n17930), .B(n36311), .Z(n17653) );
  NANDN U18461 ( .A(n17651), .B(n36309), .Z(n17652) );
  NAND U18462 ( .A(n17653), .B(n17652), .Z(n17985) );
  XOR U18463 ( .A(a[86]), .B(n968), .Z(n17933) );
  OR U18464 ( .A(n17933), .B(n29363), .Z(n17656) );
  NANDN U18465 ( .A(n17654), .B(n29864), .Z(n17655) );
  NAND U18466 ( .A(n17656), .B(n17655), .Z(n17982) );
  XOR U18467 ( .A(n34048), .B(n967), .Z(n17936) );
  NAND U18468 ( .A(n17936), .B(n28939), .Z(n17659) );
  NAND U18469 ( .A(n28938), .B(n17657), .Z(n17658) );
  AND U18470 ( .A(n17659), .B(n17658), .Z(n17983) );
  XNOR U18471 ( .A(n17982), .B(n17983), .Z(n17984) );
  XNOR U18472 ( .A(n17985), .B(n17984), .Z(n17917) );
  XOR U18473 ( .A(b[13]), .B(n31870), .Z(n17939) );
  OR U18474 ( .A(n17939), .B(n31550), .Z(n17662) );
  NANDN U18475 ( .A(n17660), .B(n31874), .Z(n17661) );
  NAND U18476 ( .A(n17662), .B(n17661), .Z(n18056) );
  NAND U18477 ( .A(n34848), .B(n17663), .Z(n17665) );
  XNOR U18478 ( .A(n35375), .B(a[64]), .Z(n17942) );
  NAND U18479 ( .A(n34618), .B(n17942), .Z(n17664) );
  NAND U18480 ( .A(n17665), .B(n17664), .Z(n18053) );
  NAND U18481 ( .A(n35188), .B(n17666), .Z(n17668) );
  XNOR U18482 ( .A(n35540), .B(a[62]), .Z(n17945) );
  NANDN U18483 ( .A(n34968), .B(n17945), .Z(n17667) );
  AND U18484 ( .A(n17668), .B(n17667), .Z(n18054) );
  XNOR U18485 ( .A(n18053), .B(n18054), .Z(n18055) );
  XNOR U18486 ( .A(n18056), .B(n18055), .Z(n17914) );
  NANDN U18487 ( .A(n17670), .B(n17669), .Z(n17674) );
  NAND U18488 ( .A(n17672), .B(n17671), .Z(n17673) );
  NAND U18489 ( .A(n17674), .B(n17673), .Z(n17915) );
  XNOR U18490 ( .A(n17914), .B(n17915), .Z(n17916) );
  XOR U18491 ( .A(n17917), .B(n17916), .Z(n17921) );
  XOR U18492 ( .A(n17920), .B(n17921), .Z(n17923) );
  XNOR U18493 ( .A(n17922), .B(n17923), .Z(n18118) );
  NANDN U18494 ( .A(n17676), .B(n17675), .Z(n17680) );
  NANDN U18495 ( .A(n17678), .B(n17677), .Z(n17679) );
  NAND U18496 ( .A(n17680), .B(n17679), .Z(n18117) );
  NANDN U18497 ( .A(n17682), .B(n17681), .Z(n17686) );
  NAND U18498 ( .A(n17684), .B(n17683), .Z(n17685) );
  NAND U18499 ( .A(n17686), .B(n17685), .Z(n17911) );
  XNOR U18500 ( .A(b[41]), .B(a[50]), .Z(n17988) );
  OR U18501 ( .A(n17988), .B(n36905), .Z(n17689) );
  NANDN U18502 ( .A(n17687), .B(n36807), .Z(n17688) );
  NAND U18503 ( .A(n17689), .B(n17688), .Z(n18016) );
  XOR U18504 ( .A(b[57]), .B(n19513), .Z(n17991) );
  OR U18505 ( .A(n17991), .B(n965), .Z(n17692) );
  NANDN U18506 ( .A(n17690), .B(n38194), .Z(n17691) );
  NAND U18507 ( .A(n17692), .B(n17691), .Z(n18013) );
  NAND U18508 ( .A(n38326), .B(n17693), .Z(n17695) );
  XOR U18509 ( .A(n38400), .B(n18841), .Z(n17994) );
  NANDN U18510 ( .A(n38273), .B(n17994), .Z(n17694) );
  AND U18511 ( .A(n17695), .B(n17694), .Z(n18014) );
  XNOR U18512 ( .A(n18013), .B(n18014), .Z(n18015) );
  XOR U18513 ( .A(n18016), .B(n18015), .Z(n18025) );
  XOR U18514 ( .A(b[33]), .B(n26347), .Z(n17997) );
  NANDN U18515 ( .A(n17997), .B(n35620), .Z(n17698) );
  NANDN U18516 ( .A(n17696), .B(n35621), .Z(n17697) );
  NAND U18517 ( .A(n17698), .B(n17697), .Z(n18032) );
  NANDN U18518 ( .A(n966), .B(a[90]), .Z(n17699) );
  XOR U18519 ( .A(n29232), .B(n17699), .Z(n17701) );
  NANDN U18520 ( .A(b[0]), .B(a[89]), .Z(n17700) );
  AND U18521 ( .A(n17701), .B(n17700), .Z(n18029) );
  XOR U18522 ( .A(b[63]), .B(n17702), .Z(n18004) );
  NANDN U18523 ( .A(n18004), .B(n38422), .Z(n17705) );
  NANDN U18524 ( .A(n17703), .B(n38423), .Z(n17704) );
  AND U18525 ( .A(n17705), .B(n17704), .Z(n18030) );
  XNOR U18526 ( .A(n18029), .B(n18030), .Z(n18031) );
  XOR U18527 ( .A(n18032), .B(n18031), .Z(n18026) );
  XNOR U18528 ( .A(n18025), .B(n18026), .Z(n18028) );
  NANDN U18529 ( .A(n17707), .B(n17706), .Z(n17711) );
  NAND U18530 ( .A(n17709), .B(n17708), .Z(n17710) );
  AND U18531 ( .A(n17711), .B(n17710), .Z(n18027) );
  XNOR U18532 ( .A(n18028), .B(n18027), .Z(n17908) );
  NANDN U18533 ( .A(n17713), .B(n17712), .Z(n17717) );
  NAND U18534 ( .A(n17715), .B(n17714), .Z(n17716) );
  AND U18535 ( .A(n17717), .B(n17716), .Z(n17909) );
  XOR U18536 ( .A(n17908), .B(n17909), .Z(n17910) );
  XNOR U18537 ( .A(n17911), .B(n17910), .Z(n18116) );
  XNOR U18538 ( .A(n18117), .B(n18116), .Z(n18119) );
  XNOR U18539 ( .A(n18118), .B(n18119), .Z(n18125) );
  XNOR U18540 ( .A(n18124), .B(n18125), .Z(n18135) );
  NAND U18541 ( .A(n17719), .B(n17718), .Z(n17723) );
  NANDN U18542 ( .A(n17721), .B(n17720), .Z(n17722) );
  NAND U18543 ( .A(n17723), .B(n17722), .Z(n17900) );
  OR U18544 ( .A(n17725), .B(n17724), .Z(n17729) );
  OR U18545 ( .A(n17727), .B(n17726), .Z(n17728) );
  NAND U18546 ( .A(n17729), .B(n17728), .Z(n17883) );
  XOR U18547 ( .A(a[80]), .B(n970), .Z(n18092) );
  OR U18548 ( .A(n18092), .B(n31369), .Z(n17732) );
  NANDN U18549 ( .A(n17730), .B(n31119), .Z(n17731) );
  NAND U18550 ( .A(n17732), .B(n17731), .Z(n18113) );
  XOR U18551 ( .A(b[43]), .B(n23447), .Z(n18095) );
  NANDN U18552 ( .A(n18095), .B(n37068), .Z(n17735) );
  NANDN U18553 ( .A(n17733), .B(n37069), .Z(n17734) );
  NAND U18554 ( .A(n17735), .B(n17734), .Z(n18110) );
  XNOR U18555 ( .A(b[45]), .B(a[46]), .Z(n18098) );
  NANDN U18556 ( .A(n18098), .B(n37261), .Z(n17738) );
  NANDN U18557 ( .A(n17736), .B(n37262), .Z(n17737) );
  AND U18558 ( .A(n17738), .B(n17737), .Z(n18111) );
  XNOR U18559 ( .A(n18110), .B(n18111), .Z(n18112) );
  XNOR U18560 ( .A(n18113), .B(n18112), .Z(n17929) );
  XOR U18561 ( .A(b[49]), .B(n22246), .Z(n18101) );
  OR U18562 ( .A(n18101), .B(n37756), .Z(n17741) );
  NANDN U18563 ( .A(n17739), .B(n37652), .Z(n17740) );
  NAND U18564 ( .A(n17741), .B(n17740), .Z(n18083) );
  NAND U18565 ( .A(n37469), .B(n17742), .Z(n17744) );
  XOR U18566 ( .A(n978), .B(n22289), .Z(n18104) );
  NAND U18567 ( .A(n18104), .B(n37471), .Z(n17743) );
  NAND U18568 ( .A(n17744), .B(n17743), .Z(n18080) );
  XOR U18569 ( .A(a[82]), .B(n969), .Z(n18107) );
  NANDN U18570 ( .A(n18107), .B(n30509), .Z(n17747) );
  NANDN U18571 ( .A(n17745), .B(n30846), .Z(n17746) );
  AND U18572 ( .A(n17747), .B(n17746), .Z(n18081) );
  XNOR U18573 ( .A(n18080), .B(n18081), .Z(n18082) );
  XNOR U18574 ( .A(n18083), .B(n18082), .Z(n17926) );
  NANDN U18575 ( .A(n17749), .B(n17748), .Z(n17753) );
  NAND U18576 ( .A(n17751), .B(n17750), .Z(n17752) );
  NAND U18577 ( .A(n17753), .B(n17752), .Z(n17927) );
  XNOR U18578 ( .A(n17926), .B(n17927), .Z(n17928) );
  XOR U18579 ( .A(n17929), .B(n17928), .Z(n17882) );
  XNOR U18580 ( .A(n17883), .B(n17882), .Z(n17885) );
  XNOR U18581 ( .A(b[35]), .B(a[56]), .Z(n18065) );
  NANDN U18582 ( .A(n18065), .B(n35985), .Z(n17756) );
  NANDN U18583 ( .A(n17754), .B(n35986), .Z(n17755) );
  NAND U18584 ( .A(n17756), .B(n17755), .Z(n18062) );
  XOR U18585 ( .A(n33185), .B(n31123), .Z(n18068) );
  NAND U18586 ( .A(n18068), .B(n29949), .Z(n17759) );
  NAND U18587 ( .A(n29948), .B(n17757), .Z(n17758) );
  NAND U18588 ( .A(n17759), .B(n17758), .Z(n18059) );
  XOR U18589 ( .A(b[55]), .B(n19980), .Z(n18071) );
  NANDN U18590 ( .A(n18071), .B(n38075), .Z(n17762) );
  NANDN U18591 ( .A(n17760), .B(n38073), .Z(n17761) );
  AND U18592 ( .A(n17762), .B(n17761), .Z(n18060) );
  XNOR U18593 ( .A(n18059), .B(n18060), .Z(n18061) );
  XNOR U18594 ( .A(n18062), .B(n18061), .Z(n17905) );
  NANDN U18595 ( .A(n17764), .B(n17763), .Z(n17768) );
  NAND U18596 ( .A(n17766), .B(n17765), .Z(n17767) );
  NAND U18597 ( .A(n17768), .B(n17767), .Z(n17902) );
  NANDN U18598 ( .A(n17770), .B(n17769), .Z(n17774) );
  NAND U18599 ( .A(n17772), .B(n17771), .Z(n17773) );
  NAND U18600 ( .A(n17774), .B(n17773), .Z(n17903) );
  XNOR U18601 ( .A(n17902), .B(n17903), .Z(n17904) );
  XOR U18602 ( .A(n17905), .B(n17904), .Z(n17884) );
  XNOR U18603 ( .A(n17885), .B(n17884), .Z(n17899) );
  NANDN U18604 ( .A(n17780), .B(n17779), .Z(n17784) );
  NAND U18605 ( .A(n17782), .B(n17781), .Z(n17783) );
  NAND U18606 ( .A(n17784), .B(n17783), .Z(n17889) );
  XNOR U18607 ( .A(n17888), .B(n17889), .Z(n17890) );
  NANDN U18608 ( .A(n17786), .B(n17785), .Z(n17790) );
  NAND U18609 ( .A(n17788), .B(n17787), .Z(n17789) );
  NAND U18610 ( .A(n17790), .B(n17789), .Z(n18022) );
  XOR U18611 ( .A(b[15]), .B(n31363), .Z(n18035) );
  OR U18612 ( .A(n18035), .B(n32010), .Z(n17793) );
  NANDN U18613 ( .A(n17791), .B(n32011), .Z(n17792) );
  NAND U18614 ( .A(n17793), .B(n17792), .Z(n17957) );
  XNOR U18615 ( .A(b[25]), .B(n28701), .Z(n18038) );
  NANDN U18616 ( .A(n34219), .B(n18038), .Z(n17796) );
  NAND U18617 ( .A(n34217), .B(n17794), .Z(n17795) );
  NAND U18618 ( .A(n17796), .B(n17795), .Z(n17954) );
  XNOR U18619 ( .A(b[17]), .B(a[74]), .Z(n18041) );
  NANDN U18620 ( .A(n18041), .B(n32543), .Z(n17799) );
  NAND U18621 ( .A(n17797), .B(n32541), .Z(n17798) );
  AND U18622 ( .A(n17799), .B(n17798), .Z(n17955) );
  XNOR U18623 ( .A(n17954), .B(n17955), .Z(n17956) );
  XNOR U18624 ( .A(n17957), .B(n17956), .Z(n17978) );
  XOR U18625 ( .A(b[39]), .B(n25134), .Z(n18044) );
  NANDN U18626 ( .A(n18044), .B(n36553), .Z(n17802) );
  NANDN U18627 ( .A(n17800), .B(n36643), .Z(n17801) );
  NAND U18628 ( .A(n17802), .B(n17801), .Z(n17951) );
  XOR U18629 ( .A(b[51]), .B(n21149), .Z(n18047) );
  NANDN U18630 ( .A(n18047), .B(n37803), .Z(n17805) );
  NANDN U18631 ( .A(n17803), .B(n37802), .Z(n17804) );
  NAND U18632 ( .A(n17805), .B(n17804), .Z(n17948) );
  XOR U18633 ( .A(b[53]), .B(n20686), .Z(n18050) );
  NANDN U18634 ( .A(n18050), .B(n37940), .Z(n17808) );
  NANDN U18635 ( .A(n17806), .B(n37941), .Z(n17807) );
  AND U18636 ( .A(n17808), .B(n17807), .Z(n17949) );
  XNOR U18637 ( .A(n17948), .B(n17949), .Z(n17950) );
  XNOR U18638 ( .A(n17951), .B(n17950), .Z(n17976) );
  NANDN U18639 ( .A(n17810), .B(n17809), .Z(n17814) );
  NAND U18640 ( .A(n17812), .B(n17811), .Z(n17813) );
  NAND U18641 ( .A(n17814), .B(n17813), .Z(n17977) );
  XOR U18642 ( .A(n17976), .B(n17977), .Z(n17979) );
  XNOR U18643 ( .A(n17978), .B(n17979), .Z(n18019) );
  NANDN U18644 ( .A(n17816), .B(n17815), .Z(n17820) );
  NAND U18645 ( .A(n17818), .B(n17817), .Z(n17819) );
  AND U18646 ( .A(n17820), .B(n17819), .Z(n18020) );
  XOR U18647 ( .A(n18019), .B(n18020), .Z(n18021) );
  XOR U18648 ( .A(n18022), .B(n18021), .Z(n17891) );
  XNOR U18649 ( .A(n17890), .B(n17891), .Z(n17898) );
  XOR U18650 ( .A(n17899), .B(n17898), .Z(n17901) );
  XNOR U18651 ( .A(n17900), .B(n17901), .Z(n18134) );
  XNOR U18652 ( .A(n18135), .B(n18134), .Z(n18137) );
  OR U18653 ( .A(n17822), .B(n17821), .Z(n17826) );
  NAND U18654 ( .A(n17824), .B(n17823), .Z(n17825) );
  AND U18655 ( .A(n17826), .B(n17825), .Z(n18136) );
  XNOR U18656 ( .A(n18137), .B(n18136), .Z(n17878) );
  XOR U18657 ( .A(n17879), .B(n17878), .Z(n17874) );
  NANDN U18658 ( .A(n17832), .B(n17831), .Z(n17836) );
  NANDN U18659 ( .A(n17834), .B(n17833), .Z(n17835) );
  AND U18660 ( .A(n17836), .B(n17835), .Z(n17872) );
  XNOR U18661 ( .A(n17873), .B(n17872), .Z(n17875) );
  XNOR U18662 ( .A(n17874), .B(n17875), .Z(n17866) );
  OR U18663 ( .A(n17838), .B(n17837), .Z(n17842) );
  NANDN U18664 ( .A(n17840), .B(n17839), .Z(n17841) );
  AND U18665 ( .A(n17842), .B(n17841), .Z(n17867) );
  XOR U18666 ( .A(n17866), .B(n17867), .Z(n17869) );
  NANDN U18667 ( .A(n17844), .B(n17843), .Z(n17848) );
  NAND U18668 ( .A(n17846), .B(n17845), .Z(n17847) );
  NAND U18669 ( .A(n17848), .B(n17847), .Z(n17868) );
  XNOR U18670 ( .A(n17869), .B(n17868), .Z(n17860) );
  NANDN U18671 ( .A(n17850), .B(n17849), .Z(n17854) );
  NAND U18672 ( .A(n17852), .B(n17851), .Z(n17853) );
  NAND U18673 ( .A(n17854), .B(n17853), .Z(n17861) );
  XNOR U18674 ( .A(n17860), .B(n17861), .Z(n17862) );
  XNOR U18675 ( .A(n17863), .B(n17862), .Z(n18140) );
  XNOR U18676 ( .A(n18140), .B(sreg[154]), .Z(n18142) );
  NAND U18677 ( .A(n17855), .B(sreg[153]), .Z(n17859) );
  OR U18678 ( .A(n17857), .B(n17856), .Z(n17858) );
  AND U18679 ( .A(n17859), .B(n17858), .Z(n18141) );
  XOR U18680 ( .A(n18142), .B(n18141), .Z(c[154]) );
  NANDN U18681 ( .A(n17861), .B(n17860), .Z(n17865) );
  NAND U18682 ( .A(n17863), .B(n17862), .Z(n17864) );
  NAND U18683 ( .A(n17865), .B(n17864), .Z(n18148) );
  NANDN U18684 ( .A(n17867), .B(n17866), .Z(n17871) );
  OR U18685 ( .A(n17869), .B(n17868), .Z(n17870) );
  NAND U18686 ( .A(n17871), .B(n17870), .Z(n18146) );
  NANDN U18687 ( .A(n17877), .B(n17876), .Z(n17881) );
  NANDN U18688 ( .A(n17879), .B(n17878), .Z(n17880) );
  NAND U18689 ( .A(n17881), .B(n17880), .Z(n18150) );
  XNOR U18690 ( .A(n18149), .B(n18150), .Z(n18151) );
  NAND U18691 ( .A(n17883), .B(n17882), .Z(n17887) );
  NANDN U18692 ( .A(n17885), .B(n17884), .Z(n17886) );
  NAND U18693 ( .A(n17887), .B(n17886), .Z(n18158) );
  NANDN U18694 ( .A(n17889), .B(n17888), .Z(n17893) );
  NANDN U18695 ( .A(n17891), .B(n17890), .Z(n17892) );
  NAND U18696 ( .A(n17893), .B(n17892), .Z(n18155) );
  XNOR U18697 ( .A(n18155), .B(n18156), .Z(n18157) );
  XOR U18698 ( .A(n18158), .B(n18157), .Z(n18415) );
  XNOR U18699 ( .A(n18415), .B(n18416), .Z(n18418) );
  NANDN U18700 ( .A(n17903), .B(n17902), .Z(n17907) );
  NAND U18701 ( .A(n17905), .B(n17904), .Z(n17906) );
  AND U18702 ( .A(n17907), .B(n17906), .Z(n18402) );
  NAND U18703 ( .A(n17909), .B(n17908), .Z(n17913) );
  NANDN U18704 ( .A(n17911), .B(n17910), .Z(n17912) );
  NAND U18705 ( .A(n17913), .B(n17912), .Z(n18399) );
  NANDN U18706 ( .A(n17915), .B(n17914), .Z(n17919) );
  NAND U18707 ( .A(n17917), .B(n17916), .Z(n17918) );
  AND U18708 ( .A(n17919), .B(n17918), .Z(n18400) );
  XNOR U18709 ( .A(n18399), .B(n18400), .Z(n18401) );
  XNOR U18710 ( .A(n18402), .B(n18401), .Z(n18387) );
  NANDN U18711 ( .A(n17921), .B(n17920), .Z(n17925) );
  OR U18712 ( .A(n17923), .B(n17922), .Z(n17924) );
  AND U18713 ( .A(n17925), .B(n17924), .Z(n18388) );
  XNOR U18714 ( .A(n18387), .B(n18388), .Z(n18390) );
  XOR U18715 ( .A(b[37]), .B(n25466), .Z(n18195) );
  NANDN U18716 ( .A(n18195), .B(n36311), .Z(n17932) );
  NANDN U18717 ( .A(n17930), .B(n36309), .Z(n17931) );
  NAND U18718 ( .A(n17932), .B(n17931), .Z(n18273) );
  XNOR U18719 ( .A(a[87]), .B(b[5]), .Z(n18198) );
  OR U18720 ( .A(n18198), .B(n29363), .Z(n17935) );
  NANDN U18721 ( .A(n17933), .B(n29864), .Z(n17934) );
  NAND U18722 ( .A(n17935), .B(n17934), .Z(n18270) );
  XNOR U18723 ( .A(a[89]), .B(n967), .Z(n18201) );
  NAND U18724 ( .A(n18201), .B(n28939), .Z(n17938) );
  NAND U18725 ( .A(n28938), .B(n17936), .Z(n17937) );
  AND U18726 ( .A(n17938), .B(n17937), .Z(n18271) );
  XNOR U18727 ( .A(n18270), .B(n18271), .Z(n18272) );
  XNOR U18728 ( .A(n18273), .B(n18272), .Z(n18182) );
  XNOR U18729 ( .A(b[13]), .B(a[79]), .Z(n18204) );
  OR U18730 ( .A(n18204), .B(n31550), .Z(n17941) );
  NANDN U18731 ( .A(n17939), .B(n31874), .Z(n17940) );
  NAND U18732 ( .A(n17941), .B(n17940), .Z(n18378) );
  NAND U18733 ( .A(n34848), .B(n17942), .Z(n17944) );
  XOR U18734 ( .A(n35375), .B(n28403), .Z(n18207) );
  NAND U18735 ( .A(n34618), .B(n18207), .Z(n17943) );
  NAND U18736 ( .A(n17944), .B(n17943), .Z(n18375) );
  NAND U18737 ( .A(n35188), .B(n17945), .Z(n17947) );
  XNOR U18738 ( .A(n35540), .B(a[63]), .Z(n18210) );
  NANDN U18739 ( .A(n34968), .B(n18210), .Z(n17946) );
  AND U18740 ( .A(n17947), .B(n17946), .Z(n18376) );
  XNOR U18741 ( .A(n18375), .B(n18376), .Z(n18377) );
  XNOR U18742 ( .A(n18378), .B(n18377), .Z(n18179) );
  NANDN U18743 ( .A(n17949), .B(n17948), .Z(n17953) );
  NAND U18744 ( .A(n17951), .B(n17950), .Z(n17952) );
  NAND U18745 ( .A(n17953), .B(n17952), .Z(n18180) );
  XNOR U18746 ( .A(n18179), .B(n18180), .Z(n18181) );
  XOR U18747 ( .A(n18182), .B(n18181), .Z(n18185) );
  NANDN U18748 ( .A(n17955), .B(n17954), .Z(n17959) );
  NAND U18749 ( .A(n17957), .B(n17956), .Z(n17958) );
  NAND U18750 ( .A(n17959), .B(n17958), .Z(n18336) );
  ANDN U18751 ( .B(b[63]), .A(n17960), .Z(n18300) );
  NANDN U18752 ( .A(n17961), .B(n38369), .Z(n17963) );
  XOR U18753 ( .A(b[61]), .B(n18639), .Z(n18225) );
  OR U18754 ( .A(n18225), .B(n38371), .Z(n17962) );
  NAND U18755 ( .A(n17963), .B(n17962), .Z(n18298) );
  NANDN U18756 ( .A(n17964), .B(n35311), .Z(n17966) );
  XOR U18757 ( .A(b[31]), .B(n27773), .Z(n18228) );
  NANDN U18758 ( .A(n18228), .B(n35313), .Z(n17965) );
  AND U18759 ( .A(n17966), .B(n17965), .Z(n18297) );
  XNOR U18760 ( .A(n18298), .B(n18297), .Z(n18299) );
  XOR U18761 ( .A(n18300), .B(n18299), .Z(n18333) );
  NAND U18762 ( .A(n33283), .B(n17967), .Z(n17969) );
  XNOR U18763 ( .A(n33020), .B(a[73]), .Z(n18231) );
  NANDN U18764 ( .A(n33021), .B(n18231), .Z(n17968) );
  NAND U18765 ( .A(n17969), .B(n17968), .Z(n18261) );
  XNOR U18766 ( .A(b[21]), .B(a[71]), .Z(n18234) );
  OR U18767 ( .A(n18234), .B(n33634), .Z(n17972) );
  NANDN U18768 ( .A(n17970), .B(n33464), .Z(n17971) );
  NAND U18769 ( .A(n17972), .B(n17971), .Z(n18258) );
  NAND U18770 ( .A(n34044), .B(n17973), .Z(n17975) );
  XNOR U18771 ( .A(n34510), .B(a[69]), .Z(n18237) );
  NANDN U18772 ( .A(n33867), .B(n18237), .Z(n17974) );
  AND U18773 ( .A(n17975), .B(n17974), .Z(n18259) );
  XNOR U18774 ( .A(n18258), .B(n18259), .Z(n18260) );
  XNOR U18775 ( .A(n18261), .B(n18260), .Z(n18334) );
  XNOR U18776 ( .A(n18333), .B(n18334), .Z(n18335) );
  XNOR U18777 ( .A(n18336), .B(n18335), .Z(n18186) );
  XOR U18778 ( .A(n18185), .B(n18186), .Z(n18187) );
  XOR U18779 ( .A(n18188), .B(n18187), .Z(n18284) );
  NANDN U18780 ( .A(n17977), .B(n17976), .Z(n17981) );
  NANDN U18781 ( .A(n17979), .B(n17978), .Z(n17980) );
  NAND U18782 ( .A(n17981), .B(n17980), .Z(n18283) );
  NANDN U18783 ( .A(n17983), .B(n17982), .Z(n17987) );
  NAND U18784 ( .A(n17985), .B(n17984), .Z(n17986) );
  NAND U18785 ( .A(n17987), .B(n17986), .Z(n18176) );
  XNOR U18786 ( .A(b[41]), .B(a[51]), .Z(n18249) );
  OR U18787 ( .A(n18249), .B(n36905), .Z(n17990) );
  NANDN U18788 ( .A(n17988), .B(n36807), .Z(n17989) );
  NAND U18789 ( .A(n17990), .B(n17989), .Z(n18267) );
  XOR U18790 ( .A(b[57]), .B(n20315), .Z(n18252) );
  OR U18791 ( .A(n18252), .B(n965), .Z(n17993) );
  NANDN U18792 ( .A(n17991), .B(n38194), .Z(n17992) );
  NAND U18793 ( .A(n17993), .B(n17992), .Z(n18264) );
  NAND U18794 ( .A(n38326), .B(n17994), .Z(n17996) );
  XOR U18795 ( .A(n38400), .B(n19656), .Z(n18255) );
  NANDN U18796 ( .A(n38273), .B(n18255), .Z(n17995) );
  AND U18797 ( .A(n17996), .B(n17995), .Z(n18265) );
  XNOR U18798 ( .A(n18264), .B(n18265), .Z(n18266) );
  XNOR U18799 ( .A(n18267), .B(n18266), .Z(n18345) );
  XNOR U18800 ( .A(b[33]), .B(a[59]), .Z(n18240) );
  NANDN U18801 ( .A(n18240), .B(n35620), .Z(n17999) );
  NANDN U18802 ( .A(n17997), .B(n35621), .Z(n17998) );
  NAND U18803 ( .A(n17999), .B(n17998), .Z(n18354) );
  NANDN U18804 ( .A(n966), .B(a[91]), .Z(n18000) );
  XOR U18805 ( .A(n29232), .B(n18000), .Z(n18002) );
  IV U18806 ( .A(a[90]), .Z(n34851) );
  NANDN U18807 ( .A(n34851), .B(n966), .Z(n18001) );
  AND U18808 ( .A(n18002), .B(n18001), .Z(n18351) );
  XOR U18809 ( .A(b[63]), .B(n18003), .Z(n18246) );
  NANDN U18810 ( .A(n18246), .B(n38422), .Z(n18006) );
  NANDN U18811 ( .A(n18004), .B(n38423), .Z(n18005) );
  AND U18812 ( .A(n18006), .B(n18005), .Z(n18352) );
  XNOR U18813 ( .A(n18351), .B(n18352), .Z(n18353) );
  XOR U18814 ( .A(n18354), .B(n18353), .Z(n18346) );
  XNOR U18815 ( .A(n18345), .B(n18346), .Z(n18347) );
  NANDN U18816 ( .A(n18008), .B(n18007), .Z(n18012) );
  NAND U18817 ( .A(n18010), .B(n18009), .Z(n18011) );
  AND U18818 ( .A(n18012), .B(n18011), .Z(n18348) );
  XNOR U18819 ( .A(n18347), .B(n18348), .Z(n18174) );
  NANDN U18820 ( .A(n18014), .B(n18013), .Z(n18018) );
  NAND U18821 ( .A(n18016), .B(n18015), .Z(n18017) );
  AND U18822 ( .A(n18018), .B(n18017), .Z(n18173) );
  XNOR U18823 ( .A(n18174), .B(n18173), .Z(n18175) );
  XNOR U18824 ( .A(n18176), .B(n18175), .Z(n18282) );
  XNOR U18825 ( .A(n18283), .B(n18282), .Z(n18285) );
  XNOR U18826 ( .A(n18284), .B(n18285), .Z(n18389) );
  XOR U18827 ( .A(n18390), .B(n18389), .Z(n18161) );
  NAND U18828 ( .A(n18020), .B(n18019), .Z(n18024) );
  NANDN U18829 ( .A(n18022), .B(n18021), .Z(n18023) );
  NAND U18830 ( .A(n18024), .B(n18023), .Z(n18403) );
  XNOR U18831 ( .A(n18403), .B(n18404), .Z(n18405) );
  NANDN U18832 ( .A(n18030), .B(n18029), .Z(n18034) );
  NAND U18833 ( .A(n18032), .B(n18031), .Z(n18033) );
  NAND U18834 ( .A(n18034), .B(n18033), .Z(n18342) );
  XNOR U18835 ( .A(b[15]), .B(a[77]), .Z(n18366) );
  OR U18836 ( .A(n18366), .B(n32010), .Z(n18037) );
  NANDN U18837 ( .A(n18035), .B(n32011), .Z(n18036) );
  NAND U18838 ( .A(n18037), .B(n18036), .Z(n18222) );
  XNOR U18839 ( .A(b[25]), .B(n29372), .Z(n18369) );
  NANDN U18840 ( .A(n34219), .B(n18369), .Z(n18040) );
  NAND U18841 ( .A(n34217), .B(n18038), .Z(n18039) );
  NAND U18842 ( .A(n18040), .B(n18039), .Z(n18219) );
  XOR U18843 ( .A(b[17]), .B(a[75]), .Z(n18372) );
  NAND U18844 ( .A(n18372), .B(n32543), .Z(n18043) );
  NANDN U18845 ( .A(n18041), .B(n32541), .Z(n18042) );
  AND U18846 ( .A(n18043), .B(n18042), .Z(n18220) );
  XNOR U18847 ( .A(n18219), .B(n18220), .Z(n18221) );
  XNOR U18848 ( .A(n18222), .B(n18221), .Z(n18276) );
  XOR U18849 ( .A(b[39]), .B(n25001), .Z(n18357) );
  NANDN U18850 ( .A(n18357), .B(n36553), .Z(n18046) );
  NANDN U18851 ( .A(n18044), .B(n36643), .Z(n18045) );
  NAND U18852 ( .A(n18046), .B(n18045), .Z(n18216) );
  XOR U18853 ( .A(b[51]), .B(n21441), .Z(n18360) );
  NANDN U18854 ( .A(n18360), .B(n37803), .Z(n18049) );
  NANDN U18855 ( .A(n18047), .B(n37802), .Z(n18048) );
  NAND U18856 ( .A(n18049), .B(n18048), .Z(n18213) );
  XOR U18857 ( .A(b[53]), .B(n20867), .Z(n18363) );
  NANDN U18858 ( .A(n18363), .B(n37940), .Z(n18052) );
  NANDN U18859 ( .A(n18050), .B(n37941), .Z(n18051) );
  AND U18860 ( .A(n18052), .B(n18051), .Z(n18214) );
  XNOR U18861 ( .A(n18213), .B(n18214), .Z(n18215) );
  XOR U18862 ( .A(n18216), .B(n18215), .Z(n18277) );
  XOR U18863 ( .A(n18276), .B(n18277), .Z(n18279) );
  NANDN U18864 ( .A(n18054), .B(n18053), .Z(n18058) );
  NAND U18865 ( .A(n18056), .B(n18055), .Z(n18057) );
  AND U18866 ( .A(n18058), .B(n18057), .Z(n18278) );
  XOR U18867 ( .A(n18279), .B(n18278), .Z(n18340) );
  NANDN U18868 ( .A(n18060), .B(n18059), .Z(n18064) );
  NAND U18869 ( .A(n18062), .B(n18061), .Z(n18063) );
  AND U18870 ( .A(n18064), .B(n18063), .Z(n18339) );
  XNOR U18871 ( .A(n18340), .B(n18339), .Z(n18341) );
  XOR U18872 ( .A(n18342), .B(n18341), .Z(n18406) );
  XNOR U18873 ( .A(n18405), .B(n18406), .Z(n18409) );
  XNOR U18874 ( .A(b[35]), .B(a[57]), .Z(n18288) );
  NANDN U18875 ( .A(n18288), .B(n35985), .Z(n18067) );
  NANDN U18876 ( .A(n18065), .B(n35986), .Z(n18066) );
  NAND U18877 ( .A(n18067), .B(n18066), .Z(n18384) );
  XNOR U18878 ( .A(a[85]), .B(n31123), .Z(n18291) );
  NAND U18879 ( .A(n18291), .B(n29949), .Z(n18070) );
  NAND U18880 ( .A(n29948), .B(n18068), .Z(n18069) );
  NAND U18881 ( .A(n18070), .B(n18069), .Z(n18381) );
  XOR U18882 ( .A(b[55]), .B(n20352), .Z(n18294) );
  NANDN U18883 ( .A(n18294), .B(n38075), .Z(n18073) );
  NANDN U18884 ( .A(n18071), .B(n38073), .Z(n18072) );
  AND U18885 ( .A(n18073), .B(n18072), .Z(n18382) );
  XNOR U18886 ( .A(n18381), .B(n18382), .Z(n18383) );
  XNOR U18887 ( .A(n18384), .B(n18383), .Z(n18170) );
  NANDN U18888 ( .A(n18075), .B(n18074), .Z(n18079) );
  NAND U18889 ( .A(n18077), .B(n18076), .Z(n18078) );
  NAND U18890 ( .A(n18079), .B(n18078), .Z(n18167) );
  NANDN U18891 ( .A(n18081), .B(n18080), .Z(n18085) );
  NAND U18892 ( .A(n18083), .B(n18082), .Z(n18084) );
  NAND U18893 ( .A(n18085), .B(n18084), .Z(n18168) );
  XNOR U18894 ( .A(n18167), .B(n18168), .Z(n18169) );
  XOR U18895 ( .A(n18170), .B(n18169), .Z(n18395) );
  OR U18896 ( .A(n18087), .B(n18086), .Z(n18091) );
  OR U18897 ( .A(n18089), .B(n18088), .Z(n18090) );
  NAND U18898 ( .A(n18091), .B(n18090), .Z(n18394) );
  XNOR U18899 ( .A(a[81]), .B(b[11]), .Z(n18309) );
  OR U18900 ( .A(n18309), .B(n31369), .Z(n18094) );
  NANDN U18901 ( .A(n18092), .B(n31119), .Z(n18093) );
  NAND U18902 ( .A(n18094), .B(n18093), .Z(n18330) );
  XOR U18903 ( .A(b[43]), .B(n23852), .Z(n18312) );
  NANDN U18904 ( .A(n18312), .B(n37068), .Z(n18097) );
  NANDN U18905 ( .A(n18095), .B(n37069), .Z(n18096) );
  NAND U18906 ( .A(n18097), .B(n18096), .Z(n18327) );
  XNOR U18907 ( .A(b[45]), .B(a[47]), .Z(n18315) );
  NANDN U18908 ( .A(n18315), .B(n37261), .Z(n18100) );
  NANDN U18909 ( .A(n18098), .B(n37262), .Z(n18099) );
  AND U18910 ( .A(n18100), .B(n18099), .Z(n18328) );
  XNOR U18911 ( .A(n18327), .B(n18328), .Z(n18329) );
  XNOR U18912 ( .A(n18330), .B(n18329), .Z(n18194) );
  XOR U18913 ( .A(b[49]), .B(n21996), .Z(n18318) );
  OR U18914 ( .A(n18318), .B(n37756), .Z(n18103) );
  NANDN U18915 ( .A(n18101), .B(n37652), .Z(n18102) );
  NAND U18916 ( .A(n18103), .B(n18102), .Z(n18306) );
  NAND U18917 ( .A(n37469), .B(n18104), .Z(n18106) );
  XOR U18918 ( .A(n978), .B(n22579), .Z(n18321) );
  NAND U18919 ( .A(n18321), .B(n37471), .Z(n18105) );
  NAND U18920 ( .A(n18106), .B(n18105), .Z(n18303) );
  XNOR U18921 ( .A(a[83]), .B(b[9]), .Z(n18324) );
  NANDN U18922 ( .A(n18324), .B(n30509), .Z(n18109) );
  NANDN U18923 ( .A(n18107), .B(n30846), .Z(n18108) );
  AND U18924 ( .A(n18109), .B(n18108), .Z(n18304) );
  XNOR U18925 ( .A(n18303), .B(n18304), .Z(n18305) );
  XNOR U18926 ( .A(n18306), .B(n18305), .Z(n18191) );
  NANDN U18927 ( .A(n18111), .B(n18110), .Z(n18115) );
  NAND U18928 ( .A(n18113), .B(n18112), .Z(n18114) );
  NAND U18929 ( .A(n18115), .B(n18114), .Z(n18192) );
  XNOR U18930 ( .A(n18191), .B(n18192), .Z(n18193) );
  XOR U18931 ( .A(n18194), .B(n18193), .Z(n18393) );
  XNOR U18932 ( .A(n18394), .B(n18393), .Z(n18396) );
  XNOR U18933 ( .A(n18395), .B(n18396), .Z(n18410) );
  NAND U18934 ( .A(n18117), .B(n18116), .Z(n18121) );
  NANDN U18935 ( .A(n18119), .B(n18118), .Z(n18120) );
  AND U18936 ( .A(n18121), .B(n18120), .Z(n18412) );
  XNOR U18937 ( .A(n18411), .B(n18412), .Z(n18162) );
  XNOR U18938 ( .A(n18161), .B(n18162), .Z(n18163) );
  OR U18939 ( .A(n18123), .B(n18122), .Z(n18127) );
  NAND U18940 ( .A(n18125), .B(n18124), .Z(n18126) );
  AND U18941 ( .A(n18127), .B(n18126), .Z(n18164) );
  XNOR U18942 ( .A(n18163), .B(n18164), .Z(n18417) );
  XNOR U18943 ( .A(n18418), .B(n18417), .Z(n18424) );
  NANDN U18944 ( .A(n18129), .B(n18128), .Z(n18133) );
  NAND U18945 ( .A(n18131), .B(n18130), .Z(n18132) );
  NAND U18946 ( .A(n18133), .B(n18132), .Z(n18421) );
  NAND U18947 ( .A(n18135), .B(n18134), .Z(n18139) );
  NANDN U18948 ( .A(n18137), .B(n18136), .Z(n18138) );
  NAND U18949 ( .A(n18139), .B(n18138), .Z(n18422) );
  XNOR U18950 ( .A(n18421), .B(n18422), .Z(n18423) );
  XOR U18951 ( .A(n18424), .B(n18423), .Z(n18152) );
  XOR U18952 ( .A(n18151), .B(n18152), .Z(n18145) );
  XNOR U18953 ( .A(n18146), .B(n18145), .Z(n18147) );
  XNOR U18954 ( .A(n18148), .B(n18147), .Z(n18427) );
  XNOR U18955 ( .A(n18427), .B(sreg[155]), .Z(n18429) );
  NAND U18956 ( .A(n18140), .B(sreg[154]), .Z(n18144) );
  OR U18957 ( .A(n18142), .B(n18141), .Z(n18143) );
  AND U18958 ( .A(n18144), .B(n18143), .Z(n18428) );
  XOR U18959 ( .A(n18429), .B(n18428), .Z(c[155]) );
  NANDN U18960 ( .A(n18150), .B(n18149), .Z(n18154) );
  NAND U18961 ( .A(n18152), .B(n18151), .Z(n18153) );
  NAND U18962 ( .A(n18154), .B(n18153), .Z(n18432) );
  NANDN U18963 ( .A(n18156), .B(n18155), .Z(n18160) );
  NAND U18964 ( .A(n18158), .B(n18157), .Z(n18159) );
  NAND U18965 ( .A(n18160), .B(n18159), .Z(n18701) );
  NANDN U18966 ( .A(n18162), .B(n18161), .Z(n18166) );
  NAND U18967 ( .A(n18164), .B(n18163), .Z(n18165) );
  NAND U18968 ( .A(n18166), .B(n18165), .Z(n18702) );
  XNOR U18969 ( .A(n18701), .B(n18702), .Z(n18703) );
  NANDN U18970 ( .A(n18168), .B(n18167), .Z(n18172) );
  NAND U18971 ( .A(n18170), .B(n18169), .Z(n18171) );
  NAND U18972 ( .A(n18172), .B(n18171), .Z(n18674) );
  NANDN U18973 ( .A(n18174), .B(n18173), .Z(n18178) );
  NANDN U18974 ( .A(n18176), .B(n18175), .Z(n18177) );
  NAND U18975 ( .A(n18178), .B(n18177), .Z(n18671) );
  NANDN U18976 ( .A(n18180), .B(n18179), .Z(n18184) );
  NAND U18977 ( .A(n18182), .B(n18181), .Z(n18183) );
  AND U18978 ( .A(n18184), .B(n18183), .Z(n18672) );
  XNOR U18979 ( .A(n18671), .B(n18672), .Z(n18673) );
  XNOR U18980 ( .A(n18674), .B(n18673), .Z(n18439) );
  OR U18981 ( .A(n18186), .B(n18185), .Z(n18190) );
  NANDN U18982 ( .A(n18188), .B(n18187), .Z(n18189) );
  AND U18983 ( .A(n18190), .B(n18189), .Z(n18438) );
  XNOR U18984 ( .A(n18439), .B(n18438), .Z(n18440) );
  XOR U18985 ( .A(b[37]), .B(n25860), .Z(n18573) );
  NANDN U18986 ( .A(n18573), .B(n36311), .Z(n18197) );
  NANDN U18987 ( .A(n18195), .B(n36309), .Z(n18196) );
  NAND U18988 ( .A(n18197), .B(n18196), .Z(n18652) );
  XOR U18989 ( .A(a[88]), .B(n968), .Z(n18576) );
  OR U18990 ( .A(n18576), .B(n29363), .Z(n18200) );
  NANDN U18991 ( .A(n18198), .B(n29864), .Z(n18199) );
  NAND U18992 ( .A(n18200), .B(n18199), .Z(n18649) );
  XOR U18993 ( .A(n34851), .B(n967), .Z(n18579) );
  NAND U18994 ( .A(n18579), .B(n28939), .Z(n18203) );
  NAND U18995 ( .A(n28938), .B(n18201), .Z(n18202) );
  AND U18996 ( .A(n18203), .B(n18202), .Z(n18650) );
  XNOR U18997 ( .A(n18649), .B(n18650), .Z(n18651) );
  XNOR U18998 ( .A(n18652), .B(n18651), .Z(n18554) );
  XOR U18999 ( .A(a[80]), .B(n971), .Z(n18582) );
  OR U19000 ( .A(n18582), .B(n31550), .Z(n18206) );
  NANDN U19001 ( .A(n18204), .B(n31874), .Z(n18205) );
  NAND U19002 ( .A(n18206), .B(n18205), .Z(n18477) );
  NAND U19003 ( .A(n34848), .B(n18207), .Z(n18209) );
  XOR U19004 ( .A(n35375), .B(n28701), .Z(n18585) );
  NAND U19005 ( .A(n34618), .B(n18585), .Z(n18208) );
  NAND U19006 ( .A(n18209), .B(n18208), .Z(n18474) );
  NAND U19007 ( .A(n35188), .B(n18210), .Z(n18212) );
  XNOR U19008 ( .A(n35540), .B(a[64]), .Z(n18588) );
  NANDN U19009 ( .A(n34968), .B(n18588), .Z(n18211) );
  AND U19010 ( .A(n18212), .B(n18211), .Z(n18475) );
  XNOR U19011 ( .A(n18474), .B(n18475), .Z(n18476) );
  XNOR U19012 ( .A(n18477), .B(n18476), .Z(n18551) );
  NANDN U19013 ( .A(n18214), .B(n18213), .Z(n18218) );
  NAND U19014 ( .A(n18216), .B(n18215), .Z(n18217) );
  NAND U19015 ( .A(n18218), .B(n18217), .Z(n18552) );
  XNOR U19016 ( .A(n18551), .B(n18552), .Z(n18553) );
  XOR U19017 ( .A(n18554), .B(n18553), .Z(n18564) );
  NANDN U19018 ( .A(n18220), .B(n18219), .Z(n18224) );
  NAND U19019 ( .A(n18222), .B(n18221), .Z(n18223) );
  NAND U19020 ( .A(n18224), .B(n18223), .Z(n18516) );
  NAND U19021 ( .A(a[28]), .B(b[63]), .Z(n18530) );
  NANDN U19022 ( .A(n18225), .B(n38369), .Z(n18227) );
  XOR U19023 ( .A(b[61]), .B(n18841), .Z(n18603) );
  OR U19024 ( .A(n18603), .B(n38371), .Z(n18226) );
  NAND U19025 ( .A(n18227), .B(n18226), .Z(n18528) );
  NANDN U19026 ( .A(n18228), .B(n35311), .Z(n18230) );
  XNOR U19027 ( .A(b[31]), .B(a[62]), .Z(n18606) );
  NANDN U19028 ( .A(n18606), .B(n35313), .Z(n18229) );
  AND U19029 ( .A(n18230), .B(n18229), .Z(n18527) );
  XNOR U19030 ( .A(n18528), .B(n18527), .Z(n18529) );
  XOR U19031 ( .A(n18530), .B(n18529), .Z(n18514) );
  NAND U19032 ( .A(n33283), .B(n18231), .Z(n18233) );
  XOR U19033 ( .A(n33020), .B(n31372), .Z(n18609) );
  NANDN U19034 ( .A(n33021), .B(n18609), .Z(n18232) );
  NAND U19035 ( .A(n18233), .B(n18232), .Z(n18621) );
  XNOR U19036 ( .A(b[21]), .B(a[72]), .Z(n18612) );
  OR U19037 ( .A(n18612), .B(n33634), .Z(n18236) );
  NANDN U19038 ( .A(n18234), .B(n33464), .Z(n18235) );
  NAND U19039 ( .A(n18236), .B(n18235), .Z(n18618) );
  NAND U19040 ( .A(n34044), .B(n18237), .Z(n18239) );
  XOR U19041 ( .A(n34510), .B(n30379), .Z(n18615) );
  NANDN U19042 ( .A(n33867), .B(n18615), .Z(n18238) );
  AND U19043 ( .A(n18239), .B(n18238), .Z(n18619) );
  XNOR U19044 ( .A(n18618), .B(n18619), .Z(n18620) );
  XNOR U19045 ( .A(n18621), .B(n18620), .Z(n18515) );
  XNOR U19046 ( .A(n18514), .B(n18515), .Z(n18517) );
  XNOR U19047 ( .A(n18516), .B(n18517), .Z(n18563) );
  XOR U19048 ( .A(n18564), .B(n18563), .Z(n18566) );
  XNOR U19049 ( .A(n18565), .B(n18566), .Z(n18542) );
  XOR U19050 ( .A(b[33]), .B(n27436), .Z(n18633) );
  NANDN U19051 ( .A(n18633), .B(n35620), .Z(n18242) );
  NANDN U19052 ( .A(n18240), .B(n35621), .Z(n18241) );
  NAND U19053 ( .A(n18242), .B(n18241), .Z(n18489) );
  NANDN U19054 ( .A(n966), .B(a[92]), .Z(n18243) );
  XOR U19055 ( .A(n29232), .B(n18243), .Z(n18245) );
  NANDN U19056 ( .A(b[0]), .B(a[91]), .Z(n18244) );
  AND U19057 ( .A(n18245), .B(n18244), .Z(n18486) );
  XOR U19058 ( .A(b[63]), .B(n18804), .Z(n18640) );
  NANDN U19059 ( .A(n18640), .B(n38422), .Z(n18248) );
  NANDN U19060 ( .A(n18246), .B(n38423), .Z(n18247) );
  AND U19061 ( .A(n18248), .B(n18247), .Z(n18487) );
  XNOR U19062 ( .A(n18486), .B(n18487), .Z(n18488) );
  XNOR U19063 ( .A(n18489), .B(n18488), .Z(n18452) );
  XNOR U19064 ( .A(b[41]), .B(a[52]), .Z(n18624) );
  OR U19065 ( .A(n18624), .B(n36905), .Z(n18251) );
  NANDN U19066 ( .A(n18249), .B(n36807), .Z(n18250) );
  NAND U19067 ( .A(n18251), .B(n18250), .Z(n18646) );
  XOR U19068 ( .A(b[57]), .B(n19980), .Z(n18627) );
  OR U19069 ( .A(n18627), .B(n965), .Z(n18254) );
  NANDN U19070 ( .A(n18252), .B(n38194), .Z(n18253) );
  NAND U19071 ( .A(n18254), .B(n18253), .Z(n18643) );
  NAND U19072 ( .A(n38326), .B(n18255), .Z(n18257) );
  XOR U19073 ( .A(n38400), .B(n19513), .Z(n18630) );
  NANDN U19074 ( .A(n38273), .B(n18630), .Z(n18256) );
  AND U19075 ( .A(n18257), .B(n18256), .Z(n18644) );
  XNOR U19076 ( .A(n18643), .B(n18644), .Z(n18645) );
  XOR U19077 ( .A(n18646), .B(n18645), .Z(n18451) );
  NANDN U19078 ( .A(n18259), .B(n18258), .Z(n18263) );
  NAND U19079 ( .A(n18261), .B(n18260), .Z(n18262) );
  AND U19080 ( .A(n18263), .B(n18262), .Z(n18450) );
  XOR U19081 ( .A(n18451), .B(n18450), .Z(n18453) );
  XNOR U19082 ( .A(n18452), .B(n18453), .Z(n18560) );
  NANDN U19083 ( .A(n18265), .B(n18264), .Z(n18269) );
  NAND U19084 ( .A(n18267), .B(n18266), .Z(n18268) );
  NAND U19085 ( .A(n18269), .B(n18268), .Z(n18557) );
  NANDN U19086 ( .A(n18271), .B(n18270), .Z(n18275) );
  NAND U19087 ( .A(n18273), .B(n18272), .Z(n18274) );
  AND U19088 ( .A(n18275), .B(n18274), .Z(n18558) );
  XNOR U19089 ( .A(n18557), .B(n18558), .Z(n18559) );
  XNOR U19090 ( .A(n18560), .B(n18559), .Z(n18540) );
  NANDN U19091 ( .A(n18277), .B(n18276), .Z(n18281) );
  NANDN U19092 ( .A(n18279), .B(n18278), .Z(n18280) );
  AND U19093 ( .A(n18281), .B(n18280), .Z(n18539) );
  XOR U19094 ( .A(n18540), .B(n18539), .Z(n18541) );
  XNOR U19095 ( .A(n18542), .B(n18541), .Z(n18441) );
  XOR U19096 ( .A(n18440), .B(n18441), .Z(n18683) );
  NAND U19097 ( .A(n18283), .B(n18282), .Z(n18287) );
  NANDN U19098 ( .A(n18285), .B(n18284), .Z(n18286) );
  NAND U19099 ( .A(n18287), .B(n18286), .Z(n18680) );
  XNOR U19100 ( .A(b[35]), .B(a[58]), .Z(n18518) );
  NANDN U19101 ( .A(n18518), .B(n35985), .Z(n18290) );
  NANDN U19102 ( .A(n18288), .B(n35986), .Z(n18289) );
  NAND U19103 ( .A(n18290), .B(n18289), .Z(n18483) );
  XOR U19104 ( .A(n33628), .B(n31123), .Z(n18521) );
  NAND U19105 ( .A(n18521), .B(n29949), .Z(n18293) );
  NAND U19106 ( .A(n29948), .B(n18291), .Z(n18292) );
  NAND U19107 ( .A(n18293), .B(n18292), .Z(n18480) );
  XOR U19108 ( .A(b[55]), .B(n20686), .Z(n18524) );
  NANDN U19109 ( .A(n18524), .B(n38075), .Z(n18296) );
  NANDN U19110 ( .A(n18294), .B(n38073), .Z(n18295) );
  AND U19111 ( .A(n18296), .B(n18295), .Z(n18481) );
  XNOR U19112 ( .A(n18480), .B(n18481), .Z(n18482) );
  XNOR U19113 ( .A(n18483), .B(n18482), .Z(n18548) );
  NANDN U19114 ( .A(n18298), .B(n18297), .Z(n18302) );
  NANDN U19115 ( .A(n18300), .B(n18299), .Z(n18301) );
  NAND U19116 ( .A(n18302), .B(n18301), .Z(n18545) );
  NANDN U19117 ( .A(n18304), .B(n18303), .Z(n18308) );
  NAND U19118 ( .A(n18306), .B(n18305), .Z(n18307) );
  NAND U19119 ( .A(n18308), .B(n18307), .Z(n18546) );
  XNOR U19120 ( .A(n18545), .B(n18546), .Z(n18547) );
  XOR U19121 ( .A(n18548), .B(n18547), .Z(n18661) );
  XOR U19122 ( .A(a[82]), .B(n970), .Z(n18490) );
  OR U19123 ( .A(n18490), .B(n31369), .Z(n18311) );
  NANDN U19124 ( .A(n18309), .B(n31119), .Z(n18310) );
  NAND U19125 ( .A(n18311), .B(n18310), .Z(n18511) );
  XOR U19126 ( .A(b[43]), .B(n24671), .Z(n18493) );
  NANDN U19127 ( .A(n18493), .B(n37068), .Z(n18314) );
  NANDN U19128 ( .A(n18312), .B(n37069), .Z(n18313) );
  NAND U19129 ( .A(n18314), .B(n18313), .Z(n18508) );
  XNOR U19130 ( .A(b[45]), .B(a[48]), .Z(n18496) );
  NANDN U19131 ( .A(n18496), .B(n37261), .Z(n18317) );
  NANDN U19132 ( .A(n18315), .B(n37262), .Z(n18316) );
  AND U19133 ( .A(n18317), .B(n18316), .Z(n18509) );
  XNOR U19134 ( .A(n18508), .B(n18509), .Z(n18510) );
  XNOR U19135 ( .A(n18511), .B(n18510), .Z(n18572) );
  XOR U19136 ( .A(b[49]), .B(n22289), .Z(n18499) );
  OR U19137 ( .A(n18499), .B(n37756), .Z(n18320) );
  NANDN U19138 ( .A(n18318), .B(n37652), .Z(n18319) );
  NAND U19139 ( .A(n18320), .B(n18319), .Z(n18536) );
  NAND U19140 ( .A(n37469), .B(n18321), .Z(n18323) );
  XOR U19141 ( .A(n978), .B(n22964), .Z(n18502) );
  NAND U19142 ( .A(n18502), .B(n37471), .Z(n18322) );
  NAND U19143 ( .A(n18323), .B(n18322), .Z(n18533) );
  XOR U19144 ( .A(a[84]), .B(n969), .Z(n18505) );
  NANDN U19145 ( .A(n18505), .B(n30509), .Z(n18326) );
  NANDN U19146 ( .A(n18324), .B(n30846), .Z(n18325) );
  AND U19147 ( .A(n18326), .B(n18325), .Z(n18534) );
  XNOR U19148 ( .A(n18533), .B(n18534), .Z(n18535) );
  XNOR U19149 ( .A(n18536), .B(n18535), .Z(n18569) );
  NANDN U19150 ( .A(n18328), .B(n18327), .Z(n18332) );
  NAND U19151 ( .A(n18330), .B(n18329), .Z(n18331) );
  NAND U19152 ( .A(n18332), .B(n18331), .Z(n18570) );
  XNOR U19153 ( .A(n18569), .B(n18570), .Z(n18571) );
  XOR U19154 ( .A(n18572), .B(n18571), .Z(n18659) );
  NANDN U19155 ( .A(n18334), .B(n18333), .Z(n18338) );
  NAND U19156 ( .A(n18336), .B(n18335), .Z(n18337) );
  AND U19157 ( .A(n18338), .B(n18337), .Z(n18660) );
  XOR U19158 ( .A(n18659), .B(n18660), .Z(n18662) );
  XNOR U19159 ( .A(n18661), .B(n18662), .Z(n18678) );
  NANDN U19160 ( .A(n18340), .B(n18339), .Z(n18344) );
  NANDN U19161 ( .A(n18342), .B(n18341), .Z(n18343) );
  NAND U19162 ( .A(n18344), .B(n18343), .Z(n18665) );
  NANDN U19163 ( .A(n18346), .B(n18345), .Z(n18350) );
  NAND U19164 ( .A(n18348), .B(n18347), .Z(n18349) );
  AND U19165 ( .A(n18350), .B(n18349), .Z(n18666) );
  XNOR U19166 ( .A(n18665), .B(n18666), .Z(n18667) );
  NANDN U19167 ( .A(n18352), .B(n18351), .Z(n18356) );
  NAND U19168 ( .A(n18354), .B(n18353), .Z(n18355) );
  NAND U19169 ( .A(n18356), .B(n18355), .Z(n18447) );
  XOR U19170 ( .A(b[39]), .B(n25177), .Z(n18465) );
  NANDN U19171 ( .A(n18465), .B(n36553), .Z(n18359) );
  NANDN U19172 ( .A(n18357), .B(n36643), .Z(n18358) );
  NAND U19173 ( .A(n18359), .B(n18358), .Z(n18594) );
  XOR U19174 ( .A(b[51]), .B(n22246), .Z(n18468) );
  NANDN U19175 ( .A(n18468), .B(n37803), .Z(n18362) );
  NANDN U19176 ( .A(n18360), .B(n37802), .Z(n18361) );
  NAND U19177 ( .A(n18362), .B(n18361), .Z(n18591) );
  XOR U19178 ( .A(b[53]), .B(n21149), .Z(n18471) );
  NANDN U19179 ( .A(n18471), .B(n37940), .Z(n18365) );
  NANDN U19180 ( .A(n18363), .B(n37941), .Z(n18364) );
  AND U19181 ( .A(n18365), .B(n18364), .Z(n18592) );
  XNOR U19182 ( .A(n18591), .B(n18592), .Z(n18593) );
  XNOR U19183 ( .A(n18594), .B(n18593), .Z(n18658) );
  XOR U19184 ( .A(b[15]), .B(n31870), .Z(n18456) );
  OR U19185 ( .A(n18456), .B(n32010), .Z(n18368) );
  NANDN U19186 ( .A(n18366), .B(n32011), .Z(n18367) );
  NAND U19187 ( .A(n18368), .B(n18367), .Z(n18600) );
  XNOR U19188 ( .A(b[25]), .B(n29868), .Z(n18459) );
  NANDN U19189 ( .A(n34219), .B(n18459), .Z(n18371) );
  NAND U19190 ( .A(n34217), .B(n18369), .Z(n18370) );
  NAND U19191 ( .A(n18371), .B(n18370), .Z(n18597) );
  XNOR U19192 ( .A(b[17]), .B(a[76]), .Z(n18462) );
  NANDN U19193 ( .A(n18462), .B(n32543), .Z(n18374) );
  NAND U19194 ( .A(n18372), .B(n32541), .Z(n18373) );
  AND U19195 ( .A(n18374), .B(n18373), .Z(n18598) );
  XNOR U19196 ( .A(n18597), .B(n18598), .Z(n18599) );
  XNOR U19197 ( .A(n18600), .B(n18599), .Z(n18655) );
  NANDN U19198 ( .A(n18376), .B(n18375), .Z(n18380) );
  NAND U19199 ( .A(n18378), .B(n18377), .Z(n18379) );
  NAND U19200 ( .A(n18380), .B(n18379), .Z(n18656) );
  XNOR U19201 ( .A(n18655), .B(n18656), .Z(n18657) );
  XOR U19202 ( .A(n18658), .B(n18657), .Z(n18444) );
  NANDN U19203 ( .A(n18382), .B(n18381), .Z(n18386) );
  NAND U19204 ( .A(n18384), .B(n18383), .Z(n18385) );
  AND U19205 ( .A(n18386), .B(n18385), .Z(n18445) );
  XOR U19206 ( .A(n18444), .B(n18445), .Z(n18446) );
  XOR U19207 ( .A(n18447), .B(n18446), .Z(n18668) );
  XNOR U19208 ( .A(n18667), .B(n18668), .Z(n18677) );
  XOR U19209 ( .A(n18680), .B(n18679), .Z(n18684) );
  XNOR U19210 ( .A(n18683), .B(n18684), .Z(n18685) );
  NAND U19211 ( .A(n18388), .B(n18387), .Z(n18392) );
  NANDN U19212 ( .A(n18390), .B(n18389), .Z(n18391) );
  NAND U19213 ( .A(n18392), .B(n18391), .Z(n18686) );
  XOR U19214 ( .A(n18685), .B(n18686), .Z(n18698) );
  NAND U19215 ( .A(n18394), .B(n18393), .Z(n18398) );
  NANDN U19216 ( .A(n18396), .B(n18395), .Z(n18397) );
  NAND U19217 ( .A(n18398), .B(n18397), .Z(n18692) );
  NANDN U19218 ( .A(n18404), .B(n18403), .Z(n18408) );
  NANDN U19219 ( .A(n18406), .B(n18405), .Z(n18407) );
  AND U19220 ( .A(n18408), .B(n18407), .Z(n18689) );
  XNOR U19221 ( .A(n18690), .B(n18689), .Z(n18691) );
  XNOR U19222 ( .A(n18692), .B(n18691), .Z(n18695) );
  OR U19223 ( .A(n18410), .B(n18409), .Z(n18414) );
  NAND U19224 ( .A(n18412), .B(n18411), .Z(n18413) );
  NAND U19225 ( .A(n18414), .B(n18413), .Z(n18696) );
  XNOR U19226 ( .A(n18698), .B(n18697), .Z(n18704) );
  XOR U19227 ( .A(n18703), .B(n18704), .Z(n18710) );
  OR U19228 ( .A(n18416), .B(n18415), .Z(n18420) );
  OR U19229 ( .A(n18418), .B(n18417), .Z(n18419) );
  NAND U19230 ( .A(n18420), .B(n18419), .Z(n18707) );
  NANDN U19231 ( .A(n18422), .B(n18421), .Z(n18426) );
  NAND U19232 ( .A(n18424), .B(n18423), .Z(n18425) );
  NAND U19233 ( .A(n18426), .B(n18425), .Z(n18708) );
  XNOR U19234 ( .A(n18707), .B(n18708), .Z(n18709) );
  XOR U19235 ( .A(n18710), .B(n18709), .Z(n18433) );
  XNOR U19236 ( .A(n18432), .B(n18433), .Z(n18434) );
  XNOR U19237 ( .A(n18435), .B(n18434), .Z(n18713) );
  XNOR U19238 ( .A(n18713), .B(sreg[156]), .Z(n18715) );
  NAND U19239 ( .A(n18427), .B(sreg[155]), .Z(n18431) );
  OR U19240 ( .A(n18429), .B(n18428), .Z(n18430) );
  AND U19241 ( .A(n18431), .B(n18430), .Z(n18714) );
  XOR U19242 ( .A(n18715), .B(n18714), .Z(c[156]) );
  NANDN U19243 ( .A(n18433), .B(n18432), .Z(n18437) );
  NAND U19244 ( .A(n18435), .B(n18434), .Z(n18436) );
  NAND U19245 ( .A(n18437), .B(n18436), .Z(n18721) );
  NANDN U19246 ( .A(n18439), .B(n18438), .Z(n18443) );
  NANDN U19247 ( .A(n18441), .B(n18440), .Z(n18442) );
  NAND U19248 ( .A(n18443), .B(n18442), .Z(n18745) );
  NAND U19249 ( .A(n18445), .B(n18444), .Z(n18449) );
  NANDN U19250 ( .A(n18447), .B(n18446), .Z(n18448) );
  NAND U19251 ( .A(n18449), .B(n18448), .Z(n18987) );
  NANDN U19252 ( .A(n18451), .B(n18450), .Z(n18455) );
  NANDN U19253 ( .A(n18453), .B(n18452), .Z(n18454) );
  NAND U19254 ( .A(n18455), .B(n18454), .Z(n18984) );
  XNOR U19255 ( .A(b[15]), .B(a[79]), .Z(n18918) );
  OR U19256 ( .A(n18918), .B(n32010), .Z(n18458) );
  NANDN U19257 ( .A(n18456), .B(n32011), .Z(n18457) );
  NAND U19258 ( .A(n18458), .B(n18457), .Z(n18801) );
  XOR U19259 ( .A(b[25]), .B(a[69]), .Z(n18921) );
  NANDN U19260 ( .A(n34219), .B(n18921), .Z(n18461) );
  NAND U19261 ( .A(n34217), .B(n18459), .Z(n18460) );
  NAND U19262 ( .A(n18461), .B(n18460), .Z(n18798) );
  XOR U19263 ( .A(b[17]), .B(a[77]), .Z(n18924) );
  NAND U19264 ( .A(n18924), .B(n32543), .Z(n18464) );
  NANDN U19265 ( .A(n18462), .B(n32541), .Z(n18463) );
  AND U19266 ( .A(n18464), .B(n18463), .Z(n18799) );
  XNOR U19267 ( .A(n18798), .B(n18799), .Z(n18800) );
  XNOR U19268 ( .A(n18801), .B(n18800), .Z(n18857) );
  XOR U19269 ( .A(b[39]), .B(n25466), .Z(n18927) );
  NANDN U19270 ( .A(n18927), .B(n36553), .Z(n18467) );
  NANDN U19271 ( .A(n18465), .B(n36643), .Z(n18466) );
  NAND U19272 ( .A(n18467), .B(n18466), .Z(n18795) );
  XOR U19273 ( .A(b[51]), .B(n21996), .Z(n18930) );
  NANDN U19274 ( .A(n18930), .B(n37803), .Z(n18470) );
  NANDN U19275 ( .A(n18468), .B(n37802), .Z(n18469) );
  NAND U19276 ( .A(n18470), .B(n18469), .Z(n18792) );
  XOR U19277 ( .A(b[53]), .B(n21441), .Z(n18933) );
  NANDN U19278 ( .A(n18933), .B(n37940), .Z(n18473) );
  NANDN U19279 ( .A(n18471), .B(n37941), .Z(n18472) );
  AND U19280 ( .A(n18473), .B(n18472), .Z(n18793) );
  XNOR U19281 ( .A(n18792), .B(n18793), .Z(n18794) );
  XOR U19282 ( .A(n18795), .B(n18794), .Z(n18858) );
  XOR U19283 ( .A(n18857), .B(n18858), .Z(n18860) );
  NANDN U19284 ( .A(n18475), .B(n18474), .Z(n18479) );
  NAND U19285 ( .A(n18477), .B(n18476), .Z(n18478) );
  NAND U19286 ( .A(n18479), .B(n18478), .Z(n18859) );
  XNOR U19287 ( .A(n18860), .B(n18859), .Z(n18963) );
  NANDN U19288 ( .A(n18481), .B(n18480), .Z(n18485) );
  NAND U19289 ( .A(n18483), .B(n18482), .Z(n18484) );
  NAND U19290 ( .A(n18485), .B(n18484), .Z(n18960) );
  XNOR U19291 ( .A(n18960), .B(n18961), .Z(n18962) );
  XOR U19292 ( .A(n18963), .B(n18962), .Z(n18985) );
  XNOR U19293 ( .A(n18984), .B(n18985), .Z(n18986) );
  XNOR U19294 ( .A(n18987), .B(n18986), .Z(n18972) );
  XNOR U19295 ( .A(a[83]), .B(b[11]), .Z(n18869) );
  OR U19296 ( .A(n18869), .B(n31369), .Z(n18492) );
  NANDN U19297 ( .A(n18490), .B(n31119), .Z(n18491) );
  NAND U19298 ( .A(n18492), .B(n18491), .Z(n18890) );
  XOR U19299 ( .A(b[43]), .B(n24288), .Z(n18872) );
  NANDN U19300 ( .A(n18872), .B(n37068), .Z(n18495) );
  NANDN U19301 ( .A(n18493), .B(n37069), .Z(n18494) );
  NAND U19302 ( .A(n18495), .B(n18494), .Z(n18887) );
  XNOR U19303 ( .A(b[45]), .B(a[49]), .Z(n18875) );
  NANDN U19304 ( .A(n18875), .B(n37261), .Z(n18498) );
  NANDN U19305 ( .A(n18496), .B(n37262), .Z(n18497) );
  AND U19306 ( .A(n18498), .B(n18497), .Z(n18888) );
  XNOR U19307 ( .A(n18887), .B(n18888), .Z(n18889) );
  XNOR U19308 ( .A(n18890), .B(n18889), .Z(n18773) );
  XOR U19309 ( .A(b[49]), .B(n22579), .Z(n18878) );
  OR U19310 ( .A(n18878), .B(n37756), .Z(n18501) );
  NANDN U19311 ( .A(n18499), .B(n37652), .Z(n18500) );
  NAND U19312 ( .A(n18501), .B(n18500), .Z(n18914) );
  NAND U19313 ( .A(n37469), .B(n18502), .Z(n18504) );
  XOR U19314 ( .A(n978), .B(n23149), .Z(n18881) );
  NAND U19315 ( .A(n18881), .B(n37471), .Z(n18503) );
  AND U19316 ( .A(n18504), .B(n18503), .Z(n18912) );
  XNOR U19317 ( .A(a[85]), .B(b[9]), .Z(n18884) );
  NANDN U19318 ( .A(n18884), .B(n30509), .Z(n18507) );
  NANDN U19319 ( .A(n18505), .B(n30846), .Z(n18506) );
  AND U19320 ( .A(n18507), .B(n18506), .Z(n18913) );
  XOR U19321 ( .A(n18914), .B(n18915), .Z(n18770) );
  NANDN U19322 ( .A(n18509), .B(n18508), .Z(n18513) );
  NAND U19323 ( .A(n18511), .B(n18510), .Z(n18512) );
  NAND U19324 ( .A(n18513), .B(n18512), .Z(n18771) );
  XNOR U19325 ( .A(n18770), .B(n18771), .Z(n18772) );
  XOR U19326 ( .A(n18773), .B(n18772), .Z(n18978) );
  XNOR U19327 ( .A(n18978), .B(n18979), .Z(n18981) );
  XOR U19328 ( .A(b[35]), .B(a[59]), .Z(n18897) );
  NAND U19329 ( .A(n35985), .B(n18897), .Z(n18520) );
  NANDN U19330 ( .A(n18518), .B(n35986), .Z(n18519) );
  NAND U19331 ( .A(n18520), .B(n18519), .Z(n18945) );
  XNOR U19332 ( .A(a[87]), .B(n31123), .Z(n18900) );
  NAND U19333 ( .A(n18900), .B(n29949), .Z(n18523) );
  NAND U19334 ( .A(n29948), .B(n18521), .Z(n18522) );
  NAND U19335 ( .A(n18523), .B(n18522), .Z(n18942) );
  XOR U19336 ( .A(b[55]), .B(n20867), .Z(n18903) );
  NANDN U19337 ( .A(n18903), .B(n38075), .Z(n18526) );
  NANDN U19338 ( .A(n18524), .B(n38073), .Z(n18525) );
  AND U19339 ( .A(n18526), .B(n18525), .Z(n18943) );
  XNOR U19340 ( .A(n18942), .B(n18943), .Z(n18944) );
  XNOR U19341 ( .A(n18945), .B(n18944), .Z(n18749) );
  NANDN U19342 ( .A(n18528), .B(n18527), .Z(n18532) );
  NAND U19343 ( .A(n18530), .B(n18529), .Z(n18531) );
  NAND U19344 ( .A(n18532), .B(n18531), .Z(n18746) );
  NANDN U19345 ( .A(n18534), .B(n18533), .Z(n18538) );
  NAND U19346 ( .A(n18536), .B(n18535), .Z(n18537) );
  NAND U19347 ( .A(n18538), .B(n18537), .Z(n18747) );
  XNOR U19348 ( .A(n18746), .B(n18747), .Z(n18748) );
  XOR U19349 ( .A(n18749), .B(n18748), .Z(n18980) );
  XNOR U19350 ( .A(n18981), .B(n18980), .Z(n18973) );
  XNOR U19351 ( .A(n18972), .B(n18973), .Z(n18974) );
  OR U19352 ( .A(n18540), .B(n18539), .Z(n18544) );
  NAND U19353 ( .A(n18542), .B(n18541), .Z(n18543) );
  NAND U19354 ( .A(n18544), .B(n18543), .Z(n18975) );
  XOR U19355 ( .A(n18974), .B(n18975), .Z(n18743) );
  NANDN U19356 ( .A(n18546), .B(n18545), .Z(n18550) );
  NAND U19357 ( .A(n18548), .B(n18547), .Z(n18549) );
  AND U19358 ( .A(n18550), .B(n18549), .Z(n18993) );
  NANDN U19359 ( .A(n18552), .B(n18551), .Z(n18556) );
  NAND U19360 ( .A(n18554), .B(n18553), .Z(n18555) );
  NAND U19361 ( .A(n18556), .B(n18555), .Z(n18990) );
  NANDN U19362 ( .A(n18558), .B(n18557), .Z(n18562) );
  NANDN U19363 ( .A(n18560), .B(n18559), .Z(n18561) );
  NAND U19364 ( .A(n18562), .B(n18561), .Z(n18991) );
  XNOR U19365 ( .A(n18990), .B(n18991), .Z(n18992) );
  XNOR U19366 ( .A(n18993), .B(n18992), .Z(n18966) );
  NANDN U19367 ( .A(n18564), .B(n18563), .Z(n18568) );
  OR U19368 ( .A(n18566), .B(n18565), .Z(n18567) );
  AND U19369 ( .A(n18568), .B(n18567), .Z(n18967) );
  XNOR U19370 ( .A(n18966), .B(n18967), .Z(n18969) );
  XOR U19371 ( .A(b[37]), .B(n26122), .Z(n18783) );
  NANDN U19372 ( .A(n18783), .B(n36311), .Z(n18575) );
  NANDN U19373 ( .A(n18573), .B(n36309), .Z(n18574) );
  NAND U19374 ( .A(n18575), .B(n18574), .Z(n18854) );
  XNOR U19375 ( .A(a[89]), .B(b[5]), .Z(n18786) );
  OR U19376 ( .A(n18786), .B(n29363), .Z(n18578) );
  NANDN U19377 ( .A(n18576), .B(n29864), .Z(n18577) );
  NAND U19378 ( .A(n18578), .B(n18577), .Z(n18851) );
  XNOR U19379 ( .A(a[91]), .B(n967), .Z(n18789) );
  NAND U19380 ( .A(n18789), .B(n28939), .Z(n18581) );
  NAND U19381 ( .A(n28938), .B(n18579), .Z(n18580) );
  AND U19382 ( .A(n18581), .B(n18580), .Z(n18852) );
  XNOR U19383 ( .A(n18851), .B(n18852), .Z(n18853) );
  XNOR U19384 ( .A(n18854), .B(n18853), .Z(n18752) );
  XNOR U19385 ( .A(a[81]), .B(b[13]), .Z(n18774) );
  OR U19386 ( .A(n18774), .B(n31550), .Z(n18584) );
  NANDN U19387 ( .A(n18582), .B(n31874), .Z(n18583) );
  NAND U19388 ( .A(n18584), .B(n18583), .Z(n18939) );
  NAND U19389 ( .A(n34848), .B(n18585), .Z(n18587) );
  XOR U19390 ( .A(n35375), .B(n29372), .Z(n18777) );
  NAND U19391 ( .A(n34618), .B(n18777), .Z(n18586) );
  NAND U19392 ( .A(n18587), .B(n18586), .Z(n18936) );
  NAND U19393 ( .A(n35188), .B(n18588), .Z(n18590) );
  XOR U19394 ( .A(n35540), .B(n28403), .Z(n18780) );
  NANDN U19395 ( .A(n34968), .B(n18780), .Z(n18589) );
  AND U19396 ( .A(n18590), .B(n18589), .Z(n18937) );
  XNOR U19397 ( .A(n18936), .B(n18937), .Z(n18938) );
  XOR U19398 ( .A(n18939), .B(n18938), .Z(n18753) );
  XOR U19399 ( .A(n18752), .B(n18753), .Z(n18755) );
  NANDN U19400 ( .A(n18592), .B(n18591), .Z(n18596) );
  NAND U19401 ( .A(n18594), .B(n18593), .Z(n18595) );
  NAND U19402 ( .A(n18596), .B(n18595), .Z(n18754) );
  XNOR U19403 ( .A(n18755), .B(n18754), .Z(n18765) );
  NANDN U19404 ( .A(n18598), .B(n18597), .Z(n18602) );
  NAND U19405 ( .A(n18600), .B(n18599), .Z(n18601) );
  NAND U19406 ( .A(n18602), .B(n18601), .Z(n18895) );
  NAND U19407 ( .A(a[29]), .B(b[63]), .Z(n18909) );
  NANDN U19408 ( .A(n18603), .B(n38369), .Z(n18605) );
  XOR U19409 ( .A(b[61]), .B(n19656), .Z(n18805) );
  OR U19410 ( .A(n18805), .B(n38371), .Z(n18604) );
  NAND U19411 ( .A(n18605), .B(n18604), .Z(n18907) );
  NANDN U19412 ( .A(n18606), .B(n35311), .Z(n18608) );
  XNOR U19413 ( .A(b[31]), .B(a[63]), .Z(n18808) );
  NANDN U19414 ( .A(n18808), .B(n35313), .Z(n18607) );
  AND U19415 ( .A(n18608), .B(n18607), .Z(n18906) );
  XNOR U19416 ( .A(n18907), .B(n18906), .Z(n18908) );
  XOR U19417 ( .A(n18909), .B(n18908), .Z(n18893) );
  NAND U19418 ( .A(n33283), .B(n18609), .Z(n18611) );
  XNOR U19419 ( .A(n33020), .B(a[75]), .Z(n18811) );
  NANDN U19420 ( .A(n33021), .B(n18811), .Z(n18610) );
  NAND U19421 ( .A(n18611), .B(n18610), .Z(n18823) );
  XOR U19422 ( .A(b[21]), .B(a[73]), .Z(n18814) );
  NANDN U19423 ( .A(n33634), .B(n18814), .Z(n18614) );
  NANDN U19424 ( .A(n18612), .B(n33464), .Z(n18613) );
  NAND U19425 ( .A(n18614), .B(n18613), .Z(n18820) );
  NAND U19426 ( .A(n34044), .B(n18615), .Z(n18617) );
  XOR U19427 ( .A(n34510), .B(n30543), .Z(n18817) );
  NANDN U19428 ( .A(n33867), .B(n18817), .Z(n18616) );
  AND U19429 ( .A(n18617), .B(n18616), .Z(n18821) );
  XNOR U19430 ( .A(n18820), .B(n18821), .Z(n18822) );
  XNOR U19431 ( .A(n18823), .B(n18822), .Z(n18894) );
  XNOR U19432 ( .A(n18893), .B(n18894), .Z(n18896) );
  XNOR U19433 ( .A(n18895), .B(n18896), .Z(n18764) );
  XNOR U19434 ( .A(n18765), .B(n18764), .Z(n18766) );
  XNOR U19435 ( .A(n18767), .B(n18766), .Z(n18866) );
  NANDN U19436 ( .A(n18619), .B(n18618), .Z(n18623) );
  NAND U19437 ( .A(n18621), .B(n18620), .Z(n18622) );
  NAND U19438 ( .A(n18623), .B(n18622), .Z(n18957) );
  XNOR U19439 ( .A(b[41]), .B(a[53]), .Z(n18826) );
  OR U19440 ( .A(n18826), .B(n36905), .Z(n18626) );
  NANDN U19441 ( .A(n18624), .B(n36807), .Z(n18625) );
  NAND U19442 ( .A(n18626), .B(n18625), .Z(n18848) );
  XOR U19443 ( .A(b[57]), .B(n20352), .Z(n18829) );
  OR U19444 ( .A(n18829), .B(n965), .Z(n18629) );
  NANDN U19445 ( .A(n18627), .B(n38194), .Z(n18628) );
  NAND U19446 ( .A(n18629), .B(n18628), .Z(n18845) );
  NAND U19447 ( .A(n38326), .B(n18630), .Z(n18632) );
  XOR U19448 ( .A(n38400), .B(n20315), .Z(n18832) );
  NANDN U19449 ( .A(n38273), .B(n18832), .Z(n18631) );
  AND U19450 ( .A(n18632), .B(n18631), .Z(n18846) );
  XNOR U19451 ( .A(n18845), .B(n18846), .Z(n18847) );
  XOR U19452 ( .A(n18848), .B(n18847), .Z(n18954) );
  XOR U19453 ( .A(b[33]), .B(n27773), .Z(n18835) );
  NANDN U19454 ( .A(n18835), .B(n35620), .Z(n18635) );
  NANDN U19455 ( .A(n18633), .B(n35621), .Z(n18634) );
  NAND U19456 ( .A(n18635), .B(n18634), .Z(n18951) );
  NANDN U19457 ( .A(n966), .B(a[93]), .Z(n18636) );
  XOR U19458 ( .A(n29232), .B(n18636), .Z(n18638) );
  IV U19459 ( .A(a[92]), .Z(n34852) );
  NANDN U19460 ( .A(n34852), .B(n966), .Z(n18637) );
  AND U19461 ( .A(n18638), .B(n18637), .Z(n18948) );
  XOR U19462 ( .A(b[63]), .B(n18639), .Z(n18842) );
  NANDN U19463 ( .A(n18842), .B(n38422), .Z(n18642) );
  NANDN U19464 ( .A(n18640), .B(n38423), .Z(n18641) );
  AND U19465 ( .A(n18642), .B(n18641), .Z(n18949) );
  XNOR U19466 ( .A(n18948), .B(n18949), .Z(n18950) );
  XOR U19467 ( .A(n18951), .B(n18950), .Z(n18955) );
  XNOR U19468 ( .A(n18954), .B(n18955), .Z(n18956) );
  XNOR U19469 ( .A(n18957), .B(n18956), .Z(n18761) );
  NANDN U19470 ( .A(n18644), .B(n18643), .Z(n18648) );
  NAND U19471 ( .A(n18646), .B(n18645), .Z(n18647) );
  NAND U19472 ( .A(n18648), .B(n18647), .Z(n18758) );
  NANDN U19473 ( .A(n18650), .B(n18649), .Z(n18654) );
  NAND U19474 ( .A(n18652), .B(n18651), .Z(n18653) );
  AND U19475 ( .A(n18654), .B(n18653), .Z(n18759) );
  XNOR U19476 ( .A(n18758), .B(n18759), .Z(n18760) );
  XOR U19477 ( .A(n18761), .B(n18760), .Z(n18864) );
  XOR U19478 ( .A(n18864), .B(n18863), .Z(n18865) );
  XOR U19479 ( .A(n18866), .B(n18865), .Z(n18968) );
  XNOR U19480 ( .A(n18969), .B(n18968), .Z(n18742) );
  XOR U19481 ( .A(n18743), .B(n18742), .Z(n18744) );
  XNOR U19482 ( .A(n18745), .B(n18744), .Z(n18732) );
  NAND U19483 ( .A(n18660), .B(n18659), .Z(n18664) );
  NAND U19484 ( .A(n18662), .B(n18661), .Z(n18663) );
  NAND U19485 ( .A(n18664), .B(n18663), .Z(n18739) );
  NANDN U19486 ( .A(n18666), .B(n18665), .Z(n18670) );
  NANDN U19487 ( .A(n18668), .B(n18667), .Z(n18669) );
  NAND U19488 ( .A(n18670), .B(n18669), .Z(n18736) );
  NANDN U19489 ( .A(n18672), .B(n18671), .Z(n18676) );
  NAND U19490 ( .A(n18674), .B(n18673), .Z(n18675) );
  AND U19491 ( .A(n18676), .B(n18675), .Z(n18737) );
  XNOR U19492 ( .A(n18736), .B(n18737), .Z(n18738) );
  XNOR U19493 ( .A(n18739), .B(n18738), .Z(n18730) );
  NANDN U19494 ( .A(n18678), .B(n18677), .Z(n18682) );
  NAND U19495 ( .A(n18680), .B(n18679), .Z(n18681) );
  NAND U19496 ( .A(n18682), .B(n18681), .Z(n18731) );
  XOR U19497 ( .A(n18730), .B(n18731), .Z(n18733) );
  XNOR U19498 ( .A(n18732), .B(n18733), .Z(n18727) );
  NANDN U19499 ( .A(n18684), .B(n18683), .Z(n18688) );
  NANDN U19500 ( .A(n18686), .B(n18685), .Z(n18687) );
  NAND U19501 ( .A(n18688), .B(n18687), .Z(n18725) );
  NANDN U19502 ( .A(n18690), .B(n18689), .Z(n18694) );
  NANDN U19503 ( .A(n18692), .B(n18691), .Z(n18693) );
  AND U19504 ( .A(n18694), .B(n18693), .Z(n18724) );
  XNOR U19505 ( .A(n18725), .B(n18724), .Z(n18726) );
  XNOR U19506 ( .A(n18727), .B(n18726), .Z(n18997) );
  OR U19507 ( .A(n18696), .B(n18695), .Z(n18700) );
  NAND U19508 ( .A(n18698), .B(n18697), .Z(n18699) );
  NAND U19509 ( .A(n18700), .B(n18699), .Z(n18995) );
  NANDN U19510 ( .A(n18702), .B(n18701), .Z(n18706) );
  NANDN U19511 ( .A(n18704), .B(n18703), .Z(n18705) );
  AND U19512 ( .A(n18706), .B(n18705), .Z(n18994) );
  XNOR U19513 ( .A(n18995), .B(n18994), .Z(n18996) );
  XNOR U19514 ( .A(n18997), .B(n18996), .Z(n18718) );
  NANDN U19515 ( .A(n18708), .B(n18707), .Z(n18712) );
  NAND U19516 ( .A(n18710), .B(n18709), .Z(n18711) );
  NAND U19517 ( .A(n18712), .B(n18711), .Z(n18719) );
  XOR U19518 ( .A(n18718), .B(n18719), .Z(n18720) );
  XNOR U19519 ( .A(n18721), .B(n18720), .Z(n19000) );
  XNOR U19520 ( .A(n19000), .B(sreg[157]), .Z(n19002) );
  NAND U19521 ( .A(n18713), .B(sreg[156]), .Z(n18717) );
  OR U19522 ( .A(n18715), .B(n18714), .Z(n18716) );
  AND U19523 ( .A(n18717), .B(n18716), .Z(n19001) );
  XOR U19524 ( .A(n19002), .B(n19001), .Z(c[157]) );
  OR U19525 ( .A(n18719), .B(n18718), .Z(n18723) );
  NAND U19526 ( .A(n18721), .B(n18720), .Z(n18722) );
  NAND U19527 ( .A(n18723), .B(n18722), .Z(n19008) );
  NANDN U19528 ( .A(n18725), .B(n18724), .Z(n18729) );
  NANDN U19529 ( .A(n18727), .B(n18726), .Z(n18728) );
  NAND U19530 ( .A(n18729), .B(n18728), .Z(n19283) );
  NANDN U19531 ( .A(n18731), .B(n18730), .Z(n18735) );
  NANDN U19532 ( .A(n18733), .B(n18732), .Z(n18734) );
  NAND U19533 ( .A(n18735), .B(n18734), .Z(n19284) );
  XNOR U19534 ( .A(n19283), .B(n19284), .Z(n19285) );
  NANDN U19535 ( .A(n18737), .B(n18736), .Z(n18741) );
  NAND U19536 ( .A(n18739), .B(n18738), .Z(n18740) );
  NAND U19537 ( .A(n18741), .B(n18740), .Z(n19277) );
  XNOR U19538 ( .A(n19277), .B(n19278), .Z(n19279) );
  NANDN U19539 ( .A(n18747), .B(n18746), .Z(n18751) );
  NAND U19540 ( .A(n18749), .B(n18748), .Z(n18750) );
  AND U19541 ( .A(n18751), .B(n18750), .Z(n19264) );
  NANDN U19542 ( .A(n18753), .B(n18752), .Z(n18757) );
  OR U19543 ( .A(n18755), .B(n18754), .Z(n18756) );
  NAND U19544 ( .A(n18757), .B(n18756), .Z(n19261) );
  NANDN U19545 ( .A(n18759), .B(n18758), .Z(n18763) );
  NAND U19546 ( .A(n18761), .B(n18760), .Z(n18762) );
  NAND U19547 ( .A(n18763), .B(n18762), .Z(n19262) );
  XNOR U19548 ( .A(n19261), .B(n19262), .Z(n19263) );
  XNOR U19549 ( .A(n19264), .B(n19263), .Z(n19245) );
  NAND U19550 ( .A(n18765), .B(n18764), .Z(n18769) );
  OR U19551 ( .A(n18767), .B(n18766), .Z(n18768) );
  AND U19552 ( .A(n18769), .B(n18768), .Z(n19246) );
  XNOR U19553 ( .A(n19245), .B(n19246), .Z(n19248) );
  XOR U19554 ( .A(a[82]), .B(n971), .Z(n19062) );
  OR U19555 ( .A(n19062), .B(n31550), .Z(n18776) );
  NANDN U19556 ( .A(n18774), .B(n31874), .Z(n18775) );
  NAND U19557 ( .A(n18776), .B(n18775), .Z(n19218) );
  NAND U19558 ( .A(n34848), .B(n18777), .Z(n18779) );
  XOR U19559 ( .A(n35375), .B(n29868), .Z(n19065) );
  NAND U19560 ( .A(n34618), .B(n19065), .Z(n18778) );
  NAND U19561 ( .A(n18779), .B(n18778), .Z(n19215) );
  NAND U19562 ( .A(n35188), .B(n18780), .Z(n18782) );
  XOR U19563 ( .A(n35540), .B(n28701), .Z(n19068) );
  NANDN U19564 ( .A(n34968), .B(n19068), .Z(n18781) );
  AND U19565 ( .A(n18782), .B(n18781), .Z(n19216) );
  XNOR U19566 ( .A(n19215), .B(n19216), .Z(n19217) );
  XNOR U19567 ( .A(n19218), .B(n19217), .Z(n19025) );
  XOR U19568 ( .A(b[37]), .B(n26347), .Z(n19053) );
  NANDN U19569 ( .A(n19053), .B(n36311), .Z(n18785) );
  NANDN U19570 ( .A(n18783), .B(n36309), .Z(n18784) );
  NAND U19571 ( .A(n18785), .B(n18784), .Z(n19131) );
  XOR U19572 ( .A(a[90]), .B(n968), .Z(n19056) );
  OR U19573 ( .A(n19056), .B(n29363), .Z(n18788) );
  NANDN U19574 ( .A(n18786), .B(n29864), .Z(n18787) );
  NAND U19575 ( .A(n18788), .B(n18787), .Z(n19128) );
  XOR U19576 ( .A(n34852), .B(n967), .Z(n19059) );
  NAND U19577 ( .A(n19059), .B(n28939), .Z(n18791) );
  NAND U19578 ( .A(n28938), .B(n18789), .Z(n18790) );
  AND U19579 ( .A(n18791), .B(n18790), .Z(n19129) );
  XNOR U19580 ( .A(n19128), .B(n19129), .Z(n19130) );
  XNOR U19581 ( .A(n19131), .B(n19130), .Z(n19023) );
  NANDN U19582 ( .A(n18793), .B(n18792), .Z(n18797) );
  NAND U19583 ( .A(n18795), .B(n18794), .Z(n18796) );
  NAND U19584 ( .A(n18797), .B(n18796), .Z(n19024) );
  XOR U19585 ( .A(n19023), .B(n19024), .Z(n19026) );
  XNOR U19586 ( .A(n19025), .B(n19026), .Z(n19041) );
  NANDN U19587 ( .A(n18799), .B(n18798), .Z(n18803) );
  NAND U19588 ( .A(n18801), .B(n18800), .Z(n18802) );
  NAND U19589 ( .A(n18803), .B(n18802), .Z(n19172) );
  ANDN U19590 ( .B(b[63]), .A(n18804), .Z(n19188) );
  NANDN U19591 ( .A(n18805), .B(n38369), .Z(n18807) );
  XOR U19592 ( .A(b[61]), .B(n19513), .Z(n19083) );
  OR U19593 ( .A(n19083), .B(n38371), .Z(n18806) );
  NAND U19594 ( .A(n18807), .B(n18806), .Z(n19186) );
  NANDN U19595 ( .A(n18808), .B(n35311), .Z(n18810) );
  XNOR U19596 ( .A(b[31]), .B(a[64]), .Z(n19086) );
  NANDN U19597 ( .A(n19086), .B(n35313), .Z(n18809) );
  AND U19598 ( .A(n18810), .B(n18809), .Z(n19185) );
  XNOR U19599 ( .A(n19186), .B(n19185), .Z(n19187) );
  XOR U19600 ( .A(n19188), .B(n19187), .Z(n19170) );
  NAND U19601 ( .A(n33283), .B(n18811), .Z(n18813) );
  XOR U19602 ( .A(n33020), .B(n31363), .Z(n19089) );
  NANDN U19603 ( .A(n33021), .B(n19089), .Z(n18812) );
  NAND U19604 ( .A(n18813), .B(n18812), .Z(n19119) );
  XNOR U19605 ( .A(b[21]), .B(a[74]), .Z(n19092) );
  OR U19606 ( .A(n19092), .B(n33634), .Z(n18816) );
  NAND U19607 ( .A(n18814), .B(n33464), .Z(n18815) );
  NAND U19608 ( .A(n18816), .B(n18815), .Z(n19116) );
  NAND U19609 ( .A(n34044), .B(n18817), .Z(n18819) );
  XOR U19610 ( .A(n34510), .B(n30210), .Z(n19095) );
  NANDN U19611 ( .A(n33867), .B(n19095), .Z(n18818) );
  AND U19612 ( .A(n18819), .B(n18818), .Z(n19117) );
  XNOR U19613 ( .A(n19116), .B(n19117), .Z(n19118) );
  XNOR U19614 ( .A(n19119), .B(n19118), .Z(n19171) );
  XOR U19615 ( .A(n19170), .B(n19171), .Z(n19173) );
  XOR U19616 ( .A(n19172), .B(n19173), .Z(n19042) );
  XOR U19617 ( .A(n19041), .B(n19042), .Z(n19043) );
  XOR U19618 ( .A(n19044), .B(n19043), .Z(n19143) );
  NANDN U19619 ( .A(n18821), .B(n18820), .Z(n18825) );
  NAND U19620 ( .A(n18823), .B(n18822), .Z(n18824) );
  NAND U19621 ( .A(n18825), .B(n18824), .Z(n19236) );
  XNOR U19622 ( .A(b[41]), .B(a[54]), .Z(n19098) );
  OR U19623 ( .A(n19098), .B(n36905), .Z(n18828) );
  NANDN U19624 ( .A(n18826), .B(n36807), .Z(n18827) );
  NAND U19625 ( .A(n18828), .B(n18827), .Z(n19125) );
  XOR U19626 ( .A(b[57]), .B(n20686), .Z(n19101) );
  OR U19627 ( .A(n19101), .B(n965), .Z(n18831) );
  NANDN U19628 ( .A(n18829), .B(n38194), .Z(n18830) );
  NAND U19629 ( .A(n18831), .B(n18830), .Z(n19122) );
  NAND U19630 ( .A(n38326), .B(n18832), .Z(n18834) );
  XOR U19631 ( .A(n38400), .B(n19980), .Z(n19104) );
  NANDN U19632 ( .A(n38273), .B(n19104), .Z(n18833) );
  AND U19633 ( .A(n18834), .B(n18833), .Z(n19123) );
  XNOR U19634 ( .A(n19122), .B(n19123), .Z(n19124) );
  XNOR U19635 ( .A(n19125), .B(n19124), .Z(n19233) );
  XNOR U19636 ( .A(b[33]), .B(a[62]), .Z(n19107) );
  NANDN U19637 ( .A(n19107), .B(n35620), .Z(n18837) );
  NANDN U19638 ( .A(n18835), .B(n35621), .Z(n18836) );
  NAND U19639 ( .A(n18837), .B(n18836), .Z(n19230) );
  NANDN U19640 ( .A(n966), .B(a[94]), .Z(n18838) );
  XOR U19641 ( .A(n29232), .B(n18838), .Z(n18840) );
  IV U19642 ( .A(a[93]), .Z(n35377) );
  NANDN U19643 ( .A(n35377), .B(n966), .Z(n18839) );
  AND U19644 ( .A(n18840), .B(n18839), .Z(n19227) );
  XOR U19645 ( .A(b[63]), .B(n18841), .Z(n19113) );
  NANDN U19646 ( .A(n19113), .B(n38422), .Z(n18844) );
  NANDN U19647 ( .A(n18842), .B(n38423), .Z(n18843) );
  AND U19648 ( .A(n18844), .B(n18843), .Z(n19228) );
  XNOR U19649 ( .A(n19227), .B(n19228), .Z(n19229) );
  XOR U19650 ( .A(n19230), .B(n19229), .Z(n19234) );
  XNOR U19651 ( .A(n19233), .B(n19234), .Z(n19235) );
  XOR U19652 ( .A(n19236), .B(n19235), .Z(n19038) );
  NANDN U19653 ( .A(n18846), .B(n18845), .Z(n18850) );
  NAND U19654 ( .A(n18848), .B(n18847), .Z(n18849) );
  NAND U19655 ( .A(n18850), .B(n18849), .Z(n19035) );
  NANDN U19656 ( .A(n18852), .B(n18851), .Z(n18856) );
  NAND U19657 ( .A(n18854), .B(n18853), .Z(n18855) );
  AND U19658 ( .A(n18856), .B(n18855), .Z(n19036) );
  XNOR U19659 ( .A(n19035), .B(n19036), .Z(n19037) );
  XNOR U19660 ( .A(n19038), .B(n19037), .Z(n19140) );
  NANDN U19661 ( .A(n18858), .B(n18857), .Z(n18862) );
  OR U19662 ( .A(n18860), .B(n18859), .Z(n18861) );
  AND U19663 ( .A(n18862), .B(n18861), .Z(n19141) );
  XNOR U19664 ( .A(n19140), .B(n19141), .Z(n19142) );
  XNOR U19665 ( .A(n19143), .B(n19142), .Z(n19247) );
  XNOR U19666 ( .A(n19248), .B(n19247), .Z(n19017) );
  OR U19667 ( .A(n18864), .B(n18863), .Z(n18868) );
  NAND U19668 ( .A(n18866), .B(n18865), .Z(n18867) );
  NAND U19669 ( .A(n18868), .B(n18867), .Z(n19268) );
  XOR U19670 ( .A(a[84]), .B(n970), .Z(n19146) );
  OR U19671 ( .A(n19146), .B(n31369), .Z(n18871) );
  NANDN U19672 ( .A(n18869), .B(n31119), .Z(n18870) );
  NAND U19673 ( .A(n18871), .B(n18870), .Z(n19167) );
  XOR U19674 ( .A(b[43]), .B(n25134), .Z(n19149) );
  NANDN U19675 ( .A(n19149), .B(n37068), .Z(n18874) );
  NANDN U19676 ( .A(n18872), .B(n37069), .Z(n18873) );
  NAND U19677 ( .A(n18874), .B(n18873), .Z(n19164) );
  XNOR U19678 ( .A(b[45]), .B(a[50]), .Z(n19152) );
  NANDN U19679 ( .A(n19152), .B(n37261), .Z(n18877) );
  NANDN U19680 ( .A(n18875), .B(n37262), .Z(n18876) );
  AND U19681 ( .A(n18877), .B(n18876), .Z(n19165) );
  XNOR U19682 ( .A(n19164), .B(n19165), .Z(n19166) );
  XNOR U19683 ( .A(n19167), .B(n19166), .Z(n19047) );
  XOR U19684 ( .A(n979), .B(n22964), .Z(n19155) );
  NANDN U19685 ( .A(n37756), .B(n19155), .Z(n18880) );
  NANDN U19686 ( .A(n18878), .B(n37652), .Z(n18879) );
  NAND U19687 ( .A(n18880), .B(n18879), .Z(n19194) );
  NAND U19688 ( .A(n37469), .B(n18881), .Z(n18883) );
  XOR U19689 ( .A(b[47]), .B(n23447), .Z(n19158) );
  NANDN U19690 ( .A(n19158), .B(n37471), .Z(n18882) );
  NAND U19691 ( .A(n18883), .B(n18882), .Z(n19191) );
  XOR U19692 ( .A(n33628), .B(n969), .Z(n19161) );
  NAND U19693 ( .A(n30509), .B(n19161), .Z(n18886) );
  NANDN U19694 ( .A(n18884), .B(n30846), .Z(n18885) );
  AND U19695 ( .A(n18886), .B(n18885), .Z(n19192) );
  XNOR U19696 ( .A(n19191), .B(n19192), .Z(n19193) );
  XOR U19697 ( .A(n19194), .B(n19193), .Z(n19048) );
  XNOR U19698 ( .A(n19047), .B(n19048), .Z(n19049) );
  NANDN U19699 ( .A(n18888), .B(n18887), .Z(n18892) );
  NAND U19700 ( .A(n18890), .B(n18889), .Z(n18891) );
  AND U19701 ( .A(n18892), .B(n18891), .Z(n19050) );
  XNOR U19702 ( .A(n19049), .B(n19050), .Z(n19252) );
  XNOR U19703 ( .A(n19252), .B(n19251), .Z(n19253) );
  XNOR U19704 ( .A(b[35]), .B(a[60]), .Z(n19176) );
  NANDN U19705 ( .A(n19176), .B(n35985), .Z(n18899) );
  NAND U19706 ( .A(n18897), .B(n35986), .Z(n18898) );
  NAND U19707 ( .A(n18899), .B(n18898), .Z(n19224) );
  XOR U19708 ( .A(n34048), .B(n31123), .Z(n19179) );
  NAND U19709 ( .A(n19179), .B(n29949), .Z(n18902) );
  NAND U19710 ( .A(n29948), .B(n18900), .Z(n18901) );
  NAND U19711 ( .A(n18902), .B(n18901), .Z(n19221) );
  XOR U19712 ( .A(b[55]), .B(n21149), .Z(n19182) );
  NANDN U19713 ( .A(n19182), .B(n38075), .Z(n18905) );
  NANDN U19714 ( .A(n18903), .B(n38073), .Z(n18904) );
  AND U19715 ( .A(n18905), .B(n18904), .Z(n19222) );
  XNOR U19716 ( .A(n19221), .B(n19222), .Z(n19223) );
  XNOR U19717 ( .A(n19224), .B(n19223), .Z(n19032) );
  NANDN U19718 ( .A(n18907), .B(n18906), .Z(n18911) );
  NAND U19719 ( .A(n18909), .B(n18908), .Z(n18910) );
  NAND U19720 ( .A(n18911), .B(n18910), .Z(n19029) );
  OR U19721 ( .A(n18913), .B(n18912), .Z(n18917) );
  NANDN U19722 ( .A(n18915), .B(n18914), .Z(n18916) );
  NAND U19723 ( .A(n18917), .B(n18916), .Z(n19030) );
  XNOR U19724 ( .A(n19029), .B(n19030), .Z(n19031) );
  XOR U19725 ( .A(n19032), .B(n19031), .Z(n19254) );
  XOR U19726 ( .A(n19253), .B(n19254), .Z(n19265) );
  XOR U19727 ( .A(a[80]), .B(n972), .Z(n19206) );
  OR U19728 ( .A(n19206), .B(n32010), .Z(n18920) );
  NANDN U19729 ( .A(n18918), .B(n32011), .Z(n18919) );
  NAND U19730 ( .A(n18920), .B(n18919), .Z(n19080) );
  XNOR U19731 ( .A(b[25]), .B(n30379), .Z(n19209) );
  NANDN U19732 ( .A(n34219), .B(n19209), .Z(n18923) );
  NAND U19733 ( .A(n34217), .B(n18921), .Z(n18922) );
  NAND U19734 ( .A(n18923), .B(n18922), .Z(n19077) );
  XNOR U19735 ( .A(b[17]), .B(a[78]), .Z(n19212) );
  NANDN U19736 ( .A(n19212), .B(n32543), .Z(n18926) );
  NAND U19737 ( .A(n18924), .B(n32541), .Z(n18925) );
  AND U19738 ( .A(n18926), .B(n18925), .Z(n19078) );
  XNOR U19739 ( .A(n19077), .B(n19078), .Z(n19079) );
  XNOR U19740 ( .A(n19080), .B(n19079), .Z(n19134) );
  XOR U19741 ( .A(b[39]), .B(n25860), .Z(n19197) );
  NANDN U19742 ( .A(n19197), .B(n36553), .Z(n18929) );
  NANDN U19743 ( .A(n18927), .B(n36643), .Z(n18928) );
  NAND U19744 ( .A(n18929), .B(n18928), .Z(n19074) );
  XOR U19745 ( .A(b[51]), .B(n22289), .Z(n19200) );
  NANDN U19746 ( .A(n19200), .B(n37803), .Z(n18932) );
  NANDN U19747 ( .A(n18930), .B(n37802), .Z(n18931) );
  NAND U19748 ( .A(n18932), .B(n18931), .Z(n19071) );
  XOR U19749 ( .A(b[53]), .B(n22246), .Z(n19203) );
  NANDN U19750 ( .A(n19203), .B(n37940), .Z(n18935) );
  NANDN U19751 ( .A(n18933), .B(n37941), .Z(n18934) );
  AND U19752 ( .A(n18935), .B(n18934), .Z(n19072) );
  XNOR U19753 ( .A(n19071), .B(n19072), .Z(n19073) );
  XOR U19754 ( .A(n19074), .B(n19073), .Z(n19135) );
  XOR U19755 ( .A(n19134), .B(n19135), .Z(n19137) );
  NANDN U19756 ( .A(n18937), .B(n18936), .Z(n18941) );
  NAND U19757 ( .A(n18939), .B(n18938), .Z(n18940) );
  NAND U19758 ( .A(n18941), .B(n18940), .Z(n19136) );
  XNOR U19759 ( .A(n19137), .B(n19136), .Z(n19242) );
  NANDN U19760 ( .A(n18943), .B(n18942), .Z(n18947) );
  NAND U19761 ( .A(n18945), .B(n18944), .Z(n18946) );
  NAND U19762 ( .A(n18947), .B(n18946), .Z(n19239) );
  NANDN U19763 ( .A(n18949), .B(n18948), .Z(n18953) );
  NAND U19764 ( .A(n18951), .B(n18950), .Z(n18952) );
  AND U19765 ( .A(n18953), .B(n18952), .Z(n19240) );
  XNOR U19766 ( .A(n19239), .B(n19240), .Z(n19241) );
  XNOR U19767 ( .A(n19242), .B(n19241), .Z(n19257) );
  OR U19768 ( .A(n18955), .B(n18954), .Z(n18959) );
  OR U19769 ( .A(n18957), .B(n18956), .Z(n18958) );
  AND U19770 ( .A(n18959), .B(n18958), .Z(n19258) );
  XNOR U19771 ( .A(n19257), .B(n19258), .Z(n19259) );
  NANDN U19772 ( .A(n18961), .B(n18960), .Z(n18965) );
  NAND U19773 ( .A(n18963), .B(n18962), .Z(n18964) );
  AND U19774 ( .A(n18965), .B(n18964), .Z(n19260) );
  XNOR U19775 ( .A(n19259), .B(n19260), .Z(n19266) );
  XNOR U19776 ( .A(n19265), .B(n19266), .Z(n19267) );
  XOR U19777 ( .A(n19268), .B(n19267), .Z(n19018) );
  XNOR U19778 ( .A(n19017), .B(n19018), .Z(n19019) );
  NAND U19779 ( .A(n18967), .B(n18966), .Z(n18971) );
  NANDN U19780 ( .A(n18969), .B(n18968), .Z(n18970) );
  NAND U19781 ( .A(n18971), .B(n18970), .Z(n19020) );
  XNOR U19782 ( .A(n19019), .B(n19020), .Z(n19273) );
  NANDN U19783 ( .A(n18973), .B(n18972), .Z(n18977) );
  NANDN U19784 ( .A(n18975), .B(n18974), .Z(n18976) );
  NAND U19785 ( .A(n18977), .B(n18976), .Z(n19272) );
  NAND U19786 ( .A(n18979), .B(n18978), .Z(n18983) );
  NANDN U19787 ( .A(n18981), .B(n18980), .Z(n18982) );
  NAND U19788 ( .A(n18983), .B(n18982), .Z(n19014) );
  NANDN U19789 ( .A(n18985), .B(n18984), .Z(n18989) );
  NAND U19790 ( .A(n18987), .B(n18986), .Z(n18988) );
  NAND U19791 ( .A(n18989), .B(n18988), .Z(n19011) );
  XNOR U19792 ( .A(n19011), .B(n19012), .Z(n19013) );
  XOR U19793 ( .A(n19014), .B(n19013), .Z(n19271) );
  XOR U19794 ( .A(n19272), .B(n19271), .Z(n19274) );
  XNOR U19795 ( .A(n19279), .B(n19280), .Z(n19286) );
  XOR U19796 ( .A(n19285), .B(n19286), .Z(n19005) );
  NANDN U19797 ( .A(n18995), .B(n18994), .Z(n18999) );
  NANDN U19798 ( .A(n18997), .B(n18996), .Z(n18998) );
  AND U19799 ( .A(n18999), .B(n18998), .Z(n19006) );
  XOR U19800 ( .A(n19005), .B(n19006), .Z(n19007) );
  XNOR U19801 ( .A(n19008), .B(n19007), .Z(n19289) );
  XNOR U19802 ( .A(n19289), .B(sreg[158]), .Z(n19291) );
  NAND U19803 ( .A(n19000), .B(sreg[157]), .Z(n19004) );
  OR U19804 ( .A(n19002), .B(n19001), .Z(n19003) );
  AND U19805 ( .A(n19004), .B(n19003), .Z(n19290) );
  XOR U19806 ( .A(n19291), .B(n19290), .Z(c[158]) );
  NAND U19807 ( .A(n19006), .B(n19005), .Z(n19010) );
  NAND U19808 ( .A(n19008), .B(n19007), .Z(n19009) );
  NAND U19809 ( .A(n19010), .B(n19009), .Z(n19297) );
  NANDN U19810 ( .A(n19012), .B(n19011), .Z(n19016) );
  NAND U19811 ( .A(n19014), .B(n19013), .Z(n19015) );
  NAND U19812 ( .A(n19016), .B(n19015), .Z(n19563) );
  NANDN U19813 ( .A(n19018), .B(n19017), .Z(n19022) );
  NANDN U19814 ( .A(n19020), .B(n19019), .Z(n19021) );
  NAND U19815 ( .A(n19022), .B(n19021), .Z(n19564) );
  XNOR U19816 ( .A(n19563), .B(n19564), .Z(n19565) );
  NANDN U19817 ( .A(n19024), .B(n19023), .Z(n19028) );
  NANDN U19818 ( .A(n19026), .B(n19025), .Z(n19027) );
  NAND U19819 ( .A(n19028), .B(n19027), .Z(n19550) );
  NANDN U19820 ( .A(n19030), .B(n19029), .Z(n19034) );
  NAND U19821 ( .A(n19032), .B(n19031), .Z(n19033) );
  AND U19822 ( .A(n19034), .B(n19033), .Z(n19547) );
  NANDN U19823 ( .A(n19036), .B(n19035), .Z(n19040) );
  NAND U19824 ( .A(n19038), .B(n19037), .Z(n19039) );
  NAND U19825 ( .A(n19040), .B(n19039), .Z(n19548) );
  XNOR U19826 ( .A(n19550), .B(n19549), .Z(n19311) );
  OR U19827 ( .A(n19042), .B(n19041), .Z(n19046) );
  NANDN U19828 ( .A(n19044), .B(n19043), .Z(n19045) );
  AND U19829 ( .A(n19046), .B(n19045), .Z(n19310) );
  XNOR U19830 ( .A(n19311), .B(n19310), .Z(n19312) );
  NANDN U19831 ( .A(n19048), .B(n19047), .Z(n19052) );
  NAND U19832 ( .A(n19050), .B(n19049), .Z(n19051) );
  NAND U19833 ( .A(n19052), .B(n19051), .Z(n19438) );
  XNOR U19834 ( .A(b[37]), .B(a[59]), .Z(n19447) );
  NANDN U19835 ( .A(n19447), .B(n36311), .Z(n19055) );
  NANDN U19836 ( .A(n19053), .B(n36309), .Z(n19054) );
  NAND U19837 ( .A(n19055), .B(n19054), .Z(n19526) );
  XNOR U19838 ( .A(a[91]), .B(b[5]), .Z(n19450) );
  OR U19839 ( .A(n19450), .B(n29363), .Z(n19058) );
  NANDN U19840 ( .A(n19056), .B(n29864), .Z(n19057) );
  NAND U19841 ( .A(n19058), .B(n19057), .Z(n19523) );
  XOR U19842 ( .A(n35377), .B(n967), .Z(n19453) );
  NAND U19843 ( .A(n19453), .B(n28939), .Z(n19061) );
  NAND U19844 ( .A(n28938), .B(n19059), .Z(n19060) );
  AND U19845 ( .A(n19061), .B(n19060), .Z(n19524) );
  XNOR U19846 ( .A(n19523), .B(n19524), .Z(n19525) );
  XNOR U19847 ( .A(n19526), .B(n19525), .Z(n19423) );
  XNOR U19848 ( .A(a[83]), .B(b[13]), .Z(n19456) );
  OR U19849 ( .A(n19456), .B(n31550), .Z(n19064) );
  NANDN U19850 ( .A(n19062), .B(n31874), .Z(n19063) );
  NAND U19851 ( .A(n19064), .B(n19063), .Z(n19337) );
  NAND U19852 ( .A(n34848), .B(n19065), .Z(n19067) );
  XNOR U19853 ( .A(n35375), .B(a[69]), .Z(n19459) );
  NAND U19854 ( .A(n34618), .B(n19459), .Z(n19066) );
  NAND U19855 ( .A(n19067), .B(n19066), .Z(n19334) );
  NAND U19856 ( .A(n35188), .B(n19068), .Z(n19070) );
  XOR U19857 ( .A(n35540), .B(n29372), .Z(n19462) );
  NANDN U19858 ( .A(n34968), .B(n19462), .Z(n19069) );
  AND U19859 ( .A(n19070), .B(n19069), .Z(n19335) );
  XNOR U19860 ( .A(n19334), .B(n19335), .Z(n19336) );
  XOR U19861 ( .A(n19337), .B(n19336), .Z(n19424) );
  XOR U19862 ( .A(n19423), .B(n19424), .Z(n19426) );
  NANDN U19863 ( .A(n19072), .B(n19071), .Z(n19076) );
  NAND U19864 ( .A(n19074), .B(n19073), .Z(n19075) );
  NAND U19865 ( .A(n19076), .B(n19075), .Z(n19425) );
  XNOR U19866 ( .A(n19426), .B(n19425), .Z(n19436) );
  NANDN U19867 ( .A(n19078), .B(n19077), .Z(n19082) );
  NAND U19868 ( .A(n19080), .B(n19079), .Z(n19081) );
  NAND U19869 ( .A(n19082), .B(n19081), .Z(n19409) );
  NAND U19870 ( .A(a[31]), .B(b[63]), .Z(n19376) );
  NANDN U19871 ( .A(n19083), .B(n38369), .Z(n19085) );
  XOR U19872 ( .A(b[61]), .B(n20315), .Z(n19477) );
  OR U19873 ( .A(n19477), .B(n38371), .Z(n19084) );
  NAND U19874 ( .A(n19085), .B(n19084), .Z(n19374) );
  NANDN U19875 ( .A(n19086), .B(n35311), .Z(n19088) );
  XOR U19876 ( .A(b[31]), .B(n28403), .Z(n19480) );
  NANDN U19877 ( .A(n19480), .B(n35313), .Z(n19087) );
  AND U19878 ( .A(n19088), .B(n19087), .Z(n19373) );
  XNOR U19879 ( .A(n19374), .B(n19373), .Z(n19375) );
  XOR U19880 ( .A(n19376), .B(n19375), .Z(n19407) );
  NAND U19881 ( .A(n33283), .B(n19089), .Z(n19091) );
  XNOR U19882 ( .A(n33020), .B(a[77]), .Z(n19483) );
  NANDN U19883 ( .A(n33021), .B(n19483), .Z(n19090) );
  NAND U19884 ( .A(n19091), .B(n19090), .Z(n19495) );
  XOR U19885 ( .A(b[21]), .B(a[75]), .Z(n19486) );
  NANDN U19886 ( .A(n33634), .B(n19486), .Z(n19094) );
  NANDN U19887 ( .A(n19092), .B(n33464), .Z(n19093) );
  NAND U19888 ( .A(n19094), .B(n19093), .Z(n19492) );
  NAND U19889 ( .A(n34044), .B(n19095), .Z(n19097) );
  XNOR U19890 ( .A(n34510), .B(a[73]), .Z(n19489) );
  NANDN U19891 ( .A(n33867), .B(n19489), .Z(n19096) );
  AND U19892 ( .A(n19097), .B(n19096), .Z(n19493) );
  XNOR U19893 ( .A(n19492), .B(n19493), .Z(n19494) );
  XNOR U19894 ( .A(n19495), .B(n19494), .Z(n19408) );
  XNOR U19895 ( .A(n19407), .B(n19408), .Z(n19410) );
  XNOR U19896 ( .A(n19409), .B(n19410), .Z(n19435) );
  XNOR U19897 ( .A(n19436), .B(n19435), .Z(n19437) );
  XNOR U19898 ( .A(n19438), .B(n19437), .Z(n19414) );
  XNOR U19899 ( .A(b[41]), .B(a[55]), .Z(n19498) );
  OR U19900 ( .A(n19498), .B(n36905), .Z(n19100) );
  NANDN U19901 ( .A(n19098), .B(n36807), .Z(n19099) );
  NAND U19902 ( .A(n19100), .B(n19099), .Z(n19520) );
  XOR U19903 ( .A(b[57]), .B(n20867), .Z(n19501) );
  OR U19904 ( .A(n19501), .B(n965), .Z(n19103) );
  NANDN U19905 ( .A(n19101), .B(n38194), .Z(n19102) );
  NAND U19906 ( .A(n19103), .B(n19102), .Z(n19517) );
  NAND U19907 ( .A(n38326), .B(n19104), .Z(n19106) );
  XOR U19908 ( .A(n38400), .B(n20352), .Z(n19504) );
  NANDN U19909 ( .A(n38273), .B(n19504), .Z(n19105) );
  AND U19910 ( .A(n19106), .B(n19105), .Z(n19518) );
  XNOR U19911 ( .A(n19517), .B(n19518), .Z(n19519) );
  XOR U19912 ( .A(n19520), .B(n19519), .Z(n19352) );
  XNOR U19913 ( .A(b[33]), .B(a[63]), .Z(n19507) );
  NANDN U19914 ( .A(n19507), .B(n35620), .Z(n19109) );
  NANDN U19915 ( .A(n19107), .B(n35621), .Z(n19108) );
  NAND U19916 ( .A(n19109), .B(n19108), .Z(n19349) );
  NANDN U19917 ( .A(n966), .B(a[95]), .Z(n19110) );
  XOR U19918 ( .A(n29232), .B(n19110), .Z(n19112) );
  IV U19919 ( .A(a[94]), .Z(n35191) );
  NANDN U19920 ( .A(n35191), .B(n966), .Z(n19111) );
  AND U19921 ( .A(n19112), .B(n19111), .Z(n19346) );
  XOR U19922 ( .A(b[63]), .B(n19656), .Z(n19514) );
  NANDN U19923 ( .A(n19514), .B(n38422), .Z(n19115) );
  NANDN U19924 ( .A(n19113), .B(n38423), .Z(n19114) );
  AND U19925 ( .A(n19115), .B(n19114), .Z(n19347) );
  XNOR U19926 ( .A(n19346), .B(n19347), .Z(n19348) );
  XOR U19927 ( .A(n19349), .B(n19348), .Z(n19353) );
  XNOR U19928 ( .A(n19352), .B(n19353), .Z(n19355) );
  NANDN U19929 ( .A(n19117), .B(n19116), .Z(n19121) );
  NAND U19930 ( .A(n19119), .B(n19118), .Z(n19120) );
  NAND U19931 ( .A(n19121), .B(n19120), .Z(n19354) );
  XNOR U19932 ( .A(n19355), .B(n19354), .Z(n19432) );
  NANDN U19933 ( .A(n19123), .B(n19122), .Z(n19127) );
  NAND U19934 ( .A(n19125), .B(n19124), .Z(n19126) );
  NAND U19935 ( .A(n19127), .B(n19126), .Z(n19429) );
  NANDN U19936 ( .A(n19129), .B(n19128), .Z(n19133) );
  NAND U19937 ( .A(n19131), .B(n19130), .Z(n19132) );
  AND U19938 ( .A(n19133), .B(n19132), .Z(n19430) );
  XNOR U19939 ( .A(n19429), .B(n19430), .Z(n19431) );
  XOR U19940 ( .A(n19432), .B(n19431), .Z(n19412) );
  NANDN U19941 ( .A(n19135), .B(n19134), .Z(n19139) );
  OR U19942 ( .A(n19137), .B(n19136), .Z(n19138) );
  AND U19943 ( .A(n19139), .B(n19138), .Z(n19411) );
  XOR U19944 ( .A(n19412), .B(n19411), .Z(n19413) );
  XNOR U19945 ( .A(n19414), .B(n19413), .Z(n19313) );
  XOR U19946 ( .A(n19312), .B(n19313), .Z(n19298) );
  NANDN U19947 ( .A(n19141), .B(n19140), .Z(n19145) );
  NAND U19948 ( .A(n19143), .B(n19142), .Z(n19144) );
  NAND U19949 ( .A(n19145), .B(n19144), .Z(n19556) );
  XNOR U19950 ( .A(a[85]), .B(b[11]), .Z(n19383) );
  OR U19951 ( .A(n19383), .B(n31369), .Z(n19148) );
  NANDN U19952 ( .A(n19146), .B(n31119), .Z(n19147) );
  NAND U19953 ( .A(n19148), .B(n19147), .Z(n19404) );
  XOR U19954 ( .A(b[43]), .B(n25001), .Z(n19386) );
  NANDN U19955 ( .A(n19386), .B(n37068), .Z(n19151) );
  NANDN U19956 ( .A(n19149), .B(n37069), .Z(n19150) );
  NAND U19957 ( .A(n19151), .B(n19150), .Z(n19401) );
  XNOR U19958 ( .A(b[45]), .B(a[51]), .Z(n19389) );
  NANDN U19959 ( .A(n19389), .B(n37261), .Z(n19154) );
  NANDN U19960 ( .A(n19152), .B(n37262), .Z(n19153) );
  AND U19961 ( .A(n19154), .B(n19153), .Z(n19402) );
  XNOR U19962 ( .A(n19401), .B(n19402), .Z(n19403) );
  XNOR U19963 ( .A(n19404), .B(n19403), .Z(n19444) );
  NAND U19964 ( .A(n37652), .B(n19155), .Z(n19157) );
  XOR U19965 ( .A(b[49]), .B(n23149), .Z(n19392) );
  OR U19966 ( .A(n19392), .B(n37756), .Z(n19156) );
  NAND U19967 ( .A(n19157), .B(n19156), .Z(n19381) );
  NANDN U19968 ( .A(n19158), .B(n37469), .Z(n19160) );
  XNOR U19969 ( .A(n978), .B(a[49]), .Z(n19395) );
  NAND U19970 ( .A(n19395), .B(n37471), .Z(n19159) );
  NAND U19971 ( .A(n19160), .B(n19159), .Z(n19379) );
  NAND U19972 ( .A(n30846), .B(n19161), .Z(n19163) );
  XNOR U19973 ( .A(a[87]), .B(n969), .Z(n19398) );
  NAND U19974 ( .A(n30509), .B(n19398), .Z(n19162) );
  NAND U19975 ( .A(n19163), .B(n19162), .Z(n19380) );
  XNOR U19976 ( .A(n19379), .B(n19380), .Z(n19382) );
  XOR U19977 ( .A(n19381), .B(n19382), .Z(n19441) );
  NANDN U19978 ( .A(n19165), .B(n19164), .Z(n19169) );
  NAND U19979 ( .A(n19167), .B(n19166), .Z(n19168) );
  NAND U19980 ( .A(n19169), .B(n19168), .Z(n19442) );
  XNOR U19981 ( .A(n19441), .B(n19442), .Z(n19443) );
  XOR U19982 ( .A(n19444), .B(n19443), .Z(n19535) );
  NANDN U19983 ( .A(n19171), .B(n19170), .Z(n19175) );
  NANDN U19984 ( .A(n19173), .B(n19172), .Z(n19174) );
  AND U19985 ( .A(n19175), .B(n19174), .Z(n19536) );
  XNOR U19986 ( .A(n19535), .B(n19536), .Z(n19538) );
  XNOR U19987 ( .A(b[35]), .B(a[61]), .Z(n19364) );
  NANDN U19988 ( .A(n19364), .B(n35985), .Z(n19178) );
  NANDN U19989 ( .A(n19176), .B(n35986), .Z(n19177) );
  NAND U19990 ( .A(n19178), .B(n19177), .Z(n19343) );
  XNOR U19991 ( .A(a[89]), .B(n31123), .Z(n19367) );
  NAND U19992 ( .A(n19367), .B(n29949), .Z(n19181) );
  NAND U19993 ( .A(n29948), .B(n19179), .Z(n19180) );
  NAND U19994 ( .A(n19181), .B(n19180), .Z(n19340) );
  XOR U19995 ( .A(b[55]), .B(n21441), .Z(n19370) );
  NANDN U19996 ( .A(n19370), .B(n38075), .Z(n19184) );
  NANDN U19997 ( .A(n19182), .B(n38073), .Z(n19183) );
  AND U19998 ( .A(n19184), .B(n19183), .Z(n19341) );
  XNOR U19999 ( .A(n19340), .B(n19341), .Z(n19342) );
  XNOR U20000 ( .A(n19343), .B(n19342), .Z(n19420) );
  NANDN U20001 ( .A(n19186), .B(n19185), .Z(n19190) );
  NANDN U20002 ( .A(n19188), .B(n19187), .Z(n19189) );
  NAND U20003 ( .A(n19190), .B(n19189), .Z(n19417) );
  NANDN U20004 ( .A(n19192), .B(n19191), .Z(n19196) );
  NAND U20005 ( .A(n19194), .B(n19193), .Z(n19195) );
  NAND U20006 ( .A(n19196), .B(n19195), .Z(n19418) );
  XNOR U20007 ( .A(n19417), .B(n19418), .Z(n19419) );
  XOR U20008 ( .A(n19420), .B(n19419), .Z(n19537) );
  XNOR U20009 ( .A(n19538), .B(n19537), .Z(n19553) );
  XOR U20010 ( .A(b[39]), .B(n26122), .Z(n19325) );
  NANDN U20011 ( .A(n19325), .B(n36553), .Z(n19199) );
  NANDN U20012 ( .A(n19197), .B(n36643), .Z(n19198) );
  NAND U20013 ( .A(n19199), .B(n19198), .Z(n19468) );
  XOR U20014 ( .A(b[51]), .B(n22579), .Z(n19328) );
  NANDN U20015 ( .A(n19328), .B(n37803), .Z(n19202) );
  NANDN U20016 ( .A(n19200), .B(n37802), .Z(n19201) );
  NAND U20017 ( .A(n19202), .B(n19201), .Z(n19465) );
  XOR U20018 ( .A(b[53]), .B(n21996), .Z(n19331) );
  NANDN U20019 ( .A(n19331), .B(n37940), .Z(n19205) );
  NANDN U20020 ( .A(n19203), .B(n37941), .Z(n19204) );
  AND U20021 ( .A(n19205), .B(n19204), .Z(n19466) );
  XNOR U20022 ( .A(n19465), .B(n19466), .Z(n19467) );
  XNOR U20023 ( .A(n19468), .B(n19467), .Z(n19532) );
  XNOR U20024 ( .A(a[81]), .B(b[15]), .Z(n19316) );
  OR U20025 ( .A(n19316), .B(n32010), .Z(n19208) );
  NANDN U20026 ( .A(n19206), .B(n32011), .Z(n19207) );
  NAND U20027 ( .A(n19208), .B(n19207), .Z(n19474) );
  XNOR U20028 ( .A(b[25]), .B(n30543), .Z(n19319) );
  NANDN U20029 ( .A(n34219), .B(n19319), .Z(n19211) );
  NAND U20030 ( .A(n34217), .B(n19209), .Z(n19210) );
  NAND U20031 ( .A(n19211), .B(n19210), .Z(n19471) );
  XOR U20032 ( .A(b[17]), .B(a[79]), .Z(n19322) );
  NAND U20033 ( .A(n19322), .B(n32543), .Z(n19214) );
  NANDN U20034 ( .A(n19212), .B(n32541), .Z(n19213) );
  AND U20035 ( .A(n19214), .B(n19213), .Z(n19472) );
  XNOR U20036 ( .A(n19471), .B(n19472), .Z(n19473) );
  XNOR U20037 ( .A(n19474), .B(n19473), .Z(n19529) );
  NANDN U20038 ( .A(n19216), .B(n19215), .Z(n19220) );
  NAND U20039 ( .A(n19218), .B(n19217), .Z(n19219) );
  NAND U20040 ( .A(n19220), .B(n19219), .Z(n19530) );
  XNOR U20041 ( .A(n19529), .B(n19530), .Z(n19531) );
  XOR U20042 ( .A(n19532), .B(n19531), .Z(n19361) );
  NANDN U20043 ( .A(n19222), .B(n19221), .Z(n19226) );
  NAND U20044 ( .A(n19224), .B(n19223), .Z(n19225) );
  NAND U20045 ( .A(n19226), .B(n19225), .Z(n19358) );
  NANDN U20046 ( .A(n19228), .B(n19227), .Z(n19232) );
  NAND U20047 ( .A(n19230), .B(n19229), .Z(n19231) );
  AND U20048 ( .A(n19232), .B(n19231), .Z(n19359) );
  XNOR U20049 ( .A(n19358), .B(n19359), .Z(n19360) );
  XNOR U20050 ( .A(n19361), .B(n19360), .Z(n19542) );
  NANDN U20051 ( .A(n19234), .B(n19233), .Z(n19238) );
  NANDN U20052 ( .A(n19236), .B(n19235), .Z(n19237) );
  AND U20053 ( .A(n19238), .B(n19237), .Z(n19541) );
  XOR U20054 ( .A(n19542), .B(n19541), .Z(n19543) );
  NANDN U20055 ( .A(n19240), .B(n19239), .Z(n19244) );
  NAND U20056 ( .A(n19242), .B(n19241), .Z(n19243) );
  AND U20057 ( .A(n19244), .B(n19243), .Z(n19544) );
  XOR U20058 ( .A(n19543), .B(n19544), .Z(n19554) );
  XOR U20059 ( .A(n19553), .B(n19554), .Z(n19555) );
  XOR U20060 ( .A(n19556), .B(n19555), .Z(n19299) );
  XNOR U20061 ( .A(n19298), .B(n19299), .Z(n19300) );
  NAND U20062 ( .A(n19246), .B(n19245), .Z(n19250) );
  OR U20063 ( .A(n19248), .B(n19247), .Z(n19249) );
  NAND U20064 ( .A(n19250), .B(n19249), .Z(n19301) );
  XOR U20065 ( .A(n19300), .B(n19301), .Z(n19560) );
  NANDN U20066 ( .A(n19252), .B(n19251), .Z(n19256) );
  NAND U20067 ( .A(n19254), .B(n19253), .Z(n19255) );
  NAND U20068 ( .A(n19256), .B(n19255), .Z(n19307) );
  XNOR U20069 ( .A(n19305), .B(n19304), .Z(n19306) );
  XOR U20070 ( .A(n19307), .B(n19306), .Z(n19557) );
  NANDN U20071 ( .A(n19266), .B(n19265), .Z(n19270) );
  NAND U20072 ( .A(n19268), .B(n19267), .Z(n19269) );
  AND U20073 ( .A(n19270), .B(n19269), .Z(n19558) );
  XNOR U20074 ( .A(n19557), .B(n19558), .Z(n19559) );
  XNOR U20075 ( .A(n19560), .B(n19559), .Z(n19566) );
  XOR U20076 ( .A(n19565), .B(n19566), .Z(n19572) );
  NANDN U20077 ( .A(n19272), .B(n19271), .Z(n19276) );
  OR U20078 ( .A(n19274), .B(n19273), .Z(n19275) );
  NAND U20079 ( .A(n19276), .B(n19275), .Z(n19570) );
  NANDN U20080 ( .A(n19278), .B(n19277), .Z(n19282) );
  NANDN U20081 ( .A(n19280), .B(n19279), .Z(n19281) );
  AND U20082 ( .A(n19282), .B(n19281), .Z(n19569) );
  XNOR U20083 ( .A(n19570), .B(n19569), .Z(n19571) );
  XNOR U20084 ( .A(n19572), .B(n19571), .Z(n19294) );
  NANDN U20085 ( .A(n19284), .B(n19283), .Z(n19288) );
  NAND U20086 ( .A(n19286), .B(n19285), .Z(n19287) );
  AND U20087 ( .A(n19288), .B(n19287), .Z(n19295) );
  XNOR U20088 ( .A(n19294), .B(n19295), .Z(n19296) );
  XNOR U20089 ( .A(n19297), .B(n19296), .Z(n19575) );
  XNOR U20090 ( .A(n19575), .B(sreg[159]), .Z(n19577) );
  NAND U20091 ( .A(n19289), .B(sreg[158]), .Z(n19293) );
  OR U20092 ( .A(n19291), .B(n19290), .Z(n19292) );
  AND U20093 ( .A(n19293), .B(n19292), .Z(n19576) );
  XOR U20094 ( .A(n19577), .B(n19576), .Z(c[159]) );
  NANDN U20095 ( .A(n19299), .B(n19298), .Z(n19303) );
  NANDN U20096 ( .A(n19301), .B(n19300), .Z(n19302) );
  NAND U20097 ( .A(n19303), .B(n19302), .Z(n19852) );
  NANDN U20098 ( .A(n19305), .B(n19304), .Z(n19309) );
  NANDN U20099 ( .A(n19307), .B(n19306), .Z(n19308) );
  AND U20100 ( .A(n19309), .B(n19308), .Z(n19851) );
  XNOR U20101 ( .A(n19852), .B(n19851), .Z(n19853) );
  NANDN U20102 ( .A(n19311), .B(n19310), .Z(n19315) );
  NANDN U20103 ( .A(n19313), .B(n19312), .Z(n19314) );
  NAND U20104 ( .A(n19315), .B(n19314), .Z(n19588) );
  XOR U20105 ( .A(a[82]), .B(n972), .Z(n19769) );
  OR U20106 ( .A(n19769), .B(n32010), .Z(n19318) );
  NANDN U20107 ( .A(n19316), .B(n32011), .Z(n19317) );
  NAND U20108 ( .A(n19318), .B(n19317), .Z(n19653) );
  XNOR U20109 ( .A(b[25]), .B(n30210), .Z(n19772) );
  NANDN U20110 ( .A(n34219), .B(n19772), .Z(n19321) );
  NAND U20111 ( .A(n34217), .B(n19319), .Z(n19320) );
  NAND U20112 ( .A(n19321), .B(n19320), .Z(n19650) );
  XNOR U20113 ( .A(b[17]), .B(a[80]), .Z(n19775) );
  NANDN U20114 ( .A(n19775), .B(n32543), .Z(n19324) );
  NAND U20115 ( .A(n19322), .B(n32541), .Z(n19323) );
  AND U20116 ( .A(n19324), .B(n19323), .Z(n19651) );
  XNOR U20117 ( .A(n19650), .B(n19651), .Z(n19652) );
  XNOR U20118 ( .A(n19653), .B(n19652), .Z(n19708) );
  XOR U20119 ( .A(b[39]), .B(n26347), .Z(n19778) );
  NANDN U20120 ( .A(n19778), .B(n36553), .Z(n19327) );
  NANDN U20121 ( .A(n19325), .B(n36643), .Z(n19326) );
  NAND U20122 ( .A(n19327), .B(n19326), .Z(n19647) );
  XOR U20123 ( .A(b[51]), .B(n22964), .Z(n19781) );
  NANDN U20124 ( .A(n19781), .B(n37803), .Z(n19330) );
  NANDN U20125 ( .A(n19328), .B(n37802), .Z(n19329) );
  NAND U20126 ( .A(n19330), .B(n19329), .Z(n19644) );
  XOR U20127 ( .A(b[53]), .B(n22289), .Z(n19784) );
  NANDN U20128 ( .A(n19784), .B(n37940), .Z(n19333) );
  NANDN U20129 ( .A(n19331), .B(n37941), .Z(n19332) );
  AND U20130 ( .A(n19333), .B(n19332), .Z(n19645) );
  XNOR U20131 ( .A(n19644), .B(n19645), .Z(n19646) );
  XOR U20132 ( .A(n19647), .B(n19646), .Z(n19709) );
  XOR U20133 ( .A(n19708), .B(n19709), .Z(n19711) );
  NANDN U20134 ( .A(n19335), .B(n19334), .Z(n19339) );
  NAND U20135 ( .A(n19337), .B(n19336), .Z(n19338) );
  NAND U20136 ( .A(n19339), .B(n19338), .Z(n19710) );
  XNOR U20137 ( .A(n19711), .B(n19710), .Z(n19814) );
  NANDN U20138 ( .A(n19341), .B(n19340), .Z(n19345) );
  NAND U20139 ( .A(n19343), .B(n19342), .Z(n19344) );
  NAND U20140 ( .A(n19345), .B(n19344), .Z(n19811) );
  NANDN U20141 ( .A(n19347), .B(n19346), .Z(n19351) );
  NAND U20142 ( .A(n19349), .B(n19348), .Z(n19350) );
  AND U20143 ( .A(n19351), .B(n19350), .Z(n19812) );
  XNOR U20144 ( .A(n19811), .B(n19812), .Z(n19813) );
  XNOR U20145 ( .A(n19814), .B(n19813), .Z(n19836) );
  OR U20146 ( .A(n19353), .B(n19352), .Z(n19357) );
  OR U20147 ( .A(n19355), .B(n19354), .Z(n19356) );
  NAND U20148 ( .A(n19357), .B(n19356), .Z(n19833) );
  NANDN U20149 ( .A(n19359), .B(n19358), .Z(n19363) );
  NANDN U20150 ( .A(n19361), .B(n19360), .Z(n19362) );
  NAND U20151 ( .A(n19363), .B(n19362), .Z(n19834) );
  XNOR U20152 ( .A(n19833), .B(n19834), .Z(n19835) );
  XOR U20153 ( .A(n19836), .B(n19835), .Z(n19840) );
  XOR U20154 ( .A(b[35]), .B(a[62]), .Z(n19748) );
  NAND U20155 ( .A(n35985), .B(n19748), .Z(n19366) );
  NANDN U20156 ( .A(n19364), .B(n35986), .Z(n19365) );
  NAND U20157 ( .A(n19366), .B(n19365), .Z(n19796) );
  XOR U20158 ( .A(n34851), .B(n31123), .Z(n19751) );
  NAND U20159 ( .A(n19751), .B(n29949), .Z(n19369) );
  NAND U20160 ( .A(n29948), .B(n19367), .Z(n19368) );
  NAND U20161 ( .A(n19369), .B(n19368), .Z(n19793) );
  XOR U20162 ( .A(b[55]), .B(n22246), .Z(n19754) );
  NANDN U20163 ( .A(n19754), .B(n38075), .Z(n19372) );
  NANDN U20164 ( .A(n19370), .B(n38073), .Z(n19371) );
  AND U20165 ( .A(n19372), .B(n19371), .Z(n19794) );
  XNOR U20166 ( .A(n19793), .B(n19794), .Z(n19795) );
  XNOR U20167 ( .A(n19796), .B(n19795), .Z(n19613) );
  NANDN U20168 ( .A(n19374), .B(n19373), .Z(n19378) );
  NAND U20169 ( .A(n19376), .B(n19375), .Z(n19377) );
  NAND U20170 ( .A(n19378), .B(n19377), .Z(n19610) );
  XNOR U20171 ( .A(n19610), .B(n19611), .Z(n19612) );
  XOR U20172 ( .A(n19613), .B(n19612), .Z(n19825) );
  XOR U20173 ( .A(a[86]), .B(n970), .Z(n19729) );
  OR U20174 ( .A(n19729), .B(n31369), .Z(n19385) );
  NANDN U20175 ( .A(n19383), .B(n31119), .Z(n19384) );
  NAND U20176 ( .A(n19385), .B(n19384), .Z(n19741) );
  XOR U20177 ( .A(b[43]), .B(n25177), .Z(n19732) );
  NANDN U20178 ( .A(n19732), .B(n37068), .Z(n19388) );
  NANDN U20179 ( .A(n19386), .B(n37069), .Z(n19387) );
  NAND U20180 ( .A(n19388), .B(n19387), .Z(n19738) );
  XNOR U20181 ( .A(b[45]), .B(a[52]), .Z(n19735) );
  NANDN U20182 ( .A(n19735), .B(n37261), .Z(n19391) );
  NANDN U20183 ( .A(n19389), .B(n37262), .Z(n19390) );
  AND U20184 ( .A(n19391), .B(n19390), .Z(n19739) );
  XNOR U20185 ( .A(n19738), .B(n19739), .Z(n19740) );
  XNOR U20186 ( .A(n19741), .B(n19740), .Z(n19625) );
  XOR U20187 ( .A(b[49]), .B(n23447), .Z(n19720) );
  OR U20188 ( .A(n19720), .B(n37756), .Z(n19394) );
  NANDN U20189 ( .A(n19392), .B(n37652), .Z(n19393) );
  NAND U20190 ( .A(n19394), .B(n19393), .Z(n19765) );
  NAND U20191 ( .A(n19395), .B(n37469), .Z(n19397) );
  XOR U20192 ( .A(n978), .B(n24671), .Z(n19723) );
  NAND U20193 ( .A(n19723), .B(n37471), .Z(n19396) );
  AND U20194 ( .A(n19397), .B(n19396), .Z(n19763) );
  XOR U20195 ( .A(a[88]), .B(n969), .Z(n19726) );
  NANDN U20196 ( .A(n19726), .B(n30509), .Z(n19400) );
  NAND U20197 ( .A(n19398), .B(n30846), .Z(n19399) );
  AND U20198 ( .A(n19400), .B(n19399), .Z(n19764) );
  XOR U20199 ( .A(n19765), .B(n19766), .Z(n19622) );
  NANDN U20200 ( .A(n19402), .B(n19401), .Z(n19406) );
  NAND U20201 ( .A(n19404), .B(n19403), .Z(n19405) );
  NAND U20202 ( .A(n19406), .B(n19405), .Z(n19623) );
  XNOR U20203 ( .A(n19622), .B(n19623), .Z(n19624) );
  XOR U20204 ( .A(n19625), .B(n19624), .Z(n19823) );
  XNOR U20205 ( .A(n19823), .B(n19824), .Z(n19826) );
  XNOR U20206 ( .A(n19825), .B(n19826), .Z(n19839) );
  XOR U20207 ( .A(n19840), .B(n19839), .Z(n19841) );
  OR U20208 ( .A(n19412), .B(n19411), .Z(n19416) );
  NAND U20209 ( .A(n19414), .B(n19413), .Z(n19415) );
  NAND U20210 ( .A(n19416), .B(n19415), .Z(n19842) );
  XOR U20211 ( .A(n19841), .B(n19842), .Z(n19587) );
  NANDN U20212 ( .A(n19418), .B(n19417), .Z(n19422) );
  NAND U20213 ( .A(n19420), .B(n19419), .Z(n19421) );
  AND U20214 ( .A(n19422), .B(n19421), .Z(n19832) );
  NANDN U20215 ( .A(n19424), .B(n19423), .Z(n19428) );
  OR U20216 ( .A(n19426), .B(n19425), .Z(n19427) );
  NAND U20217 ( .A(n19428), .B(n19427), .Z(n19829) );
  NANDN U20218 ( .A(n19430), .B(n19429), .Z(n19434) );
  NAND U20219 ( .A(n19432), .B(n19431), .Z(n19433) );
  NAND U20220 ( .A(n19434), .B(n19433), .Z(n19830) );
  XNOR U20221 ( .A(n19829), .B(n19830), .Z(n19831) );
  XNOR U20222 ( .A(n19832), .B(n19831), .Z(n19817) );
  NAND U20223 ( .A(n19436), .B(n19435), .Z(n19440) );
  OR U20224 ( .A(n19438), .B(n19437), .Z(n19439) );
  AND U20225 ( .A(n19440), .B(n19439), .Z(n19818) );
  XNOR U20226 ( .A(n19817), .B(n19818), .Z(n19820) );
  NANDN U20227 ( .A(n19442), .B(n19441), .Z(n19446) );
  NAND U20228 ( .A(n19444), .B(n19443), .Z(n19445) );
  NAND U20229 ( .A(n19446), .B(n19445), .Z(n19600) );
  XOR U20230 ( .A(b[37]), .B(n27436), .Z(n19626) );
  NANDN U20231 ( .A(n19626), .B(n36311), .Z(n19449) );
  NANDN U20232 ( .A(n19447), .B(n36309), .Z(n19448) );
  NAND U20233 ( .A(n19449), .B(n19448), .Z(n19705) );
  XOR U20234 ( .A(a[92]), .B(n968), .Z(n19629) );
  OR U20235 ( .A(n19629), .B(n29363), .Z(n19452) );
  NANDN U20236 ( .A(n19450), .B(n29864), .Z(n19451) );
  NAND U20237 ( .A(n19452), .B(n19451), .Z(n19702) );
  XOR U20238 ( .A(n35191), .B(n967), .Z(n19632) );
  NAND U20239 ( .A(n19632), .B(n28939), .Z(n19455) );
  NAND U20240 ( .A(n28938), .B(n19453), .Z(n19454) );
  AND U20241 ( .A(n19455), .B(n19454), .Z(n19703) );
  XNOR U20242 ( .A(n19702), .B(n19703), .Z(n19704) );
  XOR U20243 ( .A(n19705), .B(n19704), .Z(n19607) );
  XOR U20244 ( .A(a[84]), .B(n971), .Z(n19635) );
  OR U20245 ( .A(n19635), .B(n31550), .Z(n19458) );
  NANDN U20246 ( .A(n19456), .B(n31874), .Z(n19457) );
  NAND U20247 ( .A(n19458), .B(n19457), .Z(n19790) );
  NAND U20248 ( .A(n34848), .B(n19459), .Z(n19461) );
  XOR U20249 ( .A(n35375), .B(n30379), .Z(n19638) );
  NAND U20250 ( .A(n34618), .B(n19638), .Z(n19460) );
  NAND U20251 ( .A(n19461), .B(n19460), .Z(n19787) );
  NAND U20252 ( .A(n35188), .B(n19462), .Z(n19464) );
  XOR U20253 ( .A(n35540), .B(n29868), .Z(n19641) );
  NANDN U20254 ( .A(n34968), .B(n19641), .Z(n19463) );
  AND U20255 ( .A(n19464), .B(n19463), .Z(n19788) );
  XNOR U20256 ( .A(n19787), .B(n19788), .Z(n19789) );
  XOR U20257 ( .A(n19790), .B(n19789), .Z(n19605) );
  NANDN U20258 ( .A(n19466), .B(n19465), .Z(n19470) );
  NAND U20259 ( .A(n19468), .B(n19467), .Z(n19469) );
  AND U20260 ( .A(n19470), .B(n19469), .Z(n19604) );
  XOR U20261 ( .A(n19605), .B(n19604), .Z(n19606) );
  XOR U20262 ( .A(n19607), .B(n19606), .Z(n19599) );
  NANDN U20263 ( .A(n19472), .B(n19471), .Z(n19476) );
  NAND U20264 ( .A(n19474), .B(n19473), .Z(n19475) );
  NAND U20265 ( .A(n19476), .B(n19475), .Z(n19746) );
  NAND U20266 ( .A(a[32]), .B(b[63]), .Z(n19760) );
  NANDN U20267 ( .A(n19477), .B(n38369), .Z(n19479) );
  XOR U20268 ( .A(b[61]), .B(n19980), .Z(n19657) );
  OR U20269 ( .A(n19657), .B(n38371), .Z(n19478) );
  NAND U20270 ( .A(n19479), .B(n19478), .Z(n19758) );
  NANDN U20271 ( .A(n19480), .B(n35311), .Z(n19482) );
  XOR U20272 ( .A(b[31]), .B(n28701), .Z(n19660) );
  NANDN U20273 ( .A(n19660), .B(n35313), .Z(n19481) );
  AND U20274 ( .A(n19482), .B(n19481), .Z(n19757) );
  XNOR U20275 ( .A(n19758), .B(n19757), .Z(n19759) );
  XOR U20276 ( .A(n19760), .B(n19759), .Z(n19744) );
  NAND U20277 ( .A(n33283), .B(n19483), .Z(n19485) );
  XOR U20278 ( .A(n33020), .B(n31870), .Z(n19663) );
  NANDN U20279 ( .A(n33021), .B(n19663), .Z(n19484) );
  NAND U20280 ( .A(n19485), .B(n19484), .Z(n19675) );
  XNOR U20281 ( .A(b[21]), .B(a[76]), .Z(n19666) );
  OR U20282 ( .A(n19666), .B(n33634), .Z(n19488) );
  NAND U20283 ( .A(n19486), .B(n33464), .Z(n19487) );
  NAND U20284 ( .A(n19488), .B(n19487), .Z(n19672) );
  NAND U20285 ( .A(n34044), .B(n19489), .Z(n19491) );
  XOR U20286 ( .A(n34510), .B(n31372), .Z(n19669) );
  NANDN U20287 ( .A(n33867), .B(n19669), .Z(n19490) );
  AND U20288 ( .A(n19491), .B(n19490), .Z(n19673) );
  XNOR U20289 ( .A(n19672), .B(n19673), .Z(n19674) );
  XNOR U20290 ( .A(n19675), .B(n19674), .Z(n19745) );
  XNOR U20291 ( .A(n19744), .B(n19745), .Z(n19747) );
  XNOR U20292 ( .A(n19746), .B(n19747), .Z(n19598) );
  XOR U20293 ( .A(n19599), .B(n19598), .Z(n19601) );
  XNOR U20294 ( .A(n19600), .B(n19601), .Z(n19717) );
  NANDN U20295 ( .A(n19493), .B(n19492), .Z(n19497) );
  NAND U20296 ( .A(n19495), .B(n19494), .Z(n19496) );
  NAND U20297 ( .A(n19497), .B(n19496), .Z(n19808) );
  XNOR U20298 ( .A(b[41]), .B(a[56]), .Z(n19678) );
  OR U20299 ( .A(n19678), .B(n36905), .Z(n19500) );
  NANDN U20300 ( .A(n19498), .B(n36807), .Z(n19499) );
  NAND U20301 ( .A(n19500), .B(n19499), .Z(n19699) );
  XOR U20302 ( .A(b[57]), .B(n21149), .Z(n19681) );
  OR U20303 ( .A(n19681), .B(n965), .Z(n19503) );
  NANDN U20304 ( .A(n19501), .B(n38194), .Z(n19502) );
  NAND U20305 ( .A(n19503), .B(n19502), .Z(n19696) );
  NAND U20306 ( .A(n38326), .B(n19504), .Z(n19506) );
  XOR U20307 ( .A(n38400), .B(n20686), .Z(n19684) );
  NANDN U20308 ( .A(n38273), .B(n19684), .Z(n19505) );
  AND U20309 ( .A(n19506), .B(n19505), .Z(n19697) );
  XNOR U20310 ( .A(n19696), .B(n19697), .Z(n19698) );
  XOR U20311 ( .A(n19699), .B(n19698), .Z(n19805) );
  XNOR U20312 ( .A(b[33]), .B(a[64]), .Z(n19687) );
  NANDN U20313 ( .A(n19687), .B(n35620), .Z(n19509) );
  NANDN U20314 ( .A(n19507), .B(n35621), .Z(n19508) );
  NAND U20315 ( .A(n19509), .B(n19508), .Z(n19802) );
  NANDN U20316 ( .A(n966), .B(a[96]), .Z(n19510) );
  XOR U20317 ( .A(n29232), .B(n19510), .Z(n19512) );
  IV U20318 ( .A(a[95]), .Z(n35628) );
  NANDN U20319 ( .A(n35628), .B(n966), .Z(n19511) );
  AND U20320 ( .A(n19512), .B(n19511), .Z(n19799) );
  XOR U20321 ( .A(b[63]), .B(n19513), .Z(n19693) );
  NANDN U20322 ( .A(n19693), .B(n38422), .Z(n19516) );
  NANDN U20323 ( .A(n19514), .B(n38423), .Z(n19515) );
  AND U20324 ( .A(n19516), .B(n19515), .Z(n19800) );
  XNOR U20325 ( .A(n19799), .B(n19800), .Z(n19801) );
  XOR U20326 ( .A(n19802), .B(n19801), .Z(n19806) );
  XNOR U20327 ( .A(n19805), .B(n19806), .Z(n19807) );
  XNOR U20328 ( .A(n19808), .B(n19807), .Z(n19619) );
  NANDN U20329 ( .A(n19518), .B(n19517), .Z(n19522) );
  NAND U20330 ( .A(n19520), .B(n19519), .Z(n19521) );
  NAND U20331 ( .A(n19522), .B(n19521), .Z(n19616) );
  NANDN U20332 ( .A(n19524), .B(n19523), .Z(n19528) );
  NAND U20333 ( .A(n19526), .B(n19525), .Z(n19527) );
  AND U20334 ( .A(n19528), .B(n19527), .Z(n19617) );
  XNOR U20335 ( .A(n19616), .B(n19617), .Z(n19618) );
  XOR U20336 ( .A(n19619), .B(n19618), .Z(n19715) );
  NANDN U20337 ( .A(n19530), .B(n19529), .Z(n19534) );
  NAND U20338 ( .A(n19532), .B(n19531), .Z(n19533) );
  AND U20339 ( .A(n19534), .B(n19533), .Z(n19714) );
  XOR U20340 ( .A(n19715), .B(n19714), .Z(n19716) );
  XOR U20341 ( .A(n19717), .B(n19716), .Z(n19819) );
  XNOR U20342 ( .A(n19820), .B(n19819), .Z(n19586) );
  XNOR U20343 ( .A(n19587), .B(n19586), .Z(n19589) );
  XNOR U20344 ( .A(n19588), .B(n19589), .Z(n19847) );
  NAND U20345 ( .A(n19536), .B(n19535), .Z(n19540) );
  NANDN U20346 ( .A(n19538), .B(n19537), .Z(n19539) );
  NAND U20347 ( .A(n19540), .B(n19539), .Z(n19595) );
  OR U20348 ( .A(n19542), .B(n19541), .Z(n19546) );
  NAND U20349 ( .A(n19544), .B(n19543), .Z(n19545) );
  NAND U20350 ( .A(n19546), .B(n19545), .Z(n19593) );
  OR U20351 ( .A(n19548), .B(n19547), .Z(n19552) );
  NAND U20352 ( .A(n19550), .B(n19549), .Z(n19551) );
  AND U20353 ( .A(n19552), .B(n19551), .Z(n19592) );
  XNOR U20354 ( .A(n19593), .B(n19592), .Z(n19594) );
  XOR U20355 ( .A(n19595), .B(n19594), .Z(n19845) );
  XNOR U20356 ( .A(n19845), .B(n19846), .Z(n19848) );
  XOR U20357 ( .A(n19847), .B(n19848), .Z(n19854) );
  XNOR U20358 ( .A(n19853), .B(n19854), .Z(n19857) );
  NANDN U20359 ( .A(n19558), .B(n19557), .Z(n19562) );
  NAND U20360 ( .A(n19560), .B(n19559), .Z(n19561) );
  NAND U20361 ( .A(n19562), .B(n19561), .Z(n19858) );
  XNOR U20362 ( .A(n19857), .B(n19858), .Z(n19859) );
  NANDN U20363 ( .A(n19564), .B(n19563), .Z(n19568) );
  NANDN U20364 ( .A(n19566), .B(n19565), .Z(n19567) );
  NAND U20365 ( .A(n19568), .B(n19567), .Z(n19860) );
  XOR U20366 ( .A(n19859), .B(n19860), .Z(n19580) );
  NANDN U20367 ( .A(n19570), .B(n19569), .Z(n19574) );
  NAND U20368 ( .A(n19572), .B(n19571), .Z(n19573) );
  NAND U20369 ( .A(n19574), .B(n19573), .Z(n19581) );
  XNOR U20370 ( .A(n19580), .B(n19581), .Z(n19582) );
  XNOR U20371 ( .A(n19583), .B(n19582), .Z(n19861) );
  XNOR U20372 ( .A(n19861), .B(sreg[160]), .Z(n19863) );
  NAND U20373 ( .A(n19575), .B(sreg[159]), .Z(n19579) );
  OR U20374 ( .A(n19577), .B(n19576), .Z(n19578) );
  AND U20375 ( .A(n19579), .B(n19578), .Z(n19862) );
  XOR U20376 ( .A(n19863), .B(n19862), .Z(c[160]) );
  NANDN U20377 ( .A(n19581), .B(n19580), .Z(n19585) );
  NAND U20378 ( .A(n19583), .B(n19582), .Z(n19584) );
  NAND U20379 ( .A(n19585), .B(n19584), .Z(n19869) );
  NAND U20380 ( .A(n19587), .B(n19586), .Z(n19591) );
  NANDN U20381 ( .A(n19589), .B(n19588), .Z(n19590) );
  NAND U20382 ( .A(n19591), .B(n19590), .Z(n20139) );
  NANDN U20383 ( .A(n19593), .B(n19592), .Z(n19597) );
  NANDN U20384 ( .A(n19595), .B(n19594), .Z(n19596) );
  NAND U20385 ( .A(n19597), .B(n19596), .Z(n20140) );
  XNOR U20386 ( .A(n20139), .B(n20140), .Z(n20141) );
  NANDN U20387 ( .A(n19599), .B(n19598), .Z(n19603) );
  OR U20388 ( .A(n19601), .B(n19600), .Z(n19602) );
  NAND U20389 ( .A(n19603), .B(n19602), .Z(n20107) );
  NANDN U20390 ( .A(n19605), .B(n19604), .Z(n19609) );
  OR U20391 ( .A(n19607), .B(n19606), .Z(n19608) );
  NAND U20392 ( .A(n19609), .B(n19608), .Z(n20125) );
  NANDN U20393 ( .A(n19611), .B(n19610), .Z(n19615) );
  NAND U20394 ( .A(n19613), .B(n19612), .Z(n19614) );
  NAND U20395 ( .A(n19615), .B(n19614), .Z(n20123) );
  NANDN U20396 ( .A(n19617), .B(n19616), .Z(n19621) );
  NAND U20397 ( .A(n19619), .B(n19618), .Z(n19620) );
  NAND U20398 ( .A(n19621), .B(n19620), .Z(n20124) );
  XNOR U20399 ( .A(n20123), .B(n20124), .Z(n20126) );
  XNOR U20400 ( .A(n20125), .B(n20126), .Z(n20108) );
  XOR U20401 ( .A(n20107), .B(n20108), .Z(n20109) );
  XOR U20402 ( .A(b[37]), .B(n27773), .Z(n19935) );
  NANDN U20403 ( .A(n19935), .B(n36311), .Z(n19628) );
  NANDN U20404 ( .A(n19626), .B(n36309), .Z(n19627) );
  NAND U20405 ( .A(n19628), .B(n19627), .Z(n19993) );
  XOR U20406 ( .A(a[93]), .B(n968), .Z(n19938) );
  OR U20407 ( .A(n19938), .B(n29363), .Z(n19631) );
  NANDN U20408 ( .A(n19629), .B(n29864), .Z(n19630) );
  NAND U20409 ( .A(n19631), .B(n19630), .Z(n19990) );
  XOR U20410 ( .A(n35628), .B(n967), .Z(n19941) );
  NAND U20411 ( .A(n19941), .B(n28939), .Z(n19634) );
  NAND U20412 ( .A(n28938), .B(n19632), .Z(n19633) );
  AND U20413 ( .A(n19634), .B(n19633), .Z(n19991) );
  XNOR U20414 ( .A(n19990), .B(n19991), .Z(n19992) );
  XNOR U20415 ( .A(n19993), .B(n19992), .Z(n19884) );
  XNOR U20416 ( .A(a[85]), .B(b[13]), .Z(n19944) );
  OR U20417 ( .A(n19944), .B(n31550), .Z(n19637) );
  NANDN U20418 ( .A(n19635), .B(n31874), .Z(n19636) );
  NAND U20419 ( .A(n19637), .B(n19636), .Z(n20098) );
  NAND U20420 ( .A(n34848), .B(n19638), .Z(n19640) );
  XOR U20421 ( .A(n35375), .B(n30543), .Z(n19947) );
  NAND U20422 ( .A(n34618), .B(n19947), .Z(n19639) );
  NAND U20423 ( .A(n19640), .B(n19639), .Z(n20095) );
  NAND U20424 ( .A(n35188), .B(n19641), .Z(n19643) );
  XNOR U20425 ( .A(n35540), .B(a[69]), .Z(n19950) );
  NANDN U20426 ( .A(n34968), .B(n19950), .Z(n19642) );
  AND U20427 ( .A(n19643), .B(n19642), .Z(n20096) );
  XNOR U20428 ( .A(n20095), .B(n20096), .Z(n20097) );
  XOR U20429 ( .A(n20098), .B(n20097), .Z(n19885) );
  XNOR U20430 ( .A(n19884), .B(n19885), .Z(n19886) );
  NANDN U20431 ( .A(n19645), .B(n19644), .Z(n19649) );
  NAND U20432 ( .A(n19647), .B(n19646), .Z(n19648) );
  NAND U20433 ( .A(n19649), .B(n19648), .Z(n19887) );
  XOR U20434 ( .A(n19886), .B(n19887), .Z(n19902) );
  NANDN U20435 ( .A(n19651), .B(n19650), .Z(n19655) );
  NAND U20436 ( .A(n19653), .B(n19652), .Z(n19654) );
  NAND U20437 ( .A(n19655), .B(n19654), .Z(n20055) );
  ANDN U20438 ( .B(b[63]), .A(n19656), .Z(n20020) );
  NANDN U20439 ( .A(n19657), .B(n38369), .Z(n19659) );
  XOR U20440 ( .A(b[61]), .B(n20352), .Z(n19929) );
  OR U20441 ( .A(n19929), .B(n38371), .Z(n19658) );
  NAND U20442 ( .A(n19659), .B(n19658), .Z(n20018) );
  NANDN U20443 ( .A(n19660), .B(n35311), .Z(n19662) );
  XOR U20444 ( .A(b[31]), .B(n29372), .Z(n19932) );
  NANDN U20445 ( .A(n19932), .B(n35313), .Z(n19661) );
  AND U20446 ( .A(n19662), .B(n19661), .Z(n20017) );
  XNOR U20447 ( .A(n20018), .B(n20017), .Z(n20019) );
  XOR U20448 ( .A(n20020), .B(n20019), .Z(n20053) );
  NAND U20449 ( .A(n33283), .B(n19663), .Z(n19665) );
  XNOR U20450 ( .A(n33020), .B(a[79]), .Z(n19914) );
  NANDN U20451 ( .A(n33021), .B(n19914), .Z(n19664) );
  NAND U20452 ( .A(n19665), .B(n19664), .Z(n19962) );
  XOR U20453 ( .A(b[21]), .B(a[77]), .Z(n19917) );
  NANDN U20454 ( .A(n33634), .B(n19917), .Z(n19668) );
  NANDN U20455 ( .A(n19666), .B(n33464), .Z(n19667) );
  NAND U20456 ( .A(n19668), .B(n19667), .Z(n19959) );
  NAND U20457 ( .A(n34044), .B(n19669), .Z(n19671) );
  XNOR U20458 ( .A(n34510), .B(a[75]), .Z(n19920) );
  NANDN U20459 ( .A(n33867), .B(n19920), .Z(n19670) );
  AND U20460 ( .A(n19671), .B(n19670), .Z(n19960) );
  XNOR U20461 ( .A(n19959), .B(n19960), .Z(n19961) );
  XNOR U20462 ( .A(n19962), .B(n19961), .Z(n20054) );
  XOR U20463 ( .A(n20053), .B(n20054), .Z(n20056) );
  XOR U20464 ( .A(n20055), .B(n20056), .Z(n19903) );
  XNOR U20465 ( .A(n19902), .B(n19903), .Z(n19904) );
  XOR U20466 ( .A(n19905), .B(n19904), .Z(n20005) );
  NANDN U20467 ( .A(n19673), .B(n19672), .Z(n19677) );
  NAND U20468 ( .A(n19675), .B(n19674), .Z(n19676) );
  NAND U20469 ( .A(n19677), .B(n19676), .Z(n20062) );
  XNOR U20470 ( .A(b[41]), .B(a[57]), .Z(n19965) );
  OR U20471 ( .A(n19965), .B(n36905), .Z(n19680) );
  NANDN U20472 ( .A(n19678), .B(n36807), .Z(n19679) );
  NAND U20473 ( .A(n19680), .B(n19679), .Z(n19987) );
  XOR U20474 ( .A(b[57]), .B(n21441), .Z(n19968) );
  OR U20475 ( .A(n19968), .B(n965), .Z(n19683) );
  NANDN U20476 ( .A(n19681), .B(n38194), .Z(n19682) );
  NAND U20477 ( .A(n19683), .B(n19682), .Z(n19984) );
  NAND U20478 ( .A(n38326), .B(n19684), .Z(n19686) );
  XOR U20479 ( .A(n38400), .B(n20867), .Z(n19971) );
  NANDN U20480 ( .A(n38273), .B(n19971), .Z(n19685) );
  AND U20481 ( .A(n19686), .B(n19685), .Z(n19985) );
  XNOR U20482 ( .A(n19984), .B(n19985), .Z(n19986) );
  XOR U20483 ( .A(n19987), .B(n19986), .Z(n20059) );
  XOR U20484 ( .A(b[33]), .B(n28403), .Z(n19974) );
  NANDN U20485 ( .A(n19974), .B(n35620), .Z(n19689) );
  NANDN U20486 ( .A(n19687), .B(n35621), .Z(n19688) );
  NAND U20487 ( .A(n19689), .B(n19688), .Z(n20074) );
  NANDN U20488 ( .A(n966), .B(a[97]), .Z(n19690) );
  XOR U20489 ( .A(n29232), .B(n19690), .Z(n19692) );
  IV U20490 ( .A(a[96]), .Z(n35545) );
  NANDN U20491 ( .A(n35545), .B(n966), .Z(n19691) );
  AND U20492 ( .A(n19692), .B(n19691), .Z(n20071) );
  XOR U20493 ( .A(b[63]), .B(n20315), .Z(n19981) );
  NANDN U20494 ( .A(n19981), .B(n38422), .Z(n19695) );
  NANDN U20495 ( .A(n19693), .B(n38423), .Z(n19694) );
  AND U20496 ( .A(n19695), .B(n19694), .Z(n20072) );
  XNOR U20497 ( .A(n20071), .B(n20072), .Z(n20073) );
  XOR U20498 ( .A(n20074), .B(n20073), .Z(n20060) );
  XNOR U20499 ( .A(n20059), .B(n20060), .Z(n20061) );
  XNOR U20500 ( .A(n20062), .B(n20061), .Z(n19899) );
  NANDN U20501 ( .A(n19697), .B(n19696), .Z(n19701) );
  NAND U20502 ( .A(n19699), .B(n19698), .Z(n19700) );
  NAND U20503 ( .A(n19701), .B(n19700), .Z(n19896) );
  NANDN U20504 ( .A(n19703), .B(n19702), .Z(n19707) );
  NAND U20505 ( .A(n19705), .B(n19704), .Z(n19706) );
  AND U20506 ( .A(n19707), .B(n19706), .Z(n19897) );
  XNOR U20507 ( .A(n19896), .B(n19897), .Z(n19898) );
  XOR U20508 ( .A(n19899), .B(n19898), .Z(n20003) );
  NANDN U20509 ( .A(n19709), .B(n19708), .Z(n19713) );
  OR U20510 ( .A(n19711), .B(n19710), .Z(n19712) );
  AND U20511 ( .A(n19713), .B(n19712), .Z(n20002) );
  XOR U20512 ( .A(n20003), .B(n20002), .Z(n20004) );
  XNOR U20513 ( .A(n20005), .B(n20004), .Z(n20110) );
  XOR U20514 ( .A(n20109), .B(n20110), .Z(n19872) );
  OR U20515 ( .A(n19715), .B(n19714), .Z(n19719) );
  NAND U20516 ( .A(n19717), .B(n19716), .Z(n19718) );
  NAND U20517 ( .A(n19719), .B(n19718), .Z(n20130) );
  XOR U20518 ( .A(b[49]), .B(n23852), .Z(n20038) );
  OR U20519 ( .A(n20038), .B(n37756), .Z(n19722) );
  NANDN U20520 ( .A(n19720), .B(n37652), .Z(n19721) );
  NAND U20521 ( .A(n19722), .B(n19721), .Z(n20025) );
  NAND U20522 ( .A(n37469), .B(n19723), .Z(n19725) );
  XOR U20523 ( .A(n978), .B(n24288), .Z(n20041) );
  NAND U20524 ( .A(n20041), .B(n37471), .Z(n19724) );
  AND U20525 ( .A(n19725), .B(n19724), .Z(n20023) );
  XNOR U20526 ( .A(a[89]), .B(b[9]), .Z(n20044) );
  NANDN U20527 ( .A(n20044), .B(n30509), .Z(n19728) );
  NANDN U20528 ( .A(n19726), .B(n30846), .Z(n19727) );
  AND U20529 ( .A(n19728), .B(n19727), .Z(n20024) );
  XOR U20530 ( .A(n20025), .B(n20026), .Z(n19908) );
  XNOR U20531 ( .A(a[87]), .B(b[11]), .Z(n20029) );
  OR U20532 ( .A(n20029), .B(n31369), .Z(n19731) );
  NANDN U20533 ( .A(n19729), .B(n31119), .Z(n19730) );
  NAND U20534 ( .A(n19731), .B(n19730), .Z(n20050) );
  XOR U20535 ( .A(b[43]), .B(n25466), .Z(n20032) );
  NANDN U20536 ( .A(n20032), .B(n37068), .Z(n19734) );
  NANDN U20537 ( .A(n19732), .B(n37069), .Z(n19733) );
  NAND U20538 ( .A(n19734), .B(n19733), .Z(n20047) );
  XNOR U20539 ( .A(b[45]), .B(a[53]), .Z(n20035) );
  NANDN U20540 ( .A(n20035), .B(n37261), .Z(n19737) );
  NANDN U20541 ( .A(n19735), .B(n37262), .Z(n19736) );
  AND U20542 ( .A(n19737), .B(n19736), .Z(n20048) );
  XNOR U20543 ( .A(n20047), .B(n20048), .Z(n20049) );
  XOR U20544 ( .A(n20050), .B(n20049), .Z(n19909) );
  XNOR U20545 ( .A(n19908), .B(n19909), .Z(n19910) );
  NANDN U20546 ( .A(n19739), .B(n19738), .Z(n19743) );
  NAND U20547 ( .A(n19741), .B(n19740), .Z(n19742) );
  AND U20548 ( .A(n19743), .B(n19742), .Z(n19911) );
  XNOR U20549 ( .A(n19910), .B(n19911), .Z(n20114) );
  XNOR U20550 ( .A(n20114), .B(n20113), .Z(n20115) );
  XOR U20551 ( .A(b[35]), .B(a[63]), .Z(n20008) );
  NAND U20552 ( .A(n35985), .B(n20008), .Z(n19750) );
  NAND U20553 ( .A(n19748), .B(n35986), .Z(n19749) );
  NAND U20554 ( .A(n19750), .B(n19749), .Z(n20104) );
  XNOR U20555 ( .A(a[91]), .B(n31123), .Z(n20011) );
  NAND U20556 ( .A(n20011), .B(n29949), .Z(n19753) );
  NAND U20557 ( .A(n29948), .B(n19751), .Z(n19752) );
  NAND U20558 ( .A(n19753), .B(n19752), .Z(n20101) );
  XOR U20559 ( .A(b[55]), .B(n21996), .Z(n20014) );
  NANDN U20560 ( .A(n20014), .B(n38075), .Z(n19756) );
  NANDN U20561 ( .A(n19754), .B(n38073), .Z(n19755) );
  AND U20562 ( .A(n19756), .B(n19755), .Z(n20102) );
  XNOR U20563 ( .A(n20101), .B(n20102), .Z(n20103) );
  XNOR U20564 ( .A(n20104), .B(n20103), .Z(n19893) );
  NANDN U20565 ( .A(n19758), .B(n19757), .Z(n19762) );
  NAND U20566 ( .A(n19760), .B(n19759), .Z(n19761) );
  NAND U20567 ( .A(n19762), .B(n19761), .Z(n19890) );
  OR U20568 ( .A(n19764), .B(n19763), .Z(n19768) );
  NANDN U20569 ( .A(n19766), .B(n19765), .Z(n19767) );
  NAND U20570 ( .A(n19768), .B(n19767), .Z(n19891) );
  XNOR U20571 ( .A(n19890), .B(n19891), .Z(n19892) );
  XOR U20572 ( .A(n19893), .B(n19892), .Z(n20116) );
  XOR U20573 ( .A(n20115), .B(n20116), .Z(n20127) );
  XNOR U20574 ( .A(a[83]), .B(b[15]), .Z(n20086) );
  OR U20575 ( .A(n20086), .B(n32010), .Z(n19771) );
  NANDN U20576 ( .A(n19769), .B(n32011), .Z(n19770) );
  NAND U20577 ( .A(n19771), .B(n19770), .Z(n19926) );
  XOR U20578 ( .A(b[25]), .B(a[73]), .Z(n20089) );
  NANDN U20579 ( .A(n34219), .B(n20089), .Z(n19774) );
  NAND U20580 ( .A(n34217), .B(n19772), .Z(n19773) );
  NAND U20581 ( .A(n19774), .B(n19773), .Z(n19923) );
  XOR U20582 ( .A(b[17]), .B(a[81]), .Z(n20092) );
  NAND U20583 ( .A(n20092), .B(n32543), .Z(n19777) );
  NANDN U20584 ( .A(n19775), .B(n32541), .Z(n19776) );
  AND U20585 ( .A(n19777), .B(n19776), .Z(n19924) );
  XNOR U20586 ( .A(n19923), .B(n19924), .Z(n19925) );
  XNOR U20587 ( .A(n19926), .B(n19925), .Z(n19996) );
  XNOR U20588 ( .A(b[39]), .B(a[59]), .Z(n20077) );
  NANDN U20589 ( .A(n20077), .B(n36553), .Z(n19780) );
  NANDN U20590 ( .A(n19778), .B(n36643), .Z(n19779) );
  NAND U20591 ( .A(n19780), .B(n19779), .Z(n19956) );
  XOR U20592 ( .A(b[51]), .B(n23149), .Z(n20080) );
  NANDN U20593 ( .A(n20080), .B(n37803), .Z(n19783) );
  NANDN U20594 ( .A(n19781), .B(n37802), .Z(n19782) );
  NAND U20595 ( .A(n19783), .B(n19782), .Z(n19953) );
  XOR U20596 ( .A(b[53]), .B(n22579), .Z(n20083) );
  NANDN U20597 ( .A(n20083), .B(n37940), .Z(n19786) );
  NANDN U20598 ( .A(n19784), .B(n37941), .Z(n19785) );
  AND U20599 ( .A(n19786), .B(n19785), .Z(n19954) );
  XNOR U20600 ( .A(n19953), .B(n19954), .Z(n19955) );
  XOR U20601 ( .A(n19956), .B(n19955), .Z(n19997) );
  XOR U20602 ( .A(n19996), .B(n19997), .Z(n19999) );
  NANDN U20603 ( .A(n19788), .B(n19787), .Z(n19792) );
  NAND U20604 ( .A(n19790), .B(n19789), .Z(n19791) );
  NAND U20605 ( .A(n19792), .B(n19791), .Z(n19998) );
  XNOR U20606 ( .A(n19999), .B(n19998), .Z(n20068) );
  NANDN U20607 ( .A(n19794), .B(n19793), .Z(n19798) );
  NAND U20608 ( .A(n19796), .B(n19795), .Z(n19797) );
  NAND U20609 ( .A(n19798), .B(n19797), .Z(n20065) );
  NANDN U20610 ( .A(n19800), .B(n19799), .Z(n19804) );
  NAND U20611 ( .A(n19802), .B(n19801), .Z(n19803) );
  AND U20612 ( .A(n19804), .B(n19803), .Z(n20066) );
  XNOR U20613 ( .A(n20065), .B(n20066), .Z(n20067) );
  XNOR U20614 ( .A(n20068), .B(n20067), .Z(n20119) );
  OR U20615 ( .A(n19806), .B(n19805), .Z(n19810) );
  OR U20616 ( .A(n19808), .B(n19807), .Z(n19809) );
  AND U20617 ( .A(n19810), .B(n19809), .Z(n20120) );
  XNOR U20618 ( .A(n20119), .B(n20120), .Z(n20121) );
  NANDN U20619 ( .A(n19812), .B(n19811), .Z(n19816) );
  NAND U20620 ( .A(n19814), .B(n19813), .Z(n19815) );
  AND U20621 ( .A(n19816), .B(n19815), .Z(n20122) );
  XNOR U20622 ( .A(n20121), .B(n20122), .Z(n20128) );
  XNOR U20623 ( .A(n20127), .B(n20128), .Z(n20129) );
  XOR U20624 ( .A(n20130), .B(n20129), .Z(n19873) );
  XNOR U20625 ( .A(n19872), .B(n19873), .Z(n19874) );
  NAND U20626 ( .A(n19818), .B(n19817), .Z(n19822) );
  NANDN U20627 ( .A(n19820), .B(n19819), .Z(n19821) );
  NAND U20628 ( .A(n19822), .B(n19821), .Z(n19875) );
  XOR U20629 ( .A(n19874), .B(n19875), .Z(n20136) );
  NAND U20630 ( .A(n19824), .B(n19823), .Z(n19828) );
  NANDN U20631 ( .A(n19826), .B(n19825), .Z(n19827) );
  NAND U20632 ( .A(n19828), .B(n19827), .Z(n19881) );
  NANDN U20633 ( .A(n19834), .B(n19833), .Z(n19838) );
  NAND U20634 ( .A(n19836), .B(n19835), .Z(n19837) );
  AND U20635 ( .A(n19838), .B(n19837), .Z(n19878) );
  XNOR U20636 ( .A(n19879), .B(n19878), .Z(n19880) );
  XOR U20637 ( .A(n19881), .B(n19880), .Z(n20133) );
  OR U20638 ( .A(n19840), .B(n19839), .Z(n19844) );
  NANDN U20639 ( .A(n19842), .B(n19841), .Z(n19843) );
  NAND U20640 ( .A(n19844), .B(n19843), .Z(n20134) );
  XNOR U20641 ( .A(n20133), .B(n20134), .Z(n20135) );
  XNOR U20642 ( .A(n20136), .B(n20135), .Z(n20142) );
  XOR U20643 ( .A(n20141), .B(n20142), .Z(n20145) );
  NANDN U20644 ( .A(n19846), .B(n19845), .Z(n19850) );
  NAND U20645 ( .A(n19848), .B(n19847), .Z(n19849) );
  NAND U20646 ( .A(n19850), .B(n19849), .Z(n20146) );
  XNOR U20647 ( .A(n20145), .B(n20146), .Z(n20147) );
  NANDN U20648 ( .A(n19852), .B(n19851), .Z(n19856) );
  NAND U20649 ( .A(n19854), .B(n19853), .Z(n19855) );
  NAND U20650 ( .A(n19856), .B(n19855), .Z(n20148) );
  XOR U20651 ( .A(n20147), .B(n20148), .Z(n19866) );
  XNOR U20652 ( .A(n19866), .B(n19867), .Z(n19868) );
  XNOR U20653 ( .A(n19869), .B(n19868), .Z(n20151) );
  XNOR U20654 ( .A(n20151), .B(sreg[161]), .Z(n20153) );
  NAND U20655 ( .A(n19861), .B(sreg[160]), .Z(n19865) );
  OR U20656 ( .A(n19863), .B(n19862), .Z(n19864) );
  AND U20657 ( .A(n19865), .B(n19864), .Z(n20152) );
  XOR U20658 ( .A(n20153), .B(n20152), .Z(c[161]) );
  NANDN U20659 ( .A(n19867), .B(n19866), .Z(n19871) );
  NAND U20660 ( .A(n19869), .B(n19868), .Z(n19870) );
  NAND U20661 ( .A(n19871), .B(n19870), .Z(n20159) );
  NANDN U20662 ( .A(n19873), .B(n19872), .Z(n19877) );
  NANDN U20663 ( .A(n19875), .B(n19874), .Z(n19876) );
  NAND U20664 ( .A(n19877), .B(n19876), .Z(n20435) );
  NANDN U20665 ( .A(n19879), .B(n19878), .Z(n19883) );
  NANDN U20666 ( .A(n19881), .B(n19880), .Z(n19882) );
  AND U20667 ( .A(n19883), .B(n19882), .Z(n20434) );
  XNOR U20668 ( .A(n20435), .B(n20434), .Z(n20436) );
  NANDN U20669 ( .A(n19885), .B(n19884), .Z(n19889) );
  NANDN U20670 ( .A(n19887), .B(n19886), .Z(n19888) );
  NAND U20671 ( .A(n19889), .B(n19888), .Z(n20407) );
  NANDN U20672 ( .A(n19891), .B(n19890), .Z(n19895) );
  NAND U20673 ( .A(n19893), .B(n19892), .Z(n19894) );
  AND U20674 ( .A(n19895), .B(n19894), .Z(n20404) );
  NANDN U20675 ( .A(n19897), .B(n19896), .Z(n19901) );
  NAND U20676 ( .A(n19899), .B(n19898), .Z(n19900) );
  NAND U20677 ( .A(n19901), .B(n19900), .Z(n20405) );
  XNOR U20678 ( .A(n20407), .B(n20406), .Z(n20163) );
  NANDN U20679 ( .A(n19903), .B(n19902), .Z(n19907) );
  NANDN U20680 ( .A(n19905), .B(n19904), .Z(n19906) );
  AND U20681 ( .A(n19907), .B(n19906), .Z(n20162) );
  XNOR U20682 ( .A(n20163), .B(n20162), .Z(n20164) );
  NANDN U20683 ( .A(n19909), .B(n19908), .Z(n19913) );
  NAND U20684 ( .A(n19911), .B(n19910), .Z(n19912) );
  NAND U20685 ( .A(n19913), .B(n19912), .Z(n20276) );
  NAND U20686 ( .A(n33283), .B(n19914), .Z(n19916) );
  XOR U20687 ( .A(n33020), .B(n32814), .Z(n20322) );
  NANDN U20688 ( .A(n33021), .B(n20322), .Z(n19915) );
  NAND U20689 ( .A(n19916), .B(n19915), .Z(n20334) );
  XNOR U20690 ( .A(b[21]), .B(a[78]), .Z(n20325) );
  OR U20691 ( .A(n20325), .B(n33634), .Z(n19919) );
  NAND U20692 ( .A(n19917), .B(n33464), .Z(n19918) );
  NAND U20693 ( .A(n19919), .B(n19918), .Z(n20331) );
  NAND U20694 ( .A(n34044), .B(n19920), .Z(n19922) );
  XOR U20695 ( .A(n34510), .B(n31363), .Z(n20328) );
  NANDN U20696 ( .A(n33867), .B(n20328), .Z(n19921) );
  AND U20697 ( .A(n19922), .B(n19921), .Z(n20332) );
  XNOR U20698 ( .A(n20331), .B(n20332), .Z(n20333) );
  XNOR U20699 ( .A(n20334), .B(n20333), .Z(n20216) );
  NANDN U20700 ( .A(n19924), .B(n19923), .Z(n19928) );
  NAND U20701 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U20702 ( .A(n19928), .B(n19927), .Z(n20217) );
  XNOR U20703 ( .A(n20216), .B(n20217), .Z(n20218) );
  NAND U20704 ( .A(a[34]), .B(b[63]), .Z(n20258) );
  NANDN U20705 ( .A(n19929), .B(n38369), .Z(n19931) );
  XOR U20706 ( .A(b[61]), .B(n20686), .Z(n20316) );
  OR U20707 ( .A(n20316), .B(n38371), .Z(n19930) );
  NAND U20708 ( .A(n19931), .B(n19930), .Z(n20256) );
  NANDN U20709 ( .A(n19932), .B(n35311), .Z(n19934) );
  XOR U20710 ( .A(b[31]), .B(n29868), .Z(n20319) );
  NANDN U20711 ( .A(n20319), .B(n35313), .Z(n19933) );
  AND U20712 ( .A(n19934), .B(n19933), .Z(n20255) );
  XNOR U20713 ( .A(n20256), .B(n20255), .Z(n20257) );
  XNOR U20714 ( .A(n20258), .B(n20257), .Z(n20219) );
  XOR U20715 ( .A(n20218), .B(n20219), .Z(n20273) );
  XNOR U20716 ( .A(b[37]), .B(a[62]), .Z(n20285) );
  NANDN U20717 ( .A(n20285), .B(n36311), .Z(n19937) );
  NANDN U20718 ( .A(n19935), .B(n36309), .Z(n19936) );
  NAND U20719 ( .A(n19937), .B(n19936), .Z(n20365) );
  XOR U20720 ( .A(a[94]), .B(n968), .Z(n20288) );
  OR U20721 ( .A(n20288), .B(n29363), .Z(n19940) );
  NANDN U20722 ( .A(n19938), .B(n29864), .Z(n19939) );
  NAND U20723 ( .A(n19940), .B(n19939), .Z(n20362) );
  XOR U20724 ( .A(n35545), .B(n967), .Z(n20291) );
  NAND U20725 ( .A(n20291), .B(n28939), .Z(n19943) );
  NAND U20726 ( .A(n28938), .B(n19941), .Z(n19942) );
  AND U20727 ( .A(n19943), .B(n19942), .Z(n20363) );
  XNOR U20728 ( .A(n20362), .B(n20363), .Z(n20364) );
  XNOR U20729 ( .A(n20365), .B(n20364), .Z(n20374) );
  XOR U20730 ( .A(a[86]), .B(n971), .Z(n20294) );
  OR U20731 ( .A(n20294), .B(n31550), .Z(n19946) );
  NANDN U20732 ( .A(n19944), .B(n31874), .Z(n19945) );
  NAND U20733 ( .A(n19946), .B(n19945), .Z(n20207) );
  NAND U20734 ( .A(n34848), .B(n19947), .Z(n19949) );
  XOR U20735 ( .A(n35375), .B(n30210), .Z(n20297) );
  NAND U20736 ( .A(n34618), .B(n20297), .Z(n19948) );
  NAND U20737 ( .A(n19949), .B(n19948), .Z(n20204) );
  NAND U20738 ( .A(n35188), .B(n19950), .Z(n19952) );
  XOR U20739 ( .A(n35540), .B(n30379), .Z(n20300) );
  NANDN U20740 ( .A(n34968), .B(n20300), .Z(n19951) );
  AND U20741 ( .A(n19952), .B(n19951), .Z(n20205) );
  XNOR U20742 ( .A(n20204), .B(n20205), .Z(n20206) );
  XOR U20743 ( .A(n20207), .B(n20206), .Z(n20375) );
  XOR U20744 ( .A(n20374), .B(n20375), .Z(n20377) );
  NANDN U20745 ( .A(n19954), .B(n19953), .Z(n19958) );
  NAND U20746 ( .A(n19956), .B(n19955), .Z(n19957) );
  NAND U20747 ( .A(n19958), .B(n19957), .Z(n20376) );
  XOR U20748 ( .A(n20377), .B(n20376), .Z(n20274) );
  XNOR U20749 ( .A(n20273), .B(n20274), .Z(n20275) );
  XOR U20750 ( .A(n20276), .B(n20275), .Z(n20270) );
  NANDN U20751 ( .A(n19960), .B(n19959), .Z(n19964) );
  NAND U20752 ( .A(n19962), .B(n19961), .Z(n19963) );
  NAND U20753 ( .A(n19964), .B(n19963), .Z(n20177) );
  XNOR U20754 ( .A(b[41]), .B(a[58]), .Z(n20337) );
  OR U20755 ( .A(n20337), .B(n36905), .Z(n19967) );
  NANDN U20756 ( .A(n19965), .B(n36807), .Z(n19966) );
  NAND U20757 ( .A(n19967), .B(n19966), .Z(n20359) );
  XOR U20758 ( .A(b[57]), .B(n22246), .Z(n20340) );
  OR U20759 ( .A(n20340), .B(n965), .Z(n19970) );
  NANDN U20760 ( .A(n19968), .B(n38194), .Z(n19969) );
  NAND U20761 ( .A(n19970), .B(n19969), .Z(n20356) );
  NAND U20762 ( .A(n38326), .B(n19971), .Z(n19973) );
  XOR U20763 ( .A(n38400), .B(n21149), .Z(n20343) );
  NANDN U20764 ( .A(n38273), .B(n20343), .Z(n19972) );
  AND U20765 ( .A(n19973), .B(n19972), .Z(n20357) );
  XNOR U20766 ( .A(n20356), .B(n20357), .Z(n20358) );
  XNOR U20767 ( .A(n20359), .B(n20358), .Z(n20174) );
  XOR U20768 ( .A(b[33]), .B(n28701), .Z(n20346) );
  NANDN U20769 ( .A(n20346), .B(n35620), .Z(n19976) );
  NANDN U20770 ( .A(n19974), .B(n35621), .Z(n19975) );
  NAND U20771 ( .A(n19976), .B(n19975), .Z(n20183) );
  NANDN U20772 ( .A(n966), .B(a[98]), .Z(n19977) );
  XOR U20773 ( .A(n29232), .B(n19977), .Z(n19979) );
  NANDN U20774 ( .A(b[0]), .B(a[97]), .Z(n19978) );
  AND U20775 ( .A(n19979), .B(n19978), .Z(n20180) );
  XOR U20776 ( .A(b[63]), .B(n19980), .Z(n20353) );
  NANDN U20777 ( .A(n20353), .B(n38422), .Z(n19983) );
  NANDN U20778 ( .A(n19981), .B(n38423), .Z(n19982) );
  AND U20779 ( .A(n19983), .B(n19982), .Z(n20181) );
  XNOR U20780 ( .A(n20180), .B(n20181), .Z(n20182) );
  XOR U20781 ( .A(n20183), .B(n20182), .Z(n20175) );
  XNOR U20782 ( .A(n20174), .B(n20175), .Z(n20176) );
  XOR U20783 ( .A(n20177), .B(n20176), .Z(n20389) );
  NANDN U20784 ( .A(n19985), .B(n19984), .Z(n19989) );
  NAND U20785 ( .A(n19987), .B(n19986), .Z(n19988) );
  NAND U20786 ( .A(n19989), .B(n19988), .Z(n20386) );
  NANDN U20787 ( .A(n19991), .B(n19990), .Z(n19995) );
  NAND U20788 ( .A(n19993), .B(n19992), .Z(n19994) );
  AND U20789 ( .A(n19995), .B(n19994), .Z(n20387) );
  XNOR U20790 ( .A(n20386), .B(n20387), .Z(n20388) );
  XNOR U20791 ( .A(n20389), .B(n20388), .Z(n20267) );
  NANDN U20792 ( .A(n19997), .B(n19996), .Z(n20001) );
  OR U20793 ( .A(n19999), .B(n19998), .Z(n20000) );
  AND U20794 ( .A(n20001), .B(n20000), .Z(n20268) );
  XNOR U20795 ( .A(n20267), .B(n20268), .Z(n20269) );
  XNOR U20796 ( .A(n20270), .B(n20269), .Z(n20165) );
  XOR U20797 ( .A(n20164), .B(n20165), .Z(n20416) );
  OR U20798 ( .A(n20003), .B(n20002), .Z(n20007) );
  NAND U20799 ( .A(n20005), .B(n20004), .Z(n20006) );
  NAND U20800 ( .A(n20007), .B(n20006), .Z(n20395) );
  XOR U20801 ( .A(b[35]), .B(a[64]), .Z(n20246) );
  NAND U20802 ( .A(n35985), .B(n20246), .Z(n20010) );
  NAND U20803 ( .A(n20008), .B(n35986), .Z(n20009) );
  NAND U20804 ( .A(n20010), .B(n20009), .Z(n20213) );
  XOR U20805 ( .A(n34852), .B(n31123), .Z(n20249) );
  NAND U20806 ( .A(n20249), .B(n29949), .Z(n20013) );
  NAND U20807 ( .A(n29948), .B(n20011), .Z(n20012) );
  NAND U20808 ( .A(n20013), .B(n20012), .Z(n20210) );
  XOR U20809 ( .A(b[55]), .B(n22289), .Z(n20252) );
  NANDN U20810 ( .A(n20252), .B(n38075), .Z(n20016) );
  NANDN U20811 ( .A(n20014), .B(n38073), .Z(n20015) );
  AND U20812 ( .A(n20016), .B(n20015), .Z(n20211) );
  XNOR U20813 ( .A(n20210), .B(n20211), .Z(n20212) );
  XNOR U20814 ( .A(n20213), .B(n20212), .Z(n20383) );
  NANDN U20815 ( .A(n20018), .B(n20017), .Z(n20022) );
  NANDN U20816 ( .A(n20020), .B(n20019), .Z(n20021) );
  NAND U20817 ( .A(n20022), .B(n20021), .Z(n20380) );
  OR U20818 ( .A(n20024), .B(n20023), .Z(n20028) );
  NANDN U20819 ( .A(n20026), .B(n20025), .Z(n20027) );
  NAND U20820 ( .A(n20028), .B(n20027), .Z(n20381) );
  XNOR U20821 ( .A(n20380), .B(n20381), .Z(n20382) );
  XOR U20822 ( .A(n20383), .B(n20382), .Z(n20400) );
  XOR U20823 ( .A(a[88]), .B(n970), .Z(n20222) );
  OR U20824 ( .A(n20222), .B(n31369), .Z(n20031) );
  NANDN U20825 ( .A(n20029), .B(n31119), .Z(n20030) );
  NAND U20826 ( .A(n20031), .B(n20030), .Z(n20243) );
  XOR U20827 ( .A(b[43]), .B(n25860), .Z(n20225) );
  NANDN U20828 ( .A(n20225), .B(n37068), .Z(n20034) );
  NANDN U20829 ( .A(n20032), .B(n37069), .Z(n20033) );
  NAND U20830 ( .A(n20034), .B(n20033), .Z(n20240) );
  XNOR U20831 ( .A(b[45]), .B(a[54]), .Z(n20228) );
  NANDN U20832 ( .A(n20228), .B(n37261), .Z(n20037) );
  NANDN U20833 ( .A(n20035), .B(n37262), .Z(n20036) );
  AND U20834 ( .A(n20037), .B(n20036), .Z(n20241) );
  XNOR U20835 ( .A(n20240), .B(n20241), .Z(n20242) );
  XNOR U20836 ( .A(n20243), .B(n20242), .Z(n20279) );
  XOR U20837 ( .A(b[49]), .B(n24671), .Z(n20231) );
  OR U20838 ( .A(n20231), .B(n37756), .Z(n20040) );
  NANDN U20839 ( .A(n20038), .B(n37652), .Z(n20039) );
  NAND U20840 ( .A(n20040), .B(n20039), .Z(n20264) );
  NAND U20841 ( .A(n37469), .B(n20041), .Z(n20043) );
  XOR U20842 ( .A(n978), .B(n25134), .Z(n20234) );
  NAND U20843 ( .A(n20234), .B(n37471), .Z(n20042) );
  AND U20844 ( .A(n20043), .B(n20042), .Z(n20261) );
  XOR U20845 ( .A(a[90]), .B(n969), .Z(n20237) );
  NANDN U20846 ( .A(n20237), .B(n30509), .Z(n20046) );
  NANDN U20847 ( .A(n20044), .B(n30846), .Z(n20045) );
  AND U20848 ( .A(n20046), .B(n20045), .Z(n20262) );
  XOR U20849 ( .A(n20264), .B(n20263), .Z(n20280) );
  XNOR U20850 ( .A(n20279), .B(n20280), .Z(n20281) );
  NANDN U20851 ( .A(n20048), .B(n20047), .Z(n20052) );
  NAND U20852 ( .A(n20050), .B(n20049), .Z(n20051) );
  AND U20853 ( .A(n20052), .B(n20051), .Z(n20282) );
  XNOR U20854 ( .A(n20281), .B(n20282), .Z(n20399) );
  NANDN U20855 ( .A(n20054), .B(n20053), .Z(n20058) );
  NANDN U20856 ( .A(n20056), .B(n20055), .Z(n20057) );
  AND U20857 ( .A(n20058), .B(n20057), .Z(n20398) );
  XNOR U20858 ( .A(n20399), .B(n20398), .Z(n20401) );
  XOR U20859 ( .A(n20400), .B(n20401), .Z(n20392) );
  OR U20860 ( .A(n20060), .B(n20059), .Z(n20064) );
  OR U20861 ( .A(n20062), .B(n20061), .Z(n20063) );
  NAND U20862 ( .A(n20064), .B(n20063), .Z(n20410) );
  NANDN U20863 ( .A(n20066), .B(n20065), .Z(n20070) );
  NAND U20864 ( .A(n20068), .B(n20067), .Z(n20069) );
  NAND U20865 ( .A(n20070), .B(n20069), .Z(n20411) );
  XNOR U20866 ( .A(n20410), .B(n20411), .Z(n20412) );
  NANDN U20867 ( .A(n20072), .B(n20071), .Z(n20076) );
  NAND U20868 ( .A(n20074), .B(n20073), .Z(n20075) );
  NAND U20869 ( .A(n20076), .B(n20075), .Z(n20171) );
  XOR U20870 ( .A(b[39]), .B(n27436), .Z(n20195) );
  NANDN U20871 ( .A(n20195), .B(n36553), .Z(n20079) );
  NANDN U20872 ( .A(n20077), .B(n36643), .Z(n20078) );
  NAND U20873 ( .A(n20079), .B(n20078), .Z(n20306) );
  XOR U20874 ( .A(b[51]), .B(n23447), .Z(n20198) );
  NANDN U20875 ( .A(n20198), .B(n37803), .Z(n20082) );
  NANDN U20876 ( .A(n20080), .B(n37802), .Z(n20081) );
  NAND U20877 ( .A(n20082), .B(n20081), .Z(n20303) );
  XOR U20878 ( .A(b[53]), .B(n22964), .Z(n20201) );
  NANDN U20879 ( .A(n20201), .B(n37940), .Z(n20085) );
  NANDN U20880 ( .A(n20083), .B(n37941), .Z(n20084) );
  AND U20881 ( .A(n20085), .B(n20084), .Z(n20304) );
  XNOR U20882 ( .A(n20303), .B(n20304), .Z(n20305) );
  XNOR U20883 ( .A(n20306), .B(n20305), .Z(n20368) );
  XOR U20884 ( .A(a[84]), .B(n972), .Z(n20186) );
  OR U20885 ( .A(n20186), .B(n32010), .Z(n20088) );
  NANDN U20886 ( .A(n20086), .B(n32011), .Z(n20087) );
  NAND U20887 ( .A(n20088), .B(n20087), .Z(n20312) );
  XNOR U20888 ( .A(b[25]), .B(n31372), .Z(n20189) );
  NANDN U20889 ( .A(n34219), .B(n20189), .Z(n20091) );
  NAND U20890 ( .A(n34217), .B(n20089), .Z(n20090) );
  NAND U20891 ( .A(n20091), .B(n20090), .Z(n20309) );
  XNOR U20892 ( .A(a[82]), .B(b[17]), .Z(n20192) );
  NANDN U20893 ( .A(n20192), .B(n32543), .Z(n20094) );
  NAND U20894 ( .A(n20092), .B(n32541), .Z(n20093) );
  AND U20895 ( .A(n20094), .B(n20093), .Z(n20310) );
  XNOR U20896 ( .A(n20309), .B(n20310), .Z(n20311) );
  XOR U20897 ( .A(n20312), .B(n20311), .Z(n20369) );
  XNOR U20898 ( .A(n20368), .B(n20369), .Z(n20370) );
  NANDN U20899 ( .A(n20096), .B(n20095), .Z(n20100) );
  NAND U20900 ( .A(n20098), .B(n20097), .Z(n20099) );
  AND U20901 ( .A(n20100), .B(n20099), .Z(n20371) );
  XNOR U20902 ( .A(n20370), .B(n20371), .Z(n20169) );
  NANDN U20903 ( .A(n20102), .B(n20101), .Z(n20106) );
  NAND U20904 ( .A(n20104), .B(n20103), .Z(n20105) );
  AND U20905 ( .A(n20106), .B(n20105), .Z(n20168) );
  XNOR U20906 ( .A(n20169), .B(n20168), .Z(n20170) );
  XOR U20907 ( .A(n20171), .B(n20170), .Z(n20413) );
  XNOR U20908 ( .A(n20412), .B(n20413), .Z(n20393) );
  XOR U20909 ( .A(n20392), .B(n20393), .Z(n20394) );
  XOR U20910 ( .A(n20395), .B(n20394), .Z(n20417) );
  XNOR U20911 ( .A(n20416), .B(n20417), .Z(n20418) );
  OR U20912 ( .A(n20108), .B(n20107), .Z(n20112) );
  NANDN U20913 ( .A(n20110), .B(n20109), .Z(n20111) );
  NAND U20914 ( .A(n20112), .B(n20111), .Z(n20419) );
  XOR U20915 ( .A(n20418), .B(n20419), .Z(n20431) );
  NANDN U20916 ( .A(n20114), .B(n20113), .Z(n20118) );
  NAND U20917 ( .A(n20116), .B(n20115), .Z(n20117) );
  NAND U20918 ( .A(n20118), .B(n20117), .Z(n20425) );
  XNOR U20919 ( .A(n20423), .B(n20422), .Z(n20424) );
  XOR U20920 ( .A(n20425), .B(n20424), .Z(n20428) );
  NANDN U20921 ( .A(n20128), .B(n20127), .Z(n20132) );
  NAND U20922 ( .A(n20130), .B(n20129), .Z(n20131) );
  AND U20923 ( .A(n20132), .B(n20131), .Z(n20429) );
  XNOR U20924 ( .A(n20428), .B(n20429), .Z(n20430) );
  XNOR U20925 ( .A(n20431), .B(n20430), .Z(n20437) );
  XOR U20926 ( .A(n20436), .B(n20437), .Z(n20440) );
  NANDN U20927 ( .A(n20134), .B(n20133), .Z(n20138) );
  NAND U20928 ( .A(n20136), .B(n20135), .Z(n20137) );
  NAND U20929 ( .A(n20138), .B(n20137), .Z(n20441) );
  XNOR U20930 ( .A(n20440), .B(n20441), .Z(n20442) );
  NANDN U20931 ( .A(n20140), .B(n20139), .Z(n20144) );
  NANDN U20932 ( .A(n20142), .B(n20141), .Z(n20143) );
  NAND U20933 ( .A(n20144), .B(n20143), .Z(n20443) );
  XOR U20934 ( .A(n20442), .B(n20443), .Z(n20156) );
  NANDN U20935 ( .A(n20146), .B(n20145), .Z(n20150) );
  NANDN U20936 ( .A(n20148), .B(n20147), .Z(n20149) );
  NAND U20937 ( .A(n20150), .B(n20149), .Z(n20157) );
  XNOR U20938 ( .A(n20156), .B(n20157), .Z(n20158) );
  XNOR U20939 ( .A(n20159), .B(n20158), .Z(n20446) );
  XNOR U20940 ( .A(n20446), .B(sreg[162]), .Z(n20448) );
  NAND U20941 ( .A(n20151), .B(sreg[161]), .Z(n20155) );
  OR U20942 ( .A(n20153), .B(n20152), .Z(n20154) );
  AND U20943 ( .A(n20155), .B(n20154), .Z(n20447) );
  XOR U20944 ( .A(n20448), .B(n20447), .Z(c[162]) );
  NANDN U20945 ( .A(n20157), .B(n20156), .Z(n20161) );
  NAND U20946 ( .A(n20159), .B(n20158), .Z(n20160) );
  NAND U20947 ( .A(n20161), .B(n20160), .Z(n20454) );
  NANDN U20948 ( .A(n20163), .B(n20162), .Z(n20167) );
  NANDN U20949 ( .A(n20165), .B(n20164), .Z(n20166) );
  NAND U20950 ( .A(n20167), .B(n20166), .Z(n20460) );
  NANDN U20951 ( .A(n20169), .B(n20168), .Z(n20173) );
  NANDN U20952 ( .A(n20171), .B(n20170), .Z(n20172) );
  NAND U20953 ( .A(n20173), .B(n20172), .Z(n20702) );
  NANDN U20954 ( .A(n20175), .B(n20174), .Z(n20179) );
  NANDN U20955 ( .A(n20177), .B(n20176), .Z(n20178) );
  AND U20956 ( .A(n20179), .B(n20178), .Z(n20703) );
  XNOR U20957 ( .A(n20702), .B(n20703), .Z(n20704) );
  NANDN U20958 ( .A(n20181), .B(n20180), .Z(n20185) );
  NAND U20959 ( .A(n20183), .B(n20182), .Z(n20184) );
  NAND U20960 ( .A(n20185), .B(n20184), .Z(n20529) );
  XNOR U20961 ( .A(a[85]), .B(b[15]), .Z(n20541) );
  OR U20962 ( .A(n20541), .B(n32010), .Z(n20188) );
  NANDN U20963 ( .A(n20186), .B(n32011), .Z(n20187) );
  NAND U20964 ( .A(n20188), .B(n20187), .Z(n20635) );
  XOR U20965 ( .A(b[25]), .B(a[75]), .Z(n20544) );
  NANDN U20966 ( .A(n34219), .B(n20544), .Z(n20191) );
  NAND U20967 ( .A(n34217), .B(n20189), .Z(n20190) );
  NAND U20968 ( .A(n20191), .B(n20190), .Z(n20632) );
  XOR U20969 ( .A(a[83]), .B(b[17]), .Z(n20547) );
  NAND U20970 ( .A(n20547), .B(n32543), .Z(n20194) );
  NANDN U20971 ( .A(n20192), .B(n32541), .Z(n20193) );
  AND U20972 ( .A(n20194), .B(n20193), .Z(n20633) );
  XNOR U20973 ( .A(n20632), .B(n20633), .Z(n20634) );
  XNOR U20974 ( .A(n20635), .B(n20634), .Z(n20653) );
  XOR U20975 ( .A(b[39]), .B(n27773), .Z(n20532) );
  NANDN U20976 ( .A(n20532), .B(n36553), .Z(n20197) );
  NANDN U20977 ( .A(n20195), .B(n36643), .Z(n20196) );
  NAND U20978 ( .A(n20197), .B(n20196), .Z(n20629) );
  XOR U20979 ( .A(b[51]), .B(n23852), .Z(n20535) );
  NANDN U20980 ( .A(n20535), .B(n37803), .Z(n20200) );
  NANDN U20981 ( .A(n20198), .B(n37802), .Z(n20199) );
  NAND U20982 ( .A(n20200), .B(n20199), .Z(n20626) );
  XOR U20983 ( .A(b[53]), .B(n23149), .Z(n20538) );
  NANDN U20984 ( .A(n20538), .B(n37940), .Z(n20203) );
  NANDN U20985 ( .A(n20201), .B(n37941), .Z(n20202) );
  AND U20986 ( .A(n20203), .B(n20202), .Z(n20627) );
  XNOR U20987 ( .A(n20626), .B(n20627), .Z(n20628) );
  XOR U20988 ( .A(n20629), .B(n20628), .Z(n20654) );
  XNOR U20989 ( .A(n20653), .B(n20654), .Z(n20655) );
  NANDN U20990 ( .A(n20205), .B(n20204), .Z(n20209) );
  NAND U20991 ( .A(n20207), .B(n20206), .Z(n20208) );
  AND U20992 ( .A(n20209), .B(n20208), .Z(n20656) );
  XNOR U20993 ( .A(n20655), .B(n20656), .Z(n20527) );
  NANDN U20994 ( .A(n20211), .B(n20210), .Z(n20215) );
  NAND U20995 ( .A(n20213), .B(n20212), .Z(n20214) );
  AND U20996 ( .A(n20215), .B(n20214), .Z(n20526) );
  XNOR U20997 ( .A(n20527), .B(n20526), .Z(n20528) );
  XOR U20998 ( .A(n20529), .B(n20528), .Z(n20705) );
  XOR U20999 ( .A(n20704), .B(n20705), .Z(n20714) );
  NANDN U21000 ( .A(n20217), .B(n20216), .Z(n20221) );
  NANDN U21001 ( .A(n20219), .B(n20218), .Z(n20220) );
  NAND U21002 ( .A(n20221), .B(n20220), .Z(n20696) );
  XNOR U21003 ( .A(a[89]), .B(b[11]), .Z(n20475) );
  OR U21004 ( .A(n20475), .B(n31369), .Z(n20224) );
  NANDN U21005 ( .A(n20222), .B(n31119), .Z(n20223) );
  NAND U21006 ( .A(n20224), .B(n20223), .Z(n20496) );
  XOR U21007 ( .A(b[43]), .B(n26122), .Z(n20478) );
  NANDN U21008 ( .A(n20478), .B(n37068), .Z(n20227) );
  NANDN U21009 ( .A(n20225), .B(n37069), .Z(n20226) );
  NAND U21010 ( .A(n20227), .B(n20226), .Z(n20493) );
  XNOR U21011 ( .A(b[45]), .B(a[55]), .Z(n20481) );
  NANDN U21012 ( .A(n20481), .B(n37261), .Z(n20230) );
  NANDN U21013 ( .A(n20228), .B(n37262), .Z(n20229) );
  AND U21014 ( .A(n20230), .B(n20229), .Z(n20494) );
  XNOR U21015 ( .A(n20493), .B(n20494), .Z(n20495) );
  XNOR U21016 ( .A(n20496), .B(n20495), .Z(n20602) );
  XOR U21017 ( .A(b[49]), .B(n24288), .Z(n20484) );
  OR U21018 ( .A(n20484), .B(n37756), .Z(n20233) );
  NANDN U21019 ( .A(n20231), .B(n37652), .Z(n20232) );
  NAND U21020 ( .A(n20233), .B(n20232), .Z(n20523) );
  NAND U21021 ( .A(n37469), .B(n20234), .Z(n20236) );
  XOR U21022 ( .A(n978), .B(n25001), .Z(n20487) );
  NAND U21023 ( .A(n20487), .B(n37471), .Z(n20235) );
  NAND U21024 ( .A(n20236), .B(n20235), .Z(n20520) );
  XNOR U21025 ( .A(a[91]), .B(b[9]), .Z(n20490) );
  NANDN U21026 ( .A(n20490), .B(n30509), .Z(n20239) );
  NANDN U21027 ( .A(n20237), .B(n30846), .Z(n20238) );
  AND U21028 ( .A(n20239), .B(n20238), .Z(n20521) );
  XNOR U21029 ( .A(n20520), .B(n20521), .Z(n20522) );
  XOR U21030 ( .A(n20523), .B(n20522), .Z(n20603) );
  XNOR U21031 ( .A(n20602), .B(n20603), .Z(n20604) );
  NANDN U21032 ( .A(n20241), .B(n20240), .Z(n20245) );
  NAND U21033 ( .A(n20243), .B(n20242), .Z(n20244) );
  AND U21034 ( .A(n20245), .B(n20244), .Z(n20605) );
  XNOR U21035 ( .A(n20604), .B(n20605), .Z(n20697) );
  XNOR U21036 ( .A(n20696), .B(n20697), .Z(n20698) );
  XNOR U21037 ( .A(b[35]), .B(a[65]), .Z(n20505) );
  NANDN U21038 ( .A(n20505), .B(n35985), .Z(n20248) );
  NAND U21039 ( .A(n20246), .B(n35986), .Z(n20247) );
  NAND U21040 ( .A(n20248), .B(n20247), .Z(n20559) );
  XOR U21041 ( .A(n35377), .B(n31123), .Z(n20508) );
  NAND U21042 ( .A(n20508), .B(n29949), .Z(n20251) );
  NAND U21043 ( .A(n29948), .B(n20249), .Z(n20250) );
  NAND U21044 ( .A(n20251), .B(n20250), .Z(n20556) );
  XOR U21045 ( .A(b[55]), .B(n22579), .Z(n20511) );
  NANDN U21046 ( .A(n20511), .B(n38075), .Z(n20254) );
  NANDN U21047 ( .A(n20252), .B(n38073), .Z(n20253) );
  AND U21048 ( .A(n20254), .B(n20253), .Z(n20557) );
  XNOR U21049 ( .A(n20556), .B(n20557), .Z(n20558) );
  XNOR U21050 ( .A(n20559), .B(n20558), .Z(n20587) );
  NANDN U21051 ( .A(n20256), .B(n20255), .Z(n20260) );
  NAND U21052 ( .A(n20258), .B(n20257), .Z(n20259) );
  NAND U21053 ( .A(n20260), .B(n20259), .Z(n20584) );
  OR U21054 ( .A(n20262), .B(n20261), .Z(n20266) );
  NAND U21055 ( .A(n20264), .B(n20263), .Z(n20265) );
  NAND U21056 ( .A(n20266), .B(n20265), .Z(n20585) );
  XNOR U21057 ( .A(n20584), .B(n20585), .Z(n20586) );
  XOR U21058 ( .A(n20587), .B(n20586), .Z(n20699) );
  XOR U21059 ( .A(n20698), .B(n20699), .Z(n20715) );
  XNOR U21060 ( .A(n20714), .B(n20715), .Z(n20716) );
  NANDN U21061 ( .A(n20268), .B(n20267), .Z(n20272) );
  NAND U21062 ( .A(n20270), .B(n20269), .Z(n20271) );
  NAND U21063 ( .A(n20272), .B(n20271), .Z(n20717) );
  XOR U21064 ( .A(n20716), .B(n20717), .Z(n20458) );
  NANDN U21065 ( .A(n20274), .B(n20273), .Z(n20278) );
  NANDN U21066 ( .A(n20276), .B(n20275), .Z(n20277) );
  NAND U21067 ( .A(n20278), .B(n20277), .Z(n20469) );
  NANDN U21068 ( .A(n20280), .B(n20279), .Z(n20284) );
  NAND U21069 ( .A(n20282), .B(n20281), .Z(n20283) );
  NAND U21070 ( .A(n20284), .B(n20283), .Z(n20599) );
  XNOR U21071 ( .A(b[37]), .B(a[63]), .Z(n20608) );
  NANDN U21072 ( .A(n20608), .B(n36311), .Z(n20287) );
  NANDN U21073 ( .A(n20285), .B(n36309), .Z(n20286) );
  NAND U21074 ( .A(n20287), .B(n20286), .Z(n20662) );
  XOR U21075 ( .A(a[95]), .B(n968), .Z(n20611) );
  OR U21076 ( .A(n20611), .B(n29363), .Z(n20290) );
  NANDN U21077 ( .A(n20288), .B(n29864), .Z(n20289) );
  NAND U21078 ( .A(n20290), .B(n20289), .Z(n20659) );
  XNOR U21079 ( .A(a[97]), .B(n967), .Z(n20614) );
  NAND U21080 ( .A(n20614), .B(n28939), .Z(n20293) );
  NAND U21081 ( .A(n28938), .B(n20291), .Z(n20292) );
  AND U21082 ( .A(n20293), .B(n20292), .Z(n20660) );
  XNOR U21083 ( .A(n20659), .B(n20660), .Z(n20661) );
  XNOR U21084 ( .A(n20662), .B(n20661), .Z(n20578) );
  XNOR U21085 ( .A(a[87]), .B(b[13]), .Z(n20617) );
  OR U21086 ( .A(n20617), .B(n31550), .Z(n20296) );
  NANDN U21087 ( .A(n20294), .B(n31874), .Z(n20295) );
  NAND U21088 ( .A(n20296), .B(n20295), .Z(n20553) );
  NAND U21089 ( .A(n34848), .B(n20297), .Z(n20299) );
  XNOR U21090 ( .A(n35375), .B(a[73]), .Z(n20620) );
  NAND U21091 ( .A(n34618), .B(n20620), .Z(n20298) );
  NAND U21092 ( .A(n20299), .B(n20298), .Z(n20550) );
  NAND U21093 ( .A(n35188), .B(n20300), .Z(n20302) );
  XOR U21094 ( .A(n35540), .B(n30543), .Z(n20623) );
  NANDN U21095 ( .A(n34968), .B(n20623), .Z(n20301) );
  AND U21096 ( .A(n20302), .B(n20301), .Z(n20551) );
  XNOR U21097 ( .A(n20550), .B(n20551), .Z(n20552) );
  XOR U21098 ( .A(n20553), .B(n20552), .Z(n20579) );
  XNOR U21099 ( .A(n20578), .B(n20579), .Z(n20580) );
  NANDN U21100 ( .A(n20304), .B(n20303), .Z(n20308) );
  NAND U21101 ( .A(n20306), .B(n20305), .Z(n20307) );
  NAND U21102 ( .A(n20308), .B(n20307), .Z(n20581) );
  XOR U21103 ( .A(n20580), .B(n20581), .Z(n20596) );
  NANDN U21104 ( .A(n20310), .B(n20309), .Z(n20314) );
  NAND U21105 ( .A(n20312), .B(n20311), .Z(n20313) );
  NAND U21106 ( .A(n20314), .B(n20313), .Z(n20501) );
  ANDN U21107 ( .B(b[63]), .A(n20315), .Z(n20517) );
  NANDN U21108 ( .A(n20316), .B(n38369), .Z(n20318) );
  XOR U21109 ( .A(b[61]), .B(n20867), .Z(n20638) );
  OR U21110 ( .A(n20638), .B(n38371), .Z(n20317) );
  NAND U21111 ( .A(n20318), .B(n20317), .Z(n20515) );
  NANDN U21112 ( .A(n20319), .B(n35311), .Z(n20321) );
  XNOR U21113 ( .A(b[31]), .B(a[69]), .Z(n20641) );
  NANDN U21114 ( .A(n20641), .B(n35313), .Z(n20320) );
  AND U21115 ( .A(n20321), .B(n20320), .Z(n20514) );
  XNOR U21116 ( .A(n20515), .B(n20514), .Z(n20516) );
  XOR U21117 ( .A(n20517), .B(n20516), .Z(n20499) );
  NAND U21118 ( .A(n33283), .B(n20322), .Z(n20324) );
  XNOR U21119 ( .A(n33020), .B(a[81]), .Z(n20644) );
  NANDN U21120 ( .A(n33021), .B(n20644), .Z(n20323) );
  NAND U21121 ( .A(n20324), .B(n20323), .Z(n20668) );
  XOR U21122 ( .A(b[21]), .B(a[79]), .Z(n20647) );
  NANDN U21123 ( .A(n33634), .B(n20647), .Z(n20327) );
  NANDN U21124 ( .A(n20325), .B(n33464), .Z(n20326) );
  NAND U21125 ( .A(n20327), .B(n20326), .Z(n20665) );
  NAND U21126 ( .A(n34044), .B(n20328), .Z(n20330) );
  XNOR U21127 ( .A(n34510), .B(a[77]), .Z(n20650) );
  NANDN U21128 ( .A(n33867), .B(n20650), .Z(n20329) );
  AND U21129 ( .A(n20330), .B(n20329), .Z(n20666) );
  XNOR U21130 ( .A(n20665), .B(n20666), .Z(n20667) );
  XNOR U21131 ( .A(n20668), .B(n20667), .Z(n20500) );
  XOR U21132 ( .A(n20499), .B(n20500), .Z(n20502) );
  XOR U21133 ( .A(n20501), .B(n20502), .Z(n20597) );
  XNOR U21134 ( .A(n20596), .B(n20597), .Z(n20598) );
  XOR U21135 ( .A(n20599), .B(n20598), .Z(n20577) );
  NANDN U21136 ( .A(n20332), .B(n20331), .Z(n20336) );
  NAND U21137 ( .A(n20334), .B(n20333), .Z(n20335) );
  NAND U21138 ( .A(n20336), .B(n20335), .Z(n20571) );
  XOR U21139 ( .A(b[41]), .B(a[59]), .Z(n20671) );
  NANDN U21140 ( .A(n36905), .B(n20671), .Z(n20339) );
  NANDN U21141 ( .A(n20337), .B(n36807), .Z(n20338) );
  NAND U21142 ( .A(n20339), .B(n20338), .Z(n20693) );
  XOR U21143 ( .A(b[57]), .B(n21996), .Z(n20674) );
  OR U21144 ( .A(n20674), .B(n965), .Z(n20342) );
  NANDN U21145 ( .A(n20340), .B(n38194), .Z(n20341) );
  NAND U21146 ( .A(n20342), .B(n20341), .Z(n20690) );
  NAND U21147 ( .A(n38326), .B(n20343), .Z(n20345) );
  XOR U21148 ( .A(n38400), .B(n21441), .Z(n20677) );
  NANDN U21149 ( .A(n38273), .B(n20677), .Z(n20344) );
  AND U21150 ( .A(n20345), .B(n20344), .Z(n20691) );
  XNOR U21151 ( .A(n20690), .B(n20691), .Z(n20692) );
  XNOR U21152 ( .A(n20693), .B(n20692), .Z(n20568) );
  XOR U21153 ( .A(b[33]), .B(n29372), .Z(n20680) );
  NANDN U21154 ( .A(n20680), .B(n35620), .Z(n20348) );
  NANDN U21155 ( .A(n20346), .B(n35621), .Z(n20347) );
  NAND U21156 ( .A(n20348), .B(n20347), .Z(n20565) );
  NANDN U21157 ( .A(n966), .B(a[99]), .Z(n20349) );
  XOR U21158 ( .A(n29232), .B(n20349), .Z(n20351) );
  IV U21159 ( .A(a[98]), .Z(n35783) );
  NANDN U21160 ( .A(n35783), .B(n966), .Z(n20350) );
  AND U21161 ( .A(n20351), .B(n20350), .Z(n20562) );
  XOR U21162 ( .A(b[63]), .B(n20352), .Z(n20687) );
  NANDN U21163 ( .A(n20687), .B(n38422), .Z(n20355) );
  NANDN U21164 ( .A(n20353), .B(n38423), .Z(n20354) );
  AND U21165 ( .A(n20355), .B(n20354), .Z(n20563) );
  XNOR U21166 ( .A(n20562), .B(n20563), .Z(n20564) );
  XOR U21167 ( .A(n20565), .B(n20564), .Z(n20569) );
  XNOR U21168 ( .A(n20568), .B(n20569), .Z(n20570) );
  XOR U21169 ( .A(n20571), .B(n20570), .Z(n20593) );
  NANDN U21170 ( .A(n20357), .B(n20356), .Z(n20361) );
  NAND U21171 ( .A(n20359), .B(n20358), .Z(n20360) );
  NAND U21172 ( .A(n20361), .B(n20360), .Z(n20590) );
  NANDN U21173 ( .A(n20363), .B(n20362), .Z(n20367) );
  NAND U21174 ( .A(n20365), .B(n20364), .Z(n20366) );
  AND U21175 ( .A(n20367), .B(n20366), .Z(n20591) );
  XNOR U21176 ( .A(n20590), .B(n20591), .Z(n20592) );
  XNOR U21177 ( .A(n20593), .B(n20592), .Z(n20574) );
  NANDN U21178 ( .A(n20369), .B(n20368), .Z(n20373) );
  NAND U21179 ( .A(n20371), .B(n20370), .Z(n20372) );
  AND U21180 ( .A(n20373), .B(n20372), .Z(n20575) );
  XNOR U21181 ( .A(n20574), .B(n20575), .Z(n20576) );
  XNOR U21182 ( .A(n20577), .B(n20576), .Z(n20470) );
  XOR U21183 ( .A(n20469), .B(n20470), .Z(n20471) );
  NANDN U21184 ( .A(n20375), .B(n20374), .Z(n20379) );
  OR U21185 ( .A(n20377), .B(n20376), .Z(n20378) );
  NAND U21186 ( .A(n20379), .B(n20378), .Z(n20710) );
  NANDN U21187 ( .A(n20381), .B(n20380), .Z(n20385) );
  NAND U21188 ( .A(n20383), .B(n20382), .Z(n20384) );
  AND U21189 ( .A(n20385), .B(n20384), .Z(n20708) );
  NANDN U21190 ( .A(n20387), .B(n20386), .Z(n20391) );
  NAND U21191 ( .A(n20389), .B(n20388), .Z(n20390) );
  NAND U21192 ( .A(n20391), .B(n20390), .Z(n20709) );
  XOR U21193 ( .A(n20710), .B(n20711), .Z(n20472) );
  XNOR U21194 ( .A(n20471), .B(n20472), .Z(n20457) );
  XOR U21195 ( .A(n20458), .B(n20457), .Z(n20459) );
  XNOR U21196 ( .A(n20460), .B(n20459), .Z(n20723) );
  NAND U21197 ( .A(n20393), .B(n20392), .Z(n20397) );
  NAND U21198 ( .A(n20395), .B(n20394), .Z(n20396) );
  NAND U21199 ( .A(n20397), .B(n20396), .Z(n20720) );
  NANDN U21200 ( .A(n20399), .B(n20398), .Z(n20403) );
  NAND U21201 ( .A(n20401), .B(n20400), .Z(n20402) );
  NAND U21202 ( .A(n20403), .B(n20402), .Z(n20466) );
  OR U21203 ( .A(n20405), .B(n20404), .Z(n20409) );
  NAND U21204 ( .A(n20407), .B(n20406), .Z(n20408) );
  NAND U21205 ( .A(n20409), .B(n20408), .Z(n20464) );
  NANDN U21206 ( .A(n20411), .B(n20410), .Z(n20415) );
  NANDN U21207 ( .A(n20413), .B(n20412), .Z(n20414) );
  AND U21208 ( .A(n20415), .B(n20414), .Z(n20463) );
  XNOR U21209 ( .A(n20464), .B(n20463), .Z(n20465) );
  XOR U21210 ( .A(n20466), .B(n20465), .Z(n20721) );
  XOR U21211 ( .A(n20720), .B(n20721), .Z(n20722) );
  XOR U21212 ( .A(n20723), .B(n20722), .Z(n20729) );
  NANDN U21213 ( .A(n20417), .B(n20416), .Z(n20421) );
  NANDN U21214 ( .A(n20419), .B(n20418), .Z(n20420) );
  NAND U21215 ( .A(n20421), .B(n20420), .Z(n20727) );
  NANDN U21216 ( .A(n20423), .B(n20422), .Z(n20427) );
  NANDN U21217 ( .A(n20425), .B(n20424), .Z(n20426) );
  AND U21218 ( .A(n20427), .B(n20426), .Z(n20726) );
  XNOR U21219 ( .A(n20727), .B(n20726), .Z(n20728) );
  XNOR U21220 ( .A(n20729), .B(n20728), .Z(n20732) );
  NANDN U21221 ( .A(n20429), .B(n20428), .Z(n20433) );
  NAND U21222 ( .A(n20431), .B(n20430), .Z(n20432) );
  NAND U21223 ( .A(n20433), .B(n20432), .Z(n20733) );
  XOR U21224 ( .A(n20732), .B(n20733), .Z(n20734) );
  NANDN U21225 ( .A(n20435), .B(n20434), .Z(n20439) );
  NANDN U21226 ( .A(n20437), .B(n20436), .Z(n20438) );
  NAND U21227 ( .A(n20439), .B(n20438), .Z(n20735) );
  XOR U21228 ( .A(n20734), .B(n20735), .Z(n20451) );
  NANDN U21229 ( .A(n20441), .B(n20440), .Z(n20445) );
  NANDN U21230 ( .A(n20443), .B(n20442), .Z(n20444) );
  NAND U21231 ( .A(n20445), .B(n20444), .Z(n20452) );
  XNOR U21232 ( .A(n20451), .B(n20452), .Z(n20453) );
  XNOR U21233 ( .A(n20454), .B(n20453), .Z(n20738) );
  XNOR U21234 ( .A(n20738), .B(sreg[163]), .Z(n20740) );
  NAND U21235 ( .A(n20446), .B(sreg[162]), .Z(n20450) );
  OR U21236 ( .A(n20448), .B(n20447), .Z(n20449) );
  AND U21237 ( .A(n20450), .B(n20449), .Z(n20739) );
  XOR U21238 ( .A(n20740), .B(n20739), .Z(c[163]) );
  NANDN U21239 ( .A(n20452), .B(n20451), .Z(n20456) );
  NAND U21240 ( .A(n20454), .B(n20453), .Z(n20455) );
  NAND U21241 ( .A(n20456), .B(n20455), .Z(n20746) );
  NAND U21242 ( .A(n20458), .B(n20457), .Z(n20462) );
  NAND U21243 ( .A(n20460), .B(n20459), .Z(n20461) );
  NAND U21244 ( .A(n20462), .B(n20461), .Z(n21014) );
  NANDN U21245 ( .A(n20464), .B(n20463), .Z(n20468) );
  NANDN U21246 ( .A(n20466), .B(n20465), .Z(n20467) );
  NAND U21247 ( .A(n20468), .B(n20467), .Z(n21015) );
  XNOR U21248 ( .A(n21014), .B(n21015), .Z(n21016) );
  OR U21249 ( .A(n20470), .B(n20469), .Z(n20474) );
  NANDN U21250 ( .A(n20472), .B(n20471), .Z(n20473) );
  NAND U21251 ( .A(n20474), .B(n20473), .Z(n20751) );
  XOR U21252 ( .A(a[90]), .B(n970), .Z(n20892) );
  OR U21253 ( .A(n20892), .B(n31369), .Z(n20477) );
  NANDN U21254 ( .A(n20475), .B(n31119), .Z(n20476) );
  NAND U21255 ( .A(n20477), .B(n20476), .Z(n20904) );
  XOR U21256 ( .A(b[43]), .B(n26347), .Z(n20895) );
  NANDN U21257 ( .A(n20895), .B(n37068), .Z(n20480) );
  NANDN U21258 ( .A(n20478), .B(n37069), .Z(n20479) );
  NAND U21259 ( .A(n20480), .B(n20479), .Z(n20901) );
  XNOR U21260 ( .A(b[45]), .B(a[56]), .Z(n20898) );
  NANDN U21261 ( .A(n20898), .B(n37261), .Z(n20483) );
  NANDN U21262 ( .A(n20481), .B(n37262), .Z(n20482) );
  AND U21263 ( .A(n20483), .B(n20482), .Z(n20902) );
  XNOR U21264 ( .A(n20901), .B(n20902), .Z(n20903) );
  XNOR U21265 ( .A(n20904), .B(n20903), .Z(n20788) );
  XOR U21266 ( .A(n979), .B(n25134), .Z(n20883) );
  NANDN U21267 ( .A(n37756), .B(n20883), .Z(n20486) );
  NANDN U21268 ( .A(n20484), .B(n37652), .Z(n20485) );
  NAND U21269 ( .A(n20486), .B(n20485), .Z(n20929) );
  NAND U21270 ( .A(n37469), .B(n20487), .Z(n20489) );
  XOR U21271 ( .A(b[47]), .B(n25177), .Z(n20886) );
  NANDN U21272 ( .A(n20886), .B(n37471), .Z(n20488) );
  NAND U21273 ( .A(n20489), .B(n20488), .Z(n20926) );
  XOR U21274 ( .A(n34852), .B(n969), .Z(n20889) );
  NAND U21275 ( .A(n30509), .B(n20889), .Z(n20492) );
  NANDN U21276 ( .A(n20490), .B(n30846), .Z(n20491) );
  AND U21277 ( .A(n20492), .B(n20491), .Z(n20927) );
  XNOR U21278 ( .A(n20926), .B(n20927), .Z(n20928) );
  XNOR U21279 ( .A(n20929), .B(n20928), .Z(n20785) );
  NANDN U21280 ( .A(n20494), .B(n20493), .Z(n20498) );
  NAND U21281 ( .A(n20496), .B(n20495), .Z(n20497) );
  NAND U21282 ( .A(n20498), .B(n20497), .Z(n20786) );
  XNOR U21283 ( .A(n20785), .B(n20786), .Z(n20787) );
  XOR U21284 ( .A(n20788), .B(n20787), .Z(n20996) );
  NANDN U21285 ( .A(n20500), .B(n20499), .Z(n20504) );
  NANDN U21286 ( .A(n20502), .B(n20501), .Z(n20503) );
  AND U21287 ( .A(n20504), .B(n20503), .Z(n20997) );
  XNOR U21288 ( .A(n20996), .B(n20997), .Z(n20999) );
  XNOR U21289 ( .A(b[35]), .B(a[66]), .Z(n20911) );
  NANDN U21290 ( .A(n20911), .B(n35985), .Z(n20507) );
  NANDN U21291 ( .A(n20505), .B(n35986), .Z(n20506) );
  NAND U21292 ( .A(n20507), .B(n20506), .Z(n20959) );
  XOR U21293 ( .A(n35191), .B(n31123), .Z(n20914) );
  NAND U21294 ( .A(n20914), .B(n29949), .Z(n20510) );
  NAND U21295 ( .A(n29948), .B(n20508), .Z(n20509) );
  NAND U21296 ( .A(n20510), .B(n20509), .Z(n20956) );
  XOR U21297 ( .A(b[55]), .B(n22964), .Z(n20917) );
  NANDN U21298 ( .A(n20917), .B(n38075), .Z(n20513) );
  NANDN U21299 ( .A(n20511), .B(n38073), .Z(n20512) );
  AND U21300 ( .A(n20513), .B(n20512), .Z(n20957) );
  XNOR U21301 ( .A(n20956), .B(n20957), .Z(n20958) );
  XNOR U21302 ( .A(n20959), .B(n20958), .Z(n20764) );
  NANDN U21303 ( .A(n20515), .B(n20514), .Z(n20519) );
  NANDN U21304 ( .A(n20517), .B(n20516), .Z(n20518) );
  NAND U21305 ( .A(n20519), .B(n20518), .Z(n20761) );
  NANDN U21306 ( .A(n20521), .B(n20520), .Z(n20525) );
  NAND U21307 ( .A(n20523), .B(n20522), .Z(n20524) );
  NAND U21308 ( .A(n20525), .B(n20524), .Z(n20762) );
  XNOR U21309 ( .A(n20761), .B(n20762), .Z(n20763) );
  XOR U21310 ( .A(n20764), .B(n20763), .Z(n20998) );
  XOR U21311 ( .A(n20999), .B(n20998), .Z(n21002) );
  NANDN U21312 ( .A(n20527), .B(n20526), .Z(n20531) );
  NANDN U21313 ( .A(n20529), .B(n20528), .Z(n20530) );
  NAND U21314 ( .A(n20531), .B(n20530), .Z(n20987) );
  XNOR U21315 ( .A(b[39]), .B(a[62]), .Z(n20941) );
  NANDN U21316 ( .A(n20941), .B(n36553), .Z(n20534) );
  NANDN U21317 ( .A(n20532), .B(n36643), .Z(n20533) );
  NAND U21318 ( .A(n20534), .B(n20533), .Z(n20831) );
  XOR U21319 ( .A(b[51]), .B(n24671), .Z(n20944) );
  NANDN U21320 ( .A(n20944), .B(n37803), .Z(n20537) );
  NANDN U21321 ( .A(n20535), .B(n37802), .Z(n20536) );
  NAND U21322 ( .A(n20537), .B(n20536), .Z(n20828) );
  XOR U21323 ( .A(b[53]), .B(n23447), .Z(n20947) );
  NANDN U21324 ( .A(n20947), .B(n37940), .Z(n20540) );
  NANDN U21325 ( .A(n20538), .B(n37941), .Z(n20539) );
  AND U21326 ( .A(n20540), .B(n20539), .Z(n20829) );
  XNOR U21327 ( .A(n20828), .B(n20829), .Z(n20830) );
  XNOR U21328 ( .A(n20831), .B(n20830), .Z(n20836) );
  XOR U21329 ( .A(a[86]), .B(n972), .Z(n20932) );
  OR U21330 ( .A(n20932), .B(n32010), .Z(n20543) );
  NANDN U21331 ( .A(n20541), .B(n32011), .Z(n20542) );
  NAND U21332 ( .A(n20543), .B(n20542), .Z(n20801) );
  XNOR U21333 ( .A(b[25]), .B(n31363), .Z(n20935) );
  NANDN U21334 ( .A(n34219), .B(n20935), .Z(n20546) );
  NAND U21335 ( .A(n34217), .B(n20544), .Z(n20545) );
  NAND U21336 ( .A(n20546), .B(n20545), .Z(n20798) );
  XNOR U21337 ( .A(a[84]), .B(b[17]), .Z(n20938) );
  NANDN U21338 ( .A(n20938), .B(n32543), .Z(n20549) );
  NAND U21339 ( .A(n20547), .B(n32541), .Z(n20548) );
  AND U21340 ( .A(n20549), .B(n20548), .Z(n20799) );
  XNOR U21341 ( .A(n20798), .B(n20799), .Z(n20800) );
  XNOR U21342 ( .A(n20801), .B(n20800), .Z(n20834) );
  NANDN U21343 ( .A(n20551), .B(n20550), .Z(n20555) );
  NAND U21344 ( .A(n20553), .B(n20552), .Z(n20554) );
  NAND U21345 ( .A(n20555), .B(n20554), .Z(n20835) );
  XOR U21346 ( .A(n20834), .B(n20835), .Z(n20837) );
  XNOR U21347 ( .A(n20836), .B(n20837), .Z(n20975) );
  NANDN U21348 ( .A(n20557), .B(n20556), .Z(n20561) );
  NAND U21349 ( .A(n20559), .B(n20558), .Z(n20560) );
  NAND U21350 ( .A(n20561), .B(n20560), .Z(n20972) );
  NANDN U21351 ( .A(n20563), .B(n20562), .Z(n20567) );
  NAND U21352 ( .A(n20565), .B(n20564), .Z(n20566) );
  AND U21353 ( .A(n20567), .B(n20566), .Z(n20973) );
  XNOR U21354 ( .A(n20972), .B(n20973), .Z(n20974) );
  XNOR U21355 ( .A(n20975), .B(n20974), .Z(n20985) );
  NANDN U21356 ( .A(n20569), .B(n20568), .Z(n20573) );
  NANDN U21357 ( .A(n20571), .B(n20570), .Z(n20572) );
  AND U21358 ( .A(n20573), .B(n20572), .Z(n20984) );
  XOR U21359 ( .A(n20985), .B(n20984), .Z(n20986) );
  XOR U21360 ( .A(n20987), .B(n20986), .Z(n21003) );
  XNOR U21361 ( .A(n21002), .B(n21003), .Z(n21004) );
  XOR U21362 ( .A(n21004), .B(n21005), .Z(n20750) );
  NANDN U21363 ( .A(n20579), .B(n20578), .Z(n20583) );
  NANDN U21364 ( .A(n20581), .B(n20580), .Z(n20582) );
  NAND U21365 ( .A(n20583), .B(n20582), .Z(n20993) );
  NANDN U21366 ( .A(n20585), .B(n20584), .Z(n20589) );
  NAND U21367 ( .A(n20587), .B(n20586), .Z(n20588) );
  AND U21368 ( .A(n20589), .B(n20588), .Z(n20990) );
  NANDN U21369 ( .A(n20591), .B(n20590), .Z(n20595) );
  NAND U21370 ( .A(n20593), .B(n20592), .Z(n20594) );
  NAND U21371 ( .A(n20595), .B(n20594), .Z(n20991) );
  XNOR U21372 ( .A(n20993), .B(n20992), .Z(n20979) );
  NANDN U21373 ( .A(n20597), .B(n20596), .Z(n20601) );
  NANDN U21374 ( .A(n20599), .B(n20598), .Z(n20600) );
  AND U21375 ( .A(n20601), .B(n20600), .Z(n20978) );
  XNOR U21376 ( .A(n20979), .B(n20978), .Z(n20980) );
  NANDN U21377 ( .A(n20603), .B(n20602), .Z(n20607) );
  NAND U21378 ( .A(n20605), .B(n20604), .Z(n20606) );
  NAND U21379 ( .A(n20607), .B(n20606), .Z(n20781) );
  XNOR U21380 ( .A(b[37]), .B(a[64]), .Z(n20810) );
  NANDN U21381 ( .A(n20810), .B(n36311), .Z(n20610) );
  NANDN U21382 ( .A(n20608), .B(n36309), .Z(n20609) );
  NAND U21383 ( .A(n20610), .B(n20609), .Z(n20843) );
  XOR U21384 ( .A(a[96]), .B(n968), .Z(n20813) );
  OR U21385 ( .A(n20813), .B(n29363), .Z(n20613) );
  NANDN U21386 ( .A(n20611), .B(n29864), .Z(n20612) );
  NAND U21387 ( .A(n20613), .B(n20612), .Z(n20840) );
  XOR U21388 ( .A(n35783), .B(n967), .Z(n20816) );
  NAND U21389 ( .A(n20816), .B(n28939), .Z(n20616) );
  NAND U21390 ( .A(n28938), .B(n20614), .Z(n20615) );
  AND U21391 ( .A(n20616), .B(n20615), .Z(n20841) );
  XNOR U21392 ( .A(n20840), .B(n20841), .Z(n20842) );
  XNOR U21393 ( .A(n20843), .B(n20842), .Z(n20776) );
  XOR U21394 ( .A(a[88]), .B(n971), .Z(n20819) );
  OR U21395 ( .A(n20819), .B(n31550), .Z(n20619) );
  NANDN U21396 ( .A(n20617), .B(n31874), .Z(n20618) );
  NAND U21397 ( .A(n20619), .B(n20618), .Z(n20953) );
  NAND U21398 ( .A(n34848), .B(n20620), .Z(n20622) );
  XOR U21399 ( .A(n35375), .B(n31372), .Z(n20822) );
  NAND U21400 ( .A(n34618), .B(n20822), .Z(n20621) );
  NAND U21401 ( .A(n20622), .B(n20621), .Z(n20950) );
  NAND U21402 ( .A(n35188), .B(n20623), .Z(n20625) );
  XOR U21403 ( .A(n35540), .B(n30210), .Z(n20825) );
  NANDN U21404 ( .A(n34968), .B(n20825), .Z(n20624) );
  AND U21405 ( .A(n20625), .B(n20624), .Z(n20951) );
  XNOR U21406 ( .A(n20950), .B(n20951), .Z(n20952) );
  XNOR U21407 ( .A(n20953), .B(n20952), .Z(n20773) );
  NANDN U21408 ( .A(n20627), .B(n20626), .Z(n20631) );
  NAND U21409 ( .A(n20629), .B(n20628), .Z(n20630) );
  NAND U21410 ( .A(n20631), .B(n20630), .Z(n20774) );
  XNOR U21411 ( .A(n20773), .B(n20774), .Z(n20775) );
  XOR U21412 ( .A(n20776), .B(n20775), .Z(n20780) );
  NANDN U21413 ( .A(n20633), .B(n20632), .Z(n20637) );
  NAND U21414 ( .A(n20635), .B(n20634), .Z(n20636) );
  NAND U21415 ( .A(n20637), .B(n20636), .Z(n20909) );
  NAND U21416 ( .A(a[36]), .B(b[63]), .Z(n20923) );
  NANDN U21417 ( .A(n20638), .B(n38369), .Z(n20640) );
  XOR U21418 ( .A(b[61]), .B(n21149), .Z(n20804) );
  OR U21419 ( .A(n20804), .B(n38371), .Z(n20639) );
  NAND U21420 ( .A(n20640), .B(n20639), .Z(n20921) );
  NANDN U21421 ( .A(n20641), .B(n35311), .Z(n20643) );
  XOR U21422 ( .A(b[31]), .B(n30379), .Z(n20807) );
  NANDN U21423 ( .A(n20807), .B(n35313), .Z(n20642) );
  AND U21424 ( .A(n20643), .B(n20642), .Z(n20920) );
  XNOR U21425 ( .A(n20921), .B(n20920), .Z(n20922) );
  XOR U21426 ( .A(n20923), .B(n20922), .Z(n20907) );
  NAND U21427 ( .A(n33283), .B(n20644), .Z(n20646) );
  XOR U21428 ( .A(n33020), .B(n32815), .Z(n20789) );
  NANDN U21429 ( .A(n33021), .B(n20789), .Z(n20645) );
  NAND U21430 ( .A(n20646), .B(n20645), .Z(n20849) );
  XNOR U21431 ( .A(b[21]), .B(a[80]), .Z(n20792) );
  OR U21432 ( .A(n20792), .B(n33634), .Z(n20649) );
  NAND U21433 ( .A(n20647), .B(n33464), .Z(n20648) );
  NAND U21434 ( .A(n20649), .B(n20648), .Z(n20846) );
  NAND U21435 ( .A(n34044), .B(n20650), .Z(n20652) );
  XOR U21436 ( .A(n34510), .B(n31870), .Z(n20795) );
  NANDN U21437 ( .A(n33867), .B(n20795), .Z(n20651) );
  AND U21438 ( .A(n20652), .B(n20651), .Z(n20847) );
  XNOR U21439 ( .A(n20846), .B(n20847), .Z(n20848) );
  XNOR U21440 ( .A(n20849), .B(n20848), .Z(n20908) );
  XNOR U21441 ( .A(n20907), .B(n20908), .Z(n20910) );
  XNOR U21442 ( .A(n20909), .B(n20910), .Z(n20779) );
  XOR U21443 ( .A(n20780), .B(n20779), .Z(n20782) );
  XNOR U21444 ( .A(n20781), .B(n20782), .Z(n20879) );
  NANDN U21445 ( .A(n20654), .B(n20653), .Z(n20658) );
  NAND U21446 ( .A(n20656), .B(n20655), .Z(n20657) );
  NAND U21447 ( .A(n20658), .B(n20657), .Z(n20878) );
  NANDN U21448 ( .A(n20660), .B(n20659), .Z(n20664) );
  NAND U21449 ( .A(n20662), .B(n20661), .Z(n20663) );
  NAND U21450 ( .A(n20664), .B(n20663), .Z(n20770) );
  NANDN U21451 ( .A(n20666), .B(n20665), .Z(n20670) );
  NAND U21452 ( .A(n20668), .B(n20667), .Z(n20669) );
  NAND U21453 ( .A(n20670), .B(n20669), .Z(n20969) );
  XNOR U21454 ( .A(b[41]), .B(a[60]), .Z(n20852) );
  OR U21455 ( .A(n20852), .B(n36905), .Z(n20673) );
  NAND U21456 ( .A(n20671), .B(n36807), .Z(n20672) );
  NAND U21457 ( .A(n20673), .B(n20672), .Z(n20874) );
  XOR U21458 ( .A(b[57]), .B(n22289), .Z(n20855) );
  OR U21459 ( .A(n20855), .B(n965), .Z(n20676) );
  NANDN U21460 ( .A(n20674), .B(n38194), .Z(n20675) );
  NAND U21461 ( .A(n20676), .B(n20675), .Z(n20871) );
  NAND U21462 ( .A(n38326), .B(n20677), .Z(n20679) );
  XOR U21463 ( .A(n38400), .B(n22246), .Z(n20858) );
  NANDN U21464 ( .A(n38273), .B(n20858), .Z(n20678) );
  AND U21465 ( .A(n20679), .B(n20678), .Z(n20872) );
  XNOR U21466 ( .A(n20871), .B(n20872), .Z(n20873) );
  XOR U21467 ( .A(n20874), .B(n20873), .Z(n20967) );
  XOR U21468 ( .A(b[33]), .B(n29868), .Z(n20861) );
  NANDN U21469 ( .A(n20861), .B(n35620), .Z(n20682) );
  NANDN U21470 ( .A(n20680), .B(n35621), .Z(n20681) );
  NAND U21471 ( .A(n20682), .B(n20681), .Z(n20965) );
  NANDN U21472 ( .A(n966), .B(a[100]), .Z(n20683) );
  XOR U21473 ( .A(n29232), .B(n20683), .Z(n20685) );
  NANDN U21474 ( .A(b[0]), .B(a[99]), .Z(n20684) );
  AND U21475 ( .A(n20685), .B(n20684), .Z(n20962) );
  XOR U21476 ( .A(b[63]), .B(n20686), .Z(n20868) );
  NANDN U21477 ( .A(n20868), .B(n38422), .Z(n20689) );
  NANDN U21478 ( .A(n20687), .B(n38423), .Z(n20688) );
  AND U21479 ( .A(n20689), .B(n20688), .Z(n20963) );
  XNOR U21480 ( .A(n20962), .B(n20963), .Z(n20964) );
  XNOR U21481 ( .A(n20965), .B(n20964), .Z(n20966) );
  XNOR U21482 ( .A(n20967), .B(n20966), .Z(n20968) );
  XOR U21483 ( .A(n20969), .B(n20968), .Z(n20768) );
  NANDN U21484 ( .A(n20691), .B(n20690), .Z(n20695) );
  NAND U21485 ( .A(n20693), .B(n20692), .Z(n20694) );
  AND U21486 ( .A(n20695), .B(n20694), .Z(n20767) );
  XNOR U21487 ( .A(n20768), .B(n20767), .Z(n20769) );
  XNOR U21488 ( .A(n20770), .B(n20769), .Z(n20877) );
  XNOR U21489 ( .A(n20878), .B(n20877), .Z(n20880) );
  XNOR U21490 ( .A(n20879), .B(n20880), .Z(n20981) );
  XOR U21491 ( .A(n20980), .B(n20981), .Z(n20749) );
  XNOR U21492 ( .A(n20750), .B(n20749), .Z(n20752) );
  XNOR U21493 ( .A(n20751), .B(n20752), .Z(n21010) );
  NANDN U21494 ( .A(n20697), .B(n20696), .Z(n20701) );
  NAND U21495 ( .A(n20699), .B(n20698), .Z(n20700) );
  NAND U21496 ( .A(n20701), .B(n20700), .Z(n20758) );
  NANDN U21497 ( .A(n20703), .B(n20702), .Z(n20707) );
  NANDN U21498 ( .A(n20705), .B(n20704), .Z(n20706) );
  NAND U21499 ( .A(n20707), .B(n20706), .Z(n20756) );
  OR U21500 ( .A(n20709), .B(n20708), .Z(n20713) );
  NANDN U21501 ( .A(n20711), .B(n20710), .Z(n20712) );
  AND U21502 ( .A(n20713), .B(n20712), .Z(n20755) );
  XNOR U21503 ( .A(n20756), .B(n20755), .Z(n20757) );
  XOR U21504 ( .A(n20758), .B(n20757), .Z(n21008) );
  NANDN U21505 ( .A(n20715), .B(n20714), .Z(n20719) );
  NANDN U21506 ( .A(n20717), .B(n20716), .Z(n20718) );
  NAND U21507 ( .A(n20719), .B(n20718), .Z(n21009) );
  XNOR U21508 ( .A(n21008), .B(n21009), .Z(n21011) );
  XOR U21509 ( .A(n21010), .B(n21011), .Z(n21017) );
  XNOR U21510 ( .A(n21016), .B(n21017), .Z(n21020) );
  OR U21511 ( .A(n20721), .B(n20720), .Z(n20725) );
  NAND U21512 ( .A(n20723), .B(n20722), .Z(n20724) );
  AND U21513 ( .A(n20725), .B(n20724), .Z(n21021) );
  XNOR U21514 ( .A(n21020), .B(n21021), .Z(n21022) );
  NANDN U21515 ( .A(n20727), .B(n20726), .Z(n20731) );
  NANDN U21516 ( .A(n20729), .B(n20728), .Z(n20730) );
  NAND U21517 ( .A(n20731), .B(n20730), .Z(n21023) );
  XOR U21518 ( .A(n21022), .B(n21023), .Z(n20743) );
  OR U21519 ( .A(n20733), .B(n20732), .Z(n20737) );
  NANDN U21520 ( .A(n20735), .B(n20734), .Z(n20736) );
  NAND U21521 ( .A(n20737), .B(n20736), .Z(n20744) );
  XNOR U21522 ( .A(n20743), .B(n20744), .Z(n20745) );
  XNOR U21523 ( .A(n20746), .B(n20745), .Z(n21024) );
  XNOR U21524 ( .A(n21024), .B(sreg[164]), .Z(n21026) );
  NAND U21525 ( .A(n20738), .B(sreg[163]), .Z(n20742) );
  OR U21526 ( .A(n20740), .B(n20739), .Z(n20741) );
  AND U21527 ( .A(n20742), .B(n20741), .Z(n21025) );
  XOR U21528 ( .A(n21026), .B(n21025), .Z(c[164]) );
  NANDN U21529 ( .A(n20744), .B(n20743), .Z(n20748) );
  NAND U21530 ( .A(n20746), .B(n20745), .Z(n20747) );
  NAND U21531 ( .A(n20748), .B(n20747), .Z(n21032) );
  NAND U21532 ( .A(n20750), .B(n20749), .Z(n20754) );
  NANDN U21533 ( .A(n20752), .B(n20751), .Z(n20753) );
  NAND U21534 ( .A(n20754), .B(n20753), .Z(n21300) );
  NANDN U21535 ( .A(n20756), .B(n20755), .Z(n20760) );
  NANDN U21536 ( .A(n20758), .B(n20757), .Z(n20759) );
  NAND U21537 ( .A(n20760), .B(n20759), .Z(n21301) );
  XNOR U21538 ( .A(n21300), .B(n21301), .Z(n21302) );
  NANDN U21539 ( .A(n20762), .B(n20761), .Z(n20766) );
  NAND U21540 ( .A(n20764), .B(n20763), .Z(n20765) );
  AND U21541 ( .A(n20766), .B(n20765), .Z(n21293) );
  NANDN U21542 ( .A(n20768), .B(n20767), .Z(n20772) );
  NANDN U21543 ( .A(n20770), .B(n20769), .Z(n20771) );
  NAND U21544 ( .A(n20772), .B(n20771), .Z(n21290) );
  NANDN U21545 ( .A(n20774), .B(n20773), .Z(n20778) );
  NAND U21546 ( .A(n20776), .B(n20775), .Z(n20777) );
  AND U21547 ( .A(n20778), .B(n20777), .Z(n21291) );
  XNOR U21548 ( .A(n21290), .B(n21291), .Z(n21292) );
  XNOR U21549 ( .A(n21293), .B(n21292), .Z(n21266) );
  NANDN U21550 ( .A(n20780), .B(n20779), .Z(n20784) );
  OR U21551 ( .A(n20782), .B(n20781), .Z(n20783) );
  AND U21552 ( .A(n20784), .B(n20783), .Z(n21267) );
  XNOR U21553 ( .A(n21266), .B(n21267), .Z(n21269) );
  NAND U21554 ( .A(n33283), .B(n20789), .Z(n20791) );
  XNOR U21555 ( .A(n33020), .B(a[83]), .Z(n21071) );
  NANDN U21556 ( .A(n33021), .B(n21071), .Z(n20790) );
  NAND U21557 ( .A(n20791), .B(n20790), .Z(n21156) );
  XOR U21558 ( .A(b[21]), .B(a[81]), .Z(n21074) );
  NANDN U21559 ( .A(n33634), .B(n21074), .Z(n20794) );
  NANDN U21560 ( .A(n20792), .B(n33464), .Z(n20793) );
  NAND U21561 ( .A(n20794), .B(n20793), .Z(n21153) );
  NAND U21562 ( .A(n34044), .B(n20795), .Z(n20797) );
  XNOR U21563 ( .A(n34510), .B(a[79]), .Z(n21077) );
  NANDN U21564 ( .A(n33867), .B(n21077), .Z(n20796) );
  AND U21565 ( .A(n20797), .B(n20796), .Z(n21154) );
  XNOR U21566 ( .A(n21153), .B(n21154), .Z(n21155) );
  XOR U21567 ( .A(n21156), .B(n21155), .Z(n21217) );
  NANDN U21568 ( .A(n20799), .B(n20798), .Z(n20803) );
  NAND U21569 ( .A(n20801), .B(n20800), .Z(n20802) );
  NAND U21570 ( .A(n20803), .B(n20802), .Z(n21218) );
  XNOR U21571 ( .A(n21217), .B(n21218), .Z(n21220) );
  NAND U21572 ( .A(a[37]), .B(b[63]), .Z(n21259) );
  NANDN U21573 ( .A(n20804), .B(n38369), .Z(n20806) );
  XOR U21574 ( .A(b[61]), .B(n21441), .Z(n21086) );
  OR U21575 ( .A(n21086), .B(n38371), .Z(n20805) );
  NAND U21576 ( .A(n20806), .B(n20805), .Z(n21257) );
  NANDN U21577 ( .A(n20807), .B(n35311), .Z(n20809) );
  XOR U21578 ( .A(b[31]), .B(n30543), .Z(n21089) );
  NANDN U21579 ( .A(n21089), .B(n35313), .Z(n20808) );
  AND U21580 ( .A(n20809), .B(n20808), .Z(n21256) );
  XNOR U21581 ( .A(n21257), .B(n21256), .Z(n21258) );
  XNOR U21582 ( .A(n21259), .B(n21258), .Z(n21219) );
  XNOR U21583 ( .A(n21220), .B(n21219), .Z(n21065) );
  XOR U21584 ( .A(b[37]), .B(n28403), .Z(n21092) );
  NANDN U21585 ( .A(n21092), .B(n36311), .Z(n20812) );
  NANDN U21586 ( .A(n20810), .B(n36309), .Z(n20811) );
  NAND U21587 ( .A(n20812), .B(n20811), .Z(n21131) );
  XNOR U21588 ( .A(a[97]), .B(b[5]), .Z(n21095) );
  OR U21589 ( .A(n21095), .B(n29363), .Z(n20815) );
  NANDN U21590 ( .A(n20813), .B(n29864), .Z(n20814) );
  NAND U21591 ( .A(n20815), .B(n20814), .Z(n21128) );
  XNOR U21592 ( .A(a[99]), .B(n967), .Z(n21098) );
  NAND U21593 ( .A(n21098), .B(n28939), .Z(n20818) );
  NAND U21594 ( .A(n28938), .B(n20816), .Z(n20817) );
  AND U21595 ( .A(n20818), .B(n20817), .Z(n21129) );
  XNOR U21596 ( .A(n21128), .B(n21129), .Z(n21130) );
  XNOR U21597 ( .A(n21131), .B(n21130), .Z(n21062) );
  XNOR U21598 ( .A(a[89]), .B(b[13]), .Z(n21101) );
  OR U21599 ( .A(n21101), .B(n31550), .Z(n20821) );
  NANDN U21600 ( .A(n20819), .B(n31874), .Z(n20820) );
  NAND U21601 ( .A(n20821), .B(n20820), .Z(n21204) );
  NAND U21602 ( .A(n34848), .B(n20822), .Z(n20824) );
  XNOR U21603 ( .A(n35375), .B(a[75]), .Z(n21104) );
  NAND U21604 ( .A(n34618), .B(n21104), .Z(n20823) );
  NAND U21605 ( .A(n20824), .B(n20823), .Z(n21201) );
  NAND U21606 ( .A(n35188), .B(n20825), .Z(n20827) );
  XNOR U21607 ( .A(n35540), .B(a[73]), .Z(n21107) );
  NANDN U21608 ( .A(n34968), .B(n21107), .Z(n20826) );
  AND U21609 ( .A(n20827), .B(n20826), .Z(n21202) );
  XNOR U21610 ( .A(n21201), .B(n21202), .Z(n21203) );
  XNOR U21611 ( .A(n21204), .B(n21203), .Z(n21059) );
  NANDN U21612 ( .A(n20829), .B(n20828), .Z(n20833) );
  NAND U21613 ( .A(n20831), .B(n20830), .Z(n20832) );
  NAND U21614 ( .A(n20833), .B(n20832), .Z(n21060) );
  XNOR U21615 ( .A(n21059), .B(n21060), .Z(n21061) );
  XOR U21616 ( .A(n21062), .B(n21061), .Z(n21066) );
  XOR U21617 ( .A(n21065), .B(n21066), .Z(n21068) );
  XNOR U21618 ( .A(n21067), .B(n21068), .Z(n21167) );
  NANDN U21619 ( .A(n20835), .B(n20834), .Z(n20839) );
  NANDN U21620 ( .A(n20837), .B(n20836), .Z(n20838) );
  NAND U21621 ( .A(n20839), .B(n20838), .Z(n21166) );
  NANDN U21622 ( .A(n20841), .B(n20840), .Z(n20845) );
  NAND U21623 ( .A(n20843), .B(n20842), .Z(n20844) );
  NAND U21624 ( .A(n20845), .B(n20844), .Z(n21056) );
  NANDN U21625 ( .A(n20847), .B(n20846), .Z(n20851) );
  NAND U21626 ( .A(n20849), .B(n20848), .Z(n20850) );
  NAND U21627 ( .A(n20851), .B(n20850), .Z(n21180) );
  XNOR U21628 ( .A(b[41]), .B(a[61]), .Z(n21134) );
  OR U21629 ( .A(n21134), .B(n36905), .Z(n20854) );
  NANDN U21630 ( .A(n20852), .B(n36807), .Z(n20853) );
  NAND U21631 ( .A(n20854), .B(n20853), .Z(n21162) );
  XOR U21632 ( .A(b[57]), .B(n22579), .Z(n21137) );
  OR U21633 ( .A(n21137), .B(n965), .Z(n20857) );
  NANDN U21634 ( .A(n20855), .B(n38194), .Z(n20856) );
  NAND U21635 ( .A(n20857), .B(n20856), .Z(n21159) );
  NAND U21636 ( .A(n38326), .B(n20858), .Z(n20860) );
  XOR U21637 ( .A(n38400), .B(n21996), .Z(n21140) );
  NANDN U21638 ( .A(n38273), .B(n21140), .Z(n20859) );
  AND U21639 ( .A(n20860), .B(n20859), .Z(n21160) );
  XNOR U21640 ( .A(n21159), .B(n21160), .Z(n21161) );
  XOR U21641 ( .A(n21162), .B(n21161), .Z(n21178) );
  XNOR U21642 ( .A(b[33]), .B(a[69]), .Z(n21143) );
  NANDN U21643 ( .A(n21143), .B(n35620), .Z(n20863) );
  NANDN U21644 ( .A(n20861), .B(n35621), .Z(n20862) );
  NAND U21645 ( .A(n20863), .B(n20862), .Z(n21216) );
  NANDN U21646 ( .A(n966), .B(a[101]), .Z(n20864) );
  XOR U21647 ( .A(n29232), .B(n20864), .Z(n20866) );
  IV U21648 ( .A(a[100]), .Z(n36100) );
  NANDN U21649 ( .A(n36100), .B(n966), .Z(n20865) );
  AND U21650 ( .A(n20866), .B(n20865), .Z(n21213) );
  XOR U21651 ( .A(b[63]), .B(n20867), .Z(n21150) );
  NANDN U21652 ( .A(n21150), .B(n38422), .Z(n20870) );
  NANDN U21653 ( .A(n20868), .B(n38423), .Z(n20869) );
  AND U21654 ( .A(n20870), .B(n20869), .Z(n21214) );
  XNOR U21655 ( .A(n21213), .B(n21214), .Z(n21215) );
  XNOR U21656 ( .A(n21216), .B(n21215), .Z(n21177) );
  XOR U21657 ( .A(n21178), .B(n21177), .Z(n21179) );
  XNOR U21658 ( .A(n21180), .B(n21179), .Z(n21054) );
  NANDN U21659 ( .A(n20872), .B(n20871), .Z(n20876) );
  NAND U21660 ( .A(n20874), .B(n20873), .Z(n20875) );
  AND U21661 ( .A(n20876), .B(n20875), .Z(n21053) );
  XNOR U21662 ( .A(n21054), .B(n21053), .Z(n21055) );
  XNOR U21663 ( .A(n21056), .B(n21055), .Z(n21165) );
  XNOR U21664 ( .A(n21166), .B(n21165), .Z(n21168) );
  XNOR U21665 ( .A(n21167), .B(n21168), .Z(n21268) );
  XOR U21666 ( .A(n21269), .B(n21268), .Z(n21041) );
  NAND U21667 ( .A(n20878), .B(n20877), .Z(n20882) );
  NANDN U21668 ( .A(n20880), .B(n20879), .Z(n20881) );
  NAND U21669 ( .A(n20882), .B(n20881), .Z(n21275) );
  NAND U21670 ( .A(n37652), .B(n20883), .Z(n20885) );
  XOR U21671 ( .A(b[49]), .B(n25001), .Z(n21232) );
  OR U21672 ( .A(n21232), .B(n37756), .Z(n20884) );
  NAND U21673 ( .A(n20885), .B(n20884), .Z(n21264) );
  NANDN U21674 ( .A(n20886), .B(n37469), .Z(n20888) );
  XNOR U21675 ( .A(n978), .B(a[55]), .Z(n21235) );
  NAND U21676 ( .A(n21235), .B(n37471), .Z(n20887) );
  NAND U21677 ( .A(n20888), .B(n20887), .Z(n21262) );
  NAND U21678 ( .A(n30846), .B(n20889), .Z(n20891) );
  XNOR U21679 ( .A(n35377), .B(b[9]), .Z(n21238) );
  NAND U21680 ( .A(n30509), .B(n21238), .Z(n20890) );
  NAND U21681 ( .A(n20891), .B(n20890), .Z(n21263) );
  XNOR U21682 ( .A(n21262), .B(n21263), .Z(n21265) );
  XOR U21683 ( .A(n21264), .B(n21265), .Z(n21116) );
  XNOR U21684 ( .A(a[91]), .B(b[11]), .Z(n21223) );
  OR U21685 ( .A(n21223), .B(n31369), .Z(n20894) );
  NANDN U21686 ( .A(n20892), .B(n31119), .Z(n20893) );
  NAND U21687 ( .A(n20894), .B(n20893), .Z(n21244) );
  XNOR U21688 ( .A(b[43]), .B(a[59]), .Z(n21226) );
  NANDN U21689 ( .A(n21226), .B(n37068), .Z(n20897) );
  NANDN U21690 ( .A(n20895), .B(n37069), .Z(n20896) );
  NAND U21691 ( .A(n20897), .B(n20896), .Z(n21241) );
  XNOR U21692 ( .A(b[45]), .B(a[57]), .Z(n21229) );
  NANDN U21693 ( .A(n21229), .B(n37261), .Z(n20900) );
  NANDN U21694 ( .A(n20898), .B(n37262), .Z(n20899) );
  AND U21695 ( .A(n20900), .B(n20899), .Z(n21242) );
  XNOR U21696 ( .A(n21241), .B(n21242), .Z(n21243) );
  XOR U21697 ( .A(n21244), .B(n21243), .Z(n21117) );
  XNOR U21698 ( .A(n21116), .B(n21117), .Z(n21118) );
  NANDN U21699 ( .A(n20902), .B(n20901), .Z(n20906) );
  NAND U21700 ( .A(n20904), .B(n20903), .Z(n20905) );
  AND U21701 ( .A(n20906), .B(n20905), .Z(n21119) );
  XNOR U21702 ( .A(n21118), .B(n21119), .Z(n21279) );
  XNOR U21703 ( .A(n21279), .B(n21278), .Z(n21280) );
  XNOR U21704 ( .A(b[35]), .B(a[67]), .Z(n21247) );
  NANDN U21705 ( .A(n21247), .B(n35985), .Z(n20913) );
  NANDN U21706 ( .A(n20911), .B(n35986), .Z(n20912) );
  NAND U21707 ( .A(n20913), .B(n20912), .Z(n21210) );
  XOR U21708 ( .A(n35628), .B(n31123), .Z(n21250) );
  NAND U21709 ( .A(n21250), .B(n29949), .Z(n20916) );
  NAND U21710 ( .A(n29948), .B(n20914), .Z(n20915) );
  NAND U21711 ( .A(n20916), .B(n20915), .Z(n21207) );
  XOR U21712 ( .A(b[55]), .B(n23149), .Z(n21253) );
  NANDN U21713 ( .A(n21253), .B(n38075), .Z(n20919) );
  NANDN U21714 ( .A(n20917), .B(n38073), .Z(n20918) );
  AND U21715 ( .A(n20919), .B(n20918), .Z(n21208) );
  XNOR U21716 ( .A(n21207), .B(n21208), .Z(n21209) );
  XNOR U21717 ( .A(n21210), .B(n21209), .Z(n21050) );
  NANDN U21718 ( .A(n20921), .B(n20920), .Z(n20925) );
  NAND U21719 ( .A(n20923), .B(n20922), .Z(n20924) );
  NAND U21720 ( .A(n20925), .B(n20924), .Z(n21047) );
  NANDN U21721 ( .A(n20927), .B(n20926), .Z(n20931) );
  NAND U21722 ( .A(n20929), .B(n20928), .Z(n20930) );
  NAND U21723 ( .A(n20931), .B(n20930), .Z(n21048) );
  XNOR U21724 ( .A(n21047), .B(n21048), .Z(n21049) );
  XOR U21725 ( .A(n21050), .B(n21049), .Z(n21281) );
  XNOR U21726 ( .A(n21280), .B(n21281), .Z(n21273) );
  XNOR U21727 ( .A(a[87]), .B(b[15]), .Z(n21183) );
  OR U21728 ( .A(n21183), .B(n32010), .Z(n20934) );
  NANDN U21729 ( .A(n20932), .B(n32011), .Z(n20933) );
  NAND U21730 ( .A(n20934), .B(n20933), .Z(n21083) );
  XOR U21731 ( .A(b[25]), .B(a[77]), .Z(n21186) );
  NANDN U21732 ( .A(n34219), .B(n21186), .Z(n20937) );
  NAND U21733 ( .A(n34217), .B(n20935), .Z(n20936) );
  NAND U21734 ( .A(n20937), .B(n20936), .Z(n21080) );
  XOR U21735 ( .A(a[85]), .B(b[17]), .Z(n21189) );
  NAND U21736 ( .A(n21189), .B(n32543), .Z(n20940) );
  NANDN U21737 ( .A(n20938), .B(n32541), .Z(n20939) );
  AND U21738 ( .A(n20940), .B(n20939), .Z(n21081) );
  XNOR U21739 ( .A(n21080), .B(n21081), .Z(n21082) );
  XNOR U21740 ( .A(n21083), .B(n21082), .Z(n21122) );
  XNOR U21741 ( .A(b[39]), .B(a[63]), .Z(n21192) );
  NANDN U21742 ( .A(n21192), .B(n36553), .Z(n20943) );
  NANDN U21743 ( .A(n20941), .B(n36643), .Z(n20942) );
  NAND U21744 ( .A(n20943), .B(n20942), .Z(n21113) );
  XOR U21745 ( .A(b[51]), .B(n24288), .Z(n21195) );
  NANDN U21746 ( .A(n21195), .B(n37803), .Z(n20946) );
  NANDN U21747 ( .A(n20944), .B(n37802), .Z(n20945) );
  NAND U21748 ( .A(n20946), .B(n20945), .Z(n21110) );
  XOR U21749 ( .A(b[53]), .B(n23852), .Z(n21198) );
  NANDN U21750 ( .A(n21198), .B(n37940), .Z(n20949) );
  NANDN U21751 ( .A(n20947), .B(n37941), .Z(n20948) );
  AND U21752 ( .A(n20949), .B(n20948), .Z(n21111) );
  XNOR U21753 ( .A(n21110), .B(n21111), .Z(n21112) );
  XOR U21754 ( .A(n21113), .B(n21112), .Z(n21123) );
  XNOR U21755 ( .A(n21122), .B(n21123), .Z(n21124) );
  NANDN U21756 ( .A(n20951), .B(n20950), .Z(n20955) );
  NAND U21757 ( .A(n20953), .B(n20952), .Z(n20954) );
  NAND U21758 ( .A(n20955), .B(n20954), .Z(n21125) );
  XOR U21759 ( .A(n21124), .B(n21125), .Z(n21174) );
  NANDN U21760 ( .A(n20957), .B(n20956), .Z(n20961) );
  NAND U21761 ( .A(n20959), .B(n20958), .Z(n20960) );
  NAND U21762 ( .A(n20961), .B(n20960), .Z(n21171) );
  XNOR U21763 ( .A(n21171), .B(n21172), .Z(n21173) );
  XNOR U21764 ( .A(n21174), .B(n21173), .Z(n21284) );
  NANDN U21765 ( .A(n20967), .B(n20966), .Z(n20971) );
  NANDN U21766 ( .A(n20969), .B(n20968), .Z(n20970) );
  AND U21767 ( .A(n20971), .B(n20970), .Z(n21285) );
  XOR U21768 ( .A(n21284), .B(n21285), .Z(n21287) );
  NANDN U21769 ( .A(n20973), .B(n20972), .Z(n20977) );
  NANDN U21770 ( .A(n20975), .B(n20974), .Z(n20976) );
  AND U21771 ( .A(n20977), .B(n20976), .Z(n21286) );
  XNOR U21772 ( .A(n21287), .B(n21286), .Z(n21272) );
  XOR U21773 ( .A(n21275), .B(n21274), .Z(n21042) );
  XNOR U21774 ( .A(n21041), .B(n21042), .Z(n21043) );
  NANDN U21775 ( .A(n20979), .B(n20978), .Z(n20983) );
  NAND U21776 ( .A(n20981), .B(n20980), .Z(n20982) );
  NAND U21777 ( .A(n20983), .B(n20982), .Z(n21044) );
  XOR U21778 ( .A(n21043), .B(n21044), .Z(n21297) );
  OR U21779 ( .A(n20985), .B(n20984), .Z(n20989) );
  NAND U21780 ( .A(n20987), .B(n20986), .Z(n20988) );
  NAND U21781 ( .A(n20989), .B(n20988), .Z(n21036) );
  OR U21782 ( .A(n20991), .B(n20990), .Z(n20995) );
  NAND U21783 ( .A(n20993), .B(n20992), .Z(n20994) );
  AND U21784 ( .A(n20995), .B(n20994), .Z(n21035) );
  XNOR U21785 ( .A(n21036), .B(n21035), .Z(n21037) );
  NAND U21786 ( .A(n20997), .B(n20996), .Z(n21001) );
  NANDN U21787 ( .A(n20999), .B(n20998), .Z(n21000) );
  NAND U21788 ( .A(n21001), .B(n21000), .Z(n21038) );
  XOR U21789 ( .A(n21037), .B(n21038), .Z(n21294) );
  NANDN U21790 ( .A(n21003), .B(n21002), .Z(n21007) );
  NANDN U21791 ( .A(n21005), .B(n21004), .Z(n21006) );
  NAND U21792 ( .A(n21007), .B(n21006), .Z(n21295) );
  XNOR U21793 ( .A(n21294), .B(n21295), .Z(n21296) );
  XNOR U21794 ( .A(n21297), .B(n21296), .Z(n21303) );
  XOR U21795 ( .A(n21302), .B(n21303), .Z(n21306) );
  NANDN U21796 ( .A(n21009), .B(n21008), .Z(n21013) );
  NAND U21797 ( .A(n21011), .B(n21010), .Z(n21012) );
  NAND U21798 ( .A(n21013), .B(n21012), .Z(n21307) );
  XNOR U21799 ( .A(n21306), .B(n21307), .Z(n21308) );
  NANDN U21800 ( .A(n21015), .B(n21014), .Z(n21019) );
  NAND U21801 ( .A(n21017), .B(n21016), .Z(n21018) );
  NAND U21802 ( .A(n21019), .B(n21018), .Z(n21309) );
  XOR U21803 ( .A(n21308), .B(n21309), .Z(n21029) );
  XNOR U21804 ( .A(n21029), .B(n21030), .Z(n21031) );
  XNOR U21805 ( .A(n21032), .B(n21031), .Z(n21312) );
  XNOR U21806 ( .A(n21312), .B(sreg[165]), .Z(n21314) );
  NAND U21807 ( .A(n21024), .B(sreg[164]), .Z(n21028) );
  OR U21808 ( .A(n21026), .B(n21025), .Z(n21027) );
  AND U21809 ( .A(n21028), .B(n21027), .Z(n21313) );
  XOR U21810 ( .A(n21314), .B(n21313), .Z(c[165]) );
  NANDN U21811 ( .A(n21030), .B(n21029), .Z(n21034) );
  NAND U21812 ( .A(n21032), .B(n21031), .Z(n21033) );
  NAND U21813 ( .A(n21034), .B(n21033), .Z(n21320) );
  NANDN U21814 ( .A(n21036), .B(n21035), .Z(n21040) );
  NANDN U21815 ( .A(n21038), .B(n21037), .Z(n21039) );
  NAND U21816 ( .A(n21040), .B(n21039), .Z(n21587) );
  NANDN U21817 ( .A(n21042), .B(n21041), .Z(n21046) );
  NANDN U21818 ( .A(n21044), .B(n21043), .Z(n21045) );
  AND U21819 ( .A(n21046), .B(n21045), .Z(n21586) );
  XNOR U21820 ( .A(n21587), .B(n21586), .Z(n21588) );
  NANDN U21821 ( .A(n21048), .B(n21047), .Z(n21052) );
  NAND U21822 ( .A(n21050), .B(n21049), .Z(n21051) );
  AND U21823 ( .A(n21052), .B(n21051), .Z(n21575) );
  NANDN U21824 ( .A(n21054), .B(n21053), .Z(n21058) );
  NANDN U21825 ( .A(n21056), .B(n21055), .Z(n21057) );
  NAND U21826 ( .A(n21058), .B(n21057), .Z(n21572) );
  NANDN U21827 ( .A(n21060), .B(n21059), .Z(n21064) );
  NAND U21828 ( .A(n21062), .B(n21061), .Z(n21063) );
  AND U21829 ( .A(n21064), .B(n21063), .Z(n21573) );
  XNOR U21830 ( .A(n21572), .B(n21573), .Z(n21574) );
  XNOR U21831 ( .A(n21575), .B(n21574), .Z(n21554) );
  NANDN U21832 ( .A(n21066), .B(n21065), .Z(n21070) );
  OR U21833 ( .A(n21068), .B(n21067), .Z(n21069) );
  AND U21834 ( .A(n21070), .B(n21069), .Z(n21555) );
  XNOR U21835 ( .A(n21554), .B(n21555), .Z(n21557) );
  NAND U21836 ( .A(n33283), .B(n21071), .Z(n21073) );
  XOR U21837 ( .A(n33020), .B(n33185), .Z(n21399) );
  NANDN U21838 ( .A(n33021), .B(n21399), .Z(n21072) );
  NAND U21839 ( .A(n21073), .B(n21072), .Z(n21423) );
  XNOR U21840 ( .A(b[21]), .B(a[82]), .Z(n21402) );
  OR U21841 ( .A(n21402), .B(n33634), .Z(n21076) );
  NAND U21842 ( .A(n21074), .B(n33464), .Z(n21075) );
  NAND U21843 ( .A(n21076), .B(n21075), .Z(n21420) );
  NAND U21844 ( .A(n34044), .B(n21077), .Z(n21079) );
  XOR U21845 ( .A(n34510), .B(n32814), .Z(n21405) );
  NANDN U21846 ( .A(n33867), .B(n21405), .Z(n21078) );
  AND U21847 ( .A(n21079), .B(n21078), .Z(n21421) );
  XNOR U21848 ( .A(n21420), .B(n21421), .Z(n21422) );
  XOR U21849 ( .A(n21423), .B(n21422), .Z(n21457) );
  NANDN U21850 ( .A(n21081), .B(n21080), .Z(n21085) );
  NAND U21851 ( .A(n21083), .B(n21082), .Z(n21084) );
  NAND U21852 ( .A(n21085), .B(n21084), .Z(n21458) );
  XNOR U21853 ( .A(n21457), .B(n21458), .Z(n21460) );
  NAND U21854 ( .A(a[38]), .B(b[63]), .Z(n21499) );
  NANDN U21855 ( .A(n21086), .B(n38369), .Z(n21088) );
  XOR U21856 ( .A(b[61]), .B(n22246), .Z(n21393) );
  OR U21857 ( .A(n21393), .B(n38371), .Z(n21087) );
  NAND U21858 ( .A(n21088), .B(n21087), .Z(n21497) );
  NANDN U21859 ( .A(n21089), .B(n35311), .Z(n21091) );
  XOR U21860 ( .A(b[31]), .B(n30210), .Z(n21396) );
  NANDN U21861 ( .A(n21396), .B(n35313), .Z(n21090) );
  AND U21862 ( .A(n21091), .B(n21090), .Z(n21496) );
  XNOR U21863 ( .A(n21497), .B(n21496), .Z(n21498) );
  XNOR U21864 ( .A(n21499), .B(n21498), .Z(n21459) );
  XNOR U21865 ( .A(n21460), .B(n21459), .Z(n21335) );
  XOR U21866 ( .A(b[37]), .B(n28701), .Z(n21363) );
  NANDN U21867 ( .A(n21363), .B(n36311), .Z(n21094) );
  NANDN U21868 ( .A(n21092), .B(n36309), .Z(n21093) );
  NAND U21869 ( .A(n21094), .B(n21093), .Z(n21417) );
  XOR U21870 ( .A(a[98]), .B(n968), .Z(n21366) );
  OR U21871 ( .A(n21366), .B(n29363), .Z(n21097) );
  NANDN U21872 ( .A(n21095), .B(n29864), .Z(n21096) );
  NAND U21873 ( .A(n21097), .B(n21096), .Z(n21414) );
  XOR U21874 ( .A(n36100), .B(n967), .Z(n21369) );
  NAND U21875 ( .A(n21369), .B(n28939), .Z(n21100) );
  NAND U21876 ( .A(n28938), .B(n21098), .Z(n21099) );
  AND U21877 ( .A(n21100), .B(n21099), .Z(n21415) );
  XNOR U21878 ( .A(n21414), .B(n21415), .Z(n21416) );
  XOR U21879 ( .A(n21417), .B(n21416), .Z(n21356) );
  XOR U21880 ( .A(a[90]), .B(n971), .Z(n21372) );
  OR U21881 ( .A(n21372), .B(n31550), .Z(n21103) );
  NANDN U21882 ( .A(n21101), .B(n31874), .Z(n21102) );
  NAND U21883 ( .A(n21103), .B(n21102), .Z(n21545) );
  NAND U21884 ( .A(n34848), .B(n21104), .Z(n21106) );
  XOR U21885 ( .A(n35375), .B(n31363), .Z(n21375) );
  NAND U21886 ( .A(n34618), .B(n21375), .Z(n21105) );
  NAND U21887 ( .A(n21106), .B(n21105), .Z(n21542) );
  NAND U21888 ( .A(n35188), .B(n21107), .Z(n21109) );
  XOR U21889 ( .A(n35540), .B(n31372), .Z(n21378) );
  NANDN U21890 ( .A(n34968), .B(n21378), .Z(n21108) );
  AND U21891 ( .A(n21109), .B(n21108), .Z(n21543) );
  XNOR U21892 ( .A(n21542), .B(n21543), .Z(n21544) );
  XOR U21893 ( .A(n21545), .B(n21544), .Z(n21354) );
  NANDN U21894 ( .A(n21111), .B(n21110), .Z(n21115) );
  NAND U21895 ( .A(n21113), .B(n21112), .Z(n21114) );
  AND U21896 ( .A(n21115), .B(n21114), .Z(n21353) );
  XOR U21897 ( .A(n21354), .B(n21353), .Z(n21355) );
  XOR U21898 ( .A(n21356), .B(n21355), .Z(n21336) );
  XOR U21899 ( .A(n21335), .B(n21336), .Z(n21338) );
  NANDN U21900 ( .A(n21117), .B(n21116), .Z(n21121) );
  NAND U21901 ( .A(n21119), .B(n21118), .Z(n21120) );
  NAND U21902 ( .A(n21121), .B(n21120), .Z(n21337) );
  XNOR U21903 ( .A(n21338), .B(n21337), .Z(n21453) );
  NANDN U21904 ( .A(n21123), .B(n21122), .Z(n21127) );
  NANDN U21905 ( .A(n21125), .B(n21124), .Z(n21126) );
  NAND U21906 ( .A(n21127), .B(n21126), .Z(n21452) );
  NANDN U21907 ( .A(n21129), .B(n21128), .Z(n21133) );
  NAND U21908 ( .A(n21131), .B(n21130), .Z(n21132) );
  NAND U21909 ( .A(n21133), .B(n21132), .Z(n21350) );
  XOR U21910 ( .A(b[41]), .B(a[62]), .Z(n21426) );
  NANDN U21911 ( .A(n36905), .B(n21426), .Z(n21136) );
  NANDN U21912 ( .A(n21134), .B(n36807), .Z(n21135) );
  NAND U21913 ( .A(n21136), .B(n21135), .Z(n21448) );
  XOR U21914 ( .A(b[57]), .B(n22964), .Z(n21429) );
  OR U21915 ( .A(n21429), .B(n965), .Z(n21139) );
  NANDN U21916 ( .A(n21137), .B(n38194), .Z(n21138) );
  NAND U21917 ( .A(n21139), .B(n21138), .Z(n21445) );
  NAND U21918 ( .A(n38326), .B(n21140), .Z(n21142) );
  XOR U21919 ( .A(n38400), .B(n22289), .Z(n21432) );
  NANDN U21920 ( .A(n38273), .B(n21432), .Z(n21141) );
  AND U21921 ( .A(n21142), .B(n21141), .Z(n21446) );
  XNOR U21922 ( .A(n21445), .B(n21446), .Z(n21447) );
  XOR U21923 ( .A(n21448), .B(n21447), .Z(n21508) );
  XOR U21924 ( .A(b[33]), .B(n30379), .Z(n21435) );
  NANDN U21925 ( .A(n21435), .B(n35620), .Z(n21145) );
  NANDN U21926 ( .A(n21143), .B(n35621), .Z(n21144) );
  NAND U21927 ( .A(n21145), .B(n21144), .Z(n21521) );
  NANDN U21928 ( .A(n966), .B(a[102]), .Z(n21146) );
  XOR U21929 ( .A(n29232), .B(n21146), .Z(n21148) );
  NANDN U21930 ( .A(b[0]), .B(a[101]), .Z(n21147) );
  AND U21931 ( .A(n21148), .B(n21147), .Z(n21518) );
  XOR U21932 ( .A(b[63]), .B(n21149), .Z(n21442) );
  NANDN U21933 ( .A(n21442), .B(n38422), .Z(n21152) );
  NANDN U21934 ( .A(n21150), .B(n38423), .Z(n21151) );
  AND U21935 ( .A(n21152), .B(n21151), .Z(n21519) );
  XNOR U21936 ( .A(n21518), .B(n21519), .Z(n21520) );
  XOR U21937 ( .A(n21521), .B(n21520), .Z(n21509) );
  XNOR U21938 ( .A(n21508), .B(n21509), .Z(n21511) );
  NANDN U21939 ( .A(n21154), .B(n21153), .Z(n21158) );
  NAND U21940 ( .A(n21156), .B(n21155), .Z(n21157) );
  AND U21941 ( .A(n21158), .B(n21157), .Z(n21510) );
  XNOR U21942 ( .A(n21511), .B(n21510), .Z(n21347) );
  NANDN U21943 ( .A(n21160), .B(n21159), .Z(n21164) );
  NAND U21944 ( .A(n21162), .B(n21161), .Z(n21163) );
  AND U21945 ( .A(n21164), .B(n21163), .Z(n21348) );
  XOR U21946 ( .A(n21347), .B(n21348), .Z(n21349) );
  XNOR U21947 ( .A(n21350), .B(n21349), .Z(n21451) );
  XNOR U21948 ( .A(n21452), .B(n21451), .Z(n21454) );
  XNOR U21949 ( .A(n21453), .B(n21454), .Z(n21556) );
  XOR U21950 ( .A(n21557), .B(n21556), .Z(n21329) );
  NAND U21951 ( .A(n21166), .B(n21165), .Z(n21170) );
  NANDN U21952 ( .A(n21168), .B(n21167), .Z(n21169) );
  NAND U21953 ( .A(n21170), .B(n21169), .Z(n21563) );
  NANDN U21954 ( .A(n21172), .B(n21171), .Z(n21176) );
  NAND U21955 ( .A(n21174), .B(n21173), .Z(n21175) );
  NAND U21956 ( .A(n21176), .B(n21175), .Z(n21579) );
  NANDN U21957 ( .A(n21178), .B(n21177), .Z(n21182) );
  OR U21958 ( .A(n21180), .B(n21179), .Z(n21181) );
  NAND U21959 ( .A(n21182), .B(n21181), .Z(n21577) );
  XOR U21960 ( .A(a[88]), .B(n972), .Z(n21524) );
  OR U21961 ( .A(n21524), .B(n32010), .Z(n21185) );
  NANDN U21962 ( .A(n21183), .B(n32011), .Z(n21184) );
  NAND U21963 ( .A(n21185), .B(n21184), .Z(n21390) );
  XNOR U21964 ( .A(b[25]), .B(n31870), .Z(n21527) );
  NANDN U21965 ( .A(n34219), .B(n21527), .Z(n21188) );
  NAND U21966 ( .A(n34217), .B(n21186), .Z(n21187) );
  NAND U21967 ( .A(n21188), .B(n21187), .Z(n21387) );
  XNOR U21968 ( .A(a[86]), .B(b[17]), .Z(n21530) );
  NANDN U21969 ( .A(n21530), .B(n32543), .Z(n21191) );
  NAND U21970 ( .A(n21189), .B(n32541), .Z(n21190) );
  AND U21971 ( .A(n21191), .B(n21190), .Z(n21388) );
  XNOR U21972 ( .A(n21387), .B(n21388), .Z(n21389) );
  XNOR U21973 ( .A(n21390), .B(n21389), .Z(n21408) );
  XNOR U21974 ( .A(b[39]), .B(a[64]), .Z(n21533) );
  NANDN U21975 ( .A(n21533), .B(n36553), .Z(n21194) );
  NANDN U21976 ( .A(n21192), .B(n36643), .Z(n21193) );
  NAND U21977 ( .A(n21194), .B(n21193), .Z(n21384) );
  XOR U21978 ( .A(b[51]), .B(n25134), .Z(n21536) );
  NANDN U21979 ( .A(n21536), .B(n37803), .Z(n21197) );
  NANDN U21980 ( .A(n21195), .B(n37802), .Z(n21196) );
  NAND U21981 ( .A(n21197), .B(n21196), .Z(n21381) );
  XOR U21982 ( .A(b[53]), .B(n24671), .Z(n21539) );
  NANDN U21983 ( .A(n21539), .B(n37940), .Z(n21200) );
  NANDN U21984 ( .A(n21198), .B(n37941), .Z(n21199) );
  AND U21985 ( .A(n21200), .B(n21199), .Z(n21382) );
  XNOR U21986 ( .A(n21381), .B(n21382), .Z(n21383) );
  XOR U21987 ( .A(n21384), .B(n21383), .Z(n21409) );
  XOR U21988 ( .A(n21408), .B(n21409), .Z(n21411) );
  NANDN U21989 ( .A(n21202), .B(n21201), .Z(n21206) );
  NAND U21990 ( .A(n21204), .B(n21203), .Z(n21205) );
  NAND U21991 ( .A(n21206), .B(n21205), .Z(n21410) );
  XNOR U21992 ( .A(n21411), .B(n21410), .Z(n21515) );
  NANDN U21993 ( .A(n21208), .B(n21207), .Z(n21212) );
  NAND U21994 ( .A(n21210), .B(n21209), .Z(n21211) );
  NAND U21995 ( .A(n21212), .B(n21211), .Z(n21512) );
  XNOR U21996 ( .A(n21512), .B(n21513), .Z(n21514) );
  XOR U21997 ( .A(n21515), .B(n21514), .Z(n21576) );
  XNOR U21998 ( .A(n21577), .B(n21576), .Z(n21578) );
  XNOR U21999 ( .A(n21579), .B(n21578), .Z(n21560) );
  OR U22000 ( .A(n21218), .B(n21217), .Z(n21222) );
  OR U22001 ( .A(n21220), .B(n21219), .Z(n21221) );
  NAND U22002 ( .A(n21222), .B(n21221), .Z(n21567) );
  XOR U22003 ( .A(a[92]), .B(n970), .Z(n21463) );
  OR U22004 ( .A(n21463), .B(n31369), .Z(n21225) );
  NANDN U22005 ( .A(n21223), .B(n31119), .Z(n21224) );
  NAND U22006 ( .A(n21225), .B(n21224), .Z(n21484) );
  XOR U22007 ( .A(b[43]), .B(n27436), .Z(n21466) );
  NANDN U22008 ( .A(n21466), .B(n37068), .Z(n21228) );
  NANDN U22009 ( .A(n21226), .B(n37069), .Z(n21227) );
  NAND U22010 ( .A(n21228), .B(n21227), .Z(n21481) );
  XNOR U22011 ( .A(b[45]), .B(a[58]), .Z(n21469) );
  NANDN U22012 ( .A(n21469), .B(n37261), .Z(n21231) );
  NANDN U22013 ( .A(n21229), .B(n37262), .Z(n21230) );
  AND U22014 ( .A(n21231), .B(n21230), .Z(n21482) );
  XNOR U22015 ( .A(n21481), .B(n21482), .Z(n21483) );
  XNOR U22016 ( .A(n21484), .B(n21483), .Z(n21362) );
  XOR U22017 ( .A(n979), .B(n25177), .Z(n21472) );
  NANDN U22018 ( .A(n37756), .B(n21472), .Z(n21234) );
  NANDN U22019 ( .A(n21232), .B(n37652), .Z(n21233) );
  NAND U22020 ( .A(n21234), .B(n21233), .Z(n21505) );
  NAND U22021 ( .A(n21235), .B(n37469), .Z(n21237) );
  XOR U22022 ( .A(b[47]), .B(n25860), .Z(n21475) );
  NANDN U22023 ( .A(n21475), .B(n37471), .Z(n21236) );
  NAND U22024 ( .A(n21237), .B(n21236), .Z(n21502) );
  XOR U22025 ( .A(n35191), .B(n969), .Z(n21478) );
  NAND U22026 ( .A(n30509), .B(n21478), .Z(n21240) );
  NAND U22027 ( .A(n21238), .B(n30846), .Z(n21239) );
  AND U22028 ( .A(n21240), .B(n21239), .Z(n21503) );
  XNOR U22029 ( .A(n21502), .B(n21503), .Z(n21504) );
  XNOR U22030 ( .A(n21505), .B(n21504), .Z(n21359) );
  NANDN U22031 ( .A(n21242), .B(n21241), .Z(n21246) );
  NAND U22032 ( .A(n21244), .B(n21243), .Z(n21245) );
  NAND U22033 ( .A(n21246), .B(n21245), .Z(n21360) );
  XNOR U22034 ( .A(n21359), .B(n21360), .Z(n21361) );
  XOR U22035 ( .A(n21362), .B(n21361), .Z(n21566) );
  XNOR U22036 ( .A(n21567), .B(n21566), .Z(n21569) );
  XNOR U22037 ( .A(b[35]), .B(a[68]), .Z(n21487) );
  NANDN U22038 ( .A(n21487), .B(n35985), .Z(n21249) );
  NANDN U22039 ( .A(n21247), .B(n35986), .Z(n21248) );
  NAND U22040 ( .A(n21249), .B(n21248), .Z(n21551) );
  XOR U22041 ( .A(n35545), .B(n31123), .Z(n21490) );
  NAND U22042 ( .A(n21490), .B(n29949), .Z(n21252) );
  NAND U22043 ( .A(n29948), .B(n21250), .Z(n21251) );
  NAND U22044 ( .A(n21252), .B(n21251), .Z(n21548) );
  XOR U22045 ( .A(b[55]), .B(n23447), .Z(n21493) );
  NANDN U22046 ( .A(n21493), .B(n38075), .Z(n21255) );
  NANDN U22047 ( .A(n21253), .B(n38073), .Z(n21254) );
  AND U22048 ( .A(n21255), .B(n21254), .Z(n21549) );
  XNOR U22049 ( .A(n21548), .B(n21549), .Z(n21550) );
  XNOR U22050 ( .A(n21551), .B(n21550), .Z(n21344) );
  NANDN U22051 ( .A(n21257), .B(n21256), .Z(n21261) );
  NAND U22052 ( .A(n21259), .B(n21258), .Z(n21260) );
  NAND U22053 ( .A(n21261), .B(n21260), .Z(n21341) );
  XNOR U22054 ( .A(n21341), .B(n21342), .Z(n21343) );
  XOR U22055 ( .A(n21344), .B(n21343), .Z(n21568) );
  XOR U22056 ( .A(n21569), .B(n21568), .Z(n21561) );
  XNOR U22057 ( .A(n21560), .B(n21561), .Z(n21562) );
  XOR U22058 ( .A(n21563), .B(n21562), .Z(n21330) );
  XNOR U22059 ( .A(n21329), .B(n21330), .Z(n21331) );
  NAND U22060 ( .A(n21267), .B(n21266), .Z(n21271) );
  NANDN U22061 ( .A(n21269), .B(n21268), .Z(n21270) );
  NAND U22062 ( .A(n21271), .B(n21270), .Z(n21332) );
  XOR U22063 ( .A(n21331), .B(n21332), .Z(n21583) );
  NANDN U22064 ( .A(n21273), .B(n21272), .Z(n21277) );
  NAND U22065 ( .A(n21275), .B(n21274), .Z(n21276) );
  AND U22066 ( .A(n21277), .B(n21276), .Z(n21580) );
  NANDN U22067 ( .A(n21279), .B(n21278), .Z(n21283) );
  NAND U22068 ( .A(n21281), .B(n21280), .Z(n21282) );
  NAND U22069 ( .A(n21283), .B(n21282), .Z(n21326) );
  NANDN U22070 ( .A(n21285), .B(n21284), .Z(n21289) );
  NANDN U22071 ( .A(n21287), .B(n21286), .Z(n21288) );
  NAND U22072 ( .A(n21289), .B(n21288), .Z(n21323) );
  XNOR U22073 ( .A(n21323), .B(n21324), .Z(n21325) );
  XNOR U22074 ( .A(n21326), .B(n21325), .Z(n21581) );
  XNOR U22075 ( .A(n21583), .B(n21582), .Z(n21589) );
  XOR U22076 ( .A(n21588), .B(n21589), .Z(n21592) );
  NANDN U22077 ( .A(n21295), .B(n21294), .Z(n21299) );
  NAND U22078 ( .A(n21297), .B(n21296), .Z(n21298) );
  NAND U22079 ( .A(n21299), .B(n21298), .Z(n21593) );
  XNOR U22080 ( .A(n21592), .B(n21593), .Z(n21594) );
  NANDN U22081 ( .A(n21301), .B(n21300), .Z(n21305) );
  NANDN U22082 ( .A(n21303), .B(n21302), .Z(n21304) );
  NAND U22083 ( .A(n21305), .B(n21304), .Z(n21595) );
  XOR U22084 ( .A(n21594), .B(n21595), .Z(n21317) );
  NANDN U22085 ( .A(n21307), .B(n21306), .Z(n21311) );
  NANDN U22086 ( .A(n21309), .B(n21308), .Z(n21310) );
  NAND U22087 ( .A(n21311), .B(n21310), .Z(n21318) );
  XNOR U22088 ( .A(n21317), .B(n21318), .Z(n21319) );
  XNOR U22089 ( .A(n21320), .B(n21319), .Z(n21598) );
  XNOR U22090 ( .A(n21598), .B(sreg[166]), .Z(n21600) );
  NAND U22091 ( .A(n21312), .B(sreg[165]), .Z(n21316) );
  OR U22092 ( .A(n21314), .B(n21313), .Z(n21315) );
  AND U22093 ( .A(n21316), .B(n21315), .Z(n21599) );
  XOR U22094 ( .A(n21600), .B(n21599), .Z(c[166]) );
  NANDN U22095 ( .A(n21318), .B(n21317), .Z(n21322) );
  NAND U22096 ( .A(n21320), .B(n21319), .Z(n21321) );
  NAND U22097 ( .A(n21322), .B(n21321), .Z(n21606) );
  NANDN U22098 ( .A(n21324), .B(n21323), .Z(n21328) );
  NAND U22099 ( .A(n21326), .B(n21325), .Z(n21327) );
  NAND U22100 ( .A(n21328), .B(n21327), .Z(n21867) );
  NANDN U22101 ( .A(n21330), .B(n21329), .Z(n21334) );
  NANDN U22102 ( .A(n21332), .B(n21331), .Z(n21333) );
  NAND U22103 ( .A(n21334), .B(n21333), .Z(n21868) );
  XNOR U22104 ( .A(n21867), .B(n21868), .Z(n21869) );
  NANDN U22105 ( .A(n21336), .B(n21335), .Z(n21340) );
  OR U22106 ( .A(n21338), .B(n21337), .Z(n21339) );
  NAND U22107 ( .A(n21340), .B(n21339), .Z(n21833) );
  NANDN U22108 ( .A(n21342), .B(n21341), .Z(n21346) );
  NAND U22109 ( .A(n21344), .B(n21343), .Z(n21345) );
  NAND U22110 ( .A(n21346), .B(n21345), .Z(n21859) );
  NAND U22111 ( .A(n21348), .B(n21347), .Z(n21352) );
  NANDN U22112 ( .A(n21350), .B(n21349), .Z(n21351) );
  NAND U22113 ( .A(n21352), .B(n21351), .Z(n21857) );
  NANDN U22114 ( .A(n21354), .B(n21353), .Z(n21358) );
  OR U22115 ( .A(n21356), .B(n21355), .Z(n21357) );
  AND U22116 ( .A(n21358), .B(n21357), .Z(n21858) );
  XNOR U22117 ( .A(n21857), .B(n21858), .Z(n21860) );
  XNOR U22118 ( .A(n21859), .B(n21860), .Z(n21834) );
  XOR U22119 ( .A(n21833), .B(n21834), .Z(n21835) );
  XOR U22120 ( .A(b[37]), .B(n29372), .Z(n21662) );
  NANDN U22121 ( .A(n21662), .B(n36311), .Z(n21365) );
  NANDN U22122 ( .A(n21363), .B(n36309), .Z(n21364) );
  NAND U22123 ( .A(n21365), .B(n21364), .Z(n21701) );
  XNOR U22124 ( .A(a[99]), .B(b[5]), .Z(n21665) );
  OR U22125 ( .A(n21665), .B(n29363), .Z(n21368) );
  NANDN U22126 ( .A(n21366), .B(n29864), .Z(n21367) );
  NAND U22127 ( .A(n21368), .B(n21367), .Z(n21698) );
  XNOR U22128 ( .A(a[101]), .B(n967), .Z(n21668) );
  NAND U22129 ( .A(n21668), .B(n28939), .Z(n21371) );
  NAND U22130 ( .A(n28938), .B(n21369), .Z(n21370) );
  AND U22131 ( .A(n21371), .B(n21370), .Z(n21699) );
  XNOR U22132 ( .A(n21698), .B(n21699), .Z(n21700) );
  XNOR U22133 ( .A(n21701), .B(n21700), .Z(n21632) );
  XNOR U22134 ( .A(a[91]), .B(b[13]), .Z(n21671) );
  OR U22135 ( .A(n21671), .B(n31550), .Z(n21374) );
  NANDN U22136 ( .A(n21372), .B(n31874), .Z(n21373) );
  NAND U22137 ( .A(n21374), .B(n21373), .Z(n21814) );
  NAND U22138 ( .A(n34848), .B(n21375), .Z(n21377) );
  XNOR U22139 ( .A(n35375), .B(a[77]), .Z(n21674) );
  NAND U22140 ( .A(n34618), .B(n21674), .Z(n21376) );
  NAND U22141 ( .A(n21377), .B(n21376), .Z(n21811) );
  NAND U22142 ( .A(n35188), .B(n21378), .Z(n21380) );
  XNOR U22143 ( .A(n35540), .B(a[75]), .Z(n21677) );
  NANDN U22144 ( .A(n34968), .B(n21677), .Z(n21379) );
  AND U22145 ( .A(n21380), .B(n21379), .Z(n21812) );
  XNOR U22146 ( .A(n21811), .B(n21812), .Z(n21813) );
  XNOR U22147 ( .A(n21814), .B(n21813), .Z(n21629) );
  NANDN U22148 ( .A(n21382), .B(n21381), .Z(n21386) );
  NAND U22149 ( .A(n21384), .B(n21383), .Z(n21385) );
  NAND U22150 ( .A(n21386), .B(n21385), .Z(n21630) );
  XNOR U22151 ( .A(n21629), .B(n21630), .Z(n21631) );
  XOR U22152 ( .A(n21632), .B(n21631), .Z(n21636) );
  NANDN U22153 ( .A(n21388), .B(n21387), .Z(n21392) );
  NAND U22154 ( .A(n21390), .B(n21389), .Z(n21391) );
  NAND U22155 ( .A(n21392), .B(n21391), .Z(n21766) );
  NAND U22156 ( .A(a[39]), .B(b[63]), .Z(n21780) );
  NANDN U22157 ( .A(n21393), .B(n38369), .Z(n21395) );
  XOR U22158 ( .A(b[61]), .B(n21996), .Z(n21656) );
  OR U22159 ( .A(n21656), .B(n38371), .Z(n21394) );
  NAND U22160 ( .A(n21395), .B(n21394), .Z(n21778) );
  NANDN U22161 ( .A(n21396), .B(n35311), .Z(n21398) );
  XNOR U22162 ( .A(b[31]), .B(a[73]), .Z(n21659) );
  NANDN U22163 ( .A(n21659), .B(n35313), .Z(n21397) );
  AND U22164 ( .A(n21398), .B(n21397), .Z(n21777) );
  XNOR U22165 ( .A(n21778), .B(n21777), .Z(n21779) );
  XOR U22166 ( .A(n21780), .B(n21779), .Z(n21764) );
  NAND U22167 ( .A(n33283), .B(n21399), .Z(n21401) );
  XNOR U22168 ( .A(n33020), .B(a[85]), .Z(n21641) );
  NANDN U22169 ( .A(n33021), .B(n21641), .Z(n21400) );
  NAND U22170 ( .A(n21401), .B(n21400), .Z(n21725) );
  XOR U22171 ( .A(b[21]), .B(a[83]), .Z(n21644) );
  NANDN U22172 ( .A(n33634), .B(n21644), .Z(n21404) );
  NANDN U22173 ( .A(n21402), .B(n33464), .Z(n21403) );
  NAND U22174 ( .A(n21404), .B(n21403), .Z(n21722) );
  NAND U22175 ( .A(n34044), .B(n21405), .Z(n21407) );
  XNOR U22176 ( .A(n34510), .B(a[81]), .Z(n21647) );
  NANDN U22177 ( .A(n33867), .B(n21647), .Z(n21406) );
  AND U22178 ( .A(n21407), .B(n21406), .Z(n21723) );
  XNOR U22179 ( .A(n21722), .B(n21723), .Z(n21724) );
  XNOR U22180 ( .A(n21725), .B(n21724), .Z(n21765) );
  XNOR U22181 ( .A(n21764), .B(n21765), .Z(n21767) );
  XNOR U22182 ( .A(n21766), .B(n21767), .Z(n21635) );
  XOR U22183 ( .A(n21636), .B(n21635), .Z(n21638) );
  XNOR U22184 ( .A(n21637), .B(n21638), .Z(n21736) );
  NANDN U22185 ( .A(n21409), .B(n21408), .Z(n21413) );
  OR U22186 ( .A(n21411), .B(n21410), .Z(n21412) );
  NAND U22187 ( .A(n21413), .B(n21412), .Z(n21735) );
  NANDN U22188 ( .A(n21415), .B(n21414), .Z(n21419) );
  NAND U22189 ( .A(n21417), .B(n21416), .Z(n21418) );
  NAND U22190 ( .A(n21419), .B(n21418), .Z(n21626) );
  NANDN U22191 ( .A(n21421), .B(n21420), .Z(n21425) );
  NAND U22192 ( .A(n21423), .B(n21422), .Z(n21424) );
  NAND U22193 ( .A(n21425), .B(n21424), .Z(n21830) );
  XOR U22194 ( .A(b[41]), .B(a[63]), .Z(n21704) );
  NANDN U22195 ( .A(n36905), .B(n21704), .Z(n21428) );
  NAND U22196 ( .A(n21426), .B(n36807), .Z(n21427) );
  NAND U22197 ( .A(n21428), .B(n21427), .Z(n21731) );
  XOR U22198 ( .A(b[57]), .B(n23149), .Z(n21707) );
  OR U22199 ( .A(n21707), .B(n965), .Z(n21431) );
  NANDN U22200 ( .A(n21429), .B(n38194), .Z(n21430) );
  NAND U22201 ( .A(n21431), .B(n21430), .Z(n21728) );
  NAND U22202 ( .A(n38326), .B(n21432), .Z(n21434) );
  XOR U22203 ( .A(n38400), .B(n22579), .Z(n21710) );
  NANDN U22204 ( .A(n38273), .B(n21710), .Z(n21433) );
  AND U22205 ( .A(n21434), .B(n21433), .Z(n21729) );
  XNOR U22206 ( .A(n21728), .B(n21729), .Z(n21730) );
  XOR U22207 ( .A(n21731), .B(n21730), .Z(n21828) );
  XOR U22208 ( .A(b[33]), .B(n30543), .Z(n21713) );
  NANDN U22209 ( .A(n21713), .B(n35620), .Z(n21437) );
  NANDN U22210 ( .A(n21435), .B(n35621), .Z(n21436) );
  NAND U22211 ( .A(n21437), .B(n21436), .Z(n21826) );
  NANDN U22212 ( .A(n966), .B(a[103]), .Z(n21438) );
  XOR U22213 ( .A(n29232), .B(n21438), .Z(n21440) );
  IV U22214 ( .A(a[102]), .Z(n36420) );
  NANDN U22215 ( .A(n36420), .B(n966), .Z(n21439) );
  AND U22216 ( .A(n21440), .B(n21439), .Z(n21823) );
  XOR U22217 ( .A(b[63]), .B(n21441), .Z(n21719) );
  NANDN U22218 ( .A(n21719), .B(n38422), .Z(n21444) );
  NANDN U22219 ( .A(n21442), .B(n38423), .Z(n21443) );
  AND U22220 ( .A(n21444), .B(n21443), .Z(n21824) );
  XNOR U22221 ( .A(n21823), .B(n21824), .Z(n21825) );
  XNOR U22222 ( .A(n21826), .B(n21825), .Z(n21827) );
  XOR U22223 ( .A(n21828), .B(n21827), .Z(n21829) );
  XNOR U22224 ( .A(n21830), .B(n21829), .Z(n21624) );
  NANDN U22225 ( .A(n21446), .B(n21445), .Z(n21450) );
  NAND U22226 ( .A(n21448), .B(n21447), .Z(n21449) );
  AND U22227 ( .A(n21450), .B(n21449), .Z(n21623) );
  XNOR U22228 ( .A(n21624), .B(n21623), .Z(n21625) );
  XNOR U22229 ( .A(n21626), .B(n21625), .Z(n21734) );
  XNOR U22230 ( .A(n21735), .B(n21734), .Z(n21737) );
  XNOR U22231 ( .A(n21736), .B(n21737), .Z(n21836) );
  XNOR U22232 ( .A(n21835), .B(n21836), .Z(n21613) );
  NAND U22233 ( .A(n21452), .B(n21451), .Z(n21456) );
  NANDN U22234 ( .A(n21454), .B(n21453), .Z(n21455) );
  NAND U22235 ( .A(n21456), .B(n21455), .Z(n21842) );
  OR U22236 ( .A(n21458), .B(n21457), .Z(n21462) );
  OR U22237 ( .A(n21460), .B(n21459), .Z(n21461) );
  NAND U22238 ( .A(n21462), .B(n21461), .Z(n21846) );
  XOR U22239 ( .A(a[93]), .B(n970), .Z(n21740) );
  OR U22240 ( .A(n21740), .B(n31369), .Z(n21465) );
  NANDN U22241 ( .A(n21463), .B(n31119), .Z(n21464) );
  NAND U22242 ( .A(n21465), .B(n21464), .Z(n21761) );
  XOR U22243 ( .A(b[43]), .B(n27773), .Z(n21743) );
  NANDN U22244 ( .A(n21743), .B(n37068), .Z(n21468) );
  NANDN U22245 ( .A(n21466), .B(n37069), .Z(n21467) );
  NAND U22246 ( .A(n21468), .B(n21467), .Z(n21758) );
  XOR U22247 ( .A(b[45]), .B(a[59]), .Z(n21746) );
  NAND U22248 ( .A(n21746), .B(n37261), .Z(n21471) );
  NANDN U22249 ( .A(n21469), .B(n37262), .Z(n21470) );
  AND U22250 ( .A(n21471), .B(n21470), .Z(n21759) );
  XNOR U22251 ( .A(n21758), .B(n21759), .Z(n21760) );
  XNOR U22252 ( .A(n21761), .B(n21760), .Z(n21689) );
  NAND U22253 ( .A(n37652), .B(n21472), .Z(n21474) );
  XOR U22254 ( .A(b[49]), .B(n25466), .Z(n21749) );
  OR U22255 ( .A(n21749), .B(n37756), .Z(n21473) );
  NAND U22256 ( .A(n21474), .B(n21473), .Z(n21785) );
  NANDN U22257 ( .A(n21475), .B(n37469), .Z(n21477) );
  XNOR U22258 ( .A(n978), .B(a[57]), .Z(n21752) );
  NAND U22259 ( .A(n21752), .B(n37471), .Z(n21476) );
  NAND U22260 ( .A(n21477), .B(n21476), .Z(n21783) );
  NAND U22261 ( .A(n30846), .B(n21478), .Z(n21480) );
  XNOR U22262 ( .A(n35628), .B(b[9]), .Z(n21755) );
  NAND U22263 ( .A(n30509), .B(n21755), .Z(n21479) );
  NAND U22264 ( .A(n21480), .B(n21479), .Z(n21784) );
  XNOR U22265 ( .A(n21783), .B(n21784), .Z(n21786) );
  XOR U22266 ( .A(n21785), .B(n21786), .Z(n21686) );
  NANDN U22267 ( .A(n21482), .B(n21481), .Z(n21486) );
  NAND U22268 ( .A(n21484), .B(n21483), .Z(n21485) );
  NAND U22269 ( .A(n21486), .B(n21485), .Z(n21687) );
  XNOR U22270 ( .A(n21686), .B(n21687), .Z(n21688) );
  XOR U22271 ( .A(n21689), .B(n21688), .Z(n21845) );
  XNOR U22272 ( .A(n21846), .B(n21845), .Z(n21848) );
  XOR U22273 ( .A(b[35]), .B(a[69]), .Z(n21768) );
  NAND U22274 ( .A(n35985), .B(n21768), .Z(n21489) );
  NANDN U22275 ( .A(n21487), .B(n35986), .Z(n21488) );
  NAND U22276 ( .A(n21489), .B(n21488), .Z(n21820) );
  XNOR U22277 ( .A(a[97]), .B(n31123), .Z(n21771) );
  NAND U22278 ( .A(n21771), .B(n29949), .Z(n21492) );
  NAND U22279 ( .A(n29948), .B(n21490), .Z(n21491) );
  NAND U22280 ( .A(n21492), .B(n21491), .Z(n21817) );
  XOR U22281 ( .A(b[55]), .B(n23852), .Z(n21774) );
  NANDN U22282 ( .A(n21774), .B(n38075), .Z(n21495) );
  NANDN U22283 ( .A(n21493), .B(n38073), .Z(n21494) );
  AND U22284 ( .A(n21495), .B(n21494), .Z(n21818) );
  XNOR U22285 ( .A(n21817), .B(n21818), .Z(n21819) );
  XNOR U22286 ( .A(n21820), .B(n21819), .Z(n21620) );
  NANDN U22287 ( .A(n21497), .B(n21496), .Z(n21501) );
  NAND U22288 ( .A(n21499), .B(n21498), .Z(n21500) );
  NAND U22289 ( .A(n21501), .B(n21500), .Z(n21617) );
  NANDN U22290 ( .A(n21503), .B(n21502), .Z(n21507) );
  NAND U22291 ( .A(n21505), .B(n21504), .Z(n21506) );
  NAND U22292 ( .A(n21507), .B(n21506), .Z(n21618) );
  XNOR U22293 ( .A(n21617), .B(n21618), .Z(n21619) );
  XOR U22294 ( .A(n21620), .B(n21619), .Z(n21847) );
  XOR U22295 ( .A(n21848), .B(n21847), .Z(n21840) );
  NANDN U22296 ( .A(n21513), .B(n21512), .Z(n21517) );
  NAND U22297 ( .A(n21515), .B(n21514), .Z(n21516) );
  NAND U22298 ( .A(n21517), .B(n21516), .Z(n21852) );
  XNOR U22299 ( .A(n21851), .B(n21852), .Z(n21853) );
  NANDN U22300 ( .A(n21519), .B(n21518), .Z(n21523) );
  NAND U22301 ( .A(n21521), .B(n21520), .Z(n21522) );
  NAND U22302 ( .A(n21523), .B(n21522), .Z(n21790) );
  XNOR U22303 ( .A(a[89]), .B(b[15]), .Z(n21793) );
  OR U22304 ( .A(n21793), .B(n32010), .Z(n21526) );
  NANDN U22305 ( .A(n21524), .B(n32011), .Z(n21525) );
  NAND U22306 ( .A(n21526), .B(n21525), .Z(n21653) );
  XOR U22307 ( .A(b[25]), .B(a[79]), .Z(n21796) );
  NANDN U22308 ( .A(n34219), .B(n21796), .Z(n21529) );
  NAND U22309 ( .A(n34217), .B(n21527), .Z(n21528) );
  NAND U22310 ( .A(n21529), .B(n21528), .Z(n21650) );
  XOR U22311 ( .A(a[87]), .B(b[17]), .Z(n21799) );
  NAND U22312 ( .A(n21799), .B(n32543), .Z(n21532) );
  NANDN U22313 ( .A(n21530), .B(n32541), .Z(n21531) );
  AND U22314 ( .A(n21532), .B(n21531), .Z(n21651) );
  XNOR U22315 ( .A(n21650), .B(n21651), .Z(n21652) );
  XNOR U22316 ( .A(n21653), .B(n21652), .Z(n21692) );
  XOR U22317 ( .A(b[39]), .B(n28403), .Z(n21802) );
  NANDN U22318 ( .A(n21802), .B(n36553), .Z(n21535) );
  NANDN U22319 ( .A(n21533), .B(n36643), .Z(n21534) );
  NAND U22320 ( .A(n21535), .B(n21534), .Z(n21683) );
  XOR U22321 ( .A(b[51]), .B(n25001), .Z(n21805) );
  NANDN U22322 ( .A(n21805), .B(n37803), .Z(n21538) );
  NANDN U22323 ( .A(n21536), .B(n37802), .Z(n21537) );
  NAND U22324 ( .A(n21538), .B(n21537), .Z(n21680) );
  XOR U22325 ( .A(b[53]), .B(n24288), .Z(n21808) );
  NANDN U22326 ( .A(n21808), .B(n37940), .Z(n21541) );
  NANDN U22327 ( .A(n21539), .B(n37941), .Z(n21540) );
  AND U22328 ( .A(n21541), .B(n21540), .Z(n21681) );
  XNOR U22329 ( .A(n21680), .B(n21681), .Z(n21682) );
  XOR U22330 ( .A(n21683), .B(n21682), .Z(n21693) );
  XOR U22331 ( .A(n21692), .B(n21693), .Z(n21695) );
  NANDN U22332 ( .A(n21543), .B(n21542), .Z(n21547) );
  NAND U22333 ( .A(n21545), .B(n21544), .Z(n21546) );
  AND U22334 ( .A(n21547), .B(n21546), .Z(n21694) );
  XOR U22335 ( .A(n21695), .B(n21694), .Z(n21788) );
  NANDN U22336 ( .A(n21549), .B(n21548), .Z(n21553) );
  NAND U22337 ( .A(n21551), .B(n21550), .Z(n21552) );
  AND U22338 ( .A(n21553), .B(n21552), .Z(n21787) );
  XNOR U22339 ( .A(n21788), .B(n21787), .Z(n21789) );
  XOR U22340 ( .A(n21790), .B(n21789), .Z(n21854) );
  XNOR U22341 ( .A(n21853), .B(n21854), .Z(n21839) );
  XNOR U22342 ( .A(n21840), .B(n21839), .Z(n21841) );
  XOR U22343 ( .A(n21842), .B(n21841), .Z(n21614) );
  XNOR U22344 ( .A(n21613), .B(n21614), .Z(n21615) );
  NAND U22345 ( .A(n21555), .B(n21554), .Z(n21559) );
  NANDN U22346 ( .A(n21557), .B(n21556), .Z(n21558) );
  NAND U22347 ( .A(n21559), .B(n21558), .Z(n21616) );
  XOR U22348 ( .A(n21615), .B(n21616), .Z(n21864) );
  NANDN U22349 ( .A(n21561), .B(n21560), .Z(n21565) );
  NAND U22350 ( .A(n21563), .B(n21562), .Z(n21564) );
  AND U22351 ( .A(n21565), .B(n21564), .Z(n21861) );
  NAND U22352 ( .A(n21567), .B(n21566), .Z(n21571) );
  NANDN U22353 ( .A(n21569), .B(n21568), .Z(n21570) );
  NAND U22354 ( .A(n21571), .B(n21570), .Z(n21610) );
  XNOR U22355 ( .A(n21607), .B(n21608), .Z(n21609) );
  XNOR U22356 ( .A(n21610), .B(n21609), .Z(n21862) );
  XNOR U22357 ( .A(n21864), .B(n21863), .Z(n21870) );
  XOR U22358 ( .A(n21869), .B(n21870), .Z(n21876) );
  OR U22359 ( .A(n21581), .B(n21580), .Z(n21585) );
  NAND U22360 ( .A(n21583), .B(n21582), .Z(n21584) );
  NAND U22361 ( .A(n21585), .B(n21584), .Z(n21874) );
  NANDN U22362 ( .A(n21587), .B(n21586), .Z(n21591) );
  NANDN U22363 ( .A(n21589), .B(n21588), .Z(n21590) );
  AND U22364 ( .A(n21591), .B(n21590), .Z(n21873) );
  XNOR U22365 ( .A(n21874), .B(n21873), .Z(n21875) );
  XNOR U22366 ( .A(n21876), .B(n21875), .Z(n21603) );
  NANDN U22367 ( .A(n21593), .B(n21592), .Z(n21597) );
  NANDN U22368 ( .A(n21595), .B(n21594), .Z(n21596) );
  NAND U22369 ( .A(n21597), .B(n21596), .Z(n21604) );
  XNOR U22370 ( .A(n21603), .B(n21604), .Z(n21605) );
  XNOR U22371 ( .A(n21606), .B(n21605), .Z(n21879) );
  XNOR U22372 ( .A(n21879), .B(sreg[167]), .Z(n21881) );
  NAND U22373 ( .A(n21598), .B(sreg[166]), .Z(n21602) );
  OR U22374 ( .A(n21600), .B(n21599), .Z(n21601) );
  AND U22375 ( .A(n21602), .B(n21601), .Z(n21880) );
  XOR U22376 ( .A(n21881), .B(n21880), .Z(c[167]) );
  NANDN U22377 ( .A(n21608), .B(n21607), .Z(n21612) );
  NAND U22378 ( .A(n21610), .B(n21609), .Z(n21611) );
  NAND U22379 ( .A(n21612), .B(n21611), .Z(n22155) );
  XNOR U22380 ( .A(n22155), .B(n22156), .Z(n22157) );
  NANDN U22381 ( .A(n21618), .B(n21617), .Z(n21622) );
  NAND U22382 ( .A(n21620), .B(n21619), .Z(n21621) );
  AND U22383 ( .A(n21622), .B(n21621), .Z(n22126) );
  NANDN U22384 ( .A(n21624), .B(n21623), .Z(n21628) );
  NANDN U22385 ( .A(n21626), .B(n21625), .Z(n21627) );
  NAND U22386 ( .A(n21628), .B(n21627), .Z(n22123) );
  NANDN U22387 ( .A(n21630), .B(n21629), .Z(n21634) );
  NAND U22388 ( .A(n21632), .B(n21631), .Z(n21633) );
  AND U22389 ( .A(n21634), .B(n21633), .Z(n22124) );
  XNOR U22390 ( .A(n22123), .B(n22124), .Z(n22125) );
  XNOR U22391 ( .A(n22126), .B(n22125), .Z(n22111) );
  NANDN U22392 ( .A(n21636), .B(n21635), .Z(n21640) );
  OR U22393 ( .A(n21638), .B(n21637), .Z(n21639) );
  AND U22394 ( .A(n21640), .B(n21639), .Z(n22112) );
  XNOR U22395 ( .A(n22111), .B(n22112), .Z(n22114) );
  NAND U22396 ( .A(n33283), .B(n21641), .Z(n21643) );
  XOR U22397 ( .A(n33628), .B(n33020), .Z(n21954) );
  NANDN U22398 ( .A(n33021), .B(n21954), .Z(n21642) );
  NAND U22399 ( .A(n21643), .B(n21642), .Z(n21978) );
  XNOR U22400 ( .A(b[21]), .B(a[84]), .Z(n21957) );
  OR U22401 ( .A(n21957), .B(n33634), .Z(n21646) );
  NAND U22402 ( .A(n21644), .B(n33464), .Z(n21645) );
  NAND U22403 ( .A(n21646), .B(n21645), .Z(n21975) );
  NAND U22404 ( .A(n34044), .B(n21647), .Z(n21649) );
  XOR U22405 ( .A(n34510), .B(n32815), .Z(n21960) );
  NANDN U22406 ( .A(n33867), .B(n21960), .Z(n21648) );
  AND U22407 ( .A(n21649), .B(n21648), .Z(n21976) );
  XNOR U22408 ( .A(n21975), .B(n21976), .Z(n21977) );
  XOR U22409 ( .A(n21978), .B(n21977), .Z(n22012) );
  NANDN U22410 ( .A(n21651), .B(n21650), .Z(n21655) );
  NAND U22411 ( .A(n21653), .B(n21652), .Z(n21654) );
  NAND U22412 ( .A(n21655), .B(n21654), .Z(n22013) );
  XNOR U22413 ( .A(n22012), .B(n22013), .Z(n22015) );
  NAND U22414 ( .A(a[40]), .B(b[63]), .Z(n22054) );
  NANDN U22415 ( .A(n21656), .B(n38369), .Z(n21658) );
  XOR U22416 ( .A(b[61]), .B(n22289), .Z(n21948) );
  OR U22417 ( .A(n21948), .B(n38371), .Z(n21657) );
  NAND U22418 ( .A(n21658), .B(n21657), .Z(n22052) );
  NANDN U22419 ( .A(n21659), .B(n35311), .Z(n21661) );
  XOR U22420 ( .A(b[31]), .B(n31372), .Z(n21951) );
  NANDN U22421 ( .A(n21951), .B(n35313), .Z(n21660) );
  AND U22422 ( .A(n21661), .B(n21660), .Z(n22051) );
  XNOR U22423 ( .A(n22052), .B(n22051), .Z(n22053) );
  XNOR U22424 ( .A(n22054), .B(n22053), .Z(n22014) );
  XNOR U22425 ( .A(n22015), .B(n22014), .Z(n21888) );
  XOR U22426 ( .A(b[37]), .B(n29868), .Z(n21918) );
  NANDN U22427 ( .A(n21918), .B(n36311), .Z(n21664) );
  NANDN U22428 ( .A(n21662), .B(n36309), .Z(n21663) );
  NAND U22429 ( .A(n21664), .B(n21663), .Z(n21972) );
  XOR U22430 ( .A(a[100]), .B(n968), .Z(n21921) );
  OR U22431 ( .A(n21921), .B(n29363), .Z(n21667) );
  NANDN U22432 ( .A(n21665), .B(n29864), .Z(n21666) );
  NAND U22433 ( .A(n21667), .B(n21666), .Z(n21969) );
  XOR U22434 ( .A(n36420), .B(n967), .Z(n21924) );
  NAND U22435 ( .A(n21924), .B(n28939), .Z(n21670) );
  NAND U22436 ( .A(n28938), .B(n21668), .Z(n21669) );
  AND U22437 ( .A(n21670), .B(n21669), .Z(n21970) );
  XNOR U22438 ( .A(n21969), .B(n21970), .Z(n21971) );
  XOR U22439 ( .A(n21972), .B(n21971), .Z(n21909) );
  XOR U22440 ( .A(a[92]), .B(n971), .Z(n21927) );
  OR U22441 ( .A(n21927), .B(n31550), .Z(n21673) );
  NANDN U22442 ( .A(n21671), .B(n31874), .Z(n21672) );
  NAND U22443 ( .A(n21673), .B(n21672), .Z(n22084) );
  NAND U22444 ( .A(n34848), .B(n21674), .Z(n21676) );
  XOR U22445 ( .A(n35375), .B(n31870), .Z(n21930) );
  NAND U22446 ( .A(n34618), .B(n21930), .Z(n21675) );
  NAND U22447 ( .A(n21676), .B(n21675), .Z(n22081) );
  NAND U22448 ( .A(n35188), .B(n21677), .Z(n21679) );
  XOR U22449 ( .A(n35540), .B(n31363), .Z(n21933) );
  NANDN U22450 ( .A(n34968), .B(n21933), .Z(n21678) );
  AND U22451 ( .A(n21679), .B(n21678), .Z(n22082) );
  XNOR U22452 ( .A(n22081), .B(n22082), .Z(n22083) );
  XOR U22453 ( .A(n22084), .B(n22083), .Z(n21907) );
  NANDN U22454 ( .A(n21681), .B(n21680), .Z(n21685) );
  NAND U22455 ( .A(n21683), .B(n21682), .Z(n21684) );
  AND U22456 ( .A(n21685), .B(n21684), .Z(n21906) );
  XOR U22457 ( .A(n21907), .B(n21906), .Z(n21908) );
  XOR U22458 ( .A(n21909), .B(n21908), .Z(n21889) );
  XOR U22459 ( .A(n21888), .B(n21889), .Z(n21891) );
  NANDN U22460 ( .A(n21687), .B(n21686), .Z(n21691) );
  NAND U22461 ( .A(n21689), .B(n21688), .Z(n21690) );
  NAND U22462 ( .A(n21691), .B(n21690), .Z(n21890) );
  XNOR U22463 ( .A(n21891), .B(n21890), .Z(n22008) );
  NANDN U22464 ( .A(n21693), .B(n21692), .Z(n21697) );
  NANDN U22465 ( .A(n21695), .B(n21694), .Z(n21696) );
  NAND U22466 ( .A(n21697), .B(n21696), .Z(n22007) );
  NANDN U22467 ( .A(n21699), .B(n21698), .Z(n21703) );
  NAND U22468 ( .A(n21701), .B(n21700), .Z(n21702) );
  NAND U22469 ( .A(n21703), .B(n21702), .Z(n21903) );
  XOR U22470 ( .A(b[41]), .B(a[64]), .Z(n21981) );
  NANDN U22471 ( .A(n36905), .B(n21981), .Z(n21706) );
  NAND U22472 ( .A(n21704), .B(n36807), .Z(n21705) );
  NAND U22473 ( .A(n21706), .B(n21705), .Z(n22003) );
  XOR U22474 ( .A(b[57]), .B(n23447), .Z(n21984) );
  OR U22475 ( .A(n21984), .B(n965), .Z(n21709) );
  NANDN U22476 ( .A(n21707), .B(n38194), .Z(n21708) );
  NAND U22477 ( .A(n21709), .B(n21708), .Z(n22000) );
  NAND U22478 ( .A(n38326), .B(n21710), .Z(n21712) );
  XOR U22479 ( .A(n38400), .B(n22964), .Z(n21987) );
  NANDN U22480 ( .A(n38273), .B(n21987), .Z(n21711) );
  AND U22481 ( .A(n21712), .B(n21711), .Z(n22001) );
  XNOR U22482 ( .A(n22000), .B(n22001), .Z(n22002) );
  XOR U22483 ( .A(n22003), .B(n22002), .Z(n22099) );
  XOR U22484 ( .A(b[33]), .B(n30210), .Z(n21990) );
  NANDN U22485 ( .A(n21990), .B(n35620), .Z(n21715) );
  NANDN U22486 ( .A(n21713), .B(n35621), .Z(n21714) );
  NAND U22487 ( .A(n21715), .B(n21714), .Z(n22096) );
  NANDN U22488 ( .A(n966), .B(a[104]), .Z(n21716) );
  XOR U22489 ( .A(n29232), .B(n21716), .Z(n21718) );
  NANDN U22490 ( .A(b[0]), .B(a[103]), .Z(n21717) );
  AND U22491 ( .A(n21718), .B(n21717), .Z(n22093) );
  XOR U22492 ( .A(b[63]), .B(n22246), .Z(n21997) );
  NANDN U22493 ( .A(n21997), .B(n38422), .Z(n21721) );
  NANDN U22494 ( .A(n21719), .B(n38423), .Z(n21720) );
  AND U22495 ( .A(n21721), .B(n21720), .Z(n22094) );
  XNOR U22496 ( .A(n22093), .B(n22094), .Z(n22095) );
  XOR U22497 ( .A(n22096), .B(n22095), .Z(n22100) );
  XNOR U22498 ( .A(n22099), .B(n22100), .Z(n22102) );
  NANDN U22499 ( .A(n21723), .B(n21722), .Z(n21727) );
  NAND U22500 ( .A(n21725), .B(n21724), .Z(n21726) );
  NAND U22501 ( .A(n21727), .B(n21726), .Z(n22101) );
  XOR U22502 ( .A(n22102), .B(n22101), .Z(n21900) );
  NANDN U22503 ( .A(n21729), .B(n21728), .Z(n21733) );
  NAND U22504 ( .A(n21731), .B(n21730), .Z(n21732) );
  AND U22505 ( .A(n21733), .B(n21732), .Z(n21901) );
  XOR U22506 ( .A(n21900), .B(n21901), .Z(n21902) );
  XNOR U22507 ( .A(n21903), .B(n21902), .Z(n22006) );
  XNOR U22508 ( .A(n22007), .B(n22006), .Z(n22009) );
  XNOR U22509 ( .A(n22008), .B(n22009), .Z(n22113) );
  XOR U22510 ( .A(n22114), .B(n22113), .Z(n22143) );
  NAND U22511 ( .A(n21735), .B(n21734), .Z(n21739) );
  NANDN U22512 ( .A(n21737), .B(n21736), .Z(n21738) );
  NAND U22513 ( .A(n21739), .B(n21738), .Z(n22134) );
  XOR U22514 ( .A(a[94]), .B(n970), .Z(n22018) );
  OR U22515 ( .A(n22018), .B(n31369), .Z(n21742) );
  NANDN U22516 ( .A(n21740), .B(n31119), .Z(n21741) );
  NAND U22517 ( .A(n21742), .B(n21741), .Z(n22039) );
  XNOR U22518 ( .A(b[43]), .B(a[62]), .Z(n22021) );
  NANDN U22519 ( .A(n22021), .B(n37068), .Z(n21745) );
  NANDN U22520 ( .A(n21743), .B(n37069), .Z(n21744) );
  NAND U22521 ( .A(n21745), .B(n21744), .Z(n22036) );
  XNOR U22522 ( .A(b[45]), .B(a[60]), .Z(n22024) );
  NANDN U22523 ( .A(n22024), .B(n37261), .Z(n21748) );
  NAND U22524 ( .A(n21746), .B(n37262), .Z(n21747) );
  AND U22525 ( .A(n21748), .B(n21747), .Z(n22037) );
  XNOR U22526 ( .A(n22036), .B(n22037), .Z(n22038) );
  XNOR U22527 ( .A(n22039), .B(n22038), .Z(n21912) );
  XOR U22528 ( .A(b[49]), .B(n25860), .Z(n22027) );
  OR U22529 ( .A(n22027), .B(n37756), .Z(n21751) );
  NANDN U22530 ( .A(n21749), .B(n37652), .Z(n21750) );
  NAND U22531 ( .A(n21751), .B(n21750), .Z(n22060) );
  NAND U22532 ( .A(n21752), .B(n37469), .Z(n21754) );
  XOR U22533 ( .A(n978), .B(n26347), .Z(n22030) );
  NAND U22534 ( .A(n22030), .B(n37471), .Z(n21753) );
  NAND U22535 ( .A(n21754), .B(n21753), .Z(n22057) );
  XOR U22536 ( .A(a[96]), .B(n969), .Z(n22033) );
  NANDN U22537 ( .A(n22033), .B(n30509), .Z(n21757) );
  NAND U22538 ( .A(n21755), .B(n30846), .Z(n21756) );
  AND U22539 ( .A(n21757), .B(n21756), .Z(n22058) );
  XNOR U22540 ( .A(n22057), .B(n22058), .Z(n22059) );
  XOR U22541 ( .A(n22060), .B(n22059), .Z(n21913) );
  XNOR U22542 ( .A(n21912), .B(n21913), .Z(n21914) );
  NANDN U22543 ( .A(n21759), .B(n21758), .Z(n21763) );
  NAND U22544 ( .A(n21761), .B(n21760), .Z(n21762) );
  AND U22545 ( .A(n21763), .B(n21762), .Z(n21915) );
  XNOR U22546 ( .A(n21914), .B(n21915), .Z(n22118) );
  XNOR U22547 ( .A(n22118), .B(n22117), .Z(n22119) );
  XNOR U22548 ( .A(b[35]), .B(a[70]), .Z(n22042) );
  NANDN U22549 ( .A(n22042), .B(n35985), .Z(n21770) );
  NAND U22550 ( .A(n21768), .B(n35986), .Z(n21769) );
  NAND U22551 ( .A(n21770), .B(n21769), .Z(n22090) );
  XOR U22552 ( .A(n35783), .B(n31123), .Z(n22045) );
  NAND U22553 ( .A(n22045), .B(n29949), .Z(n21773) );
  NAND U22554 ( .A(n29948), .B(n21771), .Z(n21772) );
  NAND U22555 ( .A(n21773), .B(n21772), .Z(n22087) );
  XOR U22556 ( .A(b[55]), .B(n24671), .Z(n22048) );
  NANDN U22557 ( .A(n22048), .B(n38075), .Z(n21776) );
  NANDN U22558 ( .A(n21774), .B(n38073), .Z(n21775) );
  AND U22559 ( .A(n21776), .B(n21775), .Z(n22088) );
  XNOR U22560 ( .A(n22087), .B(n22088), .Z(n22089) );
  XNOR U22561 ( .A(n22090), .B(n22089), .Z(n21897) );
  NANDN U22562 ( .A(n21778), .B(n21777), .Z(n21782) );
  NAND U22563 ( .A(n21780), .B(n21779), .Z(n21781) );
  NAND U22564 ( .A(n21782), .B(n21781), .Z(n21894) );
  XNOR U22565 ( .A(n21894), .B(n21895), .Z(n21896) );
  XOR U22566 ( .A(n21897), .B(n21896), .Z(n22120) );
  XOR U22567 ( .A(n22119), .B(n22120), .Z(n22131) );
  NANDN U22568 ( .A(n21788), .B(n21787), .Z(n21792) );
  NANDN U22569 ( .A(n21790), .B(n21789), .Z(n21791) );
  NAND U22570 ( .A(n21792), .B(n21791), .Z(n22130) );
  XOR U22571 ( .A(a[90]), .B(n972), .Z(n22063) );
  OR U22572 ( .A(n22063), .B(n32010), .Z(n21795) );
  NANDN U22573 ( .A(n21793), .B(n32011), .Z(n21794) );
  NAND U22574 ( .A(n21795), .B(n21794), .Z(n21945) );
  XNOR U22575 ( .A(b[25]), .B(n32814), .Z(n22066) );
  NANDN U22576 ( .A(n34219), .B(n22066), .Z(n21798) );
  NAND U22577 ( .A(n34217), .B(n21796), .Z(n21797) );
  NAND U22578 ( .A(n21798), .B(n21797), .Z(n21942) );
  XNOR U22579 ( .A(a[88]), .B(b[17]), .Z(n22069) );
  NANDN U22580 ( .A(n22069), .B(n32543), .Z(n21801) );
  NAND U22581 ( .A(n21799), .B(n32541), .Z(n21800) );
  AND U22582 ( .A(n21801), .B(n21800), .Z(n21943) );
  XNOR U22583 ( .A(n21942), .B(n21943), .Z(n21944) );
  XNOR U22584 ( .A(n21945), .B(n21944), .Z(n21963) );
  XOR U22585 ( .A(b[39]), .B(n28701), .Z(n22072) );
  NANDN U22586 ( .A(n22072), .B(n36553), .Z(n21804) );
  NANDN U22587 ( .A(n21802), .B(n36643), .Z(n21803) );
  NAND U22588 ( .A(n21804), .B(n21803), .Z(n21939) );
  XOR U22589 ( .A(b[51]), .B(n25177), .Z(n22075) );
  NANDN U22590 ( .A(n22075), .B(n37803), .Z(n21807) );
  NANDN U22591 ( .A(n21805), .B(n37802), .Z(n21806) );
  NAND U22592 ( .A(n21807), .B(n21806), .Z(n21936) );
  XOR U22593 ( .A(b[53]), .B(n25134), .Z(n22078) );
  NANDN U22594 ( .A(n22078), .B(n37940), .Z(n21810) );
  NANDN U22595 ( .A(n21808), .B(n37941), .Z(n21809) );
  AND U22596 ( .A(n21810), .B(n21809), .Z(n21937) );
  XNOR U22597 ( .A(n21936), .B(n21937), .Z(n21938) );
  XOR U22598 ( .A(n21939), .B(n21938), .Z(n21964) );
  XOR U22599 ( .A(n21963), .B(n21964), .Z(n21966) );
  NANDN U22600 ( .A(n21812), .B(n21811), .Z(n21816) );
  NAND U22601 ( .A(n21814), .B(n21813), .Z(n21815) );
  NAND U22602 ( .A(n21816), .B(n21815), .Z(n21965) );
  XNOR U22603 ( .A(n21966), .B(n21965), .Z(n22108) );
  NANDN U22604 ( .A(n21818), .B(n21817), .Z(n21822) );
  NAND U22605 ( .A(n21820), .B(n21819), .Z(n21821) );
  NAND U22606 ( .A(n21822), .B(n21821), .Z(n22105) );
  XNOR U22607 ( .A(n22105), .B(n22106), .Z(n22107) );
  XNOR U22608 ( .A(n22108), .B(n22107), .Z(n22127) );
  NANDN U22609 ( .A(n21828), .B(n21827), .Z(n21832) );
  OR U22610 ( .A(n21830), .B(n21829), .Z(n21831) );
  AND U22611 ( .A(n21832), .B(n21831), .Z(n22128) );
  XNOR U22612 ( .A(n22127), .B(n22128), .Z(n22129) );
  XNOR U22613 ( .A(n22130), .B(n22129), .Z(n22132) );
  XNOR U22614 ( .A(n22131), .B(n22132), .Z(n22133) );
  XOR U22615 ( .A(n22134), .B(n22133), .Z(n22144) );
  XNOR U22616 ( .A(n22143), .B(n22144), .Z(n22145) );
  OR U22617 ( .A(n21834), .B(n21833), .Z(n21838) );
  NAND U22618 ( .A(n21836), .B(n21835), .Z(n21837) );
  NAND U22619 ( .A(n21838), .B(n21837), .Z(n22146) );
  XOR U22620 ( .A(n22145), .B(n22146), .Z(n22152) );
  NANDN U22621 ( .A(n21840), .B(n21839), .Z(n21844) );
  NAND U22622 ( .A(n21842), .B(n21841), .Z(n21843) );
  AND U22623 ( .A(n21844), .B(n21843), .Z(n22149) );
  NAND U22624 ( .A(n21846), .B(n21845), .Z(n21850) );
  NANDN U22625 ( .A(n21848), .B(n21847), .Z(n21849) );
  NAND U22626 ( .A(n21850), .B(n21849), .Z(n22140) );
  NANDN U22627 ( .A(n21852), .B(n21851), .Z(n21856) );
  NANDN U22628 ( .A(n21854), .B(n21853), .Z(n21855) );
  NAND U22629 ( .A(n21856), .B(n21855), .Z(n22137) );
  XNOR U22630 ( .A(n22137), .B(n22138), .Z(n22139) );
  XNOR U22631 ( .A(n22140), .B(n22139), .Z(n22150) );
  XNOR U22632 ( .A(n22152), .B(n22151), .Z(n22158) );
  XOR U22633 ( .A(n22157), .B(n22158), .Z(n22164) );
  OR U22634 ( .A(n21862), .B(n21861), .Z(n21866) );
  NAND U22635 ( .A(n21864), .B(n21863), .Z(n21865) );
  NAND U22636 ( .A(n21866), .B(n21865), .Z(n22162) );
  NANDN U22637 ( .A(n21868), .B(n21867), .Z(n21872) );
  NANDN U22638 ( .A(n21870), .B(n21869), .Z(n21871) );
  AND U22639 ( .A(n21872), .B(n21871), .Z(n22161) );
  XNOR U22640 ( .A(n22162), .B(n22161), .Z(n22163) );
  XNOR U22641 ( .A(n22164), .B(n22163), .Z(n21884) );
  NANDN U22642 ( .A(n21874), .B(n21873), .Z(n21878) );
  NAND U22643 ( .A(n21876), .B(n21875), .Z(n21877) );
  NAND U22644 ( .A(n21878), .B(n21877), .Z(n21885) );
  XNOR U22645 ( .A(n21884), .B(n21885), .Z(n21886) );
  XNOR U22646 ( .A(n21887), .B(n21886), .Z(n22167) );
  XNOR U22647 ( .A(n22167), .B(sreg[168]), .Z(n22169) );
  NAND U22648 ( .A(n21879), .B(sreg[167]), .Z(n21883) );
  OR U22649 ( .A(n21881), .B(n21880), .Z(n21882) );
  AND U22650 ( .A(n21883), .B(n21882), .Z(n22168) );
  XOR U22651 ( .A(n22169), .B(n22168), .Z(c[168]) );
  NANDN U22652 ( .A(n21889), .B(n21888), .Z(n21893) );
  OR U22653 ( .A(n21891), .B(n21890), .Z(n21892) );
  NAND U22654 ( .A(n21893), .B(n21892), .Z(n22406) );
  NANDN U22655 ( .A(n21895), .B(n21894), .Z(n21899) );
  NAND U22656 ( .A(n21897), .B(n21896), .Z(n21898) );
  NAND U22657 ( .A(n21899), .B(n21898), .Z(n22426) );
  NAND U22658 ( .A(n21901), .B(n21900), .Z(n21905) );
  NANDN U22659 ( .A(n21903), .B(n21902), .Z(n21904) );
  NAND U22660 ( .A(n21905), .B(n21904), .Z(n22424) );
  NANDN U22661 ( .A(n21907), .B(n21906), .Z(n21911) );
  OR U22662 ( .A(n21909), .B(n21908), .Z(n21910) );
  AND U22663 ( .A(n21911), .B(n21910), .Z(n22425) );
  XNOR U22664 ( .A(n22424), .B(n22425), .Z(n22427) );
  XNOR U22665 ( .A(n22426), .B(n22427), .Z(n22407) );
  XOR U22666 ( .A(n22406), .B(n22407), .Z(n22408) );
  NANDN U22667 ( .A(n21913), .B(n21912), .Z(n21917) );
  NAND U22668 ( .A(n21915), .B(n21914), .Z(n21916) );
  NAND U22669 ( .A(n21917), .B(n21916), .Z(n22208) );
  XNOR U22670 ( .A(b[37]), .B(a[69]), .Z(n22216) );
  NANDN U22671 ( .A(n22216), .B(n36311), .Z(n21920) );
  NANDN U22672 ( .A(n21918), .B(n36309), .Z(n21919) );
  NAND U22673 ( .A(n21920), .B(n21919), .Z(n22271) );
  XNOR U22674 ( .A(a[101]), .B(b[5]), .Z(n22219) );
  OR U22675 ( .A(n22219), .B(n29363), .Z(n21923) );
  NANDN U22676 ( .A(n21921), .B(n29864), .Z(n21922) );
  NAND U22677 ( .A(n21923), .B(n21922), .Z(n22268) );
  XNOR U22678 ( .A(a[103]), .B(n967), .Z(n22222) );
  NAND U22679 ( .A(n22222), .B(n28939), .Z(n21926) );
  NAND U22680 ( .A(n28938), .B(n21924), .Z(n21925) );
  AND U22681 ( .A(n21926), .B(n21925), .Z(n22269) );
  XNOR U22682 ( .A(n22268), .B(n22269), .Z(n22270) );
  XNOR U22683 ( .A(n22271), .B(n22270), .Z(n22203) );
  XOR U22684 ( .A(a[93]), .B(n971), .Z(n22225) );
  OR U22685 ( .A(n22225), .B(n31550), .Z(n21929) );
  NANDN U22686 ( .A(n21927), .B(n31874), .Z(n21928) );
  NAND U22687 ( .A(n21929), .B(n21928), .Z(n22344) );
  NAND U22688 ( .A(n34848), .B(n21930), .Z(n21932) );
  XNOR U22689 ( .A(n35375), .B(a[79]), .Z(n22228) );
  NAND U22690 ( .A(n34618), .B(n22228), .Z(n21931) );
  NAND U22691 ( .A(n21932), .B(n21931), .Z(n22341) );
  NAND U22692 ( .A(n35188), .B(n21933), .Z(n21935) );
  XNOR U22693 ( .A(n35540), .B(a[77]), .Z(n22231) );
  NANDN U22694 ( .A(n34968), .B(n22231), .Z(n21934) );
  AND U22695 ( .A(n21935), .B(n21934), .Z(n22342) );
  XNOR U22696 ( .A(n22341), .B(n22342), .Z(n22343) );
  XNOR U22697 ( .A(n22344), .B(n22343), .Z(n22200) );
  NANDN U22698 ( .A(n21937), .B(n21936), .Z(n21941) );
  NAND U22699 ( .A(n21939), .B(n21938), .Z(n21940) );
  NAND U22700 ( .A(n21941), .B(n21940), .Z(n22201) );
  XNOR U22701 ( .A(n22200), .B(n22201), .Z(n22202) );
  XOR U22702 ( .A(n22203), .B(n22202), .Z(n22207) );
  NANDN U22703 ( .A(n21943), .B(n21942), .Z(n21947) );
  NAND U22704 ( .A(n21945), .B(n21944), .Z(n21946) );
  NAND U22705 ( .A(n21947), .B(n21946), .Z(n22383) );
  NAND U22706 ( .A(a[41]), .B(b[63]), .Z(n22397) );
  NANDN U22707 ( .A(n21948), .B(n38369), .Z(n21950) );
  XOR U22708 ( .A(b[61]), .B(n22579), .Z(n22247) );
  OR U22709 ( .A(n22247), .B(n38371), .Z(n21949) );
  NAND U22710 ( .A(n21950), .B(n21949), .Z(n22395) );
  NANDN U22711 ( .A(n21951), .B(n35311), .Z(n21953) );
  XNOR U22712 ( .A(b[31]), .B(a[75]), .Z(n22250) );
  NANDN U22713 ( .A(n22250), .B(n35313), .Z(n21952) );
  AND U22714 ( .A(n21953), .B(n21952), .Z(n22394) );
  XNOR U22715 ( .A(n22395), .B(n22394), .Z(n22396) );
  XOR U22716 ( .A(n22397), .B(n22396), .Z(n22381) );
  NAND U22717 ( .A(n33283), .B(n21954), .Z(n21956) );
  XNOR U22718 ( .A(a[87]), .B(n33020), .Z(n22253) );
  NANDN U22719 ( .A(n33021), .B(n22253), .Z(n21955) );
  NAND U22720 ( .A(n21956), .B(n21955), .Z(n22296) );
  XOR U22721 ( .A(b[21]), .B(a[85]), .Z(n22256) );
  NANDN U22722 ( .A(n33634), .B(n22256), .Z(n21959) );
  NANDN U22723 ( .A(n21957), .B(n33464), .Z(n21958) );
  NAND U22724 ( .A(n21959), .B(n21958), .Z(n22293) );
  NAND U22725 ( .A(n34044), .B(n21960), .Z(n21962) );
  XNOR U22726 ( .A(n34510), .B(a[83]), .Z(n22259) );
  NANDN U22727 ( .A(n33867), .B(n22259), .Z(n21961) );
  AND U22728 ( .A(n21962), .B(n21961), .Z(n22294) );
  XNOR U22729 ( .A(n22293), .B(n22294), .Z(n22295) );
  XNOR U22730 ( .A(n22296), .B(n22295), .Z(n22382) );
  XNOR U22731 ( .A(n22381), .B(n22382), .Z(n22384) );
  XNOR U22732 ( .A(n22383), .B(n22384), .Z(n22206) );
  XOR U22733 ( .A(n22207), .B(n22206), .Z(n22209) );
  XNOR U22734 ( .A(n22208), .B(n22209), .Z(n22307) );
  NANDN U22735 ( .A(n21964), .B(n21963), .Z(n21968) );
  OR U22736 ( .A(n21966), .B(n21965), .Z(n21967) );
  NAND U22737 ( .A(n21968), .B(n21967), .Z(n22306) );
  NANDN U22738 ( .A(n21970), .B(n21969), .Z(n21974) );
  NAND U22739 ( .A(n21972), .B(n21971), .Z(n21973) );
  NAND U22740 ( .A(n21974), .B(n21973), .Z(n22197) );
  NANDN U22741 ( .A(n21976), .B(n21975), .Z(n21980) );
  NAND U22742 ( .A(n21978), .B(n21977), .Z(n21979) );
  NAND U22743 ( .A(n21980), .B(n21979), .Z(n22320) );
  XNOR U22744 ( .A(b[41]), .B(a[65]), .Z(n22274) );
  OR U22745 ( .A(n22274), .B(n36905), .Z(n21983) );
  NAND U22746 ( .A(n21981), .B(n36807), .Z(n21982) );
  NAND U22747 ( .A(n21983), .B(n21982), .Z(n22302) );
  XOR U22748 ( .A(b[57]), .B(n23852), .Z(n22277) );
  OR U22749 ( .A(n22277), .B(n965), .Z(n21986) );
  NANDN U22750 ( .A(n21984), .B(n38194), .Z(n21985) );
  NAND U22751 ( .A(n21986), .B(n21985), .Z(n22299) );
  NAND U22752 ( .A(n38326), .B(n21987), .Z(n21989) );
  XOR U22753 ( .A(n38400), .B(n23149), .Z(n22280) );
  NANDN U22754 ( .A(n38273), .B(n22280), .Z(n21988) );
  AND U22755 ( .A(n21989), .B(n21988), .Z(n22300) );
  XNOR U22756 ( .A(n22299), .B(n22300), .Z(n22301) );
  XOR U22757 ( .A(n22302), .B(n22301), .Z(n22318) );
  XNOR U22758 ( .A(b[33]), .B(a[73]), .Z(n22283) );
  NANDN U22759 ( .A(n22283), .B(n35620), .Z(n21992) );
  NANDN U22760 ( .A(n21990), .B(n35621), .Z(n21991) );
  NAND U22761 ( .A(n21992), .B(n21991), .Z(n22356) );
  NANDN U22762 ( .A(n966), .B(a[105]), .Z(n21993) );
  XOR U22763 ( .A(n29232), .B(n21993), .Z(n21995) );
  IV U22764 ( .A(a[104]), .Z(n36647) );
  NANDN U22765 ( .A(n36647), .B(n966), .Z(n21994) );
  AND U22766 ( .A(n21995), .B(n21994), .Z(n22353) );
  XOR U22767 ( .A(b[63]), .B(n21996), .Z(n22290) );
  NANDN U22768 ( .A(n22290), .B(n38422), .Z(n21999) );
  NANDN U22769 ( .A(n21997), .B(n38423), .Z(n21998) );
  AND U22770 ( .A(n21999), .B(n21998), .Z(n22354) );
  XNOR U22771 ( .A(n22353), .B(n22354), .Z(n22355) );
  XNOR U22772 ( .A(n22356), .B(n22355), .Z(n22317) );
  XOR U22773 ( .A(n22318), .B(n22317), .Z(n22319) );
  XNOR U22774 ( .A(n22320), .B(n22319), .Z(n22195) );
  NANDN U22775 ( .A(n22001), .B(n22000), .Z(n22005) );
  NAND U22776 ( .A(n22003), .B(n22002), .Z(n22004) );
  AND U22777 ( .A(n22005), .B(n22004), .Z(n22194) );
  XNOR U22778 ( .A(n22195), .B(n22194), .Z(n22196) );
  XNOR U22779 ( .A(n22197), .B(n22196), .Z(n22305) );
  XNOR U22780 ( .A(n22306), .B(n22305), .Z(n22308) );
  XNOR U22781 ( .A(n22307), .B(n22308), .Z(n22409) );
  XNOR U22782 ( .A(n22408), .B(n22409), .Z(n22184) );
  NAND U22783 ( .A(n22007), .B(n22006), .Z(n22011) );
  NANDN U22784 ( .A(n22009), .B(n22008), .Z(n22010) );
  NAND U22785 ( .A(n22011), .B(n22010), .Z(n22415) );
  OR U22786 ( .A(n22013), .B(n22012), .Z(n22017) );
  OR U22787 ( .A(n22015), .B(n22014), .Z(n22016) );
  NAND U22788 ( .A(n22017), .B(n22016), .Z(n22419) );
  XOR U22789 ( .A(a[95]), .B(n970), .Z(n22357) );
  OR U22790 ( .A(n22357), .B(n31369), .Z(n22020) );
  NANDN U22791 ( .A(n22018), .B(n31119), .Z(n22019) );
  NAND U22792 ( .A(n22020), .B(n22019), .Z(n22378) );
  XNOR U22793 ( .A(b[43]), .B(a[63]), .Z(n22360) );
  NANDN U22794 ( .A(n22360), .B(n37068), .Z(n22023) );
  NANDN U22795 ( .A(n22021), .B(n37069), .Z(n22022) );
  NAND U22796 ( .A(n22023), .B(n22022), .Z(n22375) );
  XNOR U22797 ( .A(b[45]), .B(a[61]), .Z(n22363) );
  NANDN U22798 ( .A(n22363), .B(n37261), .Z(n22026) );
  NANDN U22799 ( .A(n22024), .B(n37262), .Z(n22025) );
  AND U22800 ( .A(n22026), .B(n22025), .Z(n22376) );
  XNOR U22801 ( .A(n22375), .B(n22376), .Z(n22377) );
  XNOR U22802 ( .A(n22378), .B(n22377), .Z(n22215) );
  XOR U22803 ( .A(n979), .B(n26122), .Z(n22366) );
  NANDN U22804 ( .A(n37756), .B(n22366), .Z(n22029) );
  NANDN U22805 ( .A(n22027), .B(n37652), .Z(n22028) );
  NAND U22806 ( .A(n22029), .B(n22028), .Z(n22403) );
  NAND U22807 ( .A(n37469), .B(n22030), .Z(n22032) );
  XNOR U22808 ( .A(b[47]), .B(a[59]), .Z(n22369) );
  NANDN U22809 ( .A(n22369), .B(n37471), .Z(n22031) );
  NAND U22810 ( .A(n22032), .B(n22031), .Z(n22400) );
  XNOR U22811 ( .A(a[97]), .B(n969), .Z(n22372) );
  NAND U22812 ( .A(n30509), .B(n22372), .Z(n22035) );
  NANDN U22813 ( .A(n22033), .B(n30846), .Z(n22034) );
  AND U22814 ( .A(n22035), .B(n22034), .Z(n22401) );
  XNOR U22815 ( .A(n22400), .B(n22401), .Z(n22402) );
  XNOR U22816 ( .A(n22403), .B(n22402), .Z(n22212) );
  NANDN U22817 ( .A(n22037), .B(n22036), .Z(n22041) );
  NAND U22818 ( .A(n22039), .B(n22038), .Z(n22040) );
  NAND U22819 ( .A(n22041), .B(n22040), .Z(n22213) );
  XNOR U22820 ( .A(n22212), .B(n22213), .Z(n22214) );
  XOR U22821 ( .A(n22215), .B(n22214), .Z(n22418) );
  XNOR U22822 ( .A(n22419), .B(n22418), .Z(n22421) );
  XNOR U22823 ( .A(b[35]), .B(a[71]), .Z(n22385) );
  NANDN U22824 ( .A(n22385), .B(n35985), .Z(n22044) );
  NANDN U22825 ( .A(n22042), .B(n35986), .Z(n22043) );
  NAND U22826 ( .A(n22044), .B(n22043), .Z(n22350) );
  XNOR U22827 ( .A(a[99]), .B(n31123), .Z(n22388) );
  NAND U22828 ( .A(n22388), .B(n29949), .Z(n22047) );
  NAND U22829 ( .A(n29948), .B(n22045), .Z(n22046) );
  NAND U22830 ( .A(n22047), .B(n22046), .Z(n22347) );
  XOR U22831 ( .A(b[55]), .B(n24288), .Z(n22391) );
  NANDN U22832 ( .A(n22391), .B(n38075), .Z(n22050) );
  NANDN U22833 ( .A(n22048), .B(n38073), .Z(n22049) );
  AND U22834 ( .A(n22050), .B(n22049), .Z(n22348) );
  XNOR U22835 ( .A(n22347), .B(n22348), .Z(n22349) );
  XNOR U22836 ( .A(n22350), .B(n22349), .Z(n22191) );
  NANDN U22837 ( .A(n22052), .B(n22051), .Z(n22056) );
  NAND U22838 ( .A(n22054), .B(n22053), .Z(n22055) );
  NAND U22839 ( .A(n22056), .B(n22055), .Z(n22188) );
  NANDN U22840 ( .A(n22058), .B(n22057), .Z(n22062) );
  NAND U22841 ( .A(n22060), .B(n22059), .Z(n22061) );
  NAND U22842 ( .A(n22062), .B(n22061), .Z(n22189) );
  XNOR U22843 ( .A(n22188), .B(n22189), .Z(n22190) );
  XOR U22844 ( .A(n22191), .B(n22190), .Z(n22420) );
  XOR U22845 ( .A(n22421), .B(n22420), .Z(n22413) );
  XNOR U22846 ( .A(a[91]), .B(b[15]), .Z(n22323) );
  OR U22847 ( .A(n22323), .B(n32010), .Z(n22065) );
  NANDN U22848 ( .A(n22063), .B(n32011), .Z(n22064) );
  NAND U22849 ( .A(n22065), .B(n22064), .Z(n22243) );
  XOR U22850 ( .A(b[25]), .B(a[81]), .Z(n22326) );
  NANDN U22851 ( .A(n34219), .B(n22326), .Z(n22068) );
  NAND U22852 ( .A(n34217), .B(n22066), .Z(n22067) );
  NAND U22853 ( .A(n22068), .B(n22067), .Z(n22240) );
  XOR U22854 ( .A(a[89]), .B(b[17]), .Z(n22329) );
  NAND U22855 ( .A(n22329), .B(n32543), .Z(n22071) );
  NANDN U22856 ( .A(n22069), .B(n32541), .Z(n22070) );
  AND U22857 ( .A(n22071), .B(n22070), .Z(n22241) );
  XNOR U22858 ( .A(n22240), .B(n22241), .Z(n22242) );
  XNOR U22859 ( .A(n22243), .B(n22242), .Z(n22262) );
  XOR U22860 ( .A(b[39]), .B(n29372), .Z(n22332) );
  NANDN U22861 ( .A(n22332), .B(n36553), .Z(n22074) );
  NANDN U22862 ( .A(n22072), .B(n36643), .Z(n22073) );
  NAND U22863 ( .A(n22074), .B(n22073), .Z(n22237) );
  XOR U22864 ( .A(b[51]), .B(n25466), .Z(n22335) );
  NANDN U22865 ( .A(n22335), .B(n37803), .Z(n22077) );
  NANDN U22866 ( .A(n22075), .B(n37802), .Z(n22076) );
  NAND U22867 ( .A(n22077), .B(n22076), .Z(n22234) );
  XOR U22868 ( .A(b[53]), .B(n25001), .Z(n22338) );
  NANDN U22869 ( .A(n22338), .B(n37940), .Z(n22080) );
  NANDN U22870 ( .A(n22078), .B(n37941), .Z(n22079) );
  AND U22871 ( .A(n22080), .B(n22079), .Z(n22235) );
  XNOR U22872 ( .A(n22234), .B(n22235), .Z(n22236) );
  XOR U22873 ( .A(n22237), .B(n22236), .Z(n22263) );
  XOR U22874 ( .A(n22262), .B(n22263), .Z(n22265) );
  NANDN U22875 ( .A(n22082), .B(n22081), .Z(n22086) );
  NAND U22876 ( .A(n22084), .B(n22083), .Z(n22085) );
  NAND U22877 ( .A(n22086), .B(n22085), .Z(n22264) );
  XNOR U22878 ( .A(n22265), .B(n22264), .Z(n22314) );
  NANDN U22879 ( .A(n22088), .B(n22087), .Z(n22092) );
  NAND U22880 ( .A(n22090), .B(n22089), .Z(n22091) );
  NAND U22881 ( .A(n22092), .B(n22091), .Z(n22311) );
  NANDN U22882 ( .A(n22094), .B(n22093), .Z(n22098) );
  NAND U22883 ( .A(n22096), .B(n22095), .Z(n22097) );
  AND U22884 ( .A(n22098), .B(n22097), .Z(n22312) );
  XNOR U22885 ( .A(n22311), .B(n22312), .Z(n22313) );
  XNOR U22886 ( .A(n22314), .B(n22313), .Z(n22428) );
  OR U22887 ( .A(n22100), .B(n22099), .Z(n22104) );
  OR U22888 ( .A(n22102), .B(n22101), .Z(n22103) );
  AND U22889 ( .A(n22104), .B(n22103), .Z(n22429) );
  XOR U22890 ( .A(n22428), .B(n22429), .Z(n22431) );
  NANDN U22891 ( .A(n22106), .B(n22105), .Z(n22110) );
  NAND U22892 ( .A(n22108), .B(n22107), .Z(n22109) );
  AND U22893 ( .A(n22110), .B(n22109), .Z(n22430) );
  XNOR U22894 ( .A(n22431), .B(n22430), .Z(n22412) );
  XNOR U22895 ( .A(n22413), .B(n22412), .Z(n22414) );
  XOR U22896 ( .A(n22415), .B(n22414), .Z(n22185) );
  XNOR U22897 ( .A(n22184), .B(n22185), .Z(n22186) );
  NAND U22898 ( .A(n22112), .B(n22111), .Z(n22116) );
  NANDN U22899 ( .A(n22114), .B(n22113), .Z(n22115) );
  AND U22900 ( .A(n22116), .B(n22115), .Z(n22187) );
  XNOR U22901 ( .A(n22186), .B(n22187), .Z(n22436) );
  NANDN U22902 ( .A(n22118), .B(n22117), .Z(n22122) );
  NAND U22903 ( .A(n22120), .B(n22119), .Z(n22121) );
  NAND U22904 ( .A(n22122), .B(n22121), .Z(n22181) );
  XNOR U22905 ( .A(n22178), .B(n22179), .Z(n22180) );
  XNOR U22906 ( .A(n22181), .B(n22180), .Z(n22434) );
  NANDN U22907 ( .A(n22132), .B(n22131), .Z(n22136) );
  NAND U22908 ( .A(n22134), .B(n22133), .Z(n22135) );
  NAND U22909 ( .A(n22136), .B(n22135), .Z(n22435) );
  XOR U22910 ( .A(n22434), .B(n22435), .Z(n22437) );
  XNOR U22911 ( .A(n22436), .B(n22437), .Z(n22443) );
  NANDN U22912 ( .A(n22138), .B(n22137), .Z(n22142) );
  NAND U22913 ( .A(n22140), .B(n22139), .Z(n22141) );
  NAND U22914 ( .A(n22142), .B(n22141), .Z(n22440) );
  NANDN U22915 ( .A(n22144), .B(n22143), .Z(n22148) );
  NANDN U22916 ( .A(n22146), .B(n22145), .Z(n22147) );
  NAND U22917 ( .A(n22148), .B(n22147), .Z(n22441) );
  XNOR U22918 ( .A(n22440), .B(n22441), .Z(n22442) );
  XNOR U22919 ( .A(n22443), .B(n22442), .Z(n22449) );
  OR U22920 ( .A(n22150), .B(n22149), .Z(n22154) );
  NAND U22921 ( .A(n22152), .B(n22151), .Z(n22153) );
  NAND U22922 ( .A(n22154), .B(n22153), .Z(n22447) );
  NANDN U22923 ( .A(n22156), .B(n22155), .Z(n22160) );
  NANDN U22924 ( .A(n22158), .B(n22157), .Z(n22159) );
  AND U22925 ( .A(n22160), .B(n22159), .Z(n22446) );
  XNOR U22926 ( .A(n22447), .B(n22446), .Z(n22448) );
  XOR U22927 ( .A(n22449), .B(n22448), .Z(n22172) );
  NANDN U22928 ( .A(n22162), .B(n22161), .Z(n22166) );
  NAND U22929 ( .A(n22164), .B(n22163), .Z(n22165) );
  NAND U22930 ( .A(n22166), .B(n22165), .Z(n22173) );
  XOR U22931 ( .A(n22172), .B(n22173), .Z(n22174) );
  XNOR U22932 ( .A(n22175), .B(n22174), .Z(n22452) );
  XNOR U22933 ( .A(n22452), .B(sreg[169]), .Z(n22454) );
  NAND U22934 ( .A(n22167), .B(sreg[168]), .Z(n22171) );
  OR U22935 ( .A(n22169), .B(n22168), .Z(n22170) );
  AND U22936 ( .A(n22171), .B(n22170), .Z(n22453) );
  XOR U22937 ( .A(n22454), .B(n22453), .Z(c[169]) );
  OR U22938 ( .A(n22173), .B(n22172), .Z(n22177) );
  NAND U22939 ( .A(n22175), .B(n22174), .Z(n22176) );
  NAND U22940 ( .A(n22177), .B(n22176), .Z(n22460) );
  NANDN U22941 ( .A(n22179), .B(n22178), .Z(n22183) );
  NAND U22942 ( .A(n22181), .B(n22180), .Z(n22182) );
  NAND U22943 ( .A(n22183), .B(n22182), .Z(n22730) );
  XNOR U22944 ( .A(n22730), .B(n22731), .Z(n22732) );
  NANDN U22945 ( .A(n22189), .B(n22188), .Z(n22193) );
  NAND U22946 ( .A(n22191), .B(n22190), .Z(n22192) );
  AND U22947 ( .A(n22193), .B(n22192), .Z(n22472) );
  NANDN U22948 ( .A(n22195), .B(n22194), .Z(n22199) );
  NANDN U22949 ( .A(n22197), .B(n22196), .Z(n22198) );
  NAND U22950 ( .A(n22199), .B(n22198), .Z(n22469) );
  NANDN U22951 ( .A(n22201), .B(n22200), .Z(n22205) );
  NAND U22952 ( .A(n22203), .B(n22202), .Z(n22204) );
  AND U22953 ( .A(n22205), .B(n22204), .Z(n22470) );
  XNOR U22954 ( .A(n22469), .B(n22470), .Z(n22471) );
  XNOR U22955 ( .A(n22472), .B(n22471), .Z(n22706) );
  NANDN U22956 ( .A(n22207), .B(n22206), .Z(n22211) );
  OR U22957 ( .A(n22209), .B(n22208), .Z(n22210) );
  AND U22958 ( .A(n22211), .B(n22210), .Z(n22707) );
  XNOR U22959 ( .A(n22706), .B(n22707), .Z(n22709) );
  XOR U22960 ( .A(b[37]), .B(n30379), .Z(n22513) );
  NANDN U22961 ( .A(n22513), .B(n36311), .Z(n22218) );
  NANDN U22962 ( .A(n22216), .B(n36309), .Z(n22217) );
  NAND U22963 ( .A(n22218), .B(n22217), .Z(n22592) );
  XOR U22964 ( .A(a[102]), .B(n968), .Z(n22516) );
  OR U22965 ( .A(n22516), .B(n29363), .Z(n22221) );
  NANDN U22966 ( .A(n22219), .B(n29864), .Z(n22220) );
  NAND U22967 ( .A(n22221), .B(n22220), .Z(n22589) );
  XOR U22968 ( .A(n36647), .B(n967), .Z(n22519) );
  NAND U22969 ( .A(n22519), .B(n28939), .Z(n22224) );
  NAND U22970 ( .A(n28938), .B(n22222), .Z(n22223) );
  AND U22971 ( .A(n22224), .B(n22223), .Z(n22590) );
  XNOR U22972 ( .A(n22589), .B(n22590), .Z(n22591) );
  XNOR U22973 ( .A(n22592), .B(n22591), .Z(n22498) );
  XOR U22974 ( .A(a[94]), .B(n971), .Z(n22522) );
  OR U22975 ( .A(n22522), .B(n31550), .Z(n22227) );
  NANDN U22976 ( .A(n22225), .B(n31874), .Z(n22226) );
  NAND U22977 ( .A(n22227), .B(n22226), .Z(n22679) );
  NAND U22978 ( .A(n34848), .B(n22228), .Z(n22230) );
  XOR U22979 ( .A(n35375), .B(n32814), .Z(n22525) );
  NAND U22980 ( .A(n34618), .B(n22525), .Z(n22229) );
  NAND U22981 ( .A(n22230), .B(n22229), .Z(n22676) );
  NAND U22982 ( .A(n35188), .B(n22231), .Z(n22233) );
  XOR U22983 ( .A(n35540), .B(n31870), .Z(n22528) );
  NANDN U22984 ( .A(n34968), .B(n22528), .Z(n22232) );
  AND U22985 ( .A(n22233), .B(n22232), .Z(n22677) );
  XNOR U22986 ( .A(n22676), .B(n22677), .Z(n22678) );
  XNOR U22987 ( .A(n22679), .B(n22678), .Z(n22495) );
  NANDN U22988 ( .A(n22235), .B(n22234), .Z(n22239) );
  NAND U22989 ( .A(n22237), .B(n22236), .Z(n22238) );
  NAND U22990 ( .A(n22239), .B(n22238), .Z(n22496) );
  XNOR U22991 ( .A(n22495), .B(n22496), .Z(n22497) );
  XOR U22992 ( .A(n22498), .B(n22497), .Z(n22501) );
  NANDN U22993 ( .A(n22241), .B(n22240), .Z(n22245) );
  NAND U22994 ( .A(n22243), .B(n22242), .Z(n22244) );
  NAND U22995 ( .A(n22245), .B(n22244), .Z(n22634) );
  ANDN U22996 ( .B(b[63]), .A(n22246), .Z(n22649) );
  NANDN U22997 ( .A(n22247), .B(n38369), .Z(n22249) );
  XOR U22998 ( .A(b[61]), .B(n22964), .Z(n22543) );
  OR U22999 ( .A(n22543), .B(n38371), .Z(n22248) );
  NAND U23000 ( .A(n22249), .B(n22248), .Z(n22647) );
  NANDN U23001 ( .A(n22250), .B(n35311), .Z(n22252) );
  XOR U23002 ( .A(b[31]), .B(n31363), .Z(n22546) );
  NANDN U23003 ( .A(n22546), .B(n35313), .Z(n22251) );
  AND U23004 ( .A(n22252), .B(n22251), .Z(n22646) );
  XNOR U23005 ( .A(n22647), .B(n22646), .Z(n22648) );
  XOR U23006 ( .A(n22649), .B(n22648), .Z(n22631) );
  NAND U23007 ( .A(n33283), .B(n22253), .Z(n22255) );
  XOR U23008 ( .A(n34048), .B(n33020), .Z(n22549) );
  NANDN U23009 ( .A(n33021), .B(n22549), .Z(n22254) );
  NAND U23010 ( .A(n22255), .B(n22254), .Z(n22561) );
  XNOR U23011 ( .A(b[21]), .B(a[86]), .Z(n22552) );
  OR U23012 ( .A(n22552), .B(n33634), .Z(n22258) );
  NAND U23013 ( .A(n22256), .B(n33464), .Z(n22257) );
  NAND U23014 ( .A(n22258), .B(n22257), .Z(n22558) );
  NAND U23015 ( .A(n34044), .B(n22259), .Z(n22261) );
  XOR U23016 ( .A(n34510), .B(n33185), .Z(n22555) );
  NANDN U23017 ( .A(n33867), .B(n22555), .Z(n22260) );
  AND U23018 ( .A(n22261), .B(n22260), .Z(n22559) );
  XNOR U23019 ( .A(n22558), .B(n22559), .Z(n22560) );
  XNOR U23020 ( .A(n22561), .B(n22560), .Z(n22632) );
  XNOR U23021 ( .A(n22631), .B(n22632), .Z(n22633) );
  XNOR U23022 ( .A(n22634), .B(n22633), .Z(n22502) );
  XOR U23023 ( .A(n22501), .B(n22502), .Z(n22503) );
  XOR U23024 ( .A(n22504), .B(n22503), .Z(n22603) );
  NANDN U23025 ( .A(n22263), .B(n22262), .Z(n22267) );
  OR U23026 ( .A(n22265), .B(n22264), .Z(n22266) );
  NAND U23027 ( .A(n22267), .B(n22266), .Z(n22602) );
  NANDN U23028 ( .A(n22269), .B(n22268), .Z(n22273) );
  NAND U23029 ( .A(n22271), .B(n22270), .Z(n22272) );
  NAND U23030 ( .A(n22273), .B(n22272), .Z(n22492) );
  XNOR U23031 ( .A(b[41]), .B(a[66]), .Z(n22564) );
  OR U23032 ( .A(n22564), .B(n36905), .Z(n22276) );
  NANDN U23033 ( .A(n22274), .B(n36807), .Z(n22275) );
  NAND U23034 ( .A(n22276), .B(n22275), .Z(n22586) );
  XOR U23035 ( .A(b[57]), .B(n24671), .Z(n22567) );
  OR U23036 ( .A(n22567), .B(n965), .Z(n22279) );
  NANDN U23037 ( .A(n22277), .B(n38194), .Z(n22278) );
  NAND U23038 ( .A(n22279), .B(n22278), .Z(n22583) );
  NAND U23039 ( .A(n38326), .B(n22280), .Z(n22282) );
  XOR U23040 ( .A(n38400), .B(n23447), .Z(n22570) );
  NANDN U23041 ( .A(n38273), .B(n22570), .Z(n22281) );
  AND U23042 ( .A(n22282), .B(n22281), .Z(n22584) );
  XNOR U23043 ( .A(n22583), .B(n22584), .Z(n22585) );
  XOR U23044 ( .A(n22586), .B(n22585), .Z(n22694) );
  XOR U23045 ( .A(b[33]), .B(n31372), .Z(n22573) );
  NANDN U23046 ( .A(n22573), .B(n35620), .Z(n22285) );
  NANDN U23047 ( .A(n22283), .B(n35621), .Z(n22284) );
  NAND U23048 ( .A(n22285), .B(n22284), .Z(n22691) );
  NANDN U23049 ( .A(n966), .B(a[106]), .Z(n22286) );
  XOR U23050 ( .A(n29232), .B(n22286), .Z(n22288) );
  NANDN U23051 ( .A(b[0]), .B(a[105]), .Z(n22287) );
  AND U23052 ( .A(n22288), .B(n22287), .Z(n22688) );
  XOR U23053 ( .A(b[63]), .B(n22289), .Z(n22580) );
  NANDN U23054 ( .A(n22580), .B(n38422), .Z(n22292) );
  NANDN U23055 ( .A(n22290), .B(n38423), .Z(n22291) );
  AND U23056 ( .A(n22292), .B(n22291), .Z(n22689) );
  XNOR U23057 ( .A(n22688), .B(n22689), .Z(n22690) );
  XOR U23058 ( .A(n22691), .B(n22690), .Z(n22695) );
  XNOR U23059 ( .A(n22694), .B(n22695), .Z(n22697) );
  NANDN U23060 ( .A(n22294), .B(n22293), .Z(n22298) );
  NAND U23061 ( .A(n22296), .B(n22295), .Z(n22297) );
  NAND U23062 ( .A(n22298), .B(n22297), .Z(n22696) );
  XOR U23063 ( .A(n22697), .B(n22696), .Z(n22489) );
  NANDN U23064 ( .A(n22300), .B(n22299), .Z(n22304) );
  NAND U23065 ( .A(n22302), .B(n22301), .Z(n22303) );
  AND U23066 ( .A(n22304), .B(n22303), .Z(n22490) );
  XOR U23067 ( .A(n22489), .B(n22490), .Z(n22491) );
  XNOR U23068 ( .A(n22492), .B(n22491), .Z(n22601) );
  XNOR U23069 ( .A(n22602), .B(n22601), .Z(n22604) );
  XNOR U23070 ( .A(n22603), .B(n22604), .Z(n22708) );
  XOR U23071 ( .A(n22709), .B(n22708), .Z(n22718) );
  NAND U23072 ( .A(n22306), .B(n22305), .Z(n22310) );
  NANDN U23073 ( .A(n22308), .B(n22307), .Z(n22309) );
  NAND U23074 ( .A(n22310), .B(n22309), .Z(n22480) );
  NANDN U23075 ( .A(n22312), .B(n22311), .Z(n22316) );
  NAND U23076 ( .A(n22314), .B(n22313), .Z(n22315) );
  NAND U23077 ( .A(n22316), .B(n22315), .Z(n22476) );
  NANDN U23078 ( .A(n22318), .B(n22317), .Z(n22322) );
  OR U23079 ( .A(n22320), .B(n22319), .Z(n22321) );
  NAND U23080 ( .A(n22322), .B(n22321), .Z(n22474) );
  XOR U23081 ( .A(a[92]), .B(n972), .Z(n22658) );
  OR U23082 ( .A(n22658), .B(n32010), .Z(n22325) );
  NANDN U23083 ( .A(n22323), .B(n32011), .Z(n22324) );
  NAND U23084 ( .A(n22325), .B(n22324), .Z(n22540) );
  XNOR U23085 ( .A(b[25]), .B(n32815), .Z(n22661) );
  NANDN U23086 ( .A(n34219), .B(n22661), .Z(n22328) );
  NAND U23087 ( .A(n34217), .B(n22326), .Z(n22327) );
  NAND U23088 ( .A(n22328), .B(n22327), .Z(n22537) );
  XNOR U23089 ( .A(a[90]), .B(b[17]), .Z(n22664) );
  NANDN U23090 ( .A(n22664), .B(n32543), .Z(n22331) );
  NAND U23091 ( .A(n22329), .B(n32541), .Z(n22330) );
  AND U23092 ( .A(n22331), .B(n22330), .Z(n22538) );
  XNOR U23093 ( .A(n22537), .B(n22538), .Z(n22539) );
  XOR U23094 ( .A(n22540), .B(n22539), .Z(n22595) );
  XOR U23095 ( .A(b[39]), .B(n29868), .Z(n22667) );
  NANDN U23096 ( .A(n22667), .B(n36553), .Z(n22334) );
  NANDN U23097 ( .A(n22332), .B(n36643), .Z(n22333) );
  NAND U23098 ( .A(n22334), .B(n22333), .Z(n22534) );
  XOR U23099 ( .A(b[51]), .B(n25860), .Z(n22670) );
  NANDN U23100 ( .A(n22670), .B(n37803), .Z(n22337) );
  NANDN U23101 ( .A(n22335), .B(n37802), .Z(n22336) );
  NAND U23102 ( .A(n22337), .B(n22336), .Z(n22531) );
  XOR U23103 ( .A(b[53]), .B(n25177), .Z(n22673) );
  NANDN U23104 ( .A(n22673), .B(n37940), .Z(n22340) );
  NANDN U23105 ( .A(n22338), .B(n37941), .Z(n22339) );
  AND U23106 ( .A(n22340), .B(n22339), .Z(n22532) );
  XNOR U23107 ( .A(n22531), .B(n22532), .Z(n22533) );
  XOR U23108 ( .A(n22534), .B(n22533), .Z(n22596) );
  XNOR U23109 ( .A(n22595), .B(n22596), .Z(n22598) );
  NANDN U23110 ( .A(n22342), .B(n22341), .Z(n22346) );
  NAND U23111 ( .A(n22344), .B(n22343), .Z(n22345) );
  NAND U23112 ( .A(n22346), .B(n22345), .Z(n22597) );
  XNOR U23113 ( .A(n22598), .B(n22597), .Z(n22703) );
  NANDN U23114 ( .A(n22348), .B(n22347), .Z(n22352) );
  NAND U23115 ( .A(n22350), .B(n22349), .Z(n22351) );
  NAND U23116 ( .A(n22352), .B(n22351), .Z(n22700) );
  XNOR U23117 ( .A(n22700), .B(n22701), .Z(n22702) );
  XOR U23118 ( .A(n22703), .B(n22702), .Z(n22473) );
  XNOR U23119 ( .A(n22474), .B(n22473), .Z(n22475) );
  XNOR U23120 ( .A(n22476), .B(n22475), .Z(n22478) );
  XOR U23121 ( .A(a[96]), .B(n970), .Z(n22607) );
  OR U23122 ( .A(n22607), .B(n31369), .Z(n22359) );
  NANDN U23123 ( .A(n22357), .B(n31119), .Z(n22358) );
  NAND U23124 ( .A(n22359), .B(n22358), .Z(n22628) );
  XNOR U23125 ( .A(b[43]), .B(a[64]), .Z(n22610) );
  NANDN U23126 ( .A(n22610), .B(n37068), .Z(n22362) );
  NANDN U23127 ( .A(n22360), .B(n37069), .Z(n22361) );
  NAND U23128 ( .A(n22362), .B(n22361), .Z(n22625) );
  XOR U23129 ( .A(b[45]), .B(a[62]), .Z(n22613) );
  NAND U23130 ( .A(n22613), .B(n37261), .Z(n22365) );
  NANDN U23131 ( .A(n22363), .B(n37262), .Z(n22364) );
  AND U23132 ( .A(n22365), .B(n22364), .Z(n22626) );
  XNOR U23133 ( .A(n22625), .B(n22626), .Z(n22627) );
  XNOR U23134 ( .A(n22628), .B(n22627), .Z(n22507) );
  NAND U23135 ( .A(n37652), .B(n22366), .Z(n22368) );
  XOR U23136 ( .A(b[49]), .B(n26347), .Z(n22616) );
  OR U23137 ( .A(n22616), .B(n37756), .Z(n22367) );
  NAND U23138 ( .A(n22368), .B(n22367), .Z(n22654) );
  NANDN U23139 ( .A(n22369), .B(n37469), .Z(n22371) );
  XNOR U23140 ( .A(n978), .B(a[60]), .Z(n22619) );
  NAND U23141 ( .A(n22619), .B(n37471), .Z(n22370) );
  AND U23142 ( .A(n22371), .B(n22370), .Z(n22653) );
  NAND U23143 ( .A(n30846), .B(n22372), .Z(n22374) );
  XNOR U23144 ( .A(n35783), .B(b[9]), .Z(n22622) );
  NAND U23145 ( .A(n30509), .B(n22622), .Z(n22373) );
  NAND U23146 ( .A(n22374), .B(n22373), .Z(n22652) );
  XNOR U23147 ( .A(n22653), .B(n22652), .Z(n22655) );
  XOR U23148 ( .A(n22654), .B(n22655), .Z(n22508) );
  XNOR U23149 ( .A(n22507), .B(n22508), .Z(n22509) );
  NANDN U23150 ( .A(n22376), .B(n22375), .Z(n22380) );
  NAND U23151 ( .A(n22378), .B(n22377), .Z(n22379) );
  AND U23152 ( .A(n22380), .B(n22379), .Z(n22510) );
  XNOR U23153 ( .A(n22509), .B(n22510), .Z(n22464) );
  XNOR U23154 ( .A(n22464), .B(n22463), .Z(n22465) );
  XNOR U23155 ( .A(b[35]), .B(a[72]), .Z(n22637) );
  NANDN U23156 ( .A(n22637), .B(n35985), .Z(n22387) );
  NANDN U23157 ( .A(n22385), .B(n35986), .Z(n22386) );
  NAND U23158 ( .A(n22387), .B(n22386), .Z(n22685) );
  XOR U23159 ( .A(n36100), .B(n31123), .Z(n22640) );
  NAND U23160 ( .A(n22640), .B(n29949), .Z(n22390) );
  NAND U23161 ( .A(n29948), .B(n22388), .Z(n22389) );
  NAND U23162 ( .A(n22390), .B(n22389), .Z(n22682) );
  XOR U23163 ( .A(b[55]), .B(n25134), .Z(n22643) );
  NANDN U23164 ( .A(n22643), .B(n38075), .Z(n22393) );
  NANDN U23165 ( .A(n22391), .B(n38073), .Z(n22392) );
  AND U23166 ( .A(n22393), .B(n22392), .Z(n22683) );
  XNOR U23167 ( .A(n22682), .B(n22683), .Z(n22684) );
  XNOR U23168 ( .A(n22685), .B(n22684), .Z(n22486) );
  NANDN U23169 ( .A(n22395), .B(n22394), .Z(n22399) );
  NAND U23170 ( .A(n22397), .B(n22396), .Z(n22398) );
  NAND U23171 ( .A(n22399), .B(n22398), .Z(n22483) );
  NANDN U23172 ( .A(n22401), .B(n22400), .Z(n22405) );
  NAND U23173 ( .A(n22403), .B(n22402), .Z(n22404) );
  NAND U23174 ( .A(n22405), .B(n22404), .Z(n22484) );
  XNOR U23175 ( .A(n22483), .B(n22484), .Z(n22485) );
  XOR U23176 ( .A(n22486), .B(n22485), .Z(n22466) );
  XOR U23177 ( .A(n22465), .B(n22466), .Z(n22477) );
  XOR U23178 ( .A(n22478), .B(n22477), .Z(n22479) );
  XOR U23179 ( .A(n22480), .B(n22479), .Z(n22719) );
  XNOR U23180 ( .A(n22718), .B(n22719), .Z(n22720) );
  OR U23181 ( .A(n22407), .B(n22406), .Z(n22411) );
  NAND U23182 ( .A(n22409), .B(n22408), .Z(n22410) );
  NAND U23183 ( .A(n22411), .B(n22410), .Z(n22721) );
  XOR U23184 ( .A(n22720), .B(n22721), .Z(n22727) );
  NANDN U23185 ( .A(n22413), .B(n22412), .Z(n22417) );
  NAND U23186 ( .A(n22415), .B(n22414), .Z(n22416) );
  AND U23187 ( .A(n22417), .B(n22416), .Z(n22724) );
  NAND U23188 ( .A(n22419), .B(n22418), .Z(n22423) );
  NANDN U23189 ( .A(n22421), .B(n22420), .Z(n22422) );
  NAND U23190 ( .A(n22423), .B(n22422), .Z(n22715) );
  NANDN U23191 ( .A(n22429), .B(n22428), .Z(n22433) );
  NANDN U23192 ( .A(n22431), .B(n22430), .Z(n22432) );
  AND U23193 ( .A(n22433), .B(n22432), .Z(n22713) );
  XNOR U23194 ( .A(n22712), .B(n22713), .Z(n22714) );
  XNOR U23195 ( .A(n22715), .B(n22714), .Z(n22725) );
  XNOR U23196 ( .A(n22727), .B(n22726), .Z(n22733) );
  XOR U23197 ( .A(n22732), .B(n22733), .Z(n22736) );
  NANDN U23198 ( .A(n22435), .B(n22434), .Z(n22439) );
  OR U23199 ( .A(n22437), .B(n22436), .Z(n22438) );
  AND U23200 ( .A(n22439), .B(n22438), .Z(n22737) );
  XNOR U23201 ( .A(n22736), .B(n22737), .Z(n22738) );
  NANDN U23202 ( .A(n22441), .B(n22440), .Z(n22445) );
  NAND U23203 ( .A(n22443), .B(n22442), .Z(n22444) );
  NAND U23204 ( .A(n22445), .B(n22444), .Z(n22739) );
  XOR U23205 ( .A(n22738), .B(n22739), .Z(n22457) );
  NANDN U23206 ( .A(n22447), .B(n22446), .Z(n22451) );
  NAND U23207 ( .A(n22449), .B(n22448), .Z(n22450) );
  NAND U23208 ( .A(n22451), .B(n22450), .Z(n22458) );
  XNOR U23209 ( .A(n22457), .B(n22458), .Z(n22459) );
  XNOR U23210 ( .A(n22460), .B(n22459), .Z(n22742) );
  XNOR U23211 ( .A(n22742), .B(sreg[170]), .Z(n22744) );
  NAND U23212 ( .A(n22452), .B(sreg[169]), .Z(n22456) );
  OR U23213 ( .A(n22454), .B(n22453), .Z(n22455) );
  AND U23214 ( .A(n22456), .B(n22455), .Z(n22743) );
  XOR U23215 ( .A(n22744), .B(n22743), .Z(c[170]) );
  NANDN U23216 ( .A(n22458), .B(n22457), .Z(n22462) );
  NAND U23217 ( .A(n22460), .B(n22459), .Z(n22461) );
  NAND U23218 ( .A(n22462), .B(n22461), .Z(n22750) );
  NANDN U23219 ( .A(n22464), .B(n22463), .Z(n22468) );
  NAND U23220 ( .A(n22466), .B(n22465), .Z(n22467) );
  NAND U23221 ( .A(n22468), .B(n22467), .Z(n23005) );
  XNOR U23222 ( .A(n23002), .B(n23003), .Z(n23004) );
  XNOR U23223 ( .A(n23005), .B(n23004), .Z(n23014) );
  NAND U23224 ( .A(n22478), .B(n22477), .Z(n22482) );
  NAND U23225 ( .A(n22480), .B(n22479), .Z(n22481) );
  NAND U23226 ( .A(n22482), .B(n22481), .Z(n23015) );
  XNOR U23227 ( .A(n23014), .B(n23015), .Z(n23016) );
  NANDN U23228 ( .A(n22484), .B(n22483), .Z(n22488) );
  NAND U23229 ( .A(n22486), .B(n22485), .Z(n22487) );
  NAND U23230 ( .A(n22488), .B(n22487), .Z(n22989) );
  NAND U23231 ( .A(n22490), .B(n22489), .Z(n22494) );
  NANDN U23232 ( .A(n22492), .B(n22491), .Z(n22493) );
  NAND U23233 ( .A(n22494), .B(n22493), .Z(n22986) );
  NANDN U23234 ( .A(n22496), .B(n22495), .Z(n22500) );
  NAND U23235 ( .A(n22498), .B(n22497), .Z(n22499) );
  AND U23236 ( .A(n22500), .B(n22499), .Z(n22987) );
  XNOR U23237 ( .A(n22986), .B(n22987), .Z(n22988) );
  XNOR U23238 ( .A(n22989), .B(n22988), .Z(n22754) );
  OR U23239 ( .A(n22502), .B(n22501), .Z(n22506) );
  NANDN U23240 ( .A(n22504), .B(n22503), .Z(n22505) );
  AND U23241 ( .A(n22506), .B(n22505), .Z(n22753) );
  XNOR U23242 ( .A(n22754), .B(n22753), .Z(n22755) );
  NANDN U23243 ( .A(n22508), .B(n22507), .Z(n22512) );
  NAND U23244 ( .A(n22510), .B(n22509), .Z(n22511) );
  NAND U23245 ( .A(n22512), .B(n22511), .Z(n22864) );
  XOR U23246 ( .A(b[37]), .B(n30543), .Z(n22892) );
  NANDN U23247 ( .A(n22892), .B(n36311), .Z(n22515) );
  NANDN U23248 ( .A(n22513), .B(n36309), .Z(n22514) );
  NAND U23249 ( .A(n22515), .B(n22514), .Z(n22946) );
  XNOR U23250 ( .A(a[103]), .B(b[5]), .Z(n22895) );
  OR U23251 ( .A(n22895), .B(n29363), .Z(n22518) );
  NANDN U23252 ( .A(n22516), .B(n29864), .Z(n22517) );
  NAND U23253 ( .A(n22518), .B(n22517), .Z(n22943) );
  XNOR U23254 ( .A(a[105]), .B(n967), .Z(n22898) );
  NAND U23255 ( .A(n22898), .B(n28939), .Z(n22521) );
  NAND U23256 ( .A(n28938), .B(n22519), .Z(n22520) );
  AND U23257 ( .A(n22521), .B(n22520), .Z(n22944) );
  XNOR U23258 ( .A(n22943), .B(n22944), .Z(n22945) );
  XOR U23259 ( .A(n22946), .B(n22945), .Z(n22871) );
  XOR U23260 ( .A(a[95]), .B(n971), .Z(n22901) );
  OR U23261 ( .A(n22901), .B(n31550), .Z(n22524) );
  NANDN U23262 ( .A(n22522), .B(n31874), .Z(n22523) );
  NAND U23263 ( .A(n22524), .B(n22523), .Z(n22835) );
  NAND U23264 ( .A(n34848), .B(n22525), .Z(n22527) );
  XNOR U23265 ( .A(n35375), .B(a[81]), .Z(n22904) );
  NAND U23266 ( .A(n34618), .B(n22904), .Z(n22526) );
  NAND U23267 ( .A(n22527), .B(n22526), .Z(n22832) );
  NAND U23268 ( .A(n35188), .B(n22528), .Z(n22530) );
  XNOR U23269 ( .A(n35540), .B(a[79]), .Z(n22907) );
  NANDN U23270 ( .A(n34968), .B(n22907), .Z(n22529) );
  AND U23271 ( .A(n22530), .B(n22529), .Z(n22833) );
  XNOR U23272 ( .A(n22832), .B(n22833), .Z(n22834) );
  XOR U23273 ( .A(n22835), .B(n22834), .Z(n22869) );
  NANDN U23274 ( .A(n22532), .B(n22531), .Z(n22536) );
  NAND U23275 ( .A(n22534), .B(n22533), .Z(n22535) );
  AND U23276 ( .A(n22536), .B(n22535), .Z(n22868) );
  XOR U23277 ( .A(n22869), .B(n22868), .Z(n22870) );
  XOR U23278 ( .A(n22871), .B(n22870), .Z(n22863) );
  NANDN U23279 ( .A(n22538), .B(n22537), .Z(n22542) );
  NAND U23280 ( .A(n22540), .B(n22539), .Z(n22541) );
  NAND U23281 ( .A(n22542), .B(n22541), .Z(n22791) );
  NAND U23282 ( .A(a[43]), .B(b[63]), .Z(n22805) );
  NANDN U23283 ( .A(n22543), .B(n38369), .Z(n22545) );
  XOR U23284 ( .A(b[61]), .B(n23149), .Z(n22922) );
  OR U23285 ( .A(n22922), .B(n38371), .Z(n22544) );
  NAND U23286 ( .A(n22545), .B(n22544), .Z(n22803) );
  NANDN U23287 ( .A(n22546), .B(n35311), .Z(n22548) );
  XNOR U23288 ( .A(b[31]), .B(a[77]), .Z(n22925) );
  NANDN U23289 ( .A(n22925), .B(n35313), .Z(n22547) );
  AND U23290 ( .A(n22548), .B(n22547), .Z(n22802) );
  XNOR U23291 ( .A(n22803), .B(n22802), .Z(n22804) );
  XOR U23292 ( .A(n22805), .B(n22804), .Z(n22789) );
  NAND U23293 ( .A(n33283), .B(n22549), .Z(n22551) );
  XNOR U23294 ( .A(a[89]), .B(n33020), .Z(n22928) );
  NANDN U23295 ( .A(n33021), .B(n22928), .Z(n22550) );
  NAND U23296 ( .A(n22551), .B(n22550), .Z(n22971) );
  XOR U23297 ( .A(b[21]), .B(a[87]), .Z(n22931) );
  NANDN U23298 ( .A(n33634), .B(n22931), .Z(n22554) );
  NANDN U23299 ( .A(n22552), .B(n33464), .Z(n22553) );
  NAND U23300 ( .A(n22554), .B(n22553), .Z(n22968) );
  NAND U23301 ( .A(n34044), .B(n22555), .Z(n22557) );
  XNOR U23302 ( .A(n34510), .B(a[85]), .Z(n22934) );
  NANDN U23303 ( .A(n33867), .B(n22934), .Z(n22556) );
  AND U23304 ( .A(n22557), .B(n22556), .Z(n22969) );
  XNOR U23305 ( .A(n22968), .B(n22969), .Z(n22970) );
  XNOR U23306 ( .A(n22971), .B(n22970), .Z(n22790) );
  XNOR U23307 ( .A(n22789), .B(n22790), .Z(n22792) );
  XNOR U23308 ( .A(n22791), .B(n22792), .Z(n22862) );
  XOR U23309 ( .A(n22863), .B(n22862), .Z(n22865) );
  XNOR U23310 ( .A(n22864), .B(n22865), .Z(n22762) );
  NANDN U23311 ( .A(n22559), .B(n22558), .Z(n22563) );
  NAND U23312 ( .A(n22561), .B(n22560), .Z(n22562) );
  NAND U23313 ( .A(n22563), .B(n22562), .Z(n22853) );
  XNOR U23314 ( .A(b[41]), .B(a[67]), .Z(n22949) );
  OR U23315 ( .A(n22949), .B(n36905), .Z(n22566) );
  NANDN U23316 ( .A(n22564), .B(n36807), .Z(n22565) );
  NAND U23317 ( .A(n22566), .B(n22565), .Z(n22977) );
  XOR U23318 ( .A(b[57]), .B(n24288), .Z(n22952) );
  OR U23319 ( .A(n22952), .B(n965), .Z(n22569) );
  NANDN U23320 ( .A(n22567), .B(n38194), .Z(n22568) );
  NAND U23321 ( .A(n22569), .B(n22568), .Z(n22974) );
  NAND U23322 ( .A(n38326), .B(n22570), .Z(n22572) );
  XOR U23323 ( .A(n38400), .B(n23852), .Z(n22955) );
  NANDN U23324 ( .A(n38273), .B(n22955), .Z(n22571) );
  AND U23325 ( .A(n22572), .B(n22571), .Z(n22975) );
  XNOR U23326 ( .A(n22974), .B(n22975), .Z(n22976) );
  XOR U23327 ( .A(n22977), .B(n22976), .Z(n22850) );
  XNOR U23328 ( .A(b[33]), .B(a[75]), .Z(n22958) );
  NANDN U23329 ( .A(n22958), .B(n35620), .Z(n22575) );
  NANDN U23330 ( .A(n22573), .B(n35621), .Z(n22574) );
  NAND U23331 ( .A(n22575), .B(n22574), .Z(n22847) );
  NANDN U23332 ( .A(n966), .B(a[107]), .Z(n22576) );
  XOR U23333 ( .A(n29232), .B(n22576), .Z(n22578) );
  IV U23334 ( .A(a[106]), .Z(n36909) );
  NANDN U23335 ( .A(n36909), .B(n966), .Z(n22577) );
  AND U23336 ( .A(n22578), .B(n22577), .Z(n22844) );
  XOR U23337 ( .A(b[63]), .B(n22579), .Z(n22965) );
  NANDN U23338 ( .A(n22965), .B(n38422), .Z(n22582) );
  NANDN U23339 ( .A(n22580), .B(n38423), .Z(n22581) );
  AND U23340 ( .A(n22582), .B(n22581), .Z(n22845) );
  XNOR U23341 ( .A(n22844), .B(n22845), .Z(n22846) );
  XOR U23342 ( .A(n22847), .B(n22846), .Z(n22851) );
  XNOR U23343 ( .A(n22850), .B(n22851), .Z(n22852) );
  XNOR U23344 ( .A(n22853), .B(n22852), .Z(n22883) );
  NANDN U23345 ( .A(n22584), .B(n22583), .Z(n22588) );
  NAND U23346 ( .A(n22586), .B(n22585), .Z(n22587) );
  NAND U23347 ( .A(n22588), .B(n22587), .Z(n22880) );
  NANDN U23348 ( .A(n22590), .B(n22589), .Z(n22594) );
  NAND U23349 ( .A(n22592), .B(n22591), .Z(n22593) );
  AND U23350 ( .A(n22594), .B(n22593), .Z(n22881) );
  XNOR U23351 ( .A(n22880), .B(n22881), .Z(n22882) );
  XOR U23352 ( .A(n22883), .B(n22882), .Z(n22760) );
  OR U23353 ( .A(n22596), .B(n22595), .Z(n22600) );
  OR U23354 ( .A(n22598), .B(n22597), .Z(n22599) );
  AND U23355 ( .A(n22600), .B(n22599), .Z(n22759) );
  XOR U23356 ( .A(n22760), .B(n22759), .Z(n22761) );
  XNOR U23357 ( .A(n22762), .B(n22761), .Z(n22756) );
  XOR U23358 ( .A(n22755), .B(n22756), .Z(n23009) );
  NAND U23359 ( .A(n22602), .B(n22601), .Z(n22606) );
  NANDN U23360 ( .A(n22604), .B(n22603), .Z(n22605) );
  NAND U23361 ( .A(n22606), .B(n22605), .Z(n23000) );
  XNOR U23362 ( .A(a[97]), .B(b[11]), .Z(n22765) );
  OR U23363 ( .A(n22765), .B(n31369), .Z(n22609) );
  NANDN U23364 ( .A(n22607), .B(n31119), .Z(n22608) );
  NAND U23365 ( .A(n22609), .B(n22608), .Z(n22786) );
  XOR U23366 ( .A(b[43]), .B(n28403), .Z(n22768) );
  NANDN U23367 ( .A(n22768), .B(n37068), .Z(n22612) );
  NANDN U23368 ( .A(n22610), .B(n37069), .Z(n22611) );
  NAND U23369 ( .A(n22612), .B(n22611), .Z(n22783) );
  XOR U23370 ( .A(b[45]), .B(a[63]), .Z(n22771) );
  NAND U23371 ( .A(n22771), .B(n37261), .Z(n22615) );
  NAND U23372 ( .A(n22613), .B(n37262), .Z(n22614) );
  AND U23373 ( .A(n22615), .B(n22614), .Z(n22784) );
  XNOR U23374 ( .A(n22783), .B(n22784), .Z(n22785) );
  XNOR U23375 ( .A(n22786), .B(n22785), .Z(n22886) );
  XNOR U23376 ( .A(b[49]), .B(a[59]), .Z(n22774) );
  OR U23377 ( .A(n22774), .B(n37756), .Z(n22618) );
  NANDN U23378 ( .A(n22616), .B(n37652), .Z(n22617) );
  NAND U23379 ( .A(n22618), .B(n22617), .Z(n22811) );
  NAND U23380 ( .A(n22619), .B(n37469), .Z(n22621) );
  XOR U23381 ( .A(n978), .B(n27773), .Z(n22777) );
  NAND U23382 ( .A(n22777), .B(n37471), .Z(n22620) );
  NAND U23383 ( .A(n22621), .B(n22620), .Z(n22808) );
  XNOR U23384 ( .A(a[99]), .B(b[9]), .Z(n22780) );
  NANDN U23385 ( .A(n22780), .B(n30509), .Z(n22624) );
  NAND U23386 ( .A(n22622), .B(n30846), .Z(n22623) );
  AND U23387 ( .A(n22624), .B(n22623), .Z(n22809) );
  XNOR U23388 ( .A(n22808), .B(n22809), .Z(n22810) );
  XOR U23389 ( .A(n22811), .B(n22810), .Z(n22887) );
  XNOR U23390 ( .A(n22886), .B(n22887), .Z(n22888) );
  NANDN U23391 ( .A(n22626), .B(n22625), .Z(n22630) );
  NAND U23392 ( .A(n22628), .B(n22627), .Z(n22629) );
  AND U23393 ( .A(n22630), .B(n22629), .Z(n22889) );
  XNOR U23394 ( .A(n22888), .B(n22889), .Z(n22981) );
  NANDN U23395 ( .A(n22632), .B(n22631), .Z(n22636) );
  NAND U23396 ( .A(n22634), .B(n22633), .Z(n22635) );
  AND U23397 ( .A(n22636), .B(n22635), .Z(n22980) );
  XNOR U23398 ( .A(n22981), .B(n22980), .Z(n22982) );
  XOR U23399 ( .A(b[35]), .B(a[73]), .Z(n22793) );
  NAND U23400 ( .A(n35985), .B(n22793), .Z(n22639) );
  NANDN U23401 ( .A(n22637), .B(n35986), .Z(n22638) );
  NAND U23402 ( .A(n22639), .B(n22638), .Z(n22841) );
  XNOR U23403 ( .A(a[101]), .B(n31123), .Z(n22796) );
  NAND U23404 ( .A(n22796), .B(n29949), .Z(n22642) );
  NAND U23405 ( .A(n29948), .B(n22640), .Z(n22641) );
  NAND U23406 ( .A(n22642), .B(n22641), .Z(n22838) );
  XOR U23407 ( .A(b[55]), .B(n25001), .Z(n22799) );
  NANDN U23408 ( .A(n22799), .B(n38075), .Z(n22645) );
  NANDN U23409 ( .A(n22643), .B(n38073), .Z(n22644) );
  AND U23410 ( .A(n22645), .B(n22644), .Z(n22839) );
  XNOR U23411 ( .A(n22838), .B(n22839), .Z(n22840) );
  XNOR U23412 ( .A(n22841), .B(n22840), .Z(n22877) );
  NANDN U23413 ( .A(n22647), .B(n22646), .Z(n22651) );
  NANDN U23414 ( .A(n22649), .B(n22648), .Z(n22650) );
  NAND U23415 ( .A(n22651), .B(n22650), .Z(n22874) );
  NANDN U23416 ( .A(n22653), .B(n22652), .Z(n22657) );
  NAND U23417 ( .A(n22655), .B(n22654), .Z(n22656) );
  NAND U23418 ( .A(n22657), .B(n22656), .Z(n22875) );
  XNOR U23419 ( .A(n22874), .B(n22875), .Z(n22876) );
  XOR U23420 ( .A(n22877), .B(n22876), .Z(n22983) );
  XOR U23421 ( .A(n22982), .B(n22983), .Z(n22998) );
  XOR U23422 ( .A(a[93]), .B(n972), .Z(n22823) );
  OR U23423 ( .A(n22823), .B(n32010), .Z(n22660) );
  NANDN U23424 ( .A(n22658), .B(n32011), .Z(n22659) );
  NAND U23425 ( .A(n22660), .B(n22659), .Z(n22919) );
  XOR U23426 ( .A(b[25]), .B(a[83]), .Z(n22826) );
  NANDN U23427 ( .A(n34219), .B(n22826), .Z(n22663) );
  NAND U23428 ( .A(n34217), .B(n22661), .Z(n22662) );
  NAND U23429 ( .A(n22663), .B(n22662), .Z(n22916) );
  XOR U23430 ( .A(a[91]), .B(b[17]), .Z(n22829) );
  NAND U23431 ( .A(n22829), .B(n32543), .Z(n22666) );
  NANDN U23432 ( .A(n22664), .B(n32541), .Z(n22665) );
  AND U23433 ( .A(n22666), .B(n22665), .Z(n22917) );
  XNOR U23434 ( .A(n22916), .B(n22917), .Z(n22918) );
  XNOR U23435 ( .A(n22919), .B(n22918), .Z(n22937) );
  XNOR U23436 ( .A(b[39]), .B(a[69]), .Z(n22814) );
  NANDN U23437 ( .A(n22814), .B(n36553), .Z(n22669) );
  NANDN U23438 ( .A(n22667), .B(n36643), .Z(n22668) );
  NAND U23439 ( .A(n22669), .B(n22668), .Z(n22913) );
  XOR U23440 ( .A(b[51]), .B(n26122), .Z(n22817) );
  NANDN U23441 ( .A(n22817), .B(n37803), .Z(n22672) );
  NANDN U23442 ( .A(n22670), .B(n37802), .Z(n22671) );
  NAND U23443 ( .A(n22672), .B(n22671), .Z(n22910) );
  XOR U23444 ( .A(b[53]), .B(n25466), .Z(n22820) );
  NANDN U23445 ( .A(n22820), .B(n37940), .Z(n22675) );
  NANDN U23446 ( .A(n22673), .B(n37941), .Z(n22674) );
  AND U23447 ( .A(n22675), .B(n22674), .Z(n22911) );
  XNOR U23448 ( .A(n22910), .B(n22911), .Z(n22912) );
  XOR U23449 ( .A(n22913), .B(n22912), .Z(n22938) );
  XNOR U23450 ( .A(n22937), .B(n22938), .Z(n22939) );
  NANDN U23451 ( .A(n22677), .B(n22676), .Z(n22681) );
  NAND U23452 ( .A(n22679), .B(n22678), .Z(n22680) );
  NAND U23453 ( .A(n22681), .B(n22680), .Z(n22940) );
  XOR U23454 ( .A(n22939), .B(n22940), .Z(n22859) );
  NANDN U23455 ( .A(n22683), .B(n22682), .Z(n22687) );
  NAND U23456 ( .A(n22685), .B(n22684), .Z(n22686) );
  NAND U23457 ( .A(n22687), .B(n22686), .Z(n22856) );
  NANDN U23458 ( .A(n22689), .B(n22688), .Z(n22693) );
  NAND U23459 ( .A(n22691), .B(n22690), .Z(n22692) );
  AND U23460 ( .A(n22693), .B(n22692), .Z(n22857) );
  XNOR U23461 ( .A(n22856), .B(n22857), .Z(n22858) );
  XNOR U23462 ( .A(n22859), .B(n22858), .Z(n22992) );
  OR U23463 ( .A(n22695), .B(n22694), .Z(n22699) );
  OR U23464 ( .A(n22697), .B(n22696), .Z(n22698) );
  AND U23465 ( .A(n22699), .B(n22698), .Z(n22993) );
  XNOR U23466 ( .A(n22992), .B(n22993), .Z(n22994) );
  NANDN U23467 ( .A(n22701), .B(n22700), .Z(n22705) );
  NAND U23468 ( .A(n22703), .B(n22702), .Z(n22704) );
  AND U23469 ( .A(n22705), .B(n22704), .Z(n22995) );
  XNOR U23470 ( .A(n22994), .B(n22995), .Z(n22999) );
  XNOR U23471 ( .A(n22998), .B(n22999), .Z(n23001) );
  XNOR U23472 ( .A(n23000), .B(n23001), .Z(n23008) );
  XNOR U23473 ( .A(n23009), .B(n23008), .Z(n23011) );
  NAND U23474 ( .A(n22707), .B(n22706), .Z(n22711) );
  NANDN U23475 ( .A(n22709), .B(n22708), .Z(n22710) );
  AND U23476 ( .A(n22711), .B(n22710), .Z(n23010) );
  XNOR U23477 ( .A(n23011), .B(n23010), .Z(n23017) );
  XOR U23478 ( .A(n23016), .B(n23017), .Z(n23021) );
  NANDN U23479 ( .A(n22713), .B(n22712), .Z(n22717) );
  NAND U23480 ( .A(n22715), .B(n22714), .Z(n22716) );
  NAND U23481 ( .A(n22717), .B(n22716), .Z(n23018) );
  NANDN U23482 ( .A(n22719), .B(n22718), .Z(n22723) );
  NANDN U23483 ( .A(n22721), .B(n22720), .Z(n22722) );
  NAND U23484 ( .A(n22723), .B(n22722), .Z(n23019) );
  XNOR U23485 ( .A(n23018), .B(n23019), .Z(n23020) );
  XOR U23486 ( .A(n23021), .B(n23020), .Z(n23027) );
  OR U23487 ( .A(n22725), .B(n22724), .Z(n22729) );
  NAND U23488 ( .A(n22727), .B(n22726), .Z(n22728) );
  NAND U23489 ( .A(n22729), .B(n22728), .Z(n23025) );
  NANDN U23490 ( .A(n22731), .B(n22730), .Z(n22735) );
  NANDN U23491 ( .A(n22733), .B(n22732), .Z(n22734) );
  AND U23492 ( .A(n22735), .B(n22734), .Z(n23024) );
  XNOR U23493 ( .A(n23025), .B(n23024), .Z(n23026) );
  XOR U23494 ( .A(n23027), .B(n23026), .Z(n22747) );
  NANDN U23495 ( .A(n22737), .B(n22736), .Z(n22741) );
  NANDN U23496 ( .A(n22739), .B(n22738), .Z(n22740) );
  NAND U23497 ( .A(n22741), .B(n22740), .Z(n22748) );
  XOR U23498 ( .A(n22747), .B(n22748), .Z(n22749) );
  XNOR U23499 ( .A(n22750), .B(n22749), .Z(n23030) );
  XNOR U23500 ( .A(n23030), .B(sreg[171]), .Z(n23032) );
  NAND U23501 ( .A(n22742), .B(sreg[170]), .Z(n22746) );
  OR U23502 ( .A(n22744), .B(n22743), .Z(n22745) );
  AND U23503 ( .A(n22746), .B(n22745), .Z(n23031) );
  XOR U23504 ( .A(n23032), .B(n23031), .Z(c[171]) );
  OR U23505 ( .A(n22748), .B(n22747), .Z(n22752) );
  NAND U23506 ( .A(n22750), .B(n22749), .Z(n22751) );
  NAND U23507 ( .A(n22752), .B(n22751), .Z(n23038) );
  NANDN U23508 ( .A(n22754), .B(n22753), .Z(n22758) );
  NANDN U23509 ( .A(n22756), .B(n22755), .Z(n22757) );
  NAND U23510 ( .A(n22758), .B(n22757), .Z(n23297) );
  OR U23511 ( .A(n22760), .B(n22759), .Z(n22764) );
  NAND U23512 ( .A(n22762), .B(n22761), .Z(n22763) );
  NAND U23513 ( .A(n22764), .B(n22763), .Z(n23271) );
  XOR U23514 ( .A(a[98]), .B(n970), .Z(n23186) );
  OR U23515 ( .A(n23186), .B(n31369), .Z(n22767) );
  NANDN U23516 ( .A(n22765), .B(n31119), .Z(n22766) );
  NAND U23517 ( .A(n22767), .B(n22766), .Z(n23207) );
  XOR U23518 ( .A(b[43]), .B(n28701), .Z(n23189) );
  NANDN U23519 ( .A(n23189), .B(n37068), .Z(n22770) );
  NANDN U23520 ( .A(n22768), .B(n37069), .Z(n22769) );
  NAND U23521 ( .A(n22770), .B(n22769), .Z(n23204) );
  XOR U23522 ( .A(b[45]), .B(a[64]), .Z(n23192) );
  NAND U23523 ( .A(n23192), .B(n37261), .Z(n22773) );
  NAND U23524 ( .A(n22771), .B(n37262), .Z(n22772) );
  AND U23525 ( .A(n22773), .B(n22772), .Z(n23205) );
  XNOR U23526 ( .A(n23204), .B(n23205), .Z(n23206) );
  XNOR U23527 ( .A(n23207), .B(n23206), .Z(n23065) );
  XOR U23528 ( .A(b[49]), .B(n27436), .Z(n23195) );
  OR U23529 ( .A(n23195), .B(n37756), .Z(n22776) );
  NANDN U23530 ( .A(n22774), .B(n37652), .Z(n22775) );
  NAND U23531 ( .A(n22776), .B(n22775), .Z(n23183) );
  NAND U23532 ( .A(n37469), .B(n22777), .Z(n22779) );
  XNOR U23533 ( .A(n978), .B(a[62]), .Z(n23198) );
  NAND U23534 ( .A(n23198), .B(n37471), .Z(n22778) );
  AND U23535 ( .A(n22779), .B(n22778), .Z(n23180) );
  XOR U23536 ( .A(a[100]), .B(n969), .Z(n23201) );
  NANDN U23537 ( .A(n23201), .B(n30509), .Z(n22782) );
  NANDN U23538 ( .A(n22780), .B(n30846), .Z(n22781) );
  AND U23539 ( .A(n22782), .B(n22781), .Z(n23181) );
  XOR U23540 ( .A(n23183), .B(n23182), .Z(n23066) );
  XNOR U23541 ( .A(n23065), .B(n23066), .Z(n23067) );
  NANDN U23542 ( .A(n22784), .B(n22783), .Z(n22788) );
  NAND U23543 ( .A(n22786), .B(n22785), .Z(n22787) );
  AND U23544 ( .A(n22788), .B(n22787), .Z(n23068) );
  XNOR U23545 ( .A(n23067), .B(n23068), .Z(n23273) );
  XNOR U23546 ( .A(n23273), .B(n23272), .Z(n23274) );
  XNOR U23547 ( .A(b[35]), .B(a[74]), .Z(n23165) );
  NANDN U23548 ( .A(n23165), .B(n35985), .Z(n22795) );
  NAND U23549 ( .A(n22793), .B(n35986), .Z(n22794) );
  NAND U23550 ( .A(n22795), .B(n22794), .Z(n23241) );
  XOR U23551 ( .A(n36420), .B(n31123), .Z(n23168) );
  NAND U23552 ( .A(n23168), .B(n29949), .Z(n22798) );
  NAND U23553 ( .A(n29948), .B(n22796), .Z(n22797) );
  NAND U23554 ( .A(n22798), .B(n22797), .Z(n23238) );
  XOR U23555 ( .A(b[55]), .B(n25177), .Z(n23171) );
  NANDN U23556 ( .A(n23171), .B(n38075), .Z(n22801) );
  NANDN U23557 ( .A(n22799), .B(n38073), .Z(n22800) );
  AND U23558 ( .A(n22801), .B(n22800), .Z(n23239) );
  XNOR U23559 ( .A(n23238), .B(n23239), .Z(n23240) );
  XNOR U23560 ( .A(n23241), .B(n23240), .Z(n23044) );
  NANDN U23561 ( .A(n22803), .B(n22802), .Z(n22807) );
  NAND U23562 ( .A(n22805), .B(n22804), .Z(n22806) );
  NAND U23563 ( .A(n22807), .B(n22806), .Z(n23041) );
  NANDN U23564 ( .A(n22809), .B(n22808), .Z(n22813) );
  NAND U23565 ( .A(n22811), .B(n22810), .Z(n22812) );
  NAND U23566 ( .A(n22813), .B(n22812), .Z(n23042) );
  XNOR U23567 ( .A(n23041), .B(n23042), .Z(n23043) );
  XOR U23568 ( .A(n23044), .B(n23043), .Z(n23275) );
  XOR U23569 ( .A(n23274), .B(n23275), .Z(n23269) );
  XOR U23570 ( .A(b[39]), .B(n30379), .Z(n23223) );
  NANDN U23571 ( .A(n23223), .B(n36553), .Z(n22816) );
  NANDN U23572 ( .A(n22814), .B(n36643), .Z(n22815) );
  NAND U23573 ( .A(n22816), .B(n22815), .Z(n23092) );
  XOR U23574 ( .A(b[51]), .B(n26347), .Z(n23226) );
  NANDN U23575 ( .A(n23226), .B(n37803), .Z(n22819) );
  NANDN U23576 ( .A(n22817), .B(n37802), .Z(n22818) );
  NAND U23577 ( .A(n22819), .B(n22818), .Z(n23089) );
  XOR U23578 ( .A(b[53]), .B(n25860), .Z(n23229) );
  NANDN U23579 ( .A(n23229), .B(n37940), .Z(n22822) );
  NANDN U23580 ( .A(n22820), .B(n37941), .Z(n22821) );
  AND U23581 ( .A(n22822), .B(n22821), .Z(n23090) );
  XNOR U23582 ( .A(n23089), .B(n23090), .Z(n23091) );
  XNOR U23583 ( .A(n23092), .B(n23091), .Z(n23116) );
  XOR U23584 ( .A(a[94]), .B(n972), .Z(n23214) );
  OR U23585 ( .A(n23214), .B(n32010), .Z(n22825) );
  NANDN U23586 ( .A(n22823), .B(n32011), .Z(n22824) );
  NAND U23587 ( .A(n22825), .B(n22824), .Z(n23098) );
  XNOR U23588 ( .A(b[25]), .B(n33185), .Z(n23217) );
  NANDN U23589 ( .A(n34219), .B(n23217), .Z(n22828) );
  NAND U23590 ( .A(n34217), .B(n22826), .Z(n22827) );
  NAND U23591 ( .A(n22828), .B(n22827), .Z(n23095) );
  XNOR U23592 ( .A(a[92]), .B(b[17]), .Z(n23220) );
  NANDN U23593 ( .A(n23220), .B(n32543), .Z(n22831) );
  NAND U23594 ( .A(n22829), .B(n32541), .Z(n22830) );
  AND U23595 ( .A(n22831), .B(n22830), .Z(n23096) );
  XNOR U23596 ( .A(n23095), .B(n23096), .Z(n23097) );
  XOR U23597 ( .A(n23098), .B(n23097), .Z(n23117) );
  XOR U23598 ( .A(n23116), .B(n23117), .Z(n23119) );
  NANDN U23599 ( .A(n22833), .B(n22832), .Z(n22837) );
  NAND U23600 ( .A(n22835), .B(n22834), .Z(n22836) );
  NAND U23601 ( .A(n22837), .B(n22836), .Z(n23118) );
  XNOR U23602 ( .A(n23119), .B(n23118), .Z(n23259) );
  NANDN U23603 ( .A(n22839), .B(n22838), .Z(n22843) );
  NAND U23604 ( .A(n22841), .B(n22840), .Z(n22842) );
  NAND U23605 ( .A(n22843), .B(n22842), .Z(n23256) );
  NANDN U23606 ( .A(n22845), .B(n22844), .Z(n22849) );
  NAND U23607 ( .A(n22847), .B(n22846), .Z(n22848) );
  AND U23608 ( .A(n22849), .B(n22848), .Z(n23257) );
  XNOR U23609 ( .A(n23256), .B(n23257), .Z(n23258) );
  XNOR U23610 ( .A(n23259), .B(n23258), .Z(n23278) );
  OR U23611 ( .A(n22851), .B(n22850), .Z(n22855) );
  OR U23612 ( .A(n22853), .B(n22852), .Z(n22854) );
  AND U23613 ( .A(n22855), .B(n22854), .Z(n23279) );
  XOR U23614 ( .A(n23278), .B(n23279), .Z(n23281) );
  NANDN U23615 ( .A(n22857), .B(n22856), .Z(n22861) );
  NAND U23616 ( .A(n22859), .B(n22858), .Z(n22860) );
  NAND U23617 ( .A(n22861), .B(n22860), .Z(n23280) );
  XOR U23618 ( .A(n23281), .B(n23280), .Z(n23268) );
  XOR U23619 ( .A(n23269), .B(n23268), .Z(n23270) );
  XNOR U23620 ( .A(n23271), .B(n23270), .Z(n23295) );
  NANDN U23621 ( .A(n22863), .B(n22862), .Z(n22867) );
  OR U23622 ( .A(n22865), .B(n22864), .Z(n22866) );
  NAND U23623 ( .A(n22867), .B(n22866), .Z(n23262) );
  NANDN U23624 ( .A(n22869), .B(n22868), .Z(n22873) );
  OR U23625 ( .A(n22871), .B(n22870), .Z(n22872) );
  NAND U23626 ( .A(n22873), .B(n22872), .Z(n23286) );
  NANDN U23627 ( .A(n22875), .B(n22874), .Z(n22879) );
  NAND U23628 ( .A(n22877), .B(n22876), .Z(n22878) );
  NAND U23629 ( .A(n22879), .B(n22878), .Z(n23284) );
  NANDN U23630 ( .A(n22881), .B(n22880), .Z(n22885) );
  NAND U23631 ( .A(n22883), .B(n22882), .Z(n22884) );
  NAND U23632 ( .A(n22885), .B(n22884), .Z(n23285) );
  XNOR U23633 ( .A(n23284), .B(n23285), .Z(n23287) );
  XNOR U23634 ( .A(n23286), .B(n23287), .Z(n23263) );
  XOR U23635 ( .A(n23262), .B(n23263), .Z(n23264) );
  NANDN U23636 ( .A(n22887), .B(n22886), .Z(n22891) );
  NAND U23637 ( .A(n22889), .B(n22888), .Z(n22890) );
  NAND U23638 ( .A(n22891), .B(n22890), .Z(n23061) );
  XOR U23639 ( .A(b[37]), .B(n30210), .Z(n23071) );
  NANDN U23640 ( .A(n23071), .B(n36311), .Z(n22894) );
  NANDN U23641 ( .A(n22892), .B(n36309), .Z(n22893) );
  NAND U23642 ( .A(n22894), .B(n22893), .Z(n23125) );
  XOR U23643 ( .A(a[104]), .B(n968), .Z(n23074) );
  OR U23644 ( .A(n23074), .B(n29363), .Z(n22897) );
  NANDN U23645 ( .A(n22895), .B(n29864), .Z(n22896) );
  NAND U23646 ( .A(n22897), .B(n22896), .Z(n23122) );
  XOR U23647 ( .A(n36909), .B(n967), .Z(n23077) );
  NAND U23648 ( .A(n23077), .B(n28939), .Z(n22900) );
  NAND U23649 ( .A(n28938), .B(n22898), .Z(n22899) );
  AND U23650 ( .A(n22900), .B(n22899), .Z(n23123) );
  XNOR U23651 ( .A(n23122), .B(n23123), .Z(n23124) );
  XNOR U23652 ( .A(n23125), .B(n23124), .Z(n23056) );
  XOR U23653 ( .A(a[96]), .B(n971), .Z(n23080) );
  OR U23654 ( .A(n23080), .B(n31550), .Z(n22903) );
  NANDN U23655 ( .A(n22901), .B(n31874), .Z(n22902) );
  NAND U23656 ( .A(n22903), .B(n22902), .Z(n23235) );
  NAND U23657 ( .A(n34848), .B(n22904), .Z(n22906) );
  XOR U23658 ( .A(n35375), .B(n32815), .Z(n23083) );
  NAND U23659 ( .A(n34618), .B(n23083), .Z(n22905) );
  NAND U23660 ( .A(n22906), .B(n22905), .Z(n23232) );
  NAND U23661 ( .A(n35188), .B(n22907), .Z(n22909) );
  XOR U23662 ( .A(n35540), .B(n32814), .Z(n23086) );
  NANDN U23663 ( .A(n34968), .B(n23086), .Z(n22908) );
  AND U23664 ( .A(n22909), .B(n22908), .Z(n23233) );
  XNOR U23665 ( .A(n23232), .B(n23233), .Z(n23234) );
  XNOR U23666 ( .A(n23235), .B(n23234), .Z(n23053) );
  NANDN U23667 ( .A(n22911), .B(n22910), .Z(n22915) );
  NAND U23668 ( .A(n22913), .B(n22912), .Z(n22914) );
  NAND U23669 ( .A(n22915), .B(n22914), .Z(n23054) );
  XNOR U23670 ( .A(n23053), .B(n23054), .Z(n23055) );
  XOR U23671 ( .A(n23056), .B(n23055), .Z(n23060) );
  NANDN U23672 ( .A(n22917), .B(n22916), .Z(n22921) );
  NAND U23673 ( .A(n22919), .B(n22918), .Z(n22920) );
  NAND U23674 ( .A(n22921), .B(n22920), .Z(n23212) );
  NAND U23675 ( .A(a[44]), .B(b[63]), .Z(n23177) );
  NANDN U23676 ( .A(n22922), .B(n38369), .Z(n22924) );
  XOR U23677 ( .A(b[61]), .B(n23447), .Z(n23101) );
  OR U23678 ( .A(n23101), .B(n38371), .Z(n22923) );
  NAND U23679 ( .A(n22924), .B(n22923), .Z(n23175) );
  NANDN U23680 ( .A(n22925), .B(n35311), .Z(n22927) );
  XOR U23681 ( .A(b[31]), .B(n31870), .Z(n23104) );
  NANDN U23682 ( .A(n23104), .B(n35313), .Z(n22926) );
  AND U23683 ( .A(n22927), .B(n22926), .Z(n23174) );
  XNOR U23684 ( .A(n23175), .B(n23174), .Z(n23176) );
  XOR U23685 ( .A(n23177), .B(n23176), .Z(n23210) );
  NAND U23686 ( .A(n33283), .B(n22928), .Z(n22930) );
  XOR U23687 ( .A(n34851), .B(n33020), .Z(n23107) );
  NANDN U23688 ( .A(n33021), .B(n23107), .Z(n22929) );
  NAND U23689 ( .A(n22930), .B(n22929), .Z(n23131) );
  XNOR U23690 ( .A(a[88]), .B(b[21]), .Z(n23110) );
  OR U23691 ( .A(n23110), .B(n33634), .Z(n22933) );
  NAND U23692 ( .A(n22931), .B(n33464), .Z(n22932) );
  NAND U23693 ( .A(n22933), .B(n22932), .Z(n23128) );
  NAND U23694 ( .A(n34044), .B(n22934), .Z(n22936) );
  XOR U23695 ( .A(n34510), .B(n33628), .Z(n23113) );
  NANDN U23696 ( .A(n33867), .B(n23113), .Z(n22935) );
  AND U23697 ( .A(n22936), .B(n22935), .Z(n23129) );
  XNOR U23698 ( .A(n23128), .B(n23129), .Z(n23130) );
  XNOR U23699 ( .A(n23131), .B(n23130), .Z(n23211) );
  XNOR U23700 ( .A(n23210), .B(n23211), .Z(n23213) );
  XNOR U23701 ( .A(n23212), .B(n23213), .Z(n23059) );
  XOR U23702 ( .A(n23060), .B(n23059), .Z(n23062) );
  XNOR U23703 ( .A(n23061), .B(n23062), .Z(n23161) );
  NANDN U23704 ( .A(n22938), .B(n22937), .Z(n22942) );
  NANDN U23705 ( .A(n22940), .B(n22939), .Z(n22941) );
  NAND U23706 ( .A(n22942), .B(n22941), .Z(n23160) );
  NANDN U23707 ( .A(n22944), .B(n22943), .Z(n22948) );
  NAND U23708 ( .A(n22946), .B(n22945), .Z(n22947) );
  NAND U23709 ( .A(n22948), .B(n22947), .Z(n23050) );
  XNOR U23710 ( .A(b[41]), .B(a[68]), .Z(n23134) );
  OR U23711 ( .A(n23134), .B(n36905), .Z(n22951) );
  NANDN U23712 ( .A(n22949), .B(n36807), .Z(n22950) );
  NAND U23713 ( .A(n22951), .B(n22950), .Z(n23156) );
  XOR U23714 ( .A(b[57]), .B(n25134), .Z(n23137) );
  OR U23715 ( .A(n23137), .B(n965), .Z(n22954) );
  NANDN U23716 ( .A(n22952), .B(n38194), .Z(n22953) );
  NAND U23717 ( .A(n22954), .B(n22953), .Z(n23153) );
  NAND U23718 ( .A(n38326), .B(n22955), .Z(n22957) );
  XOR U23719 ( .A(n38400), .B(n24671), .Z(n23140) );
  NANDN U23720 ( .A(n38273), .B(n23140), .Z(n22956) );
  AND U23721 ( .A(n22957), .B(n22956), .Z(n23154) );
  XNOR U23722 ( .A(n23153), .B(n23154), .Z(n23155) );
  XOR U23723 ( .A(n23156), .B(n23155), .Z(n23250) );
  XOR U23724 ( .A(b[33]), .B(n31363), .Z(n23143) );
  NANDN U23725 ( .A(n23143), .B(n35620), .Z(n22960) );
  NANDN U23726 ( .A(n22958), .B(n35621), .Z(n22959) );
  NAND U23727 ( .A(n22960), .B(n22959), .Z(n23247) );
  NANDN U23728 ( .A(n966), .B(a[108]), .Z(n22961) );
  XOR U23729 ( .A(n29232), .B(n22961), .Z(n22963) );
  NANDN U23730 ( .A(b[0]), .B(a[107]), .Z(n22962) );
  AND U23731 ( .A(n22963), .B(n22962), .Z(n23244) );
  XOR U23732 ( .A(b[63]), .B(n22964), .Z(n23150) );
  NANDN U23733 ( .A(n23150), .B(n38422), .Z(n22967) );
  NANDN U23734 ( .A(n22965), .B(n38423), .Z(n22966) );
  AND U23735 ( .A(n22967), .B(n22966), .Z(n23245) );
  XNOR U23736 ( .A(n23244), .B(n23245), .Z(n23246) );
  XOR U23737 ( .A(n23247), .B(n23246), .Z(n23251) );
  XNOR U23738 ( .A(n23250), .B(n23251), .Z(n23253) );
  NANDN U23739 ( .A(n22969), .B(n22968), .Z(n22973) );
  NAND U23740 ( .A(n22971), .B(n22970), .Z(n22972) );
  NAND U23741 ( .A(n22973), .B(n22972), .Z(n23252) );
  XOR U23742 ( .A(n23253), .B(n23252), .Z(n23047) );
  NANDN U23743 ( .A(n22975), .B(n22974), .Z(n22979) );
  NAND U23744 ( .A(n22977), .B(n22976), .Z(n22978) );
  AND U23745 ( .A(n22979), .B(n22978), .Z(n23048) );
  XOR U23746 ( .A(n23047), .B(n23048), .Z(n23049) );
  XNOR U23747 ( .A(n23050), .B(n23049), .Z(n23159) );
  XNOR U23748 ( .A(n23160), .B(n23159), .Z(n23162) );
  XNOR U23749 ( .A(n23161), .B(n23162), .Z(n23265) );
  XOR U23750 ( .A(n23264), .B(n23265), .Z(n23294) );
  XNOR U23751 ( .A(n23295), .B(n23294), .Z(n23296) );
  XOR U23752 ( .A(n23297), .B(n23296), .Z(n23303) );
  NANDN U23753 ( .A(n22981), .B(n22980), .Z(n22985) );
  NAND U23754 ( .A(n22983), .B(n22982), .Z(n22984) );
  NAND U23755 ( .A(n22985), .B(n22984), .Z(n23291) );
  NANDN U23756 ( .A(n22987), .B(n22986), .Z(n22991) );
  NAND U23757 ( .A(n22989), .B(n22988), .Z(n22990) );
  NAND U23758 ( .A(n22991), .B(n22990), .Z(n23288) );
  NANDN U23759 ( .A(n22993), .B(n22992), .Z(n22997) );
  NAND U23760 ( .A(n22995), .B(n22994), .Z(n22996) );
  AND U23761 ( .A(n22997), .B(n22996), .Z(n23289) );
  XNOR U23762 ( .A(n23288), .B(n23289), .Z(n23290) );
  XOR U23763 ( .A(n23291), .B(n23290), .Z(n23301) );
  XOR U23764 ( .A(n23301), .B(n23300), .Z(n23302) );
  XOR U23765 ( .A(n23303), .B(n23302), .Z(n23309) );
  NANDN U23766 ( .A(n23003), .B(n23002), .Z(n23007) );
  NAND U23767 ( .A(n23005), .B(n23004), .Z(n23006) );
  NAND U23768 ( .A(n23007), .B(n23006), .Z(n23306) );
  NAND U23769 ( .A(n23009), .B(n23008), .Z(n23013) );
  NANDN U23770 ( .A(n23011), .B(n23010), .Z(n23012) );
  NAND U23771 ( .A(n23013), .B(n23012), .Z(n23307) );
  XNOR U23772 ( .A(n23306), .B(n23307), .Z(n23308) );
  XNOR U23773 ( .A(n23309), .B(n23308), .Z(n23313) );
  XOR U23774 ( .A(n23313), .B(n23312), .Z(n23314) );
  NANDN U23775 ( .A(n23019), .B(n23018), .Z(n23023) );
  NANDN U23776 ( .A(n23021), .B(n23020), .Z(n23022) );
  NAND U23777 ( .A(n23023), .B(n23022), .Z(n23315) );
  XOR U23778 ( .A(n23314), .B(n23315), .Z(n23035) );
  NANDN U23779 ( .A(n23025), .B(n23024), .Z(n23029) );
  NAND U23780 ( .A(n23027), .B(n23026), .Z(n23028) );
  NAND U23781 ( .A(n23029), .B(n23028), .Z(n23036) );
  XNOR U23782 ( .A(n23035), .B(n23036), .Z(n23037) );
  XNOR U23783 ( .A(n23038), .B(n23037), .Z(n23318) );
  XNOR U23784 ( .A(n23318), .B(sreg[172]), .Z(n23320) );
  NAND U23785 ( .A(n23030), .B(sreg[171]), .Z(n23034) );
  OR U23786 ( .A(n23032), .B(n23031), .Z(n23033) );
  AND U23787 ( .A(n23034), .B(n23033), .Z(n23319) );
  XOR U23788 ( .A(n23320), .B(n23319), .Z(c[172]) );
  NANDN U23789 ( .A(n23036), .B(n23035), .Z(n23040) );
  NAND U23790 ( .A(n23038), .B(n23037), .Z(n23039) );
  NAND U23791 ( .A(n23040), .B(n23039), .Z(n23326) );
  NANDN U23792 ( .A(n23042), .B(n23041), .Z(n23046) );
  NAND U23793 ( .A(n23044), .B(n23043), .Z(n23045) );
  AND U23794 ( .A(n23046), .B(n23045), .Z(n23581) );
  NAND U23795 ( .A(n23048), .B(n23047), .Z(n23052) );
  NANDN U23796 ( .A(n23050), .B(n23049), .Z(n23051) );
  NAND U23797 ( .A(n23052), .B(n23051), .Z(n23578) );
  NANDN U23798 ( .A(n23054), .B(n23053), .Z(n23058) );
  NAND U23799 ( .A(n23056), .B(n23055), .Z(n23057) );
  AND U23800 ( .A(n23058), .B(n23057), .Z(n23579) );
  XNOR U23801 ( .A(n23578), .B(n23579), .Z(n23580) );
  XNOR U23802 ( .A(n23581), .B(n23580), .Z(n23560) );
  NANDN U23803 ( .A(n23060), .B(n23059), .Z(n23064) );
  OR U23804 ( .A(n23062), .B(n23061), .Z(n23063) );
  AND U23805 ( .A(n23064), .B(n23063), .Z(n23561) );
  XNOR U23806 ( .A(n23560), .B(n23561), .Z(n23563) );
  NANDN U23807 ( .A(n23066), .B(n23065), .Z(n23070) );
  NAND U23808 ( .A(n23068), .B(n23067), .Z(n23069) );
  NAND U23809 ( .A(n23070), .B(n23069), .Z(n23361) );
  XNOR U23810 ( .A(b[37]), .B(a[73]), .Z(n23369) );
  NANDN U23811 ( .A(n23369), .B(n36311), .Z(n23073) );
  NANDN U23812 ( .A(n23071), .B(n36309), .Z(n23072) );
  NAND U23813 ( .A(n23073), .B(n23072), .Z(n23423) );
  XNOR U23814 ( .A(a[105]), .B(b[5]), .Z(n23372) );
  OR U23815 ( .A(n23372), .B(n29363), .Z(n23076) );
  NANDN U23816 ( .A(n23074), .B(n29864), .Z(n23075) );
  NAND U23817 ( .A(n23076), .B(n23075), .Z(n23420) );
  XNOR U23818 ( .A(a[107]), .B(n967), .Z(n23375) );
  NAND U23819 ( .A(n23375), .B(n28939), .Z(n23079) );
  NAND U23820 ( .A(n28938), .B(n23077), .Z(n23078) );
  AND U23821 ( .A(n23079), .B(n23078), .Z(n23421) );
  XNOR U23822 ( .A(n23420), .B(n23421), .Z(n23422) );
  XNOR U23823 ( .A(n23423), .B(n23422), .Z(n23355) );
  XNOR U23824 ( .A(a[97]), .B(b[13]), .Z(n23378) );
  OR U23825 ( .A(n23378), .B(n31550), .Z(n23082) );
  NANDN U23826 ( .A(n23080), .B(n31874), .Z(n23081) );
  NAND U23827 ( .A(n23082), .B(n23081), .Z(n23551) );
  NAND U23828 ( .A(n34848), .B(n23083), .Z(n23085) );
  XNOR U23829 ( .A(n35375), .B(a[83]), .Z(n23381) );
  NAND U23830 ( .A(n34618), .B(n23381), .Z(n23084) );
  NAND U23831 ( .A(n23085), .B(n23084), .Z(n23548) );
  NAND U23832 ( .A(n35188), .B(n23086), .Z(n23088) );
  XNOR U23833 ( .A(n35540), .B(a[81]), .Z(n23384) );
  NANDN U23834 ( .A(n34968), .B(n23384), .Z(n23087) );
  AND U23835 ( .A(n23088), .B(n23087), .Z(n23549) );
  XNOR U23836 ( .A(n23548), .B(n23549), .Z(n23550) );
  XNOR U23837 ( .A(n23551), .B(n23550), .Z(n23353) );
  NANDN U23838 ( .A(n23090), .B(n23089), .Z(n23094) );
  NAND U23839 ( .A(n23092), .B(n23091), .Z(n23093) );
  NAND U23840 ( .A(n23094), .B(n23093), .Z(n23354) );
  XOR U23841 ( .A(n23353), .B(n23354), .Z(n23356) );
  XNOR U23842 ( .A(n23355), .B(n23356), .Z(n23360) );
  NANDN U23843 ( .A(n23096), .B(n23095), .Z(n23100) );
  NAND U23844 ( .A(n23098), .B(n23097), .Z(n23099) );
  AND U23845 ( .A(n23100), .B(n23099), .Z(n23489) );
  NAND U23846 ( .A(a[45]), .B(b[63]), .Z(n23505) );
  NANDN U23847 ( .A(n23101), .B(n38369), .Z(n23103) );
  XOR U23848 ( .A(b[61]), .B(n23852), .Z(n23399) );
  OR U23849 ( .A(n23399), .B(n38371), .Z(n23102) );
  NAND U23850 ( .A(n23103), .B(n23102), .Z(n23503) );
  NANDN U23851 ( .A(n23104), .B(n35311), .Z(n23106) );
  XNOR U23852 ( .A(b[31]), .B(a[79]), .Z(n23402) );
  NANDN U23853 ( .A(n23402), .B(n35313), .Z(n23105) );
  AND U23854 ( .A(n23106), .B(n23105), .Z(n23502) );
  XNOR U23855 ( .A(n23503), .B(n23502), .Z(n23504) );
  XOR U23856 ( .A(n23505), .B(n23504), .Z(n23487) );
  NAND U23857 ( .A(n33283), .B(n23107), .Z(n23109) );
  XNOR U23858 ( .A(a[91]), .B(n33020), .Z(n23405) );
  NANDN U23859 ( .A(n33021), .B(n23405), .Z(n23108) );
  NAND U23860 ( .A(n23109), .B(n23108), .Z(n23429) );
  XOR U23861 ( .A(a[89]), .B(b[21]), .Z(n23408) );
  NANDN U23862 ( .A(n33634), .B(n23408), .Z(n23112) );
  NANDN U23863 ( .A(n23110), .B(n33464), .Z(n23111) );
  NAND U23864 ( .A(n23112), .B(n23111), .Z(n23426) );
  NAND U23865 ( .A(n34044), .B(n23113), .Z(n23115) );
  XNOR U23866 ( .A(n34510), .B(a[87]), .Z(n23411) );
  NANDN U23867 ( .A(n33867), .B(n23411), .Z(n23114) );
  AND U23868 ( .A(n23115), .B(n23114), .Z(n23427) );
  XNOR U23869 ( .A(n23426), .B(n23427), .Z(n23428) );
  XNOR U23870 ( .A(n23429), .B(n23428), .Z(n23488) );
  XNOR U23871 ( .A(n23487), .B(n23488), .Z(n23490) );
  XOR U23872 ( .A(n23489), .B(n23490), .Z(n23359) );
  XOR U23873 ( .A(n23360), .B(n23359), .Z(n23362) );
  XNOR U23874 ( .A(n23361), .B(n23362), .Z(n23459) );
  NANDN U23875 ( .A(n23117), .B(n23116), .Z(n23121) );
  OR U23876 ( .A(n23119), .B(n23118), .Z(n23120) );
  NAND U23877 ( .A(n23121), .B(n23120), .Z(n23458) );
  NANDN U23878 ( .A(n23123), .B(n23122), .Z(n23127) );
  NAND U23879 ( .A(n23125), .B(n23124), .Z(n23126) );
  NAND U23880 ( .A(n23127), .B(n23126), .Z(n23350) );
  NANDN U23881 ( .A(n23129), .B(n23128), .Z(n23133) );
  NAND U23882 ( .A(n23131), .B(n23130), .Z(n23132) );
  NAND U23883 ( .A(n23133), .B(n23132), .Z(n23517) );
  XOR U23884 ( .A(b[41]), .B(a[69]), .Z(n23432) );
  NANDN U23885 ( .A(n36905), .B(n23432), .Z(n23136) );
  NANDN U23886 ( .A(n23134), .B(n36807), .Z(n23135) );
  NAND U23887 ( .A(n23136), .B(n23135), .Z(n23454) );
  XOR U23888 ( .A(b[57]), .B(n25001), .Z(n23435) );
  OR U23889 ( .A(n23435), .B(n965), .Z(n23139) );
  NANDN U23890 ( .A(n23137), .B(n38194), .Z(n23138) );
  NAND U23891 ( .A(n23139), .B(n23138), .Z(n23451) );
  NAND U23892 ( .A(n38326), .B(n23140), .Z(n23142) );
  XOR U23893 ( .A(n38400), .B(n24288), .Z(n23438) );
  NANDN U23894 ( .A(n38273), .B(n23438), .Z(n23141) );
  AND U23895 ( .A(n23142), .B(n23141), .Z(n23452) );
  XNOR U23896 ( .A(n23451), .B(n23452), .Z(n23453) );
  XOR U23897 ( .A(n23454), .B(n23453), .Z(n23515) );
  XNOR U23898 ( .A(b[33]), .B(a[77]), .Z(n23441) );
  NANDN U23899 ( .A(n23441), .B(n35620), .Z(n23145) );
  NANDN U23900 ( .A(n23143), .B(n35621), .Z(n23144) );
  NAND U23901 ( .A(n23145), .B(n23144), .Z(n23529) );
  NANDN U23902 ( .A(n966), .B(a[109]), .Z(n23146) );
  XOR U23903 ( .A(n29232), .B(n23146), .Z(n23148) );
  IV U23904 ( .A(a[108]), .Z(n37139) );
  NANDN U23905 ( .A(n37139), .B(n966), .Z(n23147) );
  AND U23906 ( .A(n23148), .B(n23147), .Z(n23526) );
  XOR U23907 ( .A(b[63]), .B(n23149), .Z(n23448) );
  NANDN U23908 ( .A(n23448), .B(n38422), .Z(n23152) );
  NANDN U23909 ( .A(n23150), .B(n38423), .Z(n23151) );
  AND U23910 ( .A(n23152), .B(n23151), .Z(n23527) );
  XNOR U23911 ( .A(n23526), .B(n23527), .Z(n23528) );
  XNOR U23912 ( .A(n23529), .B(n23528), .Z(n23514) );
  XOR U23913 ( .A(n23515), .B(n23514), .Z(n23516) );
  XNOR U23914 ( .A(n23517), .B(n23516), .Z(n23348) );
  NANDN U23915 ( .A(n23154), .B(n23153), .Z(n23158) );
  NAND U23916 ( .A(n23156), .B(n23155), .Z(n23157) );
  AND U23917 ( .A(n23158), .B(n23157), .Z(n23347) );
  XNOR U23918 ( .A(n23348), .B(n23347), .Z(n23349) );
  XNOR U23919 ( .A(n23350), .B(n23349), .Z(n23457) );
  XNOR U23920 ( .A(n23458), .B(n23457), .Z(n23460) );
  XNOR U23921 ( .A(n23459), .B(n23460), .Z(n23562) );
  XOR U23922 ( .A(n23563), .B(n23562), .Z(n23329) );
  NAND U23923 ( .A(n23160), .B(n23159), .Z(n23164) );
  NANDN U23924 ( .A(n23162), .B(n23161), .Z(n23163) );
  NAND U23925 ( .A(n23164), .B(n23163), .Z(n23569) );
  XOR U23926 ( .A(b[35]), .B(a[75]), .Z(n23493) );
  NAND U23927 ( .A(n35985), .B(n23493), .Z(n23167) );
  NANDN U23928 ( .A(n23165), .B(n35986), .Z(n23166) );
  NAND U23929 ( .A(n23167), .B(n23166), .Z(n23557) );
  XNOR U23930 ( .A(a[103]), .B(n31123), .Z(n23496) );
  NAND U23931 ( .A(n23496), .B(n29949), .Z(n23170) );
  NAND U23932 ( .A(n29948), .B(n23168), .Z(n23169) );
  NAND U23933 ( .A(n23170), .B(n23169), .Z(n23554) );
  XOR U23934 ( .A(b[55]), .B(n25466), .Z(n23499) );
  NANDN U23935 ( .A(n23499), .B(n38075), .Z(n23173) );
  NANDN U23936 ( .A(n23171), .B(n38073), .Z(n23172) );
  AND U23937 ( .A(n23173), .B(n23172), .Z(n23555) );
  XNOR U23938 ( .A(n23554), .B(n23555), .Z(n23556) );
  XNOR U23939 ( .A(n23557), .B(n23556), .Z(n23344) );
  NANDN U23940 ( .A(n23175), .B(n23174), .Z(n23179) );
  NAND U23941 ( .A(n23177), .B(n23176), .Z(n23178) );
  NAND U23942 ( .A(n23179), .B(n23178), .Z(n23341) );
  OR U23943 ( .A(n23181), .B(n23180), .Z(n23185) );
  NAND U23944 ( .A(n23183), .B(n23182), .Z(n23184) );
  NAND U23945 ( .A(n23185), .B(n23184), .Z(n23342) );
  XNOR U23946 ( .A(n23341), .B(n23342), .Z(n23343) );
  XOR U23947 ( .A(n23344), .B(n23343), .Z(n23574) );
  XNOR U23948 ( .A(a[99]), .B(b[11]), .Z(n23463) );
  OR U23949 ( .A(n23463), .B(n31369), .Z(n23188) );
  NANDN U23950 ( .A(n23186), .B(n31119), .Z(n23187) );
  NAND U23951 ( .A(n23188), .B(n23187), .Z(n23484) );
  XOR U23952 ( .A(b[43]), .B(n29372), .Z(n23466) );
  NANDN U23953 ( .A(n23466), .B(n37068), .Z(n23191) );
  NANDN U23954 ( .A(n23189), .B(n37069), .Z(n23190) );
  NAND U23955 ( .A(n23191), .B(n23190), .Z(n23481) );
  XNOR U23956 ( .A(b[45]), .B(a[65]), .Z(n23469) );
  NANDN U23957 ( .A(n23469), .B(n37261), .Z(n23194) );
  NAND U23958 ( .A(n23192), .B(n37262), .Z(n23193) );
  AND U23959 ( .A(n23194), .B(n23193), .Z(n23482) );
  XNOR U23960 ( .A(n23481), .B(n23482), .Z(n23483) );
  XNOR U23961 ( .A(n23484), .B(n23483), .Z(n23368) );
  XOR U23962 ( .A(b[49]), .B(n27773), .Z(n23472) );
  OR U23963 ( .A(n23472), .B(n37756), .Z(n23197) );
  NANDN U23964 ( .A(n23195), .B(n37652), .Z(n23196) );
  NAND U23965 ( .A(n23197), .B(n23196), .Z(n23511) );
  NAND U23966 ( .A(n37469), .B(n23198), .Z(n23200) );
  XNOR U23967 ( .A(n978), .B(a[63]), .Z(n23475) );
  NAND U23968 ( .A(n23475), .B(n37471), .Z(n23199) );
  NAND U23969 ( .A(n23200), .B(n23199), .Z(n23508) );
  XNOR U23970 ( .A(a[101]), .B(b[9]), .Z(n23478) );
  NANDN U23971 ( .A(n23478), .B(n30509), .Z(n23203) );
  NANDN U23972 ( .A(n23201), .B(n30846), .Z(n23202) );
  AND U23973 ( .A(n23203), .B(n23202), .Z(n23509) );
  XNOR U23974 ( .A(n23508), .B(n23509), .Z(n23510) );
  XNOR U23975 ( .A(n23511), .B(n23510), .Z(n23365) );
  NANDN U23976 ( .A(n23205), .B(n23204), .Z(n23209) );
  NAND U23977 ( .A(n23207), .B(n23206), .Z(n23208) );
  NAND U23978 ( .A(n23209), .B(n23208), .Z(n23366) );
  XNOR U23979 ( .A(n23365), .B(n23366), .Z(n23367) );
  XOR U23980 ( .A(n23368), .B(n23367), .Z(n23572) );
  XOR U23981 ( .A(n23572), .B(n23573), .Z(n23575) );
  XNOR U23982 ( .A(n23574), .B(n23575), .Z(n23567) );
  XOR U23983 ( .A(a[95]), .B(n972), .Z(n23530) );
  OR U23984 ( .A(n23530), .B(n32010), .Z(n23216) );
  NANDN U23985 ( .A(n23214), .B(n32011), .Z(n23215) );
  NAND U23986 ( .A(n23216), .B(n23215), .Z(n23396) );
  XOR U23987 ( .A(b[25]), .B(a[85]), .Z(n23533) );
  NANDN U23988 ( .A(n34219), .B(n23533), .Z(n23219) );
  NAND U23989 ( .A(n34217), .B(n23217), .Z(n23218) );
  NAND U23990 ( .A(n23219), .B(n23218), .Z(n23393) );
  XNOR U23991 ( .A(a[93]), .B(b[17]), .Z(n23536) );
  NANDN U23992 ( .A(n23536), .B(n32543), .Z(n23222) );
  NANDN U23993 ( .A(n23220), .B(n32541), .Z(n23221) );
  AND U23994 ( .A(n23222), .B(n23221), .Z(n23394) );
  XNOR U23995 ( .A(n23393), .B(n23394), .Z(n23395) );
  XNOR U23996 ( .A(n23396), .B(n23395), .Z(n23414) );
  XOR U23997 ( .A(b[39]), .B(n30543), .Z(n23539) );
  NANDN U23998 ( .A(n23539), .B(n36553), .Z(n23225) );
  NANDN U23999 ( .A(n23223), .B(n36643), .Z(n23224) );
  NAND U24000 ( .A(n23225), .B(n23224), .Z(n23390) );
  XNOR U24001 ( .A(b[51]), .B(a[59]), .Z(n23542) );
  NANDN U24002 ( .A(n23542), .B(n37803), .Z(n23228) );
  NANDN U24003 ( .A(n23226), .B(n37802), .Z(n23227) );
  NAND U24004 ( .A(n23228), .B(n23227), .Z(n23387) );
  XOR U24005 ( .A(b[53]), .B(n26122), .Z(n23545) );
  NANDN U24006 ( .A(n23545), .B(n37940), .Z(n23231) );
  NANDN U24007 ( .A(n23229), .B(n37941), .Z(n23230) );
  AND U24008 ( .A(n23231), .B(n23230), .Z(n23388) );
  XNOR U24009 ( .A(n23387), .B(n23388), .Z(n23389) );
  XOR U24010 ( .A(n23390), .B(n23389), .Z(n23415) );
  XOR U24011 ( .A(n23414), .B(n23415), .Z(n23417) );
  NANDN U24012 ( .A(n23233), .B(n23232), .Z(n23237) );
  NAND U24013 ( .A(n23235), .B(n23234), .Z(n23236) );
  NAND U24014 ( .A(n23237), .B(n23236), .Z(n23416) );
  XNOR U24015 ( .A(n23417), .B(n23416), .Z(n23523) );
  NANDN U24016 ( .A(n23239), .B(n23238), .Z(n23243) );
  NAND U24017 ( .A(n23241), .B(n23240), .Z(n23242) );
  NAND U24018 ( .A(n23243), .B(n23242), .Z(n23520) );
  NANDN U24019 ( .A(n23245), .B(n23244), .Z(n23249) );
  NAND U24020 ( .A(n23247), .B(n23246), .Z(n23248) );
  AND U24021 ( .A(n23249), .B(n23248), .Z(n23521) );
  XNOR U24022 ( .A(n23520), .B(n23521), .Z(n23522) );
  XNOR U24023 ( .A(n23523), .B(n23522), .Z(n23582) );
  OR U24024 ( .A(n23251), .B(n23250), .Z(n23255) );
  OR U24025 ( .A(n23253), .B(n23252), .Z(n23254) );
  AND U24026 ( .A(n23255), .B(n23254), .Z(n23583) );
  XOR U24027 ( .A(n23582), .B(n23583), .Z(n23585) );
  NANDN U24028 ( .A(n23257), .B(n23256), .Z(n23261) );
  NAND U24029 ( .A(n23259), .B(n23258), .Z(n23260) );
  AND U24030 ( .A(n23261), .B(n23260), .Z(n23584) );
  XNOR U24031 ( .A(n23585), .B(n23584), .Z(n23566) );
  XOR U24032 ( .A(n23569), .B(n23568), .Z(n23330) );
  XNOR U24033 ( .A(n23329), .B(n23330), .Z(n23331) );
  OR U24034 ( .A(n23263), .B(n23262), .Z(n23267) );
  NAND U24035 ( .A(n23265), .B(n23264), .Z(n23266) );
  AND U24036 ( .A(n23267), .B(n23266), .Z(n23332) );
  XNOR U24037 ( .A(n23331), .B(n23332), .Z(n23591) );
  NANDN U24038 ( .A(n23273), .B(n23272), .Z(n23277) );
  NAND U24039 ( .A(n23275), .B(n23274), .Z(n23276) );
  NAND U24040 ( .A(n23277), .B(n23276), .Z(n23338) );
  NANDN U24041 ( .A(n23279), .B(n23278), .Z(n23283) );
  OR U24042 ( .A(n23281), .B(n23280), .Z(n23282) );
  NAND U24043 ( .A(n23283), .B(n23282), .Z(n23336) );
  XNOR U24044 ( .A(n23336), .B(n23335), .Z(n23337) );
  XNOR U24045 ( .A(n23338), .B(n23337), .Z(n23588) );
  XNOR U24046 ( .A(n23589), .B(n23588), .Z(n23590) );
  XNOR U24047 ( .A(n23591), .B(n23590), .Z(n23595) );
  NANDN U24048 ( .A(n23289), .B(n23288), .Z(n23293) );
  NAND U24049 ( .A(n23291), .B(n23290), .Z(n23292) );
  NAND U24050 ( .A(n23293), .B(n23292), .Z(n23592) );
  NANDN U24051 ( .A(n23295), .B(n23294), .Z(n23299) );
  NAND U24052 ( .A(n23297), .B(n23296), .Z(n23298) );
  AND U24053 ( .A(n23299), .B(n23298), .Z(n23593) );
  XNOR U24054 ( .A(n23592), .B(n23593), .Z(n23594) );
  XNOR U24055 ( .A(n23595), .B(n23594), .Z(n23601) );
  NANDN U24056 ( .A(n23301), .B(n23300), .Z(n23305) );
  OR U24057 ( .A(n23303), .B(n23302), .Z(n23304) );
  NAND U24058 ( .A(n23305), .B(n23304), .Z(n23598) );
  NANDN U24059 ( .A(n23307), .B(n23306), .Z(n23311) );
  NANDN U24060 ( .A(n23309), .B(n23308), .Z(n23310) );
  NAND U24061 ( .A(n23311), .B(n23310), .Z(n23599) );
  XNOR U24062 ( .A(n23598), .B(n23599), .Z(n23600) );
  XNOR U24063 ( .A(n23601), .B(n23600), .Z(n23323) );
  OR U24064 ( .A(n23313), .B(n23312), .Z(n23317) );
  NANDN U24065 ( .A(n23315), .B(n23314), .Z(n23316) );
  NAND U24066 ( .A(n23317), .B(n23316), .Z(n23324) );
  XOR U24067 ( .A(n23323), .B(n23324), .Z(n23325) );
  XNOR U24068 ( .A(n23326), .B(n23325), .Z(n23604) );
  XNOR U24069 ( .A(n23604), .B(sreg[173]), .Z(n23606) );
  NAND U24070 ( .A(n23318), .B(sreg[172]), .Z(n23322) );
  OR U24071 ( .A(n23320), .B(n23319), .Z(n23321) );
  AND U24072 ( .A(n23322), .B(n23321), .Z(n23605) );
  XOR U24073 ( .A(n23606), .B(n23605), .Z(c[173]) );
  OR U24074 ( .A(n23324), .B(n23323), .Z(n23328) );
  NAND U24075 ( .A(n23326), .B(n23325), .Z(n23327) );
  NAND U24076 ( .A(n23328), .B(n23327), .Z(n23612) );
  NANDN U24077 ( .A(n23330), .B(n23329), .Z(n23334) );
  NAND U24078 ( .A(n23332), .B(n23331), .Z(n23333) );
  NAND U24079 ( .A(n23334), .B(n23333), .Z(n23881) );
  NANDN U24080 ( .A(n23336), .B(n23335), .Z(n23340) );
  NANDN U24081 ( .A(n23338), .B(n23337), .Z(n23339) );
  AND U24082 ( .A(n23340), .B(n23339), .Z(n23880) );
  XNOR U24083 ( .A(n23881), .B(n23880), .Z(n23882) );
  NANDN U24084 ( .A(n23342), .B(n23341), .Z(n23346) );
  NAND U24085 ( .A(n23344), .B(n23343), .Z(n23345) );
  AND U24086 ( .A(n23346), .B(n23345), .Z(n23622) );
  NANDN U24087 ( .A(n23348), .B(n23347), .Z(n23352) );
  NANDN U24088 ( .A(n23350), .B(n23349), .Z(n23351) );
  AND U24089 ( .A(n23352), .B(n23351), .Z(n23619) );
  NANDN U24090 ( .A(n23354), .B(n23353), .Z(n23358) );
  NANDN U24091 ( .A(n23356), .B(n23355), .Z(n23357) );
  AND U24092 ( .A(n23358), .B(n23357), .Z(n23620) );
  XNOR U24093 ( .A(n23619), .B(n23620), .Z(n23621) );
  XOR U24094 ( .A(n23622), .B(n23621), .Z(n23637) );
  NANDN U24095 ( .A(n23360), .B(n23359), .Z(n23364) );
  OR U24096 ( .A(n23362), .B(n23361), .Z(n23363) );
  AND U24097 ( .A(n23364), .B(n23363), .Z(n23638) );
  XNOR U24098 ( .A(n23637), .B(n23638), .Z(n23640) );
  XOR U24099 ( .A(b[37]), .B(n31372), .Z(n23795) );
  NANDN U24100 ( .A(n23795), .B(n36311), .Z(n23371) );
  NANDN U24101 ( .A(n23369), .B(n36309), .Z(n23370) );
  NAND U24102 ( .A(n23371), .B(n23370), .Z(n23828) );
  XOR U24103 ( .A(a[106]), .B(n968), .Z(n23798) );
  OR U24104 ( .A(n23798), .B(n29363), .Z(n23374) );
  NANDN U24105 ( .A(n23372), .B(n29864), .Z(n23373) );
  NAND U24106 ( .A(n23374), .B(n23373), .Z(n23825) );
  XOR U24107 ( .A(n37139), .B(n967), .Z(n23801) );
  NAND U24108 ( .A(n23801), .B(n28939), .Z(n23377) );
  NAND U24109 ( .A(n28938), .B(n23375), .Z(n23376) );
  AND U24110 ( .A(n23377), .B(n23376), .Z(n23826) );
  XNOR U24111 ( .A(n23825), .B(n23826), .Z(n23827) );
  XNOR U24112 ( .A(n23828), .B(n23827), .Z(n23756) );
  XOR U24113 ( .A(a[98]), .B(n971), .Z(n23804) );
  OR U24114 ( .A(n23804), .B(n31550), .Z(n23380) );
  NANDN U24115 ( .A(n23378), .B(n31874), .Z(n23379) );
  NAND U24116 ( .A(n23380), .B(n23379), .Z(n23719) );
  NAND U24117 ( .A(n34848), .B(n23381), .Z(n23383) );
  XOR U24118 ( .A(n35375), .B(n33185), .Z(n23807) );
  NAND U24119 ( .A(n34618), .B(n23807), .Z(n23382) );
  NAND U24120 ( .A(n23383), .B(n23382), .Z(n23716) );
  NAND U24121 ( .A(n35188), .B(n23384), .Z(n23386) );
  XOR U24122 ( .A(n35540), .B(n32815), .Z(n23810) );
  NANDN U24123 ( .A(n34968), .B(n23810), .Z(n23385) );
  AND U24124 ( .A(n23386), .B(n23385), .Z(n23717) );
  XNOR U24125 ( .A(n23716), .B(n23717), .Z(n23718) );
  XOR U24126 ( .A(n23719), .B(n23718), .Z(n23757) );
  XOR U24127 ( .A(n23756), .B(n23757), .Z(n23759) );
  NANDN U24128 ( .A(n23388), .B(n23387), .Z(n23392) );
  NAND U24129 ( .A(n23390), .B(n23389), .Z(n23391) );
  NAND U24130 ( .A(n23392), .B(n23391), .Z(n23758) );
  XNOR U24131 ( .A(n23759), .B(n23758), .Z(n23763) );
  NANDN U24132 ( .A(n23394), .B(n23393), .Z(n23398) );
  NAND U24133 ( .A(n23396), .B(n23395), .Z(n23397) );
  NAND U24134 ( .A(n23398), .B(n23397), .Z(n23669) );
  NAND U24135 ( .A(a[46]), .B(b[63]), .Z(n23683) );
  NANDN U24136 ( .A(n23399), .B(n38369), .Z(n23401) );
  XOR U24137 ( .A(b[61]), .B(n24671), .Z(n23789) );
  OR U24138 ( .A(n23789), .B(n38371), .Z(n23400) );
  NAND U24139 ( .A(n23401), .B(n23400), .Z(n23681) );
  NANDN U24140 ( .A(n23402), .B(n35311), .Z(n23404) );
  XOR U24141 ( .A(b[31]), .B(n32814), .Z(n23792) );
  NANDN U24142 ( .A(n23792), .B(n35313), .Z(n23403) );
  AND U24143 ( .A(n23404), .B(n23403), .Z(n23680) );
  XNOR U24144 ( .A(n23681), .B(n23680), .Z(n23682) );
  XOR U24145 ( .A(n23683), .B(n23682), .Z(n23667) );
  NAND U24146 ( .A(n33283), .B(n23405), .Z(n23407) );
  XOR U24147 ( .A(n34852), .B(n33020), .Z(n23774) );
  NANDN U24148 ( .A(n33021), .B(n23774), .Z(n23406) );
  NAND U24149 ( .A(n23407), .B(n23406), .Z(n23834) );
  XNOR U24150 ( .A(a[90]), .B(b[21]), .Z(n23777) );
  OR U24151 ( .A(n23777), .B(n33634), .Z(n23410) );
  NAND U24152 ( .A(n23408), .B(n33464), .Z(n23409) );
  NAND U24153 ( .A(n23410), .B(n23409), .Z(n23831) );
  NAND U24154 ( .A(n34044), .B(n23411), .Z(n23413) );
  XOR U24155 ( .A(n34510), .B(n34048), .Z(n23780) );
  NANDN U24156 ( .A(n33867), .B(n23780), .Z(n23412) );
  AND U24157 ( .A(n23413), .B(n23412), .Z(n23832) );
  XNOR U24158 ( .A(n23831), .B(n23832), .Z(n23833) );
  XNOR U24159 ( .A(n23834), .B(n23833), .Z(n23668) );
  XNOR U24160 ( .A(n23667), .B(n23668), .Z(n23670) );
  XNOR U24161 ( .A(n23669), .B(n23670), .Z(n23762) );
  XNOR U24162 ( .A(n23763), .B(n23762), .Z(n23764) );
  XNOR U24163 ( .A(n23765), .B(n23764), .Z(n23740) );
  NANDN U24164 ( .A(n23415), .B(n23414), .Z(n23419) );
  OR U24165 ( .A(n23417), .B(n23416), .Z(n23418) );
  NAND U24166 ( .A(n23419), .B(n23418), .Z(n23739) );
  NANDN U24167 ( .A(n23421), .B(n23420), .Z(n23425) );
  NAND U24168 ( .A(n23423), .B(n23422), .Z(n23424) );
  NAND U24169 ( .A(n23425), .B(n23424), .Z(n23753) );
  NANDN U24170 ( .A(n23427), .B(n23426), .Z(n23431) );
  NAND U24171 ( .A(n23429), .B(n23428), .Z(n23430) );
  NAND U24172 ( .A(n23431), .B(n23430), .Z(n23735) );
  XNOR U24173 ( .A(b[41]), .B(a[70]), .Z(n23837) );
  OR U24174 ( .A(n23837), .B(n36905), .Z(n23434) );
  NAND U24175 ( .A(n23432), .B(n36807), .Z(n23433) );
  NAND U24176 ( .A(n23434), .B(n23433), .Z(n23859) );
  XOR U24177 ( .A(b[57]), .B(n25177), .Z(n23840) );
  OR U24178 ( .A(n23840), .B(n965), .Z(n23437) );
  NANDN U24179 ( .A(n23435), .B(n38194), .Z(n23436) );
  NAND U24180 ( .A(n23437), .B(n23436), .Z(n23856) );
  NAND U24181 ( .A(n38326), .B(n23438), .Z(n23440) );
  XOR U24182 ( .A(n38400), .B(n25134), .Z(n23843) );
  NANDN U24183 ( .A(n38273), .B(n23843), .Z(n23439) );
  AND U24184 ( .A(n23440), .B(n23439), .Z(n23857) );
  XNOR U24185 ( .A(n23856), .B(n23857), .Z(n23858) );
  XOR U24186 ( .A(n23859), .B(n23858), .Z(n23733) );
  XOR U24187 ( .A(b[33]), .B(n31870), .Z(n23846) );
  NANDN U24188 ( .A(n23846), .B(n35620), .Z(n23443) );
  NANDN U24189 ( .A(n23441), .B(n35621), .Z(n23442) );
  NAND U24190 ( .A(n23443), .B(n23442), .Z(n23731) );
  NANDN U24191 ( .A(n966), .B(a[110]), .Z(n23444) );
  XOR U24192 ( .A(n29232), .B(n23444), .Z(n23446) );
  NANDN U24193 ( .A(b[0]), .B(a[109]), .Z(n23445) );
  AND U24194 ( .A(n23446), .B(n23445), .Z(n23728) );
  XOR U24195 ( .A(b[63]), .B(n23447), .Z(n23853) );
  NANDN U24196 ( .A(n23853), .B(n38422), .Z(n23450) );
  NANDN U24197 ( .A(n23448), .B(n38423), .Z(n23449) );
  AND U24198 ( .A(n23450), .B(n23449), .Z(n23729) );
  XNOR U24199 ( .A(n23728), .B(n23729), .Z(n23730) );
  XNOR U24200 ( .A(n23731), .B(n23730), .Z(n23732) );
  XOR U24201 ( .A(n23733), .B(n23732), .Z(n23734) );
  XNOR U24202 ( .A(n23735), .B(n23734), .Z(n23751) );
  NANDN U24203 ( .A(n23452), .B(n23451), .Z(n23456) );
  NAND U24204 ( .A(n23454), .B(n23453), .Z(n23455) );
  AND U24205 ( .A(n23456), .B(n23455), .Z(n23750) );
  XNOR U24206 ( .A(n23751), .B(n23750), .Z(n23752) );
  XNOR U24207 ( .A(n23753), .B(n23752), .Z(n23738) );
  XNOR U24208 ( .A(n23739), .B(n23738), .Z(n23741) );
  XNOR U24209 ( .A(n23740), .B(n23741), .Z(n23639) );
  XOR U24210 ( .A(n23640), .B(n23639), .Z(n23868) );
  NAND U24211 ( .A(n23458), .B(n23457), .Z(n23462) );
  NANDN U24212 ( .A(n23460), .B(n23459), .Z(n23461) );
  NAND U24213 ( .A(n23462), .B(n23461), .Z(n23616) );
  XOR U24214 ( .A(a[100]), .B(n970), .Z(n23643) );
  OR U24215 ( .A(n23643), .B(n31369), .Z(n23465) );
  NANDN U24216 ( .A(n23463), .B(n31119), .Z(n23464) );
  NAND U24217 ( .A(n23465), .B(n23464), .Z(n23664) );
  XOR U24218 ( .A(b[43]), .B(n29868), .Z(n23646) );
  NANDN U24219 ( .A(n23646), .B(n37068), .Z(n23468) );
  NANDN U24220 ( .A(n23466), .B(n37069), .Z(n23467) );
  NAND U24221 ( .A(n23468), .B(n23467), .Z(n23661) );
  XNOR U24222 ( .A(b[45]), .B(a[66]), .Z(n23649) );
  NANDN U24223 ( .A(n23649), .B(n37261), .Z(n23471) );
  NANDN U24224 ( .A(n23469), .B(n37262), .Z(n23470) );
  AND U24225 ( .A(n23471), .B(n23470), .Z(n23662) );
  XNOR U24226 ( .A(n23661), .B(n23662), .Z(n23663) );
  XNOR U24227 ( .A(n23664), .B(n23663), .Z(n23768) );
  XNOR U24228 ( .A(b[49]), .B(a[62]), .Z(n23652) );
  OR U24229 ( .A(n23652), .B(n37756), .Z(n23474) );
  NANDN U24230 ( .A(n23472), .B(n37652), .Z(n23473) );
  NAND U24231 ( .A(n23474), .B(n23473), .Z(n23689) );
  NAND U24232 ( .A(n37469), .B(n23475), .Z(n23477) );
  XNOR U24233 ( .A(n978), .B(a[64]), .Z(n23655) );
  NAND U24234 ( .A(n23655), .B(n37471), .Z(n23476) );
  NAND U24235 ( .A(n23477), .B(n23476), .Z(n23686) );
  XOR U24236 ( .A(a[102]), .B(n969), .Z(n23658) );
  NANDN U24237 ( .A(n23658), .B(n30509), .Z(n23480) );
  NANDN U24238 ( .A(n23478), .B(n30846), .Z(n23479) );
  AND U24239 ( .A(n23480), .B(n23479), .Z(n23687) );
  XNOR U24240 ( .A(n23686), .B(n23687), .Z(n23688) );
  XOR U24241 ( .A(n23689), .B(n23688), .Z(n23769) );
  XNOR U24242 ( .A(n23768), .B(n23769), .Z(n23770) );
  NANDN U24243 ( .A(n23482), .B(n23481), .Z(n23486) );
  NAND U24244 ( .A(n23484), .B(n23483), .Z(n23485) );
  AND U24245 ( .A(n23486), .B(n23485), .Z(n23771) );
  XNOR U24246 ( .A(n23770), .B(n23771), .Z(n23632) );
  OR U24247 ( .A(n23488), .B(n23487), .Z(n23492) );
  OR U24248 ( .A(n23490), .B(n23489), .Z(n23491) );
  AND U24249 ( .A(n23492), .B(n23491), .Z(n23631) );
  XNOR U24250 ( .A(n23632), .B(n23631), .Z(n23633) );
  XNOR U24251 ( .A(b[35]), .B(a[76]), .Z(n23671) );
  NANDN U24252 ( .A(n23671), .B(n35985), .Z(n23495) );
  NAND U24253 ( .A(n23493), .B(n35986), .Z(n23494) );
  NAND U24254 ( .A(n23495), .B(n23494), .Z(n23725) );
  XOR U24255 ( .A(n36647), .B(n31123), .Z(n23674) );
  NAND U24256 ( .A(n23674), .B(n29949), .Z(n23498) );
  NAND U24257 ( .A(n29948), .B(n23496), .Z(n23497) );
  NAND U24258 ( .A(n23498), .B(n23497), .Z(n23722) );
  XOR U24259 ( .A(b[55]), .B(n25860), .Z(n23677) );
  NANDN U24260 ( .A(n23677), .B(n38075), .Z(n23501) );
  NANDN U24261 ( .A(n23499), .B(n38073), .Z(n23500) );
  AND U24262 ( .A(n23501), .B(n23500), .Z(n23723) );
  XNOR U24263 ( .A(n23722), .B(n23723), .Z(n23724) );
  XNOR U24264 ( .A(n23725), .B(n23724), .Z(n23747) );
  NANDN U24265 ( .A(n23503), .B(n23502), .Z(n23507) );
  NAND U24266 ( .A(n23505), .B(n23504), .Z(n23506) );
  NAND U24267 ( .A(n23507), .B(n23506), .Z(n23744) );
  NANDN U24268 ( .A(n23509), .B(n23508), .Z(n23513) );
  NAND U24269 ( .A(n23511), .B(n23510), .Z(n23512) );
  NAND U24270 ( .A(n23513), .B(n23512), .Z(n23745) );
  XNOR U24271 ( .A(n23744), .B(n23745), .Z(n23746) );
  XOR U24272 ( .A(n23747), .B(n23746), .Z(n23634) );
  XOR U24273 ( .A(n23633), .B(n23634), .Z(n23613) );
  NANDN U24274 ( .A(n23515), .B(n23514), .Z(n23519) );
  OR U24275 ( .A(n23517), .B(n23516), .Z(n23518) );
  NAND U24276 ( .A(n23519), .B(n23518), .Z(n23625) );
  NANDN U24277 ( .A(n23521), .B(n23520), .Z(n23525) );
  NAND U24278 ( .A(n23523), .B(n23522), .Z(n23524) );
  NAND U24279 ( .A(n23525), .B(n23524), .Z(n23626) );
  XNOR U24280 ( .A(n23625), .B(n23626), .Z(n23627) );
  XOR U24281 ( .A(a[96]), .B(n972), .Z(n23698) );
  OR U24282 ( .A(n23698), .B(n32010), .Z(n23532) );
  NANDN U24283 ( .A(n23530), .B(n32011), .Z(n23531) );
  NAND U24284 ( .A(n23532), .B(n23531), .Z(n23786) );
  XNOR U24285 ( .A(b[25]), .B(n33628), .Z(n23701) );
  NANDN U24286 ( .A(n34219), .B(n23701), .Z(n23535) );
  NAND U24287 ( .A(n34217), .B(n23533), .Z(n23534) );
  NAND U24288 ( .A(n23535), .B(n23534), .Z(n23783) );
  XNOR U24289 ( .A(a[94]), .B(b[17]), .Z(n23704) );
  NANDN U24290 ( .A(n23704), .B(n32543), .Z(n23538) );
  NANDN U24291 ( .A(n23536), .B(n32541), .Z(n23537) );
  AND U24292 ( .A(n23538), .B(n23537), .Z(n23784) );
  XNOR U24293 ( .A(n23783), .B(n23784), .Z(n23785) );
  XNOR U24294 ( .A(n23786), .B(n23785), .Z(n23819) );
  XOR U24295 ( .A(b[39]), .B(n30210), .Z(n23707) );
  NANDN U24296 ( .A(n23707), .B(n36553), .Z(n23541) );
  NANDN U24297 ( .A(n23539), .B(n36643), .Z(n23540) );
  NAND U24298 ( .A(n23541), .B(n23540), .Z(n23816) );
  XOR U24299 ( .A(b[51]), .B(n27436), .Z(n23710) );
  NANDN U24300 ( .A(n23710), .B(n37803), .Z(n23544) );
  NANDN U24301 ( .A(n23542), .B(n37802), .Z(n23543) );
  NAND U24302 ( .A(n23544), .B(n23543), .Z(n23813) );
  XOR U24303 ( .A(b[53]), .B(n26347), .Z(n23713) );
  NANDN U24304 ( .A(n23713), .B(n37940), .Z(n23547) );
  NANDN U24305 ( .A(n23545), .B(n37941), .Z(n23546) );
  AND U24306 ( .A(n23547), .B(n23546), .Z(n23814) );
  XNOR U24307 ( .A(n23813), .B(n23814), .Z(n23815) );
  XOR U24308 ( .A(n23816), .B(n23815), .Z(n23820) );
  XOR U24309 ( .A(n23819), .B(n23820), .Z(n23822) );
  NANDN U24310 ( .A(n23549), .B(n23548), .Z(n23553) );
  NAND U24311 ( .A(n23551), .B(n23550), .Z(n23552) );
  AND U24312 ( .A(n23553), .B(n23552), .Z(n23821) );
  XOR U24313 ( .A(n23822), .B(n23821), .Z(n23693) );
  NANDN U24314 ( .A(n23555), .B(n23554), .Z(n23559) );
  NAND U24315 ( .A(n23557), .B(n23556), .Z(n23558) );
  AND U24316 ( .A(n23559), .B(n23558), .Z(n23692) );
  XNOR U24317 ( .A(n23693), .B(n23692), .Z(n23694) );
  XOR U24318 ( .A(n23695), .B(n23694), .Z(n23628) );
  XNOR U24319 ( .A(n23627), .B(n23628), .Z(n23614) );
  XOR U24320 ( .A(n23613), .B(n23614), .Z(n23615) );
  XOR U24321 ( .A(n23616), .B(n23615), .Z(n23869) );
  XNOR U24322 ( .A(n23868), .B(n23869), .Z(n23870) );
  NAND U24323 ( .A(n23561), .B(n23560), .Z(n23565) );
  NANDN U24324 ( .A(n23563), .B(n23562), .Z(n23564) );
  NAND U24325 ( .A(n23565), .B(n23564), .Z(n23871) );
  XOR U24326 ( .A(n23870), .B(n23871), .Z(n23877) );
  NANDN U24327 ( .A(n23567), .B(n23566), .Z(n23571) );
  NAND U24328 ( .A(n23569), .B(n23568), .Z(n23570) );
  AND U24329 ( .A(n23571), .B(n23570), .Z(n23874) );
  NAND U24330 ( .A(n23573), .B(n23572), .Z(n23577) );
  NAND U24331 ( .A(n23575), .B(n23574), .Z(n23576) );
  NAND U24332 ( .A(n23577), .B(n23576), .Z(n23865) );
  NANDN U24333 ( .A(n23583), .B(n23582), .Z(n23587) );
  NANDN U24334 ( .A(n23585), .B(n23584), .Z(n23586) );
  AND U24335 ( .A(n23587), .B(n23586), .Z(n23863) );
  XNOR U24336 ( .A(n23862), .B(n23863), .Z(n23864) );
  XNOR U24337 ( .A(n23865), .B(n23864), .Z(n23875) );
  XNOR U24338 ( .A(n23877), .B(n23876), .Z(n23883) );
  XOR U24339 ( .A(n23882), .B(n23883), .Z(n23889) );
  NANDN U24340 ( .A(n23593), .B(n23592), .Z(n23597) );
  NANDN U24341 ( .A(n23595), .B(n23594), .Z(n23596) );
  NAND U24342 ( .A(n23597), .B(n23596), .Z(n23887) );
  XNOR U24343 ( .A(n23886), .B(n23887), .Z(n23888) );
  XNOR U24344 ( .A(n23889), .B(n23888), .Z(n23609) );
  NANDN U24345 ( .A(n23599), .B(n23598), .Z(n23603) );
  NANDN U24346 ( .A(n23601), .B(n23600), .Z(n23602) );
  NAND U24347 ( .A(n23603), .B(n23602), .Z(n23610) );
  XNOR U24348 ( .A(n23609), .B(n23610), .Z(n23611) );
  XNOR U24349 ( .A(n23612), .B(n23611), .Z(n23892) );
  XNOR U24350 ( .A(n23892), .B(sreg[174]), .Z(n23894) );
  NAND U24351 ( .A(n23604), .B(sreg[173]), .Z(n23608) );
  OR U24352 ( .A(n23606), .B(n23605), .Z(n23607) );
  AND U24353 ( .A(n23608), .B(n23607), .Z(n23893) );
  XOR U24354 ( .A(n23894), .B(n23893), .Z(c[174]) );
  NAND U24355 ( .A(n23614), .B(n23613), .Z(n23618) );
  NAND U24356 ( .A(n23616), .B(n23615), .Z(n23617) );
  NAND U24357 ( .A(n23618), .B(n23617), .Z(n24159) );
  OR U24358 ( .A(n23620), .B(n23619), .Z(n23624) );
  OR U24359 ( .A(n23622), .B(n23621), .Z(n23623) );
  NAND U24360 ( .A(n23624), .B(n23623), .Z(n23910) );
  NANDN U24361 ( .A(n23626), .B(n23625), .Z(n23630) );
  NANDN U24362 ( .A(n23628), .B(n23627), .Z(n23629) );
  NAND U24363 ( .A(n23630), .B(n23629), .Z(n23907) );
  NANDN U24364 ( .A(n23632), .B(n23631), .Z(n23636) );
  NAND U24365 ( .A(n23634), .B(n23633), .Z(n23635) );
  AND U24366 ( .A(n23636), .B(n23635), .Z(n23908) );
  XNOR U24367 ( .A(n23907), .B(n23908), .Z(n23909) );
  XNOR U24368 ( .A(n23910), .B(n23909), .Z(n24160) );
  XNOR U24369 ( .A(n24159), .B(n24160), .Z(n24161) );
  NAND U24370 ( .A(n23638), .B(n23637), .Z(n23642) );
  NANDN U24371 ( .A(n23640), .B(n23639), .Z(n23641) );
  NAND U24372 ( .A(n23642), .B(n23641), .Z(n23903) );
  XNOR U24373 ( .A(a[101]), .B(b[11]), .Z(n24116) );
  OR U24374 ( .A(n24116), .B(n31369), .Z(n23645) );
  NANDN U24375 ( .A(n23643), .B(n31119), .Z(n23644) );
  NAND U24376 ( .A(n23645), .B(n23644), .Z(n24128) );
  XNOR U24377 ( .A(b[43]), .B(a[69]), .Z(n24119) );
  NANDN U24378 ( .A(n24119), .B(n37068), .Z(n23648) );
  NANDN U24379 ( .A(n23646), .B(n37069), .Z(n23647) );
  NAND U24380 ( .A(n23648), .B(n23647), .Z(n24125) );
  XNOR U24381 ( .A(b[45]), .B(a[67]), .Z(n24122) );
  NANDN U24382 ( .A(n24122), .B(n37261), .Z(n23651) );
  NANDN U24383 ( .A(n23649), .B(n37262), .Z(n23650) );
  AND U24384 ( .A(n23651), .B(n23650), .Z(n24126) );
  XNOR U24385 ( .A(n24125), .B(n24126), .Z(n24127) );
  XNOR U24386 ( .A(n24128), .B(n24127), .Z(n23940) );
  XNOR U24387 ( .A(b[49]), .B(a[63]), .Z(n24107) );
  OR U24388 ( .A(n24107), .B(n37756), .Z(n23654) );
  NANDN U24389 ( .A(n23652), .B(n37652), .Z(n23653) );
  NAND U24390 ( .A(n23654), .B(n23653), .Z(n24097) );
  NAND U24391 ( .A(n37469), .B(n23655), .Z(n23657) );
  XOR U24392 ( .A(n978), .B(n28403), .Z(n24110) );
  NAND U24393 ( .A(n24110), .B(n37471), .Z(n23656) );
  AND U24394 ( .A(n23657), .B(n23656), .Z(n24095) );
  XNOR U24395 ( .A(a[103]), .B(b[9]), .Z(n24113) );
  NANDN U24396 ( .A(n24113), .B(n30509), .Z(n23660) );
  NANDN U24397 ( .A(n23658), .B(n30846), .Z(n23659) );
  AND U24398 ( .A(n23660), .B(n23659), .Z(n24096) );
  XOR U24399 ( .A(n24097), .B(n24098), .Z(n23937) );
  NANDN U24400 ( .A(n23662), .B(n23661), .Z(n23666) );
  NAND U24401 ( .A(n23664), .B(n23663), .Z(n23665) );
  NAND U24402 ( .A(n23666), .B(n23665), .Z(n23938) );
  XNOR U24403 ( .A(n23937), .B(n23938), .Z(n23939) );
  XOR U24404 ( .A(n23940), .B(n23939), .Z(n24137) );
  XNOR U24405 ( .A(n24137), .B(n24138), .Z(n24140) );
  XOR U24406 ( .A(b[35]), .B(a[77]), .Z(n24080) );
  NAND U24407 ( .A(n35985), .B(n24080), .Z(n23673) );
  NANDN U24408 ( .A(n23671), .B(n35986), .Z(n23672) );
  NAND U24409 ( .A(n23673), .B(n23672), .Z(n24073) );
  XNOR U24410 ( .A(a[105]), .B(n31123), .Z(n24083) );
  NAND U24411 ( .A(n24083), .B(n29949), .Z(n23676) );
  NAND U24412 ( .A(n29948), .B(n23674), .Z(n23675) );
  NAND U24413 ( .A(n23676), .B(n23675), .Z(n24070) );
  XOR U24414 ( .A(b[55]), .B(n26122), .Z(n24086) );
  NANDN U24415 ( .A(n24086), .B(n38075), .Z(n23679) );
  NANDN U24416 ( .A(n23677), .B(n38073), .Z(n23678) );
  AND U24417 ( .A(n23679), .B(n23678), .Z(n24071) );
  XNOR U24418 ( .A(n24070), .B(n24071), .Z(n24072) );
  XNOR U24419 ( .A(n24073), .B(n24072), .Z(n23916) );
  NANDN U24420 ( .A(n23681), .B(n23680), .Z(n23685) );
  NAND U24421 ( .A(n23683), .B(n23682), .Z(n23684) );
  NAND U24422 ( .A(n23685), .B(n23684), .Z(n23913) );
  NANDN U24423 ( .A(n23687), .B(n23686), .Z(n23691) );
  NAND U24424 ( .A(n23689), .B(n23688), .Z(n23690) );
  NAND U24425 ( .A(n23691), .B(n23690), .Z(n23914) );
  XNOR U24426 ( .A(n23913), .B(n23914), .Z(n23915) );
  XOR U24427 ( .A(n23916), .B(n23915), .Z(n24139) );
  XOR U24428 ( .A(n24140), .B(n24139), .Z(n24153) );
  NANDN U24429 ( .A(n23693), .B(n23692), .Z(n23697) );
  NANDN U24430 ( .A(n23695), .B(n23694), .Z(n23696) );
  NAND U24431 ( .A(n23697), .B(n23696), .Z(n24146) );
  XNOR U24432 ( .A(a[97]), .B(b[15]), .Z(n24055) );
  OR U24433 ( .A(n24055), .B(n32010), .Z(n23700) );
  NANDN U24434 ( .A(n23698), .B(n32011), .Z(n23699) );
  NAND U24435 ( .A(n23700), .B(n23699), .Z(n23953) );
  XOR U24436 ( .A(b[25]), .B(a[87]), .Z(n24058) );
  NANDN U24437 ( .A(n34219), .B(n24058), .Z(n23703) );
  NAND U24438 ( .A(n34217), .B(n23701), .Z(n23702) );
  NAND U24439 ( .A(n23703), .B(n23702), .Z(n23950) );
  XNOR U24440 ( .A(a[95]), .B(b[17]), .Z(n24061) );
  NANDN U24441 ( .A(n24061), .B(n32543), .Z(n23706) );
  NANDN U24442 ( .A(n23704), .B(n32541), .Z(n23705) );
  AND U24443 ( .A(n23706), .B(n23705), .Z(n23951) );
  XNOR U24444 ( .A(n23950), .B(n23951), .Z(n23952) );
  XNOR U24445 ( .A(n23953), .B(n23952), .Z(n23986) );
  XNOR U24446 ( .A(b[39]), .B(a[73]), .Z(n24046) );
  NANDN U24447 ( .A(n24046), .B(n36553), .Z(n23709) );
  NANDN U24448 ( .A(n23707), .B(n36643), .Z(n23708) );
  NAND U24449 ( .A(n23709), .B(n23708), .Z(n23983) );
  XOR U24450 ( .A(b[51]), .B(n27773), .Z(n24049) );
  NANDN U24451 ( .A(n24049), .B(n37803), .Z(n23712) );
  NANDN U24452 ( .A(n23710), .B(n37802), .Z(n23711) );
  NAND U24453 ( .A(n23712), .B(n23711), .Z(n23980) );
  XNOR U24454 ( .A(b[53]), .B(a[59]), .Z(n24052) );
  NANDN U24455 ( .A(n24052), .B(n37940), .Z(n23715) );
  NANDN U24456 ( .A(n23713), .B(n37941), .Z(n23714) );
  AND U24457 ( .A(n23715), .B(n23714), .Z(n23981) );
  XNOR U24458 ( .A(n23980), .B(n23981), .Z(n23982) );
  XOR U24459 ( .A(n23983), .B(n23982), .Z(n23987) );
  XNOR U24460 ( .A(n23986), .B(n23987), .Z(n23988) );
  NANDN U24461 ( .A(n23717), .B(n23716), .Z(n23721) );
  NAND U24462 ( .A(n23719), .B(n23718), .Z(n23720) );
  NAND U24463 ( .A(n23721), .B(n23720), .Z(n23989) );
  XOR U24464 ( .A(n23988), .B(n23989), .Z(n24037) );
  NANDN U24465 ( .A(n23723), .B(n23722), .Z(n23727) );
  NAND U24466 ( .A(n23725), .B(n23724), .Z(n23726) );
  NAND U24467 ( .A(n23727), .B(n23726), .Z(n24034) );
  XNOR U24468 ( .A(n24034), .B(n24035), .Z(n24036) );
  XNOR U24469 ( .A(n24037), .B(n24036), .Z(n24143) );
  NANDN U24470 ( .A(n23733), .B(n23732), .Z(n23737) );
  OR U24471 ( .A(n23735), .B(n23734), .Z(n23736) );
  AND U24472 ( .A(n23737), .B(n23736), .Z(n24144) );
  XNOR U24473 ( .A(n24143), .B(n24144), .Z(n24145) );
  XOR U24474 ( .A(n24146), .B(n24145), .Z(n24154) );
  XNOR U24475 ( .A(n24153), .B(n24154), .Z(n24155) );
  NAND U24476 ( .A(n23739), .B(n23738), .Z(n23743) );
  NANDN U24477 ( .A(n23741), .B(n23740), .Z(n23742) );
  NAND U24478 ( .A(n23743), .B(n23742), .Z(n24156) );
  XOR U24479 ( .A(n24155), .B(n24156), .Z(n23902) );
  NANDN U24480 ( .A(n23745), .B(n23744), .Z(n23749) );
  NAND U24481 ( .A(n23747), .B(n23746), .Z(n23748) );
  AND U24482 ( .A(n23749), .B(n23748), .Z(n24152) );
  NANDN U24483 ( .A(n23751), .B(n23750), .Z(n23755) );
  NANDN U24484 ( .A(n23753), .B(n23752), .Z(n23754) );
  NAND U24485 ( .A(n23755), .B(n23754), .Z(n24149) );
  NANDN U24486 ( .A(n23757), .B(n23756), .Z(n23761) );
  OR U24487 ( .A(n23759), .B(n23758), .Z(n23760) );
  AND U24488 ( .A(n23761), .B(n23760), .Z(n24150) );
  XNOR U24489 ( .A(n24149), .B(n24150), .Z(n24151) );
  XNOR U24490 ( .A(n24152), .B(n24151), .Z(n24131) );
  NAND U24491 ( .A(n23763), .B(n23762), .Z(n23767) );
  OR U24492 ( .A(n23765), .B(n23764), .Z(n23766) );
  AND U24493 ( .A(n23767), .B(n23766), .Z(n24132) );
  XNOR U24494 ( .A(n24131), .B(n24132), .Z(n24134) );
  NANDN U24495 ( .A(n23769), .B(n23768), .Z(n23773) );
  NAND U24496 ( .A(n23771), .B(n23770), .Z(n23772) );
  NAND U24497 ( .A(n23773), .B(n23772), .Z(n23933) );
  NAND U24498 ( .A(n33283), .B(n23774), .Z(n23776) );
  XOR U24499 ( .A(n35377), .B(n33020), .Z(n23941) );
  NANDN U24500 ( .A(n33021), .B(n23941), .Z(n23775) );
  NAND U24501 ( .A(n23776), .B(n23775), .Z(n24019) );
  XOR U24502 ( .A(a[91]), .B(b[21]), .Z(n23944) );
  NANDN U24503 ( .A(n33634), .B(n23944), .Z(n23779) );
  NANDN U24504 ( .A(n23777), .B(n33464), .Z(n23778) );
  NAND U24505 ( .A(n23779), .B(n23778), .Z(n24016) );
  NAND U24506 ( .A(n34044), .B(n23780), .Z(n23782) );
  XNOR U24507 ( .A(n34510), .B(a[89]), .Z(n23947) );
  NANDN U24508 ( .A(n33867), .B(n23947), .Z(n23781) );
  AND U24509 ( .A(n23782), .B(n23781), .Z(n24017) );
  XNOR U24510 ( .A(n24016), .B(n24017), .Z(n24018) );
  XOR U24511 ( .A(n24019), .B(n24018), .Z(n24101) );
  NANDN U24512 ( .A(n23784), .B(n23783), .Z(n23788) );
  NAND U24513 ( .A(n23786), .B(n23785), .Z(n23787) );
  NAND U24514 ( .A(n23788), .B(n23787), .Z(n24102) );
  XNOR U24515 ( .A(n24101), .B(n24102), .Z(n24104) );
  NAND U24516 ( .A(a[47]), .B(b[63]), .Z(n24092) );
  NANDN U24517 ( .A(n23789), .B(n38369), .Z(n23791) );
  XOR U24518 ( .A(b[61]), .B(n24288), .Z(n23956) );
  OR U24519 ( .A(n23956), .B(n38371), .Z(n23790) );
  NAND U24520 ( .A(n23791), .B(n23790), .Z(n24090) );
  NANDN U24521 ( .A(n23792), .B(n35311), .Z(n23794) );
  XNOR U24522 ( .A(b[31]), .B(a[81]), .Z(n23959) );
  NANDN U24523 ( .A(n23959), .B(n35313), .Z(n23793) );
  AND U24524 ( .A(n23794), .B(n23793), .Z(n24089) );
  XNOR U24525 ( .A(n24090), .B(n24089), .Z(n24091) );
  XNOR U24526 ( .A(n24092), .B(n24091), .Z(n24103) );
  XNOR U24527 ( .A(n24104), .B(n24103), .Z(n23931) );
  XNOR U24528 ( .A(b[37]), .B(a[75]), .Z(n23962) );
  NANDN U24529 ( .A(n23962), .B(n36311), .Z(n23797) );
  NANDN U24530 ( .A(n23795), .B(n36309), .Z(n23796) );
  NAND U24531 ( .A(n23797), .B(n23796), .Z(n23995) );
  XNOR U24532 ( .A(a[107]), .B(b[5]), .Z(n23965) );
  OR U24533 ( .A(n23965), .B(n29363), .Z(n23800) );
  NANDN U24534 ( .A(n23798), .B(n29864), .Z(n23799) );
  NAND U24535 ( .A(n23800), .B(n23799), .Z(n23992) );
  XNOR U24536 ( .A(a[109]), .B(n967), .Z(n23968) );
  NAND U24537 ( .A(n23968), .B(n28939), .Z(n23803) );
  NAND U24538 ( .A(n28938), .B(n23801), .Z(n23802) );
  AND U24539 ( .A(n23803), .B(n23802), .Z(n23993) );
  XNOR U24540 ( .A(n23992), .B(n23993), .Z(n23994) );
  XNOR U24541 ( .A(n23995), .B(n23994), .Z(n23925) );
  XNOR U24542 ( .A(a[99]), .B(b[13]), .Z(n23971) );
  OR U24543 ( .A(n23971), .B(n31550), .Z(n23806) );
  NANDN U24544 ( .A(n23804), .B(n31874), .Z(n23805) );
  NAND U24545 ( .A(n23806), .B(n23805), .Z(n24067) );
  NAND U24546 ( .A(n34848), .B(n23807), .Z(n23809) );
  XNOR U24547 ( .A(n35375), .B(a[85]), .Z(n23974) );
  NAND U24548 ( .A(n34618), .B(n23974), .Z(n23808) );
  NAND U24549 ( .A(n23809), .B(n23808), .Z(n24064) );
  NAND U24550 ( .A(n35188), .B(n23810), .Z(n23812) );
  XNOR U24551 ( .A(n35540), .B(a[83]), .Z(n23977) );
  NANDN U24552 ( .A(n34968), .B(n23977), .Z(n23811) );
  AND U24553 ( .A(n23812), .B(n23811), .Z(n24065) );
  XNOR U24554 ( .A(n24064), .B(n24065), .Z(n24066) );
  XOR U24555 ( .A(n24067), .B(n24066), .Z(n23926) );
  XOR U24556 ( .A(n23925), .B(n23926), .Z(n23928) );
  NANDN U24557 ( .A(n23814), .B(n23813), .Z(n23818) );
  NAND U24558 ( .A(n23816), .B(n23815), .Z(n23817) );
  NAND U24559 ( .A(n23818), .B(n23817), .Z(n23927) );
  XOR U24560 ( .A(n23928), .B(n23927), .Z(n23932) );
  XOR U24561 ( .A(n23931), .B(n23932), .Z(n23934) );
  XNOR U24562 ( .A(n23933), .B(n23934), .Z(n24030) );
  NANDN U24563 ( .A(n23820), .B(n23819), .Z(n23824) );
  NANDN U24564 ( .A(n23822), .B(n23821), .Z(n23823) );
  NAND U24565 ( .A(n23824), .B(n23823), .Z(n24029) );
  NANDN U24566 ( .A(n23826), .B(n23825), .Z(n23830) );
  NAND U24567 ( .A(n23828), .B(n23827), .Z(n23829) );
  NAND U24568 ( .A(n23830), .B(n23829), .Z(n23922) );
  NANDN U24569 ( .A(n23832), .B(n23831), .Z(n23836) );
  NAND U24570 ( .A(n23834), .B(n23833), .Z(n23835) );
  NAND U24571 ( .A(n23836), .B(n23835), .Z(n24043) );
  XNOR U24572 ( .A(b[41]), .B(a[71]), .Z(n24007) );
  OR U24573 ( .A(n24007), .B(n36905), .Z(n23839) );
  NANDN U24574 ( .A(n23837), .B(n36807), .Z(n23838) );
  NAND U24575 ( .A(n23839), .B(n23838), .Z(n24025) );
  XOR U24576 ( .A(b[57]), .B(n25466), .Z(n24010) );
  OR U24577 ( .A(n24010), .B(n965), .Z(n23842) );
  NANDN U24578 ( .A(n23840), .B(n38194), .Z(n23841) );
  NAND U24579 ( .A(n23842), .B(n23841), .Z(n24022) );
  NAND U24580 ( .A(n38326), .B(n23843), .Z(n23845) );
  XOR U24581 ( .A(n38400), .B(n25001), .Z(n24013) );
  NANDN U24582 ( .A(n38273), .B(n24013), .Z(n23844) );
  AND U24583 ( .A(n23845), .B(n23844), .Z(n24023) );
  XNOR U24584 ( .A(n24022), .B(n24023), .Z(n24024) );
  XOR U24585 ( .A(n24025), .B(n24024), .Z(n24041) );
  XNOR U24586 ( .A(b[33]), .B(a[79]), .Z(n23998) );
  NANDN U24587 ( .A(n23998), .B(n35620), .Z(n23848) );
  NANDN U24588 ( .A(n23846), .B(n35621), .Z(n23847) );
  NAND U24589 ( .A(n23848), .B(n23847), .Z(n24079) );
  NANDN U24590 ( .A(n966), .B(a[111]), .Z(n23849) );
  XOR U24591 ( .A(n29232), .B(n23849), .Z(n23851) );
  IV U24592 ( .A(a[110]), .Z(n37336) );
  NANDN U24593 ( .A(n37336), .B(n966), .Z(n23850) );
  AND U24594 ( .A(n23851), .B(n23850), .Z(n24076) );
  XOR U24595 ( .A(b[63]), .B(n23852), .Z(n24004) );
  NANDN U24596 ( .A(n24004), .B(n38422), .Z(n23855) );
  NANDN U24597 ( .A(n23853), .B(n38423), .Z(n23854) );
  AND U24598 ( .A(n23855), .B(n23854), .Z(n24077) );
  XNOR U24599 ( .A(n24076), .B(n24077), .Z(n24078) );
  XNOR U24600 ( .A(n24079), .B(n24078), .Z(n24040) );
  XOR U24601 ( .A(n24041), .B(n24040), .Z(n24042) );
  XNOR U24602 ( .A(n24043), .B(n24042), .Z(n23920) );
  NANDN U24603 ( .A(n23857), .B(n23856), .Z(n23861) );
  NAND U24604 ( .A(n23859), .B(n23858), .Z(n23860) );
  AND U24605 ( .A(n23861), .B(n23860), .Z(n23919) );
  XNOR U24606 ( .A(n23920), .B(n23919), .Z(n23921) );
  XNOR U24607 ( .A(n23922), .B(n23921), .Z(n24028) );
  XNOR U24608 ( .A(n24029), .B(n24028), .Z(n24031) );
  XNOR U24609 ( .A(n24030), .B(n24031), .Z(n24133) );
  XNOR U24610 ( .A(n24134), .B(n24133), .Z(n23901) );
  XNOR U24611 ( .A(n23902), .B(n23901), .Z(n23904) );
  XNOR U24612 ( .A(n23903), .B(n23904), .Z(n24162) );
  XOR U24613 ( .A(n24161), .B(n24162), .Z(n24167) );
  NANDN U24614 ( .A(n23863), .B(n23862), .Z(n23867) );
  NAND U24615 ( .A(n23865), .B(n23864), .Z(n23866) );
  NAND U24616 ( .A(n23867), .B(n23866), .Z(n24165) );
  NANDN U24617 ( .A(n23869), .B(n23868), .Z(n23873) );
  NANDN U24618 ( .A(n23871), .B(n23870), .Z(n23872) );
  NAND U24619 ( .A(n23873), .B(n23872), .Z(n24166) );
  XNOR U24620 ( .A(n24165), .B(n24166), .Z(n24168) );
  XNOR U24621 ( .A(n24167), .B(n24168), .Z(n24173) );
  OR U24622 ( .A(n23875), .B(n23874), .Z(n23879) );
  NAND U24623 ( .A(n23877), .B(n23876), .Z(n23878) );
  NAND U24624 ( .A(n23879), .B(n23878), .Z(n24172) );
  NANDN U24625 ( .A(n23881), .B(n23880), .Z(n23885) );
  NANDN U24626 ( .A(n23883), .B(n23882), .Z(n23884) );
  AND U24627 ( .A(n23885), .B(n23884), .Z(n24171) );
  XNOR U24628 ( .A(n24172), .B(n24171), .Z(n24174) );
  XNOR U24629 ( .A(n24173), .B(n24174), .Z(n23897) );
  NANDN U24630 ( .A(n23887), .B(n23886), .Z(n23891) );
  NAND U24631 ( .A(n23889), .B(n23888), .Z(n23890) );
  NAND U24632 ( .A(n23891), .B(n23890), .Z(n23898) );
  XNOR U24633 ( .A(n23897), .B(n23898), .Z(n23899) );
  XNOR U24634 ( .A(n23900), .B(n23899), .Z(n24175) );
  XNOR U24635 ( .A(n24175), .B(sreg[175]), .Z(n24177) );
  NAND U24636 ( .A(n23892), .B(sreg[174]), .Z(n23896) );
  OR U24637 ( .A(n23894), .B(n23893), .Z(n23895) );
  AND U24638 ( .A(n23896), .B(n23895), .Z(n24176) );
  XOR U24639 ( .A(n24177), .B(n24176), .Z(c[175]) );
  NAND U24640 ( .A(n23902), .B(n23901), .Z(n23906) );
  NANDN U24641 ( .A(n23904), .B(n23903), .Z(n23905) );
  NAND U24642 ( .A(n23906), .B(n23905), .Z(n24455) );
  NANDN U24643 ( .A(n23908), .B(n23907), .Z(n23912) );
  NAND U24644 ( .A(n23910), .B(n23909), .Z(n23911) );
  AND U24645 ( .A(n23912), .B(n23911), .Z(n24456) );
  XNOR U24646 ( .A(n24455), .B(n24456), .Z(n24457) );
  NANDN U24647 ( .A(n23914), .B(n23913), .Z(n23918) );
  NAND U24648 ( .A(n23916), .B(n23915), .Z(n23917) );
  AND U24649 ( .A(n23918), .B(n23917), .Z(n24442) );
  NANDN U24650 ( .A(n23920), .B(n23919), .Z(n23924) );
  NANDN U24651 ( .A(n23922), .B(n23921), .Z(n23923) );
  NAND U24652 ( .A(n23924), .B(n23923), .Z(n24439) );
  NANDN U24653 ( .A(n23926), .B(n23925), .Z(n23930) );
  OR U24654 ( .A(n23928), .B(n23927), .Z(n23929) );
  AND U24655 ( .A(n23930), .B(n23929), .Z(n24440) );
  XNOR U24656 ( .A(n24439), .B(n24440), .Z(n24441) );
  XNOR U24657 ( .A(n24442), .B(n24441), .Z(n24421) );
  NANDN U24658 ( .A(n23932), .B(n23931), .Z(n23936) );
  OR U24659 ( .A(n23934), .B(n23933), .Z(n23935) );
  AND U24660 ( .A(n23936), .B(n23935), .Z(n24422) );
  XNOR U24661 ( .A(n24421), .B(n24422), .Z(n24424) );
  NAND U24662 ( .A(n33283), .B(n23941), .Z(n23943) );
  XOR U24663 ( .A(n35191), .B(n33020), .Z(n24228) );
  NANDN U24664 ( .A(n33021), .B(n24228), .Z(n23942) );
  NAND U24665 ( .A(n23943), .B(n23942), .Z(n24295) );
  XNOR U24666 ( .A(a[92]), .B(b[21]), .Z(n24231) );
  OR U24667 ( .A(n24231), .B(n33634), .Z(n23946) );
  NAND U24668 ( .A(n23944), .B(n33464), .Z(n23945) );
  NAND U24669 ( .A(n23946), .B(n23945), .Z(n24292) );
  NAND U24670 ( .A(n34044), .B(n23947), .Z(n23949) );
  XOR U24671 ( .A(n34851), .B(n34510), .Z(n24234) );
  NANDN U24672 ( .A(n33867), .B(n24234), .Z(n23948) );
  AND U24673 ( .A(n23949), .B(n23948), .Z(n24293) );
  XNOR U24674 ( .A(n24292), .B(n24293), .Z(n24294) );
  XNOR U24675 ( .A(n24295), .B(n24294), .Z(n24322) );
  NANDN U24676 ( .A(n23951), .B(n23950), .Z(n23955) );
  NAND U24677 ( .A(n23953), .B(n23952), .Z(n23954) );
  NAND U24678 ( .A(n23955), .B(n23954), .Z(n24323) );
  XNOR U24679 ( .A(n24322), .B(n24323), .Z(n24324) );
  NAND U24680 ( .A(a[48]), .B(b[63]), .Z(n24364) );
  NANDN U24681 ( .A(n23956), .B(n38369), .Z(n23958) );
  XOR U24682 ( .A(b[61]), .B(n25134), .Z(n24243) );
  OR U24683 ( .A(n24243), .B(n38371), .Z(n23957) );
  NAND U24684 ( .A(n23958), .B(n23957), .Z(n24362) );
  NANDN U24685 ( .A(n23959), .B(n35311), .Z(n23961) );
  XOR U24686 ( .A(b[31]), .B(n32815), .Z(n24246) );
  NANDN U24687 ( .A(n24246), .B(n35313), .Z(n23960) );
  AND U24688 ( .A(n23961), .B(n23960), .Z(n24361) );
  XNOR U24689 ( .A(n24362), .B(n24361), .Z(n24363) );
  XNOR U24690 ( .A(n24364), .B(n24363), .Z(n24325) );
  XOR U24691 ( .A(n24324), .B(n24325), .Z(n24216) );
  XOR U24692 ( .A(b[37]), .B(n31363), .Z(n24249) );
  NANDN U24693 ( .A(n24249), .B(n36311), .Z(n23964) );
  NANDN U24694 ( .A(n23962), .B(n36309), .Z(n23963) );
  NAND U24695 ( .A(n23964), .B(n23963), .Z(n24307) );
  XOR U24696 ( .A(a[108]), .B(n968), .Z(n24252) );
  OR U24697 ( .A(n24252), .B(n29363), .Z(n23967) );
  NANDN U24698 ( .A(n23965), .B(n29864), .Z(n23966) );
  NAND U24699 ( .A(n23967), .B(n23966), .Z(n24304) );
  XOR U24700 ( .A(n37336), .B(n967), .Z(n24255) );
  NAND U24701 ( .A(n24255), .B(n28939), .Z(n23970) );
  NAND U24702 ( .A(n28938), .B(n23968), .Z(n23969) );
  AND U24703 ( .A(n23970), .B(n23969), .Z(n24305) );
  XNOR U24704 ( .A(n24304), .B(n24305), .Z(n24306) );
  XNOR U24705 ( .A(n24307), .B(n24306), .Z(n24210) );
  XOR U24706 ( .A(a[100]), .B(n971), .Z(n24258) );
  OR U24707 ( .A(n24258), .B(n31550), .Z(n23973) );
  NANDN U24708 ( .A(n23971), .B(n31874), .Z(n23972) );
  NAND U24709 ( .A(n23973), .B(n23972), .Z(n24394) );
  NAND U24710 ( .A(n34848), .B(n23974), .Z(n23976) );
  XOR U24711 ( .A(n35375), .B(n33628), .Z(n24261) );
  NAND U24712 ( .A(n34618), .B(n24261), .Z(n23975) );
  NAND U24713 ( .A(n23976), .B(n23975), .Z(n24391) );
  NAND U24714 ( .A(n35188), .B(n23977), .Z(n23979) );
  XOR U24715 ( .A(n35540), .B(n33185), .Z(n24264) );
  NANDN U24716 ( .A(n34968), .B(n24264), .Z(n23978) );
  AND U24717 ( .A(n23979), .B(n23978), .Z(n24392) );
  XNOR U24718 ( .A(n24391), .B(n24392), .Z(n24393) );
  XOR U24719 ( .A(n24394), .B(n24393), .Z(n24211) );
  XOR U24720 ( .A(n24210), .B(n24211), .Z(n24213) );
  NANDN U24721 ( .A(n23981), .B(n23980), .Z(n23985) );
  NAND U24722 ( .A(n23983), .B(n23982), .Z(n23984) );
  NAND U24723 ( .A(n23985), .B(n23984), .Z(n24212) );
  XOR U24724 ( .A(n24213), .B(n24212), .Z(n24217) );
  XNOR U24725 ( .A(n24216), .B(n24217), .Z(n24218) );
  XOR U24726 ( .A(n24219), .B(n24218), .Z(n24318) );
  NANDN U24727 ( .A(n23987), .B(n23986), .Z(n23991) );
  NANDN U24728 ( .A(n23989), .B(n23988), .Z(n23990) );
  NAND U24729 ( .A(n23991), .B(n23990), .Z(n24317) );
  NANDN U24730 ( .A(n23993), .B(n23992), .Z(n23997) );
  NAND U24731 ( .A(n23995), .B(n23994), .Z(n23996) );
  NAND U24732 ( .A(n23997), .B(n23996), .Z(n24207) );
  XOR U24733 ( .A(b[33]), .B(n32814), .Z(n24282) );
  NANDN U24734 ( .A(n24282), .B(n35620), .Z(n24000) );
  NANDN U24735 ( .A(n23998), .B(n35621), .Z(n23999) );
  NAND U24736 ( .A(n24000), .B(n23999), .Z(n24406) );
  NANDN U24737 ( .A(n966), .B(a[112]), .Z(n24001) );
  XOR U24738 ( .A(n29232), .B(n24001), .Z(n24003) );
  NANDN U24739 ( .A(b[0]), .B(a[111]), .Z(n24002) );
  AND U24740 ( .A(n24003), .B(n24002), .Z(n24403) );
  XOR U24741 ( .A(b[63]), .B(n24671), .Z(n24289) );
  NANDN U24742 ( .A(n24289), .B(n38422), .Z(n24006) );
  NANDN U24743 ( .A(n24004), .B(n38423), .Z(n24005) );
  AND U24744 ( .A(n24006), .B(n24005), .Z(n24404) );
  XNOR U24745 ( .A(n24403), .B(n24404), .Z(n24405) );
  XOR U24746 ( .A(n24406), .B(n24405), .Z(n24411) );
  XNOR U24747 ( .A(b[41]), .B(a[72]), .Z(n24273) );
  OR U24748 ( .A(n24273), .B(n36905), .Z(n24009) );
  NANDN U24749 ( .A(n24007), .B(n36807), .Z(n24008) );
  NAND U24750 ( .A(n24009), .B(n24008), .Z(n24301) );
  XOR U24751 ( .A(b[57]), .B(n25860), .Z(n24276) );
  OR U24752 ( .A(n24276), .B(n965), .Z(n24012) );
  NANDN U24753 ( .A(n24010), .B(n38194), .Z(n24011) );
  NAND U24754 ( .A(n24012), .B(n24011), .Z(n24298) );
  NAND U24755 ( .A(n38326), .B(n24013), .Z(n24015) );
  XOR U24756 ( .A(n38400), .B(n25177), .Z(n24279) );
  NANDN U24757 ( .A(n38273), .B(n24279), .Z(n24014) );
  AND U24758 ( .A(n24015), .B(n24014), .Z(n24299) );
  XNOR U24759 ( .A(n24298), .B(n24299), .Z(n24300) );
  XOR U24760 ( .A(n24301), .B(n24300), .Z(n24409) );
  NANDN U24761 ( .A(n24017), .B(n24016), .Z(n24021) );
  NAND U24762 ( .A(n24019), .B(n24018), .Z(n24020) );
  NAND U24763 ( .A(n24021), .B(n24020), .Z(n24410) );
  XNOR U24764 ( .A(n24409), .B(n24410), .Z(n24412) );
  XNOR U24765 ( .A(n24411), .B(n24412), .Z(n24205) );
  NANDN U24766 ( .A(n24023), .B(n24022), .Z(n24027) );
  NAND U24767 ( .A(n24025), .B(n24024), .Z(n24026) );
  AND U24768 ( .A(n24027), .B(n24026), .Z(n24204) );
  XNOR U24769 ( .A(n24205), .B(n24204), .Z(n24206) );
  XNOR U24770 ( .A(n24207), .B(n24206), .Z(n24316) );
  XNOR U24771 ( .A(n24317), .B(n24316), .Z(n24319) );
  XNOR U24772 ( .A(n24318), .B(n24319), .Z(n24423) );
  XOR U24773 ( .A(n24424), .B(n24423), .Z(n24186) );
  NAND U24774 ( .A(n24029), .B(n24028), .Z(n24033) );
  NANDN U24775 ( .A(n24031), .B(n24030), .Z(n24032) );
  NAND U24776 ( .A(n24033), .B(n24032), .Z(n24430) );
  NANDN U24777 ( .A(n24035), .B(n24034), .Z(n24039) );
  NAND U24778 ( .A(n24037), .B(n24036), .Z(n24038) );
  NAND U24779 ( .A(n24039), .B(n24038), .Z(n24446) );
  NANDN U24780 ( .A(n24041), .B(n24040), .Z(n24045) );
  OR U24781 ( .A(n24043), .B(n24042), .Z(n24044) );
  NAND U24782 ( .A(n24045), .B(n24044), .Z(n24443) );
  XOR U24783 ( .A(b[39]), .B(n31372), .Z(n24382) );
  NANDN U24784 ( .A(n24382), .B(n36553), .Z(n24048) );
  NANDN U24785 ( .A(n24046), .B(n36643), .Z(n24047) );
  NAND U24786 ( .A(n24048), .B(n24047), .Z(n24270) );
  XNOR U24787 ( .A(b[51]), .B(a[62]), .Z(n24385) );
  NANDN U24788 ( .A(n24385), .B(n37803), .Z(n24051) );
  NANDN U24789 ( .A(n24049), .B(n37802), .Z(n24050) );
  NAND U24790 ( .A(n24051), .B(n24050), .Z(n24267) );
  XOR U24791 ( .A(b[53]), .B(n27436), .Z(n24388) );
  NANDN U24792 ( .A(n24388), .B(n37940), .Z(n24054) );
  NANDN U24793 ( .A(n24052), .B(n37941), .Z(n24053) );
  AND U24794 ( .A(n24054), .B(n24053), .Z(n24268) );
  XNOR U24795 ( .A(n24267), .B(n24268), .Z(n24269) );
  XNOR U24796 ( .A(n24270), .B(n24269), .Z(n24313) );
  XOR U24797 ( .A(a[98]), .B(n972), .Z(n24373) );
  OR U24798 ( .A(n24373), .B(n32010), .Z(n24057) );
  NANDN U24799 ( .A(n24055), .B(n32011), .Z(n24056) );
  NAND U24800 ( .A(n24057), .B(n24056), .Z(n24240) );
  XNOR U24801 ( .A(b[25]), .B(n34048), .Z(n24376) );
  NANDN U24802 ( .A(n34219), .B(n24376), .Z(n24060) );
  NAND U24803 ( .A(n34217), .B(n24058), .Z(n24059) );
  NAND U24804 ( .A(n24060), .B(n24059), .Z(n24237) );
  XNOR U24805 ( .A(a[96]), .B(b[17]), .Z(n24379) );
  NANDN U24806 ( .A(n24379), .B(n32543), .Z(n24063) );
  NANDN U24807 ( .A(n24061), .B(n32541), .Z(n24062) );
  AND U24808 ( .A(n24063), .B(n24062), .Z(n24238) );
  XNOR U24809 ( .A(n24237), .B(n24238), .Z(n24239) );
  XNOR U24810 ( .A(n24240), .B(n24239), .Z(n24310) );
  NANDN U24811 ( .A(n24065), .B(n24064), .Z(n24069) );
  NAND U24812 ( .A(n24067), .B(n24066), .Z(n24068) );
  NAND U24813 ( .A(n24069), .B(n24068), .Z(n24311) );
  XNOR U24814 ( .A(n24310), .B(n24311), .Z(n24312) );
  XOR U24815 ( .A(n24313), .B(n24312), .Z(n24418) );
  NANDN U24816 ( .A(n24071), .B(n24070), .Z(n24075) );
  NAND U24817 ( .A(n24073), .B(n24072), .Z(n24074) );
  NAND U24818 ( .A(n24075), .B(n24074), .Z(n24415) );
  XNOR U24819 ( .A(n24415), .B(n24416), .Z(n24417) );
  XOR U24820 ( .A(n24418), .B(n24417), .Z(n24444) );
  XOR U24821 ( .A(n24443), .B(n24444), .Z(n24445) );
  XNOR U24822 ( .A(n24446), .B(n24445), .Z(n24427) );
  XNOR U24823 ( .A(b[35]), .B(a[78]), .Z(n24352) );
  NANDN U24824 ( .A(n24352), .B(n35985), .Z(n24082) );
  NAND U24825 ( .A(n24080), .B(n35986), .Z(n24081) );
  NAND U24826 ( .A(n24082), .B(n24081), .Z(n24400) );
  XOR U24827 ( .A(n36909), .B(n31123), .Z(n24355) );
  NAND U24828 ( .A(n24355), .B(n29949), .Z(n24085) );
  NAND U24829 ( .A(n29948), .B(n24083), .Z(n24084) );
  NAND U24830 ( .A(n24085), .B(n24084), .Z(n24397) );
  XOR U24831 ( .A(b[55]), .B(n26347), .Z(n24358) );
  NANDN U24832 ( .A(n24358), .B(n38075), .Z(n24088) );
  NANDN U24833 ( .A(n24086), .B(n38073), .Z(n24087) );
  AND U24834 ( .A(n24088), .B(n24087), .Z(n24398) );
  XNOR U24835 ( .A(n24397), .B(n24398), .Z(n24399) );
  XNOR U24836 ( .A(n24400), .B(n24399), .Z(n24201) );
  NANDN U24837 ( .A(n24090), .B(n24089), .Z(n24094) );
  NAND U24838 ( .A(n24092), .B(n24091), .Z(n24093) );
  NAND U24839 ( .A(n24094), .B(n24093), .Z(n24198) );
  OR U24840 ( .A(n24096), .B(n24095), .Z(n24100) );
  NANDN U24841 ( .A(n24098), .B(n24097), .Z(n24099) );
  NAND U24842 ( .A(n24100), .B(n24099), .Z(n24199) );
  XNOR U24843 ( .A(n24198), .B(n24199), .Z(n24200) );
  XOR U24844 ( .A(n24201), .B(n24200), .Z(n24435) );
  OR U24845 ( .A(n24102), .B(n24101), .Z(n24106) );
  OR U24846 ( .A(n24104), .B(n24103), .Z(n24105) );
  NAND U24847 ( .A(n24106), .B(n24105), .Z(n24433) );
  XNOR U24848 ( .A(b[49]), .B(a[64]), .Z(n24337) );
  OR U24849 ( .A(n24337), .B(n37756), .Z(n24109) );
  NANDN U24850 ( .A(n24107), .B(n37652), .Z(n24108) );
  NAND U24851 ( .A(n24109), .B(n24108), .Z(n24369) );
  NAND U24852 ( .A(n37469), .B(n24110), .Z(n24112) );
  XOR U24853 ( .A(n978), .B(n28701), .Z(n24340) );
  NAND U24854 ( .A(n24340), .B(n37471), .Z(n24111) );
  AND U24855 ( .A(n24112), .B(n24111), .Z(n24367) );
  XOR U24856 ( .A(a[104]), .B(n969), .Z(n24343) );
  NANDN U24857 ( .A(n24343), .B(n30509), .Z(n24115) );
  NANDN U24858 ( .A(n24113), .B(n30846), .Z(n24114) );
  AND U24859 ( .A(n24115), .B(n24114), .Z(n24368) );
  XOR U24860 ( .A(n24369), .B(n24370), .Z(n24222) );
  XOR U24861 ( .A(a[102]), .B(n970), .Z(n24328) );
  OR U24862 ( .A(n24328), .B(n31369), .Z(n24118) );
  NANDN U24863 ( .A(n24116), .B(n31119), .Z(n24117) );
  NAND U24864 ( .A(n24118), .B(n24117), .Z(n24349) );
  XOR U24865 ( .A(b[43]), .B(n30379), .Z(n24331) );
  NANDN U24866 ( .A(n24331), .B(n37068), .Z(n24121) );
  NANDN U24867 ( .A(n24119), .B(n37069), .Z(n24120) );
  NAND U24868 ( .A(n24121), .B(n24120), .Z(n24346) );
  XNOR U24869 ( .A(b[45]), .B(a[68]), .Z(n24334) );
  NANDN U24870 ( .A(n24334), .B(n37261), .Z(n24124) );
  NANDN U24871 ( .A(n24122), .B(n37262), .Z(n24123) );
  AND U24872 ( .A(n24124), .B(n24123), .Z(n24347) );
  XNOR U24873 ( .A(n24346), .B(n24347), .Z(n24348) );
  XOR U24874 ( .A(n24349), .B(n24348), .Z(n24223) );
  XNOR U24875 ( .A(n24222), .B(n24223), .Z(n24224) );
  NANDN U24876 ( .A(n24126), .B(n24125), .Z(n24130) );
  NAND U24877 ( .A(n24128), .B(n24127), .Z(n24129) );
  AND U24878 ( .A(n24130), .B(n24129), .Z(n24225) );
  XNOR U24879 ( .A(n24224), .B(n24225), .Z(n24434) );
  XNOR U24880 ( .A(n24433), .B(n24434), .Z(n24436) );
  XNOR U24881 ( .A(n24435), .B(n24436), .Z(n24428) );
  XOR U24882 ( .A(n24430), .B(n24429), .Z(n24187) );
  XNOR U24883 ( .A(n24186), .B(n24187), .Z(n24188) );
  NAND U24884 ( .A(n24132), .B(n24131), .Z(n24136) );
  NANDN U24885 ( .A(n24134), .B(n24133), .Z(n24135) );
  NAND U24886 ( .A(n24136), .B(n24135), .Z(n24189) );
  XOR U24887 ( .A(n24188), .B(n24189), .Z(n24452) );
  NAND U24888 ( .A(n24138), .B(n24137), .Z(n24142) );
  NANDN U24889 ( .A(n24140), .B(n24139), .Z(n24141) );
  NAND U24890 ( .A(n24142), .B(n24141), .Z(n24195) );
  NANDN U24891 ( .A(n24144), .B(n24143), .Z(n24148) );
  NAND U24892 ( .A(n24146), .B(n24145), .Z(n24147) );
  NAND U24893 ( .A(n24148), .B(n24147), .Z(n24193) );
  XNOR U24894 ( .A(n24193), .B(n24192), .Z(n24194) );
  XOR U24895 ( .A(n24195), .B(n24194), .Z(n24449) );
  NANDN U24896 ( .A(n24154), .B(n24153), .Z(n24158) );
  NANDN U24897 ( .A(n24156), .B(n24155), .Z(n24157) );
  NAND U24898 ( .A(n24158), .B(n24157), .Z(n24450) );
  XNOR U24899 ( .A(n24449), .B(n24450), .Z(n24451) );
  XNOR U24900 ( .A(n24452), .B(n24451), .Z(n24458) );
  XOR U24901 ( .A(n24457), .B(n24458), .Z(n24461) );
  NANDN U24902 ( .A(n24160), .B(n24159), .Z(n24164) );
  NAND U24903 ( .A(n24162), .B(n24161), .Z(n24163) );
  NAND U24904 ( .A(n24164), .B(n24163), .Z(n24462) );
  XNOR U24905 ( .A(n24461), .B(n24462), .Z(n24463) );
  NANDN U24906 ( .A(n24166), .B(n24165), .Z(n24170) );
  NAND U24907 ( .A(n24168), .B(n24167), .Z(n24169) );
  NAND U24908 ( .A(n24170), .B(n24169), .Z(n24464) );
  XOR U24909 ( .A(n24463), .B(n24464), .Z(n24180) );
  XNOR U24910 ( .A(n24180), .B(n24181), .Z(n24182) );
  XNOR U24911 ( .A(n24183), .B(n24182), .Z(n24467) );
  XNOR U24912 ( .A(n24467), .B(sreg[176]), .Z(n24469) );
  NAND U24913 ( .A(n24175), .B(sreg[175]), .Z(n24179) );
  OR U24914 ( .A(n24177), .B(n24176), .Z(n24178) );
  AND U24915 ( .A(n24179), .B(n24178), .Z(n24468) );
  XOR U24916 ( .A(n24469), .B(n24468), .Z(c[176]) );
  NANDN U24917 ( .A(n24181), .B(n24180), .Z(n24185) );
  NAND U24918 ( .A(n24183), .B(n24182), .Z(n24184) );
  NAND U24919 ( .A(n24185), .B(n24184), .Z(n24475) );
  NANDN U24920 ( .A(n24187), .B(n24186), .Z(n24191) );
  NANDN U24921 ( .A(n24189), .B(n24188), .Z(n24190) );
  NAND U24922 ( .A(n24191), .B(n24190), .Z(n24748) );
  NANDN U24923 ( .A(n24193), .B(n24192), .Z(n24197) );
  NANDN U24924 ( .A(n24195), .B(n24194), .Z(n24196) );
  AND U24925 ( .A(n24197), .B(n24196), .Z(n24747) );
  XNOR U24926 ( .A(n24748), .B(n24747), .Z(n24749) );
  NANDN U24927 ( .A(n24199), .B(n24198), .Z(n24203) );
  NAND U24928 ( .A(n24201), .B(n24200), .Z(n24202) );
  NAND U24929 ( .A(n24203), .B(n24202), .Z(n24505) );
  NANDN U24930 ( .A(n24205), .B(n24204), .Z(n24209) );
  NANDN U24931 ( .A(n24207), .B(n24206), .Z(n24208) );
  AND U24932 ( .A(n24209), .B(n24208), .Z(n24502) );
  NANDN U24933 ( .A(n24211), .B(n24210), .Z(n24215) );
  OR U24934 ( .A(n24213), .B(n24212), .Z(n24214) );
  AND U24935 ( .A(n24215), .B(n24214), .Z(n24503) );
  XNOR U24936 ( .A(n24505), .B(n24504), .Z(n24736) );
  NANDN U24937 ( .A(n24217), .B(n24216), .Z(n24221) );
  NANDN U24938 ( .A(n24219), .B(n24218), .Z(n24220) );
  AND U24939 ( .A(n24221), .B(n24220), .Z(n24735) );
  XNOR U24940 ( .A(n24736), .B(n24735), .Z(n24737) );
  NANDN U24941 ( .A(n24223), .B(n24222), .Z(n24227) );
  NAND U24942 ( .A(n24225), .B(n24224), .Z(n24226) );
  NAND U24943 ( .A(n24227), .B(n24226), .Z(n24732) );
  NAND U24944 ( .A(n33283), .B(n24228), .Z(n24230) );
  XOR U24945 ( .A(n35628), .B(n33020), .Z(n24678) );
  NANDN U24946 ( .A(n33021), .B(n24678), .Z(n24229) );
  NAND U24947 ( .A(n24230), .B(n24229), .Z(n24708) );
  XNOR U24948 ( .A(a[93]), .B(b[21]), .Z(n24681) );
  OR U24949 ( .A(n24681), .B(n33634), .Z(n24233) );
  NANDN U24950 ( .A(n24231), .B(n33464), .Z(n24232) );
  NAND U24951 ( .A(n24233), .B(n24232), .Z(n24705) );
  NAND U24952 ( .A(n34044), .B(n24234), .Z(n24236) );
  XNOR U24953 ( .A(a[91]), .B(n34510), .Z(n24684) );
  NANDN U24954 ( .A(n33867), .B(n24684), .Z(n24235) );
  AND U24955 ( .A(n24236), .B(n24235), .Z(n24706) );
  XNOR U24956 ( .A(n24705), .B(n24706), .Z(n24707) );
  XNOR U24957 ( .A(n24708), .B(n24707), .Z(n24589) );
  NANDN U24958 ( .A(n24238), .B(n24237), .Z(n24242) );
  NAND U24959 ( .A(n24240), .B(n24239), .Z(n24241) );
  NAND U24960 ( .A(n24242), .B(n24241), .Z(n24590) );
  XNOR U24961 ( .A(n24589), .B(n24590), .Z(n24591) );
  NAND U24962 ( .A(a[49]), .B(b[63]), .Z(n24580) );
  NANDN U24963 ( .A(n24243), .B(n38369), .Z(n24245) );
  XOR U24964 ( .A(b[61]), .B(n25001), .Z(n24672) );
  OR U24965 ( .A(n24672), .B(n38371), .Z(n24244) );
  NAND U24966 ( .A(n24245), .B(n24244), .Z(n24578) );
  NANDN U24967 ( .A(n24246), .B(n35311), .Z(n24248) );
  XNOR U24968 ( .A(b[31]), .B(a[83]), .Z(n24675) );
  NANDN U24969 ( .A(n24675), .B(n35313), .Z(n24247) );
  AND U24970 ( .A(n24248), .B(n24247), .Z(n24577) );
  XNOR U24971 ( .A(n24578), .B(n24577), .Z(n24579) );
  XNOR U24972 ( .A(n24580), .B(n24579), .Z(n24592) );
  XOR U24973 ( .A(n24591), .B(n24592), .Z(n24729) );
  XNOR U24974 ( .A(b[37]), .B(a[77]), .Z(n24641) );
  NANDN U24975 ( .A(n24641), .B(n36311), .Z(n24251) );
  NANDN U24976 ( .A(n24249), .B(n36309), .Z(n24250) );
  NAND U24977 ( .A(n24251), .B(n24250), .Z(n24720) );
  XNOR U24978 ( .A(a[109]), .B(b[5]), .Z(n24644) );
  OR U24979 ( .A(n24644), .B(n29363), .Z(n24254) );
  NANDN U24980 ( .A(n24252), .B(n29864), .Z(n24253) );
  NAND U24981 ( .A(n24254), .B(n24253), .Z(n24717) );
  XNOR U24982 ( .A(a[111]), .B(n967), .Z(n24647) );
  NAND U24983 ( .A(n24647), .B(n28939), .Z(n24257) );
  NAND U24984 ( .A(n28938), .B(n24255), .Z(n24256) );
  AND U24985 ( .A(n24257), .B(n24256), .Z(n24718) );
  XNOR U24986 ( .A(n24717), .B(n24718), .Z(n24719) );
  XNOR U24987 ( .A(n24720), .B(n24719), .Z(n24621) );
  XNOR U24988 ( .A(a[101]), .B(b[13]), .Z(n24650) );
  OR U24989 ( .A(n24650), .B(n31550), .Z(n24260) );
  NANDN U24990 ( .A(n24258), .B(n31874), .Z(n24259) );
  NAND U24991 ( .A(n24260), .B(n24259), .Z(n24541) );
  NAND U24992 ( .A(n34848), .B(n24261), .Z(n24263) );
  XNOR U24993 ( .A(n35375), .B(a[87]), .Z(n24653) );
  NAND U24994 ( .A(n34618), .B(n24653), .Z(n24262) );
  NAND U24995 ( .A(n24263), .B(n24262), .Z(n24538) );
  NAND U24996 ( .A(n35188), .B(n24264), .Z(n24266) );
  XNOR U24997 ( .A(n35540), .B(a[85]), .Z(n24656) );
  NANDN U24998 ( .A(n34968), .B(n24656), .Z(n24265) );
  AND U24999 ( .A(n24266), .B(n24265), .Z(n24539) );
  XNOR U25000 ( .A(n24538), .B(n24539), .Z(n24540) );
  XNOR U25001 ( .A(n24541), .B(n24540), .Z(n24619) );
  NANDN U25002 ( .A(n24268), .B(n24267), .Z(n24272) );
  NAND U25003 ( .A(n24270), .B(n24269), .Z(n24271) );
  NAND U25004 ( .A(n24272), .B(n24271), .Z(n24620) );
  XOR U25005 ( .A(n24619), .B(n24620), .Z(n24622) );
  XNOR U25006 ( .A(n24621), .B(n24622), .Z(n24730) );
  XNOR U25007 ( .A(n24729), .B(n24730), .Z(n24731) );
  XOR U25008 ( .A(n24732), .B(n24731), .Z(n24517) );
  XOR U25009 ( .A(b[41]), .B(a[73]), .Z(n24696) );
  NANDN U25010 ( .A(n36905), .B(n24696), .Z(n24275) );
  NANDN U25011 ( .A(n24273), .B(n36807), .Z(n24274) );
  NAND U25012 ( .A(n24275), .B(n24274), .Z(n24714) );
  XOR U25013 ( .A(b[57]), .B(n26122), .Z(n24699) );
  OR U25014 ( .A(n24699), .B(n965), .Z(n24278) );
  NANDN U25015 ( .A(n24276), .B(n38194), .Z(n24277) );
  NAND U25016 ( .A(n24278), .B(n24277), .Z(n24711) );
  NAND U25017 ( .A(n38326), .B(n24279), .Z(n24281) );
  XOR U25018 ( .A(n38400), .B(n25466), .Z(n24702) );
  NANDN U25019 ( .A(n38273), .B(n24702), .Z(n24280) );
  AND U25020 ( .A(n24281), .B(n24280), .Z(n24712) );
  XNOR U25021 ( .A(n24711), .B(n24712), .Z(n24713) );
  XNOR U25022 ( .A(n24714), .B(n24713), .Z(n24556) );
  XNOR U25023 ( .A(b[33]), .B(a[81]), .Z(n24687) );
  NANDN U25024 ( .A(n24687), .B(n35620), .Z(n24284) );
  NANDN U25025 ( .A(n24282), .B(n35621), .Z(n24283) );
  NAND U25026 ( .A(n24284), .B(n24283), .Z(n24553) );
  NANDN U25027 ( .A(n966), .B(a[113]), .Z(n24285) );
  XOR U25028 ( .A(n29232), .B(n24285), .Z(n24287) );
  IV U25029 ( .A(a[112]), .Z(n37583) );
  NANDN U25030 ( .A(n37583), .B(n966), .Z(n24286) );
  AND U25031 ( .A(n24287), .B(n24286), .Z(n24550) );
  XOR U25032 ( .A(b[63]), .B(n24288), .Z(n24693) );
  NANDN U25033 ( .A(n24693), .B(n38422), .Z(n24291) );
  NANDN U25034 ( .A(n24289), .B(n38423), .Z(n24290) );
  AND U25035 ( .A(n24291), .B(n24290), .Z(n24551) );
  XNOR U25036 ( .A(n24550), .B(n24551), .Z(n24552) );
  XOR U25037 ( .A(n24553), .B(n24552), .Z(n24557) );
  XNOR U25038 ( .A(n24556), .B(n24557), .Z(n24558) );
  NANDN U25039 ( .A(n24293), .B(n24292), .Z(n24297) );
  NAND U25040 ( .A(n24295), .B(n24294), .Z(n24296) );
  NAND U25041 ( .A(n24297), .B(n24296), .Z(n24559) );
  XOR U25042 ( .A(n24558), .B(n24559), .Z(n24634) );
  NANDN U25043 ( .A(n24299), .B(n24298), .Z(n24303) );
  NAND U25044 ( .A(n24301), .B(n24300), .Z(n24302) );
  NAND U25045 ( .A(n24303), .B(n24302), .Z(n24631) );
  NANDN U25046 ( .A(n24305), .B(n24304), .Z(n24309) );
  NAND U25047 ( .A(n24307), .B(n24306), .Z(n24308) );
  AND U25048 ( .A(n24309), .B(n24308), .Z(n24632) );
  XNOR U25049 ( .A(n24631), .B(n24632), .Z(n24633) );
  XNOR U25050 ( .A(n24634), .B(n24633), .Z(n24514) );
  NANDN U25051 ( .A(n24311), .B(n24310), .Z(n24315) );
  NAND U25052 ( .A(n24313), .B(n24312), .Z(n24314) );
  AND U25053 ( .A(n24315), .B(n24314), .Z(n24515) );
  XNOR U25054 ( .A(n24514), .B(n24515), .Z(n24516) );
  XNOR U25055 ( .A(n24517), .B(n24516), .Z(n24738) );
  XOR U25056 ( .A(n24737), .B(n24738), .Z(n24484) );
  NAND U25057 ( .A(n24317), .B(n24316), .Z(n24321) );
  NANDN U25058 ( .A(n24319), .B(n24318), .Z(n24320) );
  NAND U25059 ( .A(n24321), .B(n24320), .Z(n24493) );
  NANDN U25060 ( .A(n24323), .B(n24322), .Z(n24327) );
  NANDN U25061 ( .A(n24325), .B(n24324), .Z(n24326) );
  NAND U25062 ( .A(n24327), .B(n24326), .Z(n24497) );
  XNOR U25063 ( .A(a[103]), .B(b[11]), .Z(n24595) );
  OR U25064 ( .A(n24595), .B(n31369), .Z(n24330) );
  NANDN U25065 ( .A(n24328), .B(n31119), .Z(n24329) );
  NAND U25066 ( .A(n24330), .B(n24329), .Z(n24616) );
  XOR U25067 ( .A(b[43]), .B(n30543), .Z(n24598) );
  NANDN U25068 ( .A(n24598), .B(n37068), .Z(n24333) );
  NANDN U25069 ( .A(n24331), .B(n37069), .Z(n24332) );
  NAND U25070 ( .A(n24333), .B(n24332), .Z(n24613) );
  XOR U25071 ( .A(b[45]), .B(a[69]), .Z(n24601) );
  NAND U25072 ( .A(n24601), .B(n37261), .Z(n24336) );
  NANDN U25073 ( .A(n24334), .B(n37262), .Z(n24335) );
  AND U25074 ( .A(n24336), .B(n24335), .Z(n24614) );
  XNOR U25075 ( .A(n24613), .B(n24614), .Z(n24615) );
  XNOR U25076 ( .A(n24616), .B(n24615), .Z(n24640) );
  XOR U25077 ( .A(b[49]), .B(n28403), .Z(n24604) );
  OR U25078 ( .A(n24604), .B(n37756), .Z(n24339) );
  NANDN U25079 ( .A(n24337), .B(n37652), .Z(n24338) );
  NAND U25080 ( .A(n24339), .B(n24338), .Z(n24585) );
  NAND U25081 ( .A(n37469), .B(n24340), .Z(n24342) );
  XOR U25082 ( .A(n978), .B(n29372), .Z(n24607) );
  NAND U25083 ( .A(n24607), .B(n37471), .Z(n24341) );
  AND U25084 ( .A(n24342), .B(n24341), .Z(n24583) );
  XNOR U25085 ( .A(a[105]), .B(b[9]), .Z(n24610) );
  NANDN U25086 ( .A(n24610), .B(n30509), .Z(n24345) );
  NANDN U25087 ( .A(n24343), .B(n30846), .Z(n24344) );
  AND U25088 ( .A(n24345), .B(n24344), .Z(n24584) );
  XOR U25089 ( .A(n24585), .B(n24586), .Z(n24637) );
  NANDN U25090 ( .A(n24347), .B(n24346), .Z(n24351) );
  NAND U25091 ( .A(n24349), .B(n24348), .Z(n24350) );
  NAND U25092 ( .A(n24351), .B(n24350), .Z(n24638) );
  XNOR U25093 ( .A(n24637), .B(n24638), .Z(n24639) );
  XOR U25094 ( .A(n24640), .B(n24639), .Z(n24496) );
  XNOR U25095 ( .A(n24497), .B(n24496), .Z(n24499) );
  XOR U25096 ( .A(b[35]), .B(a[79]), .Z(n24568) );
  NAND U25097 ( .A(n35985), .B(n24568), .Z(n24354) );
  NANDN U25098 ( .A(n24352), .B(n35986), .Z(n24353) );
  NAND U25099 ( .A(n24354), .B(n24353), .Z(n24547) );
  XNOR U25100 ( .A(a[107]), .B(n31123), .Z(n24571) );
  NAND U25101 ( .A(n24571), .B(n29949), .Z(n24357) );
  NAND U25102 ( .A(n29948), .B(n24355), .Z(n24356) );
  NAND U25103 ( .A(n24357), .B(n24356), .Z(n24544) );
  XNOR U25104 ( .A(b[55]), .B(a[59]), .Z(n24574) );
  NANDN U25105 ( .A(n24574), .B(n38075), .Z(n24360) );
  NANDN U25106 ( .A(n24358), .B(n38073), .Z(n24359) );
  AND U25107 ( .A(n24360), .B(n24359), .Z(n24545) );
  XNOR U25108 ( .A(n24544), .B(n24545), .Z(n24546) );
  XNOR U25109 ( .A(n24547), .B(n24546), .Z(n24628) );
  NANDN U25110 ( .A(n24362), .B(n24361), .Z(n24366) );
  NAND U25111 ( .A(n24364), .B(n24363), .Z(n24365) );
  NAND U25112 ( .A(n24366), .B(n24365), .Z(n24625) );
  OR U25113 ( .A(n24368), .B(n24367), .Z(n24372) );
  NANDN U25114 ( .A(n24370), .B(n24369), .Z(n24371) );
  NAND U25115 ( .A(n24372), .B(n24371), .Z(n24626) );
  XNOR U25116 ( .A(n24625), .B(n24626), .Z(n24627) );
  XOR U25117 ( .A(n24628), .B(n24627), .Z(n24498) );
  XNOR U25118 ( .A(n24499), .B(n24498), .Z(n24491) );
  XNOR U25119 ( .A(a[99]), .B(b[15]), .Z(n24520) );
  OR U25120 ( .A(n24520), .B(n32010), .Z(n24375) );
  NANDN U25121 ( .A(n24373), .B(n32011), .Z(n24374) );
  NAND U25122 ( .A(n24375), .B(n24374), .Z(n24668) );
  XOR U25123 ( .A(b[25]), .B(a[89]), .Z(n24523) );
  NANDN U25124 ( .A(n34219), .B(n24523), .Z(n24378) );
  NAND U25125 ( .A(n34217), .B(n24376), .Z(n24377) );
  NAND U25126 ( .A(n24378), .B(n24377), .Z(n24665) );
  XOR U25127 ( .A(a[97]), .B(b[17]), .Z(n24526) );
  NAND U25128 ( .A(n24526), .B(n32543), .Z(n24381) );
  NANDN U25129 ( .A(n24379), .B(n32541), .Z(n24380) );
  AND U25130 ( .A(n24381), .B(n24380), .Z(n24666) );
  XNOR U25131 ( .A(n24665), .B(n24666), .Z(n24667) );
  XNOR U25132 ( .A(n24668), .B(n24667), .Z(n24723) );
  XNOR U25133 ( .A(b[39]), .B(a[75]), .Z(n24529) );
  NANDN U25134 ( .A(n24529), .B(n36553), .Z(n24384) );
  NANDN U25135 ( .A(n24382), .B(n36643), .Z(n24383) );
  NAND U25136 ( .A(n24384), .B(n24383), .Z(n24662) );
  XNOR U25137 ( .A(b[51]), .B(a[63]), .Z(n24532) );
  NANDN U25138 ( .A(n24532), .B(n37803), .Z(n24387) );
  NANDN U25139 ( .A(n24385), .B(n37802), .Z(n24386) );
  NAND U25140 ( .A(n24387), .B(n24386), .Z(n24659) );
  XOR U25141 ( .A(b[53]), .B(n27773), .Z(n24535) );
  NANDN U25142 ( .A(n24535), .B(n37940), .Z(n24390) );
  NANDN U25143 ( .A(n24388), .B(n37941), .Z(n24389) );
  AND U25144 ( .A(n24390), .B(n24389), .Z(n24660) );
  XNOR U25145 ( .A(n24659), .B(n24660), .Z(n24661) );
  XOR U25146 ( .A(n24662), .B(n24661), .Z(n24724) );
  XOR U25147 ( .A(n24723), .B(n24724), .Z(n24726) );
  NANDN U25148 ( .A(n24392), .B(n24391), .Z(n24396) );
  NAND U25149 ( .A(n24394), .B(n24393), .Z(n24395) );
  NAND U25150 ( .A(n24396), .B(n24395), .Z(n24725) );
  XNOR U25151 ( .A(n24726), .B(n24725), .Z(n24565) );
  NANDN U25152 ( .A(n24398), .B(n24397), .Z(n24402) );
  NAND U25153 ( .A(n24400), .B(n24399), .Z(n24401) );
  NAND U25154 ( .A(n24402), .B(n24401), .Z(n24562) );
  NANDN U25155 ( .A(n24404), .B(n24403), .Z(n24408) );
  NAND U25156 ( .A(n24406), .B(n24405), .Z(n24407) );
  AND U25157 ( .A(n24408), .B(n24407), .Z(n24563) );
  XNOR U25158 ( .A(n24562), .B(n24563), .Z(n24564) );
  XNOR U25159 ( .A(n24565), .B(n24564), .Z(n24511) );
  OR U25160 ( .A(n24410), .B(n24409), .Z(n24414) );
  OR U25161 ( .A(n24412), .B(n24411), .Z(n24413) );
  NAND U25162 ( .A(n24414), .B(n24413), .Z(n24508) );
  NANDN U25163 ( .A(n24416), .B(n24415), .Z(n24420) );
  NANDN U25164 ( .A(n24418), .B(n24417), .Z(n24419) );
  NAND U25165 ( .A(n24420), .B(n24419), .Z(n24509) );
  XNOR U25166 ( .A(n24508), .B(n24509), .Z(n24510) );
  XNOR U25167 ( .A(n24511), .B(n24510), .Z(n24490) );
  XOR U25168 ( .A(n24491), .B(n24490), .Z(n24492) );
  XNOR U25169 ( .A(n24493), .B(n24492), .Z(n24485) );
  XNOR U25170 ( .A(n24484), .B(n24485), .Z(n24486) );
  NAND U25171 ( .A(n24422), .B(n24421), .Z(n24426) );
  NANDN U25172 ( .A(n24424), .B(n24423), .Z(n24425) );
  NAND U25173 ( .A(n24426), .B(n24425), .Z(n24487) );
  XOR U25174 ( .A(n24486), .B(n24487), .Z(n24744) );
  NANDN U25175 ( .A(n24428), .B(n24427), .Z(n24432) );
  NAND U25176 ( .A(n24430), .B(n24429), .Z(n24431) );
  AND U25177 ( .A(n24432), .B(n24431), .Z(n24741) );
  NANDN U25178 ( .A(n24434), .B(n24433), .Z(n24438) );
  NAND U25179 ( .A(n24436), .B(n24435), .Z(n24437) );
  NAND U25180 ( .A(n24438), .B(n24437), .Z(n24481) );
  OR U25181 ( .A(n24444), .B(n24443), .Z(n24448) );
  NAND U25182 ( .A(n24446), .B(n24445), .Z(n24447) );
  NAND U25183 ( .A(n24448), .B(n24447), .Z(n24479) );
  XNOR U25184 ( .A(n24478), .B(n24479), .Z(n24480) );
  XNOR U25185 ( .A(n24481), .B(n24480), .Z(n24742) );
  XNOR U25186 ( .A(n24744), .B(n24743), .Z(n24750) );
  XOR U25187 ( .A(n24749), .B(n24750), .Z(n24753) );
  NANDN U25188 ( .A(n24450), .B(n24449), .Z(n24454) );
  NAND U25189 ( .A(n24452), .B(n24451), .Z(n24453) );
  NAND U25190 ( .A(n24454), .B(n24453), .Z(n24754) );
  XNOR U25191 ( .A(n24753), .B(n24754), .Z(n24755) );
  NANDN U25192 ( .A(n24456), .B(n24455), .Z(n24460) );
  NANDN U25193 ( .A(n24458), .B(n24457), .Z(n24459) );
  NAND U25194 ( .A(n24460), .B(n24459), .Z(n24756) );
  XOR U25195 ( .A(n24755), .B(n24756), .Z(n24472) );
  NANDN U25196 ( .A(n24462), .B(n24461), .Z(n24466) );
  NANDN U25197 ( .A(n24464), .B(n24463), .Z(n24465) );
  NAND U25198 ( .A(n24466), .B(n24465), .Z(n24473) );
  XNOR U25199 ( .A(n24472), .B(n24473), .Z(n24474) );
  XNOR U25200 ( .A(n24475), .B(n24474), .Z(n24759) );
  XNOR U25201 ( .A(n24759), .B(sreg[177]), .Z(n24761) );
  NAND U25202 ( .A(n24467), .B(sreg[176]), .Z(n24471) );
  OR U25203 ( .A(n24469), .B(n24468), .Z(n24470) );
  AND U25204 ( .A(n24471), .B(n24470), .Z(n24760) );
  XOR U25205 ( .A(n24761), .B(n24760), .Z(c[177]) );
  NANDN U25206 ( .A(n24473), .B(n24472), .Z(n24477) );
  NAND U25207 ( .A(n24475), .B(n24474), .Z(n24476) );
  NAND U25208 ( .A(n24477), .B(n24476), .Z(n24767) );
  NANDN U25209 ( .A(n24479), .B(n24478), .Z(n24483) );
  NAND U25210 ( .A(n24481), .B(n24480), .Z(n24482) );
  NAND U25211 ( .A(n24483), .B(n24482), .Z(n24768) );
  NANDN U25212 ( .A(n24485), .B(n24484), .Z(n24489) );
  NANDN U25213 ( .A(n24487), .B(n24486), .Z(n24488) );
  NAND U25214 ( .A(n24489), .B(n24488), .Z(n24769) );
  XNOR U25215 ( .A(n24768), .B(n24769), .Z(n24770) );
  NANDN U25216 ( .A(n24491), .B(n24490), .Z(n24495) );
  OR U25217 ( .A(n24493), .B(n24492), .Z(n24494) );
  NAND U25218 ( .A(n24495), .B(n24494), .Z(n24775) );
  NAND U25219 ( .A(n24497), .B(n24496), .Z(n24501) );
  NANDN U25220 ( .A(n24499), .B(n24498), .Z(n24500) );
  NAND U25221 ( .A(n24501), .B(n24500), .Z(n25030) );
  OR U25222 ( .A(n24503), .B(n24502), .Z(n24507) );
  NAND U25223 ( .A(n24505), .B(n24504), .Z(n24506) );
  NAND U25224 ( .A(n24507), .B(n24506), .Z(n25028) );
  NANDN U25225 ( .A(n24509), .B(n24508), .Z(n24513) );
  NAND U25226 ( .A(n24511), .B(n24510), .Z(n24512) );
  AND U25227 ( .A(n24513), .B(n24512), .Z(n25027) );
  XNOR U25228 ( .A(n25028), .B(n25027), .Z(n25029) );
  XNOR U25229 ( .A(n25030), .B(n25029), .Z(n24774) );
  XNOR U25230 ( .A(n24775), .B(n24774), .Z(n24777) );
  NANDN U25231 ( .A(n24515), .B(n24514), .Z(n24519) );
  NAND U25232 ( .A(n24517), .B(n24516), .Z(n24518) );
  NAND U25233 ( .A(n24519), .B(n24518), .Z(n24801) );
  XOR U25234 ( .A(a[100]), .B(n972), .Z(n24814) );
  OR U25235 ( .A(n24814), .B(n32010), .Z(n24522) );
  NANDN U25236 ( .A(n24520), .B(n32011), .Z(n24521) );
  NAND U25237 ( .A(n24522), .B(n24521), .Z(n24947) );
  XNOR U25238 ( .A(n34851), .B(b[25]), .Z(n24817) );
  NANDN U25239 ( .A(n34219), .B(n24817), .Z(n24525) );
  NAND U25240 ( .A(n34217), .B(n24523), .Z(n24524) );
  NAND U25241 ( .A(n24525), .B(n24524), .Z(n24944) );
  XNOR U25242 ( .A(a[98]), .B(b[17]), .Z(n24820) );
  NANDN U25243 ( .A(n24820), .B(n32543), .Z(n24528) );
  NAND U25244 ( .A(n24526), .B(n32541), .Z(n24527) );
  AND U25245 ( .A(n24528), .B(n24527), .Z(n24945) );
  XNOR U25246 ( .A(n24944), .B(n24945), .Z(n24946) );
  XNOR U25247 ( .A(n24947), .B(n24946), .Z(n25017) );
  XOR U25248 ( .A(b[39]), .B(n31363), .Z(n24823) );
  NANDN U25249 ( .A(n24823), .B(n36553), .Z(n24531) );
  NANDN U25250 ( .A(n24529), .B(n36643), .Z(n24530) );
  NAND U25251 ( .A(n24531), .B(n24530), .Z(n24977) );
  XNOR U25252 ( .A(b[51]), .B(a[64]), .Z(n24826) );
  NANDN U25253 ( .A(n24826), .B(n37803), .Z(n24534) );
  NANDN U25254 ( .A(n24532), .B(n37802), .Z(n24533) );
  NAND U25255 ( .A(n24534), .B(n24533), .Z(n24974) );
  XNOR U25256 ( .A(b[53]), .B(a[62]), .Z(n24829) );
  NANDN U25257 ( .A(n24829), .B(n37940), .Z(n24537) );
  NANDN U25258 ( .A(n24535), .B(n37941), .Z(n24536) );
  AND U25259 ( .A(n24537), .B(n24536), .Z(n24975) );
  XNOR U25260 ( .A(n24974), .B(n24975), .Z(n24976) );
  XOR U25261 ( .A(n24977), .B(n24976), .Z(n25018) );
  XOR U25262 ( .A(n25017), .B(n25018), .Z(n25020) );
  NANDN U25263 ( .A(n24539), .B(n24538), .Z(n24543) );
  NAND U25264 ( .A(n24541), .B(n24540), .Z(n24542) );
  NAND U25265 ( .A(n24543), .B(n24542), .Z(n25019) );
  XNOR U25266 ( .A(n25020), .B(n25019), .Z(n24851) );
  NANDN U25267 ( .A(n24545), .B(n24544), .Z(n24549) );
  NAND U25268 ( .A(n24547), .B(n24546), .Z(n24548) );
  NAND U25269 ( .A(n24549), .B(n24548), .Z(n24848) );
  NANDN U25270 ( .A(n24551), .B(n24550), .Z(n24555) );
  NAND U25271 ( .A(n24553), .B(n24552), .Z(n24554) );
  AND U25272 ( .A(n24555), .B(n24554), .Z(n24849) );
  XNOR U25273 ( .A(n24848), .B(n24849), .Z(n24850) );
  XNOR U25274 ( .A(n24851), .B(n24850), .Z(n24786) );
  NANDN U25275 ( .A(n24557), .B(n24556), .Z(n24561) );
  NANDN U25276 ( .A(n24559), .B(n24558), .Z(n24560) );
  AND U25277 ( .A(n24561), .B(n24560), .Z(n24787) );
  XNOR U25278 ( .A(n24786), .B(n24787), .Z(n24788) );
  NANDN U25279 ( .A(n24563), .B(n24562), .Z(n24567) );
  NAND U25280 ( .A(n24565), .B(n24564), .Z(n24566) );
  AND U25281 ( .A(n24567), .B(n24566), .Z(n24789) );
  XNOR U25282 ( .A(n24788), .B(n24789), .Z(n24799) );
  XNOR U25283 ( .A(b[35]), .B(a[80]), .Z(n24884) );
  NANDN U25284 ( .A(n24884), .B(n35985), .Z(n24570) );
  NAND U25285 ( .A(n24568), .B(n35986), .Z(n24569) );
  NAND U25286 ( .A(n24570), .B(n24569), .Z(n24841) );
  XOR U25287 ( .A(n37139), .B(n31123), .Z(n24887) );
  NAND U25288 ( .A(n24887), .B(n29949), .Z(n24573) );
  NAND U25289 ( .A(n29948), .B(n24571), .Z(n24572) );
  NAND U25290 ( .A(n24573), .B(n24572), .Z(n24838) );
  XOR U25291 ( .A(b[55]), .B(n27436), .Z(n24890) );
  NANDN U25292 ( .A(n24890), .B(n38075), .Z(n24576) );
  NANDN U25293 ( .A(n24574), .B(n38073), .Z(n24575) );
  AND U25294 ( .A(n24576), .B(n24575), .Z(n24839) );
  XNOR U25295 ( .A(n24838), .B(n24839), .Z(n24840) );
  XNOR U25296 ( .A(n24841), .B(n24840), .Z(n24914) );
  NANDN U25297 ( .A(n24578), .B(n24577), .Z(n24582) );
  NAND U25298 ( .A(n24580), .B(n24579), .Z(n24581) );
  NAND U25299 ( .A(n24582), .B(n24581), .Z(n24911) );
  OR U25300 ( .A(n24584), .B(n24583), .Z(n24588) );
  NANDN U25301 ( .A(n24586), .B(n24585), .Z(n24587) );
  NAND U25302 ( .A(n24588), .B(n24587), .Z(n24912) );
  XNOR U25303 ( .A(n24911), .B(n24912), .Z(n24913) );
  XOR U25304 ( .A(n24914), .B(n24913), .Z(n24782) );
  NANDN U25305 ( .A(n24590), .B(n24589), .Z(n24594) );
  NANDN U25306 ( .A(n24592), .B(n24591), .Z(n24593) );
  NAND U25307 ( .A(n24594), .B(n24593), .Z(n24780) );
  XOR U25308 ( .A(a[104]), .B(n970), .Z(n24854) );
  OR U25309 ( .A(n24854), .B(n31369), .Z(n24597) );
  NANDN U25310 ( .A(n24595), .B(n31119), .Z(n24596) );
  NAND U25311 ( .A(n24597), .B(n24596), .Z(n24875) );
  XOR U25312 ( .A(b[43]), .B(n30210), .Z(n24857) );
  NANDN U25313 ( .A(n24857), .B(n37068), .Z(n24600) );
  NANDN U25314 ( .A(n24598), .B(n37069), .Z(n24599) );
  NAND U25315 ( .A(n24600), .B(n24599), .Z(n24872) );
  XNOR U25316 ( .A(b[45]), .B(a[70]), .Z(n24860) );
  NANDN U25317 ( .A(n24860), .B(n37261), .Z(n24603) );
  NAND U25318 ( .A(n24601), .B(n37262), .Z(n24602) );
  AND U25319 ( .A(n24603), .B(n24602), .Z(n24873) );
  XNOR U25320 ( .A(n24872), .B(n24873), .Z(n24874) );
  XNOR U25321 ( .A(n24875), .B(n24874), .Z(n24929) );
  XOR U25322 ( .A(b[49]), .B(n28701), .Z(n24863) );
  OR U25323 ( .A(n24863), .B(n37756), .Z(n24606) );
  NANDN U25324 ( .A(n24604), .B(n37652), .Z(n24605) );
  NAND U25325 ( .A(n24606), .B(n24605), .Z(n24902) );
  NAND U25326 ( .A(n37469), .B(n24607), .Z(n24609) );
  XOR U25327 ( .A(n978), .B(n29868), .Z(n24866) );
  NAND U25328 ( .A(n24866), .B(n37471), .Z(n24608) );
  AND U25329 ( .A(n24609), .B(n24608), .Z(n24899) );
  XOR U25330 ( .A(a[106]), .B(n969), .Z(n24869) );
  NANDN U25331 ( .A(n24869), .B(n30509), .Z(n24612) );
  NANDN U25332 ( .A(n24610), .B(n30846), .Z(n24611) );
  AND U25333 ( .A(n24612), .B(n24611), .Z(n24900) );
  XOR U25334 ( .A(n24902), .B(n24901), .Z(n24930) );
  XNOR U25335 ( .A(n24929), .B(n24930), .Z(n24931) );
  NANDN U25336 ( .A(n24614), .B(n24613), .Z(n24618) );
  NAND U25337 ( .A(n24616), .B(n24615), .Z(n24617) );
  AND U25338 ( .A(n24618), .B(n24617), .Z(n24932) );
  XNOR U25339 ( .A(n24931), .B(n24932), .Z(n24781) );
  XNOR U25340 ( .A(n24780), .B(n24781), .Z(n24783) );
  XOR U25341 ( .A(n24782), .B(n24783), .Z(n24798) );
  XNOR U25342 ( .A(n24799), .B(n24798), .Z(n24800) );
  XNOR U25343 ( .A(n24801), .B(n24800), .Z(n25034) );
  NANDN U25344 ( .A(n24620), .B(n24619), .Z(n24624) );
  NANDN U25345 ( .A(n24622), .B(n24621), .Z(n24623) );
  NAND U25346 ( .A(n24624), .B(n24623), .Z(n24794) );
  NANDN U25347 ( .A(n24626), .B(n24625), .Z(n24630) );
  NAND U25348 ( .A(n24628), .B(n24627), .Z(n24629) );
  AND U25349 ( .A(n24630), .B(n24629), .Z(n24792) );
  NANDN U25350 ( .A(n24632), .B(n24631), .Z(n24636) );
  NAND U25351 ( .A(n24634), .B(n24633), .Z(n24635) );
  NAND U25352 ( .A(n24636), .B(n24635), .Z(n24793) );
  XOR U25353 ( .A(n24794), .B(n24795), .Z(n25026) );
  XOR U25354 ( .A(b[37]), .B(n31870), .Z(n24956) );
  NANDN U25355 ( .A(n24956), .B(n36311), .Z(n24643) );
  NANDN U25356 ( .A(n24641), .B(n36309), .Z(n24642) );
  NAND U25357 ( .A(n24643), .B(n24642), .Z(n25014) );
  XOR U25358 ( .A(a[110]), .B(n968), .Z(n24959) );
  OR U25359 ( .A(n24959), .B(n29363), .Z(n24646) );
  NANDN U25360 ( .A(n24644), .B(n29864), .Z(n24645) );
  NAND U25361 ( .A(n24646), .B(n24645), .Z(n25011) );
  XOR U25362 ( .A(n37583), .B(n967), .Z(n24962) );
  NAND U25363 ( .A(n24962), .B(n28939), .Z(n24649) );
  NAND U25364 ( .A(n28938), .B(n24647), .Z(n24648) );
  AND U25365 ( .A(n24649), .B(n24648), .Z(n25012) );
  XNOR U25366 ( .A(n25011), .B(n25012), .Z(n25013) );
  XNOR U25367 ( .A(n25014), .B(n25013), .Z(n24907) );
  XOR U25368 ( .A(a[102]), .B(n971), .Z(n24965) );
  OR U25369 ( .A(n24965), .B(n31550), .Z(n24652) );
  NANDN U25370 ( .A(n24650), .B(n31874), .Z(n24651) );
  NAND U25371 ( .A(n24652), .B(n24651), .Z(n24835) );
  NAND U25372 ( .A(n34848), .B(n24653), .Z(n24655) );
  XOR U25373 ( .A(n35375), .B(n34048), .Z(n24968) );
  NAND U25374 ( .A(n34618), .B(n24968), .Z(n24654) );
  NAND U25375 ( .A(n24655), .B(n24654), .Z(n24832) );
  NAND U25376 ( .A(n35188), .B(n24656), .Z(n24658) );
  XOR U25377 ( .A(n35540), .B(n33628), .Z(n24971) );
  NANDN U25378 ( .A(n34968), .B(n24971), .Z(n24657) );
  AND U25379 ( .A(n24658), .B(n24657), .Z(n24833) );
  XNOR U25380 ( .A(n24832), .B(n24833), .Z(n24834) );
  XNOR U25381 ( .A(n24835), .B(n24834), .Z(n24905) );
  NANDN U25382 ( .A(n24660), .B(n24659), .Z(n24664) );
  NAND U25383 ( .A(n24662), .B(n24661), .Z(n24663) );
  NAND U25384 ( .A(n24664), .B(n24663), .Z(n24906) );
  XOR U25385 ( .A(n24905), .B(n24906), .Z(n24908) );
  XNOR U25386 ( .A(n24907), .B(n24908), .Z(n24923) );
  NANDN U25387 ( .A(n24666), .B(n24665), .Z(n24670) );
  NAND U25388 ( .A(n24668), .B(n24667), .Z(n24669) );
  NAND U25389 ( .A(n24670), .B(n24669), .Z(n24880) );
  ANDN U25390 ( .B(b[63]), .A(n24671), .Z(n24896) );
  NANDN U25391 ( .A(n24672), .B(n38369), .Z(n24674) );
  XOR U25392 ( .A(b[61]), .B(n25177), .Z(n24950) );
  OR U25393 ( .A(n24950), .B(n38371), .Z(n24673) );
  NAND U25394 ( .A(n24674), .B(n24673), .Z(n24894) );
  NANDN U25395 ( .A(n24675), .B(n35311), .Z(n24677) );
  XOR U25396 ( .A(b[31]), .B(n33185), .Z(n24953) );
  NANDN U25397 ( .A(n24953), .B(n35313), .Z(n24676) );
  AND U25398 ( .A(n24677), .B(n24676), .Z(n24893) );
  XNOR U25399 ( .A(n24894), .B(n24893), .Z(n24895) );
  XOR U25400 ( .A(n24896), .B(n24895), .Z(n24878) );
  NAND U25401 ( .A(n33283), .B(n24678), .Z(n24680) );
  XOR U25402 ( .A(n35545), .B(n33020), .Z(n24935) );
  NANDN U25403 ( .A(n33021), .B(n24935), .Z(n24679) );
  NAND U25404 ( .A(n24680), .B(n24679), .Z(n24983) );
  XNOR U25405 ( .A(a[94]), .B(b[21]), .Z(n24938) );
  OR U25406 ( .A(n24938), .B(n33634), .Z(n24683) );
  NANDN U25407 ( .A(n24681), .B(n33464), .Z(n24682) );
  NAND U25408 ( .A(n24683), .B(n24682), .Z(n24980) );
  NAND U25409 ( .A(n34044), .B(n24684), .Z(n24686) );
  XOR U25410 ( .A(n34852), .B(n34510), .Z(n24941) );
  NANDN U25411 ( .A(n33867), .B(n24941), .Z(n24685) );
  AND U25412 ( .A(n24686), .B(n24685), .Z(n24981) );
  XNOR U25413 ( .A(n24980), .B(n24981), .Z(n24982) );
  XNOR U25414 ( .A(n24983), .B(n24982), .Z(n24879) );
  XOR U25415 ( .A(n24878), .B(n24879), .Z(n24881) );
  XOR U25416 ( .A(n24880), .B(n24881), .Z(n24924) );
  XOR U25417 ( .A(n24923), .B(n24924), .Z(n24925) );
  XOR U25418 ( .A(n24926), .B(n24925), .Z(n24805) );
  XOR U25419 ( .A(b[33]), .B(n32815), .Z(n24995) );
  NANDN U25420 ( .A(n24995), .B(n35620), .Z(n24689) );
  NANDN U25421 ( .A(n24687), .B(n35621), .Z(n24688) );
  NAND U25422 ( .A(n24689), .B(n24688), .Z(n24847) );
  NANDN U25423 ( .A(n966), .B(a[114]), .Z(n24690) );
  XOR U25424 ( .A(n29232), .B(n24690), .Z(n24692) );
  NANDN U25425 ( .A(b[0]), .B(a[113]), .Z(n24691) );
  AND U25426 ( .A(n24692), .B(n24691), .Z(n24844) );
  XOR U25427 ( .A(b[63]), .B(n25134), .Z(n25002) );
  NANDN U25428 ( .A(n25002), .B(n38422), .Z(n24695) );
  NANDN U25429 ( .A(n24693), .B(n38423), .Z(n24694) );
  AND U25430 ( .A(n24695), .B(n24694), .Z(n24845) );
  XNOR U25431 ( .A(n24844), .B(n24845), .Z(n24846) );
  XNOR U25432 ( .A(n24847), .B(n24846), .Z(n24810) );
  XNOR U25433 ( .A(b[41]), .B(a[74]), .Z(n24986) );
  OR U25434 ( .A(n24986), .B(n36905), .Z(n24698) );
  NAND U25435 ( .A(n24696), .B(n36807), .Z(n24697) );
  NAND U25436 ( .A(n24698), .B(n24697), .Z(n25008) );
  XOR U25437 ( .A(b[57]), .B(n26347), .Z(n24989) );
  OR U25438 ( .A(n24989), .B(n965), .Z(n24701) );
  NANDN U25439 ( .A(n24699), .B(n38194), .Z(n24700) );
  NAND U25440 ( .A(n24701), .B(n24700), .Z(n25005) );
  NAND U25441 ( .A(n38326), .B(n24702), .Z(n24704) );
  XOR U25442 ( .A(n38400), .B(n25860), .Z(n24992) );
  NANDN U25443 ( .A(n38273), .B(n24992), .Z(n24703) );
  AND U25444 ( .A(n24704), .B(n24703), .Z(n25006) );
  XNOR U25445 ( .A(n25005), .B(n25006), .Z(n25007) );
  XNOR U25446 ( .A(n25008), .B(n25007), .Z(n24808) );
  NANDN U25447 ( .A(n24706), .B(n24705), .Z(n24710) );
  NAND U25448 ( .A(n24708), .B(n24707), .Z(n24709) );
  NAND U25449 ( .A(n24710), .B(n24709), .Z(n24809) );
  XOR U25450 ( .A(n24808), .B(n24809), .Z(n24811) );
  XNOR U25451 ( .A(n24810), .B(n24811), .Z(n24920) );
  NANDN U25452 ( .A(n24712), .B(n24711), .Z(n24716) );
  NAND U25453 ( .A(n24714), .B(n24713), .Z(n24715) );
  NAND U25454 ( .A(n24716), .B(n24715), .Z(n24917) );
  NANDN U25455 ( .A(n24718), .B(n24717), .Z(n24722) );
  NAND U25456 ( .A(n24720), .B(n24719), .Z(n24721) );
  AND U25457 ( .A(n24722), .B(n24721), .Z(n24918) );
  XNOR U25458 ( .A(n24917), .B(n24918), .Z(n24919) );
  XNOR U25459 ( .A(n24920), .B(n24919), .Z(n24803) );
  NANDN U25460 ( .A(n24724), .B(n24723), .Z(n24728) );
  OR U25461 ( .A(n24726), .B(n24725), .Z(n24727) );
  AND U25462 ( .A(n24728), .B(n24727), .Z(n24802) );
  XOR U25463 ( .A(n24803), .B(n24802), .Z(n24804) );
  XNOR U25464 ( .A(n24805), .B(n24804), .Z(n25023) );
  NANDN U25465 ( .A(n24730), .B(n24729), .Z(n24734) );
  NANDN U25466 ( .A(n24732), .B(n24731), .Z(n24733) );
  AND U25467 ( .A(n24734), .B(n24733), .Z(n25024) );
  XNOR U25468 ( .A(n25023), .B(n25024), .Z(n25025) );
  XOR U25469 ( .A(n25026), .B(n25025), .Z(n25033) );
  XOR U25470 ( .A(n25034), .B(n25033), .Z(n25035) );
  NANDN U25471 ( .A(n24736), .B(n24735), .Z(n24740) );
  NANDN U25472 ( .A(n24738), .B(n24737), .Z(n24739) );
  AND U25473 ( .A(n24740), .B(n24739), .Z(n25036) );
  XOR U25474 ( .A(n25035), .B(n25036), .Z(n24776) );
  XNOR U25475 ( .A(n24777), .B(n24776), .Z(n24771) );
  XOR U25476 ( .A(n24770), .B(n24771), .Z(n25042) );
  OR U25477 ( .A(n24742), .B(n24741), .Z(n24746) );
  NAND U25478 ( .A(n24744), .B(n24743), .Z(n24745) );
  NAND U25479 ( .A(n24746), .B(n24745), .Z(n25040) );
  NANDN U25480 ( .A(n24748), .B(n24747), .Z(n24752) );
  NANDN U25481 ( .A(n24750), .B(n24749), .Z(n24751) );
  AND U25482 ( .A(n24752), .B(n24751), .Z(n25039) );
  XNOR U25483 ( .A(n25040), .B(n25039), .Z(n25041) );
  XNOR U25484 ( .A(n25042), .B(n25041), .Z(n24764) );
  NANDN U25485 ( .A(n24754), .B(n24753), .Z(n24758) );
  NANDN U25486 ( .A(n24756), .B(n24755), .Z(n24757) );
  NAND U25487 ( .A(n24758), .B(n24757), .Z(n24765) );
  XNOR U25488 ( .A(n24764), .B(n24765), .Z(n24766) );
  XNOR U25489 ( .A(n24767), .B(n24766), .Z(n25045) );
  XNOR U25490 ( .A(n25045), .B(sreg[178]), .Z(n25047) );
  NAND U25491 ( .A(n24759), .B(sreg[177]), .Z(n24763) );
  OR U25492 ( .A(n24761), .B(n24760), .Z(n24762) );
  AND U25493 ( .A(n24763), .B(n24762), .Z(n25046) );
  XOR U25494 ( .A(n25047), .B(n25046), .Z(c[178]) );
  NANDN U25495 ( .A(n24769), .B(n24768), .Z(n24773) );
  NANDN U25496 ( .A(n24771), .B(n24770), .Z(n24772) );
  NAND U25497 ( .A(n24773), .B(n24772), .Z(n25056) );
  OR U25498 ( .A(n24775), .B(n24774), .Z(n24779) );
  OR U25499 ( .A(n24777), .B(n24776), .Z(n24778) );
  AND U25500 ( .A(n24779), .B(n24778), .Z(n25057) );
  XNOR U25501 ( .A(n25056), .B(n25057), .Z(n25058) );
  NANDN U25502 ( .A(n24781), .B(n24780), .Z(n24785) );
  NAND U25503 ( .A(n24783), .B(n24782), .Z(n24784) );
  NAND U25504 ( .A(n24785), .B(n24784), .Z(n25333) );
  NANDN U25505 ( .A(n24787), .B(n24786), .Z(n24791) );
  NAND U25506 ( .A(n24789), .B(n24788), .Z(n24790) );
  NAND U25507 ( .A(n24791), .B(n24790), .Z(n25331) );
  OR U25508 ( .A(n24793), .B(n24792), .Z(n24797) );
  NANDN U25509 ( .A(n24795), .B(n24794), .Z(n24796) );
  AND U25510 ( .A(n24797), .B(n24796), .Z(n25330) );
  XNOR U25511 ( .A(n25331), .B(n25330), .Z(n25332) );
  XOR U25512 ( .A(n25333), .B(n25332), .Z(n25068) );
  XNOR U25513 ( .A(n25068), .B(n25069), .Z(n25070) );
  OR U25514 ( .A(n24803), .B(n24802), .Z(n24807) );
  NAND U25515 ( .A(n24805), .B(n24804), .Z(n24806) );
  NAND U25516 ( .A(n24807), .B(n24806), .Z(n25305) );
  NANDN U25517 ( .A(n24809), .B(n24808), .Z(n24813) );
  NANDN U25518 ( .A(n24811), .B(n24810), .Z(n24812) );
  NAND U25519 ( .A(n24813), .B(n24812), .Z(n25314) );
  XNOR U25520 ( .A(a[101]), .B(b[15]), .Z(n25254) );
  OR U25521 ( .A(n25254), .B(n32010), .Z(n24816) );
  NANDN U25522 ( .A(n24814), .B(n32011), .Z(n24815) );
  NAND U25523 ( .A(n24816), .B(n24815), .Z(n25131) );
  XOR U25524 ( .A(a[91]), .B(b[25]), .Z(n25257) );
  NANDN U25525 ( .A(n34219), .B(n25257), .Z(n24819) );
  NAND U25526 ( .A(n34217), .B(n24817), .Z(n24818) );
  NAND U25527 ( .A(n24819), .B(n24818), .Z(n25128) );
  XOR U25528 ( .A(a[99]), .B(b[17]), .Z(n25260) );
  NAND U25529 ( .A(n25260), .B(n32543), .Z(n24822) );
  NANDN U25530 ( .A(n24820), .B(n32541), .Z(n24821) );
  AND U25531 ( .A(n24822), .B(n24821), .Z(n25129) );
  XNOR U25532 ( .A(n25128), .B(n25129), .Z(n25130) );
  XNOR U25533 ( .A(n25131), .B(n25130), .Z(n25150) );
  XNOR U25534 ( .A(b[39]), .B(a[77]), .Z(n25263) );
  NANDN U25535 ( .A(n25263), .B(n36553), .Z(n24825) );
  NANDN U25536 ( .A(n24823), .B(n36643), .Z(n24824) );
  NAND U25537 ( .A(n24825), .B(n24824), .Z(n25125) );
  XOR U25538 ( .A(b[51]), .B(n28403), .Z(n25266) );
  NANDN U25539 ( .A(n25266), .B(n37803), .Z(n24828) );
  NANDN U25540 ( .A(n24826), .B(n37802), .Z(n24827) );
  NAND U25541 ( .A(n24828), .B(n24827), .Z(n25122) );
  XNOR U25542 ( .A(b[53]), .B(a[63]), .Z(n25269) );
  NANDN U25543 ( .A(n25269), .B(n37940), .Z(n24831) );
  NANDN U25544 ( .A(n24829), .B(n37941), .Z(n24830) );
  AND U25545 ( .A(n24831), .B(n24830), .Z(n25123) );
  XNOR U25546 ( .A(n25122), .B(n25123), .Z(n25124) );
  XOR U25547 ( .A(n25125), .B(n25124), .Z(n25151) );
  XOR U25548 ( .A(n25150), .B(n25151), .Z(n25153) );
  NANDN U25549 ( .A(n24833), .B(n24832), .Z(n24837) );
  NAND U25550 ( .A(n24835), .B(n24834), .Z(n24836) );
  NAND U25551 ( .A(n24837), .B(n24836), .Z(n25152) );
  XNOR U25552 ( .A(n25153), .B(n25152), .Z(n25299) );
  NANDN U25553 ( .A(n24839), .B(n24838), .Z(n24843) );
  NAND U25554 ( .A(n24841), .B(n24840), .Z(n24842) );
  NAND U25555 ( .A(n24843), .B(n24842), .Z(n25296) );
  XNOR U25556 ( .A(n25296), .B(n25297), .Z(n25298) );
  XOR U25557 ( .A(n25299), .B(n25298), .Z(n25315) );
  XNOR U25558 ( .A(n25314), .B(n25315), .Z(n25316) );
  NANDN U25559 ( .A(n24849), .B(n24848), .Z(n24853) );
  NAND U25560 ( .A(n24851), .B(n24850), .Z(n24852) );
  AND U25561 ( .A(n24853), .B(n24852), .Z(n25317) );
  XNOR U25562 ( .A(n25316), .B(n25317), .Z(n25303) );
  XNOR U25563 ( .A(a[105]), .B(b[11]), .Z(n25230) );
  OR U25564 ( .A(n25230), .B(n31369), .Z(n24856) );
  NANDN U25565 ( .A(n24854), .B(n31119), .Z(n24855) );
  NAND U25566 ( .A(n24856), .B(n24855), .Z(n25251) );
  XNOR U25567 ( .A(b[43]), .B(a[73]), .Z(n25233) );
  NANDN U25568 ( .A(n25233), .B(n37068), .Z(n24859) );
  NANDN U25569 ( .A(n24857), .B(n37069), .Z(n24858) );
  NAND U25570 ( .A(n24859), .B(n24858), .Z(n25248) );
  XNOR U25571 ( .A(b[45]), .B(a[71]), .Z(n25236) );
  NANDN U25572 ( .A(n25236), .B(n37261), .Z(n24862) );
  NANDN U25573 ( .A(n24860), .B(n37262), .Z(n24861) );
  AND U25574 ( .A(n24862), .B(n24861), .Z(n25249) );
  XNOR U25575 ( .A(n25248), .B(n25249), .Z(n25250) );
  XNOR U25576 ( .A(n25251), .B(n25250), .Z(n25098) );
  XOR U25577 ( .A(b[49]), .B(n29372), .Z(n25239) );
  OR U25578 ( .A(n25239), .B(n37756), .Z(n24865) );
  NANDN U25579 ( .A(n24863), .B(n37652), .Z(n24864) );
  NAND U25580 ( .A(n24865), .B(n24864), .Z(n25221) );
  NAND U25581 ( .A(n37469), .B(n24866), .Z(n24868) );
  XNOR U25582 ( .A(n978), .B(a[69]), .Z(n25242) );
  NAND U25583 ( .A(n25242), .B(n37471), .Z(n24867) );
  NAND U25584 ( .A(n24868), .B(n24867), .Z(n25218) );
  XNOR U25585 ( .A(a[107]), .B(b[9]), .Z(n25245) );
  NANDN U25586 ( .A(n25245), .B(n30509), .Z(n24871) );
  NANDN U25587 ( .A(n24869), .B(n30846), .Z(n24870) );
  AND U25588 ( .A(n24871), .B(n24870), .Z(n25219) );
  XNOR U25589 ( .A(n25218), .B(n25219), .Z(n25220) );
  XOR U25590 ( .A(n25221), .B(n25220), .Z(n25099) );
  XNOR U25591 ( .A(n25098), .B(n25099), .Z(n25100) );
  NANDN U25592 ( .A(n24873), .B(n24872), .Z(n24877) );
  NAND U25593 ( .A(n24875), .B(n24874), .Z(n24876) );
  AND U25594 ( .A(n24877), .B(n24876), .Z(n25101) );
  XNOR U25595 ( .A(n25100), .B(n25101), .Z(n25309) );
  NANDN U25596 ( .A(n24879), .B(n24878), .Z(n24883) );
  NANDN U25597 ( .A(n24881), .B(n24880), .Z(n24882) );
  AND U25598 ( .A(n24883), .B(n24882), .Z(n25308) );
  XNOR U25599 ( .A(n25309), .B(n25308), .Z(n25310) );
  XOR U25600 ( .A(b[35]), .B(a[81]), .Z(n25203) );
  NAND U25601 ( .A(n35985), .B(n25203), .Z(n24886) );
  NANDN U25602 ( .A(n24884), .B(n35986), .Z(n24885) );
  NAND U25603 ( .A(n24886), .B(n24885), .Z(n25281) );
  XNOR U25604 ( .A(a[109]), .B(n31123), .Z(n25206) );
  NAND U25605 ( .A(n25206), .B(n29949), .Z(n24889) );
  NAND U25606 ( .A(n29948), .B(n24887), .Z(n24888) );
  NAND U25607 ( .A(n24889), .B(n24888), .Z(n25278) );
  XOR U25608 ( .A(b[55]), .B(n27773), .Z(n25209) );
  NANDN U25609 ( .A(n25209), .B(n38075), .Z(n24892) );
  NANDN U25610 ( .A(n24890), .B(n38073), .Z(n24891) );
  AND U25611 ( .A(n24892), .B(n24891), .Z(n25279) );
  XNOR U25612 ( .A(n25278), .B(n25279), .Z(n25280) );
  XNOR U25613 ( .A(n25281), .B(n25280), .Z(n25089) );
  NANDN U25614 ( .A(n24894), .B(n24893), .Z(n24898) );
  NANDN U25615 ( .A(n24896), .B(n24895), .Z(n24897) );
  NAND U25616 ( .A(n24898), .B(n24897), .Z(n25086) );
  OR U25617 ( .A(n24900), .B(n24899), .Z(n24904) );
  NAND U25618 ( .A(n24902), .B(n24901), .Z(n24903) );
  NAND U25619 ( .A(n24904), .B(n24903), .Z(n25087) );
  XNOR U25620 ( .A(n25086), .B(n25087), .Z(n25088) );
  XOR U25621 ( .A(n25089), .B(n25088), .Z(n25311) );
  XOR U25622 ( .A(n25310), .B(n25311), .Z(n25302) );
  XNOR U25623 ( .A(n25303), .B(n25302), .Z(n25304) );
  XNOR U25624 ( .A(n25305), .B(n25304), .Z(n25327) );
  NANDN U25625 ( .A(n24906), .B(n24905), .Z(n24910) );
  NANDN U25626 ( .A(n24908), .B(n24907), .Z(n24909) );
  NAND U25627 ( .A(n24910), .B(n24909), .Z(n25323) );
  NANDN U25628 ( .A(n24912), .B(n24911), .Z(n24916) );
  NAND U25629 ( .A(n24914), .B(n24913), .Z(n24915) );
  AND U25630 ( .A(n24916), .B(n24915), .Z(n25320) );
  NANDN U25631 ( .A(n24918), .B(n24917), .Z(n24922) );
  NANDN U25632 ( .A(n24920), .B(n24919), .Z(n24921) );
  NAND U25633 ( .A(n24922), .B(n24921), .Z(n25321) );
  XNOR U25634 ( .A(n25323), .B(n25322), .Z(n25075) );
  OR U25635 ( .A(n24924), .B(n24923), .Z(n24928) );
  NANDN U25636 ( .A(n24926), .B(n24925), .Z(n24927) );
  AND U25637 ( .A(n24928), .B(n24927), .Z(n25074) );
  XNOR U25638 ( .A(n25075), .B(n25074), .Z(n25076) );
  NANDN U25639 ( .A(n24930), .B(n24929), .Z(n24934) );
  NAND U25640 ( .A(n24932), .B(n24931), .Z(n24933) );
  NAND U25641 ( .A(n24934), .B(n24933), .Z(n25196) );
  NAND U25642 ( .A(n33283), .B(n24935), .Z(n24937) );
  XNOR U25643 ( .A(a[97]), .B(n33020), .Z(n25141) );
  NANDN U25644 ( .A(n33021), .B(n25141), .Z(n24936) );
  NAND U25645 ( .A(n24937), .B(n24936), .Z(n25184) );
  XNOR U25646 ( .A(a[95]), .B(b[21]), .Z(n25144) );
  OR U25647 ( .A(n25144), .B(n33634), .Z(n24940) );
  NANDN U25648 ( .A(n24938), .B(n33464), .Z(n24939) );
  NAND U25649 ( .A(n24940), .B(n24939), .Z(n25181) );
  NAND U25650 ( .A(n34044), .B(n24941), .Z(n24943) );
  XOR U25651 ( .A(n35377), .B(n34510), .Z(n25147) );
  NANDN U25652 ( .A(n33867), .B(n25147), .Z(n24942) );
  AND U25653 ( .A(n24943), .B(n24942), .Z(n25182) );
  XNOR U25654 ( .A(n25181), .B(n25182), .Z(n25183) );
  XNOR U25655 ( .A(n25184), .B(n25183), .Z(n25224) );
  NANDN U25656 ( .A(n24945), .B(n24944), .Z(n24949) );
  NAND U25657 ( .A(n24947), .B(n24946), .Z(n24948) );
  NAND U25658 ( .A(n24949), .B(n24948), .Z(n25225) );
  XNOR U25659 ( .A(n25224), .B(n25225), .Z(n25226) );
  NAND U25660 ( .A(a[51]), .B(b[63]), .Z(n25215) );
  NANDN U25661 ( .A(n24950), .B(n38369), .Z(n24952) );
  XOR U25662 ( .A(b[61]), .B(n25466), .Z(n25135) );
  OR U25663 ( .A(n25135), .B(n38371), .Z(n24951) );
  NAND U25664 ( .A(n24952), .B(n24951), .Z(n25213) );
  NANDN U25665 ( .A(n24953), .B(n35311), .Z(n24955) );
  XNOR U25666 ( .A(b[31]), .B(a[85]), .Z(n25138) );
  NANDN U25667 ( .A(n25138), .B(n35313), .Z(n24954) );
  AND U25668 ( .A(n24955), .B(n24954), .Z(n25212) );
  XNOR U25669 ( .A(n25213), .B(n25212), .Z(n25214) );
  XNOR U25670 ( .A(n25215), .B(n25214), .Z(n25227) );
  XOR U25671 ( .A(n25226), .B(n25227), .Z(n25193) );
  XNOR U25672 ( .A(b[37]), .B(a[79]), .Z(n25104) );
  NANDN U25673 ( .A(n25104), .B(n36311), .Z(n24958) );
  NANDN U25674 ( .A(n24956), .B(n36309), .Z(n24957) );
  NAND U25675 ( .A(n24958), .B(n24957), .Z(n25159) );
  XNOR U25676 ( .A(a[111]), .B(b[5]), .Z(n25107) );
  OR U25677 ( .A(n25107), .B(n29363), .Z(n24961) );
  NANDN U25678 ( .A(n24959), .B(n29864), .Z(n24960) );
  NAND U25679 ( .A(n24961), .B(n24960), .Z(n25156) );
  XNOR U25680 ( .A(a[113]), .B(n967), .Z(n25110) );
  NAND U25681 ( .A(n25110), .B(n28939), .Z(n24964) );
  NAND U25682 ( .A(n28938), .B(n24962), .Z(n24963) );
  AND U25683 ( .A(n24964), .B(n24963), .Z(n25157) );
  XNOR U25684 ( .A(n25156), .B(n25157), .Z(n25158) );
  XNOR U25685 ( .A(n25159), .B(n25158), .Z(n25082) );
  XNOR U25686 ( .A(a[103]), .B(b[13]), .Z(n25113) );
  OR U25687 ( .A(n25113), .B(n31550), .Z(n24967) );
  NANDN U25688 ( .A(n24965), .B(n31874), .Z(n24966) );
  NAND U25689 ( .A(n24967), .B(n24966), .Z(n25275) );
  NAND U25690 ( .A(n34848), .B(n24968), .Z(n24970) );
  XNOR U25691 ( .A(n35375), .B(a[89]), .Z(n25116) );
  NAND U25692 ( .A(n34618), .B(n25116), .Z(n24969) );
  NAND U25693 ( .A(n24970), .B(n24969), .Z(n25272) );
  NAND U25694 ( .A(n35188), .B(n24971), .Z(n24973) );
  XNOR U25695 ( .A(n35540), .B(a[87]), .Z(n25119) );
  NANDN U25696 ( .A(n34968), .B(n25119), .Z(n24972) );
  AND U25697 ( .A(n24973), .B(n24972), .Z(n25273) );
  XNOR U25698 ( .A(n25272), .B(n25273), .Z(n25274) );
  XNOR U25699 ( .A(n25275), .B(n25274), .Z(n25080) );
  NANDN U25700 ( .A(n24975), .B(n24974), .Z(n24979) );
  NAND U25701 ( .A(n24977), .B(n24976), .Z(n24978) );
  NAND U25702 ( .A(n24979), .B(n24978), .Z(n25081) );
  XOR U25703 ( .A(n25080), .B(n25081), .Z(n25083) );
  XNOR U25704 ( .A(n25082), .B(n25083), .Z(n25194) );
  XNOR U25705 ( .A(n25193), .B(n25194), .Z(n25195) );
  XOR U25706 ( .A(n25196), .B(n25195), .Z(n25202) );
  NANDN U25707 ( .A(n24981), .B(n24980), .Z(n24985) );
  NAND U25708 ( .A(n24983), .B(n24982), .Z(n24984) );
  NAND U25709 ( .A(n24985), .B(n24984), .Z(n25293) );
  XOR U25710 ( .A(b[41]), .B(a[75]), .Z(n25162) );
  NANDN U25711 ( .A(n36905), .B(n25162), .Z(n24988) );
  NANDN U25712 ( .A(n24986), .B(n36807), .Z(n24987) );
  NAND U25713 ( .A(n24988), .B(n24987), .Z(n25190) );
  XNOR U25714 ( .A(b[57]), .B(a[59]), .Z(n25165) );
  OR U25715 ( .A(n25165), .B(n965), .Z(n24991) );
  NANDN U25716 ( .A(n24989), .B(n38194), .Z(n24990) );
  NAND U25717 ( .A(n24991), .B(n24990), .Z(n25187) );
  NAND U25718 ( .A(n38326), .B(n24992), .Z(n24994) );
  XOR U25719 ( .A(n38400), .B(n26122), .Z(n25168) );
  NANDN U25720 ( .A(n38273), .B(n25168), .Z(n24993) );
  AND U25721 ( .A(n24994), .B(n24993), .Z(n25188) );
  XNOR U25722 ( .A(n25187), .B(n25188), .Z(n25189) );
  XNOR U25723 ( .A(n25190), .B(n25189), .Z(n25290) );
  XNOR U25724 ( .A(b[33]), .B(a[83]), .Z(n25171) );
  NANDN U25725 ( .A(n25171), .B(n35620), .Z(n24997) );
  NANDN U25726 ( .A(n24995), .B(n35621), .Z(n24996) );
  NAND U25727 ( .A(n24997), .B(n24996), .Z(n25287) );
  NANDN U25728 ( .A(n966), .B(a[115]), .Z(n24998) );
  XOR U25729 ( .A(n29232), .B(n24998), .Z(n25000) );
  IV U25730 ( .A(a[114]), .Z(n37873) );
  NANDN U25731 ( .A(n37873), .B(n966), .Z(n24999) );
  AND U25732 ( .A(n25000), .B(n24999), .Z(n25284) );
  XOR U25733 ( .A(b[63]), .B(n25001), .Z(n25178) );
  NANDN U25734 ( .A(n25178), .B(n38422), .Z(n25004) );
  NANDN U25735 ( .A(n25002), .B(n38423), .Z(n25003) );
  AND U25736 ( .A(n25004), .B(n25003), .Z(n25285) );
  XNOR U25737 ( .A(n25284), .B(n25285), .Z(n25286) );
  XOR U25738 ( .A(n25287), .B(n25286), .Z(n25291) );
  XNOR U25739 ( .A(n25290), .B(n25291), .Z(n25292) );
  XOR U25740 ( .A(n25293), .B(n25292), .Z(n25095) );
  NANDN U25741 ( .A(n25006), .B(n25005), .Z(n25010) );
  NAND U25742 ( .A(n25008), .B(n25007), .Z(n25009) );
  NAND U25743 ( .A(n25010), .B(n25009), .Z(n25092) );
  NANDN U25744 ( .A(n25012), .B(n25011), .Z(n25016) );
  NAND U25745 ( .A(n25014), .B(n25013), .Z(n25015) );
  AND U25746 ( .A(n25016), .B(n25015), .Z(n25093) );
  XNOR U25747 ( .A(n25092), .B(n25093), .Z(n25094) );
  XNOR U25748 ( .A(n25095), .B(n25094), .Z(n25199) );
  NANDN U25749 ( .A(n25018), .B(n25017), .Z(n25022) );
  OR U25750 ( .A(n25020), .B(n25019), .Z(n25021) );
  AND U25751 ( .A(n25022), .B(n25021), .Z(n25200) );
  XNOR U25752 ( .A(n25199), .B(n25200), .Z(n25201) );
  XNOR U25753 ( .A(n25202), .B(n25201), .Z(n25077) );
  XNOR U25754 ( .A(n25076), .B(n25077), .Z(n25326) );
  XNOR U25755 ( .A(n25327), .B(n25326), .Z(n25328) );
  XNOR U25756 ( .A(n25328), .B(n25329), .Z(n25071) );
  XNOR U25757 ( .A(n25070), .B(n25071), .Z(n25064) );
  NANDN U25758 ( .A(n25028), .B(n25027), .Z(n25032) );
  NANDN U25759 ( .A(n25030), .B(n25029), .Z(n25031) );
  NAND U25760 ( .A(n25032), .B(n25031), .Z(n25063) );
  NAND U25761 ( .A(n25034), .B(n25033), .Z(n25038) );
  NAND U25762 ( .A(n25036), .B(n25035), .Z(n25037) );
  AND U25763 ( .A(n25038), .B(n25037), .Z(n25062) );
  XNOR U25764 ( .A(n25063), .B(n25062), .Z(n25065) );
  XOR U25765 ( .A(n25064), .B(n25065), .Z(n25059) );
  XOR U25766 ( .A(n25058), .B(n25059), .Z(n25050) );
  NANDN U25767 ( .A(n25040), .B(n25039), .Z(n25044) );
  NAND U25768 ( .A(n25042), .B(n25041), .Z(n25043) );
  AND U25769 ( .A(n25044), .B(n25043), .Z(n25051) );
  XOR U25770 ( .A(n25050), .B(n25051), .Z(n25052) );
  XNOR U25771 ( .A(n25053), .B(n25052), .Z(n25336) );
  XNOR U25772 ( .A(n25336), .B(sreg[179]), .Z(n25338) );
  NAND U25773 ( .A(n25045), .B(sreg[178]), .Z(n25049) );
  OR U25774 ( .A(n25047), .B(n25046), .Z(n25048) );
  AND U25775 ( .A(n25049), .B(n25048), .Z(n25337) );
  XOR U25776 ( .A(n25338), .B(n25337), .Z(c[179]) );
  NAND U25777 ( .A(n25051), .B(n25050), .Z(n25055) );
  NAND U25778 ( .A(n25053), .B(n25052), .Z(n25054) );
  NAND U25779 ( .A(n25055), .B(n25054), .Z(n25344) );
  NANDN U25780 ( .A(n25057), .B(n25056), .Z(n25061) );
  NAND U25781 ( .A(n25059), .B(n25058), .Z(n25060) );
  NAND U25782 ( .A(n25061), .B(n25060), .Z(n25342) );
  NANDN U25783 ( .A(n25063), .B(n25062), .Z(n25067) );
  NAND U25784 ( .A(n25065), .B(n25064), .Z(n25066) );
  NAND U25785 ( .A(n25067), .B(n25066), .Z(n25620) );
  NANDN U25786 ( .A(n25069), .B(n25068), .Z(n25073) );
  NANDN U25787 ( .A(n25071), .B(n25070), .Z(n25072) );
  NAND U25788 ( .A(n25073), .B(n25072), .Z(n25619) );
  NANDN U25789 ( .A(n25075), .B(n25074), .Z(n25079) );
  NANDN U25790 ( .A(n25077), .B(n25076), .Z(n25078) );
  NAND U25791 ( .A(n25079), .B(n25078), .Z(n25597) );
  NANDN U25792 ( .A(n25081), .B(n25080), .Z(n25085) );
  NANDN U25793 ( .A(n25083), .B(n25082), .Z(n25084) );
  NAND U25794 ( .A(n25085), .B(n25084), .Z(n25365) );
  NANDN U25795 ( .A(n25087), .B(n25086), .Z(n25091) );
  NAND U25796 ( .A(n25089), .B(n25088), .Z(n25090) );
  AND U25797 ( .A(n25091), .B(n25090), .Z(n25363) );
  NANDN U25798 ( .A(n25093), .B(n25092), .Z(n25097) );
  NAND U25799 ( .A(n25095), .B(n25094), .Z(n25096) );
  NAND U25800 ( .A(n25097), .B(n25096), .Z(n25364) );
  XOR U25801 ( .A(n25365), .B(n25366), .Z(n25372) );
  NANDN U25802 ( .A(n25099), .B(n25098), .Z(n25103) );
  NAND U25803 ( .A(n25101), .B(n25100), .Z(n25102) );
  NAND U25804 ( .A(n25103), .B(n25102), .Z(n25396) );
  XOR U25805 ( .A(b[37]), .B(n32814), .Z(n25424) );
  NANDN U25806 ( .A(n25424), .B(n36311), .Z(n25106) );
  NANDN U25807 ( .A(n25104), .B(n36309), .Z(n25105) );
  NAND U25808 ( .A(n25106), .B(n25105), .Z(n25457) );
  XOR U25809 ( .A(a[112]), .B(n968), .Z(n25427) );
  OR U25810 ( .A(n25427), .B(n29363), .Z(n25109) );
  NANDN U25811 ( .A(n25107), .B(n29864), .Z(n25108) );
  NAND U25812 ( .A(n25109), .B(n25108), .Z(n25454) );
  XOR U25813 ( .A(n37873), .B(n967), .Z(n25430) );
  NAND U25814 ( .A(n25430), .B(n28939), .Z(n25112) );
  NAND U25815 ( .A(n28938), .B(n25110), .Z(n25111) );
  AND U25816 ( .A(n25112), .B(n25111), .Z(n25455) );
  XNOR U25817 ( .A(n25454), .B(n25455), .Z(n25456) );
  XNOR U25818 ( .A(n25457), .B(n25456), .Z(n25387) );
  XOR U25819 ( .A(a[104]), .B(n971), .Z(n25433) );
  OR U25820 ( .A(n25433), .B(n31550), .Z(n25115) );
  NANDN U25821 ( .A(n25113), .B(n31874), .Z(n25114) );
  NAND U25822 ( .A(n25115), .B(n25114), .Z(n25585) );
  NAND U25823 ( .A(n34848), .B(n25116), .Z(n25118) );
  XOR U25824 ( .A(n35375), .B(n34851), .Z(n25436) );
  NAND U25825 ( .A(n34618), .B(n25436), .Z(n25117) );
  NAND U25826 ( .A(n25118), .B(n25117), .Z(n25582) );
  NAND U25827 ( .A(n35188), .B(n25119), .Z(n25121) );
  XOR U25828 ( .A(n35540), .B(n34048), .Z(n25439) );
  NANDN U25829 ( .A(n34968), .B(n25439), .Z(n25120) );
  AND U25830 ( .A(n25121), .B(n25120), .Z(n25583) );
  XNOR U25831 ( .A(n25582), .B(n25583), .Z(n25584) );
  XOR U25832 ( .A(n25585), .B(n25584), .Z(n25388) );
  XOR U25833 ( .A(n25387), .B(n25388), .Z(n25390) );
  NANDN U25834 ( .A(n25123), .B(n25122), .Z(n25127) );
  NAND U25835 ( .A(n25125), .B(n25124), .Z(n25126) );
  NAND U25836 ( .A(n25127), .B(n25126), .Z(n25389) );
  XNOR U25837 ( .A(n25390), .B(n25389), .Z(n25393) );
  NANDN U25838 ( .A(n25129), .B(n25128), .Z(n25133) );
  NAND U25839 ( .A(n25131), .B(n25130), .Z(n25132) );
  NAND U25840 ( .A(n25133), .B(n25132), .Z(n25522) );
  ANDN U25841 ( .B(b[63]), .A(n25134), .Z(n25537) );
  NANDN U25842 ( .A(n25135), .B(n38369), .Z(n25137) );
  XOR U25843 ( .A(b[61]), .B(n25860), .Z(n25418) );
  OR U25844 ( .A(n25418), .B(n38371), .Z(n25136) );
  NAND U25845 ( .A(n25137), .B(n25136), .Z(n25535) );
  NANDN U25846 ( .A(n25138), .B(n35311), .Z(n25140) );
  XOR U25847 ( .A(b[31]), .B(n33628), .Z(n25421) );
  NANDN U25848 ( .A(n25421), .B(n35313), .Z(n25139) );
  AND U25849 ( .A(n25140), .B(n25139), .Z(n25534) );
  XNOR U25850 ( .A(n25535), .B(n25534), .Z(n25536) );
  XOR U25851 ( .A(n25537), .B(n25536), .Z(n25519) );
  NAND U25852 ( .A(n33283), .B(n25141), .Z(n25143) );
  XOR U25853 ( .A(n35783), .B(n33020), .Z(n25403) );
  NANDN U25854 ( .A(n33021), .B(n25403), .Z(n25142) );
  NAND U25855 ( .A(n25143), .B(n25142), .Z(n25482) );
  XNOR U25856 ( .A(a[96]), .B(b[21]), .Z(n25406) );
  OR U25857 ( .A(n25406), .B(n33634), .Z(n25146) );
  NANDN U25858 ( .A(n25144), .B(n33464), .Z(n25145) );
  NAND U25859 ( .A(n25146), .B(n25145), .Z(n25479) );
  NAND U25860 ( .A(n34044), .B(n25147), .Z(n25149) );
  XOR U25861 ( .A(n35191), .B(n34510), .Z(n25409) );
  NANDN U25862 ( .A(n33867), .B(n25409), .Z(n25148) );
  AND U25863 ( .A(n25149), .B(n25148), .Z(n25480) );
  XNOR U25864 ( .A(n25479), .B(n25480), .Z(n25481) );
  XNOR U25865 ( .A(n25482), .B(n25481), .Z(n25520) );
  XNOR U25866 ( .A(n25519), .B(n25520), .Z(n25521) );
  XNOR U25867 ( .A(n25522), .B(n25521), .Z(n25394) );
  XNOR U25868 ( .A(n25393), .B(n25394), .Z(n25395) );
  XOR U25869 ( .A(n25396), .B(n25395), .Z(n25494) );
  NANDN U25870 ( .A(n25151), .B(n25150), .Z(n25155) );
  OR U25871 ( .A(n25153), .B(n25152), .Z(n25154) );
  NAND U25872 ( .A(n25155), .B(n25154), .Z(n25492) );
  NANDN U25873 ( .A(n25157), .B(n25156), .Z(n25161) );
  NAND U25874 ( .A(n25159), .B(n25158), .Z(n25160) );
  NAND U25875 ( .A(n25161), .B(n25160), .Z(n25384) );
  XNOR U25876 ( .A(b[41]), .B(a[76]), .Z(n25470) );
  OR U25877 ( .A(n25470), .B(n36905), .Z(n25164) );
  NAND U25878 ( .A(n25162), .B(n36807), .Z(n25163) );
  NAND U25879 ( .A(n25164), .B(n25163), .Z(n25488) );
  XOR U25880 ( .A(b[57]), .B(n27436), .Z(n25473) );
  OR U25881 ( .A(n25473), .B(n965), .Z(n25167) );
  NANDN U25882 ( .A(n25165), .B(n38194), .Z(n25166) );
  NAND U25883 ( .A(n25167), .B(n25166), .Z(n25485) );
  NAND U25884 ( .A(n38326), .B(n25168), .Z(n25170) );
  XOR U25885 ( .A(n38400), .B(n26347), .Z(n25476) );
  NANDN U25886 ( .A(n38273), .B(n25476), .Z(n25169) );
  AND U25887 ( .A(n25170), .B(n25169), .Z(n25486) );
  XNOR U25888 ( .A(n25485), .B(n25486), .Z(n25487) );
  XNOR U25889 ( .A(n25488), .B(n25487), .Z(n25546) );
  XOR U25890 ( .A(b[33]), .B(n33185), .Z(n25460) );
  NANDN U25891 ( .A(n25460), .B(n35620), .Z(n25173) );
  NANDN U25892 ( .A(n25171), .B(n35621), .Z(n25172) );
  NAND U25893 ( .A(n25173), .B(n25172), .Z(n25561) );
  NANDN U25894 ( .A(n966), .B(a[116]), .Z(n25174) );
  XOR U25895 ( .A(n29232), .B(n25174), .Z(n25176) );
  NANDN U25896 ( .A(b[0]), .B(a[115]), .Z(n25175) );
  AND U25897 ( .A(n25176), .B(n25175), .Z(n25558) );
  XOR U25898 ( .A(b[63]), .B(n25177), .Z(n25467) );
  NANDN U25899 ( .A(n25467), .B(n38422), .Z(n25180) );
  NANDN U25900 ( .A(n25178), .B(n38423), .Z(n25179) );
  AND U25901 ( .A(n25180), .B(n25179), .Z(n25559) );
  XNOR U25902 ( .A(n25558), .B(n25559), .Z(n25560) );
  XOR U25903 ( .A(n25561), .B(n25560), .Z(n25547) );
  XNOR U25904 ( .A(n25546), .B(n25547), .Z(n25548) );
  NANDN U25905 ( .A(n25182), .B(n25181), .Z(n25186) );
  NAND U25906 ( .A(n25184), .B(n25183), .Z(n25185) );
  AND U25907 ( .A(n25186), .B(n25185), .Z(n25549) );
  XNOR U25908 ( .A(n25548), .B(n25549), .Z(n25382) );
  NANDN U25909 ( .A(n25188), .B(n25187), .Z(n25192) );
  NAND U25910 ( .A(n25190), .B(n25189), .Z(n25191) );
  AND U25911 ( .A(n25192), .B(n25191), .Z(n25381) );
  XNOR U25912 ( .A(n25382), .B(n25381), .Z(n25383) );
  XNOR U25913 ( .A(n25384), .B(n25383), .Z(n25491) );
  XOR U25914 ( .A(n25492), .B(n25491), .Z(n25493) );
  XNOR U25915 ( .A(n25494), .B(n25493), .Z(n25369) );
  NANDN U25916 ( .A(n25194), .B(n25193), .Z(n25198) );
  NANDN U25917 ( .A(n25196), .B(n25195), .Z(n25197) );
  AND U25918 ( .A(n25198), .B(n25197), .Z(n25370) );
  XNOR U25919 ( .A(n25369), .B(n25370), .Z(n25371) );
  XOR U25920 ( .A(n25372), .B(n25371), .Z(n25594) );
  XNOR U25921 ( .A(b[35]), .B(a[82]), .Z(n25525) );
  NANDN U25922 ( .A(n25525), .B(n35985), .Z(n25205) );
  NAND U25923 ( .A(n25203), .B(n35986), .Z(n25204) );
  NAND U25924 ( .A(n25205), .B(n25204), .Z(n25591) );
  XOR U25925 ( .A(n37336), .B(n31123), .Z(n25528) );
  NAND U25926 ( .A(n25528), .B(n29949), .Z(n25208) );
  NAND U25927 ( .A(n29948), .B(n25206), .Z(n25207) );
  NAND U25928 ( .A(n25208), .B(n25207), .Z(n25588) );
  XNOR U25929 ( .A(b[55]), .B(a[62]), .Z(n25531) );
  NANDN U25930 ( .A(n25531), .B(n38075), .Z(n25211) );
  NANDN U25931 ( .A(n25209), .B(n38073), .Z(n25210) );
  AND U25932 ( .A(n25211), .B(n25210), .Z(n25589) );
  XNOR U25933 ( .A(n25588), .B(n25589), .Z(n25590) );
  XNOR U25934 ( .A(n25591), .B(n25590), .Z(n25378) );
  NANDN U25935 ( .A(n25213), .B(n25212), .Z(n25217) );
  NAND U25936 ( .A(n25215), .B(n25214), .Z(n25216) );
  NAND U25937 ( .A(n25217), .B(n25216), .Z(n25375) );
  NANDN U25938 ( .A(n25219), .B(n25218), .Z(n25223) );
  NAND U25939 ( .A(n25221), .B(n25220), .Z(n25222) );
  NAND U25940 ( .A(n25223), .B(n25222), .Z(n25376) );
  XNOR U25941 ( .A(n25375), .B(n25376), .Z(n25377) );
  XOR U25942 ( .A(n25378), .B(n25377), .Z(n25355) );
  NANDN U25943 ( .A(n25225), .B(n25224), .Z(n25229) );
  NANDN U25944 ( .A(n25227), .B(n25226), .Z(n25228) );
  NAND U25945 ( .A(n25229), .B(n25228), .Z(n25354) );
  XOR U25946 ( .A(a[106]), .B(n970), .Z(n25495) );
  OR U25947 ( .A(n25495), .B(n31369), .Z(n25232) );
  NANDN U25948 ( .A(n25230), .B(n31119), .Z(n25231) );
  NAND U25949 ( .A(n25232), .B(n25231), .Z(n25516) );
  XOR U25950 ( .A(b[43]), .B(n31372), .Z(n25498) );
  NANDN U25951 ( .A(n25498), .B(n37068), .Z(n25235) );
  NANDN U25952 ( .A(n25233), .B(n37069), .Z(n25234) );
  NAND U25953 ( .A(n25235), .B(n25234), .Z(n25513) );
  XNOR U25954 ( .A(b[45]), .B(a[72]), .Z(n25501) );
  NANDN U25955 ( .A(n25501), .B(n37261), .Z(n25238) );
  NANDN U25956 ( .A(n25236), .B(n37262), .Z(n25237) );
  AND U25957 ( .A(n25238), .B(n25237), .Z(n25514) );
  XNOR U25958 ( .A(n25513), .B(n25514), .Z(n25515) );
  XNOR U25959 ( .A(n25516), .B(n25515), .Z(n25402) );
  XOR U25960 ( .A(b[49]), .B(n29868), .Z(n25504) );
  OR U25961 ( .A(n25504), .B(n37756), .Z(n25241) );
  NANDN U25962 ( .A(n25239), .B(n37652), .Z(n25240) );
  NAND U25963 ( .A(n25241), .B(n25240), .Z(n25543) );
  NAND U25964 ( .A(n37469), .B(n25242), .Z(n25244) );
  XOR U25965 ( .A(n978), .B(n30379), .Z(n25507) );
  NAND U25966 ( .A(n25507), .B(n37471), .Z(n25243) );
  NAND U25967 ( .A(n25244), .B(n25243), .Z(n25540) );
  XOR U25968 ( .A(a[108]), .B(n969), .Z(n25510) );
  NANDN U25969 ( .A(n25510), .B(n30509), .Z(n25247) );
  NANDN U25970 ( .A(n25245), .B(n30846), .Z(n25246) );
  AND U25971 ( .A(n25247), .B(n25246), .Z(n25541) );
  XNOR U25972 ( .A(n25540), .B(n25541), .Z(n25542) );
  XNOR U25973 ( .A(n25543), .B(n25542), .Z(n25399) );
  NANDN U25974 ( .A(n25249), .B(n25248), .Z(n25253) );
  NAND U25975 ( .A(n25251), .B(n25250), .Z(n25252) );
  NAND U25976 ( .A(n25253), .B(n25252), .Z(n25400) );
  XNOR U25977 ( .A(n25399), .B(n25400), .Z(n25401) );
  XOR U25978 ( .A(n25402), .B(n25401), .Z(n25353) );
  XOR U25979 ( .A(n25354), .B(n25353), .Z(n25356) );
  XOR U25980 ( .A(n25355), .B(n25356), .Z(n25347) );
  XOR U25981 ( .A(a[102]), .B(n972), .Z(n25564) );
  OR U25982 ( .A(n25564), .B(n32010), .Z(n25256) );
  NANDN U25983 ( .A(n25254), .B(n32011), .Z(n25255) );
  NAND U25984 ( .A(n25256), .B(n25255), .Z(n25415) );
  XNOR U25985 ( .A(n34852), .B(b[25]), .Z(n25567) );
  NANDN U25986 ( .A(n34219), .B(n25567), .Z(n25259) );
  NAND U25987 ( .A(n34217), .B(n25257), .Z(n25258) );
  NAND U25988 ( .A(n25259), .B(n25258), .Z(n25412) );
  XNOR U25989 ( .A(a[100]), .B(b[17]), .Z(n25570) );
  NANDN U25990 ( .A(n25570), .B(n32543), .Z(n25262) );
  NAND U25991 ( .A(n25260), .B(n32541), .Z(n25261) );
  AND U25992 ( .A(n25262), .B(n25261), .Z(n25413) );
  XNOR U25993 ( .A(n25412), .B(n25413), .Z(n25414) );
  XNOR U25994 ( .A(n25415), .B(n25414), .Z(n25448) );
  XOR U25995 ( .A(b[39]), .B(n31870), .Z(n25573) );
  NANDN U25996 ( .A(n25573), .B(n36553), .Z(n25265) );
  NANDN U25997 ( .A(n25263), .B(n36643), .Z(n25264) );
  NAND U25998 ( .A(n25265), .B(n25264), .Z(n25445) );
  XOR U25999 ( .A(b[51]), .B(n28701), .Z(n25576) );
  NANDN U26000 ( .A(n25576), .B(n37803), .Z(n25268) );
  NANDN U26001 ( .A(n25266), .B(n37802), .Z(n25267) );
  NAND U26002 ( .A(n25268), .B(n25267), .Z(n25442) );
  XNOR U26003 ( .A(b[53]), .B(a[64]), .Z(n25579) );
  NANDN U26004 ( .A(n25579), .B(n37940), .Z(n25271) );
  NANDN U26005 ( .A(n25269), .B(n37941), .Z(n25270) );
  AND U26006 ( .A(n25271), .B(n25270), .Z(n25443) );
  XNOR U26007 ( .A(n25442), .B(n25443), .Z(n25444) );
  XOR U26008 ( .A(n25445), .B(n25444), .Z(n25449) );
  XOR U26009 ( .A(n25448), .B(n25449), .Z(n25451) );
  NANDN U26010 ( .A(n25273), .B(n25272), .Z(n25277) );
  NAND U26011 ( .A(n25275), .B(n25274), .Z(n25276) );
  NAND U26012 ( .A(n25277), .B(n25276), .Z(n25450) );
  XNOR U26013 ( .A(n25451), .B(n25450), .Z(n25555) );
  NANDN U26014 ( .A(n25279), .B(n25278), .Z(n25283) );
  NAND U26015 ( .A(n25281), .B(n25280), .Z(n25282) );
  NAND U26016 ( .A(n25283), .B(n25282), .Z(n25552) );
  NANDN U26017 ( .A(n25285), .B(n25284), .Z(n25289) );
  NAND U26018 ( .A(n25287), .B(n25286), .Z(n25288) );
  AND U26019 ( .A(n25289), .B(n25288), .Z(n25553) );
  XNOR U26020 ( .A(n25552), .B(n25553), .Z(n25554) );
  XNOR U26021 ( .A(n25555), .B(n25554), .Z(n25359) );
  NANDN U26022 ( .A(n25291), .B(n25290), .Z(n25295) );
  NANDN U26023 ( .A(n25293), .B(n25292), .Z(n25294) );
  AND U26024 ( .A(n25295), .B(n25294), .Z(n25360) );
  XNOR U26025 ( .A(n25359), .B(n25360), .Z(n25361) );
  NANDN U26026 ( .A(n25297), .B(n25296), .Z(n25301) );
  NAND U26027 ( .A(n25299), .B(n25298), .Z(n25300) );
  AND U26028 ( .A(n25301), .B(n25300), .Z(n25362) );
  XNOR U26029 ( .A(n25361), .B(n25362), .Z(n25348) );
  XNOR U26030 ( .A(n25347), .B(n25348), .Z(n25349) );
  XNOR U26031 ( .A(n25350), .B(n25349), .Z(n25595) );
  XOR U26032 ( .A(n25594), .B(n25595), .Z(n25596) );
  XNOR U26033 ( .A(n25597), .B(n25596), .Z(n25609) );
  NANDN U26034 ( .A(n25303), .B(n25302), .Z(n25307) );
  NAND U26035 ( .A(n25305), .B(n25304), .Z(n25306) );
  NAND U26036 ( .A(n25307), .B(n25306), .Z(n25606) );
  NANDN U26037 ( .A(n25309), .B(n25308), .Z(n25313) );
  NAND U26038 ( .A(n25311), .B(n25310), .Z(n25312) );
  NAND U26039 ( .A(n25313), .B(n25312), .Z(n25603) );
  NANDN U26040 ( .A(n25315), .B(n25314), .Z(n25319) );
  NAND U26041 ( .A(n25317), .B(n25316), .Z(n25318) );
  NAND U26042 ( .A(n25319), .B(n25318), .Z(n25601) );
  OR U26043 ( .A(n25321), .B(n25320), .Z(n25325) );
  NAND U26044 ( .A(n25323), .B(n25322), .Z(n25324) );
  AND U26045 ( .A(n25325), .B(n25324), .Z(n25600) );
  XNOR U26046 ( .A(n25601), .B(n25600), .Z(n25602) );
  XOR U26047 ( .A(n25603), .B(n25602), .Z(n25607) );
  XOR U26048 ( .A(n25606), .B(n25607), .Z(n25608) );
  XOR U26049 ( .A(n25609), .B(n25608), .Z(n25615) );
  NANDN U26050 ( .A(n25331), .B(n25330), .Z(n25335) );
  NANDN U26051 ( .A(n25333), .B(n25332), .Z(n25334) );
  NAND U26052 ( .A(n25335), .B(n25334), .Z(n25613) );
  XNOR U26053 ( .A(n25612), .B(n25613), .Z(n25614) );
  XNOR U26054 ( .A(n25615), .B(n25614), .Z(n25618) );
  XNOR U26055 ( .A(n25619), .B(n25618), .Z(n25621) );
  XNOR U26056 ( .A(n25620), .B(n25621), .Z(n25341) );
  XOR U26057 ( .A(n25342), .B(n25341), .Z(n25343) );
  XNOR U26058 ( .A(n25344), .B(n25343), .Z(n25624) );
  XNOR U26059 ( .A(n25624), .B(sreg[180]), .Z(n25626) );
  NAND U26060 ( .A(n25336), .B(sreg[179]), .Z(n25340) );
  OR U26061 ( .A(n25338), .B(n25337), .Z(n25339) );
  AND U26062 ( .A(n25340), .B(n25339), .Z(n25625) );
  XOR U26063 ( .A(n25626), .B(n25625), .Z(c[180]) );
  NAND U26064 ( .A(n25342), .B(n25341), .Z(n25346) );
  NAND U26065 ( .A(n25344), .B(n25343), .Z(n25345) );
  NAND U26066 ( .A(n25346), .B(n25345), .Z(n25632) );
  NANDN U26067 ( .A(n25348), .B(n25347), .Z(n25352) );
  NAND U26068 ( .A(n25350), .B(n25349), .Z(n25351) );
  NAND U26069 ( .A(n25352), .B(n25351), .Z(n25647) );
  NAND U26070 ( .A(n25354), .B(n25353), .Z(n25358) );
  NAND U26071 ( .A(n25356), .B(n25355), .Z(n25357) );
  NAND U26072 ( .A(n25358), .B(n25357), .Z(n25656) );
  OR U26073 ( .A(n25364), .B(n25363), .Z(n25368) );
  NANDN U26074 ( .A(n25366), .B(n25365), .Z(n25367) );
  AND U26075 ( .A(n25368), .B(n25367), .Z(n25653) );
  XNOR U26076 ( .A(n25654), .B(n25653), .Z(n25655) );
  XOR U26077 ( .A(n25656), .B(n25655), .Z(n25648) );
  XOR U26078 ( .A(n25647), .B(n25648), .Z(n25649) );
  NANDN U26079 ( .A(n25370), .B(n25369), .Z(n25374) );
  NAND U26080 ( .A(n25372), .B(n25371), .Z(n25373) );
  NAND U26081 ( .A(n25374), .B(n25373), .Z(n25662) );
  NANDN U26082 ( .A(n25376), .B(n25375), .Z(n25380) );
  NAND U26083 ( .A(n25378), .B(n25377), .Z(n25379) );
  NAND U26084 ( .A(n25380), .B(n25379), .Z(n25905) );
  NANDN U26085 ( .A(n25382), .B(n25381), .Z(n25386) );
  NANDN U26086 ( .A(n25384), .B(n25383), .Z(n25385) );
  NAND U26087 ( .A(n25386), .B(n25385), .Z(n25902) );
  NANDN U26088 ( .A(n25388), .B(n25387), .Z(n25392) );
  OR U26089 ( .A(n25390), .B(n25389), .Z(n25391) );
  AND U26090 ( .A(n25392), .B(n25391), .Z(n25903) );
  XNOR U26091 ( .A(n25902), .B(n25903), .Z(n25904) );
  XNOR U26092 ( .A(n25905), .B(n25904), .Z(n25664) );
  NANDN U26093 ( .A(n25394), .B(n25393), .Z(n25398) );
  NANDN U26094 ( .A(n25396), .B(n25395), .Z(n25397) );
  AND U26095 ( .A(n25398), .B(n25397), .Z(n25663) );
  XNOR U26096 ( .A(n25664), .B(n25663), .Z(n25665) );
  NAND U26097 ( .A(n33283), .B(n25403), .Z(n25405) );
  XNOR U26098 ( .A(a[99]), .B(n33020), .Z(n25836) );
  NANDN U26099 ( .A(n33021), .B(n25836), .Z(n25404) );
  NAND U26100 ( .A(n25405), .B(n25404), .Z(n25867) );
  XOR U26101 ( .A(a[97]), .B(b[21]), .Z(n25839) );
  NANDN U26102 ( .A(n33634), .B(n25839), .Z(n25408) );
  NANDN U26103 ( .A(n25406), .B(n33464), .Z(n25407) );
  NAND U26104 ( .A(n25408), .B(n25407), .Z(n25864) );
  NAND U26105 ( .A(n34044), .B(n25409), .Z(n25411) );
  XOR U26106 ( .A(n35628), .B(n34510), .Z(n25842) );
  NANDN U26107 ( .A(n33867), .B(n25842), .Z(n25410) );
  AND U26108 ( .A(n25411), .B(n25410), .Z(n25865) );
  XNOR U26109 ( .A(n25864), .B(n25865), .Z(n25866) );
  XNOR U26110 ( .A(n25867), .B(n25866), .Z(n25669) );
  NANDN U26111 ( .A(n25413), .B(n25412), .Z(n25417) );
  NAND U26112 ( .A(n25415), .B(n25414), .Z(n25416) );
  NAND U26113 ( .A(n25417), .B(n25416), .Z(n25670) );
  XNOR U26114 ( .A(n25669), .B(n25670), .Z(n25671) );
  NAND U26115 ( .A(a[53]), .B(b[63]), .Z(n25711) );
  NANDN U26116 ( .A(n25418), .B(n38369), .Z(n25420) );
  XOR U26117 ( .A(b[61]), .B(n26122), .Z(n25830) );
  OR U26118 ( .A(n25830), .B(n38371), .Z(n25419) );
  NAND U26119 ( .A(n25420), .B(n25419), .Z(n25709) );
  NANDN U26120 ( .A(n25421), .B(n35311), .Z(n25423) );
  XNOR U26121 ( .A(b[31]), .B(a[87]), .Z(n25833) );
  NANDN U26122 ( .A(n25833), .B(n35313), .Z(n25422) );
  AND U26123 ( .A(n25423), .B(n25422), .Z(n25708) );
  XNOR U26124 ( .A(n25709), .B(n25708), .Z(n25710) );
  XNOR U26125 ( .A(n25711), .B(n25710), .Z(n25672) );
  XOR U26126 ( .A(n25671), .B(n25672), .Z(n25772) );
  XNOR U26127 ( .A(b[37]), .B(a[81]), .Z(n25800) );
  NANDN U26128 ( .A(n25800), .B(n36311), .Z(n25426) );
  NANDN U26129 ( .A(n25424), .B(n36309), .Z(n25425) );
  NAND U26130 ( .A(n25426), .B(n25425), .Z(n25879) );
  XNOR U26131 ( .A(a[113]), .B(b[5]), .Z(n25803) );
  OR U26132 ( .A(n25803), .B(n29363), .Z(n25429) );
  NANDN U26133 ( .A(n25427), .B(n29864), .Z(n25428) );
  NAND U26134 ( .A(n25429), .B(n25428), .Z(n25876) );
  XNOR U26135 ( .A(a[115]), .B(n967), .Z(n25806) );
  NAND U26136 ( .A(n25806), .B(n28939), .Z(n25432) );
  NAND U26137 ( .A(n28938), .B(n25430), .Z(n25431) );
  AND U26138 ( .A(n25432), .B(n25431), .Z(n25877) );
  XNOR U26139 ( .A(n25876), .B(n25877), .Z(n25878) );
  XNOR U26140 ( .A(n25879), .B(n25878), .Z(n25793) );
  XNOR U26141 ( .A(a[105]), .B(b[13]), .Z(n25809) );
  OR U26142 ( .A(n25809), .B(n31550), .Z(n25435) );
  NANDN U26143 ( .A(n25433), .B(n31874), .Z(n25434) );
  NAND U26144 ( .A(n25435), .B(n25434), .Z(n25753) );
  NAND U26145 ( .A(n34848), .B(n25436), .Z(n25438) );
  XNOR U26146 ( .A(n35375), .B(a[91]), .Z(n25812) );
  NAND U26147 ( .A(n34618), .B(n25812), .Z(n25437) );
  NAND U26148 ( .A(n25438), .B(n25437), .Z(n25750) );
  NAND U26149 ( .A(n35188), .B(n25439), .Z(n25441) );
  XNOR U26150 ( .A(n35540), .B(a[89]), .Z(n25815) );
  NANDN U26151 ( .A(n34968), .B(n25815), .Z(n25440) );
  AND U26152 ( .A(n25441), .B(n25440), .Z(n25751) );
  XNOR U26153 ( .A(n25750), .B(n25751), .Z(n25752) );
  XNOR U26154 ( .A(n25753), .B(n25752), .Z(n25790) );
  NANDN U26155 ( .A(n25443), .B(n25442), .Z(n25447) );
  NAND U26156 ( .A(n25445), .B(n25444), .Z(n25446) );
  NAND U26157 ( .A(n25447), .B(n25446), .Z(n25791) );
  XNOR U26158 ( .A(n25790), .B(n25791), .Z(n25792) );
  XOR U26159 ( .A(n25793), .B(n25792), .Z(n25773) );
  XNOR U26160 ( .A(n25772), .B(n25773), .Z(n25774) );
  XOR U26161 ( .A(n25775), .B(n25774), .Z(n25768) );
  NANDN U26162 ( .A(n25449), .B(n25448), .Z(n25453) );
  OR U26163 ( .A(n25451), .B(n25450), .Z(n25452) );
  NAND U26164 ( .A(n25453), .B(n25452), .Z(n25767) );
  NANDN U26165 ( .A(n25455), .B(n25454), .Z(n25459) );
  NAND U26166 ( .A(n25457), .B(n25456), .Z(n25458) );
  NAND U26167 ( .A(n25459), .B(n25458), .Z(n25787) );
  XNOR U26168 ( .A(b[33]), .B(a[85]), .Z(n25854) );
  NANDN U26169 ( .A(n25854), .B(n35620), .Z(n25462) );
  NANDN U26170 ( .A(n25460), .B(n35621), .Z(n25461) );
  NAND U26171 ( .A(n25462), .B(n25461), .Z(n25765) );
  NANDN U26172 ( .A(n966), .B(a[117]), .Z(n25463) );
  XOR U26173 ( .A(n29232), .B(n25463), .Z(n25465) );
  IV U26174 ( .A(a[116]), .Z(n38046) );
  NANDN U26175 ( .A(n38046), .B(n966), .Z(n25464) );
  AND U26176 ( .A(n25465), .B(n25464), .Z(n25762) );
  XOR U26177 ( .A(b[63]), .B(n25466), .Z(n25861) );
  NANDN U26178 ( .A(n25861), .B(n38422), .Z(n25469) );
  NANDN U26179 ( .A(n25467), .B(n38423), .Z(n25468) );
  AND U26180 ( .A(n25469), .B(n25468), .Z(n25763) );
  XNOR U26181 ( .A(n25762), .B(n25763), .Z(n25764) );
  XNOR U26182 ( .A(n25765), .B(n25764), .Z(n25728) );
  XOR U26183 ( .A(b[41]), .B(a[77]), .Z(n25845) );
  NANDN U26184 ( .A(n36905), .B(n25845), .Z(n25472) );
  NANDN U26185 ( .A(n25470), .B(n36807), .Z(n25471) );
  NAND U26186 ( .A(n25472), .B(n25471), .Z(n25873) );
  XOR U26187 ( .A(b[57]), .B(n27773), .Z(n25848) );
  OR U26188 ( .A(n25848), .B(n965), .Z(n25475) );
  NANDN U26189 ( .A(n25473), .B(n38194), .Z(n25474) );
  NAND U26190 ( .A(n25475), .B(n25474), .Z(n25870) );
  NAND U26191 ( .A(n38326), .B(n25476), .Z(n25478) );
  XNOR U26192 ( .A(n38400), .B(a[59]), .Z(n25851) );
  NANDN U26193 ( .A(n38273), .B(n25851), .Z(n25477) );
  AND U26194 ( .A(n25478), .B(n25477), .Z(n25871) );
  XNOR U26195 ( .A(n25870), .B(n25871), .Z(n25872) );
  XNOR U26196 ( .A(n25873), .B(n25872), .Z(n25726) );
  NANDN U26197 ( .A(n25480), .B(n25479), .Z(n25484) );
  NAND U26198 ( .A(n25482), .B(n25481), .Z(n25483) );
  NAND U26199 ( .A(n25484), .B(n25483), .Z(n25727) );
  XOR U26200 ( .A(n25726), .B(n25727), .Z(n25729) );
  XNOR U26201 ( .A(n25728), .B(n25729), .Z(n25784) );
  NANDN U26202 ( .A(n25486), .B(n25485), .Z(n25490) );
  NAND U26203 ( .A(n25488), .B(n25487), .Z(n25489) );
  AND U26204 ( .A(n25490), .B(n25489), .Z(n25785) );
  XOR U26205 ( .A(n25784), .B(n25785), .Z(n25786) );
  XNOR U26206 ( .A(n25787), .B(n25786), .Z(n25766) );
  XNOR U26207 ( .A(n25767), .B(n25766), .Z(n25769) );
  XNOR U26208 ( .A(n25768), .B(n25769), .Z(n25666) );
  XNOR U26209 ( .A(n25665), .B(n25666), .Z(n25659) );
  XNOR U26210 ( .A(a[107]), .B(b[11]), .Z(n25675) );
  OR U26211 ( .A(n25675), .B(n31369), .Z(n25497) );
  NANDN U26212 ( .A(n25495), .B(n31119), .Z(n25496) );
  NAND U26213 ( .A(n25497), .B(n25496), .Z(n25696) );
  XNOR U26214 ( .A(b[43]), .B(a[75]), .Z(n25678) );
  NANDN U26215 ( .A(n25678), .B(n37068), .Z(n25500) );
  NANDN U26216 ( .A(n25498), .B(n37069), .Z(n25499) );
  NAND U26217 ( .A(n25500), .B(n25499), .Z(n25693) );
  XOR U26218 ( .A(b[45]), .B(a[73]), .Z(n25681) );
  NAND U26219 ( .A(n25681), .B(n37261), .Z(n25503) );
  NANDN U26220 ( .A(n25501), .B(n37262), .Z(n25502) );
  AND U26221 ( .A(n25503), .B(n25502), .Z(n25694) );
  XNOR U26222 ( .A(n25693), .B(n25694), .Z(n25695) );
  XNOR U26223 ( .A(n25696), .B(n25695), .Z(n25799) );
  XNOR U26224 ( .A(b[49]), .B(a[69]), .Z(n25684) );
  OR U26225 ( .A(n25684), .B(n37756), .Z(n25506) );
  NANDN U26226 ( .A(n25504), .B(n37652), .Z(n25505) );
  NAND U26227 ( .A(n25506), .B(n25505), .Z(n25717) );
  NAND U26228 ( .A(n37469), .B(n25507), .Z(n25509) );
  XOR U26229 ( .A(n978), .B(n30543), .Z(n25687) );
  NAND U26230 ( .A(n25687), .B(n37471), .Z(n25508) );
  NAND U26231 ( .A(n25509), .B(n25508), .Z(n25714) );
  XNOR U26232 ( .A(a[109]), .B(b[9]), .Z(n25690) );
  NANDN U26233 ( .A(n25690), .B(n30509), .Z(n25512) );
  NANDN U26234 ( .A(n25510), .B(n30846), .Z(n25511) );
  AND U26235 ( .A(n25512), .B(n25511), .Z(n25715) );
  XNOR U26236 ( .A(n25714), .B(n25715), .Z(n25716) );
  XNOR U26237 ( .A(n25717), .B(n25716), .Z(n25796) );
  NANDN U26238 ( .A(n25514), .B(n25513), .Z(n25518) );
  NAND U26239 ( .A(n25516), .B(n25515), .Z(n25517) );
  NAND U26240 ( .A(n25518), .B(n25517), .Z(n25797) );
  XNOR U26241 ( .A(n25796), .B(n25797), .Z(n25798) );
  XOR U26242 ( .A(n25799), .B(n25798), .Z(n25890) );
  NANDN U26243 ( .A(n25520), .B(n25519), .Z(n25524) );
  NAND U26244 ( .A(n25522), .B(n25521), .Z(n25523) );
  AND U26245 ( .A(n25524), .B(n25523), .Z(n25891) );
  XNOR U26246 ( .A(n25890), .B(n25891), .Z(n25893) );
  XOR U26247 ( .A(b[35]), .B(a[83]), .Z(n25699) );
  NAND U26248 ( .A(n35985), .B(n25699), .Z(n25527) );
  NANDN U26249 ( .A(n25525), .B(n35986), .Z(n25526) );
  NAND U26250 ( .A(n25527), .B(n25526), .Z(n25759) );
  XNOR U26251 ( .A(a[111]), .B(n31123), .Z(n25702) );
  NAND U26252 ( .A(n25702), .B(n29949), .Z(n25530) );
  NAND U26253 ( .A(n29948), .B(n25528), .Z(n25529) );
  NAND U26254 ( .A(n25530), .B(n25529), .Z(n25756) );
  XNOR U26255 ( .A(b[55]), .B(a[63]), .Z(n25705) );
  NANDN U26256 ( .A(n25705), .B(n38075), .Z(n25533) );
  NANDN U26257 ( .A(n25531), .B(n38073), .Z(n25532) );
  AND U26258 ( .A(n25533), .B(n25532), .Z(n25757) );
  XNOR U26259 ( .A(n25756), .B(n25757), .Z(n25758) );
  XNOR U26260 ( .A(n25759), .B(n25758), .Z(n25781) );
  NANDN U26261 ( .A(n25535), .B(n25534), .Z(n25539) );
  NANDN U26262 ( .A(n25537), .B(n25536), .Z(n25538) );
  NAND U26263 ( .A(n25539), .B(n25538), .Z(n25778) );
  NANDN U26264 ( .A(n25541), .B(n25540), .Z(n25545) );
  NAND U26265 ( .A(n25543), .B(n25542), .Z(n25544) );
  NAND U26266 ( .A(n25545), .B(n25544), .Z(n25779) );
  XNOR U26267 ( .A(n25778), .B(n25779), .Z(n25780) );
  XOR U26268 ( .A(n25781), .B(n25780), .Z(n25892) );
  XNOR U26269 ( .A(n25893), .B(n25892), .Z(n25886) );
  NANDN U26270 ( .A(n25547), .B(n25546), .Z(n25551) );
  NAND U26271 ( .A(n25549), .B(n25548), .Z(n25550) );
  NAND U26272 ( .A(n25551), .B(n25550), .Z(n25896) );
  NANDN U26273 ( .A(n25553), .B(n25552), .Z(n25557) );
  NAND U26274 ( .A(n25555), .B(n25554), .Z(n25556) );
  NAND U26275 ( .A(n25557), .B(n25556), .Z(n25897) );
  XNOR U26276 ( .A(n25896), .B(n25897), .Z(n25898) );
  NANDN U26277 ( .A(n25559), .B(n25558), .Z(n25563) );
  NAND U26278 ( .A(n25561), .B(n25560), .Z(n25562) );
  NAND U26279 ( .A(n25563), .B(n25562), .Z(n25723) );
  XNOR U26280 ( .A(a[103]), .B(b[15]), .Z(n25732) );
  OR U26281 ( .A(n25732), .B(n32010), .Z(n25566) );
  NANDN U26282 ( .A(n25564), .B(n32011), .Z(n25565) );
  NAND U26283 ( .A(n25566), .B(n25565), .Z(n25827) );
  XNOR U26284 ( .A(n35377), .B(b[25]), .Z(n25735) );
  NANDN U26285 ( .A(n34219), .B(n25735), .Z(n25569) );
  NAND U26286 ( .A(n34217), .B(n25567), .Z(n25568) );
  NAND U26287 ( .A(n25569), .B(n25568), .Z(n25824) );
  XOR U26288 ( .A(a[101]), .B(b[17]), .Z(n25738) );
  NAND U26289 ( .A(n25738), .B(n32543), .Z(n25572) );
  NANDN U26290 ( .A(n25570), .B(n32541), .Z(n25571) );
  AND U26291 ( .A(n25572), .B(n25571), .Z(n25825) );
  XNOR U26292 ( .A(n25824), .B(n25825), .Z(n25826) );
  XOR U26293 ( .A(n25827), .B(n25826), .Z(n25882) );
  XNOR U26294 ( .A(b[39]), .B(a[79]), .Z(n25741) );
  NANDN U26295 ( .A(n25741), .B(n36553), .Z(n25575) );
  NANDN U26296 ( .A(n25573), .B(n36643), .Z(n25574) );
  NAND U26297 ( .A(n25575), .B(n25574), .Z(n25821) );
  XOR U26298 ( .A(b[51]), .B(n29372), .Z(n25744) );
  NANDN U26299 ( .A(n25744), .B(n37803), .Z(n25578) );
  NANDN U26300 ( .A(n25576), .B(n37802), .Z(n25577) );
  NAND U26301 ( .A(n25578), .B(n25577), .Z(n25818) );
  XOR U26302 ( .A(b[53]), .B(n28403), .Z(n25747) );
  NANDN U26303 ( .A(n25747), .B(n37940), .Z(n25581) );
  NANDN U26304 ( .A(n25579), .B(n37941), .Z(n25580) );
  AND U26305 ( .A(n25581), .B(n25580), .Z(n25819) );
  XNOR U26306 ( .A(n25818), .B(n25819), .Z(n25820) );
  XOR U26307 ( .A(n25821), .B(n25820), .Z(n25883) );
  XNOR U26308 ( .A(n25882), .B(n25883), .Z(n25885) );
  NANDN U26309 ( .A(n25583), .B(n25582), .Z(n25587) );
  NAND U26310 ( .A(n25585), .B(n25584), .Z(n25586) );
  AND U26311 ( .A(n25587), .B(n25586), .Z(n25884) );
  XNOR U26312 ( .A(n25885), .B(n25884), .Z(n25720) );
  NANDN U26313 ( .A(n25589), .B(n25588), .Z(n25593) );
  NAND U26314 ( .A(n25591), .B(n25590), .Z(n25592) );
  AND U26315 ( .A(n25593), .B(n25592), .Z(n25721) );
  XOR U26316 ( .A(n25720), .B(n25721), .Z(n25722) );
  XOR U26317 ( .A(n25723), .B(n25722), .Z(n25899) );
  XNOR U26318 ( .A(n25898), .B(n25899), .Z(n25887) );
  XOR U26319 ( .A(n25886), .B(n25887), .Z(n25888) );
  XOR U26320 ( .A(n25889), .B(n25888), .Z(n25660) );
  XNOR U26321 ( .A(n25659), .B(n25660), .Z(n25661) );
  XNOR U26322 ( .A(n25662), .B(n25661), .Z(n25650) );
  XOR U26323 ( .A(n25649), .B(n25650), .Z(n25644) );
  OR U26324 ( .A(n25595), .B(n25594), .Z(n25599) );
  NAND U26325 ( .A(n25597), .B(n25596), .Z(n25598) );
  NAND U26326 ( .A(n25599), .B(n25598), .Z(n25641) );
  NANDN U26327 ( .A(n25601), .B(n25600), .Z(n25605) );
  NANDN U26328 ( .A(n25603), .B(n25602), .Z(n25604) );
  NAND U26329 ( .A(n25605), .B(n25604), .Z(n25642) );
  XNOR U26330 ( .A(n25641), .B(n25642), .Z(n25643) );
  XNOR U26331 ( .A(n25644), .B(n25643), .Z(n25635) );
  OR U26332 ( .A(n25607), .B(n25606), .Z(n25611) );
  NAND U26333 ( .A(n25609), .B(n25608), .Z(n25610) );
  AND U26334 ( .A(n25611), .B(n25610), .Z(n25636) );
  XOR U26335 ( .A(n25635), .B(n25636), .Z(n25638) );
  NANDN U26336 ( .A(n25613), .B(n25612), .Z(n25617) );
  NANDN U26337 ( .A(n25615), .B(n25614), .Z(n25616) );
  NAND U26338 ( .A(n25617), .B(n25616), .Z(n25637) );
  XNOR U26339 ( .A(n25638), .B(n25637), .Z(n25629) );
  NAND U26340 ( .A(n25619), .B(n25618), .Z(n25623) );
  NANDN U26341 ( .A(n25621), .B(n25620), .Z(n25622) );
  AND U26342 ( .A(n25623), .B(n25622), .Z(n25630) );
  XNOR U26343 ( .A(n25629), .B(n25630), .Z(n25631) );
  XNOR U26344 ( .A(n25632), .B(n25631), .Z(n25908) );
  XNOR U26345 ( .A(n25908), .B(sreg[181]), .Z(n25910) );
  NAND U26346 ( .A(n25624), .B(sreg[180]), .Z(n25628) );
  OR U26347 ( .A(n25626), .B(n25625), .Z(n25627) );
  AND U26348 ( .A(n25628), .B(n25627), .Z(n25909) );
  XOR U26349 ( .A(n25910), .B(n25909), .Z(c[181]) );
  NANDN U26350 ( .A(n25630), .B(n25629), .Z(n25634) );
  NAND U26351 ( .A(n25632), .B(n25631), .Z(n25633) );
  NAND U26352 ( .A(n25634), .B(n25633), .Z(n25916) );
  NANDN U26353 ( .A(n25636), .B(n25635), .Z(n25640) );
  OR U26354 ( .A(n25638), .B(n25637), .Z(n25639) );
  NAND U26355 ( .A(n25640), .B(n25639), .Z(n25913) );
  NANDN U26356 ( .A(n25642), .B(n25641), .Z(n25646) );
  NAND U26357 ( .A(n25644), .B(n25643), .Z(n25645) );
  NAND U26358 ( .A(n25646), .B(n25645), .Z(n26195) );
  OR U26359 ( .A(n25648), .B(n25647), .Z(n25652) );
  NANDN U26360 ( .A(n25650), .B(n25649), .Z(n25651) );
  NAND U26361 ( .A(n25652), .B(n25651), .Z(n26193) );
  NANDN U26362 ( .A(n25654), .B(n25653), .Z(n25658) );
  NANDN U26363 ( .A(n25656), .B(n25655), .Z(n25657) );
  NAND U26364 ( .A(n25658), .B(n25657), .Z(n26187) );
  XNOR U26365 ( .A(n26187), .B(n26186), .Z(n26188) );
  NANDN U26366 ( .A(n25664), .B(n25663), .Z(n25668) );
  NAND U26367 ( .A(n25666), .B(n25665), .Z(n25667) );
  NAND U26368 ( .A(n25668), .B(n25667), .Z(n26176) );
  NANDN U26369 ( .A(n25670), .B(n25669), .Z(n25674) );
  NANDN U26370 ( .A(n25672), .B(n25671), .Z(n25673) );
  NAND U26371 ( .A(n25674), .B(n25673), .Z(n26151) );
  XOR U26372 ( .A(a[108]), .B(n970), .Z(n25946) );
  OR U26373 ( .A(n25946), .B(n31369), .Z(n25677) );
  NANDN U26374 ( .A(n25675), .B(n31119), .Z(n25676) );
  NAND U26375 ( .A(n25677), .B(n25676), .Z(n25967) );
  XOR U26376 ( .A(b[43]), .B(n31363), .Z(n25949) );
  NANDN U26377 ( .A(n25949), .B(n37068), .Z(n25680) );
  NANDN U26378 ( .A(n25678), .B(n37069), .Z(n25679) );
  NAND U26379 ( .A(n25680), .B(n25679), .Z(n25964) );
  XNOR U26380 ( .A(b[45]), .B(a[74]), .Z(n25952) );
  NANDN U26381 ( .A(n25952), .B(n37261), .Z(n25683) );
  NAND U26382 ( .A(n25681), .B(n37262), .Z(n25682) );
  AND U26383 ( .A(n25683), .B(n25682), .Z(n25965) );
  XNOR U26384 ( .A(n25964), .B(n25965), .Z(n25966) );
  XNOR U26385 ( .A(n25967), .B(n25966), .Z(n26055) );
  XOR U26386 ( .A(n979), .B(n30379), .Z(n25955) );
  NANDN U26387 ( .A(n37756), .B(n25955), .Z(n25686) );
  NANDN U26388 ( .A(n25684), .B(n37652), .Z(n25685) );
  NAND U26389 ( .A(n25686), .B(n25685), .Z(n25942) );
  NAND U26390 ( .A(n37469), .B(n25687), .Z(n25689) );
  XOR U26391 ( .A(b[47]), .B(n30210), .Z(n25958) );
  NANDN U26392 ( .A(n25958), .B(n37471), .Z(n25688) );
  AND U26393 ( .A(n25689), .B(n25688), .Z(n25940) );
  XOR U26394 ( .A(n37336), .B(n969), .Z(n25961) );
  NAND U26395 ( .A(n30509), .B(n25961), .Z(n25692) );
  NANDN U26396 ( .A(n25690), .B(n30846), .Z(n25691) );
  AND U26397 ( .A(n25692), .B(n25691), .Z(n25941) );
  XOR U26398 ( .A(n25942), .B(n25943), .Z(n26052) );
  NANDN U26399 ( .A(n25694), .B(n25693), .Z(n25698) );
  NAND U26400 ( .A(n25696), .B(n25695), .Z(n25697) );
  NAND U26401 ( .A(n25698), .B(n25697), .Z(n26053) );
  XNOR U26402 ( .A(n26052), .B(n26053), .Z(n26054) );
  XOR U26403 ( .A(n26055), .B(n26054), .Z(n26150) );
  XNOR U26404 ( .A(n26151), .B(n26150), .Z(n26153) );
  XNOR U26405 ( .A(b[35]), .B(a[84]), .Z(n25925) );
  NANDN U26406 ( .A(n25925), .B(n35985), .Z(n25701) );
  NAND U26407 ( .A(n25699), .B(n35986), .Z(n25700) );
  NAND U26408 ( .A(n25701), .B(n25700), .Z(n26001) );
  XOR U26409 ( .A(n37583), .B(n31123), .Z(n25928) );
  NAND U26410 ( .A(n25928), .B(n29949), .Z(n25704) );
  NAND U26411 ( .A(n29948), .B(n25702), .Z(n25703) );
  NAND U26412 ( .A(n25704), .B(n25703), .Z(n25998) );
  XNOR U26413 ( .A(b[55]), .B(a[64]), .Z(n25931) );
  NANDN U26414 ( .A(n25931), .B(n38075), .Z(n25707) );
  NANDN U26415 ( .A(n25705), .B(n38073), .Z(n25706) );
  AND U26416 ( .A(n25707), .B(n25706), .Z(n25999) );
  XNOR U26417 ( .A(n25998), .B(n25999), .Z(n26000) );
  XNOR U26418 ( .A(n26001), .B(n26000), .Z(n26031) );
  NANDN U26419 ( .A(n25709), .B(n25708), .Z(n25713) );
  NAND U26420 ( .A(n25711), .B(n25710), .Z(n25712) );
  NAND U26421 ( .A(n25713), .B(n25712), .Z(n26028) );
  NANDN U26422 ( .A(n25715), .B(n25714), .Z(n25719) );
  NAND U26423 ( .A(n25717), .B(n25716), .Z(n25718) );
  NAND U26424 ( .A(n25719), .B(n25718), .Z(n26029) );
  XNOR U26425 ( .A(n26028), .B(n26029), .Z(n26030) );
  XOR U26426 ( .A(n26031), .B(n26030), .Z(n26152) );
  XOR U26427 ( .A(n26153), .B(n26152), .Z(n26144) );
  NAND U26428 ( .A(n25721), .B(n25720), .Z(n25725) );
  NANDN U26429 ( .A(n25723), .B(n25722), .Z(n25724) );
  NAND U26430 ( .A(n25725), .B(n25724), .Z(n26159) );
  NANDN U26431 ( .A(n25727), .B(n25726), .Z(n25731) );
  NANDN U26432 ( .A(n25729), .B(n25728), .Z(n25730) );
  NAND U26433 ( .A(n25731), .B(n25730), .Z(n26156) );
  XOR U26434 ( .A(a[104]), .B(n972), .Z(n25974) );
  OR U26435 ( .A(n25974), .B(n32010), .Z(n25734) );
  NANDN U26436 ( .A(n25732), .B(n32011), .Z(n25733) );
  NAND U26437 ( .A(n25734), .B(n25733), .Z(n26068) );
  XNOR U26438 ( .A(n35191), .B(b[25]), .Z(n25977) );
  NANDN U26439 ( .A(n34219), .B(n25977), .Z(n25737) );
  NAND U26440 ( .A(n34217), .B(n25735), .Z(n25736) );
  NAND U26441 ( .A(n25737), .B(n25736), .Z(n26065) );
  XNOR U26442 ( .A(a[102]), .B(b[17]), .Z(n25980) );
  NANDN U26443 ( .A(n25980), .B(n32543), .Z(n25740) );
  NAND U26444 ( .A(n25738), .B(n32541), .Z(n25739) );
  AND U26445 ( .A(n25740), .B(n25739), .Z(n26066) );
  XNOR U26446 ( .A(n26065), .B(n26066), .Z(n26067) );
  XNOR U26447 ( .A(n26068), .B(n26067), .Z(n26138) );
  XOR U26448 ( .A(b[39]), .B(n32814), .Z(n25983) );
  NANDN U26449 ( .A(n25983), .B(n36553), .Z(n25743) );
  NANDN U26450 ( .A(n25741), .B(n36643), .Z(n25742) );
  NAND U26451 ( .A(n25743), .B(n25742), .Z(n26098) );
  XOR U26452 ( .A(b[51]), .B(n29868), .Z(n25986) );
  NANDN U26453 ( .A(n25986), .B(n37803), .Z(n25746) );
  NANDN U26454 ( .A(n25744), .B(n37802), .Z(n25745) );
  NAND U26455 ( .A(n25746), .B(n25745), .Z(n26095) );
  XOR U26456 ( .A(b[53]), .B(n28701), .Z(n25989) );
  NANDN U26457 ( .A(n25989), .B(n37940), .Z(n25749) );
  NANDN U26458 ( .A(n25747), .B(n37941), .Z(n25748) );
  AND U26459 ( .A(n25749), .B(n25748), .Z(n26096) );
  XNOR U26460 ( .A(n26095), .B(n26096), .Z(n26097) );
  XOR U26461 ( .A(n26098), .B(n26097), .Z(n26139) );
  XNOR U26462 ( .A(n26138), .B(n26139), .Z(n26140) );
  NANDN U26463 ( .A(n25751), .B(n25750), .Z(n25755) );
  NAND U26464 ( .A(n25753), .B(n25752), .Z(n25754) );
  NAND U26465 ( .A(n25755), .B(n25754), .Z(n26141) );
  XOR U26466 ( .A(n26140), .B(n26141), .Z(n26019) );
  NANDN U26467 ( .A(n25757), .B(n25756), .Z(n25761) );
  NAND U26468 ( .A(n25759), .B(n25758), .Z(n25760) );
  NAND U26469 ( .A(n25761), .B(n25760), .Z(n26016) );
  XNOR U26470 ( .A(n26016), .B(n26017), .Z(n26018) );
  XOR U26471 ( .A(n26019), .B(n26018), .Z(n26157) );
  XNOR U26472 ( .A(n26156), .B(n26157), .Z(n26158) );
  XOR U26473 ( .A(n26159), .B(n26158), .Z(n26145) );
  XNOR U26474 ( .A(n26144), .B(n26145), .Z(n26146) );
  NAND U26475 ( .A(n25767), .B(n25766), .Z(n25771) );
  NANDN U26476 ( .A(n25769), .B(n25768), .Z(n25770) );
  NAND U26477 ( .A(n25771), .B(n25770), .Z(n26147) );
  XOR U26478 ( .A(n26146), .B(n26147), .Z(n26175) );
  NANDN U26479 ( .A(n25773), .B(n25772), .Z(n25777) );
  NANDN U26480 ( .A(n25775), .B(n25774), .Z(n25776) );
  NAND U26481 ( .A(n25777), .B(n25776), .Z(n25919) );
  NANDN U26482 ( .A(n25779), .B(n25778), .Z(n25783) );
  NAND U26483 ( .A(n25781), .B(n25780), .Z(n25782) );
  NAND U26484 ( .A(n25783), .B(n25782), .Z(n26164) );
  NAND U26485 ( .A(n25785), .B(n25784), .Z(n25789) );
  NANDN U26486 ( .A(n25787), .B(n25786), .Z(n25788) );
  AND U26487 ( .A(n25789), .B(n25788), .Z(n26162) );
  NANDN U26488 ( .A(n25791), .B(n25790), .Z(n25795) );
  NAND U26489 ( .A(n25793), .B(n25792), .Z(n25794) );
  AND U26490 ( .A(n25795), .B(n25794), .Z(n26163) );
  XOR U26491 ( .A(n26164), .B(n26165), .Z(n25920) );
  XOR U26492 ( .A(n25919), .B(n25920), .Z(n25921) );
  XOR U26493 ( .A(b[37]), .B(n32815), .Z(n26077) );
  NANDN U26494 ( .A(n26077), .B(n36311), .Z(n25802) );
  NANDN U26495 ( .A(n25800), .B(n36309), .Z(n25801) );
  NAND U26496 ( .A(n25802), .B(n25801), .Z(n26135) );
  XOR U26497 ( .A(a[114]), .B(n968), .Z(n26080) );
  OR U26498 ( .A(n26080), .B(n29363), .Z(n25805) );
  NANDN U26499 ( .A(n25803), .B(n29864), .Z(n25804) );
  NAND U26500 ( .A(n25805), .B(n25804), .Z(n26132) );
  XOR U26501 ( .A(n38046), .B(n967), .Z(n26083) );
  NAND U26502 ( .A(n26083), .B(n28939), .Z(n25808) );
  NAND U26503 ( .A(n28938), .B(n25806), .Z(n25807) );
  AND U26504 ( .A(n25808), .B(n25807), .Z(n26133) );
  XNOR U26505 ( .A(n26132), .B(n26133), .Z(n26134) );
  XNOR U26506 ( .A(n26135), .B(n26134), .Z(n26034) );
  XOR U26507 ( .A(a[106]), .B(n971), .Z(n26086) );
  OR U26508 ( .A(n26086), .B(n31550), .Z(n25811) );
  NANDN U26509 ( .A(n25809), .B(n31874), .Z(n25810) );
  NAND U26510 ( .A(n25811), .B(n25810), .Z(n25995) );
  NAND U26511 ( .A(n34848), .B(n25812), .Z(n25814) );
  XOR U26512 ( .A(n35375), .B(n34852), .Z(n26089) );
  NAND U26513 ( .A(n34618), .B(n26089), .Z(n25813) );
  NAND U26514 ( .A(n25814), .B(n25813), .Z(n25992) );
  NAND U26515 ( .A(n35188), .B(n25815), .Z(n25817) );
  XOR U26516 ( .A(n35540), .B(n34851), .Z(n26092) );
  NANDN U26517 ( .A(n34968), .B(n26092), .Z(n25816) );
  AND U26518 ( .A(n25817), .B(n25816), .Z(n25993) );
  XNOR U26519 ( .A(n25992), .B(n25993), .Z(n25994) );
  XOR U26520 ( .A(n25995), .B(n25994), .Z(n26035) );
  XOR U26521 ( .A(n26034), .B(n26035), .Z(n26037) );
  NANDN U26522 ( .A(n25819), .B(n25818), .Z(n25823) );
  NAND U26523 ( .A(n25821), .B(n25820), .Z(n25822) );
  NAND U26524 ( .A(n25823), .B(n25822), .Z(n26036) );
  XNOR U26525 ( .A(n26037), .B(n26036), .Z(n26047) );
  NANDN U26526 ( .A(n25825), .B(n25824), .Z(n25829) );
  NAND U26527 ( .A(n25827), .B(n25826), .Z(n25828) );
  NAND U26528 ( .A(n25829), .B(n25828), .Z(n25972) );
  NAND U26529 ( .A(a[54]), .B(b[63]), .Z(n25937) );
  NANDN U26530 ( .A(n25830), .B(n38369), .Z(n25832) );
  XOR U26531 ( .A(b[61]), .B(n26347), .Z(n26071) );
  OR U26532 ( .A(n26071), .B(n38371), .Z(n25831) );
  NAND U26533 ( .A(n25832), .B(n25831), .Z(n25935) );
  NANDN U26534 ( .A(n25833), .B(n35311), .Z(n25835) );
  XOR U26535 ( .A(b[31]), .B(n34048), .Z(n26074) );
  NANDN U26536 ( .A(n26074), .B(n35313), .Z(n25834) );
  AND U26537 ( .A(n25835), .B(n25834), .Z(n25934) );
  XNOR U26538 ( .A(n25935), .B(n25934), .Z(n25936) );
  XOR U26539 ( .A(n25937), .B(n25936), .Z(n25970) );
  NAND U26540 ( .A(n33283), .B(n25836), .Z(n25838) );
  XOR U26541 ( .A(n36100), .B(n33020), .Z(n26056) );
  NANDN U26542 ( .A(n33021), .B(n26056), .Z(n25837) );
  NAND U26543 ( .A(n25838), .B(n25837), .Z(n26104) );
  XNOR U26544 ( .A(a[98]), .B(b[21]), .Z(n26059) );
  OR U26545 ( .A(n26059), .B(n33634), .Z(n25841) );
  NAND U26546 ( .A(n25839), .B(n33464), .Z(n25840) );
  NAND U26547 ( .A(n25841), .B(n25840), .Z(n26101) );
  NAND U26548 ( .A(n34044), .B(n25842), .Z(n25844) );
  XOR U26549 ( .A(n35545), .B(n34510), .Z(n26062) );
  NANDN U26550 ( .A(n33867), .B(n26062), .Z(n25843) );
  AND U26551 ( .A(n25844), .B(n25843), .Z(n26102) );
  XNOR U26552 ( .A(n26101), .B(n26102), .Z(n26103) );
  XNOR U26553 ( .A(n26104), .B(n26103), .Z(n25971) );
  XNOR U26554 ( .A(n25970), .B(n25971), .Z(n25973) );
  XNOR U26555 ( .A(n25972), .B(n25973), .Z(n26046) );
  XNOR U26556 ( .A(n26047), .B(n26046), .Z(n26048) );
  XNOR U26557 ( .A(n26049), .B(n26048), .Z(n26025) );
  XNOR U26558 ( .A(b[41]), .B(a[78]), .Z(n26107) );
  OR U26559 ( .A(n26107), .B(n36905), .Z(n25847) );
  NAND U26560 ( .A(n25845), .B(n36807), .Z(n25846) );
  NAND U26561 ( .A(n25847), .B(n25846), .Z(n26129) );
  XNOR U26562 ( .A(b[57]), .B(a[62]), .Z(n26110) );
  OR U26563 ( .A(n26110), .B(n965), .Z(n25850) );
  NANDN U26564 ( .A(n25848), .B(n38194), .Z(n25849) );
  NAND U26565 ( .A(n25850), .B(n25849), .Z(n26126) );
  NAND U26566 ( .A(n38326), .B(n25851), .Z(n25853) );
  XOR U26567 ( .A(n38400), .B(n27436), .Z(n26113) );
  NANDN U26568 ( .A(n38273), .B(n26113), .Z(n25852) );
  AND U26569 ( .A(n25853), .B(n25852), .Z(n26127) );
  XNOR U26570 ( .A(n26126), .B(n26127), .Z(n26128) );
  XOR U26571 ( .A(n26129), .B(n26128), .Z(n26010) );
  XOR U26572 ( .A(b[33]), .B(n33628), .Z(n26116) );
  NANDN U26573 ( .A(n26116), .B(n35620), .Z(n25856) );
  NANDN U26574 ( .A(n25854), .B(n35621), .Z(n25855) );
  NAND U26575 ( .A(n25856), .B(n25855), .Z(n26007) );
  NANDN U26576 ( .A(n966), .B(a[118]), .Z(n25857) );
  XOR U26577 ( .A(n29232), .B(n25857), .Z(n25859) );
  NANDN U26578 ( .A(b[0]), .B(a[117]), .Z(n25858) );
  AND U26579 ( .A(n25859), .B(n25858), .Z(n26004) );
  XOR U26580 ( .A(b[63]), .B(n25860), .Z(n26123) );
  NANDN U26581 ( .A(n26123), .B(n38422), .Z(n25863) );
  NANDN U26582 ( .A(n25861), .B(n38423), .Z(n25862) );
  AND U26583 ( .A(n25863), .B(n25862), .Z(n26005) );
  XNOR U26584 ( .A(n26004), .B(n26005), .Z(n26006) );
  XOR U26585 ( .A(n26007), .B(n26006), .Z(n26011) );
  XNOR U26586 ( .A(n26010), .B(n26011), .Z(n26013) );
  NANDN U26587 ( .A(n25865), .B(n25864), .Z(n25869) );
  NAND U26588 ( .A(n25867), .B(n25866), .Z(n25868) );
  NAND U26589 ( .A(n25869), .B(n25868), .Z(n26012) );
  XNOR U26590 ( .A(n26013), .B(n26012), .Z(n26043) );
  NANDN U26591 ( .A(n25871), .B(n25870), .Z(n25875) );
  NAND U26592 ( .A(n25873), .B(n25872), .Z(n25874) );
  NAND U26593 ( .A(n25875), .B(n25874), .Z(n26040) );
  NANDN U26594 ( .A(n25877), .B(n25876), .Z(n25881) );
  NAND U26595 ( .A(n25879), .B(n25878), .Z(n25880) );
  AND U26596 ( .A(n25881), .B(n25880), .Z(n26041) );
  XNOR U26597 ( .A(n26040), .B(n26041), .Z(n26042) );
  XOR U26598 ( .A(n26043), .B(n26042), .Z(n26023) );
  XOR U26599 ( .A(n26023), .B(n26022), .Z(n26024) );
  XOR U26600 ( .A(n26025), .B(n26024), .Z(n25922) );
  XOR U26601 ( .A(n25921), .B(n25922), .Z(n26174) );
  XNOR U26602 ( .A(n26175), .B(n26174), .Z(n26177) );
  XNOR U26603 ( .A(n26176), .B(n26177), .Z(n26182) );
  NAND U26604 ( .A(n25891), .B(n25890), .Z(n25895) );
  NANDN U26605 ( .A(n25893), .B(n25892), .Z(n25894) );
  NAND U26606 ( .A(n25895), .B(n25894), .Z(n26171) );
  NANDN U26607 ( .A(n25897), .B(n25896), .Z(n25901) );
  NANDN U26608 ( .A(n25899), .B(n25898), .Z(n25900) );
  NAND U26609 ( .A(n25901), .B(n25900), .Z(n26168) );
  NANDN U26610 ( .A(n25903), .B(n25902), .Z(n25907) );
  NAND U26611 ( .A(n25905), .B(n25904), .Z(n25906) );
  AND U26612 ( .A(n25907), .B(n25906), .Z(n26169) );
  XNOR U26613 ( .A(n26168), .B(n26169), .Z(n26170) );
  XNOR U26614 ( .A(n26171), .B(n26170), .Z(n26181) );
  XNOR U26615 ( .A(n26180), .B(n26181), .Z(n26183) );
  XOR U26616 ( .A(n26182), .B(n26183), .Z(n26189) );
  XOR U26617 ( .A(n26188), .B(n26189), .Z(n26192) );
  XNOR U26618 ( .A(n26193), .B(n26192), .Z(n26194) );
  XNOR U26619 ( .A(n26195), .B(n26194), .Z(n25914) );
  XOR U26620 ( .A(n25913), .B(n25914), .Z(n25915) );
  XNOR U26621 ( .A(n25916), .B(n25915), .Z(n26196) );
  XNOR U26622 ( .A(n26196), .B(sreg[182]), .Z(n26198) );
  NAND U26623 ( .A(n25908), .B(sreg[181]), .Z(n25912) );
  OR U26624 ( .A(n25910), .B(n25909), .Z(n25911) );
  AND U26625 ( .A(n25912), .B(n25911), .Z(n26197) );
  XOR U26626 ( .A(n26198), .B(n26197), .Z(c[182]) );
  OR U26627 ( .A(n25914), .B(n25913), .Z(n25918) );
  NAND U26628 ( .A(n25916), .B(n25915), .Z(n25917) );
  NAND U26629 ( .A(n25918), .B(n25917), .Z(n26204) );
  OR U26630 ( .A(n25920), .B(n25919), .Z(n25924) );
  NAND U26631 ( .A(n25922), .B(n25921), .Z(n25923) );
  NAND U26632 ( .A(n25924), .B(n25923), .Z(n26210) );
  XOR U26633 ( .A(b[35]), .B(a[85]), .Z(n26391) );
  NAND U26634 ( .A(n35985), .B(n26391), .Z(n25927) );
  NANDN U26635 ( .A(n25925), .B(n35986), .Z(n25926) );
  NAND U26636 ( .A(n25927), .B(n25926), .Z(n26437) );
  XNOR U26637 ( .A(a[113]), .B(n31123), .Z(n26394) );
  NAND U26638 ( .A(n26394), .B(n29949), .Z(n25930) );
  NAND U26639 ( .A(n29948), .B(n25928), .Z(n25929) );
  NAND U26640 ( .A(n25930), .B(n25929), .Z(n26434) );
  XOR U26641 ( .A(b[55]), .B(n28403), .Z(n26397) );
  NANDN U26642 ( .A(n26397), .B(n38075), .Z(n25933) );
  NANDN U26643 ( .A(n25931), .B(n38073), .Z(n25932) );
  AND U26644 ( .A(n25933), .B(n25932), .Z(n26435) );
  XNOR U26645 ( .A(n26434), .B(n26435), .Z(n26436) );
  XNOR U26646 ( .A(n26437), .B(n26436), .Z(n26248) );
  NANDN U26647 ( .A(n25935), .B(n25934), .Z(n25939) );
  NAND U26648 ( .A(n25937), .B(n25936), .Z(n25938) );
  NAND U26649 ( .A(n25939), .B(n25938), .Z(n26245) );
  OR U26650 ( .A(n25941), .B(n25940), .Z(n25945) );
  NANDN U26651 ( .A(n25943), .B(n25942), .Z(n25944) );
  NAND U26652 ( .A(n25945), .B(n25944), .Z(n26246) );
  XNOR U26653 ( .A(n26245), .B(n26246), .Z(n26247) );
  XOR U26654 ( .A(n26248), .B(n26247), .Z(n26225) );
  XNOR U26655 ( .A(a[109]), .B(b[11]), .Z(n26367) );
  OR U26656 ( .A(n26367), .B(n31369), .Z(n25948) );
  NANDN U26657 ( .A(n25946), .B(n31119), .Z(n25947) );
  NAND U26658 ( .A(n25948), .B(n25947), .Z(n26388) );
  XNOR U26659 ( .A(b[43]), .B(a[77]), .Z(n26370) );
  NANDN U26660 ( .A(n26370), .B(n37068), .Z(n25951) );
  NANDN U26661 ( .A(n25949), .B(n37069), .Z(n25950) );
  NAND U26662 ( .A(n25951), .B(n25950), .Z(n26385) );
  XOR U26663 ( .A(b[45]), .B(a[75]), .Z(n26373) );
  NAND U26664 ( .A(n26373), .B(n37261), .Z(n25954) );
  NANDN U26665 ( .A(n25952), .B(n37262), .Z(n25953) );
  AND U26666 ( .A(n25954), .B(n25953), .Z(n26386) );
  XNOR U26667 ( .A(n26385), .B(n26386), .Z(n26387) );
  XNOR U26668 ( .A(n26388), .B(n26387), .Z(n26266) );
  NAND U26669 ( .A(n37652), .B(n25955), .Z(n25957) );
  XOR U26670 ( .A(b[49]), .B(n30543), .Z(n26376) );
  OR U26671 ( .A(n26376), .B(n37756), .Z(n25956) );
  NAND U26672 ( .A(n25957), .B(n25956), .Z(n26408) );
  NANDN U26673 ( .A(n25958), .B(n37469), .Z(n25960) );
  XNOR U26674 ( .A(n978), .B(a[73]), .Z(n26379) );
  NAND U26675 ( .A(n26379), .B(n37471), .Z(n25959) );
  NAND U26676 ( .A(n25960), .B(n25959), .Z(n26406) );
  NAND U26677 ( .A(n30846), .B(n25961), .Z(n25963) );
  XNOR U26678 ( .A(a[111]), .B(n969), .Z(n26382) );
  NAND U26679 ( .A(n30509), .B(n26382), .Z(n25962) );
  NAND U26680 ( .A(n25963), .B(n25962), .Z(n26407) );
  XNOR U26681 ( .A(n26406), .B(n26407), .Z(n26409) );
  XOR U26682 ( .A(n26408), .B(n26409), .Z(n26263) );
  NANDN U26683 ( .A(n25965), .B(n25964), .Z(n25969) );
  NAND U26684 ( .A(n25967), .B(n25966), .Z(n25968) );
  NAND U26685 ( .A(n25969), .B(n25968), .Z(n26264) );
  XNOR U26686 ( .A(n26263), .B(n26264), .Z(n26265) );
  XOR U26687 ( .A(n26266), .B(n26265), .Z(n26223) );
  XOR U26688 ( .A(n26223), .B(n26224), .Z(n26226) );
  XNOR U26689 ( .A(n26225), .B(n26226), .Z(n26217) );
  XNOR U26690 ( .A(a[105]), .B(b[15]), .Z(n26416) );
  OR U26691 ( .A(n26416), .B(n32010), .Z(n25976) );
  NANDN U26692 ( .A(n25974), .B(n32011), .Z(n25975) );
  NAND U26693 ( .A(n25976), .B(n25975), .Z(n26296) );
  XNOR U26694 ( .A(n35628), .B(b[25]), .Z(n26419) );
  NANDN U26695 ( .A(n34219), .B(n26419), .Z(n25979) );
  NAND U26696 ( .A(n34217), .B(n25977), .Z(n25978) );
  NAND U26697 ( .A(n25979), .B(n25978), .Z(n26293) );
  XOR U26698 ( .A(a[103]), .B(b[17]), .Z(n26422) );
  NAND U26699 ( .A(n26422), .B(n32543), .Z(n25982) );
  NANDN U26700 ( .A(n25980), .B(n32541), .Z(n25981) );
  AND U26701 ( .A(n25982), .B(n25981), .Z(n26294) );
  XNOR U26702 ( .A(n26293), .B(n26294), .Z(n26295) );
  XNOR U26703 ( .A(n26296), .B(n26295), .Z(n26314) );
  XNOR U26704 ( .A(b[39]), .B(a[81]), .Z(n26425) );
  NANDN U26705 ( .A(n26425), .B(n36553), .Z(n25985) );
  NANDN U26706 ( .A(n25983), .B(n36643), .Z(n25984) );
  NAND U26707 ( .A(n25985), .B(n25984), .Z(n26290) );
  XNOR U26708 ( .A(b[51]), .B(a[69]), .Z(n26428) );
  NANDN U26709 ( .A(n26428), .B(n37803), .Z(n25988) );
  NANDN U26710 ( .A(n25986), .B(n37802), .Z(n25987) );
  NAND U26711 ( .A(n25988), .B(n25987), .Z(n26287) );
  XOR U26712 ( .A(b[53]), .B(n29372), .Z(n26431) );
  NANDN U26713 ( .A(n26431), .B(n37940), .Z(n25991) );
  NANDN U26714 ( .A(n25989), .B(n37941), .Z(n25990) );
  AND U26715 ( .A(n25991), .B(n25990), .Z(n26288) );
  XNOR U26716 ( .A(n26287), .B(n26288), .Z(n26289) );
  XOR U26717 ( .A(n26290), .B(n26289), .Z(n26315) );
  XOR U26718 ( .A(n26314), .B(n26315), .Z(n26317) );
  NANDN U26719 ( .A(n25993), .B(n25992), .Z(n25997) );
  NAND U26720 ( .A(n25995), .B(n25994), .Z(n25996) );
  NAND U26721 ( .A(n25997), .B(n25996), .Z(n26316) );
  XNOR U26722 ( .A(n26317), .B(n26316), .Z(n26455) );
  NANDN U26723 ( .A(n25999), .B(n25998), .Z(n26003) );
  NAND U26724 ( .A(n26001), .B(n26000), .Z(n26002) );
  NAND U26725 ( .A(n26003), .B(n26002), .Z(n26452) );
  NANDN U26726 ( .A(n26005), .B(n26004), .Z(n26009) );
  NAND U26727 ( .A(n26007), .B(n26006), .Z(n26008) );
  AND U26728 ( .A(n26009), .B(n26008), .Z(n26453) );
  XNOR U26729 ( .A(n26452), .B(n26453), .Z(n26454) );
  XNOR U26730 ( .A(n26455), .B(n26454), .Z(n26229) );
  OR U26731 ( .A(n26011), .B(n26010), .Z(n26015) );
  OR U26732 ( .A(n26013), .B(n26012), .Z(n26014) );
  AND U26733 ( .A(n26015), .B(n26014), .Z(n26230) );
  XOR U26734 ( .A(n26229), .B(n26230), .Z(n26232) );
  NANDN U26735 ( .A(n26017), .B(n26016), .Z(n26021) );
  NAND U26736 ( .A(n26019), .B(n26018), .Z(n26020) );
  NAND U26737 ( .A(n26021), .B(n26020), .Z(n26231) );
  XNOR U26738 ( .A(n26232), .B(n26231), .Z(n26218) );
  OR U26739 ( .A(n26023), .B(n26022), .Z(n26027) );
  NAND U26740 ( .A(n26025), .B(n26024), .Z(n26026) );
  AND U26741 ( .A(n26027), .B(n26026), .Z(n26219) );
  XOR U26742 ( .A(n26220), .B(n26219), .Z(n26207) );
  NANDN U26743 ( .A(n26029), .B(n26028), .Z(n26033) );
  NAND U26744 ( .A(n26031), .B(n26030), .Z(n26032) );
  AND U26745 ( .A(n26033), .B(n26032), .Z(n26238) );
  NANDN U26746 ( .A(n26035), .B(n26034), .Z(n26039) );
  OR U26747 ( .A(n26037), .B(n26036), .Z(n26038) );
  NAND U26748 ( .A(n26039), .B(n26038), .Z(n26235) );
  NANDN U26749 ( .A(n26041), .B(n26040), .Z(n26045) );
  NAND U26750 ( .A(n26043), .B(n26042), .Z(n26044) );
  NAND U26751 ( .A(n26045), .B(n26044), .Z(n26236) );
  XNOR U26752 ( .A(n26235), .B(n26236), .Z(n26237) );
  XNOR U26753 ( .A(n26238), .B(n26237), .Z(n26458) );
  NAND U26754 ( .A(n26047), .B(n26046), .Z(n26051) );
  OR U26755 ( .A(n26049), .B(n26048), .Z(n26050) );
  AND U26756 ( .A(n26051), .B(n26050), .Z(n26459) );
  XNOR U26757 ( .A(n26458), .B(n26459), .Z(n26460) );
  NAND U26758 ( .A(n33283), .B(n26056), .Z(n26058) );
  XNOR U26759 ( .A(a[101]), .B(n33020), .Z(n26305) );
  NANDN U26760 ( .A(n33021), .B(n26305), .Z(n26057) );
  NAND U26761 ( .A(n26058), .B(n26057), .Z(n26329) );
  XOR U26762 ( .A(a[99]), .B(b[21]), .Z(n26308) );
  NANDN U26763 ( .A(n33634), .B(n26308), .Z(n26061) );
  NANDN U26764 ( .A(n26059), .B(n33464), .Z(n26060) );
  NAND U26765 ( .A(n26061), .B(n26060), .Z(n26326) );
  NAND U26766 ( .A(n34044), .B(n26062), .Z(n26064) );
  XNOR U26767 ( .A(a[97]), .B(n34510), .Z(n26311) );
  NANDN U26768 ( .A(n33867), .B(n26311), .Z(n26063) );
  AND U26769 ( .A(n26064), .B(n26063), .Z(n26327) );
  XNOR U26770 ( .A(n26326), .B(n26327), .Z(n26328) );
  XNOR U26771 ( .A(n26329), .B(n26328), .Z(n26361) );
  NANDN U26772 ( .A(n26066), .B(n26065), .Z(n26070) );
  NAND U26773 ( .A(n26068), .B(n26067), .Z(n26069) );
  NAND U26774 ( .A(n26070), .B(n26069), .Z(n26362) );
  XNOR U26775 ( .A(n26361), .B(n26362), .Z(n26363) );
  NAND U26776 ( .A(a[55]), .B(b[63]), .Z(n26403) );
  NANDN U26777 ( .A(n26071), .B(n38369), .Z(n26073) );
  XNOR U26778 ( .A(b[61]), .B(a[59]), .Z(n26299) );
  OR U26779 ( .A(n26299), .B(n38371), .Z(n26072) );
  NAND U26780 ( .A(n26073), .B(n26072), .Z(n26401) );
  NANDN U26781 ( .A(n26074), .B(n35311), .Z(n26076) );
  XNOR U26782 ( .A(b[31]), .B(a[89]), .Z(n26302) );
  NANDN U26783 ( .A(n26302), .B(n35313), .Z(n26075) );
  AND U26784 ( .A(n26076), .B(n26075), .Z(n26400) );
  XNOR U26785 ( .A(n26401), .B(n26400), .Z(n26402) );
  XNOR U26786 ( .A(n26403), .B(n26402), .Z(n26364) );
  XOR U26787 ( .A(n26363), .B(n26364), .Z(n26257) );
  XNOR U26788 ( .A(b[37]), .B(a[83]), .Z(n26278) );
  NANDN U26789 ( .A(n26278), .B(n36311), .Z(n26079) );
  NANDN U26790 ( .A(n26077), .B(n36309), .Z(n26078) );
  NAND U26791 ( .A(n26079), .B(n26078), .Z(n26323) );
  XNOR U26792 ( .A(a[115]), .B(b[5]), .Z(n26281) );
  OR U26793 ( .A(n26281), .B(n29363), .Z(n26082) );
  NANDN U26794 ( .A(n26080), .B(n29864), .Z(n26081) );
  NAND U26795 ( .A(n26082), .B(n26081), .Z(n26320) );
  XNOR U26796 ( .A(a[117]), .B(n967), .Z(n26284) );
  NAND U26797 ( .A(n26284), .B(n28939), .Z(n26085) );
  NAND U26798 ( .A(n28938), .B(n26083), .Z(n26084) );
  AND U26799 ( .A(n26085), .B(n26084), .Z(n26321) );
  XNOR U26800 ( .A(n26320), .B(n26321), .Z(n26322) );
  XNOR U26801 ( .A(n26323), .B(n26322), .Z(n26241) );
  XNOR U26802 ( .A(a[107]), .B(b[13]), .Z(n26269) );
  OR U26803 ( .A(n26269), .B(n31550), .Z(n26088) );
  NANDN U26804 ( .A(n26086), .B(n31874), .Z(n26087) );
  NAND U26805 ( .A(n26088), .B(n26087), .Z(n26413) );
  NAND U26806 ( .A(n34848), .B(n26089), .Z(n26091) );
  XOR U26807 ( .A(n35375), .B(n35377), .Z(n26272) );
  NAND U26808 ( .A(n34618), .B(n26272), .Z(n26090) );
  NAND U26809 ( .A(n26091), .B(n26090), .Z(n26410) );
  NAND U26810 ( .A(n35188), .B(n26092), .Z(n26094) );
  XNOR U26811 ( .A(n35540), .B(a[91]), .Z(n26275) );
  NANDN U26812 ( .A(n34968), .B(n26275), .Z(n26093) );
  AND U26813 ( .A(n26094), .B(n26093), .Z(n26411) );
  XNOR U26814 ( .A(n26410), .B(n26411), .Z(n26412) );
  XNOR U26815 ( .A(n26413), .B(n26412), .Z(n26239) );
  NANDN U26816 ( .A(n26096), .B(n26095), .Z(n26100) );
  NAND U26817 ( .A(n26098), .B(n26097), .Z(n26099) );
  NAND U26818 ( .A(n26100), .B(n26099), .Z(n26240) );
  XOR U26819 ( .A(n26239), .B(n26240), .Z(n26242) );
  XNOR U26820 ( .A(n26241), .B(n26242), .Z(n26258) );
  XNOR U26821 ( .A(n26257), .B(n26258), .Z(n26259) );
  XOR U26822 ( .A(n26260), .B(n26259), .Z(n26360) );
  NANDN U26823 ( .A(n26102), .B(n26101), .Z(n26106) );
  NAND U26824 ( .A(n26104), .B(n26103), .Z(n26105) );
  NAND U26825 ( .A(n26106), .B(n26105), .Z(n26449) );
  XOR U26826 ( .A(b[41]), .B(a[79]), .Z(n26332) );
  NANDN U26827 ( .A(n36905), .B(n26332), .Z(n26109) );
  NANDN U26828 ( .A(n26107), .B(n36807), .Z(n26108) );
  NAND U26829 ( .A(n26109), .B(n26108), .Z(n26354) );
  XNOR U26830 ( .A(b[57]), .B(a[63]), .Z(n26335) );
  OR U26831 ( .A(n26335), .B(n965), .Z(n26112) );
  NANDN U26832 ( .A(n26110), .B(n38194), .Z(n26111) );
  NAND U26833 ( .A(n26112), .B(n26111), .Z(n26351) );
  NAND U26834 ( .A(n38326), .B(n26113), .Z(n26115) );
  XOR U26835 ( .A(n38400), .B(n27773), .Z(n26338) );
  NANDN U26836 ( .A(n38273), .B(n26338), .Z(n26114) );
  AND U26837 ( .A(n26115), .B(n26114), .Z(n26352) );
  XNOR U26838 ( .A(n26351), .B(n26352), .Z(n26353) );
  XNOR U26839 ( .A(n26354), .B(n26353), .Z(n26446) );
  XNOR U26840 ( .A(b[33]), .B(a[87]), .Z(n26341) );
  NANDN U26841 ( .A(n26341), .B(n35620), .Z(n26118) );
  NANDN U26842 ( .A(n26116), .B(n35621), .Z(n26117) );
  NAND U26843 ( .A(n26118), .B(n26117), .Z(n26443) );
  NANDN U26844 ( .A(n966), .B(a[119]), .Z(n26119) );
  XOR U26845 ( .A(n29232), .B(n26119), .Z(n26121) );
  IV U26846 ( .A(a[118]), .Z(n38143) );
  NANDN U26847 ( .A(n38143), .B(n966), .Z(n26120) );
  AND U26848 ( .A(n26121), .B(n26120), .Z(n26440) );
  XOR U26849 ( .A(b[63]), .B(n26122), .Z(n26348) );
  NANDN U26850 ( .A(n26348), .B(n38422), .Z(n26125) );
  NANDN U26851 ( .A(n26123), .B(n38423), .Z(n26124) );
  AND U26852 ( .A(n26125), .B(n26124), .Z(n26441) );
  XNOR U26853 ( .A(n26440), .B(n26441), .Z(n26442) );
  XOR U26854 ( .A(n26443), .B(n26442), .Z(n26447) );
  XNOR U26855 ( .A(n26446), .B(n26447), .Z(n26448) );
  XOR U26856 ( .A(n26449), .B(n26448), .Z(n26254) );
  NANDN U26857 ( .A(n26127), .B(n26126), .Z(n26131) );
  NAND U26858 ( .A(n26129), .B(n26128), .Z(n26130) );
  NAND U26859 ( .A(n26131), .B(n26130), .Z(n26251) );
  NANDN U26860 ( .A(n26133), .B(n26132), .Z(n26137) );
  NAND U26861 ( .A(n26135), .B(n26134), .Z(n26136) );
  AND U26862 ( .A(n26137), .B(n26136), .Z(n26252) );
  XNOR U26863 ( .A(n26251), .B(n26252), .Z(n26253) );
  XNOR U26864 ( .A(n26254), .B(n26253), .Z(n26357) );
  NANDN U26865 ( .A(n26139), .B(n26138), .Z(n26143) );
  NANDN U26866 ( .A(n26141), .B(n26140), .Z(n26142) );
  AND U26867 ( .A(n26143), .B(n26142), .Z(n26358) );
  XNOR U26868 ( .A(n26357), .B(n26358), .Z(n26359) );
  XNOR U26869 ( .A(n26360), .B(n26359), .Z(n26461) );
  XOR U26870 ( .A(n26460), .B(n26461), .Z(n26208) );
  XOR U26871 ( .A(n26207), .B(n26208), .Z(n26209) );
  XNOR U26872 ( .A(n26210), .B(n26209), .Z(n26467) );
  NANDN U26873 ( .A(n26145), .B(n26144), .Z(n26149) );
  NANDN U26874 ( .A(n26147), .B(n26146), .Z(n26148) );
  NAND U26875 ( .A(n26149), .B(n26148), .Z(n26464) );
  NAND U26876 ( .A(n26151), .B(n26150), .Z(n26155) );
  NANDN U26877 ( .A(n26153), .B(n26152), .Z(n26154) );
  NAND U26878 ( .A(n26155), .B(n26154), .Z(n26214) );
  NANDN U26879 ( .A(n26157), .B(n26156), .Z(n26161) );
  NAND U26880 ( .A(n26159), .B(n26158), .Z(n26160) );
  NAND U26881 ( .A(n26161), .B(n26160), .Z(n26212) );
  OR U26882 ( .A(n26163), .B(n26162), .Z(n26167) );
  NANDN U26883 ( .A(n26165), .B(n26164), .Z(n26166) );
  AND U26884 ( .A(n26167), .B(n26166), .Z(n26211) );
  XNOR U26885 ( .A(n26212), .B(n26211), .Z(n26213) );
  XOR U26886 ( .A(n26214), .B(n26213), .Z(n26465) );
  XNOR U26887 ( .A(n26464), .B(n26465), .Z(n26466) );
  XOR U26888 ( .A(n26467), .B(n26466), .Z(n26473) );
  NANDN U26889 ( .A(n26169), .B(n26168), .Z(n26173) );
  NAND U26890 ( .A(n26171), .B(n26170), .Z(n26172) );
  NAND U26891 ( .A(n26173), .B(n26172), .Z(n26470) );
  NAND U26892 ( .A(n26175), .B(n26174), .Z(n26179) );
  NANDN U26893 ( .A(n26177), .B(n26176), .Z(n26178) );
  AND U26894 ( .A(n26179), .B(n26178), .Z(n26471) );
  XNOR U26895 ( .A(n26470), .B(n26471), .Z(n26472) );
  XNOR U26896 ( .A(n26473), .B(n26472), .Z(n26476) );
  NANDN U26897 ( .A(n26181), .B(n26180), .Z(n26185) );
  NAND U26898 ( .A(n26183), .B(n26182), .Z(n26184) );
  NAND U26899 ( .A(n26185), .B(n26184), .Z(n26477) );
  XOR U26900 ( .A(n26476), .B(n26477), .Z(n26478) );
  NANDN U26901 ( .A(n26187), .B(n26186), .Z(n26191) );
  NAND U26902 ( .A(n26189), .B(n26188), .Z(n26190) );
  NAND U26903 ( .A(n26191), .B(n26190), .Z(n26479) );
  XOR U26904 ( .A(n26478), .B(n26479), .Z(n26201) );
  XNOR U26905 ( .A(n26201), .B(n26202), .Z(n26203) );
  XNOR U26906 ( .A(n26204), .B(n26203), .Z(n26482) );
  XNOR U26907 ( .A(n26482), .B(sreg[183]), .Z(n26484) );
  NAND U26908 ( .A(n26196), .B(sreg[182]), .Z(n26200) );
  OR U26909 ( .A(n26198), .B(n26197), .Z(n26199) );
  AND U26910 ( .A(n26200), .B(n26199), .Z(n26483) );
  XOR U26911 ( .A(n26484), .B(n26483), .Z(c[183]) );
  NANDN U26912 ( .A(n26202), .B(n26201), .Z(n26206) );
  NAND U26913 ( .A(n26204), .B(n26203), .Z(n26205) );
  NAND U26914 ( .A(n26206), .B(n26205), .Z(n26490) );
  NANDN U26915 ( .A(n26212), .B(n26211), .Z(n26216) );
  NANDN U26916 ( .A(n26214), .B(n26213), .Z(n26215) );
  NAND U26917 ( .A(n26216), .B(n26215), .Z(n26500) );
  XNOR U26918 ( .A(n26499), .B(n26500), .Z(n26501) );
  OR U26919 ( .A(n26218), .B(n26217), .Z(n26222) );
  OR U26920 ( .A(n26220), .B(n26219), .Z(n26221) );
  AND U26921 ( .A(n26222), .B(n26221), .Z(n26505) );
  NAND U26922 ( .A(n26224), .B(n26223), .Z(n26228) );
  NAND U26923 ( .A(n26226), .B(n26225), .Z(n26227) );
  NAND U26924 ( .A(n26228), .B(n26227), .Z(n26766) );
  NANDN U26925 ( .A(n26230), .B(n26229), .Z(n26234) );
  OR U26926 ( .A(n26232), .B(n26231), .Z(n26233) );
  NAND U26927 ( .A(n26234), .B(n26233), .Z(n26764) );
  XNOR U26928 ( .A(n26764), .B(n26763), .Z(n26765) );
  XNOR U26929 ( .A(n26766), .B(n26765), .Z(n26506) );
  XOR U26930 ( .A(n26505), .B(n26506), .Z(n26507) );
  NANDN U26931 ( .A(n26240), .B(n26239), .Z(n26244) );
  NANDN U26932 ( .A(n26242), .B(n26241), .Z(n26243) );
  NAND U26933 ( .A(n26244), .B(n26243), .Z(n26750) );
  NANDN U26934 ( .A(n26246), .B(n26245), .Z(n26250) );
  NAND U26935 ( .A(n26248), .B(n26247), .Z(n26249) );
  AND U26936 ( .A(n26250), .B(n26249), .Z(n26747) );
  NANDN U26937 ( .A(n26252), .B(n26251), .Z(n26256) );
  NAND U26938 ( .A(n26254), .B(n26253), .Z(n26255) );
  NAND U26939 ( .A(n26256), .B(n26255), .Z(n26748) );
  XNOR U26940 ( .A(n26750), .B(n26749), .Z(n26730) );
  NANDN U26941 ( .A(n26258), .B(n26257), .Z(n26262) );
  NANDN U26942 ( .A(n26260), .B(n26259), .Z(n26261) );
  AND U26943 ( .A(n26262), .B(n26261), .Z(n26729) );
  XNOR U26944 ( .A(n26730), .B(n26729), .Z(n26731) );
  NANDN U26945 ( .A(n26264), .B(n26263), .Z(n26268) );
  NAND U26946 ( .A(n26266), .B(n26265), .Z(n26267) );
  NAND U26947 ( .A(n26268), .B(n26267), .Z(n26726) );
  XOR U26948 ( .A(a[108]), .B(n971), .Z(n26660) );
  OR U26949 ( .A(n26660), .B(n31550), .Z(n26271) );
  NANDN U26950 ( .A(n26269), .B(n31874), .Z(n26270) );
  NAND U26951 ( .A(n26271), .B(n26270), .Z(n26538) );
  NAND U26952 ( .A(n34848), .B(n26272), .Z(n26274) );
  XOR U26953 ( .A(n35191), .B(n35375), .Z(n26663) );
  NAND U26954 ( .A(n34618), .B(n26663), .Z(n26273) );
  NAND U26955 ( .A(n26274), .B(n26273), .Z(n26535) );
  NAND U26956 ( .A(n35188), .B(n26275), .Z(n26277) );
  XOR U26957 ( .A(n35540), .B(n34852), .Z(n26666) );
  NANDN U26958 ( .A(n34968), .B(n26666), .Z(n26276) );
  AND U26959 ( .A(n26277), .B(n26276), .Z(n26536) );
  XNOR U26960 ( .A(n26535), .B(n26536), .Z(n26537) );
  XOR U26961 ( .A(n26538), .B(n26537), .Z(n26624) );
  XOR U26962 ( .A(b[37]), .B(n33185), .Z(n26651) );
  NANDN U26963 ( .A(n26651), .B(n36311), .Z(n26280) );
  NANDN U26964 ( .A(n26278), .B(n36309), .Z(n26279) );
  NAND U26965 ( .A(n26280), .B(n26279), .Z(n26714) );
  XOR U26966 ( .A(a[116]), .B(n968), .Z(n26654) );
  OR U26967 ( .A(n26654), .B(n29363), .Z(n26283) );
  NANDN U26968 ( .A(n26281), .B(n29864), .Z(n26282) );
  NAND U26969 ( .A(n26283), .B(n26282), .Z(n26711) );
  XOR U26970 ( .A(n38143), .B(n967), .Z(n26657) );
  NAND U26971 ( .A(n26657), .B(n28939), .Z(n26286) );
  NAND U26972 ( .A(n28938), .B(n26284), .Z(n26285) );
  AND U26973 ( .A(n26286), .B(n26285), .Z(n26712) );
  XNOR U26974 ( .A(n26711), .B(n26712), .Z(n26713) );
  XOR U26975 ( .A(n26714), .B(n26713), .Z(n26625) );
  XNOR U26976 ( .A(n26624), .B(n26625), .Z(n26627) );
  NANDN U26977 ( .A(n26288), .B(n26287), .Z(n26292) );
  NAND U26978 ( .A(n26290), .B(n26289), .Z(n26291) );
  NAND U26979 ( .A(n26292), .B(n26291), .Z(n26626) );
  XNOR U26980 ( .A(n26627), .B(n26626), .Z(n26724) );
  NANDN U26981 ( .A(n26294), .B(n26293), .Z(n26298) );
  NAND U26982 ( .A(n26296), .B(n26295), .Z(n26297) );
  NAND U26983 ( .A(n26298), .B(n26297), .Z(n26589) );
  NAND U26984 ( .A(a[56]), .B(b[63]), .Z(n26603) );
  NANDN U26985 ( .A(n26299), .B(n38369), .Z(n26301) );
  XOR U26986 ( .A(b[61]), .B(n27436), .Z(n26645) );
  OR U26987 ( .A(n26645), .B(n38371), .Z(n26300) );
  NAND U26988 ( .A(n26301), .B(n26300), .Z(n26601) );
  NANDN U26989 ( .A(n26302), .B(n35311), .Z(n26304) );
  XOR U26990 ( .A(b[31]), .B(n34851), .Z(n26648) );
  NANDN U26991 ( .A(n26648), .B(n35313), .Z(n26303) );
  AND U26992 ( .A(n26304), .B(n26303), .Z(n26600) );
  XNOR U26993 ( .A(n26601), .B(n26600), .Z(n26602) );
  XOR U26994 ( .A(n26603), .B(n26602), .Z(n26587) );
  NAND U26995 ( .A(n33283), .B(n26305), .Z(n26307) );
  XOR U26996 ( .A(n36420), .B(n33020), .Z(n26630) );
  NANDN U26997 ( .A(n33021), .B(n26630), .Z(n26306) );
  NAND U26998 ( .A(n26307), .B(n26306), .Z(n26702) );
  XNOR U26999 ( .A(a[100]), .B(b[21]), .Z(n26633) );
  OR U27000 ( .A(n26633), .B(n33634), .Z(n26310) );
  NAND U27001 ( .A(n26308), .B(n33464), .Z(n26309) );
  NAND U27002 ( .A(n26310), .B(n26309), .Z(n26699) );
  NAND U27003 ( .A(n34044), .B(n26311), .Z(n26313) );
  XOR U27004 ( .A(n35783), .B(n34510), .Z(n26636) );
  NANDN U27005 ( .A(n33867), .B(n26636), .Z(n26312) );
  AND U27006 ( .A(n26313), .B(n26312), .Z(n26700) );
  XNOR U27007 ( .A(n26699), .B(n26700), .Z(n26701) );
  XNOR U27008 ( .A(n26702), .B(n26701), .Z(n26588) );
  XNOR U27009 ( .A(n26587), .B(n26588), .Z(n26590) );
  XNOR U27010 ( .A(n26589), .B(n26590), .Z(n26723) );
  XOR U27011 ( .A(n26724), .B(n26723), .Z(n26725) );
  XOR U27012 ( .A(n26726), .B(n26725), .Z(n26513) );
  NANDN U27013 ( .A(n26315), .B(n26314), .Z(n26319) );
  OR U27014 ( .A(n26317), .B(n26316), .Z(n26318) );
  NAND U27015 ( .A(n26319), .B(n26318), .Z(n26512) );
  NANDN U27016 ( .A(n26321), .B(n26320), .Z(n26325) );
  NAND U27017 ( .A(n26323), .B(n26322), .Z(n26324) );
  NAND U27018 ( .A(n26325), .B(n26324), .Z(n26621) );
  NANDN U27019 ( .A(n26327), .B(n26326), .Z(n26331) );
  NAND U27020 ( .A(n26329), .B(n26328), .Z(n26330) );
  NAND U27021 ( .A(n26331), .B(n26330), .Z(n26554) );
  XNOR U27022 ( .A(b[41]), .B(a[80]), .Z(n26681) );
  OR U27023 ( .A(n26681), .B(n36905), .Z(n26334) );
  NAND U27024 ( .A(n26332), .B(n36807), .Z(n26333) );
  NAND U27025 ( .A(n26334), .B(n26333), .Z(n26708) );
  XNOR U27026 ( .A(b[57]), .B(a[64]), .Z(n26684) );
  OR U27027 ( .A(n26684), .B(n965), .Z(n26337) );
  NANDN U27028 ( .A(n26335), .B(n38194), .Z(n26336) );
  NAND U27029 ( .A(n26337), .B(n26336), .Z(n26705) );
  NAND U27030 ( .A(n38326), .B(n26338), .Z(n26340) );
  XNOR U27031 ( .A(n38400), .B(a[62]), .Z(n26687) );
  NANDN U27032 ( .A(n38273), .B(n26687), .Z(n26339) );
  AND U27033 ( .A(n26340), .B(n26339), .Z(n26706) );
  XNOR U27034 ( .A(n26705), .B(n26706), .Z(n26707) );
  XOR U27035 ( .A(n26708), .B(n26707), .Z(n26552) );
  XOR U27036 ( .A(b[33]), .B(n34048), .Z(n26690) );
  NANDN U27037 ( .A(n26690), .B(n35620), .Z(n26343) );
  NANDN U27038 ( .A(n26341), .B(n35621), .Z(n26342) );
  NAND U27039 ( .A(n26343), .B(n26342), .Z(n26550) );
  NANDN U27040 ( .A(n966), .B(a[120]), .Z(n26344) );
  XOR U27041 ( .A(n29232), .B(n26344), .Z(n26346) );
  IV U27042 ( .A(a[119]), .Z(n38193) );
  NANDN U27043 ( .A(n38193), .B(n966), .Z(n26345) );
  AND U27044 ( .A(n26346), .B(n26345), .Z(n26547) );
  XOR U27045 ( .A(b[63]), .B(n26347), .Z(n26696) );
  NANDN U27046 ( .A(n26696), .B(n38422), .Z(n26350) );
  NANDN U27047 ( .A(n26348), .B(n38423), .Z(n26349) );
  AND U27048 ( .A(n26350), .B(n26349), .Z(n26548) );
  XNOR U27049 ( .A(n26547), .B(n26548), .Z(n26549) );
  XNOR U27050 ( .A(n26550), .B(n26549), .Z(n26551) );
  XOR U27051 ( .A(n26552), .B(n26551), .Z(n26553) );
  XNOR U27052 ( .A(n26554), .B(n26553), .Z(n26619) );
  NANDN U27053 ( .A(n26352), .B(n26351), .Z(n26356) );
  NAND U27054 ( .A(n26354), .B(n26353), .Z(n26355) );
  AND U27055 ( .A(n26356), .B(n26355), .Z(n26618) );
  XNOR U27056 ( .A(n26619), .B(n26618), .Z(n26620) );
  XNOR U27057 ( .A(n26621), .B(n26620), .Z(n26511) );
  XNOR U27058 ( .A(n26512), .B(n26511), .Z(n26514) );
  XNOR U27059 ( .A(n26513), .B(n26514), .Z(n26732) );
  XNOR U27060 ( .A(n26731), .B(n26732), .Z(n26759) );
  NANDN U27061 ( .A(n26362), .B(n26361), .Z(n26366) );
  NANDN U27062 ( .A(n26364), .B(n26363), .Z(n26365) );
  NAND U27063 ( .A(n26366), .B(n26365), .Z(n26735) );
  XOR U27064 ( .A(a[110]), .B(n970), .Z(n26563) );
  OR U27065 ( .A(n26563), .B(n31369), .Z(n26369) );
  NANDN U27066 ( .A(n26367), .B(n31119), .Z(n26368) );
  NAND U27067 ( .A(n26369), .B(n26368), .Z(n26584) );
  XOR U27068 ( .A(b[43]), .B(n31870), .Z(n26566) );
  NANDN U27069 ( .A(n26566), .B(n37068), .Z(n26372) );
  NANDN U27070 ( .A(n26370), .B(n37069), .Z(n26371) );
  NAND U27071 ( .A(n26372), .B(n26371), .Z(n26581) );
  XNOR U27072 ( .A(b[45]), .B(a[76]), .Z(n26569) );
  NANDN U27073 ( .A(n26569), .B(n37261), .Z(n26375) );
  NAND U27074 ( .A(n26373), .B(n37262), .Z(n26374) );
  AND U27075 ( .A(n26375), .B(n26374), .Z(n26582) );
  XNOR U27076 ( .A(n26581), .B(n26582), .Z(n26583) );
  XNOR U27077 ( .A(n26584), .B(n26583), .Z(n26675) );
  XOR U27078 ( .A(b[49]), .B(n30210), .Z(n26572) );
  OR U27079 ( .A(n26572), .B(n37756), .Z(n26378) );
  NANDN U27080 ( .A(n26376), .B(n37652), .Z(n26377) );
  NAND U27081 ( .A(n26378), .B(n26377), .Z(n26609) );
  NAND U27082 ( .A(n26379), .B(n37469), .Z(n26381) );
  XOR U27083 ( .A(n978), .B(n31372), .Z(n26575) );
  NAND U27084 ( .A(n26575), .B(n37471), .Z(n26380) );
  AND U27085 ( .A(n26381), .B(n26380), .Z(n26606) );
  XOR U27086 ( .A(a[112]), .B(n969), .Z(n26578) );
  NANDN U27087 ( .A(n26578), .B(n30509), .Z(n26384) );
  NAND U27088 ( .A(n26382), .B(n30846), .Z(n26383) );
  AND U27089 ( .A(n26384), .B(n26383), .Z(n26607) );
  XOR U27090 ( .A(n26609), .B(n26608), .Z(n26676) );
  XNOR U27091 ( .A(n26675), .B(n26676), .Z(n26677) );
  NANDN U27092 ( .A(n26386), .B(n26385), .Z(n26390) );
  NAND U27093 ( .A(n26388), .B(n26387), .Z(n26389) );
  AND U27094 ( .A(n26390), .B(n26389), .Z(n26678) );
  XNOR U27095 ( .A(n26677), .B(n26678), .Z(n26736) );
  XNOR U27096 ( .A(n26735), .B(n26736), .Z(n26737) );
  XNOR U27097 ( .A(b[35]), .B(a[86]), .Z(n26591) );
  NANDN U27098 ( .A(n26591), .B(n35985), .Z(n26393) );
  NAND U27099 ( .A(n26391), .B(n35986), .Z(n26392) );
  NAND U27100 ( .A(n26393), .B(n26392), .Z(n26544) );
  XOR U27101 ( .A(n37873), .B(n31123), .Z(n26594) );
  NAND U27102 ( .A(n26594), .B(n29949), .Z(n26396) );
  NAND U27103 ( .A(n29948), .B(n26394), .Z(n26395) );
  NAND U27104 ( .A(n26396), .B(n26395), .Z(n26541) );
  XOR U27105 ( .A(b[55]), .B(n28701), .Z(n26597) );
  NANDN U27106 ( .A(n26597), .B(n38075), .Z(n26399) );
  NANDN U27107 ( .A(n26397), .B(n38073), .Z(n26398) );
  AND U27108 ( .A(n26399), .B(n26398), .Z(n26542) );
  XNOR U27109 ( .A(n26541), .B(n26542), .Z(n26543) );
  XNOR U27110 ( .A(n26544), .B(n26543), .Z(n26615) );
  NANDN U27111 ( .A(n26401), .B(n26400), .Z(n26405) );
  NAND U27112 ( .A(n26403), .B(n26402), .Z(n26404) );
  NAND U27113 ( .A(n26405), .B(n26404), .Z(n26612) );
  XNOR U27114 ( .A(n26612), .B(n26613), .Z(n26614) );
  XOR U27115 ( .A(n26615), .B(n26614), .Z(n26738) );
  XNOR U27116 ( .A(n26737), .B(n26738), .Z(n26754) );
  NANDN U27117 ( .A(n26411), .B(n26410), .Z(n26415) );
  NAND U27118 ( .A(n26413), .B(n26412), .Z(n26414) );
  NAND U27119 ( .A(n26415), .B(n26414), .Z(n26720) );
  XOR U27120 ( .A(a[106]), .B(n972), .Z(n26517) );
  OR U27121 ( .A(n26517), .B(n32010), .Z(n26418) );
  NANDN U27122 ( .A(n26416), .B(n32011), .Z(n26417) );
  NAND U27123 ( .A(n26418), .B(n26417), .Z(n26642) );
  XNOR U27124 ( .A(n35545), .B(b[25]), .Z(n26520) );
  NANDN U27125 ( .A(n34219), .B(n26520), .Z(n26421) );
  NAND U27126 ( .A(n34217), .B(n26419), .Z(n26420) );
  NAND U27127 ( .A(n26421), .B(n26420), .Z(n26639) );
  XNOR U27128 ( .A(a[104]), .B(b[17]), .Z(n26523) );
  NANDN U27129 ( .A(n26523), .B(n32543), .Z(n26424) );
  NAND U27130 ( .A(n26422), .B(n32541), .Z(n26423) );
  AND U27131 ( .A(n26424), .B(n26423), .Z(n26640) );
  XNOR U27132 ( .A(n26639), .B(n26640), .Z(n26641) );
  XNOR U27133 ( .A(n26642), .B(n26641), .Z(n26717) );
  XOR U27134 ( .A(b[39]), .B(n32815), .Z(n26526) );
  NANDN U27135 ( .A(n26526), .B(n36553), .Z(n26427) );
  NANDN U27136 ( .A(n26425), .B(n36643), .Z(n26426) );
  NAND U27137 ( .A(n26427), .B(n26426), .Z(n26672) );
  XOR U27138 ( .A(b[51]), .B(n30379), .Z(n26529) );
  NANDN U27139 ( .A(n26529), .B(n37803), .Z(n26430) );
  NANDN U27140 ( .A(n26428), .B(n37802), .Z(n26429) );
  NAND U27141 ( .A(n26430), .B(n26429), .Z(n26669) );
  XOR U27142 ( .A(b[53]), .B(n29868), .Z(n26532) );
  NANDN U27143 ( .A(n26532), .B(n37940), .Z(n26433) );
  NANDN U27144 ( .A(n26431), .B(n37941), .Z(n26432) );
  AND U27145 ( .A(n26433), .B(n26432), .Z(n26670) );
  XNOR U27146 ( .A(n26669), .B(n26670), .Z(n26671) );
  XOR U27147 ( .A(n26672), .B(n26671), .Z(n26718) );
  XNOR U27148 ( .A(n26717), .B(n26718), .Z(n26719) );
  XOR U27149 ( .A(n26720), .B(n26719), .Z(n26560) );
  NANDN U27150 ( .A(n26435), .B(n26434), .Z(n26439) );
  NAND U27151 ( .A(n26437), .B(n26436), .Z(n26438) );
  NAND U27152 ( .A(n26439), .B(n26438), .Z(n26557) );
  NANDN U27153 ( .A(n26441), .B(n26440), .Z(n26445) );
  NAND U27154 ( .A(n26443), .B(n26442), .Z(n26444) );
  AND U27155 ( .A(n26445), .B(n26444), .Z(n26558) );
  XNOR U27156 ( .A(n26557), .B(n26558), .Z(n26559) );
  XNOR U27157 ( .A(n26560), .B(n26559), .Z(n26741) );
  NANDN U27158 ( .A(n26447), .B(n26446), .Z(n26451) );
  NANDN U27159 ( .A(n26449), .B(n26448), .Z(n26450) );
  AND U27160 ( .A(n26451), .B(n26450), .Z(n26742) );
  XOR U27161 ( .A(n26741), .B(n26742), .Z(n26744) );
  NANDN U27162 ( .A(n26453), .B(n26452), .Z(n26457) );
  NAND U27163 ( .A(n26455), .B(n26454), .Z(n26456) );
  AND U27164 ( .A(n26457), .B(n26456), .Z(n26743) );
  XNOR U27165 ( .A(n26744), .B(n26743), .Z(n26753) );
  XOR U27166 ( .A(n26756), .B(n26755), .Z(n26760) );
  XNOR U27167 ( .A(n26759), .B(n26760), .Z(n26761) );
  NAND U27168 ( .A(n26459), .B(n26458), .Z(n26463) );
  OR U27169 ( .A(n26461), .B(n26460), .Z(n26462) );
  AND U27170 ( .A(n26463), .B(n26462), .Z(n26762) );
  XOR U27171 ( .A(n26761), .B(n26762), .Z(n26508) );
  XOR U27172 ( .A(n26507), .B(n26508), .Z(n26502) );
  XOR U27173 ( .A(n26501), .B(n26502), .Z(n26493) );
  NANDN U27174 ( .A(n26465), .B(n26464), .Z(n26469) );
  NAND U27175 ( .A(n26467), .B(n26466), .Z(n26468) );
  AND U27176 ( .A(n26469), .B(n26468), .Z(n26494) );
  XNOR U27177 ( .A(n26493), .B(n26494), .Z(n26495) );
  NANDN U27178 ( .A(n26471), .B(n26470), .Z(n26475) );
  NANDN U27179 ( .A(n26473), .B(n26472), .Z(n26474) );
  NAND U27180 ( .A(n26475), .B(n26474), .Z(n26496) );
  XOR U27181 ( .A(n26495), .B(n26496), .Z(n26487) );
  OR U27182 ( .A(n26477), .B(n26476), .Z(n26481) );
  NANDN U27183 ( .A(n26479), .B(n26478), .Z(n26480) );
  NAND U27184 ( .A(n26481), .B(n26480), .Z(n26488) );
  XNOR U27185 ( .A(n26487), .B(n26488), .Z(n26489) );
  XNOR U27186 ( .A(n26490), .B(n26489), .Z(n26769) );
  XNOR U27187 ( .A(n26769), .B(sreg[184]), .Z(n26771) );
  NAND U27188 ( .A(n26482), .B(sreg[183]), .Z(n26486) );
  OR U27189 ( .A(n26484), .B(n26483), .Z(n26485) );
  AND U27190 ( .A(n26486), .B(n26485), .Z(n26770) );
  XOR U27191 ( .A(n26771), .B(n26770), .Z(c[184]) );
  NANDN U27192 ( .A(n26488), .B(n26487), .Z(n26492) );
  NAND U27193 ( .A(n26490), .B(n26489), .Z(n26491) );
  NAND U27194 ( .A(n26492), .B(n26491), .Z(n26777) );
  NANDN U27195 ( .A(n26494), .B(n26493), .Z(n26498) );
  NANDN U27196 ( .A(n26496), .B(n26495), .Z(n26497) );
  NAND U27197 ( .A(n26498), .B(n26497), .Z(n26775) );
  NANDN U27198 ( .A(n26500), .B(n26499), .Z(n26504) );
  NANDN U27199 ( .A(n26502), .B(n26501), .Z(n26503) );
  NAND U27200 ( .A(n26504), .B(n26503), .Z(n26778) );
  OR U27201 ( .A(n26506), .B(n26505), .Z(n26510) );
  NANDN U27202 ( .A(n26508), .B(n26507), .Z(n26509) );
  AND U27203 ( .A(n26510), .B(n26509), .Z(n26779) );
  XNOR U27204 ( .A(n26778), .B(n26779), .Z(n26780) );
  NAND U27205 ( .A(n26512), .B(n26511), .Z(n26516) );
  NANDN U27206 ( .A(n26514), .B(n26513), .Z(n26515) );
  NAND U27207 ( .A(n26516), .B(n26515), .Z(n27023) );
  XNOR U27208 ( .A(a[107]), .B(b[15]), .Z(n26875) );
  OR U27209 ( .A(n26875), .B(n32010), .Z(n26519) );
  NANDN U27210 ( .A(n26517), .B(n32011), .Z(n26518) );
  NAND U27211 ( .A(n26519), .B(n26518), .Z(n26939) );
  XOR U27212 ( .A(a[97]), .B(b[25]), .Z(n26878) );
  NANDN U27213 ( .A(n34219), .B(n26878), .Z(n26522) );
  NAND U27214 ( .A(n34217), .B(n26520), .Z(n26521) );
  NAND U27215 ( .A(n26522), .B(n26521), .Z(n26936) );
  XOR U27216 ( .A(a[105]), .B(b[17]), .Z(n26881) );
  NAND U27217 ( .A(n26881), .B(n32543), .Z(n26525) );
  NANDN U27218 ( .A(n26523), .B(n32541), .Z(n26524) );
  AND U27219 ( .A(n26525), .B(n26524), .Z(n26937) );
  XNOR U27220 ( .A(n26936), .B(n26937), .Z(n26938) );
  XNOR U27221 ( .A(n26939), .B(n26938), .Z(n26972) );
  XNOR U27222 ( .A(b[39]), .B(a[83]), .Z(n26884) );
  NANDN U27223 ( .A(n26884), .B(n36553), .Z(n26528) );
  NANDN U27224 ( .A(n26526), .B(n36643), .Z(n26527) );
  NAND U27225 ( .A(n26528), .B(n26527), .Z(n26969) );
  XOR U27226 ( .A(b[51]), .B(n30543), .Z(n26887) );
  NANDN U27227 ( .A(n26887), .B(n37803), .Z(n26531) );
  NANDN U27228 ( .A(n26529), .B(n37802), .Z(n26530) );
  NAND U27229 ( .A(n26531), .B(n26530), .Z(n26966) );
  XNOR U27230 ( .A(b[53]), .B(a[69]), .Z(n26890) );
  NANDN U27231 ( .A(n26890), .B(n37940), .Z(n26534) );
  NANDN U27232 ( .A(n26532), .B(n37941), .Z(n26533) );
  AND U27233 ( .A(n26534), .B(n26533), .Z(n26967) );
  XNOR U27234 ( .A(n26966), .B(n26967), .Z(n26968) );
  XOR U27235 ( .A(n26969), .B(n26968), .Z(n26973) );
  XOR U27236 ( .A(n26972), .B(n26973), .Z(n26975) );
  NANDN U27237 ( .A(n26536), .B(n26535), .Z(n26540) );
  NAND U27238 ( .A(n26538), .B(n26537), .Z(n26539) );
  NAND U27239 ( .A(n26540), .B(n26539), .Z(n26974) );
  XNOR U27240 ( .A(n26975), .B(n26974), .Z(n26866) );
  NANDN U27241 ( .A(n26542), .B(n26541), .Z(n26546) );
  NAND U27242 ( .A(n26544), .B(n26543), .Z(n26545) );
  NAND U27243 ( .A(n26546), .B(n26545), .Z(n26863) );
  XNOR U27244 ( .A(n26863), .B(n26864), .Z(n26865) );
  XNOR U27245 ( .A(n26866), .B(n26865), .Z(n27036) );
  NANDN U27246 ( .A(n26552), .B(n26551), .Z(n26556) );
  OR U27247 ( .A(n26554), .B(n26553), .Z(n26555) );
  AND U27248 ( .A(n26556), .B(n26555), .Z(n27037) );
  XNOR U27249 ( .A(n27036), .B(n27037), .Z(n27038) );
  NANDN U27250 ( .A(n26558), .B(n26557), .Z(n26562) );
  NAND U27251 ( .A(n26560), .B(n26559), .Z(n26561) );
  AND U27252 ( .A(n26562), .B(n26561), .Z(n27039) );
  XNOR U27253 ( .A(n27038), .B(n27039), .Z(n27020) );
  XNOR U27254 ( .A(a[111]), .B(b[11]), .Z(n26812) );
  OR U27255 ( .A(n26812), .B(n31369), .Z(n26565) );
  NANDN U27256 ( .A(n26563), .B(n31119), .Z(n26564) );
  NAND U27257 ( .A(n26565), .B(n26564), .Z(n26833) );
  XNOR U27258 ( .A(b[43]), .B(a[79]), .Z(n26815) );
  NANDN U27259 ( .A(n26815), .B(n37068), .Z(n26568) );
  NANDN U27260 ( .A(n26566), .B(n37069), .Z(n26567) );
  NAND U27261 ( .A(n26568), .B(n26567), .Z(n26830) );
  XOR U27262 ( .A(b[45]), .B(a[77]), .Z(n26818) );
  NAND U27263 ( .A(n26818), .B(n37261), .Z(n26571) );
  NANDN U27264 ( .A(n26569), .B(n37262), .Z(n26570) );
  AND U27265 ( .A(n26571), .B(n26570), .Z(n26831) );
  XNOR U27266 ( .A(n26830), .B(n26831), .Z(n26832) );
  XNOR U27267 ( .A(n26833), .B(n26832), .Z(n26926) );
  XNOR U27268 ( .A(b[49]), .B(a[73]), .Z(n26821) );
  OR U27269 ( .A(n26821), .B(n37756), .Z(n26574) );
  NANDN U27270 ( .A(n26572), .B(n37652), .Z(n26573) );
  NAND U27271 ( .A(n26574), .B(n26573), .Z(n26854) );
  NAND U27272 ( .A(n37469), .B(n26575), .Z(n26577) );
  XNOR U27273 ( .A(n978), .B(a[75]), .Z(n26824) );
  NAND U27274 ( .A(n26824), .B(n37471), .Z(n26576) );
  NAND U27275 ( .A(n26577), .B(n26576), .Z(n26851) );
  XNOR U27276 ( .A(a[113]), .B(b[9]), .Z(n26827) );
  NANDN U27277 ( .A(n26827), .B(n30509), .Z(n26580) );
  NANDN U27278 ( .A(n26578), .B(n30846), .Z(n26579) );
  AND U27279 ( .A(n26580), .B(n26579), .Z(n26852) );
  XNOR U27280 ( .A(n26851), .B(n26852), .Z(n26853) );
  XNOR U27281 ( .A(n26854), .B(n26853), .Z(n26923) );
  NANDN U27282 ( .A(n26582), .B(n26581), .Z(n26586) );
  NAND U27283 ( .A(n26584), .B(n26583), .Z(n26585) );
  NAND U27284 ( .A(n26586), .B(n26585), .Z(n26924) );
  XNOR U27285 ( .A(n26923), .B(n26924), .Z(n26925) );
  XOR U27286 ( .A(n26926), .B(n26925), .Z(n27026) );
  XNOR U27287 ( .A(n27026), .B(n27027), .Z(n27029) );
  XOR U27288 ( .A(b[35]), .B(a[87]), .Z(n26836) );
  NAND U27289 ( .A(n35985), .B(n26836), .Z(n26593) );
  NANDN U27290 ( .A(n26591), .B(n35986), .Z(n26592) );
  NAND U27291 ( .A(n26593), .B(n26592), .Z(n26902) );
  XNOR U27292 ( .A(a[115]), .B(n31123), .Z(n26839) );
  NAND U27293 ( .A(n26839), .B(n29949), .Z(n26596) );
  NAND U27294 ( .A(n29948), .B(n26594), .Z(n26595) );
  NAND U27295 ( .A(n26596), .B(n26595), .Z(n26899) );
  XOR U27296 ( .A(b[55]), .B(n29372), .Z(n26842) );
  NANDN U27297 ( .A(n26842), .B(n38075), .Z(n26599) );
  NANDN U27298 ( .A(n26597), .B(n38073), .Z(n26598) );
  AND U27299 ( .A(n26599), .B(n26598), .Z(n26900) );
  XNOR U27300 ( .A(n26899), .B(n26900), .Z(n26901) );
  XNOR U27301 ( .A(n26902), .B(n26901), .Z(n26914) );
  NANDN U27302 ( .A(n26601), .B(n26600), .Z(n26605) );
  NAND U27303 ( .A(n26603), .B(n26602), .Z(n26604) );
  NAND U27304 ( .A(n26605), .B(n26604), .Z(n26911) );
  OR U27305 ( .A(n26607), .B(n26606), .Z(n26611) );
  NAND U27306 ( .A(n26609), .B(n26608), .Z(n26610) );
  NAND U27307 ( .A(n26611), .B(n26610), .Z(n26912) );
  XNOR U27308 ( .A(n26911), .B(n26912), .Z(n26913) );
  XOR U27309 ( .A(n26914), .B(n26913), .Z(n27028) );
  XOR U27310 ( .A(n27029), .B(n27028), .Z(n27021) );
  XOR U27311 ( .A(n27020), .B(n27021), .Z(n27022) );
  XNOR U27312 ( .A(n27023), .B(n27022), .Z(n26790) );
  NANDN U27313 ( .A(n26613), .B(n26612), .Z(n26617) );
  NAND U27314 ( .A(n26615), .B(n26614), .Z(n26616) );
  NAND U27315 ( .A(n26617), .B(n26616), .Z(n27034) );
  NANDN U27316 ( .A(n26619), .B(n26618), .Z(n26623) );
  NANDN U27317 ( .A(n26621), .B(n26620), .Z(n26622) );
  NAND U27318 ( .A(n26623), .B(n26622), .Z(n27032) );
  OR U27319 ( .A(n26625), .B(n26624), .Z(n26629) );
  OR U27320 ( .A(n26627), .B(n26626), .Z(n26628) );
  NAND U27321 ( .A(n26629), .B(n26628), .Z(n27033) );
  XNOR U27322 ( .A(n27032), .B(n27033), .Z(n27035) );
  XOR U27323 ( .A(n27034), .B(n27035), .Z(n26799) );
  NAND U27324 ( .A(n33283), .B(n26630), .Z(n26632) );
  XNOR U27325 ( .A(a[103]), .B(n33020), .Z(n26927) );
  NANDN U27326 ( .A(n33021), .B(n26927), .Z(n26631) );
  NAND U27327 ( .A(n26632), .B(n26631), .Z(n26987) );
  XOR U27328 ( .A(a[101]), .B(b[21]), .Z(n26930) );
  NANDN U27329 ( .A(n33634), .B(n26930), .Z(n26635) );
  NANDN U27330 ( .A(n26633), .B(n33464), .Z(n26634) );
  NAND U27331 ( .A(n26635), .B(n26634), .Z(n26984) );
  NAND U27332 ( .A(n34044), .B(n26636), .Z(n26638) );
  XNOR U27333 ( .A(a[99]), .B(n34510), .Z(n26933) );
  NANDN U27334 ( .A(n33867), .B(n26933), .Z(n26637) );
  AND U27335 ( .A(n26638), .B(n26637), .Z(n26985) );
  XNOR U27336 ( .A(n26984), .B(n26985), .Z(n26986) );
  XNOR U27337 ( .A(n26987), .B(n26986), .Z(n26806) );
  NANDN U27338 ( .A(n26640), .B(n26639), .Z(n26644) );
  NAND U27339 ( .A(n26642), .B(n26641), .Z(n26643) );
  NAND U27340 ( .A(n26644), .B(n26643), .Z(n26807) );
  XNOR U27341 ( .A(n26806), .B(n26807), .Z(n26808) );
  NAND U27342 ( .A(a[57]), .B(b[63]), .Z(n26848) );
  NANDN U27343 ( .A(n26645), .B(n38369), .Z(n26647) );
  XOR U27344 ( .A(b[61]), .B(n27773), .Z(n26942) );
  OR U27345 ( .A(n26942), .B(n38371), .Z(n26646) );
  NAND U27346 ( .A(n26647), .B(n26646), .Z(n26846) );
  NANDN U27347 ( .A(n26648), .B(n35311), .Z(n26650) );
  XNOR U27348 ( .A(b[31]), .B(a[91]), .Z(n26945) );
  NANDN U27349 ( .A(n26945), .B(n35313), .Z(n26649) );
  AND U27350 ( .A(n26650), .B(n26649), .Z(n26845) );
  XNOR U27351 ( .A(n26846), .B(n26845), .Z(n26847) );
  XNOR U27352 ( .A(n26848), .B(n26847), .Z(n26809) );
  XOR U27353 ( .A(n26808), .B(n26809), .Z(n27014) );
  XNOR U27354 ( .A(b[37]), .B(a[85]), .Z(n26948) );
  NANDN U27355 ( .A(n26948), .B(n36311), .Z(n26653) );
  NANDN U27356 ( .A(n26651), .B(n36309), .Z(n26652) );
  NAND U27357 ( .A(n26653), .B(n26652), .Z(n26981) );
  XNOR U27358 ( .A(a[117]), .B(b[5]), .Z(n26951) );
  OR U27359 ( .A(n26951), .B(n29363), .Z(n26656) );
  NANDN U27360 ( .A(n26654), .B(n29864), .Z(n26655) );
  NAND U27361 ( .A(n26656), .B(n26655), .Z(n26978) );
  XOR U27362 ( .A(n38193), .B(n967), .Z(n26954) );
  NAND U27363 ( .A(n26954), .B(n28939), .Z(n26659) );
  NAND U27364 ( .A(n28938), .B(n26657), .Z(n26658) );
  AND U27365 ( .A(n26659), .B(n26658), .Z(n26979) );
  XNOR U27366 ( .A(n26978), .B(n26979), .Z(n26980) );
  XNOR U27367 ( .A(n26981), .B(n26980), .Z(n26907) );
  XNOR U27368 ( .A(a[109]), .B(b[13]), .Z(n26957) );
  OR U27369 ( .A(n26957), .B(n31550), .Z(n26662) );
  NANDN U27370 ( .A(n26660), .B(n31874), .Z(n26661) );
  NAND U27371 ( .A(n26662), .B(n26661), .Z(n26896) );
  NAND U27372 ( .A(n34848), .B(n26663), .Z(n26665) );
  XOR U27373 ( .A(n35628), .B(n35375), .Z(n26960) );
  NAND U27374 ( .A(n34618), .B(n26960), .Z(n26664) );
  NAND U27375 ( .A(n26665), .B(n26664), .Z(n26893) );
  NAND U27376 ( .A(n35188), .B(n26666), .Z(n26668) );
  XOR U27377 ( .A(n35540), .B(n35377), .Z(n26963) );
  NANDN U27378 ( .A(n34968), .B(n26963), .Z(n26667) );
  AND U27379 ( .A(n26668), .B(n26667), .Z(n26894) );
  XNOR U27380 ( .A(n26893), .B(n26894), .Z(n26895) );
  XNOR U27381 ( .A(n26896), .B(n26895), .Z(n26905) );
  NANDN U27382 ( .A(n26670), .B(n26669), .Z(n26674) );
  NAND U27383 ( .A(n26672), .B(n26671), .Z(n26673) );
  NAND U27384 ( .A(n26674), .B(n26673), .Z(n26906) );
  XOR U27385 ( .A(n26905), .B(n26906), .Z(n26908) );
  XNOR U27386 ( .A(n26907), .B(n26908), .Z(n27015) );
  XNOR U27387 ( .A(n27014), .B(n27015), .Z(n27016) );
  NANDN U27388 ( .A(n26676), .B(n26675), .Z(n26680) );
  NAND U27389 ( .A(n26678), .B(n26677), .Z(n26679) );
  NAND U27390 ( .A(n26680), .B(n26679), .Z(n27017) );
  XOR U27391 ( .A(n27016), .B(n27017), .Z(n26805) );
  XOR U27392 ( .A(b[41]), .B(a[81]), .Z(n26990) );
  NANDN U27393 ( .A(n36905), .B(n26990), .Z(n26683) );
  NANDN U27394 ( .A(n26681), .B(n36807), .Z(n26682) );
  NAND U27395 ( .A(n26683), .B(n26682), .Z(n27011) );
  XOR U27396 ( .A(b[57]), .B(n28403), .Z(n26993) );
  OR U27397 ( .A(n26993), .B(n965), .Z(n26686) );
  NANDN U27398 ( .A(n26684), .B(n38194), .Z(n26685) );
  NAND U27399 ( .A(n26686), .B(n26685), .Z(n27008) );
  NAND U27400 ( .A(n38326), .B(n26687), .Z(n26689) );
  XNOR U27401 ( .A(n38400), .B(a[63]), .Z(n26996) );
  NANDN U27402 ( .A(n38273), .B(n26996), .Z(n26688) );
  AND U27403 ( .A(n26689), .B(n26688), .Z(n27009) );
  XNOR U27404 ( .A(n27008), .B(n27009), .Z(n27010) );
  XNOR U27405 ( .A(n27011), .B(n27010), .Z(n26857) );
  XNOR U27406 ( .A(b[33]), .B(a[89]), .Z(n26999) );
  NANDN U27407 ( .A(n26999), .B(n35620), .Z(n26692) );
  NANDN U27408 ( .A(n26690), .B(n35621), .Z(n26691) );
  NAND U27409 ( .A(n26692), .B(n26691), .Z(n26872) );
  NANDN U27410 ( .A(n966), .B(a[121]), .Z(n26693) );
  XOR U27411 ( .A(n29232), .B(n26693), .Z(n26695) );
  IV U27412 ( .A(a[120]), .Z(n38134) );
  NANDN U27413 ( .A(n38134), .B(n966), .Z(n26694) );
  AND U27414 ( .A(n26695), .B(n26694), .Z(n26869) );
  XNOR U27415 ( .A(b[63]), .B(a[59]), .Z(n27005) );
  NANDN U27416 ( .A(n27005), .B(n38422), .Z(n26698) );
  NANDN U27417 ( .A(n26696), .B(n38423), .Z(n26697) );
  AND U27418 ( .A(n26698), .B(n26697), .Z(n26870) );
  XNOR U27419 ( .A(n26869), .B(n26870), .Z(n26871) );
  XOR U27420 ( .A(n26872), .B(n26871), .Z(n26858) );
  XNOR U27421 ( .A(n26857), .B(n26858), .Z(n26859) );
  NANDN U27422 ( .A(n26700), .B(n26699), .Z(n26704) );
  NAND U27423 ( .A(n26702), .B(n26701), .Z(n26703) );
  NAND U27424 ( .A(n26704), .B(n26703), .Z(n26860) );
  XOR U27425 ( .A(n26859), .B(n26860), .Z(n26920) );
  NANDN U27426 ( .A(n26706), .B(n26705), .Z(n26710) );
  NAND U27427 ( .A(n26708), .B(n26707), .Z(n26709) );
  NAND U27428 ( .A(n26710), .B(n26709), .Z(n26917) );
  NANDN U27429 ( .A(n26712), .B(n26711), .Z(n26716) );
  NAND U27430 ( .A(n26714), .B(n26713), .Z(n26715) );
  AND U27431 ( .A(n26716), .B(n26715), .Z(n26918) );
  XNOR U27432 ( .A(n26917), .B(n26918), .Z(n26919) );
  XNOR U27433 ( .A(n26920), .B(n26919), .Z(n26802) );
  NANDN U27434 ( .A(n26718), .B(n26717), .Z(n26722) );
  NANDN U27435 ( .A(n26720), .B(n26719), .Z(n26721) );
  AND U27436 ( .A(n26722), .B(n26721), .Z(n26803) );
  XNOR U27437 ( .A(n26802), .B(n26803), .Z(n26804) );
  XNOR U27438 ( .A(n26805), .B(n26804), .Z(n26796) );
  NAND U27439 ( .A(n26724), .B(n26723), .Z(n26728) );
  NANDN U27440 ( .A(n26726), .B(n26725), .Z(n26727) );
  AND U27441 ( .A(n26728), .B(n26727), .Z(n26797) );
  XNOR U27442 ( .A(n26796), .B(n26797), .Z(n26798) );
  XNOR U27443 ( .A(n26799), .B(n26798), .Z(n26791) );
  XOR U27444 ( .A(n26790), .B(n26791), .Z(n26793) );
  NANDN U27445 ( .A(n26730), .B(n26729), .Z(n26734) );
  NAND U27446 ( .A(n26732), .B(n26731), .Z(n26733) );
  NAND U27447 ( .A(n26734), .B(n26733), .Z(n26792) );
  XNOR U27448 ( .A(n26793), .B(n26792), .Z(n27045) );
  NANDN U27449 ( .A(n26736), .B(n26735), .Z(n26740) );
  NAND U27450 ( .A(n26738), .B(n26737), .Z(n26739) );
  NAND U27451 ( .A(n26740), .B(n26739), .Z(n26787) );
  NANDN U27452 ( .A(n26742), .B(n26741), .Z(n26746) );
  NANDN U27453 ( .A(n26744), .B(n26743), .Z(n26745) );
  NAND U27454 ( .A(n26746), .B(n26745), .Z(n26785) );
  OR U27455 ( .A(n26748), .B(n26747), .Z(n26752) );
  NAND U27456 ( .A(n26750), .B(n26749), .Z(n26751) );
  AND U27457 ( .A(n26752), .B(n26751), .Z(n26784) );
  XNOR U27458 ( .A(n26785), .B(n26784), .Z(n26786) );
  XNOR U27459 ( .A(n26787), .B(n26786), .Z(n27042) );
  NANDN U27460 ( .A(n26754), .B(n26753), .Z(n26758) );
  NAND U27461 ( .A(n26756), .B(n26755), .Z(n26757) );
  AND U27462 ( .A(n26758), .B(n26757), .Z(n27043) );
  XNOR U27463 ( .A(n27045), .B(n27044), .Z(n27051) );
  NANDN U27464 ( .A(n26764), .B(n26763), .Z(n26768) );
  NANDN U27465 ( .A(n26766), .B(n26765), .Z(n26767) );
  AND U27466 ( .A(n26768), .B(n26767), .Z(n27048) );
  XNOR U27467 ( .A(n27049), .B(n27048), .Z(n27050) );
  XOR U27468 ( .A(n27051), .B(n27050), .Z(n26781) );
  XNOR U27469 ( .A(n26780), .B(n26781), .Z(n26774) );
  XNOR U27470 ( .A(n26775), .B(n26774), .Z(n26776) );
  XNOR U27471 ( .A(n26777), .B(n26776), .Z(n27054) );
  XNOR U27472 ( .A(n27054), .B(sreg[185]), .Z(n27056) );
  NAND U27473 ( .A(n26769), .B(sreg[184]), .Z(n26773) );
  OR U27474 ( .A(n26771), .B(n26770), .Z(n26772) );
  AND U27475 ( .A(n26773), .B(n26772), .Z(n27055) );
  XOR U27476 ( .A(n27056), .B(n27055), .Z(c[185]) );
  NANDN U27477 ( .A(n26779), .B(n26778), .Z(n26783) );
  NANDN U27478 ( .A(n26781), .B(n26780), .Z(n26782) );
  NAND U27479 ( .A(n26783), .B(n26782), .Z(n27059) );
  NANDN U27480 ( .A(n26785), .B(n26784), .Z(n26789) );
  NANDN U27481 ( .A(n26787), .B(n26786), .Z(n26788) );
  NAND U27482 ( .A(n26789), .B(n26788), .Z(n27330) );
  NANDN U27483 ( .A(n26791), .B(n26790), .Z(n26795) );
  OR U27484 ( .A(n26793), .B(n26792), .Z(n26794) );
  AND U27485 ( .A(n26795), .B(n26794), .Z(n27329) );
  XNOR U27486 ( .A(n27330), .B(n27329), .Z(n27331) );
  NANDN U27487 ( .A(n26797), .B(n26796), .Z(n26801) );
  NAND U27488 ( .A(n26799), .B(n26798), .Z(n26800) );
  NAND U27489 ( .A(n26801), .B(n26800), .Z(n27320) );
  NANDN U27490 ( .A(n26807), .B(n26806), .Z(n26811) );
  NANDN U27491 ( .A(n26809), .B(n26808), .Z(n26810) );
  NAND U27492 ( .A(n26811), .B(n26810), .Z(n27287) );
  XOR U27493 ( .A(a[112]), .B(n970), .Z(n27102) );
  OR U27494 ( .A(n27102), .B(n31369), .Z(n26814) );
  NANDN U27495 ( .A(n26812), .B(n31119), .Z(n26813) );
  NAND U27496 ( .A(n26814), .B(n26813), .Z(n27099) );
  XOR U27497 ( .A(b[43]), .B(n32814), .Z(n27105) );
  NANDN U27498 ( .A(n27105), .B(n37068), .Z(n26817) );
  NANDN U27499 ( .A(n26815), .B(n37069), .Z(n26816) );
  NAND U27500 ( .A(n26817), .B(n26816), .Z(n27096) );
  XNOR U27501 ( .A(b[45]), .B(a[78]), .Z(n27108) );
  NANDN U27502 ( .A(n27108), .B(n37261), .Z(n26820) );
  NAND U27503 ( .A(n26818), .B(n37262), .Z(n26819) );
  AND U27504 ( .A(n26820), .B(n26819), .Z(n27097) );
  XNOR U27505 ( .A(n27096), .B(n27097), .Z(n27098) );
  XNOR U27506 ( .A(n27099), .B(n27098), .Z(n27194) );
  XOR U27507 ( .A(n979), .B(n31372), .Z(n27111) );
  NANDN U27508 ( .A(n37756), .B(n27111), .Z(n26823) );
  NANDN U27509 ( .A(n26821), .B(n37652), .Z(n26822) );
  NAND U27510 ( .A(n26823), .B(n26822), .Z(n27072) );
  NAND U27511 ( .A(n37469), .B(n26824), .Z(n26826) );
  XOR U27512 ( .A(b[47]), .B(n31363), .Z(n27114) );
  NANDN U27513 ( .A(n27114), .B(n37471), .Z(n26825) );
  NAND U27514 ( .A(n26826), .B(n26825), .Z(n27069) );
  XOR U27515 ( .A(n37873), .B(n969), .Z(n27117) );
  NAND U27516 ( .A(n30509), .B(n27117), .Z(n26829) );
  NANDN U27517 ( .A(n26827), .B(n30846), .Z(n26828) );
  AND U27518 ( .A(n26829), .B(n26828), .Z(n27070) );
  XNOR U27519 ( .A(n27069), .B(n27070), .Z(n27071) );
  XOR U27520 ( .A(n27072), .B(n27071), .Z(n27195) );
  XNOR U27521 ( .A(n27194), .B(n27195), .Z(n27196) );
  NANDN U27522 ( .A(n26831), .B(n26830), .Z(n26835) );
  NAND U27523 ( .A(n26833), .B(n26832), .Z(n26834) );
  AND U27524 ( .A(n26835), .B(n26834), .Z(n27197) );
  XNOR U27525 ( .A(n27196), .B(n27197), .Z(n27288) );
  XNOR U27526 ( .A(n27287), .B(n27288), .Z(n27289) );
  XNOR U27527 ( .A(b[35]), .B(a[88]), .Z(n27081) );
  NANDN U27528 ( .A(n27081), .B(n35985), .Z(n26838) );
  NAND U27529 ( .A(n26836), .B(n35986), .Z(n26837) );
  NAND U27530 ( .A(n26838), .B(n26837), .Z(n27153) );
  XOR U27531 ( .A(n38046), .B(n31123), .Z(n27075) );
  NAND U27532 ( .A(n27075), .B(n29949), .Z(n26841) );
  NAND U27533 ( .A(n29948), .B(n26839), .Z(n26840) );
  NAND U27534 ( .A(n26841), .B(n26840), .Z(n27150) );
  XOR U27535 ( .A(b[55]), .B(n29868), .Z(n27078) );
  NANDN U27536 ( .A(n27078), .B(n38075), .Z(n26844) );
  NANDN U27537 ( .A(n26842), .B(n38073), .Z(n26843) );
  AND U27538 ( .A(n26844), .B(n26843), .Z(n27151) );
  XNOR U27539 ( .A(n27150), .B(n27151), .Z(n27152) );
  XNOR U27540 ( .A(n27153), .B(n27152), .Z(n27173) );
  NANDN U27541 ( .A(n26846), .B(n26845), .Z(n26850) );
  NAND U27542 ( .A(n26848), .B(n26847), .Z(n26849) );
  NAND U27543 ( .A(n26850), .B(n26849), .Z(n27170) );
  NANDN U27544 ( .A(n26852), .B(n26851), .Z(n26856) );
  NAND U27545 ( .A(n26854), .B(n26853), .Z(n26855) );
  NAND U27546 ( .A(n26856), .B(n26855), .Z(n27171) );
  XNOR U27547 ( .A(n27170), .B(n27171), .Z(n27172) );
  XOR U27548 ( .A(n27173), .B(n27172), .Z(n27290) );
  XNOR U27549 ( .A(n27289), .B(n27290), .Z(n27306) );
  NANDN U27550 ( .A(n26858), .B(n26857), .Z(n26862) );
  NANDN U27551 ( .A(n26860), .B(n26859), .Z(n26861) );
  NAND U27552 ( .A(n26862), .B(n26861), .Z(n27293) );
  NANDN U27553 ( .A(n26864), .B(n26863), .Z(n26868) );
  NAND U27554 ( .A(n26866), .B(n26865), .Z(n26867) );
  NAND U27555 ( .A(n26868), .B(n26867), .Z(n27294) );
  XNOR U27556 ( .A(n27293), .B(n27294), .Z(n27295) );
  NANDN U27557 ( .A(n26870), .B(n26869), .Z(n26874) );
  NAND U27558 ( .A(n26872), .B(n26871), .Z(n26873) );
  NAND U27559 ( .A(n26874), .B(n26873), .Z(n27123) );
  XOR U27560 ( .A(a[108]), .B(n972), .Z(n27147) );
  OR U27561 ( .A(n27147), .B(n32010), .Z(n26877) );
  NANDN U27562 ( .A(n26875), .B(n32011), .Z(n26876) );
  NAND U27563 ( .A(n26877), .B(n26876), .Z(n27218) );
  XNOR U27564 ( .A(n35783), .B(b[25]), .Z(n27141) );
  NANDN U27565 ( .A(n34219), .B(n27141), .Z(n26880) );
  NAND U27566 ( .A(n34217), .B(n26878), .Z(n26879) );
  NAND U27567 ( .A(n26880), .B(n26879), .Z(n27215) );
  XNOR U27568 ( .A(a[106]), .B(b[17]), .Z(n27144) );
  NANDN U27569 ( .A(n27144), .B(n32543), .Z(n26883) );
  NAND U27570 ( .A(n26881), .B(n32541), .Z(n26882) );
  AND U27571 ( .A(n26883), .B(n26882), .Z(n27216) );
  XNOR U27572 ( .A(n27215), .B(n27216), .Z(n27217) );
  XNOR U27573 ( .A(n27218), .B(n27217), .Z(n27245) );
  XOR U27574 ( .A(b[39]), .B(n33185), .Z(n27132) );
  NANDN U27575 ( .A(n27132), .B(n36553), .Z(n26886) );
  NANDN U27576 ( .A(n26884), .B(n36643), .Z(n26885) );
  NAND U27577 ( .A(n26886), .B(n26885), .Z(n27242) );
  XOR U27578 ( .A(b[51]), .B(n30210), .Z(n27135) );
  NANDN U27579 ( .A(n27135), .B(n37803), .Z(n26889) );
  NANDN U27580 ( .A(n26887), .B(n37802), .Z(n26888) );
  NAND U27581 ( .A(n26889), .B(n26888), .Z(n27239) );
  XOR U27582 ( .A(b[53]), .B(n30379), .Z(n27138) );
  NANDN U27583 ( .A(n27138), .B(n37940), .Z(n26892) );
  NANDN U27584 ( .A(n26890), .B(n37941), .Z(n26891) );
  AND U27585 ( .A(n26892), .B(n26891), .Z(n27240) );
  XNOR U27586 ( .A(n27239), .B(n27240), .Z(n27241) );
  XOR U27587 ( .A(n27242), .B(n27241), .Z(n27246) );
  XOR U27588 ( .A(n27245), .B(n27246), .Z(n27248) );
  NANDN U27589 ( .A(n26894), .B(n26893), .Z(n26898) );
  NAND U27590 ( .A(n26896), .B(n26895), .Z(n26897) );
  AND U27591 ( .A(n26898), .B(n26897), .Z(n27247) );
  XOR U27592 ( .A(n27248), .B(n27247), .Z(n27121) );
  NANDN U27593 ( .A(n26900), .B(n26899), .Z(n26904) );
  NAND U27594 ( .A(n26902), .B(n26901), .Z(n26903) );
  AND U27595 ( .A(n26904), .B(n26903), .Z(n27120) );
  XNOR U27596 ( .A(n27121), .B(n27120), .Z(n27122) );
  XOR U27597 ( .A(n27123), .B(n27122), .Z(n27296) );
  XNOR U27598 ( .A(n27295), .B(n27296), .Z(n27305) );
  XOR U27599 ( .A(n27308), .B(n27307), .Z(n27318) );
  NANDN U27600 ( .A(n26906), .B(n26905), .Z(n26910) );
  NANDN U27601 ( .A(n26908), .B(n26907), .Z(n26909) );
  NAND U27602 ( .A(n26910), .B(n26909), .Z(n27301) );
  NANDN U27603 ( .A(n26912), .B(n26911), .Z(n26916) );
  NAND U27604 ( .A(n26914), .B(n26913), .Z(n26915) );
  AND U27605 ( .A(n26916), .B(n26915), .Z(n27299) );
  NANDN U27606 ( .A(n26918), .B(n26917), .Z(n26922) );
  NAND U27607 ( .A(n26920), .B(n26919), .Z(n26921) );
  NAND U27608 ( .A(n26922), .B(n26921), .Z(n27300) );
  XOR U27609 ( .A(n27301), .B(n27302), .Z(n27068) );
  NAND U27610 ( .A(n33283), .B(n26927), .Z(n26929) );
  XOR U27611 ( .A(n36647), .B(n33020), .Z(n27200) );
  NANDN U27612 ( .A(n33021), .B(n27200), .Z(n26928) );
  NAND U27613 ( .A(n26929), .B(n26928), .Z(n27278) );
  XNOR U27614 ( .A(a[102]), .B(b[21]), .Z(n27203) );
  OR U27615 ( .A(n27203), .B(n33634), .Z(n26932) );
  NAND U27616 ( .A(n26930), .B(n33464), .Z(n26931) );
  NAND U27617 ( .A(n26932), .B(n26931), .Z(n27275) );
  NAND U27618 ( .A(n34044), .B(n26933), .Z(n26935) );
  XOR U27619 ( .A(n36100), .B(n34510), .Z(n27206) );
  NANDN U27620 ( .A(n33867), .B(n27206), .Z(n26934) );
  AND U27621 ( .A(n26935), .B(n26934), .Z(n27276) );
  XNOR U27622 ( .A(n27275), .B(n27276), .Z(n27277) );
  XNOR U27623 ( .A(n27278), .B(n27277), .Z(n27090) );
  NANDN U27624 ( .A(n26937), .B(n26936), .Z(n26941) );
  NAND U27625 ( .A(n26939), .B(n26938), .Z(n26940) );
  NAND U27626 ( .A(n26941), .B(n26940), .Z(n27091) );
  XOR U27627 ( .A(n27090), .B(n27091), .Z(n27093) );
  NAND U27628 ( .A(a[58]), .B(b[63]), .Z(n27087) );
  NANDN U27629 ( .A(n26942), .B(n38369), .Z(n26944) );
  XNOR U27630 ( .A(n984), .B(a[62]), .Z(n27212) );
  NANDN U27631 ( .A(n38371), .B(n27212), .Z(n26943) );
  NAND U27632 ( .A(n26944), .B(n26943), .Z(n27085) );
  NANDN U27633 ( .A(n26945), .B(n35311), .Z(n26947) );
  XNOR U27634 ( .A(n973), .B(a[92]), .Z(n27209) );
  NAND U27635 ( .A(n27209), .B(n35313), .Z(n26946) );
  AND U27636 ( .A(n26947), .B(n26946), .Z(n27084) );
  XNOR U27637 ( .A(n27085), .B(n27084), .Z(n27086) );
  XNOR U27638 ( .A(n27087), .B(n27086), .Z(n27092) );
  XNOR U27639 ( .A(n27093), .B(n27092), .Z(n27188) );
  XOR U27640 ( .A(b[37]), .B(n33628), .Z(n27221) );
  NANDN U27641 ( .A(n27221), .B(n36311), .Z(n26950) );
  NANDN U27642 ( .A(n26948), .B(n36309), .Z(n26949) );
  NAND U27643 ( .A(n26950), .B(n26949), .Z(n27254) );
  XOR U27644 ( .A(a[118]), .B(n968), .Z(n27224) );
  OR U27645 ( .A(n27224), .B(n29363), .Z(n26953) );
  NANDN U27646 ( .A(n26951), .B(n29864), .Z(n26952) );
  NAND U27647 ( .A(n26953), .B(n26952), .Z(n27251) );
  XOR U27648 ( .A(n38134), .B(n967), .Z(n27227) );
  NAND U27649 ( .A(n27227), .B(n28939), .Z(n26956) );
  NAND U27650 ( .A(n28938), .B(n26954), .Z(n26955) );
  AND U27651 ( .A(n26956), .B(n26955), .Z(n27252) );
  XNOR U27652 ( .A(n27251), .B(n27252), .Z(n27253) );
  XNOR U27653 ( .A(n27254), .B(n27253), .Z(n27185) );
  XOR U27654 ( .A(a[110]), .B(n971), .Z(n27230) );
  OR U27655 ( .A(n27230), .B(n31550), .Z(n26959) );
  NANDN U27656 ( .A(n26957), .B(n31874), .Z(n26958) );
  NAND U27657 ( .A(n26959), .B(n26958), .Z(n27129) );
  NAND U27658 ( .A(n34848), .B(n26960), .Z(n26962) );
  XOR U27659 ( .A(n35545), .B(n35375), .Z(n27233) );
  NAND U27660 ( .A(n34618), .B(n27233), .Z(n26961) );
  NAND U27661 ( .A(n26962), .B(n26961), .Z(n27126) );
  NAND U27662 ( .A(n35188), .B(n26963), .Z(n26965) );
  XOR U27663 ( .A(n35191), .B(n35540), .Z(n27236) );
  NANDN U27664 ( .A(n34968), .B(n27236), .Z(n26964) );
  AND U27665 ( .A(n26965), .B(n26964), .Z(n27127) );
  XNOR U27666 ( .A(n27126), .B(n27127), .Z(n27128) );
  XNOR U27667 ( .A(n27129), .B(n27128), .Z(n27182) );
  NANDN U27668 ( .A(n26967), .B(n26966), .Z(n26971) );
  NAND U27669 ( .A(n26969), .B(n26968), .Z(n26970) );
  NAND U27670 ( .A(n26971), .B(n26970), .Z(n27183) );
  XNOR U27671 ( .A(n27182), .B(n27183), .Z(n27184) );
  XOR U27672 ( .A(n27185), .B(n27184), .Z(n27189) );
  XNOR U27673 ( .A(n27188), .B(n27189), .Z(n27190) );
  XOR U27674 ( .A(n27191), .B(n27190), .Z(n27169) );
  NANDN U27675 ( .A(n26973), .B(n26972), .Z(n26977) );
  OR U27676 ( .A(n26975), .B(n26974), .Z(n26976) );
  NAND U27677 ( .A(n26977), .B(n26976), .Z(n27167) );
  NANDN U27678 ( .A(n26979), .B(n26978), .Z(n26983) );
  NAND U27679 ( .A(n26981), .B(n26980), .Z(n26982) );
  NAND U27680 ( .A(n26983), .B(n26982), .Z(n27179) );
  NANDN U27681 ( .A(n26985), .B(n26984), .Z(n26989) );
  NAND U27682 ( .A(n26987), .B(n26986), .Z(n26988) );
  NAND U27683 ( .A(n26989), .B(n26988), .Z(n27163) );
  XNOR U27684 ( .A(b[41]), .B(a[82]), .Z(n27272) );
  OR U27685 ( .A(n27272), .B(n36905), .Z(n26992) );
  NAND U27686 ( .A(n26990), .B(n36807), .Z(n26991) );
  NAND U27687 ( .A(n26992), .B(n26991), .Z(n27284) );
  XOR U27688 ( .A(b[57]), .B(n28701), .Z(n27266) );
  OR U27689 ( .A(n27266), .B(n965), .Z(n26995) );
  NANDN U27690 ( .A(n26993), .B(n38194), .Z(n26994) );
  NAND U27691 ( .A(n26995), .B(n26994), .Z(n27281) );
  NAND U27692 ( .A(n38326), .B(n26996), .Z(n26998) );
  XNOR U27693 ( .A(n38400), .B(a[64]), .Z(n27269) );
  NANDN U27694 ( .A(n38273), .B(n27269), .Z(n26997) );
  AND U27695 ( .A(n26998), .B(n26997), .Z(n27282) );
  XNOR U27696 ( .A(n27281), .B(n27282), .Z(n27283) );
  XOR U27697 ( .A(n27284), .B(n27283), .Z(n27161) );
  XOR U27698 ( .A(b[33]), .B(n34851), .Z(n27257) );
  NANDN U27699 ( .A(n27257), .B(n35620), .Z(n27001) );
  NANDN U27700 ( .A(n26999), .B(n35621), .Z(n27000) );
  NAND U27701 ( .A(n27001), .B(n27000), .Z(n27159) );
  NANDN U27702 ( .A(n966), .B(a[122]), .Z(n27002) );
  XOR U27703 ( .A(n29232), .B(n27002), .Z(n27004) );
  NANDN U27704 ( .A(b[0]), .B(a[121]), .Z(n27003) );
  AND U27705 ( .A(n27004), .B(n27003), .Z(n27156) );
  XOR U27706 ( .A(b[63]), .B(n27436), .Z(n27263) );
  NANDN U27707 ( .A(n27263), .B(n38422), .Z(n27007) );
  NANDN U27708 ( .A(n27005), .B(n38423), .Z(n27006) );
  AND U27709 ( .A(n27007), .B(n27006), .Z(n27157) );
  XNOR U27710 ( .A(n27156), .B(n27157), .Z(n27158) );
  XNOR U27711 ( .A(n27159), .B(n27158), .Z(n27160) );
  XOR U27712 ( .A(n27161), .B(n27160), .Z(n27162) );
  XNOR U27713 ( .A(n27163), .B(n27162), .Z(n27177) );
  NANDN U27714 ( .A(n27009), .B(n27008), .Z(n27013) );
  NAND U27715 ( .A(n27011), .B(n27010), .Z(n27012) );
  AND U27716 ( .A(n27013), .B(n27012), .Z(n27176) );
  XNOR U27717 ( .A(n27177), .B(n27176), .Z(n27178) );
  XNOR U27718 ( .A(n27179), .B(n27178), .Z(n27166) );
  XOR U27719 ( .A(n27167), .B(n27166), .Z(n27168) );
  XNOR U27720 ( .A(n27169), .B(n27168), .Z(n27065) );
  NANDN U27721 ( .A(n27015), .B(n27014), .Z(n27019) );
  NANDN U27722 ( .A(n27017), .B(n27016), .Z(n27018) );
  AND U27723 ( .A(n27019), .B(n27018), .Z(n27066) );
  XNOR U27724 ( .A(n27065), .B(n27066), .Z(n27067) );
  XOR U27725 ( .A(n27068), .B(n27067), .Z(n27317) );
  XOR U27726 ( .A(n27318), .B(n27317), .Z(n27319) );
  XNOR U27727 ( .A(n27320), .B(n27319), .Z(n27326) );
  OR U27728 ( .A(n27021), .B(n27020), .Z(n27025) );
  NAND U27729 ( .A(n27023), .B(n27022), .Z(n27024) );
  NAND U27730 ( .A(n27025), .B(n27024), .Z(n27323) );
  NAND U27731 ( .A(n27027), .B(n27026), .Z(n27031) );
  NANDN U27732 ( .A(n27029), .B(n27028), .Z(n27030) );
  NAND U27733 ( .A(n27031), .B(n27030), .Z(n27314) );
  NANDN U27734 ( .A(n27037), .B(n27036), .Z(n27041) );
  NAND U27735 ( .A(n27039), .B(n27038), .Z(n27040) );
  AND U27736 ( .A(n27041), .B(n27040), .Z(n27312) );
  XNOR U27737 ( .A(n27311), .B(n27312), .Z(n27313) );
  XNOR U27738 ( .A(n27314), .B(n27313), .Z(n27324) );
  XNOR U27739 ( .A(n27323), .B(n27324), .Z(n27325) );
  XOR U27740 ( .A(n27326), .B(n27325), .Z(n27332) );
  XNOR U27741 ( .A(n27331), .B(n27332), .Z(n27338) );
  OR U27742 ( .A(n27043), .B(n27042), .Z(n27047) );
  NAND U27743 ( .A(n27045), .B(n27044), .Z(n27046) );
  NAND U27744 ( .A(n27047), .B(n27046), .Z(n27336) );
  NANDN U27745 ( .A(n27049), .B(n27048), .Z(n27053) );
  NANDN U27746 ( .A(n27051), .B(n27050), .Z(n27052) );
  AND U27747 ( .A(n27053), .B(n27052), .Z(n27335) );
  XNOR U27748 ( .A(n27336), .B(n27335), .Z(n27337) );
  XOR U27749 ( .A(n27338), .B(n27337), .Z(n27060) );
  XNOR U27750 ( .A(n27059), .B(n27060), .Z(n27061) );
  XNOR U27751 ( .A(n27062), .B(n27061), .Z(n27341) );
  XNOR U27752 ( .A(n27341), .B(sreg[186]), .Z(n27343) );
  NAND U27753 ( .A(n27054), .B(sreg[185]), .Z(n27058) );
  OR U27754 ( .A(n27056), .B(n27055), .Z(n27057) );
  AND U27755 ( .A(n27058), .B(n27057), .Z(n27342) );
  XOR U27756 ( .A(n27343), .B(n27342), .Z(c[186]) );
  NANDN U27757 ( .A(n27060), .B(n27059), .Z(n27064) );
  NAND U27758 ( .A(n27062), .B(n27061), .Z(n27063) );
  NAND U27759 ( .A(n27064), .B(n27063), .Z(n27349) );
  NANDN U27760 ( .A(n27070), .B(n27069), .Z(n27074) );
  NAND U27761 ( .A(n27072), .B(n27071), .Z(n27073) );
  NAND U27762 ( .A(n27074), .B(n27073), .Z(n27385) );
  XNOR U27763 ( .A(a[117]), .B(n31123), .Z(n27553) );
  NAND U27764 ( .A(n27553), .B(n29949), .Z(n27077) );
  NAND U27765 ( .A(n29948), .B(n27075), .Z(n27076) );
  NAND U27766 ( .A(n27077), .B(n27076), .Z(n27535) );
  XNOR U27767 ( .A(b[55]), .B(a[69]), .Z(n27556) );
  NANDN U27768 ( .A(n27556), .B(n38075), .Z(n27080) );
  NANDN U27769 ( .A(n27078), .B(n38073), .Z(n27079) );
  NAND U27770 ( .A(n27080), .B(n27079), .Z(n27532) );
  XOR U27771 ( .A(b[35]), .B(a[89]), .Z(n27550) );
  NAND U27772 ( .A(n35985), .B(n27550), .Z(n27083) );
  NANDN U27773 ( .A(n27081), .B(n35986), .Z(n27082) );
  AND U27774 ( .A(n27083), .B(n27082), .Z(n27533) );
  XNOR U27775 ( .A(n27532), .B(n27533), .Z(n27534) );
  XNOR U27776 ( .A(n27535), .B(n27534), .Z(n27383) );
  NANDN U27777 ( .A(n27085), .B(n27084), .Z(n27089) );
  NAND U27778 ( .A(n27087), .B(n27086), .Z(n27088) );
  AND U27779 ( .A(n27089), .B(n27088), .Z(n27382) );
  XNOR U27780 ( .A(n27383), .B(n27382), .Z(n27384) );
  XNOR U27781 ( .A(n27385), .B(n27384), .Z(n27595) );
  NANDN U27782 ( .A(n27091), .B(n27090), .Z(n27095) );
  OR U27783 ( .A(n27093), .B(n27092), .Z(n27094) );
  AND U27784 ( .A(n27095), .B(n27094), .Z(n27596) );
  XNOR U27785 ( .A(n27595), .B(n27596), .Z(n27597) );
  NANDN U27786 ( .A(n27097), .B(n27096), .Z(n27101) );
  NAND U27787 ( .A(n27099), .B(n27098), .Z(n27100) );
  NAND U27788 ( .A(n27101), .B(n27100), .Z(n27454) );
  XNOR U27789 ( .A(a[113]), .B(b[11]), .Z(n27580) );
  OR U27790 ( .A(n27580), .B(n31369), .Z(n27104) );
  NANDN U27791 ( .A(n27102), .B(n31119), .Z(n27103) );
  NAND U27792 ( .A(n27104), .B(n27103), .Z(n27568) );
  XNOR U27793 ( .A(b[43]), .B(a[81]), .Z(n27583) );
  NANDN U27794 ( .A(n27583), .B(n37068), .Z(n27107) );
  NANDN U27795 ( .A(n27105), .B(n37069), .Z(n27106) );
  NAND U27796 ( .A(n27107), .B(n27106), .Z(n27565) );
  XOR U27797 ( .A(b[45]), .B(a[79]), .Z(n27586) );
  NAND U27798 ( .A(n27586), .B(n37261), .Z(n27110) );
  NANDN U27799 ( .A(n27108), .B(n37262), .Z(n27109) );
  AND U27800 ( .A(n27110), .B(n27109), .Z(n27566) );
  XNOR U27801 ( .A(n27565), .B(n27566), .Z(n27567) );
  XNOR U27802 ( .A(n27568), .B(n27567), .Z(n27452) );
  NAND U27803 ( .A(n37652), .B(n27111), .Z(n27113) );
  XOR U27804 ( .A(n979), .B(a[75]), .Z(n27571) );
  OR U27805 ( .A(n27571), .B(n37756), .Z(n27112) );
  NAND U27806 ( .A(n27113), .B(n27112), .Z(n27546) );
  NANDN U27807 ( .A(n27114), .B(n37469), .Z(n27116) );
  XNOR U27808 ( .A(b[47]), .B(a[77]), .Z(n27574) );
  NANDN U27809 ( .A(n27574), .B(n37471), .Z(n27115) );
  AND U27810 ( .A(n27116), .B(n27115), .Z(n27545) );
  NAND U27811 ( .A(n30846), .B(n27117), .Z(n27119) );
  XNOR U27812 ( .A(a[115]), .B(n969), .Z(n27577) );
  NAND U27813 ( .A(n30509), .B(n27577), .Z(n27118) );
  NAND U27814 ( .A(n27119), .B(n27118), .Z(n27544) );
  XNOR U27815 ( .A(n27545), .B(n27544), .Z(n27547) );
  XOR U27816 ( .A(n27546), .B(n27547), .Z(n27453) );
  XOR U27817 ( .A(n27452), .B(n27453), .Z(n27455) );
  XOR U27818 ( .A(n27454), .B(n27455), .Z(n27598) );
  XOR U27819 ( .A(n27597), .B(n27598), .Z(n27589) );
  NANDN U27820 ( .A(n27121), .B(n27120), .Z(n27125) );
  NANDN U27821 ( .A(n27123), .B(n27122), .Z(n27124) );
  NAND U27822 ( .A(n27125), .B(n27124), .Z(n27608) );
  NANDN U27823 ( .A(n27127), .B(n27126), .Z(n27131) );
  NAND U27824 ( .A(n27129), .B(n27128), .Z(n27130) );
  NAND U27825 ( .A(n27131), .B(n27130), .Z(n27427) );
  XNOR U27826 ( .A(b[39]), .B(a[85]), .Z(n27508) );
  NANDN U27827 ( .A(n27508), .B(n36553), .Z(n27134) );
  NANDN U27828 ( .A(n27132), .B(n36643), .Z(n27133) );
  NAND U27829 ( .A(n27134), .B(n27133), .Z(n27461) );
  XNOR U27830 ( .A(b[51]), .B(a[73]), .Z(n27511) );
  NANDN U27831 ( .A(n27511), .B(n37803), .Z(n27137) );
  NANDN U27832 ( .A(n27135), .B(n37802), .Z(n27136) );
  NAND U27833 ( .A(n27137), .B(n27136), .Z(n27458) );
  XOR U27834 ( .A(b[53]), .B(n30543), .Z(n27514) );
  NANDN U27835 ( .A(n27514), .B(n37940), .Z(n27140) );
  NANDN U27836 ( .A(n27138), .B(n37941), .Z(n27139) );
  AND U27837 ( .A(n27140), .B(n27139), .Z(n27459) );
  XNOR U27838 ( .A(n27458), .B(n27459), .Z(n27460) );
  XOR U27839 ( .A(n27461), .B(n27460), .Z(n27424) );
  XOR U27840 ( .A(a[99]), .B(b[25]), .Z(n27520) );
  NANDN U27841 ( .A(n34219), .B(n27520), .Z(n27143) );
  NAND U27842 ( .A(n34217), .B(n27141), .Z(n27142) );
  NAND U27843 ( .A(n27143), .B(n27142), .Z(n27433) );
  XOR U27844 ( .A(a[107]), .B(b[17]), .Z(n27523) );
  NAND U27845 ( .A(n27523), .B(n32543), .Z(n27146) );
  NANDN U27846 ( .A(n27144), .B(n32541), .Z(n27145) );
  NAND U27847 ( .A(n27146), .B(n27145), .Z(n27430) );
  XNOR U27848 ( .A(a[109]), .B(b[15]), .Z(n27517) );
  OR U27849 ( .A(n27517), .B(n32010), .Z(n27149) );
  NANDN U27850 ( .A(n27147), .B(n32011), .Z(n27148) );
  AND U27851 ( .A(n27149), .B(n27148), .Z(n27431) );
  XNOR U27852 ( .A(n27430), .B(n27431), .Z(n27432) );
  XOR U27853 ( .A(n27433), .B(n27432), .Z(n27425) );
  XNOR U27854 ( .A(n27424), .B(n27425), .Z(n27426) );
  XNOR U27855 ( .A(n27427), .B(n27426), .Z(n27501) );
  NANDN U27856 ( .A(n27151), .B(n27150), .Z(n27155) );
  NAND U27857 ( .A(n27153), .B(n27152), .Z(n27154) );
  NAND U27858 ( .A(n27155), .B(n27154), .Z(n27498) );
  XNOR U27859 ( .A(n27498), .B(n27499), .Z(n27500) );
  XOR U27860 ( .A(n27501), .B(n27500), .Z(n27606) );
  NANDN U27861 ( .A(n27161), .B(n27160), .Z(n27165) );
  OR U27862 ( .A(n27163), .B(n27162), .Z(n27164) );
  AND U27863 ( .A(n27165), .B(n27164), .Z(n27605) );
  XOR U27864 ( .A(n27606), .B(n27605), .Z(n27607) );
  XOR U27865 ( .A(n27608), .B(n27607), .Z(n27590) );
  XOR U27866 ( .A(n27589), .B(n27590), .Z(n27591) );
  XOR U27867 ( .A(n27591), .B(n27592), .Z(n27353) );
  NANDN U27868 ( .A(n27171), .B(n27170), .Z(n27175) );
  NAND U27869 ( .A(n27173), .B(n27172), .Z(n27174) );
  NAND U27870 ( .A(n27175), .B(n27174), .Z(n27602) );
  NANDN U27871 ( .A(n27177), .B(n27176), .Z(n27181) );
  NANDN U27872 ( .A(n27179), .B(n27178), .Z(n27180) );
  NAND U27873 ( .A(n27181), .B(n27180), .Z(n27599) );
  NANDN U27874 ( .A(n27183), .B(n27182), .Z(n27187) );
  NAND U27875 ( .A(n27185), .B(n27184), .Z(n27186) );
  AND U27876 ( .A(n27187), .B(n27186), .Z(n27600) );
  XNOR U27877 ( .A(n27599), .B(n27600), .Z(n27601) );
  XNOR U27878 ( .A(n27602), .B(n27601), .Z(n27365) );
  NANDN U27879 ( .A(n27189), .B(n27188), .Z(n27193) );
  NANDN U27880 ( .A(n27191), .B(n27190), .Z(n27192) );
  AND U27881 ( .A(n27193), .B(n27192), .Z(n27364) );
  XNOR U27882 ( .A(n27365), .B(n27364), .Z(n27366) );
  NANDN U27883 ( .A(n27195), .B(n27194), .Z(n27199) );
  NAND U27884 ( .A(n27197), .B(n27196), .Z(n27198) );
  NAND U27885 ( .A(n27199), .B(n27198), .Z(n27485) );
  NAND U27886 ( .A(n33283), .B(n27200), .Z(n27202) );
  XNOR U27887 ( .A(a[105]), .B(n33020), .Z(n27443) );
  NANDN U27888 ( .A(n33021), .B(n27443), .Z(n27201) );
  NAND U27889 ( .A(n27202), .B(n27201), .Z(n27391) );
  XOR U27890 ( .A(a[103]), .B(b[21]), .Z(n27446) );
  NANDN U27891 ( .A(n33634), .B(n27446), .Z(n27205) );
  NANDN U27892 ( .A(n27203), .B(n33464), .Z(n27204) );
  NAND U27893 ( .A(n27205), .B(n27204), .Z(n27388) );
  NAND U27894 ( .A(n34044), .B(n27206), .Z(n27208) );
  XNOR U27895 ( .A(a[101]), .B(n34510), .Z(n27449) );
  NANDN U27896 ( .A(n33867), .B(n27449), .Z(n27207) );
  AND U27897 ( .A(n27208), .B(n27207), .Z(n27389) );
  XNOR U27898 ( .A(n27388), .B(n27389), .Z(n27390) );
  XNOR U27899 ( .A(n27391), .B(n27390), .Z(n27538) );
  XOR U27900 ( .A(b[31]), .B(n35377), .Z(n27440) );
  NANDN U27901 ( .A(n27440), .B(n35313), .Z(n27211) );
  NAND U27902 ( .A(n27209), .B(n35311), .Z(n27210) );
  NAND U27903 ( .A(n27211), .B(n27210), .Z(n27562) );
  XNOR U27904 ( .A(b[61]), .B(a[63]), .Z(n27437) );
  OR U27905 ( .A(n27437), .B(n38371), .Z(n27214) );
  NAND U27906 ( .A(n27212), .B(n38369), .Z(n27213) );
  NAND U27907 ( .A(n27214), .B(n27213), .Z(n27559) );
  NANDN U27908 ( .A(n985), .B(a[59]), .Z(n27560) );
  XNOR U27909 ( .A(n27559), .B(n27560), .Z(n27561) );
  XOR U27910 ( .A(n27562), .B(n27561), .Z(n27539) );
  XOR U27911 ( .A(n27538), .B(n27539), .Z(n27541) );
  NANDN U27912 ( .A(n27216), .B(n27215), .Z(n27220) );
  NAND U27913 ( .A(n27218), .B(n27217), .Z(n27219) );
  NAND U27914 ( .A(n27220), .B(n27219), .Z(n27540) );
  XNOR U27915 ( .A(n27541), .B(n27540), .Z(n27482) );
  XNOR U27916 ( .A(b[37]), .B(a[87]), .Z(n27473) );
  NANDN U27917 ( .A(n27473), .B(n36311), .Z(n27223) );
  NANDN U27918 ( .A(n27221), .B(n36309), .Z(n27222) );
  NAND U27919 ( .A(n27223), .B(n27222), .Z(n27415) );
  XOR U27920 ( .A(a[119]), .B(n968), .Z(n27476) );
  OR U27921 ( .A(n27476), .B(n29363), .Z(n27226) );
  NANDN U27922 ( .A(n27224), .B(n29864), .Z(n27225) );
  NAND U27923 ( .A(n27226), .B(n27225), .Z(n27412) );
  XNOR U27924 ( .A(a[121]), .B(n967), .Z(n27479) );
  NAND U27925 ( .A(n27479), .B(n28939), .Z(n27229) );
  NAND U27926 ( .A(n28938), .B(n27227), .Z(n27228) );
  AND U27927 ( .A(n27229), .B(n27228), .Z(n27413) );
  XNOR U27928 ( .A(n27412), .B(n27413), .Z(n27414) );
  XNOR U27929 ( .A(n27415), .B(n27414), .Z(n27379) );
  XNOR U27930 ( .A(a[111]), .B(b[13]), .Z(n27464) );
  OR U27931 ( .A(n27464), .B(n31550), .Z(n27232) );
  NANDN U27932 ( .A(n27230), .B(n31874), .Z(n27231) );
  NAND U27933 ( .A(n27232), .B(n27231), .Z(n27529) );
  NAND U27934 ( .A(n34848), .B(n27233), .Z(n27235) );
  XNOR U27935 ( .A(a[97]), .B(n35375), .Z(n27467) );
  NAND U27936 ( .A(n34618), .B(n27467), .Z(n27234) );
  NAND U27937 ( .A(n27235), .B(n27234), .Z(n27526) );
  NAND U27938 ( .A(n35188), .B(n27236), .Z(n27238) );
  XOR U27939 ( .A(n35540), .B(n35628), .Z(n27470) );
  NANDN U27940 ( .A(n34968), .B(n27470), .Z(n27237) );
  AND U27941 ( .A(n27238), .B(n27237), .Z(n27527) );
  XNOR U27942 ( .A(n27526), .B(n27527), .Z(n27528) );
  XNOR U27943 ( .A(n27529), .B(n27528), .Z(n27376) );
  NANDN U27944 ( .A(n27240), .B(n27239), .Z(n27244) );
  NAND U27945 ( .A(n27242), .B(n27241), .Z(n27243) );
  NAND U27946 ( .A(n27244), .B(n27243), .Z(n27377) );
  XNOR U27947 ( .A(n27376), .B(n27377), .Z(n27378) );
  XOR U27948 ( .A(n27379), .B(n27378), .Z(n27483) );
  XNOR U27949 ( .A(n27482), .B(n27483), .Z(n27484) );
  XOR U27950 ( .A(n27485), .B(n27484), .Z(n27490) );
  NANDN U27951 ( .A(n27246), .B(n27245), .Z(n27250) );
  NANDN U27952 ( .A(n27248), .B(n27247), .Z(n27249) );
  NAND U27953 ( .A(n27250), .B(n27249), .Z(n27489) );
  NANDN U27954 ( .A(n27252), .B(n27251), .Z(n27256) );
  NAND U27955 ( .A(n27254), .B(n27253), .Z(n27255) );
  NAND U27956 ( .A(n27256), .B(n27255), .Z(n27373) );
  XNOR U27957 ( .A(b[33]), .B(a[91]), .Z(n27403) );
  NANDN U27958 ( .A(n27403), .B(n35620), .Z(n27259) );
  NANDN U27959 ( .A(n27257), .B(n35621), .Z(n27258) );
  NAND U27960 ( .A(n27259), .B(n27258), .Z(n27507) );
  NANDN U27961 ( .A(n966), .B(a[123]), .Z(n27260) );
  XOR U27962 ( .A(n29232), .B(n27260), .Z(n27262) );
  IV U27963 ( .A(a[122]), .Z(n38251) );
  NANDN U27964 ( .A(n38251), .B(n966), .Z(n27261) );
  AND U27965 ( .A(n27262), .B(n27261), .Z(n27504) );
  XOR U27966 ( .A(b[63]), .B(n27773), .Z(n27409) );
  NANDN U27967 ( .A(n27409), .B(n38422), .Z(n27265) );
  NANDN U27968 ( .A(n27263), .B(n38423), .Z(n27264) );
  AND U27969 ( .A(n27265), .B(n27264), .Z(n27505) );
  XNOR U27970 ( .A(n27504), .B(n27505), .Z(n27506) );
  XNOR U27971 ( .A(n27507), .B(n27506), .Z(n27497) );
  XOR U27972 ( .A(b[57]), .B(n29372), .Z(n27397) );
  OR U27973 ( .A(n27397), .B(n965), .Z(n27268) );
  NANDN U27974 ( .A(n27266), .B(n38194), .Z(n27267) );
  NAND U27975 ( .A(n27268), .B(n27267), .Z(n27421) );
  NAND U27976 ( .A(n38326), .B(n27269), .Z(n27271) );
  XOR U27977 ( .A(n38400), .B(n28403), .Z(n27400) );
  NANDN U27978 ( .A(n38273), .B(n27400), .Z(n27270) );
  NAND U27979 ( .A(n27271), .B(n27270), .Z(n27418) );
  XOR U27980 ( .A(b[41]), .B(a[83]), .Z(n27394) );
  NANDN U27981 ( .A(n36905), .B(n27394), .Z(n27274) );
  NANDN U27982 ( .A(n27272), .B(n36807), .Z(n27273) );
  AND U27983 ( .A(n27274), .B(n27273), .Z(n27419) );
  XNOR U27984 ( .A(n27418), .B(n27419), .Z(n27420) );
  XNOR U27985 ( .A(n27421), .B(n27420), .Z(n27494) );
  NANDN U27986 ( .A(n27276), .B(n27275), .Z(n27280) );
  NAND U27987 ( .A(n27278), .B(n27277), .Z(n27279) );
  NAND U27988 ( .A(n27280), .B(n27279), .Z(n27495) );
  XNOR U27989 ( .A(n27494), .B(n27495), .Z(n27496) );
  XOR U27990 ( .A(n27497), .B(n27496), .Z(n27370) );
  NANDN U27991 ( .A(n27282), .B(n27281), .Z(n27286) );
  NAND U27992 ( .A(n27284), .B(n27283), .Z(n27285) );
  AND U27993 ( .A(n27286), .B(n27285), .Z(n27371) );
  XOR U27994 ( .A(n27370), .B(n27371), .Z(n27372) );
  XNOR U27995 ( .A(n27373), .B(n27372), .Z(n27488) );
  XNOR U27996 ( .A(n27489), .B(n27488), .Z(n27491) );
  XNOR U27997 ( .A(n27490), .B(n27491), .Z(n27367) );
  XOR U27998 ( .A(n27366), .B(n27367), .Z(n27352) );
  XOR U27999 ( .A(n27353), .B(n27352), .Z(n27354) );
  XOR U28000 ( .A(n27355), .B(n27354), .Z(n27614) );
  NANDN U28001 ( .A(n27288), .B(n27287), .Z(n27292) );
  NAND U28002 ( .A(n27290), .B(n27289), .Z(n27291) );
  NAND U28003 ( .A(n27292), .B(n27291), .Z(n27361) );
  NANDN U28004 ( .A(n27294), .B(n27293), .Z(n27298) );
  NANDN U28005 ( .A(n27296), .B(n27295), .Z(n27297) );
  NAND U28006 ( .A(n27298), .B(n27297), .Z(n27359) );
  OR U28007 ( .A(n27300), .B(n27299), .Z(n27304) );
  NANDN U28008 ( .A(n27302), .B(n27301), .Z(n27303) );
  AND U28009 ( .A(n27304), .B(n27303), .Z(n27358) );
  XNOR U28010 ( .A(n27359), .B(n27358), .Z(n27360) );
  XNOR U28011 ( .A(n27361), .B(n27360), .Z(n27611) );
  NANDN U28012 ( .A(n27306), .B(n27305), .Z(n27310) );
  NANDN U28013 ( .A(n27308), .B(n27307), .Z(n27309) );
  AND U28014 ( .A(n27310), .B(n27309), .Z(n27612) );
  XNOR U28015 ( .A(n27614), .B(n27613), .Z(n27619) );
  NANDN U28016 ( .A(n27312), .B(n27311), .Z(n27316) );
  NAND U28017 ( .A(n27314), .B(n27313), .Z(n27315) );
  NAND U28018 ( .A(n27316), .B(n27315), .Z(n27617) );
  NAND U28019 ( .A(n27318), .B(n27317), .Z(n27322) );
  NAND U28020 ( .A(n27320), .B(n27319), .Z(n27321) );
  NAND U28021 ( .A(n27322), .B(n27321), .Z(n27618) );
  XNOR U28022 ( .A(n27617), .B(n27618), .Z(n27620) );
  XNOR U28023 ( .A(n27619), .B(n27620), .Z(n27623) );
  NANDN U28024 ( .A(n27324), .B(n27323), .Z(n27328) );
  NAND U28025 ( .A(n27326), .B(n27325), .Z(n27327) );
  NAND U28026 ( .A(n27328), .B(n27327), .Z(n27624) );
  XNOR U28027 ( .A(n27623), .B(n27624), .Z(n27625) );
  NANDN U28028 ( .A(n27330), .B(n27329), .Z(n27334) );
  NAND U28029 ( .A(n27332), .B(n27331), .Z(n27333) );
  NAND U28030 ( .A(n27334), .B(n27333), .Z(n27626) );
  XOR U28031 ( .A(n27625), .B(n27626), .Z(n27346) );
  NANDN U28032 ( .A(n27336), .B(n27335), .Z(n27340) );
  NAND U28033 ( .A(n27338), .B(n27337), .Z(n27339) );
  NAND U28034 ( .A(n27340), .B(n27339), .Z(n27347) );
  XNOR U28035 ( .A(n27346), .B(n27347), .Z(n27348) );
  XNOR U28036 ( .A(n27349), .B(n27348), .Z(n27627) );
  XNOR U28037 ( .A(n27627), .B(sreg[187]), .Z(n27629) );
  NAND U28038 ( .A(n27341), .B(sreg[186]), .Z(n27345) );
  OR U28039 ( .A(n27343), .B(n27342), .Z(n27344) );
  AND U28040 ( .A(n27345), .B(n27344), .Z(n27628) );
  XOR U28041 ( .A(n27629), .B(n27628), .Z(c[187]) );
  NANDN U28042 ( .A(n27347), .B(n27346), .Z(n27351) );
  NAND U28043 ( .A(n27349), .B(n27348), .Z(n27350) );
  NAND U28044 ( .A(n27351), .B(n27350), .Z(n27635) );
  NAND U28045 ( .A(n27353), .B(n27352), .Z(n27357) );
  NANDN U28046 ( .A(n27355), .B(n27354), .Z(n27356) );
  NAND U28047 ( .A(n27357), .B(n27356), .Z(n27899) );
  NANDN U28048 ( .A(n27359), .B(n27358), .Z(n27363) );
  NANDN U28049 ( .A(n27361), .B(n27360), .Z(n27362) );
  NAND U28050 ( .A(n27363), .B(n27362), .Z(n27900) );
  XNOR U28051 ( .A(n27899), .B(n27900), .Z(n27901) );
  NANDN U28052 ( .A(n27365), .B(n27364), .Z(n27369) );
  NAND U28053 ( .A(n27367), .B(n27366), .Z(n27368) );
  NAND U28054 ( .A(n27369), .B(n27368), .Z(n27892) );
  NAND U28055 ( .A(n27371), .B(n27370), .Z(n27375) );
  NANDN U28056 ( .A(n27373), .B(n27372), .Z(n27374) );
  NAND U28057 ( .A(n27375), .B(n27374), .Z(n27871) );
  NANDN U28058 ( .A(n27377), .B(n27376), .Z(n27381) );
  NAND U28059 ( .A(n27379), .B(n27378), .Z(n27380) );
  AND U28060 ( .A(n27381), .B(n27380), .Z(n27872) );
  XNOR U28061 ( .A(n27871), .B(n27872), .Z(n27873) );
  NANDN U28062 ( .A(n27383), .B(n27382), .Z(n27387) );
  NAND U28063 ( .A(n27385), .B(n27384), .Z(n27386) );
  NAND U28064 ( .A(n27387), .B(n27386), .Z(n27874) );
  XOR U28065 ( .A(n27873), .B(n27874), .Z(n27858) );
  NANDN U28066 ( .A(n27389), .B(n27388), .Z(n27393) );
  NAND U28067 ( .A(n27391), .B(n27390), .Z(n27392) );
  NAND U28068 ( .A(n27393), .B(n27392), .Z(n27687) );
  XNOR U28069 ( .A(b[41]), .B(a[84]), .Z(n27825) );
  OR U28070 ( .A(n27825), .B(n36905), .Z(n27396) );
  NAND U28071 ( .A(n27394), .B(n36807), .Z(n27395) );
  NAND U28072 ( .A(n27396), .B(n27395), .Z(n27852) );
  XOR U28073 ( .A(b[57]), .B(n29868), .Z(n27828) );
  OR U28074 ( .A(n27828), .B(n965), .Z(n27399) );
  NANDN U28075 ( .A(n27397), .B(n38194), .Z(n27398) );
  NAND U28076 ( .A(n27399), .B(n27398), .Z(n27849) );
  NAND U28077 ( .A(n38326), .B(n27400), .Z(n27402) );
  XOR U28078 ( .A(n38400), .B(n28701), .Z(n27831) );
  NANDN U28079 ( .A(n38273), .B(n27831), .Z(n27401) );
  AND U28080 ( .A(n27402), .B(n27401), .Z(n27850) );
  XNOR U28081 ( .A(n27849), .B(n27850), .Z(n27851) );
  XOR U28082 ( .A(n27852), .B(n27851), .Z(n27684) );
  XOR U28083 ( .A(b[33]), .B(n34852), .Z(n27834) );
  NANDN U28084 ( .A(n27834), .B(n35620), .Z(n27405) );
  NANDN U28085 ( .A(n27403), .B(n35621), .Z(n27404) );
  NAND U28086 ( .A(n27405), .B(n27404), .Z(n27681) );
  NANDN U28087 ( .A(n966), .B(a[124]), .Z(n27406) );
  XOR U28088 ( .A(n29232), .B(n27406), .Z(n27408) );
  NANDN U28089 ( .A(b[0]), .B(a[123]), .Z(n27407) );
  AND U28090 ( .A(n27408), .B(n27407), .Z(n27678) );
  XNOR U28091 ( .A(b[63]), .B(a[62]), .Z(n27840) );
  NANDN U28092 ( .A(n27840), .B(n38422), .Z(n27411) );
  NANDN U28093 ( .A(n27409), .B(n38423), .Z(n27410) );
  AND U28094 ( .A(n27411), .B(n27410), .Z(n27679) );
  XNOR U28095 ( .A(n27678), .B(n27679), .Z(n27680) );
  XOR U28096 ( .A(n27681), .B(n27680), .Z(n27685) );
  XNOR U28097 ( .A(n27684), .B(n27685), .Z(n27686) );
  XNOR U28098 ( .A(n27687), .B(n27686), .Z(n27752) );
  NANDN U28099 ( .A(n27413), .B(n27412), .Z(n27417) );
  NAND U28100 ( .A(n27415), .B(n27414), .Z(n27416) );
  NAND U28101 ( .A(n27417), .B(n27416), .Z(n27749) );
  NANDN U28102 ( .A(n27419), .B(n27418), .Z(n27423) );
  NAND U28103 ( .A(n27421), .B(n27420), .Z(n27422) );
  AND U28104 ( .A(n27423), .B(n27422), .Z(n27750) );
  XNOR U28105 ( .A(n27749), .B(n27750), .Z(n27751) );
  XOR U28106 ( .A(n27752), .B(n27751), .Z(n27637) );
  OR U28107 ( .A(n27425), .B(n27424), .Z(n27429) );
  OR U28108 ( .A(n27427), .B(n27426), .Z(n27428) );
  AND U28109 ( .A(n27429), .B(n27428), .Z(n27636) );
  XOR U28110 ( .A(n27637), .B(n27636), .Z(n27638) );
  NANDN U28111 ( .A(n27431), .B(n27430), .Z(n27435) );
  NAND U28112 ( .A(n27433), .B(n27432), .Z(n27434) );
  NAND U28113 ( .A(n27435), .B(n27434), .Z(n27692) );
  ANDN U28114 ( .B(b[63]), .A(n27436), .Z(n27706) );
  NANDN U28115 ( .A(n27437), .B(n38369), .Z(n27439) );
  XNOR U28116 ( .A(b[61]), .B(a[64]), .Z(n27774) );
  OR U28117 ( .A(n27774), .B(n38371), .Z(n27438) );
  NAND U28118 ( .A(n27439), .B(n27438), .Z(n27704) );
  NANDN U28119 ( .A(n27440), .B(n35311), .Z(n27442) );
  XOR U28120 ( .A(b[31]), .B(n35191), .Z(n27777) );
  NANDN U28121 ( .A(n27777), .B(n35313), .Z(n27441) );
  AND U28122 ( .A(n27442), .B(n27441), .Z(n27703) );
  XNOR U28123 ( .A(n27704), .B(n27703), .Z(n27705) );
  XOR U28124 ( .A(n27706), .B(n27705), .Z(n27690) );
  NAND U28125 ( .A(n33283), .B(n27443), .Z(n27445) );
  XOR U28126 ( .A(n36909), .B(n33020), .Z(n27780) );
  NANDN U28127 ( .A(n33021), .B(n27780), .Z(n27444) );
  NAND U28128 ( .A(n27445), .B(n27444), .Z(n27822) );
  XNOR U28129 ( .A(a[104]), .B(b[21]), .Z(n27783) );
  OR U28130 ( .A(n27783), .B(n33634), .Z(n27448) );
  NAND U28131 ( .A(n27446), .B(n33464), .Z(n27447) );
  NAND U28132 ( .A(n27448), .B(n27447), .Z(n27819) );
  NAND U28133 ( .A(n34044), .B(n27449), .Z(n27451) );
  XOR U28134 ( .A(n36420), .B(n34510), .Z(n27786) );
  NANDN U28135 ( .A(n33867), .B(n27786), .Z(n27450) );
  AND U28136 ( .A(n27451), .B(n27450), .Z(n27820) );
  XNOR U28137 ( .A(n27819), .B(n27820), .Z(n27821) );
  XNOR U28138 ( .A(n27822), .B(n27821), .Z(n27691) );
  XNOR U28139 ( .A(n27690), .B(n27691), .Z(n27693) );
  XNOR U28140 ( .A(n27692), .B(n27693), .Z(n27758) );
  NANDN U28141 ( .A(n27453), .B(n27452), .Z(n27457) );
  OR U28142 ( .A(n27455), .B(n27454), .Z(n27456) );
  NAND U28143 ( .A(n27457), .B(n27456), .Z(n27755) );
  NANDN U28144 ( .A(n27459), .B(n27458), .Z(n27463) );
  NAND U28145 ( .A(n27461), .B(n27460), .Z(n27462) );
  NAND U28146 ( .A(n27463), .B(n27462), .Z(n27746) );
  XOR U28147 ( .A(a[112]), .B(n971), .Z(n27789) );
  OR U28148 ( .A(n27789), .B(n31550), .Z(n27466) );
  NANDN U28149 ( .A(n27464), .B(n31874), .Z(n27465) );
  NAND U28150 ( .A(n27466), .B(n27465), .Z(n27669) );
  NAND U28151 ( .A(n34848), .B(n27467), .Z(n27469) );
  XOR U28152 ( .A(n35783), .B(n35375), .Z(n27792) );
  NAND U28153 ( .A(n34618), .B(n27792), .Z(n27468) );
  NAND U28154 ( .A(n27469), .B(n27468), .Z(n27666) );
  NAND U28155 ( .A(n35188), .B(n27470), .Z(n27472) );
  XOR U28156 ( .A(n35545), .B(n35540), .Z(n27795) );
  NANDN U28157 ( .A(n34968), .B(n27795), .Z(n27471) );
  AND U28158 ( .A(n27472), .B(n27471), .Z(n27667) );
  XNOR U28159 ( .A(n27666), .B(n27667), .Z(n27668) );
  XOR U28160 ( .A(n27669), .B(n27668), .Z(n27743) );
  XOR U28161 ( .A(b[37]), .B(n34048), .Z(n27798) );
  NANDN U28162 ( .A(n27798), .B(n36311), .Z(n27475) );
  NANDN U28163 ( .A(n27473), .B(n36309), .Z(n27474) );
  NAND U28164 ( .A(n27475), .B(n27474), .Z(n27846) );
  XOR U28165 ( .A(a[120]), .B(n968), .Z(n27801) );
  OR U28166 ( .A(n27801), .B(n29363), .Z(n27478) );
  NANDN U28167 ( .A(n27476), .B(n29864), .Z(n27477) );
  NAND U28168 ( .A(n27478), .B(n27477), .Z(n27843) );
  XOR U28169 ( .A(n38251), .B(n967), .Z(n27804) );
  NAND U28170 ( .A(n27804), .B(n28939), .Z(n27481) );
  NAND U28171 ( .A(n28938), .B(n27479), .Z(n27480) );
  AND U28172 ( .A(n27481), .B(n27480), .Z(n27844) );
  XNOR U28173 ( .A(n27843), .B(n27844), .Z(n27845) );
  XOR U28174 ( .A(n27846), .B(n27845), .Z(n27744) );
  XOR U28175 ( .A(n27743), .B(n27744), .Z(n27745) );
  XOR U28176 ( .A(n27746), .B(n27745), .Z(n27756) );
  XNOR U28177 ( .A(n27755), .B(n27756), .Z(n27757) );
  XOR U28178 ( .A(n27758), .B(n27757), .Z(n27639) );
  XNOR U28179 ( .A(n27638), .B(n27639), .Z(n27855) );
  NANDN U28180 ( .A(n27483), .B(n27482), .Z(n27487) );
  NANDN U28181 ( .A(n27485), .B(n27484), .Z(n27486) );
  AND U28182 ( .A(n27487), .B(n27486), .Z(n27856) );
  XNOR U28183 ( .A(n27855), .B(n27856), .Z(n27857) );
  XNOR U28184 ( .A(n27858), .B(n27857), .Z(n27890) );
  NAND U28185 ( .A(n27489), .B(n27488), .Z(n27493) );
  NANDN U28186 ( .A(n27491), .B(n27490), .Z(n27492) );
  NAND U28187 ( .A(n27493), .B(n27492), .Z(n27878) );
  NANDN U28188 ( .A(n27499), .B(n27498), .Z(n27503) );
  NAND U28189 ( .A(n27501), .B(n27500), .Z(n27502) );
  NAND U28190 ( .A(n27503), .B(n27502), .Z(n27866) );
  XNOR U28191 ( .A(n27865), .B(n27866), .Z(n27867) );
  XOR U28192 ( .A(b[39]), .B(n33628), .Z(n27657) );
  NANDN U28193 ( .A(n27657), .B(n36553), .Z(n27510) );
  NANDN U28194 ( .A(n27508), .B(n36643), .Z(n27509) );
  NAND U28195 ( .A(n27510), .B(n27509), .Z(n27810) );
  XOR U28196 ( .A(b[51]), .B(n31372), .Z(n27660) );
  NANDN U28197 ( .A(n27660), .B(n37803), .Z(n27513) );
  NANDN U28198 ( .A(n27511), .B(n37802), .Z(n27512) );
  NAND U28199 ( .A(n27513), .B(n27512), .Z(n27807) );
  XOR U28200 ( .A(b[53]), .B(n30210), .Z(n27663) );
  NANDN U28201 ( .A(n27663), .B(n37940), .Z(n27516) );
  NANDN U28202 ( .A(n27514), .B(n37941), .Z(n27515) );
  AND U28203 ( .A(n27516), .B(n27515), .Z(n27808) );
  XNOR U28204 ( .A(n27807), .B(n27808), .Z(n27809) );
  XNOR U28205 ( .A(n27810), .B(n27809), .Z(n27815) );
  XOR U28206 ( .A(a[110]), .B(n972), .Z(n27648) );
  OR U28207 ( .A(n27648), .B(n32010), .Z(n27519) );
  NANDN U28208 ( .A(n27517), .B(n32011), .Z(n27518) );
  NAND U28209 ( .A(n27519), .B(n27518), .Z(n27770) );
  XNOR U28210 ( .A(n36100), .B(b[25]), .Z(n27651) );
  NANDN U28211 ( .A(n34219), .B(n27651), .Z(n27522) );
  NAND U28212 ( .A(n34217), .B(n27520), .Z(n27521) );
  NAND U28213 ( .A(n27522), .B(n27521), .Z(n27767) );
  XNOR U28214 ( .A(a[108]), .B(b[17]), .Z(n27654) );
  NANDN U28215 ( .A(n27654), .B(n32543), .Z(n27525) );
  NAND U28216 ( .A(n27523), .B(n32541), .Z(n27524) );
  AND U28217 ( .A(n27525), .B(n27524), .Z(n27768) );
  XNOR U28218 ( .A(n27767), .B(n27768), .Z(n27769) );
  XNOR U28219 ( .A(n27770), .B(n27769), .Z(n27813) );
  NANDN U28220 ( .A(n27527), .B(n27526), .Z(n27531) );
  NAND U28221 ( .A(n27529), .B(n27528), .Z(n27530) );
  NAND U28222 ( .A(n27531), .B(n27530), .Z(n27814) );
  XOR U28223 ( .A(n27813), .B(n27814), .Z(n27816) );
  XNOR U28224 ( .A(n27815), .B(n27816), .Z(n27642) );
  NANDN U28225 ( .A(n27533), .B(n27532), .Z(n27537) );
  NAND U28226 ( .A(n27535), .B(n27534), .Z(n27536) );
  AND U28227 ( .A(n27537), .B(n27536), .Z(n27643) );
  XOR U28228 ( .A(n27642), .B(n27643), .Z(n27644) );
  XOR U28229 ( .A(n27645), .B(n27644), .Z(n27868) );
  XNOR U28230 ( .A(n27867), .B(n27868), .Z(n27877) );
  XNOR U28231 ( .A(n27878), .B(n27877), .Z(n27880) );
  NANDN U28232 ( .A(n27539), .B(n27538), .Z(n27543) );
  OR U28233 ( .A(n27541), .B(n27540), .Z(n27542) );
  NAND U28234 ( .A(n27543), .B(n27542), .Z(n27860) );
  NANDN U28235 ( .A(n27545), .B(n27544), .Z(n27549) );
  NAND U28236 ( .A(n27547), .B(n27546), .Z(n27548) );
  NAND U28237 ( .A(n27549), .B(n27548), .Z(n27739) );
  XNOR U28238 ( .A(b[35]), .B(a[90]), .Z(n27694) );
  NANDN U28239 ( .A(n27694), .B(n35985), .Z(n27552) );
  NAND U28240 ( .A(n27550), .B(n35986), .Z(n27551) );
  NAND U28241 ( .A(n27552), .B(n27551), .Z(n27675) );
  XOR U28242 ( .A(n38143), .B(n31123), .Z(n27697) );
  NAND U28243 ( .A(n27697), .B(n29949), .Z(n27555) );
  NAND U28244 ( .A(n29948), .B(n27553), .Z(n27554) );
  NAND U28245 ( .A(n27555), .B(n27554), .Z(n27672) );
  XOR U28246 ( .A(b[55]), .B(n30379), .Z(n27700) );
  NANDN U28247 ( .A(n27700), .B(n38075), .Z(n27558) );
  NANDN U28248 ( .A(n27556), .B(n38073), .Z(n27557) );
  AND U28249 ( .A(n27558), .B(n27557), .Z(n27673) );
  XNOR U28250 ( .A(n27672), .B(n27673), .Z(n27674) );
  XNOR U28251 ( .A(n27675), .B(n27674), .Z(n27737) );
  NANDN U28252 ( .A(n27560), .B(n27559), .Z(n27564) );
  NAND U28253 ( .A(n27562), .B(n27561), .Z(n27563) );
  NAND U28254 ( .A(n27564), .B(n27563), .Z(n27738) );
  XOR U28255 ( .A(n27737), .B(n27738), .Z(n27740) );
  XOR U28256 ( .A(n27739), .B(n27740), .Z(n27859) );
  XNOR U28257 ( .A(n27860), .B(n27859), .Z(n27861) );
  NANDN U28258 ( .A(n27566), .B(n27565), .Z(n27570) );
  NAND U28259 ( .A(n27568), .B(n27567), .Z(n27569) );
  NAND U28260 ( .A(n27570), .B(n27569), .Z(n27764) );
  NANDN U28261 ( .A(n27571), .B(n37652), .Z(n27573) );
  XOR U28262 ( .A(b[49]), .B(n31363), .Z(n27719) );
  OR U28263 ( .A(n27719), .B(n37756), .Z(n27572) );
  NAND U28264 ( .A(n27573), .B(n27572), .Z(n27711) );
  NANDN U28265 ( .A(n27574), .B(n37469), .Z(n27576) );
  XNOR U28266 ( .A(n978), .B(a[78]), .Z(n27722) );
  NAND U28267 ( .A(n27722), .B(n37471), .Z(n27575) );
  NAND U28268 ( .A(n27576), .B(n27575), .Z(n27709) );
  NAND U28269 ( .A(n30846), .B(n27577), .Z(n27579) );
  XNOR U28270 ( .A(n38046), .B(b[9]), .Z(n27725) );
  NAND U28271 ( .A(n30509), .B(n27725), .Z(n27578) );
  NAND U28272 ( .A(n27579), .B(n27578), .Z(n27710) );
  XNOR U28273 ( .A(n27709), .B(n27710), .Z(n27712) );
  XOR U28274 ( .A(n27711), .B(n27712), .Z(n27761) );
  XOR U28275 ( .A(a[114]), .B(n970), .Z(n27728) );
  OR U28276 ( .A(n27728), .B(n31369), .Z(n27582) );
  NANDN U28277 ( .A(n27580), .B(n31119), .Z(n27581) );
  NAND U28278 ( .A(n27582), .B(n27581), .Z(n27716) );
  XOR U28279 ( .A(b[43]), .B(n32815), .Z(n27731) );
  NANDN U28280 ( .A(n27731), .B(n37068), .Z(n27585) );
  NANDN U28281 ( .A(n27583), .B(n37069), .Z(n27584) );
  NAND U28282 ( .A(n27585), .B(n27584), .Z(n27713) );
  XNOR U28283 ( .A(b[45]), .B(a[80]), .Z(n27734) );
  NANDN U28284 ( .A(n27734), .B(n37261), .Z(n27588) );
  NAND U28285 ( .A(n27586), .B(n37262), .Z(n27587) );
  AND U28286 ( .A(n27588), .B(n27587), .Z(n27714) );
  XNOR U28287 ( .A(n27713), .B(n27714), .Z(n27715) );
  XOR U28288 ( .A(n27716), .B(n27715), .Z(n27762) );
  XNOR U28289 ( .A(n27761), .B(n27762), .Z(n27763) );
  XOR U28290 ( .A(n27764), .B(n27763), .Z(n27862) );
  XOR U28291 ( .A(n27861), .B(n27862), .Z(n27879) );
  XNOR U28292 ( .A(n27880), .B(n27879), .Z(n27889) );
  XOR U28293 ( .A(n27890), .B(n27889), .Z(n27891) );
  XNOR U28294 ( .A(n27892), .B(n27891), .Z(n27895) );
  OR U28295 ( .A(n27590), .B(n27589), .Z(n27594) );
  NANDN U28296 ( .A(n27592), .B(n27591), .Z(n27593) );
  NAND U28297 ( .A(n27594), .B(n27593), .Z(n27894) );
  NANDN U28298 ( .A(n27600), .B(n27599), .Z(n27604) );
  NAND U28299 ( .A(n27602), .B(n27601), .Z(n27603) );
  NAND U28300 ( .A(n27604), .B(n27603), .Z(n27883) );
  OR U28301 ( .A(n27606), .B(n27605), .Z(n27610) );
  NAND U28302 ( .A(n27608), .B(n27607), .Z(n27609) );
  AND U28303 ( .A(n27610), .B(n27609), .Z(n27884) );
  XNOR U28304 ( .A(n27883), .B(n27884), .Z(n27885) );
  XOR U28305 ( .A(n27886), .B(n27885), .Z(n27893) );
  XOR U28306 ( .A(n27894), .B(n27893), .Z(n27896) );
  XOR U28307 ( .A(n27895), .B(n27896), .Z(n27902) );
  XNOR U28308 ( .A(n27901), .B(n27902), .Z(n27907) );
  OR U28309 ( .A(n27612), .B(n27611), .Z(n27616) );
  NANDN U28310 ( .A(n27614), .B(n27613), .Z(n27615) );
  NAND U28311 ( .A(n27616), .B(n27615), .Z(n27906) );
  NANDN U28312 ( .A(n27618), .B(n27617), .Z(n27622) );
  NAND U28313 ( .A(n27620), .B(n27619), .Z(n27621) );
  AND U28314 ( .A(n27622), .B(n27621), .Z(n27905) );
  XNOR U28315 ( .A(n27906), .B(n27905), .Z(n27908) );
  XNOR U28316 ( .A(n27907), .B(n27908), .Z(n27632) );
  XNOR U28317 ( .A(n27632), .B(n27633), .Z(n27634) );
  XNOR U28318 ( .A(n27635), .B(n27634), .Z(n27909) );
  XNOR U28319 ( .A(n27909), .B(sreg[188]), .Z(n27911) );
  NAND U28320 ( .A(n27627), .B(sreg[187]), .Z(n27631) );
  OR U28321 ( .A(n27629), .B(n27628), .Z(n27630) );
  AND U28322 ( .A(n27631), .B(n27630), .Z(n27910) );
  XOR U28323 ( .A(n27911), .B(n27910), .Z(c[188]) );
  OR U28324 ( .A(n27637), .B(n27636), .Z(n27641) );
  NAND U28325 ( .A(n27639), .B(n27638), .Z(n27640) );
  AND U28326 ( .A(n27641), .B(n27640), .Z(n27946) );
  NAND U28327 ( .A(n27643), .B(n27642), .Z(n27647) );
  NANDN U28328 ( .A(n27645), .B(n27644), .Z(n27646) );
  NAND U28329 ( .A(n27647), .B(n27646), .Z(n27939) );
  XNOR U28330 ( .A(a[111]), .B(b[15]), .Z(n28092) );
  OR U28331 ( .A(n28092), .B(n32010), .Z(n27650) );
  NANDN U28332 ( .A(n27648), .B(n32011), .Z(n27649) );
  NAND U28333 ( .A(n27650), .B(n27649), .Z(n28038) );
  XOR U28334 ( .A(a[101]), .B(b[25]), .Z(n28086) );
  NANDN U28335 ( .A(n34219), .B(n28086), .Z(n27653) );
  NAND U28336 ( .A(n34217), .B(n27651), .Z(n27652) );
  NAND U28337 ( .A(n27653), .B(n27652), .Z(n28035) );
  XOR U28338 ( .A(a[109]), .B(b[17]), .Z(n28089) );
  NAND U28339 ( .A(n28089), .B(n32543), .Z(n27656) );
  NANDN U28340 ( .A(n27654), .B(n32541), .Z(n27655) );
  AND U28341 ( .A(n27656), .B(n27655), .Z(n28036) );
  XNOR U28342 ( .A(n28035), .B(n28036), .Z(n28037) );
  XNOR U28343 ( .A(n28038), .B(n28037), .Z(n27978) );
  XNOR U28344 ( .A(b[39]), .B(a[87]), .Z(n28077) );
  NANDN U28345 ( .A(n28077), .B(n36553), .Z(n27659) );
  NANDN U28346 ( .A(n27657), .B(n36643), .Z(n27658) );
  NAND U28347 ( .A(n27659), .B(n27658), .Z(n28068) );
  XNOR U28348 ( .A(b[51]), .B(a[75]), .Z(n28080) );
  NANDN U28349 ( .A(n28080), .B(n37803), .Z(n27662) );
  NANDN U28350 ( .A(n27660), .B(n37802), .Z(n27661) );
  NAND U28351 ( .A(n27662), .B(n27661), .Z(n28065) );
  XNOR U28352 ( .A(b[53]), .B(a[73]), .Z(n28083) );
  NANDN U28353 ( .A(n28083), .B(n37940), .Z(n27665) );
  NANDN U28354 ( .A(n27663), .B(n37941), .Z(n27664) );
  AND U28355 ( .A(n27665), .B(n27664), .Z(n28066) );
  XNOR U28356 ( .A(n28065), .B(n28066), .Z(n28067) );
  XOR U28357 ( .A(n28068), .B(n28067), .Z(n27979) );
  XOR U28358 ( .A(n27978), .B(n27979), .Z(n27981) );
  NANDN U28359 ( .A(n27667), .B(n27666), .Z(n27671) );
  NAND U28360 ( .A(n27669), .B(n27668), .Z(n27670) );
  NAND U28361 ( .A(n27671), .B(n27670), .Z(n27980) );
  XNOR U28362 ( .A(n27981), .B(n27980), .Z(n28122) );
  NANDN U28363 ( .A(n27673), .B(n27672), .Z(n27677) );
  NAND U28364 ( .A(n27675), .B(n27674), .Z(n27676) );
  NAND U28365 ( .A(n27677), .B(n27676), .Z(n28119) );
  NANDN U28366 ( .A(n27679), .B(n27678), .Z(n27683) );
  NAND U28367 ( .A(n27681), .B(n27680), .Z(n27682) );
  AND U28368 ( .A(n27683), .B(n27682), .Z(n28120) );
  XNOR U28369 ( .A(n28119), .B(n28120), .Z(n28121) );
  XNOR U28370 ( .A(n28122), .B(n28121), .Z(n27936) );
  OR U28371 ( .A(n27685), .B(n27684), .Z(n27689) );
  OR U28372 ( .A(n27687), .B(n27686), .Z(n27688) );
  AND U28373 ( .A(n27689), .B(n27688), .Z(n27937) );
  XNOR U28374 ( .A(n27936), .B(n27937), .Z(n27938) );
  XNOR U28375 ( .A(n27939), .B(n27938), .Z(n27947) );
  XNOR U28376 ( .A(n27946), .B(n27947), .Z(n27949) );
  XOR U28377 ( .A(b[35]), .B(a[91]), .Z(n28141) );
  NAND U28378 ( .A(n35985), .B(n28141), .Z(n27696) );
  NANDN U28379 ( .A(n27694), .B(n35986), .Z(n27695) );
  NAND U28380 ( .A(n27696), .B(n27695), .Z(n28104) );
  XOR U28381 ( .A(n38193), .B(n31123), .Z(n28135) );
  NAND U28382 ( .A(n28135), .B(n29949), .Z(n27699) );
  NAND U28383 ( .A(n29948), .B(n27697), .Z(n27698) );
  NAND U28384 ( .A(n27699), .B(n27698), .Z(n28101) );
  XOR U28385 ( .A(b[55]), .B(n30543), .Z(n28138) );
  NANDN U28386 ( .A(n28138), .B(n38075), .Z(n27702) );
  NANDN U28387 ( .A(n27700), .B(n38073), .Z(n27701) );
  AND U28388 ( .A(n27702), .B(n27701), .Z(n28102) );
  XNOR U28389 ( .A(n28101), .B(n28102), .Z(n28103) );
  XNOR U28390 ( .A(n28104), .B(n28103), .Z(n27959) );
  NANDN U28391 ( .A(n27704), .B(n27703), .Z(n27708) );
  NANDN U28392 ( .A(n27706), .B(n27705), .Z(n27707) );
  NAND U28393 ( .A(n27708), .B(n27707), .Z(n27956) );
  XNOR U28394 ( .A(n27956), .B(n27957), .Z(n27958) );
  XOR U28395 ( .A(n27959), .B(n27958), .Z(n27942) );
  XNOR U28396 ( .A(n27943), .B(n27942), .Z(n27944) );
  NANDN U28397 ( .A(n27714), .B(n27713), .Z(n27718) );
  NAND U28398 ( .A(n27716), .B(n27715), .Z(n27717) );
  NAND U28399 ( .A(n27718), .B(n27717), .Z(n28043) );
  XNOR U28400 ( .A(b[49]), .B(a[77]), .Z(n28156) );
  OR U28401 ( .A(n28156), .B(n37756), .Z(n27721) );
  NANDN U28402 ( .A(n27719), .B(n37652), .Z(n27720) );
  NAND U28403 ( .A(n27721), .B(n27720), .Z(n28146) );
  NAND U28404 ( .A(n27722), .B(n37469), .Z(n27724) );
  XNOR U28405 ( .A(n978), .B(a[79]), .Z(n28159) );
  NAND U28406 ( .A(n28159), .B(n37471), .Z(n27723) );
  AND U28407 ( .A(n27724), .B(n27723), .Z(n28144) );
  XNOR U28408 ( .A(a[117]), .B(b[9]), .Z(n28162) );
  NANDN U28409 ( .A(n28162), .B(n30509), .Z(n27727) );
  NAND U28410 ( .A(n27725), .B(n30846), .Z(n27726) );
  AND U28411 ( .A(n27727), .B(n27726), .Z(n28145) );
  XOR U28412 ( .A(n28146), .B(n28147), .Z(n28041) );
  XNOR U28413 ( .A(a[115]), .B(b[11]), .Z(n28165) );
  OR U28414 ( .A(n28165), .B(n31369), .Z(n27730) );
  NANDN U28415 ( .A(n27728), .B(n31119), .Z(n27729) );
  NAND U28416 ( .A(n27730), .B(n27729), .Z(n28153) );
  XNOR U28417 ( .A(b[43]), .B(a[83]), .Z(n28168) );
  NANDN U28418 ( .A(n28168), .B(n37068), .Z(n27733) );
  NANDN U28419 ( .A(n27731), .B(n37069), .Z(n27732) );
  NAND U28420 ( .A(n27733), .B(n27732), .Z(n28150) );
  XOR U28421 ( .A(b[45]), .B(a[81]), .Z(n28171) );
  NAND U28422 ( .A(n28171), .B(n37261), .Z(n27736) );
  NANDN U28423 ( .A(n27734), .B(n37262), .Z(n27735) );
  AND U28424 ( .A(n27736), .B(n27735), .Z(n28151) );
  XNOR U28425 ( .A(n28150), .B(n28151), .Z(n28152) );
  XOR U28426 ( .A(n28153), .B(n28152), .Z(n28042) );
  XOR U28427 ( .A(n28041), .B(n28042), .Z(n28044) );
  XOR U28428 ( .A(n28043), .B(n28044), .Z(n27945) );
  XOR U28429 ( .A(n27944), .B(n27945), .Z(n27948) );
  NANDN U28430 ( .A(n27738), .B(n27737), .Z(n27742) );
  OR U28431 ( .A(n27740), .B(n27739), .Z(n27741) );
  NAND U28432 ( .A(n27742), .B(n27741), .Z(n27934) );
  OR U28433 ( .A(n27744), .B(n27743), .Z(n27748) );
  NANDN U28434 ( .A(n27746), .B(n27745), .Z(n27747) );
  NAND U28435 ( .A(n27748), .B(n27747), .Z(n27932) );
  NANDN U28436 ( .A(n27750), .B(n27749), .Z(n27754) );
  NAND U28437 ( .A(n27752), .B(n27751), .Z(n27753) );
  NAND U28438 ( .A(n27754), .B(n27753), .Z(n27933) );
  XNOR U28439 ( .A(n27932), .B(n27933), .Z(n27935) );
  XOR U28440 ( .A(n27934), .B(n27935), .Z(n27954) );
  NANDN U28441 ( .A(n27756), .B(n27755), .Z(n27760) );
  NAND U28442 ( .A(n27758), .B(n27757), .Z(n27759) );
  NAND U28443 ( .A(n27760), .B(n27759), .Z(n27952) );
  NANDN U28444 ( .A(n27762), .B(n27761), .Z(n27766) );
  NANDN U28445 ( .A(n27764), .B(n27763), .Z(n27765) );
  NAND U28446 ( .A(n27766), .B(n27765), .Z(n27977) );
  NANDN U28447 ( .A(n27768), .B(n27767), .Z(n27772) );
  NAND U28448 ( .A(n27770), .B(n27769), .Z(n27771) );
  NAND U28449 ( .A(n27772), .B(n27771), .Z(n28127) );
  ANDN U28450 ( .B(b[63]), .A(n27773), .Z(n28132) );
  NANDN U28451 ( .A(n27774), .B(n38369), .Z(n27776) );
  XNOR U28452 ( .A(n984), .B(a[65]), .Z(n28023) );
  NANDN U28453 ( .A(n38371), .B(n28023), .Z(n27775) );
  NAND U28454 ( .A(n27776), .B(n27775), .Z(n28130) );
  NANDN U28455 ( .A(n27777), .B(n35311), .Z(n27779) );
  XNOR U28456 ( .A(n973), .B(a[95]), .Z(n28020) );
  NAND U28457 ( .A(n28020), .B(n35313), .Z(n27778) );
  AND U28458 ( .A(n27779), .B(n27778), .Z(n28129) );
  XNOR U28459 ( .A(n28130), .B(n28129), .Z(n28131) );
  XOR U28460 ( .A(n28132), .B(n28131), .Z(n28125) );
  NAND U28461 ( .A(n33283), .B(n27780), .Z(n27782) );
  XNOR U28462 ( .A(a[107]), .B(n33020), .Z(n28026) );
  NANDN U28463 ( .A(n33021), .B(n28026), .Z(n27781) );
  NAND U28464 ( .A(n27782), .B(n27781), .Z(n28005) );
  XOR U28465 ( .A(a[105]), .B(b[21]), .Z(n28029) );
  NANDN U28466 ( .A(n33634), .B(n28029), .Z(n27785) );
  NANDN U28467 ( .A(n27783), .B(n33464), .Z(n27784) );
  NAND U28468 ( .A(n27785), .B(n27784), .Z(n28002) );
  NAND U28469 ( .A(n34044), .B(n27786), .Z(n27788) );
  XNOR U28470 ( .A(a[103]), .B(n34510), .Z(n28032) );
  NANDN U28471 ( .A(n33867), .B(n28032), .Z(n27787) );
  AND U28472 ( .A(n27788), .B(n27787), .Z(n28003) );
  XNOR U28473 ( .A(n28002), .B(n28003), .Z(n28004) );
  XNOR U28474 ( .A(n28005), .B(n28004), .Z(n28126) );
  XNOR U28475 ( .A(n28125), .B(n28126), .Z(n28128) );
  XNOR U28476 ( .A(n28127), .B(n28128), .Z(n27974) );
  XNOR U28477 ( .A(a[113]), .B(b[13]), .Z(n28056) );
  OR U28478 ( .A(n28056), .B(n31550), .Z(n27791) );
  NANDN U28479 ( .A(n27789), .B(n31874), .Z(n27790) );
  NAND U28480 ( .A(n27791), .B(n27790), .Z(n28098) );
  NAND U28481 ( .A(n34848), .B(n27792), .Z(n27794) );
  XNOR U28482 ( .A(a[99]), .B(n35375), .Z(n28059) );
  NAND U28483 ( .A(n34618), .B(n28059), .Z(n27793) );
  NAND U28484 ( .A(n27794), .B(n27793), .Z(n28095) );
  NAND U28485 ( .A(n35188), .B(n27795), .Z(n27797) );
  XNOR U28486 ( .A(a[97]), .B(n35540), .Z(n28062) );
  NANDN U28487 ( .A(n34968), .B(n28062), .Z(n27796) );
  AND U28488 ( .A(n27797), .B(n27796), .Z(n28096) );
  XNOR U28489 ( .A(n28095), .B(n28096), .Z(n28097) );
  XOR U28490 ( .A(n28098), .B(n28097), .Z(n27964) );
  XNOR U28491 ( .A(b[37]), .B(a[89]), .Z(n28047) );
  NANDN U28492 ( .A(n28047), .B(n36311), .Z(n27800) );
  NANDN U28493 ( .A(n27798), .B(n36309), .Z(n27799) );
  NAND U28494 ( .A(n27800), .B(n27799), .Z(n28011) );
  XNOR U28495 ( .A(a[121]), .B(b[5]), .Z(n28050) );
  OR U28496 ( .A(n28050), .B(n29363), .Z(n27803) );
  NANDN U28497 ( .A(n27801), .B(n29864), .Z(n27802) );
  NAND U28498 ( .A(n27803), .B(n27802), .Z(n28008) );
  XNOR U28499 ( .A(a[123]), .B(n967), .Z(n28053) );
  NAND U28500 ( .A(n28053), .B(n28939), .Z(n27806) );
  NAND U28501 ( .A(n28938), .B(n27804), .Z(n27805) );
  AND U28502 ( .A(n27806), .B(n27805), .Z(n28009) );
  XNOR U28503 ( .A(n28008), .B(n28009), .Z(n28010) );
  XOR U28504 ( .A(n28011), .B(n28010), .Z(n27962) );
  NANDN U28505 ( .A(n27808), .B(n27807), .Z(n27812) );
  NAND U28506 ( .A(n27810), .B(n27809), .Z(n27811) );
  NAND U28507 ( .A(n27812), .B(n27811), .Z(n27963) );
  XNOR U28508 ( .A(n27962), .B(n27963), .Z(n27965) );
  XNOR U28509 ( .A(n27964), .B(n27965), .Z(n27975) );
  XNOR U28510 ( .A(n27974), .B(n27975), .Z(n27976) );
  XNOR U28511 ( .A(n27977), .B(n27976), .Z(n28074) );
  NANDN U28512 ( .A(n27814), .B(n27813), .Z(n27818) );
  NANDN U28513 ( .A(n27816), .B(n27815), .Z(n27817) );
  NAND U28514 ( .A(n27818), .B(n27817), .Z(n28072) );
  NANDN U28515 ( .A(n27820), .B(n27819), .Z(n27824) );
  NAND U28516 ( .A(n27822), .B(n27821), .Z(n27823) );
  NAND U28517 ( .A(n27824), .B(n27823), .Z(n28116) );
  XOR U28518 ( .A(b[41]), .B(a[85]), .Z(n27999) );
  NANDN U28519 ( .A(n36905), .B(n27999), .Z(n27827) );
  NANDN U28520 ( .A(n27825), .B(n36807), .Z(n27826) );
  NAND U28521 ( .A(n27827), .B(n27826), .Z(n28017) );
  XNOR U28522 ( .A(b[57]), .B(a[69]), .Z(n27993) );
  OR U28523 ( .A(n27993), .B(n965), .Z(n27830) );
  NANDN U28524 ( .A(n27828), .B(n38194), .Z(n27829) );
  NAND U28525 ( .A(n27830), .B(n27829), .Z(n28014) );
  NAND U28526 ( .A(n38326), .B(n27831), .Z(n27833) );
  XOR U28527 ( .A(n38400), .B(n29372), .Z(n27996) );
  NANDN U28528 ( .A(n38273), .B(n27996), .Z(n27832) );
  AND U28529 ( .A(n27833), .B(n27832), .Z(n28015) );
  XNOR U28530 ( .A(n28014), .B(n28015), .Z(n28016) );
  XOR U28531 ( .A(n28017), .B(n28016), .Z(n28113) );
  XOR U28532 ( .A(b[33]), .B(n35377), .Z(n27984) );
  NANDN U28533 ( .A(n27984), .B(n35620), .Z(n27836) );
  NANDN U28534 ( .A(n27834), .B(n35621), .Z(n27835) );
  NAND U28535 ( .A(n27836), .B(n27835), .Z(n28110) );
  NANDN U28536 ( .A(n966), .B(a[125]), .Z(n27837) );
  XOR U28537 ( .A(n29232), .B(n27837), .Z(n27839) );
  IV U28538 ( .A(a[124]), .Z(n38321) );
  NANDN U28539 ( .A(n38321), .B(n966), .Z(n27838) );
  AND U28540 ( .A(n27839), .B(n27838), .Z(n28107) );
  XNOR U28541 ( .A(b[63]), .B(a[63]), .Z(n27990) );
  NANDN U28542 ( .A(n27990), .B(n38422), .Z(n27842) );
  NANDN U28543 ( .A(n27840), .B(n38423), .Z(n27841) );
  AND U28544 ( .A(n27842), .B(n27841), .Z(n28108) );
  XNOR U28545 ( .A(n28107), .B(n28108), .Z(n28109) );
  XOR U28546 ( .A(n28110), .B(n28109), .Z(n28114) );
  XNOR U28547 ( .A(n28113), .B(n28114), .Z(n28115) );
  XNOR U28548 ( .A(n28116), .B(n28115), .Z(n27971) );
  NANDN U28549 ( .A(n27844), .B(n27843), .Z(n27848) );
  NAND U28550 ( .A(n27846), .B(n27845), .Z(n27847) );
  NAND U28551 ( .A(n27848), .B(n27847), .Z(n27968) );
  NANDN U28552 ( .A(n27850), .B(n27849), .Z(n27854) );
  NAND U28553 ( .A(n27852), .B(n27851), .Z(n27853) );
  AND U28554 ( .A(n27854), .B(n27853), .Z(n27969) );
  XNOR U28555 ( .A(n27968), .B(n27969), .Z(n27970) );
  XOR U28556 ( .A(n27971), .B(n27970), .Z(n28071) );
  XNOR U28557 ( .A(n28072), .B(n28071), .Z(n28073) );
  XOR U28558 ( .A(n28074), .B(n28073), .Z(n27953) );
  XNOR U28559 ( .A(n27952), .B(n27953), .Z(n27955) );
  XOR U28560 ( .A(n27954), .B(n27955), .Z(n28180) );
  XNOR U28561 ( .A(n28181), .B(n28180), .Z(n28182) );
  XNOR U28562 ( .A(n28182), .B(n28183), .Z(n27928) );
  NAND U28563 ( .A(n27860), .B(n27859), .Z(n27864) );
  OR U28564 ( .A(n27862), .B(n27861), .Z(n27863) );
  NAND U28565 ( .A(n27864), .B(n27863), .Z(n28177) );
  NANDN U28566 ( .A(n27866), .B(n27865), .Z(n27870) );
  NANDN U28567 ( .A(n27868), .B(n27867), .Z(n27869) );
  NAND U28568 ( .A(n27870), .B(n27869), .Z(n28174) );
  NANDN U28569 ( .A(n27872), .B(n27871), .Z(n27876) );
  NANDN U28570 ( .A(n27874), .B(n27873), .Z(n27875) );
  AND U28571 ( .A(n27876), .B(n27875), .Z(n28175) );
  XNOR U28572 ( .A(n28174), .B(n28175), .Z(n28176) );
  XNOR U28573 ( .A(n28177), .B(n28176), .Z(n27926) );
  NAND U28574 ( .A(n27878), .B(n27877), .Z(n27882) );
  NANDN U28575 ( .A(n27880), .B(n27879), .Z(n27881) );
  NAND U28576 ( .A(n27882), .B(n27881), .Z(n27927) );
  XOR U28577 ( .A(n27926), .B(n27927), .Z(n27929) );
  NANDN U28578 ( .A(n27884), .B(n27883), .Z(n27888) );
  NAND U28579 ( .A(n27886), .B(n27885), .Z(n27887) );
  NAND U28580 ( .A(n27888), .B(n27887), .Z(n27920) );
  XNOR U28581 ( .A(n27920), .B(n27921), .Z(n27922) );
  XOR U28582 ( .A(n27923), .B(n27922), .Z(n28186) );
  NANDN U28583 ( .A(n27894), .B(n27893), .Z(n27898) );
  OR U28584 ( .A(n27896), .B(n27895), .Z(n27897) );
  NAND U28585 ( .A(n27898), .B(n27897), .Z(n28187) );
  XOR U28586 ( .A(n28186), .B(n28187), .Z(n28188) );
  NANDN U28587 ( .A(n27900), .B(n27899), .Z(n27904) );
  NAND U28588 ( .A(n27902), .B(n27901), .Z(n27903) );
  NAND U28589 ( .A(n27904), .B(n27903), .Z(n28189) );
  XOR U28590 ( .A(n28188), .B(n28189), .Z(n27914) );
  XNOR U28591 ( .A(n27914), .B(n27915), .Z(n27916) );
  XNOR U28592 ( .A(n27917), .B(n27916), .Z(n28192) );
  XNOR U28593 ( .A(n28192), .B(sreg[189]), .Z(n28194) );
  NAND U28594 ( .A(n27909), .B(sreg[188]), .Z(n27913) );
  OR U28595 ( .A(n27911), .B(n27910), .Z(n27912) );
  AND U28596 ( .A(n27913), .B(n27912), .Z(n28193) );
  XOR U28597 ( .A(n28194), .B(n28193), .Z(c[189]) );
  NANDN U28598 ( .A(n27915), .B(n27914), .Z(n27919) );
  NAND U28599 ( .A(n27917), .B(n27916), .Z(n27918) );
  NAND U28600 ( .A(n27919), .B(n27918), .Z(n28200) );
  NANDN U28601 ( .A(n27921), .B(n27920), .Z(n27925) );
  NAND U28602 ( .A(n27923), .B(n27922), .Z(n27924) );
  NAND U28603 ( .A(n27925), .B(n27924), .Z(n28203) );
  NANDN U28604 ( .A(n27927), .B(n27926), .Z(n27931) );
  OR U28605 ( .A(n27929), .B(n27928), .Z(n27930) );
  NAND U28606 ( .A(n27931), .B(n27930), .Z(n28204) );
  XNOR U28607 ( .A(n28203), .B(n28204), .Z(n28205) );
  NANDN U28608 ( .A(n27937), .B(n27936), .Z(n27941) );
  NAND U28609 ( .A(n27939), .B(n27938), .Z(n27940) );
  AND U28610 ( .A(n27941), .B(n27940), .Z(n28454) );
  XNOR U28611 ( .A(n28455), .B(n28454), .Z(n28456) );
  XOR U28612 ( .A(n28456), .B(n28457), .Z(n28472) );
  OR U28613 ( .A(n27947), .B(n27946), .Z(n27951) );
  NANDN U28614 ( .A(n27949), .B(n27948), .Z(n27950) );
  AND U28615 ( .A(n27951), .B(n27950), .Z(n28473) );
  XNOR U28616 ( .A(n28472), .B(n28473), .Z(n28475) );
  NANDN U28617 ( .A(n27957), .B(n27956), .Z(n27961) );
  NAND U28618 ( .A(n27959), .B(n27958), .Z(n27960) );
  NAND U28619 ( .A(n27961), .B(n27960), .Z(n28442) );
  OR U28620 ( .A(n27963), .B(n27962), .Z(n27967) );
  OR U28621 ( .A(n27965), .B(n27964), .Z(n27966) );
  NAND U28622 ( .A(n27967), .B(n27966), .Z(n28440) );
  NANDN U28623 ( .A(n27969), .B(n27968), .Z(n27973) );
  NAND U28624 ( .A(n27971), .B(n27970), .Z(n27972) );
  NAND U28625 ( .A(n27973), .B(n27972), .Z(n28441) );
  XNOR U28626 ( .A(n28440), .B(n28441), .Z(n28443) );
  XOR U28627 ( .A(n28442), .B(n28443), .Z(n28211) );
  NANDN U28628 ( .A(n27979), .B(n27978), .Z(n27983) );
  OR U28629 ( .A(n27981), .B(n27980), .Z(n27982) );
  NAND U28630 ( .A(n27983), .B(n27982), .Z(n28213) );
  XOR U28631 ( .A(b[33]), .B(n35191), .Z(n28397) );
  NANDN U28632 ( .A(n28397), .B(n35620), .Z(n27986) );
  NANDN U28633 ( .A(n27984), .B(n35621), .Z(n27985) );
  NAND U28634 ( .A(n27986), .B(n27985), .Z(n28228) );
  NANDN U28635 ( .A(n966), .B(a[126]), .Z(n27987) );
  XOR U28636 ( .A(n29232), .B(n27987), .Z(n27989) );
  NANDN U28637 ( .A(b[0]), .B(a[125]), .Z(n27988) );
  AND U28638 ( .A(n27989), .B(n27988), .Z(n28225) );
  XNOR U28639 ( .A(b[63]), .B(a[64]), .Z(n28404) );
  NANDN U28640 ( .A(n28404), .B(n38422), .Z(n27992) );
  NANDN U28641 ( .A(n27990), .B(n38423), .Z(n27991) );
  AND U28642 ( .A(n27992), .B(n27991), .Z(n28226) );
  XNOR U28643 ( .A(n28225), .B(n28226), .Z(n28227) );
  XNOR U28644 ( .A(n28228), .B(n28227), .Z(n28261) );
  XOR U28645 ( .A(b[57]), .B(n30379), .Z(n28407) );
  OR U28646 ( .A(n28407), .B(n965), .Z(n27995) );
  NANDN U28647 ( .A(n27993), .B(n38194), .Z(n27994) );
  NAND U28648 ( .A(n27995), .B(n27994), .Z(n28431) );
  NAND U28649 ( .A(n38326), .B(n27996), .Z(n27998) );
  XOR U28650 ( .A(n38400), .B(n29868), .Z(n28410) );
  NANDN U28651 ( .A(n38273), .B(n28410), .Z(n27997) );
  NAND U28652 ( .A(n27998), .B(n27997), .Z(n28428) );
  XNOR U28653 ( .A(b[41]), .B(a[86]), .Z(n28413) );
  OR U28654 ( .A(n28413), .B(n36905), .Z(n28001) );
  NAND U28655 ( .A(n27999), .B(n36807), .Z(n28000) );
  AND U28656 ( .A(n28001), .B(n28000), .Z(n28429) );
  XNOR U28657 ( .A(n28428), .B(n28429), .Z(n28430) );
  XOR U28658 ( .A(n28431), .B(n28430), .Z(n28260) );
  NANDN U28659 ( .A(n28003), .B(n28002), .Z(n28007) );
  NAND U28660 ( .A(n28005), .B(n28004), .Z(n28006) );
  NAND U28661 ( .A(n28007), .B(n28006), .Z(n28259) );
  XNOR U28662 ( .A(n28260), .B(n28259), .Z(n28262) );
  XNOR U28663 ( .A(n28261), .B(n28262), .Z(n28325) );
  NANDN U28664 ( .A(n28009), .B(n28008), .Z(n28013) );
  NAND U28665 ( .A(n28011), .B(n28010), .Z(n28012) );
  NAND U28666 ( .A(n28013), .B(n28012), .Z(n28322) );
  NANDN U28667 ( .A(n28015), .B(n28014), .Z(n28019) );
  NAND U28668 ( .A(n28017), .B(n28016), .Z(n28018) );
  AND U28669 ( .A(n28019), .B(n28018), .Z(n28323) );
  XNOR U28670 ( .A(n28322), .B(n28323), .Z(n28324) );
  XNOR U28671 ( .A(n28325), .B(n28324), .Z(n28214) );
  XNOR U28672 ( .A(n28213), .B(n28214), .Z(n28215) );
  XOR U28673 ( .A(b[31]), .B(n35545), .Z(n28352) );
  NANDN U28674 ( .A(n28352), .B(n35313), .Z(n28022) );
  NAND U28675 ( .A(n28020), .B(n35311), .Z(n28021) );
  NAND U28676 ( .A(n28022), .B(n28021), .Z(n28289) );
  XOR U28677 ( .A(b[61]), .B(n28701), .Z(n28355) );
  OR U28678 ( .A(n28355), .B(n38371), .Z(n28025) );
  NAND U28679 ( .A(n28023), .B(n38369), .Z(n28024) );
  NAND U28680 ( .A(n28025), .B(n28024), .Z(n28286) );
  NANDN U28681 ( .A(n985), .B(a[62]), .Z(n28287) );
  XNOR U28682 ( .A(n28286), .B(n28287), .Z(n28288) );
  XNOR U28683 ( .A(n28289), .B(n28288), .Z(n28267) );
  NAND U28684 ( .A(n33283), .B(n28026), .Z(n28028) );
  XOR U28685 ( .A(n37139), .B(n33020), .Z(n28358) );
  NANDN U28686 ( .A(n33021), .B(n28358), .Z(n28027) );
  NAND U28687 ( .A(n28028), .B(n28027), .Z(n28419) );
  XNOR U28688 ( .A(a[106]), .B(b[21]), .Z(n28361) );
  OR U28689 ( .A(n28361), .B(n33634), .Z(n28031) );
  NAND U28690 ( .A(n28029), .B(n33464), .Z(n28030) );
  NAND U28691 ( .A(n28031), .B(n28030), .Z(n28416) );
  NAND U28692 ( .A(n34044), .B(n28032), .Z(n28034) );
  XOR U28693 ( .A(n36647), .B(n34510), .Z(n28364) );
  NANDN U28694 ( .A(n33867), .B(n28364), .Z(n28033) );
  AND U28695 ( .A(n28034), .B(n28033), .Z(n28417) );
  XNOR U28696 ( .A(n28416), .B(n28417), .Z(n28418) );
  XNOR U28697 ( .A(n28419), .B(n28418), .Z(n28265) );
  NANDN U28698 ( .A(n28036), .B(n28035), .Z(n28040) );
  NAND U28699 ( .A(n28038), .B(n28037), .Z(n28039) );
  NAND U28700 ( .A(n28040), .B(n28039), .Z(n28266) );
  XOR U28701 ( .A(n28265), .B(n28266), .Z(n28268) );
  XNOR U28702 ( .A(n28267), .B(n28268), .Z(n28336) );
  NANDN U28703 ( .A(n28042), .B(n28041), .Z(n28046) );
  OR U28704 ( .A(n28044), .B(n28043), .Z(n28045) );
  NAND U28705 ( .A(n28046), .B(n28045), .Z(n28334) );
  XOR U28706 ( .A(b[37]), .B(n34851), .Z(n28367) );
  NANDN U28707 ( .A(n28367), .B(n36311), .Z(n28049) );
  NANDN U28708 ( .A(n28047), .B(n36309), .Z(n28048) );
  NAND U28709 ( .A(n28049), .B(n28048), .Z(n28425) );
  XOR U28710 ( .A(a[122]), .B(n968), .Z(n28370) );
  OR U28711 ( .A(n28370), .B(n29363), .Z(n28052) );
  NANDN U28712 ( .A(n28050), .B(n29864), .Z(n28051) );
  NAND U28713 ( .A(n28052), .B(n28051), .Z(n28422) );
  XOR U28714 ( .A(n38321), .B(n967), .Z(n28373) );
  NAND U28715 ( .A(n28373), .B(n28939), .Z(n28055) );
  NAND U28716 ( .A(n28938), .B(n28053), .Z(n28054) );
  AND U28717 ( .A(n28055), .B(n28054), .Z(n28423) );
  XNOR U28718 ( .A(n28422), .B(n28423), .Z(n28424) );
  XNOR U28719 ( .A(n28425), .B(n28424), .Z(n28328) );
  XOR U28720 ( .A(a[114]), .B(n971), .Z(n28376) );
  OR U28721 ( .A(n28376), .B(n31550), .Z(n28058) );
  NANDN U28722 ( .A(n28056), .B(n31874), .Z(n28057) );
  NAND U28723 ( .A(n28058), .B(n28057), .Z(n28232) );
  NAND U28724 ( .A(n34848), .B(n28059), .Z(n28061) );
  XOR U28725 ( .A(n36100), .B(n35375), .Z(n28379) );
  NAND U28726 ( .A(n34618), .B(n28379), .Z(n28060) );
  NAND U28727 ( .A(n28061), .B(n28060), .Z(n28229) );
  NAND U28728 ( .A(n35188), .B(n28062), .Z(n28064) );
  XOR U28729 ( .A(n35783), .B(n35540), .Z(n28382) );
  NANDN U28730 ( .A(n34968), .B(n28382), .Z(n28063) );
  AND U28731 ( .A(n28064), .B(n28063), .Z(n28230) );
  XNOR U28732 ( .A(n28229), .B(n28230), .Z(n28231) );
  XOR U28733 ( .A(n28232), .B(n28231), .Z(n28329) );
  XOR U28734 ( .A(n28328), .B(n28329), .Z(n28331) );
  NANDN U28735 ( .A(n28066), .B(n28065), .Z(n28070) );
  NAND U28736 ( .A(n28068), .B(n28067), .Z(n28069) );
  AND U28737 ( .A(n28070), .B(n28069), .Z(n28330) );
  XOR U28738 ( .A(n28331), .B(n28330), .Z(n28335) );
  XNOR U28739 ( .A(n28334), .B(n28335), .Z(n28337) );
  XOR U28740 ( .A(n28336), .B(n28337), .Z(n28216) );
  XOR U28741 ( .A(n28215), .B(n28216), .Z(n28209) );
  XOR U28742 ( .A(n28210), .B(n28209), .Z(n28212) );
  XOR U28743 ( .A(n28211), .B(n28212), .Z(n28460) );
  NANDN U28744 ( .A(n28072), .B(n28071), .Z(n28076) );
  NAND U28745 ( .A(n28074), .B(n28073), .Z(n28075) );
  NAND U28746 ( .A(n28076), .B(n28075), .Z(n28435) );
  XOR U28747 ( .A(b[39]), .B(n34048), .Z(n28244) );
  NANDN U28748 ( .A(n28244), .B(n36553), .Z(n28079) );
  NANDN U28749 ( .A(n28077), .B(n36643), .Z(n28078) );
  NAND U28750 ( .A(n28079), .B(n28078), .Z(n28388) );
  XOR U28751 ( .A(b[51]), .B(n31363), .Z(n28247) );
  NANDN U28752 ( .A(n28247), .B(n37803), .Z(n28082) );
  NANDN U28753 ( .A(n28080), .B(n37802), .Z(n28081) );
  NAND U28754 ( .A(n28082), .B(n28081), .Z(n28385) );
  XOR U28755 ( .A(b[53]), .B(n31372), .Z(n28250) );
  NANDN U28756 ( .A(n28250), .B(n37940), .Z(n28085) );
  NANDN U28757 ( .A(n28083), .B(n37941), .Z(n28084) );
  AND U28758 ( .A(n28085), .B(n28084), .Z(n28386) );
  XNOR U28759 ( .A(n28385), .B(n28386), .Z(n28387) );
  XOR U28760 ( .A(n28388), .B(n28387), .Z(n28394) );
  XNOR U28761 ( .A(n36420), .B(b[25]), .Z(n28235) );
  NANDN U28762 ( .A(n34219), .B(n28235), .Z(n28088) );
  NAND U28763 ( .A(n34217), .B(n28086), .Z(n28087) );
  NAND U28764 ( .A(n28088), .B(n28087), .Z(n28349) );
  XNOR U28765 ( .A(a[110]), .B(b[17]), .Z(n28238) );
  NANDN U28766 ( .A(n28238), .B(n32543), .Z(n28091) );
  NAND U28767 ( .A(n28089), .B(n32541), .Z(n28090) );
  NAND U28768 ( .A(n28091), .B(n28090), .Z(n28346) );
  XOR U28769 ( .A(a[112]), .B(n972), .Z(n28241) );
  OR U28770 ( .A(n28241), .B(n32010), .Z(n28094) );
  NANDN U28771 ( .A(n28092), .B(n32011), .Z(n28093) );
  AND U28772 ( .A(n28094), .B(n28093), .Z(n28347) );
  XNOR U28773 ( .A(n28346), .B(n28347), .Z(n28348) );
  XOR U28774 ( .A(n28349), .B(n28348), .Z(n28392) );
  NANDN U28775 ( .A(n28096), .B(n28095), .Z(n28100) );
  NAND U28776 ( .A(n28098), .B(n28097), .Z(n28099) );
  AND U28777 ( .A(n28100), .B(n28099), .Z(n28391) );
  XOR U28778 ( .A(n28392), .B(n28391), .Z(n28393) );
  XOR U28779 ( .A(n28394), .B(n28393), .Z(n28222) );
  NANDN U28780 ( .A(n28102), .B(n28101), .Z(n28106) );
  NAND U28781 ( .A(n28104), .B(n28103), .Z(n28105) );
  NAND U28782 ( .A(n28106), .B(n28105), .Z(n28219) );
  NANDN U28783 ( .A(n28108), .B(n28107), .Z(n28112) );
  NAND U28784 ( .A(n28110), .B(n28109), .Z(n28111) );
  AND U28785 ( .A(n28112), .B(n28111), .Z(n28220) );
  XNOR U28786 ( .A(n28219), .B(n28220), .Z(n28221) );
  XNOR U28787 ( .A(n28222), .B(n28221), .Z(n28447) );
  OR U28788 ( .A(n28114), .B(n28113), .Z(n28118) );
  OR U28789 ( .A(n28116), .B(n28115), .Z(n28117) );
  NAND U28790 ( .A(n28118), .B(n28117), .Z(n28444) );
  NANDN U28791 ( .A(n28120), .B(n28119), .Z(n28124) );
  NAND U28792 ( .A(n28122), .B(n28121), .Z(n28123) );
  NAND U28793 ( .A(n28124), .B(n28123), .Z(n28445) );
  XNOR U28794 ( .A(n28444), .B(n28445), .Z(n28446) );
  XNOR U28795 ( .A(n28447), .B(n28446), .Z(n28434) );
  XOR U28796 ( .A(n28435), .B(n28434), .Z(n28437) );
  NANDN U28797 ( .A(n28130), .B(n28129), .Z(n28134) );
  NANDN U28798 ( .A(n28132), .B(n28131), .Z(n28133) );
  NAND U28799 ( .A(n28134), .B(n28133), .Z(n28316) );
  XOR U28800 ( .A(n38134), .B(n31123), .Z(n28277) );
  NAND U28801 ( .A(n28277), .B(n29949), .Z(n28137) );
  NAND U28802 ( .A(n29948), .B(n28135), .Z(n28136) );
  NAND U28803 ( .A(n28137), .B(n28136), .Z(n28256) );
  XOR U28804 ( .A(b[55]), .B(n30210), .Z(n28280) );
  NANDN U28805 ( .A(n28280), .B(n38075), .Z(n28140) );
  NANDN U28806 ( .A(n28138), .B(n38073), .Z(n28139) );
  NAND U28807 ( .A(n28140), .B(n28139), .Z(n28253) );
  XNOR U28808 ( .A(b[35]), .B(a[92]), .Z(n28283) );
  NANDN U28809 ( .A(n28283), .B(n35985), .Z(n28143) );
  NAND U28810 ( .A(n28141), .B(n35986), .Z(n28142) );
  AND U28811 ( .A(n28143), .B(n28142), .Z(n28254) );
  XNOR U28812 ( .A(n28253), .B(n28254), .Z(n28255) );
  XOR U28813 ( .A(n28256), .B(n28255), .Z(n28317) );
  XNOR U28814 ( .A(n28316), .B(n28317), .Z(n28318) );
  OR U28815 ( .A(n28145), .B(n28144), .Z(n28149) );
  NANDN U28816 ( .A(n28147), .B(n28146), .Z(n28148) );
  AND U28817 ( .A(n28149), .B(n28148), .Z(n28319) );
  XOR U28818 ( .A(n28318), .B(n28319), .Z(n28450) );
  XNOR U28819 ( .A(n28451), .B(n28450), .Z(n28452) );
  NANDN U28820 ( .A(n28151), .B(n28150), .Z(n28155) );
  NAND U28821 ( .A(n28153), .B(n28152), .Z(n28154) );
  NAND U28822 ( .A(n28155), .B(n28154), .Z(n28342) );
  XOR U28823 ( .A(b[49]), .B(n31870), .Z(n28298) );
  OR U28824 ( .A(n28298), .B(n37756), .Z(n28158) );
  NANDN U28825 ( .A(n28156), .B(n37652), .Z(n28157) );
  NAND U28826 ( .A(n28158), .B(n28157), .Z(n28273) );
  NAND U28827 ( .A(n37469), .B(n28159), .Z(n28161) );
  XOR U28828 ( .A(n978), .B(n32814), .Z(n28301) );
  NAND U28829 ( .A(n28301), .B(n37471), .Z(n28160) );
  AND U28830 ( .A(n28161), .B(n28160), .Z(n28271) );
  XOR U28831 ( .A(a[118]), .B(n969), .Z(n28304) );
  NANDN U28832 ( .A(n28304), .B(n30509), .Z(n28164) );
  NANDN U28833 ( .A(n28162), .B(n30846), .Z(n28163) );
  AND U28834 ( .A(n28164), .B(n28163), .Z(n28272) );
  XOR U28835 ( .A(n28273), .B(n28274), .Z(n28340) );
  XOR U28836 ( .A(a[116]), .B(n970), .Z(n28307) );
  OR U28837 ( .A(n28307), .B(n31369), .Z(n28167) );
  NANDN U28838 ( .A(n28165), .B(n31119), .Z(n28166) );
  NAND U28839 ( .A(n28167), .B(n28166), .Z(n28295) );
  XOR U28840 ( .A(b[43]), .B(n33185), .Z(n28310) );
  NANDN U28841 ( .A(n28310), .B(n37068), .Z(n28170) );
  NANDN U28842 ( .A(n28168), .B(n37069), .Z(n28169) );
  NAND U28843 ( .A(n28170), .B(n28169), .Z(n28292) );
  XNOR U28844 ( .A(b[45]), .B(a[82]), .Z(n28313) );
  NANDN U28845 ( .A(n28313), .B(n37261), .Z(n28173) );
  NAND U28846 ( .A(n28171), .B(n37262), .Z(n28172) );
  AND U28847 ( .A(n28173), .B(n28172), .Z(n28293) );
  XNOR U28848 ( .A(n28292), .B(n28293), .Z(n28294) );
  XOR U28849 ( .A(n28295), .B(n28294), .Z(n28341) );
  XOR U28850 ( .A(n28340), .B(n28341), .Z(n28343) );
  XOR U28851 ( .A(n28342), .B(n28343), .Z(n28453) );
  XOR U28852 ( .A(n28452), .B(n28453), .Z(n28436) );
  XNOR U28853 ( .A(n28437), .B(n28436), .Z(n28461) );
  XOR U28854 ( .A(n28460), .B(n28461), .Z(n28462) );
  XNOR U28855 ( .A(n28463), .B(n28462), .Z(n28474) );
  XNOR U28856 ( .A(n28475), .B(n28474), .Z(n28469) );
  NANDN U28857 ( .A(n28175), .B(n28174), .Z(n28179) );
  NAND U28858 ( .A(n28177), .B(n28176), .Z(n28178) );
  NAND U28859 ( .A(n28179), .B(n28178), .Z(n28466) );
  NANDN U28860 ( .A(n28181), .B(n28180), .Z(n28185) );
  NANDN U28861 ( .A(n28183), .B(n28182), .Z(n28184) );
  AND U28862 ( .A(n28185), .B(n28184), .Z(n28467) );
  XNOR U28863 ( .A(n28466), .B(n28467), .Z(n28468) );
  XOR U28864 ( .A(n28469), .B(n28468), .Z(n28206) );
  XNOR U28865 ( .A(n28205), .B(n28206), .Z(n28197) );
  OR U28866 ( .A(n28187), .B(n28186), .Z(n28191) );
  NANDN U28867 ( .A(n28189), .B(n28188), .Z(n28190) );
  AND U28868 ( .A(n28191), .B(n28190), .Z(n28198) );
  XOR U28869 ( .A(n28197), .B(n28198), .Z(n28199) );
  XNOR U28870 ( .A(n28200), .B(n28199), .Z(n28478) );
  XNOR U28871 ( .A(n28478), .B(sreg[190]), .Z(n28480) );
  NAND U28872 ( .A(n28192), .B(sreg[189]), .Z(n28196) );
  OR U28873 ( .A(n28194), .B(n28193), .Z(n28195) );
  AND U28874 ( .A(n28196), .B(n28195), .Z(n28479) );
  XOR U28875 ( .A(n28480), .B(n28479), .Z(c[190]) );
  NAND U28876 ( .A(n28198), .B(n28197), .Z(n28202) );
  NAND U28877 ( .A(n28200), .B(n28199), .Z(n28201) );
  NAND U28878 ( .A(n28202), .B(n28201), .Z(n28486) );
  NANDN U28879 ( .A(n28204), .B(n28203), .Z(n28208) );
  NANDN U28880 ( .A(n28206), .B(n28205), .Z(n28207) );
  NAND U28881 ( .A(n28208), .B(n28207), .Z(n28484) );
  NANDN U28882 ( .A(n28214), .B(n28213), .Z(n28218) );
  NAND U28883 ( .A(n28216), .B(n28215), .Z(n28217) );
  NAND U28884 ( .A(n28218), .B(n28217), .Z(n28726) );
  NANDN U28885 ( .A(n28220), .B(n28219), .Z(n28224) );
  NANDN U28886 ( .A(n28222), .B(n28221), .Z(n28223) );
  NAND U28887 ( .A(n28224), .B(n28223), .Z(n28737) );
  NANDN U28888 ( .A(n28230), .B(n28229), .Z(n28234) );
  NAND U28889 ( .A(n28232), .B(n28231), .Z(n28233) );
  NAND U28890 ( .A(n28234), .B(n28233), .Z(n28683) );
  XOR U28891 ( .A(a[103]), .B(b[25]), .Z(n28581) );
  NANDN U28892 ( .A(n34219), .B(n28581), .Z(n28237) );
  NAND U28893 ( .A(n34217), .B(n28235), .Z(n28236) );
  NAND U28894 ( .A(n28237), .B(n28236), .Z(n28678) );
  XOR U28895 ( .A(a[111]), .B(b[17]), .Z(n28584) );
  NAND U28896 ( .A(n28584), .B(n32543), .Z(n28240) );
  NANDN U28897 ( .A(n28238), .B(n32541), .Z(n28239) );
  NAND U28898 ( .A(n28240), .B(n28239), .Z(n28675) );
  XNOR U28899 ( .A(a[113]), .B(b[15]), .Z(n28578) );
  OR U28900 ( .A(n28578), .B(n32010), .Z(n28243) );
  NANDN U28901 ( .A(n28241), .B(n32011), .Z(n28242) );
  AND U28902 ( .A(n28243), .B(n28242), .Z(n28676) );
  XNOR U28903 ( .A(n28675), .B(n28676), .Z(n28677) );
  XNOR U28904 ( .A(n28678), .B(n28677), .Z(n28681) );
  XNOR U28905 ( .A(b[39]), .B(a[89]), .Z(n28587) );
  NANDN U28906 ( .A(n28587), .B(n36553), .Z(n28246) );
  NANDN U28907 ( .A(n28244), .B(n36643), .Z(n28245) );
  NAND U28908 ( .A(n28246), .B(n28245), .Z(n28657) );
  XNOR U28909 ( .A(b[51]), .B(a[77]), .Z(n28590) );
  NANDN U28910 ( .A(n28590), .B(n37803), .Z(n28249) );
  NANDN U28911 ( .A(n28247), .B(n37802), .Z(n28248) );
  NAND U28912 ( .A(n28249), .B(n28248), .Z(n28654) );
  XNOR U28913 ( .A(b[53]), .B(a[75]), .Z(n28593) );
  NANDN U28914 ( .A(n28593), .B(n37940), .Z(n28252) );
  NANDN U28915 ( .A(n28250), .B(n37941), .Z(n28251) );
  AND U28916 ( .A(n28252), .B(n28251), .Z(n28655) );
  XNOR U28917 ( .A(n28654), .B(n28655), .Z(n28656) );
  XOR U28918 ( .A(n28657), .B(n28656), .Z(n28682) );
  XOR U28919 ( .A(n28681), .B(n28682), .Z(n28684) );
  XNOR U28920 ( .A(n28683), .B(n28684), .Z(n28562) );
  NANDN U28921 ( .A(n28254), .B(n28253), .Z(n28258) );
  NAND U28922 ( .A(n28256), .B(n28255), .Z(n28257) );
  AND U28923 ( .A(n28258), .B(n28257), .Z(n28563) );
  XNOR U28924 ( .A(n28562), .B(n28563), .Z(n28564) );
  XNOR U28925 ( .A(n28565), .B(n28564), .Z(n28735) );
  OR U28926 ( .A(n28260), .B(n28259), .Z(n28264) );
  NANDN U28927 ( .A(n28262), .B(n28261), .Z(n28263) );
  AND U28928 ( .A(n28264), .B(n28263), .Z(n28736) );
  XOR U28929 ( .A(n28735), .B(n28736), .Z(n28738) );
  XOR U28930 ( .A(n28737), .B(n28738), .Z(n28723) );
  NANDN U28931 ( .A(n28266), .B(n28265), .Z(n28270) );
  NANDN U28932 ( .A(n28268), .B(n28267), .Z(n28269) );
  NAND U28933 ( .A(n28270), .B(n28269), .Z(n28730) );
  OR U28934 ( .A(n28272), .B(n28271), .Z(n28276) );
  NANDN U28935 ( .A(n28274), .B(n28273), .Z(n28275) );
  NAND U28936 ( .A(n28276), .B(n28275), .Z(n28614) );
  XNOR U28937 ( .A(a[121]), .B(n31123), .Z(n28517) );
  NAND U28938 ( .A(n28517), .B(n29949), .Z(n28279) );
  NAND U28939 ( .A(n29948), .B(n28277), .Z(n28278) );
  NAND U28940 ( .A(n28279), .B(n28278), .Z(n28599) );
  XNOR U28941 ( .A(b[55]), .B(a[73]), .Z(n28520) );
  NANDN U28942 ( .A(n28520), .B(n38075), .Z(n28282) );
  NANDN U28943 ( .A(n28280), .B(n38073), .Z(n28281) );
  NAND U28944 ( .A(n28282), .B(n28281), .Z(n28596) );
  XNOR U28945 ( .A(b[35]), .B(a[93]), .Z(n28523) );
  NANDN U28946 ( .A(n28523), .B(n35985), .Z(n28285) );
  NANDN U28947 ( .A(n28283), .B(n35986), .Z(n28284) );
  AND U28948 ( .A(n28285), .B(n28284), .Z(n28597) );
  XNOR U28949 ( .A(n28596), .B(n28597), .Z(n28598) );
  XNOR U28950 ( .A(n28599), .B(n28598), .Z(n28612) );
  NANDN U28951 ( .A(n28287), .B(n28286), .Z(n28291) );
  NAND U28952 ( .A(n28289), .B(n28288), .Z(n28290) );
  NAND U28953 ( .A(n28291), .B(n28290), .Z(n28613) );
  XOR U28954 ( .A(n28612), .B(n28613), .Z(n28615) );
  XOR U28955 ( .A(n28614), .B(n28615), .Z(n28729) );
  XNOR U28956 ( .A(n28730), .B(n28729), .Z(n28732) );
  NANDN U28957 ( .A(n28293), .B(n28292), .Z(n28297) );
  NAND U28958 ( .A(n28295), .B(n28294), .Z(n28296) );
  NAND U28959 ( .A(n28297), .B(n28296), .Z(n28632) );
  XNOR U28960 ( .A(b[49]), .B(a[79]), .Z(n28538) );
  OR U28961 ( .A(n28538), .B(n37756), .Z(n28300) );
  NANDN U28962 ( .A(n28298), .B(n37652), .Z(n28299) );
  NAND U28963 ( .A(n28300), .B(n28299), .Z(n28514) );
  NAND U28964 ( .A(n37469), .B(n28301), .Z(n28303) );
  XNOR U28965 ( .A(n978), .B(a[81]), .Z(n28541) );
  NAND U28966 ( .A(n28541), .B(n37471), .Z(n28302) );
  NAND U28967 ( .A(n28303), .B(n28302), .Z(n28511) );
  XOR U28968 ( .A(a[119]), .B(n969), .Z(n28544) );
  NANDN U28969 ( .A(n28544), .B(n30509), .Z(n28306) );
  NANDN U28970 ( .A(n28304), .B(n30846), .Z(n28305) );
  AND U28971 ( .A(n28306), .B(n28305), .Z(n28512) );
  XNOR U28972 ( .A(n28511), .B(n28512), .Z(n28513) );
  XNOR U28973 ( .A(n28514), .B(n28513), .Z(n28630) );
  XNOR U28974 ( .A(a[117]), .B(b[11]), .Z(n28547) );
  OR U28975 ( .A(n28547), .B(n31369), .Z(n28309) );
  NANDN U28976 ( .A(n28307), .B(n31119), .Z(n28308) );
  NAND U28977 ( .A(n28309), .B(n28308), .Z(n28535) );
  XNOR U28978 ( .A(b[43]), .B(a[85]), .Z(n28550) );
  NANDN U28979 ( .A(n28550), .B(n37068), .Z(n28312) );
  NANDN U28980 ( .A(n28310), .B(n37069), .Z(n28311) );
  NAND U28981 ( .A(n28312), .B(n28311), .Z(n28532) );
  XOR U28982 ( .A(b[45]), .B(a[83]), .Z(n28553) );
  NAND U28983 ( .A(n28553), .B(n37261), .Z(n28315) );
  NANDN U28984 ( .A(n28313), .B(n37262), .Z(n28314) );
  AND U28985 ( .A(n28315), .B(n28314), .Z(n28533) );
  XNOR U28986 ( .A(n28532), .B(n28533), .Z(n28534) );
  XOR U28987 ( .A(n28535), .B(n28534), .Z(n28631) );
  XOR U28988 ( .A(n28630), .B(n28631), .Z(n28633) );
  XOR U28989 ( .A(n28632), .B(n28633), .Z(n28731) );
  XOR U28990 ( .A(n28732), .B(n28731), .Z(n28724) );
  XNOR U28991 ( .A(n28723), .B(n28724), .Z(n28725) );
  XNOR U28992 ( .A(n28726), .B(n28725), .Z(n28493) );
  NANDN U28993 ( .A(n28317), .B(n28316), .Z(n28321) );
  NAND U28994 ( .A(n28319), .B(n28318), .Z(n28320) );
  NAND U28995 ( .A(n28321), .B(n28320), .Z(n28742) );
  NANDN U28996 ( .A(n28323), .B(n28322), .Z(n28327) );
  NANDN U28997 ( .A(n28325), .B(n28324), .Z(n28326) );
  AND U28998 ( .A(n28327), .B(n28326), .Z(n28741) );
  NANDN U28999 ( .A(n28329), .B(n28328), .Z(n28333) );
  NANDN U29000 ( .A(n28331), .B(n28330), .Z(n28332) );
  NAND U29001 ( .A(n28333), .B(n28332), .Z(n28744) );
  XOR U29002 ( .A(n28743), .B(n28744), .Z(n28502) );
  NANDN U29003 ( .A(n28335), .B(n28334), .Z(n28339) );
  NAND U29004 ( .A(n28337), .B(n28336), .Z(n28338) );
  NAND U29005 ( .A(n28339), .B(n28338), .Z(n28499) );
  NANDN U29006 ( .A(n28341), .B(n28340), .Z(n28345) );
  OR U29007 ( .A(n28343), .B(n28342), .Z(n28344) );
  NAND U29008 ( .A(n28345), .B(n28344), .Z(n28611) );
  NANDN U29009 ( .A(n28347), .B(n28346), .Z(n28351) );
  NAND U29010 ( .A(n28349), .B(n28348), .Z(n28350) );
  NAND U29011 ( .A(n28351), .B(n28350), .Z(n28508) );
  XNOR U29012 ( .A(b[31]), .B(a[97]), .Z(n28660) );
  NANDN U29013 ( .A(n28660), .B(n35313), .Z(n28354) );
  NANDN U29014 ( .A(n28352), .B(n35311), .Z(n28353) );
  NAND U29015 ( .A(n28354), .B(n28353), .Z(n28529) );
  XOR U29016 ( .A(b[61]), .B(n29372), .Z(n28663) );
  OR U29017 ( .A(n28663), .B(n38371), .Z(n28357) );
  NANDN U29018 ( .A(n28355), .B(n38369), .Z(n28356) );
  NAND U29019 ( .A(n28357), .B(n28356), .Z(n28526) );
  NANDN U29020 ( .A(n985), .B(a[63]), .Z(n28527) );
  XNOR U29021 ( .A(n28526), .B(n28527), .Z(n28528) );
  XNOR U29022 ( .A(n28529), .B(n28528), .Z(n28505) );
  NAND U29023 ( .A(n33283), .B(n28358), .Z(n28360) );
  XNOR U29024 ( .A(a[109]), .B(n33020), .Z(n28666) );
  NANDN U29025 ( .A(n33021), .B(n28666), .Z(n28359) );
  NAND U29026 ( .A(n28360), .B(n28359), .Z(n28696) );
  XOR U29027 ( .A(a[107]), .B(b[21]), .Z(n28669) );
  NANDN U29028 ( .A(n33634), .B(n28669), .Z(n28363) );
  NANDN U29029 ( .A(n28361), .B(n33464), .Z(n28362) );
  NAND U29030 ( .A(n28363), .B(n28362), .Z(n28693) );
  NAND U29031 ( .A(n34044), .B(n28364), .Z(n28366) );
  XNOR U29032 ( .A(a[105]), .B(n34510), .Z(n28672) );
  NANDN U29033 ( .A(n33867), .B(n28672), .Z(n28365) );
  AND U29034 ( .A(n28366), .B(n28365), .Z(n28694) );
  XNOR U29035 ( .A(n28693), .B(n28694), .Z(n28695) );
  XOR U29036 ( .A(n28696), .B(n28695), .Z(n28506) );
  XNOR U29037 ( .A(n28505), .B(n28506), .Z(n28507) );
  XNOR U29038 ( .A(n28508), .B(n28507), .Z(n28608) );
  XNOR U29039 ( .A(b[37]), .B(a[91]), .Z(n28636) );
  NANDN U29040 ( .A(n28636), .B(n36311), .Z(n28369) );
  NANDN U29041 ( .A(n28367), .B(n36309), .Z(n28368) );
  NAND U29042 ( .A(n28369), .B(n28368), .Z(n28690) );
  XNOR U29043 ( .A(a[123]), .B(b[5]), .Z(n28639) );
  OR U29044 ( .A(n28639), .B(n29363), .Z(n28372) );
  NANDN U29045 ( .A(n28370), .B(n29864), .Z(n28371) );
  NAND U29046 ( .A(n28372), .B(n28371), .Z(n28687) );
  XNOR U29047 ( .A(a[125]), .B(n967), .Z(n28642) );
  NAND U29048 ( .A(n28642), .B(n28939), .Z(n28375) );
  NAND U29049 ( .A(n28938), .B(n28373), .Z(n28374) );
  AND U29050 ( .A(n28375), .B(n28374), .Z(n28688) );
  XNOR U29051 ( .A(n28687), .B(n28688), .Z(n28689) );
  XNOR U29052 ( .A(n28690), .B(n28689), .Z(n28626) );
  XNOR U29053 ( .A(a[115]), .B(b[13]), .Z(n28645) );
  OR U29054 ( .A(n28645), .B(n31550), .Z(n28378) );
  NANDN U29055 ( .A(n28376), .B(n31874), .Z(n28377) );
  NAND U29056 ( .A(n28378), .B(n28377), .Z(n28575) );
  NAND U29057 ( .A(n34848), .B(n28379), .Z(n28381) );
  XNOR U29058 ( .A(a[101]), .B(n35375), .Z(n28648) );
  NAND U29059 ( .A(n34618), .B(n28648), .Z(n28380) );
  NAND U29060 ( .A(n28381), .B(n28380), .Z(n28572) );
  NAND U29061 ( .A(n35188), .B(n28382), .Z(n28384) );
  XNOR U29062 ( .A(a[99]), .B(n35540), .Z(n28651) );
  NANDN U29063 ( .A(n34968), .B(n28651), .Z(n28383) );
  AND U29064 ( .A(n28384), .B(n28383), .Z(n28573) );
  XNOR U29065 ( .A(n28572), .B(n28573), .Z(n28574) );
  XNOR U29066 ( .A(n28575), .B(n28574), .Z(n28624) );
  NANDN U29067 ( .A(n28386), .B(n28385), .Z(n28390) );
  NAND U29068 ( .A(n28388), .B(n28387), .Z(n28389) );
  NAND U29069 ( .A(n28390), .B(n28389), .Z(n28625) );
  XOR U29070 ( .A(n28624), .B(n28625), .Z(n28627) );
  XNOR U29071 ( .A(n28626), .B(n28627), .Z(n28609) );
  XOR U29072 ( .A(n28608), .B(n28609), .Z(n28610) );
  XNOR U29073 ( .A(n28611), .B(n28610), .Z(n28559) );
  NANDN U29074 ( .A(n28392), .B(n28391), .Z(n28396) );
  OR U29075 ( .A(n28394), .B(n28393), .Z(n28395) );
  NAND U29076 ( .A(n28396), .B(n28395), .Z(n28556) );
  XOR U29077 ( .A(b[33]), .B(n35628), .Z(n28705) );
  NANDN U29078 ( .A(n28705), .B(n35620), .Z(n28399) );
  NANDN U29079 ( .A(n28397), .B(n35621), .Z(n28398) );
  NAND U29080 ( .A(n28399), .B(n28398), .Z(n28571) );
  NANDN U29081 ( .A(n966), .B(a[127]), .Z(n28400) );
  XOR U29082 ( .A(n29232), .B(n28400), .Z(n28402) );
  NANDN U29083 ( .A(n987), .B(n966), .Z(n28401) );
  AND U29084 ( .A(n28402), .B(n28401), .Z(n28568) );
  XOR U29085 ( .A(b[63]), .B(n28403), .Z(n28702) );
  NANDN U29086 ( .A(n28702), .B(n38422), .Z(n28406) );
  NANDN U29087 ( .A(n28404), .B(n38423), .Z(n28405) );
  AND U29088 ( .A(n28406), .B(n28405), .Z(n28569) );
  XNOR U29089 ( .A(n28568), .B(n28569), .Z(n28570) );
  XNOR U29090 ( .A(n28571), .B(n28570), .Z(n28602) );
  XOR U29091 ( .A(b[57]), .B(n30543), .Z(n28708) );
  OR U29092 ( .A(n28708), .B(n965), .Z(n28409) );
  NANDN U29093 ( .A(n28407), .B(n38194), .Z(n28408) );
  NAND U29094 ( .A(n28409), .B(n28408), .Z(n28720) );
  NAND U29095 ( .A(n38326), .B(n28410), .Z(n28412) );
  XNOR U29096 ( .A(n38400), .B(a[69]), .Z(n28711) );
  NANDN U29097 ( .A(n38273), .B(n28711), .Z(n28411) );
  NAND U29098 ( .A(n28412), .B(n28411), .Z(n28717) );
  XOR U29099 ( .A(b[41]), .B(a[87]), .Z(n28714) );
  NANDN U29100 ( .A(n36905), .B(n28714), .Z(n28415) );
  NANDN U29101 ( .A(n28413), .B(n36807), .Z(n28414) );
  AND U29102 ( .A(n28415), .B(n28414), .Z(n28718) );
  XNOR U29103 ( .A(n28717), .B(n28718), .Z(n28719) );
  XOR U29104 ( .A(n28720), .B(n28719), .Z(n28603) );
  XNOR U29105 ( .A(n28602), .B(n28603), .Z(n28604) );
  NANDN U29106 ( .A(n28417), .B(n28416), .Z(n28421) );
  NAND U29107 ( .A(n28419), .B(n28418), .Z(n28420) );
  NAND U29108 ( .A(n28421), .B(n28420), .Z(n28605) );
  XOR U29109 ( .A(n28604), .B(n28605), .Z(n28621) );
  NANDN U29110 ( .A(n28423), .B(n28422), .Z(n28427) );
  NAND U29111 ( .A(n28425), .B(n28424), .Z(n28426) );
  NAND U29112 ( .A(n28427), .B(n28426), .Z(n28618) );
  NANDN U29113 ( .A(n28429), .B(n28428), .Z(n28433) );
  NAND U29114 ( .A(n28431), .B(n28430), .Z(n28432) );
  AND U29115 ( .A(n28433), .B(n28432), .Z(n28619) );
  XNOR U29116 ( .A(n28618), .B(n28619), .Z(n28620) );
  XOR U29117 ( .A(n28621), .B(n28620), .Z(n28557) );
  XNOR U29118 ( .A(n28556), .B(n28557), .Z(n28558) );
  XOR U29119 ( .A(n28559), .B(n28558), .Z(n28500) );
  XNOR U29120 ( .A(n28499), .B(n28500), .Z(n28501) );
  XOR U29121 ( .A(n28502), .B(n28501), .Z(n28494) );
  XOR U29122 ( .A(n28493), .B(n28494), .Z(n28496) );
  XNOR U29123 ( .A(n28495), .B(n28496), .Z(n28755) );
  NANDN U29124 ( .A(n28435), .B(n28434), .Z(n28439) );
  NANDN U29125 ( .A(n28437), .B(n28436), .Z(n28438) );
  AND U29126 ( .A(n28439), .B(n28438), .Z(n28753) );
  NANDN U29127 ( .A(n28445), .B(n28444), .Z(n28449) );
  NANDN U29128 ( .A(n28447), .B(n28446), .Z(n28448) );
  NAND U29129 ( .A(n28449), .B(n28448), .Z(n28487) );
  XNOR U29130 ( .A(n28487), .B(n28488), .Z(n28489) );
  XNOR U29131 ( .A(n28490), .B(n28489), .Z(n28754) );
  XOR U29132 ( .A(n28755), .B(n28756), .Z(n28750) );
  NANDN U29133 ( .A(n28455), .B(n28454), .Z(n28459) );
  NAND U29134 ( .A(n28457), .B(n28456), .Z(n28458) );
  NAND U29135 ( .A(n28459), .B(n28458), .Z(n28747) );
  NAND U29136 ( .A(n28461), .B(n28460), .Z(n28465) );
  NAND U29137 ( .A(n28463), .B(n28462), .Z(n28464) );
  NAND U29138 ( .A(n28465), .B(n28464), .Z(n28748) );
  XNOR U29139 ( .A(n28747), .B(n28748), .Z(n28749) );
  XOR U29140 ( .A(n28750), .B(n28749), .Z(n28762) );
  NANDN U29141 ( .A(n28467), .B(n28466), .Z(n28471) );
  NANDN U29142 ( .A(n28469), .B(n28468), .Z(n28470) );
  NAND U29143 ( .A(n28471), .B(n28470), .Z(n28759) );
  OR U29144 ( .A(n28473), .B(n28472), .Z(n28477) );
  OR U29145 ( .A(n28475), .B(n28474), .Z(n28476) );
  AND U29146 ( .A(n28477), .B(n28476), .Z(n28760) );
  XNOR U29147 ( .A(n28759), .B(n28760), .Z(n28761) );
  XNOR U29148 ( .A(n28762), .B(n28761), .Z(n28483) );
  XOR U29149 ( .A(n28484), .B(n28483), .Z(n28485) );
  XNOR U29150 ( .A(n28486), .B(n28485), .Z(n28765) );
  XNOR U29151 ( .A(n28765), .B(sreg[191]), .Z(n28767) );
  NAND U29152 ( .A(n28478), .B(sreg[190]), .Z(n28482) );
  OR U29153 ( .A(n28480), .B(n28479), .Z(n28481) );
  AND U29154 ( .A(n28482), .B(n28481), .Z(n28766) );
  XOR U29155 ( .A(n28767), .B(n28766), .Z(c[191]) );
  NANDN U29156 ( .A(n28488), .B(n28487), .Z(n28492) );
  NAND U29157 ( .A(n28490), .B(n28489), .Z(n28491) );
  NAND U29158 ( .A(n28492), .B(n28491), .Z(n29042) );
  NANDN U29159 ( .A(n28494), .B(n28493), .Z(n28498) );
  OR U29160 ( .A(n28496), .B(n28495), .Z(n28497) );
  NAND U29161 ( .A(n28498), .B(n28497), .Z(n29043) );
  XNOR U29162 ( .A(n29042), .B(n29043), .Z(n29044) );
  NANDN U29163 ( .A(n28500), .B(n28499), .Z(n28504) );
  NAND U29164 ( .A(n28502), .B(n28501), .Z(n28503) );
  NAND U29165 ( .A(n28504), .B(n28503), .Z(n29027) );
  NANDN U29166 ( .A(n28506), .B(n28505), .Z(n28510) );
  NANDN U29167 ( .A(n28508), .B(n28507), .Z(n28509) );
  NAND U29168 ( .A(n28510), .B(n28509), .Z(n29013) );
  NANDN U29169 ( .A(n28512), .B(n28511), .Z(n28516) );
  NAND U29170 ( .A(n28514), .B(n28513), .Z(n28515) );
  NAND U29171 ( .A(n28516), .B(n28515), .Z(n28903) );
  XOR U29172 ( .A(n38251), .B(n31123), .Z(n28981) );
  NAND U29173 ( .A(n28981), .B(n29949), .Z(n28519) );
  NAND U29174 ( .A(n29948), .B(n28517), .Z(n28518) );
  NAND U29175 ( .A(n28519), .B(n28518), .Z(n28809) );
  XOR U29176 ( .A(b[55]), .B(n31372), .Z(n28854) );
  NANDN U29177 ( .A(n28854), .B(n38075), .Z(n28522) );
  NANDN U29178 ( .A(n28520), .B(n38073), .Z(n28521) );
  NAND U29179 ( .A(n28522), .B(n28521), .Z(n28806) );
  XNOR U29180 ( .A(b[35]), .B(a[94]), .Z(n28848) );
  NANDN U29181 ( .A(n28848), .B(n35985), .Z(n28525) );
  NANDN U29182 ( .A(n28523), .B(n35986), .Z(n28524) );
  AND U29183 ( .A(n28525), .B(n28524), .Z(n28807) );
  XNOR U29184 ( .A(n28806), .B(n28807), .Z(n28808) );
  XNOR U29185 ( .A(n28809), .B(n28808), .Z(n28901) );
  NANDN U29186 ( .A(n28527), .B(n28526), .Z(n28531) );
  NAND U29187 ( .A(n28529), .B(n28528), .Z(n28530) );
  NAND U29188 ( .A(n28531), .B(n28530), .Z(n28902) );
  XOR U29189 ( .A(n28901), .B(n28902), .Z(n28904) );
  XOR U29190 ( .A(n28903), .B(n28904), .Z(n29012) );
  XNOR U29191 ( .A(n29013), .B(n29012), .Z(n29015) );
  NANDN U29192 ( .A(n28533), .B(n28532), .Z(n28537) );
  NAND U29193 ( .A(n28535), .B(n28534), .Z(n28536) );
  NAND U29194 ( .A(n28537), .B(n28536), .Z(n28959) );
  XOR U29195 ( .A(b[49]), .B(n32814), .Z(n28872) );
  OR U29196 ( .A(n28872), .B(n37756), .Z(n28540) );
  NANDN U29197 ( .A(n28538), .B(n37652), .Z(n28539) );
  NAND U29198 ( .A(n28540), .B(n28539), .Z(n28845) );
  NAND U29199 ( .A(n37469), .B(n28541), .Z(n28543) );
  XOR U29200 ( .A(n978), .B(n32815), .Z(n28875) );
  NAND U29201 ( .A(n28875), .B(n37471), .Z(n28542) );
  NAND U29202 ( .A(n28543), .B(n28542), .Z(n28842) );
  XOR U29203 ( .A(a[120]), .B(n969), .Z(n28851) );
  NANDN U29204 ( .A(n28851), .B(n30509), .Z(n28546) );
  NANDN U29205 ( .A(n28544), .B(n30846), .Z(n28545) );
  AND U29206 ( .A(n28546), .B(n28545), .Z(n28843) );
  XNOR U29207 ( .A(n28842), .B(n28843), .Z(n28844) );
  XNOR U29208 ( .A(n28845), .B(n28844), .Z(n28957) );
  XOR U29209 ( .A(a[118]), .B(n970), .Z(n28878) );
  OR U29210 ( .A(n28878), .B(n31369), .Z(n28549) );
  NANDN U29211 ( .A(n28547), .B(n31119), .Z(n28548) );
  NAND U29212 ( .A(n28549), .B(n28548), .Z(n28884) );
  XOR U29213 ( .A(b[43]), .B(n33628), .Z(n28866) );
  NANDN U29214 ( .A(n28866), .B(n37068), .Z(n28552) );
  NANDN U29215 ( .A(n28550), .B(n37069), .Z(n28551) );
  NAND U29216 ( .A(n28552), .B(n28551), .Z(n28881) );
  XNOR U29217 ( .A(b[45]), .B(a[84]), .Z(n28869) );
  NANDN U29218 ( .A(n28869), .B(n37261), .Z(n28555) );
  NAND U29219 ( .A(n28553), .B(n37262), .Z(n28554) );
  AND U29220 ( .A(n28555), .B(n28554), .Z(n28882) );
  XNOR U29221 ( .A(n28881), .B(n28882), .Z(n28883) );
  XOR U29222 ( .A(n28884), .B(n28883), .Z(n28958) );
  XOR U29223 ( .A(n28957), .B(n28958), .Z(n28960) );
  XOR U29224 ( .A(n28959), .B(n28960), .Z(n29014) );
  XOR U29225 ( .A(n29015), .B(n29014), .Z(n28781) );
  NANDN U29226 ( .A(n28557), .B(n28556), .Z(n28561) );
  NANDN U29227 ( .A(n28559), .B(n28558), .Z(n28560) );
  AND U29228 ( .A(n28561), .B(n28560), .Z(n28779) );
  NANDN U29229 ( .A(n28563), .B(n28562), .Z(n28567) );
  NAND U29230 ( .A(n28565), .B(n28564), .Z(n28566) );
  NAND U29231 ( .A(n28567), .B(n28566), .Z(n29008) );
  NANDN U29232 ( .A(n28573), .B(n28572), .Z(n28577) );
  NAND U29233 ( .A(n28575), .B(n28574), .Z(n28576) );
  NAND U29234 ( .A(n28577), .B(n28576), .Z(n28953) );
  XOR U29235 ( .A(a[114]), .B(n972), .Z(n28969) );
  OR U29236 ( .A(n28969), .B(n32010), .Z(n28580) );
  NANDN U29237 ( .A(n28578), .B(n32011), .Z(n28579) );
  NAND U29238 ( .A(n28580), .B(n28579), .Z(n28990) );
  XNOR U29239 ( .A(n36647), .B(b[25]), .Z(n28999) );
  NANDN U29240 ( .A(n34219), .B(n28999), .Z(n28583) );
  NAND U29241 ( .A(n34217), .B(n28581), .Z(n28582) );
  NAND U29242 ( .A(n28583), .B(n28582), .Z(n28987) );
  XNOR U29243 ( .A(a[112]), .B(b[17]), .Z(n28818) );
  NANDN U29244 ( .A(n28818), .B(n32543), .Z(n28586) );
  NAND U29245 ( .A(n28584), .B(n32541), .Z(n28585) );
  AND U29246 ( .A(n28586), .B(n28585), .Z(n28988) );
  XNOR U29247 ( .A(n28987), .B(n28988), .Z(n28989) );
  XNOR U29248 ( .A(n28990), .B(n28989), .Z(n28951) );
  XOR U29249 ( .A(n976), .B(n34851), .Z(n28833) );
  NAND U29250 ( .A(n28833), .B(n36553), .Z(n28589) );
  NANDN U29251 ( .A(n28587), .B(n36643), .Z(n28588) );
  NAND U29252 ( .A(n28589), .B(n28588), .Z(n28966) );
  XOR U29253 ( .A(n980), .B(n31870), .Z(n28827) );
  NAND U29254 ( .A(n28827), .B(n37803), .Z(n28592) );
  NANDN U29255 ( .A(n28590), .B(n37802), .Z(n28591) );
  NAND U29256 ( .A(n28592), .B(n28591), .Z(n28963) );
  XOR U29257 ( .A(n981), .B(n31363), .Z(n28830) );
  NAND U29258 ( .A(n28830), .B(n37940), .Z(n28595) );
  NANDN U29259 ( .A(n28593), .B(n37941), .Z(n28594) );
  AND U29260 ( .A(n28595), .B(n28594), .Z(n28964) );
  XNOR U29261 ( .A(n28963), .B(n28964), .Z(n28965) );
  XOR U29262 ( .A(n28966), .B(n28965), .Z(n28952) );
  XOR U29263 ( .A(n28951), .B(n28952), .Z(n28954) );
  XNOR U29264 ( .A(n28953), .B(n28954), .Z(n28794) );
  NANDN U29265 ( .A(n28597), .B(n28596), .Z(n28601) );
  NAND U29266 ( .A(n28599), .B(n28598), .Z(n28600) );
  AND U29267 ( .A(n28601), .B(n28600), .Z(n28795) );
  XNOR U29268 ( .A(n28794), .B(n28795), .Z(n28796) );
  XNOR U29269 ( .A(n28797), .B(n28796), .Z(n29006) );
  NANDN U29270 ( .A(n28603), .B(n28602), .Z(n28607) );
  NANDN U29271 ( .A(n28605), .B(n28604), .Z(n28606) );
  AND U29272 ( .A(n28607), .B(n28606), .Z(n29007) );
  XOR U29273 ( .A(n29006), .B(n29007), .Z(n29009) );
  XNOR U29274 ( .A(n29008), .B(n29009), .Z(n28778) );
  XOR U29275 ( .A(n28781), .B(n28780), .Z(n29025) );
  NANDN U29276 ( .A(n28613), .B(n28612), .Z(n28617) );
  OR U29277 ( .A(n28615), .B(n28614), .Z(n28616) );
  AND U29278 ( .A(n28617), .B(n28616), .Z(n29018) );
  NANDN U29279 ( .A(n28619), .B(n28618), .Z(n28623) );
  NAND U29280 ( .A(n28621), .B(n28620), .Z(n28622) );
  NAND U29281 ( .A(n28623), .B(n28622), .Z(n29019) );
  NANDN U29282 ( .A(n28625), .B(n28624), .Z(n28629) );
  NANDN U29283 ( .A(n28627), .B(n28626), .Z(n28628) );
  NAND U29284 ( .A(n28629), .B(n28628), .Z(n29021) );
  XNOR U29285 ( .A(n29020), .B(n29021), .Z(n28785) );
  XNOR U29286 ( .A(n28784), .B(n28785), .Z(n28786) );
  NANDN U29287 ( .A(n28631), .B(n28630), .Z(n28635) );
  OR U29288 ( .A(n28633), .B(n28632), .Z(n28634) );
  NAND U29289 ( .A(n28635), .B(n28634), .Z(n28910) );
  XOR U29290 ( .A(b[37]), .B(n34852), .Z(n28978) );
  NANDN U29291 ( .A(n28978), .B(n36311), .Z(n28638) );
  NANDN U29292 ( .A(n28636), .B(n36309), .Z(n28637) );
  NAND U29293 ( .A(n28638), .B(n28637), .Z(n28916) );
  XOR U29294 ( .A(a[124]), .B(n968), .Z(n28984) );
  OR U29295 ( .A(n28984), .B(n29363), .Z(n28641) );
  NANDN U29296 ( .A(n28639), .B(n29864), .Z(n28640) );
  NAND U29297 ( .A(n28641), .B(n28640), .Z(n28913) );
  XOR U29298 ( .A(n987), .B(n967), .Z(n28937) );
  NAND U29299 ( .A(n28937), .B(n28939), .Z(n28644) );
  NAND U29300 ( .A(n28938), .B(n28642), .Z(n28643) );
  AND U29301 ( .A(n28644), .B(n28643), .Z(n28914) );
  XNOR U29302 ( .A(n28913), .B(n28914), .Z(n28915) );
  XNOR U29303 ( .A(n28916), .B(n28915), .Z(n28894) );
  XOR U29304 ( .A(a[116]), .B(n971), .Z(n28863) );
  OR U29305 ( .A(n28863), .B(n31550), .Z(n28647) );
  NANDN U29306 ( .A(n28645), .B(n31874), .Z(n28646) );
  NAND U29307 ( .A(n28647), .B(n28646), .Z(n28815) );
  NAND U29308 ( .A(n34848), .B(n28648), .Z(n28650) );
  XOR U29309 ( .A(a[102]), .B(n35375), .Z(n28821) );
  NANDN U29310 ( .A(n28821), .B(n34618), .Z(n28649) );
  NAND U29311 ( .A(n28650), .B(n28649), .Z(n28812) );
  NAND U29312 ( .A(n35188), .B(n28651), .Z(n28653) );
  XOR U29313 ( .A(n36100), .B(n35540), .Z(n28972) );
  NANDN U29314 ( .A(n34968), .B(n28972), .Z(n28652) );
  AND U29315 ( .A(n28653), .B(n28652), .Z(n28813) );
  XNOR U29316 ( .A(n28812), .B(n28813), .Z(n28814) );
  XNOR U29317 ( .A(n28815), .B(n28814), .Z(n28891) );
  NANDN U29318 ( .A(n28655), .B(n28654), .Z(n28659) );
  NAND U29319 ( .A(n28657), .B(n28656), .Z(n28658) );
  NAND U29320 ( .A(n28659), .B(n28658), .Z(n28892) );
  XNOR U29321 ( .A(n28891), .B(n28892), .Z(n28893) );
  XOR U29322 ( .A(n28894), .B(n28893), .Z(n28907) );
  XOR U29323 ( .A(a[98]), .B(n973), .Z(n28975) );
  NANDN U29324 ( .A(n28975), .B(n35313), .Z(n28662) );
  NANDN U29325 ( .A(n28660), .B(n35311), .Z(n28661) );
  NAND U29326 ( .A(n28662), .B(n28661), .Z(n28860) );
  XOR U29327 ( .A(b[61]), .B(n29868), .Z(n29002) );
  OR U29328 ( .A(n29002), .B(n38371), .Z(n28665) );
  NANDN U29329 ( .A(n28663), .B(n38369), .Z(n28664) );
  NAND U29330 ( .A(n28665), .B(n28664), .Z(n28857) );
  NANDN U29331 ( .A(n985), .B(a[64]), .Z(n28858) );
  XNOR U29332 ( .A(n28857), .B(n28858), .Z(n28859) );
  XNOR U29333 ( .A(n28860), .B(n28859), .Z(n28887) );
  NAND U29334 ( .A(n33283), .B(n28666), .Z(n28668) );
  XOR U29335 ( .A(a[110]), .B(n33020), .Z(n28824) );
  OR U29336 ( .A(n28824), .B(n33021), .Z(n28667) );
  NAND U29337 ( .A(n28668), .B(n28667), .Z(n28922) );
  XNOR U29338 ( .A(a[108]), .B(b[21]), .Z(n28993) );
  OR U29339 ( .A(n28993), .B(n33634), .Z(n28671) );
  NAND U29340 ( .A(n28669), .B(n33464), .Z(n28670) );
  NAND U29341 ( .A(n28671), .B(n28670), .Z(n28919) );
  NAND U29342 ( .A(n34044), .B(n28672), .Z(n28674) );
  XOR U29343 ( .A(n36909), .B(n34510), .Z(n28996) );
  NANDN U29344 ( .A(n33867), .B(n28996), .Z(n28673) );
  AND U29345 ( .A(n28674), .B(n28673), .Z(n28920) );
  XNOR U29346 ( .A(n28919), .B(n28920), .Z(n28921) );
  XOR U29347 ( .A(n28922), .B(n28921), .Z(n28888) );
  XNOR U29348 ( .A(n28887), .B(n28888), .Z(n28889) );
  NANDN U29349 ( .A(n28676), .B(n28675), .Z(n28680) );
  NAND U29350 ( .A(n28678), .B(n28677), .Z(n28679) );
  AND U29351 ( .A(n28680), .B(n28679), .Z(n28890) );
  XNOR U29352 ( .A(n28889), .B(n28890), .Z(n28908) );
  XNOR U29353 ( .A(n28907), .B(n28908), .Z(n28909) );
  XNOR U29354 ( .A(n28910), .B(n28909), .Z(n28792) );
  NANDN U29355 ( .A(n28682), .B(n28681), .Z(n28686) );
  OR U29356 ( .A(n28684), .B(n28683), .Z(n28685) );
  NAND U29357 ( .A(n28686), .B(n28685), .Z(n28791) );
  NANDN U29358 ( .A(n28688), .B(n28687), .Z(n28692) );
  NAND U29359 ( .A(n28690), .B(n28689), .Z(n28691) );
  NAND U29360 ( .A(n28692), .B(n28691), .Z(n28898) );
  NANDN U29361 ( .A(n28694), .B(n28693), .Z(n28698) );
  NAND U29362 ( .A(n28696), .B(n28695), .Z(n28697) );
  AND U29363 ( .A(n28698), .B(n28697), .Z(n28839) );
  NANDN U29364 ( .A(n966), .B(b[1]), .Z(n28700) );
  IV U29365 ( .A(a[127]), .Z(n38463) );
  NANDN U29366 ( .A(n29232), .B(n38463), .Z(n28699) );
  NAND U29367 ( .A(n28700), .B(n28699), .Z(n28803) );
  XOR U29368 ( .A(b[63]), .B(n28701), .Z(n28942) );
  NANDN U29369 ( .A(n28942), .B(n38422), .Z(n28704) );
  NANDN U29370 ( .A(n28702), .B(n38423), .Z(n28703) );
  NAND U29371 ( .A(n28704), .B(n28703), .Z(n28800) );
  XOR U29372 ( .A(b[33]), .B(n35545), .Z(n28934) );
  NANDN U29373 ( .A(n28934), .B(n35620), .Z(n28707) );
  NANDN U29374 ( .A(n28705), .B(n35621), .Z(n28706) );
  AND U29375 ( .A(n28707), .B(n28706), .Z(n28801) );
  XNOR U29376 ( .A(n28800), .B(n28801), .Z(n28802) );
  XNOR U29377 ( .A(n28803), .B(n28802), .Z(n28837) );
  XOR U29378 ( .A(b[57]), .B(n30210), .Z(n28925) );
  OR U29379 ( .A(n28925), .B(n965), .Z(n28710) );
  NANDN U29380 ( .A(n28708), .B(n38194), .Z(n28709) );
  NAND U29381 ( .A(n28710), .B(n28709), .Z(n28948) );
  NAND U29382 ( .A(n38326), .B(n28711), .Z(n28713) );
  XOR U29383 ( .A(n38400), .B(n30379), .Z(n28928) );
  NANDN U29384 ( .A(n38273), .B(n28928), .Z(n28712) );
  NAND U29385 ( .A(n28713), .B(n28712), .Z(n28945) );
  XNOR U29386 ( .A(b[41]), .B(a[88]), .Z(n28931) );
  OR U29387 ( .A(n28931), .B(n36905), .Z(n28716) );
  NAND U29388 ( .A(n28714), .B(n36807), .Z(n28715) );
  AND U29389 ( .A(n28716), .B(n28715), .Z(n28946) );
  XNOR U29390 ( .A(n28945), .B(n28946), .Z(n28947) );
  XNOR U29391 ( .A(n28948), .B(n28947), .Z(n28836) );
  XOR U29392 ( .A(n28837), .B(n28836), .Z(n28838) );
  XNOR U29393 ( .A(n28839), .B(n28838), .Z(n28896) );
  NANDN U29394 ( .A(n28718), .B(n28717), .Z(n28722) );
  NAND U29395 ( .A(n28720), .B(n28719), .Z(n28721) );
  NAND U29396 ( .A(n28722), .B(n28721), .Z(n28895) );
  XOR U29397 ( .A(n28896), .B(n28895), .Z(n28897) );
  XNOR U29398 ( .A(n28898), .B(n28897), .Z(n28790) );
  XNOR U29399 ( .A(n28791), .B(n28790), .Z(n28793) );
  XOR U29400 ( .A(n28792), .B(n28793), .Z(n28787) );
  XOR U29401 ( .A(n28786), .B(n28787), .Z(n29024) );
  XOR U29402 ( .A(n29025), .B(n29024), .Z(n29026) );
  XOR U29403 ( .A(n29027), .B(n29026), .Z(n29039) );
  NANDN U29404 ( .A(n28724), .B(n28723), .Z(n28728) );
  NAND U29405 ( .A(n28726), .B(n28725), .Z(n28727) );
  NAND U29406 ( .A(n28728), .B(n28727), .Z(n29036) );
  NAND U29407 ( .A(n28730), .B(n28729), .Z(n28734) );
  NANDN U29408 ( .A(n28732), .B(n28731), .Z(n28733) );
  NAND U29409 ( .A(n28734), .B(n28733), .Z(n29033) );
  NANDN U29410 ( .A(n28736), .B(n28735), .Z(n28740) );
  OR U29411 ( .A(n28738), .B(n28737), .Z(n28739) );
  NAND U29412 ( .A(n28740), .B(n28739), .Z(n29030) );
  OR U29413 ( .A(n28742), .B(n28741), .Z(n28746) );
  NANDN U29414 ( .A(n28744), .B(n28743), .Z(n28745) );
  NAND U29415 ( .A(n28746), .B(n28745), .Z(n29031) );
  XNOR U29416 ( .A(n29030), .B(n29031), .Z(n29032) );
  XNOR U29417 ( .A(n29033), .B(n29032), .Z(n29037) );
  XNOR U29418 ( .A(n29036), .B(n29037), .Z(n29038) );
  XNOR U29419 ( .A(n29039), .B(n29038), .Z(n29045) );
  XOR U29420 ( .A(n29044), .B(n29045), .Z(n29051) );
  NANDN U29421 ( .A(n28748), .B(n28747), .Z(n28752) );
  NAND U29422 ( .A(n28750), .B(n28749), .Z(n28751) );
  NAND U29423 ( .A(n28752), .B(n28751), .Z(n29048) );
  OR U29424 ( .A(n28754), .B(n28753), .Z(n28758) );
  NANDN U29425 ( .A(n28756), .B(n28755), .Z(n28757) );
  NAND U29426 ( .A(n28758), .B(n28757), .Z(n29049) );
  XNOR U29427 ( .A(n29048), .B(n29049), .Z(n29050) );
  XNOR U29428 ( .A(n29051), .B(n29050), .Z(n28772) );
  NANDN U29429 ( .A(n28760), .B(n28759), .Z(n28764) );
  NANDN U29430 ( .A(n28762), .B(n28761), .Z(n28763) );
  AND U29431 ( .A(n28764), .B(n28763), .Z(n28773) );
  XNOR U29432 ( .A(n28772), .B(n28773), .Z(n28774) );
  XOR U29433 ( .A(n28775), .B(n28774), .Z(n28771) );
  NAND U29434 ( .A(n28765), .B(sreg[191]), .Z(n28769) );
  OR U29435 ( .A(n28767), .B(n28766), .Z(n28768) );
  AND U29436 ( .A(n28769), .B(n28768), .Z(n28770) );
  XOR U29437 ( .A(n28771), .B(n28770), .Z(c[192]) );
  OR U29438 ( .A(n28771), .B(n28770), .Z(n29335) );
  NANDN U29439 ( .A(n28773), .B(n28772), .Z(n28777) );
  NAND U29440 ( .A(n28775), .B(n28774), .Z(n28776) );
  NAND U29441 ( .A(n28777), .B(n28776), .Z(n29330) );
  OR U29442 ( .A(n28779), .B(n28778), .Z(n28783) );
  OR U29443 ( .A(n28781), .B(n28780), .Z(n28782) );
  AND U29444 ( .A(n28783), .B(n28782), .Z(n29055) );
  NANDN U29445 ( .A(n28785), .B(n28784), .Z(n28789) );
  NAND U29446 ( .A(n28787), .B(n28786), .Z(n28788) );
  NAND U29447 ( .A(n28789), .B(n28788), .Z(n29309) );
  NANDN U29448 ( .A(n28795), .B(n28794), .Z(n28799) );
  NAND U29449 ( .A(n28797), .B(n28796), .Z(n28798) );
  NAND U29450 ( .A(n28799), .B(n28798), .Z(n29300) );
  NANDN U29451 ( .A(n28801), .B(n28800), .Z(n28805) );
  NAND U29452 ( .A(n28803), .B(n28802), .Z(n28804) );
  NAND U29453 ( .A(n28805), .B(n28804), .Z(n29252) );
  NANDN U29454 ( .A(n28807), .B(n28806), .Z(n28811) );
  NAND U29455 ( .A(n28809), .B(n28808), .Z(n28810) );
  NAND U29456 ( .A(n28811), .B(n28810), .Z(n29249) );
  NANDN U29457 ( .A(n28813), .B(n28812), .Z(n28817) );
  NAND U29458 ( .A(n28815), .B(n28814), .Z(n28816) );
  NAND U29459 ( .A(n28817), .B(n28816), .Z(n29194) );
  XNOR U29460 ( .A(a[113]), .B(b[17]), .Z(n29206) );
  NANDN U29461 ( .A(n29206), .B(n32543), .Z(n28820) );
  NANDN U29462 ( .A(n28818), .B(n32541), .Z(n28819) );
  NAND U29463 ( .A(n28820), .B(n28819), .Z(n29226) );
  NANDN U29464 ( .A(n28821), .B(n34848), .Z(n28823) );
  XNOR U29465 ( .A(a[103]), .B(n35375), .Z(n29273) );
  NAND U29466 ( .A(n34618), .B(n29273), .Z(n28822) );
  NAND U29467 ( .A(n28823), .B(n28822), .Z(n29224) );
  NANDN U29468 ( .A(n28824), .B(n33283), .Z(n28826) );
  XNOR U29469 ( .A(a[111]), .B(n33020), .Z(n29200) );
  NANDN U29470 ( .A(n33021), .B(n29200), .Z(n28825) );
  NAND U29471 ( .A(n28826), .B(n28825), .Z(n29225) );
  XNOR U29472 ( .A(n29224), .B(n29225), .Z(n29227) );
  XOR U29473 ( .A(n29226), .B(n29227), .Z(n29191) );
  NAND U29474 ( .A(n37802), .B(n28827), .Z(n28829) );
  XNOR U29475 ( .A(b[51]), .B(a[79]), .Z(n29270) );
  NANDN U29476 ( .A(n29270), .B(n37803), .Z(n28828) );
  AND U29477 ( .A(n28829), .B(n28828), .Z(n29287) );
  NAND U29478 ( .A(n37941), .B(n28830), .Z(n28832) );
  XNOR U29479 ( .A(b[53]), .B(a[77]), .Z(n29240) );
  NANDN U29480 ( .A(n29240), .B(n37940), .Z(n28831) );
  AND U29481 ( .A(n28832), .B(n28831), .Z(n29286) );
  NAND U29482 ( .A(n36643), .B(n28833), .Z(n28835) );
  XNOR U29483 ( .A(n976), .B(a[91]), .Z(n29246) );
  NAND U29484 ( .A(n29246), .B(n36553), .Z(n28834) );
  AND U29485 ( .A(n28835), .B(n28834), .Z(n29285) );
  XNOR U29486 ( .A(n29286), .B(n29285), .Z(n29288) );
  XOR U29487 ( .A(n29287), .B(n29288), .Z(n29192) );
  XNOR U29488 ( .A(n29191), .B(n29192), .Z(n29193) );
  XOR U29489 ( .A(n29194), .B(n29193), .Z(n29250) );
  XOR U29490 ( .A(n29249), .B(n29250), .Z(n29251) );
  XOR U29491 ( .A(n29252), .B(n29251), .Z(n29297) );
  OR U29492 ( .A(n28837), .B(n28836), .Z(n28841) );
  NANDN U29493 ( .A(n28839), .B(n28838), .Z(n28840) );
  AND U29494 ( .A(n28841), .B(n28840), .Z(n29298) );
  XNOR U29495 ( .A(n29297), .B(n29298), .Z(n29299) );
  XNOR U29496 ( .A(n29300), .B(n29299), .Z(n29145) );
  NANDN U29497 ( .A(n28843), .B(n28842), .Z(n28847) );
  NAND U29498 ( .A(n28845), .B(n28844), .Z(n28846) );
  NAND U29499 ( .A(n28847), .B(n28846), .Z(n29074) );
  XNOR U29500 ( .A(b[35]), .B(a[95]), .Z(n29090) );
  NANDN U29501 ( .A(n29090), .B(n35985), .Z(n28850) );
  NANDN U29502 ( .A(n28848), .B(n35986), .Z(n28849) );
  NAND U29503 ( .A(n28850), .B(n28849), .Z(n29182) );
  XNOR U29504 ( .A(a[121]), .B(b[9]), .Z(n29164) );
  NANDN U29505 ( .A(n29164), .B(n30509), .Z(n28853) );
  NANDN U29506 ( .A(n28851), .B(n30846), .Z(n28852) );
  NAND U29507 ( .A(n28853), .B(n28852), .Z(n29179) );
  XNOR U29508 ( .A(b[55]), .B(a[75]), .Z(n29243) );
  NANDN U29509 ( .A(n29243), .B(n38075), .Z(n28856) );
  NANDN U29510 ( .A(n28854), .B(n38073), .Z(n28855) );
  AND U29511 ( .A(n28856), .B(n28855), .Z(n29180) );
  XNOR U29512 ( .A(n29179), .B(n29180), .Z(n29181) );
  XNOR U29513 ( .A(n29182), .B(n29181), .Z(n29072) );
  NANDN U29514 ( .A(n28858), .B(n28857), .Z(n28862) );
  NAND U29515 ( .A(n28860), .B(n28859), .Z(n28861) );
  NAND U29516 ( .A(n28862), .B(n28861), .Z(n29073) );
  XOR U29517 ( .A(n29072), .B(n29073), .Z(n29075) );
  XNOR U29518 ( .A(n29074), .B(n29075), .Z(n29136) );
  XNOR U29519 ( .A(a[117]), .B(b[13]), .Z(n29209) );
  OR U29520 ( .A(n29209), .B(n31550), .Z(n28865) );
  NANDN U29521 ( .A(n28863), .B(n31874), .Z(n28864) );
  NAND U29522 ( .A(n28865), .B(n28864), .Z(n29264) );
  XNOR U29523 ( .A(b[43]), .B(a[87]), .Z(n29279) );
  NANDN U29524 ( .A(n29279), .B(n37068), .Z(n28868) );
  NANDN U29525 ( .A(n28866), .B(n37069), .Z(n28867) );
  NAND U29526 ( .A(n28868), .B(n28867), .Z(n29261) );
  XOR U29527 ( .A(b[45]), .B(a[85]), .Z(n29282) );
  NAND U29528 ( .A(n29282), .B(n37261), .Z(n28871) );
  NANDN U29529 ( .A(n28869), .B(n37262), .Z(n28870) );
  AND U29530 ( .A(n28871), .B(n28870), .Z(n29262) );
  XNOR U29531 ( .A(n29261), .B(n29262), .Z(n29263) );
  XNOR U29532 ( .A(n29264), .B(n29263), .Z(n29118) );
  XNOR U29533 ( .A(n979), .B(a[81]), .Z(n29176) );
  NANDN U29534 ( .A(n37756), .B(n29176), .Z(n28874) );
  NANDN U29535 ( .A(n28872), .B(n37652), .Z(n28873) );
  NAND U29536 ( .A(n28874), .B(n28873), .Z(n29112) );
  NAND U29537 ( .A(n37469), .B(n28875), .Z(n28877) );
  XNOR U29538 ( .A(b[47]), .B(a[83]), .Z(n29173) );
  NANDN U29539 ( .A(n29173), .B(n37471), .Z(n28876) );
  NAND U29540 ( .A(n28877), .B(n28876), .Z(n29109) );
  XOR U29541 ( .A(a[119]), .B(n970), .Z(n29276) );
  OR U29542 ( .A(n29276), .B(n31369), .Z(n28880) );
  NANDN U29543 ( .A(n28878), .B(n31119), .Z(n28879) );
  AND U29544 ( .A(n28880), .B(n28879), .Z(n29110) );
  XNOR U29545 ( .A(n29109), .B(n29110), .Z(n29111) );
  XNOR U29546 ( .A(n29112), .B(n29111), .Z(n29115) );
  NANDN U29547 ( .A(n28882), .B(n28881), .Z(n28886) );
  NAND U29548 ( .A(n28884), .B(n28883), .Z(n28885) );
  NAND U29549 ( .A(n28886), .B(n28885), .Z(n29116) );
  XNOR U29550 ( .A(n29115), .B(n29116), .Z(n29117) );
  XOR U29551 ( .A(n29118), .B(n29117), .Z(n29133) );
  XOR U29552 ( .A(n29133), .B(n29134), .Z(n29135) );
  XOR U29553 ( .A(n29136), .B(n29135), .Z(n29146) );
  XNOR U29554 ( .A(n29145), .B(n29146), .Z(n29147) );
  XNOR U29555 ( .A(n29148), .B(n29147), .Z(n29310) );
  XNOR U29556 ( .A(n29309), .B(n29310), .Z(n29311) );
  OR U29557 ( .A(n28896), .B(n28895), .Z(n28900) );
  NANDN U29558 ( .A(n28898), .B(n28897), .Z(n28899) );
  NAND U29559 ( .A(n28900), .B(n28899), .Z(n29139) );
  NANDN U29560 ( .A(n28902), .B(n28901), .Z(n28906) );
  OR U29561 ( .A(n28904), .B(n28903), .Z(n28905) );
  AND U29562 ( .A(n28906), .B(n28905), .Z(n29140) );
  XNOR U29563 ( .A(n29139), .B(n29140), .Z(n29141) );
  XNOR U29564 ( .A(n29142), .B(n29141), .Z(n29069) );
  NANDN U29565 ( .A(n28908), .B(n28907), .Z(n28912) );
  NAND U29566 ( .A(n28910), .B(n28909), .Z(n28911) );
  NAND U29567 ( .A(n28912), .B(n28911), .Z(n29067) );
  NANDN U29568 ( .A(n28914), .B(n28913), .Z(n28918) );
  NAND U29569 ( .A(n28916), .B(n28915), .Z(n28917) );
  NAND U29570 ( .A(n28918), .B(n28917), .Z(n29130) );
  NANDN U29571 ( .A(n28920), .B(n28919), .Z(n28924) );
  NAND U29572 ( .A(n28922), .B(n28921), .Z(n28923) );
  NAND U29573 ( .A(n28924), .B(n28923), .Z(n29293) );
  XNOR U29574 ( .A(b[57]), .B(a[73]), .Z(n29237) );
  OR U29575 ( .A(n29237), .B(n965), .Z(n28927) );
  NANDN U29576 ( .A(n28925), .B(n38194), .Z(n28926) );
  NAND U29577 ( .A(n28927), .B(n28926), .Z(n29221) );
  NAND U29578 ( .A(n38326), .B(n28928), .Z(n28930) );
  XOR U29579 ( .A(n38400), .B(n30543), .Z(n29102) );
  NANDN U29580 ( .A(n38273), .B(n29102), .Z(n28929) );
  NAND U29581 ( .A(n28930), .B(n28929), .Z(n29218) );
  XOR U29582 ( .A(b[41]), .B(a[89]), .Z(n29215) );
  NANDN U29583 ( .A(n36905), .B(n29215), .Z(n28933) );
  NANDN U29584 ( .A(n28931), .B(n36807), .Z(n28932) );
  AND U29585 ( .A(n28933), .B(n28932), .Z(n29219) );
  XNOR U29586 ( .A(n29218), .B(n29219), .Z(n29220) );
  XNOR U29587 ( .A(n29221), .B(n29220), .Z(n29291) );
  XNOR U29588 ( .A(b[33]), .B(a[97]), .Z(n29084) );
  NANDN U29589 ( .A(n29084), .B(n35620), .Z(n28936) );
  NANDN U29590 ( .A(n28934), .B(n35621), .Z(n28935) );
  NAND U29591 ( .A(n28936), .B(n28935), .Z(n29258) );
  NAND U29592 ( .A(n28938), .B(n28937), .Z(n28941) );
  XNOR U29593 ( .A(n38463), .B(b[3]), .Z(n29234) );
  NAND U29594 ( .A(n29234), .B(n28939), .Z(n28940) );
  NAND U29595 ( .A(n28941), .B(n28940), .Z(n29255) );
  XOR U29596 ( .A(b[63]), .B(n29372), .Z(n29087) );
  NANDN U29597 ( .A(n29087), .B(n38422), .Z(n28944) );
  NANDN U29598 ( .A(n28942), .B(n38423), .Z(n28943) );
  AND U29599 ( .A(n28944), .B(n28943), .Z(n29256) );
  XNOR U29600 ( .A(n29255), .B(n29256), .Z(n29257) );
  XOR U29601 ( .A(n29258), .B(n29257), .Z(n29292) );
  XOR U29602 ( .A(n29291), .B(n29292), .Z(n29294) );
  XNOR U29603 ( .A(n29293), .B(n29294), .Z(n29127) );
  NANDN U29604 ( .A(n28946), .B(n28945), .Z(n28950) );
  NAND U29605 ( .A(n28948), .B(n28947), .Z(n28949) );
  AND U29606 ( .A(n28950), .B(n28949), .Z(n29128) );
  XNOR U29607 ( .A(n29127), .B(n29128), .Z(n29129) );
  XNOR U29608 ( .A(n29130), .B(n29129), .Z(n29151) );
  NANDN U29609 ( .A(n28952), .B(n28951), .Z(n28956) );
  OR U29610 ( .A(n28954), .B(n28953), .Z(n28955) );
  AND U29611 ( .A(n28956), .B(n28955), .Z(n29152) );
  XNOR U29612 ( .A(n29151), .B(n29152), .Z(n29153) );
  NANDN U29613 ( .A(n28958), .B(n28957), .Z(n28962) );
  OR U29614 ( .A(n28960), .B(n28959), .Z(n28961) );
  AND U29615 ( .A(n28962), .B(n28961), .Z(n29304) );
  NANDN U29616 ( .A(n28964), .B(n28963), .Z(n28968) );
  NAND U29617 ( .A(n28966), .B(n28965), .Z(n28967) );
  NAND U29618 ( .A(n28968), .B(n28967), .Z(n29123) );
  XNOR U29619 ( .A(a[115]), .B(b[15]), .Z(n29212) );
  OR U29620 ( .A(n29212), .B(n32010), .Z(n28971) );
  NANDN U29621 ( .A(n28969), .B(n32011), .Z(n28970) );
  NAND U29622 ( .A(n28971), .B(n28970), .Z(n29158) );
  NAND U29623 ( .A(n35188), .B(n28972), .Z(n28974) );
  XNOR U29624 ( .A(a[101]), .B(n35540), .Z(n29161) );
  NANDN U29625 ( .A(n34968), .B(n29161), .Z(n28973) );
  NAND U29626 ( .A(n28974), .B(n28973), .Z(n29155) );
  XNOR U29627 ( .A(a[99]), .B(b[31]), .Z(n29228) );
  NANDN U29628 ( .A(n29228), .B(n35313), .Z(n28977) );
  NANDN U29629 ( .A(n28975), .B(n35311), .Z(n28976) );
  AND U29630 ( .A(n28977), .B(n28976), .Z(n29156) );
  XNOR U29631 ( .A(n29155), .B(n29156), .Z(n29157) );
  XNOR U29632 ( .A(n29158), .B(n29157), .Z(n29121) );
  XOR U29633 ( .A(b[37]), .B(n35377), .Z(n29099) );
  NANDN U29634 ( .A(n29099), .B(n36311), .Z(n28980) );
  NANDN U29635 ( .A(n28978), .B(n36309), .Z(n28979) );
  NAND U29636 ( .A(n28980), .B(n28979), .Z(n29188) );
  XNOR U29637 ( .A(a[123]), .B(n31123), .Z(n29167) );
  NAND U29638 ( .A(n29167), .B(n29949), .Z(n28983) );
  NAND U29639 ( .A(n29948), .B(n28981), .Z(n28982) );
  NAND U29640 ( .A(n28983), .B(n28982), .Z(n29185) );
  XNOR U29641 ( .A(a[125]), .B(b[5]), .Z(n29267) );
  OR U29642 ( .A(n29267), .B(n29363), .Z(n28986) );
  NANDN U29643 ( .A(n28984), .B(n29864), .Z(n28985) );
  AND U29644 ( .A(n28986), .B(n28985), .Z(n29186) );
  XNOR U29645 ( .A(n29185), .B(n29186), .Z(n29187) );
  XOR U29646 ( .A(n29188), .B(n29187), .Z(n29122) );
  XOR U29647 ( .A(n29121), .B(n29122), .Z(n29124) );
  XNOR U29648 ( .A(n29123), .B(n29124), .Z(n29303) );
  NANDN U29649 ( .A(n28988), .B(n28987), .Z(n28992) );
  NAND U29650 ( .A(n28990), .B(n28989), .Z(n28991) );
  NAND U29651 ( .A(n28992), .B(n28991), .Z(n29081) );
  XOR U29652 ( .A(a[109]), .B(b[21]), .Z(n29170) );
  NANDN U29653 ( .A(n33634), .B(n29170), .Z(n28995) );
  NANDN U29654 ( .A(n28993), .B(n33464), .Z(n28994) );
  NAND U29655 ( .A(n28995), .B(n28994), .Z(n29096) );
  NAND U29656 ( .A(n34044), .B(n28996), .Z(n28998) );
  XNOR U29657 ( .A(a[107]), .B(n34510), .Z(n29197) );
  NANDN U29658 ( .A(n33867), .B(n29197), .Z(n28997) );
  NAND U29659 ( .A(n28998), .B(n28997), .Z(n29093) );
  XOR U29660 ( .A(a[105]), .B(b[25]), .Z(n29203) );
  NANDN U29661 ( .A(n34219), .B(n29203), .Z(n29001) );
  NAND U29662 ( .A(n34217), .B(n28999), .Z(n29000) );
  AND U29663 ( .A(n29001), .B(n29000), .Z(n29094) );
  XNOR U29664 ( .A(n29093), .B(n29094), .Z(n29095) );
  XNOR U29665 ( .A(n29096), .B(n29095), .Z(n29079) );
  NANDN U29666 ( .A(n29002), .B(n38369), .Z(n29004) );
  XNOR U29667 ( .A(n984), .B(a[69]), .Z(n29105) );
  NANDN U29668 ( .A(n38371), .B(n29105), .Z(n29003) );
  AND U29669 ( .A(n29004), .B(n29003), .Z(n29108) );
  AND U29670 ( .A(a[65]), .B(b[63]), .Z(n29858) );
  XOR U29671 ( .A(n29858), .B(n29232), .Z(n29005) );
  XNOR U29672 ( .A(n29108), .B(n29005), .Z(n29078) );
  XOR U29673 ( .A(n29079), .B(n29078), .Z(n29080) );
  XOR U29674 ( .A(n29081), .B(n29080), .Z(n29305) );
  XNOR U29675 ( .A(n29306), .B(n29305), .Z(n29154) );
  XNOR U29676 ( .A(n29153), .B(n29154), .Z(n29066) );
  XOR U29677 ( .A(n29067), .B(n29066), .Z(n29068) );
  XOR U29678 ( .A(n29069), .B(n29068), .Z(n29312) );
  XOR U29679 ( .A(n29311), .B(n29312), .Z(n29054) );
  NANDN U29680 ( .A(n29007), .B(n29006), .Z(n29011) );
  OR U29681 ( .A(n29009), .B(n29008), .Z(n29010) );
  NAND U29682 ( .A(n29011), .B(n29010), .Z(n29316) );
  NAND U29683 ( .A(n29013), .B(n29012), .Z(n29017) );
  NANDN U29684 ( .A(n29015), .B(n29014), .Z(n29016) );
  AND U29685 ( .A(n29017), .B(n29016), .Z(n29315) );
  XNOR U29686 ( .A(n29316), .B(n29315), .Z(n29317) );
  OR U29687 ( .A(n29019), .B(n29018), .Z(n29023) );
  NAND U29688 ( .A(n29021), .B(n29020), .Z(n29022) );
  NAND U29689 ( .A(n29023), .B(n29022), .Z(n29318) );
  XNOR U29690 ( .A(n29317), .B(n29318), .Z(n29056) );
  XOR U29691 ( .A(n29057), .B(n29056), .Z(n29063) );
  OR U29692 ( .A(n29025), .B(n29024), .Z(n29029) );
  NANDN U29693 ( .A(n29027), .B(n29026), .Z(n29028) );
  NAND U29694 ( .A(n29029), .B(n29028), .Z(n29060) );
  NANDN U29695 ( .A(n29031), .B(n29030), .Z(n29035) );
  NAND U29696 ( .A(n29033), .B(n29032), .Z(n29034) );
  NAND U29697 ( .A(n29035), .B(n29034), .Z(n29061) );
  XNOR U29698 ( .A(n29060), .B(n29061), .Z(n29062) );
  XNOR U29699 ( .A(n29063), .B(n29062), .Z(n29321) );
  NANDN U29700 ( .A(n29037), .B(n29036), .Z(n29041) );
  NAND U29701 ( .A(n29039), .B(n29038), .Z(n29040) );
  AND U29702 ( .A(n29041), .B(n29040), .Z(n29322) );
  XNOR U29703 ( .A(n29321), .B(n29322), .Z(n29324) );
  NANDN U29704 ( .A(n29043), .B(n29042), .Z(n29047) );
  NANDN U29705 ( .A(n29045), .B(n29044), .Z(n29046) );
  NAND U29706 ( .A(n29047), .B(n29046), .Z(n29323) );
  XNOR U29707 ( .A(n29324), .B(n29323), .Z(n29327) );
  NANDN U29708 ( .A(n29049), .B(n29048), .Z(n29053) );
  NAND U29709 ( .A(n29051), .B(n29050), .Z(n29052) );
  NAND U29710 ( .A(n29053), .B(n29052), .Z(n29328) );
  XNOR U29711 ( .A(n29327), .B(n29328), .Z(n29329) );
  XOR U29712 ( .A(n29330), .B(n29329), .Z(n29334) );
  XOR U29713 ( .A(n29335), .B(n29334), .Z(c[193]) );
  OR U29714 ( .A(n29055), .B(n29054), .Z(n29059) );
  OR U29715 ( .A(n29057), .B(n29056), .Z(n29058) );
  NAND U29716 ( .A(n29059), .B(n29058), .Z(n29344) );
  NANDN U29717 ( .A(n29061), .B(n29060), .Z(n29065) );
  NANDN U29718 ( .A(n29063), .B(n29062), .Z(n29064) );
  NAND U29719 ( .A(n29065), .B(n29064), .Z(n29341) );
  NAND U29720 ( .A(n29067), .B(n29066), .Z(n29071) );
  NANDN U29721 ( .A(n29069), .B(n29068), .Z(n29070) );
  NAND U29722 ( .A(n29071), .B(n29070), .Z(n29350) );
  NANDN U29723 ( .A(n29073), .B(n29072), .Z(n29077) );
  OR U29724 ( .A(n29075), .B(n29074), .Z(n29076) );
  NAND U29725 ( .A(n29077), .B(n29076), .Z(n29351) );
  NAND U29726 ( .A(n29079), .B(n29078), .Z(n29083) );
  NANDN U29727 ( .A(n29081), .B(n29080), .Z(n29082) );
  AND U29728 ( .A(n29083), .B(n29082), .Z(n29352) );
  XNOR U29729 ( .A(n29351), .B(n29352), .Z(n29353) );
  NAND U29730 ( .A(a[66]), .B(b[63]), .Z(n29374) );
  XNOR U29731 ( .A(n974), .B(a[98]), .Z(n29525) );
  NAND U29732 ( .A(n35620), .B(n29525), .Z(n29086) );
  NANDN U29733 ( .A(n29084), .B(n35621), .Z(n29085) );
  AND U29734 ( .A(n29086), .B(n29085), .Z(n29373) );
  XNOR U29735 ( .A(n29858), .B(n29373), .Z(n29375) );
  XNOR U29736 ( .A(n29374), .B(n29375), .Z(n29492) );
  XOR U29737 ( .A(b[63]), .B(n29868), .Z(n29414) );
  NANDN U29738 ( .A(n29414), .B(n38422), .Z(n29089) );
  NANDN U29739 ( .A(n29087), .B(n38423), .Z(n29088) );
  NAND U29740 ( .A(n29089), .B(n29088), .Z(n29489) );
  XNOR U29741 ( .A(b[35]), .B(a[96]), .Z(n29567) );
  NANDN U29742 ( .A(n29567), .B(n35985), .Z(n29092) );
  NANDN U29743 ( .A(n29090), .B(n35986), .Z(n29091) );
  AND U29744 ( .A(n29092), .B(n29091), .Z(n29490) );
  XNOR U29745 ( .A(n29489), .B(n29490), .Z(n29491) );
  XNOR U29746 ( .A(n29492), .B(n29491), .Z(n29467) );
  NANDN U29747 ( .A(n29094), .B(n29093), .Z(n29098) );
  NAND U29748 ( .A(n29096), .B(n29095), .Z(n29097) );
  NAND U29749 ( .A(n29098), .B(n29097), .Z(n29466) );
  XOR U29750 ( .A(b[37]), .B(n35191), .Z(n29367) );
  NANDN U29751 ( .A(n29367), .B(n36311), .Z(n29101) );
  NANDN U29752 ( .A(n29099), .B(n36309), .Z(n29100) );
  NAND U29753 ( .A(n29101), .B(n29100), .Z(n29543) );
  NAND U29754 ( .A(n38326), .B(n29102), .Z(n29104) );
  XOR U29755 ( .A(n38400), .B(n30210), .Z(n29498) );
  NANDN U29756 ( .A(n38273), .B(n29498), .Z(n29103) );
  NAND U29757 ( .A(n29104), .B(n29103), .Z(n29540) );
  XOR U29758 ( .A(b[61]), .B(n30379), .Z(n29501) );
  OR U29759 ( .A(n29501), .B(n38371), .Z(n29107) );
  NAND U29760 ( .A(n29105), .B(n38369), .Z(n29106) );
  AND U29761 ( .A(n29107), .B(n29106), .Z(n29541) );
  XNOR U29762 ( .A(n29540), .B(n29541), .Z(n29542) );
  XOR U29763 ( .A(n29543), .B(n29542), .Z(n29465) );
  XNOR U29764 ( .A(n29466), .B(n29465), .Z(n29468) );
  XNOR U29765 ( .A(n29467), .B(n29468), .Z(n29474) );
  NANDN U29766 ( .A(n29110), .B(n29109), .Z(n29114) );
  NAND U29767 ( .A(n29112), .B(n29111), .Z(n29113) );
  AND U29768 ( .A(n29114), .B(n29113), .Z(n29471) );
  XNOR U29769 ( .A(n29472), .B(n29471), .Z(n29473) );
  XOR U29770 ( .A(n29474), .B(n29473), .Z(n29354) );
  XOR U29771 ( .A(n29353), .B(n29354), .Z(n29595) );
  NANDN U29772 ( .A(n29116), .B(n29115), .Z(n29120) );
  NAND U29773 ( .A(n29118), .B(n29117), .Z(n29119) );
  NAND U29774 ( .A(n29120), .B(n29119), .Z(n29360) );
  NANDN U29775 ( .A(n29122), .B(n29121), .Z(n29126) );
  OR U29776 ( .A(n29124), .B(n29123), .Z(n29125) );
  NAND U29777 ( .A(n29126), .B(n29125), .Z(n29357) );
  NANDN U29778 ( .A(n29128), .B(n29127), .Z(n29132) );
  NAND U29779 ( .A(n29130), .B(n29129), .Z(n29131) );
  NAND U29780 ( .A(n29132), .B(n29131), .Z(n29358) );
  XNOR U29781 ( .A(n29357), .B(n29358), .Z(n29359) );
  XNOR U29782 ( .A(n29360), .B(n29359), .Z(n29592) );
  OR U29783 ( .A(n29134), .B(n29133), .Z(n29138) );
  NAND U29784 ( .A(n29136), .B(n29135), .Z(n29137) );
  AND U29785 ( .A(n29138), .B(n29137), .Z(n29593) );
  XNOR U29786 ( .A(n29592), .B(n29593), .Z(n29594) );
  XNOR U29787 ( .A(n29595), .B(n29594), .Z(n29347) );
  NANDN U29788 ( .A(n29140), .B(n29139), .Z(n29144) );
  NAND U29789 ( .A(n29142), .B(n29141), .Z(n29143) );
  AND U29790 ( .A(n29144), .B(n29143), .Z(n29348) );
  XNOR U29791 ( .A(n29347), .B(n29348), .Z(n29349) );
  XNOR U29792 ( .A(n29350), .B(n29349), .Z(n29603) );
  NANDN U29793 ( .A(n29146), .B(n29145), .Z(n29150) );
  NAND U29794 ( .A(n29148), .B(n29147), .Z(n29149) );
  NAND U29795 ( .A(n29150), .B(n29149), .Z(n29600) );
  NANDN U29796 ( .A(n29156), .B(n29155), .Z(n29160) );
  NAND U29797 ( .A(n29158), .B(n29157), .Z(n29159) );
  NAND U29798 ( .A(n29160), .B(n29159), .Z(n29404) );
  NAND U29799 ( .A(n35188), .B(n29161), .Z(n29163) );
  XOR U29800 ( .A(n36420), .B(n35540), .Z(n29450) );
  NANDN U29801 ( .A(n34968), .B(n29450), .Z(n29162) );
  NAND U29802 ( .A(n29163), .B(n29162), .Z(n29429) );
  XOR U29803 ( .A(n38251), .B(n969), .Z(n29519) );
  NAND U29804 ( .A(n30509), .B(n29519), .Z(n29166) );
  NANDN U29805 ( .A(n29164), .B(n30846), .Z(n29165) );
  NAND U29806 ( .A(n29166), .B(n29165), .Z(n29426) );
  XOR U29807 ( .A(n38321), .B(n31123), .Z(n29411) );
  NAND U29808 ( .A(n29411), .B(n29949), .Z(n29169) );
  NAND U29809 ( .A(n29948), .B(n29167), .Z(n29168) );
  AND U29810 ( .A(n29169), .B(n29168), .Z(n29427) );
  XNOR U29811 ( .A(n29426), .B(n29427), .Z(n29428) );
  XNOR U29812 ( .A(n29429), .B(n29428), .Z(n29402) );
  XNOR U29813 ( .A(n37336), .B(b[21]), .Z(n29435) );
  NANDN U29814 ( .A(n33634), .B(n29435), .Z(n29172) );
  NAND U29815 ( .A(n29170), .B(n33464), .Z(n29171) );
  AND U29816 ( .A(n29172), .B(n29171), .Z(n29485) );
  NANDN U29817 ( .A(n29173), .B(n37469), .Z(n29175) );
  XNOR U29818 ( .A(n978), .B(a[84]), .Z(n29420) );
  NAND U29819 ( .A(n29420), .B(n37471), .Z(n29174) );
  AND U29820 ( .A(n29175), .B(n29174), .Z(n29484) );
  NAND U29821 ( .A(n37652), .B(n29176), .Z(n29178) );
  XOR U29822 ( .A(b[49]), .B(n32815), .Z(n29423) );
  OR U29823 ( .A(n29423), .B(n37756), .Z(n29177) );
  AND U29824 ( .A(n29178), .B(n29177), .Z(n29483) );
  XNOR U29825 ( .A(n29484), .B(n29483), .Z(n29486) );
  XOR U29826 ( .A(n29485), .B(n29486), .Z(n29403) );
  XOR U29827 ( .A(n29402), .B(n29403), .Z(n29405) );
  XNOR U29828 ( .A(n29404), .B(n29405), .Z(n29479) );
  NANDN U29829 ( .A(n29180), .B(n29179), .Z(n29184) );
  NAND U29830 ( .A(n29182), .B(n29181), .Z(n29183) );
  AND U29831 ( .A(n29184), .B(n29183), .Z(n29478) );
  NANDN U29832 ( .A(n29186), .B(n29185), .Z(n29190) );
  NAND U29833 ( .A(n29188), .B(n29187), .Z(n29189) );
  AND U29834 ( .A(n29190), .B(n29189), .Z(n29477) );
  XNOR U29835 ( .A(n29478), .B(n29477), .Z(n29480) );
  XNOR U29836 ( .A(n29479), .B(n29480), .Z(n29462) );
  NANDN U29837 ( .A(n29192), .B(n29191), .Z(n29196) );
  NANDN U29838 ( .A(n29194), .B(n29193), .Z(n29195) );
  NAND U29839 ( .A(n29196), .B(n29195), .Z(n29459) );
  NAND U29840 ( .A(n34044), .B(n29197), .Z(n29199) );
  XOR U29841 ( .A(n37139), .B(n34510), .Z(n29417) );
  NANDN U29842 ( .A(n33867), .B(n29417), .Z(n29198) );
  NAND U29843 ( .A(n29199), .B(n29198), .Z(n29381) );
  NAND U29844 ( .A(n29200), .B(n33283), .Z(n29202) );
  XOR U29845 ( .A(n37583), .B(n33020), .Z(n29438) );
  NANDN U29846 ( .A(n33021), .B(n29438), .Z(n29201) );
  NAND U29847 ( .A(n29202), .B(n29201), .Z(n29378) );
  XNOR U29848 ( .A(n36909), .B(b[25]), .Z(n29441) );
  NANDN U29849 ( .A(n34219), .B(n29441), .Z(n29205) );
  NAND U29850 ( .A(n34217), .B(n29203), .Z(n29204) );
  AND U29851 ( .A(n29205), .B(n29204), .Z(n29379) );
  XNOR U29852 ( .A(n29378), .B(n29379), .Z(n29380) );
  XOR U29853 ( .A(n29381), .B(n29380), .Z(n29504) );
  XNOR U29854 ( .A(a[114]), .B(b[17]), .Z(n29432) );
  NANDN U29855 ( .A(n29432), .B(n32543), .Z(n29208) );
  NANDN U29856 ( .A(n29206), .B(n32541), .Z(n29207) );
  NAND U29857 ( .A(n29208), .B(n29207), .Z(n29505) );
  XNOR U29858 ( .A(n29504), .B(n29505), .Z(n29507) );
  XOR U29859 ( .A(a[118]), .B(n971), .Z(n29552) );
  OR U29860 ( .A(n29552), .B(n31550), .Z(n29211) );
  NANDN U29861 ( .A(n29209), .B(n31874), .Z(n29210) );
  NAND U29862 ( .A(n29211), .B(n29210), .Z(n29549) );
  XOR U29863 ( .A(a[116]), .B(n972), .Z(n29444) );
  OR U29864 ( .A(n29444), .B(n32010), .Z(n29214) );
  NANDN U29865 ( .A(n29212), .B(n32011), .Z(n29213) );
  NAND U29866 ( .A(n29214), .B(n29213), .Z(n29546) );
  XNOR U29867 ( .A(b[41]), .B(a[90]), .Z(n29495) );
  OR U29868 ( .A(n29495), .B(n36905), .Z(n29217) );
  NAND U29869 ( .A(n29215), .B(n36807), .Z(n29216) );
  AND U29870 ( .A(n29217), .B(n29216), .Z(n29547) );
  XNOR U29871 ( .A(n29546), .B(n29547), .Z(n29548) );
  XOR U29872 ( .A(n29549), .B(n29548), .Z(n29506) );
  XNOR U29873 ( .A(n29507), .B(n29506), .Z(n29455) );
  NANDN U29874 ( .A(n29219), .B(n29218), .Z(n29223) );
  NAND U29875 ( .A(n29221), .B(n29220), .Z(n29222) );
  NAND U29876 ( .A(n29223), .B(n29222), .Z(n29453) );
  XOR U29877 ( .A(a[100]), .B(n973), .Z(n29522) );
  NANDN U29878 ( .A(n29522), .B(n35313), .Z(n29230) );
  NANDN U29879 ( .A(n29228), .B(n35311), .Z(n29229) );
  NAND U29880 ( .A(n29230), .B(n29229), .Z(n29393) );
  NANDN U29881 ( .A(n29232), .B(b[2]), .Z(n29231) );
  XOR U29882 ( .A(n967), .B(n29231), .Z(n29236) );
  XOR U29883 ( .A(b[2]), .B(n29232), .Z(n29233) );
  NANDN U29884 ( .A(n29234), .B(n29233), .Z(n29235) );
  AND U29885 ( .A(n29236), .B(n29235), .Z(n29390) );
  XOR U29886 ( .A(b[57]), .B(n31372), .Z(n29564) );
  OR U29887 ( .A(n29564), .B(n965), .Z(n29239) );
  NANDN U29888 ( .A(n29237), .B(n38194), .Z(n29238) );
  AND U29889 ( .A(n29239), .B(n29238), .Z(n29391) );
  XNOR U29890 ( .A(n29390), .B(n29391), .Z(n29392) );
  XOR U29891 ( .A(n29393), .B(n29392), .Z(n29577) );
  XOR U29892 ( .A(n981), .B(n31870), .Z(n29516) );
  NAND U29893 ( .A(n29516), .B(n37940), .Z(n29242) );
  NANDN U29894 ( .A(n29240), .B(n37941), .Z(n29241) );
  NAND U29895 ( .A(n29242), .B(n29241), .Z(n29387) );
  XOR U29896 ( .A(b[55]), .B(n31363), .Z(n29561) );
  NANDN U29897 ( .A(n29561), .B(n38075), .Z(n29245) );
  NANDN U29898 ( .A(n29243), .B(n38073), .Z(n29244) );
  NAND U29899 ( .A(n29245), .B(n29244), .Z(n29384) );
  XOR U29900 ( .A(b[39]), .B(n34852), .Z(n29408) );
  NANDN U29901 ( .A(n29408), .B(n36553), .Z(n29248) );
  NAND U29902 ( .A(n29246), .B(n36643), .Z(n29247) );
  AND U29903 ( .A(n29248), .B(n29247), .Z(n29385) );
  XNOR U29904 ( .A(n29384), .B(n29385), .Z(n29386) );
  XNOR U29905 ( .A(n29387), .B(n29386), .Z(n29576) );
  XOR U29906 ( .A(n29577), .B(n29576), .Z(n29578) );
  XOR U29907 ( .A(n29579), .B(n29578), .Z(n29454) );
  XOR U29908 ( .A(n29453), .B(n29454), .Z(n29456) );
  XNOR U29909 ( .A(n29455), .B(n29456), .Z(n29460) );
  XNOR U29910 ( .A(n29459), .B(n29460), .Z(n29461) );
  XNOR U29911 ( .A(n29462), .B(n29461), .Z(n29586) );
  OR U29912 ( .A(n29250), .B(n29249), .Z(n29254) );
  NANDN U29913 ( .A(n29252), .B(n29251), .Z(n29253) );
  NAND U29914 ( .A(n29254), .B(n29253), .Z(n29585) );
  NANDN U29915 ( .A(n29256), .B(n29255), .Z(n29260) );
  NAND U29916 ( .A(n29258), .B(n29257), .Z(n29259) );
  NAND U29917 ( .A(n29260), .B(n29259), .Z(n29537) );
  NANDN U29918 ( .A(n29262), .B(n29261), .Z(n29266) );
  NAND U29919 ( .A(n29264), .B(n29263), .Z(n29265) );
  NAND U29920 ( .A(n29266), .B(n29265), .Z(n29398) );
  XOR U29921 ( .A(a[126]), .B(n968), .Z(n29364) );
  OR U29922 ( .A(n29364), .B(n29363), .Z(n29269) );
  NANDN U29923 ( .A(n29267), .B(n29864), .Z(n29268) );
  NAND U29924 ( .A(n29269), .B(n29268), .Z(n29573) );
  XOR U29925 ( .A(b[51]), .B(n32814), .Z(n29531) );
  NANDN U29926 ( .A(n29531), .B(n37803), .Z(n29272) );
  NANDN U29927 ( .A(n29270), .B(n37802), .Z(n29271) );
  NAND U29928 ( .A(n29272), .B(n29271), .Z(n29570) );
  NAND U29929 ( .A(n29273), .B(n34848), .Z(n29275) );
  XOR U29930 ( .A(n36647), .B(n35375), .Z(n29447) );
  NAND U29931 ( .A(n34618), .B(n29447), .Z(n29274) );
  AND U29932 ( .A(n29275), .B(n29274), .Z(n29571) );
  XNOR U29933 ( .A(n29570), .B(n29571), .Z(n29572) );
  XNOR U29934 ( .A(n29573), .B(n29572), .Z(n29396) );
  XOR U29935 ( .A(a[120]), .B(n970), .Z(n29528) );
  OR U29936 ( .A(n29528), .B(n31369), .Z(n29278) );
  NANDN U29937 ( .A(n29276), .B(n31119), .Z(n29277) );
  NAND U29938 ( .A(n29278), .B(n29277), .Z(n29513) );
  XOR U29939 ( .A(n977), .B(n34048), .Z(n29555) );
  NAND U29940 ( .A(n29555), .B(n37068), .Z(n29281) );
  NANDN U29941 ( .A(n29279), .B(n37069), .Z(n29280) );
  NAND U29942 ( .A(n29281), .B(n29280), .Z(n29510) );
  XNOR U29943 ( .A(b[45]), .B(a[86]), .Z(n29558) );
  NANDN U29944 ( .A(n29558), .B(n37261), .Z(n29284) );
  NAND U29945 ( .A(n29282), .B(n37262), .Z(n29283) );
  AND U29946 ( .A(n29284), .B(n29283), .Z(n29511) );
  XNOR U29947 ( .A(n29510), .B(n29511), .Z(n29512) );
  XOR U29948 ( .A(n29513), .B(n29512), .Z(n29397) );
  XOR U29949 ( .A(n29396), .B(n29397), .Z(n29399) );
  XNOR U29950 ( .A(n29398), .B(n29399), .Z(n29534) );
  OR U29951 ( .A(n29286), .B(n29285), .Z(n29290) );
  OR U29952 ( .A(n29288), .B(n29287), .Z(n29289) );
  AND U29953 ( .A(n29290), .B(n29289), .Z(n29535) );
  XNOR U29954 ( .A(n29534), .B(n29535), .Z(n29536) );
  XNOR U29955 ( .A(n29537), .B(n29536), .Z(n29582) );
  NANDN U29956 ( .A(n29292), .B(n29291), .Z(n29296) );
  OR U29957 ( .A(n29294), .B(n29293), .Z(n29295) );
  AND U29958 ( .A(n29296), .B(n29295), .Z(n29583) );
  XNOR U29959 ( .A(n29582), .B(n29583), .Z(n29584) );
  XNOR U29960 ( .A(n29585), .B(n29584), .Z(n29587) );
  XNOR U29961 ( .A(n29586), .B(n29587), .Z(n29588) );
  XNOR U29962 ( .A(n29589), .B(n29588), .Z(n29596) );
  NANDN U29963 ( .A(n29298), .B(n29297), .Z(n29302) );
  NAND U29964 ( .A(n29300), .B(n29299), .Z(n29301) );
  AND U29965 ( .A(n29302), .B(n29301), .Z(n29597) );
  XNOR U29966 ( .A(n29596), .B(n29597), .Z(n29598) );
  OR U29967 ( .A(n29304), .B(n29303), .Z(n29308) );
  OR U29968 ( .A(n29306), .B(n29305), .Z(n29307) );
  AND U29969 ( .A(n29308), .B(n29307), .Z(n29599) );
  XNOR U29970 ( .A(n29598), .B(n29599), .Z(n29601) );
  XOR U29971 ( .A(n29600), .B(n29601), .Z(n29602) );
  XOR U29972 ( .A(n29603), .B(n29602), .Z(n29609) );
  NANDN U29973 ( .A(n29310), .B(n29309), .Z(n29314) );
  NANDN U29974 ( .A(n29312), .B(n29311), .Z(n29313) );
  NAND U29975 ( .A(n29314), .B(n29313), .Z(n29606) );
  NANDN U29976 ( .A(n29316), .B(n29315), .Z(n29320) );
  NANDN U29977 ( .A(n29318), .B(n29317), .Z(n29319) );
  NAND U29978 ( .A(n29320), .B(n29319), .Z(n29607) );
  XNOR U29979 ( .A(n29606), .B(n29607), .Z(n29608) );
  XOR U29980 ( .A(n29609), .B(n29608), .Z(n29342) );
  XOR U29981 ( .A(n29341), .B(n29342), .Z(n29343) );
  XNOR U29982 ( .A(n29344), .B(n29343), .Z(n29338) );
  NAND U29983 ( .A(n29322), .B(n29321), .Z(n29326) );
  OR U29984 ( .A(n29324), .B(n29323), .Z(n29325) );
  NAND U29985 ( .A(n29326), .B(n29325), .Z(n29339) );
  NANDN U29986 ( .A(n29328), .B(n29327), .Z(n29332) );
  NAND U29987 ( .A(n29330), .B(n29329), .Z(n29331) );
  AND U29988 ( .A(n29332), .B(n29331), .Z(n29340) );
  XOR U29989 ( .A(n29339), .B(n29340), .Z(n29333) );
  XNOR U29990 ( .A(n29338), .B(n29333), .Z(n29337) );
  OR U29991 ( .A(n29335), .B(n29334), .Z(n29336) );
  XOR U29992 ( .A(n29337), .B(n29336), .Z(c[194]) );
  OR U29993 ( .A(n29337), .B(n29336), .Z(n29892) );
  OR U29994 ( .A(n29342), .B(n29341), .Z(n29346) );
  NAND U29995 ( .A(n29344), .B(n29343), .Z(n29345) );
  NAND U29996 ( .A(n29346), .B(n29345), .Z(n29612) );
  NANDN U29997 ( .A(n29352), .B(n29351), .Z(n29356) );
  NANDN U29998 ( .A(n29354), .B(n29353), .Z(n29355) );
  AND U29999 ( .A(n29356), .B(n29355), .Z(n29630) );
  NANDN U30000 ( .A(n29358), .B(n29357), .Z(n29362) );
  NAND U30001 ( .A(n29360), .B(n29359), .Z(n29361) );
  AND U30002 ( .A(n29362), .B(n29361), .Z(n29631) );
  XOR U30003 ( .A(n29630), .B(n29631), .Z(n29632) );
  XOR U30004 ( .A(a[127]), .B(n968), .Z(n29865) );
  OR U30005 ( .A(n29865), .B(n29363), .Z(n29366) );
  NANDN U30006 ( .A(n29364), .B(n29864), .Z(n29365) );
  NAND U30007 ( .A(n29366), .B(n29365), .Z(n29729) );
  XOR U30008 ( .A(b[37]), .B(n35628), .Z(n29810) );
  NANDN U30009 ( .A(n29810), .B(n36311), .Z(n29369) );
  NANDN U30010 ( .A(n29367), .B(n36309), .Z(n29368) );
  AND U30011 ( .A(n29369), .B(n29368), .Z(n29730) );
  XNOR U30012 ( .A(n29729), .B(n29730), .Z(n29731) );
  NOR U30013 ( .A(n29371), .B(n29370), .Z(n29859) );
  XNOR U30014 ( .A(n29858), .B(n29859), .Z(n29861) );
  NANDN U30015 ( .A(n29372), .B(b[63]), .Z(n29860) );
  XOR U30016 ( .A(n29861), .B(n29860), .Z(n29732) );
  XNOR U30017 ( .A(n29731), .B(n29732), .Z(n29708) );
  NAND U30018 ( .A(n29373), .B(n29858), .Z(n29377) );
  NANDN U30019 ( .A(n29375), .B(n29374), .Z(n29376) );
  NAND U30020 ( .A(n29377), .B(n29376), .Z(n29709) );
  NANDN U30021 ( .A(n29379), .B(n29378), .Z(n29383) );
  NAND U30022 ( .A(n29381), .B(n29380), .Z(n29382) );
  AND U30023 ( .A(n29383), .B(n29382), .Z(n29710) );
  XOR U30024 ( .A(n29711), .B(n29710), .Z(n29780) );
  NANDN U30025 ( .A(n29385), .B(n29384), .Z(n29389) );
  NAND U30026 ( .A(n29387), .B(n29386), .Z(n29388) );
  NAND U30027 ( .A(n29389), .B(n29388), .Z(n29778) );
  NANDN U30028 ( .A(n29391), .B(n29390), .Z(n29395) );
  NAND U30029 ( .A(n29393), .B(n29392), .Z(n29394) );
  AND U30030 ( .A(n29395), .B(n29394), .Z(n29777) );
  XNOR U30031 ( .A(n29778), .B(n29777), .Z(n29779) );
  XOR U30032 ( .A(n29780), .B(n29779), .Z(n29768) );
  NANDN U30033 ( .A(n29397), .B(n29396), .Z(n29401) );
  OR U30034 ( .A(n29399), .B(n29398), .Z(n29400) );
  NAND U30035 ( .A(n29401), .B(n29400), .Z(n29765) );
  NANDN U30036 ( .A(n29403), .B(n29402), .Z(n29407) );
  OR U30037 ( .A(n29405), .B(n29404), .Z(n29406) );
  NAND U30038 ( .A(n29407), .B(n29406), .Z(n29792) );
  XOR U30039 ( .A(b[39]), .B(n35377), .Z(n29726) );
  NANDN U30040 ( .A(n29726), .B(n36553), .Z(n29410) );
  NANDN U30041 ( .A(n29408), .B(n36643), .Z(n29409) );
  NAND U30042 ( .A(n29410), .B(n29409), .Z(n29677) );
  XNOR U30043 ( .A(a[125]), .B(n31123), .Z(n29813) );
  NAND U30044 ( .A(n29813), .B(n29949), .Z(n29413) );
  NAND U30045 ( .A(n29948), .B(n29411), .Z(n29412) );
  NAND U30046 ( .A(n29413), .B(n29412), .Z(n29674) );
  XNOR U30047 ( .A(b[63]), .B(a[69]), .Z(n29869) );
  NANDN U30048 ( .A(n29869), .B(n38422), .Z(n29416) );
  NANDN U30049 ( .A(n29414), .B(n38423), .Z(n29415) );
  AND U30050 ( .A(n29416), .B(n29415), .Z(n29675) );
  XNOR U30051 ( .A(n29674), .B(n29675), .Z(n29676) );
  XOR U30052 ( .A(n29677), .B(n29676), .Z(n29773) );
  NAND U30053 ( .A(n34044), .B(n29417), .Z(n29419) );
  XNOR U30054 ( .A(a[109]), .B(n34510), .Z(n29801) );
  NANDN U30055 ( .A(n33867), .B(n29801), .Z(n29418) );
  NAND U30056 ( .A(n29419), .B(n29418), .Z(n29717) );
  NAND U30057 ( .A(n29420), .B(n37469), .Z(n29422) );
  XNOR U30058 ( .A(n978), .B(a[85]), .Z(n29807) );
  NAND U30059 ( .A(n29807), .B(n37471), .Z(n29421) );
  NAND U30060 ( .A(n29422), .B(n29421), .Z(n29714) );
  XNOR U30061 ( .A(b[49]), .B(a[83]), .Z(n29756) );
  OR U30062 ( .A(n29756), .B(n37756), .Z(n29425) );
  NANDN U30063 ( .A(n29423), .B(n37652), .Z(n29424) );
  AND U30064 ( .A(n29425), .B(n29424), .Z(n29715) );
  XNOR U30065 ( .A(n29714), .B(n29715), .Z(n29716) );
  XOR U30066 ( .A(n29717), .B(n29716), .Z(n29771) );
  NANDN U30067 ( .A(n29427), .B(n29426), .Z(n29431) );
  NAND U30068 ( .A(n29429), .B(n29428), .Z(n29430) );
  NAND U30069 ( .A(n29431), .B(n29430), .Z(n29772) );
  XNOR U30070 ( .A(n29771), .B(n29772), .Z(n29774) );
  XNOR U30071 ( .A(n29773), .B(n29774), .Z(n29790) );
  XNOR U30072 ( .A(a[115]), .B(b[17]), .Z(n29825) );
  NANDN U30073 ( .A(n29825), .B(n32543), .Z(n29434) );
  NANDN U30074 ( .A(n29432), .B(n32541), .Z(n29433) );
  NAND U30075 ( .A(n29434), .B(n29433), .Z(n29760) );
  XOR U30076 ( .A(a[111]), .B(b[21]), .Z(n29828) );
  NANDN U30077 ( .A(n33634), .B(n29828), .Z(n29437) );
  NAND U30078 ( .A(n29435), .B(n33464), .Z(n29436) );
  NAND U30079 ( .A(n29437), .B(n29436), .Z(n29875) );
  NAND U30080 ( .A(n33283), .B(n29438), .Z(n29440) );
  XNOR U30081 ( .A(a[113]), .B(n33020), .Z(n29831) );
  NANDN U30082 ( .A(n33021), .B(n29831), .Z(n29439) );
  NAND U30083 ( .A(n29440), .B(n29439), .Z(n29872) );
  XOR U30084 ( .A(a[107]), .B(b[25]), .Z(n29834) );
  NANDN U30085 ( .A(n34219), .B(n29834), .Z(n29443) );
  NAND U30086 ( .A(n34217), .B(n29441), .Z(n29442) );
  AND U30087 ( .A(n29443), .B(n29442), .Z(n29873) );
  XNOR U30088 ( .A(n29872), .B(n29873), .Z(n29874) );
  XOR U30089 ( .A(n29875), .B(n29874), .Z(n29759) );
  XNOR U30090 ( .A(n29760), .B(n29759), .Z(n29762) );
  XNOR U30091 ( .A(a[117]), .B(b[15]), .Z(n29837) );
  OR U30092 ( .A(n29837), .B(n32010), .Z(n29446) );
  NANDN U30093 ( .A(n29444), .B(n32011), .Z(n29445) );
  NAND U30094 ( .A(n29446), .B(n29445), .Z(n29683) );
  NAND U30095 ( .A(n34848), .B(n29447), .Z(n29449) );
  XNOR U30096 ( .A(a[105]), .B(n35375), .Z(n29840) );
  NAND U30097 ( .A(n34618), .B(n29840), .Z(n29448) );
  NAND U30098 ( .A(n29449), .B(n29448), .Z(n29680) );
  NAND U30099 ( .A(n35188), .B(n29450), .Z(n29452) );
  XNOR U30100 ( .A(a[103]), .B(n35540), .Z(n29843) );
  NANDN U30101 ( .A(n34968), .B(n29843), .Z(n29451) );
  AND U30102 ( .A(n29452), .B(n29451), .Z(n29681) );
  XNOR U30103 ( .A(n29680), .B(n29681), .Z(n29682) );
  XOR U30104 ( .A(n29683), .B(n29682), .Z(n29761) );
  XNOR U30105 ( .A(n29762), .B(n29761), .Z(n29789) );
  XOR U30106 ( .A(n29790), .B(n29789), .Z(n29791) );
  XNOR U30107 ( .A(n29792), .B(n29791), .Z(n29766) );
  XNOR U30108 ( .A(n29765), .B(n29766), .Z(n29767) );
  XOR U30109 ( .A(n29768), .B(n29767), .Z(n29665) );
  NANDN U30110 ( .A(n29454), .B(n29453), .Z(n29458) );
  NANDN U30111 ( .A(n29456), .B(n29455), .Z(n29457) );
  NAND U30112 ( .A(n29458), .B(n29457), .Z(n29662) );
  NANDN U30113 ( .A(n29460), .B(n29459), .Z(n29464) );
  NANDN U30114 ( .A(n29462), .B(n29461), .Z(n29463) );
  NAND U30115 ( .A(n29464), .B(n29463), .Z(n29663) );
  XNOR U30116 ( .A(n29662), .B(n29663), .Z(n29664) );
  XOR U30117 ( .A(n29665), .B(n29664), .Z(n29633) );
  XNOR U30118 ( .A(n29632), .B(n29633), .Z(n29639) );
  OR U30119 ( .A(n29466), .B(n29465), .Z(n29470) );
  OR U30120 ( .A(n29468), .B(n29467), .Z(n29469) );
  NAND U30121 ( .A(n29470), .B(n29469), .Z(n29655) );
  NANDN U30122 ( .A(n29472), .B(n29471), .Z(n29476) );
  NANDN U30123 ( .A(n29474), .B(n29473), .Z(n29475) );
  NAND U30124 ( .A(n29476), .B(n29475), .Z(n29652) );
  OR U30125 ( .A(n29478), .B(n29477), .Z(n29482) );
  NANDN U30126 ( .A(n29480), .B(n29479), .Z(n29481) );
  NAND U30127 ( .A(n29482), .B(n29481), .Z(n29653) );
  XNOR U30128 ( .A(n29652), .B(n29653), .Z(n29654) );
  XNOR U30129 ( .A(n29655), .B(n29654), .Z(n29661) );
  OR U30130 ( .A(n29484), .B(n29483), .Z(n29488) );
  OR U30131 ( .A(n29486), .B(n29485), .Z(n29487) );
  NAND U30132 ( .A(n29488), .B(n29487), .Z(n29783) );
  NANDN U30133 ( .A(n29490), .B(n29489), .Z(n29494) );
  NANDN U30134 ( .A(n29492), .B(n29491), .Z(n29493) );
  AND U30135 ( .A(n29494), .B(n29493), .Z(n29784) );
  XNOR U30136 ( .A(n29783), .B(n29784), .Z(n29785) );
  XOR U30137 ( .A(b[41]), .B(a[91]), .Z(n29689) );
  NANDN U30138 ( .A(n36905), .B(n29689), .Z(n29497) );
  NANDN U30139 ( .A(n29495), .B(n36807), .Z(n29496) );
  NAND U30140 ( .A(n29497), .B(n29496), .Z(n29855) );
  NAND U30141 ( .A(n38326), .B(n29498), .Z(n29500) );
  XNOR U30142 ( .A(n38400), .B(a[73]), .Z(n29723) );
  NANDN U30143 ( .A(n38273), .B(n29723), .Z(n29499) );
  NAND U30144 ( .A(n29500), .B(n29499), .Z(n29852) );
  XOR U30145 ( .A(b[61]), .B(n30543), .Z(n29816) );
  OR U30146 ( .A(n29816), .B(n38371), .Z(n29503) );
  NANDN U30147 ( .A(n29501), .B(n38369), .Z(n29502) );
  AND U30148 ( .A(n29503), .B(n29502), .Z(n29853) );
  XNOR U30149 ( .A(n29852), .B(n29853), .Z(n29854) );
  XNOR U30150 ( .A(n29855), .B(n29854), .Z(n29786) );
  XOR U30151 ( .A(n29785), .B(n29786), .Z(n29645) );
  OR U30152 ( .A(n29505), .B(n29504), .Z(n29509) );
  OR U30153 ( .A(n29507), .B(n29506), .Z(n29508) );
  NAND U30154 ( .A(n29509), .B(n29508), .Z(n29643) );
  NANDN U30155 ( .A(n29511), .B(n29510), .Z(n29515) );
  NAND U30156 ( .A(n29513), .B(n29512), .Z(n29514) );
  NAND U30157 ( .A(n29515), .B(n29514), .Z(n29849) );
  NAND U30158 ( .A(n37941), .B(n29516), .Z(n29518) );
  XNOR U30159 ( .A(b[53]), .B(a[79]), .Z(n29695) );
  NANDN U30160 ( .A(n29695), .B(n37940), .Z(n29517) );
  NAND U30161 ( .A(n29518), .B(n29517), .Z(n29706) );
  NAND U30162 ( .A(n30846), .B(n29519), .Z(n29521) );
  XNOR U30163 ( .A(a[123]), .B(n969), .Z(n29744) );
  NAND U30164 ( .A(n30509), .B(n29744), .Z(n29520) );
  NAND U30165 ( .A(n29521), .B(n29520), .Z(n29704) );
  NANDN U30166 ( .A(n29522), .B(n35311), .Z(n29524) );
  XNOR U30167 ( .A(a[101]), .B(n973), .Z(n29747) );
  NAND U30168 ( .A(n29747), .B(n35313), .Z(n29523) );
  NAND U30169 ( .A(n29524), .B(n29523), .Z(n29705) );
  XNOR U30170 ( .A(n29704), .B(n29705), .Z(n29707) );
  XOR U30171 ( .A(n29706), .B(n29707), .Z(n29846) );
  XNOR U30172 ( .A(b[33]), .B(a[99]), .Z(n29750) );
  NANDN U30173 ( .A(n29750), .B(n35620), .Z(n29527) );
  NAND U30174 ( .A(n29525), .B(n35621), .Z(n29526) );
  NAND U30175 ( .A(n29527), .B(n29526), .Z(n29822) );
  XNOR U30176 ( .A(a[121]), .B(b[11]), .Z(n29753) );
  OR U30177 ( .A(n29753), .B(n31369), .Z(n29530) );
  NANDN U30178 ( .A(n29528), .B(n31119), .Z(n29529) );
  NAND U30179 ( .A(n29530), .B(n29529), .Z(n29819) );
  XNOR U30180 ( .A(b[51]), .B(a[81]), .Z(n29741) );
  NANDN U30181 ( .A(n29741), .B(n37803), .Z(n29533) );
  NANDN U30182 ( .A(n29531), .B(n37802), .Z(n29532) );
  AND U30183 ( .A(n29533), .B(n29532), .Z(n29820) );
  XNOR U30184 ( .A(n29819), .B(n29820), .Z(n29821) );
  XOR U30185 ( .A(n29822), .B(n29821), .Z(n29847) );
  XNOR U30186 ( .A(n29846), .B(n29847), .Z(n29848) );
  XNOR U30187 ( .A(n29849), .B(n29848), .Z(n29642) );
  XOR U30188 ( .A(n29643), .B(n29642), .Z(n29644) );
  XNOR U30189 ( .A(n29645), .B(n29644), .Z(n29658) );
  NANDN U30190 ( .A(n29535), .B(n29534), .Z(n29539) );
  NAND U30191 ( .A(n29537), .B(n29536), .Z(n29538) );
  NAND U30192 ( .A(n29539), .B(n29538), .Z(n29648) );
  NANDN U30193 ( .A(n29541), .B(n29540), .Z(n29545) );
  NAND U30194 ( .A(n29543), .B(n29542), .Z(n29544) );
  NAND U30195 ( .A(n29545), .B(n29544), .Z(n29671) );
  NANDN U30196 ( .A(n29547), .B(n29546), .Z(n29551) );
  NAND U30197 ( .A(n29549), .B(n29548), .Z(n29550) );
  NAND U30198 ( .A(n29551), .B(n29550), .Z(n29797) );
  XOR U30199 ( .A(a[119]), .B(n971), .Z(n29686) );
  OR U30200 ( .A(n29686), .B(n31550), .Z(n29554) );
  NANDN U30201 ( .A(n29552), .B(n31874), .Z(n29553) );
  NAND U30202 ( .A(n29554), .B(n29553), .Z(n29738) );
  XNOR U30203 ( .A(b[43]), .B(a[89]), .Z(n29692) );
  NANDN U30204 ( .A(n29692), .B(n37068), .Z(n29557) );
  NAND U30205 ( .A(n29555), .B(n37069), .Z(n29556) );
  NAND U30206 ( .A(n29557), .B(n29556), .Z(n29735) );
  XOR U30207 ( .A(b[45]), .B(a[87]), .Z(n29804) );
  NAND U30208 ( .A(n29804), .B(n37261), .Z(n29560) );
  NANDN U30209 ( .A(n29558), .B(n37262), .Z(n29559) );
  AND U30210 ( .A(n29560), .B(n29559), .Z(n29736) );
  XNOR U30211 ( .A(n29735), .B(n29736), .Z(n29737) );
  XNOR U30212 ( .A(n29738), .B(n29737), .Z(n29795) );
  XNOR U30213 ( .A(b[55]), .B(a[77]), .Z(n29698) );
  NANDN U30214 ( .A(n29698), .B(n38075), .Z(n29563) );
  NANDN U30215 ( .A(n29561), .B(n38073), .Z(n29562) );
  NAND U30216 ( .A(n29563), .B(n29562), .Z(n29881) );
  XNOR U30217 ( .A(b[57]), .B(a[75]), .Z(n29720) );
  OR U30218 ( .A(n29720), .B(n965), .Z(n29566) );
  NANDN U30219 ( .A(n29564), .B(n38194), .Z(n29565) );
  NAND U30220 ( .A(n29566), .B(n29565), .Z(n29878) );
  XOR U30221 ( .A(b[35]), .B(a[97]), .Z(n29701) );
  NAND U30222 ( .A(n35985), .B(n29701), .Z(n29569) );
  NANDN U30223 ( .A(n29567), .B(n35986), .Z(n29568) );
  AND U30224 ( .A(n29569), .B(n29568), .Z(n29879) );
  XNOR U30225 ( .A(n29878), .B(n29879), .Z(n29880) );
  XOR U30226 ( .A(n29881), .B(n29880), .Z(n29796) );
  XOR U30227 ( .A(n29795), .B(n29796), .Z(n29798) );
  XNOR U30228 ( .A(n29797), .B(n29798), .Z(n29668) );
  NANDN U30229 ( .A(n29571), .B(n29570), .Z(n29575) );
  NAND U30230 ( .A(n29573), .B(n29572), .Z(n29574) );
  AND U30231 ( .A(n29575), .B(n29574), .Z(n29669) );
  XNOR U30232 ( .A(n29668), .B(n29669), .Z(n29670) );
  XNOR U30233 ( .A(n29671), .B(n29670), .Z(n29646) );
  NANDN U30234 ( .A(n29577), .B(n29576), .Z(n29581) );
  OR U30235 ( .A(n29579), .B(n29578), .Z(n29580) );
  AND U30236 ( .A(n29581), .B(n29580), .Z(n29647) );
  XOR U30237 ( .A(n29646), .B(n29647), .Z(n29649) );
  XOR U30238 ( .A(n29648), .B(n29649), .Z(n29659) );
  XNOR U30239 ( .A(n29658), .B(n29659), .Z(n29660) );
  XOR U30240 ( .A(n29661), .B(n29660), .Z(n29636) );
  XOR U30241 ( .A(n29636), .B(n29637), .Z(n29638) );
  XNOR U30242 ( .A(n29639), .B(n29638), .Z(n29627) );
  NANDN U30243 ( .A(n29587), .B(n29586), .Z(n29591) );
  NAND U30244 ( .A(n29589), .B(n29588), .Z(n29590) );
  NAND U30245 ( .A(n29591), .B(n29590), .Z(n29624) );
  XNOR U30246 ( .A(n29624), .B(n29625), .Z(n29626) );
  XNOR U30247 ( .A(n29627), .B(n29626), .Z(n29618) );
  XNOR U30248 ( .A(n29619), .B(n29618), .Z(n29621) );
  XNOR U30249 ( .A(n29621), .B(n29620), .Z(n29884) );
  OR U30250 ( .A(n29601), .B(n29600), .Z(n29605) );
  NAND U30251 ( .A(n29603), .B(n29602), .Z(n29604) );
  AND U30252 ( .A(n29605), .B(n29604), .Z(n29885) );
  XNOR U30253 ( .A(n29884), .B(n29885), .Z(n29886) );
  NANDN U30254 ( .A(n29607), .B(n29606), .Z(n29611) );
  NANDN U30255 ( .A(n29609), .B(n29608), .Z(n29610) );
  NAND U30256 ( .A(n29611), .B(n29610), .Z(n29887) );
  XNOR U30257 ( .A(n29886), .B(n29887), .Z(n29613) );
  XNOR U30258 ( .A(n29612), .B(n29613), .Z(n29614) );
  XNOR U30259 ( .A(n29615), .B(n29614), .Z(n29891) );
  XOR U30260 ( .A(n29892), .B(n29891), .Z(c[195]) );
  NANDN U30261 ( .A(n29613), .B(n29612), .Z(n29617) );
  NANDN U30262 ( .A(n29615), .B(n29614), .Z(n29616) );
  NAND U30263 ( .A(n29617), .B(n29616), .Z(n29895) );
  NAND U30264 ( .A(n29619), .B(n29618), .Z(n29623) );
  OR U30265 ( .A(n29621), .B(n29620), .Z(n29622) );
  NAND U30266 ( .A(n29623), .B(n29622), .Z(n30163) );
  NANDN U30267 ( .A(n29625), .B(n29624), .Z(n29629) );
  NANDN U30268 ( .A(n29627), .B(n29626), .Z(n29628) );
  NAND U30269 ( .A(n29629), .B(n29628), .Z(n30160) );
  OR U30270 ( .A(n29631), .B(n29630), .Z(n29635) );
  NANDN U30271 ( .A(n29633), .B(n29632), .Z(n29634) );
  NAND U30272 ( .A(n29635), .B(n29634), .Z(n30157) );
  NAND U30273 ( .A(n29637), .B(n29636), .Z(n29641) );
  NANDN U30274 ( .A(n29639), .B(n29638), .Z(n29640) );
  NAND U30275 ( .A(n29641), .B(n29640), .Z(n30155) );
  NANDN U30276 ( .A(n29647), .B(n29646), .Z(n29651) );
  OR U30277 ( .A(n29649), .B(n29648), .Z(n29650) );
  NAND U30278 ( .A(n29651), .B(n29650), .Z(n30143) );
  NANDN U30279 ( .A(n29653), .B(n29652), .Z(n29657) );
  NAND U30280 ( .A(n29655), .B(n29654), .Z(n29656) );
  AND U30281 ( .A(n29657), .B(n29656), .Z(n30142) );
  XNOR U30282 ( .A(n30143), .B(n30142), .Z(n30144) );
  XOR U30283 ( .A(n30145), .B(n30144), .Z(n30148) );
  XNOR U30284 ( .A(n30148), .B(n30149), .Z(n30150) );
  NANDN U30285 ( .A(n29663), .B(n29662), .Z(n29667) );
  NAND U30286 ( .A(n29665), .B(n29664), .Z(n29666) );
  NAND U30287 ( .A(n29667), .B(n29666), .Z(n29899) );
  NANDN U30288 ( .A(n29669), .B(n29668), .Z(n29673) );
  NAND U30289 ( .A(n29671), .B(n29670), .Z(n29672) );
  NAND U30290 ( .A(n29673), .B(n29672), .Z(n29916) );
  NANDN U30291 ( .A(n29675), .B(n29674), .Z(n29679) );
  NAND U30292 ( .A(n29677), .B(n29676), .Z(n29678) );
  NAND U30293 ( .A(n29679), .B(n29678), .Z(n30109) );
  NANDN U30294 ( .A(n29681), .B(n29680), .Z(n29685) );
  NAND U30295 ( .A(n29683), .B(n29682), .Z(n29684) );
  NAND U30296 ( .A(n29685), .B(n29684), .Z(n30132) );
  XOR U30297 ( .A(a[120]), .B(n971), .Z(n29979) );
  OR U30298 ( .A(n29979), .B(n31550), .Z(n29688) );
  NANDN U30299 ( .A(n29686), .B(n31874), .Z(n29687) );
  NAND U30300 ( .A(n29688), .B(n29687), .Z(n29941) );
  XNOR U30301 ( .A(b[41]), .B(a[92]), .Z(n30021) );
  OR U30302 ( .A(n30021), .B(n36905), .Z(n29691) );
  NAND U30303 ( .A(n29689), .B(n36807), .Z(n29690) );
  NAND U30304 ( .A(n29691), .B(n29690), .Z(n29938) );
  XOR U30305 ( .A(b[43]), .B(n34851), .Z(n30056) );
  NANDN U30306 ( .A(n30056), .B(n37068), .Z(n29694) );
  NANDN U30307 ( .A(n29692), .B(n37069), .Z(n29693) );
  AND U30308 ( .A(n29694), .B(n29693), .Z(n29939) );
  XNOR U30309 ( .A(n29938), .B(n29939), .Z(n29940) );
  XNOR U30310 ( .A(n29941), .B(n29940), .Z(n30130) );
  XOR U30311 ( .A(b[53]), .B(n32814), .Z(n29985) );
  NANDN U30312 ( .A(n29985), .B(n37940), .Z(n29697) );
  NANDN U30313 ( .A(n29695), .B(n37941), .Z(n29696) );
  NAND U30314 ( .A(n29697), .B(n29696), .Z(n30033) );
  XOR U30315 ( .A(b[55]), .B(n31870), .Z(n30088) );
  NANDN U30316 ( .A(n30088), .B(n38075), .Z(n29700) );
  NANDN U30317 ( .A(n29698), .B(n38073), .Z(n29699) );
  NAND U30318 ( .A(n29700), .B(n29699), .Z(n30030) );
  XNOR U30319 ( .A(b[35]), .B(a[98]), .Z(n30047) );
  NANDN U30320 ( .A(n30047), .B(n35985), .Z(n29703) );
  NAND U30321 ( .A(n29701), .B(n35986), .Z(n29702) );
  AND U30322 ( .A(n29703), .B(n29702), .Z(n30031) );
  XNOR U30323 ( .A(n30030), .B(n30031), .Z(n30032) );
  XOR U30324 ( .A(n30033), .B(n30032), .Z(n30131) );
  XOR U30325 ( .A(n30130), .B(n30131), .Z(n30133) );
  XNOR U30326 ( .A(n30132), .B(n30133), .Z(n30106) );
  XNOR U30327 ( .A(n30106), .B(n30107), .Z(n30108) );
  XNOR U30328 ( .A(n30109), .B(n30108), .Z(n29914) );
  OR U30329 ( .A(n29709), .B(n29708), .Z(n29713) );
  OR U30330 ( .A(n29711), .B(n29710), .Z(n29712) );
  NAND U30331 ( .A(n29713), .B(n29712), .Z(n29915) );
  XOR U30332 ( .A(n29914), .B(n29915), .Z(n29917) );
  XNOR U30333 ( .A(n29916), .B(n29917), .Z(n29902) );
  NANDN U30334 ( .A(n29715), .B(n29714), .Z(n29719) );
  NAND U30335 ( .A(n29717), .B(n29716), .Z(n29718) );
  NAND U30336 ( .A(n29719), .B(n29718), .Z(n30120) );
  XOR U30337 ( .A(b[57]), .B(n31363), .Z(n30018) );
  OR U30338 ( .A(n30018), .B(n965), .Z(n29722) );
  NANDN U30339 ( .A(n29720), .B(n38194), .Z(n29721) );
  NAND U30340 ( .A(n29722), .B(n29721), .Z(n29967) );
  NAND U30341 ( .A(n38326), .B(n29723), .Z(n29725) );
  XOR U30342 ( .A(n38400), .B(n31372), .Z(n29944) );
  NANDN U30343 ( .A(n38273), .B(n29944), .Z(n29724) );
  NAND U30344 ( .A(n29725), .B(n29724), .Z(n29964) );
  XOR U30345 ( .A(b[39]), .B(n35191), .Z(n29955) );
  NANDN U30346 ( .A(n29955), .B(n36553), .Z(n29728) );
  NANDN U30347 ( .A(n29726), .B(n36643), .Z(n29727) );
  AND U30348 ( .A(n29728), .B(n29727), .Z(n29965) );
  XNOR U30349 ( .A(n29964), .B(n29965), .Z(n29966) );
  XNOR U30350 ( .A(n29967), .B(n29966), .Z(n30118) );
  NANDN U30351 ( .A(n29730), .B(n29729), .Z(n29734) );
  NAND U30352 ( .A(n29732), .B(n29731), .Z(n29733) );
  NAND U30353 ( .A(n29734), .B(n29733), .Z(n30119) );
  XOR U30354 ( .A(n30118), .B(n30119), .Z(n30121) );
  XNOR U30355 ( .A(n30120), .B(n30121), .Z(n29911) );
  NANDN U30356 ( .A(n29736), .B(n29735), .Z(n29740) );
  NAND U30357 ( .A(n29738), .B(n29737), .Z(n29739) );
  NAND U30358 ( .A(n29740), .B(n29739), .Z(n30114) );
  XOR U30359 ( .A(b[51]), .B(n32815), .Z(n30085) );
  NANDN U30360 ( .A(n30085), .B(n37803), .Z(n29743) );
  NANDN U30361 ( .A(n29741), .B(n37802), .Z(n29742) );
  NAND U30362 ( .A(n29743), .B(n29742), .Z(n30073) );
  XOR U30363 ( .A(a[124]), .B(n969), .Z(n30015) );
  NANDN U30364 ( .A(n30015), .B(n30509), .Z(n29746) );
  NAND U30365 ( .A(n29744), .B(n30846), .Z(n29745) );
  NAND U30366 ( .A(n29746), .B(n29745), .Z(n30070) );
  XOR U30367 ( .A(a[102]), .B(n973), .Z(n29976) );
  NANDN U30368 ( .A(n29976), .B(n35313), .Z(n29749) );
  NAND U30369 ( .A(n29747), .B(n35311), .Z(n29748) );
  AND U30370 ( .A(n29749), .B(n29748), .Z(n30071) );
  XNOR U30371 ( .A(n30070), .B(n30071), .Z(n30072) );
  XNOR U30372 ( .A(n30073), .B(n30072), .Z(n30112) );
  XOR U30373 ( .A(a[100]), .B(n974), .Z(n29952) );
  NANDN U30374 ( .A(n29952), .B(n35620), .Z(n29752) );
  NANDN U30375 ( .A(n29750), .B(n35621), .Z(n29751) );
  NAND U30376 ( .A(n29752), .B(n29751), .Z(n30079) );
  XOR U30377 ( .A(a[122]), .B(n970), .Z(n29982) );
  OR U30378 ( .A(n29982), .B(n31369), .Z(n29755) );
  NANDN U30379 ( .A(n29753), .B(n31119), .Z(n29754) );
  NAND U30380 ( .A(n29755), .B(n29754), .Z(n30076) );
  XOR U30381 ( .A(b[49]), .B(n33185), .Z(n30097) );
  OR U30382 ( .A(n30097), .B(n37756), .Z(n29758) );
  NANDN U30383 ( .A(n29756), .B(n37652), .Z(n29757) );
  AND U30384 ( .A(n29758), .B(n29757), .Z(n30077) );
  XNOR U30385 ( .A(n30076), .B(n30077), .Z(n30078) );
  XOR U30386 ( .A(n30079), .B(n30078), .Z(n30113) );
  XOR U30387 ( .A(n30112), .B(n30113), .Z(n30115) );
  XNOR U30388 ( .A(n30114), .B(n30115), .Z(n29908) );
  OR U30389 ( .A(n29760), .B(n29759), .Z(n29764) );
  OR U30390 ( .A(n29762), .B(n29761), .Z(n29763) );
  NAND U30391 ( .A(n29764), .B(n29763), .Z(n29909) );
  XNOR U30392 ( .A(n29908), .B(n29909), .Z(n29910) );
  XNOR U30393 ( .A(n29911), .B(n29910), .Z(n29903) );
  XNOR U30394 ( .A(n29902), .B(n29903), .Z(n29904) );
  NANDN U30395 ( .A(n29766), .B(n29765), .Z(n29770) );
  NANDN U30396 ( .A(n29768), .B(n29767), .Z(n29769) );
  NAND U30397 ( .A(n29770), .B(n29769), .Z(n29905) );
  XOR U30398 ( .A(n29904), .B(n29905), .Z(n29897) );
  OR U30399 ( .A(n29772), .B(n29771), .Z(n29776) );
  OR U30400 ( .A(n29774), .B(n29773), .Z(n29775) );
  NAND U30401 ( .A(n29776), .B(n29775), .Z(n29923) );
  NANDN U30402 ( .A(n29778), .B(n29777), .Z(n29782) );
  NANDN U30403 ( .A(n29780), .B(n29779), .Z(n29781) );
  NAND U30404 ( .A(n29782), .B(n29781), .Z(n29921) );
  NANDN U30405 ( .A(n29784), .B(n29783), .Z(n29788) );
  NANDN U30406 ( .A(n29786), .B(n29785), .Z(n29787) );
  AND U30407 ( .A(n29788), .B(n29787), .Z(n29920) );
  XOR U30408 ( .A(n29921), .B(n29920), .Z(n29922) );
  XNOR U30409 ( .A(n29923), .B(n29922), .Z(n29928) );
  OR U30410 ( .A(n29790), .B(n29789), .Z(n29794) );
  NAND U30411 ( .A(n29792), .B(n29791), .Z(n29793) );
  NAND U30412 ( .A(n29794), .B(n29793), .Z(n29927) );
  NANDN U30413 ( .A(n29796), .B(n29795), .Z(n29800) );
  OR U30414 ( .A(n29798), .B(n29797), .Z(n29799) );
  NAND U30415 ( .A(n29800), .B(n29799), .Z(n29932) );
  NAND U30416 ( .A(n34044), .B(n29801), .Z(n29803) );
  XOR U30417 ( .A(n37336), .B(n34510), .Z(n30006) );
  NANDN U30418 ( .A(n33867), .B(n30006), .Z(n29802) );
  NAND U30419 ( .A(n29803), .B(n29802), .Z(n29973) );
  XNOR U30420 ( .A(b[45]), .B(a[88]), .Z(n30009) );
  NANDN U30421 ( .A(n30009), .B(n37261), .Z(n29806) );
  NAND U30422 ( .A(n29804), .B(n37262), .Z(n29805) );
  NAND U30423 ( .A(n29806), .B(n29805), .Z(n29970) );
  NAND U30424 ( .A(n37469), .B(n29807), .Z(n29809) );
  XOR U30425 ( .A(n978), .B(n33628), .Z(n30094) );
  NAND U30426 ( .A(n30094), .B(n37471), .Z(n29808) );
  AND U30427 ( .A(n29809), .B(n29808), .Z(n29971) );
  XNOR U30428 ( .A(n29970), .B(n29971), .Z(n29972) );
  XNOR U30429 ( .A(n29973), .B(n29972), .Z(n30136) );
  XOR U30430 ( .A(b[37]), .B(n35545), .Z(n30044) );
  NANDN U30431 ( .A(n30044), .B(n36311), .Z(n29812) );
  NANDN U30432 ( .A(n29810), .B(n36309), .Z(n29811) );
  NAND U30433 ( .A(n29812), .B(n29811), .Z(n30027) );
  XOR U30434 ( .A(n987), .B(n31123), .Z(n29947) );
  NAND U30435 ( .A(n29947), .B(n29949), .Z(n29815) );
  NAND U30436 ( .A(n29948), .B(n29813), .Z(n29814) );
  NAND U30437 ( .A(n29815), .B(n29814), .Z(n30024) );
  XOR U30438 ( .A(b[61]), .B(n30210), .Z(n29958) );
  OR U30439 ( .A(n29958), .B(n38371), .Z(n29818) );
  NANDN U30440 ( .A(n29816), .B(n38369), .Z(n29817) );
  AND U30441 ( .A(n29818), .B(n29817), .Z(n30025) );
  XNOR U30442 ( .A(n30024), .B(n30025), .Z(n30026) );
  XOR U30443 ( .A(n30027), .B(n30026), .Z(n30137) );
  XOR U30444 ( .A(n30136), .B(n30137), .Z(n30139) );
  NANDN U30445 ( .A(n29820), .B(n29819), .Z(n29824) );
  NAND U30446 ( .A(n29822), .B(n29821), .Z(n29823) );
  NAND U30447 ( .A(n29824), .B(n29823), .Z(n30138) );
  XNOR U30448 ( .A(n30139), .B(n30138), .Z(n30100) );
  XNOR U30449 ( .A(n38046), .B(b[17]), .Z(n29988) );
  NAND U30450 ( .A(n29988), .B(n32543), .Z(n29827) );
  NANDN U30451 ( .A(n29825), .B(n32541), .Z(n29826) );
  NAND U30452 ( .A(n29827), .B(n29826), .Z(n30037) );
  XNOR U30453 ( .A(a[112]), .B(b[21]), .Z(n30091) );
  OR U30454 ( .A(n30091), .B(n33634), .Z(n29830) );
  NAND U30455 ( .A(n29828), .B(n33464), .Z(n29829) );
  NAND U30456 ( .A(n29830), .B(n29829), .Z(n30003) );
  NAND U30457 ( .A(n33283), .B(n29831), .Z(n29833) );
  XOR U30458 ( .A(n37873), .B(n33020), .Z(n30082) );
  NANDN U30459 ( .A(n33021), .B(n30082), .Z(n29832) );
  NAND U30460 ( .A(n29833), .B(n29832), .Z(n30000) );
  XNOR U30461 ( .A(n37139), .B(b[25]), .Z(n30012) );
  NANDN U30462 ( .A(n34219), .B(n30012), .Z(n29836) );
  NAND U30463 ( .A(n34217), .B(n29834), .Z(n29835) );
  AND U30464 ( .A(n29836), .B(n29835), .Z(n30001) );
  XNOR U30465 ( .A(n30000), .B(n30001), .Z(n30002) );
  XOR U30466 ( .A(n30003), .B(n30002), .Z(n30036) );
  XNOR U30467 ( .A(n30037), .B(n30036), .Z(n30039) );
  XOR U30468 ( .A(a[118]), .B(n972), .Z(n29991) );
  OR U30469 ( .A(n29991), .B(n32010), .Z(n29839) );
  NANDN U30470 ( .A(n29837), .B(n32011), .Z(n29838) );
  NAND U30471 ( .A(n29839), .B(n29838), .Z(n30062) );
  NAND U30472 ( .A(n34848), .B(n29840), .Z(n29842) );
  XOR U30473 ( .A(n36909), .B(n35375), .Z(n30050) );
  NAND U30474 ( .A(n34618), .B(n30050), .Z(n29841) );
  NAND U30475 ( .A(n29842), .B(n29841), .Z(n30059) );
  NAND U30476 ( .A(n35188), .B(n29843), .Z(n29845) );
  XOR U30477 ( .A(n36647), .B(n35540), .Z(n30053) );
  NANDN U30478 ( .A(n34968), .B(n30053), .Z(n29844) );
  AND U30479 ( .A(n29845), .B(n29844), .Z(n30060) );
  XNOR U30480 ( .A(n30059), .B(n30060), .Z(n30061) );
  XOR U30481 ( .A(n30062), .B(n30061), .Z(n30038) );
  XOR U30482 ( .A(n30039), .B(n30038), .Z(n30101) );
  XNOR U30483 ( .A(n30100), .B(n30101), .Z(n30102) );
  NANDN U30484 ( .A(n29847), .B(n29846), .Z(n29851) );
  NANDN U30485 ( .A(n29849), .B(n29848), .Z(n29850) );
  NAND U30486 ( .A(n29851), .B(n29850), .Z(n30103) );
  XNOR U30487 ( .A(n30102), .B(n30103), .Z(n29933) );
  XNOR U30488 ( .A(n29932), .B(n29933), .Z(n29934) );
  NANDN U30489 ( .A(n29853), .B(n29852), .Z(n29857) );
  NAND U30490 ( .A(n29855), .B(n29854), .Z(n29856) );
  NAND U30491 ( .A(n29857), .B(n29856), .Z(n30127) );
  NAND U30492 ( .A(n29859), .B(n29858), .Z(n29863) );
  OR U30493 ( .A(n29861), .B(n29860), .Z(n29862) );
  AND U30494 ( .A(n29863), .B(n29862), .Z(n29995) );
  NANDN U30495 ( .A(n29865), .B(n29864), .Z(n29867) );
  ANDN U30496 ( .B(n29867), .A(n29866), .Z(n30066) );
  ANDN U30497 ( .B(b[63]), .A(n29868), .Z(n30265) );
  XOR U30498 ( .A(b[63]), .B(n30379), .Z(n29961) );
  NANDN U30499 ( .A(n29961), .B(n38422), .Z(n29871) );
  NANDN U30500 ( .A(n29869), .B(n38423), .Z(n29870) );
  AND U30501 ( .A(n29871), .B(n29870), .Z(n30065) );
  XNOR U30502 ( .A(n30265), .B(n30065), .Z(n30067) );
  XNOR U30503 ( .A(n30066), .B(n30067), .Z(n29994) );
  NANDN U30504 ( .A(n29873), .B(n29872), .Z(n29877) );
  NAND U30505 ( .A(n29875), .B(n29874), .Z(n29876) );
  AND U30506 ( .A(n29877), .B(n29876), .Z(n29996) );
  XOR U30507 ( .A(n29997), .B(n29996), .Z(n30124) );
  NANDN U30508 ( .A(n29879), .B(n29878), .Z(n29883) );
  NAND U30509 ( .A(n29881), .B(n29880), .Z(n29882) );
  NAND U30510 ( .A(n29883), .B(n29882), .Z(n30125) );
  XOR U30511 ( .A(n30124), .B(n30125), .Z(n30126) );
  XOR U30512 ( .A(n30127), .B(n30126), .Z(n29935) );
  XNOR U30513 ( .A(n29934), .B(n29935), .Z(n29926) );
  XNOR U30514 ( .A(n29927), .B(n29926), .Z(n29929) );
  XOR U30515 ( .A(n29928), .B(n29929), .Z(n29896) );
  XOR U30516 ( .A(n29897), .B(n29896), .Z(n29898) );
  XOR U30517 ( .A(n29899), .B(n29898), .Z(n30151) );
  XNOR U30518 ( .A(n30150), .B(n30151), .Z(n30154) );
  XNOR U30519 ( .A(n30155), .B(n30154), .Z(n30156) );
  XNOR U30520 ( .A(n30157), .B(n30156), .Z(n30161) );
  XNOR U30521 ( .A(n30160), .B(n30161), .Z(n30162) );
  XNOR U30522 ( .A(n30163), .B(n30162), .Z(n29893) );
  NANDN U30523 ( .A(n29885), .B(n29884), .Z(n29889) );
  NANDN U30524 ( .A(n29887), .B(n29886), .Z(n29888) );
  AND U30525 ( .A(n29889), .B(n29888), .Z(n29894) );
  XOR U30526 ( .A(n29893), .B(n29894), .Z(n29890) );
  XNOR U30527 ( .A(n29895), .B(n29890), .Z(n30167) );
  OR U30528 ( .A(n29892), .B(n29891), .Z(n30166) );
  XOR U30529 ( .A(n30167), .B(n30166), .Z(c[196]) );
  NAND U30530 ( .A(n29897), .B(n29896), .Z(n29901) );
  NANDN U30531 ( .A(n29899), .B(n29898), .Z(n29900) );
  NAND U30532 ( .A(n29901), .B(n29900), .Z(n30436) );
  NANDN U30533 ( .A(n29903), .B(n29902), .Z(n29907) );
  NANDN U30534 ( .A(n29905), .B(n29904), .Z(n29906) );
  NAND U30535 ( .A(n29907), .B(n29906), .Z(n30429) );
  NANDN U30536 ( .A(n29909), .B(n29908), .Z(n29913) );
  NAND U30537 ( .A(n29911), .B(n29910), .Z(n29912) );
  NAND U30538 ( .A(n29913), .B(n29912), .Z(n30185) );
  NANDN U30539 ( .A(n29915), .B(n29914), .Z(n29919) );
  OR U30540 ( .A(n29917), .B(n29916), .Z(n29918) );
  NAND U30541 ( .A(n29919), .B(n29918), .Z(n30182) );
  OR U30542 ( .A(n29921), .B(n29920), .Z(n29925) );
  NANDN U30543 ( .A(n29923), .B(n29922), .Z(n29924) );
  NAND U30544 ( .A(n29925), .B(n29924), .Z(n30183) );
  XNOR U30545 ( .A(n30182), .B(n30183), .Z(n30184) );
  XOR U30546 ( .A(n30185), .B(n30184), .Z(n30430) );
  XOR U30547 ( .A(n30429), .B(n30430), .Z(n30431) );
  NAND U30548 ( .A(n29927), .B(n29926), .Z(n29931) );
  OR U30549 ( .A(n29929), .B(n29928), .Z(n29930) );
  NAND U30550 ( .A(n29931), .B(n29930), .Z(n30191) );
  NANDN U30551 ( .A(n29933), .B(n29932), .Z(n29937) );
  NANDN U30552 ( .A(n29935), .B(n29934), .Z(n29936) );
  NAND U30553 ( .A(n29937), .B(n29936), .Z(n30428) );
  NANDN U30554 ( .A(n29939), .B(n29938), .Z(n29943) );
  NAND U30555 ( .A(n29941), .B(n29940), .Z(n29942) );
  NAND U30556 ( .A(n29943), .B(n29942), .Z(n30344) );
  NAND U30557 ( .A(n38326), .B(n29944), .Z(n29946) );
  XNOR U30558 ( .A(n38400), .B(a[75]), .Z(n30302) );
  NANDN U30559 ( .A(n38273), .B(n30302), .Z(n29945) );
  NAND U30560 ( .A(n29946), .B(n29945), .Z(n30290) );
  NAND U30561 ( .A(n29948), .B(n29947), .Z(n29951) );
  XNOR U30562 ( .A(n38463), .B(b[7]), .Z(n30376) );
  NAND U30563 ( .A(n30376), .B(n29949), .Z(n29950) );
  NAND U30564 ( .A(n29951), .B(n29950), .Z(n30287) );
  XNOR U30565 ( .A(a[101]), .B(b[33]), .Z(n30241) );
  NANDN U30566 ( .A(n30241), .B(n35620), .Z(n29954) );
  NANDN U30567 ( .A(n29952), .B(n35621), .Z(n29953) );
  AND U30568 ( .A(n29954), .B(n29953), .Z(n30288) );
  XNOR U30569 ( .A(n30287), .B(n30288), .Z(n30289) );
  XOR U30570 ( .A(n30290), .B(n30289), .Z(n30342) );
  XOR U30571 ( .A(b[39]), .B(n35628), .Z(n30299) );
  NANDN U30572 ( .A(n30299), .B(n36553), .Z(n29957) );
  NANDN U30573 ( .A(n29955), .B(n36643), .Z(n29956) );
  NAND U30574 ( .A(n29957), .B(n29956), .Z(n30356) );
  XNOR U30575 ( .A(b[61]), .B(a[73]), .Z(n30207) );
  OR U30576 ( .A(n30207), .B(n38371), .Z(n29960) );
  NANDN U30577 ( .A(n29958), .B(n38369), .Z(n29959) );
  NAND U30578 ( .A(n29960), .B(n29959), .Z(n30353) );
  XOR U30579 ( .A(b[63]), .B(n30543), .Z(n30211) );
  NANDN U30580 ( .A(n30211), .B(n38422), .Z(n29963) );
  NANDN U30581 ( .A(n29961), .B(n38423), .Z(n29962) );
  AND U30582 ( .A(n29963), .B(n29962), .Z(n30354) );
  XNOR U30583 ( .A(n30353), .B(n30354), .Z(n30355) );
  XNOR U30584 ( .A(n30356), .B(n30355), .Z(n30341) );
  XOR U30585 ( .A(n30342), .B(n30341), .Z(n30343) );
  XNOR U30586 ( .A(n30344), .B(n30343), .Z(n30200) );
  NANDN U30587 ( .A(n29965), .B(n29964), .Z(n29969) );
  NAND U30588 ( .A(n29967), .B(n29966), .Z(n29968) );
  NAND U30589 ( .A(n29969), .B(n29968), .Z(n30199) );
  NANDN U30590 ( .A(n29971), .B(n29970), .Z(n29975) );
  NAND U30591 ( .A(n29973), .B(n29972), .Z(n29974) );
  NAND U30592 ( .A(n29975), .B(n29974), .Z(n30277) );
  XNOR U30593 ( .A(a[103]), .B(b[31]), .Z(n30368) );
  NANDN U30594 ( .A(n30368), .B(n35313), .Z(n29978) );
  NANDN U30595 ( .A(n29976), .B(n35311), .Z(n29977) );
  NAND U30596 ( .A(n29978), .B(n29977), .Z(n30223) );
  XNOR U30597 ( .A(a[121]), .B(b[13]), .Z(n30335) );
  OR U30598 ( .A(n30335), .B(n31550), .Z(n29981) );
  NANDN U30599 ( .A(n29979), .B(n31874), .Z(n29980) );
  NAND U30600 ( .A(n29981), .B(n29980), .Z(n30220) );
  XNOR U30601 ( .A(a[123]), .B(b[11]), .Z(n30305) );
  OR U30602 ( .A(n30305), .B(n31369), .Z(n29984) );
  NANDN U30603 ( .A(n29982), .B(n31119), .Z(n29983) );
  AND U30604 ( .A(n29984), .B(n29983), .Z(n30221) );
  XNOR U30605 ( .A(n30220), .B(n30221), .Z(n30222) );
  XNOR U30606 ( .A(n30223), .B(n30222), .Z(n30275) );
  XNOR U30607 ( .A(b[53]), .B(a[81]), .Z(n30244) );
  NANDN U30608 ( .A(n30244), .B(n37940), .Z(n29987) );
  NANDN U30609 ( .A(n29985), .B(n37941), .Z(n29986) );
  NAND U30610 ( .A(n29987), .B(n29986), .Z(n30229) );
  XOR U30611 ( .A(a[117]), .B(b[17]), .Z(n30232) );
  NAND U30612 ( .A(n30232), .B(n32543), .Z(n29990) );
  NAND U30613 ( .A(n29988), .B(n32541), .Z(n29989) );
  NAND U30614 ( .A(n29990), .B(n29989), .Z(n30226) );
  XOR U30615 ( .A(a[119]), .B(n972), .Z(n30235) );
  OR U30616 ( .A(n30235), .B(n32010), .Z(n29993) );
  NANDN U30617 ( .A(n29991), .B(n32011), .Z(n29992) );
  AND U30618 ( .A(n29993), .B(n29992), .Z(n30227) );
  XNOR U30619 ( .A(n30226), .B(n30227), .Z(n30228) );
  XOR U30620 ( .A(n30229), .B(n30228), .Z(n30276) );
  XOR U30621 ( .A(n30275), .B(n30276), .Z(n30278) );
  XOR U30622 ( .A(n30277), .B(n30278), .Z(n30198) );
  XOR U30623 ( .A(n30199), .B(n30198), .Z(n30201) );
  XNOR U30624 ( .A(n30200), .B(n30201), .Z(n30410) );
  OR U30625 ( .A(n29995), .B(n29994), .Z(n29999) );
  OR U30626 ( .A(n29997), .B(n29996), .Z(n29998) );
  NAND U30627 ( .A(n29999), .B(n29998), .Z(n30408) );
  NANDN U30628 ( .A(n30001), .B(n30000), .Z(n30005) );
  NAND U30629 ( .A(n30003), .B(n30002), .Z(n30004) );
  NAND U30630 ( .A(n30005), .B(n30004), .Z(n30284) );
  NAND U30631 ( .A(n34044), .B(n30006), .Z(n30008) );
  XNOR U30632 ( .A(a[111]), .B(n34510), .Z(n30308) );
  NANDN U30633 ( .A(n33867), .B(n30308), .Z(n30007) );
  NAND U30634 ( .A(n30008), .B(n30007), .Z(n30320) );
  XOR U30635 ( .A(b[45]), .B(a[89]), .Z(n30329) );
  NAND U30636 ( .A(n30329), .B(n37261), .Z(n30011) );
  NANDN U30637 ( .A(n30009), .B(n37262), .Z(n30010) );
  NAND U30638 ( .A(n30011), .B(n30010), .Z(n30317) );
  XOR U30639 ( .A(a[109]), .B(b[25]), .Z(n30323) );
  NANDN U30640 ( .A(n34219), .B(n30323), .Z(n30014) );
  NAND U30641 ( .A(n34217), .B(n30012), .Z(n30013) );
  AND U30642 ( .A(n30014), .B(n30013), .Z(n30318) );
  XNOR U30643 ( .A(n30317), .B(n30318), .Z(n30319) );
  XOR U30644 ( .A(n30320), .B(n30319), .Z(n30281) );
  XNOR U30645 ( .A(a[125]), .B(b[9]), .Z(n30380) );
  NANDN U30646 ( .A(n30380), .B(n30509), .Z(n30017) );
  NANDN U30647 ( .A(n30015), .B(n30846), .Z(n30016) );
  NAND U30648 ( .A(n30017), .B(n30016), .Z(n30386) );
  XNOR U30649 ( .A(b[57]), .B(a[77]), .Z(n30332) );
  OR U30650 ( .A(n30332), .B(n965), .Z(n30020) );
  NANDN U30651 ( .A(n30018), .B(n38194), .Z(n30019) );
  NAND U30652 ( .A(n30020), .B(n30019), .Z(n30383) );
  XNOR U30653 ( .A(b[41]), .B(a[93]), .Z(n30204) );
  OR U30654 ( .A(n30204), .B(n36905), .Z(n30023) );
  NANDN U30655 ( .A(n30021), .B(n36807), .Z(n30022) );
  AND U30656 ( .A(n30023), .B(n30022), .Z(n30384) );
  XNOR U30657 ( .A(n30383), .B(n30384), .Z(n30385) );
  XOR U30658 ( .A(n30386), .B(n30385), .Z(n30282) );
  XNOR U30659 ( .A(n30281), .B(n30282), .Z(n30283) );
  XNOR U30660 ( .A(n30284), .B(n30283), .Z(n30350) );
  NANDN U30661 ( .A(n30025), .B(n30024), .Z(n30029) );
  NAND U30662 ( .A(n30027), .B(n30026), .Z(n30028) );
  NAND U30663 ( .A(n30029), .B(n30028), .Z(n30347) );
  NANDN U30664 ( .A(n30031), .B(n30030), .Z(n30035) );
  NAND U30665 ( .A(n30033), .B(n30032), .Z(n30034) );
  AND U30666 ( .A(n30035), .B(n30034), .Z(n30348) );
  XNOR U30667 ( .A(n30347), .B(n30348), .Z(n30349) );
  XOR U30668 ( .A(n30350), .B(n30349), .Z(n30407) );
  XOR U30669 ( .A(n30408), .B(n30407), .Z(n30409) );
  XNOR U30670 ( .A(n30410), .B(n30409), .Z(n30426) );
  OR U30671 ( .A(n30037), .B(n30036), .Z(n30041) );
  OR U30672 ( .A(n30039), .B(n30038), .Z(n30040) );
  NAND U30673 ( .A(n30041), .B(n30040), .Z(n30420) );
  NANDN U30674 ( .A(n30042), .B(b[3]), .Z(n30043) );
  AND U30675 ( .A(n30043), .B(b[5]), .Z(n30214) );
  XNOR U30676 ( .A(b[37]), .B(a[97]), .Z(n30338) );
  NANDN U30677 ( .A(n30338), .B(n36311), .Z(n30046) );
  NANDN U30678 ( .A(n30044), .B(n36309), .Z(n30045) );
  AND U30679 ( .A(n30046), .B(n30045), .Z(n30215) );
  XOR U30680 ( .A(n30214), .B(n30215), .Z(n30216) );
  NANDN U30681 ( .A(n985), .B(a[69]), .Z(n30268) );
  XOR U30682 ( .A(b[35]), .B(a[99]), .Z(n30326) );
  NAND U30683 ( .A(n35985), .B(n30326), .Z(n30049) );
  NANDN U30684 ( .A(n30047), .B(n35986), .Z(n30048) );
  AND U30685 ( .A(n30049), .B(n30048), .Z(n30266) );
  XOR U30686 ( .A(n30265), .B(n30266), .Z(n30267) );
  XOR U30687 ( .A(n30216), .B(n30217), .Z(n30389) );
  NAND U30688 ( .A(n34848), .B(n30050), .Z(n30052) );
  XNOR U30689 ( .A(a[107]), .B(n35375), .Z(n30371) );
  NAND U30690 ( .A(n34618), .B(n30371), .Z(n30051) );
  NAND U30691 ( .A(n30052), .B(n30051), .Z(n30253) );
  NAND U30692 ( .A(n35188), .B(n30053), .Z(n30055) );
  XNOR U30693 ( .A(a[105]), .B(n35540), .Z(n30365) );
  NANDN U30694 ( .A(n34968), .B(n30365), .Z(n30054) );
  NAND U30695 ( .A(n30055), .B(n30054), .Z(n30250) );
  XNOR U30696 ( .A(b[43]), .B(a[91]), .Z(n30238) );
  NANDN U30697 ( .A(n30238), .B(n37068), .Z(n30058) );
  NANDN U30698 ( .A(n30056), .B(n37069), .Z(n30057) );
  AND U30699 ( .A(n30058), .B(n30057), .Z(n30251) );
  XNOR U30700 ( .A(n30250), .B(n30251), .Z(n30252) );
  XOR U30701 ( .A(n30253), .B(n30252), .Z(n30390) );
  XNOR U30702 ( .A(n30389), .B(n30390), .Z(n30392) );
  NANDN U30703 ( .A(n30060), .B(n30059), .Z(n30064) );
  NAND U30704 ( .A(n30062), .B(n30061), .Z(n30063) );
  NAND U30705 ( .A(n30064), .B(n30063), .Z(n30391) );
  XOR U30706 ( .A(n30392), .B(n30391), .Z(n30194) );
  OR U30707 ( .A(n30065), .B(n30265), .Z(n30069) );
  OR U30708 ( .A(n30067), .B(n30066), .Z(n30068) );
  NAND U30709 ( .A(n30069), .B(n30068), .Z(n30193) );
  NANDN U30710 ( .A(n30071), .B(n30070), .Z(n30075) );
  NAND U30711 ( .A(n30073), .B(n30072), .Z(n30074) );
  AND U30712 ( .A(n30075), .B(n30074), .Z(n30192) );
  XNOR U30713 ( .A(n30193), .B(n30192), .Z(n30195) );
  XOR U30714 ( .A(n30194), .B(n30195), .Z(n30419) );
  XNOR U30715 ( .A(n30420), .B(n30419), .Z(n30422) );
  NANDN U30716 ( .A(n30077), .B(n30076), .Z(n30081) );
  NAND U30717 ( .A(n30079), .B(n30078), .Z(n30080) );
  NAND U30718 ( .A(n30081), .B(n30080), .Z(n30271) );
  NAND U30719 ( .A(n33283), .B(n30082), .Z(n30084) );
  XNOR U30720 ( .A(a[115]), .B(n33020), .Z(n30259) );
  NANDN U30721 ( .A(n33021), .B(n30259), .Z(n30083) );
  NAND U30722 ( .A(n30084), .B(n30083), .Z(n30362) );
  XNOR U30723 ( .A(b[51]), .B(a[83]), .Z(n30314) );
  NANDN U30724 ( .A(n30314), .B(n37803), .Z(n30087) );
  NANDN U30725 ( .A(n30085), .B(n37802), .Z(n30086) );
  NAND U30726 ( .A(n30087), .B(n30086), .Z(n30359) );
  XNOR U30727 ( .A(b[55]), .B(a[79]), .Z(n30247) );
  NANDN U30728 ( .A(n30247), .B(n38075), .Z(n30090) );
  NANDN U30729 ( .A(n30088), .B(n38073), .Z(n30089) );
  AND U30730 ( .A(n30090), .B(n30089), .Z(n30360) );
  XNOR U30731 ( .A(n30359), .B(n30360), .Z(n30361) );
  XNOR U30732 ( .A(n30362), .B(n30361), .Z(n30269) );
  XOR U30733 ( .A(a[113]), .B(b[21]), .Z(n30256) );
  NANDN U30734 ( .A(n33634), .B(n30256), .Z(n30093) );
  NANDN U30735 ( .A(n30091), .B(n33464), .Z(n30092) );
  NAND U30736 ( .A(n30093), .B(n30092), .Z(n30296) );
  NAND U30737 ( .A(n37469), .B(n30094), .Z(n30096) );
  XNOR U30738 ( .A(n978), .B(a[87]), .Z(n30262) );
  NAND U30739 ( .A(n30262), .B(n37471), .Z(n30095) );
  NAND U30740 ( .A(n30096), .B(n30095), .Z(n30293) );
  XNOR U30741 ( .A(b[49]), .B(a[85]), .Z(n30311) );
  OR U30742 ( .A(n30311), .B(n37756), .Z(n30099) );
  NANDN U30743 ( .A(n30097), .B(n37652), .Z(n30098) );
  AND U30744 ( .A(n30099), .B(n30098), .Z(n30294) );
  XNOR U30745 ( .A(n30293), .B(n30294), .Z(n30295) );
  XOR U30746 ( .A(n30296), .B(n30295), .Z(n30270) );
  XOR U30747 ( .A(n30269), .B(n30270), .Z(n30272) );
  XOR U30748 ( .A(n30271), .B(n30272), .Z(n30421) );
  XNOR U30749 ( .A(n30422), .B(n30421), .Z(n30425) );
  XOR U30750 ( .A(n30426), .B(n30425), .Z(n30427) );
  XNOR U30751 ( .A(n30428), .B(n30427), .Z(n30189) );
  NANDN U30752 ( .A(n30101), .B(n30100), .Z(n30105) );
  NANDN U30753 ( .A(n30103), .B(n30102), .Z(n30104) );
  NAND U30754 ( .A(n30105), .B(n30104), .Z(n30401) );
  NANDN U30755 ( .A(n30107), .B(n30106), .Z(n30111) );
  NAND U30756 ( .A(n30109), .B(n30108), .Z(n30110) );
  NAND U30757 ( .A(n30111), .B(n30110), .Z(n30414) );
  NANDN U30758 ( .A(n30113), .B(n30112), .Z(n30117) );
  OR U30759 ( .A(n30115), .B(n30114), .Z(n30116) );
  AND U30760 ( .A(n30117), .B(n30116), .Z(n30413) );
  XNOR U30761 ( .A(n30414), .B(n30413), .Z(n30415) );
  NANDN U30762 ( .A(n30119), .B(n30118), .Z(n30123) );
  OR U30763 ( .A(n30121), .B(n30120), .Z(n30122) );
  AND U30764 ( .A(n30123), .B(n30122), .Z(n30416) );
  XOR U30765 ( .A(n30401), .B(n30402), .Z(n30403) );
  OR U30766 ( .A(n30125), .B(n30124), .Z(n30129) );
  NANDN U30767 ( .A(n30127), .B(n30126), .Z(n30128) );
  NAND U30768 ( .A(n30129), .B(n30128), .Z(n30398) );
  NANDN U30769 ( .A(n30131), .B(n30130), .Z(n30135) );
  OR U30770 ( .A(n30133), .B(n30132), .Z(n30134) );
  NAND U30771 ( .A(n30135), .B(n30134), .Z(n30395) );
  NANDN U30772 ( .A(n30137), .B(n30136), .Z(n30141) );
  OR U30773 ( .A(n30139), .B(n30138), .Z(n30140) );
  AND U30774 ( .A(n30141), .B(n30140), .Z(n30396) );
  XNOR U30775 ( .A(n30395), .B(n30396), .Z(n30397) );
  XOR U30776 ( .A(n30398), .B(n30397), .Z(n30404) );
  XOR U30777 ( .A(n30403), .B(n30404), .Z(n30188) );
  XNOR U30778 ( .A(n30189), .B(n30188), .Z(n30190) );
  XNOR U30779 ( .A(n30191), .B(n30190), .Z(n30432) );
  XNOR U30780 ( .A(n30431), .B(n30432), .Z(n30435) );
  XNOR U30781 ( .A(n30436), .B(n30435), .Z(n30438) );
  NANDN U30782 ( .A(n30143), .B(n30142), .Z(n30147) );
  NANDN U30783 ( .A(n30145), .B(n30144), .Z(n30146) );
  NAND U30784 ( .A(n30147), .B(n30146), .Z(n30437) );
  XNOR U30785 ( .A(n30438), .B(n30437), .Z(n30176) );
  NANDN U30786 ( .A(n30149), .B(n30148), .Z(n30153) );
  NANDN U30787 ( .A(n30151), .B(n30150), .Z(n30152) );
  NAND U30788 ( .A(n30153), .B(n30152), .Z(n30177) );
  XNOR U30789 ( .A(n30176), .B(n30177), .Z(n30178) );
  NANDN U30790 ( .A(n30155), .B(n30154), .Z(n30159) );
  NAND U30791 ( .A(n30157), .B(n30156), .Z(n30158) );
  AND U30792 ( .A(n30159), .B(n30158), .Z(n30179) );
  XNOR U30793 ( .A(n30178), .B(n30179), .Z(n30171) );
  NANDN U30794 ( .A(n30161), .B(n30160), .Z(n30165) );
  NAND U30795 ( .A(n30163), .B(n30162), .Z(n30164) );
  AND U30796 ( .A(n30165), .B(n30164), .Z(n30170) );
  XNOR U30797 ( .A(n30171), .B(n30170), .Z(n30173) );
  XOR U30798 ( .A(n30172), .B(n30173), .Z(n30168) );
  OR U30799 ( .A(n30167), .B(n30166), .Z(n30169) );
  XNOR U30800 ( .A(n30168), .B(n30169), .Z(c[197]) );
  NANDN U30801 ( .A(n30169), .B(n30168), .Z(n30443) );
  NANDN U30802 ( .A(n30171), .B(n30170), .Z(n30175) );
  NAND U30803 ( .A(n30173), .B(n30172), .Z(n30174) );
  NAND U30804 ( .A(n30175), .B(n30174), .Z(n30446) );
  NANDN U30805 ( .A(n30177), .B(n30176), .Z(n30181) );
  NAND U30806 ( .A(n30179), .B(n30178), .Z(n30180) );
  AND U30807 ( .A(n30181), .B(n30180), .Z(n30445) );
  NANDN U30808 ( .A(n30183), .B(n30182), .Z(n30187) );
  NANDN U30809 ( .A(n30185), .B(n30184), .Z(n30186) );
  NAND U30810 ( .A(n30187), .B(n30186), .Z(n30699) );
  NANDN U30811 ( .A(n30193), .B(n30192), .Z(n30197) );
  NAND U30812 ( .A(n30195), .B(n30194), .Z(n30196) );
  NAND U30813 ( .A(n30197), .B(n30196), .Z(n30459) );
  NANDN U30814 ( .A(n30199), .B(n30198), .Z(n30203) );
  OR U30815 ( .A(n30201), .B(n30200), .Z(n30202) );
  AND U30816 ( .A(n30203), .B(n30202), .Z(n30460) );
  XNOR U30817 ( .A(n30459), .B(n30460), .Z(n30461) );
  XNOR U30818 ( .A(b[41]), .B(a[94]), .Z(n30503) );
  OR U30819 ( .A(n30503), .B(n36905), .Z(n30206) );
  NANDN U30820 ( .A(n30204), .B(n36807), .Z(n30205) );
  NAND U30821 ( .A(n30206), .B(n30205), .Z(n30494) );
  XOR U30822 ( .A(b[61]), .B(n31372), .Z(n30574) );
  OR U30823 ( .A(n30574), .B(n38371), .Z(n30209) );
  NANDN U30824 ( .A(n30207), .B(n38369), .Z(n30208) );
  NAND U30825 ( .A(n30209), .B(n30208), .Z(n30491) );
  XOR U30826 ( .A(b[63]), .B(n30210), .Z(n30534) );
  NANDN U30827 ( .A(n30534), .B(n38422), .Z(n30213) );
  NANDN U30828 ( .A(n30211), .B(n38423), .Z(n30212) );
  AND U30829 ( .A(n30213), .B(n30212), .Z(n30492) );
  XNOR U30830 ( .A(n30491), .B(n30492), .Z(n30493) );
  XNOR U30831 ( .A(n30494), .B(n30493), .Z(n30607) );
  OR U30832 ( .A(n30215), .B(n30214), .Z(n30219) );
  NAND U30833 ( .A(n30217), .B(n30216), .Z(n30218) );
  NAND U30834 ( .A(n30219), .B(n30218), .Z(n30605) );
  NANDN U30835 ( .A(n30221), .B(n30220), .Z(n30225) );
  NAND U30836 ( .A(n30223), .B(n30222), .Z(n30224) );
  AND U30837 ( .A(n30225), .B(n30224), .Z(n30604) );
  XNOR U30838 ( .A(n30605), .B(n30604), .Z(n30606) );
  XOR U30839 ( .A(n30607), .B(n30606), .Z(n30663) );
  NANDN U30840 ( .A(n30227), .B(n30226), .Z(n30231) );
  NAND U30841 ( .A(n30229), .B(n30228), .Z(n30230) );
  NAND U30842 ( .A(n30231), .B(n30230), .Z(n30487) );
  XNOR U30843 ( .A(a[118]), .B(b[17]), .Z(n30513) );
  NANDN U30844 ( .A(n30513), .B(n32543), .Z(n30234) );
  NAND U30845 ( .A(n30232), .B(n32541), .Z(n30233) );
  NAND U30846 ( .A(n30234), .B(n30233), .Z(n30595) );
  XOR U30847 ( .A(a[120]), .B(n972), .Z(n30643) );
  OR U30848 ( .A(n30643), .B(n32010), .Z(n30237) );
  NANDN U30849 ( .A(n30235), .B(n32011), .Z(n30236) );
  NAND U30850 ( .A(n30237), .B(n30236), .Z(n30592) );
  XOR U30851 ( .A(b[43]), .B(n34852), .Z(n30637) );
  NANDN U30852 ( .A(n30637), .B(n37068), .Z(n30240) );
  NANDN U30853 ( .A(n30238), .B(n37069), .Z(n30239) );
  AND U30854 ( .A(n30240), .B(n30239), .Z(n30593) );
  XNOR U30855 ( .A(n30592), .B(n30593), .Z(n30594) );
  XNOR U30856 ( .A(n30595), .B(n30594), .Z(n30485) );
  XOR U30857 ( .A(a[102]), .B(n974), .Z(n30583) );
  NANDN U30858 ( .A(n30583), .B(n35620), .Z(n30243) );
  NANDN U30859 ( .A(n30241), .B(n35621), .Z(n30242) );
  NAND U30860 ( .A(n30243), .B(n30242), .Z(n30556) );
  XOR U30861 ( .A(b[53]), .B(n32815), .Z(n30631) );
  NANDN U30862 ( .A(n30631), .B(n37940), .Z(n30246) );
  NANDN U30863 ( .A(n30244), .B(n37941), .Z(n30245) );
  NAND U30864 ( .A(n30246), .B(n30245), .Z(n30553) );
  XOR U30865 ( .A(b[55]), .B(n32814), .Z(n30634) );
  NANDN U30866 ( .A(n30634), .B(n38075), .Z(n30249) );
  NANDN U30867 ( .A(n30247), .B(n38073), .Z(n30248) );
  AND U30868 ( .A(n30249), .B(n30248), .Z(n30554) );
  XNOR U30869 ( .A(n30553), .B(n30554), .Z(n30555) );
  XOR U30870 ( .A(n30556), .B(n30555), .Z(n30486) );
  XOR U30871 ( .A(n30485), .B(n30486), .Z(n30488) );
  XOR U30872 ( .A(n30487), .B(n30488), .Z(n30661) );
  NANDN U30873 ( .A(n30251), .B(n30250), .Z(n30255) );
  NAND U30874 ( .A(n30253), .B(n30252), .Z(n30254) );
  NAND U30875 ( .A(n30255), .B(n30254), .Z(n30600) );
  XNOR U30876 ( .A(a[114]), .B(b[21]), .Z(n30625) );
  OR U30877 ( .A(n30625), .B(n33634), .Z(n30258) );
  NAND U30878 ( .A(n30256), .B(n33464), .Z(n30257) );
  NAND U30879 ( .A(n30258), .B(n30257), .Z(n30525) );
  NAND U30880 ( .A(n33283), .B(n30259), .Z(n30261) );
  XOR U30881 ( .A(n38046), .B(n33020), .Z(n30544) );
  NANDN U30882 ( .A(n33021), .B(n30544), .Z(n30260) );
  NAND U30883 ( .A(n30261), .B(n30260), .Z(n30522) );
  NAND U30884 ( .A(n37469), .B(n30262), .Z(n30264) );
  XOR U30885 ( .A(n978), .B(n34048), .Z(n30516) );
  NAND U30886 ( .A(n30516), .B(n37471), .Z(n30263) );
  AND U30887 ( .A(n30264), .B(n30263), .Z(n30523) );
  XNOR U30888 ( .A(n30522), .B(n30523), .Z(n30524) );
  XNOR U30889 ( .A(n30525), .B(n30524), .Z(n30598) );
  XOR U30890 ( .A(n30598), .B(n30599), .Z(n30601) );
  XNOR U30891 ( .A(n30600), .B(n30601), .Z(n30660) );
  XOR U30892 ( .A(n30661), .B(n30660), .Z(n30662) );
  XOR U30893 ( .A(n30663), .B(n30662), .Z(n30468) );
  NANDN U30894 ( .A(n30270), .B(n30269), .Z(n30274) );
  OR U30895 ( .A(n30272), .B(n30271), .Z(n30273) );
  NAND U30896 ( .A(n30274), .B(n30273), .Z(n30465) );
  NANDN U30897 ( .A(n30276), .B(n30275), .Z(n30280) );
  OR U30898 ( .A(n30278), .B(n30277), .Z(n30279) );
  AND U30899 ( .A(n30280), .B(n30279), .Z(n30466) );
  XNOR U30900 ( .A(n30465), .B(n30466), .Z(n30467) );
  XOR U30901 ( .A(n30468), .B(n30467), .Z(n30462) );
  XOR U30902 ( .A(n30461), .B(n30462), .Z(n30453) );
  OR U30903 ( .A(n30282), .B(n30281), .Z(n30286) );
  OR U30904 ( .A(n30284), .B(n30283), .Z(n30285) );
  NAND U30905 ( .A(n30286), .B(n30285), .Z(n30669) );
  NANDN U30906 ( .A(n30288), .B(n30287), .Z(n30292) );
  NAND U30907 ( .A(n30290), .B(n30289), .Z(n30291) );
  NAND U30908 ( .A(n30292), .B(n30291), .Z(n30472) );
  NANDN U30909 ( .A(n30294), .B(n30293), .Z(n30298) );
  NAND U30910 ( .A(n30296), .B(n30295), .Z(n30297) );
  NAND U30911 ( .A(n30298), .B(n30297), .Z(n30481) );
  XOR U30912 ( .A(b[39]), .B(n35545), .Z(n30537) );
  NANDN U30913 ( .A(n30537), .B(n36553), .Z(n30301) );
  NANDN U30914 ( .A(n30299), .B(n36643), .Z(n30300) );
  NAND U30915 ( .A(n30301), .B(n30300), .Z(n30568) );
  NAND U30916 ( .A(n38326), .B(n30302), .Z(n30304) );
  XOR U30917 ( .A(n38400), .B(n31363), .Z(n30506) );
  NANDN U30918 ( .A(n38273), .B(n30506), .Z(n30303) );
  NAND U30919 ( .A(n30304), .B(n30303), .Z(n30565) );
  XOR U30920 ( .A(a[124]), .B(n970), .Z(n30580) );
  OR U30921 ( .A(n30580), .B(n31369), .Z(n30307) );
  NANDN U30922 ( .A(n30305), .B(n31119), .Z(n30306) );
  AND U30923 ( .A(n30307), .B(n30306), .Z(n30566) );
  XNOR U30924 ( .A(n30565), .B(n30566), .Z(n30567) );
  XNOR U30925 ( .A(n30568), .B(n30567), .Z(n30479) );
  NAND U30926 ( .A(n34044), .B(n30308), .Z(n30310) );
  XOR U30927 ( .A(a[112]), .B(n34510), .Z(n30628) );
  OR U30928 ( .A(n30628), .B(n33867), .Z(n30309) );
  NAND U30929 ( .A(n30310), .B(n30309), .Z(n30589) );
  XOR U30930 ( .A(b[49]), .B(n33628), .Z(n30519) );
  OR U30931 ( .A(n30519), .B(n37756), .Z(n30313) );
  NANDN U30932 ( .A(n30311), .B(n37652), .Z(n30312) );
  NAND U30933 ( .A(n30313), .B(n30312), .Z(n30586) );
  XOR U30934 ( .A(b[51]), .B(n33185), .Z(n30640) );
  NANDN U30935 ( .A(n30640), .B(n37803), .Z(n30316) );
  NANDN U30936 ( .A(n30314), .B(n37802), .Z(n30315) );
  AND U30937 ( .A(n30316), .B(n30315), .Z(n30587) );
  XNOR U30938 ( .A(n30586), .B(n30587), .Z(n30588) );
  XOR U30939 ( .A(n30589), .B(n30588), .Z(n30480) );
  XOR U30940 ( .A(n30479), .B(n30480), .Z(n30482) );
  XOR U30941 ( .A(n30481), .B(n30482), .Z(n30471) );
  XNOR U30942 ( .A(n30472), .B(n30471), .Z(n30473) );
  NANDN U30943 ( .A(n30318), .B(n30317), .Z(n30322) );
  NAND U30944 ( .A(n30320), .B(n30319), .Z(n30321) );
  NAND U30945 ( .A(n30322), .B(n30321), .Z(n30561) );
  XNOR U30946 ( .A(n37336), .B(b[25]), .Z(n30616) );
  NANDN U30947 ( .A(n34219), .B(n30616), .Z(n30325) );
  NAND U30948 ( .A(n34217), .B(n30323), .Z(n30324) );
  NAND U30949 ( .A(n30325), .B(n30324), .Z(n30500) );
  XNOR U30950 ( .A(b[35]), .B(n36100), .Z(n30571) );
  NAND U30951 ( .A(n35985), .B(n30571), .Z(n30328) );
  NAND U30952 ( .A(n30326), .B(n35986), .Z(n30327) );
  NAND U30953 ( .A(n30328), .B(n30327), .Z(n30497) );
  XNOR U30954 ( .A(b[45]), .B(a[90]), .Z(n30550) );
  NANDN U30955 ( .A(n30550), .B(n37261), .Z(n30331) );
  NAND U30956 ( .A(n30329), .B(n37262), .Z(n30330) );
  AND U30957 ( .A(n30331), .B(n30330), .Z(n30498) );
  XNOR U30958 ( .A(n30497), .B(n30498), .Z(n30499) );
  XNOR U30959 ( .A(n30500), .B(n30499), .Z(n30559) );
  XOR U30960 ( .A(b[57]), .B(n31870), .Z(n30577) );
  OR U30961 ( .A(n30577), .B(n965), .Z(n30334) );
  NANDN U30962 ( .A(n30332), .B(n38194), .Z(n30333) );
  NAND U30963 ( .A(n30334), .B(n30333), .Z(n30531) );
  XOR U30964 ( .A(a[122]), .B(n971), .Z(n30646) );
  OR U30965 ( .A(n30646), .B(n31550), .Z(n30337) );
  NANDN U30966 ( .A(n30335), .B(n31874), .Z(n30336) );
  NAND U30967 ( .A(n30337), .B(n30336), .Z(n30528) );
  XOR U30968 ( .A(b[37]), .B(n35783), .Z(n30540) );
  NANDN U30969 ( .A(n30540), .B(n36311), .Z(n30340) );
  NANDN U30970 ( .A(n30338), .B(n36309), .Z(n30339) );
  AND U30971 ( .A(n30340), .B(n30339), .Z(n30529) );
  XNOR U30972 ( .A(n30528), .B(n30529), .Z(n30530) );
  XOR U30973 ( .A(n30531), .B(n30530), .Z(n30560) );
  XOR U30974 ( .A(n30559), .B(n30560), .Z(n30562) );
  XOR U30975 ( .A(n30561), .B(n30562), .Z(n30474) );
  XOR U30976 ( .A(n30473), .B(n30474), .Z(n30666) );
  NANDN U30977 ( .A(n30342), .B(n30341), .Z(n30346) );
  OR U30978 ( .A(n30344), .B(n30343), .Z(n30345) );
  NAND U30979 ( .A(n30346), .B(n30345), .Z(n30667) );
  XOR U30980 ( .A(n30666), .B(n30667), .Z(n30668) );
  XNOR U30981 ( .A(n30669), .B(n30668), .Z(n30679) );
  NANDN U30982 ( .A(n30348), .B(n30347), .Z(n30352) );
  NAND U30983 ( .A(n30350), .B(n30349), .Z(n30351) );
  NAND U30984 ( .A(n30352), .B(n30351), .Z(n30674) );
  NANDN U30985 ( .A(n30354), .B(n30353), .Z(n30358) );
  NAND U30986 ( .A(n30356), .B(n30355), .Z(n30357) );
  NAND U30987 ( .A(n30358), .B(n30357), .Z(n30478) );
  NANDN U30988 ( .A(n30360), .B(n30359), .Z(n30364) );
  NAND U30989 ( .A(n30362), .B(n30361), .Z(n30363) );
  NAND U30990 ( .A(n30364), .B(n30363), .Z(n30613) );
  NAND U30991 ( .A(n35188), .B(n30365), .Z(n30367) );
  XOR U30992 ( .A(n36909), .B(n35540), .Z(n30622) );
  NANDN U30993 ( .A(n34968), .B(n30622), .Z(n30366) );
  NAND U30994 ( .A(n30367), .B(n30366), .Z(n30652) );
  XOR U30995 ( .A(a[104]), .B(n973), .Z(n30547) );
  NANDN U30996 ( .A(n30547), .B(n35313), .Z(n30370) );
  NANDN U30997 ( .A(n30368), .B(n35311), .Z(n30369) );
  NAND U30998 ( .A(n30370), .B(n30369), .Z(n30649) );
  NAND U30999 ( .A(n34848), .B(n30371), .Z(n30373) );
  XOR U31000 ( .A(n37139), .B(n35375), .Z(n30619) );
  NAND U31001 ( .A(n34618), .B(n30619), .Z(n30372) );
  AND U31002 ( .A(n30373), .B(n30372), .Z(n30650) );
  XNOR U31003 ( .A(n30649), .B(n30650), .Z(n30651) );
  XOR U31004 ( .A(n30652), .B(n30651), .Z(n30610) );
  XOR U31005 ( .A(n31123), .B(n30374), .Z(n30378) );
  XOR U31006 ( .A(n968), .B(b[6]), .Z(n30375) );
  NANDN U31007 ( .A(n30376), .B(n30375), .Z(n30377) );
  AND U31008 ( .A(n30378), .B(n30377), .Z(n30656) );
  ANDN U31009 ( .B(b[63]), .A(n30379), .Z(n30942) );
  XOR U31010 ( .A(a[126]), .B(n969), .Z(n30510) );
  NANDN U31011 ( .A(n30510), .B(n30509), .Z(n30382) );
  NANDN U31012 ( .A(n30380), .B(n30846), .Z(n30381) );
  AND U31013 ( .A(n30382), .B(n30381), .Z(n30655) );
  XNOR U31014 ( .A(n30942), .B(n30655), .Z(n30657) );
  XNOR U31015 ( .A(n30656), .B(n30657), .Z(n30611) );
  XNOR U31016 ( .A(n30610), .B(n30611), .Z(n30612) );
  XNOR U31017 ( .A(n30613), .B(n30612), .Z(n30475) );
  NANDN U31018 ( .A(n30384), .B(n30383), .Z(n30388) );
  NAND U31019 ( .A(n30386), .B(n30385), .Z(n30387) );
  AND U31020 ( .A(n30388), .B(n30387), .Z(n30476) );
  XNOR U31021 ( .A(n30475), .B(n30476), .Z(n30477) );
  XNOR U31022 ( .A(n30478), .B(n30477), .Z(n30672) );
  OR U31023 ( .A(n30390), .B(n30389), .Z(n30394) );
  OR U31024 ( .A(n30392), .B(n30391), .Z(n30393) );
  AND U31025 ( .A(n30394), .B(n30393), .Z(n30673) );
  XOR U31026 ( .A(n30672), .B(n30673), .Z(n30675) );
  XOR U31027 ( .A(n30674), .B(n30675), .Z(n30678) );
  XOR U31028 ( .A(n30679), .B(n30678), .Z(n30681) );
  NANDN U31029 ( .A(n30396), .B(n30395), .Z(n30400) );
  NAND U31030 ( .A(n30398), .B(n30397), .Z(n30399) );
  AND U31031 ( .A(n30400), .B(n30399), .Z(n30680) );
  XOR U31032 ( .A(n30681), .B(n30680), .Z(n30454) );
  XNOR U31033 ( .A(n30453), .B(n30454), .Z(n30455) );
  OR U31034 ( .A(n30402), .B(n30401), .Z(n30406) );
  NAND U31035 ( .A(n30404), .B(n30403), .Z(n30405) );
  NAND U31036 ( .A(n30406), .B(n30405), .Z(n30456) );
  XOR U31037 ( .A(n30455), .B(n30456), .Z(n30693) );
  NAND U31038 ( .A(n30408), .B(n30407), .Z(n30412) );
  NAND U31039 ( .A(n30410), .B(n30409), .Z(n30411) );
  NAND U31040 ( .A(n30412), .B(n30411), .Z(n30684) );
  OR U31041 ( .A(n30414), .B(n30413), .Z(n30418) );
  OR U31042 ( .A(n30416), .B(n30415), .Z(n30417) );
  NAND U31043 ( .A(n30418), .B(n30417), .Z(n30685) );
  XNOR U31044 ( .A(n30684), .B(n30685), .Z(n30686) );
  NAND U31045 ( .A(n30420), .B(n30419), .Z(n30424) );
  NANDN U31046 ( .A(n30422), .B(n30421), .Z(n30423) );
  NAND U31047 ( .A(n30424), .B(n30423), .Z(n30687) );
  XOR U31048 ( .A(n30686), .B(n30687), .Z(n30690) );
  XNOR U31049 ( .A(n30690), .B(n30691), .Z(n30692) );
  XNOR U31050 ( .A(n30693), .B(n30692), .Z(n30697) );
  XNOR U31051 ( .A(n30696), .B(n30697), .Z(n30698) );
  XNOR U31052 ( .A(n30699), .B(n30698), .Z(n30447) );
  OR U31053 ( .A(n30430), .B(n30429), .Z(n30434) );
  NANDN U31054 ( .A(n30432), .B(n30431), .Z(n30433) );
  NAND U31055 ( .A(n30434), .B(n30433), .Z(n30448) );
  XOR U31056 ( .A(n30447), .B(n30448), .Z(n30450) );
  NAND U31057 ( .A(n30436), .B(n30435), .Z(n30440) );
  OR U31058 ( .A(n30438), .B(n30437), .Z(n30439) );
  NAND U31059 ( .A(n30440), .B(n30439), .Z(n30449) );
  XOR U31060 ( .A(n30450), .B(n30449), .Z(n30444) );
  XNOR U31061 ( .A(n30445), .B(n30444), .Z(n30441) );
  XOR U31062 ( .A(n30446), .B(n30441), .Z(n30442) );
  XNOR U31063 ( .A(n30443), .B(n30442), .Z(c[198]) );
  NANDN U31064 ( .A(n30443), .B(n30442), .Z(n30963) );
  NANDN U31065 ( .A(n30448), .B(n30447), .Z(n30452) );
  OR U31066 ( .A(n30450), .B(n30449), .Z(n30451) );
  NAND U31067 ( .A(n30452), .B(n30451), .Z(n30706) );
  NANDN U31068 ( .A(n30454), .B(n30453), .Z(n30458) );
  NANDN U31069 ( .A(n30456), .B(n30455), .Z(n30457) );
  NAND U31070 ( .A(n30458), .B(n30457), .Z(n30716) );
  NANDN U31071 ( .A(n30460), .B(n30459), .Z(n30464) );
  NANDN U31072 ( .A(n30462), .B(n30461), .Z(n30463) );
  NAND U31073 ( .A(n30464), .B(n30463), .Z(n30730) );
  NANDN U31074 ( .A(n30466), .B(n30465), .Z(n30470) );
  NANDN U31075 ( .A(n30468), .B(n30467), .Z(n30469) );
  NAND U31076 ( .A(n30470), .B(n30469), .Z(n30741) );
  NANDN U31077 ( .A(n30480), .B(n30479), .Z(n30484) );
  OR U31078 ( .A(n30482), .B(n30481), .Z(n30483) );
  NAND U31079 ( .A(n30484), .B(n30483), .Z(n30791) );
  NANDN U31080 ( .A(n30486), .B(n30485), .Z(n30490) );
  OR U31081 ( .A(n30488), .B(n30487), .Z(n30489) );
  AND U31082 ( .A(n30490), .B(n30489), .Z(n30792) );
  XNOR U31083 ( .A(n30791), .B(n30792), .Z(n30793) );
  XNOR U31084 ( .A(n30794), .B(n30793), .Z(n30739) );
  XNOR U31085 ( .A(n30740), .B(n30739), .Z(n30742) );
  XNOR U31086 ( .A(n30741), .B(n30742), .Z(n30727) );
  NANDN U31087 ( .A(n30492), .B(n30491), .Z(n30496) );
  NAND U31088 ( .A(n30494), .B(n30493), .Z(n30495) );
  NAND U31089 ( .A(n30496), .B(n30495), .Z(n30812) );
  NANDN U31090 ( .A(n30498), .B(n30497), .Z(n30502) );
  NAND U31091 ( .A(n30500), .B(n30499), .Z(n30501) );
  NAND U31092 ( .A(n30502), .B(n30501), .Z(n30787) );
  XNOR U31093 ( .A(b[41]), .B(a[95]), .Z(n30907) );
  OR U31094 ( .A(n30907), .B(n36905), .Z(n30505) );
  NANDN U31095 ( .A(n30503), .B(n36807), .Z(n30504) );
  NAND U31096 ( .A(n30505), .B(n30504), .Z(n30892) );
  NAND U31097 ( .A(n38326), .B(n30506), .Z(n30508) );
  XNOR U31098 ( .A(n38400), .B(a[77]), .Z(n30910) );
  NANDN U31099 ( .A(n38273), .B(n30910), .Z(n30507) );
  NAND U31100 ( .A(n30508), .B(n30507), .Z(n30889) );
  XOR U31101 ( .A(a[127]), .B(n969), .Z(n30847) );
  NANDN U31102 ( .A(n30847), .B(n30509), .Z(n30512) );
  NANDN U31103 ( .A(n30510), .B(n30846), .Z(n30511) );
  AND U31104 ( .A(n30512), .B(n30511), .Z(n30890) );
  XNOR U31105 ( .A(n30889), .B(n30890), .Z(n30891) );
  XNOR U31106 ( .A(n30892), .B(n30891), .Z(n30785) );
  XNOR U31107 ( .A(a[119]), .B(b[17]), .Z(n30830) );
  NANDN U31108 ( .A(n30830), .B(n32543), .Z(n30515) );
  NANDN U31109 ( .A(n30513), .B(n32541), .Z(n30514) );
  NAND U31110 ( .A(n30515), .B(n30514), .Z(n30947) );
  NAND U31111 ( .A(n37469), .B(n30516), .Z(n30518) );
  XNOR U31112 ( .A(b[47]), .B(a[89]), .Z(n30856) );
  NANDN U31113 ( .A(n30856), .B(n37471), .Z(n30517) );
  NAND U31114 ( .A(n30518), .B(n30517), .Z(n30944) );
  XNOR U31115 ( .A(b[49]), .B(a[87]), .Z(n30934) );
  OR U31116 ( .A(n30934), .B(n37756), .Z(n30521) );
  NANDN U31117 ( .A(n30519), .B(n37652), .Z(n30520) );
  AND U31118 ( .A(n30521), .B(n30520), .Z(n30945) );
  XNOR U31119 ( .A(n30944), .B(n30945), .Z(n30946) );
  XOR U31120 ( .A(n30947), .B(n30946), .Z(n30786) );
  XOR U31121 ( .A(n30785), .B(n30786), .Z(n30788) );
  XNOR U31122 ( .A(n30787), .B(n30788), .Z(n30809) );
  NANDN U31123 ( .A(n30523), .B(n30522), .Z(n30527) );
  NAND U31124 ( .A(n30525), .B(n30524), .Z(n30526) );
  AND U31125 ( .A(n30527), .B(n30526), .Z(n30810) );
  XNOR U31126 ( .A(n30809), .B(n30810), .Z(n30811) );
  XNOR U31127 ( .A(n30812), .B(n30811), .Z(n30880) );
  NANDN U31128 ( .A(n30529), .B(n30528), .Z(n30533) );
  NAND U31129 ( .A(n30531), .B(n30530), .Z(n30532) );
  NAND U31130 ( .A(n30533), .B(n30532), .Z(n30877) );
  XNOR U31131 ( .A(b[63]), .B(a[73]), .Z(n30843) );
  NANDN U31132 ( .A(n30843), .B(n38422), .Z(n30536) );
  NANDN U31133 ( .A(n30534), .B(n38423), .Z(n30535) );
  NAND U31134 ( .A(n30536), .B(n30535), .Z(n30850) );
  XNOR U31135 ( .A(b[39]), .B(a[97]), .Z(n30770) );
  NANDN U31136 ( .A(n30770), .B(n36553), .Z(n30539) );
  NANDN U31137 ( .A(n30537), .B(n36643), .Z(n30538) );
  AND U31138 ( .A(n30539), .B(n30538), .Z(n30851) );
  XNOR U31139 ( .A(n30850), .B(n30851), .Z(n30852) );
  NANDN U31140 ( .A(n30540), .B(n36309), .Z(n30542) );
  XNOR U31141 ( .A(n975), .B(a[99]), .Z(n30859) );
  NAND U31142 ( .A(n30859), .B(n36311), .Z(n30541) );
  AND U31143 ( .A(n30542), .B(n30541), .Z(n30941) );
  ANDN U31144 ( .B(b[63]), .A(n30543), .Z(n30940) );
  XOR U31145 ( .A(n30941), .B(n30940), .Z(n30943) );
  XOR U31146 ( .A(n30942), .B(n30943), .Z(n30853) );
  XOR U31147 ( .A(n30852), .B(n30853), .Z(n30842) );
  NAND U31148 ( .A(n33283), .B(n30544), .Z(n30546) );
  XNOR U31149 ( .A(a[117]), .B(n33020), .Z(n30919) );
  NANDN U31150 ( .A(n33021), .B(n30919), .Z(n30545) );
  NAND U31151 ( .A(n30546), .B(n30545), .Z(n30928) );
  XNOR U31152 ( .A(a[105]), .B(b[31]), .Z(n30862) );
  NANDN U31153 ( .A(n30862), .B(n35313), .Z(n30549) );
  NANDN U31154 ( .A(n30547), .B(n35311), .Z(n30548) );
  NAND U31155 ( .A(n30549), .B(n30548), .Z(n30925) );
  XOR U31156 ( .A(b[45]), .B(a[91]), .Z(n30922) );
  NAND U31157 ( .A(n30922), .B(n37261), .Z(n30552) );
  NANDN U31158 ( .A(n30550), .B(n37262), .Z(n30551) );
  AND U31159 ( .A(n30552), .B(n30551), .Z(n30926) );
  XNOR U31160 ( .A(n30925), .B(n30926), .Z(n30927) );
  XNOR U31161 ( .A(n30928), .B(n30927), .Z(n30839) );
  NANDN U31162 ( .A(n30554), .B(n30553), .Z(n30558) );
  NAND U31163 ( .A(n30556), .B(n30555), .Z(n30557) );
  NAND U31164 ( .A(n30558), .B(n30557), .Z(n30840) );
  XNOR U31165 ( .A(n30839), .B(n30840), .Z(n30841) );
  XNOR U31166 ( .A(n30842), .B(n30841), .Z(n30878) );
  XOR U31167 ( .A(n30877), .B(n30878), .Z(n30879) );
  XOR U31168 ( .A(n30880), .B(n30879), .Z(n30806) );
  NANDN U31169 ( .A(n30560), .B(n30559), .Z(n30564) );
  OR U31170 ( .A(n30562), .B(n30561), .Z(n30563) );
  NAND U31171 ( .A(n30564), .B(n30563), .Z(n30803) );
  NANDN U31172 ( .A(n30566), .B(n30565), .Z(n30570) );
  NAND U31173 ( .A(n30568), .B(n30567), .Z(n30569) );
  NAND U31174 ( .A(n30570), .B(n30569), .Z(n30748) );
  NAND U31175 ( .A(n35986), .B(n30571), .Z(n30573) );
  XNOR U31176 ( .A(b[35]), .B(a[101]), .Z(n30868) );
  NANDN U31177 ( .A(n30868), .B(n35985), .Z(n30572) );
  NAND U31178 ( .A(n30573), .B(n30572), .Z(n30750) );
  NANDN U31179 ( .A(n30574), .B(n38369), .Z(n30576) );
  XNOR U31180 ( .A(n984), .B(a[75]), .Z(n30776) );
  NANDN U31181 ( .A(n38371), .B(n30776), .Z(n30575) );
  AND U31182 ( .A(n30576), .B(n30575), .Z(n30749) );
  XNOR U31183 ( .A(n30750), .B(n30749), .Z(n30752) );
  XNOR U31184 ( .A(n30751), .B(n30752), .Z(n30886) );
  XNOR U31185 ( .A(b[57]), .B(a[79]), .Z(n30761) );
  OR U31186 ( .A(n30761), .B(n965), .Z(n30579) );
  NANDN U31187 ( .A(n30577), .B(n38194), .Z(n30578) );
  NAND U31188 ( .A(n30579), .B(n30578), .Z(n30904) );
  XNOR U31189 ( .A(a[125]), .B(b[11]), .Z(n30773) );
  OR U31190 ( .A(n30773), .B(n31369), .Z(n30582) );
  NANDN U31191 ( .A(n30580), .B(n31119), .Z(n30581) );
  NAND U31192 ( .A(n30582), .B(n30581), .Z(n30901) );
  XNOR U31193 ( .A(a[103]), .B(b[33]), .Z(n30865) );
  NANDN U31194 ( .A(n30865), .B(n35620), .Z(n30585) );
  NANDN U31195 ( .A(n30583), .B(n35621), .Z(n30584) );
  AND U31196 ( .A(n30585), .B(n30584), .Z(n30902) );
  XNOR U31197 ( .A(n30901), .B(n30902), .Z(n30903) );
  XOR U31198 ( .A(n30904), .B(n30903), .Z(n30883) );
  NANDN U31199 ( .A(n30587), .B(n30586), .Z(n30591) );
  NAND U31200 ( .A(n30589), .B(n30588), .Z(n30590) );
  NAND U31201 ( .A(n30591), .B(n30590), .Z(n30884) );
  XNOR U31202 ( .A(n30883), .B(n30884), .Z(n30885) );
  XNOR U31203 ( .A(n30886), .B(n30885), .Z(n30745) );
  NANDN U31204 ( .A(n30593), .B(n30592), .Z(n30597) );
  NAND U31205 ( .A(n30595), .B(n30594), .Z(n30596) );
  AND U31206 ( .A(n30597), .B(n30596), .Z(n30746) );
  XNOR U31207 ( .A(n30745), .B(n30746), .Z(n30747) );
  XNOR U31208 ( .A(n30748), .B(n30747), .Z(n30804) );
  XOR U31209 ( .A(n30803), .B(n30804), .Z(n30805) );
  XNOR U31210 ( .A(n30806), .B(n30805), .Z(n30736) );
  NANDN U31211 ( .A(n30599), .B(n30598), .Z(n30603) );
  OR U31212 ( .A(n30601), .B(n30600), .Z(n30602) );
  NAND U31213 ( .A(n30603), .B(n30602), .Z(n30733) );
  NANDN U31214 ( .A(n30605), .B(n30604), .Z(n30609) );
  NAND U31215 ( .A(n30607), .B(n30606), .Z(n30608) );
  NAND U31216 ( .A(n30609), .B(n30608), .Z(n30800) );
  OR U31217 ( .A(n30611), .B(n30610), .Z(n30615) );
  OR U31218 ( .A(n30613), .B(n30612), .Z(n30614) );
  NAND U31219 ( .A(n30615), .B(n30614), .Z(n30797) );
  XOR U31220 ( .A(a[111]), .B(b[25]), .Z(n30764) );
  NANDN U31221 ( .A(n34219), .B(n30764), .Z(n30618) );
  NAND U31222 ( .A(n34217), .B(n30616), .Z(n30617) );
  NAND U31223 ( .A(n30618), .B(n30617), .Z(n30818) );
  NAND U31224 ( .A(n34848), .B(n30619), .Z(n30621) );
  XNOR U31225 ( .A(a[109]), .B(n35375), .Z(n30821) );
  NAND U31226 ( .A(n34618), .B(n30821), .Z(n30620) );
  NAND U31227 ( .A(n30621), .B(n30620), .Z(n30815) );
  NAND U31228 ( .A(n35188), .B(n30622), .Z(n30624) );
  XNOR U31229 ( .A(a[107]), .B(n35540), .Z(n30931) );
  NANDN U31230 ( .A(n34968), .B(n30931), .Z(n30623) );
  AND U31231 ( .A(n30624), .B(n30623), .Z(n30816) );
  XNOR U31232 ( .A(n30815), .B(n30816), .Z(n30817) );
  XNOR U31233 ( .A(n30818), .B(n30817), .Z(n30898) );
  XOR U31234 ( .A(a[115]), .B(b[21]), .Z(n30916) );
  NANDN U31235 ( .A(n33634), .B(n30916), .Z(n30627) );
  NANDN U31236 ( .A(n30625), .B(n33464), .Z(n30626) );
  NAND U31237 ( .A(n30627), .B(n30626), .Z(n30896) );
  NANDN U31238 ( .A(n30628), .B(n34044), .Z(n30630) );
  XNOR U31239 ( .A(a[113]), .B(n34510), .Z(n30767) );
  NANDN U31240 ( .A(n33867), .B(n30767), .Z(n30629) );
  AND U31241 ( .A(n30630), .B(n30629), .Z(n30895) );
  XNOR U31242 ( .A(n30896), .B(n30895), .Z(n30897) );
  XOR U31243 ( .A(n30898), .B(n30897), .Z(n30952) );
  XNOR U31244 ( .A(b[53]), .B(a[83]), .Z(n30824) );
  NANDN U31245 ( .A(n30824), .B(n37940), .Z(n30633) );
  NANDN U31246 ( .A(n30631), .B(n37941), .Z(n30632) );
  NAND U31247 ( .A(n30633), .B(n30632), .Z(n30782) );
  XNOR U31248 ( .A(b[55]), .B(a[81]), .Z(n30827) );
  NANDN U31249 ( .A(n30827), .B(n38075), .Z(n30636) );
  NANDN U31250 ( .A(n30634), .B(n38073), .Z(n30635) );
  NAND U31251 ( .A(n30636), .B(n30635), .Z(n30779) );
  XOR U31252 ( .A(b[43]), .B(n35377), .Z(n30836) );
  NANDN U31253 ( .A(n30836), .B(n37068), .Z(n30639) );
  NANDN U31254 ( .A(n30637), .B(n37069), .Z(n30638) );
  AND U31255 ( .A(n30639), .B(n30638), .Z(n30780) );
  XNOR U31256 ( .A(n30779), .B(n30780), .Z(n30781) );
  XOR U31257 ( .A(n30782), .B(n30781), .Z(n30950) );
  XNOR U31258 ( .A(b[51]), .B(a[85]), .Z(n30937) );
  NANDN U31259 ( .A(n30937), .B(n37803), .Z(n30642) );
  NANDN U31260 ( .A(n30640), .B(n37802), .Z(n30641) );
  NAND U31261 ( .A(n30642), .B(n30641), .Z(n30758) );
  XNOR U31262 ( .A(a[121]), .B(b[15]), .Z(n30833) );
  OR U31263 ( .A(n30833), .B(n32010), .Z(n30645) );
  NANDN U31264 ( .A(n30643), .B(n32011), .Z(n30644) );
  NAND U31265 ( .A(n30645), .B(n30644), .Z(n30755) );
  XNOR U31266 ( .A(a[123]), .B(b[13]), .Z(n30913) );
  OR U31267 ( .A(n30913), .B(n31550), .Z(n30648) );
  NANDN U31268 ( .A(n30646), .B(n31874), .Z(n30647) );
  AND U31269 ( .A(n30648), .B(n30647), .Z(n30756) );
  XNOR U31270 ( .A(n30755), .B(n30756), .Z(n30757) );
  XOR U31271 ( .A(n30758), .B(n30757), .Z(n30951) );
  XNOR U31272 ( .A(n30950), .B(n30951), .Z(n30953) );
  XNOR U31273 ( .A(n30952), .B(n30953), .Z(n30874) );
  NANDN U31274 ( .A(n30650), .B(n30649), .Z(n30654) );
  NAND U31275 ( .A(n30652), .B(n30651), .Z(n30653) );
  NAND U31276 ( .A(n30654), .B(n30653), .Z(n30871) );
  OR U31277 ( .A(n30655), .B(n30942), .Z(n30659) );
  NANDN U31278 ( .A(n30657), .B(n30656), .Z(n30658) );
  AND U31279 ( .A(n30659), .B(n30658), .Z(n30872) );
  XNOR U31280 ( .A(n30871), .B(n30872), .Z(n30873) );
  XNOR U31281 ( .A(n30874), .B(n30873), .Z(n30798) );
  XNOR U31282 ( .A(n30797), .B(n30798), .Z(n30799) );
  XNOR U31283 ( .A(n30800), .B(n30799), .Z(n30734) );
  XNOR U31284 ( .A(n30733), .B(n30734), .Z(n30735) );
  XOR U31285 ( .A(n30736), .B(n30735), .Z(n30728) );
  XNOR U31286 ( .A(n30727), .B(n30728), .Z(n30729) );
  XNOR U31287 ( .A(n30730), .B(n30729), .Z(n30724) );
  NANDN U31288 ( .A(n30661), .B(n30660), .Z(n30665) );
  OR U31289 ( .A(n30663), .B(n30662), .Z(n30664) );
  NAND U31290 ( .A(n30665), .B(n30664), .Z(n30959) );
  OR U31291 ( .A(n30667), .B(n30666), .Z(n30671) );
  NANDN U31292 ( .A(n30669), .B(n30668), .Z(n30670) );
  NAND U31293 ( .A(n30671), .B(n30670), .Z(n30956) );
  NANDN U31294 ( .A(n30673), .B(n30672), .Z(n30677) );
  OR U31295 ( .A(n30675), .B(n30674), .Z(n30676) );
  NAND U31296 ( .A(n30677), .B(n30676), .Z(n30957) );
  XNOR U31297 ( .A(n30956), .B(n30957), .Z(n30958) );
  XOR U31298 ( .A(n30959), .B(n30958), .Z(n30722) );
  NANDN U31299 ( .A(n30679), .B(n30678), .Z(n30683) );
  OR U31300 ( .A(n30681), .B(n30680), .Z(n30682) );
  AND U31301 ( .A(n30683), .B(n30682), .Z(n30721) );
  XNOR U31302 ( .A(n30722), .B(n30721), .Z(n30723) );
  XNOR U31303 ( .A(n30724), .B(n30723), .Z(n30715) );
  XOR U31304 ( .A(n30716), .B(n30715), .Z(n30717) );
  NANDN U31305 ( .A(n30685), .B(n30684), .Z(n30689) );
  NANDN U31306 ( .A(n30687), .B(n30686), .Z(n30688) );
  NAND U31307 ( .A(n30689), .B(n30688), .Z(n30718) );
  XOR U31308 ( .A(n30717), .B(n30718), .Z(n30709) );
  NANDN U31309 ( .A(n30691), .B(n30690), .Z(n30695) );
  NAND U31310 ( .A(n30693), .B(n30692), .Z(n30694) );
  NAND U31311 ( .A(n30695), .B(n30694), .Z(n30710) );
  XNOR U31312 ( .A(n30709), .B(n30710), .Z(n30711) );
  NANDN U31313 ( .A(n30697), .B(n30696), .Z(n30701) );
  NAND U31314 ( .A(n30699), .B(n30698), .Z(n30700) );
  NAND U31315 ( .A(n30701), .B(n30700), .Z(n30712) );
  XOR U31316 ( .A(n30711), .B(n30712), .Z(n30703) );
  XNOR U31317 ( .A(n30706), .B(n30703), .Z(n30702) );
  XNOR U31318 ( .A(n30705), .B(n30702), .Z(n30962) );
  XOR U31319 ( .A(n30963), .B(n30962), .Z(c[199]) );
  XOR U31320 ( .A(n30706), .B(n30705), .Z(n30704) );
  NAND U31321 ( .A(n30704), .B(n30703), .Z(n30708) );
  OR U31322 ( .A(n30706), .B(n30705), .Z(n30707) );
  AND U31323 ( .A(n30708), .B(n30707), .Z(n30975) );
  NANDN U31324 ( .A(n30710), .B(n30709), .Z(n30714) );
  NANDN U31325 ( .A(n30712), .B(n30711), .Z(n30713) );
  NAND U31326 ( .A(n30714), .B(n30713), .Z(n30972) );
  OR U31327 ( .A(n30716), .B(n30715), .Z(n30720) );
  NANDN U31328 ( .A(n30718), .B(n30717), .Z(n30719) );
  NAND U31329 ( .A(n30720), .B(n30719), .Z(n30966) );
  OR U31330 ( .A(n30722), .B(n30721), .Z(n30726) );
  OR U31331 ( .A(n30724), .B(n30723), .Z(n30725) );
  AND U31332 ( .A(n30726), .B(n30725), .Z(n30967) );
  XNOR U31333 ( .A(n30966), .B(n30967), .Z(n30968) );
  NANDN U31334 ( .A(n30728), .B(n30727), .Z(n30732) );
  NAND U31335 ( .A(n30730), .B(n30729), .Z(n30731) );
  NAND U31336 ( .A(n30732), .B(n30731), .Z(n30979) );
  NANDN U31337 ( .A(n30734), .B(n30733), .Z(n30738) );
  NANDN U31338 ( .A(n30736), .B(n30735), .Z(n30737) );
  NAND U31339 ( .A(n30738), .B(n30737), .Z(n30984) );
  NAND U31340 ( .A(n30740), .B(n30739), .Z(n30744) );
  NANDN U31341 ( .A(n30742), .B(n30741), .Z(n30743) );
  AND U31342 ( .A(n30744), .B(n30743), .Z(n30985) );
  XNOR U31343 ( .A(n30984), .B(n30985), .Z(n30986) );
  NANDN U31344 ( .A(n30750), .B(n30749), .Z(n30754) );
  NAND U31345 ( .A(n30752), .B(n30751), .Z(n30753) );
  NAND U31346 ( .A(n30754), .B(n30753), .Z(n31076) );
  NANDN U31347 ( .A(n30756), .B(n30755), .Z(n30760) );
  NAND U31348 ( .A(n30758), .B(n30757), .Z(n30759) );
  NAND U31349 ( .A(n30760), .B(n30759), .Z(n31139) );
  XOR U31350 ( .A(b[57]), .B(n32814), .Z(n31187) );
  OR U31351 ( .A(n31187), .B(n965), .Z(n30763) );
  NANDN U31352 ( .A(n30761), .B(n38194), .Z(n30762) );
  NAND U31353 ( .A(n30763), .B(n30762), .Z(n31208) );
  XNOR U31354 ( .A(a[112]), .B(b[25]), .Z(n31184) );
  OR U31355 ( .A(n31184), .B(n34219), .Z(n30766) );
  NAND U31356 ( .A(n34217), .B(n30764), .Z(n30765) );
  NAND U31357 ( .A(n30766), .B(n30765), .Z(n31205) );
  NAND U31358 ( .A(n30767), .B(n34044), .Z(n30769) );
  XOR U31359 ( .A(n37873), .B(n34510), .Z(n31181) );
  NANDN U31360 ( .A(n33867), .B(n31181), .Z(n30768) );
  AND U31361 ( .A(n30769), .B(n30768), .Z(n31206) );
  XNOR U31362 ( .A(n31205), .B(n31206), .Z(n31207) );
  XOR U31363 ( .A(n31208), .B(n31207), .Z(n31136) );
  XOR U31364 ( .A(b[39]), .B(n35783), .Z(n31116) );
  NANDN U31365 ( .A(n31116), .B(n36553), .Z(n30772) );
  NANDN U31366 ( .A(n30770), .B(n36643), .Z(n30771) );
  NAND U31367 ( .A(n30772), .B(n30771), .Z(n31041) );
  XOR U31368 ( .A(a[126]), .B(n970), .Z(n31120) );
  OR U31369 ( .A(n31120), .B(n31369), .Z(n30775) );
  NANDN U31370 ( .A(n30773), .B(n31119), .Z(n30774) );
  NAND U31371 ( .A(n30775), .B(n30774), .Z(n31038) );
  XOR U31372 ( .A(b[61]), .B(n31363), .Z(n31023) );
  OR U31373 ( .A(n31023), .B(n38371), .Z(n30778) );
  NAND U31374 ( .A(n30776), .B(n38369), .Z(n30777) );
  AND U31375 ( .A(n30778), .B(n30777), .Z(n31039) );
  XNOR U31376 ( .A(n31038), .B(n31039), .Z(n31040) );
  XOR U31377 ( .A(n31041), .B(n31040), .Z(n31137) );
  XNOR U31378 ( .A(n31136), .B(n31137), .Z(n31138) );
  XNOR U31379 ( .A(n31139), .B(n31138), .Z(n31074) );
  NANDN U31380 ( .A(n30780), .B(n30779), .Z(n30784) );
  NAND U31381 ( .A(n30782), .B(n30781), .Z(n30783) );
  AND U31382 ( .A(n30784), .B(n30783), .Z(n31075) );
  XOR U31383 ( .A(n31074), .B(n31075), .Z(n31077) );
  XNOR U31384 ( .A(n31076), .B(n31077), .Z(n31068) );
  NANDN U31385 ( .A(n30786), .B(n30785), .Z(n30790) );
  OR U31386 ( .A(n30788), .B(n30787), .Z(n30789) );
  AND U31387 ( .A(n30790), .B(n30789), .Z(n31069) );
  XNOR U31388 ( .A(n31068), .B(n31069), .Z(n31070) );
  XOR U31389 ( .A(n31071), .B(n31070), .Z(n31219) );
  NANDN U31390 ( .A(n30792), .B(n30791), .Z(n30796) );
  NANDN U31391 ( .A(n30794), .B(n30793), .Z(n30795) );
  NAND U31392 ( .A(n30796), .B(n30795), .Z(n31218) );
  NANDN U31393 ( .A(n30798), .B(n30797), .Z(n30802) );
  NAND U31394 ( .A(n30800), .B(n30799), .Z(n30801) );
  NAND U31395 ( .A(n30802), .B(n30801), .Z(n31217) );
  XNOR U31396 ( .A(n31218), .B(n31217), .Z(n31220) );
  XNOR U31397 ( .A(n31219), .B(n31220), .Z(n30992) );
  OR U31398 ( .A(n30804), .B(n30803), .Z(n30808) );
  NANDN U31399 ( .A(n30806), .B(n30805), .Z(n30807) );
  NAND U31400 ( .A(n30808), .B(n30807), .Z(n30991) );
  NANDN U31401 ( .A(n30810), .B(n30809), .Z(n30814) );
  NAND U31402 ( .A(n30812), .B(n30811), .Z(n30813) );
  NAND U31403 ( .A(n30814), .B(n30813), .Z(n31065) );
  NANDN U31404 ( .A(n30816), .B(n30815), .Z(n30820) );
  NAND U31405 ( .A(n30818), .B(n30817), .Z(n30819) );
  NAND U31406 ( .A(n30820), .B(n30819), .Z(n31010) );
  NAND U31407 ( .A(n34848), .B(n30821), .Z(n30823) );
  XOR U31408 ( .A(n37336), .B(n35375), .Z(n31178) );
  NAND U31409 ( .A(n34618), .B(n31178), .Z(n30822) );
  NAND U31410 ( .A(n30823), .B(n30822), .Z(n31035) );
  XOR U31411 ( .A(b[53]), .B(n33185), .Z(n31095) );
  NANDN U31412 ( .A(n31095), .B(n37940), .Z(n30826) );
  NANDN U31413 ( .A(n30824), .B(n37941), .Z(n30825) );
  NAND U31414 ( .A(n30826), .B(n30825), .Z(n31032) );
  XOR U31415 ( .A(b[55]), .B(n32815), .Z(n31098) );
  NANDN U31416 ( .A(n31098), .B(n38075), .Z(n30829) );
  NANDN U31417 ( .A(n30827), .B(n38073), .Z(n30828) );
  AND U31418 ( .A(n30829), .B(n30828), .Z(n31033) );
  XNOR U31419 ( .A(n31032), .B(n31033), .Z(n31034) );
  XNOR U31420 ( .A(n31035), .B(n31034), .Z(n31008) );
  XNOR U31421 ( .A(a[120]), .B(b[17]), .Z(n31014) );
  NANDN U31422 ( .A(n31014), .B(n32543), .Z(n30832) );
  NANDN U31423 ( .A(n30830), .B(n32541), .Z(n30831) );
  NAND U31424 ( .A(n30832), .B(n30831), .Z(n31163) );
  XOR U31425 ( .A(a[122]), .B(n972), .Z(n31026) );
  OR U31426 ( .A(n31026), .B(n32010), .Z(n30835) );
  NANDN U31427 ( .A(n30833), .B(n32011), .Z(n30834) );
  NAND U31428 ( .A(n30835), .B(n30834), .Z(n31160) );
  XOR U31429 ( .A(b[43]), .B(n35191), .Z(n31029) );
  NANDN U31430 ( .A(n31029), .B(n37068), .Z(n30838) );
  NANDN U31431 ( .A(n30836), .B(n37069), .Z(n30837) );
  AND U31432 ( .A(n30838), .B(n30837), .Z(n31161) );
  XNOR U31433 ( .A(n31160), .B(n31161), .Z(n31162) );
  XOR U31434 ( .A(n31163), .B(n31162), .Z(n31009) );
  XOR U31435 ( .A(n31008), .B(n31009), .Z(n31011) );
  XOR U31436 ( .A(n31010), .B(n31011), .Z(n31058) );
  XOR U31437 ( .A(b[63]), .B(n31372), .Z(n31092) );
  NANDN U31438 ( .A(n31092), .B(n38422), .Z(n30845) );
  NANDN U31439 ( .A(n30843), .B(n38423), .Z(n30844) );
  NAND U31440 ( .A(n30845), .B(n30844), .Z(n31126) );
  NANDN U31441 ( .A(n30847), .B(n30846), .Z(n30848) );
  NANDN U31442 ( .A(n30849), .B(n30848), .Z(n31125) );
  AND U31443 ( .A(b[63]), .B(a[72]), .Z(n31445) );
  XOR U31444 ( .A(n31125), .B(n31445), .Z(n31127) );
  XNOR U31445 ( .A(n31126), .B(n31127), .Z(n31130) );
  NANDN U31446 ( .A(n30851), .B(n30850), .Z(n30855) );
  NANDN U31447 ( .A(n30853), .B(n30852), .Z(n30854) );
  NAND U31448 ( .A(n30855), .B(n30854), .Z(n31131) );
  XOR U31449 ( .A(n31130), .B(n31131), .Z(n31132) );
  NANDN U31450 ( .A(n30856), .B(n37469), .Z(n30858) );
  XNOR U31451 ( .A(n978), .B(a[90]), .Z(n31199) );
  NAND U31452 ( .A(n31199), .B(n37471), .Z(n30857) );
  AND U31453 ( .A(n30858), .B(n30857), .Z(n31110) );
  XOR U31454 ( .A(b[37]), .B(n36100), .Z(n31193) );
  NANDN U31455 ( .A(n31193), .B(n36311), .Z(n30861) );
  NAND U31456 ( .A(n30859), .B(n36309), .Z(n30860) );
  AND U31457 ( .A(n30861), .B(n30860), .Z(n31111) );
  XOR U31458 ( .A(n31110), .B(n31111), .Z(n31112) );
  XOR U31459 ( .A(a[106]), .B(n973), .Z(n31172) );
  NANDN U31460 ( .A(n31172), .B(n35313), .Z(n30864) );
  NANDN U31461 ( .A(n30862), .B(n35311), .Z(n30863) );
  AND U31462 ( .A(n30864), .B(n30863), .Z(n31113) );
  XNOR U31463 ( .A(n31112), .B(n31113), .Z(n31157) );
  XNOR U31464 ( .A(n36647), .B(b[33]), .Z(n31017) );
  NAND U31465 ( .A(n35620), .B(n31017), .Z(n30867) );
  NANDN U31466 ( .A(n30865), .B(n35621), .Z(n30866) );
  NAND U31467 ( .A(n30867), .B(n30866), .Z(n31155) );
  NANDN U31468 ( .A(n30868), .B(n35986), .Z(n30870) );
  XNOR U31469 ( .A(a[102]), .B(b[35]), .Z(n31020) );
  NANDN U31470 ( .A(n31020), .B(n35985), .Z(n30869) );
  AND U31471 ( .A(n30870), .B(n30869), .Z(n31154) );
  XNOR U31472 ( .A(n31155), .B(n31154), .Z(n31156) );
  XOR U31473 ( .A(n31157), .B(n31156), .Z(n31133) );
  XOR U31474 ( .A(n31132), .B(n31133), .Z(n31056) );
  XNOR U31475 ( .A(n31058), .B(n31059), .Z(n31063) );
  NANDN U31476 ( .A(n30872), .B(n30871), .Z(n30876) );
  NANDN U31477 ( .A(n30874), .B(n30873), .Z(n30875) );
  AND U31478 ( .A(n30876), .B(n30875), .Z(n31062) );
  XOR U31479 ( .A(n31063), .B(n31062), .Z(n31064) );
  XNOR U31480 ( .A(n31065), .B(n31064), .Z(n30999) );
  OR U31481 ( .A(n30878), .B(n30877), .Z(n30882) );
  NAND U31482 ( .A(n30880), .B(n30879), .Z(n30881) );
  NAND U31483 ( .A(n30882), .B(n30881), .Z(n30996) );
  OR U31484 ( .A(n30884), .B(n30883), .Z(n30888) );
  OR U31485 ( .A(n30886), .B(n30885), .Z(n30887) );
  NAND U31486 ( .A(n30888), .B(n30887), .Z(n31053) );
  NANDN U31487 ( .A(n30890), .B(n30889), .Z(n30894) );
  NAND U31488 ( .A(n30892), .B(n30891), .Z(n30893) );
  NAND U31489 ( .A(n30894), .B(n30893), .Z(n31005) );
  NANDN U31490 ( .A(n30896), .B(n30895), .Z(n30900) );
  NAND U31491 ( .A(n30898), .B(n30897), .Z(n30899) );
  NAND U31492 ( .A(n30900), .B(n30899), .Z(n31002) );
  NANDN U31493 ( .A(n30902), .B(n30901), .Z(n30906) );
  NAND U31494 ( .A(n30904), .B(n30903), .Z(n30905) );
  NAND U31495 ( .A(n30906), .B(n30905), .Z(n31003) );
  XNOR U31496 ( .A(n31002), .B(n31003), .Z(n31004) );
  XOR U31497 ( .A(n31005), .B(n31004), .Z(n31214) );
  XNOR U31498 ( .A(b[41]), .B(a[96]), .Z(n31086) );
  OR U31499 ( .A(n31086), .B(n36905), .Z(n30909) );
  NANDN U31500 ( .A(n30907), .B(n36807), .Z(n30908) );
  NAND U31501 ( .A(n30909), .B(n30908), .Z(n31151) );
  NAND U31502 ( .A(n38326), .B(n30910), .Z(n30912) );
  XOR U31503 ( .A(n38400), .B(n31870), .Z(n31190) );
  NANDN U31504 ( .A(n38273), .B(n31190), .Z(n30911) );
  NAND U31505 ( .A(n30912), .B(n30911), .Z(n31148) );
  XOR U31506 ( .A(a[124]), .B(n971), .Z(n31089) );
  OR U31507 ( .A(n31089), .B(n31550), .Z(n30915) );
  NANDN U31508 ( .A(n30913), .B(n31874), .Z(n30914) );
  AND U31509 ( .A(n30915), .B(n30914), .Z(n31149) );
  XNOR U31510 ( .A(n31148), .B(n31149), .Z(n31150) );
  XNOR U31511 ( .A(n31151), .B(n31150), .Z(n31142) );
  XNOR U31512 ( .A(a[116]), .B(b[21]), .Z(n31175) );
  OR U31513 ( .A(n31175), .B(n33634), .Z(n30918) );
  NAND U31514 ( .A(n30916), .B(n33464), .Z(n30917) );
  NAND U31515 ( .A(n30918), .B(n30917), .Z(n31047) );
  NAND U31516 ( .A(n33283), .B(n30919), .Z(n30921) );
  XOR U31517 ( .A(n38143), .B(n33020), .Z(n31166) );
  NANDN U31518 ( .A(n33021), .B(n31166), .Z(n30920) );
  NAND U31519 ( .A(n30921), .B(n30920), .Z(n31044) );
  XNOR U31520 ( .A(b[45]), .B(a[92]), .Z(n31101) );
  NANDN U31521 ( .A(n31101), .B(n37261), .Z(n30924) );
  NAND U31522 ( .A(n30922), .B(n37262), .Z(n30923) );
  AND U31523 ( .A(n30924), .B(n30923), .Z(n31045) );
  XNOR U31524 ( .A(n31044), .B(n31045), .Z(n31046) );
  XOR U31525 ( .A(n31047), .B(n31046), .Z(n31143) );
  XOR U31526 ( .A(n31142), .B(n31143), .Z(n31145) );
  NANDN U31527 ( .A(n30926), .B(n30925), .Z(n30930) );
  NAND U31528 ( .A(n30928), .B(n30927), .Z(n30929) );
  NAND U31529 ( .A(n30930), .B(n30929), .Z(n31144) );
  XNOR U31530 ( .A(n31145), .B(n31144), .Z(n31211) );
  NAND U31531 ( .A(n35188), .B(n30931), .Z(n30933) );
  XOR U31532 ( .A(n37139), .B(n35540), .Z(n31169) );
  NANDN U31533 ( .A(n34968), .B(n31169), .Z(n30932) );
  NAND U31534 ( .A(n30933), .B(n30932), .Z(n31083) );
  XOR U31535 ( .A(b[49]), .B(n34048), .Z(n31202) );
  OR U31536 ( .A(n31202), .B(n37756), .Z(n30936) );
  NANDN U31537 ( .A(n30934), .B(n37652), .Z(n30935) );
  NAND U31538 ( .A(n30936), .B(n30935), .Z(n31080) );
  XOR U31539 ( .A(b[51]), .B(n33628), .Z(n31196) );
  NANDN U31540 ( .A(n31196), .B(n37803), .Z(n30939) );
  NANDN U31541 ( .A(n30937), .B(n37802), .Z(n30938) );
  AND U31542 ( .A(n30939), .B(n30938), .Z(n31081) );
  XNOR U31543 ( .A(n31080), .B(n31081), .Z(n31082) );
  XNOR U31544 ( .A(n31083), .B(n31082), .Z(n31107) );
  NANDN U31545 ( .A(n30945), .B(n30944), .Z(n30949) );
  NAND U31546 ( .A(n30947), .B(n30946), .Z(n30948) );
  AND U31547 ( .A(n30949), .B(n30948), .Z(n31104) );
  XNOR U31548 ( .A(n31105), .B(n31104), .Z(n31106) );
  XOR U31549 ( .A(n31107), .B(n31106), .Z(n31212) );
  XNOR U31550 ( .A(n31211), .B(n31212), .Z(n31213) );
  XNOR U31551 ( .A(n31214), .B(n31213), .Z(n31050) );
  OR U31552 ( .A(n30951), .B(n30950), .Z(n30955) );
  NANDN U31553 ( .A(n30953), .B(n30952), .Z(n30954) );
  AND U31554 ( .A(n30955), .B(n30954), .Z(n31051) );
  XNOR U31555 ( .A(n31050), .B(n31051), .Z(n31052) );
  XNOR U31556 ( .A(n31053), .B(n31052), .Z(n30997) );
  XNOR U31557 ( .A(n30996), .B(n30997), .Z(n30998) );
  XOR U31558 ( .A(n30999), .B(n30998), .Z(n30990) );
  XOR U31559 ( .A(n30991), .B(n30990), .Z(n30993) );
  XOR U31560 ( .A(n30992), .B(n30993), .Z(n30987) );
  XOR U31561 ( .A(n30986), .B(n30987), .Z(n30978) );
  XNOR U31562 ( .A(n30979), .B(n30978), .Z(n30981) );
  NANDN U31563 ( .A(n30957), .B(n30956), .Z(n30961) );
  NAND U31564 ( .A(n30959), .B(n30958), .Z(n30960) );
  AND U31565 ( .A(n30961), .B(n30960), .Z(n30980) );
  XNOR U31566 ( .A(n30981), .B(n30980), .Z(n30969) );
  XOR U31567 ( .A(n30968), .B(n30969), .Z(n30973) );
  XNOR U31568 ( .A(n30972), .B(n30973), .Z(n30974) );
  XNOR U31569 ( .A(n30975), .B(n30974), .Z(n30965) );
  OR U31570 ( .A(n30963), .B(n30962), .Z(n30964) );
  XOR U31571 ( .A(n30965), .B(n30964), .Z(c[200]) );
  OR U31572 ( .A(n30965), .B(n30964), .Z(n31482) );
  NANDN U31573 ( .A(n30967), .B(n30966), .Z(n30971) );
  NAND U31574 ( .A(n30969), .B(n30968), .Z(n30970) );
  NAND U31575 ( .A(n30971), .B(n30970), .Z(n31226) );
  NANDN U31576 ( .A(n30973), .B(n30972), .Z(n30977) );
  NAND U31577 ( .A(n30975), .B(n30974), .Z(n30976) );
  NAND U31578 ( .A(n30977), .B(n30976), .Z(n31227) );
  NAND U31579 ( .A(n30979), .B(n30978), .Z(n30983) );
  NANDN U31580 ( .A(n30981), .B(n30980), .Z(n30982) );
  NAND U31581 ( .A(n30983), .B(n30982), .Z(n31230) );
  NANDN U31582 ( .A(n30985), .B(n30984), .Z(n30989) );
  NAND U31583 ( .A(n30987), .B(n30986), .Z(n30988) );
  NAND U31584 ( .A(n30989), .B(n30988), .Z(n31229) );
  NANDN U31585 ( .A(n30991), .B(n30990), .Z(n30995) );
  OR U31586 ( .A(n30993), .B(n30992), .Z(n30994) );
  NAND U31587 ( .A(n30995), .B(n30994), .Z(n31476) );
  NANDN U31588 ( .A(n30997), .B(n30996), .Z(n31001) );
  NAND U31589 ( .A(n30999), .B(n30998), .Z(n31000) );
  NAND U31590 ( .A(n31001), .B(n31000), .Z(n31469) );
  NANDN U31591 ( .A(n31003), .B(n31002), .Z(n31007) );
  NANDN U31592 ( .A(n31005), .B(n31004), .Z(n31006) );
  NAND U31593 ( .A(n31007), .B(n31006), .Z(n31397) );
  NANDN U31594 ( .A(n31009), .B(n31008), .Z(n31013) );
  OR U31595 ( .A(n31011), .B(n31010), .Z(n31012) );
  NAND U31596 ( .A(n31013), .B(n31012), .Z(n31394) );
  XOR U31597 ( .A(a[121]), .B(b[17]), .Z(n31273) );
  NAND U31598 ( .A(n31273), .B(n32543), .Z(n31016) );
  NANDN U31599 ( .A(n31014), .B(n32541), .Z(n31015) );
  NAND U31600 ( .A(n31016), .B(n31015), .Z(n31342) );
  XNOR U31601 ( .A(a[105]), .B(b[33]), .Z(n31276) );
  NANDN U31602 ( .A(n31276), .B(n35620), .Z(n31019) );
  NAND U31603 ( .A(n31017), .B(n35621), .Z(n31018) );
  NAND U31604 ( .A(n31019), .B(n31018), .Z(n31339) );
  XOR U31605 ( .A(a[103]), .B(b[35]), .Z(n31279) );
  NAND U31606 ( .A(n35985), .B(n31279), .Z(n31022) );
  NANDN U31607 ( .A(n31020), .B(n35986), .Z(n31021) );
  AND U31608 ( .A(n31022), .B(n31021), .Z(n31340) );
  XNOR U31609 ( .A(n31339), .B(n31340), .Z(n31341) );
  XOR U31610 ( .A(n31342), .B(n31341), .Z(n31385) );
  XNOR U31611 ( .A(b[61]), .B(a[77]), .Z(n31360) );
  OR U31612 ( .A(n31360), .B(n38371), .Z(n31025) );
  NANDN U31613 ( .A(n31023), .B(n38369), .Z(n31024) );
  NAND U31614 ( .A(n31025), .B(n31024), .Z(n31433) );
  XNOR U31615 ( .A(a[123]), .B(b[15]), .Z(n31333) );
  OR U31616 ( .A(n31333), .B(n32010), .Z(n31028) );
  NANDN U31617 ( .A(n31026), .B(n32011), .Z(n31027) );
  NAND U31618 ( .A(n31028), .B(n31027), .Z(n31430) );
  XOR U31619 ( .A(b[43]), .B(n35628), .Z(n31321) );
  NANDN U31620 ( .A(n31321), .B(n37068), .Z(n31031) );
  NANDN U31621 ( .A(n31029), .B(n37069), .Z(n31030) );
  AND U31622 ( .A(n31031), .B(n31030), .Z(n31431) );
  XNOR U31623 ( .A(n31430), .B(n31431), .Z(n31432) );
  XOR U31624 ( .A(n31433), .B(n31432), .Z(n31383) );
  NANDN U31625 ( .A(n31033), .B(n31032), .Z(n31037) );
  NAND U31626 ( .A(n31035), .B(n31034), .Z(n31036) );
  NAND U31627 ( .A(n31037), .B(n31036), .Z(n31382) );
  XNOR U31628 ( .A(n31383), .B(n31382), .Z(n31384) );
  XOR U31629 ( .A(n31385), .B(n31384), .Z(n31249) );
  NANDN U31630 ( .A(n31039), .B(n31038), .Z(n31043) );
  NAND U31631 ( .A(n31041), .B(n31040), .Z(n31042) );
  NAND U31632 ( .A(n31043), .B(n31042), .Z(n31246) );
  NANDN U31633 ( .A(n31045), .B(n31044), .Z(n31049) );
  NAND U31634 ( .A(n31047), .B(n31046), .Z(n31048) );
  AND U31635 ( .A(n31049), .B(n31048), .Z(n31247) );
  XNOR U31636 ( .A(n31246), .B(n31247), .Z(n31248) );
  XNOR U31637 ( .A(n31249), .B(n31248), .Z(n31395) );
  XNOR U31638 ( .A(n31394), .B(n31395), .Z(n31396) );
  XNOR U31639 ( .A(n31397), .B(n31396), .Z(n31466) );
  NANDN U31640 ( .A(n31051), .B(n31050), .Z(n31055) );
  NAND U31641 ( .A(n31053), .B(n31052), .Z(n31054) );
  NAND U31642 ( .A(n31055), .B(n31054), .Z(n31464) );
  OR U31643 ( .A(n31057), .B(n31056), .Z(n31061) );
  NANDN U31644 ( .A(n31059), .B(n31058), .Z(n31060) );
  AND U31645 ( .A(n31061), .B(n31060), .Z(n31463) );
  XNOR U31646 ( .A(n31464), .B(n31463), .Z(n31465) );
  XOR U31647 ( .A(n31466), .B(n31465), .Z(n31470) );
  XNOR U31648 ( .A(n31469), .B(n31470), .Z(n31471) );
  OR U31649 ( .A(n31063), .B(n31062), .Z(n31067) );
  NAND U31650 ( .A(n31065), .B(n31064), .Z(n31066) );
  NAND U31651 ( .A(n31067), .B(n31066), .Z(n31237) );
  NANDN U31652 ( .A(n31069), .B(n31068), .Z(n31073) );
  NANDN U31653 ( .A(n31071), .B(n31070), .Z(n31072) );
  NAND U31654 ( .A(n31073), .B(n31072), .Z(n31235) );
  NANDN U31655 ( .A(n31075), .B(n31074), .Z(n31079) );
  OR U31656 ( .A(n31077), .B(n31076), .Z(n31078) );
  NAND U31657 ( .A(n31079), .B(n31078), .Z(n31243) );
  NANDN U31658 ( .A(n31081), .B(n31080), .Z(n31085) );
  NAND U31659 ( .A(n31083), .B(n31082), .Z(n31084) );
  NAND U31660 ( .A(n31085), .B(n31084), .Z(n31459) );
  XOR U31661 ( .A(b[41]), .B(a[97]), .Z(n31357) );
  NANDN U31662 ( .A(n36905), .B(n31357), .Z(n31088) );
  NANDN U31663 ( .A(n31086), .B(n36807), .Z(n31087) );
  NAND U31664 ( .A(n31088), .B(n31087), .Z(n31427) );
  XNOR U31665 ( .A(a[125]), .B(n971), .Z(n31373) );
  NANDN U31666 ( .A(n31550), .B(n31373), .Z(n31091) );
  NANDN U31667 ( .A(n31089), .B(n31874), .Z(n31090) );
  NAND U31668 ( .A(n31091), .B(n31090), .Z(n31424) );
  XNOR U31669 ( .A(b[63]), .B(a[75]), .Z(n31364) );
  NANDN U31670 ( .A(n31364), .B(n38422), .Z(n31094) );
  NANDN U31671 ( .A(n31092), .B(n38423), .Z(n31093) );
  AND U31672 ( .A(n31094), .B(n31093), .Z(n31425) );
  XNOR U31673 ( .A(n31424), .B(n31425), .Z(n31426) );
  XNOR U31674 ( .A(n31427), .B(n31426), .Z(n31457) );
  XNOR U31675 ( .A(b[53]), .B(a[85]), .Z(n31327) );
  NANDN U31676 ( .A(n31327), .B(n37940), .Z(n31097) );
  NANDN U31677 ( .A(n31095), .B(n37941), .Z(n31096) );
  NAND U31678 ( .A(n31097), .B(n31096), .Z(n31297) );
  XNOR U31679 ( .A(b[55]), .B(a[83]), .Z(n31330) );
  NANDN U31680 ( .A(n31330), .B(n38075), .Z(n31100) );
  NANDN U31681 ( .A(n31098), .B(n38073), .Z(n31099) );
  NAND U31682 ( .A(n31100), .B(n31099), .Z(n31294) );
  XNOR U31683 ( .A(b[45]), .B(a[93]), .Z(n31267) );
  NANDN U31684 ( .A(n31267), .B(n37261), .Z(n31103) );
  NANDN U31685 ( .A(n31101), .B(n37262), .Z(n31102) );
  AND U31686 ( .A(n31103), .B(n31102), .Z(n31295) );
  XNOR U31687 ( .A(n31294), .B(n31295), .Z(n31296) );
  XOR U31688 ( .A(n31297), .B(n31296), .Z(n31458) );
  XOR U31689 ( .A(n31457), .B(n31458), .Z(n31460) );
  XOR U31690 ( .A(n31459), .B(n31460), .Z(n31408) );
  NANDN U31691 ( .A(n31105), .B(n31104), .Z(n31109) );
  NAND U31692 ( .A(n31107), .B(n31106), .Z(n31108) );
  AND U31693 ( .A(n31109), .B(n31108), .Z(n31407) );
  OR U31694 ( .A(n31111), .B(n31110), .Z(n31115) );
  NANDN U31695 ( .A(n31113), .B(n31112), .Z(n31114) );
  NAND U31696 ( .A(n31115), .B(n31114), .Z(n31254) );
  XNOR U31697 ( .A(b[39]), .B(a[99]), .Z(n31454) );
  NANDN U31698 ( .A(n31454), .B(n36553), .Z(n31118) );
  NANDN U31699 ( .A(n31116), .B(n36643), .Z(n31117) );
  NAND U31700 ( .A(n31118), .B(n31117), .Z(n31291) );
  XOR U31701 ( .A(a[127]), .B(n970), .Z(n31368) );
  OR U31702 ( .A(n31368), .B(n31369), .Z(n31122) );
  NANDN U31703 ( .A(n31120), .B(n31119), .Z(n31121) );
  NAND U31704 ( .A(n31122), .B(n31121), .Z(n31288) );
  NANDN U31705 ( .A(n31123), .B(b[8]), .Z(n31124) );
  AND U31706 ( .A(n31124), .B(b[9]), .Z(n31442) );
  NANDN U31707 ( .A(n985), .B(a[73]), .Z(n31443) );
  XOR U31708 ( .A(n31442), .B(n31443), .Z(n31444) );
  XNOR U31709 ( .A(n31445), .B(n31444), .Z(n31289) );
  XNOR U31710 ( .A(n31288), .B(n31289), .Z(n31290) );
  XNOR U31711 ( .A(n31291), .B(n31290), .Z(n31252) );
  NANDN U31712 ( .A(n31445), .B(n31125), .Z(n31129) );
  NANDN U31713 ( .A(n31127), .B(n31126), .Z(n31128) );
  NAND U31714 ( .A(n31129), .B(n31128), .Z(n31253) );
  XOR U31715 ( .A(n31252), .B(n31253), .Z(n31255) );
  XNOR U31716 ( .A(n31254), .B(n31255), .Z(n31406) );
  XNOR U31717 ( .A(n31408), .B(n31409), .Z(n31240) );
  OR U31718 ( .A(n31131), .B(n31130), .Z(n31135) );
  NANDN U31719 ( .A(n31133), .B(n31132), .Z(n31134) );
  NAND U31720 ( .A(n31135), .B(n31134), .Z(n31241) );
  XOR U31721 ( .A(n31240), .B(n31241), .Z(n31242) );
  XNOR U31722 ( .A(n31243), .B(n31242), .Z(n31402) );
  OR U31723 ( .A(n31137), .B(n31136), .Z(n31141) );
  OR U31724 ( .A(n31139), .B(n31138), .Z(n31140) );
  NAND U31725 ( .A(n31141), .B(n31140), .Z(n31414) );
  NANDN U31726 ( .A(n31143), .B(n31142), .Z(n31147) );
  OR U31727 ( .A(n31145), .B(n31144), .Z(n31146) );
  NAND U31728 ( .A(n31147), .B(n31146), .Z(n31413) );
  NANDN U31729 ( .A(n31149), .B(n31148), .Z(n31153) );
  NAND U31730 ( .A(n31151), .B(n31150), .Z(n31152) );
  NAND U31731 ( .A(n31153), .B(n31152), .Z(n31421) );
  NANDN U31732 ( .A(n31155), .B(n31154), .Z(n31159) );
  NANDN U31733 ( .A(n31157), .B(n31156), .Z(n31158) );
  NAND U31734 ( .A(n31159), .B(n31158), .Z(n31418) );
  NANDN U31735 ( .A(n31161), .B(n31160), .Z(n31165) );
  NAND U31736 ( .A(n31163), .B(n31162), .Z(n31164) );
  NAND U31737 ( .A(n31165), .B(n31164), .Z(n31419) );
  XNOR U31738 ( .A(n31418), .B(n31419), .Z(n31420) );
  XOR U31739 ( .A(n31421), .B(n31420), .Z(n31391) );
  NAND U31740 ( .A(n33283), .B(n31166), .Z(n31168) );
  XOR U31741 ( .A(n38193), .B(n33020), .Z(n31300) );
  NANDN U31742 ( .A(n33021), .B(n31300), .Z(n31167) );
  NAND U31743 ( .A(n31168), .B(n31167), .Z(n31354) );
  NAND U31744 ( .A(n35188), .B(n31169), .Z(n31171) );
  XNOR U31745 ( .A(a[109]), .B(n35540), .Z(n31303) );
  NANDN U31746 ( .A(n34968), .B(n31303), .Z(n31170) );
  NAND U31747 ( .A(n31171), .B(n31170), .Z(n31351) );
  XNOR U31748 ( .A(a[107]), .B(b[31]), .Z(n31306) );
  NANDN U31749 ( .A(n31306), .B(n35313), .Z(n31174) );
  NANDN U31750 ( .A(n31172), .B(n35311), .Z(n31173) );
  AND U31751 ( .A(n31174), .B(n31173), .Z(n31352) );
  XNOR U31752 ( .A(n31351), .B(n31352), .Z(n31353) );
  XNOR U31753 ( .A(n31354), .B(n31353), .Z(n31285) );
  XOR U31754 ( .A(a[117]), .B(b[21]), .Z(n31309) );
  NANDN U31755 ( .A(n33634), .B(n31309), .Z(n31177) );
  NANDN U31756 ( .A(n31175), .B(n33464), .Z(n31176) );
  NAND U31757 ( .A(n31177), .B(n31176), .Z(n31439) );
  NAND U31758 ( .A(n34848), .B(n31178), .Z(n31180) );
  XNOR U31759 ( .A(a[111]), .B(n35375), .Z(n31318) );
  NAND U31760 ( .A(n34618), .B(n31318), .Z(n31179) );
  NAND U31761 ( .A(n31180), .B(n31179), .Z(n31436) );
  NAND U31762 ( .A(n34044), .B(n31181), .Z(n31183) );
  XNOR U31763 ( .A(a[115]), .B(n34510), .Z(n31315) );
  NANDN U31764 ( .A(n33867), .B(n31315), .Z(n31182) );
  AND U31765 ( .A(n31183), .B(n31182), .Z(n31437) );
  XNOR U31766 ( .A(n31436), .B(n31437), .Z(n31438) );
  XNOR U31767 ( .A(n31439), .B(n31438), .Z(n31282) );
  XOR U31768 ( .A(a[113]), .B(b[25]), .Z(n31312) );
  NANDN U31769 ( .A(n34219), .B(n31312), .Z(n31186) );
  NANDN U31770 ( .A(n31184), .B(n34217), .Z(n31185) );
  NAND U31771 ( .A(n31186), .B(n31185), .Z(n31283) );
  XNOR U31772 ( .A(n31282), .B(n31283), .Z(n31284) );
  XOR U31773 ( .A(n31285), .B(n31284), .Z(n31389) );
  XNOR U31774 ( .A(b[57]), .B(a[81]), .Z(n31448) );
  OR U31775 ( .A(n31448), .B(n965), .Z(n31189) );
  NANDN U31776 ( .A(n31187), .B(n38194), .Z(n31188) );
  NAND U31777 ( .A(n31189), .B(n31188), .Z(n31348) );
  NAND U31778 ( .A(n38326), .B(n31190), .Z(n31192) );
  XNOR U31779 ( .A(n38400), .B(a[79]), .Z(n31451) );
  NANDN U31780 ( .A(n38273), .B(n31451), .Z(n31191) );
  NAND U31781 ( .A(n31192), .B(n31191), .Z(n31345) );
  XNOR U31782 ( .A(b[37]), .B(a[101]), .Z(n31336) );
  NANDN U31783 ( .A(n31336), .B(n36311), .Z(n31195) );
  NANDN U31784 ( .A(n31193), .B(n36309), .Z(n31194) );
  AND U31785 ( .A(n31195), .B(n31194), .Z(n31346) );
  XNOR U31786 ( .A(n31345), .B(n31346), .Z(n31347) );
  XNOR U31787 ( .A(n31348), .B(n31347), .Z(n31376) );
  XNOR U31788 ( .A(b[51]), .B(a[87]), .Z(n31324) );
  NANDN U31789 ( .A(n31324), .B(n37803), .Z(n31198) );
  NANDN U31790 ( .A(n31196), .B(n37802), .Z(n31197) );
  NAND U31791 ( .A(n31198), .B(n31197), .Z(n31261) );
  NAND U31792 ( .A(n31199), .B(n37469), .Z(n31201) );
  XNOR U31793 ( .A(n978), .B(a[91]), .Z(n31270) );
  NAND U31794 ( .A(n31270), .B(n37471), .Z(n31200) );
  NAND U31795 ( .A(n31201), .B(n31200), .Z(n31258) );
  XNOR U31796 ( .A(b[49]), .B(a[89]), .Z(n31264) );
  OR U31797 ( .A(n31264), .B(n37756), .Z(n31204) );
  NANDN U31798 ( .A(n31202), .B(n37652), .Z(n31203) );
  AND U31799 ( .A(n31204), .B(n31203), .Z(n31259) );
  XNOR U31800 ( .A(n31258), .B(n31259), .Z(n31260) );
  XOR U31801 ( .A(n31261), .B(n31260), .Z(n31377) );
  XOR U31802 ( .A(n31376), .B(n31377), .Z(n31379) );
  NANDN U31803 ( .A(n31206), .B(n31205), .Z(n31210) );
  NAND U31804 ( .A(n31208), .B(n31207), .Z(n31209) );
  NAND U31805 ( .A(n31210), .B(n31209), .Z(n31378) );
  XOR U31806 ( .A(n31379), .B(n31378), .Z(n31388) );
  XOR U31807 ( .A(n31389), .B(n31388), .Z(n31390) );
  XOR U31808 ( .A(n31391), .B(n31390), .Z(n31412) );
  XOR U31809 ( .A(n31413), .B(n31412), .Z(n31415) );
  XOR U31810 ( .A(n31414), .B(n31415), .Z(n31400) );
  NANDN U31811 ( .A(n31212), .B(n31211), .Z(n31216) );
  NAND U31812 ( .A(n31214), .B(n31213), .Z(n31215) );
  NAND U31813 ( .A(n31216), .B(n31215), .Z(n31401) );
  XOR U31814 ( .A(n31235), .B(n31234), .Z(n31236) );
  XOR U31815 ( .A(n31237), .B(n31236), .Z(n31472) );
  XNOR U31816 ( .A(n31471), .B(n31472), .Z(n31475) );
  XNOR U31817 ( .A(n31476), .B(n31475), .Z(n31478) );
  OR U31818 ( .A(n31218), .B(n31217), .Z(n31222) );
  NANDN U31819 ( .A(n31220), .B(n31219), .Z(n31221) );
  AND U31820 ( .A(n31222), .B(n31221), .Z(n31477) );
  XNOR U31821 ( .A(n31478), .B(n31477), .Z(n31228) );
  XNOR U31822 ( .A(n31229), .B(n31228), .Z(n31231) );
  XOR U31823 ( .A(n31230), .B(n31231), .Z(n31225) );
  IV U31824 ( .A(n31225), .Z(n31224) );
  XNOR U31825 ( .A(n31227), .B(n31224), .Z(n31223) );
  XNOR U31826 ( .A(n31226), .B(n31223), .Z(n31481) );
  XNOR U31827 ( .A(n31482), .B(n31481), .Z(c[201]) );
  NAND U31828 ( .A(n31229), .B(n31228), .Z(n31233) );
  NANDN U31829 ( .A(n31231), .B(n31230), .Z(n31232) );
  NAND U31830 ( .A(n31233), .B(n31232), .Z(n31486) );
  NAND U31831 ( .A(n31235), .B(n31234), .Z(n31239) );
  NANDN U31832 ( .A(n31237), .B(n31236), .Z(n31238) );
  NAND U31833 ( .A(n31239), .B(n31238), .Z(n31723) );
  OR U31834 ( .A(n31241), .B(n31240), .Z(n31245) );
  NAND U31835 ( .A(n31243), .B(n31242), .Z(n31244) );
  NAND U31836 ( .A(n31245), .B(n31244), .Z(n31713) );
  NANDN U31837 ( .A(n31247), .B(n31246), .Z(n31251) );
  NANDN U31838 ( .A(n31249), .B(n31248), .Z(n31250) );
  NAND U31839 ( .A(n31251), .B(n31250), .Z(n31506) );
  NANDN U31840 ( .A(n31253), .B(n31252), .Z(n31257) );
  OR U31841 ( .A(n31255), .B(n31254), .Z(n31256) );
  NAND U31842 ( .A(n31257), .B(n31256), .Z(n31504) );
  NANDN U31843 ( .A(n31259), .B(n31258), .Z(n31263) );
  NAND U31844 ( .A(n31261), .B(n31260), .Z(n31262) );
  NAND U31845 ( .A(n31263), .B(n31262), .Z(n31515) );
  XOR U31846 ( .A(b[49]), .B(n34851), .Z(n31568) );
  OR U31847 ( .A(n31568), .B(n37756), .Z(n31266) );
  NANDN U31848 ( .A(n31264), .B(n37652), .Z(n31265) );
  NAND U31849 ( .A(n31266), .B(n31265), .Z(n31683) );
  XNOR U31850 ( .A(b[45]), .B(a[94]), .Z(n31565) );
  NANDN U31851 ( .A(n31565), .B(n37261), .Z(n31269) );
  NANDN U31852 ( .A(n31267), .B(n37262), .Z(n31268) );
  NAND U31853 ( .A(n31269), .B(n31268), .Z(n31680) );
  NAND U31854 ( .A(n37469), .B(n31270), .Z(n31272) );
  XOR U31855 ( .A(n978), .B(n34852), .Z(n31698) );
  NAND U31856 ( .A(n31698), .B(n37471), .Z(n31271) );
  AND U31857 ( .A(n31272), .B(n31271), .Z(n31681) );
  XNOR U31858 ( .A(n31680), .B(n31681), .Z(n31682) );
  XNOR U31859 ( .A(n31683), .B(n31682), .Z(n31513) );
  XNOR U31860 ( .A(a[122]), .B(b[17]), .Z(n31562) );
  NANDN U31861 ( .A(n31562), .B(n32543), .Z(n31275) );
  NAND U31862 ( .A(n31273), .B(n32541), .Z(n31274) );
  NAND U31863 ( .A(n31275), .B(n31274), .Z(n31662) );
  XOR U31864 ( .A(a[106]), .B(n974), .Z(n31617) );
  NANDN U31865 ( .A(n31617), .B(n35620), .Z(n31278) );
  NANDN U31866 ( .A(n31276), .B(n35621), .Z(n31277) );
  NAND U31867 ( .A(n31278), .B(n31277), .Z(n31659) );
  XNOR U31868 ( .A(n36647), .B(b[35]), .Z(n31546) );
  NAND U31869 ( .A(n35985), .B(n31546), .Z(n31281) );
  NAND U31870 ( .A(n31279), .B(n35986), .Z(n31280) );
  AND U31871 ( .A(n31281), .B(n31280), .Z(n31660) );
  XNOR U31872 ( .A(n31659), .B(n31660), .Z(n31661) );
  XOR U31873 ( .A(n31662), .B(n31661), .Z(n31514) );
  XOR U31874 ( .A(n31513), .B(n31514), .Z(n31516) );
  XOR U31875 ( .A(n31515), .B(n31516), .Z(n31647) );
  NANDN U31876 ( .A(n31283), .B(n31282), .Z(n31287) );
  NAND U31877 ( .A(n31285), .B(n31284), .Z(n31286) );
  NAND U31878 ( .A(n31287), .B(n31286), .Z(n31648) );
  XNOR U31879 ( .A(n31647), .B(n31648), .Z(n31650) );
  NANDN U31880 ( .A(n31289), .B(n31288), .Z(n31293) );
  NAND U31881 ( .A(n31291), .B(n31290), .Z(n31292) );
  NAND U31882 ( .A(n31293), .B(n31292), .Z(n31520) );
  NANDN U31883 ( .A(n31295), .B(n31294), .Z(n31299) );
  NAND U31884 ( .A(n31297), .B(n31296), .Z(n31298) );
  AND U31885 ( .A(n31299), .B(n31298), .Z(n31519) );
  XNOR U31886 ( .A(n31520), .B(n31519), .Z(n31521) );
  NAND U31887 ( .A(n33283), .B(n31300), .Z(n31302) );
  XOR U31888 ( .A(n38134), .B(n33020), .Z(n31559) );
  NANDN U31889 ( .A(n33021), .B(n31559), .Z(n31301) );
  NAND U31890 ( .A(n31302), .B(n31301), .Z(n31608) );
  NAND U31891 ( .A(n35188), .B(n31303), .Z(n31305) );
  XOR U31892 ( .A(n37336), .B(n35540), .Z(n31695) );
  NANDN U31893 ( .A(n34968), .B(n31695), .Z(n31304) );
  NAND U31894 ( .A(n31305), .B(n31304), .Z(n31605) );
  XOR U31895 ( .A(a[108]), .B(n973), .Z(n31614) );
  NANDN U31896 ( .A(n31614), .B(n35313), .Z(n31308) );
  NANDN U31897 ( .A(n31306), .B(n35311), .Z(n31307) );
  AND U31898 ( .A(n31308), .B(n31307), .Z(n31606) );
  XNOR U31899 ( .A(n31605), .B(n31606), .Z(n31607) );
  XOR U31900 ( .A(n31608), .B(n31607), .Z(n31655) );
  XNOR U31901 ( .A(a[118]), .B(b[21]), .Z(n31574) );
  OR U31902 ( .A(n31574), .B(n33634), .Z(n31311) );
  NAND U31903 ( .A(n31309), .B(n33464), .Z(n31310) );
  NAND U31904 ( .A(n31311), .B(n31310), .Z(n31556) );
  XNOR U31905 ( .A(n37873), .B(b[25]), .Z(n31689) );
  NANDN U31906 ( .A(n34219), .B(n31689), .Z(n31314) );
  NAND U31907 ( .A(n31312), .B(n34217), .Z(n31313) );
  NAND U31908 ( .A(n31314), .B(n31313), .Z(n31553) );
  NAND U31909 ( .A(n34044), .B(n31315), .Z(n31317) );
  XOR U31910 ( .A(n38046), .B(n34510), .Z(n31692) );
  NANDN U31911 ( .A(n33867), .B(n31692), .Z(n31316) );
  AND U31912 ( .A(n31317), .B(n31316), .Z(n31554) );
  XNOR U31913 ( .A(n31553), .B(n31554), .Z(n31555) );
  XOR U31914 ( .A(n31556), .B(n31555), .Z(n31653) );
  NAND U31915 ( .A(n31318), .B(n34848), .Z(n31320) );
  XNOR U31916 ( .A(n37583), .B(b[27]), .Z(n31665) );
  NAND U31917 ( .A(n34618), .B(n31665), .Z(n31319) );
  NAND U31918 ( .A(n31320), .B(n31319), .Z(n31654) );
  XNOR U31919 ( .A(n31653), .B(n31654), .Z(n31656) );
  XNOR U31920 ( .A(n31655), .B(n31656), .Z(n31522) );
  XNOR U31921 ( .A(n31521), .B(n31522), .Z(n31649) );
  XNOR U31922 ( .A(n31650), .B(n31649), .Z(n31503) );
  XOR U31923 ( .A(n31504), .B(n31503), .Z(n31505) );
  XNOR U31924 ( .A(n31506), .B(n31505), .Z(n31644) );
  XOR U31925 ( .A(b[43]), .B(n35545), .Z(n31537) );
  NANDN U31926 ( .A(n31537), .B(n37068), .Z(n31323) );
  NANDN U31927 ( .A(n31321), .B(n37069), .Z(n31322) );
  NAND U31928 ( .A(n31323), .B(n31322), .Z(n31534) );
  XOR U31929 ( .A(b[51]), .B(n34048), .Z(n31701) );
  NANDN U31930 ( .A(n31701), .B(n37803), .Z(n31326) );
  NANDN U31931 ( .A(n31324), .B(n37802), .Z(n31325) );
  NAND U31932 ( .A(n31326), .B(n31325), .Z(n31531) );
  XOR U31933 ( .A(b[53]), .B(n33628), .Z(n31668) );
  NANDN U31934 ( .A(n31668), .B(n37940), .Z(n31329) );
  NANDN U31935 ( .A(n31327), .B(n37941), .Z(n31328) );
  AND U31936 ( .A(n31329), .B(n31328), .Z(n31532) );
  XNOR U31937 ( .A(n31531), .B(n31532), .Z(n31533) );
  XNOR U31938 ( .A(n31534), .B(n31533), .Z(n31586) );
  XOR U31939 ( .A(b[55]), .B(n33185), .Z(n31671) );
  NANDN U31940 ( .A(n31671), .B(n38075), .Z(n31332) );
  NANDN U31941 ( .A(n31330), .B(n38073), .Z(n31331) );
  NAND U31942 ( .A(n31332), .B(n31331), .Z(n31602) );
  XOR U31943 ( .A(a[124]), .B(n972), .Z(n31540) );
  OR U31944 ( .A(n31540), .B(n32010), .Z(n31335) );
  NANDN U31945 ( .A(n31333), .B(n32011), .Z(n31334) );
  NAND U31946 ( .A(n31335), .B(n31334), .Z(n31599) );
  XOR U31947 ( .A(b[37]), .B(n36420), .Z(n31620) );
  NANDN U31948 ( .A(n31620), .B(n36311), .Z(n31338) );
  NANDN U31949 ( .A(n31336), .B(n36309), .Z(n31337) );
  AND U31950 ( .A(n31338), .B(n31337), .Z(n31600) );
  XNOR U31951 ( .A(n31599), .B(n31600), .Z(n31601) );
  XNOR U31952 ( .A(n31602), .B(n31601), .Z(n31583) );
  NANDN U31953 ( .A(n31340), .B(n31339), .Z(n31344) );
  NAND U31954 ( .A(n31342), .B(n31341), .Z(n31343) );
  NAND U31955 ( .A(n31344), .B(n31343), .Z(n31584) );
  XNOR U31956 ( .A(n31583), .B(n31584), .Z(n31585) );
  XOR U31957 ( .A(n31586), .B(n31585), .Z(n31637) );
  NANDN U31958 ( .A(n31346), .B(n31345), .Z(n31350) );
  NAND U31959 ( .A(n31348), .B(n31347), .Z(n31349) );
  NAND U31960 ( .A(n31350), .B(n31349), .Z(n31636) );
  NANDN U31961 ( .A(n31352), .B(n31351), .Z(n31356) );
  NAND U31962 ( .A(n31354), .B(n31353), .Z(n31355) );
  NAND U31963 ( .A(n31356), .B(n31355), .Z(n31579) );
  XNOR U31964 ( .A(b[41]), .B(a[98]), .Z(n31611) );
  OR U31965 ( .A(n31611), .B(n36905), .Z(n31359) );
  NAND U31966 ( .A(n31357), .B(n36807), .Z(n31358) );
  NAND U31967 ( .A(n31359), .B(n31358), .Z(n31596) );
  XOR U31968 ( .A(b[61]), .B(n31870), .Z(n31543) );
  OR U31969 ( .A(n31543), .B(n38371), .Z(n31362) );
  NANDN U31970 ( .A(n31360), .B(n38369), .Z(n31361) );
  NAND U31971 ( .A(n31362), .B(n31361), .Z(n31593) );
  XOR U31972 ( .A(b[63]), .B(n31363), .Z(n31623) );
  NANDN U31973 ( .A(n31623), .B(n38422), .Z(n31366) );
  NANDN U31974 ( .A(n31364), .B(n38423), .Z(n31365) );
  AND U31975 ( .A(n31366), .B(n31365), .Z(n31594) );
  XNOR U31976 ( .A(n31593), .B(n31594), .Z(n31595) );
  XNOR U31977 ( .A(n31596), .B(n31595), .Z(n31577) );
  XOR U31978 ( .A(n970), .B(n31367), .Z(n31371) );
  NAND U31979 ( .A(n31369), .B(n31368), .Z(n31370) );
  AND U31980 ( .A(n31371), .B(n31370), .Z(n31675) );
  ANDN U31981 ( .B(b[63]), .A(n31372), .Z(n31674) );
  XNOR U31982 ( .A(n31675), .B(n31674), .Z(n31676) );
  NAND U31983 ( .A(n31874), .B(n31373), .Z(n31375) );
  XOR U31984 ( .A(n987), .B(n971), .Z(n31549) );
  NANDN U31985 ( .A(n31550), .B(n31549), .Z(n31374) );
  AND U31986 ( .A(n31375), .B(n31374), .Z(n31677) );
  XNOR U31987 ( .A(n31676), .B(n31677), .Z(n31578) );
  XOR U31988 ( .A(n31577), .B(n31578), .Z(n31580) );
  XOR U31989 ( .A(n31579), .B(n31580), .Z(n31635) );
  XOR U31990 ( .A(n31636), .B(n31635), .Z(n31638) );
  XOR U31991 ( .A(n31637), .B(n31638), .Z(n31704) );
  NANDN U31992 ( .A(n31377), .B(n31376), .Z(n31381) );
  OR U31993 ( .A(n31379), .B(n31378), .Z(n31380) );
  NAND U31994 ( .A(n31381), .B(n31380), .Z(n31705) );
  XNOR U31995 ( .A(n31704), .B(n31705), .Z(n31706) );
  OR U31996 ( .A(n31383), .B(n31382), .Z(n31387) );
  OR U31997 ( .A(n31385), .B(n31384), .Z(n31386) );
  NAND U31998 ( .A(n31387), .B(n31386), .Z(n31707) );
  XOR U31999 ( .A(n31706), .B(n31707), .Z(n31641) );
  OR U32000 ( .A(n31389), .B(n31388), .Z(n31393) );
  NAND U32001 ( .A(n31391), .B(n31390), .Z(n31392) );
  NAND U32002 ( .A(n31393), .B(n31392), .Z(n31642) );
  XNOR U32003 ( .A(n31641), .B(n31642), .Z(n31643) );
  XOR U32004 ( .A(n31644), .B(n31643), .Z(n31710) );
  NANDN U32005 ( .A(n31395), .B(n31394), .Z(n31399) );
  NAND U32006 ( .A(n31397), .B(n31396), .Z(n31398) );
  NAND U32007 ( .A(n31399), .B(n31398), .Z(n31711) );
  XOR U32008 ( .A(n31710), .B(n31711), .Z(n31712) );
  XNOR U32009 ( .A(n31713), .B(n31712), .Z(n31718) );
  OR U32010 ( .A(n31401), .B(n31400), .Z(n31405) );
  NANDN U32011 ( .A(n31403), .B(n31402), .Z(n31404) );
  NAND U32012 ( .A(n31405), .B(n31404), .Z(n31717) );
  OR U32013 ( .A(n31407), .B(n31406), .Z(n31411) );
  NANDN U32014 ( .A(n31409), .B(n31408), .Z(n31410) );
  NAND U32015 ( .A(n31411), .B(n31410), .Z(n31497) );
  NANDN U32016 ( .A(n31413), .B(n31412), .Z(n31417) );
  OR U32017 ( .A(n31415), .B(n31414), .Z(n31416) );
  NAND U32018 ( .A(n31417), .B(n31416), .Z(n31498) );
  XNOR U32019 ( .A(n31497), .B(n31498), .Z(n31499) );
  NANDN U32020 ( .A(n31419), .B(n31418), .Z(n31423) );
  NANDN U32021 ( .A(n31421), .B(n31420), .Z(n31422) );
  NAND U32022 ( .A(n31423), .B(n31422), .Z(n31512) );
  NANDN U32023 ( .A(n31425), .B(n31424), .Z(n31429) );
  NAND U32024 ( .A(n31427), .B(n31426), .Z(n31428) );
  NAND U32025 ( .A(n31429), .B(n31428), .Z(n31632) );
  NANDN U32026 ( .A(n31431), .B(n31430), .Z(n31435) );
  NAND U32027 ( .A(n31433), .B(n31432), .Z(n31434) );
  NAND U32028 ( .A(n31435), .B(n31434), .Z(n31629) );
  NANDN U32029 ( .A(n31437), .B(n31436), .Z(n31441) );
  NAND U32030 ( .A(n31439), .B(n31438), .Z(n31440) );
  NAND U32031 ( .A(n31441), .B(n31440), .Z(n31590) );
  OR U32032 ( .A(n31443), .B(n31442), .Z(n31447) );
  NAND U32033 ( .A(n31445), .B(n31444), .Z(n31446) );
  NAND U32034 ( .A(n31447), .B(n31446), .Z(n31587) );
  XOR U32035 ( .A(b[57]), .B(n32815), .Z(n31686) );
  OR U32036 ( .A(n31686), .B(n965), .Z(n31450) );
  NANDN U32037 ( .A(n31448), .B(n38194), .Z(n31449) );
  NAND U32038 ( .A(n31450), .B(n31449), .Z(n31528) );
  NAND U32039 ( .A(n38326), .B(n31451), .Z(n31453) );
  XOR U32040 ( .A(n38400), .B(n32814), .Z(n31571) );
  NANDN U32041 ( .A(n38273), .B(n31571), .Z(n31452) );
  NAND U32042 ( .A(n31453), .B(n31452), .Z(n31525) );
  XOR U32043 ( .A(n976), .B(n36100), .Z(n31626) );
  NAND U32044 ( .A(n31626), .B(n36553), .Z(n31456) );
  NANDN U32045 ( .A(n31454), .B(n36643), .Z(n31455) );
  AND U32046 ( .A(n31456), .B(n31455), .Z(n31526) );
  XNOR U32047 ( .A(n31525), .B(n31526), .Z(n31527) );
  XNOR U32048 ( .A(n31528), .B(n31527), .Z(n31588) );
  XNOR U32049 ( .A(n31587), .B(n31588), .Z(n31589) );
  XNOR U32050 ( .A(n31590), .B(n31589), .Z(n31630) );
  XNOR U32051 ( .A(n31629), .B(n31630), .Z(n31631) );
  XNOR U32052 ( .A(n31632), .B(n31631), .Z(n31509) );
  NANDN U32053 ( .A(n31458), .B(n31457), .Z(n31462) );
  OR U32054 ( .A(n31460), .B(n31459), .Z(n31461) );
  AND U32055 ( .A(n31462), .B(n31461), .Z(n31510) );
  XNOR U32056 ( .A(n31509), .B(n31510), .Z(n31511) );
  XNOR U32057 ( .A(n31512), .B(n31511), .Z(n31500) );
  XNOR U32058 ( .A(n31499), .B(n31500), .Z(n31716) );
  XNOR U32059 ( .A(n31717), .B(n31716), .Z(n31719) );
  XNOR U32060 ( .A(n31718), .B(n31719), .Z(n31722) );
  XNOR U32061 ( .A(n31723), .B(n31722), .Z(n31725) );
  NANDN U32062 ( .A(n31464), .B(n31463), .Z(n31468) );
  NAND U32063 ( .A(n31466), .B(n31465), .Z(n31467) );
  NAND U32064 ( .A(n31468), .B(n31467), .Z(n31724) );
  XNOR U32065 ( .A(n31725), .B(n31724), .Z(n31491) );
  NANDN U32066 ( .A(n31470), .B(n31469), .Z(n31474) );
  NANDN U32067 ( .A(n31472), .B(n31471), .Z(n31473) );
  NAND U32068 ( .A(n31474), .B(n31473), .Z(n31492) );
  XNOR U32069 ( .A(n31491), .B(n31492), .Z(n31493) );
  NAND U32070 ( .A(n31476), .B(n31475), .Z(n31480) );
  NANDN U32071 ( .A(n31478), .B(n31477), .Z(n31479) );
  AND U32072 ( .A(n31480), .B(n31479), .Z(n31494) );
  XOR U32073 ( .A(n31493), .B(n31494), .Z(n31485) );
  XOR U32074 ( .A(n31486), .B(n31485), .Z(n31488) );
  XNOR U32075 ( .A(n31487), .B(n31488), .Z(n31483) );
  NANDN U32076 ( .A(n31482), .B(n31481), .Z(n31484) );
  XNOR U32077 ( .A(n31483), .B(n31484), .Z(c[202]) );
  NANDN U32078 ( .A(n31484), .B(n31483), .Z(n31730) );
  NANDN U32079 ( .A(n31486), .B(n31485), .Z(n31490) );
  NANDN U32080 ( .A(n31488), .B(n31487), .Z(n31489) );
  NAND U32081 ( .A(n31490), .B(n31489), .Z(n31733) );
  NANDN U32082 ( .A(n31492), .B(n31491), .Z(n31496) );
  NAND U32083 ( .A(n31494), .B(n31493), .Z(n31495) );
  AND U32084 ( .A(n31496), .B(n31495), .Z(n31732) );
  NANDN U32085 ( .A(n31498), .B(n31497), .Z(n31502) );
  NANDN U32086 ( .A(n31500), .B(n31499), .Z(n31501) );
  NAND U32087 ( .A(n31502), .B(n31501), .Z(n31969) );
  OR U32088 ( .A(n31504), .B(n31503), .Z(n31508) );
  NAND U32089 ( .A(n31506), .B(n31505), .Z(n31507) );
  NAND U32090 ( .A(n31508), .B(n31507), .Z(n31749) );
  NANDN U32091 ( .A(n31514), .B(n31513), .Z(n31518) );
  OR U32092 ( .A(n31516), .B(n31515), .Z(n31517) );
  NAND U32093 ( .A(n31518), .B(n31517), .Z(n31807) );
  NANDN U32094 ( .A(n31520), .B(n31519), .Z(n31524) );
  NANDN U32095 ( .A(n31522), .B(n31521), .Z(n31523) );
  NAND U32096 ( .A(n31524), .B(n31523), .Z(n31804) );
  NANDN U32097 ( .A(n31526), .B(n31525), .Z(n31530) );
  NAND U32098 ( .A(n31528), .B(n31527), .Z(n31529) );
  AND U32099 ( .A(n31530), .B(n31529), .Z(n31816) );
  NANDN U32100 ( .A(n31532), .B(n31531), .Z(n31536) );
  NAND U32101 ( .A(n31534), .B(n31533), .Z(n31535) );
  NAND U32102 ( .A(n31536), .B(n31535), .Z(n31959) );
  XNOR U32103 ( .A(b[43]), .B(a[97]), .Z(n31864) );
  NANDN U32104 ( .A(n31864), .B(n37068), .Z(n31539) );
  NANDN U32105 ( .A(n31537), .B(n37069), .Z(n31538) );
  NAND U32106 ( .A(n31539), .B(n31538), .Z(n31887) );
  XNOR U32107 ( .A(a[125]), .B(b[15]), .Z(n31941) );
  OR U32108 ( .A(n31941), .B(n32010), .Z(n31542) );
  NANDN U32109 ( .A(n31540), .B(n32011), .Z(n31541) );
  NAND U32110 ( .A(n31542), .B(n31541), .Z(n31884) );
  XNOR U32111 ( .A(b[61]), .B(a[79]), .Z(n31932) );
  OR U32112 ( .A(n31932), .B(n38371), .Z(n31545) );
  NANDN U32113 ( .A(n31543), .B(n38369), .Z(n31544) );
  AND U32114 ( .A(n31545), .B(n31544), .Z(n31885) );
  XNOR U32115 ( .A(n31884), .B(n31885), .Z(n31886) );
  XNOR U32116 ( .A(n31887), .B(n31886), .Z(n31957) );
  NAND U32117 ( .A(n35986), .B(n31546), .Z(n31548) );
  XOR U32118 ( .A(a[105]), .B(b[35]), .Z(n31831) );
  NAND U32119 ( .A(n35985), .B(n31831), .Z(n31547) );
  AND U32120 ( .A(n31548), .B(n31547), .Z(n31891) );
  XNOR U32121 ( .A(n31890), .B(n31891), .Z(n31893) );
  NAND U32122 ( .A(n31874), .B(n31549), .Z(n31552) );
  XOR U32123 ( .A(a[127]), .B(n971), .Z(n31875) );
  OR U32124 ( .A(n31875), .B(n31550), .Z(n31551) );
  AND U32125 ( .A(n31552), .B(n31551), .Z(n31892) );
  XNOR U32126 ( .A(n31893), .B(n31892), .Z(n31956) );
  XOR U32127 ( .A(n31957), .B(n31956), .Z(n31958) );
  XNOR U32128 ( .A(n31959), .B(n31958), .Z(n31817) );
  NANDN U32129 ( .A(n31554), .B(n31553), .Z(n31558) );
  NAND U32130 ( .A(n31556), .B(n31555), .Z(n31557) );
  NAND U32131 ( .A(n31558), .B(n31557), .Z(n31776) );
  NAND U32132 ( .A(n33283), .B(n31559), .Z(n31561) );
  XNOR U32133 ( .A(a[121]), .B(n33020), .Z(n31929) );
  NANDN U32134 ( .A(n33021), .B(n31929), .Z(n31560) );
  NAND U32135 ( .A(n31561), .B(n31560), .Z(n31846) );
  XOR U32136 ( .A(a[123]), .B(b[17]), .Z(n31938) );
  NAND U32137 ( .A(n31938), .B(n32543), .Z(n31564) );
  NANDN U32138 ( .A(n31562), .B(n32541), .Z(n31563) );
  NAND U32139 ( .A(n31564), .B(n31563), .Z(n31843) );
  XNOR U32140 ( .A(b[45]), .B(a[95]), .Z(n31926) );
  NANDN U32141 ( .A(n31926), .B(n37261), .Z(n31567) );
  NANDN U32142 ( .A(n31565), .B(n37262), .Z(n31566) );
  AND U32143 ( .A(n31567), .B(n31566), .Z(n31844) );
  XNOR U32144 ( .A(n31843), .B(n31844), .Z(n31845) );
  XNOR U32145 ( .A(n31846), .B(n31845), .Z(n31774) );
  XNOR U32146 ( .A(b[49]), .B(a[91]), .Z(n31867) );
  OR U32147 ( .A(n31867), .B(n37756), .Z(n31570) );
  NANDN U32148 ( .A(n31568), .B(n37652), .Z(n31569) );
  NAND U32149 ( .A(n31570), .B(n31569), .Z(n31917) );
  NAND U32150 ( .A(n38326), .B(n31571), .Z(n31573) );
  XNOR U32151 ( .A(n38400), .B(a[81]), .Z(n31795) );
  NANDN U32152 ( .A(n38273), .B(n31795), .Z(n31572) );
  NAND U32153 ( .A(n31573), .B(n31572), .Z(n31914) );
  XNOR U32154 ( .A(a[119]), .B(b[21]), .Z(n31911) );
  OR U32155 ( .A(n31911), .B(n33634), .Z(n31576) );
  NANDN U32156 ( .A(n31574), .B(n33464), .Z(n31575) );
  AND U32157 ( .A(n31576), .B(n31575), .Z(n31915) );
  XNOR U32158 ( .A(n31914), .B(n31915), .Z(n31916) );
  XOR U32159 ( .A(n31917), .B(n31916), .Z(n31775) );
  XOR U32160 ( .A(n31774), .B(n31775), .Z(n31777) );
  XNOR U32161 ( .A(n31776), .B(n31777), .Z(n31819) );
  XOR U32162 ( .A(n31818), .B(n31819), .Z(n31767) );
  NANDN U32163 ( .A(n31578), .B(n31577), .Z(n31582) );
  OR U32164 ( .A(n31580), .B(n31579), .Z(n31581) );
  NAND U32165 ( .A(n31582), .B(n31581), .Z(n31764) );
  XNOR U32166 ( .A(n31764), .B(n31765), .Z(n31766) );
  XOR U32167 ( .A(n31767), .B(n31766), .Z(n31805) );
  XNOR U32168 ( .A(n31804), .B(n31805), .Z(n31806) );
  XNOR U32169 ( .A(n31807), .B(n31806), .Z(n31755) );
  NANDN U32170 ( .A(n31588), .B(n31587), .Z(n31592) );
  NAND U32171 ( .A(n31590), .B(n31589), .Z(n31591) );
  NAND U32172 ( .A(n31592), .B(n31591), .Z(n31811) );
  NANDN U32173 ( .A(n31594), .B(n31593), .Z(n31598) );
  NAND U32174 ( .A(n31596), .B(n31595), .Z(n31597) );
  NAND U32175 ( .A(n31598), .B(n31597), .Z(n31946) );
  NANDN U32176 ( .A(n31600), .B(n31599), .Z(n31604) );
  NAND U32177 ( .A(n31602), .B(n31601), .Z(n31603) );
  NAND U32178 ( .A(n31604), .B(n31603), .Z(n31945) );
  NANDN U32179 ( .A(n31606), .B(n31605), .Z(n31610) );
  NAND U32180 ( .A(n31608), .B(n31607), .Z(n31609) );
  NAND U32181 ( .A(n31610), .B(n31609), .Z(n31770) );
  XOR U32182 ( .A(b[41]), .B(a[99]), .Z(n31935) );
  NANDN U32183 ( .A(n36905), .B(n31935), .Z(n31613) );
  NANDN U32184 ( .A(n31611), .B(n36807), .Z(n31612) );
  NAND U32185 ( .A(n31613), .B(n31612), .Z(n31881) );
  XNOR U32186 ( .A(a[109]), .B(b[31]), .Z(n31861) );
  NANDN U32187 ( .A(n31861), .B(n35313), .Z(n31616) );
  NANDN U32188 ( .A(n31614), .B(n35311), .Z(n31615) );
  NAND U32189 ( .A(n31616), .B(n31615), .Z(n31878) );
  XNOR U32190 ( .A(a[107]), .B(n974), .Z(n31834) );
  NAND U32191 ( .A(n35620), .B(n31834), .Z(n31619) );
  NANDN U32192 ( .A(n31617), .B(n35621), .Z(n31618) );
  AND U32193 ( .A(n31619), .B(n31618), .Z(n31879) );
  XNOR U32194 ( .A(n31878), .B(n31879), .Z(n31880) );
  XNOR U32195 ( .A(n31881), .B(n31880), .Z(n31768) );
  XNOR U32196 ( .A(b[37]), .B(a[103]), .Z(n31902) );
  NANDN U32197 ( .A(n31902), .B(n36311), .Z(n31622) );
  NANDN U32198 ( .A(n31620), .B(n36309), .Z(n31621) );
  NAND U32199 ( .A(n31622), .B(n31621), .Z(n31837) );
  NANDN U32200 ( .A(n985), .B(a[75]), .Z(n31838) );
  XNOR U32201 ( .A(n31837), .B(n31838), .Z(n31839) );
  XOR U32202 ( .A(n31674), .B(n31839), .Z(n31850) );
  XNOR U32203 ( .A(n985), .B(a[77]), .Z(n31871) );
  NAND U32204 ( .A(n31871), .B(n38422), .Z(n31625) );
  NANDN U32205 ( .A(n31623), .B(n38423), .Z(n31624) );
  NAND U32206 ( .A(n31625), .B(n31624), .Z(n31849) );
  XOR U32207 ( .A(n31850), .B(n31849), .Z(n31851) );
  NAND U32208 ( .A(n36643), .B(n31626), .Z(n31628) );
  XNOR U32209 ( .A(n976), .B(a[101]), .Z(n31828) );
  NAND U32210 ( .A(n31828), .B(n36553), .Z(n31627) );
  AND U32211 ( .A(n31628), .B(n31627), .Z(n31852) );
  XNOR U32212 ( .A(n31851), .B(n31852), .Z(n31769) );
  XOR U32213 ( .A(n31768), .B(n31769), .Z(n31771) );
  XOR U32214 ( .A(n31770), .B(n31771), .Z(n31944) );
  XOR U32215 ( .A(n31945), .B(n31944), .Z(n31947) );
  XOR U32216 ( .A(n31946), .B(n31947), .Z(n31810) );
  XOR U32217 ( .A(n31811), .B(n31810), .Z(n31813) );
  NANDN U32218 ( .A(n31630), .B(n31629), .Z(n31634) );
  NAND U32219 ( .A(n31632), .B(n31631), .Z(n31633) );
  NAND U32220 ( .A(n31634), .B(n31633), .Z(n31812) );
  XNOR U32221 ( .A(n31813), .B(n31812), .Z(n31752) );
  NANDN U32222 ( .A(n31636), .B(n31635), .Z(n31640) );
  NANDN U32223 ( .A(n31638), .B(n31637), .Z(n31639) );
  NAND U32224 ( .A(n31640), .B(n31639), .Z(n31753) );
  XNOR U32225 ( .A(n31752), .B(n31753), .Z(n31754) );
  XOR U32226 ( .A(n31755), .B(n31754), .Z(n31747) );
  XNOR U32227 ( .A(n31746), .B(n31747), .Z(n31748) );
  XOR U32228 ( .A(n31749), .B(n31748), .Z(n31965) );
  NANDN U32229 ( .A(n31642), .B(n31641), .Z(n31646) );
  NAND U32230 ( .A(n31644), .B(n31643), .Z(n31645) );
  NAND U32231 ( .A(n31646), .B(n31645), .Z(n31963) );
  OR U32232 ( .A(n31648), .B(n31647), .Z(n31652) );
  OR U32233 ( .A(n31650), .B(n31649), .Z(n31651) );
  NAND U32234 ( .A(n31652), .B(n31651), .Z(n31743) );
  OR U32235 ( .A(n31654), .B(n31653), .Z(n31658) );
  OR U32236 ( .A(n31656), .B(n31655), .Z(n31657) );
  NAND U32237 ( .A(n31658), .B(n31657), .Z(n31759) );
  NANDN U32238 ( .A(n31660), .B(n31659), .Z(n31664) );
  NAND U32239 ( .A(n31662), .B(n31661), .Z(n31663) );
  NAND U32240 ( .A(n31664), .B(n31663), .Z(n31952) );
  NAND U32241 ( .A(n31665), .B(n34848), .Z(n31667) );
  XNOR U32242 ( .A(a[113]), .B(n35375), .Z(n31899) );
  NAND U32243 ( .A(n34618), .B(n31899), .Z(n31666) );
  NAND U32244 ( .A(n31667), .B(n31666), .Z(n31783) );
  XNOR U32245 ( .A(b[53]), .B(a[87]), .Z(n31789) );
  NANDN U32246 ( .A(n31789), .B(n37940), .Z(n31670) );
  NANDN U32247 ( .A(n31668), .B(n37941), .Z(n31669) );
  NAND U32248 ( .A(n31670), .B(n31669), .Z(n31780) );
  XNOR U32249 ( .A(b[55]), .B(a[85]), .Z(n31792) );
  NANDN U32250 ( .A(n31792), .B(n38075), .Z(n31673) );
  NANDN U32251 ( .A(n31671), .B(n38073), .Z(n31672) );
  AND U32252 ( .A(n31673), .B(n31672), .Z(n31781) );
  XNOR U32253 ( .A(n31780), .B(n31781), .Z(n31782) );
  XNOR U32254 ( .A(n31783), .B(n31782), .Z(n31950) );
  IV U32255 ( .A(n31674), .Z(n31840) );
  OR U32256 ( .A(n31675), .B(n31840), .Z(n31679) );
  NAND U32257 ( .A(n31677), .B(n31676), .Z(n31678) );
  AND U32258 ( .A(n31679), .B(n31678), .Z(n31951) );
  XOR U32259 ( .A(n31950), .B(n31951), .Z(n31953) );
  XOR U32260 ( .A(n31952), .B(n31953), .Z(n31758) );
  XNOR U32261 ( .A(n31759), .B(n31758), .Z(n31761) );
  NANDN U32262 ( .A(n31681), .B(n31680), .Z(n31685) );
  NAND U32263 ( .A(n31683), .B(n31682), .Z(n31684) );
  NAND U32264 ( .A(n31685), .B(n31684), .Z(n31857) );
  XNOR U32265 ( .A(b[57]), .B(a[83]), .Z(n31896) );
  OR U32266 ( .A(n31896), .B(n965), .Z(n31688) );
  NANDN U32267 ( .A(n31686), .B(n38194), .Z(n31687) );
  NAND U32268 ( .A(n31688), .B(n31687), .Z(n31923) );
  XOR U32269 ( .A(a[115]), .B(b[25]), .Z(n31798) );
  NANDN U32270 ( .A(n34219), .B(n31798), .Z(n31691) );
  NAND U32271 ( .A(n34217), .B(n31689), .Z(n31690) );
  NAND U32272 ( .A(n31691), .B(n31690), .Z(n31920) );
  NAND U32273 ( .A(n34044), .B(n31692), .Z(n31694) );
  XNOR U32274 ( .A(a[117]), .B(n34510), .Z(n31908) );
  NANDN U32275 ( .A(n33867), .B(n31908), .Z(n31693) );
  AND U32276 ( .A(n31694), .B(n31693), .Z(n31921) );
  XNOR U32277 ( .A(n31920), .B(n31921), .Z(n31922) );
  XNOR U32278 ( .A(n31923), .B(n31922), .Z(n31855) );
  NAND U32279 ( .A(n35188), .B(n31695), .Z(n31697) );
  XNOR U32280 ( .A(a[111]), .B(n35540), .Z(n31786) );
  NANDN U32281 ( .A(n34968), .B(n31786), .Z(n31696) );
  NAND U32282 ( .A(n31697), .B(n31696), .Z(n31825) );
  NAND U32283 ( .A(n37469), .B(n31698), .Z(n31700) );
  XOR U32284 ( .A(n978), .B(n35377), .Z(n31905) );
  NAND U32285 ( .A(n31905), .B(n37471), .Z(n31699) );
  NAND U32286 ( .A(n31700), .B(n31699), .Z(n31822) );
  XNOR U32287 ( .A(b[51]), .B(a[89]), .Z(n31801) );
  NANDN U32288 ( .A(n31801), .B(n37803), .Z(n31703) );
  NANDN U32289 ( .A(n31701), .B(n37802), .Z(n31702) );
  AND U32290 ( .A(n31703), .B(n31702), .Z(n31823) );
  XNOR U32291 ( .A(n31822), .B(n31823), .Z(n31824) );
  XOR U32292 ( .A(n31825), .B(n31824), .Z(n31856) );
  XOR U32293 ( .A(n31855), .B(n31856), .Z(n31858) );
  XOR U32294 ( .A(n31857), .B(n31858), .Z(n31760) );
  XOR U32295 ( .A(n31761), .B(n31760), .Z(n31740) );
  NANDN U32296 ( .A(n31705), .B(n31704), .Z(n31709) );
  NANDN U32297 ( .A(n31707), .B(n31706), .Z(n31708) );
  AND U32298 ( .A(n31709), .B(n31708), .Z(n31741) );
  XNOR U32299 ( .A(n31740), .B(n31741), .Z(n31742) );
  XOR U32300 ( .A(n31743), .B(n31742), .Z(n31962) );
  XNOR U32301 ( .A(n31963), .B(n31962), .Z(n31964) );
  XNOR U32302 ( .A(n31965), .B(n31964), .Z(n31966) );
  OR U32303 ( .A(n31711), .B(n31710), .Z(n31715) );
  NAND U32304 ( .A(n31713), .B(n31712), .Z(n31714) );
  NAND U32305 ( .A(n31715), .B(n31714), .Z(n31967) );
  XNOR U32306 ( .A(n31966), .B(n31967), .Z(n31968) );
  XNOR U32307 ( .A(n31969), .B(n31968), .Z(n31737) );
  NAND U32308 ( .A(n31717), .B(n31716), .Z(n31721) );
  NANDN U32309 ( .A(n31719), .B(n31718), .Z(n31720) );
  NAND U32310 ( .A(n31721), .B(n31720), .Z(n31735) );
  NAND U32311 ( .A(n31723), .B(n31722), .Z(n31727) );
  OR U32312 ( .A(n31725), .B(n31724), .Z(n31726) );
  AND U32313 ( .A(n31727), .B(n31726), .Z(n31734) );
  XNOR U32314 ( .A(n31735), .B(n31734), .Z(n31736) );
  XOR U32315 ( .A(n31737), .B(n31736), .Z(n31731) );
  XNOR U32316 ( .A(n31732), .B(n31731), .Z(n31728) );
  XOR U32317 ( .A(n31733), .B(n31728), .Z(n31729) );
  XNOR U32318 ( .A(n31730), .B(n31729), .Z(c[203]) );
  NANDN U32319 ( .A(n31730), .B(n31729), .Z(n32209) );
  NANDN U32320 ( .A(n31735), .B(n31734), .Z(n31739) );
  NAND U32321 ( .A(n31737), .B(n31736), .Z(n31738) );
  NAND U32322 ( .A(n31739), .B(n31738), .Z(n31974) );
  NANDN U32323 ( .A(n31741), .B(n31740), .Z(n31745) );
  NAND U32324 ( .A(n31743), .B(n31742), .Z(n31744) );
  NAND U32325 ( .A(n31745), .B(n31744), .Z(n32205) );
  NANDN U32326 ( .A(n31747), .B(n31746), .Z(n31751) );
  NANDN U32327 ( .A(n31749), .B(n31748), .Z(n31750) );
  NAND U32328 ( .A(n31751), .B(n31750), .Z(n32203) );
  NANDN U32329 ( .A(n31753), .B(n31752), .Z(n31757) );
  NAND U32330 ( .A(n31755), .B(n31754), .Z(n31756) );
  NAND U32331 ( .A(n31757), .B(n31756), .Z(n32199) );
  NAND U32332 ( .A(n31759), .B(n31758), .Z(n31763) );
  NANDN U32333 ( .A(n31761), .B(n31760), .Z(n31762) );
  NAND U32334 ( .A(n31763), .B(n31762), .Z(n32050) );
  XNOR U32335 ( .A(n32050), .B(n32051), .Z(n32052) );
  NANDN U32336 ( .A(n31769), .B(n31768), .Z(n31773) );
  OR U32337 ( .A(n31771), .B(n31770), .Z(n31772) );
  NAND U32338 ( .A(n31773), .B(n31772), .Z(n32041) );
  NANDN U32339 ( .A(n31775), .B(n31774), .Z(n31779) );
  OR U32340 ( .A(n31777), .B(n31776), .Z(n31778) );
  NAND U32341 ( .A(n31779), .B(n31778), .Z(n32038) );
  NANDN U32342 ( .A(n31781), .B(n31780), .Z(n31785) );
  NAND U32343 ( .A(n31783), .B(n31782), .Z(n31784) );
  NAND U32344 ( .A(n31785), .B(n31784), .Z(n32065) );
  NAND U32345 ( .A(n35188), .B(n31786), .Z(n31788) );
  XOR U32346 ( .A(n37583), .B(n35540), .Z(n32026) );
  NANDN U32347 ( .A(n34968), .B(n32026), .Z(n31787) );
  NAND U32348 ( .A(n31788), .B(n31787), .Z(n32077) );
  XOR U32349 ( .A(b[53]), .B(n34048), .Z(n32165) );
  NANDN U32350 ( .A(n32165), .B(n37940), .Z(n31791) );
  NANDN U32351 ( .A(n31789), .B(n37941), .Z(n31790) );
  NAND U32352 ( .A(n31791), .B(n31790), .Z(n32074) );
  XOR U32353 ( .A(b[55]), .B(n33628), .Z(n32107) );
  NANDN U32354 ( .A(n32107), .B(n38075), .Z(n31794) );
  NANDN U32355 ( .A(n31792), .B(n38073), .Z(n31793) );
  AND U32356 ( .A(n31794), .B(n31793), .Z(n32075) );
  XNOR U32357 ( .A(n32074), .B(n32075), .Z(n32076) );
  XOR U32358 ( .A(n32077), .B(n32076), .Z(n32063) );
  NAND U32359 ( .A(n38326), .B(n31795), .Z(n31797) );
  XOR U32360 ( .A(n38400), .B(n32815), .Z(n32092) );
  NANDN U32361 ( .A(n38273), .B(n32092), .Z(n31796) );
  NAND U32362 ( .A(n31797), .B(n31796), .Z(n32101) );
  XNOR U32363 ( .A(n38046), .B(b[25]), .Z(n32159) );
  NANDN U32364 ( .A(n34219), .B(n32159), .Z(n31800) );
  NAND U32365 ( .A(n34217), .B(n31798), .Z(n31799) );
  NAND U32366 ( .A(n31800), .B(n31799), .Z(n32098) );
  XOR U32367 ( .A(b[51]), .B(n34851), .Z(n32095) );
  NANDN U32368 ( .A(n32095), .B(n37803), .Z(n31803) );
  NANDN U32369 ( .A(n31801), .B(n37802), .Z(n31802) );
  AND U32370 ( .A(n31803), .B(n31802), .Z(n32099) );
  XNOR U32371 ( .A(n32098), .B(n32099), .Z(n32100) );
  XNOR U32372 ( .A(n32101), .B(n32100), .Z(n32062) );
  XOR U32373 ( .A(n32063), .B(n32062), .Z(n32064) );
  XNOR U32374 ( .A(n32065), .B(n32064), .Z(n32039) );
  XNOR U32375 ( .A(n32038), .B(n32039), .Z(n32040) );
  XOR U32376 ( .A(n32041), .B(n32040), .Z(n32053) );
  XOR U32377 ( .A(n32052), .B(n32053), .Z(n32198) );
  XNOR U32378 ( .A(n32199), .B(n32198), .Z(n32200) );
  NANDN U32379 ( .A(n31805), .B(n31804), .Z(n31809) );
  NAND U32380 ( .A(n31807), .B(n31806), .Z(n31808) );
  NAND U32381 ( .A(n31809), .B(n31808), .Z(n32195) );
  NANDN U32382 ( .A(n31811), .B(n31810), .Z(n31815) );
  OR U32383 ( .A(n31813), .B(n31812), .Z(n31814) );
  NAND U32384 ( .A(n31815), .B(n31814), .Z(n32192) );
  OR U32385 ( .A(n31817), .B(n31816), .Z(n31821) );
  NAND U32386 ( .A(n31819), .B(n31818), .Z(n31820) );
  NAND U32387 ( .A(n31821), .B(n31820), .Z(n32057) );
  NANDN U32388 ( .A(n31823), .B(n31822), .Z(n31827) );
  NAND U32389 ( .A(n31825), .B(n31824), .Z(n31826) );
  NAND U32390 ( .A(n31827), .B(n31826), .Z(n32003) );
  XOR U32391 ( .A(b[39]), .B(n36420), .Z(n32156) );
  NANDN U32392 ( .A(n32156), .B(n36553), .Z(n31830) );
  NAND U32393 ( .A(n31828), .B(n36643), .Z(n31829) );
  NAND U32394 ( .A(n31830), .B(n31829), .Z(n32131) );
  XNOR U32395 ( .A(a[106]), .B(b[35]), .Z(n32104) );
  NANDN U32396 ( .A(n32104), .B(n35985), .Z(n31833) );
  NAND U32397 ( .A(n31831), .B(n35986), .Z(n31832) );
  NAND U32398 ( .A(n31833), .B(n31832), .Z(n32128) );
  XOR U32399 ( .A(a[108]), .B(n974), .Z(n32035) );
  NANDN U32400 ( .A(n32035), .B(n35620), .Z(n31836) );
  NAND U32401 ( .A(n31834), .B(n35621), .Z(n31835) );
  AND U32402 ( .A(n31836), .B(n31835), .Z(n32129) );
  XNOR U32403 ( .A(n32128), .B(n32129), .Z(n32130) );
  XNOR U32404 ( .A(n32131), .B(n32130), .Z(n32001) );
  NANDN U32405 ( .A(n31838), .B(n31837), .Z(n31842) );
  NANDN U32406 ( .A(n31840), .B(n31839), .Z(n31841) );
  NAND U32407 ( .A(n31842), .B(n31841), .Z(n32002) );
  XOR U32408 ( .A(n32001), .B(n32002), .Z(n32004) );
  XNOR U32409 ( .A(n32003), .B(n32004), .Z(n31995) );
  NANDN U32410 ( .A(n31844), .B(n31843), .Z(n31848) );
  NAND U32411 ( .A(n31846), .B(n31845), .Z(n31847) );
  AND U32412 ( .A(n31848), .B(n31847), .Z(n31996) );
  XNOR U32413 ( .A(n31995), .B(n31996), .Z(n31997) );
  OR U32414 ( .A(n31850), .B(n31849), .Z(n31854) );
  NAND U32415 ( .A(n31852), .B(n31851), .Z(n31853) );
  NAND U32416 ( .A(n31854), .B(n31853), .Z(n31998) );
  XOR U32417 ( .A(n31997), .B(n31998), .Z(n31989) );
  NANDN U32418 ( .A(n31856), .B(n31855), .Z(n31860) );
  OR U32419 ( .A(n31858), .B(n31857), .Z(n31859) );
  AND U32420 ( .A(n31860), .B(n31859), .Z(n31990) );
  XNOR U32421 ( .A(n31989), .B(n31990), .Z(n31991) );
  XOR U32422 ( .A(a[110]), .B(n973), .Z(n32032) );
  NANDN U32423 ( .A(n32032), .B(n35313), .Z(n31863) );
  NANDN U32424 ( .A(n31861), .B(n35311), .Z(n31862) );
  NAND U32425 ( .A(n31863), .B(n31862), .Z(n32125) );
  XOR U32426 ( .A(b[43]), .B(n35783), .Z(n32007) );
  NANDN U32427 ( .A(n32007), .B(n37068), .Z(n31866) );
  NANDN U32428 ( .A(n31864), .B(n37069), .Z(n31865) );
  NAND U32429 ( .A(n31866), .B(n31865), .Z(n32122) );
  XOR U32430 ( .A(b[49]), .B(n34852), .Z(n32086) );
  OR U32431 ( .A(n32086), .B(n37756), .Z(n31869) );
  NANDN U32432 ( .A(n31867), .B(n37652), .Z(n31868) );
  AND U32433 ( .A(n31869), .B(n31868), .Z(n32123) );
  XNOR U32434 ( .A(n32122), .B(n32123), .Z(n32124) );
  XNOR U32435 ( .A(n32125), .B(n32124), .Z(n32068) );
  XOR U32436 ( .A(b[63]), .B(n31870), .Z(n32015) );
  NANDN U32437 ( .A(n32015), .B(n38422), .Z(n31873) );
  NAND U32438 ( .A(n31871), .B(n38423), .Z(n31872) );
  NAND U32439 ( .A(n31873), .B(n31872), .Z(n32019) );
  NANDN U32440 ( .A(n31875), .B(n31874), .Z(n31876) );
  NANDN U32441 ( .A(n31877), .B(n31876), .Z(n32018) );
  AND U32442 ( .A(b[63]), .B(a[76]), .Z(n32282) );
  XOR U32443 ( .A(n32018), .B(n32282), .Z(n32020) );
  XNOR U32444 ( .A(n32019), .B(n32020), .Z(n32069) );
  XOR U32445 ( .A(n32068), .B(n32069), .Z(n32071) );
  NANDN U32446 ( .A(n31879), .B(n31878), .Z(n31883) );
  NAND U32447 ( .A(n31881), .B(n31880), .Z(n31882) );
  NAND U32448 ( .A(n31883), .B(n31882), .Z(n32070) );
  XNOR U32449 ( .A(n32071), .B(n32070), .Z(n32177) );
  NANDN U32450 ( .A(n31885), .B(n31884), .Z(n31889) );
  NAND U32451 ( .A(n31887), .B(n31886), .Z(n31888) );
  NAND U32452 ( .A(n31889), .B(n31888), .Z(n32174) );
  NAND U32453 ( .A(n31891), .B(n31890), .Z(n31895) );
  NANDN U32454 ( .A(n31893), .B(n31892), .Z(n31894) );
  NAND U32455 ( .A(n31895), .B(n31894), .Z(n32175) );
  XNOR U32456 ( .A(n32174), .B(n32175), .Z(n32176) );
  XNOR U32457 ( .A(n32177), .B(n32176), .Z(n32046) );
  XOR U32458 ( .A(b[57]), .B(n33185), .Z(n32110) );
  OR U32459 ( .A(n32110), .B(n965), .Z(n31898) );
  NANDN U32460 ( .A(n31896), .B(n38194), .Z(n31897) );
  NAND U32461 ( .A(n31898), .B(n31897), .Z(n32171) );
  NAND U32462 ( .A(n34848), .B(n31899), .Z(n31901) );
  XOR U32463 ( .A(n37873), .B(n35375), .Z(n32023) );
  NAND U32464 ( .A(n34618), .B(n32023), .Z(n31900) );
  NAND U32465 ( .A(n31901), .B(n31900), .Z(n32168) );
  XOR U32466 ( .A(a[104]), .B(n975), .Z(n32029) );
  NANDN U32467 ( .A(n32029), .B(n36311), .Z(n31904) );
  NANDN U32468 ( .A(n31902), .B(n36309), .Z(n31903) );
  AND U32469 ( .A(n31904), .B(n31903), .Z(n32169) );
  XNOR U32470 ( .A(n32168), .B(n32169), .Z(n32170) );
  XNOR U32471 ( .A(n32171), .B(n32170), .Z(n32186) );
  NAND U32472 ( .A(n37469), .B(n31905), .Z(n31907) );
  XOR U32473 ( .A(n978), .B(n35191), .Z(n32162) );
  NAND U32474 ( .A(n32162), .B(n37471), .Z(n31906) );
  NAND U32475 ( .A(n31907), .B(n31906), .Z(n32149) );
  NAND U32476 ( .A(n34044), .B(n31908), .Z(n31910) );
  XOR U32477 ( .A(n38143), .B(n34510), .Z(n32089) );
  NANDN U32478 ( .A(n33867), .B(n32089), .Z(n31909) );
  NAND U32479 ( .A(n31910), .B(n31909), .Z(n32146) );
  XNOR U32480 ( .A(a[120]), .B(b[21]), .Z(n32083) );
  OR U32481 ( .A(n32083), .B(n33634), .Z(n31913) );
  NANDN U32482 ( .A(n31911), .B(n33464), .Z(n31912) );
  AND U32483 ( .A(n31913), .B(n31912), .Z(n32147) );
  XNOR U32484 ( .A(n32146), .B(n32147), .Z(n32148) );
  XOR U32485 ( .A(n32149), .B(n32148), .Z(n32187) );
  XNOR U32486 ( .A(n32186), .B(n32187), .Z(n32188) );
  NANDN U32487 ( .A(n31915), .B(n31914), .Z(n31919) );
  NAND U32488 ( .A(n31917), .B(n31916), .Z(n31918) );
  AND U32489 ( .A(n31919), .B(n31918), .Z(n32189) );
  XNOR U32490 ( .A(n32188), .B(n32189), .Z(n32045) );
  NANDN U32491 ( .A(n31921), .B(n31920), .Z(n31925) );
  NAND U32492 ( .A(n31923), .B(n31922), .Z(n31924) );
  NAND U32493 ( .A(n31925), .B(n31924), .Z(n32182) );
  XNOR U32494 ( .A(b[45]), .B(a[96]), .Z(n32119) );
  NANDN U32495 ( .A(n32119), .B(n37261), .Z(n31928) );
  NANDN U32496 ( .A(n31926), .B(n37262), .Z(n31927) );
  NAND U32497 ( .A(n31928), .B(n31927), .Z(n32143) );
  NAND U32498 ( .A(n33283), .B(n31929), .Z(n31931) );
  XOR U32499 ( .A(n38251), .B(n33020), .Z(n32113) );
  NANDN U32500 ( .A(n33021), .B(n32113), .Z(n31930) );
  NAND U32501 ( .A(n31931), .B(n31930), .Z(n32140) );
  XOR U32502 ( .A(b[61]), .B(n32814), .Z(n32080) );
  OR U32503 ( .A(n32080), .B(n38371), .Z(n31934) );
  NANDN U32504 ( .A(n31932), .B(n38369), .Z(n31933) );
  AND U32505 ( .A(n31934), .B(n31933), .Z(n32141) );
  XNOR U32506 ( .A(n32140), .B(n32141), .Z(n32142) );
  XNOR U32507 ( .A(n32143), .B(n32142), .Z(n32180) );
  XNOR U32508 ( .A(b[41]), .B(a[100]), .Z(n32153) );
  OR U32509 ( .A(n32153), .B(n36905), .Z(n31937) );
  NAND U32510 ( .A(n31935), .B(n36807), .Z(n31936) );
  NAND U32511 ( .A(n31937), .B(n31936), .Z(n32137) );
  XNOR U32512 ( .A(a[124]), .B(b[17]), .Z(n32116) );
  NANDN U32513 ( .A(n32116), .B(n32543), .Z(n31940) );
  NAND U32514 ( .A(n31938), .B(n32541), .Z(n31939) );
  NAND U32515 ( .A(n31940), .B(n31939), .Z(n32134) );
  XOR U32516 ( .A(a[126]), .B(n972), .Z(n32012) );
  OR U32517 ( .A(n32012), .B(n32010), .Z(n31943) );
  NANDN U32518 ( .A(n31941), .B(n32011), .Z(n31942) );
  AND U32519 ( .A(n31943), .B(n31942), .Z(n32135) );
  XNOR U32520 ( .A(n32134), .B(n32135), .Z(n32136) );
  XOR U32521 ( .A(n32137), .B(n32136), .Z(n32181) );
  XOR U32522 ( .A(n32180), .B(n32181), .Z(n32183) );
  XOR U32523 ( .A(n32182), .B(n32183), .Z(n32044) );
  XOR U32524 ( .A(n32045), .B(n32044), .Z(n32047) );
  XNOR U32525 ( .A(n32046), .B(n32047), .Z(n31992) );
  XOR U32526 ( .A(n31991), .B(n31992), .Z(n32056) );
  XNOR U32527 ( .A(n32057), .B(n32056), .Z(n32058) );
  NANDN U32528 ( .A(n31945), .B(n31944), .Z(n31949) );
  OR U32529 ( .A(n31947), .B(n31946), .Z(n31948) );
  NAND U32530 ( .A(n31949), .B(n31948), .Z(n31986) );
  NANDN U32531 ( .A(n31951), .B(n31950), .Z(n31955) );
  OR U32532 ( .A(n31953), .B(n31952), .Z(n31954) );
  NAND U32533 ( .A(n31955), .B(n31954), .Z(n31983) );
  NAND U32534 ( .A(n31957), .B(n31956), .Z(n31961) );
  NANDN U32535 ( .A(n31959), .B(n31958), .Z(n31960) );
  AND U32536 ( .A(n31961), .B(n31960), .Z(n31984) );
  XNOR U32537 ( .A(n31983), .B(n31984), .Z(n31985) );
  XNOR U32538 ( .A(n31986), .B(n31985), .Z(n32059) );
  XOR U32539 ( .A(n32058), .B(n32059), .Z(n32193) );
  XNOR U32540 ( .A(n32192), .B(n32193), .Z(n32194) );
  XOR U32541 ( .A(n32195), .B(n32194), .Z(n32201) );
  XOR U32542 ( .A(n32200), .B(n32201), .Z(n32202) );
  XNOR U32543 ( .A(n32203), .B(n32202), .Z(n32204) );
  XNOR U32544 ( .A(n32205), .B(n32204), .Z(n31977) );
  XNOR U32545 ( .A(n31977), .B(n31978), .Z(n31979) );
  XOR U32546 ( .A(n31979), .B(n31980), .Z(n31971) );
  XNOR U32547 ( .A(n31974), .B(n31971), .Z(n31970) );
  XNOR U32548 ( .A(n31973), .B(n31970), .Z(n32208) );
  XOR U32549 ( .A(n32209), .B(n32208), .Z(c[204]) );
  XOR U32550 ( .A(n31974), .B(n31973), .Z(n31972) );
  NAND U32551 ( .A(n31972), .B(n31971), .Z(n31976) );
  OR U32552 ( .A(n31974), .B(n31973), .Z(n31975) );
  AND U32553 ( .A(n31976), .B(n31975), .Z(n32214) );
  NANDN U32554 ( .A(n31978), .B(n31977), .Z(n31982) );
  NANDN U32555 ( .A(n31980), .B(n31979), .Z(n31981) );
  NAND U32556 ( .A(n31982), .B(n31981), .Z(n32213) );
  NANDN U32557 ( .A(n31984), .B(n31983), .Z(n31988) );
  NAND U32558 ( .A(n31986), .B(n31985), .Z(n31987) );
  NAND U32559 ( .A(n31988), .B(n31987), .Z(n32239) );
  NANDN U32560 ( .A(n31990), .B(n31989), .Z(n31994) );
  NAND U32561 ( .A(n31992), .B(n31991), .Z(n31993) );
  NAND U32562 ( .A(n31994), .B(n31993), .Z(n32237) );
  NANDN U32563 ( .A(n31996), .B(n31995), .Z(n32000) );
  NANDN U32564 ( .A(n31998), .B(n31997), .Z(n31999) );
  NAND U32565 ( .A(n32000), .B(n31999), .Z(n32251) );
  NANDN U32566 ( .A(n32002), .B(n32001), .Z(n32006) );
  OR U32567 ( .A(n32004), .B(n32003), .Z(n32005) );
  NAND U32568 ( .A(n32006), .B(n32005), .Z(n32249) );
  XNOR U32569 ( .A(b[43]), .B(a[99]), .Z(n32377) );
  NANDN U32570 ( .A(n32377), .B(n37068), .Z(n32009) );
  NANDN U32571 ( .A(n32007), .B(n37069), .Z(n32008) );
  NAND U32572 ( .A(n32009), .B(n32008), .Z(n32328) );
  XNOR U32573 ( .A(n38463), .B(b[15]), .Z(n32347) );
  NANDN U32574 ( .A(n32010), .B(n32347), .Z(n32014) );
  NANDN U32575 ( .A(n32012), .B(n32011), .Z(n32013) );
  NAND U32576 ( .A(n32014), .B(n32013), .Z(n32325) );
  XNOR U32577 ( .A(b[63]), .B(a[79]), .Z(n32350) );
  NANDN U32578 ( .A(n32350), .B(n38422), .Z(n32017) );
  NANDN U32579 ( .A(n32015), .B(n38423), .Z(n32016) );
  AND U32580 ( .A(n32017), .B(n32016), .Z(n32326) );
  XNOR U32581 ( .A(n32325), .B(n32326), .Z(n32327) );
  XNOR U32582 ( .A(n32328), .B(n32327), .Z(n32285) );
  NANDN U32583 ( .A(n32282), .B(n32018), .Z(n32022) );
  NANDN U32584 ( .A(n32020), .B(n32019), .Z(n32021) );
  NAND U32585 ( .A(n32022), .B(n32021), .Z(n32286) );
  XNOR U32586 ( .A(n32285), .B(n32286), .Z(n32287) );
  NAND U32587 ( .A(n34848), .B(n32023), .Z(n32025) );
  XNOR U32588 ( .A(a[115]), .B(b[27]), .Z(n32386) );
  NANDN U32589 ( .A(n32386), .B(n34618), .Z(n32024) );
  NAND U32590 ( .A(n32025), .B(n32024), .Z(n32334) );
  NAND U32591 ( .A(n35188), .B(n32026), .Z(n32028) );
  XNOR U32592 ( .A(a[113]), .B(n35540), .Z(n32270) );
  NANDN U32593 ( .A(n34968), .B(n32270), .Z(n32027) );
  NAND U32594 ( .A(n32028), .B(n32027), .Z(n32331) );
  XNOR U32595 ( .A(a[105]), .B(n975), .Z(n32380) );
  NAND U32596 ( .A(n32380), .B(n36311), .Z(n32031) );
  NANDN U32597 ( .A(n32029), .B(n36309), .Z(n32030) );
  AND U32598 ( .A(n32031), .B(n32030), .Z(n32332) );
  XNOR U32599 ( .A(n32331), .B(n32332), .Z(n32333) );
  XNOR U32600 ( .A(n32334), .B(n32333), .Z(n32292) );
  NANDN U32601 ( .A(n32032), .B(n35311), .Z(n32034) );
  XNOR U32602 ( .A(a[111]), .B(n973), .Z(n32371) );
  NAND U32603 ( .A(n32371), .B(n35313), .Z(n32033) );
  NAND U32604 ( .A(n32034), .B(n32033), .Z(n32290) );
  XNOR U32605 ( .A(a[109]), .B(n974), .Z(n32374) );
  NAND U32606 ( .A(n35620), .B(n32374), .Z(n32037) );
  NANDN U32607 ( .A(n32035), .B(n35621), .Z(n32036) );
  AND U32608 ( .A(n32037), .B(n32036), .Z(n32289) );
  XNOR U32609 ( .A(n32290), .B(n32289), .Z(n32291) );
  XOR U32610 ( .A(n32292), .B(n32291), .Z(n32288) );
  XOR U32611 ( .A(n32287), .B(n32288), .Z(n32248) );
  XOR U32612 ( .A(n32249), .B(n32248), .Z(n32250) );
  XOR U32613 ( .A(n32251), .B(n32250), .Z(n32245) );
  NANDN U32614 ( .A(n32039), .B(n32038), .Z(n32043) );
  NAND U32615 ( .A(n32041), .B(n32040), .Z(n32042) );
  AND U32616 ( .A(n32043), .B(n32042), .Z(n32242) );
  NANDN U32617 ( .A(n32045), .B(n32044), .Z(n32049) );
  NANDN U32618 ( .A(n32047), .B(n32046), .Z(n32048) );
  AND U32619 ( .A(n32049), .B(n32048), .Z(n32243) );
  XNOR U32620 ( .A(n32245), .B(n32244), .Z(n32236) );
  XOR U32621 ( .A(n32237), .B(n32236), .Z(n32238) );
  XNOR U32622 ( .A(n32239), .B(n32238), .Z(n32227) );
  NANDN U32623 ( .A(n32051), .B(n32050), .Z(n32055) );
  NAND U32624 ( .A(n32053), .B(n32052), .Z(n32054) );
  AND U32625 ( .A(n32055), .B(n32054), .Z(n32220) );
  NANDN U32626 ( .A(n32057), .B(n32056), .Z(n32061) );
  NANDN U32627 ( .A(n32059), .B(n32058), .Z(n32060) );
  AND U32628 ( .A(n32061), .B(n32060), .Z(n32218) );
  NANDN U32629 ( .A(n32063), .B(n32062), .Z(n32067) );
  OR U32630 ( .A(n32065), .B(n32064), .Z(n32066) );
  NAND U32631 ( .A(n32067), .B(n32066), .Z(n32231) );
  NANDN U32632 ( .A(n32069), .B(n32068), .Z(n32073) );
  OR U32633 ( .A(n32071), .B(n32070), .Z(n32072) );
  NAND U32634 ( .A(n32073), .B(n32072), .Z(n32428) );
  NANDN U32635 ( .A(n32075), .B(n32074), .Z(n32079) );
  NAND U32636 ( .A(n32077), .B(n32076), .Z(n32078) );
  NAND U32637 ( .A(n32079), .B(n32078), .Z(n32406) );
  XNOR U32638 ( .A(b[61]), .B(a[81]), .Z(n32319) );
  OR U32639 ( .A(n32319), .B(n38371), .Z(n32082) );
  NANDN U32640 ( .A(n32080), .B(n38369), .Z(n32081) );
  NAND U32641 ( .A(n32082), .B(n32081), .Z(n32356) );
  XOR U32642 ( .A(a[121]), .B(b[21]), .Z(n32398) );
  NANDN U32643 ( .A(n33634), .B(n32398), .Z(n32085) );
  NANDN U32644 ( .A(n32083), .B(n33464), .Z(n32084) );
  NAND U32645 ( .A(n32085), .B(n32084), .Z(n32353) );
  XOR U32646 ( .A(b[49]), .B(n35377), .Z(n32322) );
  OR U32647 ( .A(n32322), .B(n37756), .Z(n32088) );
  NANDN U32648 ( .A(n32086), .B(n37652), .Z(n32087) );
  AND U32649 ( .A(n32088), .B(n32087), .Z(n32354) );
  XNOR U32650 ( .A(n32353), .B(n32354), .Z(n32355) );
  XNOR U32651 ( .A(n32356), .B(n32355), .Z(n32404) );
  NAND U32652 ( .A(n34044), .B(n32089), .Z(n32091) );
  XOR U32653 ( .A(n38193), .B(n34510), .Z(n32395) );
  NANDN U32654 ( .A(n33867), .B(n32395), .Z(n32090) );
  NAND U32655 ( .A(n32091), .B(n32090), .Z(n32368) );
  NAND U32656 ( .A(n38326), .B(n32092), .Z(n32094) );
  XNOR U32657 ( .A(n38400), .B(a[83]), .Z(n32389) );
  NANDN U32658 ( .A(n38273), .B(n32389), .Z(n32093) );
  NAND U32659 ( .A(n32094), .B(n32093), .Z(n32365) );
  XNOR U32660 ( .A(b[51]), .B(a[91]), .Z(n32392) );
  NANDN U32661 ( .A(n32392), .B(n37803), .Z(n32097) );
  NANDN U32662 ( .A(n32095), .B(n37802), .Z(n32096) );
  AND U32663 ( .A(n32097), .B(n32096), .Z(n32366) );
  XNOR U32664 ( .A(n32365), .B(n32366), .Z(n32367) );
  XOR U32665 ( .A(n32368), .B(n32367), .Z(n32405) );
  XOR U32666 ( .A(n32404), .B(n32405), .Z(n32407) );
  XOR U32667 ( .A(n32406), .B(n32407), .Z(n32419) );
  NANDN U32668 ( .A(n32099), .B(n32098), .Z(n32103) );
  NAND U32669 ( .A(n32101), .B(n32100), .Z(n32102) );
  NAND U32670 ( .A(n32103), .B(n32102), .Z(n32417) );
  XOR U32671 ( .A(a[107]), .B(b[35]), .Z(n32383) );
  NAND U32672 ( .A(n35985), .B(n32383), .Z(n32106) );
  NANDN U32673 ( .A(n32104), .B(n35986), .Z(n32105) );
  NAND U32674 ( .A(n32106), .B(n32105), .Z(n32304) );
  XNOR U32675 ( .A(b[55]), .B(a[87]), .Z(n32310) );
  NANDN U32676 ( .A(n32310), .B(n38075), .Z(n32109) );
  NANDN U32677 ( .A(n32107), .B(n38073), .Z(n32108) );
  NAND U32678 ( .A(n32109), .B(n32108), .Z(n32301) );
  XNOR U32679 ( .A(b[57]), .B(a[85]), .Z(n32313) );
  OR U32680 ( .A(n32313), .B(n965), .Z(n32112) );
  NANDN U32681 ( .A(n32110), .B(n38194), .Z(n32111) );
  AND U32682 ( .A(n32112), .B(n32111), .Z(n32302) );
  XNOR U32683 ( .A(n32301), .B(n32302), .Z(n32303) );
  XNOR U32684 ( .A(n32304), .B(n32303), .Z(n32257) );
  NAND U32685 ( .A(n33283), .B(n32113), .Z(n32115) );
  XNOR U32686 ( .A(a[123]), .B(n33020), .Z(n32340) );
  NANDN U32687 ( .A(n33021), .B(n32340), .Z(n32114) );
  NAND U32688 ( .A(n32115), .B(n32114), .Z(n32298) );
  XOR U32689 ( .A(a[125]), .B(b[17]), .Z(n32343) );
  NAND U32690 ( .A(n32343), .B(n32543), .Z(n32118) );
  NANDN U32691 ( .A(n32116), .B(n32541), .Z(n32117) );
  NAND U32692 ( .A(n32118), .B(n32117), .Z(n32295) );
  XOR U32693 ( .A(b[45]), .B(a[97]), .Z(n32401) );
  NAND U32694 ( .A(n32401), .B(n37261), .Z(n32121) );
  NANDN U32695 ( .A(n32119), .B(n37262), .Z(n32120) );
  AND U32696 ( .A(n32121), .B(n32120), .Z(n32296) );
  XNOR U32697 ( .A(n32295), .B(n32296), .Z(n32297) );
  XNOR U32698 ( .A(n32298), .B(n32297), .Z(n32254) );
  NANDN U32699 ( .A(n32123), .B(n32122), .Z(n32127) );
  NAND U32700 ( .A(n32125), .B(n32124), .Z(n32126) );
  NAND U32701 ( .A(n32127), .B(n32126), .Z(n32255) );
  XNOR U32702 ( .A(n32254), .B(n32255), .Z(n32256) );
  XOR U32703 ( .A(n32257), .B(n32256), .Z(n32422) );
  NANDN U32704 ( .A(n32129), .B(n32128), .Z(n32133) );
  NAND U32705 ( .A(n32131), .B(n32130), .Z(n32132) );
  NAND U32706 ( .A(n32133), .B(n32132), .Z(n32423) );
  XOR U32707 ( .A(n32422), .B(n32423), .Z(n32425) );
  NANDN U32708 ( .A(n32135), .B(n32134), .Z(n32139) );
  NAND U32709 ( .A(n32137), .B(n32136), .Z(n32138) );
  NAND U32710 ( .A(n32139), .B(n32138), .Z(n32424) );
  XNOR U32711 ( .A(n32425), .B(n32424), .Z(n32416) );
  XOR U32712 ( .A(n32417), .B(n32416), .Z(n32418) );
  XNOR U32713 ( .A(n32419), .B(n32418), .Z(n32429) );
  XNOR U32714 ( .A(n32428), .B(n32429), .Z(n32430) );
  NANDN U32715 ( .A(n32141), .B(n32140), .Z(n32145) );
  NAND U32716 ( .A(n32143), .B(n32142), .Z(n32144) );
  NAND U32717 ( .A(n32145), .B(n32144), .Z(n32413) );
  NANDN U32718 ( .A(n32147), .B(n32146), .Z(n32151) );
  NAND U32719 ( .A(n32149), .B(n32148), .Z(n32150) );
  NAND U32720 ( .A(n32151), .B(n32150), .Z(n32261) );
  NANDN U32721 ( .A(n970), .B(b[12]), .Z(n32152) );
  AND U32722 ( .A(n32152), .B(b[13]), .Z(n32359) );
  XOR U32723 ( .A(b[41]), .B(a[101]), .Z(n32337) );
  NANDN U32724 ( .A(n36905), .B(n32337), .Z(n32155) );
  NANDN U32725 ( .A(n32153), .B(n36807), .Z(n32154) );
  AND U32726 ( .A(n32155), .B(n32154), .Z(n32360) );
  XOR U32727 ( .A(n32359), .B(n32360), .Z(n32361) );
  XNOR U32728 ( .A(b[39]), .B(a[103]), .Z(n32307) );
  NANDN U32729 ( .A(n32307), .B(n36553), .Z(n32158) );
  NANDN U32730 ( .A(n32156), .B(n36643), .Z(n32157) );
  NAND U32731 ( .A(n32158), .B(n32157), .Z(n32279) );
  NANDN U32732 ( .A(n985), .B(a[77]), .Z(n32280) );
  XNOR U32733 ( .A(n32279), .B(n32280), .Z(n32281) );
  XNOR U32734 ( .A(n32282), .B(n32281), .Z(n32362) );
  XNOR U32735 ( .A(n32361), .B(n32362), .Z(n32259) );
  XOR U32736 ( .A(a[117]), .B(b[25]), .Z(n32316) );
  NANDN U32737 ( .A(n34219), .B(n32316), .Z(n32161) );
  NAND U32738 ( .A(n34217), .B(n32159), .Z(n32160) );
  NAND U32739 ( .A(n32161), .B(n32160), .Z(n32267) );
  NAND U32740 ( .A(n37469), .B(n32162), .Z(n32164) );
  XOR U32741 ( .A(n978), .B(n35628), .Z(n32273) );
  NAND U32742 ( .A(n32273), .B(n37471), .Z(n32163) );
  NAND U32743 ( .A(n32164), .B(n32163), .Z(n32264) );
  XNOR U32744 ( .A(b[53]), .B(a[89]), .Z(n32276) );
  NANDN U32745 ( .A(n32276), .B(n37940), .Z(n32167) );
  NANDN U32746 ( .A(n32165), .B(n37941), .Z(n32166) );
  AND U32747 ( .A(n32167), .B(n32166), .Z(n32265) );
  XNOR U32748 ( .A(n32264), .B(n32265), .Z(n32266) );
  XNOR U32749 ( .A(n32267), .B(n32266), .Z(n32258) );
  XOR U32750 ( .A(n32259), .B(n32258), .Z(n32260) );
  XNOR U32751 ( .A(n32261), .B(n32260), .Z(n32411) );
  NANDN U32752 ( .A(n32169), .B(n32168), .Z(n32173) );
  NAND U32753 ( .A(n32171), .B(n32170), .Z(n32172) );
  AND U32754 ( .A(n32173), .B(n32172), .Z(n32410) );
  XNOR U32755 ( .A(n32411), .B(n32410), .Z(n32412) );
  XOR U32756 ( .A(n32413), .B(n32412), .Z(n32431) );
  XNOR U32757 ( .A(n32430), .B(n32431), .Z(n32230) );
  XNOR U32758 ( .A(n32231), .B(n32230), .Z(n32232) );
  NANDN U32759 ( .A(n32175), .B(n32174), .Z(n32179) );
  NAND U32760 ( .A(n32177), .B(n32176), .Z(n32178) );
  NAND U32761 ( .A(n32179), .B(n32178), .Z(n32437) );
  NANDN U32762 ( .A(n32181), .B(n32180), .Z(n32185) );
  OR U32763 ( .A(n32183), .B(n32182), .Z(n32184) );
  NAND U32764 ( .A(n32185), .B(n32184), .Z(n32434) );
  NANDN U32765 ( .A(n32187), .B(n32186), .Z(n32191) );
  NAND U32766 ( .A(n32189), .B(n32188), .Z(n32190) );
  AND U32767 ( .A(n32191), .B(n32190), .Z(n32435) );
  XNOR U32768 ( .A(n32434), .B(n32435), .Z(n32436) );
  XOR U32769 ( .A(n32437), .B(n32436), .Z(n32233) );
  XNOR U32770 ( .A(n32232), .B(n32233), .Z(n32219) );
  XNOR U32771 ( .A(n32218), .B(n32219), .Z(n32221) );
  XNOR U32772 ( .A(n32220), .B(n32221), .Z(n32224) );
  NANDN U32773 ( .A(n32193), .B(n32192), .Z(n32197) );
  NAND U32774 ( .A(n32195), .B(n32194), .Z(n32196) );
  NAND U32775 ( .A(n32197), .B(n32196), .Z(n32225) );
  XNOR U32776 ( .A(n32224), .B(n32225), .Z(n32226) );
  XOR U32777 ( .A(n32227), .B(n32226), .Z(n32440) );
  XNOR U32778 ( .A(n32440), .B(n32441), .Z(n32443) );
  NAND U32779 ( .A(n32203), .B(n32202), .Z(n32207) );
  OR U32780 ( .A(n32205), .B(n32204), .Z(n32206) );
  AND U32781 ( .A(n32207), .B(n32206), .Z(n32442) );
  XNOR U32782 ( .A(n32443), .B(n32442), .Z(n32212) );
  XNOR U32783 ( .A(n32213), .B(n32212), .Z(n32215) );
  XNOR U32784 ( .A(n32214), .B(n32215), .Z(n32210) );
  OR U32785 ( .A(n32209), .B(n32208), .Z(n32211) );
  XNOR U32786 ( .A(n32210), .B(n32211), .Z(c[205]) );
  NANDN U32787 ( .A(n32211), .B(n32210), .Z(n32671) );
  NAND U32788 ( .A(n32213), .B(n32212), .Z(n32217) );
  NANDN U32789 ( .A(n32215), .B(n32214), .Z(n32216) );
  AND U32790 ( .A(n32217), .B(n32216), .Z(n32449) );
  OR U32791 ( .A(n32219), .B(n32218), .Z(n32223) );
  OR U32792 ( .A(n32221), .B(n32220), .Z(n32222) );
  NAND U32793 ( .A(n32223), .B(n32222), .Z(n32669) );
  NANDN U32794 ( .A(n32225), .B(n32224), .Z(n32229) );
  NAND U32795 ( .A(n32227), .B(n32226), .Z(n32228) );
  NAND U32796 ( .A(n32229), .B(n32228), .Z(n32667) );
  NAND U32797 ( .A(n32231), .B(n32230), .Z(n32235) );
  OR U32798 ( .A(n32233), .B(n32232), .Z(n32234) );
  NAND U32799 ( .A(n32235), .B(n32234), .Z(n32459) );
  NAND U32800 ( .A(n32237), .B(n32236), .Z(n32241) );
  NAND U32801 ( .A(n32239), .B(n32238), .Z(n32240) );
  NAND U32802 ( .A(n32241), .B(n32240), .Z(n32456) );
  OR U32803 ( .A(n32243), .B(n32242), .Z(n32247) );
  NANDN U32804 ( .A(n32245), .B(n32244), .Z(n32246) );
  NAND U32805 ( .A(n32247), .B(n32246), .Z(n32453) );
  NAND U32806 ( .A(n32249), .B(n32248), .Z(n32253) );
  NANDN U32807 ( .A(n32251), .B(n32250), .Z(n32252) );
  NAND U32808 ( .A(n32253), .B(n32252), .Z(n32493) );
  NANDN U32809 ( .A(n32259), .B(n32258), .Z(n32263) );
  OR U32810 ( .A(n32261), .B(n32260), .Z(n32262) );
  AND U32811 ( .A(n32263), .B(n32262), .Z(n32577) );
  XNOR U32812 ( .A(n32576), .B(n32577), .Z(n32578) );
  NANDN U32813 ( .A(n32265), .B(n32264), .Z(n32269) );
  NAND U32814 ( .A(n32267), .B(n32266), .Z(n32268) );
  NAND U32815 ( .A(n32269), .B(n32268), .Z(n32572) );
  NAND U32816 ( .A(n35188), .B(n32270), .Z(n32272) );
  XNOR U32817 ( .A(n37873), .B(b[29]), .Z(n32532) );
  NANDN U32818 ( .A(n34968), .B(n32532), .Z(n32271) );
  NAND U32819 ( .A(n32272), .B(n32271), .Z(n32657) );
  NAND U32820 ( .A(n37469), .B(n32273), .Z(n32275) );
  XOR U32821 ( .A(n978), .B(n35545), .Z(n32621) );
  NAND U32822 ( .A(n32621), .B(n37471), .Z(n32274) );
  NAND U32823 ( .A(n32275), .B(n32274), .Z(n32654) );
  XOR U32824 ( .A(b[53]), .B(n34851), .Z(n32645) );
  NANDN U32825 ( .A(n32645), .B(n37940), .Z(n32278) );
  NANDN U32826 ( .A(n32276), .B(n37941), .Z(n32277) );
  AND U32827 ( .A(n32278), .B(n32277), .Z(n32655) );
  XNOR U32828 ( .A(n32654), .B(n32655), .Z(n32656) );
  XNOR U32829 ( .A(n32657), .B(n32656), .Z(n32570) );
  NANDN U32830 ( .A(n32280), .B(n32279), .Z(n32284) );
  NAND U32831 ( .A(n32282), .B(n32281), .Z(n32283) );
  NAND U32832 ( .A(n32284), .B(n32283), .Z(n32571) );
  XOR U32833 ( .A(n32570), .B(n32571), .Z(n32573) );
  XOR U32834 ( .A(n32572), .B(n32573), .Z(n32579) );
  XOR U32835 ( .A(n32578), .B(n32579), .Z(n32492) );
  XNOR U32836 ( .A(n32493), .B(n32492), .Z(n32495) );
  NANDN U32837 ( .A(n32290), .B(n32289), .Z(n32294) );
  NAND U32838 ( .A(n32292), .B(n32291), .Z(n32293) );
  NAND U32839 ( .A(n32294), .B(n32293), .Z(n32462) );
  NANDN U32840 ( .A(n32296), .B(n32295), .Z(n32300) );
  NAND U32841 ( .A(n32298), .B(n32297), .Z(n32299) );
  NAND U32842 ( .A(n32300), .B(n32299), .Z(n32463) );
  XNOR U32843 ( .A(n32462), .B(n32463), .Z(n32464) );
  NANDN U32844 ( .A(n32302), .B(n32301), .Z(n32306) );
  NAND U32845 ( .A(n32304), .B(n32303), .Z(n32305) );
  NAND U32846 ( .A(n32306), .B(n32305), .Z(n32488) );
  XOR U32847 ( .A(n36647), .B(n976), .Z(n32520) );
  NAND U32848 ( .A(n32520), .B(n36553), .Z(n32309) );
  NANDN U32849 ( .A(n32307), .B(n36643), .Z(n32308) );
  NAND U32850 ( .A(n32309), .B(n32308), .Z(n32603) );
  XOR U32851 ( .A(b[55]), .B(n34048), .Z(n32651) );
  NANDN U32852 ( .A(n32651), .B(n38075), .Z(n32312) );
  NANDN U32853 ( .A(n32310), .B(n38073), .Z(n32311) );
  NAND U32854 ( .A(n32312), .B(n32311), .Z(n32600) );
  XOR U32855 ( .A(b[57]), .B(n33628), .Z(n32615) );
  OR U32856 ( .A(n32615), .B(n965), .Z(n32315) );
  NANDN U32857 ( .A(n32313), .B(n38194), .Z(n32314) );
  AND U32858 ( .A(n32315), .B(n32314), .Z(n32601) );
  XNOR U32859 ( .A(n32600), .B(n32601), .Z(n32602) );
  XNOR U32860 ( .A(n32603), .B(n32602), .Z(n32486) );
  XNOR U32861 ( .A(n38143), .B(b[25]), .Z(n32550) );
  NANDN U32862 ( .A(n34219), .B(n32550), .Z(n32318) );
  NAND U32863 ( .A(n34217), .B(n32316), .Z(n32317) );
  NAND U32864 ( .A(n32318), .B(n32317), .Z(n32633) );
  XOR U32865 ( .A(b[61]), .B(n32815), .Z(n32609) );
  OR U32866 ( .A(n32609), .B(n38371), .Z(n32321) );
  NANDN U32867 ( .A(n32319), .B(n38369), .Z(n32320) );
  NAND U32868 ( .A(n32321), .B(n32320), .Z(n32630) );
  XOR U32869 ( .A(b[49]), .B(n35191), .Z(n32553) );
  OR U32870 ( .A(n32553), .B(n37756), .Z(n32324) );
  NANDN U32871 ( .A(n32322), .B(n37652), .Z(n32323) );
  AND U32872 ( .A(n32324), .B(n32323), .Z(n32631) );
  XNOR U32873 ( .A(n32630), .B(n32631), .Z(n32632) );
  XOR U32874 ( .A(n32633), .B(n32632), .Z(n32487) );
  XOR U32875 ( .A(n32486), .B(n32487), .Z(n32489) );
  XOR U32876 ( .A(n32488), .B(n32489), .Z(n32465) );
  XOR U32877 ( .A(n32464), .B(n32465), .Z(n32504) );
  XNOR U32878 ( .A(n32505), .B(n32504), .Z(n32506) );
  NANDN U32879 ( .A(n32326), .B(n32325), .Z(n32330) );
  NAND U32880 ( .A(n32328), .B(n32327), .Z(n32329) );
  NAND U32881 ( .A(n32330), .B(n32329), .Z(n32477) );
  NANDN U32882 ( .A(n32332), .B(n32331), .Z(n32336) );
  NAND U32883 ( .A(n32334), .B(n32333), .Z(n32335) );
  NAND U32884 ( .A(n32336), .B(n32335), .Z(n32584) );
  XNOR U32885 ( .A(b[41]), .B(a[102]), .Z(n32546) );
  OR U32886 ( .A(n32546), .B(n36905), .Z(n32339) );
  NAND U32887 ( .A(n32337), .B(n36807), .Z(n32338) );
  NAND U32888 ( .A(n32339), .B(n32338), .Z(n32627) );
  NAND U32889 ( .A(n33283), .B(n32340), .Z(n32342) );
  XOR U32890 ( .A(n38321), .B(n33020), .Z(n32639) );
  NANDN U32891 ( .A(n33021), .B(n32639), .Z(n32341) );
  NAND U32892 ( .A(n32342), .B(n32341), .Z(n32624) );
  XNOR U32893 ( .A(a[126]), .B(b[17]), .Z(n32542) );
  NANDN U32894 ( .A(n32542), .B(n32543), .Z(n32345) );
  NAND U32895 ( .A(n32343), .B(n32541), .Z(n32344) );
  AND U32896 ( .A(n32345), .B(n32344), .Z(n32625) );
  XNOR U32897 ( .A(n32624), .B(n32625), .Z(n32626) );
  XNOR U32898 ( .A(n32627), .B(n32626), .Z(n32582) );
  NANDN U32899 ( .A(n971), .B(b[14]), .Z(n32549) );
  XOR U32900 ( .A(n972), .B(n32549), .Z(n32349) );
  XOR U32901 ( .A(b[14]), .B(n971), .Z(n32346) );
  NANDN U32902 ( .A(n32347), .B(n32346), .Z(n32348) );
  AND U32903 ( .A(n32349), .B(n32348), .Z(n32566) );
  AND U32904 ( .A(b[63]), .B(a[78]), .Z(n32806) );
  XOR U32905 ( .A(b[63]), .B(n32814), .Z(n32642) );
  NANDN U32906 ( .A(n32642), .B(n38422), .Z(n32352) );
  NANDN U32907 ( .A(n32350), .B(n38423), .Z(n32351) );
  AND U32908 ( .A(n32352), .B(n32351), .Z(n32565) );
  XNOR U32909 ( .A(n32806), .B(n32565), .Z(n32567) );
  XNOR U32910 ( .A(n32566), .B(n32567), .Z(n32583) );
  XOR U32911 ( .A(n32582), .B(n32583), .Z(n32585) );
  XOR U32912 ( .A(n32584), .B(n32585), .Z(n32474) );
  NANDN U32913 ( .A(n32354), .B(n32353), .Z(n32358) );
  NAND U32914 ( .A(n32356), .B(n32355), .Z(n32357) );
  AND U32915 ( .A(n32358), .B(n32357), .Z(n32475) );
  XOR U32916 ( .A(n32474), .B(n32475), .Z(n32476) );
  XOR U32917 ( .A(n32477), .B(n32476), .Z(n32507) );
  XOR U32918 ( .A(n32506), .B(n32507), .Z(n32494) );
  XOR U32919 ( .A(n32495), .B(n32494), .Z(n32451) );
  OR U32920 ( .A(n32360), .B(n32359), .Z(n32364) );
  NANDN U32921 ( .A(n32362), .B(n32361), .Z(n32363) );
  NAND U32922 ( .A(n32364), .B(n32363), .Z(n32469) );
  NANDN U32923 ( .A(n32366), .B(n32365), .Z(n32370) );
  NAND U32924 ( .A(n32368), .B(n32367), .Z(n32369) );
  AND U32925 ( .A(n32370), .B(n32369), .Z(n32468) );
  XNOR U32926 ( .A(n32469), .B(n32468), .Z(n32470) );
  XOR U32927 ( .A(a[112]), .B(n973), .Z(n32526) );
  NANDN U32928 ( .A(n32526), .B(n35313), .Z(n32373) );
  NAND U32929 ( .A(n32371), .B(n35311), .Z(n32372) );
  NAND U32930 ( .A(n32373), .B(n32372), .Z(n32538) );
  XOR U32931 ( .A(a[110]), .B(n974), .Z(n32523) );
  NANDN U32932 ( .A(n32523), .B(n35620), .Z(n32376) );
  NAND U32933 ( .A(n32374), .B(n35621), .Z(n32375) );
  NAND U32934 ( .A(n32376), .B(n32375), .Z(n32535) );
  XOR U32935 ( .A(b[43]), .B(n36100), .Z(n32636) );
  NANDN U32936 ( .A(n32636), .B(n37068), .Z(n32379) );
  NANDN U32937 ( .A(n32377), .B(n37069), .Z(n32378) );
  AND U32938 ( .A(n32379), .B(n32378), .Z(n32536) );
  XNOR U32939 ( .A(n32535), .B(n32536), .Z(n32537) );
  XNOR U32940 ( .A(n32538), .B(n32537), .Z(n32591) );
  NAND U32941 ( .A(n32380), .B(n36309), .Z(n32382) );
  XOR U32942 ( .A(a[106]), .B(n975), .Z(n32517) );
  NANDN U32943 ( .A(n32517), .B(n36311), .Z(n32381) );
  NAND U32944 ( .A(n32382), .B(n32381), .Z(n32589) );
  NAND U32945 ( .A(n35986), .B(n32383), .Z(n32385) );
  XNOR U32946 ( .A(a[108]), .B(b[35]), .Z(n32529) );
  NANDN U32947 ( .A(n32529), .B(n35985), .Z(n32384) );
  AND U32948 ( .A(n32385), .B(n32384), .Z(n32588) );
  XNOR U32949 ( .A(n32589), .B(n32588), .Z(n32590) );
  XOR U32950 ( .A(n32591), .B(n32590), .Z(n32482) );
  NANDN U32951 ( .A(n32386), .B(n34848), .Z(n32388) );
  XOR U32952 ( .A(a[116]), .B(n35375), .Z(n32514) );
  NANDN U32953 ( .A(n32514), .B(n34618), .Z(n32387) );
  NAND U32954 ( .A(n32388), .B(n32387), .Z(n32561) );
  NAND U32955 ( .A(n38326), .B(n32389), .Z(n32391) );
  XOR U32956 ( .A(n38400), .B(n33185), .Z(n32618) );
  NANDN U32957 ( .A(n38273), .B(n32618), .Z(n32390) );
  AND U32958 ( .A(n32391), .B(n32390), .Z(n32559) );
  XOR U32959 ( .A(b[51]), .B(n34852), .Z(n32556) );
  NANDN U32960 ( .A(n32556), .B(n37803), .Z(n32394) );
  NANDN U32961 ( .A(n32392), .B(n37802), .Z(n32393) );
  AND U32962 ( .A(n32394), .B(n32393), .Z(n32560) );
  XOR U32963 ( .A(n32561), .B(n32562), .Z(n32480) );
  NAND U32964 ( .A(n34044), .B(n32395), .Z(n32397) );
  XOR U32965 ( .A(n38134), .B(n34510), .Z(n32648) );
  NANDN U32966 ( .A(n33867), .B(n32648), .Z(n32396) );
  NAND U32967 ( .A(n32397), .B(n32396), .Z(n32597) );
  XNOR U32968 ( .A(a[122]), .B(b[21]), .Z(n32606) );
  OR U32969 ( .A(n32606), .B(n33634), .Z(n32400) );
  NAND U32970 ( .A(n32398), .B(n33464), .Z(n32399) );
  NAND U32971 ( .A(n32400), .B(n32399), .Z(n32594) );
  XNOR U32972 ( .A(b[45]), .B(a[98]), .Z(n32612) );
  NANDN U32973 ( .A(n32612), .B(n37261), .Z(n32403) );
  NAND U32974 ( .A(n32401), .B(n37262), .Z(n32402) );
  AND U32975 ( .A(n32403), .B(n32402), .Z(n32595) );
  XNOR U32976 ( .A(n32594), .B(n32595), .Z(n32596) );
  XOR U32977 ( .A(n32597), .B(n32596), .Z(n32481) );
  XOR U32978 ( .A(n32480), .B(n32481), .Z(n32483) );
  XNOR U32979 ( .A(n32482), .B(n32483), .Z(n32471) );
  XNOR U32980 ( .A(n32470), .B(n32471), .Z(n32510) );
  NANDN U32981 ( .A(n32405), .B(n32404), .Z(n32409) );
  OR U32982 ( .A(n32407), .B(n32406), .Z(n32408) );
  NAND U32983 ( .A(n32409), .B(n32408), .Z(n32511) );
  XNOR U32984 ( .A(n32510), .B(n32511), .Z(n32512) );
  NANDN U32985 ( .A(n32411), .B(n32410), .Z(n32415) );
  NANDN U32986 ( .A(n32413), .B(n32412), .Z(n32414) );
  AND U32987 ( .A(n32415), .B(n32414), .Z(n32513) );
  XOR U32988 ( .A(n32512), .B(n32513), .Z(n32501) );
  OR U32989 ( .A(n32417), .B(n32416), .Z(n32421) );
  NAND U32990 ( .A(n32419), .B(n32418), .Z(n32420) );
  AND U32991 ( .A(n32421), .B(n32420), .Z(n32498) );
  NANDN U32992 ( .A(n32423), .B(n32422), .Z(n32427) );
  OR U32993 ( .A(n32425), .B(n32424), .Z(n32426) );
  AND U32994 ( .A(n32427), .B(n32426), .Z(n32499) );
  XOR U32995 ( .A(n32498), .B(n32499), .Z(n32500) );
  XOR U32996 ( .A(n32501), .B(n32500), .Z(n32663) );
  NANDN U32997 ( .A(n32429), .B(n32428), .Z(n32433) );
  NANDN U32998 ( .A(n32431), .B(n32430), .Z(n32432) );
  NAND U32999 ( .A(n32433), .B(n32432), .Z(n32660) );
  NANDN U33000 ( .A(n32435), .B(n32434), .Z(n32439) );
  NANDN U33001 ( .A(n32437), .B(n32436), .Z(n32438) );
  AND U33002 ( .A(n32439), .B(n32438), .Z(n32661) );
  XNOR U33003 ( .A(n32660), .B(n32661), .Z(n32662) );
  XNOR U33004 ( .A(n32663), .B(n32662), .Z(n32450) );
  XNOR U33005 ( .A(n32451), .B(n32450), .Z(n32452) );
  XNOR U33006 ( .A(n32453), .B(n32452), .Z(n32457) );
  XNOR U33007 ( .A(n32456), .B(n32457), .Z(n32458) );
  XOR U33008 ( .A(n32459), .B(n32458), .Z(n32666) );
  XNOR U33009 ( .A(n32667), .B(n32666), .Z(n32668) );
  XNOR U33010 ( .A(n32669), .B(n32668), .Z(n32447) );
  NAND U33011 ( .A(n32441), .B(n32440), .Z(n32445) );
  NANDN U33012 ( .A(n32443), .B(n32442), .Z(n32444) );
  AND U33013 ( .A(n32445), .B(n32444), .Z(n32448) );
  XOR U33014 ( .A(n32447), .B(n32448), .Z(n32446) );
  XNOR U33015 ( .A(n32449), .B(n32446), .Z(n32670) );
  XOR U33016 ( .A(n32671), .B(n32670), .Z(c[206]) );
  NANDN U33017 ( .A(n32451), .B(n32450), .Z(n32455) );
  NAND U33018 ( .A(n32453), .B(n32452), .Z(n32454) );
  NAND U33019 ( .A(n32455), .B(n32454), .Z(n32895) );
  NANDN U33020 ( .A(n32457), .B(n32456), .Z(n32461) );
  NAND U33021 ( .A(n32459), .B(n32458), .Z(n32460) );
  AND U33022 ( .A(n32461), .B(n32460), .Z(n32894) );
  XNOR U33023 ( .A(n32895), .B(n32894), .Z(n32896) );
  NANDN U33024 ( .A(n32463), .B(n32462), .Z(n32467) );
  NAND U33025 ( .A(n32465), .B(n32464), .Z(n32466) );
  NAND U33026 ( .A(n32467), .B(n32466), .Z(n32873) );
  NANDN U33027 ( .A(n32469), .B(n32468), .Z(n32473) );
  NAND U33028 ( .A(n32471), .B(n32470), .Z(n32472) );
  NAND U33029 ( .A(n32473), .B(n32472), .Z(n32870) );
  NAND U33030 ( .A(n32475), .B(n32474), .Z(n32479) );
  NANDN U33031 ( .A(n32477), .B(n32476), .Z(n32478) );
  NAND U33032 ( .A(n32479), .B(n32478), .Z(n32695) );
  NANDN U33033 ( .A(n32481), .B(n32480), .Z(n32485) );
  NANDN U33034 ( .A(n32483), .B(n32482), .Z(n32484) );
  NAND U33035 ( .A(n32485), .B(n32484), .Z(n32692) );
  NANDN U33036 ( .A(n32487), .B(n32486), .Z(n32491) );
  OR U33037 ( .A(n32489), .B(n32488), .Z(n32490) );
  AND U33038 ( .A(n32491), .B(n32490), .Z(n32693) );
  XNOR U33039 ( .A(n32692), .B(n32693), .Z(n32694) );
  XNOR U33040 ( .A(n32695), .B(n32694), .Z(n32871) );
  XNOR U33041 ( .A(n32870), .B(n32871), .Z(n32872) );
  XOR U33042 ( .A(n32873), .B(n32872), .Z(n32891) );
  NAND U33043 ( .A(n32493), .B(n32492), .Z(n32497) );
  NANDN U33044 ( .A(n32495), .B(n32494), .Z(n32496) );
  NAND U33045 ( .A(n32497), .B(n32496), .Z(n32889) );
  OR U33046 ( .A(n32499), .B(n32498), .Z(n32503) );
  NANDN U33047 ( .A(n32501), .B(n32500), .Z(n32502) );
  NAND U33048 ( .A(n32503), .B(n32502), .Z(n32888) );
  XOR U33049 ( .A(n32889), .B(n32888), .Z(n32890) );
  XOR U33050 ( .A(n32891), .B(n32890), .Z(n32884) );
  NAND U33051 ( .A(n32505), .B(n32504), .Z(n32509) );
  OR U33052 ( .A(n32507), .B(n32506), .Z(n32508) );
  NAND U33053 ( .A(n32509), .B(n32508), .Z(n32683) );
  NANDN U33054 ( .A(n32514), .B(n34848), .Z(n32516) );
  XNOR U33055 ( .A(a[117]), .B(n35375), .Z(n32755) );
  NAND U33056 ( .A(n34618), .B(n32755), .Z(n32515) );
  NAND U33057 ( .A(n32516), .B(n32515), .Z(n32827) );
  NANDN U33058 ( .A(n32517), .B(n36309), .Z(n32519) );
  XNOR U33059 ( .A(a[107]), .B(n975), .Z(n32857) );
  NAND U33060 ( .A(n32857), .B(n36311), .Z(n32518) );
  NAND U33061 ( .A(n32519), .B(n32518), .Z(n32825) );
  NAND U33062 ( .A(n36643), .B(n32520), .Z(n32522) );
  XNOR U33063 ( .A(n976), .B(a[105]), .Z(n32752) );
  NAND U33064 ( .A(n32752), .B(n36553), .Z(n32521) );
  NAND U33065 ( .A(n32522), .B(n32521), .Z(n32826) );
  XNOR U33066 ( .A(n32825), .B(n32826), .Z(n32828) );
  XOR U33067 ( .A(n32827), .B(n32828), .Z(n32869) );
  XNOR U33068 ( .A(a[111]), .B(b[33]), .Z(n32758) );
  NANDN U33069 ( .A(n32758), .B(n35620), .Z(n32525) );
  NANDN U33070 ( .A(n32523), .B(n35621), .Z(n32524) );
  NAND U33071 ( .A(n32525), .B(n32524), .Z(n32800) );
  XNOR U33072 ( .A(a[113]), .B(n973), .Z(n32764) );
  NAND U33073 ( .A(n32764), .B(n35313), .Z(n32528) );
  NANDN U33074 ( .A(n32526), .B(n35311), .Z(n32527) );
  NAND U33075 ( .A(n32528), .B(n32527), .Z(n32797) );
  XOR U33076 ( .A(a[109]), .B(b[35]), .Z(n32749) );
  NAND U33077 ( .A(n35985), .B(n32749), .Z(n32531) );
  NANDN U33078 ( .A(n32529), .B(n35986), .Z(n32530) );
  AND U33079 ( .A(n32531), .B(n32530), .Z(n32798) );
  XNOR U33080 ( .A(n32797), .B(n32798), .Z(n32799) );
  XNOR U33081 ( .A(n32800), .B(n32799), .Z(n32866) );
  NAND U33082 ( .A(n32532), .B(n35188), .Z(n32534) );
  XNOR U33083 ( .A(a[115]), .B(n35540), .Z(n32761) );
  NANDN U33084 ( .A(n34968), .B(n32761), .Z(n32533) );
  NAND U33085 ( .A(n32534), .B(n32533), .Z(n32867) );
  XNOR U33086 ( .A(n32866), .B(n32867), .Z(n32868) );
  XNOR U33087 ( .A(n32869), .B(n32868), .Z(n32730) );
  NANDN U33088 ( .A(n32536), .B(n32535), .Z(n32540) );
  NAND U33089 ( .A(n32538), .B(n32537), .Z(n32539) );
  NAND U33090 ( .A(n32540), .B(n32539), .Z(n32725) );
  NANDN U33091 ( .A(n32542), .B(n32541), .Z(n32545) );
  XNOR U33092 ( .A(a[127]), .B(b[17]), .Z(n32810) );
  NANDN U33093 ( .A(n32810), .B(n32543), .Z(n32544) );
  NAND U33094 ( .A(n32545), .B(n32544), .Z(n32838) );
  XOR U33095 ( .A(b[41]), .B(a[103]), .Z(n32829) );
  NANDN U33096 ( .A(n36905), .B(n32829), .Z(n32548) );
  NANDN U33097 ( .A(n32546), .B(n36807), .Z(n32547) );
  AND U33098 ( .A(n32548), .B(n32547), .Z(n32839) );
  XNOR U33099 ( .A(n32838), .B(n32839), .Z(n32840) );
  AND U33100 ( .A(n32549), .B(b[15]), .Z(n32803) );
  NANDN U33101 ( .A(n985), .B(a[79]), .Z(n32804) );
  XOR U33102 ( .A(n32803), .B(n32804), .Z(n32805) );
  XNOR U33103 ( .A(n32806), .B(n32805), .Z(n32841) );
  XOR U33104 ( .A(n32840), .B(n32841), .Z(n32723) );
  XNOR U33105 ( .A(n38193), .B(b[25]), .Z(n32746) );
  NANDN U33106 ( .A(n34219), .B(n32746), .Z(n32552) );
  NAND U33107 ( .A(n34217), .B(n32550), .Z(n32551) );
  NAND U33108 ( .A(n32552), .B(n32551), .Z(n32845) );
  XOR U33109 ( .A(b[49]), .B(n35628), .Z(n32854) );
  OR U33110 ( .A(n32854), .B(n37756), .Z(n32555) );
  NANDN U33111 ( .A(n32553), .B(n37652), .Z(n32554) );
  NAND U33112 ( .A(n32555), .B(n32554), .Z(n32842) );
  XOR U33113 ( .A(b[51]), .B(n35377), .Z(n32863) );
  NANDN U33114 ( .A(n32863), .B(n37803), .Z(n32558) );
  NANDN U33115 ( .A(n32556), .B(n37802), .Z(n32557) );
  AND U33116 ( .A(n32558), .B(n32557), .Z(n32843) );
  XNOR U33117 ( .A(n32842), .B(n32843), .Z(n32844) );
  XOR U33118 ( .A(n32845), .B(n32844), .Z(n32722) );
  XNOR U33119 ( .A(n32723), .B(n32722), .Z(n32724) );
  XNOR U33120 ( .A(n32725), .B(n32724), .Z(n32707) );
  OR U33121 ( .A(n32560), .B(n32559), .Z(n32564) );
  NANDN U33122 ( .A(n32562), .B(n32561), .Z(n32563) );
  NAND U33123 ( .A(n32564), .B(n32563), .Z(n32704) );
  OR U33124 ( .A(n32565), .B(n32806), .Z(n32569) );
  NANDN U33125 ( .A(n32567), .B(n32566), .Z(n32568) );
  AND U33126 ( .A(n32569), .B(n32568), .Z(n32705) );
  XNOR U33127 ( .A(n32704), .B(n32705), .Z(n32706) );
  XNOR U33128 ( .A(n32707), .B(n32706), .Z(n32728) );
  NANDN U33129 ( .A(n32571), .B(n32570), .Z(n32575) );
  OR U33130 ( .A(n32573), .B(n32572), .Z(n32574) );
  AND U33131 ( .A(n32575), .B(n32574), .Z(n32729) );
  XNOR U33132 ( .A(n32728), .B(n32729), .Z(n32731) );
  XNOR U33133 ( .A(n32730), .B(n32731), .Z(n32878) );
  NANDN U33134 ( .A(n32577), .B(n32576), .Z(n32581) );
  NAND U33135 ( .A(n32579), .B(n32578), .Z(n32580) );
  AND U33136 ( .A(n32581), .B(n32580), .Z(n32877) );
  NANDN U33137 ( .A(n32583), .B(n32582), .Z(n32587) );
  OR U33138 ( .A(n32585), .B(n32584), .Z(n32586) );
  NAND U33139 ( .A(n32587), .B(n32586), .Z(n32687) );
  NANDN U33140 ( .A(n32589), .B(n32588), .Z(n32593) );
  NAND U33141 ( .A(n32591), .B(n32590), .Z(n32592) );
  AND U33142 ( .A(n32593), .B(n32592), .Z(n32698) );
  NANDN U33143 ( .A(n32595), .B(n32594), .Z(n32599) );
  NAND U33144 ( .A(n32597), .B(n32596), .Z(n32598) );
  NAND U33145 ( .A(n32599), .B(n32598), .Z(n32699) );
  NANDN U33146 ( .A(n32601), .B(n32600), .Z(n32605) );
  NAND U33147 ( .A(n32603), .B(n32602), .Z(n32604) );
  NAND U33148 ( .A(n32605), .B(n32604), .Z(n32718) );
  XOR U33149 ( .A(a[123]), .B(b[21]), .Z(n32860) );
  NANDN U33150 ( .A(n33634), .B(n32860), .Z(n32608) );
  NANDN U33151 ( .A(n32606), .B(n33464), .Z(n32607) );
  NAND U33152 ( .A(n32608), .B(n32607), .Z(n32742) );
  XNOR U33153 ( .A(b[61]), .B(a[83]), .Z(n32776) );
  OR U33154 ( .A(n32776), .B(n38371), .Z(n32611) );
  NANDN U33155 ( .A(n32609), .B(n38369), .Z(n32610) );
  AND U33156 ( .A(n32611), .B(n32610), .Z(n32740) );
  XOR U33157 ( .A(b[45]), .B(a[99]), .Z(n32788) );
  NAND U33158 ( .A(n32788), .B(n37261), .Z(n32614) );
  NANDN U33159 ( .A(n32612), .B(n37262), .Z(n32613) );
  AND U33160 ( .A(n32614), .B(n32613), .Z(n32741) );
  XOR U33161 ( .A(n32742), .B(n32743), .Z(n32716) );
  XNOR U33162 ( .A(b[57]), .B(a[87]), .Z(n32782) );
  OR U33163 ( .A(n32782), .B(n965), .Z(n32617) );
  NANDN U33164 ( .A(n32615), .B(n38194), .Z(n32616) );
  NAND U33165 ( .A(n32617), .B(n32616), .Z(n32822) );
  NAND U33166 ( .A(n38326), .B(n32618), .Z(n32620) );
  XNOR U33167 ( .A(n38400), .B(a[85]), .Z(n32785) );
  NANDN U33168 ( .A(n38273), .B(n32785), .Z(n32619) );
  NAND U33169 ( .A(n32620), .B(n32619), .Z(n32819) );
  NAND U33170 ( .A(n37469), .B(n32621), .Z(n32623) );
  XNOR U33171 ( .A(n978), .B(a[97]), .Z(n32851) );
  NAND U33172 ( .A(n32851), .B(n37471), .Z(n32622) );
  AND U33173 ( .A(n32623), .B(n32622), .Z(n32820) );
  XNOR U33174 ( .A(n32819), .B(n32820), .Z(n32821) );
  XOR U33175 ( .A(n32822), .B(n32821), .Z(n32717) );
  XOR U33176 ( .A(n32716), .B(n32717), .Z(n32719) );
  XOR U33177 ( .A(n32718), .B(n32719), .Z(n32700) );
  XNOR U33178 ( .A(n32687), .B(n32686), .Z(n32688) );
  NANDN U33179 ( .A(n32625), .B(n32624), .Z(n32629) );
  NAND U33180 ( .A(n32627), .B(n32626), .Z(n32628) );
  NAND U33181 ( .A(n32629), .B(n32628), .Z(n32713) );
  NANDN U33182 ( .A(n32631), .B(n32630), .Z(n32635) );
  NAND U33183 ( .A(n32633), .B(n32632), .Z(n32634) );
  NAND U33184 ( .A(n32635), .B(n32634), .Z(n32710) );
  XNOR U33185 ( .A(b[43]), .B(a[101]), .Z(n32773) );
  NANDN U33186 ( .A(n32773), .B(n37068), .Z(n32638) );
  NANDN U33187 ( .A(n32636), .B(n37069), .Z(n32637) );
  NAND U33188 ( .A(n32638), .B(n32637), .Z(n32794) );
  NAND U33189 ( .A(n33283), .B(n32639), .Z(n32641) );
  XNOR U33190 ( .A(a[125]), .B(n33020), .Z(n32779) );
  NANDN U33191 ( .A(n33021), .B(n32779), .Z(n32640) );
  NAND U33192 ( .A(n32641), .B(n32640), .Z(n32791) );
  XNOR U33193 ( .A(b[63]), .B(a[81]), .Z(n32816) );
  NANDN U33194 ( .A(n32816), .B(n38422), .Z(n32644) );
  NANDN U33195 ( .A(n32642), .B(n38423), .Z(n32643) );
  AND U33196 ( .A(n32644), .B(n32643), .Z(n32792) );
  XNOR U33197 ( .A(n32791), .B(n32792), .Z(n32793) );
  XNOR U33198 ( .A(n32794), .B(n32793), .Z(n32734) );
  XNOR U33199 ( .A(b[53]), .B(a[91]), .Z(n32832) );
  NANDN U33200 ( .A(n32832), .B(n37940), .Z(n32647) );
  NANDN U33201 ( .A(n32645), .B(n37941), .Z(n32646) );
  NAND U33202 ( .A(n32647), .B(n32646), .Z(n32770) );
  NAND U33203 ( .A(n34044), .B(n32648), .Z(n32650) );
  XNOR U33204 ( .A(a[121]), .B(n34510), .Z(n32848) );
  NANDN U33205 ( .A(n33867), .B(n32848), .Z(n32649) );
  NAND U33206 ( .A(n32650), .B(n32649), .Z(n32767) );
  XNOR U33207 ( .A(b[55]), .B(a[89]), .Z(n32835) );
  NANDN U33208 ( .A(n32835), .B(n38075), .Z(n32653) );
  NANDN U33209 ( .A(n32651), .B(n38073), .Z(n32652) );
  AND U33210 ( .A(n32653), .B(n32652), .Z(n32768) );
  XNOR U33211 ( .A(n32767), .B(n32768), .Z(n32769) );
  XOR U33212 ( .A(n32770), .B(n32769), .Z(n32735) );
  XOR U33213 ( .A(n32734), .B(n32735), .Z(n32737) );
  NANDN U33214 ( .A(n32655), .B(n32654), .Z(n32659) );
  NAND U33215 ( .A(n32657), .B(n32656), .Z(n32658) );
  NAND U33216 ( .A(n32659), .B(n32658), .Z(n32736) );
  XOR U33217 ( .A(n32710), .B(n32711), .Z(n32712) );
  XOR U33218 ( .A(n32713), .B(n32712), .Z(n32689) );
  XNOR U33219 ( .A(n32688), .B(n32689), .Z(n32876) );
  XNOR U33220 ( .A(n32878), .B(n32879), .Z(n32680) );
  XOR U33221 ( .A(n32681), .B(n32680), .Z(n32682) );
  XNOR U33222 ( .A(n32683), .B(n32682), .Z(n32882) );
  NANDN U33223 ( .A(n32661), .B(n32660), .Z(n32665) );
  NANDN U33224 ( .A(n32663), .B(n32662), .Z(n32664) );
  NAND U33225 ( .A(n32665), .B(n32664), .Z(n32883) );
  XOR U33226 ( .A(n32882), .B(n32883), .Z(n32885) );
  XOR U33227 ( .A(n32884), .B(n32885), .Z(n32897) );
  XOR U33228 ( .A(n32896), .B(n32897), .Z(n32674) );
  XNOR U33229 ( .A(n32674), .B(n32675), .Z(n32677) );
  XNOR U33230 ( .A(n32676), .B(n32677), .Z(n32672) );
  OR U33231 ( .A(n32671), .B(n32670), .Z(n32673) );
  XNOR U33232 ( .A(n32672), .B(n32673), .Z(c[207]) );
  NANDN U33233 ( .A(n32673), .B(n32672), .Z(n33115) );
  NAND U33234 ( .A(n32675), .B(n32674), .Z(n32679) );
  NANDN U33235 ( .A(n32677), .B(n32676), .Z(n32678) );
  AND U33236 ( .A(n32679), .B(n32678), .Z(n32903) );
  OR U33237 ( .A(n32681), .B(n32680), .Z(n32685) );
  NAND U33238 ( .A(n32683), .B(n32682), .Z(n32684) );
  NAND U33239 ( .A(n32685), .B(n32684), .Z(n32905) );
  NAND U33240 ( .A(n32687), .B(n32686), .Z(n32691) );
  OR U33241 ( .A(n32689), .B(n32688), .Z(n32690) );
  NAND U33242 ( .A(n32691), .B(n32690), .Z(n32986) );
  NANDN U33243 ( .A(n32693), .B(n32692), .Z(n32697) );
  NAND U33244 ( .A(n32695), .B(n32694), .Z(n32696) );
  AND U33245 ( .A(n32697), .B(n32696), .Z(n32987) );
  XNOR U33246 ( .A(n32986), .B(n32987), .Z(n32988) );
  OR U33247 ( .A(n32699), .B(n32698), .Z(n32703) );
  NANDN U33248 ( .A(n32701), .B(n32700), .Z(n32702) );
  NAND U33249 ( .A(n32703), .B(n32702), .Z(n32982) );
  NANDN U33250 ( .A(n32705), .B(n32704), .Z(n32709) );
  NANDN U33251 ( .A(n32707), .B(n32706), .Z(n32708) );
  NAND U33252 ( .A(n32709), .B(n32708), .Z(n32981) );
  OR U33253 ( .A(n32711), .B(n32710), .Z(n32715) );
  NANDN U33254 ( .A(n32713), .B(n32712), .Z(n32714) );
  NAND U33255 ( .A(n32715), .B(n32714), .Z(n33105) );
  NANDN U33256 ( .A(n32717), .B(n32716), .Z(n32721) );
  OR U33257 ( .A(n32719), .B(n32718), .Z(n32720) );
  NAND U33258 ( .A(n32721), .B(n32720), .Z(n33102) );
  NANDN U33259 ( .A(n32723), .B(n32722), .Z(n32727) );
  NAND U33260 ( .A(n32725), .B(n32724), .Z(n32726) );
  NAND U33261 ( .A(n32727), .B(n32726), .Z(n33103) );
  XNOR U33262 ( .A(n33102), .B(n33103), .Z(n33104) );
  XOR U33263 ( .A(n33105), .B(n33104), .Z(n32980) );
  XOR U33264 ( .A(n32981), .B(n32980), .Z(n32983) );
  XOR U33265 ( .A(n32982), .B(n32983), .Z(n32989) );
  XOR U33266 ( .A(n32988), .B(n32989), .Z(n32912) );
  NAND U33267 ( .A(n32729), .B(n32728), .Z(n32733) );
  NANDN U33268 ( .A(n32731), .B(n32730), .Z(n32732) );
  NAND U33269 ( .A(n32733), .B(n32732), .Z(n32918) );
  NANDN U33270 ( .A(n32735), .B(n32734), .Z(n32739) );
  OR U33271 ( .A(n32737), .B(n32736), .Z(n32738) );
  NAND U33272 ( .A(n32739), .B(n32738), .Z(n33096) );
  OR U33273 ( .A(n32741), .B(n32740), .Z(n32745) );
  NANDN U33274 ( .A(n32743), .B(n32742), .Z(n32744) );
  NAND U33275 ( .A(n32745), .B(n32744), .Z(n33085) );
  XNOR U33276 ( .A(n38134), .B(b[25]), .Z(n33036) );
  NANDN U33277 ( .A(n34219), .B(n33036), .Z(n32748) );
  NAND U33278 ( .A(n34217), .B(n32746), .Z(n32747) );
  NAND U33279 ( .A(n32748), .B(n32747), .Z(n33016) );
  XNOR U33280 ( .A(a[110]), .B(b[35]), .Z(n32953) );
  NANDN U33281 ( .A(n32953), .B(n35985), .Z(n32751) );
  NAND U33282 ( .A(n32749), .B(n35986), .Z(n32750) );
  NAND U33283 ( .A(n32751), .B(n32750), .Z(n33013) );
  XOR U33284 ( .A(n36909), .B(n976), .Z(n33030) );
  NAND U33285 ( .A(n33030), .B(n36553), .Z(n32754) );
  NAND U33286 ( .A(n32752), .B(n36643), .Z(n32753) );
  AND U33287 ( .A(n32754), .B(n32753), .Z(n33014) );
  XNOR U33288 ( .A(n33013), .B(n33014), .Z(n33015) );
  XNOR U33289 ( .A(n33016), .B(n33015), .Z(n32995) );
  NAND U33290 ( .A(n32755), .B(n34848), .Z(n32757) );
  XOR U33291 ( .A(n38143), .B(n35375), .Z(n32947) );
  NAND U33292 ( .A(n34618), .B(n32947), .Z(n32756) );
  NAND U33293 ( .A(n32757), .B(n32756), .Z(n33057) );
  XOR U33294 ( .A(a[112]), .B(n974), .Z(n33075) );
  NANDN U33295 ( .A(n33075), .B(n35620), .Z(n32760) );
  NANDN U33296 ( .A(n32758), .B(n35621), .Z(n32759) );
  NAND U33297 ( .A(n32760), .B(n32759), .Z(n33054) );
  NAND U33298 ( .A(n32761), .B(n35188), .Z(n32763) );
  XOR U33299 ( .A(n38046), .B(n35540), .Z(n33051) );
  NANDN U33300 ( .A(n34968), .B(n33051), .Z(n32762) );
  AND U33301 ( .A(n32763), .B(n32762), .Z(n33055) );
  XNOR U33302 ( .A(n33054), .B(n33055), .Z(n33056) );
  XNOR U33303 ( .A(n33057), .B(n33056), .Z(n32992) );
  NAND U33304 ( .A(n32764), .B(n35311), .Z(n32766) );
  XNOR U33305 ( .A(n37873), .B(b[31]), .Z(n33048) );
  NAND U33306 ( .A(n33048), .B(n35313), .Z(n32765) );
  NAND U33307 ( .A(n32766), .B(n32765), .Z(n32993) );
  XNOR U33308 ( .A(n32992), .B(n32993), .Z(n32994) );
  XOR U33309 ( .A(n32995), .B(n32994), .Z(n33084) );
  XOR U33310 ( .A(n33085), .B(n33084), .Z(n33087) );
  NANDN U33311 ( .A(n32768), .B(n32767), .Z(n32772) );
  NAND U33312 ( .A(n32770), .B(n32769), .Z(n32771) );
  NAND U33313 ( .A(n32772), .B(n32771), .Z(n32931) );
  XOR U33314 ( .A(b[43]), .B(n36420), .Z(n33024) );
  NANDN U33315 ( .A(n33024), .B(n37068), .Z(n32775) );
  NANDN U33316 ( .A(n32773), .B(n37069), .Z(n32774) );
  NAND U33317 ( .A(n32775), .B(n32774), .Z(n32971) );
  XOR U33318 ( .A(b[61]), .B(n33185), .Z(n32950) );
  OR U33319 ( .A(n32950), .B(n38371), .Z(n32778) );
  NANDN U33320 ( .A(n32776), .B(n38369), .Z(n32777) );
  NAND U33321 ( .A(n32778), .B(n32777), .Z(n32968) );
  NAND U33322 ( .A(n33283), .B(n32779), .Z(n32781) );
  XOR U33323 ( .A(n987), .B(n33020), .Z(n33019) );
  NANDN U33324 ( .A(n33021), .B(n33019), .Z(n32780) );
  AND U33325 ( .A(n32781), .B(n32780), .Z(n32969) );
  XNOR U33326 ( .A(n32968), .B(n32969), .Z(n32970) );
  XOR U33327 ( .A(n32971), .B(n32970), .Z(n32928) );
  XOR U33328 ( .A(b[57]), .B(n34048), .Z(n33045) );
  OR U33329 ( .A(n33045), .B(n965), .Z(n32784) );
  NANDN U33330 ( .A(n32782), .B(n38194), .Z(n32783) );
  NAND U33331 ( .A(n32784), .B(n32783), .Z(n32977) );
  NAND U33332 ( .A(n38326), .B(n32785), .Z(n32787) );
  XOR U33333 ( .A(n38400), .B(n33628), .Z(n33081) );
  NANDN U33334 ( .A(n38273), .B(n33081), .Z(n32786) );
  NAND U33335 ( .A(n32787), .B(n32786), .Z(n32974) );
  XNOR U33336 ( .A(b[45]), .B(a[100]), .Z(n33066) );
  NANDN U33337 ( .A(n33066), .B(n37261), .Z(n32790) );
  NAND U33338 ( .A(n32788), .B(n37262), .Z(n32789) );
  AND U33339 ( .A(n32790), .B(n32789), .Z(n32975) );
  XNOR U33340 ( .A(n32974), .B(n32975), .Z(n32976) );
  XOR U33341 ( .A(n32977), .B(n32976), .Z(n32929) );
  XNOR U33342 ( .A(n32928), .B(n32929), .Z(n32930) );
  XNOR U33343 ( .A(n32931), .B(n32930), .Z(n33086) );
  XNOR U33344 ( .A(n33087), .B(n33086), .Z(n33097) );
  XNOR U33345 ( .A(n33096), .B(n33097), .Z(n33098) );
  NANDN U33346 ( .A(n32792), .B(n32791), .Z(n32796) );
  NAND U33347 ( .A(n32794), .B(n32793), .Z(n32795) );
  NAND U33348 ( .A(n32796), .B(n32795), .Z(n32937) );
  NANDN U33349 ( .A(n32798), .B(n32797), .Z(n32802) );
  NAND U33350 ( .A(n32800), .B(n32799), .Z(n32801) );
  NAND U33351 ( .A(n32802), .B(n32801), .Z(n32996) );
  OR U33352 ( .A(n32804), .B(n32803), .Z(n32808) );
  NAND U33353 ( .A(n32806), .B(n32805), .Z(n32807) );
  AND U33354 ( .A(n32808), .B(n32807), .Z(n32997) );
  XNOR U33355 ( .A(n32996), .B(n32997), .Z(n32998) );
  XNOR U33356 ( .A(b[17]), .B(n32809), .Z(n32813) );
  NAND U33357 ( .A(n32811), .B(n32810), .Z(n32812) );
  NAND U33358 ( .A(n32813), .B(n32812), .Z(n33004) );
  ANDN U33359 ( .B(b[63]), .A(n32814), .Z(n33152) );
  XOR U33360 ( .A(b[63]), .B(n32815), .Z(n33072) );
  NANDN U33361 ( .A(n33072), .B(n38422), .Z(n32818) );
  NANDN U33362 ( .A(n32816), .B(n38423), .Z(n32817) );
  AND U33363 ( .A(n32818), .B(n32817), .Z(n33002) );
  XNOR U33364 ( .A(n32998), .B(n32999), .Z(n32934) );
  NANDN U33365 ( .A(n32820), .B(n32819), .Z(n32824) );
  NAND U33366 ( .A(n32822), .B(n32821), .Z(n32823) );
  NAND U33367 ( .A(n32824), .B(n32823), .Z(n32935) );
  XNOR U33368 ( .A(n32934), .B(n32935), .Z(n32936) );
  XOR U33369 ( .A(n32937), .B(n32936), .Z(n33099) );
  XOR U33370 ( .A(n33098), .B(n33099), .Z(n32917) );
  XNOR U33371 ( .A(b[41]), .B(a[104]), .Z(n33033) );
  OR U33372 ( .A(n33033), .B(n36905), .Z(n32831) );
  NAND U33373 ( .A(n32829), .B(n36807), .Z(n32830) );
  NAND U33374 ( .A(n32831), .B(n32830), .Z(n33010) );
  XOR U33375 ( .A(b[53]), .B(n34852), .Z(n32959) );
  NANDN U33376 ( .A(n32959), .B(n37940), .Z(n32834) );
  NANDN U33377 ( .A(n32832), .B(n37941), .Z(n32833) );
  NAND U33378 ( .A(n32834), .B(n32833), .Z(n33007) );
  XOR U33379 ( .A(b[55]), .B(n34851), .Z(n33078) );
  NANDN U33380 ( .A(n33078), .B(n38075), .Z(n32837) );
  NANDN U33381 ( .A(n32835), .B(n38073), .Z(n32836) );
  AND U33382 ( .A(n32837), .B(n32836), .Z(n33008) );
  XNOR U33383 ( .A(n33007), .B(n33008), .Z(n33009) );
  XOR U33384 ( .A(n33010), .B(n33009), .Z(n32922) );
  XNOR U33385 ( .A(n32922), .B(n32923), .Z(n32924) );
  XNOR U33386 ( .A(n32925), .B(n32924), .Z(n33093) );
  NANDN U33387 ( .A(n32843), .B(n32842), .Z(n32847) );
  NAND U33388 ( .A(n32845), .B(n32844), .Z(n32846) );
  NAND U33389 ( .A(n32847), .B(n32846), .Z(n32940) );
  NAND U33390 ( .A(n34044), .B(n32848), .Z(n32850) );
  XOR U33391 ( .A(n38251), .B(n34510), .Z(n33039) );
  NANDN U33392 ( .A(n33867), .B(n33039), .Z(n32849) );
  NAND U33393 ( .A(n32850), .B(n32849), .Z(n32965) );
  NAND U33394 ( .A(n37469), .B(n32851), .Z(n32853) );
  XOR U33395 ( .A(n978), .B(n35783), .Z(n33042) );
  NAND U33396 ( .A(n33042), .B(n37471), .Z(n32852) );
  NAND U33397 ( .A(n32853), .B(n32852), .Z(n32962) );
  XOR U33398 ( .A(b[49]), .B(n35545), .Z(n32956) );
  OR U33399 ( .A(n32956), .B(n37756), .Z(n32856) );
  NANDN U33400 ( .A(n32854), .B(n37652), .Z(n32855) );
  AND U33401 ( .A(n32856), .B(n32855), .Z(n32963) );
  XNOR U33402 ( .A(n32962), .B(n32963), .Z(n32964) );
  XNOR U33403 ( .A(n32965), .B(n32964), .Z(n32938) );
  XOR U33404 ( .A(a[108]), .B(n975), .Z(n33027) );
  NANDN U33405 ( .A(n33027), .B(n36311), .Z(n32859) );
  NAND U33406 ( .A(n32857), .B(n36309), .Z(n32858) );
  NAND U33407 ( .A(n32859), .B(n32858), .Z(n33063) );
  XNOR U33408 ( .A(a[124]), .B(b[21]), .Z(n33069) );
  OR U33409 ( .A(n33069), .B(n33634), .Z(n32862) );
  NAND U33410 ( .A(n32860), .B(n33464), .Z(n32861) );
  NAND U33411 ( .A(n32862), .B(n32861), .Z(n33060) );
  XOR U33412 ( .A(b[51]), .B(n35191), .Z(n32944) );
  NANDN U33413 ( .A(n32944), .B(n37803), .Z(n32865) );
  NANDN U33414 ( .A(n32863), .B(n37802), .Z(n32864) );
  AND U33415 ( .A(n32865), .B(n32864), .Z(n33061) );
  XNOR U33416 ( .A(n33060), .B(n33061), .Z(n33062) );
  XOR U33417 ( .A(n33063), .B(n33062), .Z(n32939) );
  XOR U33418 ( .A(n32938), .B(n32939), .Z(n32941) );
  XNOR U33419 ( .A(n32940), .B(n32941), .Z(n33090) );
  XNOR U33420 ( .A(n33090), .B(n33091), .Z(n33092) );
  XOR U33421 ( .A(n33093), .B(n33092), .Z(n32916) );
  XNOR U33422 ( .A(n32917), .B(n32916), .Z(n32919) );
  XNOR U33423 ( .A(n32918), .B(n32919), .Z(n32910) );
  NANDN U33424 ( .A(n32871), .B(n32870), .Z(n32875) );
  NAND U33425 ( .A(n32873), .B(n32872), .Z(n32874) );
  AND U33426 ( .A(n32875), .B(n32874), .Z(n32911) );
  XNOR U33427 ( .A(n32910), .B(n32911), .Z(n32913) );
  XNOR U33428 ( .A(n32912), .B(n32913), .Z(n32904) );
  XOR U33429 ( .A(n32905), .B(n32904), .Z(n32907) );
  OR U33430 ( .A(n32877), .B(n32876), .Z(n32881) );
  OR U33431 ( .A(n32879), .B(n32878), .Z(n32880) );
  NAND U33432 ( .A(n32881), .B(n32880), .Z(n32906) );
  XNOR U33433 ( .A(n32907), .B(n32906), .Z(n33108) );
  NANDN U33434 ( .A(n32883), .B(n32882), .Z(n32887) );
  OR U33435 ( .A(n32885), .B(n32884), .Z(n32886) );
  NAND U33436 ( .A(n32887), .B(n32886), .Z(n33109) );
  XNOR U33437 ( .A(n33108), .B(n33109), .Z(n33110) );
  OR U33438 ( .A(n32889), .B(n32888), .Z(n32893) );
  NANDN U33439 ( .A(n32891), .B(n32890), .Z(n32892) );
  AND U33440 ( .A(n32893), .B(n32892), .Z(n33111) );
  XNOR U33441 ( .A(n33110), .B(n33111), .Z(n32901) );
  NANDN U33442 ( .A(n32895), .B(n32894), .Z(n32899) );
  NAND U33443 ( .A(n32897), .B(n32896), .Z(n32898) );
  AND U33444 ( .A(n32899), .B(n32898), .Z(n32902) );
  XOR U33445 ( .A(n32901), .B(n32902), .Z(n32900) );
  XNOR U33446 ( .A(n32903), .B(n32900), .Z(n33114) );
  XOR U33447 ( .A(n33115), .B(n33114), .Z(c[208]) );
  NANDN U33448 ( .A(n32905), .B(n32904), .Z(n32909) );
  OR U33449 ( .A(n32907), .B(n32906), .Z(n32908) );
  NAND U33450 ( .A(n32909), .B(n32908), .Z(n33124) );
  NAND U33451 ( .A(n32911), .B(n32910), .Z(n32915) );
  NANDN U33452 ( .A(n32913), .B(n32912), .Z(n32914) );
  NAND U33453 ( .A(n32915), .B(n32914), .Z(n33123) );
  NAND U33454 ( .A(n32917), .B(n32916), .Z(n32921) );
  NANDN U33455 ( .A(n32919), .B(n32918), .Z(n32920) );
  NAND U33456 ( .A(n32921), .B(n32920), .Z(n33131) );
  OR U33457 ( .A(n32923), .B(n32922), .Z(n32927) );
  OR U33458 ( .A(n32925), .B(n32924), .Z(n32926) );
  NAND U33459 ( .A(n32927), .B(n32926), .Z(n33325) );
  OR U33460 ( .A(n32929), .B(n32928), .Z(n32933) );
  OR U33461 ( .A(n32931), .B(n32930), .Z(n32932) );
  AND U33462 ( .A(n32933), .B(n32932), .Z(n33326) );
  XNOR U33463 ( .A(n33325), .B(n33326), .Z(n33327) );
  NANDN U33464 ( .A(n32939), .B(n32938), .Z(n32943) );
  OR U33465 ( .A(n32941), .B(n32940), .Z(n32942) );
  NAND U33466 ( .A(n32943), .B(n32942), .Z(n33201) );
  XOR U33467 ( .A(b[51]), .B(n35628), .Z(n33252) );
  NANDN U33468 ( .A(n33252), .B(n37803), .Z(n32946) );
  NANDN U33469 ( .A(n32944), .B(n37802), .Z(n32945) );
  NAND U33470 ( .A(n32946), .B(n32945), .Z(n33176) );
  NAND U33471 ( .A(n34848), .B(n32947), .Z(n32949) );
  XOR U33472 ( .A(n38193), .B(n35375), .Z(n33228) );
  NAND U33473 ( .A(n34618), .B(n33228), .Z(n32948) );
  NAND U33474 ( .A(n32949), .B(n32948), .Z(n33173) );
  XNOR U33475 ( .A(b[61]), .B(a[85]), .Z(n33182) );
  OR U33476 ( .A(n33182), .B(n38371), .Z(n32952) );
  NANDN U33477 ( .A(n32950), .B(n38369), .Z(n32951) );
  AND U33478 ( .A(n32952), .B(n32951), .Z(n33174) );
  XNOR U33479 ( .A(n33173), .B(n33174), .Z(n33175) );
  XNOR U33480 ( .A(n33176), .B(n33175), .Z(n33210) );
  XOR U33481 ( .A(a[111]), .B(b[35]), .Z(n33213) );
  NAND U33482 ( .A(n35985), .B(n33213), .Z(n32955) );
  NANDN U33483 ( .A(n32953), .B(n35986), .Z(n32954) );
  NAND U33484 ( .A(n32955), .B(n32954), .Z(n33279) );
  XNOR U33485 ( .A(b[49]), .B(a[97]), .Z(n33222) );
  OR U33486 ( .A(n33222), .B(n37756), .Z(n32958) );
  NANDN U33487 ( .A(n32956), .B(n37652), .Z(n32957) );
  NAND U33488 ( .A(n32958), .B(n32957), .Z(n33276) );
  XOR U33489 ( .A(b[53]), .B(n35377), .Z(n33219) );
  NANDN U33490 ( .A(n33219), .B(n37940), .Z(n32961) );
  NANDN U33491 ( .A(n32959), .B(n37941), .Z(n32960) );
  AND U33492 ( .A(n32961), .B(n32960), .Z(n33277) );
  XNOR U33493 ( .A(n33276), .B(n33277), .Z(n33278) );
  XNOR U33494 ( .A(n33279), .B(n33278), .Z(n33207) );
  NANDN U33495 ( .A(n32963), .B(n32962), .Z(n32967) );
  NAND U33496 ( .A(n32965), .B(n32964), .Z(n32966) );
  NAND U33497 ( .A(n32967), .B(n32966), .Z(n33208) );
  XNOR U33498 ( .A(n33207), .B(n33208), .Z(n33209) );
  XOR U33499 ( .A(n33210), .B(n33209), .Z(n33322) );
  NANDN U33500 ( .A(n32969), .B(n32968), .Z(n32973) );
  NAND U33501 ( .A(n32971), .B(n32970), .Z(n32972) );
  AND U33502 ( .A(n32973), .B(n32972), .Z(n33319) );
  NANDN U33503 ( .A(n32975), .B(n32974), .Z(n32979) );
  NAND U33504 ( .A(n32977), .B(n32976), .Z(n32978) );
  AND U33505 ( .A(n32979), .B(n32978), .Z(n33320) );
  XNOR U33506 ( .A(n33322), .B(n33321), .Z(n33202) );
  XNOR U33507 ( .A(n33201), .B(n33202), .Z(n33203) );
  XNOR U33508 ( .A(n33204), .B(n33203), .Z(n33328) );
  XNOR U33509 ( .A(n33327), .B(n33328), .Z(n33128) );
  NANDN U33510 ( .A(n32981), .B(n32980), .Z(n32985) );
  NANDN U33511 ( .A(n32983), .B(n32982), .Z(n32984) );
  NAND U33512 ( .A(n32985), .B(n32984), .Z(n33129) );
  XNOR U33513 ( .A(n33131), .B(n33130), .Z(n33135) );
  NANDN U33514 ( .A(n32987), .B(n32986), .Z(n32991) );
  NANDN U33515 ( .A(n32989), .B(n32988), .Z(n32990) );
  AND U33516 ( .A(n32991), .B(n32990), .Z(n33134) );
  XNOR U33517 ( .A(n33135), .B(n33134), .Z(n33136) );
  NANDN U33518 ( .A(n32997), .B(n32996), .Z(n33001) );
  NAND U33519 ( .A(n32999), .B(n32998), .Z(n33000) );
  NAND U33520 ( .A(n33001), .B(n33000), .Z(n33196) );
  XNOR U33521 ( .A(n33195), .B(n33196), .Z(n33197) );
  OR U33522 ( .A(n33002), .B(n33152), .Z(n33006) );
  NANDN U33523 ( .A(n33004), .B(n33003), .Z(n33005) );
  NAND U33524 ( .A(n33006), .B(n33005), .Z(n33309) );
  NANDN U33525 ( .A(n33008), .B(n33007), .Z(n33012) );
  NAND U33526 ( .A(n33010), .B(n33009), .Z(n33011) );
  AND U33527 ( .A(n33012), .B(n33011), .Z(n33307) );
  NANDN U33528 ( .A(n33014), .B(n33013), .Z(n33018) );
  NAND U33529 ( .A(n33016), .B(n33015), .Z(n33017) );
  NAND U33530 ( .A(n33018), .B(n33017), .Z(n33170) );
  NAND U33531 ( .A(n33283), .B(n33019), .Z(n33023) );
  XOR U33532 ( .A(n38463), .B(n33020), .Z(n33282) );
  NANDN U33533 ( .A(n33021), .B(n33282), .Z(n33022) );
  NAND U33534 ( .A(n33023), .B(n33022), .Z(n33189) );
  XNOR U33535 ( .A(b[43]), .B(a[103]), .Z(n33158) );
  NANDN U33536 ( .A(n33158), .B(n37068), .Z(n33026) );
  NANDN U33537 ( .A(n33024), .B(n37069), .Z(n33025) );
  AND U33538 ( .A(n33026), .B(n33025), .Z(n33190) );
  XNOR U33539 ( .A(n33189), .B(n33190), .Z(n33191) );
  NANDN U33540 ( .A(n985), .B(a[81]), .Z(n33155) );
  XOR U33541 ( .A(n33152), .B(n33153), .Z(n33154) );
  XOR U33542 ( .A(n33155), .B(n33154), .Z(n33192) );
  XOR U33543 ( .A(n33191), .B(n33192), .Z(n33167) );
  NANDN U33544 ( .A(n33027), .B(n36309), .Z(n33029) );
  XNOR U33545 ( .A(a[109]), .B(n975), .Z(n33267) );
  NAND U33546 ( .A(n33267), .B(n36311), .Z(n33028) );
  AND U33547 ( .A(n33029), .B(n33028), .Z(n33149) );
  NAND U33548 ( .A(n36643), .B(n33030), .Z(n33032) );
  XNOR U33549 ( .A(a[107]), .B(n976), .Z(n33270) );
  NAND U33550 ( .A(n33270), .B(n36553), .Z(n33031) );
  AND U33551 ( .A(n33032), .B(n33031), .Z(n33146) );
  XOR U33552 ( .A(b[41]), .B(a[105]), .Z(n33273) );
  NANDN U33553 ( .A(n36905), .B(n33273), .Z(n33035) );
  NANDN U33554 ( .A(n33033), .B(n36807), .Z(n33034) );
  AND U33555 ( .A(n33035), .B(n33034), .Z(n33147) );
  XNOR U33556 ( .A(n33146), .B(n33147), .Z(n33148) );
  XNOR U33557 ( .A(n33167), .B(n33168), .Z(n33169) );
  XNOR U33558 ( .A(n33170), .B(n33169), .Z(n33308) );
  XOR U33559 ( .A(n33309), .B(n33310), .Z(n33303) );
  XOR U33560 ( .A(a[121]), .B(b[25]), .Z(n33161) );
  NANDN U33561 ( .A(n34219), .B(n33161), .Z(n33038) );
  NAND U33562 ( .A(n34217), .B(n33036), .Z(n33037) );
  NAND U33563 ( .A(n33038), .B(n33037), .Z(n33292) );
  NAND U33564 ( .A(n34044), .B(n33039), .Z(n33041) );
  XNOR U33565 ( .A(a[123]), .B(n34510), .Z(n33164) );
  NANDN U33566 ( .A(n33867), .B(n33164), .Z(n33040) );
  NAND U33567 ( .A(n33041), .B(n33040), .Z(n33289) );
  NAND U33568 ( .A(n37469), .B(n33042), .Z(n33044) );
  XNOR U33569 ( .A(n978), .B(a[99]), .Z(n33216) );
  NAND U33570 ( .A(n33216), .B(n37471), .Z(n33043) );
  AND U33571 ( .A(n33044), .B(n33043), .Z(n33290) );
  XNOR U33572 ( .A(n33289), .B(n33290), .Z(n33291) );
  XNOR U33573 ( .A(n33292), .B(n33291), .Z(n33295) );
  XNOR U33574 ( .A(b[57]), .B(a[89]), .Z(n33243) );
  OR U33575 ( .A(n33243), .B(n965), .Z(n33047) );
  NANDN U33576 ( .A(n33045), .B(n38194), .Z(n33046) );
  NAND U33577 ( .A(n33047), .B(n33046), .Z(n33258) );
  XNOR U33578 ( .A(a[115]), .B(b[31]), .Z(n33246) );
  NANDN U33579 ( .A(n33246), .B(n35313), .Z(n33050) );
  NAND U33580 ( .A(n33048), .B(n35311), .Z(n33049) );
  NAND U33581 ( .A(n33050), .B(n33049), .Z(n33255) );
  NAND U33582 ( .A(n35188), .B(n33051), .Z(n33053) );
  XNOR U33583 ( .A(a[117]), .B(n35540), .Z(n33249) );
  NANDN U33584 ( .A(n34968), .B(n33249), .Z(n33052) );
  AND U33585 ( .A(n33053), .B(n33052), .Z(n33256) );
  XNOR U33586 ( .A(n33255), .B(n33256), .Z(n33257) );
  XOR U33587 ( .A(n33258), .B(n33257), .Z(n33296) );
  XNOR U33588 ( .A(n33295), .B(n33296), .Z(n33297) );
  NANDN U33589 ( .A(n33055), .B(n33054), .Z(n33059) );
  NAND U33590 ( .A(n33057), .B(n33056), .Z(n33058) );
  AND U33591 ( .A(n33059), .B(n33058), .Z(n33298) );
  XNOR U33592 ( .A(n33297), .B(n33298), .Z(n33302) );
  NANDN U33593 ( .A(n33061), .B(n33060), .Z(n33065) );
  NAND U33594 ( .A(n33063), .B(n33062), .Z(n33064) );
  NAND U33595 ( .A(n33065), .B(n33064), .Z(n33316) );
  XOR U33596 ( .A(b[45]), .B(a[101]), .Z(n33179) );
  NAND U33597 ( .A(n33179), .B(n37261), .Z(n33068) );
  NANDN U33598 ( .A(n33066), .B(n37262), .Z(n33067) );
  NAND U33599 ( .A(n33068), .B(n33067), .Z(n33264) );
  XOR U33600 ( .A(a[125]), .B(b[21]), .Z(n33286) );
  NANDN U33601 ( .A(n33634), .B(n33286), .Z(n33071) );
  NANDN U33602 ( .A(n33069), .B(n33464), .Z(n33070) );
  NAND U33603 ( .A(n33071), .B(n33070), .Z(n33261) );
  XNOR U33604 ( .A(b[63]), .B(a[83]), .Z(n33186) );
  NANDN U33605 ( .A(n33186), .B(n38422), .Z(n33074) );
  NANDN U33606 ( .A(n33072), .B(n38423), .Z(n33073) );
  AND U33607 ( .A(n33074), .B(n33073), .Z(n33262) );
  XNOR U33608 ( .A(n33261), .B(n33262), .Z(n33263) );
  XNOR U33609 ( .A(n33264), .B(n33263), .Z(n33313) );
  XNOR U33610 ( .A(a[113]), .B(b[33]), .Z(n33237) );
  NANDN U33611 ( .A(n33237), .B(n35620), .Z(n33077) );
  NANDN U33612 ( .A(n33075), .B(n35621), .Z(n33076) );
  NAND U33613 ( .A(n33077), .B(n33076), .Z(n33234) );
  XNOR U33614 ( .A(b[55]), .B(a[91]), .Z(n33240) );
  NANDN U33615 ( .A(n33240), .B(n38075), .Z(n33080) );
  NANDN U33616 ( .A(n33078), .B(n38073), .Z(n33079) );
  NAND U33617 ( .A(n33080), .B(n33079), .Z(n33231) );
  NAND U33618 ( .A(n38326), .B(n33081), .Z(n33083) );
  XNOR U33619 ( .A(n38400), .B(a[87]), .Z(n33225) );
  NANDN U33620 ( .A(n38273), .B(n33225), .Z(n33082) );
  AND U33621 ( .A(n33083), .B(n33082), .Z(n33232) );
  XNOR U33622 ( .A(n33231), .B(n33232), .Z(n33233) );
  XOR U33623 ( .A(n33234), .B(n33233), .Z(n33314) );
  XNOR U33624 ( .A(n33313), .B(n33314), .Z(n33315) );
  XNOR U33625 ( .A(n33316), .B(n33315), .Z(n33301) );
  XOR U33626 ( .A(n33302), .B(n33301), .Z(n33304) );
  XNOR U33627 ( .A(n33303), .B(n33304), .Z(n33198) );
  XNOR U33628 ( .A(n33197), .B(n33198), .Z(n33140) );
  NANDN U33629 ( .A(n33085), .B(n33084), .Z(n33089) );
  OR U33630 ( .A(n33087), .B(n33086), .Z(n33088) );
  AND U33631 ( .A(n33089), .B(n33088), .Z(n33141) );
  NANDN U33632 ( .A(n33091), .B(n33090), .Z(n33095) );
  NAND U33633 ( .A(n33093), .B(n33092), .Z(n33094) );
  NAND U33634 ( .A(n33095), .B(n33094), .Z(n33142) );
  XOR U33635 ( .A(n33143), .B(n33142), .Z(n33334) );
  NANDN U33636 ( .A(n33097), .B(n33096), .Z(n33101) );
  NANDN U33637 ( .A(n33099), .B(n33098), .Z(n33100) );
  NAND U33638 ( .A(n33101), .B(n33100), .Z(n33332) );
  NANDN U33639 ( .A(n33103), .B(n33102), .Z(n33107) );
  NAND U33640 ( .A(n33105), .B(n33104), .Z(n33106) );
  AND U33641 ( .A(n33107), .B(n33106), .Z(n33331) );
  XNOR U33642 ( .A(n33332), .B(n33331), .Z(n33333) );
  XOR U33643 ( .A(n33334), .B(n33333), .Z(n33137) );
  XNOR U33644 ( .A(n33136), .B(n33137), .Z(n33122) );
  XNOR U33645 ( .A(n33123), .B(n33122), .Z(n33125) );
  XNOR U33646 ( .A(n33124), .B(n33125), .Z(n33116) );
  NANDN U33647 ( .A(n33109), .B(n33108), .Z(n33113) );
  NAND U33648 ( .A(n33111), .B(n33110), .Z(n33112) );
  AND U33649 ( .A(n33113), .B(n33112), .Z(n33117) );
  XNOR U33650 ( .A(n33116), .B(n33117), .Z(n33119) );
  XNOR U33651 ( .A(n33118), .B(n33119), .Z(n33337) );
  OR U33652 ( .A(n33115), .B(n33114), .Z(n33338) );
  XNOR U33653 ( .A(n33337), .B(n33338), .Z(c[209]) );
  NAND U33654 ( .A(n33117), .B(n33116), .Z(n33121) );
  NANDN U33655 ( .A(n33119), .B(n33118), .Z(n33120) );
  NAND U33656 ( .A(n33121), .B(n33120), .Z(n33342) );
  NAND U33657 ( .A(n33123), .B(n33122), .Z(n33127) );
  NANDN U33658 ( .A(n33125), .B(n33124), .Z(n33126) );
  NAND U33659 ( .A(n33127), .B(n33126), .Z(n33339) );
  OR U33660 ( .A(n33129), .B(n33128), .Z(n33133) );
  NAND U33661 ( .A(n33131), .B(n33130), .Z(n33132) );
  NAND U33662 ( .A(n33133), .B(n33132), .Z(n33346) );
  NANDN U33663 ( .A(n33135), .B(n33134), .Z(n33139) );
  NANDN U33664 ( .A(n33137), .B(n33136), .Z(n33138) );
  AND U33665 ( .A(n33139), .B(n33138), .Z(n33345) );
  XNOR U33666 ( .A(n33346), .B(n33345), .Z(n33347) );
  OR U33667 ( .A(n33141), .B(n33140), .Z(n33145) );
  OR U33668 ( .A(n33143), .B(n33142), .Z(n33144) );
  NAND U33669 ( .A(n33145), .B(n33144), .Z(n33360) );
  OR U33670 ( .A(n33147), .B(n33146), .Z(n33151) );
  OR U33671 ( .A(n33149), .B(n33148), .Z(n33150) );
  AND U33672 ( .A(n33151), .B(n33150), .Z(n33391) );
  NANDN U33673 ( .A(n33153), .B(n33152), .Z(n33157) );
  OR U33674 ( .A(n33155), .B(n33154), .Z(n33156) );
  AND U33675 ( .A(n33157), .B(n33156), .Z(n33392) );
  XOR U33676 ( .A(n33391), .B(n33392), .Z(n33393) );
  XOR U33677 ( .A(b[43]), .B(n36647), .Z(n33443) );
  NANDN U33678 ( .A(n33443), .B(n37068), .Z(n33160) );
  NANDN U33679 ( .A(n33158), .B(n37069), .Z(n33159) );
  NAND U33680 ( .A(n33160), .B(n33159), .Z(n33428) );
  XNOR U33681 ( .A(n38251), .B(b[25]), .Z(n33513) );
  NANDN U33682 ( .A(n34219), .B(n33513), .Z(n33163) );
  NAND U33683 ( .A(n34217), .B(n33161), .Z(n33162) );
  NAND U33684 ( .A(n33163), .B(n33162), .Z(n33425) );
  NAND U33685 ( .A(n34044), .B(n33164), .Z(n33166) );
  XNOR U33686 ( .A(n38321), .B(b[23]), .Z(n33510) );
  NANDN U33687 ( .A(n33867), .B(n33510), .Z(n33165) );
  AND U33688 ( .A(n33166), .B(n33165), .Z(n33426) );
  XNOR U33689 ( .A(n33425), .B(n33426), .Z(n33427) );
  XNOR U33690 ( .A(n33428), .B(n33427), .Z(n33394) );
  XNOR U33691 ( .A(n33393), .B(n33394), .Z(n33409) );
  NANDN U33692 ( .A(n33168), .B(n33167), .Z(n33172) );
  NAND U33693 ( .A(n33170), .B(n33169), .Z(n33171) );
  NAND U33694 ( .A(n33172), .B(n33171), .Z(n33408) );
  NANDN U33695 ( .A(n33174), .B(n33173), .Z(n33178) );
  NAND U33696 ( .A(n33176), .B(n33175), .Z(n33177) );
  NAND U33697 ( .A(n33178), .B(n33177), .Z(n33542) );
  XNOR U33698 ( .A(b[45]), .B(a[102]), .Z(n33478) );
  NANDN U33699 ( .A(n33478), .B(n37261), .Z(n33181) );
  NAND U33700 ( .A(n33179), .B(n37262), .Z(n33180) );
  NAND U33701 ( .A(n33181), .B(n33180), .Z(n33422) );
  XOR U33702 ( .A(b[61]), .B(n33628), .Z(n33522) );
  OR U33703 ( .A(n33522), .B(n38371), .Z(n33184) );
  NANDN U33704 ( .A(n33182), .B(n38369), .Z(n33183) );
  NAND U33705 ( .A(n33184), .B(n33183), .Z(n33419) );
  XOR U33706 ( .A(b[63]), .B(n33185), .Z(n33440) );
  NANDN U33707 ( .A(n33440), .B(n38422), .Z(n33188) );
  NANDN U33708 ( .A(n33186), .B(n38423), .Z(n33187) );
  AND U33709 ( .A(n33188), .B(n33187), .Z(n33420) );
  XNOR U33710 ( .A(n33419), .B(n33420), .Z(n33421) );
  XNOR U33711 ( .A(n33422), .B(n33421), .Z(n33540) );
  NANDN U33712 ( .A(n33190), .B(n33189), .Z(n33194) );
  NAND U33713 ( .A(n33192), .B(n33191), .Z(n33193) );
  NAND U33714 ( .A(n33194), .B(n33193), .Z(n33541) );
  XOR U33715 ( .A(n33540), .B(n33541), .Z(n33543) );
  XOR U33716 ( .A(n33542), .B(n33543), .Z(n33407) );
  XOR U33717 ( .A(n33408), .B(n33407), .Z(n33410) );
  XOR U33718 ( .A(n33409), .B(n33410), .Z(n33369) );
  NANDN U33719 ( .A(n33196), .B(n33195), .Z(n33200) );
  NAND U33720 ( .A(n33198), .B(n33197), .Z(n33199) );
  NAND U33721 ( .A(n33200), .B(n33199), .Z(n33370) );
  XOR U33722 ( .A(n33369), .B(n33370), .Z(n33371) );
  NANDN U33723 ( .A(n33202), .B(n33201), .Z(n33206) );
  NAND U33724 ( .A(n33204), .B(n33203), .Z(n33205) );
  AND U33725 ( .A(n33206), .B(n33205), .Z(n33372) );
  XNOR U33726 ( .A(n33371), .B(n33372), .Z(n33354) );
  NANDN U33727 ( .A(n33208), .B(n33207), .Z(n33212) );
  NAND U33728 ( .A(n33210), .B(n33209), .Z(n33211) );
  NAND U33729 ( .A(n33212), .B(n33211), .Z(n33384) );
  XNOR U33730 ( .A(a[112]), .B(b[35]), .Z(n33484) );
  NANDN U33731 ( .A(n33484), .B(n35985), .Z(n33215) );
  NAND U33732 ( .A(n33213), .B(n35986), .Z(n33214) );
  NAND U33733 ( .A(n33215), .B(n33214), .Z(n33507) );
  NAND U33734 ( .A(n37469), .B(n33216), .Z(n33218) );
  XOR U33735 ( .A(n978), .B(n36100), .Z(n33434) );
  NAND U33736 ( .A(n33434), .B(n37471), .Z(n33217) );
  NAND U33737 ( .A(n33218), .B(n33217), .Z(n33504) );
  XOR U33738 ( .A(b[53]), .B(n35191), .Z(n33437) );
  NANDN U33739 ( .A(n33437), .B(n37940), .Z(n33221) );
  NANDN U33740 ( .A(n33219), .B(n37941), .Z(n33220) );
  AND U33741 ( .A(n33221), .B(n33220), .Z(n33505) );
  XNOR U33742 ( .A(n33504), .B(n33505), .Z(n33506) );
  XOR U33743 ( .A(n33507), .B(n33506), .Z(n33397) );
  XOR U33744 ( .A(b[49]), .B(n35783), .Z(n33516) );
  OR U33745 ( .A(n33516), .B(n37756), .Z(n33224) );
  NANDN U33746 ( .A(n33222), .B(n37652), .Z(n33223) );
  NAND U33747 ( .A(n33224), .B(n33223), .Z(n33501) );
  NAND U33748 ( .A(n38326), .B(n33225), .Z(n33227) );
  XOR U33749 ( .A(n38400), .B(n34048), .Z(n33519) );
  NANDN U33750 ( .A(n38273), .B(n33519), .Z(n33226) );
  NAND U33751 ( .A(n33227), .B(n33226), .Z(n33498) );
  NAND U33752 ( .A(n34848), .B(n33228), .Z(n33230) );
  XOR U33753 ( .A(n38134), .B(n35375), .Z(n33461) );
  NAND U33754 ( .A(n34618), .B(n33461), .Z(n33229) );
  AND U33755 ( .A(n33230), .B(n33229), .Z(n33499) );
  XNOR U33756 ( .A(n33498), .B(n33499), .Z(n33500) );
  XOR U33757 ( .A(n33501), .B(n33500), .Z(n33398) );
  XNOR U33758 ( .A(n33397), .B(n33398), .Z(n33400) );
  NANDN U33759 ( .A(n33232), .B(n33231), .Z(n33236) );
  NAND U33760 ( .A(n33234), .B(n33233), .Z(n33235) );
  NAND U33761 ( .A(n33236), .B(n33235), .Z(n33399) );
  XOR U33762 ( .A(n33400), .B(n33399), .Z(n33403) );
  XOR U33763 ( .A(a[114]), .B(n974), .Z(n33481) );
  NANDN U33764 ( .A(n33481), .B(n35620), .Z(n33239) );
  NANDN U33765 ( .A(n33237), .B(n35621), .Z(n33238) );
  NAND U33766 ( .A(n33239), .B(n33238), .Z(n33452) );
  XOR U33767 ( .A(b[55]), .B(n34852), .Z(n33458) );
  NANDN U33768 ( .A(n33458), .B(n38075), .Z(n33242) );
  NANDN U33769 ( .A(n33240), .B(n38073), .Z(n33241) );
  NAND U33770 ( .A(n33242), .B(n33241), .Z(n33449) );
  XOR U33771 ( .A(b[57]), .B(n34851), .Z(n33455) );
  OR U33772 ( .A(n33455), .B(n965), .Z(n33245) );
  NANDN U33773 ( .A(n33243), .B(n38194), .Z(n33244) );
  AND U33774 ( .A(n33245), .B(n33244), .Z(n33450) );
  XNOR U33775 ( .A(n33449), .B(n33450), .Z(n33451) );
  XOR U33776 ( .A(n33452), .B(n33451), .Z(n33387) );
  XOR U33777 ( .A(a[116]), .B(n973), .Z(n33472) );
  NANDN U33778 ( .A(n33472), .B(n35313), .Z(n33248) );
  NANDN U33779 ( .A(n33246), .B(n35311), .Z(n33247) );
  NAND U33780 ( .A(n33248), .B(n33247), .Z(n33531) );
  NAND U33781 ( .A(n35188), .B(n33249), .Z(n33251) );
  XOR U33782 ( .A(n38143), .B(n35540), .Z(n33431) );
  NANDN U33783 ( .A(n34968), .B(n33431), .Z(n33250) );
  NAND U33784 ( .A(n33251), .B(n33250), .Z(n33528) );
  XOR U33785 ( .A(b[51]), .B(n35545), .Z(n33525) );
  NANDN U33786 ( .A(n33525), .B(n37803), .Z(n33254) );
  NANDN U33787 ( .A(n33252), .B(n37802), .Z(n33253) );
  AND U33788 ( .A(n33254), .B(n33253), .Z(n33529) );
  XNOR U33789 ( .A(n33528), .B(n33529), .Z(n33530) );
  XOR U33790 ( .A(n33531), .B(n33530), .Z(n33385) );
  NANDN U33791 ( .A(n33256), .B(n33255), .Z(n33260) );
  NAND U33792 ( .A(n33258), .B(n33257), .Z(n33259) );
  NAND U33793 ( .A(n33260), .B(n33259), .Z(n33386) );
  XNOR U33794 ( .A(n33385), .B(n33386), .Z(n33388) );
  XNOR U33795 ( .A(n33387), .B(n33388), .Z(n33404) );
  XNOR U33796 ( .A(n33403), .B(n33404), .Z(n33405) );
  NANDN U33797 ( .A(n33262), .B(n33261), .Z(n33266) );
  NAND U33798 ( .A(n33264), .B(n33263), .Z(n33265) );
  NAND U33799 ( .A(n33266), .B(n33265), .Z(n33416) );
  XOR U33800 ( .A(a[110]), .B(n975), .Z(n33475) );
  NANDN U33801 ( .A(n33475), .B(n36311), .Z(n33269) );
  NAND U33802 ( .A(n33267), .B(n36309), .Z(n33268) );
  NAND U33803 ( .A(n33269), .B(n33268), .Z(n33495) );
  XOR U33804 ( .A(a[108]), .B(n976), .Z(n33469) );
  NANDN U33805 ( .A(n33469), .B(n36553), .Z(n33272) );
  NAND U33806 ( .A(n33270), .B(n36643), .Z(n33271) );
  NAND U33807 ( .A(n33272), .B(n33271), .Z(n33492) );
  XNOR U33808 ( .A(b[41]), .B(a[106]), .Z(n33446) );
  OR U33809 ( .A(n33446), .B(n36905), .Z(n33275) );
  NAND U33810 ( .A(n33273), .B(n36807), .Z(n33274) );
  AND U33811 ( .A(n33275), .B(n33274), .Z(n33493) );
  XNOR U33812 ( .A(n33492), .B(n33493), .Z(n33494) );
  XOR U33813 ( .A(n33495), .B(n33494), .Z(n33534) );
  NANDN U33814 ( .A(n33277), .B(n33276), .Z(n33281) );
  NAND U33815 ( .A(n33279), .B(n33278), .Z(n33280) );
  NAND U33816 ( .A(n33281), .B(n33280), .Z(n33535) );
  XNOR U33817 ( .A(n33534), .B(n33535), .Z(n33537) );
  NAND U33818 ( .A(n33283), .B(n33282), .Z(n33285) );
  ANDN U33819 ( .B(n33285), .A(n33284), .Z(n33489) );
  AND U33820 ( .A(a[82]), .B(b[63]), .Z(n33609) );
  XNOR U33821 ( .A(a[126]), .B(b[21]), .Z(n33465) );
  OR U33822 ( .A(n33465), .B(n33634), .Z(n33288) );
  NAND U33823 ( .A(n33286), .B(n33464), .Z(n33287) );
  NAND U33824 ( .A(n33288), .B(n33287), .Z(n33487) );
  XNOR U33825 ( .A(n33609), .B(n33487), .Z(n33488) );
  XNOR U33826 ( .A(n33489), .B(n33488), .Z(n33536) );
  XNOR U33827 ( .A(n33537), .B(n33536), .Z(n33414) );
  NANDN U33828 ( .A(n33290), .B(n33289), .Z(n33294) );
  NAND U33829 ( .A(n33292), .B(n33291), .Z(n33293) );
  AND U33830 ( .A(n33294), .B(n33293), .Z(n33413) );
  XNOR U33831 ( .A(n33414), .B(n33413), .Z(n33415) );
  XOR U33832 ( .A(n33416), .B(n33415), .Z(n33406) );
  XOR U33833 ( .A(n33405), .B(n33406), .Z(n33381) );
  NANDN U33834 ( .A(n33296), .B(n33295), .Z(n33300) );
  NAND U33835 ( .A(n33298), .B(n33297), .Z(n33299) );
  NAND U33836 ( .A(n33300), .B(n33299), .Z(n33382) );
  XNOR U33837 ( .A(n33381), .B(n33382), .Z(n33383) );
  XOR U33838 ( .A(n33384), .B(n33383), .Z(n33377) );
  NANDN U33839 ( .A(n33302), .B(n33301), .Z(n33306) );
  NANDN U33840 ( .A(n33304), .B(n33303), .Z(n33305) );
  NAND U33841 ( .A(n33306), .B(n33305), .Z(n33376) );
  OR U33842 ( .A(n33308), .B(n33307), .Z(n33312) );
  NANDN U33843 ( .A(n33310), .B(n33309), .Z(n33311) );
  NAND U33844 ( .A(n33312), .B(n33311), .Z(n33364) );
  NANDN U33845 ( .A(n33314), .B(n33313), .Z(n33318) );
  NANDN U33846 ( .A(n33316), .B(n33315), .Z(n33317) );
  AND U33847 ( .A(n33318), .B(n33317), .Z(n33363) );
  XNOR U33848 ( .A(n33364), .B(n33363), .Z(n33365) );
  OR U33849 ( .A(n33320), .B(n33319), .Z(n33324) );
  NANDN U33850 ( .A(n33322), .B(n33321), .Z(n33323) );
  NAND U33851 ( .A(n33324), .B(n33323), .Z(n33366) );
  XOR U33852 ( .A(n33365), .B(n33366), .Z(n33375) );
  XNOR U33853 ( .A(n33376), .B(n33375), .Z(n33378) );
  XNOR U33854 ( .A(n33377), .B(n33378), .Z(n33351) );
  NANDN U33855 ( .A(n33326), .B(n33325), .Z(n33330) );
  NANDN U33856 ( .A(n33328), .B(n33327), .Z(n33329) );
  NAND U33857 ( .A(n33330), .B(n33329), .Z(n33352) );
  XNOR U33858 ( .A(n33351), .B(n33352), .Z(n33353) );
  XNOR U33859 ( .A(n33354), .B(n33353), .Z(n33357) );
  NANDN U33860 ( .A(n33332), .B(n33331), .Z(n33336) );
  NANDN U33861 ( .A(n33334), .B(n33333), .Z(n33335) );
  NAND U33862 ( .A(n33336), .B(n33335), .Z(n33358) );
  XNOR U33863 ( .A(n33357), .B(n33358), .Z(n33359) );
  XNOR U33864 ( .A(n33360), .B(n33359), .Z(n33348) );
  XNOR U33865 ( .A(n33347), .B(n33348), .Z(n33340) );
  XNOR U33866 ( .A(n33339), .B(n33340), .Z(n33341) );
  XNOR U33867 ( .A(n33342), .B(n33341), .Z(n33547) );
  NANDN U33868 ( .A(n33338), .B(n33337), .Z(n33546) );
  XOR U33869 ( .A(n33547), .B(n33546), .Z(c[210]) );
  NANDN U33870 ( .A(n33340), .B(n33339), .Z(n33344) );
  NAND U33871 ( .A(n33342), .B(n33341), .Z(n33343) );
  NAND U33872 ( .A(n33344), .B(n33343), .Z(n33553) );
  NANDN U33873 ( .A(n33346), .B(n33345), .Z(n33350) );
  NANDN U33874 ( .A(n33348), .B(n33347), .Z(n33349) );
  NAND U33875 ( .A(n33350), .B(n33349), .Z(n33551) );
  OR U33876 ( .A(n33352), .B(n33351), .Z(n33356) );
  OR U33877 ( .A(n33354), .B(n33353), .Z(n33355) );
  NAND U33878 ( .A(n33356), .B(n33355), .Z(n33755) );
  NANDN U33879 ( .A(n33358), .B(n33357), .Z(n33362) );
  NAND U33880 ( .A(n33360), .B(n33359), .Z(n33361) );
  NAND U33881 ( .A(n33362), .B(n33361), .Z(n33756) );
  XNOR U33882 ( .A(n33755), .B(n33756), .Z(n33757) );
  OR U33883 ( .A(n33364), .B(n33363), .Z(n33368) );
  OR U33884 ( .A(n33366), .B(n33365), .Z(n33367) );
  NAND U33885 ( .A(n33368), .B(n33367), .Z(n33753) );
  OR U33886 ( .A(n33370), .B(n33369), .Z(n33374) );
  NAND U33887 ( .A(n33372), .B(n33371), .Z(n33373) );
  NAND U33888 ( .A(n33374), .B(n33373), .Z(n33752) );
  NAND U33889 ( .A(n33376), .B(n33375), .Z(n33380) );
  NANDN U33890 ( .A(n33378), .B(n33377), .Z(n33379) );
  NAND U33891 ( .A(n33380), .B(n33379), .Z(n33748) );
  OR U33892 ( .A(n33386), .B(n33385), .Z(n33390) );
  OR U33893 ( .A(n33388), .B(n33387), .Z(n33389) );
  AND U33894 ( .A(n33390), .B(n33389), .Z(n33568) );
  OR U33895 ( .A(n33392), .B(n33391), .Z(n33396) );
  NANDN U33896 ( .A(n33394), .B(n33393), .Z(n33395) );
  NAND U33897 ( .A(n33396), .B(n33395), .Z(n33569) );
  XOR U33898 ( .A(n33568), .B(n33569), .Z(n33570) );
  OR U33899 ( .A(n33398), .B(n33397), .Z(n33402) );
  OR U33900 ( .A(n33400), .B(n33399), .Z(n33401) );
  AND U33901 ( .A(n33402), .B(n33401), .Z(n33571) );
  XNOR U33902 ( .A(n33570), .B(n33571), .Z(n33562) );
  XOR U33903 ( .A(n33562), .B(n33563), .Z(n33564) );
  XNOR U33904 ( .A(n33565), .B(n33564), .Z(n33746) );
  NANDN U33905 ( .A(n33408), .B(n33407), .Z(n33412) );
  OR U33906 ( .A(n33410), .B(n33409), .Z(n33411) );
  NAND U33907 ( .A(n33412), .B(n33411), .Z(n33741) );
  NANDN U33908 ( .A(n33414), .B(n33413), .Z(n33418) );
  NANDN U33909 ( .A(n33416), .B(n33415), .Z(n33417) );
  NAND U33910 ( .A(n33418), .B(n33417), .Z(n33736) );
  NANDN U33911 ( .A(n33420), .B(n33419), .Z(n33424) );
  NAND U33912 ( .A(n33422), .B(n33421), .Z(n33423) );
  AND U33913 ( .A(n33424), .B(n33423), .Z(n33577) );
  NANDN U33914 ( .A(n33426), .B(n33425), .Z(n33430) );
  NAND U33915 ( .A(n33428), .B(n33427), .Z(n33429) );
  NAND U33916 ( .A(n33430), .B(n33429), .Z(n33588) );
  NAND U33917 ( .A(n35188), .B(n33431), .Z(n33433) );
  XNOR U33918 ( .A(n38193), .B(b[29]), .Z(n33676) );
  NANDN U33919 ( .A(n34968), .B(n33676), .Z(n33432) );
  NAND U33920 ( .A(n33433), .B(n33432), .Z(n33595) );
  NAND U33921 ( .A(n37469), .B(n33434), .Z(n33436) );
  XNOR U33922 ( .A(n978), .B(a[101]), .Z(n33667) );
  NAND U33923 ( .A(n33667), .B(n37471), .Z(n33435) );
  NAND U33924 ( .A(n33436), .B(n33435), .Z(n33592) );
  XOR U33925 ( .A(b[53]), .B(n35628), .Z(n33601) );
  NANDN U33926 ( .A(n33601), .B(n37940), .Z(n33439) );
  NANDN U33927 ( .A(n33437), .B(n37941), .Z(n33438) );
  AND U33928 ( .A(n33439), .B(n33438), .Z(n33593) );
  XNOR U33929 ( .A(n33592), .B(n33593), .Z(n33594) );
  XNOR U33930 ( .A(n33595), .B(n33594), .Z(n33586) );
  XNOR U33931 ( .A(b[63]), .B(a[85]), .Z(n33629) );
  NANDN U33932 ( .A(n33629), .B(n38422), .Z(n33442) );
  NANDN U33933 ( .A(n33440), .B(n38423), .Z(n33441) );
  NAND U33934 ( .A(n33442), .B(n33441), .Z(n33637) );
  XNOR U33935 ( .A(b[43]), .B(a[105]), .Z(n33709) );
  NANDN U33936 ( .A(n33709), .B(n37068), .Z(n33445) );
  NANDN U33937 ( .A(n33443), .B(n37069), .Z(n33444) );
  AND U33938 ( .A(n33445), .B(n33444), .Z(n33638) );
  XNOR U33939 ( .A(n33637), .B(n33638), .Z(n33639) );
  XOR U33940 ( .A(b[41]), .B(a[107]), .Z(n33625) );
  NANDN U33941 ( .A(n36905), .B(n33625), .Z(n33448) );
  NANDN U33942 ( .A(n33446), .B(n36807), .Z(n33447) );
  NAND U33943 ( .A(n33448), .B(n33447), .Z(n33607) );
  NANDN U33944 ( .A(n985), .B(a[83]), .Z(n33608) );
  XNOR U33945 ( .A(n33607), .B(n33608), .Z(n33610) );
  XNOR U33946 ( .A(n33609), .B(n33610), .Z(n33640) );
  XNOR U33947 ( .A(n33639), .B(n33640), .Z(n33587) );
  XOR U33948 ( .A(n33586), .B(n33587), .Z(n33589) );
  XNOR U33949 ( .A(n33588), .B(n33589), .Z(n33574) );
  NANDN U33950 ( .A(n33450), .B(n33449), .Z(n33454) );
  NAND U33951 ( .A(n33452), .B(n33451), .Z(n33453) );
  AND U33952 ( .A(n33454), .B(n33453), .Z(n33575) );
  XNOR U33953 ( .A(n33574), .B(n33575), .Z(n33576) );
  XNOR U33954 ( .A(n33577), .B(n33576), .Z(n33734) );
  XNOR U33955 ( .A(b[57]), .B(a[91]), .Z(n33724) );
  OR U33956 ( .A(n33724), .B(n965), .Z(n33457) );
  NANDN U33957 ( .A(n33455), .B(n38194), .Z(n33456) );
  NAND U33958 ( .A(n33457), .B(n33456), .Z(n33664) );
  XOR U33959 ( .A(b[55]), .B(n35377), .Z(n33604) );
  NANDN U33960 ( .A(n33604), .B(n38075), .Z(n33460) );
  NANDN U33961 ( .A(n33458), .B(n38073), .Z(n33459) );
  NAND U33962 ( .A(n33460), .B(n33459), .Z(n33661) );
  NAND U33963 ( .A(n34848), .B(n33461), .Z(n33463) );
  XNOR U33964 ( .A(a[121]), .B(b[27]), .Z(n33670) );
  NANDN U33965 ( .A(n33670), .B(n34618), .Z(n33462) );
  AND U33966 ( .A(n33463), .B(n33462), .Z(n33662) );
  XNOR U33967 ( .A(n33661), .B(n33662), .Z(n33663) );
  XNOR U33968 ( .A(n33664), .B(n33663), .Z(n33643) );
  XNOR U33969 ( .A(a[127]), .B(b[21]), .Z(n33633) );
  OR U33970 ( .A(n33633), .B(n33634), .Z(n33467) );
  NANDN U33971 ( .A(n33465), .B(n33464), .Z(n33466) );
  NAND U33972 ( .A(n33467), .B(n33466), .Z(n33700) );
  NAND U33973 ( .A(b[18]), .B(b[17]), .Z(n33468) );
  AND U33974 ( .A(n33468), .B(b[19]), .Z(n33697) );
  XNOR U33975 ( .A(a[109]), .B(n976), .Z(n33622) );
  NAND U33976 ( .A(n33622), .B(n36553), .Z(n33471) );
  NANDN U33977 ( .A(n33469), .B(n36643), .Z(n33470) );
  AND U33978 ( .A(n33471), .B(n33470), .Z(n33698) );
  XOR U33979 ( .A(n33697), .B(n33698), .Z(n33699) );
  XOR U33980 ( .A(n33700), .B(n33699), .Z(n33644) );
  XOR U33981 ( .A(n33643), .B(n33644), .Z(n33646) );
  XNOR U33982 ( .A(a[117]), .B(b[31]), .Z(n33721) );
  NANDN U33983 ( .A(n33721), .B(n35313), .Z(n33474) );
  NANDN U33984 ( .A(n33472), .B(n35311), .Z(n33473) );
  NAND U33985 ( .A(n33474), .B(n33473), .Z(n33730) );
  XNOR U33986 ( .A(a[111]), .B(b[37]), .Z(n33613) );
  NANDN U33987 ( .A(n33613), .B(n36311), .Z(n33477) );
  NANDN U33988 ( .A(n33475), .B(n36309), .Z(n33476) );
  NAND U33989 ( .A(n33477), .B(n33476), .Z(n33727) );
  XOR U33990 ( .A(b[45]), .B(a[103]), .Z(n33616) );
  NAND U33991 ( .A(n33616), .B(n37261), .Z(n33480) );
  NANDN U33992 ( .A(n33478), .B(n37262), .Z(n33479) );
  AND U33993 ( .A(n33480), .B(n33479), .Z(n33728) );
  XNOR U33994 ( .A(n33727), .B(n33728), .Z(n33729) );
  XNOR U33995 ( .A(n33730), .B(n33729), .Z(n33651) );
  XNOR U33996 ( .A(a[115]), .B(n974), .Z(n33718) );
  NAND U33997 ( .A(n35620), .B(n33718), .Z(n33483) );
  NANDN U33998 ( .A(n33481), .B(n35621), .Z(n33482) );
  NAND U33999 ( .A(n33483), .B(n33482), .Z(n33650) );
  NANDN U34000 ( .A(n33484), .B(n35986), .Z(n33486) );
  XOR U34001 ( .A(a[113]), .B(b[35]), .Z(n33598) );
  NAND U34002 ( .A(n35985), .B(n33598), .Z(n33485) );
  NAND U34003 ( .A(n33486), .B(n33485), .Z(n33649) );
  XOR U34004 ( .A(n33646), .B(n33645), .Z(n33694) );
  NANDN U34005 ( .A(n33609), .B(n33487), .Z(n33491) );
  NANDN U34006 ( .A(n33489), .B(n33488), .Z(n33490) );
  NAND U34007 ( .A(n33491), .B(n33490), .Z(n33691) );
  NANDN U34008 ( .A(n33493), .B(n33492), .Z(n33497) );
  NAND U34009 ( .A(n33495), .B(n33494), .Z(n33496) );
  AND U34010 ( .A(n33497), .B(n33496), .Z(n33692) );
  XNOR U34011 ( .A(n33691), .B(n33692), .Z(n33693) );
  XOR U34012 ( .A(n33694), .B(n33693), .Z(n33733) );
  XOR U34013 ( .A(n33734), .B(n33733), .Z(n33735) );
  XNOR U34014 ( .A(n33736), .B(n33735), .Z(n33739) );
  NANDN U34015 ( .A(n33499), .B(n33498), .Z(n33503) );
  NAND U34016 ( .A(n33501), .B(n33500), .Z(n33502) );
  NAND U34017 ( .A(n33503), .B(n33502), .Z(n33688) );
  NANDN U34018 ( .A(n33505), .B(n33504), .Z(n33509) );
  NAND U34019 ( .A(n33507), .B(n33506), .Z(n33508) );
  NAND U34020 ( .A(n33509), .B(n33508), .Z(n33583) );
  NAND U34021 ( .A(n33510), .B(n34044), .Z(n33512) );
  XNOR U34022 ( .A(a[125]), .B(n34510), .Z(n33712) );
  NANDN U34023 ( .A(n33867), .B(n33712), .Z(n33511) );
  AND U34024 ( .A(n33512), .B(n33511), .Z(n33655) );
  XOR U34025 ( .A(a[123]), .B(b[25]), .Z(n33673) );
  NANDN U34026 ( .A(n34219), .B(n33673), .Z(n33515) );
  NAND U34027 ( .A(n33513), .B(n34217), .Z(n33514) );
  AND U34028 ( .A(n33515), .B(n33514), .Z(n33656) );
  XOR U34029 ( .A(n33655), .B(n33656), .Z(n33657) );
  XNOR U34030 ( .A(n979), .B(a[99]), .Z(n33682) );
  NANDN U34031 ( .A(n37756), .B(n33682), .Z(n33518) );
  NANDN U34032 ( .A(n33516), .B(n37652), .Z(n33517) );
  AND U34033 ( .A(n33518), .B(n33517), .Z(n33658) );
  XNOR U34034 ( .A(n33657), .B(n33658), .Z(n33581) );
  NAND U34035 ( .A(n38326), .B(n33519), .Z(n33521) );
  XNOR U34036 ( .A(n38400), .B(a[89]), .Z(n33679) );
  NANDN U34037 ( .A(n38273), .B(n33679), .Z(n33520) );
  NAND U34038 ( .A(n33521), .B(n33520), .Z(n33706) );
  XNOR U34039 ( .A(b[61]), .B(a[87]), .Z(n33715) );
  OR U34040 ( .A(n33715), .B(n38371), .Z(n33524) );
  NANDN U34041 ( .A(n33522), .B(n38369), .Z(n33523) );
  NAND U34042 ( .A(n33524), .B(n33523), .Z(n33703) );
  XNOR U34043 ( .A(b[51]), .B(a[97]), .Z(n33619) );
  NANDN U34044 ( .A(n33619), .B(n37803), .Z(n33527) );
  NANDN U34045 ( .A(n33525), .B(n37802), .Z(n33526) );
  AND U34046 ( .A(n33527), .B(n33526), .Z(n33704) );
  XNOR U34047 ( .A(n33703), .B(n33704), .Z(n33705) );
  XOR U34048 ( .A(n33706), .B(n33705), .Z(n33580) );
  XOR U34049 ( .A(n33581), .B(n33580), .Z(n33582) );
  XOR U34050 ( .A(n33583), .B(n33582), .Z(n33685) );
  NANDN U34051 ( .A(n33529), .B(n33528), .Z(n33533) );
  NAND U34052 ( .A(n33531), .B(n33530), .Z(n33532) );
  AND U34053 ( .A(n33533), .B(n33532), .Z(n33686) );
  XNOR U34054 ( .A(n33685), .B(n33686), .Z(n33687) );
  XOR U34055 ( .A(n33688), .B(n33687), .Z(n33556) );
  OR U34056 ( .A(n33535), .B(n33534), .Z(n33539) );
  OR U34057 ( .A(n33537), .B(n33536), .Z(n33538) );
  AND U34058 ( .A(n33539), .B(n33538), .Z(n33557) );
  XNOR U34059 ( .A(n33556), .B(n33557), .Z(n33559) );
  NANDN U34060 ( .A(n33541), .B(n33540), .Z(n33545) );
  OR U34061 ( .A(n33543), .B(n33542), .Z(n33544) );
  AND U34062 ( .A(n33545), .B(n33544), .Z(n33558) );
  XOR U34063 ( .A(n33559), .B(n33558), .Z(n33740) );
  XOR U34064 ( .A(n33739), .B(n33740), .Z(n33742) );
  XOR U34065 ( .A(n33741), .B(n33742), .Z(n33745) );
  XNOR U34066 ( .A(n33746), .B(n33745), .Z(n33747) );
  XNOR U34067 ( .A(n33748), .B(n33747), .Z(n33751) );
  XNOR U34068 ( .A(n33752), .B(n33751), .Z(n33754) );
  XOR U34069 ( .A(n33753), .B(n33754), .Z(n33758) );
  XOR U34070 ( .A(n33757), .B(n33758), .Z(n33550) );
  XNOR U34071 ( .A(n33551), .B(n33550), .Z(n33552) );
  XNOR U34072 ( .A(n33553), .B(n33552), .Z(n33549) );
  OR U34073 ( .A(n33547), .B(n33546), .Z(n33548) );
  XOR U34074 ( .A(n33549), .B(n33548), .Z(c[211]) );
  OR U34075 ( .A(n33549), .B(n33548), .Z(n33763) );
  NANDN U34076 ( .A(n33551), .B(n33550), .Z(n33555) );
  NAND U34077 ( .A(n33553), .B(n33552), .Z(n33554) );
  AND U34078 ( .A(n33555), .B(n33554), .Z(n33957) );
  OR U34079 ( .A(n33557), .B(n33556), .Z(n33561) );
  OR U34080 ( .A(n33559), .B(n33558), .Z(n33560) );
  NAND U34081 ( .A(n33561), .B(n33560), .Z(n33771) );
  OR U34082 ( .A(n33563), .B(n33562), .Z(n33567) );
  NAND U34083 ( .A(n33565), .B(n33564), .Z(n33566) );
  AND U34084 ( .A(n33567), .B(n33566), .Z(n33768) );
  OR U34085 ( .A(n33569), .B(n33568), .Z(n33573) );
  NANDN U34086 ( .A(n33571), .B(n33570), .Z(n33572) );
  NAND U34087 ( .A(n33573), .B(n33572), .Z(n33769) );
  XOR U34088 ( .A(n33768), .B(n33769), .Z(n33770) );
  XNOR U34089 ( .A(n33771), .B(n33770), .Z(n33777) );
  NANDN U34090 ( .A(n33575), .B(n33574), .Z(n33579) );
  NANDN U34091 ( .A(n33577), .B(n33576), .Z(n33578) );
  NAND U34092 ( .A(n33579), .B(n33578), .Z(n33950) );
  OR U34093 ( .A(n33581), .B(n33580), .Z(n33585) );
  NANDN U34094 ( .A(n33583), .B(n33582), .Z(n33584) );
  NAND U34095 ( .A(n33585), .B(n33584), .Z(n33827) );
  NANDN U34096 ( .A(n33587), .B(n33586), .Z(n33591) );
  OR U34097 ( .A(n33589), .B(n33588), .Z(n33590) );
  NAND U34098 ( .A(n33591), .B(n33590), .Z(n33825) );
  NANDN U34099 ( .A(n33593), .B(n33592), .Z(n33597) );
  NAND U34100 ( .A(n33595), .B(n33594), .Z(n33596) );
  NAND U34101 ( .A(n33597), .B(n33596), .Z(n33820) );
  XNOR U34102 ( .A(a[114]), .B(b[35]), .Z(n33928) );
  NANDN U34103 ( .A(n33928), .B(n35985), .Z(n33600) );
  NAND U34104 ( .A(n33598), .B(n35986), .Z(n33599) );
  NAND U34105 ( .A(n33600), .B(n33599), .Z(n33876) );
  XOR U34106 ( .A(b[53]), .B(n35545), .Z(n33922) );
  NANDN U34107 ( .A(n33922), .B(n37940), .Z(n33603) );
  NANDN U34108 ( .A(n33601), .B(n37941), .Z(n33602) );
  NAND U34109 ( .A(n33603), .B(n33602), .Z(n33873) );
  XOR U34110 ( .A(b[55]), .B(n35191), .Z(n33916) );
  NANDN U34111 ( .A(n33916), .B(n38075), .Z(n33606) );
  NANDN U34112 ( .A(n33604), .B(n38073), .Z(n33605) );
  AND U34113 ( .A(n33606), .B(n33605), .Z(n33874) );
  XNOR U34114 ( .A(n33873), .B(n33874), .Z(n33875) );
  XNOR U34115 ( .A(n33876), .B(n33875), .Z(n33818) );
  NANDN U34116 ( .A(n33608), .B(n33607), .Z(n33612) );
  NAND U34117 ( .A(n33610), .B(n33609), .Z(n33611) );
  NAND U34118 ( .A(n33612), .B(n33611), .Z(n33819) );
  XOR U34119 ( .A(n33818), .B(n33819), .Z(n33821) );
  XOR U34120 ( .A(n33820), .B(n33821), .Z(n33824) );
  XOR U34121 ( .A(n33825), .B(n33824), .Z(n33826) );
  XNOR U34122 ( .A(n33827), .B(n33826), .Z(n33949) );
  XNOR U34123 ( .A(n33950), .B(n33949), .Z(n33952) );
  XOR U34124 ( .A(a[112]), .B(n975), .Z(n33815) );
  NANDN U34125 ( .A(n33815), .B(n36311), .Z(n33615) );
  NANDN U34126 ( .A(n33613), .B(n36309), .Z(n33614) );
  NAND U34127 ( .A(n33615), .B(n33614), .Z(n33783) );
  XNOR U34128 ( .A(b[45]), .B(a[104]), .Z(n33863) );
  NANDN U34129 ( .A(n33863), .B(n37261), .Z(n33618) );
  NAND U34130 ( .A(n33616), .B(n37262), .Z(n33617) );
  NAND U34131 ( .A(n33618), .B(n33617), .Z(n33780) );
  XOR U34132 ( .A(b[51]), .B(n35783), .Z(n33803) );
  NANDN U34133 ( .A(n33803), .B(n37803), .Z(n33621) );
  NANDN U34134 ( .A(n33619), .B(n37802), .Z(n33620) );
  AND U34135 ( .A(n33621), .B(n33620), .Z(n33781) );
  XNOR U34136 ( .A(n33780), .B(n33781), .Z(n33782) );
  XNOR U34137 ( .A(n33783), .B(n33782), .Z(n33900) );
  NAND U34138 ( .A(n36643), .B(n33622), .Z(n33624) );
  XNOR U34139 ( .A(n37336), .B(b[39]), .Z(n33809) );
  NAND U34140 ( .A(n33809), .B(n36553), .Z(n33623) );
  NAND U34141 ( .A(n33624), .B(n33623), .Z(n33898) );
  NAND U34142 ( .A(n36807), .B(n33625), .Z(n33627) );
  XNOR U34143 ( .A(n37139), .B(b[41]), .Z(n33913) );
  NANDN U34144 ( .A(n36905), .B(n33913), .Z(n33626) );
  AND U34145 ( .A(n33627), .B(n33626), .Z(n33897) );
  XNOR U34146 ( .A(n33898), .B(n33897), .Z(n33899) );
  XOR U34147 ( .A(n33900), .B(n33899), .Z(n33893) );
  XOR U34148 ( .A(b[63]), .B(n33628), .Z(n33791) );
  NANDN U34149 ( .A(n33791), .B(n38422), .Z(n33631) );
  NANDN U34150 ( .A(n33629), .B(n38423), .Z(n33630) );
  NAND U34151 ( .A(n33631), .B(n33630), .Z(n33787) );
  XNOR U34152 ( .A(b[21]), .B(n33632), .Z(n33636) );
  NAND U34153 ( .A(n33634), .B(n33633), .Z(n33635) );
  AND U34154 ( .A(n33636), .B(n33635), .Z(n33786) );
  AND U34155 ( .A(b[63]), .B(a[84]), .Z(n33985) );
  XOR U34156 ( .A(n33786), .B(n33985), .Z(n33788) );
  XNOR U34157 ( .A(n33787), .B(n33788), .Z(n33891) );
  NANDN U34158 ( .A(n33638), .B(n33637), .Z(n33642) );
  NANDN U34159 ( .A(n33640), .B(n33639), .Z(n33641) );
  NAND U34160 ( .A(n33642), .B(n33641), .Z(n33892) );
  XOR U34161 ( .A(n33891), .B(n33892), .Z(n33894) );
  XOR U34162 ( .A(n33893), .B(n33894), .Z(n33832) );
  NANDN U34163 ( .A(n33644), .B(n33643), .Z(n33648) );
  NANDN U34164 ( .A(n33646), .B(n33645), .Z(n33647) );
  NAND U34165 ( .A(n33648), .B(n33647), .Z(n33830) );
  OR U34166 ( .A(n33650), .B(n33649), .Z(n33654) );
  NANDN U34167 ( .A(n33652), .B(n33651), .Z(n33653) );
  AND U34168 ( .A(n33654), .B(n33653), .Z(n33931) );
  OR U34169 ( .A(n33656), .B(n33655), .Z(n33660) );
  NANDN U34170 ( .A(n33658), .B(n33657), .Z(n33659) );
  NAND U34171 ( .A(n33660), .B(n33659), .Z(n33932) );
  XNOR U34172 ( .A(n33931), .B(n33932), .Z(n33933) );
  NANDN U34173 ( .A(n33662), .B(n33661), .Z(n33666) );
  NAND U34174 ( .A(n33664), .B(n33663), .Z(n33665) );
  NAND U34175 ( .A(n33666), .B(n33665), .Z(n33851) );
  NAND U34176 ( .A(n33667), .B(n37469), .Z(n33669) );
  XNOR U34177 ( .A(n978), .B(a[102]), .Z(n33860) );
  NAND U34178 ( .A(n33860), .B(n37471), .Z(n33668) );
  NAND U34179 ( .A(n33669), .B(n33668), .Z(n33911) );
  NANDN U34180 ( .A(n33670), .B(n34848), .Z(n33672) );
  XNOR U34181 ( .A(n38251), .B(b[27]), .Z(n33925) );
  NAND U34182 ( .A(n34618), .B(n33925), .Z(n33671) );
  NAND U34183 ( .A(n33672), .B(n33671), .Z(n33909) );
  XNOR U34184 ( .A(n38321), .B(b[25]), .Z(n33857) );
  NANDN U34185 ( .A(n34219), .B(n33857), .Z(n33675) );
  NAND U34186 ( .A(n33673), .B(n34217), .Z(n33674) );
  NAND U34187 ( .A(n33675), .B(n33674), .Z(n33910) );
  XNOR U34188 ( .A(n33909), .B(n33910), .Z(n33912) );
  XOR U34189 ( .A(n33911), .B(n33912), .Z(n33848) );
  NAND U34190 ( .A(n33676), .B(n35188), .Z(n33678) );
  XNOR U34191 ( .A(n38134), .B(b[29]), .Z(n33797) );
  NANDN U34192 ( .A(n34968), .B(n33797), .Z(n33677) );
  NAND U34193 ( .A(n33678), .B(n33677), .Z(n33905) );
  NAND U34194 ( .A(n33679), .B(n38326), .Z(n33681) );
  XNOR U34195 ( .A(n38400), .B(a[90]), .Z(n33854) );
  NANDN U34196 ( .A(n38273), .B(n33854), .Z(n33680) );
  AND U34197 ( .A(n33681), .B(n33680), .Z(n33904) );
  NAND U34198 ( .A(n37652), .B(n33682), .Z(n33684) );
  XOR U34199 ( .A(b[49]), .B(n36100), .Z(n33800) );
  OR U34200 ( .A(n33800), .B(n37756), .Z(n33683) );
  NAND U34201 ( .A(n33684), .B(n33683), .Z(n33903) );
  XNOR U34202 ( .A(n33904), .B(n33903), .Z(n33906) );
  XOR U34203 ( .A(n33905), .B(n33906), .Z(n33849) );
  XNOR U34204 ( .A(n33848), .B(n33849), .Z(n33850) );
  XOR U34205 ( .A(n33851), .B(n33850), .Z(n33934) );
  XOR U34206 ( .A(n33830), .B(n33831), .Z(n33833) );
  XNOR U34207 ( .A(n33832), .B(n33833), .Z(n33951) );
  XNOR U34208 ( .A(n33952), .B(n33951), .Z(n33946) );
  NANDN U34209 ( .A(n33686), .B(n33685), .Z(n33690) );
  NAND U34210 ( .A(n33688), .B(n33687), .Z(n33689) );
  NAND U34211 ( .A(n33690), .B(n33689), .Z(n33940) );
  NANDN U34212 ( .A(n33692), .B(n33691), .Z(n33696) );
  NAND U34213 ( .A(n33694), .B(n33693), .Z(n33695) );
  NAND U34214 ( .A(n33696), .B(n33695), .Z(n33937) );
  OR U34215 ( .A(n33698), .B(n33697), .Z(n33702) );
  NAND U34216 ( .A(n33700), .B(n33699), .Z(n33701) );
  NAND U34217 ( .A(n33702), .B(n33701), .Z(n33845) );
  NANDN U34218 ( .A(n33704), .B(n33703), .Z(n33708) );
  NAND U34219 ( .A(n33706), .B(n33705), .Z(n33707) );
  NAND U34220 ( .A(n33708), .B(n33707), .Z(n33843) );
  XOR U34221 ( .A(n977), .B(n36909), .Z(n33794) );
  NAND U34222 ( .A(n33794), .B(n37068), .Z(n33711) );
  NANDN U34223 ( .A(n33709), .B(n37069), .Z(n33710) );
  NAND U34224 ( .A(n33711), .B(n33710), .Z(n33882) );
  NAND U34225 ( .A(n33712), .B(n34044), .Z(n33714) );
  XOR U34226 ( .A(a[126]), .B(n34510), .Z(n33866) );
  OR U34227 ( .A(n33866), .B(n33867), .Z(n33713) );
  NAND U34228 ( .A(n33714), .B(n33713), .Z(n33879) );
  XOR U34229 ( .A(b[61]), .B(n34048), .Z(n33870) );
  OR U34230 ( .A(n33870), .B(n38371), .Z(n33717) );
  NANDN U34231 ( .A(n33715), .B(n38369), .Z(n33716) );
  AND U34232 ( .A(n33717), .B(n33716), .Z(n33880) );
  XNOR U34233 ( .A(n33879), .B(n33880), .Z(n33881) );
  XOR U34234 ( .A(n33882), .B(n33881), .Z(n33838) );
  XOR U34235 ( .A(a[116]), .B(n974), .Z(n33812) );
  NANDN U34236 ( .A(n33812), .B(n35620), .Z(n33720) );
  NAND U34237 ( .A(n33718), .B(n35621), .Z(n33719) );
  NAND U34238 ( .A(n33720), .B(n33719), .Z(n33888) );
  XOR U34239 ( .A(a[118]), .B(n973), .Z(n33806) );
  NANDN U34240 ( .A(n33806), .B(n35313), .Z(n33723) );
  NANDN U34241 ( .A(n33721), .B(n35311), .Z(n33722) );
  NAND U34242 ( .A(n33723), .B(n33722), .Z(n33885) );
  XOR U34243 ( .A(b[57]), .B(n34852), .Z(n33919) );
  OR U34244 ( .A(n33919), .B(n965), .Z(n33726) );
  NANDN U34245 ( .A(n33724), .B(n38194), .Z(n33725) );
  AND U34246 ( .A(n33726), .B(n33725), .Z(n33886) );
  XNOR U34247 ( .A(n33885), .B(n33886), .Z(n33887) );
  XOR U34248 ( .A(n33888), .B(n33887), .Z(n33836) );
  NANDN U34249 ( .A(n33728), .B(n33727), .Z(n33732) );
  NAND U34250 ( .A(n33730), .B(n33729), .Z(n33731) );
  NAND U34251 ( .A(n33732), .B(n33731), .Z(n33837) );
  XNOR U34252 ( .A(n33836), .B(n33837), .Z(n33839) );
  XNOR U34253 ( .A(n33838), .B(n33839), .Z(n33842) );
  XOR U34254 ( .A(n33843), .B(n33842), .Z(n33844) );
  XOR U34255 ( .A(n33845), .B(n33844), .Z(n33938) );
  XOR U34256 ( .A(n33937), .B(n33938), .Z(n33939) );
  XOR U34257 ( .A(n33940), .B(n33939), .Z(n33943) );
  OR U34258 ( .A(n33734), .B(n33733), .Z(n33738) );
  NAND U34259 ( .A(n33736), .B(n33735), .Z(n33737) );
  NAND U34260 ( .A(n33738), .B(n33737), .Z(n33944) );
  XNOR U34261 ( .A(n33943), .B(n33944), .Z(n33945) );
  XNOR U34262 ( .A(n33946), .B(n33945), .Z(n33774) );
  NANDN U34263 ( .A(n33740), .B(n33739), .Z(n33744) );
  OR U34264 ( .A(n33742), .B(n33741), .Z(n33743) );
  NAND U34265 ( .A(n33744), .B(n33743), .Z(n33775) );
  XOR U34266 ( .A(n33774), .B(n33775), .Z(n33776) );
  XNOR U34267 ( .A(n33777), .B(n33776), .Z(n33766) );
  NANDN U34268 ( .A(n33746), .B(n33745), .Z(n33750) );
  NANDN U34269 ( .A(n33748), .B(n33747), .Z(n33749) );
  NAND U34270 ( .A(n33750), .B(n33749), .Z(n33765) );
  XNOR U34271 ( .A(n33765), .B(n33764), .Z(n33767) );
  XOR U34272 ( .A(n33766), .B(n33767), .Z(n33955) );
  NANDN U34273 ( .A(n33756), .B(n33755), .Z(n33760) );
  NAND U34274 ( .A(n33758), .B(n33757), .Z(n33759) );
  AND U34275 ( .A(n33760), .B(n33759), .Z(n33956) );
  XNOR U34276 ( .A(n33955), .B(n33956), .Z(n33761) );
  XNOR U34277 ( .A(n33957), .B(n33761), .Z(n33762) );
  XOR U34278 ( .A(n33763), .B(n33762), .Z(c[212]) );
  OR U34279 ( .A(n33763), .B(n33762), .Z(n34154) );
  OR U34280 ( .A(n33769), .B(n33768), .Z(n33773) );
  NANDN U34281 ( .A(n33771), .B(n33770), .Z(n33772) );
  NAND U34282 ( .A(n33773), .B(n33772), .Z(n33965) );
  OR U34283 ( .A(n33775), .B(n33774), .Z(n33779) );
  NANDN U34284 ( .A(n33777), .B(n33776), .Z(n33778) );
  NAND U34285 ( .A(n33779), .B(n33778), .Z(n33962) );
  NANDN U34286 ( .A(n33781), .B(n33780), .Z(n33785) );
  NAND U34287 ( .A(n33783), .B(n33782), .Z(n33784) );
  NAND U34288 ( .A(n33785), .B(n33784), .Z(n34118) );
  NANDN U34289 ( .A(n33985), .B(n33786), .Z(n33790) );
  NANDN U34290 ( .A(n33788), .B(n33787), .Z(n33789) );
  NAND U34291 ( .A(n33790), .B(n33789), .Z(n34116) );
  XNOR U34292 ( .A(n33984), .B(n33985), .Z(n33987) );
  NANDN U34293 ( .A(n985), .B(a[85]), .Z(n33986) );
  XNOR U34294 ( .A(n33987), .B(n33986), .Z(n34109) );
  XNOR U34295 ( .A(n985), .B(a[87]), .Z(n34049) );
  NAND U34296 ( .A(n34049), .B(n38422), .Z(n33793) );
  NANDN U34297 ( .A(n33791), .B(n38423), .Z(n33792) );
  NAND U34298 ( .A(n33793), .B(n33792), .Z(n34110) );
  XNOR U34299 ( .A(n34109), .B(n34110), .Z(n34111) );
  NAND U34300 ( .A(n37069), .B(n33794), .Z(n33796) );
  XNOR U34301 ( .A(n977), .B(a[107]), .Z(n34097) );
  NAND U34302 ( .A(n34097), .B(n37068), .Z(n33795) );
  NAND U34303 ( .A(n33796), .B(n33795), .Z(n34112) );
  XNOR U34304 ( .A(n34111), .B(n34112), .Z(n34115) );
  XNOR U34305 ( .A(n34116), .B(n34115), .Z(n34117) );
  XNOR U34306 ( .A(n34118), .B(n34117), .Z(n34020) );
  NAND U34307 ( .A(n33797), .B(n35188), .Z(n33799) );
  XNOR U34308 ( .A(a[121]), .B(n35540), .Z(n33999) );
  NANDN U34309 ( .A(n34968), .B(n33999), .Z(n33798) );
  NAND U34310 ( .A(n33799), .B(n33798), .Z(n33993) );
  XNOR U34311 ( .A(b[49]), .B(a[101]), .Z(n34091) );
  OR U34312 ( .A(n34091), .B(n37756), .Z(n33802) );
  NANDN U34313 ( .A(n33800), .B(n37652), .Z(n33801) );
  NAND U34314 ( .A(n33802), .B(n33801), .Z(n33990) );
  XNOR U34315 ( .A(b[51]), .B(a[99]), .Z(n34067) );
  NANDN U34316 ( .A(n34067), .B(n37803), .Z(n33805) );
  NANDN U34317 ( .A(n33803), .B(n37802), .Z(n33804) );
  AND U34318 ( .A(n33805), .B(n33804), .Z(n33991) );
  XNOR U34319 ( .A(n33990), .B(n33991), .Z(n33992) );
  XNOR U34320 ( .A(n33993), .B(n33992), .Z(n34008) );
  XOR U34321 ( .A(a[119]), .B(n973), .Z(n34041) );
  NANDN U34322 ( .A(n34041), .B(n35313), .Z(n33808) );
  NANDN U34323 ( .A(n33806), .B(n35311), .Z(n33807) );
  NAND U34324 ( .A(n33808), .B(n33807), .Z(n34079) );
  XNOR U34325 ( .A(a[111]), .B(b[39]), .Z(n34035) );
  NANDN U34326 ( .A(n34035), .B(n36553), .Z(n33811) );
  NAND U34327 ( .A(n33809), .B(n36643), .Z(n33810) );
  NAND U34328 ( .A(n33811), .B(n33810), .Z(n34076) );
  XNOR U34329 ( .A(a[117]), .B(b[33]), .Z(n34088) );
  NANDN U34330 ( .A(n34088), .B(n35620), .Z(n33814) );
  NANDN U34331 ( .A(n33812), .B(n35621), .Z(n33813) );
  AND U34332 ( .A(n33814), .B(n33813), .Z(n34077) );
  XNOR U34333 ( .A(n34076), .B(n34077), .Z(n34078) );
  XNOR U34334 ( .A(n34079), .B(n34078), .Z(n34005) );
  NANDN U34335 ( .A(n33815), .B(n36309), .Z(n33817) );
  XNOR U34336 ( .A(a[113]), .B(n975), .Z(n34100) );
  NAND U34337 ( .A(n34100), .B(n36311), .Z(n33816) );
  NAND U34338 ( .A(n33817), .B(n33816), .Z(n34006) );
  XNOR U34339 ( .A(n34005), .B(n34006), .Z(n34007) );
  XOR U34340 ( .A(n34008), .B(n34007), .Z(n34017) );
  NANDN U34341 ( .A(n33819), .B(n33818), .Z(n33823) );
  OR U34342 ( .A(n33821), .B(n33820), .Z(n33822) );
  NAND U34343 ( .A(n33823), .B(n33822), .Z(n34018) );
  XOR U34344 ( .A(n34017), .B(n34018), .Z(n34019) );
  XNOR U34345 ( .A(n34020), .B(n34019), .Z(n34137) );
  NAND U34346 ( .A(n33825), .B(n33824), .Z(n33829) );
  NAND U34347 ( .A(n33827), .B(n33826), .Z(n33828) );
  AND U34348 ( .A(n33829), .B(n33828), .Z(n34138) );
  XNOR U34349 ( .A(n34137), .B(n34138), .Z(n34140) );
  NANDN U34350 ( .A(n33831), .B(n33830), .Z(n33835) );
  NANDN U34351 ( .A(n33833), .B(n33832), .Z(n33834) );
  NAND U34352 ( .A(n33835), .B(n33834), .Z(n34139) );
  XNOR U34353 ( .A(n34140), .B(n34139), .Z(n34150) );
  OR U34354 ( .A(n33837), .B(n33836), .Z(n33841) );
  OR U34355 ( .A(n33839), .B(n33838), .Z(n33840) );
  NAND U34356 ( .A(n33841), .B(n33840), .Z(n34026) );
  OR U34357 ( .A(n33843), .B(n33842), .Z(n33847) );
  NANDN U34358 ( .A(n33845), .B(n33844), .Z(n33846) );
  NAND U34359 ( .A(n33847), .B(n33846), .Z(n34023) );
  NANDN U34360 ( .A(n33849), .B(n33848), .Z(n33853) );
  NANDN U34361 ( .A(n33851), .B(n33850), .Z(n33852) );
  AND U34362 ( .A(n33853), .B(n33852), .Z(n34024) );
  XNOR U34363 ( .A(n34023), .B(n34024), .Z(n34025) );
  XNOR U34364 ( .A(n34026), .B(n34025), .Z(n34146) );
  NAND U34365 ( .A(n33854), .B(n38326), .Z(n33856) );
  XNOR U34366 ( .A(n38400), .B(a[91]), .Z(n34073) );
  NANDN U34367 ( .A(n38273), .B(n34073), .Z(n33855) );
  NAND U34368 ( .A(n33856), .B(n33855), .Z(n33981) );
  XOR U34369 ( .A(a[125]), .B(b[25]), .Z(n34064) );
  NANDN U34370 ( .A(n34219), .B(n34064), .Z(n33859) );
  NAND U34371 ( .A(n33857), .B(n34217), .Z(n33858) );
  NAND U34372 ( .A(n33859), .B(n33858), .Z(n33978) );
  NAND U34373 ( .A(n33860), .B(n37469), .Z(n33862) );
  XNOR U34374 ( .A(n978), .B(a[103]), .Z(n34002) );
  NAND U34375 ( .A(n37471), .B(n34002), .Z(n33861) );
  AND U34376 ( .A(n33862), .B(n33861), .Z(n33979) );
  XNOR U34377 ( .A(n33978), .B(n33979), .Z(n33980) );
  XOR U34378 ( .A(n33981), .B(n33980), .Z(n34125) );
  XOR U34379 ( .A(b[45]), .B(a[105]), .Z(n34058) );
  NAND U34380 ( .A(n37261), .B(n34058), .Z(n33865) );
  NANDN U34381 ( .A(n33863), .B(n37262), .Z(n33864) );
  NAND U34382 ( .A(n33865), .B(n33864), .Z(n33975) );
  NANDN U34383 ( .A(n33866), .B(n34044), .Z(n33869) );
  XNOR U34384 ( .A(n38463), .B(b[23]), .Z(n34045) );
  NANDN U34385 ( .A(n33867), .B(n34045), .Z(n33868) );
  NAND U34386 ( .A(n33869), .B(n33868), .Z(n33972) );
  XNOR U34387 ( .A(b[61]), .B(a[89]), .Z(n34061) );
  OR U34388 ( .A(n34061), .B(n38371), .Z(n33872) );
  NANDN U34389 ( .A(n33870), .B(n38369), .Z(n33871) );
  AND U34390 ( .A(n33872), .B(n33871), .Z(n33973) );
  XNOR U34391 ( .A(n33972), .B(n33973), .Z(n33974) );
  XOR U34392 ( .A(n33975), .B(n33974), .Z(n34126) );
  XNOR U34393 ( .A(n34125), .B(n34126), .Z(n34128) );
  NANDN U34394 ( .A(n33874), .B(n33873), .Z(n33878) );
  NAND U34395 ( .A(n33876), .B(n33875), .Z(n33877) );
  NAND U34396 ( .A(n33878), .B(n33877), .Z(n34127) );
  XNOR U34397 ( .A(n34128), .B(n34127), .Z(n34014) );
  NANDN U34398 ( .A(n33880), .B(n33879), .Z(n33884) );
  NAND U34399 ( .A(n33882), .B(n33881), .Z(n33883) );
  NAND U34400 ( .A(n33884), .B(n33883), .Z(n34011) );
  NANDN U34401 ( .A(n33886), .B(n33885), .Z(n33890) );
  NAND U34402 ( .A(n33888), .B(n33887), .Z(n33889) );
  AND U34403 ( .A(n33890), .B(n33889), .Z(n34012) );
  XNOR U34404 ( .A(n34011), .B(n34012), .Z(n34013) );
  XOR U34405 ( .A(n34014), .B(n34013), .Z(n34132) );
  OR U34406 ( .A(n33892), .B(n33891), .Z(n33896) );
  NAND U34407 ( .A(n33894), .B(n33893), .Z(n33895) );
  AND U34408 ( .A(n33896), .B(n33895), .Z(n34131) );
  XOR U34409 ( .A(n34132), .B(n34131), .Z(n34133) );
  NANDN U34410 ( .A(n33898), .B(n33897), .Z(n33902) );
  NAND U34411 ( .A(n33900), .B(n33899), .Z(n33901) );
  NAND U34412 ( .A(n33902), .B(n33901), .Z(n34029) );
  NANDN U34413 ( .A(n33904), .B(n33903), .Z(n33908) );
  NAND U34414 ( .A(n33906), .B(n33905), .Z(n33907) );
  NAND U34415 ( .A(n33908), .B(n33907), .Z(n34030) );
  XNOR U34416 ( .A(n34029), .B(n34030), .Z(n34031) );
  XOR U34417 ( .A(a[109]), .B(b[41]), .Z(n34106) );
  NANDN U34418 ( .A(n36905), .B(n34106), .Z(n33915) );
  NAND U34419 ( .A(n33913), .B(n36807), .Z(n33914) );
  NAND U34420 ( .A(n33915), .B(n33914), .Z(n34085) );
  XOR U34421 ( .A(b[55]), .B(n35628), .Z(n34038) );
  NANDN U34422 ( .A(n34038), .B(n38075), .Z(n33918) );
  NANDN U34423 ( .A(n33916), .B(n38073), .Z(n33917) );
  NAND U34424 ( .A(n33918), .B(n33917), .Z(n34082) );
  XOR U34425 ( .A(b[57]), .B(n35377), .Z(n34070) );
  OR U34426 ( .A(n34070), .B(n965), .Z(n33921) );
  NANDN U34427 ( .A(n33919), .B(n38194), .Z(n33920) );
  AND U34428 ( .A(n33921), .B(n33920), .Z(n34083) );
  XNOR U34429 ( .A(n34082), .B(n34083), .Z(n34084) );
  XNOR U34430 ( .A(n34085), .B(n34084), .Z(n34119) );
  XNOR U34431 ( .A(b[53]), .B(a[97]), .Z(n34094) );
  NANDN U34432 ( .A(n34094), .B(n37940), .Z(n33924) );
  NANDN U34433 ( .A(n33922), .B(n37941), .Z(n33923) );
  NAND U34434 ( .A(n33924), .B(n33923), .Z(n34055) );
  NAND U34435 ( .A(n33925), .B(n34848), .Z(n33927) );
  XNOR U34436 ( .A(a[123]), .B(b[27]), .Z(n33996) );
  NANDN U34437 ( .A(n33996), .B(n34618), .Z(n33926) );
  NAND U34438 ( .A(n33927), .B(n33926), .Z(n34052) );
  XOR U34439 ( .A(a[115]), .B(b[35]), .Z(n34103) );
  NAND U34440 ( .A(n35985), .B(n34103), .Z(n33930) );
  NANDN U34441 ( .A(n33928), .B(n35986), .Z(n33929) );
  AND U34442 ( .A(n33930), .B(n33929), .Z(n34053) );
  XNOR U34443 ( .A(n34052), .B(n34053), .Z(n34054) );
  XOR U34444 ( .A(n34055), .B(n34054), .Z(n34120) );
  XOR U34445 ( .A(n34119), .B(n34120), .Z(n34122) );
  XOR U34446 ( .A(n34121), .B(n34122), .Z(n34032) );
  XOR U34447 ( .A(n34031), .B(n34032), .Z(n34134) );
  XNOR U34448 ( .A(n34133), .B(n34134), .Z(n34143) );
  OR U34449 ( .A(n33932), .B(n33931), .Z(n33936) );
  OR U34450 ( .A(n33934), .B(n33933), .Z(n33935) );
  NAND U34451 ( .A(n33936), .B(n33935), .Z(n34144) );
  XNOR U34452 ( .A(n34143), .B(n34144), .Z(n34145) );
  XOR U34453 ( .A(n34146), .B(n34145), .Z(n34148) );
  OR U34454 ( .A(n33938), .B(n33937), .Z(n33942) );
  NANDN U34455 ( .A(n33940), .B(n33939), .Z(n33941) );
  AND U34456 ( .A(n33942), .B(n33941), .Z(n34147) );
  XOR U34457 ( .A(n34148), .B(n34147), .Z(n34149) );
  XNOR U34458 ( .A(n34150), .B(n34149), .Z(n33968) );
  NANDN U34459 ( .A(n33944), .B(n33943), .Z(n33948) );
  NANDN U34460 ( .A(n33946), .B(n33945), .Z(n33947) );
  AND U34461 ( .A(n33948), .B(n33947), .Z(n33969) );
  XNOR U34462 ( .A(n33968), .B(n33969), .Z(n33970) );
  OR U34463 ( .A(n33950), .B(n33949), .Z(n33954) );
  NANDN U34464 ( .A(n33952), .B(n33951), .Z(n33953) );
  AND U34465 ( .A(n33954), .B(n33953), .Z(n33971) );
  XNOR U34466 ( .A(n33970), .B(n33971), .Z(n33963) );
  XOR U34467 ( .A(n33962), .B(n33963), .Z(n33964) );
  XOR U34468 ( .A(n33965), .B(n33964), .Z(n33959) );
  XOR U34469 ( .A(n33959), .B(n33961), .Z(n33958) );
  XNOR U34470 ( .A(n33960), .B(n33958), .Z(n34153) );
  XNOR U34471 ( .A(n34154), .B(n34153), .Z(c[213]) );
  OR U34472 ( .A(n33963), .B(n33962), .Z(n33967) );
  NAND U34473 ( .A(n33965), .B(n33964), .Z(n33966) );
  NAND U34474 ( .A(n33967), .B(n33966), .Z(n34155) );
  NANDN U34475 ( .A(n33973), .B(n33972), .Z(n33977) );
  NAND U34476 ( .A(n33975), .B(n33974), .Z(n33976) );
  NAND U34477 ( .A(n33977), .B(n33976), .Z(n34177) );
  NANDN U34478 ( .A(n33979), .B(n33978), .Z(n33983) );
  NAND U34479 ( .A(n33981), .B(n33980), .Z(n33982) );
  AND U34480 ( .A(n33983), .B(n33982), .Z(n34178) );
  XNOR U34481 ( .A(n34177), .B(n34178), .Z(n34179) );
  NAND U34482 ( .A(n33985), .B(n33984), .Z(n33989) );
  OR U34483 ( .A(n33987), .B(n33986), .Z(n33988) );
  AND U34484 ( .A(n33989), .B(n33988), .Z(n34315) );
  NANDN U34485 ( .A(n33991), .B(n33990), .Z(n33995) );
  NAND U34486 ( .A(n33993), .B(n33992), .Z(n33994) );
  AND U34487 ( .A(n33995), .B(n33994), .Z(n34316) );
  XOR U34488 ( .A(n34315), .B(n34316), .Z(n34318) );
  NANDN U34489 ( .A(n33996), .B(n34848), .Z(n33998) );
  XNOR U34490 ( .A(n38321), .B(b[27]), .Z(n34276) );
  NAND U34491 ( .A(n34618), .B(n34276), .Z(n33997) );
  AND U34492 ( .A(n33998), .B(n33997), .Z(n34195) );
  NAND U34493 ( .A(n33999), .B(n35188), .Z(n34001) );
  XOR U34494 ( .A(n38251), .B(n35540), .Z(n34294) );
  NANDN U34495 ( .A(n34968), .B(n34294), .Z(n34000) );
  AND U34496 ( .A(n34001), .B(n34000), .Z(n34196) );
  XNOR U34497 ( .A(n34195), .B(n34196), .Z(n34197) );
  NAND U34498 ( .A(n34002), .B(n37469), .Z(n34004) );
  XOR U34499 ( .A(n978), .B(n36647), .Z(n34297) );
  NAND U34500 ( .A(n34297), .B(n37471), .Z(n34003) );
  AND U34501 ( .A(n34004), .B(n34003), .Z(n34198) );
  XNOR U34502 ( .A(n34318), .B(n34317), .Z(n34180) );
  XOR U34503 ( .A(n34179), .B(n34180), .Z(n34228) );
  NANDN U34504 ( .A(n34006), .B(n34005), .Z(n34010) );
  NAND U34505 ( .A(n34008), .B(n34007), .Z(n34009) );
  NAND U34506 ( .A(n34010), .B(n34009), .Z(n34225) );
  NANDN U34507 ( .A(n34012), .B(n34011), .Z(n34016) );
  NAND U34508 ( .A(n34014), .B(n34013), .Z(n34015) );
  NAND U34509 ( .A(n34016), .B(n34015), .Z(n34226) );
  XNOR U34510 ( .A(n34225), .B(n34226), .Z(n34227) );
  XNOR U34511 ( .A(n34228), .B(n34227), .Z(n34331) );
  OR U34512 ( .A(n34018), .B(n34017), .Z(n34022) );
  NANDN U34513 ( .A(n34020), .B(n34019), .Z(n34021) );
  AND U34514 ( .A(n34022), .B(n34021), .Z(n34332) );
  XNOR U34515 ( .A(n34331), .B(n34332), .Z(n34333) );
  NANDN U34516 ( .A(n34024), .B(n34023), .Z(n34028) );
  NAND U34517 ( .A(n34026), .B(n34025), .Z(n34027) );
  AND U34518 ( .A(n34028), .B(n34027), .Z(n34334) );
  XNOR U34519 ( .A(n34333), .B(n34334), .Z(n34169) );
  NANDN U34520 ( .A(n34030), .B(n34029), .Z(n34034) );
  NAND U34521 ( .A(n34032), .B(n34031), .Z(n34033) );
  NAND U34522 ( .A(n34034), .B(n34033), .Z(n34329) );
  XOR U34523 ( .A(a[112]), .B(n976), .Z(n34207) );
  NANDN U34524 ( .A(n34207), .B(n36553), .Z(n34037) );
  NANDN U34525 ( .A(n34035), .B(n36643), .Z(n34036) );
  NAND U34526 ( .A(n34037), .B(n34036), .Z(n34204) );
  XOR U34527 ( .A(b[55]), .B(n35545), .Z(n34261) );
  NANDN U34528 ( .A(n34261), .B(n38075), .Z(n34040) );
  NANDN U34529 ( .A(n34038), .B(n38073), .Z(n34039) );
  NAND U34530 ( .A(n34040), .B(n34039), .Z(n34201) );
  XOR U34531 ( .A(a[120]), .B(n973), .Z(n34291) );
  NANDN U34532 ( .A(n34291), .B(n35313), .Z(n34043) );
  NANDN U34533 ( .A(n34041), .B(n35311), .Z(n34042) );
  AND U34534 ( .A(n34043), .B(n34042), .Z(n34202) );
  XNOR U34535 ( .A(n34201), .B(n34202), .Z(n34203) );
  XOR U34536 ( .A(n34204), .B(n34203), .Z(n34235) );
  NAND U34537 ( .A(n34045), .B(n34044), .Z(n34047) );
  ANDN U34538 ( .B(n34047), .A(n34046), .Z(n34255) );
  AND U34539 ( .A(a[86]), .B(b[63]), .Z(n34467) );
  XOR U34540 ( .A(b[63]), .B(n34048), .Z(n34279) );
  NANDN U34541 ( .A(n34279), .B(n38422), .Z(n34051) );
  NAND U34542 ( .A(n34049), .B(n38423), .Z(n34050) );
  NAND U34543 ( .A(n34051), .B(n34050), .Z(n34253) );
  XNOR U34544 ( .A(n34467), .B(n34253), .Z(n34254) );
  XNOR U34545 ( .A(n34255), .B(n34254), .Z(n34236) );
  XNOR U34546 ( .A(n34235), .B(n34236), .Z(n34238) );
  NANDN U34547 ( .A(n34053), .B(n34052), .Z(n34057) );
  NAND U34548 ( .A(n34055), .B(n34054), .Z(n34056) );
  NAND U34549 ( .A(n34057), .B(n34056), .Z(n34237) );
  XNOR U34550 ( .A(n34238), .B(n34237), .Z(n34173) );
  XNOR U34551 ( .A(b[45]), .B(n36909), .Z(n34222) );
  NAND U34552 ( .A(n34222), .B(n37261), .Z(n34060) );
  NAND U34553 ( .A(n34058), .B(n37262), .Z(n34059) );
  NAND U34554 ( .A(n34060), .B(n34059), .Z(n34192) );
  XOR U34555 ( .A(b[61]), .B(n34851), .Z(n34273) );
  OR U34556 ( .A(n34273), .B(n38371), .Z(n34063) );
  NANDN U34557 ( .A(n34061), .B(n38369), .Z(n34062) );
  NAND U34558 ( .A(n34063), .B(n34062), .Z(n34189) );
  XNOR U34559 ( .A(a[126]), .B(b[25]), .Z(n34218) );
  OR U34560 ( .A(n34218), .B(n34219), .Z(n34066) );
  NAND U34561 ( .A(n34064), .B(n34217), .Z(n34065) );
  AND U34562 ( .A(n34066), .B(n34065), .Z(n34190) );
  XNOR U34563 ( .A(n34189), .B(n34190), .Z(n34191) );
  XNOR U34564 ( .A(n34192), .B(n34191), .Z(n34321) );
  XOR U34565 ( .A(b[51]), .B(n36100), .Z(n34267) );
  NANDN U34566 ( .A(n34267), .B(n37803), .Z(n34069) );
  NANDN U34567 ( .A(n34067), .B(n37802), .Z(n34068) );
  NAND U34568 ( .A(n34069), .B(n34068), .Z(n34312) );
  XOR U34569 ( .A(b[57]), .B(n35191), .Z(n34264) );
  OR U34570 ( .A(n34264), .B(n965), .Z(n34072) );
  NANDN U34571 ( .A(n34070), .B(n38194), .Z(n34071) );
  NAND U34572 ( .A(n34072), .B(n34071), .Z(n34309) );
  NAND U34573 ( .A(n38326), .B(n34073), .Z(n34075) );
  XOR U34574 ( .A(n38400), .B(n34852), .Z(n34270) );
  NANDN U34575 ( .A(n38273), .B(n34270), .Z(n34074) );
  AND U34576 ( .A(n34075), .B(n34074), .Z(n34310) );
  XNOR U34577 ( .A(n34309), .B(n34310), .Z(n34311) );
  XOR U34578 ( .A(n34312), .B(n34311), .Z(n34322) );
  XOR U34579 ( .A(n34321), .B(n34322), .Z(n34324) );
  NANDN U34580 ( .A(n34077), .B(n34076), .Z(n34081) );
  NAND U34581 ( .A(n34079), .B(n34078), .Z(n34080) );
  NAND U34582 ( .A(n34081), .B(n34080), .Z(n34323) );
  XOR U34583 ( .A(n34324), .B(n34323), .Z(n34174) );
  XNOR U34584 ( .A(n34173), .B(n34174), .Z(n34175) );
  NANDN U34585 ( .A(n34083), .B(n34082), .Z(n34087) );
  NAND U34586 ( .A(n34085), .B(n34084), .Z(n34086) );
  AND U34587 ( .A(n34087), .B(n34086), .Z(n34241) );
  XOR U34588 ( .A(a[118]), .B(n974), .Z(n34306) );
  NANDN U34589 ( .A(n34306), .B(n35620), .Z(n34090) );
  NANDN U34590 ( .A(n34088), .B(n35621), .Z(n34089) );
  NAND U34591 ( .A(n34090), .B(n34089), .Z(n34288) );
  XOR U34592 ( .A(b[49]), .B(n36420), .Z(n34282) );
  OR U34593 ( .A(n34282), .B(n37756), .Z(n34093) );
  NANDN U34594 ( .A(n34091), .B(n37652), .Z(n34092) );
  NAND U34595 ( .A(n34093), .B(n34092), .Z(n34285) );
  XOR U34596 ( .A(b[53]), .B(n35783), .Z(n34300) );
  NANDN U34597 ( .A(n34300), .B(n37940), .Z(n34096) );
  NANDN U34598 ( .A(n34094), .B(n37941), .Z(n34095) );
  AND U34599 ( .A(n34096), .B(n34095), .Z(n34286) );
  XNOR U34600 ( .A(n34285), .B(n34286), .Z(n34287) );
  XNOR U34601 ( .A(n34288), .B(n34287), .Z(n34186) );
  NAND U34602 ( .A(n37069), .B(n34097), .Z(n34099) );
  XNOR U34603 ( .A(n977), .B(a[108]), .Z(n34210) );
  NAND U34604 ( .A(n34210), .B(n37068), .Z(n34098) );
  AND U34605 ( .A(n34099), .B(n34098), .Z(n34247) );
  XOR U34606 ( .A(a[114]), .B(n975), .Z(n34258) );
  NANDN U34607 ( .A(n34258), .B(n36311), .Z(n34102) );
  NAND U34608 ( .A(n34100), .B(n36309), .Z(n34101) );
  AND U34609 ( .A(n34102), .B(n34101), .Z(n34248) );
  XOR U34610 ( .A(n34247), .B(n34248), .Z(n34249) );
  XNOR U34611 ( .A(a[116]), .B(b[35]), .Z(n34303) );
  NANDN U34612 ( .A(n34303), .B(n35985), .Z(n34105) );
  NAND U34613 ( .A(n34103), .B(n35986), .Z(n34104) );
  AND U34614 ( .A(n34105), .B(n34104), .Z(n34250) );
  XNOR U34615 ( .A(n34249), .B(n34250), .Z(n34183) );
  NAND U34616 ( .A(n36807), .B(n34106), .Z(n34108) );
  XNOR U34617 ( .A(n37336), .B(b[41]), .Z(n34213) );
  NANDN U34618 ( .A(n36905), .B(n34213), .Z(n34107) );
  NAND U34619 ( .A(n34108), .B(n34107), .Z(n34184) );
  XOR U34620 ( .A(n34183), .B(n34184), .Z(n34185) );
  XOR U34621 ( .A(n34186), .B(n34185), .Z(n34242) );
  XNOR U34622 ( .A(n34241), .B(n34242), .Z(n34243) );
  NANDN U34623 ( .A(n34110), .B(n34109), .Z(n34114) );
  NANDN U34624 ( .A(n34112), .B(n34111), .Z(n34113) );
  NAND U34625 ( .A(n34114), .B(n34113), .Z(n34244) );
  XOR U34626 ( .A(n34175), .B(n34176), .Z(n34327) );
  NANDN U34627 ( .A(n34120), .B(n34119), .Z(n34124) );
  OR U34628 ( .A(n34122), .B(n34121), .Z(n34123) );
  NAND U34629 ( .A(n34124), .B(n34123), .Z(n34231) );
  OR U34630 ( .A(n34126), .B(n34125), .Z(n34130) );
  OR U34631 ( .A(n34128), .B(n34127), .Z(n34129) );
  AND U34632 ( .A(n34130), .B(n34129), .Z(n34232) );
  XNOR U34633 ( .A(n34231), .B(n34232), .Z(n34234) );
  XOR U34634 ( .A(n34233), .B(n34234), .Z(n34328) );
  XNOR U34635 ( .A(n34327), .B(n34328), .Z(n34330) );
  XOR U34636 ( .A(n34329), .B(n34330), .Z(n34167) );
  OR U34637 ( .A(n34132), .B(n34131), .Z(n34136) );
  NAND U34638 ( .A(n34134), .B(n34133), .Z(n34135) );
  NAND U34639 ( .A(n34136), .B(n34135), .Z(n34168) );
  XOR U34640 ( .A(n34167), .B(n34168), .Z(n34170) );
  XNOR U34641 ( .A(n34169), .B(n34170), .Z(n34161) );
  NAND U34642 ( .A(n34138), .B(n34137), .Z(n34142) );
  OR U34643 ( .A(n34140), .B(n34139), .Z(n34141) );
  NAND U34644 ( .A(n34142), .B(n34141), .Z(n34162) );
  XNOR U34645 ( .A(n34161), .B(n34162), .Z(n34163) );
  XOR U34646 ( .A(n34163), .B(n34164), .Z(n34337) );
  OR U34647 ( .A(n34148), .B(n34147), .Z(n34152) );
  NAND U34648 ( .A(n34150), .B(n34149), .Z(n34151) );
  NAND U34649 ( .A(n34152), .B(n34151), .Z(n34338) );
  XNOR U34650 ( .A(n34337), .B(n34338), .Z(n34339) );
  XNOR U34651 ( .A(n34340), .B(n34339), .Z(n34156) );
  XNOR U34652 ( .A(n34155), .B(n34156), .Z(n34158) );
  XOR U34653 ( .A(n34157), .B(n34158), .Z(n34343) );
  NANDN U34654 ( .A(n34154), .B(n34153), .Z(n34344) );
  XNOR U34655 ( .A(n34343), .B(n34344), .Z(c[214]) );
  NANDN U34656 ( .A(n34156), .B(n34155), .Z(n34160) );
  NAND U34657 ( .A(n34158), .B(n34157), .Z(n34159) );
  NAND U34658 ( .A(n34160), .B(n34159), .Z(n34350) );
  NANDN U34659 ( .A(n34162), .B(n34161), .Z(n34166) );
  NANDN U34660 ( .A(n34164), .B(n34163), .Z(n34165) );
  NAND U34661 ( .A(n34166), .B(n34165), .Z(n34356) );
  NANDN U34662 ( .A(n34168), .B(n34167), .Z(n34172) );
  OR U34663 ( .A(n34170), .B(n34169), .Z(n34171) );
  NAND U34664 ( .A(n34172), .B(n34171), .Z(n34353) );
  NANDN U34665 ( .A(n34178), .B(n34177), .Z(n34182) );
  NANDN U34666 ( .A(n34180), .B(n34179), .Z(n34181) );
  NAND U34667 ( .A(n34182), .B(n34181), .Z(n34389) );
  OR U34668 ( .A(n34184), .B(n34183), .Z(n34188) );
  NAND U34669 ( .A(n34186), .B(n34185), .Z(n34187) );
  NAND U34670 ( .A(n34188), .B(n34187), .Z(n34390) );
  XNOR U34671 ( .A(n34389), .B(n34390), .Z(n34391) );
  NANDN U34672 ( .A(n34190), .B(n34189), .Z(n34194) );
  NAND U34673 ( .A(n34192), .B(n34191), .Z(n34193) );
  AND U34674 ( .A(n34194), .B(n34193), .Z(n34374) );
  OR U34675 ( .A(n34196), .B(n34195), .Z(n34200) );
  OR U34676 ( .A(n34198), .B(n34197), .Z(n34199) );
  AND U34677 ( .A(n34200), .B(n34199), .Z(n34371) );
  NANDN U34678 ( .A(n34202), .B(n34201), .Z(n34206) );
  NAND U34679 ( .A(n34204), .B(n34203), .Z(n34205) );
  NAND U34680 ( .A(n34206), .B(n34205), .Z(n34496) );
  XNOR U34681 ( .A(a[113]), .B(b[39]), .Z(n34479) );
  NANDN U34682 ( .A(n34479), .B(n36553), .Z(n34209) );
  NANDN U34683 ( .A(n34207), .B(n36643), .Z(n34208) );
  NAND U34684 ( .A(n34209), .B(n34208), .Z(n34485) );
  XNOR U34685 ( .A(b[43]), .B(a[109]), .Z(n34473) );
  NANDN U34686 ( .A(n34473), .B(n37068), .Z(n34212) );
  NAND U34687 ( .A(n34210), .B(n37069), .Z(n34211) );
  NAND U34688 ( .A(n34212), .B(n34211), .Z(n34482) );
  XOR U34689 ( .A(a[111]), .B(b[41]), .Z(n34476) );
  NANDN U34690 ( .A(n36905), .B(n34476), .Z(n34215) );
  NAND U34691 ( .A(n34213), .B(n36807), .Z(n34214) );
  AND U34692 ( .A(n34215), .B(n34214), .Z(n34483) );
  XNOR U34693 ( .A(n34482), .B(n34483), .Z(n34484) );
  XNOR U34694 ( .A(n34485), .B(n34484), .Z(n34494) );
  NAND U34695 ( .A(b[22]), .B(b[21]), .Z(n34216) );
  NAND U34696 ( .A(b[23]), .B(n34216), .Z(n34468) );
  XNOR U34697 ( .A(n34468), .B(n34467), .Z(n34470) );
  NANDN U34698 ( .A(n985), .B(a[87]), .Z(n34469) );
  XNOR U34699 ( .A(n34470), .B(n34469), .Z(n34488) );
  NANDN U34700 ( .A(n34218), .B(n34217), .Z(n34221) );
  XNOR U34701 ( .A(a[127]), .B(b[25]), .Z(n34511) );
  OR U34702 ( .A(n34511), .B(n34219), .Z(n34220) );
  NAND U34703 ( .A(n34221), .B(n34220), .Z(n34489) );
  XNOR U34704 ( .A(n34488), .B(n34489), .Z(n34490) );
  NAND U34705 ( .A(n37262), .B(n34222), .Z(n34224) );
  XOR U34706 ( .A(b[45]), .B(a[107]), .Z(n34440) );
  NAND U34707 ( .A(n37261), .B(n34440), .Z(n34223) );
  AND U34708 ( .A(n34224), .B(n34223), .Z(n34491) );
  XNOR U34709 ( .A(n34490), .B(n34491), .Z(n34495) );
  XOR U34710 ( .A(n34494), .B(n34495), .Z(n34497) );
  XOR U34711 ( .A(n34496), .B(n34497), .Z(n34372) );
  XNOR U34712 ( .A(n34371), .B(n34372), .Z(n34373) );
  XNOR U34713 ( .A(n34391), .B(n34392), .Z(n34359) );
  XNOR U34714 ( .A(n34360), .B(n34359), .Z(n34362) );
  NANDN U34715 ( .A(n34226), .B(n34225), .Z(n34230) );
  NAND U34716 ( .A(n34228), .B(n34227), .Z(n34229) );
  AND U34717 ( .A(n34230), .B(n34229), .Z(n34361) );
  XNOR U34718 ( .A(n34362), .B(n34361), .Z(n34533) );
  OR U34719 ( .A(n34236), .B(n34235), .Z(n34240) );
  OR U34720 ( .A(n34238), .B(n34237), .Z(n34239) );
  NAND U34721 ( .A(n34240), .B(n34239), .Z(n34527) );
  OR U34722 ( .A(n34242), .B(n34241), .Z(n34246) );
  OR U34723 ( .A(n34244), .B(n34243), .Z(n34245) );
  NAND U34724 ( .A(n34246), .B(n34245), .Z(n34525) );
  OR U34725 ( .A(n34248), .B(n34247), .Z(n34252) );
  NANDN U34726 ( .A(n34250), .B(n34249), .Z(n34251) );
  NAND U34727 ( .A(n34252), .B(n34251), .Z(n34368) );
  NANDN U34728 ( .A(n34467), .B(n34253), .Z(n34257) );
  NANDN U34729 ( .A(n34255), .B(n34254), .Z(n34256) );
  NAND U34730 ( .A(n34257), .B(n34256), .Z(n34366) );
  XNOR U34731 ( .A(a[115]), .B(b[37]), .Z(n34401) );
  NANDN U34732 ( .A(n34401), .B(n36311), .Z(n34260) );
  NANDN U34733 ( .A(n34258), .B(n36309), .Z(n34259) );
  NAND U34734 ( .A(n34260), .B(n34259), .Z(n34398) );
  XNOR U34735 ( .A(b[55]), .B(a[97]), .Z(n34407) );
  NANDN U34736 ( .A(n34407), .B(n38075), .Z(n34263) );
  NANDN U34737 ( .A(n34261), .B(n38073), .Z(n34262) );
  NAND U34738 ( .A(n34263), .B(n34262), .Z(n34395) );
  XOR U34739 ( .A(b[57]), .B(n35628), .Z(n34434) );
  OR U34740 ( .A(n34434), .B(n965), .Z(n34266) );
  NANDN U34741 ( .A(n34264), .B(n38194), .Z(n34265) );
  AND U34742 ( .A(n34266), .B(n34265), .Z(n34396) );
  XNOR U34743 ( .A(n34395), .B(n34396), .Z(n34397) );
  XOR U34744 ( .A(n34398), .B(n34397), .Z(n34365) );
  XNOR U34745 ( .A(n34366), .B(n34365), .Z(n34367) );
  XNOR U34746 ( .A(n34368), .B(n34367), .Z(n34380) );
  XNOR U34747 ( .A(b[51]), .B(a[101]), .Z(n34425) );
  NANDN U34748 ( .A(n34425), .B(n37803), .Z(n34269) );
  NANDN U34749 ( .A(n34267), .B(n37802), .Z(n34268) );
  NAND U34750 ( .A(n34269), .B(n34268), .Z(n34503) );
  NAND U34751 ( .A(n38326), .B(n34270), .Z(n34272) );
  XOR U34752 ( .A(n38400), .B(n35377), .Z(n34437) );
  NANDN U34753 ( .A(n38273), .B(n34437), .Z(n34271) );
  NAND U34754 ( .A(n34272), .B(n34271), .Z(n34500) );
  XNOR U34755 ( .A(b[61]), .B(a[91]), .Z(n34413) );
  OR U34756 ( .A(n34413), .B(n38371), .Z(n34275) );
  NANDN U34757 ( .A(n34273), .B(n38369), .Z(n34274) );
  AND U34758 ( .A(n34275), .B(n34274), .Z(n34501) );
  XNOR U34759 ( .A(n34500), .B(n34501), .Z(n34502) );
  XNOR U34760 ( .A(n34503), .B(n34502), .Z(n34452) );
  NAND U34761 ( .A(n34276), .B(n34848), .Z(n34278) );
  XNOR U34762 ( .A(a[125]), .B(n35375), .Z(n34416) );
  NAND U34763 ( .A(n34618), .B(n34416), .Z(n34277) );
  NAND U34764 ( .A(n34278), .B(n34277), .Z(n34446) );
  XNOR U34765 ( .A(b[63]), .B(a[89]), .Z(n34506) );
  NANDN U34766 ( .A(n34506), .B(n38422), .Z(n34281) );
  NANDN U34767 ( .A(n34279), .B(n38423), .Z(n34280) );
  NAND U34768 ( .A(n34281), .B(n34280), .Z(n34443) );
  XNOR U34769 ( .A(b[49]), .B(a[103]), .Z(n34515) );
  OR U34770 ( .A(n34515), .B(n37756), .Z(n34284) );
  NANDN U34771 ( .A(n34282), .B(n37652), .Z(n34283) );
  AND U34772 ( .A(n34284), .B(n34283), .Z(n34444) );
  XNOR U34773 ( .A(n34443), .B(n34444), .Z(n34445) );
  XNOR U34774 ( .A(n34446), .B(n34445), .Z(n34449) );
  NANDN U34775 ( .A(n34286), .B(n34285), .Z(n34290) );
  NAND U34776 ( .A(n34288), .B(n34287), .Z(n34289) );
  NAND U34777 ( .A(n34290), .B(n34289), .Z(n34450) );
  XNOR U34778 ( .A(n34449), .B(n34450), .Z(n34451) );
  XOR U34779 ( .A(n34452), .B(n34451), .Z(n34378) );
  XNOR U34780 ( .A(a[121]), .B(b[31]), .Z(n34518) );
  NANDN U34781 ( .A(n34518), .B(n35313), .Z(n34293) );
  NANDN U34782 ( .A(n34291), .B(n35311), .Z(n34292) );
  NAND U34783 ( .A(n34293), .B(n34292), .Z(n34464) );
  NAND U34784 ( .A(n35188), .B(n34294), .Z(n34296) );
  XNOR U34785 ( .A(a[123]), .B(n35540), .Z(n34521) );
  NANDN U34786 ( .A(n34968), .B(n34521), .Z(n34295) );
  NAND U34787 ( .A(n34296), .B(n34295), .Z(n34461) );
  NAND U34788 ( .A(n37469), .B(n34297), .Z(n34299) );
  XNOR U34789 ( .A(n978), .B(a[105]), .Z(n34410) );
  NAND U34790 ( .A(n34410), .B(n37471), .Z(n34298) );
  AND U34791 ( .A(n34299), .B(n34298), .Z(n34462) );
  XNOR U34792 ( .A(n34461), .B(n34462), .Z(n34463) );
  XNOR U34793 ( .A(n34464), .B(n34463), .Z(n34455) );
  XNOR U34794 ( .A(b[53]), .B(a[99]), .Z(n34404) );
  NANDN U34795 ( .A(n34404), .B(n37940), .Z(n34302) );
  NANDN U34796 ( .A(n34300), .B(n37941), .Z(n34301) );
  NAND U34797 ( .A(n34302), .B(n34301), .Z(n34422) );
  XOR U34798 ( .A(a[117]), .B(b[35]), .Z(n34428) );
  NAND U34799 ( .A(n35985), .B(n34428), .Z(n34305) );
  NANDN U34800 ( .A(n34303), .B(n35986), .Z(n34304) );
  NAND U34801 ( .A(n34305), .B(n34304), .Z(n34419) );
  XOR U34802 ( .A(a[119]), .B(n974), .Z(n34431) );
  NANDN U34803 ( .A(n34431), .B(n35620), .Z(n34308) );
  NANDN U34804 ( .A(n34306), .B(n35621), .Z(n34307) );
  AND U34805 ( .A(n34308), .B(n34307), .Z(n34420) );
  XNOR U34806 ( .A(n34419), .B(n34420), .Z(n34421) );
  XOR U34807 ( .A(n34422), .B(n34421), .Z(n34456) );
  XOR U34808 ( .A(n34455), .B(n34456), .Z(n34458) );
  NANDN U34809 ( .A(n34310), .B(n34309), .Z(n34314) );
  NAND U34810 ( .A(n34312), .B(n34311), .Z(n34313) );
  NAND U34811 ( .A(n34314), .B(n34313), .Z(n34457) );
  XOR U34812 ( .A(n34458), .B(n34457), .Z(n34377) );
  XOR U34813 ( .A(n34378), .B(n34377), .Z(n34379) );
  XOR U34814 ( .A(n34380), .B(n34379), .Z(n34385) );
  OR U34815 ( .A(n34316), .B(n34315), .Z(n34320) );
  NAND U34816 ( .A(n34318), .B(n34317), .Z(n34319) );
  NAND U34817 ( .A(n34320), .B(n34319), .Z(n34383) );
  NANDN U34818 ( .A(n34322), .B(n34321), .Z(n34326) );
  OR U34819 ( .A(n34324), .B(n34323), .Z(n34325) );
  NAND U34820 ( .A(n34326), .B(n34325), .Z(n34384) );
  XNOR U34821 ( .A(n34383), .B(n34384), .Z(n34386) );
  XOR U34822 ( .A(n34385), .B(n34386), .Z(n34524) );
  XNOR U34823 ( .A(n34525), .B(n34524), .Z(n34526) );
  XOR U34824 ( .A(n34527), .B(n34526), .Z(n34530) );
  XNOR U34825 ( .A(n34531), .B(n34530), .Z(n34532) );
  XOR U34826 ( .A(n34533), .B(n34532), .Z(n34537) );
  NANDN U34827 ( .A(n34332), .B(n34331), .Z(n34336) );
  NAND U34828 ( .A(n34334), .B(n34333), .Z(n34335) );
  NAND U34829 ( .A(n34336), .B(n34335), .Z(n34535) );
  XNOR U34830 ( .A(n34534), .B(n34535), .Z(n34536) );
  XOR U34831 ( .A(n34537), .B(n34536), .Z(n34354) );
  XOR U34832 ( .A(n34353), .B(n34354), .Z(n34355) );
  XNOR U34833 ( .A(n34356), .B(n34355), .Z(n34347) );
  NANDN U34834 ( .A(n34338), .B(n34337), .Z(n34342) );
  NAND U34835 ( .A(n34340), .B(n34339), .Z(n34341) );
  AND U34836 ( .A(n34342), .B(n34341), .Z(n34348) );
  XNOR U34837 ( .A(n34347), .B(n34348), .Z(n34349) );
  XNOR U34838 ( .A(n34350), .B(n34349), .Z(n34346) );
  NANDN U34839 ( .A(n34344), .B(n34343), .Z(n34345) );
  XOR U34840 ( .A(n34346), .B(n34345), .Z(c[215]) );
  OR U34841 ( .A(n34346), .B(n34345), .Z(n34726) );
  NANDN U34842 ( .A(n34348), .B(n34347), .Z(n34352) );
  NAND U34843 ( .A(n34350), .B(n34349), .Z(n34351) );
  AND U34844 ( .A(n34352), .B(n34351), .Z(n34545) );
  OR U34845 ( .A(n34354), .B(n34353), .Z(n34358) );
  NAND U34846 ( .A(n34356), .B(n34355), .Z(n34357) );
  AND U34847 ( .A(n34358), .B(n34357), .Z(n34542) );
  NAND U34848 ( .A(n34360), .B(n34359), .Z(n34364) );
  NANDN U34849 ( .A(n34362), .B(n34361), .Z(n34363) );
  NAND U34850 ( .A(n34364), .B(n34363), .Z(n34549) );
  OR U34851 ( .A(n34366), .B(n34365), .Z(n34370) );
  OR U34852 ( .A(n34368), .B(n34367), .Z(n34369) );
  NAND U34853 ( .A(n34370), .B(n34369), .Z(n34716) );
  OR U34854 ( .A(n34372), .B(n34371), .Z(n34376) );
  OR U34855 ( .A(n34374), .B(n34373), .Z(n34375) );
  NAND U34856 ( .A(n34376), .B(n34375), .Z(n34713) );
  OR U34857 ( .A(n34378), .B(n34377), .Z(n34382) );
  NAND U34858 ( .A(n34380), .B(n34379), .Z(n34381) );
  AND U34859 ( .A(n34382), .B(n34381), .Z(n34714) );
  XNOR U34860 ( .A(n34713), .B(n34714), .Z(n34715) );
  XOR U34861 ( .A(n34716), .B(n34715), .Z(n34554) );
  NANDN U34862 ( .A(n34384), .B(n34383), .Z(n34388) );
  NAND U34863 ( .A(n34386), .B(n34385), .Z(n34387) );
  NAND U34864 ( .A(n34388), .B(n34387), .Z(n34555) );
  XNOR U34865 ( .A(n34554), .B(n34555), .Z(n34556) );
  NANDN U34866 ( .A(n34390), .B(n34389), .Z(n34394) );
  NANDN U34867 ( .A(n34392), .B(n34391), .Z(n34393) );
  NAND U34868 ( .A(n34394), .B(n34393), .Z(n34563) );
  NANDN U34869 ( .A(n34396), .B(n34395), .Z(n34400) );
  NAND U34870 ( .A(n34398), .B(n34397), .Z(n34399) );
  NAND U34871 ( .A(n34400), .B(n34399), .Z(n34586) );
  XOR U34872 ( .A(a[116]), .B(n975), .Z(n34692) );
  NANDN U34873 ( .A(n34692), .B(n36311), .Z(n34403) );
  NANDN U34874 ( .A(n34401), .B(n36309), .Z(n34402) );
  NAND U34875 ( .A(n34403), .B(n34402), .Z(n34639) );
  XOR U34876 ( .A(b[53]), .B(n36100), .Z(n34686) );
  NANDN U34877 ( .A(n34686), .B(n37940), .Z(n34406) );
  NANDN U34878 ( .A(n34404), .B(n37941), .Z(n34405) );
  NAND U34879 ( .A(n34406), .B(n34405), .Z(n34636) );
  XOR U34880 ( .A(b[55]), .B(n35783), .Z(n34611) );
  NANDN U34881 ( .A(n34611), .B(n38075), .Z(n34409) );
  NANDN U34882 ( .A(n34407), .B(n38073), .Z(n34408) );
  AND U34883 ( .A(n34409), .B(n34408), .Z(n34637) );
  XNOR U34884 ( .A(n34636), .B(n34637), .Z(n34638) );
  XNOR U34885 ( .A(n34639), .B(n34638), .Z(n34584) );
  NAND U34886 ( .A(n37469), .B(n34410), .Z(n34412) );
  XOR U34887 ( .A(b[47]), .B(n36909), .Z(n34621) );
  NANDN U34888 ( .A(n34621), .B(n37471), .Z(n34411) );
  NAND U34889 ( .A(n34412), .B(n34411), .Z(n34599) );
  XOR U34890 ( .A(b[61]), .B(n34852), .Z(n34642) );
  OR U34891 ( .A(n34642), .B(n38371), .Z(n34415) );
  NANDN U34892 ( .A(n34413), .B(n38369), .Z(n34414) );
  NAND U34893 ( .A(n34415), .B(n34414), .Z(n34596) );
  NAND U34894 ( .A(n34848), .B(n34416), .Z(n34418) );
  XOR U34895 ( .A(a[126]), .B(n35375), .Z(n34617) );
  NANDN U34896 ( .A(n34617), .B(n34618), .Z(n34417) );
  AND U34897 ( .A(n34418), .B(n34417), .Z(n34597) );
  XNOR U34898 ( .A(n34596), .B(n34597), .Z(n34598) );
  XOR U34899 ( .A(n34599), .B(n34598), .Z(n34585) );
  XOR U34900 ( .A(n34584), .B(n34585), .Z(n34587) );
  XNOR U34901 ( .A(n34586), .B(n34587), .Z(n34575) );
  NANDN U34902 ( .A(n34420), .B(n34419), .Z(n34424) );
  NAND U34903 ( .A(n34422), .B(n34421), .Z(n34423) );
  NAND U34904 ( .A(n34424), .B(n34423), .Z(n34632) );
  XOR U34905 ( .A(b[51]), .B(n36420), .Z(n34648) );
  NANDN U34906 ( .A(n34648), .B(n37803), .Z(n34427) );
  NANDN U34907 ( .A(n34425), .B(n37802), .Z(n34426) );
  NAND U34908 ( .A(n34427), .B(n34426), .Z(n34605) );
  XNOR U34909 ( .A(a[118]), .B(b[35]), .Z(n34608) );
  NANDN U34910 ( .A(n34608), .B(n35985), .Z(n34430) );
  NAND U34911 ( .A(n34428), .B(n35986), .Z(n34429) );
  NAND U34912 ( .A(n34430), .B(n34429), .Z(n34602) );
  XOR U34913 ( .A(a[120]), .B(n974), .Z(n34651) );
  NANDN U34914 ( .A(n34651), .B(n35620), .Z(n34433) );
  NANDN U34915 ( .A(n34431), .B(n35621), .Z(n34432) );
  AND U34916 ( .A(n34433), .B(n34432), .Z(n34603) );
  XNOR U34917 ( .A(n34602), .B(n34603), .Z(n34604) );
  XNOR U34918 ( .A(n34605), .B(n34604), .Z(n34630) );
  XOR U34919 ( .A(b[57]), .B(n35545), .Z(n34614) );
  OR U34920 ( .A(n34614), .B(n965), .Z(n34436) );
  NANDN U34921 ( .A(n34434), .B(n38194), .Z(n34435) );
  NAND U34922 ( .A(n34436), .B(n34435), .Z(n34669) );
  NAND U34923 ( .A(n38326), .B(n34437), .Z(n34439) );
  XOR U34924 ( .A(n38400), .B(n35191), .Z(n34654) );
  NANDN U34925 ( .A(n38273), .B(n34654), .Z(n34438) );
  NAND U34926 ( .A(n34439), .B(n34438), .Z(n34666) );
  XNOR U34927 ( .A(b[45]), .B(a[108]), .Z(n34657) );
  NANDN U34928 ( .A(n34657), .B(n37261), .Z(n34442) );
  NAND U34929 ( .A(n34440), .B(n37262), .Z(n34441) );
  AND U34930 ( .A(n34442), .B(n34441), .Z(n34667) );
  XNOR U34931 ( .A(n34666), .B(n34667), .Z(n34668) );
  XOR U34932 ( .A(n34669), .B(n34668), .Z(n34631) );
  XOR U34933 ( .A(n34630), .B(n34631), .Z(n34633) );
  XNOR U34934 ( .A(n34632), .B(n34633), .Z(n34572) );
  NANDN U34935 ( .A(n34444), .B(n34443), .Z(n34448) );
  NAND U34936 ( .A(n34446), .B(n34445), .Z(n34447) );
  AND U34937 ( .A(n34448), .B(n34447), .Z(n34573) );
  XNOR U34938 ( .A(n34572), .B(n34573), .Z(n34574) );
  XNOR U34939 ( .A(n34575), .B(n34574), .Z(n34627) );
  NANDN U34940 ( .A(n34450), .B(n34449), .Z(n34454) );
  NAND U34941 ( .A(n34452), .B(n34451), .Z(n34453) );
  NAND U34942 ( .A(n34454), .B(n34453), .Z(n34624) );
  NANDN U34943 ( .A(n34456), .B(n34455), .Z(n34460) );
  OR U34944 ( .A(n34458), .B(n34457), .Z(n34459) );
  AND U34945 ( .A(n34460), .B(n34459), .Z(n34625) );
  XNOR U34946 ( .A(n34624), .B(n34625), .Z(n34626) );
  XOR U34947 ( .A(n34627), .B(n34626), .Z(n34560) );
  NANDN U34948 ( .A(n34462), .B(n34461), .Z(n34466) );
  NAND U34949 ( .A(n34464), .B(n34463), .Z(n34465) );
  NAND U34950 ( .A(n34466), .B(n34465), .Z(n34579) );
  NAND U34951 ( .A(n34468), .B(n34467), .Z(n34472) );
  OR U34952 ( .A(n34470), .B(n34469), .Z(n34471) );
  AND U34953 ( .A(n34472), .B(n34471), .Z(n34701) );
  XOR U34954 ( .A(n37336), .B(n977), .Z(n34698) );
  NAND U34955 ( .A(n34698), .B(n37068), .Z(n34475) );
  NANDN U34956 ( .A(n34473), .B(n37069), .Z(n34474) );
  NAND U34957 ( .A(n34475), .B(n34474), .Z(n34593) );
  XNOR U34958 ( .A(n37583), .B(b[41]), .Z(n34695) );
  NANDN U34959 ( .A(n36905), .B(n34695), .Z(n34478) );
  NAND U34960 ( .A(n34476), .B(n36807), .Z(n34477) );
  NAND U34961 ( .A(n34478), .B(n34477), .Z(n34590) );
  XOR U34962 ( .A(a[114]), .B(n976), .Z(n34689) );
  NANDN U34963 ( .A(n34689), .B(n36553), .Z(n34481) );
  NANDN U34964 ( .A(n34479), .B(n36643), .Z(n34480) );
  AND U34965 ( .A(n34481), .B(n34480), .Z(n34591) );
  XNOR U34966 ( .A(n34590), .B(n34591), .Z(n34592) );
  XNOR U34967 ( .A(n34593), .B(n34592), .Z(n34702) );
  XNOR U34968 ( .A(n34701), .B(n34702), .Z(n34703) );
  NANDN U34969 ( .A(n34483), .B(n34482), .Z(n34487) );
  NAND U34970 ( .A(n34485), .B(n34484), .Z(n34486) );
  AND U34971 ( .A(n34487), .B(n34486), .Z(n34704) );
  XOR U34972 ( .A(n34703), .B(n34704), .Z(n34578) );
  XNOR U34973 ( .A(n34579), .B(n34578), .Z(n34581) );
  NANDN U34974 ( .A(n34489), .B(n34488), .Z(n34493) );
  NAND U34975 ( .A(n34491), .B(n34490), .Z(n34492) );
  NAND U34976 ( .A(n34493), .B(n34492), .Z(n34580) );
  XNOR U34977 ( .A(n34581), .B(n34580), .Z(n34569) );
  NANDN U34978 ( .A(n34495), .B(n34494), .Z(n34499) );
  OR U34979 ( .A(n34497), .B(n34496), .Z(n34498) );
  NAND U34980 ( .A(n34499), .B(n34498), .Z(n34566) );
  NANDN U34981 ( .A(n34501), .B(n34500), .Z(n34505) );
  NAND U34982 ( .A(n34503), .B(n34502), .Z(n34504) );
  NAND U34983 ( .A(n34505), .B(n34504), .Z(n34710) );
  XOR U34984 ( .A(b[63]), .B(n34851), .Z(n34678) );
  NANDN U34985 ( .A(n34678), .B(n38422), .Z(n34508) );
  NANDN U34986 ( .A(n34506), .B(n38423), .Z(n34507) );
  NAND U34987 ( .A(n34508), .B(n34507), .Z(n34682) );
  XNOR U34988 ( .A(b[25]), .B(n34509), .Z(n34514) );
  XOR U34989 ( .A(n34510), .B(b[24]), .Z(n34512) );
  NAND U34990 ( .A(n34512), .B(n34511), .Z(n34513) );
  AND U34991 ( .A(n34514), .B(n34513), .Z(n34681) );
  AND U34992 ( .A(b[63]), .B(a[88]), .Z(n34816) );
  XOR U34993 ( .A(n34681), .B(n34816), .Z(n34683) );
  XNOR U34994 ( .A(n34682), .B(n34683), .Z(n34708) );
  XOR U34995 ( .A(b[49]), .B(n36647), .Z(n34672) );
  OR U34996 ( .A(n34672), .B(n37756), .Z(n34517) );
  NANDN U34997 ( .A(n34515), .B(n37652), .Z(n34516) );
  NAND U34998 ( .A(n34517), .B(n34516), .Z(n34663) );
  XOR U34999 ( .A(a[122]), .B(n973), .Z(n34645) );
  NANDN U35000 ( .A(n34645), .B(n35313), .Z(n34520) );
  NANDN U35001 ( .A(n34518), .B(n35311), .Z(n34519) );
  NAND U35002 ( .A(n34520), .B(n34519), .Z(n34660) );
  NAND U35003 ( .A(n35188), .B(n34521), .Z(n34523) );
  XOR U35004 ( .A(n38321), .B(n35540), .Z(n34675) );
  NANDN U35005 ( .A(n34968), .B(n34675), .Z(n34522) );
  AND U35006 ( .A(n34523), .B(n34522), .Z(n34661) );
  XNOR U35007 ( .A(n34660), .B(n34661), .Z(n34662) );
  XNOR U35008 ( .A(n34663), .B(n34662), .Z(n34707) );
  XOR U35009 ( .A(n34708), .B(n34707), .Z(n34709) );
  XNOR U35010 ( .A(n34710), .B(n34709), .Z(n34567) );
  XNOR U35011 ( .A(n34566), .B(n34567), .Z(n34568) );
  XOR U35012 ( .A(n34569), .B(n34568), .Z(n34561) );
  XOR U35013 ( .A(n34560), .B(n34561), .Z(n34562) );
  XOR U35014 ( .A(n34563), .B(n34562), .Z(n34557) );
  XNOR U35015 ( .A(n34556), .B(n34557), .Z(n34548) );
  XOR U35016 ( .A(n34549), .B(n34548), .Z(n34551) );
  NAND U35017 ( .A(n34525), .B(n34524), .Z(n34529) );
  OR U35018 ( .A(n34527), .B(n34526), .Z(n34528) );
  NAND U35019 ( .A(n34529), .B(n34528), .Z(n34550) );
  XNOR U35020 ( .A(n34551), .B(n34550), .Z(n34722) );
  NANDN U35021 ( .A(n34535), .B(n34534), .Z(n34539) );
  NANDN U35022 ( .A(n34537), .B(n34536), .Z(n34538) );
  NAND U35023 ( .A(n34539), .B(n34538), .Z(n34720) );
  XNOR U35024 ( .A(n34719), .B(n34720), .Z(n34721) );
  XOR U35025 ( .A(n34722), .B(n34721), .Z(n34543) );
  IV U35026 ( .A(n34543), .Z(n34541) );
  XOR U35027 ( .A(n34542), .B(n34541), .Z(n34540) );
  XNOR U35028 ( .A(n34545), .B(n34540), .Z(n34725) );
  XOR U35029 ( .A(n34726), .B(n34725), .Z(c[216]) );
  NANDN U35030 ( .A(n34541), .B(n34542), .Z(n34547) );
  NOR U35031 ( .A(n34543), .B(n34542), .Z(n34544) );
  OR U35032 ( .A(n34545), .B(n34544), .Z(n34546) );
  NAND U35033 ( .A(n34547), .B(n34546), .Z(n34731) );
  NANDN U35034 ( .A(n34549), .B(n34548), .Z(n34553) );
  OR U35035 ( .A(n34551), .B(n34550), .Z(n34552) );
  NAND U35036 ( .A(n34553), .B(n34552), .Z(n34910) );
  NANDN U35037 ( .A(n34555), .B(n34554), .Z(n34559) );
  NANDN U35038 ( .A(n34557), .B(n34556), .Z(n34558) );
  NAND U35039 ( .A(n34559), .B(n34558), .Z(n34907) );
  NAND U35040 ( .A(n34561), .B(n34560), .Z(n34565) );
  NANDN U35041 ( .A(n34563), .B(n34562), .Z(n34564) );
  NAND U35042 ( .A(n34565), .B(n34564), .Z(n34901) );
  NANDN U35043 ( .A(n34567), .B(n34566), .Z(n34571) );
  NAND U35044 ( .A(n34569), .B(n34568), .Z(n34570) );
  NAND U35045 ( .A(n34571), .B(n34570), .Z(n34738) );
  NANDN U35046 ( .A(n34573), .B(n34572), .Z(n34577) );
  NAND U35047 ( .A(n34575), .B(n34574), .Z(n34576) );
  NAND U35048 ( .A(n34577), .B(n34576), .Z(n34735) );
  NAND U35049 ( .A(n34579), .B(n34578), .Z(n34583) );
  OR U35050 ( .A(n34581), .B(n34580), .Z(n34582) );
  NAND U35051 ( .A(n34583), .B(n34582), .Z(n34880) );
  NANDN U35052 ( .A(n34585), .B(n34584), .Z(n34589) );
  OR U35053 ( .A(n34587), .B(n34586), .Z(n34588) );
  NAND U35054 ( .A(n34589), .B(n34588), .Z(n34878) );
  NANDN U35055 ( .A(n34591), .B(n34590), .Z(n34595) );
  NAND U35056 ( .A(n34593), .B(n34592), .Z(n34594) );
  NAND U35057 ( .A(n34595), .B(n34594), .Z(n34872) );
  NANDN U35058 ( .A(n34597), .B(n34596), .Z(n34601) );
  NAND U35059 ( .A(n34599), .B(n34598), .Z(n34600) );
  AND U35060 ( .A(n34601), .B(n34600), .Z(n34871) );
  XNOR U35061 ( .A(n34872), .B(n34871), .Z(n34873) );
  NANDN U35062 ( .A(n34603), .B(n34602), .Z(n34607) );
  NAND U35063 ( .A(n34605), .B(n34604), .Z(n34606) );
  NAND U35064 ( .A(n34607), .B(n34606), .Z(n34804) );
  XNOR U35065 ( .A(a[119]), .B(b[35]), .Z(n34762) );
  NANDN U35066 ( .A(n34762), .B(n35985), .Z(n34610) );
  NANDN U35067 ( .A(n34608), .B(n35986), .Z(n34609) );
  NAND U35068 ( .A(n34610), .B(n34609), .Z(n34811) );
  XNOR U35069 ( .A(b[55]), .B(a[99]), .Z(n34820) );
  NANDN U35070 ( .A(n34820), .B(n38075), .Z(n34613) );
  NANDN U35071 ( .A(n34611), .B(n38073), .Z(n34612) );
  NAND U35072 ( .A(n34613), .B(n34612), .Z(n34808) );
  XNOR U35073 ( .A(b[57]), .B(a[97]), .Z(n34823) );
  OR U35074 ( .A(n34823), .B(n965), .Z(n34616) );
  NANDN U35075 ( .A(n34614), .B(n38194), .Z(n34615) );
  AND U35076 ( .A(n34616), .B(n34615), .Z(n34809) );
  XNOR U35077 ( .A(n34808), .B(n34809), .Z(n34810) );
  XNOR U35078 ( .A(n34811), .B(n34810), .Z(n34802) );
  NANDN U35079 ( .A(n985), .B(a[89]), .Z(n34815) );
  XOR U35080 ( .A(n34814), .B(n34815), .Z(n34817) );
  XNOR U35081 ( .A(n34816), .B(n34817), .Z(n34741) );
  NANDN U35082 ( .A(n34617), .B(n34848), .Z(n34620) );
  XOR U35083 ( .A(n38463), .B(n35375), .Z(n34847) );
  NAND U35084 ( .A(n34618), .B(n34847), .Z(n34619) );
  NAND U35085 ( .A(n34620), .B(n34619), .Z(n34742) );
  XOR U35086 ( .A(n34741), .B(n34742), .Z(n34743) );
  NANDN U35087 ( .A(n34621), .B(n37469), .Z(n34623) );
  XNOR U35088 ( .A(n978), .B(a[107]), .Z(n34856) );
  NAND U35089 ( .A(n34856), .B(n37471), .Z(n34622) );
  AND U35090 ( .A(n34623), .B(n34622), .Z(n34744) );
  XNOR U35091 ( .A(n34743), .B(n34744), .Z(n34803) );
  XOR U35092 ( .A(n34802), .B(n34803), .Z(n34805) );
  XOR U35093 ( .A(n34804), .B(n34805), .Z(n34874) );
  XOR U35094 ( .A(n34873), .B(n34874), .Z(n34877) );
  XOR U35095 ( .A(n34878), .B(n34877), .Z(n34879) );
  XOR U35096 ( .A(n34880), .B(n34879), .Z(n34736) );
  XOR U35097 ( .A(n34735), .B(n34736), .Z(n34737) );
  XNOR U35098 ( .A(n34738), .B(n34737), .Z(n34898) );
  NANDN U35099 ( .A(n34625), .B(n34624), .Z(n34629) );
  NAND U35100 ( .A(n34627), .B(n34626), .Z(n34628) );
  NAND U35101 ( .A(n34629), .B(n34628), .Z(n34896) );
  NANDN U35102 ( .A(n34631), .B(n34630), .Z(n34635) );
  OR U35103 ( .A(n34633), .B(n34632), .Z(n34634) );
  NAND U35104 ( .A(n34635), .B(n34634), .Z(n34886) );
  NANDN U35105 ( .A(n34637), .B(n34636), .Z(n34641) );
  NAND U35106 ( .A(n34639), .B(n34638), .Z(n34640) );
  NAND U35107 ( .A(n34641), .B(n34640), .Z(n34798) );
  XOR U35108 ( .A(b[61]), .B(n35377), .Z(n34862) );
  OR U35109 ( .A(n34862), .B(n38371), .Z(n34644) );
  NANDN U35110 ( .A(n34642), .B(n38369), .Z(n34643) );
  NAND U35111 ( .A(n34644), .B(n34643), .Z(n34832) );
  XNOR U35112 ( .A(a[123]), .B(b[31]), .Z(n34753) );
  NANDN U35113 ( .A(n34753), .B(n35313), .Z(n34647) );
  NANDN U35114 ( .A(n34645), .B(n35311), .Z(n34646) );
  NAND U35115 ( .A(n34647), .B(n34646), .Z(n34829) );
  XNOR U35116 ( .A(b[51]), .B(a[103]), .Z(n34768) );
  NANDN U35117 ( .A(n34768), .B(n37803), .Z(n34650) );
  NANDN U35118 ( .A(n34648), .B(n37802), .Z(n34649) );
  AND U35119 ( .A(n34650), .B(n34649), .Z(n34830) );
  XNOR U35120 ( .A(n34829), .B(n34830), .Z(n34831) );
  XNOR U35121 ( .A(n34832), .B(n34831), .Z(n34796) );
  XNOR U35122 ( .A(a[121]), .B(b[33]), .Z(n34765) );
  NANDN U35123 ( .A(n34765), .B(n35620), .Z(n34653) );
  NANDN U35124 ( .A(n34651), .B(n35621), .Z(n34652) );
  NAND U35125 ( .A(n34653), .B(n34652), .Z(n34750) );
  NAND U35126 ( .A(n38326), .B(n34654), .Z(n34656) );
  XOR U35127 ( .A(n38400), .B(n35628), .Z(n34756) );
  NANDN U35128 ( .A(n38273), .B(n34756), .Z(n34655) );
  NAND U35129 ( .A(n34656), .B(n34655), .Z(n34747) );
  XOR U35130 ( .A(b[45]), .B(a[109]), .Z(n34826) );
  NAND U35131 ( .A(n34826), .B(n37261), .Z(n34659) );
  NANDN U35132 ( .A(n34657), .B(n37262), .Z(n34658) );
  AND U35133 ( .A(n34659), .B(n34658), .Z(n34748) );
  XNOR U35134 ( .A(n34747), .B(n34748), .Z(n34749) );
  XOR U35135 ( .A(n34750), .B(n34749), .Z(n34797) );
  XOR U35136 ( .A(n34796), .B(n34797), .Z(n34799) );
  XNOR U35137 ( .A(n34798), .B(n34799), .Z(n34793) );
  NANDN U35138 ( .A(n34661), .B(n34660), .Z(n34665) );
  NAND U35139 ( .A(n34663), .B(n34662), .Z(n34664) );
  NAND U35140 ( .A(n34665), .B(n34664), .Z(n34790) );
  NANDN U35141 ( .A(n34667), .B(n34666), .Z(n34671) );
  NAND U35142 ( .A(n34669), .B(n34668), .Z(n34670) );
  AND U35143 ( .A(n34671), .B(n34670), .Z(n34791) );
  XNOR U35144 ( .A(n34790), .B(n34791), .Z(n34792) );
  XNOR U35145 ( .A(n34793), .B(n34792), .Z(n34884) );
  XNOR U35146 ( .A(b[49]), .B(a[105]), .Z(n34759) );
  OR U35147 ( .A(n34759), .B(n37756), .Z(n34674) );
  NANDN U35148 ( .A(n34672), .B(n37652), .Z(n34673) );
  NAND U35149 ( .A(n34674), .B(n34673), .Z(n34838) );
  NAND U35150 ( .A(n35188), .B(n34675), .Z(n34677) );
  XNOR U35151 ( .A(a[125]), .B(n35540), .Z(n34859) );
  NANDN U35152 ( .A(n34968), .B(n34859), .Z(n34676) );
  NAND U35153 ( .A(n34677), .B(n34676), .Z(n34835) );
  XNOR U35154 ( .A(b[63]), .B(a[91]), .Z(n34853) );
  NANDN U35155 ( .A(n34853), .B(n38422), .Z(n34680) );
  NANDN U35156 ( .A(n34678), .B(n38423), .Z(n34679) );
  AND U35157 ( .A(n34680), .B(n34679), .Z(n34836) );
  XNOR U35158 ( .A(n34835), .B(n34836), .Z(n34837) );
  XNOR U35159 ( .A(n34838), .B(n34837), .Z(n34789) );
  NANDN U35160 ( .A(n34816), .B(n34681), .Z(n34685) );
  NANDN U35161 ( .A(n34683), .B(n34682), .Z(n34684) );
  NAND U35162 ( .A(n34685), .B(n34684), .Z(n34787) );
  XNOR U35163 ( .A(b[53]), .B(a[101]), .Z(n34771) );
  NANDN U35164 ( .A(n34771), .B(n37940), .Z(n34688) );
  NANDN U35165 ( .A(n34686), .B(n37941), .Z(n34687) );
  AND U35166 ( .A(n34688), .B(n34687), .Z(n34865) );
  XNOR U35167 ( .A(a[115]), .B(n976), .Z(n34783) );
  NAND U35168 ( .A(n34783), .B(n36553), .Z(n34691) );
  NANDN U35169 ( .A(n34689), .B(n36643), .Z(n34690) );
  AND U35170 ( .A(n34691), .B(n34690), .Z(n34866) );
  XNOR U35171 ( .A(a[117]), .B(b[37]), .Z(n34777) );
  NANDN U35172 ( .A(n34777), .B(n36311), .Z(n34694) );
  NANDN U35173 ( .A(n34692), .B(n36309), .Z(n34693) );
  AND U35174 ( .A(n34694), .B(n34693), .Z(n34868) );
  XOR U35175 ( .A(n34867), .B(n34868), .Z(n34844) );
  NAND U35176 ( .A(n36807), .B(n34695), .Z(n34697) );
  XOR U35177 ( .A(a[113]), .B(b[41]), .Z(n34780) );
  NANDN U35178 ( .A(n36905), .B(n34780), .Z(n34696) );
  NAND U35179 ( .A(n34697), .B(n34696), .Z(n34842) );
  NAND U35180 ( .A(n37069), .B(n34698), .Z(n34700) );
  XNOR U35181 ( .A(a[111]), .B(n977), .Z(n34774) );
  NAND U35182 ( .A(n34774), .B(n37068), .Z(n34699) );
  AND U35183 ( .A(n34700), .B(n34699), .Z(n34841) );
  XNOR U35184 ( .A(n34842), .B(n34841), .Z(n34843) );
  XOR U35185 ( .A(n34844), .B(n34843), .Z(n34786) );
  XNOR U35186 ( .A(n34787), .B(n34786), .Z(n34788) );
  XOR U35187 ( .A(n34789), .B(n34788), .Z(n34883) );
  XOR U35188 ( .A(n34884), .B(n34883), .Z(n34885) );
  XNOR U35189 ( .A(n34886), .B(n34885), .Z(n34892) );
  OR U35190 ( .A(n34702), .B(n34701), .Z(n34706) );
  OR U35191 ( .A(n34704), .B(n34703), .Z(n34705) );
  NAND U35192 ( .A(n34706), .B(n34705), .Z(n34889) );
  NANDN U35193 ( .A(n34708), .B(n34707), .Z(n34712) );
  OR U35194 ( .A(n34710), .B(n34709), .Z(n34711) );
  NAND U35195 ( .A(n34712), .B(n34711), .Z(n34890) );
  XNOR U35196 ( .A(n34889), .B(n34890), .Z(n34891) );
  XOR U35197 ( .A(n34892), .B(n34891), .Z(n34895) );
  XNOR U35198 ( .A(n34896), .B(n34895), .Z(n34897) );
  XOR U35199 ( .A(n34898), .B(n34897), .Z(n34902) );
  XNOR U35200 ( .A(n34901), .B(n34902), .Z(n34903) );
  NANDN U35201 ( .A(n34714), .B(n34713), .Z(n34718) );
  NANDN U35202 ( .A(n34716), .B(n34715), .Z(n34717) );
  AND U35203 ( .A(n34718), .B(n34717), .Z(n34904) );
  XNOR U35204 ( .A(n34903), .B(n34904), .Z(n34908) );
  XNOR U35205 ( .A(n34907), .B(n34908), .Z(n34909) );
  XNOR U35206 ( .A(n34910), .B(n34909), .Z(n34729) );
  NANDN U35207 ( .A(n34720), .B(n34719), .Z(n34724) );
  NAND U35208 ( .A(n34722), .B(n34721), .Z(n34723) );
  AND U35209 ( .A(n34724), .B(n34723), .Z(n34730) );
  XOR U35210 ( .A(n34729), .B(n34730), .Z(n34732) );
  XNOR U35211 ( .A(n34731), .B(n34732), .Z(n34727) );
  OR U35212 ( .A(n34726), .B(n34725), .Z(n34728) );
  XNOR U35213 ( .A(n34727), .B(n34728), .Z(c[217]) );
  NANDN U35214 ( .A(n34728), .B(n34727), .Z(n35083) );
  NANDN U35215 ( .A(n34730), .B(n34729), .Z(n34734) );
  NANDN U35216 ( .A(n34732), .B(n34731), .Z(n34733) );
  AND U35217 ( .A(n34734), .B(n34733), .Z(n34918) );
  OR U35218 ( .A(n34736), .B(n34735), .Z(n34740) );
  NAND U35219 ( .A(n34738), .B(n34737), .Z(n34739) );
  NAND U35220 ( .A(n34740), .B(n34739), .Z(n34922) );
  OR U35221 ( .A(n34742), .B(n34741), .Z(n34746) );
  NAND U35222 ( .A(n34744), .B(n34743), .Z(n34745) );
  NAND U35223 ( .A(n34746), .B(n34745), .Z(n34946) );
  NANDN U35224 ( .A(n34748), .B(n34747), .Z(n34752) );
  NAND U35225 ( .A(n34750), .B(n34749), .Z(n34751) );
  NAND U35226 ( .A(n34752), .B(n34751), .Z(n34944) );
  XOR U35227 ( .A(a[124]), .B(n973), .Z(n34964) );
  NANDN U35228 ( .A(n34964), .B(n35313), .Z(n34755) );
  NANDN U35229 ( .A(n34753), .B(n35311), .Z(n34754) );
  NAND U35230 ( .A(n34755), .B(n34754), .Z(n34989) );
  NAND U35231 ( .A(n38326), .B(n34756), .Z(n34758) );
  XOR U35232 ( .A(n38400), .B(n35545), .Z(n34971) );
  NANDN U35233 ( .A(n38273), .B(n34971), .Z(n34757) );
  NAND U35234 ( .A(n34758), .B(n34757), .Z(n34986) );
  XOR U35235 ( .A(b[49]), .B(n36909), .Z(n35013) );
  OR U35236 ( .A(n35013), .B(n37756), .Z(n34761) );
  NANDN U35237 ( .A(n34759), .B(n37652), .Z(n34760) );
  AND U35238 ( .A(n34761), .B(n34760), .Z(n34987) );
  XNOR U35239 ( .A(n34986), .B(n34987), .Z(n34988) );
  XOR U35240 ( .A(n34989), .B(n34988), .Z(n34949) );
  XNOR U35241 ( .A(a[120]), .B(b[35]), .Z(n35010) );
  NANDN U35242 ( .A(n35010), .B(n35985), .Z(n34764) );
  NANDN U35243 ( .A(n34762), .B(n35986), .Z(n34763) );
  NAND U35244 ( .A(n34764), .B(n34763), .Z(n35073) );
  XOR U35245 ( .A(a[122]), .B(n974), .Z(n35067) );
  NANDN U35246 ( .A(n35067), .B(n35620), .Z(n34767) );
  NANDN U35247 ( .A(n34765), .B(n35621), .Z(n34766) );
  NAND U35248 ( .A(n34767), .B(n34766), .Z(n35070) );
  XOR U35249 ( .A(b[51]), .B(n36647), .Z(n34977) );
  NANDN U35250 ( .A(n34977), .B(n37803), .Z(n34770) );
  NANDN U35251 ( .A(n34768), .B(n37802), .Z(n34769) );
  AND U35252 ( .A(n34770), .B(n34769), .Z(n35071) );
  XNOR U35253 ( .A(n35070), .B(n35071), .Z(n35072) );
  XOR U35254 ( .A(n35073), .B(n35072), .Z(n34950) );
  XNOR U35255 ( .A(n34949), .B(n34950), .Z(n34952) );
  XOR U35256 ( .A(b[53]), .B(n36420), .Z(n35016) );
  NANDN U35257 ( .A(n35016), .B(n37940), .Z(n34773) );
  NANDN U35258 ( .A(n34771), .B(n37941), .Z(n34772) );
  AND U35259 ( .A(n34773), .B(n34772), .Z(n35048) );
  XOR U35260 ( .A(a[112]), .B(n977), .Z(n35007) );
  NANDN U35261 ( .A(n35007), .B(n37068), .Z(n34776) );
  NAND U35262 ( .A(n34774), .B(n37069), .Z(n34775) );
  AND U35263 ( .A(n34776), .B(n34775), .Z(n35049) );
  XNOR U35264 ( .A(n35048), .B(n35049), .Z(n35051) );
  XOR U35265 ( .A(a[118]), .B(n975), .Z(n35001) );
  NANDN U35266 ( .A(n35001), .B(n36311), .Z(n34779) );
  NANDN U35267 ( .A(n34777), .B(n36309), .Z(n34778) );
  AND U35268 ( .A(n34779), .B(n34778), .Z(n35050) );
  XNOR U35269 ( .A(n35051), .B(n35050), .Z(n34983) );
  NAND U35270 ( .A(n36807), .B(n34780), .Z(n34782) );
  XNOR U35271 ( .A(n37873), .B(b[41]), .Z(n35004) );
  NANDN U35272 ( .A(n36905), .B(n35004), .Z(n34781) );
  NAND U35273 ( .A(n34782), .B(n34781), .Z(n34981) );
  NAND U35274 ( .A(n36643), .B(n34783), .Z(n34785) );
  XOR U35275 ( .A(n38046), .B(n976), .Z(n34998) );
  NAND U35276 ( .A(n34998), .B(n36553), .Z(n34784) );
  AND U35277 ( .A(n34785), .B(n34784), .Z(n34980) );
  XNOR U35278 ( .A(n34981), .B(n34980), .Z(n34982) );
  XOR U35279 ( .A(n34983), .B(n34982), .Z(n34951) );
  XNOR U35280 ( .A(n34952), .B(n34951), .Z(n34943) );
  XNOR U35281 ( .A(n34944), .B(n34943), .Z(n34945) );
  XNOR U35282 ( .A(n34946), .B(n34945), .Z(n35026) );
  NANDN U35283 ( .A(n34791), .B(n34790), .Z(n34795) );
  NAND U35284 ( .A(n34793), .B(n34792), .Z(n34794) );
  NAND U35285 ( .A(n34795), .B(n34794), .Z(n35024) );
  XNOR U35286 ( .A(n35023), .B(n35024), .Z(n35025) );
  XOR U35287 ( .A(n35026), .B(n35025), .Z(n35022) );
  NANDN U35288 ( .A(n34797), .B(n34796), .Z(n34801) );
  OR U35289 ( .A(n34799), .B(n34798), .Z(n34800) );
  NAND U35290 ( .A(n34801), .B(n34800), .Z(n35029) );
  NANDN U35291 ( .A(n34803), .B(n34802), .Z(n34807) );
  OR U35292 ( .A(n34805), .B(n34804), .Z(n34806) );
  AND U35293 ( .A(n34807), .B(n34806), .Z(n35030) );
  XNOR U35294 ( .A(n35029), .B(n35030), .Z(n35031) );
  NANDN U35295 ( .A(n34809), .B(n34808), .Z(n34813) );
  NAND U35296 ( .A(n34811), .B(n34810), .Z(n34812) );
  NAND U35297 ( .A(n34813), .B(n34812), .Z(n35041) );
  NANDN U35298 ( .A(n34815), .B(n34814), .Z(n34819) );
  NANDN U35299 ( .A(n34817), .B(n34816), .Z(n34818) );
  NAND U35300 ( .A(n34819), .B(n34818), .Z(n35039) );
  XOR U35301 ( .A(b[55]), .B(n36100), .Z(n35061) );
  NANDN U35302 ( .A(n35061), .B(n38075), .Z(n34822) );
  NANDN U35303 ( .A(n34820), .B(n38073), .Z(n34821) );
  NAND U35304 ( .A(n34822), .B(n34821), .Z(n34958) );
  XOR U35305 ( .A(b[57]), .B(n35783), .Z(n35064) );
  OR U35306 ( .A(n35064), .B(n965), .Z(n34825) );
  NANDN U35307 ( .A(n34823), .B(n38194), .Z(n34824) );
  NAND U35308 ( .A(n34825), .B(n34824), .Z(n34955) );
  XNOR U35309 ( .A(b[45]), .B(a[110]), .Z(n34961) );
  NANDN U35310 ( .A(n34961), .B(n37261), .Z(n34828) );
  NAND U35311 ( .A(n34826), .B(n37262), .Z(n34827) );
  AND U35312 ( .A(n34828), .B(n34827), .Z(n34956) );
  XNOR U35313 ( .A(n34955), .B(n34956), .Z(n34957) );
  XNOR U35314 ( .A(n34958), .B(n34957), .Z(n35040) );
  XNOR U35315 ( .A(n35039), .B(n35040), .Z(n35042) );
  XOR U35316 ( .A(n35041), .B(n35042), .Z(n34936) );
  NANDN U35317 ( .A(n34830), .B(n34829), .Z(n34834) );
  NAND U35318 ( .A(n34832), .B(n34831), .Z(n34833) );
  NAND U35319 ( .A(n34834), .B(n34833), .Z(n35035) );
  NANDN U35320 ( .A(n34836), .B(n34835), .Z(n34840) );
  NAND U35321 ( .A(n34838), .B(n34837), .Z(n34839) );
  AND U35322 ( .A(n34840), .B(n34839), .Z(n35036) );
  XNOR U35323 ( .A(n35035), .B(n35036), .Z(n35037) );
  NANDN U35324 ( .A(n34842), .B(n34841), .Z(n34846) );
  NAND U35325 ( .A(n34844), .B(n34843), .Z(n34845) );
  NAND U35326 ( .A(n34846), .B(n34845), .Z(n35038) );
  XNOR U35327 ( .A(n35037), .B(n35038), .Z(n34934) );
  NAND U35328 ( .A(n34848), .B(n34847), .Z(n34850) );
  ANDN U35329 ( .B(n34850), .A(n34849), .Z(n35045) );
  ANDN U35330 ( .B(b[63]), .A(n34851), .Z(n35183) );
  XOR U35331 ( .A(b[63]), .B(n34852), .Z(n35054) );
  NANDN U35332 ( .A(n35054), .B(n38422), .Z(n34855) );
  NANDN U35333 ( .A(n34853), .B(n38423), .Z(n34854) );
  NAND U35334 ( .A(n34855), .B(n34854), .Z(n35043) );
  XNOR U35335 ( .A(n35183), .B(n35043), .Z(n35044) );
  XNOR U35336 ( .A(n35045), .B(n35044), .Z(n34939) );
  NAND U35337 ( .A(n34856), .B(n37469), .Z(n34858) );
  XOR U35338 ( .A(n978), .B(n37139), .Z(n35057) );
  NAND U35339 ( .A(n35057), .B(n37471), .Z(n34857) );
  NAND U35340 ( .A(n34858), .B(n34857), .Z(n34995) );
  NAND U35341 ( .A(n35188), .B(n34859), .Z(n34861) );
  XOR U35342 ( .A(n987), .B(n35540), .Z(n34967) );
  NANDN U35343 ( .A(n34968), .B(n34967), .Z(n34860) );
  NAND U35344 ( .A(n34861), .B(n34860), .Z(n34992) );
  XOR U35345 ( .A(b[61]), .B(n35191), .Z(n34974) );
  OR U35346 ( .A(n34974), .B(n38371), .Z(n34864) );
  NANDN U35347 ( .A(n34862), .B(n38369), .Z(n34863) );
  AND U35348 ( .A(n34864), .B(n34863), .Z(n34993) );
  XNOR U35349 ( .A(n34992), .B(n34993), .Z(n34994) );
  XNOR U35350 ( .A(n34995), .B(n34994), .Z(n34937) );
  OR U35351 ( .A(n34866), .B(n34865), .Z(n34870) );
  NANDN U35352 ( .A(n34868), .B(n34867), .Z(n34869) );
  NAND U35353 ( .A(n34870), .B(n34869), .Z(n34938) );
  XOR U35354 ( .A(n34937), .B(n34938), .Z(n34940) );
  XOR U35355 ( .A(n34939), .B(n34940), .Z(n34933) );
  XNOR U35356 ( .A(n34934), .B(n34933), .Z(n34935) );
  XNOR U35357 ( .A(n34936), .B(n34935), .Z(n35032) );
  XNOR U35358 ( .A(n35031), .B(n35032), .Z(n35019) );
  NANDN U35359 ( .A(n34872), .B(n34871), .Z(n34876) );
  NAND U35360 ( .A(n34874), .B(n34873), .Z(n34875) );
  NAND U35361 ( .A(n34876), .B(n34875), .Z(n35020) );
  XNOR U35362 ( .A(n35019), .B(n35020), .Z(n35021) );
  XNOR U35363 ( .A(n35022), .B(n35021), .Z(n34930) );
  NAND U35364 ( .A(n34878), .B(n34877), .Z(n34882) );
  NANDN U35365 ( .A(n34880), .B(n34879), .Z(n34881) );
  NAND U35366 ( .A(n34882), .B(n34881), .Z(n34927) );
  NAND U35367 ( .A(n34884), .B(n34883), .Z(n34888) );
  NAND U35368 ( .A(n34886), .B(n34885), .Z(n34887) );
  AND U35369 ( .A(n34888), .B(n34887), .Z(n34928) );
  XNOR U35370 ( .A(n34927), .B(n34928), .Z(n34929) );
  XOR U35371 ( .A(n34930), .B(n34929), .Z(n34921) );
  XNOR U35372 ( .A(n34922), .B(n34921), .Z(n34924) );
  NANDN U35373 ( .A(n34890), .B(n34889), .Z(n34894) );
  NAND U35374 ( .A(n34892), .B(n34891), .Z(n34893) );
  NAND U35375 ( .A(n34894), .B(n34893), .Z(n34923) );
  XNOR U35376 ( .A(n34924), .B(n34923), .Z(n35076) );
  NANDN U35377 ( .A(n34896), .B(n34895), .Z(n34900) );
  NAND U35378 ( .A(n34898), .B(n34897), .Z(n34899) );
  AND U35379 ( .A(n34900), .B(n34899), .Z(n35077) );
  XNOR U35380 ( .A(n35076), .B(n35077), .Z(n35078) );
  NANDN U35381 ( .A(n34902), .B(n34901), .Z(n34906) );
  NAND U35382 ( .A(n34904), .B(n34903), .Z(n34905) );
  NAND U35383 ( .A(n34906), .B(n34905), .Z(n35079) );
  XNOR U35384 ( .A(n35078), .B(n35079), .Z(n34916) );
  IV U35385 ( .A(n34916), .Z(n34914) );
  NANDN U35386 ( .A(n34908), .B(n34907), .Z(n34912) );
  NAND U35387 ( .A(n34910), .B(n34909), .Z(n34911) );
  AND U35388 ( .A(n34912), .B(n34911), .Z(n34915) );
  XOR U35389 ( .A(n34914), .B(n34915), .Z(n34913) );
  XNOR U35390 ( .A(n34918), .B(n34913), .Z(n35082) );
  XOR U35391 ( .A(n35083), .B(n35082), .Z(c[218]) );
  NANDN U35392 ( .A(n34914), .B(n34915), .Z(n34920) );
  NOR U35393 ( .A(n34916), .B(n34915), .Z(n34917) );
  OR U35394 ( .A(n34918), .B(n34917), .Z(n34919) );
  NAND U35395 ( .A(n34920), .B(n34919), .Z(n35086) );
  NAND U35396 ( .A(n34922), .B(n34921), .Z(n34926) );
  OR U35397 ( .A(n34924), .B(n34923), .Z(n34925) );
  NAND U35398 ( .A(n34926), .B(n34925), .Z(n35249) );
  NANDN U35399 ( .A(n34928), .B(n34927), .Z(n34932) );
  NAND U35400 ( .A(n34930), .B(n34929), .Z(n34931) );
  NAND U35401 ( .A(n34932), .B(n34931), .Z(n35247) );
  NANDN U35402 ( .A(n34938), .B(n34937), .Z(n34942) );
  OR U35403 ( .A(n34940), .B(n34939), .Z(n34941) );
  NAND U35404 ( .A(n34942), .B(n34941), .Z(n35145) );
  NANDN U35405 ( .A(n34944), .B(n34943), .Z(n34948) );
  NAND U35406 ( .A(n34946), .B(n34945), .Z(n34947) );
  NAND U35407 ( .A(n34948), .B(n34947), .Z(n35143) );
  OR U35408 ( .A(n34950), .B(n34949), .Z(n34954) );
  NANDN U35409 ( .A(n34952), .B(n34951), .Z(n34953) );
  AND U35410 ( .A(n34954), .B(n34953), .Z(n35144) );
  XNOR U35411 ( .A(n35143), .B(n35144), .Z(n35146) );
  XOR U35412 ( .A(n35145), .B(n35146), .Z(n35102) );
  NANDN U35413 ( .A(n34956), .B(n34955), .Z(n34960) );
  NAND U35414 ( .A(n34958), .B(n34957), .Z(n34959) );
  NAND U35415 ( .A(n34960), .B(n34959), .Z(n35242) );
  XOR U35416 ( .A(b[45]), .B(a[111]), .Z(n35159) );
  NAND U35417 ( .A(n35159), .B(n37261), .Z(n34963) );
  NANDN U35418 ( .A(n34961), .B(n37262), .Z(n34962) );
  NAND U35419 ( .A(n34963), .B(n34962), .Z(n35198) );
  XNOR U35420 ( .A(a[125]), .B(b[31]), .Z(n35122) );
  NANDN U35421 ( .A(n35122), .B(n35313), .Z(n34966) );
  NANDN U35422 ( .A(n34964), .B(n35311), .Z(n34965) );
  NAND U35423 ( .A(n34966), .B(n34965), .Z(n35195) );
  NAND U35424 ( .A(n35188), .B(n34967), .Z(n34970) );
  XOR U35425 ( .A(n38463), .B(n35540), .Z(n35187) );
  NANDN U35426 ( .A(n34968), .B(n35187), .Z(n34969) );
  AND U35427 ( .A(n34970), .B(n34969), .Z(n35196) );
  XNOR U35428 ( .A(n35195), .B(n35196), .Z(n35197) );
  XNOR U35429 ( .A(n35198), .B(n35197), .Z(n35240) );
  NAND U35430 ( .A(n38326), .B(n34971), .Z(n34973) );
  XNOR U35431 ( .A(n38400), .B(a[97]), .Z(n35165) );
  NANDN U35432 ( .A(n38273), .B(n35165), .Z(n34972) );
  NAND U35433 ( .A(n34973), .B(n34972), .Z(n35225) );
  XOR U35434 ( .A(b[61]), .B(n35628), .Z(n35168) );
  OR U35435 ( .A(n35168), .B(n38371), .Z(n34976) );
  NANDN U35436 ( .A(n34974), .B(n38369), .Z(n34975) );
  NAND U35437 ( .A(n34976), .B(n34975), .Z(n35222) );
  XNOR U35438 ( .A(b[51]), .B(a[105]), .Z(n35204) );
  NANDN U35439 ( .A(n35204), .B(n37803), .Z(n34979) );
  NANDN U35440 ( .A(n34977), .B(n37802), .Z(n34978) );
  AND U35441 ( .A(n34979), .B(n34978), .Z(n35223) );
  XNOR U35442 ( .A(n35222), .B(n35223), .Z(n35224) );
  XOR U35443 ( .A(n35225), .B(n35224), .Z(n35241) );
  XOR U35444 ( .A(n35240), .B(n35241), .Z(n35243) );
  XOR U35445 ( .A(n35242), .B(n35243), .Z(n35147) );
  NANDN U35446 ( .A(n34981), .B(n34980), .Z(n34985) );
  NAND U35447 ( .A(n34983), .B(n34982), .Z(n34984) );
  NAND U35448 ( .A(n34985), .B(n34984), .Z(n35231) );
  NANDN U35449 ( .A(n34987), .B(n34986), .Z(n34991) );
  NAND U35450 ( .A(n34989), .B(n34988), .Z(n34990) );
  NAND U35451 ( .A(n34991), .B(n34990), .Z(n35229) );
  NANDN U35452 ( .A(n34993), .B(n34992), .Z(n34997) );
  NAND U35453 ( .A(n34995), .B(n34994), .Z(n34996) );
  AND U35454 ( .A(n34997), .B(n34996), .Z(n35228) );
  XNOR U35455 ( .A(n35229), .B(n35228), .Z(n35230) );
  XOR U35456 ( .A(n35231), .B(n35230), .Z(n35148) );
  XOR U35457 ( .A(n35147), .B(n35148), .Z(n35149) );
  NAND U35458 ( .A(n36643), .B(n34998), .Z(n35000) );
  XNOR U35459 ( .A(a[117]), .B(n976), .Z(n35213) );
  NAND U35460 ( .A(n35213), .B(n36553), .Z(n34999) );
  NAND U35461 ( .A(n35000), .B(n34999), .Z(n35113) );
  XOR U35462 ( .A(a[119]), .B(n975), .Z(n35219) );
  NANDN U35463 ( .A(n35219), .B(n36311), .Z(n35003) );
  NANDN U35464 ( .A(n35001), .B(n36309), .Z(n35002) );
  NAND U35465 ( .A(n35003), .B(n35002), .Z(n35119) );
  XOR U35466 ( .A(a[115]), .B(b[41]), .Z(n35216) );
  NANDN U35467 ( .A(n36905), .B(n35216), .Z(n35006) );
  NAND U35468 ( .A(n35004), .B(n36807), .Z(n35005) );
  NAND U35469 ( .A(n35006), .B(n35005), .Z(n35116) );
  XNOR U35470 ( .A(a[113]), .B(b[43]), .Z(n35201) );
  NANDN U35471 ( .A(n35201), .B(n37068), .Z(n35009) );
  NANDN U35472 ( .A(n35007), .B(n37069), .Z(n35008) );
  AND U35473 ( .A(n35009), .B(n35008), .Z(n35117) );
  XNOR U35474 ( .A(n35116), .B(n35117), .Z(n35118) );
  XNOR U35475 ( .A(n35119), .B(n35118), .Z(n35112) );
  XNOR U35476 ( .A(n35113), .B(n35112), .Z(n35115) );
  XOR U35477 ( .A(a[121]), .B(b[35]), .Z(n35210) );
  NAND U35478 ( .A(n35985), .B(n35210), .Z(n35012) );
  NANDN U35479 ( .A(n35010), .B(n35986), .Z(n35011) );
  NAND U35480 ( .A(n35012), .B(n35011), .Z(n35180) );
  XNOR U35481 ( .A(b[49]), .B(a[107]), .Z(n35162) );
  OR U35482 ( .A(n35162), .B(n37756), .Z(n35015) );
  NANDN U35483 ( .A(n35013), .B(n37652), .Z(n35014) );
  NAND U35484 ( .A(n35015), .B(n35014), .Z(n35177) );
  XNOR U35485 ( .A(b[53]), .B(a[103]), .Z(n35153) );
  NANDN U35486 ( .A(n35153), .B(n37940), .Z(n35018) );
  NANDN U35487 ( .A(n35016), .B(n37941), .Z(n35017) );
  AND U35488 ( .A(n35018), .B(n35017), .Z(n35178) );
  XNOR U35489 ( .A(n35177), .B(n35178), .Z(n35179) );
  XNOR U35490 ( .A(n35180), .B(n35179), .Z(n35114) );
  XNOR U35491 ( .A(n35115), .B(n35114), .Z(n35150) );
  XNOR U35492 ( .A(n35149), .B(n35150), .Z(n35103) );
  XOR U35493 ( .A(n35102), .B(n35103), .Z(n35104) );
  XNOR U35494 ( .A(n35105), .B(n35104), .Z(n35092) );
  NANDN U35495 ( .A(n35024), .B(n35023), .Z(n35028) );
  NANDN U35496 ( .A(n35026), .B(n35025), .Z(n35027) );
  NAND U35497 ( .A(n35028), .B(n35027), .Z(n35098) );
  NANDN U35498 ( .A(n35030), .B(n35029), .Z(n35034) );
  NAND U35499 ( .A(n35032), .B(n35031), .Z(n35033) );
  NAND U35500 ( .A(n35034), .B(n35033), .Z(n35097) );
  NANDN U35501 ( .A(n35183), .B(n35043), .Z(n35047) );
  NANDN U35502 ( .A(n35045), .B(n35044), .Z(n35046) );
  NAND U35503 ( .A(n35047), .B(n35046), .Z(n35109) );
  OR U35504 ( .A(n35049), .B(n35048), .Z(n35053) );
  OR U35505 ( .A(n35051), .B(n35050), .Z(n35052) );
  NAND U35506 ( .A(n35053), .B(n35052), .Z(n35236) );
  XOR U35507 ( .A(b[63]), .B(n35377), .Z(n35192) );
  NANDN U35508 ( .A(n35192), .B(n38422), .Z(n35056) );
  NANDN U35509 ( .A(n35054), .B(n38423), .Z(n35055) );
  NAND U35510 ( .A(n35056), .B(n35055), .Z(n35131) );
  NAND U35511 ( .A(n37469), .B(n35057), .Z(n35059) );
  XNOR U35512 ( .A(n978), .B(a[109]), .Z(n35128) );
  NAND U35513 ( .A(n35128), .B(n37471), .Z(n35058) );
  AND U35514 ( .A(n35059), .B(n35058), .Z(n35132) );
  XNOR U35515 ( .A(n35131), .B(n35132), .Z(n35133) );
  NANDN U35516 ( .A(n985), .B(a[91]), .Z(n35186) );
  NAND U35517 ( .A(b[26]), .B(b[25]), .Z(n35060) );
  AND U35518 ( .A(n35060), .B(b[27]), .Z(n35184) );
  XOR U35519 ( .A(n35183), .B(n35184), .Z(n35185) );
  XOR U35520 ( .A(n35186), .B(n35185), .Z(n35134) );
  XOR U35521 ( .A(n35133), .B(n35134), .Z(n35234) );
  XNOR U35522 ( .A(b[55]), .B(a[101]), .Z(n35156) );
  NANDN U35523 ( .A(n35156), .B(n38075), .Z(n35063) );
  NANDN U35524 ( .A(n35061), .B(n38073), .Z(n35062) );
  NAND U35525 ( .A(n35063), .B(n35062), .Z(n35174) );
  XNOR U35526 ( .A(b[57]), .B(a[99]), .Z(n35125) );
  OR U35527 ( .A(n35125), .B(n965), .Z(n35066) );
  NANDN U35528 ( .A(n35064), .B(n38194), .Z(n35065) );
  NAND U35529 ( .A(n35066), .B(n35065), .Z(n35171) );
  XNOR U35530 ( .A(a[123]), .B(b[33]), .Z(n35207) );
  NANDN U35531 ( .A(n35207), .B(n35620), .Z(n35069) );
  NANDN U35532 ( .A(n35067), .B(n35621), .Z(n35068) );
  AND U35533 ( .A(n35069), .B(n35068), .Z(n35172) );
  XNOR U35534 ( .A(n35171), .B(n35172), .Z(n35173) );
  XNOR U35535 ( .A(n35174), .B(n35173), .Z(n35235) );
  XOR U35536 ( .A(n35234), .B(n35235), .Z(n35237) );
  XNOR U35537 ( .A(n35236), .B(n35237), .Z(n35106) );
  NANDN U35538 ( .A(n35071), .B(n35070), .Z(n35075) );
  NAND U35539 ( .A(n35073), .B(n35072), .Z(n35074) );
  NAND U35540 ( .A(n35075), .B(n35074), .Z(n35107) );
  XOR U35541 ( .A(n35106), .B(n35107), .Z(n35108) );
  XOR U35542 ( .A(n35109), .B(n35108), .Z(n35138) );
  XOR U35543 ( .A(n35137), .B(n35138), .Z(n35139) );
  XNOR U35544 ( .A(n35140), .B(n35139), .Z(n35096) );
  XNOR U35545 ( .A(n35097), .B(n35096), .Z(n35099) );
  XNOR U35546 ( .A(n35098), .B(n35099), .Z(n35090) );
  XOR U35547 ( .A(n35091), .B(n35090), .Z(n35093) );
  XOR U35548 ( .A(n35092), .B(n35093), .Z(n35246) );
  XOR U35549 ( .A(n35247), .B(n35246), .Z(n35248) );
  XNOR U35550 ( .A(n35249), .B(n35248), .Z(n35084) );
  NANDN U35551 ( .A(n35077), .B(n35076), .Z(n35081) );
  NANDN U35552 ( .A(n35079), .B(n35078), .Z(n35080) );
  AND U35553 ( .A(n35081), .B(n35080), .Z(n35085) );
  XOR U35554 ( .A(n35084), .B(n35085), .Z(n35087) );
  XNOR U35555 ( .A(n35086), .B(n35087), .Z(n35252) );
  OR U35556 ( .A(n35083), .B(n35082), .Z(n35253) );
  XNOR U35557 ( .A(n35252), .B(n35253), .Z(c[219]) );
  NANDN U35558 ( .A(n35085), .B(n35084), .Z(n35089) );
  NANDN U35559 ( .A(n35087), .B(n35086), .Z(n35088) );
  NAND U35560 ( .A(n35089), .B(n35088), .Z(n35259) );
  NANDN U35561 ( .A(n35091), .B(n35090), .Z(n35095) );
  OR U35562 ( .A(n35093), .B(n35092), .Z(n35094) );
  NAND U35563 ( .A(n35095), .B(n35094), .Z(n35420) );
  NAND U35564 ( .A(n35097), .B(n35096), .Z(n35101) );
  NANDN U35565 ( .A(n35099), .B(n35098), .Z(n35100) );
  NAND U35566 ( .A(n35101), .B(n35100), .Z(n35418) );
  OR U35567 ( .A(n35107), .B(n35106), .Z(n35111) );
  NANDN U35568 ( .A(n35109), .B(n35108), .Z(n35110) );
  NAND U35569 ( .A(n35111), .B(n35110), .Z(n35401) );
  NANDN U35570 ( .A(n35117), .B(n35116), .Z(n35121) );
  NAND U35571 ( .A(n35119), .B(n35118), .Z(n35120) );
  NAND U35572 ( .A(n35121), .B(n35120), .Z(n35354) );
  XOR U35573 ( .A(a[126]), .B(n973), .Z(n35312) );
  NANDN U35574 ( .A(n35312), .B(n35313), .Z(n35124) );
  NANDN U35575 ( .A(n35122), .B(n35311), .Z(n35123) );
  NAND U35576 ( .A(n35124), .B(n35123), .Z(n35275) );
  XOR U35577 ( .A(b[57]), .B(n36100), .Z(n35296) );
  OR U35578 ( .A(n35296), .B(n965), .Z(n35127) );
  NANDN U35579 ( .A(n35125), .B(n38194), .Z(n35126) );
  NAND U35580 ( .A(n35127), .B(n35126), .Z(n35272) );
  NAND U35581 ( .A(n37469), .B(n35128), .Z(n35130) );
  XOR U35582 ( .A(n978), .B(n37336), .Z(n35316) );
  NAND U35583 ( .A(n35316), .B(n37471), .Z(n35129) );
  AND U35584 ( .A(n35130), .B(n35129), .Z(n35273) );
  XNOR U35585 ( .A(n35272), .B(n35273), .Z(n35274) );
  XNOR U35586 ( .A(n35275), .B(n35274), .Z(n35352) );
  NANDN U35587 ( .A(n35132), .B(n35131), .Z(n35136) );
  NAND U35588 ( .A(n35134), .B(n35133), .Z(n35135) );
  NAND U35589 ( .A(n35136), .B(n35135), .Z(n35353) );
  XOR U35590 ( .A(n35352), .B(n35353), .Z(n35355) );
  XOR U35591 ( .A(n35354), .B(n35355), .Z(n35399) );
  XNOR U35592 ( .A(n35400), .B(n35399), .Z(n35402) );
  XNOR U35593 ( .A(n35401), .B(n35402), .Z(n35411) );
  OR U35594 ( .A(n35138), .B(n35137), .Z(n35142) );
  NANDN U35595 ( .A(n35140), .B(n35139), .Z(n35141) );
  NAND U35596 ( .A(n35142), .B(n35141), .Z(n35412) );
  XNOR U35597 ( .A(n35411), .B(n35412), .Z(n35414) );
  XOR U35598 ( .A(n35414), .B(n35413), .Z(n35263) );
  XNOR U35599 ( .A(n35262), .B(n35263), .Z(n35265) );
  NAND U35600 ( .A(n35148), .B(n35147), .Z(n35152) );
  NANDN U35601 ( .A(n35150), .B(n35149), .Z(n35151) );
  NAND U35602 ( .A(n35152), .B(n35151), .Z(n35349) );
  XOR U35603 ( .A(b[53]), .B(n36647), .Z(n35287) );
  NANDN U35604 ( .A(n35287), .B(n37940), .Z(n35155) );
  NANDN U35605 ( .A(n35153), .B(n37941), .Z(n35154) );
  NAND U35606 ( .A(n35155), .B(n35154), .Z(n35366) );
  XOR U35607 ( .A(b[55]), .B(n36420), .Z(n35290) );
  NANDN U35608 ( .A(n35290), .B(n38075), .Z(n35158) );
  NANDN U35609 ( .A(n35156), .B(n38073), .Z(n35157) );
  NAND U35610 ( .A(n35158), .B(n35157), .Z(n35363) );
  XNOR U35611 ( .A(a[112]), .B(b[45]), .Z(n35319) );
  NANDN U35612 ( .A(n35319), .B(n37261), .Z(n35161) );
  NAND U35613 ( .A(n35159), .B(n37262), .Z(n35160) );
  AND U35614 ( .A(n35161), .B(n35160), .Z(n35364) );
  XNOR U35615 ( .A(n35363), .B(n35364), .Z(n35365) );
  XNOR U35616 ( .A(n35366), .B(n35365), .Z(n35340) );
  XOR U35617 ( .A(b[49]), .B(n37139), .Z(n35372) );
  OR U35618 ( .A(n35372), .B(n37756), .Z(n35164) );
  NANDN U35619 ( .A(n35162), .B(n37652), .Z(n35163) );
  NAND U35620 ( .A(n35164), .B(n35163), .Z(n35390) );
  NAND U35621 ( .A(n38326), .B(n35165), .Z(n35167) );
  XOR U35622 ( .A(n38400), .B(n35783), .Z(n35293) );
  NANDN U35623 ( .A(n38273), .B(n35293), .Z(n35166) );
  NAND U35624 ( .A(n35167), .B(n35166), .Z(n35387) );
  XOR U35625 ( .A(b[61]), .B(n35545), .Z(n35308) );
  OR U35626 ( .A(n35308), .B(n38371), .Z(n35170) );
  NANDN U35627 ( .A(n35168), .B(n38369), .Z(n35169) );
  AND U35628 ( .A(n35170), .B(n35169), .Z(n35388) );
  XNOR U35629 ( .A(n35387), .B(n35388), .Z(n35389) );
  XOR U35630 ( .A(n35390), .B(n35389), .Z(n35341) );
  XOR U35631 ( .A(n35340), .B(n35341), .Z(n35343) );
  NANDN U35632 ( .A(n35172), .B(n35171), .Z(n35176) );
  NAND U35633 ( .A(n35174), .B(n35173), .Z(n35175) );
  NAND U35634 ( .A(n35176), .B(n35175), .Z(n35342) );
  XNOR U35635 ( .A(n35343), .B(n35342), .Z(n35267) );
  NANDN U35636 ( .A(n35178), .B(n35177), .Z(n35182) );
  NAND U35637 ( .A(n35180), .B(n35179), .Z(n35181) );
  NAND U35638 ( .A(n35182), .B(n35181), .Z(n35328) );
  XNOR U35639 ( .A(n35328), .B(n35329), .Z(n35330) );
  NAND U35640 ( .A(n35188), .B(n35187), .Z(n35190) );
  ANDN U35641 ( .B(n35190), .A(n35189), .Z(n35360) );
  AND U35642 ( .A(a[92]), .B(b[63]), .Z(n35524) );
  XOR U35643 ( .A(b[63]), .B(n35191), .Z(n35369) );
  NANDN U35644 ( .A(n35369), .B(n38422), .Z(n35194) );
  NANDN U35645 ( .A(n35192), .B(n38423), .Z(n35193) );
  NAND U35646 ( .A(n35194), .B(n35193), .Z(n35358) );
  XNOR U35647 ( .A(n35524), .B(n35358), .Z(n35359) );
  XNOR U35648 ( .A(n35360), .B(n35359), .Z(n35331) );
  XOR U35649 ( .A(n35330), .B(n35331), .Z(n35266) );
  XNOR U35650 ( .A(n35267), .B(n35266), .Z(n35269) );
  NANDN U35651 ( .A(n35196), .B(n35195), .Z(n35200) );
  NAND U35652 ( .A(n35198), .B(n35197), .Z(n35199) );
  NAND U35653 ( .A(n35200), .B(n35199), .Z(n35337) );
  XOR U35654 ( .A(a[114]), .B(n977), .Z(n35381) );
  NANDN U35655 ( .A(n35381), .B(n37068), .Z(n35203) );
  NANDN U35656 ( .A(n35201), .B(n37069), .Z(n35202) );
  NAND U35657 ( .A(n35203), .B(n35202), .Z(n35281) );
  XOR U35658 ( .A(b[51]), .B(n36909), .Z(n35384) );
  NANDN U35659 ( .A(n35384), .B(n37803), .Z(n35206) );
  NANDN U35660 ( .A(n35204), .B(n37802), .Z(n35205) );
  NAND U35661 ( .A(n35206), .B(n35205), .Z(n35278) );
  XOR U35662 ( .A(a[124]), .B(n974), .Z(n35325) );
  NANDN U35663 ( .A(n35325), .B(n35620), .Z(n35209) );
  NANDN U35664 ( .A(n35207), .B(n35621), .Z(n35208) );
  AND U35665 ( .A(n35209), .B(n35208), .Z(n35279) );
  XNOR U35666 ( .A(n35278), .B(n35279), .Z(n35280) );
  XNOR U35667 ( .A(n35281), .B(n35280), .Z(n35396) );
  XNOR U35668 ( .A(a[122]), .B(b[35]), .Z(n35322) );
  NANDN U35669 ( .A(n35322), .B(n35985), .Z(n35212) );
  NAND U35670 ( .A(n35210), .B(n35986), .Z(n35211) );
  NAND U35671 ( .A(n35212), .B(n35211), .Z(n35305) );
  XOR U35672 ( .A(a[118]), .B(n976), .Z(n35284) );
  NANDN U35673 ( .A(n35284), .B(n36553), .Z(n35215) );
  NAND U35674 ( .A(n35213), .B(n36643), .Z(n35214) );
  NAND U35675 ( .A(n35215), .B(n35214), .Z(n35302) );
  XNOR U35676 ( .A(a[116]), .B(b[41]), .Z(n35378) );
  OR U35677 ( .A(n35378), .B(n36905), .Z(n35218) );
  NAND U35678 ( .A(n35216), .B(n36807), .Z(n35217) );
  AND U35679 ( .A(n35218), .B(n35217), .Z(n35303) );
  XNOR U35680 ( .A(n35302), .B(n35303), .Z(n35304) );
  XNOR U35681 ( .A(n35305), .B(n35304), .Z(n35393) );
  NANDN U35682 ( .A(n35219), .B(n36309), .Z(n35221) );
  XNOR U35683 ( .A(n38134), .B(b[37]), .Z(n35299) );
  NAND U35684 ( .A(n35299), .B(n36311), .Z(n35220) );
  NAND U35685 ( .A(n35221), .B(n35220), .Z(n35394) );
  XNOR U35686 ( .A(n35393), .B(n35394), .Z(n35395) );
  XOR U35687 ( .A(n35396), .B(n35395), .Z(n35335) );
  NANDN U35688 ( .A(n35223), .B(n35222), .Z(n35227) );
  NAND U35689 ( .A(n35225), .B(n35224), .Z(n35226) );
  AND U35690 ( .A(n35227), .B(n35226), .Z(n35334) );
  XOR U35691 ( .A(n35335), .B(n35334), .Z(n35336) );
  XNOR U35692 ( .A(n35337), .B(n35336), .Z(n35268) );
  XNOR U35693 ( .A(n35269), .B(n35268), .Z(n35346) );
  NANDN U35694 ( .A(n35229), .B(n35228), .Z(n35233) );
  NAND U35695 ( .A(n35231), .B(n35230), .Z(n35232) );
  AND U35696 ( .A(n35233), .B(n35232), .Z(n35407) );
  NANDN U35697 ( .A(n35235), .B(n35234), .Z(n35239) );
  NANDN U35698 ( .A(n35237), .B(n35236), .Z(n35238) );
  NAND U35699 ( .A(n35239), .B(n35238), .Z(n35406) );
  NANDN U35700 ( .A(n35241), .B(n35240), .Z(n35245) );
  OR U35701 ( .A(n35243), .B(n35242), .Z(n35244) );
  AND U35702 ( .A(n35245), .B(n35244), .Z(n35405) );
  XNOR U35703 ( .A(n35406), .B(n35405), .Z(n35408) );
  XNOR U35704 ( .A(n35407), .B(n35408), .Z(n35347) );
  XNOR U35705 ( .A(n35346), .B(n35347), .Z(n35348) );
  XOR U35706 ( .A(n35349), .B(n35348), .Z(n35264) );
  XNOR U35707 ( .A(n35265), .B(n35264), .Z(n35417) );
  XOR U35708 ( .A(n35418), .B(n35417), .Z(n35419) );
  XNOR U35709 ( .A(n35420), .B(n35419), .Z(n35256) );
  NAND U35710 ( .A(n35247), .B(n35246), .Z(n35251) );
  NAND U35711 ( .A(n35249), .B(n35248), .Z(n35250) );
  NAND U35712 ( .A(n35251), .B(n35250), .Z(n35257) );
  XNOR U35713 ( .A(n35256), .B(n35257), .Z(n35258) );
  XNOR U35714 ( .A(n35259), .B(n35258), .Z(n35255) );
  NANDN U35715 ( .A(n35253), .B(n35252), .Z(n35254) );
  XOR U35716 ( .A(n35255), .B(n35254), .Z(c[220]) );
  OR U35717 ( .A(n35255), .B(n35254), .Z(n35425) );
  NANDN U35718 ( .A(n35257), .B(n35256), .Z(n35261) );
  NAND U35719 ( .A(n35259), .B(n35258), .Z(n35260) );
  NAND U35720 ( .A(n35261), .B(n35260), .Z(n35429) );
  NAND U35721 ( .A(n35267), .B(n35266), .Z(n35271) );
  OR U35722 ( .A(n35269), .B(n35268), .Z(n35270) );
  NAND U35723 ( .A(n35271), .B(n35270), .Z(n35454) );
  NANDN U35724 ( .A(n35273), .B(n35272), .Z(n35277) );
  NAND U35725 ( .A(n35275), .B(n35274), .Z(n35276) );
  NAND U35726 ( .A(n35277), .B(n35276), .Z(n35589) );
  NANDN U35727 ( .A(n35279), .B(n35278), .Z(n35283) );
  NAND U35728 ( .A(n35281), .B(n35280), .Z(n35282) );
  NAND U35729 ( .A(n35283), .B(n35282), .Z(n35578) );
  XOR U35730 ( .A(a[119]), .B(n976), .Z(n35536) );
  NANDN U35731 ( .A(n35536), .B(n36553), .Z(n35286) );
  NANDN U35732 ( .A(n35284), .B(n36643), .Z(n35285) );
  NAND U35733 ( .A(n35286), .B(n35285), .Z(n35561) );
  XNOR U35734 ( .A(b[53]), .B(a[105]), .Z(n35473) );
  NANDN U35735 ( .A(n35473), .B(n37940), .Z(n35289) );
  NANDN U35736 ( .A(n35287), .B(n37941), .Z(n35288) );
  NAND U35737 ( .A(n35289), .B(n35288), .Z(n35558) );
  XNOR U35738 ( .A(b[55]), .B(a[103]), .Z(n35530) );
  NANDN U35739 ( .A(n35530), .B(n38075), .Z(n35292) );
  NANDN U35740 ( .A(n35290), .B(n38073), .Z(n35291) );
  AND U35741 ( .A(n35292), .B(n35291), .Z(n35559) );
  XNOR U35742 ( .A(n35558), .B(n35559), .Z(n35560) );
  XNOR U35743 ( .A(n35561), .B(n35560), .Z(n35576) );
  NAND U35744 ( .A(n38326), .B(n35293), .Z(n35295) );
  XNOR U35745 ( .A(n38400), .B(a[99]), .Z(n35533) );
  NANDN U35746 ( .A(n38273), .B(n35533), .Z(n35294) );
  NAND U35747 ( .A(n35295), .B(n35294), .Z(n35470) );
  XNOR U35748 ( .A(b[57]), .B(a[101]), .Z(n35476) );
  OR U35749 ( .A(n35476), .B(n965), .Z(n35298) );
  NANDN U35750 ( .A(n35296), .B(n38194), .Z(n35297) );
  NAND U35751 ( .A(n35298), .B(n35297), .Z(n35467) );
  XNOR U35752 ( .A(a[121]), .B(b[37]), .Z(n35500) );
  NANDN U35753 ( .A(n35500), .B(n36311), .Z(n35301) );
  NAND U35754 ( .A(n35299), .B(n36309), .Z(n35300) );
  AND U35755 ( .A(n35301), .B(n35300), .Z(n35468) );
  XNOR U35756 ( .A(n35467), .B(n35468), .Z(n35469) );
  XOR U35757 ( .A(n35470), .B(n35469), .Z(n35577) );
  XOR U35758 ( .A(n35576), .B(n35577), .Z(n35579) );
  XOR U35759 ( .A(n35578), .B(n35579), .Z(n35588) );
  XNOR U35760 ( .A(n35589), .B(n35588), .Z(n35590) );
  NANDN U35761 ( .A(n35303), .B(n35302), .Z(n35307) );
  NAND U35762 ( .A(n35305), .B(n35304), .Z(n35306) );
  NAND U35763 ( .A(n35307), .B(n35306), .Z(n35584) );
  XNOR U35764 ( .A(b[61]), .B(a[97]), .Z(n35482) );
  OR U35765 ( .A(n35482), .B(n38371), .Z(n35310) );
  NANDN U35766 ( .A(n35308), .B(n38369), .Z(n35309) );
  NAND U35767 ( .A(n35310), .B(n35309), .Z(n35567) );
  NANDN U35768 ( .A(n35312), .B(n35311), .Z(n35315) );
  XNOR U35769 ( .A(n38463), .B(b[31]), .Z(n35542) );
  NAND U35770 ( .A(n35542), .B(n35313), .Z(n35314) );
  NAND U35771 ( .A(n35315), .B(n35314), .Z(n35564) );
  NAND U35772 ( .A(n37469), .B(n35316), .Z(n35318) );
  XNOR U35773 ( .A(n978), .B(a[111]), .Z(n35552) );
  NAND U35774 ( .A(n35552), .B(n37471), .Z(n35317) );
  AND U35775 ( .A(n35318), .B(n35317), .Z(n35565) );
  XNOR U35776 ( .A(n35564), .B(n35565), .Z(n35566) );
  XNOR U35777 ( .A(n35567), .B(n35566), .Z(n35582) );
  XOR U35778 ( .A(a[113]), .B(b[45]), .Z(n35549) );
  NAND U35779 ( .A(n35549), .B(n37261), .Z(n35321) );
  NANDN U35780 ( .A(n35319), .B(n37262), .Z(n35320) );
  NAND U35781 ( .A(n35321), .B(n35320), .Z(n35494) );
  XOR U35782 ( .A(a[123]), .B(b[35]), .Z(n35503) );
  NAND U35783 ( .A(n35985), .B(n35503), .Z(n35324) );
  NANDN U35784 ( .A(n35322), .B(n35986), .Z(n35323) );
  NAND U35785 ( .A(n35324), .B(n35323), .Z(n35491) );
  XNOR U35786 ( .A(a[125]), .B(b[33]), .Z(n35485) );
  NANDN U35787 ( .A(n35485), .B(n35620), .Z(n35327) );
  NANDN U35788 ( .A(n35325), .B(n35621), .Z(n35326) );
  AND U35789 ( .A(n35327), .B(n35326), .Z(n35492) );
  XNOR U35790 ( .A(n35491), .B(n35492), .Z(n35493) );
  XOR U35791 ( .A(n35494), .B(n35493), .Z(n35583) );
  XOR U35792 ( .A(n35582), .B(n35583), .Z(n35585) );
  XOR U35793 ( .A(n35584), .B(n35585), .Z(n35591) );
  XOR U35794 ( .A(n35590), .B(n35591), .Z(n35451) );
  NANDN U35795 ( .A(n35329), .B(n35328), .Z(n35333) );
  NAND U35796 ( .A(n35331), .B(n35330), .Z(n35332) );
  NAND U35797 ( .A(n35333), .B(n35332), .Z(n35460) );
  OR U35798 ( .A(n35335), .B(n35334), .Z(n35339) );
  NAND U35799 ( .A(n35337), .B(n35336), .Z(n35338) );
  NAND U35800 ( .A(n35339), .B(n35338), .Z(n35457) );
  NANDN U35801 ( .A(n35341), .B(n35340), .Z(n35345) );
  OR U35802 ( .A(n35343), .B(n35342), .Z(n35344) );
  NAND U35803 ( .A(n35345), .B(n35344), .Z(n35458) );
  XNOR U35804 ( .A(n35457), .B(n35458), .Z(n35459) );
  XNOR U35805 ( .A(n35460), .B(n35459), .Z(n35452) );
  XOR U35806 ( .A(n35451), .B(n35452), .Z(n35453) );
  XNOR U35807 ( .A(n35454), .B(n35453), .Z(n35447) );
  NANDN U35808 ( .A(n35347), .B(n35346), .Z(n35351) );
  NAND U35809 ( .A(n35349), .B(n35348), .Z(n35350) );
  NAND U35810 ( .A(n35351), .B(n35350), .Z(n35446) );
  NANDN U35811 ( .A(n35353), .B(n35352), .Z(n35357) );
  OR U35812 ( .A(n35355), .B(n35354), .Z(n35356) );
  NAND U35813 ( .A(n35357), .B(n35356), .Z(n35515) );
  NANDN U35814 ( .A(n35524), .B(n35358), .Z(n35362) );
  NANDN U35815 ( .A(n35360), .B(n35359), .Z(n35361) );
  NAND U35816 ( .A(n35362), .B(n35361), .Z(n35573) );
  NANDN U35817 ( .A(n35364), .B(n35363), .Z(n35368) );
  NAND U35818 ( .A(n35366), .B(n35365), .Z(n35367) );
  NAND U35819 ( .A(n35368), .B(n35367), .Z(n35571) );
  XOR U35820 ( .A(b[63]), .B(n35628), .Z(n35546) );
  NANDN U35821 ( .A(n35546), .B(n38422), .Z(n35371) );
  NANDN U35822 ( .A(n35369), .B(n38423), .Z(n35370) );
  NAND U35823 ( .A(n35371), .B(n35370), .Z(n35506) );
  XNOR U35824 ( .A(b[49]), .B(a[109]), .Z(n35488) );
  OR U35825 ( .A(n35488), .B(n37756), .Z(n35374) );
  NANDN U35826 ( .A(n35372), .B(n37652), .Z(n35373) );
  AND U35827 ( .A(n35374), .B(n35373), .Z(n35507) );
  XNOR U35828 ( .A(n35506), .B(n35507), .Z(n35508) );
  NANDN U35829 ( .A(n35375), .B(b[28]), .Z(n35376) );
  NANDN U35830 ( .A(n35540), .B(n35376), .Z(n35525) );
  XNOR U35831 ( .A(n35525), .B(n35524), .Z(n35527) );
  ANDN U35832 ( .B(b[63]), .A(n35377), .Z(n35526) );
  XNOR U35833 ( .A(n35527), .B(n35526), .Z(n35509) );
  XOR U35834 ( .A(n35508), .B(n35509), .Z(n35463) );
  XOR U35835 ( .A(a[117]), .B(b[41]), .Z(n35479) );
  NANDN U35836 ( .A(n36905), .B(n35479), .Z(n35380) );
  NANDN U35837 ( .A(n35378), .B(n36807), .Z(n35379) );
  NAND U35838 ( .A(n35380), .B(n35379), .Z(n35521) );
  XNOR U35839 ( .A(a[115]), .B(b[43]), .Z(n35555) );
  NANDN U35840 ( .A(n35555), .B(n37068), .Z(n35383) );
  NANDN U35841 ( .A(n35381), .B(n37069), .Z(n35382) );
  NAND U35842 ( .A(n35383), .B(n35382), .Z(n35518) );
  XNOR U35843 ( .A(b[51]), .B(a[107]), .Z(n35497) );
  NANDN U35844 ( .A(n35497), .B(n37803), .Z(n35386) );
  NANDN U35845 ( .A(n35384), .B(n37802), .Z(n35385) );
  AND U35846 ( .A(n35386), .B(n35385), .Z(n35519) );
  XNOR U35847 ( .A(n35518), .B(n35519), .Z(n35520) );
  XNOR U35848 ( .A(n35521), .B(n35520), .Z(n35464) );
  XOR U35849 ( .A(n35463), .B(n35464), .Z(n35466) );
  NANDN U35850 ( .A(n35388), .B(n35387), .Z(n35392) );
  NAND U35851 ( .A(n35390), .B(n35389), .Z(n35391) );
  NAND U35852 ( .A(n35392), .B(n35391), .Z(n35465) );
  XNOR U35853 ( .A(n35466), .B(n35465), .Z(n35570) );
  XOR U35854 ( .A(n35571), .B(n35570), .Z(n35572) );
  XNOR U35855 ( .A(n35573), .B(n35572), .Z(n35512) );
  NANDN U35856 ( .A(n35394), .B(n35393), .Z(n35398) );
  NAND U35857 ( .A(n35396), .B(n35395), .Z(n35397) );
  AND U35858 ( .A(n35398), .B(n35397), .Z(n35513) );
  XNOR U35859 ( .A(n35512), .B(n35513), .Z(n35514) );
  XNOR U35860 ( .A(n35515), .B(n35514), .Z(n35440) );
  NAND U35861 ( .A(n35400), .B(n35399), .Z(n35404) );
  NANDN U35862 ( .A(n35402), .B(n35401), .Z(n35403) );
  AND U35863 ( .A(n35404), .B(n35403), .Z(n35439) );
  XNOR U35864 ( .A(n35440), .B(n35439), .Z(n35442) );
  OR U35865 ( .A(n35406), .B(n35405), .Z(n35410) );
  OR U35866 ( .A(n35408), .B(n35407), .Z(n35409) );
  AND U35867 ( .A(n35410), .B(n35409), .Z(n35441) );
  XNOR U35868 ( .A(n35442), .B(n35441), .Z(n35445) );
  XOR U35869 ( .A(n35446), .B(n35445), .Z(n35448) );
  XOR U35870 ( .A(n35447), .B(n35448), .Z(n35433) );
  OR U35871 ( .A(n35412), .B(n35411), .Z(n35416) );
  OR U35872 ( .A(n35414), .B(n35413), .Z(n35415) );
  NAND U35873 ( .A(n35416), .B(n35415), .Z(n35434) );
  XNOR U35874 ( .A(n35433), .B(n35434), .Z(n35436) );
  XNOR U35875 ( .A(n35435), .B(n35436), .Z(n35428) );
  IV U35876 ( .A(n35428), .Z(n35426) );
  NAND U35877 ( .A(n35418), .B(n35417), .Z(n35422) );
  NAND U35878 ( .A(n35420), .B(n35419), .Z(n35421) );
  AND U35879 ( .A(n35422), .B(n35421), .Z(n35427) );
  XNOR U35880 ( .A(n35426), .B(n35427), .Z(n35423) );
  XOR U35881 ( .A(n35429), .B(n35423), .Z(n35424) );
  XNOR U35882 ( .A(n35425), .B(n35424), .Z(c[221]) );
  NANDN U35883 ( .A(n35425), .B(n35424), .Z(n35750) );
  NANDN U35884 ( .A(n35426), .B(n35427), .Z(n35432) );
  NOR U35885 ( .A(n35428), .B(n35427), .Z(n35430) );
  NANDN U35886 ( .A(n35430), .B(n35429), .Z(n35431) );
  NAND U35887 ( .A(n35432), .B(n35431), .Z(n35601) );
  OR U35888 ( .A(n35434), .B(n35433), .Z(n35438) );
  OR U35889 ( .A(n35436), .B(n35435), .Z(n35437) );
  NAND U35890 ( .A(n35438), .B(n35437), .Z(n35599) );
  OR U35891 ( .A(n35440), .B(n35439), .Z(n35444) );
  OR U35892 ( .A(n35442), .B(n35441), .Z(n35443) );
  NAND U35893 ( .A(n35444), .B(n35443), .Z(n35593) );
  NANDN U35894 ( .A(n35446), .B(n35445), .Z(n35450) );
  OR U35895 ( .A(n35448), .B(n35447), .Z(n35449) );
  NAND U35896 ( .A(n35450), .B(n35449), .Z(n35594) );
  XOR U35897 ( .A(n35593), .B(n35594), .Z(n35595) );
  OR U35898 ( .A(n35452), .B(n35451), .Z(n35456) );
  NAND U35899 ( .A(n35454), .B(n35453), .Z(n35455) );
  NAND U35900 ( .A(n35456), .B(n35455), .Z(n35742) );
  NANDN U35901 ( .A(n35458), .B(n35457), .Z(n35462) );
  NAND U35902 ( .A(n35460), .B(n35459), .Z(n35461) );
  NAND U35903 ( .A(n35462), .B(n35461), .Z(n35739) );
  NANDN U35904 ( .A(n35468), .B(n35467), .Z(n35472) );
  NAND U35905 ( .A(n35470), .B(n35469), .Z(n35471) );
  NAND U35906 ( .A(n35472), .B(n35471), .Z(n35694) );
  XOR U35907 ( .A(b[53]), .B(n36909), .Z(n35669) );
  NANDN U35908 ( .A(n35669), .B(n37940), .Z(n35475) );
  NANDN U35909 ( .A(n35473), .B(n37941), .Z(n35474) );
  NAND U35910 ( .A(n35475), .B(n35474), .Z(n35608) );
  XOR U35911 ( .A(n983), .B(n36420), .Z(n35642) );
  NANDN U35912 ( .A(n965), .B(n35642), .Z(n35478) );
  NANDN U35913 ( .A(n35476), .B(n38194), .Z(n35477) );
  NAND U35914 ( .A(n35478), .B(n35477), .Z(n35605) );
  XNOR U35915 ( .A(a[118]), .B(b[41]), .Z(n35614) );
  OR U35916 ( .A(n35614), .B(n36905), .Z(n35481) );
  NAND U35917 ( .A(n35479), .B(n36807), .Z(n35480) );
  AND U35918 ( .A(n35481), .B(n35480), .Z(n35606) );
  XNOR U35919 ( .A(n35605), .B(n35606), .Z(n35607) );
  XNOR U35920 ( .A(n35608), .B(n35607), .Z(n35692) );
  XOR U35921 ( .A(b[61]), .B(n35783), .Z(n35663) );
  OR U35922 ( .A(n35663), .B(n38371), .Z(n35484) );
  NANDN U35923 ( .A(n35482), .B(n38369), .Z(n35483) );
  NAND U35924 ( .A(n35484), .B(n35483), .Z(n35639) );
  XOR U35925 ( .A(a[126]), .B(n974), .Z(n35622) );
  NANDN U35926 ( .A(n35622), .B(n35620), .Z(n35487) );
  NANDN U35927 ( .A(n35485), .B(n35621), .Z(n35486) );
  NAND U35928 ( .A(n35487), .B(n35486), .Z(n35636) );
  XOR U35929 ( .A(b[49]), .B(n37336), .Z(n35625) );
  OR U35930 ( .A(n35625), .B(n37756), .Z(n35490) );
  NANDN U35931 ( .A(n35488), .B(n37652), .Z(n35489) );
  AND U35932 ( .A(n35490), .B(n35489), .Z(n35637) );
  XNOR U35933 ( .A(n35636), .B(n35637), .Z(n35638) );
  XOR U35934 ( .A(n35639), .B(n35638), .Z(n35693) );
  XOR U35935 ( .A(n35692), .B(n35693), .Z(n35695) );
  XOR U35936 ( .A(n35694), .B(n35695), .Z(n35722) );
  XNOR U35937 ( .A(n35723), .B(n35722), .Z(n35724) );
  NANDN U35938 ( .A(n35492), .B(n35491), .Z(n35496) );
  NAND U35939 ( .A(n35494), .B(n35493), .Z(n35495) );
  NAND U35940 ( .A(n35496), .B(n35495), .Z(n35706) );
  XOR U35941 ( .A(b[51]), .B(n37139), .Z(n35677) );
  NANDN U35942 ( .A(n35677), .B(n37803), .Z(n35499) );
  NANDN U35943 ( .A(n35497), .B(n37802), .Z(n35498) );
  NAND U35944 ( .A(n35499), .B(n35498), .Z(n35633) );
  XOR U35945 ( .A(a[122]), .B(n975), .Z(n35666) );
  NANDN U35946 ( .A(n35666), .B(n36311), .Z(n35502) );
  NANDN U35947 ( .A(n35500), .B(n36309), .Z(n35501) );
  NAND U35948 ( .A(n35502), .B(n35501), .Z(n35630) );
  XNOR U35949 ( .A(a[124]), .B(b[35]), .Z(n35680) );
  NANDN U35950 ( .A(n35680), .B(n35985), .Z(n35505) );
  NAND U35951 ( .A(n35503), .B(n35986), .Z(n35504) );
  AND U35952 ( .A(n35505), .B(n35504), .Z(n35631) );
  XNOR U35953 ( .A(n35630), .B(n35631), .Z(n35632) );
  XNOR U35954 ( .A(n35633), .B(n35632), .Z(n35704) );
  NANDN U35955 ( .A(n35507), .B(n35506), .Z(n35511) );
  NAND U35956 ( .A(n35509), .B(n35508), .Z(n35510) );
  NAND U35957 ( .A(n35511), .B(n35510), .Z(n35705) );
  XOR U35958 ( .A(n35704), .B(n35705), .Z(n35707) );
  XOR U35959 ( .A(n35706), .B(n35707), .Z(n35725) );
  XOR U35960 ( .A(n35724), .B(n35725), .Z(n35736) );
  NANDN U35961 ( .A(n35513), .B(n35512), .Z(n35517) );
  NAND U35962 ( .A(n35515), .B(n35514), .Z(n35516) );
  NAND U35963 ( .A(n35517), .B(n35516), .Z(n35737) );
  XOR U35964 ( .A(n35736), .B(n35737), .Z(n35738) );
  XNOR U35965 ( .A(n35739), .B(n35738), .Z(n35743) );
  XNOR U35966 ( .A(n35742), .B(n35743), .Z(n35744) );
  NANDN U35967 ( .A(n35519), .B(n35518), .Z(n35523) );
  NAND U35968 ( .A(n35521), .B(n35520), .Z(n35522) );
  NAND U35969 ( .A(n35523), .B(n35522), .Z(n35710) );
  NAND U35970 ( .A(n35525), .B(n35524), .Z(n35529) );
  NANDN U35971 ( .A(n35527), .B(n35526), .Z(n35528) );
  AND U35972 ( .A(n35529), .B(n35528), .Z(n35711) );
  XNOR U35973 ( .A(n35710), .B(n35711), .Z(n35712) );
  XOR U35974 ( .A(b[55]), .B(n36647), .Z(n35645) );
  NANDN U35975 ( .A(n35645), .B(n38075), .Z(n35532) );
  NANDN U35976 ( .A(n35530), .B(n38073), .Z(n35531) );
  NAND U35977 ( .A(n35532), .B(n35531), .Z(n35660) );
  NAND U35978 ( .A(n38326), .B(n35533), .Z(n35535) );
  XOR U35979 ( .A(n38400), .B(n36100), .Z(n35611) );
  NANDN U35980 ( .A(n38273), .B(n35611), .Z(n35534) );
  NAND U35981 ( .A(n35535), .B(n35534), .Z(n35657) );
  XOR U35982 ( .A(a[120]), .B(n976), .Z(n35617) );
  NANDN U35983 ( .A(n35617), .B(n36553), .Z(n35538) );
  NANDN U35984 ( .A(n35536), .B(n36643), .Z(n35537) );
  AND U35985 ( .A(n35538), .B(n35537), .Z(n35658) );
  XNOR U35986 ( .A(n35657), .B(n35658), .Z(n35659) );
  XOR U35987 ( .A(n35660), .B(n35659), .Z(n35713) );
  XOR U35988 ( .A(n35712), .B(n35713), .Z(n35729) );
  XOR U35989 ( .A(n973), .B(n35539), .Z(n35544) );
  XOR U35990 ( .A(n35540), .B(b[30]), .Z(n35541) );
  NANDN U35991 ( .A(n35542), .B(n35541), .Z(n35543) );
  AND U35992 ( .A(n35544), .B(n35543), .Z(n35673) );
  AND U35993 ( .A(a[94]), .B(b[63]), .Z(n35819) );
  XOR U35994 ( .A(b[63]), .B(n35545), .Z(n35683) );
  NANDN U35995 ( .A(n35683), .B(n38422), .Z(n35548) );
  NANDN U35996 ( .A(n35546), .B(n38423), .Z(n35547) );
  AND U35997 ( .A(n35548), .B(n35547), .Z(n35672) );
  XOR U35998 ( .A(n35819), .B(n35672), .Z(n35674) );
  XOR U35999 ( .A(n35673), .B(n35674), .Z(n35700) );
  XNOR U36000 ( .A(n37873), .B(b[45]), .Z(n35651) );
  NAND U36001 ( .A(n35651), .B(n37261), .Z(n35551) );
  NAND U36002 ( .A(n35549), .B(n37262), .Z(n35550) );
  NAND U36003 ( .A(n35551), .B(n35550), .Z(n35689) );
  NAND U36004 ( .A(n37469), .B(n35552), .Z(n35554) );
  XOR U36005 ( .A(b[47]), .B(n37583), .Z(n35654) );
  NANDN U36006 ( .A(n35654), .B(n37471), .Z(n35553) );
  NAND U36007 ( .A(n35554), .B(n35553), .Z(n35686) );
  XOR U36008 ( .A(a[116]), .B(n977), .Z(n35648) );
  NANDN U36009 ( .A(n35648), .B(n37068), .Z(n35557) );
  NANDN U36010 ( .A(n35555), .B(n37069), .Z(n35556) );
  AND U36011 ( .A(n35557), .B(n35556), .Z(n35687) );
  XNOR U36012 ( .A(n35686), .B(n35687), .Z(n35688) );
  XNOR U36013 ( .A(n35689), .B(n35688), .Z(n35698) );
  NANDN U36014 ( .A(n35559), .B(n35558), .Z(n35563) );
  NAND U36015 ( .A(n35561), .B(n35560), .Z(n35562) );
  NAND U36016 ( .A(n35563), .B(n35562), .Z(n35699) );
  XOR U36017 ( .A(n35698), .B(n35699), .Z(n35701) );
  XOR U36018 ( .A(n35700), .B(n35701), .Z(n35726) );
  NANDN U36019 ( .A(n35565), .B(n35564), .Z(n35569) );
  NAND U36020 ( .A(n35567), .B(n35566), .Z(n35568) );
  NAND U36021 ( .A(n35569), .B(n35568), .Z(n35727) );
  XNOR U36022 ( .A(n35726), .B(n35727), .Z(n35728) );
  XNOR U36023 ( .A(n35729), .B(n35728), .Z(n35717) );
  NAND U36024 ( .A(n35571), .B(n35570), .Z(n35575) );
  NAND U36025 ( .A(n35573), .B(n35572), .Z(n35574) );
  NAND U36026 ( .A(n35575), .B(n35574), .Z(n35735) );
  NANDN U36027 ( .A(n35577), .B(n35576), .Z(n35581) );
  OR U36028 ( .A(n35579), .B(n35578), .Z(n35580) );
  NAND U36029 ( .A(n35581), .B(n35580), .Z(n35732) );
  NANDN U36030 ( .A(n35583), .B(n35582), .Z(n35587) );
  OR U36031 ( .A(n35585), .B(n35584), .Z(n35586) );
  AND U36032 ( .A(n35587), .B(n35586), .Z(n35733) );
  XNOR U36033 ( .A(n35732), .B(n35733), .Z(n35734) );
  XNOR U36034 ( .A(n35735), .B(n35734), .Z(n35716) );
  XOR U36035 ( .A(n35717), .B(n35716), .Z(n35718) );
  XOR U36036 ( .A(n35718), .B(n35719), .Z(n35745) );
  XOR U36037 ( .A(n35744), .B(n35745), .Z(n35596) );
  XNOR U36038 ( .A(n35595), .B(n35596), .Z(n35602) );
  XNOR U36039 ( .A(n35599), .B(n35602), .Z(n35592) );
  XNOR U36040 ( .A(n35601), .B(n35592), .Z(n35749) );
  XOR U36041 ( .A(n35750), .B(n35749), .Z(c[222]) );
  NANDN U36042 ( .A(n35594), .B(n35593), .Z(n35598) );
  OR U36043 ( .A(n35596), .B(n35595), .Z(n35597) );
  NAND U36044 ( .A(n35598), .B(n35597), .Z(n35752) );
  XOR U36045 ( .A(n35602), .B(n35601), .Z(n35600) );
  NAND U36046 ( .A(n35600), .B(n35599), .Z(n35604) );
  OR U36047 ( .A(n35602), .B(n35601), .Z(n35603) );
  NAND U36048 ( .A(n35604), .B(n35603), .Z(n35751) );
  NANDN U36049 ( .A(n35606), .B(n35605), .Z(n35610) );
  NAND U36050 ( .A(n35608), .B(n35607), .Z(n35609) );
  NAND U36051 ( .A(n35610), .B(n35609), .Z(n35880) );
  NAND U36052 ( .A(n38326), .B(n35611), .Z(n35613) );
  XNOR U36053 ( .A(n38400), .B(a[101]), .Z(n35844) );
  NANDN U36054 ( .A(n38273), .B(n35844), .Z(n35612) );
  NAND U36055 ( .A(n35613), .B(n35612), .Z(n35814) );
  XNOR U36056 ( .A(a[119]), .B(b[41]), .Z(n35766) );
  OR U36057 ( .A(n35766), .B(n36905), .Z(n35616) );
  NANDN U36058 ( .A(n35614), .B(n36807), .Z(n35615) );
  NAND U36059 ( .A(n35616), .B(n35615), .Z(n35811) );
  XNOR U36060 ( .A(a[121]), .B(b[39]), .Z(n35763) );
  NANDN U36061 ( .A(n35763), .B(n36553), .Z(n35619) );
  NANDN U36062 ( .A(n35617), .B(n36643), .Z(n35618) );
  AND U36063 ( .A(n35619), .B(n35618), .Z(n35812) );
  XNOR U36064 ( .A(n35811), .B(n35812), .Z(n35813) );
  XNOR U36065 ( .A(n35814), .B(n35813), .Z(n35806) );
  XOR U36066 ( .A(a[127]), .B(n974), .Z(n35779) );
  NANDN U36067 ( .A(n35779), .B(n35620), .Z(n35624) );
  NANDN U36068 ( .A(n35622), .B(n35621), .Z(n35623) );
  NAND U36069 ( .A(n35624), .B(n35623), .Z(n35787) );
  XNOR U36070 ( .A(b[49]), .B(a[111]), .Z(n35838) );
  OR U36071 ( .A(n35838), .B(n37756), .Z(n35627) );
  NANDN U36072 ( .A(n35625), .B(n37652), .Z(n35626) );
  AND U36073 ( .A(n35627), .B(n35626), .Z(n35788) );
  XNOR U36074 ( .A(n35787), .B(n35788), .Z(n35789) );
  ANDN U36075 ( .B(b[63]), .A(n35628), .Z(n35817) );
  XOR U36076 ( .A(n35629), .B(n35817), .Z(n35820) );
  XNOR U36077 ( .A(n35819), .B(n35820), .Z(n35790) );
  XOR U36078 ( .A(n35789), .B(n35790), .Z(n35805) );
  XOR U36079 ( .A(n35806), .B(n35805), .Z(n35807) );
  NANDN U36080 ( .A(n35631), .B(n35630), .Z(n35635) );
  NAND U36081 ( .A(n35633), .B(n35632), .Z(n35634) );
  AND U36082 ( .A(n35635), .B(n35634), .Z(n35808) );
  XNOR U36083 ( .A(n35807), .B(n35808), .Z(n35796) );
  NANDN U36084 ( .A(n35637), .B(n35636), .Z(n35641) );
  NAND U36085 ( .A(n35639), .B(n35638), .Z(n35640) );
  NAND U36086 ( .A(n35641), .B(n35640), .Z(n35793) );
  NAND U36087 ( .A(n38194), .B(n35642), .Z(n35644) );
  XNOR U36088 ( .A(n983), .B(a[103]), .Z(n35841) );
  NANDN U36089 ( .A(n965), .B(n35841), .Z(n35643) );
  AND U36090 ( .A(n35644), .B(n35643), .Z(n35832) );
  XNOR U36091 ( .A(b[55]), .B(a[105]), .Z(n35829) );
  NANDN U36092 ( .A(n35829), .B(n38075), .Z(n35647) );
  NANDN U36093 ( .A(n35645), .B(n38073), .Z(n35646) );
  AND U36094 ( .A(n35647), .B(n35646), .Z(n35833) );
  XOR U36095 ( .A(n35832), .B(n35833), .Z(n35834) );
  XNOR U36096 ( .A(a[117]), .B(n977), .Z(n35772) );
  NAND U36097 ( .A(n35772), .B(n37068), .Z(n35650) );
  NANDN U36098 ( .A(n35648), .B(n37069), .Z(n35649) );
  AND U36099 ( .A(n35650), .B(n35649), .Z(n35835) );
  XNOR U36100 ( .A(n35834), .B(n35835), .Z(n35865) );
  NAND U36101 ( .A(n37262), .B(n35651), .Z(n35653) );
  XNOR U36102 ( .A(a[115]), .B(b[45]), .Z(n35775) );
  NANDN U36103 ( .A(n35775), .B(n37261), .Z(n35652) );
  NAND U36104 ( .A(n35653), .B(n35652), .Z(n35863) );
  NANDN U36105 ( .A(n35654), .B(n37469), .Z(n35656) );
  XNOR U36106 ( .A(n978), .B(a[113]), .Z(n35769) );
  NAND U36107 ( .A(n35769), .B(n37471), .Z(n35655) );
  AND U36108 ( .A(n35656), .B(n35655), .Z(n35862) );
  XNOR U36109 ( .A(n35863), .B(n35862), .Z(n35864) );
  XOR U36110 ( .A(n35865), .B(n35864), .Z(n35794) );
  XOR U36111 ( .A(n35793), .B(n35794), .Z(n35795) );
  XOR U36112 ( .A(n35796), .B(n35795), .Z(n35881) );
  XOR U36113 ( .A(n35880), .B(n35881), .Z(n35882) );
  NANDN U36114 ( .A(n35658), .B(n35657), .Z(n35662) );
  NAND U36115 ( .A(n35660), .B(n35659), .Z(n35661) );
  NAND U36116 ( .A(n35662), .B(n35661), .Z(n35802) );
  XNOR U36117 ( .A(b[61]), .B(a[99]), .Z(n35850) );
  OR U36118 ( .A(n35850), .B(n38371), .Z(n35665) );
  NANDN U36119 ( .A(n35663), .B(n38369), .Z(n35664) );
  NAND U36120 ( .A(n35665), .B(n35664), .Z(n35871) );
  XNOR U36121 ( .A(a[123]), .B(b[37]), .Z(n35826) );
  NANDN U36122 ( .A(n35826), .B(n36311), .Z(n35668) );
  NANDN U36123 ( .A(n35666), .B(n36309), .Z(n35667) );
  NAND U36124 ( .A(n35668), .B(n35667), .Z(n35868) );
  XNOR U36125 ( .A(b[53]), .B(a[107]), .Z(n35823) );
  NANDN U36126 ( .A(n35823), .B(n37940), .Z(n35671) );
  NANDN U36127 ( .A(n35669), .B(n37941), .Z(n35670) );
  AND U36128 ( .A(n35671), .B(n35670), .Z(n35869) );
  XNOR U36129 ( .A(n35868), .B(n35869), .Z(n35870) );
  XOR U36130 ( .A(n35871), .B(n35870), .Z(n35874) );
  OR U36131 ( .A(n35819), .B(n35672), .Z(n35676) );
  NAND U36132 ( .A(n35674), .B(n35673), .Z(n35675) );
  NAND U36133 ( .A(n35676), .B(n35675), .Z(n35875) );
  XNOR U36134 ( .A(n35874), .B(n35875), .Z(n35877) );
  XNOR U36135 ( .A(b[51]), .B(a[109]), .Z(n35853) );
  NANDN U36136 ( .A(n35853), .B(n37803), .Z(n35679) );
  NANDN U36137 ( .A(n35677), .B(n37802), .Z(n35678) );
  NAND U36138 ( .A(n35679), .B(n35678), .Z(n35859) );
  XOR U36139 ( .A(a[125]), .B(b[35]), .Z(n35847) );
  NAND U36140 ( .A(n35985), .B(n35847), .Z(n35682) );
  NANDN U36141 ( .A(n35680), .B(n35986), .Z(n35681) );
  NAND U36142 ( .A(n35682), .B(n35681), .Z(n35856) );
  XNOR U36143 ( .A(b[63]), .B(a[97]), .Z(n35784) );
  NANDN U36144 ( .A(n35784), .B(n38422), .Z(n35685) );
  NANDN U36145 ( .A(n35683), .B(n38423), .Z(n35684) );
  AND U36146 ( .A(n35685), .B(n35684), .Z(n35857) );
  XNOR U36147 ( .A(n35856), .B(n35857), .Z(n35858) );
  XOR U36148 ( .A(n35859), .B(n35858), .Z(n35876) );
  XNOR U36149 ( .A(n35877), .B(n35876), .Z(n35800) );
  NANDN U36150 ( .A(n35687), .B(n35686), .Z(n35691) );
  NAND U36151 ( .A(n35689), .B(n35688), .Z(n35690) );
  AND U36152 ( .A(n35691), .B(n35690), .Z(n35799) );
  XNOR U36153 ( .A(n35800), .B(n35799), .Z(n35801) );
  XOR U36154 ( .A(n35802), .B(n35801), .Z(n35883) );
  XOR U36155 ( .A(n35882), .B(n35883), .Z(n35760) );
  NANDN U36156 ( .A(n35693), .B(n35692), .Z(n35697) );
  OR U36157 ( .A(n35695), .B(n35694), .Z(n35696) );
  NAND U36158 ( .A(n35697), .B(n35696), .Z(n35757) );
  NANDN U36159 ( .A(n35699), .B(n35698), .Z(n35703) );
  OR U36160 ( .A(n35701), .B(n35700), .Z(n35702) );
  NAND U36161 ( .A(n35703), .B(n35702), .Z(n35887) );
  NANDN U36162 ( .A(n35705), .B(n35704), .Z(n35709) );
  OR U36163 ( .A(n35707), .B(n35706), .Z(n35708) );
  NAND U36164 ( .A(n35709), .B(n35708), .Z(n35886) );
  XNOR U36165 ( .A(n35887), .B(n35886), .Z(n35888) );
  NANDN U36166 ( .A(n35711), .B(n35710), .Z(n35715) );
  NAND U36167 ( .A(n35713), .B(n35712), .Z(n35714) );
  AND U36168 ( .A(n35715), .B(n35714), .Z(n35889) );
  XOR U36169 ( .A(n35757), .B(n35758), .Z(n35759) );
  XNOR U36170 ( .A(n35760), .B(n35759), .Z(n35895) );
  OR U36171 ( .A(n35717), .B(n35716), .Z(n35721) );
  NAND U36172 ( .A(n35719), .B(n35718), .Z(n35720) );
  NAND U36173 ( .A(n35721), .B(n35720), .Z(n35892) );
  NANDN U36174 ( .A(n35727), .B(n35726), .Z(n35731) );
  NANDN U36175 ( .A(n35729), .B(n35728), .Z(n35730) );
  AND U36176 ( .A(n35731), .B(n35730), .Z(n35899) );
  XNOR U36177 ( .A(n35898), .B(n35899), .Z(n35901) );
  XNOR U36178 ( .A(n35901), .B(n35900), .Z(n35893) );
  XOR U36179 ( .A(n35892), .B(n35893), .Z(n35894) );
  XOR U36180 ( .A(n35895), .B(n35894), .Z(n35902) );
  OR U36181 ( .A(n35737), .B(n35736), .Z(n35741) );
  NAND U36182 ( .A(n35739), .B(n35738), .Z(n35740) );
  AND U36183 ( .A(n35741), .B(n35740), .Z(n35903) );
  XNOR U36184 ( .A(n35902), .B(n35903), .Z(n35905) );
  NANDN U36185 ( .A(n35743), .B(n35742), .Z(n35747) );
  NAND U36186 ( .A(n35745), .B(n35744), .Z(n35746) );
  NAND U36187 ( .A(n35747), .B(n35746), .Z(n35904) );
  XNOR U36188 ( .A(n35905), .B(n35904), .Z(n35753) );
  XNOR U36189 ( .A(n35751), .B(n35753), .Z(n35748) );
  XNOR U36190 ( .A(n35752), .B(n35748), .Z(n35908) );
  OR U36191 ( .A(n35750), .B(n35749), .Z(n35909) );
  XNOR U36192 ( .A(n35908), .B(n35909), .Z(c[223]) );
  OR U36193 ( .A(n35751), .B(n35752), .Z(n35756) );
  XOR U36194 ( .A(n35752), .B(n35751), .Z(n35754) );
  NAND U36195 ( .A(n35754), .B(n35753), .Z(n35755) );
  AND U36196 ( .A(n35756), .B(n35755), .Z(n35915) );
  OR U36197 ( .A(n35758), .B(n35757), .Z(n35762) );
  NAND U36198 ( .A(n35760), .B(n35759), .Z(n35761) );
  NAND U36199 ( .A(n35762), .B(n35761), .Z(n35918) );
  XOR U36200 ( .A(a[122]), .B(n976), .Z(n35965) );
  NANDN U36201 ( .A(n35965), .B(n36553), .Z(n35765) );
  NANDN U36202 ( .A(n35763), .B(n36643), .Z(n35764) );
  NAND U36203 ( .A(n35765), .B(n35764), .Z(n36029) );
  XNOR U36204 ( .A(n38134), .B(b[41]), .Z(n35974) );
  NANDN U36205 ( .A(n36905), .B(n35974), .Z(n35768) );
  NANDN U36206 ( .A(n35766), .B(n36807), .Z(n35767) );
  NAND U36207 ( .A(n35768), .B(n35767), .Z(n36026) );
  NAND U36208 ( .A(n35769), .B(n37469), .Z(n35771) );
  XOR U36209 ( .A(n37873), .B(n978), .Z(n35999) );
  NAND U36210 ( .A(n35999), .B(n37471), .Z(n35770) );
  AND U36211 ( .A(n35771), .B(n35770), .Z(n36027) );
  XNOR U36212 ( .A(n36026), .B(n36027), .Z(n36028) );
  XNOR U36213 ( .A(n36029), .B(n36028), .Z(n35941) );
  NAND U36214 ( .A(n37069), .B(n35772), .Z(n35774) );
  XNOR U36215 ( .A(n38143), .B(b[43]), .Z(n35968) );
  NAND U36216 ( .A(n35968), .B(n37068), .Z(n35773) );
  NAND U36217 ( .A(n35774), .B(n35773), .Z(n35939) );
  NANDN U36218 ( .A(n35775), .B(n37262), .Z(n35777) );
  XNOR U36219 ( .A(a[116]), .B(b[45]), .Z(n35956) );
  NANDN U36220 ( .A(n35956), .B(n37261), .Z(n35776) );
  AND U36221 ( .A(n35777), .B(n35776), .Z(n35938) );
  XNOR U36222 ( .A(n35939), .B(n35938), .Z(n35940) );
  XOR U36223 ( .A(n35941), .B(n35940), .Z(n36022) );
  XOR U36224 ( .A(n974), .B(n35778), .Z(n35782) );
  XOR U36225 ( .A(b[32]), .B(n973), .Z(n35780) );
  NAND U36226 ( .A(n35780), .B(n35779), .Z(n35781) );
  AND U36227 ( .A(n35782), .B(n35781), .Z(n35978) );
  AND U36228 ( .A(b[63]), .B(a[96]), .Z(n36132) );
  XOR U36229 ( .A(b[63]), .B(n35783), .Z(n36038) );
  NANDN U36230 ( .A(n36038), .B(n38422), .Z(n35786) );
  NANDN U36231 ( .A(n35784), .B(n38423), .Z(n35785) );
  AND U36232 ( .A(n35786), .B(n35785), .Z(n35977) );
  XNOR U36233 ( .A(n36132), .B(n35977), .Z(n35979) );
  XNOR U36234 ( .A(n35978), .B(n35979), .Z(n36020) );
  NANDN U36235 ( .A(n35788), .B(n35787), .Z(n35792) );
  NANDN U36236 ( .A(n35790), .B(n35789), .Z(n35791) );
  NAND U36237 ( .A(n35792), .B(n35791), .Z(n36021) );
  XOR U36238 ( .A(n36020), .B(n36021), .Z(n36023) );
  XNOR U36239 ( .A(n36022), .B(n36023), .Z(n35928) );
  OR U36240 ( .A(n35794), .B(n35793), .Z(n35798) );
  NANDN U36241 ( .A(n35796), .B(n35795), .Z(n35797) );
  NAND U36242 ( .A(n35798), .B(n35797), .Z(n35929) );
  XNOR U36243 ( .A(n35928), .B(n35929), .Z(n35930) );
  NANDN U36244 ( .A(n35800), .B(n35799), .Z(n35804) );
  NANDN U36245 ( .A(n35802), .B(n35801), .Z(n35803) );
  NAND U36246 ( .A(n35804), .B(n35803), .Z(n35931) );
  XOR U36247 ( .A(n35930), .B(n35931), .Z(n35927) );
  OR U36248 ( .A(n35806), .B(n35805), .Z(n35810) );
  NANDN U36249 ( .A(n35808), .B(n35807), .Z(n35809) );
  NAND U36250 ( .A(n35810), .B(n35809), .Z(n36047) );
  NANDN U36251 ( .A(n35812), .B(n35811), .Z(n35816) );
  NAND U36252 ( .A(n35814), .B(n35813), .Z(n35815) );
  NAND U36253 ( .A(n35816), .B(n35815), .Z(n35935) );
  NANDN U36254 ( .A(n35818), .B(n35817), .Z(n35822) );
  NAND U36255 ( .A(n35820), .B(n35819), .Z(n35821) );
  NAND U36256 ( .A(n35822), .B(n35821), .Z(n35932) );
  XOR U36257 ( .A(b[53]), .B(n37139), .Z(n35971) );
  NANDN U36258 ( .A(n35971), .B(n37940), .Z(n35825) );
  NANDN U36259 ( .A(n35823), .B(n37941), .Z(n35824) );
  NAND U36260 ( .A(n35825), .B(n35824), .Z(n35947) );
  XOR U36261 ( .A(a[124]), .B(n975), .Z(n35993) );
  NANDN U36262 ( .A(n35993), .B(n36311), .Z(n35828) );
  NANDN U36263 ( .A(n35826), .B(n36309), .Z(n35827) );
  NAND U36264 ( .A(n35828), .B(n35827), .Z(n35944) );
  XOR U36265 ( .A(b[55]), .B(n36909), .Z(n35959) );
  NANDN U36266 ( .A(n35959), .B(n38075), .Z(n35831) );
  NANDN U36267 ( .A(n35829), .B(n38073), .Z(n35830) );
  AND U36268 ( .A(n35831), .B(n35830), .Z(n35945) );
  XNOR U36269 ( .A(n35944), .B(n35945), .Z(n35946) );
  XNOR U36270 ( .A(n35947), .B(n35946), .Z(n35933) );
  XNOR U36271 ( .A(n35932), .B(n35933), .Z(n35934) );
  XNOR U36272 ( .A(n35935), .B(n35934), .Z(n36009) );
  OR U36273 ( .A(n35833), .B(n35832), .Z(n35837) );
  NANDN U36274 ( .A(n35835), .B(n35834), .Z(n35836) );
  NAND U36275 ( .A(n35837), .B(n35836), .Z(n36004) );
  XOR U36276 ( .A(b[49]), .B(n37583), .Z(n35990) );
  OR U36277 ( .A(n35990), .B(n37756), .Z(n35840) );
  NANDN U36278 ( .A(n35838), .B(n37652), .Z(n35839) );
  NAND U36279 ( .A(n35840), .B(n35839), .Z(n35953) );
  XOR U36280 ( .A(b[57]), .B(n36647), .Z(n35962) );
  OR U36281 ( .A(n35962), .B(n965), .Z(n35843) );
  NAND U36282 ( .A(n35841), .B(n38194), .Z(n35842) );
  NAND U36283 ( .A(n35843), .B(n35842), .Z(n35950) );
  NAND U36284 ( .A(n38326), .B(n35844), .Z(n35846) );
  XOR U36285 ( .A(n38400), .B(n36420), .Z(n35996) );
  NANDN U36286 ( .A(n38273), .B(n35996), .Z(n35845) );
  AND U36287 ( .A(n35846), .B(n35845), .Z(n35951) );
  XNOR U36288 ( .A(n35950), .B(n35951), .Z(n35952) );
  XNOR U36289 ( .A(n35953), .B(n35952), .Z(n36002) );
  XNOR U36290 ( .A(a[126]), .B(b[35]), .Z(n35987) );
  NANDN U36291 ( .A(n35987), .B(n35985), .Z(n35849) );
  NAND U36292 ( .A(n35847), .B(n35986), .Z(n35848) );
  NAND U36293 ( .A(n35849), .B(n35848), .Z(n36035) );
  XOR U36294 ( .A(b[61]), .B(n36100), .Z(n35982) );
  OR U36295 ( .A(n35982), .B(n38371), .Z(n35852) );
  NANDN U36296 ( .A(n35850), .B(n38369), .Z(n35851) );
  NAND U36297 ( .A(n35852), .B(n35851), .Z(n36032) );
  XOR U36298 ( .A(n980), .B(n37336), .Z(n36041) );
  NAND U36299 ( .A(n36041), .B(n37803), .Z(n35855) );
  NANDN U36300 ( .A(n35853), .B(n37802), .Z(n35854) );
  AND U36301 ( .A(n35855), .B(n35854), .Z(n36033) );
  XNOR U36302 ( .A(n36032), .B(n36033), .Z(n36034) );
  XOR U36303 ( .A(n36035), .B(n36034), .Z(n36003) );
  XOR U36304 ( .A(n36002), .B(n36003), .Z(n36005) );
  XOR U36305 ( .A(n36004), .B(n36005), .Z(n36008) );
  XOR U36306 ( .A(n36009), .B(n36008), .Z(n36010) );
  NANDN U36307 ( .A(n35857), .B(n35856), .Z(n35861) );
  NAND U36308 ( .A(n35859), .B(n35858), .Z(n35860) );
  NAND U36309 ( .A(n35861), .B(n35860), .Z(n36017) );
  NANDN U36310 ( .A(n35863), .B(n35862), .Z(n35867) );
  NANDN U36311 ( .A(n35865), .B(n35864), .Z(n35866) );
  NAND U36312 ( .A(n35867), .B(n35866), .Z(n36014) );
  NANDN U36313 ( .A(n35869), .B(n35868), .Z(n35873) );
  NAND U36314 ( .A(n35871), .B(n35870), .Z(n35872) );
  NAND U36315 ( .A(n35873), .B(n35872), .Z(n36015) );
  XNOR U36316 ( .A(n36014), .B(n36015), .Z(n36016) );
  XOR U36317 ( .A(n36017), .B(n36016), .Z(n36011) );
  XOR U36318 ( .A(n36010), .B(n36011), .Z(n36044) );
  OR U36319 ( .A(n35875), .B(n35874), .Z(n35879) );
  OR U36320 ( .A(n35877), .B(n35876), .Z(n35878) );
  NAND U36321 ( .A(n35879), .B(n35878), .Z(n36045) );
  XNOR U36322 ( .A(n36044), .B(n36045), .Z(n36046) );
  XNOR U36323 ( .A(n36047), .B(n36046), .Z(n35924) );
  OR U36324 ( .A(n35881), .B(n35880), .Z(n35885) );
  NANDN U36325 ( .A(n35883), .B(n35882), .Z(n35884) );
  AND U36326 ( .A(n35885), .B(n35884), .Z(n35925) );
  XNOR U36327 ( .A(n35924), .B(n35925), .Z(n35926) );
  XNOR U36328 ( .A(n35927), .B(n35926), .Z(n35919) );
  XOR U36329 ( .A(n35918), .B(n35919), .Z(n35920) );
  OR U36330 ( .A(n35887), .B(n35886), .Z(n35891) );
  OR U36331 ( .A(n35889), .B(n35888), .Z(n35890) );
  NAND U36332 ( .A(n35891), .B(n35890), .Z(n35921) );
  XOR U36333 ( .A(n35920), .B(n35921), .Z(n36053) );
  OR U36334 ( .A(n35893), .B(n35892), .Z(n35897) );
  NAND U36335 ( .A(n35895), .B(n35894), .Z(n35896) );
  NAND U36336 ( .A(n35897), .B(n35896), .Z(n36051) );
  XNOR U36337 ( .A(n36051), .B(n36050), .Z(n36052) );
  XNOR U36338 ( .A(n36053), .B(n36052), .Z(n35913) );
  NAND U36339 ( .A(n35903), .B(n35902), .Z(n35907) );
  OR U36340 ( .A(n35905), .B(n35904), .Z(n35906) );
  AND U36341 ( .A(n35907), .B(n35906), .Z(n35912) );
  XNOR U36342 ( .A(n35913), .B(n35912), .Z(n35914) );
  XNOR U36343 ( .A(n35915), .B(n35914), .Z(n35910) );
  NANDN U36344 ( .A(n35909), .B(n35908), .Z(n35911) );
  XNOR U36345 ( .A(n35910), .B(n35911), .Z(c[224]) );
  NANDN U36346 ( .A(n35911), .B(n35910), .Z(n36203) );
  NANDN U36347 ( .A(n35913), .B(n35912), .Z(n35917) );
  NANDN U36348 ( .A(n35915), .B(n35914), .Z(n35916) );
  AND U36349 ( .A(n35917), .B(n35916), .Z(n36059) );
  OR U36350 ( .A(n35919), .B(n35918), .Z(n35923) );
  NANDN U36351 ( .A(n35921), .B(n35920), .Z(n35922) );
  NAND U36352 ( .A(n35923), .B(n35922), .Z(n36199) );
  NANDN U36353 ( .A(n35933), .B(n35932), .Z(n35937) );
  NAND U36354 ( .A(n35935), .B(n35934), .Z(n35936) );
  NAND U36355 ( .A(n35937), .B(n35936), .Z(n36193) );
  NANDN U36356 ( .A(n35939), .B(n35938), .Z(n35943) );
  NAND U36357 ( .A(n35941), .B(n35940), .Z(n35942) );
  NAND U36358 ( .A(n35943), .B(n35942), .Z(n36148) );
  NANDN U36359 ( .A(n35945), .B(n35944), .Z(n35949) );
  NAND U36360 ( .A(n35947), .B(n35946), .Z(n35948) );
  NAND U36361 ( .A(n35949), .B(n35948), .Z(n36146) );
  NANDN U36362 ( .A(n35951), .B(n35950), .Z(n35955) );
  NAND U36363 ( .A(n35953), .B(n35952), .Z(n35954) );
  AND U36364 ( .A(n35955), .B(n35954), .Z(n36145) );
  XNOR U36365 ( .A(n36146), .B(n36145), .Z(n36147) );
  XNOR U36366 ( .A(n36148), .B(n36147), .Z(n36079) );
  XOR U36367 ( .A(a[117]), .B(b[45]), .Z(n36172) );
  NAND U36368 ( .A(n36172), .B(n37261), .Z(n35958) );
  NANDN U36369 ( .A(n35956), .B(n37262), .Z(n35957) );
  NAND U36370 ( .A(n35958), .B(n35957), .Z(n36127) );
  XNOR U36371 ( .A(b[55]), .B(a[107]), .Z(n36136) );
  NANDN U36372 ( .A(n36136), .B(n38075), .Z(n35961) );
  NANDN U36373 ( .A(n35959), .B(n38073), .Z(n35960) );
  NAND U36374 ( .A(n35961), .B(n35960), .Z(n36124) );
  XNOR U36375 ( .A(b[57]), .B(a[105]), .Z(n36181) );
  OR U36376 ( .A(n36181), .B(n965), .Z(n35964) );
  NANDN U36377 ( .A(n35962), .B(n38194), .Z(n35963) );
  AND U36378 ( .A(n35964), .B(n35963), .Z(n36125) );
  XNOR U36379 ( .A(n36124), .B(n36125), .Z(n36126) );
  XNOR U36380 ( .A(n36127), .B(n36126), .Z(n36085) );
  XNOR U36381 ( .A(a[123]), .B(b[39]), .Z(n36112) );
  NANDN U36382 ( .A(n36112), .B(n36553), .Z(n35967) );
  NANDN U36383 ( .A(n35965), .B(n36643), .Z(n35966) );
  NAND U36384 ( .A(n35967), .B(n35966), .Z(n36097) );
  XOR U36385 ( .A(a[119]), .B(n977), .Z(n36187) );
  NANDN U36386 ( .A(n36187), .B(n37068), .Z(n35970) );
  NAND U36387 ( .A(n35968), .B(n37069), .Z(n35969) );
  NAND U36388 ( .A(n35970), .B(n35969), .Z(n36094) );
  XNOR U36389 ( .A(b[53]), .B(a[109]), .Z(n36178) );
  NANDN U36390 ( .A(n36178), .B(n37940), .Z(n35973) );
  NANDN U36391 ( .A(n35971), .B(n37941), .Z(n35972) );
  AND U36392 ( .A(n35973), .B(n35972), .Z(n36095) );
  XNOR U36393 ( .A(n36094), .B(n36095), .Z(n36096) );
  XNOR U36394 ( .A(n36097), .B(n36096), .Z(n36082) );
  NAND U36395 ( .A(n36807), .B(n35974), .Z(n35976) );
  XOR U36396 ( .A(a[121]), .B(b[41]), .Z(n36169) );
  NANDN U36397 ( .A(n36905), .B(n36169), .Z(n35975) );
  NAND U36398 ( .A(n35976), .B(n35975), .Z(n36083) );
  XNOR U36399 ( .A(n36082), .B(n36083), .Z(n36084) );
  XOR U36400 ( .A(n36085), .B(n36084), .Z(n36077) );
  OR U36401 ( .A(n35977), .B(n36132), .Z(n35981) );
  NANDN U36402 ( .A(n35979), .B(n35978), .Z(n35980) );
  NAND U36403 ( .A(n35981), .B(n35980), .Z(n36091) );
  NANDN U36404 ( .A(n35982), .B(n38369), .Z(n35984) );
  XNOR U36405 ( .A(n984), .B(a[101]), .Z(n36142) );
  NANDN U36406 ( .A(n38371), .B(n36142), .Z(n35983) );
  AND U36407 ( .A(n35984), .B(n35983), .Z(n36118) );
  XNOR U36408 ( .A(a[127]), .B(b[35]), .Z(n36105) );
  NANDN U36409 ( .A(n36105), .B(n35985), .Z(n35989) );
  NANDN U36410 ( .A(n35987), .B(n35986), .Z(n35988) );
  AND U36411 ( .A(n35989), .B(n35988), .Z(n36119) );
  XOR U36412 ( .A(n36118), .B(n36119), .Z(n36120) );
  XNOR U36413 ( .A(b[49]), .B(a[113]), .Z(n36175) );
  OR U36414 ( .A(n36175), .B(n37756), .Z(n35992) );
  NANDN U36415 ( .A(n35990), .B(n37652), .Z(n35991) );
  AND U36416 ( .A(n35992), .B(n35991), .Z(n36121) );
  XNOR U36417 ( .A(n36120), .B(n36121), .Z(n36089) );
  XNOR U36418 ( .A(a[125]), .B(b[37]), .Z(n36115) );
  NANDN U36419 ( .A(n36115), .B(n36311), .Z(n35995) );
  NANDN U36420 ( .A(n35993), .B(n36309), .Z(n35994) );
  NAND U36421 ( .A(n35995), .B(n35994), .Z(n36166) );
  NAND U36422 ( .A(n38326), .B(n35996), .Z(n35998) );
  XNOR U36423 ( .A(n38400), .B(a[103]), .Z(n36139) );
  NANDN U36424 ( .A(n38273), .B(n36139), .Z(n35997) );
  NAND U36425 ( .A(n35998), .B(n35997), .Z(n36163) );
  NAND U36426 ( .A(n37469), .B(n35999), .Z(n36001) );
  XNOR U36427 ( .A(a[115]), .B(n978), .Z(n36184) );
  NAND U36428 ( .A(n36184), .B(n37471), .Z(n36000) );
  AND U36429 ( .A(n36001), .B(n36000), .Z(n36164) );
  XNOR U36430 ( .A(n36163), .B(n36164), .Z(n36165) );
  XOR U36431 ( .A(n36166), .B(n36165), .Z(n36088) );
  XOR U36432 ( .A(n36089), .B(n36088), .Z(n36090) );
  XNOR U36433 ( .A(n36091), .B(n36090), .Z(n36076) );
  XOR U36434 ( .A(n36077), .B(n36076), .Z(n36078) );
  XOR U36435 ( .A(n36079), .B(n36078), .Z(n36190) );
  NANDN U36436 ( .A(n36003), .B(n36002), .Z(n36007) );
  OR U36437 ( .A(n36005), .B(n36004), .Z(n36006) );
  AND U36438 ( .A(n36007), .B(n36006), .Z(n36191) );
  XOR U36439 ( .A(n36190), .B(n36191), .Z(n36192) );
  XNOR U36440 ( .A(n36193), .B(n36192), .Z(n36066) );
  NAND U36441 ( .A(n36009), .B(n36008), .Z(n36013) );
  NANDN U36442 ( .A(n36011), .B(n36010), .Z(n36012) );
  AND U36443 ( .A(n36013), .B(n36012), .Z(n36067) );
  XNOR U36444 ( .A(n36066), .B(n36067), .Z(n36068) );
  NANDN U36445 ( .A(n36015), .B(n36014), .Z(n36019) );
  NANDN U36446 ( .A(n36017), .B(n36016), .Z(n36018) );
  NAND U36447 ( .A(n36019), .B(n36018), .Z(n36072) );
  OR U36448 ( .A(n36021), .B(n36020), .Z(n36025) );
  NAND U36449 ( .A(n36023), .B(n36022), .Z(n36024) );
  NAND U36450 ( .A(n36025), .B(n36024), .Z(n36071) );
  NANDN U36451 ( .A(n36027), .B(n36026), .Z(n36031) );
  NAND U36452 ( .A(n36029), .B(n36028), .Z(n36030) );
  NAND U36453 ( .A(n36031), .B(n36030), .Z(n36153) );
  NANDN U36454 ( .A(n36033), .B(n36032), .Z(n36037) );
  NAND U36455 ( .A(n36035), .B(n36034), .Z(n36036) );
  NAND U36456 ( .A(n36037), .B(n36036), .Z(n36152) );
  NANDN U36457 ( .A(n985), .B(a[97]), .Z(n36131) );
  XNOR U36458 ( .A(n36130), .B(n36131), .Z(n36133) );
  XNOR U36459 ( .A(n36132), .B(n36133), .Z(n36158) );
  XNOR U36460 ( .A(n985), .B(a[99]), .Z(n36101) );
  NAND U36461 ( .A(n36101), .B(n38422), .Z(n36040) );
  NANDN U36462 ( .A(n36038), .B(n38423), .Z(n36039) );
  NAND U36463 ( .A(n36040), .B(n36039), .Z(n36157) );
  XOR U36464 ( .A(n36158), .B(n36157), .Z(n36159) );
  NAND U36465 ( .A(n37802), .B(n36041), .Z(n36043) );
  XNOR U36466 ( .A(b[51]), .B(a[111]), .Z(n36109) );
  NANDN U36467 ( .A(n36109), .B(n37803), .Z(n36042) );
  AND U36468 ( .A(n36043), .B(n36042), .Z(n36160) );
  XOR U36469 ( .A(n36159), .B(n36160), .Z(n36151) );
  XOR U36470 ( .A(n36152), .B(n36151), .Z(n36154) );
  XOR U36471 ( .A(n36153), .B(n36154), .Z(n36070) );
  XNOR U36472 ( .A(n36071), .B(n36070), .Z(n36073) );
  XNOR U36473 ( .A(n36072), .B(n36073), .Z(n36069) );
  XOR U36474 ( .A(n36068), .B(n36069), .Z(n36060) );
  XNOR U36475 ( .A(n36061), .B(n36060), .Z(n36062) );
  NANDN U36476 ( .A(n36045), .B(n36044), .Z(n36049) );
  NAND U36477 ( .A(n36047), .B(n36046), .Z(n36048) );
  AND U36478 ( .A(n36049), .B(n36048), .Z(n36063) );
  XNOR U36479 ( .A(n36062), .B(n36063), .Z(n36197) );
  XNOR U36480 ( .A(n36196), .B(n36197), .Z(n36198) );
  XNOR U36481 ( .A(n36199), .B(n36198), .Z(n36057) );
  NANDN U36482 ( .A(n36051), .B(n36050), .Z(n36055) );
  NAND U36483 ( .A(n36053), .B(n36052), .Z(n36054) );
  AND U36484 ( .A(n36055), .B(n36054), .Z(n36058) );
  XOR U36485 ( .A(n36057), .B(n36058), .Z(n36056) );
  XNOR U36486 ( .A(n36059), .B(n36056), .Z(n36202) );
  XOR U36487 ( .A(n36203), .B(n36202), .Z(c[225]) );
  NANDN U36488 ( .A(n36061), .B(n36060), .Z(n36065) );
  NAND U36489 ( .A(n36063), .B(n36062), .Z(n36064) );
  NAND U36490 ( .A(n36065), .B(n36064), .Z(n36338) );
  NAND U36491 ( .A(n36071), .B(n36070), .Z(n36075) );
  NANDN U36492 ( .A(n36073), .B(n36072), .Z(n36074) );
  NAND U36493 ( .A(n36075), .B(n36074), .Z(n36213) );
  OR U36494 ( .A(n36077), .B(n36076), .Z(n36081) );
  NAND U36495 ( .A(n36079), .B(n36078), .Z(n36080) );
  NAND U36496 ( .A(n36081), .B(n36080), .Z(n36219) );
  NANDN U36497 ( .A(n36083), .B(n36082), .Z(n36087) );
  NAND U36498 ( .A(n36085), .B(n36084), .Z(n36086) );
  NAND U36499 ( .A(n36087), .B(n36086), .Z(n36332) );
  OR U36500 ( .A(n36089), .B(n36088), .Z(n36093) );
  NANDN U36501 ( .A(n36091), .B(n36090), .Z(n36092) );
  NAND U36502 ( .A(n36093), .B(n36092), .Z(n36329) );
  NANDN U36503 ( .A(n36095), .B(n36094), .Z(n36099) );
  NAND U36504 ( .A(n36097), .B(n36096), .Z(n36098) );
  NAND U36505 ( .A(n36099), .B(n36098), .Z(n36326) );
  XOR U36506 ( .A(b[63]), .B(n36100), .Z(n36250) );
  NANDN U36507 ( .A(n36250), .B(n38422), .Z(n36103) );
  NAND U36508 ( .A(n36101), .B(n38423), .Z(n36102) );
  NAND U36509 ( .A(n36103), .B(n36102), .Z(n36254) );
  XNOR U36510 ( .A(b[35]), .B(n36104), .Z(n36108) );
  XOR U36511 ( .A(b[34]), .B(n974), .Z(n36106) );
  NAND U36512 ( .A(n36106), .B(n36105), .Z(n36107) );
  AND U36513 ( .A(n36108), .B(n36107), .Z(n36253) );
  AND U36514 ( .A(b[63]), .B(a[98]), .Z(n36384) );
  XOR U36515 ( .A(n36253), .B(n36384), .Z(n36255) );
  XNOR U36516 ( .A(n36254), .B(n36255), .Z(n36324) );
  XOR U36517 ( .A(n980), .B(n37583), .Z(n36314) );
  NAND U36518 ( .A(n36314), .B(n37803), .Z(n36111) );
  NANDN U36519 ( .A(n36109), .B(n37802), .Z(n36110) );
  NAND U36520 ( .A(n36111), .B(n36110), .Z(n36297) );
  XOR U36521 ( .A(a[124]), .B(n976), .Z(n36279) );
  NANDN U36522 ( .A(n36279), .B(n36553), .Z(n36114) );
  NANDN U36523 ( .A(n36112), .B(n36643), .Z(n36113) );
  NAND U36524 ( .A(n36114), .B(n36113), .Z(n36294) );
  XOR U36525 ( .A(a[126]), .B(n975), .Z(n36310) );
  NANDN U36526 ( .A(n36310), .B(n36311), .Z(n36117) );
  NANDN U36527 ( .A(n36115), .B(n36309), .Z(n36116) );
  AND U36528 ( .A(n36117), .B(n36116), .Z(n36295) );
  XNOR U36529 ( .A(n36294), .B(n36295), .Z(n36296) );
  XOR U36530 ( .A(n36297), .B(n36296), .Z(n36323) );
  XOR U36531 ( .A(n36324), .B(n36323), .Z(n36325) );
  XNOR U36532 ( .A(n36326), .B(n36325), .Z(n36222) );
  OR U36533 ( .A(n36119), .B(n36118), .Z(n36123) );
  NANDN U36534 ( .A(n36121), .B(n36120), .Z(n36122) );
  AND U36535 ( .A(n36123), .B(n36122), .Z(n36223) );
  XNOR U36536 ( .A(n36222), .B(n36223), .Z(n36225) );
  NANDN U36537 ( .A(n36125), .B(n36124), .Z(n36129) );
  NAND U36538 ( .A(n36127), .B(n36126), .Z(n36128) );
  NAND U36539 ( .A(n36129), .B(n36128), .Z(n36317) );
  OR U36540 ( .A(n36131), .B(n36130), .Z(n36135) );
  NANDN U36541 ( .A(n36133), .B(n36132), .Z(n36134) );
  AND U36542 ( .A(n36135), .B(n36134), .Z(n36318) );
  XNOR U36543 ( .A(n36317), .B(n36318), .Z(n36319) );
  XOR U36544 ( .A(b[55]), .B(n37139), .Z(n36303) );
  NANDN U36545 ( .A(n36303), .B(n38075), .Z(n36138) );
  NANDN U36546 ( .A(n36136), .B(n38073), .Z(n36137) );
  NAND U36547 ( .A(n36138), .B(n36137), .Z(n36273) );
  NAND U36548 ( .A(n38326), .B(n36139), .Z(n36141) );
  XOR U36549 ( .A(n38400), .B(n36647), .Z(n36306) );
  NANDN U36550 ( .A(n38273), .B(n36306), .Z(n36140) );
  NAND U36551 ( .A(n36141), .B(n36140), .Z(n36270) );
  XOR U36552 ( .A(b[61]), .B(n36420), .Z(n36247) );
  OR U36553 ( .A(n36247), .B(n38371), .Z(n36144) );
  NAND U36554 ( .A(n36142), .B(n38369), .Z(n36143) );
  AND U36555 ( .A(n36144), .B(n36143), .Z(n36271) );
  XNOR U36556 ( .A(n36270), .B(n36271), .Z(n36272) );
  XOR U36557 ( .A(n36273), .B(n36272), .Z(n36320) );
  XOR U36558 ( .A(n36319), .B(n36320), .Z(n36224) );
  XNOR U36559 ( .A(n36225), .B(n36224), .Z(n36330) );
  XNOR U36560 ( .A(n36329), .B(n36330), .Z(n36331) );
  XOR U36561 ( .A(n36332), .B(n36331), .Z(n36218) );
  XNOR U36562 ( .A(n36219), .B(n36218), .Z(n36220) );
  NANDN U36563 ( .A(n36146), .B(n36145), .Z(n36150) );
  NAND U36564 ( .A(n36148), .B(n36147), .Z(n36149) );
  NAND U36565 ( .A(n36150), .B(n36149), .Z(n36231) );
  NANDN U36566 ( .A(n36152), .B(n36151), .Z(n36156) );
  OR U36567 ( .A(n36154), .B(n36153), .Z(n36155) );
  NAND U36568 ( .A(n36156), .B(n36155), .Z(n36228) );
  OR U36569 ( .A(n36158), .B(n36157), .Z(n36162) );
  NAND U36570 ( .A(n36160), .B(n36159), .Z(n36161) );
  NAND U36571 ( .A(n36162), .B(n36161), .Z(n36237) );
  NANDN U36572 ( .A(n36164), .B(n36163), .Z(n36168) );
  NAND U36573 ( .A(n36166), .B(n36165), .Z(n36167) );
  NAND U36574 ( .A(n36168), .B(n36167), .Z(n36235) );
  XNOR U36575 ( .A(a[122]), .B(b[41]), .Z(n36276) );
  OR U36576 ( .A(n36276), .B(n36905), .Z(n36171) );
  NAND U36577 ( .A(n36169), .B(n36807), .Z(n36170) );
  NAND U36578 ( .A(n36171), .B(n36170), .Z(n36261) );
  XNOR U36579 ( .A(a[118]), .B(b[45]), .Z(n36288) );
  NANDN U36580 ( .A(n36288), .B(n37261), .Z(n36174) );
  NAND U36581 ( .A(n36172), .B(n37262), .Z(n36173) );
  NAND U36582 ( .A(n36174), .B(n36173), .Z(n36258) );
  XOR U36583 ( .A(a[114]), .B(n979), .Z(n36300) );
  OR U36584 ( .A(n36300), .B(n37756), .Z(n36177) );
  NANDN U36585 ( .A(n36175), .B(n37652), .Z(n36176) );
  AND U36586 ( .A(n36177), .B(n36176), .Z(n36259) );
  XNOR U36587 ( .A(n36258), .B(n36259), .Z(n36260) );
  XNOR U36588 ( .A(n36261), .B(n36260), .Z(n36243) );
  XOR U36589 ( .A(b[53]), .B(n37336), .Z(n36282) );
  NANDN U36590 ( .A(n36282), .B(n37940), .Z(n36180) );
  NANDN U36591 ( .A(n36178), .B(n37941), .Z(n36179) );
  NAND U36592 ( .A(n36180), .B(n36179), .Z(n36267) );
  XOR U36593 ( .A(b[57]), .B(n36909), .Z(n36285) );
  OR U36594 ( .A(n36285), .B(n965), .Z(n36183) );
  NANDN U36595 ( .A(n36181), .B(n38194), .Z(n36182) );
  NAND U36596 ( .A(n36183), .B(n36182), .Z(n36264) );
  NAND U36597 ( .A(n37469), .B(n36184), .Z(n36186) );
  XOR U36598 ( .A(n38046), .B(n978), .Z(n36244) );
  NAND U36599 ( .A(n36244), .B(n37471), .Z(n36185) );
  AND U36600 ( .A(n36186), .B(n36185), .Z(n36265) );
  XNOR U36601 ( .A(n36264), .B(n36265), .Z(n36266) );
  XNOR U36602 ( .A(n36267), .B(n36266), .Z(n36240) );
  NANDN U36603 ( .A(n36187), .B(n37069), .Z(n36189) );
  XNOR U36604 ( .A(n38134), .B(b[43]), .Z(n36291) );
  NAND U36605 ( .A(n36291), .B(n37068), .Z(n36188) );
  NAND U36606 ( .A(n36189), .B(n36188), .Z(n36241) );
  XNOR U36607 ( .A(n36240), .B(n36241), .Z(n36242) );
  XOR U36608 ( .A(n36243), .B(n36242), .Z(n36234) );
  XNOR U36609 ( .A(n36235), .B(n36234), .Z(n36236) );
  XNOR U36610 ( .A(n36237), .B(n36236), .Z(n36229) );
  XNOR U36611 ( .A(n36228), .B(n36229), .Z(n36230) );
  XOR U36612 ( .A(n36231), .B(n36230), .Z(n36221) );
  XOR U36613 ( .A(n36220), .B(n36221), .Z(n36212) );
  XNOR U36614 ( .A(n36213), .B(n36212), .Z(n36215) );
  NAND U36615 ( .A(n36191), .B(n36190), .Z(n36195) );
  NAND U36616 ( .A(n36193), .B(n36192), .Z(n36194) );
  AND U36617 ( .A(n36195), .B(n36194), .Z(n36214) );
  XNOR U36618 ( .A(n36215), .B(n36214), .Z(n36335) );
  XOR U36619 ( .A(n36336), .B(n36335), .Z(n36337) );
  XNOR U36620 ( .A(n36338), .B(n36337), .Z(n36206) );
  NANDN U36621 ( .A(n36197), .B(n36196), .Z(n36201) );
  NAND U36622 ( .A(n36199), .B(n36198), .Z(n36200) );
  NAND U36623 ( .A(n36201), .B(n36200), .Z(n36207) );
  XOR U36624 ( .A(n36206), .B(n36207), .Z(n36209) );
  XNOR U36625 ( .A(n36208), .B(n36209), .Z(n36204) );
  OR U36626 ( .A(n36203), .B(n36202), .Z(n36205) );
  XNOR U36627 ( .A(n36204), .B(n36205), .Z(c[226]) );
  NANDN U36628 ( .A(n36205), .B(n36204), .Z(n36343) );
  NANDN U36629 ( .A(n36207), .B(n36206), .Z(n36211) );
  NANDN U36630 ( .A(n36209), .B(n36208), .Z(n36210) );
  NAND U36631 ( .A(n36211), .B(n36210), .Z(n36346) );
  NAND U36632 ( .A(n36213), .B(n36212), .Z(n36217) );
  NANDN U36633 ( .A(n36215), .B(n36214), .Z(n36216) );
  NAND U36634 ( .A(n36217), .B(n36216), .Z(n36477) );
  OR U36635 ( .A(n36223), .B(n36222), .Z(n36227) );
  NANDN U36636 ( .A(n36225), .B(n36224), .Z(n36226) );
  NAND U36637 ( .A(n36227), .B(n36226), .Z(n36350) );
  NANDN U36638 ( .A(n36229), .B(n36228), .Z(n36233) );
  NAND U36639 ( .A(n36231), .B(n36230), .Z(n36232) );
  NAND U36640 ( .A(n36233), .B(n36232), .Z(n36347) );
  NANDN U36641 ( .A(n36235), .B(n36234), .Z(n36239) );
  NAND U36642 ( .A(n36237), .B(n36236), .Z(n36238) );
  NAND U36643 ( .A(n36239), .B(n36238), .Z(n36362) );
  NAND U36644 ( .A(n37469), .B(n36244), .Z(n36246) );
  XNOR U36645 ( .A(a[117]), .B(n978), .Z(n36395) );
  NAND U36646 ( .A(n36395), .B(n37471), .Z(n36245) );
  NAND U36647 ( .A(n36246), .B(n36245), .Z(n36442) );
  XNOR U36648 ( .A(b[61]), .B(a[103]), .Z(n36457) );
  OR U36649 ( .A(n36457), .B(n38371), .Z(n36249) );
  NANDN U36650 ( .A(n36247), .B(n38369), .Z(n36248) );
  NAND U36651 ( .A(n36249), .B(n36248), .Z(n36439) );
  XNOR U36652 ( .A(b[63]), .B(a[101]), .Z(n36421) );
  NANDN U36653 ( .A(n36421), .B(n38422), .Z(n36252) );
  NANDN U36654 ( .A(n36250), .B(n38423), .Z(n36251) );
  AND U36655 ( .A(n36252), .B(n36251), .Z(n36440) );
  XNOR U36656 ( .A(n36439), .B(n36440), .Z(n36441) );
  XNOR U36657 ( .A(n36442), .B(n36441), .Z(n36368) );
  NANDN U36658 ( .A(n36384), .B(n36253), .Z(n36257) );
  NANDN U36659 ( .A(n36255), .B(n36254), .Z(n36256) );
  NAND U36660 ( .A(n36257), .B(n36256), .Z(n36366) );
  NANDN U36661 ( .A(n36259), .B(n36258), .Z(n36263) );
  NAND U36662 ( .A(n36261), .B(n36260), .Z(n36262) );
  AND U36663 ( .A(n36263), .B(n36262), .Z(n36365) );
  XNOR U36664 ( .A(n36366), .B(n36365), .Z(n36367) );
  XOR U36665 ( .A(n36368), .B(n36367), .Z(n36359) );
  XOR U36666 ( .A(n36360), .B(n36359), .Z(n36361) );
  XNOR U36667 ( .A(n36362), .B(n36361), .Z(n36353) );
  NANDN U36668 ( .A(n36265), .B(n36264), .Z(n36269) );
  NAND U36669 ( .A(n36267), .B(n36266), .Z(n36268) );
  NAND U36670 ( .A(n36269), .B(n36268), .Z(n36464) );
  NANDN U36671 ( .A(n36271), .B(n36270), .Z(n36275) );
  NAND U36672 ( .A(n36273), .B(n36272), .Z(n36274) );
  NAND U36673 ( .A(n36275), .B(n36274), .Z(n36373) );
  XOR U36674 ( .A(a[123]), .B(b[41]), .Z(n36424) );
  NANDN U36675 ( .A(n36905), .B(n36424), .Z(n36278) );
  NANDN U36676 ( .A(n36276), .B(n36807), .Z(n36277) );
  NAND U36677 ( .A(n36278), .B(n36277), .Z(n36407) );
  XNOR U36678 ( .A(a[125]), .B(b[39]), .Z(n36454) );
  NANDN U36679 ( .A(n36454), .B(n36553), .Z(n36281) );
  NANDN U36680 ( .A(n36279), .B(n36643), .Z(n36280) );
  NAND U36681 ( .A(n36281), .B(n36280), .Z(n36404) );
  XNOR U36682 ( .A(b[53]), .B(a[111]), .Z(n36430) );
  NANDN U36683 ( .A(n36430), .B(n37940), .Z(n36284) );
  NANDN U36684 ( .A(n36282), .B(n37941), .Z(n36283) );
  AND U36685 ( .A(n36284), .B(n36283), .Z(n36405) );
  XNOR U36686 ( .A(n36404), .B(n36405), .Z(n36406) );
  XNOR U36687 ( .A(n36407), .B(n36406), .Z(n36371) );
  XNOR U36688 ( .A(n983), .B(a[107]), .Z(n36445) );
  NANDN U36689 ( .A(n965), .B(n36445), .Z(n36287) );
  NANDN U36690 ( .A(n36285), .B(n38194), .Z(n36286) );
  NAND U36691 ( .A(n36287), .B(n36286), .Z(n36436) );
  XNOR U36692 ( .A(a[119]), .B(b[45]), .Z(n36392) );
  NANDN U36693 ( .A(n36392), .B(n37261), .Z(n36290) );
  NANDN U36694 ( .A(n36288), .B(n37262), .Z(n36289) );
  NAND U36695 ( .A(n36290), .B(n36289), .Z(n36433) );
  XNOR U36696 ( .A(a[121]), .B(b[43]), .Z(n36448) );
  NANDN U36697 ( .A(n36448), .B(n37068), .Z(n36293) );
  NAND U36698 ( .A(n36291), .B(n37069), .Z(n36292) );
  AND U36699 ( .A(n36293), .B(n36292), .Z(n36434) );
  XNOR U36700 ( .A(n36433), .B(n36434), .Z(n36435) );
  XOR U36701 ( .A(n36436), .B(n36435), .Z(n36372) );
  XOR U36702 ( .A(n36371), .B(n36372), .Z(n36374) );
  XOR U36703 ( .A(n36373), .B(n36374), .Z(n36463) );
  XOR U36704 ( .A(n36464), .B(n36463), .Z(n36466) );
  NANDN U36705 ( .A(n36295), .B(n36294), .Z(n36299) );
  NAND U36706 ( .A(n36297), .B(n36296), .Z(n36298) );
  NAND U36707 ( .A(n36299), .B(n36298), .Z(n36412) );
  XNOR U36708 ( .A(a[115]), .B(n979), .Z(n36389) );
  NANDN U36709 ( .A(n37756), .B(n36389), .Z(n36302) );
  NANDN U36710 ( .A(n36300), .B(n37652), .Z(n36301) );
  NAND U36711 ( .A(n36302), .B(n36301), .Z(n36401) );
  XNOR U36712 ( .A(b[55]), .B(a[109]), .Z(n36451) );
  NANDN U36713 ( .A(n36451), .B(n38075), .Z(n36305) );
  NANDN U36714 ( .A(n36303), .B(n38073), .Z(n36304) );
  NAND U36715 ( .A(n36305), .B(n36304), .Z(n36398) );
  NAND U36716 ( .A(n38326), .B(n36306), .Z(n36308) );
  XNOR U36717 ( .A(n38400), .B(a[105]), .Z(n36427) );
  NANDN U36718 ( .A(n38273), .B(n36427), .Z(n36307) );
  AND U36719 ( .A(n36308), .B(n36307), .Z(n36399) );
  XNOR U36720 ( .A(n36398), .B(n36399), .Z(n36400) );
  XNOR U36721 ( .A(n36401), .B(n36400), .Z(n36410) );
  XNOR U36722 ( .A(n36383), .B(n36384), .Z(n36386) );
  NANDN U36723 ( .A(n985), .B(a[99]), .Z(n36385) );
  XNOR U36724 ( .A(n36386), .B(n36385), .Z(n36377) );
  NANDN U36725 ( .A(n36310), .B(n36309), .Z(n36313) );
  XNOR U36726 ( .A(n38463), .B(b[37]), .Z(n36417) );
  NAND U36727 ( .A(n36417), .B(n36311), .Z(n36312) );
  NAND U36728 ( .A(n36313), .B(n36312), .Z(n36378) );
  XNOR U36729 ( .A(n36377), .B(n36378), .Z(n36379) );
  NAND U36730 ( .A(n37802), .B(n36314), .Z(n36316) );
  XNOR U36731 ( .A(b[51]), .B(a[113]), .Z(n36460) );
  NANDN U36732 ( .A(n36460), .B(n37803), .Z(n36315) );
  AND U36733 ( .A(n36316), .B(n36315), .Z(n36380) );
  XNOR U36734 ( .A(n36379), .B(n36380), .Z(n36411) );
  XOR U36735 ( .A(n36410), .B(n36411), .Z(n36413) );
  XOR U36736 ( .A(n36412), .B(n36413), .Z(n36465) );
  XOR U36737 ( .A(n36466), .B(n36465), .Z(n36472) );
  NANDN U36738 ( .A(n36318), .B(n36317), .Z(n36322) );
  NAND U36739 ( .A(n36320), .B(n36319), .Z(n36321) );
  NAND U36740 ( .A(n36322), .B(n36321), .Z(n36469) );
  OR U36741 ( .A(n36324), .B(n36323), .Z(n36328) );
  NANDN U36742 ( .A(n36326), .B(n36325), .Z(n36327) );
  NAND U36743 ( .A(n36328), .B(n36327), .Z(n36470) );
  XNOR U36744 ( .A(n36469), .B(n36470), .Z(n36471) );
  XNOR U36745 ( .A(n36472), .B(n36471), .Z(n36354) );
  XOR U36746 ( .A(n36353), .B(n36354), .Z(n36356) );
  NANDN U36747 ( .A(n36330), .B(n36329), .Z(n36334) );
  NAND U36748 ( .A(n36332), .B(n36331), .Z(n36333) );
  NAND U36749 ( .A(n36334), .B(n36333), .Z(n36355) );
  XOR U36750 ( .A(n36356), .B(n36355), .Z(n36348) );
  XNOR U36751 ( .A(n36347), .B(n36348), .Z(n36349) );
  XNOR U36752 ( .A(n36350), .B(n36349), .Z(n36475) );
  XNOR U36753 ( .A(n36476), .B(n36475), .Z(n36478) );
  XOR U36754 ( .A(n36477), .B(n36478), .Z(n36344) );
  NAND U36755 ( .A(n36336), .B(n36335), .Z(n36340) );
  NAND U36756 ( .A(n36338), .B(n36337), .Z(n36339) );
  AND U36757 ( .A(n36340), .B(n36339), .Z(n36345) );
  XOR U36758 ( .A(n36344), .B(n36345), .Z(n36341) );
  XOR U36759 ( .A(n36346), .B(n36341), .Z(n36342) );
  XNOR U36760 ( .A(n36343), .B(n36342), .Z(c[227]) );
  NANDN U36761 ( .A(n36343), .B(n36342), .Z(n36600) );
  NANDN U36762 ( .A(n36348), .B(n36347), .Z(n36352) );
  NANDN U36763 ( .A(n36350), .B(n36349), .Z(n36351) );
  NAND U36764 ( .A(n36352), .B(n36351), .Z(n36598) );
  NANDN U36765 ( .A(n36354), .B(n36353), .Z(n36358) );
  OR U36766 ( .A(n36356), .B(n36355), .Z(n36357) );
  NAND U36767 ( .A(n36358), .B(n36357), .Z(n36596) );
  NAND U36768 ( .A(n36360), .B(n36359), .Z(n36364) );
  NAND U36769 ( .A(n36362), .B(n36361), .Z(n36363) );
  NAND U36770 ( .A(n36364), .B(n36363), .Z(n36488) );
  NANDN U36771 ( .A(n36366), .B(n36365), .Z(n36370) );
  NAND U36772 ( .A(n36368), .B(n36367), .Z(n36369) );
  NAND U36773 ( .A(n36370), .B(n36369), .Z(n36518) );
  NANDN U36774 ( .A(n36372), .B(n36371), .Z(n36376) );
  OR U36775 ( .A(n36374), .B(n36373), .Z(n36375) );
  NAND U36776 ( .A(n36376), .B(n36375), .Z(n36515) );
  NANDN U36777 ( .A(n36378), .B(n36377), .Z(n36382) );
  NAND U36778 ( .A(n36380), .B(n36379), .Z(n36381) );
  NAND U36779 ( .A(n36382), .B(n36381), .Z(n36500) );
  NAND U36780 ( .A(n36384), .B(n36383), .Z(n36388) );
  OR U36781 ( .A(n36386), .B(n36385), .Z(n36387) );
  AND U36782 ( .A(n36388), .B(n36387), .Z(n36525) );
  NAND U36783 ( .A(n37652), .B(n36389), .Z(n36391) );
  XOR U36784 ( .A(a[116]), .B(n979), .Z(n36535) );
  OR U36785 ( .A(n36535), .B(n37756), .Z(n36390) );
  NAND U36786 ( .A(n36391), .B(n36390), .Z(n36591) );
  XNOR U36787 ( .A(n38134), .B(b[45]), .Z(n36544) );
  NAND U36788 ( .A(n36544), .B(n37261), .Z(n36394) );
  NANDN U36789 ( .A(n36392), .B(n37262), .Z(n36393) );
  AND U36790 ( .A(n36394), .B(n36393), .Z(n36592) );
  XNOR U36791 ( .A(n36591), .B(n36592), .Z(n36594) );
  NAND U36792 ( .A(n36395), .B(n37469), .Z(n36397) );
  XOR U36793 ( .A(a[118]), .B(n978), .Z(n36547) );
  NANDN U36794 ( .A(n36547), .B(n37471), .Z(n36396) );
  NAND U36795 ( .A(n36397), .B(n36396), .Z(n36593) );
  XNOR U36796 ( .A(n36594), .B(n36593), .Z(n36526) );
  XNOR U36797 ( .A(n36525), .B(n36526), .Z(n36528) );
  NANDN U36798 ( .A(n36399), .B(n36398), .Z(n36403) );
  NAND U36799 ( .A(n36401), .B(n36400), .Z(n36402) );
  AND U36800 ( .A(n36403), .B(n36402), .Z(n36527) );
  XOR U36801 ( .A(n36528), .B(n36527), .Z(n36497) );
  NANDN U36802 ( .A(n36405), .B(n36404), .Z(n36409) );
  NAND U36803 ( .A(n36407), .B(n36406), .Z(n36408) );
  NAND U36804 ( .A(n36409), .B(n36408), .Z(n36498) );
  XOR U36805 ( .A(n36497), .B(n36498), .Z(n36499) );
  XNOR U36806 ( .A(n36500), .B(n36499), .Z(n36516) );
  XNOR U36807 ( .A(n36515), .B(n36516), .Z(n36517) );
  XNOR U36808 ( .A(n36518), .B(n36517), .Z(n36494) );
  NANDN U36809 ( .A(n36411), .B(n36410), .Z(n36415) );
  OR U36810 ( .A(n36413), .B(n36412), .Z(n36414) );
  NAND U36811 ( .A(n36415), .B(n36414), .Z(n36524) );
  XOR U36812 ( .A(n975), .B(n36580), .Z(n36419) );
  XNOR U36813 ( .A(b[36]), .B(b[35]), .Z(n36416) );
  NANDN U36814 ( .A(n36417), .B(n36416), .Z(n36418) );
  AND U36815 ( .A(n36419), .B(n36418), .Z(n36567) );
  AND U36816 ( .A(a[100]), .B(b[63]), .Z(n36687) );
  XOR U36817 ( .A(b[63]), .B(n36420), .Z(n36581) );
  NANDN U36818 ( .A(n36581), .B(n38422), .Z(n36423) );
  NANDN U36819 ( .A(n36421), .B(n38423), .Z(n36422) );
  AND U36820 ( .A(n36423), .B(n36422), .Z(n36566) );
  XOR U36821 ( .A(n36687), .B(n36566), .Z(n36568) );
  XOR U36822 ( .A(n36567), .B(n36568), .Z(n36512) );
  NAND U36823 ( .A(n36807), .B(n36424), .Z(n36426) );
  XNOR U36824 ( .A(n38321), .B(b[41]), .Z(n36574) );
  NANDN U36825 ( .A(n36905), .B(n36574), .Z(n36425) );
  NAND U36826 ( .A(n36426), .B(n36425), .Z(n36587) );
  NAND U36827 ( .A(n38326), .B(n36427), .Z(n36429) );
  XOR U36828 ( .A(n38400), .B(n36909), .Z(n36577) );
  NANDN U36829 ( .A(n38273), .B(n36577), .Z(n36428) );
  AND U36830 ( .A(n36429), .B(n36428), .Z(n36588) );
  XNOR U36831 ( .A(n36587), .B(n36588), .Z(n36589) );
  XOR U36832 ( .A(b[53]), .B(n37583), .Z(n36557) );
  NANDN U36833 ( .A(n36557), .B(n37940), .Z(n36432) );
  NANDN U36834 ( .A(n36430), .B(n37941), .Z(n36431) );
  AND U36835 ( .A(n36432), .B(n36431), .Z(n36590) );
  XNOR U36836 ( .A(n36589), .B(n36590), .Z(n36509) );
  NANDN U36837 ( .A(n36434), .B(n36433), .Z(n36438) );
  NAND U36838 ( .A(n36436), .B(n36435), .Z(n36437) );
  NAND U36839 ( .A(n36438), .B(n36437), .Z(n36510) );
  XOR U36840 ( .A(n36509), .B(n36510), .Z(n36511) );
  XNOR U36841 ( .A(n36512), .B(n36511), .Z(n36521) );
  NANDN U36842 ( .A(n36440), .B(n36439), .Z(n36444) );
  NAND U36843 ( .A(n36442), .B(n36441), .Z(n36443) );
  NAND U36844 ( .A(n36444), .B(n36443), .Z(n36506) );
  NAND U36845 ( .A(n38194), .B(n36445), .Z(n36447) );
  XNOR U36846 ( .A(n983), .B(a[108]), .Z(n36538) );
  NANDN U36847 ( .A(n965), .B(n36538), .Z(n36446) );
  NAND U36848 ( .A(n36447), .B(n36446), .Z(n36531) );
  XOR U36849 ( .A(a[122]), .B(n977), .Z(n36541) );
  NANDN U36850 ( .A(n36541), .B(n37068), .Z(n36450) );
  NANDN U36851 ( .A(n36448), .B(n37069), .Z(n36449) );
  AND U36852 ( .A(n36450), .B(n36449), .Z(n36532) );
  XNOR U36853 ( .A(n36531), .B(n36532), .Z(n36533) );
  XOR U36854 ( .A(b[55]), .B(n37336), .Z(n36571) );
  NANDN U36855 ( .A(n36571), .B(n38075), .Z(n36453) );
  NANDN U36856 ( .A(n36451), .B(n38073), .Z(n36452) );
  AND U36857 ( .A(n36453), .B(n36452), .Z(n36534) );
  XNOR U36858 ( .A(n36533), .B(n36534), .Z(n36504) );
  XOR U36859 ( .A(a[126]), .B(n976), .Z(n36554) );
  NANDN U36860 ( .A(n36554), .B(n36553), .Z(n36456) );
  NANDN U36861 ( .A(n36454), .B(n36643), .Z(n36455) );
  NAND U36862 ( .A(n36456), .B(n36455), .Z(n36563) );
  XOR U36863 ( .A(b[61]), .B(n36647), .Z(n36550) );
  OR U36864 ( .A(n36550), .B(n38371), .Z(n36459) );
  NANDN U36865 ( .A(n36457), .B(n38369), .Z(n36458) );
  NAND U36866 ( .A(n36459), .B(n36458), .Z(n36560) );
  XOR U36867 ( .A(n980), .B(n37873), .Z(n36584) );
  NAND U36868 ( .A(n36584), .B(n37803), .Z(n36462) );
  NANDN U36869 ( .A(n36460), .B(n37802), .Z(n36461) );
  AND U36870 ( .A(n36462), .B(n36461), .Z(n36561) );
  XNOR U36871 ( .A(n36560), .B(n36561), .Z(n36562) );
  XOR U36872 ( .A(n36563), .B(n36562), .Z(n36503) );
  XOR U36873 ( .A(n36504), .B(n36503), .Z(n36505) );
  XOR U36874 ( .A(n36506), .B(n36505), .Z(n36522) );
  XNOR U36875 ( .A(n36521), .B(n36522), .Z(n36523) );
  XNOR U36876 ( .A(n36524), .B(n36523), .Z(n36491) );
  NANDN U36877 ( .A(n36464), .B(n36463), .Z(n36468) );
  NANDN U36878 ( .A(n36466), .B(n36465), .Z(n36467) );
  NAND U36879 ( .A(n36468), .B(n36467), .Z(n36492) );
  XNOR U36880 ( .A(n36491), .B(n36492), .Z(n36493) );
  XOR U36881 ( .A(n36494), .B(n36493), .Z(n36485) );
  NANDN U36882 ( .A(n36470), .B(n36469), .Z(n36474) );
  NAND U36883 ( .A(n36472), .B(n36471), .Z(n36473) );
  NAND U36884 ( .A(n36474), .B(n36473), .Z(n36486) );
  XOR U36885 ( .A(n36485), .B(n36486), .Z(n36487) );
  XOR U36886 ( .A(n36488), .B(n36487), .Z(n36595) );
  XNOR U36887 ( .A(n36596), .B(n36595), .Z(n36597) );
  XNOR U36888 ( .A(n36598), .B(n36597), .Z(n36482) );
  NAND U36889 ( .A(n36476), .B(n36475), .Z(n36480) );
  NANDN U36890 ( .A(n36478), .B(n36477), .Z(n36479) );
  AND U36891 ( .A(n36480), .B(n36479), .Z(n36483) );
  XOR U36892 ( .A(n36482), .B(n36483), .Z(n36481) );
  XOR U36893 ( .A(n36484), .B(n36481), .Z(n36599) );
  XNOR U36894 ( .A(n36600), .B(n36599), .Z(c[228]) );
  OR U36895 ( .A(n36486), .B(n36485), .Z(n36490) );
  NAND U36896 ( .A(n36488), .B(n36487), .Z(n36489) );
  NAND U36897 ( .A(n36490), .B(n36489), .Z(n36729) );
  NANDN U36898 ( .A(n36492), .B(n36491), .Z(n36496) );
  NAND U36899 ( .A(n36494), .B(n36493), .Z(n36495) );
  NAND U36900 ( .A(n36496), .B(n36495), .Z(n36726) );
  OR U36901 ( .A(n36498), .B(n36497), .Z(n36502) );
  NAND U36902 ( .A(n36500), .B(n36499), .Z(n36501) );
  NAND U36903 ( .A(n36502), .B(n36501), .Z(n36711) );
  OR U36904 ( .A(n36504), .B(n36503), .Z(n36508) );
  NANDN U36905 ( .A(n36506), .B(n36505), .Z(n36507) );
  NAND U36906 ( .A(n36508), .B(n36507), .Z(n36708) );
  OR U36907 ( .A(n36510), .B(n36509), .Z(n36514) );
  NANDN U36908 ( .A(n36512), .B(n36511), .Z(n36513) );
  AND U36909 ( .A(n36514), .B(n36513), .Z(n36709) );
  XNOR U36910 ( .A(n36708), .B(n36709), .Z(n36710) );
  XNOR U36911 ( .A(n36711), .B(n36710), .Z(n36723) );
  NANDN U36912 ( .A(n36516), .B(n36515), .Z(n36520) );
  NAND U36913 ( .A(n36518), .B(n36517), .Z(n36519) );
  NAND U36914 ( .A(n36520), .B(n36519), .Z(n36720) );
  OR U36915 ( .A(n36526), .B(n36525), .Z(n36530) );
  OR U36916 ( .A(n36528), .B(n36527), .Z(n36529) );
  NAND U36917 ( .A(n36530), .B(n36529), .Z(n36608) );
  XNOR U36918 ( .A(a[117]), .B(b[49]), .Z(n36625) );
  OR U36919 ( .A(n36625), .B(n37756), .Z(n36537) );
  NANDN U36920 ( .A(n36535), .B(n37652), .Z(n36536) );
  NAND U36921 ( .A(n36537), .B(n36536), .Z(n36654) );
  XNOR U36922 ( .A(b[57]), .B(a[109]), .Z(n36699) );
  OR U36923 ( .A(n36699), .B(n965), .Z(n36540) );
  NAND U36924 ( .A(n36538), .B(n38194), .Z(n36539) );
  NAND U36925 ( .A(n36540), .B(n36539), .Z(n36651) );
  XNOR U36926 ( .A(a[123]), .B(b[43]), .Z(n36637) );
  NANDN U36927 ( .A(n36637), .B(n37068), .Z(n36543) );
  NANDN U36928 ( .A(n36541), .B(n37069), .Z(n36542) );
  AND U36929 ( .A(n36543), .B(n36542), .Z(n36652) );
  XNOR U36930 ( .A(n36651), .B(n36652), .Z(n36653) );
  XNOR U36931 ( .A(n36654), .B(n36653), .Z(n36678) );
  NAND U36932 ( .A(n37262), .B(n36544), .Z(n36546) );
  XOR U36933 ( .A(a[121]), .B(b[45]), .Z(n36696) );
  NAND U36934 ( .A(n37261), .B(n36696), .Z(n36545) );
  NAND U36935 ( .A(n36546), .B(n36545), .Z(n36676) );
  NANDN U36936 ( .A(n36547), .B(n37469), .Z(n36549) );
  XNOR U36937 ( .A(n38193), .B(b[47]), .Z(n36693) );
  NAND U36938 ( .A(n36693), .B(n37471), .Z(n36548) );
  AND U36939 ( .A(n36549), .B(n36548), .Z(n36675) );
  XNOR U36940 ( .A(n36676), .B(n36675), .Z(n36677) );
  XOR U36941 ( .A(n36678), .B(n36677), .Z(n36615) );
  XNOR U36942 ( .A(b[61]), .B(a[105]), .Z(n36622) );
  OR U36943 ( .A(n36622), .B(n38371), .Z(n36552) );
  NANDN U36944 ( .A(n36550), .B(n38369), .Z(n36551) );
  NAND U36945 ( .A(n36552), .B(n36551), .Z(n36672) );
  XOR U36946 ( .A(a[127]), .B(n976), .Z(n36644) );
  NANDN U36947 ( .A(n36644), .B(n36553), .Z(n36556) );
  NANDN U36948 ( .A(n36554), .B(n36643), .Z(n36555) );
  NAND U36949 ( .A(n36556), .B(n36555), .Z(n36669) );
  XNOR U36950 ( .A(b[53]), .B(a[113]), .Z(n36634) );
  NANDN U36951 ( .A(n36634), .B(n37940), .Z(n36559) );
  NANDN U36952 ( .A(n36557), .B(n37941), .Z(n36558) );
  AND U36953 ( .A(n36559), .B(n36558), .Z(n36670) );
  XNOR U36954 ( .A(n36669), .B(n36670), .Z(n36671) );
  XNOR U36955 ( .A(n36672), .B(n36671), .Z(n36613) );
  NANDN U36956 ( .A(n36561), .B(n36560), .Z(n36565) );
  NAND U36957 ( .A(n36563), .B(n36562), .Z(n36564) );
  NAND U36958 ( .A(n36565), .B(n36564), .Z(n36614) );
  XOR U36959 ( .A(n36613), .B(n36614), .Z(n36616) );
  XNOR U36960 ( .A(n36615), .B(n36616), .Z(n36714) );
  XOR U36961 ( .A(n36715), .B(n36714), .Z(n36717) );
  OR U36962 ( .A(n36687), .B(n36566), .Z(n36570) );
  NAND U36963 ( .A(n36568), .B(n36567), .Z(n36569) );
  NAND U36964 ( .A(n36570), .B(n36569), .Z(n36665) );
  XNOR U36965 ( .A(b[55]), .B(a[111]), .Z(n36631) );
  NANDN U36966 ( .A(n36631), .B(n38075), .Z(n36573) );
  NANDN U36967 ( .A(n36571), .B(n38073), .Z(n36572) );
  NAND U36968 ( .A(n36573), .B(n36572), .Z(n36684) );
  XOR U36969 ( .A(a[125]), .B(b[41]), .Z(n36640) );
  NANDN U36970 ( .A(n36905), .B(n36640), .Z(n36576) );
  NAND U36971 ( .A(n36574), .B(n36807), .Z(n36575) );
  NAND U36972 ( .A(n36576), .B(n36575), .Z(n36681) );
  NAND U36973 ( .A(n38326), .B(n36577), .Z(n36579) );
  XNOR U36974 ( .A(n38400), .B(a[107]), .Z(n36619) );
  NANDN U36975 ( .A(n38273), .B(n36619), .Z(n36578) );
  AND U36976 ( .A(n36579), .B(n36578), .Z(n36682) );
  XNOR U36977 ( .A(n36681), .B(n36682), .Z(n36683) );
  XNOR U36978 ( .A(n36684), .B(n36683), .Z(n36663) );
  NAND U36979 ( .A(b[37]), .B(n36580), .Z(n36688) );
  XNOR U36980 ( .A(n36688), .B(n36687), .Z(n36690) );
  NANDN U36981 ( .A(n985), .B(a[101]), .Z(n36689) );
  XNOR U36982 ( .A(n36690), .B(n36689), .Z(n36657) );
  XNOR U36983 ( .A(n985), .B(a[103]), .Z(n36648) );
  NAND U36984 ( .A(n36648), .B(n38422), .Z(n36583) );
  NANDN U36985 ( .A(n36581), .B(n38423), .Z(n36582) );
  NAND U36986 ( .A(n36583), .B(n36582), .Z(n36658) );
  XNOR U36987 ( .A(n36657), .B(n36658), .Z(n36659) );
  NAND U36988 ( .A(n37802), .B(n36584), .Z(n36586) );
  XOR U36989 ( .A(n980), .B(a[115]), .Z(n36628) );
  NANDN U36990 ( .A(n36628), .B(n37803), .Z(n36585) );
  AND U36991 ( .A(n36586), .B(n36585), .Z(n36660) );
  XNOR U36992 ( .A(n36659), .B(n36660), .Z(n36664) );
  XOR U36993 ( .A(n36663), .B(n36664), .Z(n36666) );
  XOR U36994 ( .A(n36665), .B(n36666), .Z(n36704) );
  XNOR U36995 ( .A(n36703), .B(n36702), .Z(n36705) );
  XOR U36996 ( .A(n36704), .B(n36705), .Z(n36716) );
  XOR U36997 ( .A(n36717), .B(n36716), .Z(n36607) );
  XNOR U36998 ( .A(n36608), .B(n36607), .Z(n36609) );
  XNOR U36999 ( .A(n36610), .B(n36609), .Z(n36721) );
  XNOR U37000 ( .A(n36720), .B(n36721), .Z(n36722) );
  XOR U37001 ( .A(n36723), .B(n36722), .Z(n36727) );
  XOR U37002 ( .A(n36726), .B(n36727), .Z(n36728) );
  XNOR U37003 ( .A(n36729), .B(n36728), .Z(n36601) );
  XOR U37004 ( .A(n36601), .B(n36602), .Z(n36604) );
  XNOR U37005 ( .A(n36603), .B(n36604), .Z(n36732) );
  NANDN U37006 ( .A(n36600), .B(n36599), .Z(n36733) );
  XNOR U37007 ( .A(n36732), .B(n36733), .Z(c[229]) );
  NANDN U37008 ( .A(n36602), .B(n36601), .Z(n36606) );
  NANDN U37009 ( .A(n36604), .B(n36603), .Z(n36605) );
  NAND U37010 ( .A(n36606), .B(n36605), .Z(n36737) );
  NANDN U37011 ( .A(n36608), .B(n36607), .Z(n36612) );
  NAND U37012 ( .A(n36610), .B(n36609), .Z(n36611) );
  NAND U37013 ( .A(n36612), .B(n36611), .Z(n36850) );
  NANDN U37014 ( .A(n36614), .B(n36613), .Z(n36618) );
  NANDN U37015 ( .A(n36616), .B(n36615), .Z(n36617) );
  NAND U37016 ( .A(n36618), .B(n36617), .Z(n36822) );
  NAND U37017 ( .A(n38326), .B(n36619), .Z(n36621) );
  XOR U37018 ( .A(n38400), .B(n37139), .Z(n36764) );
  NANDN U37019 ( .A(n38273), .B(n36764), .Z(n36620) );
  NAND U37020 ( .A(n36621), .B(n36620), .Z(n36794) );
  XOR U37021 ( .A(b[61]), .B(n36909), .Z(n36810) );
  OR U37022 ( .A(n36810), .B(n38371), .Z(n36624) );
  NANDN U37023 ( .A(n36622), .B(n38369), .Z(n36623) );
  NAND U37024 ( .A(n36624), .B(n36623), .Z(n36791) );
  XOR U37025 ( .A(n38143), .B(n979), .Z(n36773) );
  NANDN U37026 ( .A(n37756), .B(n36773), .Z(n36627) );
  NANDN U37027 ( .A(n36625), .B(n37652), .Z(n36626) );
  AND U37028 ( .A(n36627), .B(n36626), .Z(n36792) );
  XNOR U37029 ( .A(n36791), .B(n36792), .Z(n36793) );
  XNOR U37030 ( .A(n36794), .B(n36793), .Z(n36782) );
  NANDN U37031 ( .A(n36628), .B(n37802), .Z(n36630) );
  XOR U37032 ( .A(a[116]), .B(n980), .Z(n36776) );
  NANDN U37033 ( .A(n36776), .B(n37803), .Z(n36629) );
  NAND U37034 ( .A(n36630), .B(n36629), .Z(n36780) );
  XNOR U37035 ( .A(n982), .B(a[112]), .Z(n36816) );
  NAND U37036 ( .A(n38075), .B(n36816), .Z(n36633) );
  NANDN U37037 ( .A(n36631), .B(n38073), .Z(n36632) );
  AND U37038 ( .A(n36633), .B(n36632), .Z(n36779) );
  XNOR U37039 ( .A(n36780), .B(n36779), .Z(n36781) );
  XOR U37040 ( .A(n36782), .B(n36781), .Z(n36839) );
  XOR U37041 ( .A(n981), .B(n37873), .Z(n36803) );
  NAND U37042 ( .A(n36803), .B(n37940), .Z(n36636) );
  NANDN U37043 ( .A(n36634), .B(n37941), .Z(n36635) );
  NAND U37044 ( .A(n36636), .B(n36635), .Z(n36788) );
  XOR U37045 ( .A(a[124]), .B(n977), .Z(n36767) );
  NANDN U37046 ( .A(n36767), .B(n37068), .Z(n36639) );
  NANDN U37047 ( .A(n36637), .B(n37069), .Z(n36638) );
  NAND U37048 ( .A(n36639), .B(n36638), .Z(n36785) );
  XNOR U37049 ( .A(n987), .B(b[41]), .Z(n36806) );
  NANDN U37050 ( .A(n36905), .B(n36806), .Z(n36642) );
  NAND U37051 ( .A(n36640), .B(n36807), .Z(n36641) );
  AND U37052 ( .A(n36642), .B(n36641), .Z(n36786) );
  XNOR U37053 ( .A(n36785), .B(n36786), .Z(n36787) );
  XNOR U37054 ( .A(n36788), .B(n36787), .Z(n36837) );
  NANDN U37055 ( .A(n36644), .B(n36643), .Z(n36645) );
  NANDN U37056 ( .A(n36646), .B(n36645), .Z(n36798) );
  AND U37057 ( .A(a[102]), .B(b[63]), .Z(n36901) );
  XOR U37058 ( .A(b[63]), .B(n36647), .Z(n36813) );
  NANDN U37059 ( .A(n36813), .B(n38422), .Z(n36650) );
  NAND U37060 ( .A(n36648), .B(n38423), .Z(n36649) );
  AND U37061 ( .A(n36650), .B(n36649), .Z(n36797) );
  XOR U37062 ( .A(n36901), .B(n36797), .Z(n36799) );
  XOR U37063 ( .A(n36798), .B(n36799), .Z(n36838) );
  XOR U37064 ( .A(n36837), .B(n36838), .Z(n36840) );
  XOR U37065 ( .A(n36839), .B(n36840), .Z(n36825) );
  NANDN U37066 ( .A(n36652), .B(n36651), .Z(n36656) );
  NAND U37067 ( .A(n36654), .B(n36653), .Z(n36655) );
  AND U37068 ( .A(n36656), .B(n36655), .Z(n36826) );
  XNOR U37069 ( .A(n36825), .B(n36826), .Z(n36827) );
  NANDN U37070 ( .A(n36658), .B(n36657), .Z(n36662) );
  NAND U37071 ( .A(n36660), .B(n36659), .Z(n36661) );
  NAND U37072 ( .A(n36662), .B(n36661), .Z(n36828) );
  XOR U37073 ( .A(n36827), .B(n36828), .Z(n36819) );
  NANDN U37074 ( .A(n36664), .B(n36663), .Z(n36668) );
  OR U37075 ( .A(n36666), .B(n36665), .Z(n36667) );
  AND U37076 ( .A(n36668), .B(n36667), .Z(n36820) );
  XNOR U37077 ( .A(n36819), .B(n36820), .Z(n36821) );
  XNOR U37078 ( .A(n36822), .B(n36821), .Z(n36743) );
  NANDN U37079 ( .A(n36670), .B(n36669), .Z(n36674) );
  NAND U37080 ( .A(n36672), .B(n36671), .Z(n36673) );
  NAND U37081 ( .A(n36674), .B(n36673), .Z(n36746) );
  NANDN U37082 ( .A(n36676), .B(n36675), .Z(n36680) );
  NAND U37083 ( .A(n36678), .B(n36677), .Z(n36679) );
  NAND U37084 ( .A(n36680), .B(n36679), .Z(n36747) );
  XNOR U37085 ( .A(n36746), .B(n36747), .Z(n36748) );
  NANDN U37086 ( .A(n36682), .B(n36681), .Z(n36686) );
  NAND U37087 ( .A(n36684), .B(n36683), .Z(n36685) );
  NAND U37088 ( .A(n36686), .B(n36685), .Z(n36831) );
  NAND U37089 ( .A(n36688), .B(n36687), .Z(n36692) );
  OR U37090 ( .A(n36690), .B(n36689), .Z(n36691) );
  AND U37091 ( .A(n36692), .B(n36691), .Z(n36832) );
  XNOR U37092 ( .A(n36831), .B(n36832), .Z(n36833) );
  NAND U37093 ( .A(n36693), .B(n37469), .Z(n36695) );
  XOR U37094 ( .A(n38134), .B(n978), .Z(n36758) );
  NAND U37095 ( .A(n36758), .B(n37471), .Z(n36694) );
  NAND U37096 ( .A(n36695), .B(n36694), .Z(n36755) );
  XNOR U37097 ( .A(n38251), .B(b[45]), .Z(n36770) );
  NAND U37098 ( .A(n36770), .B(n37261), .Z(n36698) );
  NAND U37099 ( .A(n36696), .B(n37262), .Z(n36697) );
  NAND U37100 ( .A(n36698), .B(n36697), .Z(n36752) );
  XOR U37101 ( .A(b[57]), .B(n37336), .Z(n36761) );
  OR U37102 ( .A(n36761), .B(n965), .Z(n36701) );
  NANDN U37103 ( .A(n36699), .B(n38194), .Z(n36700) );
  AND U37104 ( .A(n36701), .B(n36700), .Z(n36753) );
  XNOR U37105 ( .A(n36752), .B(n36753), .Z(n36754) );
  XOR U37106 ( .A(n36755), .B(n36754), .Z(n36834) );
  XOR U37107 ( .A(n36833), .B(n36834), .Z(n36749) );
  XOR U37108 ( .A(n36748), .B(n36749), .Z(n36740) );
  OR U37109 ( .A(n36703), .B(n36702), .Z(n36707) );
  NANDN U37110 ( .A(n36705), .B(n36704), .Z(n36706) );
  AND U37111 ( .A(n36707), .B(n36706), .Z(n36741) );
  XNOR U37112 ( .A(n36740), .B(n36741), .Z(n36742) );
  XNOR U37113 ( .A(n36743), .B(n36742), .Z(n36846) );
  NANDN U37114 ( .A(n36709), .B(n36708), .Z(n36713) );
  NAND U37115 ( .A(n36711), .B(n36710), .Z(n36712) );
  NAND U37116 ( .A(n36713), .B(n36712), .Z(n36844) );
  NANDN U37117 ( .A(n36715), .B(n36714), .Z(n36719) );
  OR U37118 ( .A(n36717), .B(n36716), .Z(n36718) );
  AND U37119 ( .A(n36719), .B(n36718), .Z(n36843) );
  XNOR U37120 ( .A(n36844), .B(n36843), .Z(n36845) );
  XOR U37121 ( .A(n36846), .B(n36845), .Z(n36849) );
  XNOR U37122 ( .A(n36850), .B(n36849), .Z(n36851) );
  NANDN U37123 ( .A(n36721), .B(n36720), .Z(n36725) );
  NANDN U37124 ( .A(n36723), .B(n36722), .Z(n36724) );
  AND U37125 ( .A(n36725), .B(n36724), .Z(n36852) );
  XNOR U37126 ( .A(n36851), .B(n36852), .Z(n36735) );
  OR U37127 ( .A(n36727), .B(n36726), .Z(n36731) );
  NAND U37128 ( .A(n36729), .B(n36728), .Z(n36730) );
  AND U37129 ( .A(n36731), .B(n36730), .Z(n36734) );
  XNOR U37130 ( .A(n36735), .B(n36734), .Z(n36736) );
  XNOR U37131 ( .A(n36737), .B(n36736), .Z(n36856) );
  NANDN U37132 ( .A(n36733), .B(n36732), .Z(n36855) );
  XOR U37133 ( .A(n36856), .B(n36855), .Z(c[230]) );
  NANDN U37134 ( .A(n36735), .B(n36734), .Z(n36739) );
  NAND U37135 ( .A(n36737), .B(n36736), .Z(n36738) );
  NAND U37136 ( .A(n36739), .B(n36738), .Z(n36860) );
  OR U37137 ( .A(n36741), .B(n36740), .Z(n36745) );
  OR U37138 ( .A(n36743), .B(n36742), .Z(n36744) );
  NAND U37139 ( .A(n36745), .B(n36744), .Z(n36970) );
  NANDN U37140 ( .A(n36747), .B(n36746), .Z(n36751) );
  NAND U37141 ( .A(n36749), .B(n36748), .Z(n36750) );
  NAND U37142 ( .A(n36751), .B(n36750), .Z(n36964) );
  NANDN U37143 ( .A(n36753), .B(n36752), .Z(n36757) );
  NAND U37144 ( .A(n36755), .B(n36754), .Z(n36756) );
  NAND U37145 ( .A(n36757), .B(n36756), .Z(n36888) );
  NAND U37146 ( .A(n37469), .B(n36758), .Z(n36760) );
  XNOR U37147 ( .A(a[121]), .B(n978), .Z(n36916) );
  NAND U37148 ( .A(n36916), .B(n37471), .Z(n36759) );
  NAND U37149 ( .A(n36760), .B(n36759), .Z(n36875) );
  XNOR U37150 ( .A(n983), .B(a[111]), .Z(n36922) );
  NANDN U37151 ( .A(n965), .B(n36922), .Z(n36763) );
  NANDN U37152 ( .A(n36761), .B(n38194), .Z(n36762) );
  NAND U37153 ( .A(n36763), .B(n36762), .Z(n36896) );
  NAND U37154 ( .A(n38326), .B(n36764), .Z(n36766) );
  XNOR U37155 ( .A(b[59]), .B(a[109]), .Z(n36925) );
  OR U37156 ( .A(n36925), .B(n38273), .Z(n36765) );
  NAND U37157 ( .A(n36766), .B(n36765), .Z(n36893) );
  XNOR U37158 ( .A(a[125]), .B(b[43]), .Z(n36945) );
  NANDN U37159 ( .A(n36945), .B(n37068), .Z(n36769) );
  NANDN U37160 ( .A(n36767), .B(n37069), .Z(n36768) );
  AND U37161 ( .A(n36769), .B(n36768), .Z(n36894) );
  XNOR U37162 ( .A(n36893), .B(n36894), .Z(n36895) );
  XNOR U37163 ( .A(n36896), .B(n36895), .Z(n36876) );
  XNOR U37164 ( .A(n36875), .B(n36876), .Z(n36877) );
  NAND U37165 ( .A(n37262), .B(n36770), .Z(n36772) );
  XOR U37166 ( .A(a[123]), .B(b[45]), .Z(n36913) );
  NAND U37167 ( .A(n37261), .B(n36913), .Z(n36771) );
  NAND U37168 ( .A(n36772), .B(n36771), .Z(n36940) );
  NAND U37169 ( .A(n37652), .B(n36773), .Z(n36775) );
  XOR U37170 ( .A(n38193), .B(b[49]), .Z(n36931) );
  OR U37171 ( .A(n36931), .B(n37756), .Z(n36774) );
  NAND U37172 ( .A(n36775), .B(n36774), .Z(n36938) );
  XNOR U37173 ( .A(b[51]), .B(a[117]), .Z(n36919) );
  NANDN U37174 ( .A(n36919), .B(n37803), .Z(n36778) );
  NANDN U37175 ( .A(n36776), .B(n37802), .Z(n36777) );
  AND U37176 ( .A(n36778), .B(n36777), .Z(n36939) );
  XNOR U37177 ( .A(n36938), .B(n36939), .Z(n36941) );
  XNOR U37178 ( .A(n36940), .B(n36941), .Z(n36878) );
  XNOR U37179 ( .A(n36877), .B(n36878), .Z(n36887) );
  XNOR U37180 ( .A(n36888), .B(n36887), .Z(n36890) );
  NANDN U37181 ( .A(n36780), .B(n36779), .Z(n36784) );
  NAND U37182 ( .A(n36782), .B(n36781), .Z(n36783) );
  AND U37183 ( .A(n36784), .B(n36783), .Z(n36889) );
  XNOR U37184 ( .A(n36890), .B(n36889), .Z(n36961) );
  NANDN U37185 ( .A(n36786), .B(n36785), .Z(n36790) );
  NAND U37186 ( .A(n36788), .B(n36787), .Z(n36789) );
  NAND U37187 ( .A(n36790), .B(n36789), .Z(n36872) );
  NANDN U37188 ( .A(n36792), .B(n36791), .Z(n36796) );
  NAND U37189 ( .A(n36794), .B(n36793), .Z(n36795) );
  NAND U37190 ( .A(n36796), .B(n36795), .Z(n36869) );
  OR U37191 ( .A(n36901), .B(n36797), .Z(n36801) );
  NAND U37192 ( .A(n36799), .B(n36798), .Z(n36800) );
  NAND U37193 ( .A(n36801), .B(n36800), .Z(n36884) );
  NANDN U37194 ( .A(n975), .B(b[38]), .Z(n36802) );
  AND U37195 ( .A(n36802), .B(b[39]), .Z(n36899) );
  NANDN U37196 ( .A(n985), .B(a[103]), .Z(n36900) );
  XOR U37197 ( .A(n36899), .B(n36900), .Z(n36902) );
  XNOR U37198 ( .A(n36901), .B(n36902), .Z(n36954) );
  NAND U37199 ( .A(n37941), .B(n36803), .Z(n36805) );
  XNOR U37200 ( .A(b[53]), .B(a[115]), .Z(n36942) );
  NANDN U37201 ( .A(n36942), .B(n37940), .Z(n36804) );
  NAND U37202 ( .A(n36805), .B(n36804), .Z(n36951) );
  NAND U37203 ( .A(n36807), .B(n36806), .Z(n36809) );
  XNOR U37204 ( .A(n38463), .B(b[41]), .Z(n36906) );
  NANDN U37205 ( .A(n36905), .B(n36906), .Z(n36808) );
  NAND U37206 ( .A(n36809), .B(n36808), .Z(n36952) );
  XNOR U37207 ( .A(n36951), .B(n36952), .Z(n36953) );
  XOR U37208 ( .A(n36954), .B(n36953), .Z(n36881) );
  NANDN U37209 ( .A(n36810), .B(n38369), .Z(n36812) );
  XNOR U37210 ( .A(n984), .B(a[107]), .Z(n36948) );
  NANDN U37211 ( .A(n38371), .B(n36948), .Z(n36811) );
  NAND U37212 ( .A(n36812), .B(n36811), .Z(n36936) );
  XNOR U37213 ( .A(n985), .B(a[105]), .Z(n36910) );
  NAND U37214 ( .A(n36910), .B(n38422), .Z(n36815) );
  NANDN U37215 ( .A(n36813), .B(n38423), .Z(n36814) );
  NAND U37216 ( .A(n36815), .B(n36814), .Z(n36934) );
  XNOR U37217 ( .A(b[55]), .B(a[113]), .Z(n36928) );
  NANDN U37218 ( .A(n36928), .B(n38075), .Z(n36818) );
  NAND U37219 ( .A(n36816), .B(n38073), .Z(n36817) );
  AND U37220 ( .A(n36818), .B(n36817), .Z(n36935) );
  XNOR U37221 ( .A(n36934), .B(n36935), .Z(n36937) );
  XNOR U37222 ( .A(n36936), .B(n36937), .Z(n36882) );
  XNOR U37223 ( .A(n36881), .B(n36882), .Z(n36883) );
  XNOR U37224 ( .A(n36884), .B(n36883), .Z(n36870) );
  XNOR U37225 ( .A(n36869), .B(n36870), .Z(n36871) );
  XOR U37226 ( .A(n36872), .B(n36871), .Z(n36962) );
  XOR U37227 ( .A(n36961), .B(n36962), .Z(n36963) );
  XNOR U37228 ( .A(n36964), .B(n36963), .Z(n36864) );
  NANDN U37229 ( .A(n36820), .B(n36819), .Z(n36824) );
  NAND U37230 ( .A(n36822), .B(n36821), .Z(n36823) );
  AND U37231 ( .A(n36824), .B(n36823), .Z(n36863) );
  XNOR U37232 ( .A(n36864), .B(n36863), .Z(n36865) );
  NANDN U37233 ( .A(n36826), .B(n36825), .Z(n36830) );
  NANDN U37234 ( .A(n36828), .B(n36827), .Z(n36829) );
  NAND U37235 ( .A(n36830), .B(n36829), .Z(n36958) );
  NANDN U37236 ( .A(n36832), .B(n36831), .Z(n36836) );
  NAND U37237 ( .A(n36834), .B(n36833), .Z(n36835) );
  NAND U37238 ( .A(n36836), .B(n36835), .Z(n36955) );
  NANDN U37239 ( .A(n36838), .B(n36837), .Z(n36842) );
  NANDN U37240 ( .A(n36840), .B(n36839), .Z(n36841) );
  NAND U37241 ( .A(n36842), .B(n36841), .Z(n36956) );
  XNOR U37242 ( .A(n36955), .B(n36956), .Z(n36957) );
  XNOR U37243 ( .A(n36958), .B(n36957), .Z(n36866) );
  XOR U37244 ( .A(n36865), .B(n36866), .Z(n36967) );
  NANDN U37245 ( .A(n36844), .B(n36843), .Z(n36848) );
  NAND U37246 ( .A(n36846), .B(n36845), .Z(n36847) );
  NAND U37247 ( .A(n36848), .B(n36847), .Z(n36968) );
  XNOR U37248 ( .A(n36967), .B(n36968), .Z(n36969) );
  XNOR U37249 ( .A(n36970), .B(n36969), .Z(n36857) );
  NANDN U37250 ( .A(n36850), .B(n36849), .Z(n36854) );
  NAND U37251 ( .A(n36852), .B(n36851), .Z(n36853) );
  AND U37252 ( .A(n36854), .B(n36853), .Z(n36858) );
  XNOR U37253 ( .A(n36857), .B(n36858), .Z(n36859) );
  XNOR U37254 ( .A(n36860), .B(n36859), .Z(n36974) );
  OR U37255 ( .A(n36856), .B(n36855), .Z(n36973) );
  XOR U37256 ( .A(n36974), .B(n36973), .Z(c[231]) );
  NANDN U37257 ( .A(n36858), .B(n36857), .Z(n36862) );
  NAND U37258 ( .A(n36860), .B(n36859), .Z(n36861) );
  NAND U37259 ( .A(n36862), .B(n36861), .Z(n36980) );
  NANDN U37260 ( .A(n36864), .B(n36863), .Z(n36868) );
  NANDN U37261 ( .A(n36866), .B(n36865), .Z(n36867) );
  NAND U37262 ( .A(n36868), .B(n36867), .Z(n36986) );
  NANDN U37263 ( .A(n36870), .B(n36869), .Z(n36874) );
  NAND U37264 ( .A(n36872), .B(n36871), .Z(n36873) );
  NAND U37265 ( .A(n36874), .B(n36873), .Z(n36998) );
  NANDN U37266 ( .A(n36876), .B(n36875), .Z(n36880) );
  NANDN U37267 ( .A(n36878), .B(n36877), .Z(n36879) );
  NAND U37268 ( .A(n36880), .B(n36879), .Z(n36995) );
  NANDN U37269 ( .A(n36882), .B(n36881), .Z(n36886) );
  NAND U37270 ( .A(n36884), .B(n36883), .Z(n36885) );
  AND U37271 ( .A(n36886), .B(n36885), .Z(n36996) );
  XNOR U37272 ( .A(n36995), .B(n36996), .Z(n36997) );
  XNOR U37273 ( .A(n36998), .B(n36997), .Z(n36992) );
  NAND U37274 ( .A(n36888), .B(n36887), .Z(n36892) );
  NANDN U37275 ( .A(n36890), .B(n36889), .Z(n36891) );
  NAND U37276 ( .A(n36892), .B(n36891), .Z(n37085) );
  NANDN U37277 ( .A(n36894), .B(n36893), .Z(n36898) );
  NAND U37278 ( .A(n36896), .B(n36895), .Z(n36897) );
  NAND U37279 ( .A(n36898), .B(n36897), .Z(n37053) );
  OR U37280 ( .A(n36900), .B(n36899), .Z(n36904) );
  NAND U37281 ( .A(n36902), .B(n36901), .Z(n36903) );
  NAND U37282 ( .A(n36904), .B(n36903), .Z(n37051) );
  NANDN U37283 ( .A(n976), .B(b[40]), .Z(n37032) );
  XNOR U37284 ( .A(b[41]), .B(n37032), .Z(n36908) );
  NANDN U37285 ( .A(n36906), .B(n36905), .Z(n36907) );
  AND U37286 ( .A(n36908), .B(n36907), .Z(n37045) );
  AND U37287 ( .A(b[63]), .B(a[104]), .Z(n37106) );
  XOR U37288 ( .A(n37045), .B(n37106), .Z(n37047) );
  XOR U37289 ( .A(b[63]), .B(n36909), .Z(n37033) );
  NANDN U37290 ( .A(n37033), .B(n38422), .Z(n36912) );
  NAND U37291 ( .A(n36910), .B(n38423), .Z(n36911) );
  AND U37292 ( .A(n36912), .B(n36911), .Z(n37046) );
  XOR U37293 ( .A(n37051), .B(n37050), .Z(n37052) );
  XNOR U37294 ( .A(n37053), .B(n37052), .Z(n37014) );
  XNOR U37295 ( .A(a[124]), .B(b[45]), .Z(n37065) );
  NANDN U37296 ( .A(n37065), .B(n37261), .Z(n36915) );
  NAND U37297 ( .A(n36913), .B(n37262), .Z(n36914) );
  NAND U37298 ( .A(n36915), .B(n36914), .Z(n37059) );
  NAND U37299 ( .A(n37469), .B(n36916), .Z(n36918) );
  XOR U37300 ( .A(n38251), .B(n978), .Z(n37079) );
  NAND U37301 ( .A(n37079), .B(n37471), .Z(n36917) );
  NAND U37302 ( .A(n36918), .B(n36917), .Z(n37056) );
  XOR U37303 ( .A(a[118]), .B(n980), .Z(n37023) );
  NANDN U37304 ( .A(n37023), .B(n37803), .Z(n36921) );
  NANDN U37305 ( .A(n36919), .B(n37802), .Z(n36920) );
  AND U37306 ( .A(n36921), .B(n36920), .Z(n37057) );
  XNOR U37307 ( .A(n37056), .B(n37057), .Z(n37058) );
  XNOR U37308 ( .A(n37059), .B(n37058), .Z(n37010) );
  XOR U37309 ( .A(b[57]), .B(n37583), .Z(n37026) );
  OR U37310 ( .A(n37026), .B(n965), .Z(n36924) );
  NAND U37311 ( .A(n36922), .B(n38194), .Z(n36923) );
  NAND U37312 ( .A(n36924), .B(n36923), .Z(n37042) );
  NANDN U37313 ( .A(n36925), .B(n38326), .Z(n36927) );
  XOR U37314 ( .A(n38400), .B(n37336), .Z(n37029) );
  NANDN U37315 ( .A(n38273), .B(n37029), .Z(n36926) );
  NAND U37316 ( .A(n36927), .B(n36926), .Z(n37039) );
  XOR U37317 ( .A(b[55]), .B(n37873), .Z(n37062) );
  NANDN U37318 ( .A(n37062), .B(n38075), .Z(n36930) );
  NANDN U37319 ( .A(n36928), .B(n38073), .Z(n36929) );
  AND U37320 ( .A(n36930), .B(n36929), .Z(n37040) );
  XNOR U37321 ( .A(n37039), .B(n37040), .Z(n37041) );
  XNOR U37322 ( .A(n37042), .B(n37041), .Z(n37007) );
  NANDN U37323 ( .A(n36931), .B(n37652), .Z(n36933) );
  XOR U37324 ( .A(a[120]), .B(n979), .Z(n37076) );
  OR U37325 ( .A(n37076), .B(n37756), .Z(n36932) );
  NAND U37326 ( .A(n36933), .B(n36932), .Z(n37008) );
  XNOR U37327 ( .A(n37007), .B(n37008), .Z(n37009) );
  XOR U37328 ( .A(n37010), .B(n37009), .Z(n37011) );
  XOR U37329 ( .A(n37011), .B(n37012), .Z(n37013) );
  XOR U37330 ( .A(n37014), .B(n37013), .Z(n37083) );
  XOR U37331 ( .A(n981), .B(n38046), .Z(n37036) );
  NAND U37332 ( .A(n37036), .B(n37940), .Z(n36944) );
  NANDN U37333 ( .A(n36942), .B(n37941), .Z(n36943) );
  NAND U37334 ( .A(n36944), .B(n36943), .Z(n37020) );
  XOR U37335 ( .A(a[126]), .B(n977), .Z(n37070) );
  NANDN U37336 ( .A(n37070), .B(n37068), .Z(n36947) );
  NANDN U37337 ( .A(n36945), .B(n37069), .Z(n36946) );
  NAND U37338 ( .A(n36947), .B(n36946), .Z(n37017) );
  XOR U37339 ( .A(b[61]), .B(n37139), .Z(n37073) );
  OR U37340 ( .A(n37073), .B(n38371), .Z(n36950) );
  NAND U37341 ( .A(n36948), .B(n38369), .Z(n36949) );
  AND U37342 ( .A(n36950), .B(n36949), .Z(n37018) );
  XNOR U37343 ( .A(n37017), .B(n37018), .Z(n37019) );
  XNOR U37344 ( .A(n37020), .B(n37019), .Z(n37001) );
  XOR U37345 ( .A(n37001), .B(n37002), .Z(n37004) );
  XOR U37346 ( .A(n37003), .B(n37004), .Z(n37082) );
  XOR U37347 ( .A(n37083), .B(n37082), .Z(n37084) );
  XNOR U37348 ( .A(n37085), .B(n37084), .Z(n36989) );
  NANDN U37349 ( .A(n36956), .B(n36955), .Z(n36960) );
  NAND U37350 ( .A(n36958), .B(n36957), .Z(n36959) );
  NAND U37351 ( .A(n36960), .B(n36959), .Z(n36990) );
  XNOR U37352 ( .A(n36989), .B(n36990), .Z(n36991) );
  XOR U37353 ( .A(n36992), .B(n36991), .Z(n36984) );
  NAND U37354 ( .A(n36962), .B(n36961), .Z(n36966) );
  NAND U37355 ( .A(n36964), .B(n36963), .Z(n36965) );
  AND U37356 ( .A(n36966), .B(n36965), .Z(n36983) );
  XOR U37357 ( .A(n36984), .B(n36983), .Z(n36985) );
  XNOR U37358 ( .A(n36986), .B(n36985), .Z(n36978) );
  NANDN U37359 ( .A(n36968), .B(n36967), .Z(n36972) );
  NAND U37360 ( .A(n36970), .B(n36969), .Z(n36971) );
  AND U37361 ( .A(n36972), .B(n36971), .Z(n36977) );
  XNOR U37362 ( .A(n36978), .B(n36977), .Z(n36979) );
  XNOR U37363 ( .A(n36980), .B(n36979), .Z(n36976) );
  OR U37364 ( .A(n36974), .B(n36973), .Z(n36975) );
  XOR U37365 ( .A(n36976), .B(n36975), .Z(c[232]) );
  OR U37366 ( .A(n36976), .B(n36975), .Z(n37197) );
  NANDN U37367 ( .A(n36978), .B(n36977), .Z(n36982) );
  NAND U37368 ( .A(n36980), .B(n36979), .Z(n36981) );
  NAND U37369 ( .A(n36982), .B(n36981), .Z(n37091) );
  OR U37370 ( .A(n36984), .B(n36983), .Z(n36988) );
  NAND U37371 ( .A(n36986), .B(n36985), .Z(n36987) );
  AND U37372 ( .A(n36988), .B(n36987), .Z(n37090) );
  NANDN U37373 ( .A(n36990), .B(n36989), .Z(n36994) );
  NAND U37374 ( .A(n36992), .B(n36991), .Z(n36993) );
  NAND U37375 ( .A(n36994), .B(n36993), .Z(n37195) );
  NANDN U37376 ( .A(n36996), .B(n36995), .Z(n37000) );
  NAND U37377 ( .A(n36998), .B(n36997), .Z(n36999) );
  NAND U37378 ( .A(n37000), .B(n36999), .Z(n37092) );
  NANDN U37379 ( .A(n37002), .B(n37001), .Z(n37006) );
  OR U37380 ( .A(n37004), .B(n37003), .Z(n37005) );
  AND U37381 ( .A(n37006), .B(n37005), .Z(n37098) );
  XNOR U37382 ( .A(n37098), .B(n37099), .Z(n37100) );
  NAND U37383 ( .A(n37012), .B(n37011), .Z(n37016) );
  NAND U37384 ( .A(n37014), .B(n37013), .Z(n37015) );
  AND U37385 ( .A(n37016), .B(n37015), .Z(n37101) );
  XOR U37386 ( .A(n37092), .B(n37093), .Z(n37094) );
  NANDN U37387 ( .A(n37018), .B(n37017), .Z(n37022) );
  NAND U37388 ( .A(n37020), .B(n37019), .Z(n37021) );
  NAND U37389 ( .A(n37022), .B(n37021), .Z(n37130) );
  XOR U37390 ( .A(a[119]), .B(n980), .Z(n37149) );
  NANDN U37391 ( .A(n37149), .B(n37803), .Z(n37025) );
  NANDN U37392 ( .A(n37023), .B(n37802), .Z(n37024) );
  NAND U37393 ( .A(n37025), .B(n37024), .Z(n37179) );
  XNOR U37394 ( .A(b[57]), .B(a[113]), .Z(n37152) );
  OR U37395 ( .A(n37152), .B(n965), .Z(n37028) );
  NANDN U37396 ( .A(n37026), .B(n38194), .Z(n37027) );
  NAND U37397 ( .A(n37028), .B(n37027), .Z(n37176) );
  NAND U37398 ( .A(n38326), .B(n37029), .Z(n37031) );
  XNOR U37399 ( .A(n38400), .B(a[111]), .Z(n37158) );
  NANDN U37400 ( .A(n38273), .B(n37158), .Z(n37030) );
  AND U37401 ( .A(n37031), .B(n37030), .Z(n37177) );
  XNOR U37402 ( .A(n37176), .B(n37177), .Z(n37178) );
  XNOR U37403 ( .A(n37179), .B(n37178), .Z(n37128) );
  NAND U37404 ( .A(n37032), .B(b[41]), .Z(n37104) );
  NANDN U37405 ( .A(n985), .B(a[105]), .Z(n37105) );
  XOR U37406 ( .A(n37104), .B(n37105), .Z(n37107) );
  XNOR U37407 ( .A(n37106), .B(n37107), .Z(n37143) );
  XNOR U37408 ( .A(n985), .B(a[107]), .Z(n37140) );
  NAND U37409 ( .A(n37140), .B(n38422), .Z(n37035) );
  NANDN U37410 ( .A(n37033), .B(n38423), .Z(n37034) );
  NAND U37411 ( .A(n37035), .B(n37034), .Z(n37144) );
  XOR U37412 ( .A(n37143), .B(n37144), .Z(n37145) );
  NAND U37413 ( .A(n37941), .B(n37036), .Z(n37038) );
  XNOR U37414 ( .A(b[53]), .B(a[117]), .Z(n37155) );
  NANDN U37415 ( .A(n37155), .B(n37940), .Z(n37037) );
  AND U37416 ( .A(n37038), .B(n37037), .Z(n37146) );
  XNOR U37417 ( .A(n37145), .B(n37146), .Z(n37129) );
  XOR U37418 ( .A(n37128), .B(n37129), .Z(n37131) );
  XNOR U37419 ( .A(n37130), .B(n37131), .Z(n37188) );
  NANDN U37420 ( .A(n37040), .B(n37039), .Z(n37044) );
  NAND U37421 ( .A(n37042), .B(n37041), .Z(n37043) );
  AND U37422 ( .A(n37044), .B(n37043), .Z(n37186) );
  NANDN U37423 ( .A(n37106), .B(n37045), .Z(n37049) );
  OR U37424 ( .A(n37047), .B(n37046), .Z(n37048) );
  AND U37425 ( .A(n37049), .B(n37048), .Z(n37187) );
  XOR U37426 ( .A(n37188), .B(n37189), .Z(n37185) );
  NAND U37427 ( .A(n37051), .B(n37050), .Z(n37055) );
  NAND U37428 ( .A(n37053), .B(n37052), .Z(n37054) );
  NAND U37429 ( .A(n37055), .B(n37054), .Z(n37183) );
  NANDN U37430 ( .A(n37057), .B(n37056), .Z(n37061) );
  NAND U37431 ( .A(n37059), .B(n37058), .Z(n37060) );
  NAND U37432 ( .A(n37061), .B(n37060), .Z(n37125) );
  XNOR U37433 ( .A(b[55]), .B(a[115]), .Z(n37167) );
  NANDN U37434 ( .A(n37167), .B(n38075), .Z(n37064) );
  NANDN U37435 ( .A(n37062), .B(n38073), .Z(n37063) );
  NAND U37436 ( .A(n37064), .B(n37063), .Z(n37113) );
  XOR U37437 ( .A(a[125]), .B(b[45]), .Z(n37173) );
  NAND U37438 ( .A(n37173), .B(n37261), .Z(n37067) );
  NANDN U37439 ( .A(n37065), .B(n37262), .Z(n37066) );
  NAND U37440 ( .A(n37067), .B(n37066), .Z(n37110) );
  XNOR U37441 ( .A(n38463), .B(b[43]), .Z(n37136) );
  NAND U37442 ( .A(n37136), .B(n37068), .Z(n37072) );
  NANDN U37443 ( .A(n37070), .B(n37069), .Z(n37071) );
  AND U37444 ( .A(n37072), .B(n37071), .Z(n37111) );
  XNOR U37445 ( .A(n37110), .B(n37111), .Z(n37112) );
  XOR U37446 ( .A(n37113), .B(n37112), .Z(n37123) );
  XNOR U37447 ( .A(b[61]), .B(a[109]), .Z(n37161) );
  OR U37448 ( .A(n37161), .B(n38371), .Z(n37075) );
  NANDN U37449 ( .A(n37073), .B(n38369), .Z(n37074) );
  NAND U37450 ( .A(n37075), .B(n37074), .Z(n37119) );
  XNOR U37451 ( .A(a[121]), .B(b[49]), .Z(n37164) );
  OR U37452 ( .A(n37164), .B(n37756), .Z(n37078) );
  NANDN U37453 ( .A(n37076), .B(n37652), .Z(n37077) );
  NAND U37454 ( .A(n37078), .B(n37077), .Z(n37116) );
  NAND U37455 ( .A(n37469), .B(n37079), .Z(n37081) );
  XNOR U37456 ( .A(a[123]), .B(n978), .Z(n37170) );
  NAND U37457 ( .A(n37170), .B(n37471), .Z(n37080) );
  AND U37458 ( .A(n37081), .B(n37080), .Z(n37117) );
  XNOR U37459 ( .A(n37116), .B(n37117), .Z(n37118) );
  XNOR U37460 ( .A(n37119), .B(n37118), .Z(n37122) );
  XOR U37461 ( .A(n37123), .B(n37122), .Z(n37124) );
  XOR U37462 ( .A(n37125), .B(n37124), .Z(n37182) );
  XNOR U37463 ( .A(n37183), .B(n37182), .Z(n37184) );
  XOR U37464 ( .A(n37185), .B(n37184), .Z(n37095) );
  XNOR U37465 ( .A(n37094), .B(n37095), .Z(n37192) );
  OR U37466 ( .A(n37083), .B(n37082), .Z(n37087) );
  NAND U37467 ( .A(n37085), .B(n37084), .Z(n37086) );
  AND U37468 ( .A(n37087), .B(n37086), .Z(n37193) );
  XNOR U37469 ( .A(n37192), .B(n37193), .Z(n37194) );
  XNOR U37470 ( .A(n37195), .B(n37194), .Z(n37089) );
  XNOR U37471 ( .A(n37090), .B(n37089), .Z(n37088) );
  XOR U37472 ( .A(n37091), .B(n37088), .Z(n37196) );
  XNOR U37473 ( .A(n37197), .B(n37196), .Z(c[233]) );
  OR U37474 ( .A(n37093), .B(n37092), .Z(n37097) );
  NAND U37475 ( .A(n37095), .B(n37094), .Z(n37096) );
  NAND U37476 ( .A(n37097), .B(n37096), .Z(n37291) );
  OR U37477 ( .A(n37099), .B(n37098), .Z(n37103) );
  OR U37478 ( .A(n37101), .B(n37100), .Z(n37102) );
  AND U37479 ( .A(n37103), .B(n37102), .Z(n37292) );
  XNOR U37480 ( .A(n37291), .B(n37292), .Z(n37293) );
  NANDN U37481 ( .A(n37105), .B(n37104), .Z(n37109) );
  NANDN U37482 ( .A(n37107), .B(n37106), .Z(n37108) );
  NAND U37483 ( .A(n37109), .B(n37108), .Z(n37219) );
  NANDN U37484 ( .A(n37111), .B(n37110), .Z(n37115) );
  NAND U37485 ( .A(n37113), .B(n37112), .Z(n37114) );
  NAND U37486 ( .A(n37115), .B(n37114), .Z(n37217) );
  NANDN U37487 ( .A(n37117), .B(n37116), .Z(n37121) );
  NAND U37488 ( .A(n37119), .B(n37118), .Z(n37120) );
  AND U37489 ( .A(n37121), .B(n37120), .Z(n37216) );
  XNOR U37490 ( .A(n37217), .B(n37216), .Z(n37218) );
  XOR U37491 ( .A(n37219), .B(n37218), .Z(n37211) );
  NANDN U37492 ( .A(n37123), .B(n37122), .Z(n37127) );
  OR U37493 ( .A(n37125), .B(n37124), .Z(n37126) );
  AND U37494 ( .A(n37127), .B(n37126), .Z(n37210) );
  XNOR U37495 ( .A(n37211), .B(n37210), .Z(n37213) );
  NANDN U37496 ( .A(n37129), .B(n37128), .Z(n37133) );
  OR U37497 ( .A(n37131), .B(n37130), .Z(n37132) );
  NAND U37498 ( .A(n37133), .B(n37132), .Z(n37225) );
  XOR U37499 ( .A(n977), .B(n37134), .Z(n37138) );
  XNOR U37500 ( .A(b[42]), .B(b[41]), .Z(n37135) );
  NANDN U37501 ( .A(n37136), .B(n37135), .Z(n37137) );
  AND U37502 ( .A(n37138), .B(n37137), .Z(n37248) );
  AND U37503 ( .A(a[106]), .B(b[63]), .Z(n37367) );
  XOR U37504 ( .A(b[63]), .B(n37139), .Z(n37252) );
  NANDN U37505 ( .A(n37252), .B(n38422), .Z(n37142) );
  NAND U37506 ( .A(n37140), .B(n38423), .Z(n37141) );
  AND U37507 ( .A(n37142), .B(n37141), .Z(n37247) );
  XOR U37508 ( .A(n37367), .B(n37247), .Z(n37249) );
  XOR U37509 ( .A(n37248), .B(n37249), .Z(n37288) );
  OR U37510 ( .A(n37144), .B(n37143), .Z(n37148) );
  NAND U37511 ( .A(n37146), .B(n37145), .Z(n37147) );
  NAND U37512 ( .A(n37148), .B(n37147), .Z(n37285) );
  XOR U37513 ( .A(a[120]), .B(n980), .Z(n37232) );
  NANDN U37514 ( .A(n37232), .B(n37803), .Z(n37151) );
  NANDN U37515 ( .A(n37149), .B(n37802), .Z(n37150) );
  NAND U37516 ( .A(n37151), .B(n37150), .Z(n37272) );
  XOR U37517 ( .A(b[57]), .B(n37873), .Z(n37229) );
  OR U37518 ( .A(n37229), .B(n965), .Z(n37154) );
  NANDN U37519 ( .A(n37152), .B(n38194), .Z(n37153) );
  NAND U37520 ( .A(n37154), .B(n37153), .Z(n37269) );
  XOR U37521 ( .A(b[53]), .B(n38143), .Z(n37266) );
  NANDN U37522 ( .A(n37266), .B(n37940), .Z(n37157) );
  NANDN U37523 ( .A(n37155), .B(n37941), .Z(n37156) );
  AND U37524 ( .A(n37157), .B(n37156), .Z(n37270) );
  XNOR U37525 ( .A(n37269), .B(n37270), .Z(n37271) );
  XOR U37526 ( .A(n37272), .B(n37271), .Z(n37286) );
  XNOR U37527 ( .A(n37285), .B(n37286), .Z(n37287) );
  XNOR U37528 ( .A(n37288), .B(n37287), .Z(n37222) );
  NAND U37529 ( .A(n38326), .B(n37158), .Z(n37160) );
  XOR U37530 ( .A(b[59]), .B(n37583), .Z(n37226) );
  OR U37531 ( .A(n37226), .B(n38273), .Z(n37159) );
  NAND U37532 ( .A(n37160), .B(n37159), .Z(n37278) );
  XOR U37533 ( .A(b[61]), .B(n37336), .Z(n37258) );
  OR U37534 ( .A(n37258), .B(n38371), .Z(n37163) );
  NANDN U37535 ( .A(n37161), .B(n38369), .Z(n37162) );
  NAND U37536 ( .A(n37163), .B(n37162), .Z(n37275) );
  XOR U37537 ( .A(n38251), .B(n979), .Z(n37238) );
  NANDN U37538 ( .A(n37756), .B(n37238), .Z(n37166) );
  NANDN U37539 ( .A(n37164), .B(n37652), .Z(n37165) );
  AND U37540 ( .A(n37166), .B(n37165), .Z(n37276) );
  XNOR U37541 ( .A(n37275), .B(n37276), .Z(n37277) );
  XNOR U37542 ( .A(n37278), .B(n37277), .Z(n37281) );
  XOR U37543 ( .A(b[55]), .B(n38046), .Z(n37255) );
  NANDN U37544 ( .A(n37255), .B(n38075), .Z(n37169) );
  NANDN U37545 ( .A(n37167), .B(n38073), .Z(n37168) );
  NAND U37546 ( .A(n37169), .B(n37168), .Z(n37244) );
  NAND U37547 ( .A(n37469), .B(n37170), .Z(n37172) );
  XOR U37548 ( .A(a[124]), .B(n978), .Z(n37235) );
  NANDN U37549 ( .A(n37235), .B(n37471), .Z(n37171) );
  NAND U37550 ( .A(n37172), .B(n37171), .Z(n37241) );
  XNOR U37551 ( .A(a[126]), .B(b[45]), .Z(n37263) );
  NANDN U37552 ( .A(n37263), .B(n37261), .Z(n37175) );
  NAND U37553 ( .A(n37173), .B(n37262), .Z(n37174) );
  AND U37554 ( .A(n37175), .B(n37174), .Z(n37242) );
  XNOR U37555 ( .A(n37241), .B(n37242), .Z(n37243) );
  XOR U37556 ( .A(n37244), .B(n37243), .Z(n37282) );
  XNOR U37557 ( .A(n37281), .B(n37282), .Z(n37283) );
  NANDN U37558 ( .A(n37177), .B(n37176), .Z(n37181) );
  NAND U37559 ( .A(n37179), .B(n37178), .Z(n37180) );
  AND U37560 ( .A(n37181), .B(n37180), .Z(n37284) );
  XNOR U37561 ( .A(n37283), .B(n37284), .Z(n37223) );
  XNOR U37562 ( .A(n37222), .B(n37223), .Z(n37224) );
  XNOR U37563 ( .A(n37225), .B(n37224), .Z(n37212) );
  XNOR U37564 ( .A(n37213), .B(n37212), .Z(n37207) );
  OR U37565 ( .A(n37187), .B(n37186), .Z(n37191) );
  NANDN U37566 ( .A(n37189), .B(n37188), .Z(n37190) );
  NAND U37567 ( .A(n37191), .B(n37190), .Z(n37205) );
  XNOR U37568 ( .A(n37204), .B(n37205), .Z(n37206) );
  XOR U37569 ( .A(n37207), .B(n37206), .Z(n37294) );
  XOR U37570 ( .A(n37293), .B(n37294), .Z(n37198) );
  XNOR U37571 ( .A(n37198), .B(n37199), .Z(n37201) );
  XOR U37572 ( .A(n37200), .B(n37201), .Z(n37297) );
  NANDN U37573 ( .A(n37197), .B(n37196), .Z(n37298) );
  XNOR U37574 ( .A(n37297), .B(n37298), .Z(c[234]) );
  NANDN U37575 ( .A(n37199), .B(n37198), .Z(n37203) );
  NAND U37576 ( .A(n37201), .B(n37200), .Z(n37202) );
  NAND U37577 ( .A(n37203), .B(n37202), .Z(n37304) );
  NANDN U37578 ( .A(n37205), .B(n37204), .Z(n37209) );
  NANDN U37579 ( .A(n37207), .B(n37206), .Z(n37208) );
  NAND U37580 ( .A(n37209), .B(n37208), .Z(n37307) );
  OR U37581 ( .A(n37211), .B(n37210), .Z(n37215) );
  OR U37582 ( .A(n37213), .B(n37212), .Z(n37214) );
  AND U37583 ( .A(n37215), .B(n37214), .Z(n37308) );
  XNOR U37584 ( .A(n37307), .B(n37308), .Z(n37309) );
  NANDN U37585 ( .A(n37217), .B(n37216), .Z(n37221) );
  NANDN U37586 ( .A(n37219), .B(n37218), .Z(n37220) );
  NAND U37587 ( .A(n37221), .B(n37220), .Z(n37401) );
  NANDN U37588 ( .A(n37226), .B(n38326), .Z(n37228) );
  XNOR U37589 ( .A(b[59]), .B(a[113]), .Z(n37353) );
  OR U37590 ( .A(n37353), .B(n38273), .Z(n37227) );
  AND U37591 ( .A(n37228), .B(n37227), .Z(n37319) );
  XNOR U37592 ( .A(b[57]), .B(a[115]), .Z(n37377) );
  OR U37593 ( .A(n37377), .B(n965), .Z(n37231) );
  NANDN U37594 ( .A(n37229), .B(n38194), .Z(n37230) );
  AND U37595 ( .A(n37231), .B(n37230), .Z(n37320) );
  XOR U37596 ( .A(n37319), .B(n37320), .Z(n37321) );
  XNOR U37597 ( .A(a[121]), .B(n980), .Z(n37362) );
  NAND U37598 ( .A(n37362), .B(n37803), .Z(n37234) );
  NANDN U37599 ( .A(n37232), .B(n37802), .Z(n37233) );
  AND U37600 ( .A(n37234), .B(n37233), .Z(n37322) );
  XNOR U37601 ( .A(n37321), .B(n37322), .Z(n37347) );
  NANDN U37602 ( .A(n37235), .B(n37469), .Z(n37237) );
  XNOR U37603 ( .A(a[125]), .B(n978), .Z(n37374) );
  NAND U37604 ( .A(n37374), .B(n37471), .Z(n37236) );
  NAND U37605 ( .A(n37237), .B(n37236), .Z(n37345) );
  NAND U37606 ( .A(n37652), .B(n37238), .Z(n37240) );
  XNOR U37607 ( .A(a[123]), .B(b[49]), .Z(n37371) );
  OR U37608 ( .A(n37371), .B(n37756), .Z(n37239) );
  AND U37609 ( .A(n37240), .B(n37239), .Z(n37344) );
  XNOR U37610 ( .A(n37345), .B(n37344), .Z(n37346) );
  XOR U37611 ( .A(n37347), .B(n37346), .Z(n37388) );
  NANDN U37612 ( .A(n37242), .B(n37241), .Z(n37246) );
  NAND U37613 ( .A(n37244), .B(n37243), .Z(n37245) );
  AND U37614 ( .A(n37246), .B(n37245), .Z(n37386) );
  OR U37615 ( .A(n37367), .B(n37247), .Z(n37251) );
  NAND U37616 ( .A(n37249), .B(n37248), .Z(n37250) );
  NAND U37617 ( .A(n37251), .B(n37250), .Z(n37343) );
  XNOR U37618 ( .A(b[63]), .B(a[109]), .Z(n37337) );
  NANDN U37619 ( .A(n37337), .B(n38422), .Z(n37254) );
  NANDN U37620 ( .A(n37252), .B(n38423), .Z(n37253) );
  NAND U37621 ( .A(n37254), .B(n37253), .Z(n37325) );
  XNOR U37622 ( .A(b[55]), .B(a[117]), .Z(n37350) );
  NANDN U37623 ( .A(n37350), .B(n38075), .Z(n37257) );
  NANDN U37624 ( .A(n37255), .B(n38073), .Z(n37256) );
  AND U37625 ( .A(n37257), .B(n37256), .Z(n37326) );
  XNOR U37626 ( .A(n37325), .B(n37326), .Z(n37327) );
  NANDN U37627 ( .A(n985), .B(a[107]), .Z(n37366) );
  XOR U37628 ( .A(n37365), .B(n37366), .Z(n37368) );
  XOR U37629 ( .A(n37367), .B(n37368), .Z(n37328) );
  XNOR U37630 ( .A(n37327), .B(n37328), .Z(n37340) );
  XNOR U37631 ( .A(b[61]), .B(a[111]), .Z(n37356) );
  OR U37632 ( .A(n37356), .B(n38371), .Z(n37260) );
  NANDN U37633 ( .A(n37258), .B(n38369), .Z(n37259) );
  NAND U37634 ( .A(n37260), .B(n37259), .Z(n37383) );
  XNOR U37635 ( .A(n38463), .B(b[45]), .Z(n37333) );
  NAND U37636 ( .A(n37333), .B(n37261), .Z(n37265) );
  NANDN U37637 ( .A(n37263), .B(n37262), .Z(n37264) );
  NAND U37638 ( .A(n37265), .B(n37264), .Z(n37380) );
  XOR U37639 ( .A(n981), .B(n38193), .Z(n37359) );
  NAND U37640 ( .A(n37359), .B(n37940), .Z(n37268) );
  NANDN U37641 ( .A(n37266), .B(n37941), .Z(n37267) );
  AND U37642 ( .A(n37268), .B(n37267), .Z(n37381) );
  XNOR U37643 ( .A(n37380), .B(n37381), .Z(n37382) );
  XOR U37644 ( .A(n37383), .B(n37382), .Z(n37341) );
  XOR U37645 ( .A(n37340), .B(n37341), .Z(n37342) );
  XNOR U37646 ( .A(n37343), .B(n37342), .Z(n37387) );
  XNOR U37647 ( .A(n37386), .B(n37387), .Z(n37389) );
  XNOR U37648 ( .A(n37388), .B(n37389), .Z(n37313) );
  NANDN U37649 ( .A(n37270), .B(n37269), .Z(n37274) );
  NAND U37650 ( .A(n37272), .B(n37271), .Z(n37273) );
  NAND U37651 ( .A(n37274), .B(n37273), .Z(n37314) );
  XOR U37652 ( .A(n37313), .B(n37314), .Z(n37315) );
  NANDN U37653 ( .A(n37276), .B(n37275), .Z(n37280) );
  NAND U37654 ( .A(n37278), .B(n37277), .Z(n37279) );
  NAND U37655 ( .A(n37280), .B(n37279), .Z(n37316) );
  XOR U37656 ( .A(n37315), .B(n37316), .Z(n37395) );
  NANDN U37657 ( .A(n37286), .B(n37285), .Z(n37290) );
  NANDN U37658 ( .A(n37288), .B(n37287), .Z(n37289) );
  AND U37659 ( .A(n37290), .B(n37289), .Z(n37392) );
  XNOR U37660 ( .A(n37393), .B(n37392), .Z(n37394) );
  XOR U37661 ( .A(n37395), .B(n37394), .Z(n37399) );
  XNOR U37662 ( .A(n37398), .B(n37399), .Z(n37400) );
  XNOR U37663 ( .A(n37401), .B(n37400), .Z(n37310) );
  XOR U37664 ( .A(n37309), .B(n37310), .Z(n37301) );
  NANDN U37665 ( .A(n37292), .B(n37291), .Z(n37296) );
  NANDN U37666 ( .A(n37294), .B(n37293), .Z(n37295) );
  NAND U37667 ( .A(n37296), .B(n37295), .Z(n37302) );
  XNOR U37668 ( .A(n37301), .B(n37302), .Z(n37303) );
  XNOR U37669 ( .A(n37304), .B(n37303), .Z(n37300) );
  NANDN U37670 ( .A(n37298), .B(n37297), .Z(n37299) );
  XOR U37671 ( .A(n37300), .B(n37299), .Z(c[235]) );
  OR U37672 ( .A(n37300), .B(n37299), .Z(n37499) );
  NANDN U37673 ( .A(n37302), .B(n37301), .Z(n37306) );
  NAND U37674 ( .A(n37304), .B(n37303), .Z(n37305) );
  AND U37675 ( .A(n37306), .B(n37305), .Z(n37409) );
  NANDN U37676 ( .A(n37308), .B(n37307), .Z(n37312) );
  NANDN U37677 ( .A(n37310), .B(n37309), .Z(n37311) );
  AND U37678 ( .A(n37312), .B(n37311), .Z(n37406) );
  OR U37679 ( .A(n37314), .B(n37313), .Z(n37318) );
  NANDN U37680 ( .A(n37316), .B(n37315), .Z(n37317) );
  NAND U37681 ( .A(n37318), .B(n37317), .Z(n37493) );
  OR U37682 ( .A(n37320), .B(n37319), .Z(n37324) );
  NANDN U37683 ( .A(n37322), .B(n37321), .Z(n37323) );
  NAND U37684 ( .A(n37324), .B(n37323), .Z(n37482) );
  NANDN U37685 ( .A(n37326), .B(n37325), .Z(n37330) );
  NANDN U37686 ( .A(n37328), .B(n37327), .Z(n37329) );
  AND U37687 ( .A(n37330), .B(n37329), .Z(n37483) );
  XNOR U37688 ( .A(n37482), .B(n37483), .Z(n37484) );
  XNOR U37689 ( .A(b[45]), .B(n37331), .Z(n37335) );
  XOR U37690 ( .A(b[44]), .B(n977), .Z(n37332) );
  NANDN U37691 ( .A(n37333), .B(n37332), .Z(n37334) );
  AND U37692 ( .A(n37335), .B(n37334), .Z(n37478) );
  AND U37693 ( .A(a[108]), .B(b[63]), .Z(n37569) );
  XOR U37694 ( .A(b[63]), .B(n37336), .Z(n37430) );
  NANDN U37695 ( .A(n37430), .B(n38422), .Z(n37339) );
  NANDN U37696 ( .A(n37337), .B(n38423), .Z(n37338) );
  AND U37697 ( .A(n37339), .B(n37338), .Z(n37477) );
  XOR U37698 ( .A(n37569), .B(n37477), .Z(n37479) );
  XOR U37699 ( .A(n37478), .B(n37479), .Z(n37485) );
  XNOR U37700 ( .A(n37484), .B(n37485), .Z(n37488) );
  XNOR U37701 ( .A(n37488), .B(n37489), .Z(n37490) );
  NANDN U37702 ( .A(n37345), .B(n37344), .Z(n37349) );
  NANDN U37703 ( .A(n37347), .B(n37346), .Z(n37348) );
  NAND U37704 ( .A(n37349), .B(n37348), .Z(n37421) );
  XNOR U37705 ( .A(n982), .B(a[118]), .Z(n37424) );
  NAND U37706 ( .A(n38075), .B(n37424), .Z(n37352) );
  NANDN U37707 ( .A(n37350), .B(n38073), .Z(n37351) );
  AND U37708 ( .A(n37352), .B(n37351), .Z(n37465) );
  NANDN U37709 ( .A(n37353), .B(n38326), .Z(n37355) );
  XNOR U37710 ( .A(n38400), .B(a[114]), .Z(n37433) );
  NANDN U37711 ( .A(n38273), .B(n37433), .Z(n37354) );
  AND U37712 ( .A(n37355), .B(n37354), .Z(n37464) );
  NANDN U37713 ( .A(n37356), .B(n38369), .Z(n37358) );
  XNOR U37714 ( .A(n984), .B(a[112]), .Z(n37436) );
  NANDN U37715 ( .A(n38371), .B(n37436), .Z(n37357) );
  AND U37716 ( .A(n37358), .B(n37357), .Z(n37463) );
  XNOR U37717 ( .A(n37464), .B(n37463), .Z(n37466) );
  XNOR U37718 ( .A(n37465), .B(n37466), .Z(n37454) );
  NAND U37719 ( .A(n37941), .B(n37359), .Z(n37361) );
  XOR U37720 ( .A(n38134), .B(b[53]), .Z(n37442) );
  NANDN U37721 ( .A(n37442), .B(n37940), .Z(n37360) );
  NAND U37722 ( .A(n37361), .B(n37360), .Z(n37452) );
  NAND U37723 ( .A(n37802), .B(n37362), .Z(n37364) );
  XOR U37724 ( .A(a[122]), .B(n980), .Z(n37439) );
  NANDN U37725 ( .A(n37439), .B(n37803), .Z(n37363) );
  AND U37726 ( .A(n37364), .B(n37363), .Z(n37451) );
  XNOR U37727 ( .A(n37452), .B(n37451), .Z(n37453) );
  XNOR U37728 ( .A(n37454), .B(n37453), .Z(n37460) );
  NANDN U37729 ( .A(n37366), .B(n37365), .Z(n37370) );
  NANDN U37730 ( .A(n37368), .B(n37367), .Z(n37369) );
  NAND U37731 ( .A(n37370), .B(n37369), .Z(n37457) );
  XOR U37732 ( .A(a[124]), .B(n979), .Z(n37427) );
  OR U37733 ( .A(n37427), .B(n37756), .Z(n37373) );
  NANDN U37734 ( .A(n37371), .B(n37652), .Z(n37372) );
  NAND U37735 ( .A(n37373), .B(n37372), .Z(n37448) );
  NAND U37736 ( .A(n37374), .B(n37469), .Z(n37376) );
  XOR U37737 ( .A(a[126]), .B(n978), .Z(n37470) );
  NANDN U37738 ( .A(n37470), .B(n37471), .Z(n37375) );
  NAND U37739 ( .A(n37376), .B(n37375), .Z(n37445) );
  XOR U37740 ( .A(n983), .B(n38046), .Z(n37474) );
  NANDN U37741 ( .A(n965), .B(n37474), .Z(n37379) );
  NANDN U37742 ( .A(n37377), .B(n38194), .Z(n37378) );
  AND U37743 ( .A(n37379), .B(n37378), .Z(n37446) );
  XNOR U37744 ( .A(n37445), .B(n37446), .Z(n37447) );
  XNOR U37745 ( .A(n37448), .B(n37447), .Z(n37458) );
  XNOR U37746 ( .A(n37457), .B(n37458), .Z(n37459) );
  XOR U37747 ( .A(n37460), .B(n37459), .Z(n37418) );
  NANDN U37748 ( .A(n37381), .B(n37380), .Z(n37385) );
  NAND U37749 ( .A(n37383), .B(n37382), .Z(n37384) );
  NAND U37750 ( .A(n37385), .B(n37384), .Z(n37419) );
  XOR U37751 ( .A(n37418), .B(n37419), .Z(n37420) );
  XOR U37752 ( .A(n37421), .B(n37420), .Z(n37491) );
  XOR U37753 ( .A(n37490), .B(n37491), .Z(n37492) );
  XNOR U37754 ( .A(n37493), .B(n37492), .Z(n37495) );
  OR U37755 ( .A(n37387), .B(n37386), .Z(n37391) );
  NANDN U37756 ( .A(n37389), .B(n37388), .Z(n37390) );
  NAND U37757 ( .A(n37391), .B(n37390), .Z(n37494) );
  XNOR U37758 ( .A(n37495), .B(n37494), .Z(n37412) );
  NANDN U37759 ( .A(n37393), .B(n37392), .Z(n37397) );
  NAND U37760 ( .A(n37395), .B(n37394), .Z(n37396) );
  AND U37761 ( .A(n37397), .B(n37396), .Z(n37413) );
  XNOR U37762 ( .A(n37412), .B(n37413), .Z(n37414) );
  NANDN U37763 ( .A(n37399), .B(n37398), .Z(n37403) );
  NAND U37764 ( .A(n37401), .B(n37400), .Z(n37402) );
  NAND U37765 ( .A(n37403), .B(n37402), .Z(n37415) );
  XNOR U37766 ( .A(n37414), .B(n37415), .Z(n37407) );
  IV U37767 ( .A(n37407), .Z(n37405) );
  XOR U37768 ( .A(n37406), .B(n37405), .Z(n37404) );
  XNOR U37769 ( .A(n37409), .B(n37404), .Z(n37498) );
  XOR U37770 ( .A(n37499), .B(n37498), .Z(c[236]) );
  NANDN U37771 ( .A(n37405), .B(n37406), .Z(n37411) );
  NOR U37772 ( .A(n37407), .B(n37406), .Z(n37408) );
  OR U37773 ( .A(n37409), .B(n37408), .Z(n37410) );
  NAND U37774 ( .A(n37411), .B(n37410), .Z(n37502) );
  NANDN U37775 ( .A(n37413), .B(n37412), .Z(n37417) );
  NANDN U37776 ( .A(n37415), .B(n37414), .Z(n37416) );
  NAND U37777 ( .A(n37417), .B(n37416), .Z(n37500) );
  OR U37778 ( .A(n37419), .B(n37418), .Z(n37423) );
  NAND U37779 ( .A(n37421), .B(n37420), .Z(n37422) );
  NAND U37780 ( .A(n37423), .B(n37422), .Z(n37512) );
  XOR U37781 ( .A(b[55]), .B(n38193), .Z(n37545) );
  NANDN U37782 ( .A(n37545), .B(n38075), .Z(n37426) );
  NAND U37783 ( .A(n37424), .B(n38073), .Z(n37425) );
  NAND U37784 ( .A(n37426), .B(n37425), .Z(n37554) );
  XNOR U37785 ( .A(a[125]), .B(b[49]), .Z(n37539) );
  OR U37786 ( .A(n37539), .B(n37756), .Z(n37429) );
  NANDN U37787 ( .A(n37427), .B(n37652), .Z(n37428) );
  NAND U37788 ( .A(n37429), .B(n37428), .Z(n37551) );
  XNOR U37789 ( .A(b[63]), .B(a[111]), .Z(n37584) );
  NANDN U37790 ( .A(n37584), .B(n38422), .Z(n37432) );
  NANDN U37791 ( .A(n37430), .B(n38423), .Z(n37431) );
  AND U37792 ( .A(n37432), .B(n37431), .Z(n37552) );
  XNOR U37793 ( .A(n37551), .B(n37552), .Z(n37553) );
  XNOR U37794 ( .A(n37554), .B(n37553), .Z(n37566) );
  NAND U37795 ( .A(n37433), .B(n38326), .Z(n37435) );
  XNOR U37796 ( .A(n38400), .B(a[115]), .Z(n37530) );
  NANDN U37797 ( .A(n38273), .B(n37530), .Z(n37434) );
  NAND U37798 ( .A(n37435), .B(n37434), .Z(n37560) );
  XNOR U37799 ( .A(b[61]), .B(a[113]), .Z(n37533) );
  OR U37800 ( .A(n37533), .B(n38371), .Z(n37438) );
  NAND U37801 ( .A(n37436), .B(n38369), .Z(n37437) );
  NAND U37802 ( .A(n37438), .B(n37437), .Z(n37557) );
  XNOR U37803 ( .A(a[123]), .B(n980), .Z(n37548) );
  NAND U37804 ( .A(n37548), .B(n37803), .Z(n37441) );
  NANDN U37805 ( .A(n37439), .B(n37802), .Z(n37440) );
  AND U37806 ( .A(n37441), .B(n37440), .Z(n37558) );
  XNOR U37807 ( .A(n37557), .B(n37558), .Z(n37559) );
  XNOR U37808 ( .A(n37560), .B(n37559), .Z(n37563) );
  NANDN U37809 ( .A(n37442), .B(n37941), .Z(n37444) );
  XNOR U37810 ( .A(a[121]), .B(b[53]), .Z(n37542) );
  NANDN U37811 ( .A(n37542), .B(n37940), .Z(n37443) );
  NAND U37812 ( .A(n37444), .B(n37443), .Z(n37564) );
  XNOR U37813 ( .A(n37563), .B(n37564), .Z(n37565) );
  XOR U37814 ( .A(n37566), .B(n37565), .Z(n37525) );
  NANDN U37815 ( .A(n37446), .B(n37445), .Z(n37450) );
  NAND U37816 ( .A(n37448), .B(n37447), .Z(n37449) );
  AND U37817 ( .A(n37450), .B(n37449), .Z(n37524) );
  XOR U37818 ( .A(n37525), .B(n37524), .Z(n37526) );
  NANDN U37819 ( .A(n37452), .B(n37451), .Z(n37456) );
  NAND U37820 ( .A(n37454), .B(n37453), .Z(n37455) );
  NAND U37821 ( .A(n37456), .B(n37455), .Z(n37527) );
  XOR U37822 ( .A(n37526), .B(n37527), .Z(n37590) );
  NANDN U37823 ( .A(n37458), .B(n37457), .Z(n37462) );
  NAND U37824 ( .A(n37460), .B(n37459), .Z(n37461) );
  NAND U37825 ( .A(n37462), .B(n37461), .Z(n37588) );
  OR U37826 ( .A(n37464), .B(n37463), .Z(n37468) );
  OR U37827 ( .A(n37466), .B(n37465), .Z(n37467) );
  NAND U37828 ( .A(n37468), .B(n37467), .Z(n37518) );
  XNOR U37829 ( .A(n37570), .B(n37569), .Z(n37572) );
  NANDN U37830 ( .A(n985), .B(a[109]), .Z(n37571) );
  XNOR U37831 ( .A(n37572), .B(n37571), .Z(n37575) );
  NANDN U37832 ( .A(n37470), .B(n37469), .Z(n37473) );
  XNOR U37833 ( .A(n38463), .B(b[47]), .Z(n37580) );
  NAND U37834 ( .A(n37580), .B(n37471), .Z(n37472) );
  NAND U37835 ( .A(n37473), .B(n37472), .Z(n37576) );
  XNOR U37836 ( .A(n37575), .B(n37576), .Z(n37577) );
  NAND U37837 ( .A(n38194), .B(n37474), .Z(n37476) );
  XNOR U37838 ( .A(n983), .B(a[117]), .Z(n37536) );
  NANDN U37839 ( .A(n965), .B(n37536), .Z(n37475) );
  AND U37840 ( .A(n37476), .B(n37475), .Z(n37578) );
  XNOR U37841 ( .A(n37577), .B(n37578), .Z(n37519) );
  XOR U37842 ( .A(n37518), .B(n37519), .Z(n37520) );
  OR U37843 ( .A(n37569), .B(n37477), .Z(n37481) );
  NAND U37844 ( .A(n37479), .B(n37478), .Z(n37480) );
  AND U37845 ( .A(n37481), .B(n37480), .Z(n37521) );
  XOR U37846 ( .A(n37520), .B(n37521), .Z(n37587) );
  XNOR U37847 ( .A(n37588), .B(n37587), .Z(n37589) );
  XNOR U37848 ( .A(n37590), .B(n37589), .Z(n37513) );
  XNOR U37849 ( .A(n37512), .B(n37513), .Z(n37514) );
  NANDN U37850 ( .A(n37483), .B(n37482), .Z(n37487) );
  NAND U37851 ( .A(n37485), .B(n37484), .Z(n37486) );
  NAND U37852 ( .A(n37487), .B(n37486), .Z(n37515) );
  XOR U37853 ( .A(n37514), .B(n37515), .Z(n37506) );
  XNOR U37854 ( .A(n37506), .B(n37507), .Z(n37508) );
  NAND U37855 ( .A(n37493), .B(n37492), .Z(n37497) );
  OR U37856 ( .A(n37495), .B(n37494), .Z(n37496) );
  AND U37857 ( .A(n37497), .B(n37496), .Z(n37509) );
  XNOR U37858 ( .A(n37508), .B(n37509), .Z(n37501) );
  XNOR U37859 ( .A(n37500), .B(n37501), .Z(n37503) );
  XOR U37860 ( .A(n37502), .B(n37503), .Z(n37593) );
  OR U37861 ( .A(n37499), .B(n37498), .Z(n37594) );
  XNOR U37862 ( .A(n37593), .B(n37594), .Z(c[237]) );
  NANDN U37863 ( .A(n37501), .B(n37500), .Z(n37505) );
  NAND U37864 ( .A(n37503), .B(n37502), .Z(n37504) );
  NAND U37865 ( .A(n37505), .B(n37504), .Z(n37598) );
  NANDN U37866 ( .A(n37507), .B(n37506), .Z(n37511) );
  NAND U37867 ( .A(n37509), .B(n37508), .Z(n37510) );
  NAND U37868 ( .A(n37511), .B(n37510), .Z(n37595) );
  NANDN U37869 ( .A(n37513), .B(n37512), .Z(n37517) );
  NANDN U37870 ( .A(n37515), .B(n37514), .Z(n37516) );
  NAND U37871 ( .A(n37517), .B(n37516), .Z(n37675) );
  OR U37872 ( .A(n37519), .B(n37518), .Z(n37523) );
  NAND U37873 ( .A(n37521), .B(n37520), .Z(n37522) );
  NAND U37874 ( .A(n37523), .B(n37522), .Z(n37604) );
  OR U37875 ( .A(n37525), .B(n37524), .Z(n37529) );
  NANDN U37876 ( .A(n37527), .B(n37526), .Z(n37528) );
  NAND U37877 ( .A(n37529), .B(n37528), .Z(n37602) );
  NAND U37878 ( .A(n38326), .B(n37530), .Z(n37532) );
  XOR U37879 ( .A(n38400), .B(n38046), .Z(n37627) );
  NANDN U37880 ( .A(n38273), .B(n37627), .Z(n37531) );
  NAND U37881 ( .A(n37532), .B(n37531), .Z(n37659) );
  XOR U37882 ( .A(b[61]), .B(n37873), .Z(n37630) );
  OR U37883 ( .A(n37630), .B(n38371), .Z(n37535) );
  NANDN U37884 ( .A(n37533), .B(n38369), .Z(n37534) );
  NAND U37885 ( .A(n37535), .B(n37534), .Z(n37656) );
  XOR U37886 ( .A(b[57]), .B(n38143), .Z(n37637) );
  OR U37887 ( .A(n37637), .B(n965), .Z(n37538) );
  NAND U37888 ( .A(n37536), .B(n38194), .Z(n37537) );
  AND U37889 ( .A(n37538), .B(n37537), .Z(n37657) );
  XNOR U37890 ( .A(n37656), .B(n37657), .Z(n37658) );
  XNOR U37891 ( .A(n37659), .B(n37658), .Z(n37616) );
  XOR U37892 ( .A(a[126]), .B(n979), .Z(n37653) );
  OR U37893 ( .A(n37653), .B(n37756), .Z(n37541) );
  NANDN U37894 ( .A(n37539), .B(n37652), .Z(n37540) );
  NAND U37895 ( .A(n37541), .B(n37540), .Z(n37643) );
  XOR U37896 ( .A(a[122]), .B(n981), .Z(n37624) );
  NANDN U37897 ( .A(n37624), .B(n37940), .Z(n37544) );
  NANDN U37898 ( .A(n37542), .B(n37941), .Z(n37543) );
  NAND U37899 ( .A(n37544), .B(n37543), .Z(n37640) );
  XOR U37900 ( .A(b[55]), .B(n38134), .Z(n37646) );
  NANDN U37901 ( .A(n37646), .B(n38075), .Z(n37547) );
  NANDN U37902 ( .A(n37545), .B(n38073), .Z(n37546) );
  AND U37903 ( .A(n37547), .B(n37546), .Z(n37641) );
  XNOR U37904 ( .A(n37640), .B(n37641), .Z(n37642) );
  XNOR U37905 ( .A(n37643), .B(n37642), .Z(n37613) );
  NAND U37906 ( .A(n37802), .B(n37548), .Z(n37550) );
  XOR U37907 ( .A(a[124]), .B(n980), .Z(n37649) );
  NANDN U37908 ( .A(n37649), .B(n37803), .Z(n37549) );
  NAND U37909 ( .A(n37550), .B(n37549), .Z(n37614) );
  XNOR U37910 ( .A(n37613), .B(n37614), .Z(n37615) );
  XOR U37911 ( .A(n37616), .B(n37615), .Z(n37610) );
  NANDN U37912 ( .A(n37552), .B(n37551), .Z(n37556) );
  NAND U37913 ( .A(n37554), .B(n37553), .Z(n37555) );
  NAND U37914 ( .A(n37556), .B(n37555), .Z(n37607) );
  NANDN U37915 ( .A(n37558), .B(n37557), .Z(n37562) );
  NAND U37916 ( .A(n37560), .B(n37559), .Z(n37561) );
  AND U37917 ( .A(n37562), .B(n37561), .Z(n37608) );
  XNOR U37918 ( .A(n37607), .B(n37608), .Z(n37609) );
  XNOR U37919 ( .A(n37610), .B(n37609), .Z(n37670) );
  NANDN U37920 ( .A(n37564), .B(n37563), .Z(n37568) );
  NAND U37921 ( .A(n37566), .B(n37565), .Z(n37567) );
  NAND U37922 ( .A(n37568), .B(n37567), .Z(n37669) );
  NAND U37923 ( .A(n37570), .B(n37569), .Z(n37574) );
  OR U37924 ( .A(n37572), .B(n37571), .Z(n37573) );
  NAND U37925 ( .A(n37574), .B(n37573), .Z(n37662) );
  XNOR U37926 ( .A(n37662), .B(n37663), .Z(n37664) );
  NAND U37927 ( .A(b[45]), .B(b[46]), .Z(n37633) );
  XOR U37928 ( .A(n978), .B(n37633), .Z(n37582) );
  XNOR U37929 ( .A(b[46]), .B(b[45]), .Z(n37579) );
  NANDN U37930 ( .A(n37580), .B(n37579), .Z(n37581) );
  AND U37931 ( .A(n37582), .B(n37581), .Z(n37620) );
  AND U37932 ( .A(a[110]), .B(b[63]), .Z(n37720) );
  XOR U37933 ( .A(b[63]), .B(n37583), .Z(n37634) );
  NANDN U37934 ( .A(n37634), .B(n38422), .Z(n37586) );
  NANDN U37935 ( .A(n37584), .B(n38423), .Z(n37585) );
  AND U37936 ( .A(n37586), .B(n37585), .Z(n37619) );
  XOR U37937 ( .A(n37720), .B(n37619), .Z(n37621) );
  XOR U37938 ( .A(n37620), .B(n37621), .Z(n37665) );
  XOR U37939 ( .A(n37664), .B(n37665), .Z(n37668) );
  XOR U37940 ( .A(n37669), .B(n37668), .Z(n37671) );
  XNOR U37941 ( .A(n37670), .B(n37671), .Z(n37601) );
  XNOR U37942 ( .A(n37602), .B(n37601), .Z(n37603) );
  XNOR U37943 ( .A(n37604), .B(n37603), .Z(n37672) );
  NANDN U37944 ( .A(n37588), .B(n37587), .Z(n37592) );
  NAND U37945 ( .A(n37590), .B(n37589), .Z(n37591) );
  AND U37946 ( .A(n37592), .B(n37591), .Z(n37673) );
  XNOR U37947 ( .A(n37672), .B(n37673), .Z(n37674) );
  XOR U37948 ( .A(n37675), .B(n37674), .Z(n37596) );
  XNOR U37949 ( .A(n37595), .B(n37596), .Z(n37597) );
  XNOR U37950 ( .A(n37598), .B(n37597), .Z(n37679) );
  NANDN U37951 ( .A(n37594), .B(n37593), .Z(n37678) );
  XOR U37952 ( .A(n37679), .B(n37678), .Z(c[238]) );
  NANDN U37953 ( .A(n37596), .B(n37595), .Z(n37600) );
  NAND U37954 ( .A(n37598), .B(n37597), .Z(n37599) );
  NAND U37955 ( .A(n37600), .B(n37599), .Z(n37685) );
  NAND U37956 ( .A(n37602), .B(n37601), .Z(n37606) );
  OR U37957 ( .A(n37604), .B(n37603), .Z(n37605) );
  NAND U37958 ( .A(n37606), .B(n37605), .Z(n37765) );
  NANDN U37959 ( .A(n37608), .B(n37607), .Z(n37612) );
  NANDN U37960 ( .A(n37610), .B(n37609), .Z(n37611) );
  NAND U37961 ( .A(n37612), .B(n37611), .Z(n37688) );
  NANDN U37962 ( .A(n37614), .B(n37613), .Z(n37618) );
  NAND U37963 ( .A(n37616), .B(n37615), .Z(n37617) );
  NAND U37964 ( .A(n37618), .B(n37617), .Z(n37695) );
  OR U37965 ( .A(n37720), .B(n37619), .Z(n37623) );
  NAND U37966 ( .A(n37621), .B(n37620), .Z(n37622) );
  NAND U37967 ( .A(n37623), .B(n37622), .Z(n37702) );
  XNOR U37968 ( .A(a[123]), .B(n981), .Z(n37745) );
  NAND U37969 ( .A(n37940), .B(n37745), .Z(n37626) );
  NANDN U37970 ( .A(n37624), .B(n37941), .Z(n37625) );
  NAND U37971 ( .A(n37626), .B(n37625), .Z(n37715) );
  NAND U37972 ( .A(n38326), .B(n37627), .Z(n37629) );
  XNOR U37973 ( .A(n38400), .B(a[117]), .Z(n37751) );
  NANDN U37974 ( .A(n38273), .B(n37751), .Z(n37628) );
  NAND U37975 ( .A(n37629), .B(n37628), .Z(n37712) );
  XNOR U37976 ( .A(b[61]), .B(a[115]), .Z(n37730) );
  OR U37977 ( .A(n37730), .B(n38371), .Z(n37632) );
  NANDN U37978 ( .A(n37630), .B(n38369), .Z(n37631) );
  AND U37979 ( .A(n37632), .B(n37631), .Z(n37713) );
  XNOR U37980 ( .A(n37712), .B(n37713), .Z(n37714) );
  XNOR U37981 ( .A(n37715), .B(n37714), .Z(n37700) );
  AND U37982 ( .A(n37633), .B(b[47]), .Z(n37718) );
  NANDN U37983 ( .A(n985), .B(a[111]), .Z(n37719) );
  XOR U37984 ( .A(n37718), .B(n37719), .Z(n37721) );
  XNOR U37985 ( .A(n37720), .B(n37721), .Z(n37736) );
  XNOR U37986 ( .A(b[63]), .B(a[113]), .Z(n37759) );
  NANDN U37987 ( .A(n37759), .B(n38422), .Z(n37636) );
  NANDN U37988 ( .A(n37634), .B(n38423), .Z(n37635) );
  NAND U37989 ( .A(n37636), .B(n37635), .Z(n37733) );
  XOR U37990 ( .A(b[57]), .B(n38193), .Z(n37727) );
  OR U37991 ( .A(n37727), .B(n965), .Z(n37639) );
  NANDN U37992 ( .A(n37637), .B(n38194), .Z(n37638) );
  AND U37993 ( .A(n37639), .B(n37638), .Z(n37734) );
  XNOR U37994 ( .A(n37733), .B(n37734), .Z(n37735) );
  XNOR U37995 ( .A(n37736), .B(n37735), .Z(n37701) );
  XOR U37996 ( .A(n37700), .B(n37701), .Z(n37703) );
  XOR U37997 ( .A(n37702), .B(n37703), .Z(n37694) );
  XNOR U37998 ( .A(n37695), .B(n37694), .Z(n37697) );
  NANDN U37999 ( .A(n37641), .B(n37640), .Z(n37645) );
  NAND U38000 ( .A(n37643), .B(n37642), .Z(n37644) );
  NAND U38001 ( .A(n37645), .B(n37644), .Z(n37708) );
  XNOR U38002 ( .A(b[55]), .B(a[121]), .Z(n37724) );
  NANDN U38003 ( .A(n37724), .B(n38075), .Z(n37648) );
  NANDN U38004 ( .A(n37646), .B(n38073), .Z(n37647) );
  NAND U38005 ( .A(n37648), .B(n37647), .Z(n37742) );
  XNOR U38006 ( .A(a[125]), .B(b[51]), .Z(n37748) );
  NANDN U38007 ( .A(n37748), .B(n37803), .Z(n37651) );
  NANDN U38008 ( .A(n37649), .B(n37802), .Z(n37650) );
  NAND U38009 ( .A(n37651), .B(n37650), .Z(n37739) );
  XOR U38010 ( .A(a[127]), .B(n979), .Z(n37755) );
  OR U38011 ( .A(n37755), .B(n37756), .Z(n37655) );
  NANDN U38012 ( .A(n37653), .B(n37652), .Z(n37654) );
  AND U38013 ( .A(n37655), .B(n37654), .Z(n37740) );
  XNOR U38014 ( .A(n37739), .B(n37740), .Z(n37741) );
  XNOR U38015 ( .A(n37742), .B(n37741), .Z(n37706) );
  NANDN U38016 ( .A(n37657), .B(n37656), .Z(n37661) );
  NAND U38017 ( .A(n37659), .B(n37658), .Z(n37660) );
  NAND U38018 ( .A(n37661), .B(n37660), .Z(n37707) );
  XOR U38019 ( .A(n37706), .B(n37707), .Z(n37709) );
  XOR U38020 ( .A(n37708), .B(n37709), .Z(n37696) );
  XOR U38021 ( .A(n37697), .B(n37696), .Z(n37689) );
  XOR U38022 ( .A(n37688), .B(n37689), .Z(n37690) );
  NANDN U38023 ( .A(n37663), .B(n37662), .Z(n37667) );
  NAND U38024 ( .A(n37665), .B(n37664), .Z(n37666) );
  NAND U38025 ( .A(n37667), .B(n37666), .Z(n37691) );
  XOR U38026 ( .A(n37690), .B(n37691), .Z(n37762) );
  XNOR U38027 ( .A(n37762), .B(n37763), .Z(n37764) );
  XNOR U38028 ( .A(n37765), .B(n37764), .Z(n37683) );
  NANDN U38029 ( .A(n37673), .B(n37672), .Z(n37677) );
  NAND U38030 ( .A(n37675), .B(n37674), .Z(n37676) );
  AND U38031 ( .A(n37677), .B(n37676), .Z(n37682) );
  XNOR U38032 ( .A(n37683), .B(n37682), .Z(n37684) );
  XNOR U38033 ( .A(n37685), .B(n37684), .Z(n37681) );
  OR U38034 ( .A(n37679), .B(n37678), .Z(n37680) );
  XOR U38035 ( .A(n37681), .B(n37680), .Z(c[239]) );
  OR U38036 ( .A(n37681), .B(n37680), .Z(n37843) );
  NANDN U38037 ( .A(n37683), .B(n37682), .Z(n37687) );
  NAND U38038 ( .A(n37685), .B(n37684), .Z(n37686) );
  AND U38039 ( .A(n37687), .B(n37686), .Z(n37771) );
  OR U38040 ( .A(n37689), .B(n37688), .Z(n37693) );
  NANDN U38041 ( .A(n37691), .B(n37690), .Z(n37692) );
  NAND U38042 ( .A(n37693), .B(n37692), .Z(n37839) );
  NAND U38043 ( .A(n37695), .B(n37694), .Z(n37699) );
  NANDN U38044 ( .A(n37697), .B(n37696), .Z(n37698) );
  NAND U38045 ( .A(n37699), .B(n37698), .Z(n37836) );
  NANDN U38046 ( .A(n37701), .B(n37700), .Z(n37705) );
  OR U38047 ( .A(n37703), .B(n37702), .Z(n37704) );
  NAND U38048 ( .A(n37705), .B(n37704), .Z(n37775) );
  NANDN U38049 ( .A(n37707), .B(n37706), .Z(n37711) );
  OR U38050 ( .A(n37709), .B(n37708), .Z(n37710) );
  NAND U38051 ( .A(n37711), .B(n37710), .Z(n37772) );
  NANDN U38052 ( .A(n37713), .B(n37712), .Z(n37717) );
  NAND U38053 ( .A(n37715), .B(n37714), .Z(n37716) );
  NAND U38054 ( .A(n37717), .B(n37716), .Z(n37778) );
  OR U38055 ( .A(n37719), .B(n37718), .Z(n37723) );
  NAND U38056 ( .A(n37721), .B(n37720), .Z(n37722) );
  AND U38057 ( .A(n37723), .B(n37722), .Z(n37779) );
  XNOR U38058 ( .A(n37778), .B(n37779), .Z(n37780) );
  XNOR U38059 ( .A(n38251), .B(b[55]), .Z(n37815) );
  NAND U38060 ( .A(n38075), .B(n37815), .Z(n37726) );
  NANDN U38061 ( .A(n37724), .B(n38073), .Z(n37725) );
  NAND U38062 ( .A(n37726), .B(n37725), .Z(n37812) );
  XOR U38063 ( .A(b[57]), .B(n38134), .Z(n37824) );
  OR U38064 ( .A(n37824), .B(n965), .Z(n37729) );
  NANDN U38065 ( .A(n37727), .B(n38194), .Z(n37728) );
  NAND U38066 ( .A(n37729), .B(n37728), .Z(n37809) );
  XNOR U38067 ( .A(n984), .B(a[116]), .Z(n37827) );
  NANDN U38068 ( .A(n38371), .B(n37827), .Z(n37732) );
  NANDN U38069 ( .A(n37730), .B(n38369), .Z(n37731) );
  AND U38070 ( .A(n37732), .B(n37731), .Z(n37810) );
  XNOR U38071 ( .A(n37809), .B(n37810), .Z(n37811) );
  XNOR U38072 ( .A(n37812), .B(n37811), .Z(n37781) );
  XOR U38073 ( .A(n37780), .B(n37781), .Z(n37833) );
  NANDN U38074 ( .A(n37734), .B(n37733), .Z(n37738) );
  NANDN U38075 ( .A(n37736), .B(n37735), .Z(n37737) );
  NAND U38076 ( .A(n37738), .B(n37737), .Z(n37831) );
  NANDN U38077 ( .A(n37740), .B(n37739), .Z(n37744) );
  NAND U38078 ( .A(n37742), .B(n37741), .Z(n37743) );
  NAND U38079 ( .A(n37744), .B(n37743), .Z(n37797) );
  XOR U38080 ( .A(a[124]), .B(n981), .Z(n37818) );
  NANDN U38081 ( .A(n37818), .B(n37940), .Z(n37747) );
  NAND U38082 ( .A(n37745), .B(n37941), .Z(n37746) );
  NAND U38083 ( .A(n37747), .B(n37746), .Z(n37787) );
  XOR U38084 ( .A(n987), .B(n980), .Z(n37801) );
  NAND U38085 ( .A(n37801), .B(n37803), .Z(n37750) );
  NANDN U38086 ( .A(n37748), .B(n37802), .Z(n37749) );
  NAND U38087 ( .A(n37750), .B(n37749), .Z(n37784) );
  NAND U38088 ( .A(n37751), .B(n38326), .Z(n37753) );
  XOR U38089 ( .A(b[59]), .B(n38143), .Z(n37806) );
  OR U38090 ( .A(n37806), .B(n38273), .Z(n37752) );
  AND U38091 ( .A(n37753), .B(n37752), .Z(n37785) );
  XNOR U38092 ( .A(n37784), .B(n37785), .Z(n37786) );
  XNOR U38093 ( .A(n37787), .B(n37786), .Z(n37795) );
  XOR U38094 ( .A(n979), .B(n37754), .Z(n37758) );
  NAND U38095 ( .A(n37756), .B(n37755), .Z(n37757) );
  AND U38096 ( .A(n37758), .B(n37757), .Z(n37791) );
  AND U38097 ( .A(b[63]), .B(a[112]), .Z(n37864) );
  XOR U38098 ( .A(b[63]), .B(n37873), .Z(n37821) );
  NANDN U38099 ( .A(n37821), .B(n38422), .Z(n37761) );
  NANDN U38100 ( .A(n37759), .B(n38423), .Z(n37760) );
  AND U38101 ( .A(n37761), .B(n37760), .Z(n37790) );
  XNOR U38102 ( .A(n37864), .B(n37790), .Z(n37792) );
  XNOR U38103 ( .A(n37791), .B(n37792), .Z(n37796) );
  XOR U38104 ( .A(n37795), .B(n37796), .Z(n37798) );
  XOR U38105 ( .A(n37797), .B(n37798), .Z(n37830) );
  XNOR U38106 ( .A(n37831), .B(n37830), .Z(n37832) );
  XNOR U38107 ( .A(n37833), .B(n37832), .Z(n37773) );
  XNOR U38108 ( .A(n37772), .B(n37773), .Z(n37774) );
  XNOR U38109 ( .A(n37775), .B(n37774), .Z(n37837) );
  XNOR U38110 ( .A(n37836), .B(n37837), .Z(n37838) );
  XNOR U38111 ( .A(n37839), .B(n37838), .Z(n37769) );
  NANDN U38112 ( .A(n37763), .B(n37762), .Z(n37767) );
  NAND U38113 ( .A(n37765), .B(n37764), .Z(n37766) );
  AND U38114 ( .A(n37767), .B(n37766), .Z(n37770) );
  XOR U38115 ( .A(n37769), .B(n37770), .Z(n37768) );
  XNOR U38116 ( .A(n37771), .B(n37768), .Z(n37842) );
  XOR U38117 ( .A(n37843), .B(n37842), .Z(c[240]) );
  NANDN U38118 ( .A(n37773), .B(n37772), .Z(n37777) );
  NAND U38119 ( .A(n37775), .B(n37774), .Z(n37776) );
  NAND U38120 ( .A(n37777), .B(n37776), .Z(n37917) );
  NANDN U38121 ( .A(n37779), .B(n37778), .Z(n37783) );
  NANDN U38122 ( .A(n37781), .B(n37780), .Z(n37782) );
  AND U38123 ( .A(n37783), .B(n37782), .Z(n37853) );
  NANDN U38124 ( .A(n37785), .B(n37784), .Z(n37789) );
  NAND U38125 ( .A(n37787), .B(n37786), .Z(n37788) );
  AND U38126 ( .A(n37789), .B(n37788), .Z(n37850) );
  OR U38127 ( .A(n37790), .B(n37864), .Z(n37794) );
  NANDN U38128 ( .A(n37792), .B(n37791), .Z(n37793) );
  AND U38129 ( .A(n37794), .B(n37793), .Z(n37851) );
  XNOR U38130 ( .A(n37850), .B(n37851), .Z(n37852) );
  NANDN U38131 ( .A(n37796), .B(n37795), .Z(n37800) );
  OR U38132 ( .A(n37798), .B(n37797), .Z(n37799) );
  NAND U38133 ( .A(n37800), .B(n37799), .Z(n37856) );
  XNOR U38134 ( .A(n37857), .B(n37856), .Z(n37859) );
  NANDN U38135 ( .A(n985), .B(a[113]), .Z(n37863) );
  XNOR U38136 ( .A(n37862), .B(n37863), .Z(n37865) );
  XNOR U38137 ( .A(n37864), .B(n37865), .Z(n37878) );
  NAND U38138 ( .A(n37802), .B(n37801), .Z(n37805) );
  XOR U38139 ( .A(a[127]), .B(n980), .Z(n37869) );
  NANDN U38140 ( .A(n37869), .B(n37803), .Z(n37804) );
  NAND U38141 ( .A(n37805), .B(n37804), .Z(n37877) );
  XOR U38142 ( .A(n37878), .B(n37877), .Z(n37879) );
  NANDN U38143 ( .A(n37806), .B(n38326), .Z(n37808) );
  XNOR U38144 ( .A(n38400), .B(a[119]), .Z(n37895) );
  NANDN U38145 ( .A(n38273), .B(n37895), .Z(n37807) );
  NAND U38146 ( .A(n37808), .B(n37807), .Z(n37880) );
  XOR U38147 ( .A(n37879), .B(n37880), .Z(n37904) );
  NANDN U38148 ( .A(n37810), .B(n37809), .Z(n37814) );
  NAND U38149 ( .A(n37812), .B(n37811), .Z(n37813) );
  AND U38150 ( .A(n37814), .B(n37813), .Z(n37905) );
  XNOR U38151 ( .A(n37904), .B(n37905), .Z(n37906) );
  XNOR U38152 ( .A(a[123]), .B(n982), .Z(n37901) );
  NAND U38153 ( .A(n38075), .B(n37901), .Z(n37817) );
  NAND U38154 ( .A(n37815), .B(n38073), .Z(n37816) );
  NAND U38155 ( .A(n37817), .B(n37816), .Z(n37910) );
  XNOR U38156 ( .A(a[125]), .B(b[53]), .Z(n37898) );
  NANDN U38157 ( .A(n37898), .B(n37940), .Z(n37820) );
  NANDN U38158 ( .A(n37818), .B(n37941), .Z(n37819) );
  NAND U38159 ( .A(n37820), .B(n37819), .Z(n37886) );
  XNOR U38160 ( .A(b[63]), .B(a[115]), .Z(n37874) );
  NANDN U38161 ( .A(n37874), .B(n38422), .Z(n37823) );
  NANDN U38162 ( .A(n37821), .B(n38423), .Z(n37822) );
  NAND U38163 ( .A(n37823), .B(n37822), .Z(n37883) );
  XNOR U38164 ( .A(b[57]), .B(a[121]), .Z(n37889) );
  OR U38165 ( .A(n37889), .B(n965), .Z(n37826) );
  NANDN U38166 ( .A(n37824), .B(n38194), .Z(n37825) );
  AND U38167 ( .A(n37826), .B(n37825), .Z(n37884) );
  XNOR U38168 ( .A(n37883), .B(n37884), .Z(n37885) );
  XNOR U38169 ( .A(n37886), .B(n37885), .Z(n37911) );
  XNOR U38170 ( .A(n37910), .B(n37911), .Z(n37913) );
  NAND U38171 ( .A(n37827), .B(n38369), .Z(n37829) );
  XNOR U38172 ( .A(n984), .B(a[117]), .Z(n37892) );
  NANDN U38173 ( .A(n38371), .B(n37892), .Z(n37828) );
  NAND U38174 ( .A(n37829), .B(n37828), .Z(n37912) );
  XNOR U38175 ( .A(n37913), .B(n37912), .Z(n37907) );
  XNOR U38176 ( .A(n37906), .B(n37907), .Z(n37858) );
  XNOR U38177 ( .A(n37859), .B(n37858), .Z(n37915) );
  NANDN U38178 ( .A(n37831), .B(n37830), .Z(n37835) );
  NAND U38179 ( .A(n37833), .B(n37832), .Z(n37834) );
  AND U38180 ( .A(n37835), .B(n37834), .Z(n37914) );
  XOR U38181 ( .A(n37915), .B(n37914), .Z(n37916) );
  XNOR U38182 ( .A(n37917), .B(n37916), .Z(n37844) );
  NANDN U38183 ( .A(n37837), .B(n37836), .Z(n37841) );
  NAND U38184 ( .A(n37839), .B(n37838), .Z(n37840) );
  NAND U38185 ( .A(n37841), .B(n37840), .Z(n37845) );
  XOR U38186 ( .A(n37844), .B(n37845), .Z(n37847) );
  XNOR U38187 ( .A(n37846), .B(n37847), .Z(n37920) );
  OR U38188 ( .A(n37843), .B(n37842), .Z(n37921) );
  XNOR U38189 ( .A(n37920), .B(n37921), .Z(c[241]) );
  NANDN U38190 ( .A(n37845), .B(n37844), .Z(n37849) );
  NANDN U38191 ( .A(n37847), .B(n37846), .Z(n37848) );
  NAND U38192 ( .A(n37849), .B(n37848), .Z(n37986) );
  OR U38193 ( .A(n37851), .B(n37850), .Z(n37855) );
  OR U38194 ( .A(n37853), .B(n37852), .Z(n37854) );
  NAND U38195 ( .A(n37855), .B(n37854), .Z(n37923) );
  OR U38196 ( .A(n37857), .B(n37856), .Z(n37861) );
  NANDN U38197 ( .A(n37859), .B(n37858), .Z(n37860) );
  NAND U38198 ( .A(n37861), .B(n37860), .Z(n37922) );
  XOR U38199 ( .A(n37923), .B(n37922), .Z(n37924) );
  OR U38200 ( .A(n37863), .B(n37862), .Z(n37867) );
  NANDN U38201 ( .A(n37865), .B(n37864), .Z(n37866) );
  NAND U38202 ( .A(n37867), .B(n37866), .Z(n37972) );
  XOR U38203 ( .A(n980), .B(n37868), .Z(n37872) );
  XOR U38204 ( .A(b[50]), .B(n979), .Z(n37870) );
  NAND U38205 ( .A(n37870), .B(n37869), .Z(n37871) );
  AND U38206 ( .A(n37872), .B(n37871), .Z(n37961) );
  ANDN U38207 ( .B(b[63]), .A(n37873), .Z(n38023) );
  XOR U38208 ( .A(b[63]), .B(n38046), .Z(n37951) );
  NANDN U38209 ( .A(n37951), .B(n38422), .Z(n37876) );
  NANDN U38210 ( .A(n37874), .B(n38423), .Z(n37875) );
  AND U38211 ( .A(n37876), .B(n37875), .Z(n37960) );
  XNOR U38212 ( .A(n38023), .B(n37960), .Z(n37962) );
  XNOR U38213 ( .A(n37961), .B(n37962), .Z(n37971) );
  XNOR U38214 ( .A(n37972), .B(n37971), .Z(n37974) );
  OR U38215 ( .A(n37878), .B(n37877), .Z(n37882) );
  NANDN U38216 ( .A(n37880), .B(n37879), .Z(n37881) );
  AND U38217 ( .A(n37882), .B(n37881), .Z(n37973) );
  XNOR U38218 ( .A(n37974), .B(n37973), .Z(n37936) );
  NANDN U38219 ( .A(n37884), .B(n37883), .Z(n37888) );
  NAND U38220 ( .A(n37886), .B(n37885), .Z(n37887) );
  NAND U38221 ( .A(n37888), .B(n37887), .Z(n37935) );
  XOR U38222 ( .A(b[57]), .B(n38251), .Z(n37954) );
  OR U38223 ( .A(n37954), .B(n965), .Z(n37891) );
  NANDN U38224 ( .A(n37889), .B(n38194), .Z(n37890) );
  NAND U38225 ( .A(n37891), .B(n37890), .Z(n37968) );
  XOR U38226 ( .A(b[61]), .B(n38143), .Z(n37948) );
  OR U38227 ( .A(n37948), .B(n38371), .Z(n37894) );
  NAND U38228 ( .A(n37892), .B(n38369), .Z(n37893) );
  NAND U38229 ( .A(n37894), .B(n37893), .Z(n37965) );
  NAND U38230 ( .A(n37895), .B(n38326), .Z(n37897) );
  XOR U38231 ( .A(n38400), .B(n38134), .Z(n37945) );
  NANDN U38232 ( .A(n38273), .B(n37945), .Z(n37896) );
  AND U38233 ( .A(n37897), .B(n37896), .Z(n37966) );
  XNOR U38234 ( .A(n37965), .B(n37966), .Z(n37967) );
  XNOR U38235 ( .A(n37968), .B(n37967), .Z(n37980) );
  XOR U38236 ( .A(a[126]), .B(n981), .Z(n37942) );
  NANDN U38237 ( .A(n37942), .B(n37940), .Z(n37900) );
  NANDN U38238 ( .A(n37898), .B(n37941), .Z(n37899) );
  NAND U38239 ( .A(n37900), .B(n37899), .Z(n37977) );
  XOR U38240 ( .A(a[124]), .B(n982), .Z(n37957) );
  NANDN U38241 ( .A(n37957), .B(n38075), .Z(n37903) );
  NAND U38242 ( .A(n37901), .B(n38073), .Z(n37902) );
  AND U38243 ( .A(n37903), .B(n37902), .Z(n37978) );
  XNOR U38244 ( .A(n37977), .B(n37978), .Z(n37979) );
  XNOR U38245 ( .A(n37980), .B(n37979), .Z(n37934) );
  XNOR U38246 ( .A(n37935), .B(n37934), .Z(n37937) );
  XOR U38247 ( .A(n37936), .B(n37937), .Z(n37931) );
  NANDN U38248 ( .A(n37905), .B(n37904), .Z(n37909) );
  NANDN U38249 ( .A(n37907), .B(n37906), .Z(n37908) );
  NAND U38250 ( .A(n37909), .B(n37908), .Z(n37929) );
  XNOR U38251 ( .A(n37929), .B(n37928), .Z(n37930) );
  XNOR U38252 ( .A(n37931), .B(n37930), .Z(n37925) );
  XNOR U38253 ( .A(n37924), .B(n37925), .Z(n37983) );
  OR U38254 ( .A(n37915), .B(n37914), .Z(n37919) );
  NAND U38255 ( .A(n37917), .B(n37916), .Z(n37918) );
  NAND U38256 ( .A(n37919), .B(n37918), .Z(n37984) );
  XOR U38257 ( .A(n37983), .B(n37984), .Z(n37985) );
  XNOR U38258 ( .A(n37986), .B(n37985), .Z(n37991) );
  NANDN U38259 ( .A(n37921), .B(n37920), .Z(n37990) );
  XOR U38260 ( .A(n37991), .B(n37990), .Z(c[242]) );
  OR U38261 ( .A(n37923), .B(n37922), .Z(n37927) );
  NANDN U38262 ( .A(n37925), .B(n37924), .Z(n37926) );
  NAND U38263 ( .A(n37927), .B(n37926), .Z(n37994) );
  NANDN U38264 ( .A(n37929), .B(n37928), .Z(n37933) );
  NAND U38265 ( .A(n37931), .B(n37930), .Z(n37932) );
  NAND U38266 ( .A(n37933), .B(n37932), .Z(n38053) );
  NAND U38267 ( .A(n37935), .B(n37934), .Z(n37939) );
  NANDN U38268 ( .A(n37937), .B(n37936), .Z(n37938) );
  NAND U38269 ( .A(n37939), .B(n37938), .Z(n38051) );
  XNOR U38270 ( .A(n38463), .B(b[53]), .Z(n38043) );
  NAND U38271 ( .A(n38043), .B(n37940), .Z(n37944) );
  NANDN U38272 ( .A(n37942), .B(n37941), .Z(n37943) );
  NAND U38273 ( .A(n37944), .B(n37943), .Z(n38017) );
  NAND U38274 ( .A(n38326), .B(n37945), .Z(n37947) );
  XNOR U38275 ( .A(b[59]), .B(a[121]), .Z(n38029) );
  OR U38276 ( .A(n38029), .B(n38273), .Z(n37946) );
  AND U38277 ( .A(n37947), .B(n37946), .Z(n38018) );
  XNOR U38278 ( .A(n38017), .B(n38018), .Z(n38019) );
  NANDN U38279 ( .A(n985), .B(a[115]), .Z(n38026) );
  XOR U38280 ( .A(n38023), .B(n38024), .Z(n38025) );
  XOR U38281 ( .A(n38026), .B(n38025), .Z(n38020) );
  XOR U38282 ( .A(n38019), .B(n38020), .Z(n38007) );
  XOR U38283 ( .A(b[61]), .B(n38193), .Z(n38047) );
  OR U38284 ( .A(n38047), .B(n38371), .Z(n37950) );
  NANDN U38285 ( .A(n37948), .B(n38369), .Z(n37949) );
  NAND U38286 ( .A(n37950), .B(n37949), .Z(n38005) );
  XNOR U38287 ( .A(b[63]), .B(a[117]), .Z(n38038) );
  NANDN U38288 ( .A(n38038), .B(n38422), .Z(n37953) );
  NANDN U38289 ( .A(n37951), .B(n38423), .Z(n37952) );
  NAND U38290 ( .A(n37953), .B(n37952), .Z(n38014) );
  XNOR U38291 ( .A(n983), .B(a[123]), .Z(n38032) );
  NANDN U38292 ( .A(n965), .B(n38032), .Z(n37956) );
  NANDN U38293 ( .A(n37954), .B(n38194), .Z(n37955) );
  NAND U38294 ( .A(n37956), .B(n37955), .Z(n38011) );
  XNOR U38295 ( .A(a[125]), .B(b[55]), .Z(n38035) );
  NANDN U38296 ( .A(n38035), .B(n38075), .Z(n37959) );
  NANDN U38297 ( .A(n37957), .B(n38073), .Z(n37958) );
  AND U38298 ( .A(n37959), .B(n37958), .Z(n38012) );
  XNOR U38299 ( .A(n38011), .B(n38012), .Z(n38013) );
  XNOR U38300 ( .A(n38014), .B(n38013), .Z(n38006) );
  XNOR U38301 ( .A(n38005), .B(n38006), .Z(n38008) );
  XOR U38302 ( .A(n38007), .B(n38008), .Z(n38001) );
  OR U38303 ( .A(n37960), .B(n38023), .Z(n37964) );
  NANDN U38304 ( .A(n37962), .B(n37961), .Z(n37963) );
  NAND U38305 ( .A(n37964), .B(n37963), .Z(n37999) );
  NANDN U38306 ( .A(n37966), .B(n37965), .Z(n37970) );
  NAND U38307 ( .A(n37968), .B(n37967), .Z(n37969) );
  AND U38308 ( .A(n37970), .B(n37969), .Z(n38000) );
  XNOR U38309 ( .A(n37999), .B(n38000), .Z(n38002) );
  XNOR U38310 ( .A(n38001), .B(n38002), .Z(n37995) );
  NAND U38311 ( .A(n37972), .B(n37971), .Z(n37976) );
  NANDN U38312 ( .A(n37974), .B(n37973), .Z(n37975) );
  NAND U38313 ( .A(n37976), .B(n37975), .Z(n37996) );
  XNOR U38314 ( .A(n37995), .B(n37996), .Z(n37997) );
  NANDN U38315 ( .A(n37978), .B(n37977), .Z(n37982) );
  NANDN U38316 ( .A(n37980), .B(n37979), .Z(n37981) );
  AND U38317 ( .A(n37982), .B(n37981), .Z(n37998) );
  XOR U38318 ( .A(n37997), .B(n37998), .Z(n38050) );
  XNOR U38319 ( .A(n38051), .B(n38050), .Z(n38052) );
  XNOR U38320 ( .A(n38053), .B(n38052), .Z(n37992) );
  OR U38321 ( .A(n37984), .B(n37983), .Z(n37988) );
  NAND U38322 ( .A(n37986), .B(n37985), .Z(n37987) );
  AND U38323 ( .A(n37988), .B(n37987), .Z(n37993) );
  XOR U38324 ( .A(n37992), .B(n37993), .Z(n37989) );
  XNOR U38325 ( .A(n37994), .B(n37989), .Z(n38055) );
  OR U38326 ( .A(n37991), .B(n37990), .Z(n38054) );
  XOR U38327 ( .A(n38055), .B(n38054), .Z(c[243]) );
  NANDN U38328 ( .A(n38000), .B(n37999), .Z(n38004) );
  NAND U38329 ( .A(n38002), .B(n38001), .Z(n38003) );
  NAND U38330 ( .A(n38004), .B(n38003), .Z(n38110) );
  NANDN U38331 ( .A(n38006), .B(n38005), .Z(n38010) );
  NAND U38332 ( .A(n38008), .B(n38007), .Z(n38009) );
  NAND U38333 ( .A(n38010), .B(n38009), .Z(n38103) );
  NANDN U38334 ( .A(n38012), .B(n38011), .Z(n38016) );
  NAND U38335 ( .A(n38014), .B(n38013), .Z(n38015) );
  NAND U38336 ( .A(n38016), .B(n38015), .Z(n38100) );
  NANDN U38337 ( .A(n38018), .B(n38017), .Z(n38022) );
  NAND U38338 ( .A(n38020), .B(n38019), .Z(n38021) );
  NAND U38339 ( .A(n38022), .B(n38021), .Z(n38098) );
  NANDN U38340 ( .A(n38024), .B(n38023), .Z(n38028) );
  OR U38341 ( .A(n38026), .B(n38025), .Z(n38027) );
  AND U38342 ( .A(n38028), .B(n38027), .Z(n38097) );
  XNOR U38343 ( .A(n38098), .B(n38097), .Z(n38099) );
  XOR U38344 ( .A(n38100), .B(n38099), .Z(n38104) );
  XOR U38345 ( .A(n38103), .B(n38104), .Z(n38105) );
  NANDN U38346 ( .A(n38029), .B(n38326), .Z(n38031) );
  XOR U38347 ( .A(n38400), .B(n38251), .Z(n38078) );
  NANDN U38348 ( .A(n38273), .B(n38078), .Z(n38030) );
  NAND U38349 ( .A(n38031), .B(n38030), .Z(n38072) );
  NAND U38350 ( .A(n38194), .B(n38032), .Z(n38034) );
  XOR U38351 ( .A(n38321), .B(n983), .Z(n38085) );
  NANDN U38352 ( .A(n965), .B(n38085), .Z(n38033) );
  NAND U38353 ( .A(n38034), .B(n38033), .Z(n38069) );
  XNOR U38354 ( .A(n987), .B(b[55]), .Z(n38074) );
  NAND U38355 ( .A(n38075), .B(n38074), .Z(n38037) );
  NANDN U38356 ( .A(n38035), .B(n38073), .Z(n38036) );
  AND U38357 ( .A(n38037), .B(n38036), .Z(n38070) );
  XNOR U38358 ( .A(n38069), .B(n38070), .Z(n38071) );
  XOR U38359 ( .A(n38072), .B(n38071), .Z(n38094) );
  XOR U38360 ( .A(b[63]), .B(n38143), .Z(n38082) );
  NANDN U38361 ( .A(n38082), .B(n38422), .Z(n38040) );
  NANDN U38362 ( .A(n38038), .B(n38423), .Z(n38039) );
  NAND U38363 ( .A(n38040), .B(n38039), .Z(n38065) );
  XOR U38364 ( .A(n981), .B(n38041), .Z(n38045) );
  XOR U38365 ( .A(b[52]), .B(n980), .Z(n38042) );
  NANDN U38366 ( .A(n38043), .B(n38042), .Z(n38044) );
  AND U38367 ( .A(n38045), .B(n38044), .Z(n38064) );
  ANDN U38368 ( .B(b[63]), .A(n38046), .Z(n38119) );
  XOR U38369 ( .A(n38064), .B(n38119), .Z(n38066) );
  XOR U38370 ( .A(n38065), .B(n38066), .Z(n38091) );
  NANDN U38371 ( .A(n38047), .B(n38369), .Z(n38049) );
  XOR U38372 ( .A(b[61]), .B(n38134), .Z(n38088) );
  OR U38373 ( .A(n38088), .B(n38371), .Z(n38048) );
  NAND U38374 ( .A(n38049), .B(n38048), .Z(n38092) );
  XNOR U38375 ( .A(n38091), .B(n38092), .Z(n38093) );
  XOR U38376 ( .A(n38094), .B(n38093), .Z(n38106) );
  XNOR U38377 ( .A(n38105), .B(n38106), .Z(n38109) );
  XNOR U38378 ( .A(n38110), .B(n38109), .Z(n38111) );
  XNOR U38379 ( .A(n38112), .B(n38111), .Z(n38058) );
  XOR U38380 ( .A(n38058), .B(n38059), .Z(n38061) );
  XNOR U38381 ( .A(n38060), .B(n38061), .Z(n38056) );
  OR U38382 ( .A(n38055), .B(n38054), .Z(n38057) );
  XNOR U38383 ( .A(n38056), .B(n38057), .Z(c[244]) );
  NANDN U38384 ( .A(n38057), .B(n38056), .Z(n38167) );
  NANDN U38385 ( .A(n38059), .B(n38058), .Z(n38063) );
  NANDN U38386 ( .A(n38061), .B(n38060), .Z(n38062) );
  NAND U38387 ( .A(n38063), .B(n38062), .Z(n38116) );
  NANDN U38388 ( .A(n38119), .B(n38064), .Z(n38068) );
  NANDN U38389 ( .A(n38066), .B(n38065), .Z(n38067) );
  NAND U38390 ( .A(n38068), .B(n38067), .Z(n38148) );
  NAND U38391 ( .A(n38074), .B(n38073), .Z(n38077) );
  XOR U38392 ( .A(a[127]), .B(n982), .Z(n38139) );
  NANDN U38393 ( .A(n38139), .B(n38075), .Z(n38076) );
  NAND U38394 ( .A(n38077), .B(n38076), .Z(n38144) );
  NAND U38395 ( .A(n38078), .B(n38326), .Z(n38080) );
  XNOR U38396 ( .A(n38400), .B(a[123]), .Z(n38128) );
  NANDN U38397 ( .A(n38273), .B(n38128), .Z(n38079) );
  AND U38398 ( .A(n38080), .B(n38079), .Z(n38145) );
  XNOR U38399 ( .A(n38144), .B(n38145), .Z(n38147) );
  NANDN U38400 ( .A(n985), .B(a[117]), .Z(n38118) );
  XOR U38401 ( .A(n38081), .B(n38118), .Z(n38120) );
  XNOR U38402 ( .A(n38119), .B(n38120), .Z(n38146) );
  XNOR U38403 ( .A(n38147), .B(n38146), .Z(n38155) );
  XNOR U38404 ( .A(n985), .B(a[119]), .Z(n38135) );
  NAND U38405 ( .A(n38135), .B(n38422), .Z(n38084) );
  NANDN U38406 ( .A(n38082), .B(n38423), .Z(n38083) );
  NAND U38407 ( .A(n38084), .B(n38083), .Z(n38123) );
  NAND U38408 ( .A(n38194), .B(n38085), .Z(n38087) );
  XNOR U38409 ( .A(a[125]), .B(n983), .Z(n38131) );
  NANDN U38410 ( .A(n965), .B(n38131), .Z(n38086) );
  NAND U38411 ( .A(n38087), .B(n38086), .Z(n38121) );
  NANDN U38412 ( .A(n38088), .B(n38369), .Z(n38090) );
  XNOR U38413 ( .A(n984), .B(a[121]), .Z(n38125) );
  NANDN U38414 ( .A(n38371), .B(n38125), .Z(n38089) );
  NAND U38415 ( .A(n38090), .B(n38089), .Z(n38122) );
  XNOR U38416 ( .A(n38121), .B(n38122), .Z(n38124) );
  XOR U38417 ( .A(n38123), .B(n38124), .Z(n38154) );
  XNOR U38418 ( .A(n38155), .B(n38154), .Z(n38156) );
  XNOR U38419 ( .A(n38148), .B(n38149), .Z(n38150) );
  NANDN U38420 ( .A(n38092), .B(n38091), .Z(n38096) );
  NANDN U38421 ( .A(n38094), .B(n38093), .Z(n38095) );
  NAND U38422 ( .A(n38096), .B(n38095), .Z(n38151) );
  XOR U38423 ( .A(n38150), .B(n38151), .Z(n38163) );
  NANDN U38424 ( .A(n38098), .B(n38097), .Z(n38102) );
  NANDN U38425 ( .A(n38100), .B(n38099), .Z(n38101) );
  NAND U38426 ( .A(n38102), .B(n38101), .Z(n38160) );
  OR U38427 ( .A(n38104), .B(n38103), .Z(n38108) );
  NANDN U38428 ( .A(n38106), .B(n38105), .Z(n38107) );
  AND U38429 ( .A(n38108), .B(n38107), .Z(n38161) );
  XNOR U38430 ( .A(n38160), .B(n38161), .Z(n38162) );
  XNOR U38431 ( .A(n38163), .B(n38162), .Z(n38114) );
  XOR U38432 ( .A(n38114), .B(n38115), .Z(n38113) );
  XOR U38433 ( .A(n38116), .B(n38113), .Z(n38166) );
  XNOR U38434 ( .A(n38167), .B(n38166), .Z(c[245]) );
  XOR U38435 ( .A(b[61]), .B(n38251), .Z(n38198) );
  OR U38436 ( .A(n38198), .B(n38371), .Z(n38127) );
  NAND U38437 ( .A(n38125), .B(n38369), .Z(n38126) );
  NAND U38438 ( .A(n38127), .B(n38126), .Z(n38209) );
  NAND U38439 ( .A(n38326), .B(n38128), .Z(n38130) );
  XOR U38440 ( .A(n38400), .B(n38321), .Z(n38189) );
  NANDN U38441 ( .A(n38273), .B(n38189), .Z(n38129) );
  NAND U38442 ( .A(n38130), .B(n38129), .Z(n38206) );
  XOR U38443 ( .A(a[126]), .B(n983), .Z(n38195) );
  OR U38444 ( .A(n38195), .B(n965), .Z(n38133) );
  NAND U38445 ( .A(n38131), .B(n38194), .Z(n38132) );
  AND U38446 ( .A(n38133), .B(n38132), .Z(n38207) );
  XNOR U38447 ( .A(n38206), .B(n38207), .Z(n38208) );
  XOR U38448 ( .A(n38209), .B(n38208), .Z(n38176) );
  XOR U38449 ( .A(b[63]), .B(n38134), .Z(n38186) );
  NANDN U38450 ( .A(n38186), .B(n38422), .Z(n38137) );
  NAND U38451 ( .A(n38135), .B(n38423), .Z(n38136) );
  NAND U38452 ( .A(n38137), .B(n38136), .Z(n38202) );
  XOR U38453 ( .A(n982), .B(n38138), .Z(n38142) );
  XOR U38454 ( .A(b[54]), .B(n981), .Z(n38140) );
  NAND U38455 ( .A(n38140), .B(n38139), .Z(n38141) );
  AND U38456 ( .A(n38142), .B(n38141), .Z(n38201) );
  ANDN U38457 ( .B(b[63]), .A(n38143), .Z(n38235) );
  XOR U38458 ( .A(n38201), .B(n38235), .Z(n38203) );
  XNOR U38459 ( .A(n38202), .B(n38203), .Z(n38177) );
  XOR U38460 ( .A(n38176), .B(n38177), .Z(n38178) );
  XNOR U38461 ( .A(n38179), .B(n38178), .Z(n38182) );
  XNOR U38462 ( .A(n38182), .B(n38183), .Z(n38185) );
  XOR U38463 ( .A(n38184), .B(n38185), .Z(n38212) );
  NANDN U38464 ( .A(n38149), .B(n38148), .Z(n38153) );
  NANDN U38465 ( .A(n38151), .B(n38150), .Z(n38152) );
  NAND U38466 ( .A(n38153), .B(n38152), .Z(n38213) );
  XNOR U38467 ( .A(n38212), .B(n38213), .Z(n38214) );
  OR U38468 ( .A(n38155), .B(n38154), .Z(n38159) );
  OR U38469 ( .A(n38157), .B(n38156), .Z(n38158) );
  NAND U38470 ( .A(n38159), .B(n38158), .Z(n38215) );
  XOR U38471 ( .A(n38214), .B(n38215), .Z(n38170) );
  NANDN U38472 ( .A(n38161), .B(n38160), .Z(n38165) );
  NAND U38473 ( .A(n38163), .B(n38162), .Z(n38164) );
  NAND U38474 ( .A(n38165), .B(n38164), .Z(n38171) );
  XNOR U38475 ( .A(n38170), .B(n38171), .Z(n38173) );
  XOR U38476 ( .A(n38172), .B(n38173), .Z(n38168) );
  NANDN U38477 ( .A(n38167), .B(n38166), .Z(n38169) );
  XNOR U38478 ( .A(n38168), .B(n38169), .Z(c[246]) );
  NANDN U38479 ( .A(n38169), .B(n38168), .Z(n38266) );
  NANDN U38480 ( .A(n38171), .B(n38170), .Z(n38175) );
  NAND U38481 ( .A(n38173), .B(n38172), .Z(n38174) );
  NAND U38482 ( .A(n38175), .B(n38174), .Z(n38263) );
  OR U38483 ( .A(n38177), .B(n38176), .Z(n38181) );
  NANDN U38484 ( .A(n38179), .B(n38178), .Z(n38180) );
  AND U38485 ( .A(n38181), .B(n38180), .Z(n38217) );
  XOR U38486 ( .A(n38217), .B(n38218), .Z(n38219) );
  XNOR U38487 ( .A(b[63]), .B(a[121]), .Z(n38252) );
  NANDN U38488 ( .A(n38252), .B(n38422), .Z(n38188) );
  NANDN U38489 ( .A(n38186), .B(n38423), .Z(n38187) );
  NAND U38490 ( .A(n38188), .B(n38187), .Z(n38258) );
  NAND U38491 ( .A(n38326), .B(n38189), .Z(n38191) );
  XNOR U38492 ( .A(n38400), .B(a[125]), .Z(n38244) );
  NANDN U38493 ( .A(n38273), .B(n38244), .Z(n38190) );
  NAND U38494 ( .A(n38191), .B(n38190), .Z(n38256) );
  XNOR U38495 ( .A(n38192), .B(n38235), .Z(n38238) );
  NANDN U38496 ( .A(n38193), .B(b[63]), .Z(n38237) );
  XOR U38497 ( .A(n38238), .B(n38237), .Z(n38231) );
  XNOR U38498 ( .A(n38463), .B(b[57]), .Z(n38248) );
  NANDN U38499 ( .A(n965), .B(n38248), .Z(n38197) );
  NANDN U38500 ( .A(n38195), .B(n38194), .Z(n38196) );
  NAND U38501 ( .A(n38197), .B(n38196), .Z(n38229) );
  XNOR U38502 ( .A(n984), .B(a[123]), .Z(n38241) );
  NANDN U38503 ( .A(n38371), .B(n38241), .Z(n38200) );
  NANDN U38504 ( .A(n38198), .B(n38369), .Z(n38199) );
  AND U38505 ( .A(n38200), .B(n38199), .Z(n38230) );
  XNOR U38506 ( .A(n38229), .B(n38230), .Z(n38232) );
  XOR U38507 ( .A(n38231), .B(n38232), .Z(n38255) );
  XOR U38508 ( .A(n38256), .B(n38255), .Z(n38257) );
  XNOR U38509 ( .A(n38258), .B(n38257), .Z(n38226) );
  NANDN U38510 ( .A(n38235), .B(n38201), .Z(n38205) );
  NANDN U38511 ( .A(n38203), .B(n38202), .Z(n38204) );
  NAND U38512 ( .A(n38205), .B(n38204), .Z(n38224) );
  NANDN U38513 ( .A(n38207), .B(n38206), .Z(n38211) );
  NAND U38514 ( .A(n38209), .B(n38208), .Z(n38210) );
  AND U38515 ( .A(n38211), .B(n38210), .Z(n38223) );
  XNOR U38516 ( .A(n38224), .B(n38223), .Z(n38225) );
  XNOR U38517 ( .A(n38226), .B(n38225), .Z(n38220) );
  XOR U38518 ( .A(n38219), .B(n38220), .Z(n38261) );
  XOR U38519 ( .A(n38261), .B(n38262), .Z(n38216) );
  XOR U38520 ( .A(n38263), .B(n38216), .Z(n38265) );
  XNOR U38521 ( .A(n38266), .B(n38265), .Z(c[247]) );
  OR U38522 ( .A(n38218), .B(n38217), .Z(n38222) );
  NANDN U38523 ( .A(n38220), .B(n38219), .Z(n38221) );
  NAND U38524 ( .A(n38222), .B(n38221), .Z(n38271) );
  NANDN U38525 ( .A(n38224), .B(n38223), .Z(n38228) );
  NAND U38526 ( .A(n38226), .B(n38225), .Z(n38227) );
  NAND U38527 ( .A(n38228), .B(n38227), .Z(n38302) );
  NANDN U38528 ( .A(n38230), .B(n38229), .Z(n38234) );
  NAND U38529 ( .A(n38232), .B(n38231), .Z(n38233) );
  NAND U38530 ( .A(n38234), .B(n38233), .Z(n38293) );
  NANDN U38531 ( .A(n38236), .B(n38235), .Z(n38240) );
  OR U38532 ( .A(n38238), .B(n38237), .Z(n38239) );
  NAND U38533 ( .A(n38240), .B(n38239), .Z(n38290) );
  XOR U38534 ( .A(b[61]), .B(n38321), .Z(n38281) );
  OR U38535 ( .A(n38281), .B(n38371), .Z(n38243) );
  NAND U38536 ( .A(n38241), .B(n38369), .Z(n38242) );
  AND U38537 ( .A(n38243), .B(n38242), .Z(n38287) );
  NAND U38538 ( .A(n38326), .B(n38244), .Z(n38246) );
  XOR U38539 ( .A(n38400), .B(n987), .Z(n38272) );
  NANDN U38540 ( .A(n38273), .B(n38272), .Z(n38245) );
  AND U38541 ( .A(n38246), .B(n38245), .Z(n38288) );
  XNOR U38542 ( .A(n38290), .B(n38289), .Z(n38294) );
  XNOR U38543 ( .A(n38293), .B(n38294), .Z(n38295) );
  XNOR U38544 ( .A(n983), .B(n38247), .Z(n38250) );
  OR U38545 ( .A(n38248), .B(n964), .Z(n38249) );
  NAND U38546 ( .A(n38250), .B(n38249), .Z(n38278) );
  AND U38547 ( .A(a[120]), .B(b[63]), .Z(n38331) );
  XOR U38548 ( .A(n985), .B(n38251), .Z(n38284) );
  NAND U38549 ( .A(n38422), .B(n38284), .Z(n38254) );
  NANDN U38550 ( .A(n38252), .B(n38423), .Z(n38253) );
  AND U38551 ( .A(n38254), .B(n38253), .Z(n38276) );
  XOR U38552 ( .A(n38331), .B(n38276), .Z(n38277) );
  XOR U38553 ( .A(n38278), .B(n38277), .Z(n38296) );
  XOR U38554 ( .A(n38295), .B(n38296), .Z(n38299) );
  NAND U38555 ( .A(n38256), .B(n38255), .Z(n38260) );
  NAND U38556 ( .A(n38258), .B(n38257), .Z(n38259) );
  NAND U38557 ( .A(n38260), .B(n38259), .Z(n38300) );
  XNOR U38558 ( .A(n38299), .B(n38300), .Z(n38301) );
  XNOR U38559 ( .A(n38302), .B(n38301), .Z(n38269) );
  XOR U38560 ( .A(n38269), .B(n38270), .Z(n38264) );
  XNOR U38561 ( .A(n38271), .B(n38264), .Z(n38268) );
  NANDN U38562 ( .A(n38266), .B(n38265), .Z(n38267) );
  XOR U38563 ( .A(n38268), .B(n38267), .Z(c[248]) );
  OR U38564 ( .A(n38268), .B(n38267), .Z(n38345) );
  NAND U38565 ( .A(n38326), .B(n38272), .Z(n38275) );
  XOR U38566 ( .A(n38463), .B(n38400), .Z(n38325) );
  NANDN U38567 ( .A(n38273), .B(n38325), .Z(n38274) );
  NAND U38568 ( .A(n38275), .B(n38274), .Z(n38338) );
  OR U38569 ( .A(n38331), .B(n38276), .Z(n38280) );
  NANDN U38570 ( .A(n38278), .B(n38277), .Z(n38279) );
  AND U38571 ( .A(n38280), .B(n38279), .Z(n38339) );
  XNOR U38572 ( .A(n38338), .B(n38339), .Z(n38340) );
  NANDN U38573 ( .A(n38281), .B(n38369), .Z(n38283) );
  XNOR U38574 ( .A(b[61]), .B(a[125]), .Z(n38335) );
  OR U38575 ( .A(n38335), .B(n38371), .Z(n38282) );
  AND U38576 ( .A(n38283), .B(n38282), .Z(n38315) );
  XNOR U38577 ( .A(b[63]), .B(a[123]), .Z(n38322) );
  NANDN U38578 ( .A(n38322), .B(n38422), .Z(n38286) );
  NAND U38579 ( .A(n38284), .B(n38423), .Z(n38285) );
  AND U38580 ( .A(n38286), .B(n38285), .Z(n38316) );
  XOR U38581 ( .A(n38315), .B(n38316), .Z(n38317) );
  NANDN U38582 ( .A(n985), .B(a[121]), .Z(n38330) );
  XNOR U38583 ( .A(n38329), .B(n38330), .Z(n38332) );
  XOR U38584 ( .A(n38331), .B(n38332), .Z(n38318) );
  XOR U38585 ( .A(n38317), .B(n38318), .Z(n38341) );
  XOR U38586 ( .A(n38340), .B(n38341), .Z(n38312) );
  OR U38587 ( .A(n38288), .B(n38287), .Z(n38292) );
  NAND U38588 ( .A(n38290), .B(n38289), .Z(n38291) );
  NAND U38589 ( .A(n38292), .B(n38291), .Z(n38310) );
  NANDN U38590 ( .A(n38294), .B(n38293), .Z(n38298) );
  NANDN U38591 ( .A(n38296), .B(n38295), .Z(n38297) );
  AND U38592 ( .A(n38298), .B(n38297), .Z(n38309) );
  XNOR U38593 ( .A(n38310), .B(n38309), .Z(n38311) );
  XNOR U38594 ( .A(n38312), .B(n38311), .Z(n38306) );
  NANDN U38595 ( .A(n38300), .B(n38299), .Z(n38304) );
  NAND U38596 ( .A(n38302), .B(n38301), .Z(n38303) );
  AND U38597 ( .A(n38304), .B(n38303), .Z(n38307) );
  XOR U38598 ( .A(n38306), .B(n38307), .Z(n38305) );
  XOR U38599 ( .A(n38308), .B(n38305), .Z(n38344) );
  XNOR U38600 ( .A(n38345), .B(n38344), .Z(c[249]) );
  NANDN U38601 ( .A(n38310), .B(n38309), .Z(n38314) );
  NAND U38602 ( .A(n38312), .B(n38311), .Z(n38313) );
  NAND U38603 ( .A(n38314), .B(n38313), .Z(n38349) );
  OR U38604 ( .A(n38316), .B(n38315), .Z(n38320) );
  NANDN U38605 ( .A(n38318), .B(n38317), .Z(n38319) );
  NAND U38606 ( .A(n38320), .B(n38319), .Z(n38377) );
  XOR U38607 ( .A(b[63]), .B(n38321), .Z(n38366) );
  NANDN U38608 ( .A(n38366), .B(n38422), .Z(n38324) );
  NANDN U38609 ( .A(n38322), .B(n38423), .Z(n38323) );
  NAND U38610 ( .A(n38324), .B(n38323), .Z(n38361) );
  NAND U38611 ( .A(n38326), .B(n38325), .Z(n38328) );
  ANDN U38612 ( .B(n38328), .A(n38327), .Z(n38360) );
  AND U38613 ( .A(b[63]), .B(a[122]), .Z(n38393) );
  XNOR U38614 ( .A(n38360), .B(n38393), .Z(n38362) );
  XNOR U38615 ( .A(n38361), .B(n38362), .Z(n38354) );
  OR U38616 ( .A(n38330), .B(n38329), .Z(n38334) );
  NANDN U38617 ( .A(n38332), .B(n38331), .Z(n38333) );
  NAND U38618 ( .A(n38334), .B(n38333), .Z(n38355) );
  XOR U38619 ( .A(n38354), .B(n38355), .Z(n38356) );
  NANDN U38620 ( .A(n38335), .B(n38369), .Z(n38337) );
  XOR U38621 ( .A(b[61]), .B(n987), .Z(n38370) );
  OR U38622 ( .A(n38370), .B(n38371), .Z(n38336) );
  NAND U38623 ( .A(n38337), .B(n38336), .Z(n38357) );
  XOR U38624 ( .A(n38356), .B(n38357), .Z(n38374) );
  NANDN U38625 ( .A(n38339), .B(n38338), .Z(n38343) );
  NANDN U38626 ( .A(n38341), .B(n38340), .Z(n38342) );
  AND U38627 ( .A(n38343), .B(n38342), .Z(n38375) );
  XNOR U38628 ( .A(n38374), .B(n38375), .Z(n38376) );
  XOR U38629 ( .A(n38377), .B(n38376), .Z(n38348) );
  XOR U38630 ( .A(n38349), .B(n38348), .Z(n38351) );
  XNOR U38631 ( .A(n38350), .B(n38351), .Z(n38346) );
  NANDN U38632 ( .A(n38345), .B(n38344), .Z(n38347) );
  XNOR U38633 ( .A(n38346), .B(n38347), .Z(c[250]) );
  NANDN U38634 ( .A(n38347), .B(n38346), .Z(n38382) );
  NANDN U38635 ( .A(n38349), .B(n38348), .Z(n38353) );
  NANDN U38636 ( .A(n38351), .B(n38350), .Z(n38352) );
  AND U38637 ( .A(n38353), .B(n38352), .Z(n38385) );
  OR U38638 ( .A(n38355), .B(n38354), .Z(n38359) );
  NANDN U38639 ( .A(n38357), .B(n38356), .Z(n38358) );
  NAND U38640 ( .A(n38359), .B(n38358), .Z(n38389) );
  OR U38641 ( .A(n38360), .B(n38393), .Z(n38364) );
  NANDN U38642 ( .A(n38362), .B(n38361), .Z(n38363) );
  NAND U38643 ( .A(n38364), .B(n38363), .Z(n38387) );
  NANDN U38644 ( .A(n983), .B(b[58]), .Z(n38365) );
  AND U38645 ( .A(n38365), .B(b[59]), .Z(n38390) );
  NANDN U38646 ( .A(n985), .B(a[123]), .Z(n38391) );
  XOR U38647 ( .A(n38390), .B(n38391), .Z(n38392) );
  XOR U38648 ( .A(n38393), .B(n38392), .Z(n38406) );
  XNOR U38649 ( .A(n985), .B(a[125]), .Z(n38396) );
  NAND U38650 ( .A(n38396), .B(n38422), .Z(n38368) );
  NANDN U38651 ( .A(n38366), .B(n38423), .Z(n38367) );
  NAND U38652 ( .A(n38368), .B(n38367), .Z(n38405) );
  XOR U38653 ( .A(n38406), .B(n38405), .Z(n38407) );
  NANDN U38654 ( .A(n38370), .B(n38369), .Z(n38373) );
  XOR U38655 ( .A(b[61]), .B(n38463), .Z(n38401) );
  OR U38656 ( .A(n38401), .B(n38371), .Z(n38372) );
  AND U38657 ( .A(n38373), .B(n38372), .Z(n38408) );
  XOR U38658 ( .A(n38407), .B(n38408), .Z(n38386) );
  XNOR U38659 ( .A(n38387), .B(n38386), .Z(n38388) );
  XNOR U38660 ( .A(n38389), .B(n38388), .Z(n38383) );
  NANDN U38661 ( .A(n38375), .B(n38374), .Z(n38379) );
  NAND U38662 ( .A(n38377), .B(n38376), .Z(n38378) );
  AND U38663 ( .A(n38379), .B(n38378), .Z(n38384) );
  XOR U38664 ( .A(n38383), .B(n38384), .Z(n38380) );
  XNOR U38665 ( .A(n38385), .B(n38380), .Z(n38381) );
  XOR U38666 ( .A(n38382), .B(n38381), .Z(c[251]) );
  OR U38667 ( .A(n38382), .B(n38381), .Z(n38413) );
  OR U38668 ( .A(n38391), .B(n38390), .Z(n38395) );
  NAND U38669 ( .A(n38393), .B(n38392), .Z(n38394) );
  NAND U38670 ( .A(n38395), .B(n38394), .Z(n38427) );
  XNOR U38671 ( .A(n985), .B(a[126]), .Z(n38424) );
  NAND U38672 ( .A(n38424), .B(n38422), .Z(n38398) );
  NAND U38673 ( .A(n38396), .B(n38423), .Z(n38397) );
  NAND U38674 ( .A(n38398), .B(n38397), .Z(n38419) );
  XOR U38675 ( .A(n984), .B(n38399), .Z(n38404) );
  XOR U38676 ( .A(b[60]), .B(n38400), .Z(n38402) );
  NAND U38677 ( .A(n38402), .B(n38401), .Z(n38403) );
  AND U38678 ( .A(n38404), .B(n38403), .Z(n38417) );
  AND U38679 ( .A(a[124]), .B(b[63]), .Z(n38439) );
  XNOR U38680 ( .A(n38417), .B(n38439), .Z(n38418) );
  XNOR U38681 ( .A(n38419), .B(n38418), .Z(n38428) );
  XNOR U38682 ( .A(n38427), .B(n38428), .Z(n38429) );
  OR U38683 ( .A(n38406), .B(n38405), .Z(n38410) );
  NAND U38684 ( .A(n38408), .B(n38407), .Z(n38409) );
  NAND U38685 ( .A(n38410), .B(n38409), .Z(n38430) );
  XOR U38686 ( .A(n38429), .B(n38430), .Z(n38415) );
  XNOR U38687 ( .A(n38414), .B(n38415), .Z(n38411) );
  XOR U38688 ( .A(n38416), .B(n38411), .Z(n38412) );
  XNOR U38689 ( .A(n38413), .B(n38412), .Z(c[252]) );
  NANDN U38690 ( .A(n38413), .B(n38412), .Z(n38460) );
  XOR U38691 ( .A(n38440), .B(n38439), .Z(n38442) );
  NANDN U38692 ( .A(n985), .B(a[125]), .Z(n38441) );
  XNOR U38693 ( .A(n38442), .B(n38441), .Z(n38449) );
  NANDN U38694 ( .A(n38439), .B(n38417), .Z(n38421) );
  NAND U38695 ( .A(n38419), .B(n38418), .Z(n38420) );
  NAND U38696 ( .A(n38421), .B(n38420), .Z(n38447) );
  XOR U38697 ( .A(b[63]), .B(n38463), .Z(n38435) );
  NANDN U38698 ( .A(n38435), .B(n38422), .Z(n38426) );
  NAND U38699 ( .A(n38424), .B(n38423), .Z(n38425) );
  AND U38700 ( .A(n38426), .B(n38425), .Z(n38446) );
  XNOR U38701 ( .A(n38447), .B(n38446), .Z(n38448) );
  XOR U38702 ( .A(n38449), .B(n38448), .Z(n38452) );
  NANDN U38703 ( .A(n38428), .B(n38427), .Z(n38432) );
  NANDN U38704 ( .A(n38430), .B(n38429), .Z(n38431) );
  AND U38705 ( .A(n38432), .B(n38431), .Z(n38453) );
  XNOR U38706 ( .A(n38452), .B(n38453), .Z(n38454) );
  XOR U38707 ( .A(n38455), .B(n38454), .Z(n38459) );
  XOR U38708 ( .A(n38460), .B(n38459), .Z(c[253]) );
  NANDN U38709 ( .A(n38433), .B(b[61]), .Z(n38434) );
  XOR U38710 ( .A(n985), .B(n38434), .Z(n38438) );
  XOR U38711 ( .A(n984), .B(b[62]), .Z(n38436) );
  NAND U38712 ( .A(n38436), .B(n38435), .Z(n38437) );
  NAND U38713 ( .A(n38438), .B(n38437), .Z(n38468) );
  NANDN U38714 ( .A(n38440), .B(n38439), .Z(n38444) );
  OR U38715 ( .A(n38442), .B(n38441), .Z(n38443) );
  NAND U38716 ( .A(n38444), .B(n38443), .Z(n38469) );
  AND U38717 ( .A(a[126]), .B(b[63]), .Z(n38467) );
  XNOR U38718 ( .A(n38469), .B(n38467), .Z(n38445) );
  XOR U38719 ( .A(n38468), .B(n38445), .Z(n38465) );
  NANDN U38720 ( .A(n38447), .B(n38446), .Z(n38451) );
  NAND U38721 ( .A(n38449), .B(n38448), .Z(n38450) );
  AND U38722 ( .A(n38451), .B(n38450), .Z(n38464) );
  NAND U38723 ( .A(n38453), .B(n38452), .Z(n38457) );
  OR U38724 ( .A(n38455), .B(n38454), .Z(n38456) );
  AND U38725 ( .A(n38457), .B(n38456), .Z(n38466) );
  XOR U38726 ( .A(n38464), .B(n38466), .Z(n38458) );
  XNOR U38727 ( .A(n38465), .B(n38458), .Z(n38471) );
  OR U38728 ( .A(n38460), .B(n38459), .Z(n38470) );
  XNOR U38729 ( .A(n38471), .B(n38470), .Z(c[254]) );
endmodule

