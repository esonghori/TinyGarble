
module mult_N64_CC32 ( clk, rst, a, b, c );
  input [63:0] a;
  input [1:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822;
  wire   [127:0] sreg;

  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U5 ( .A(n800), .B(n798), .Z(n1) );
  XOR U6 ( .A(n800), .B(n798), .Z(n2) );
  NANDN U7 ( .A(n799), .B(n2), .Z(n3) );
  NAND U8 ( .A(n1), .B(n3), .Z(n807) );
  NAND U9 ( .A(n807), .B(n805), .Z(n4) );
  XOR U10 ( .A(n807), .B(n805), .Z(n5) );
  NANDN U11 ( .A(n806), .B(n5), .Z(n6) );
  NAND U12 ( .A(n4), .B(n6), .Z(n815) );
  OR U13 ( .A(n392), .B(n394), .Z(n7) );
  NANDN U14 ( .A(n393), .B(n7), .Z(n8) );
  NANDN U15 ( .A(n394), .B(n393), .Z(n9) );
  NAND U16 ( .A(n391), .B(n9), .Z(n10) );
  NAND U17 ( .A(n8), .B(n10), .Z(n401) );
  NAND U18 ( .A(n415), .B(n413), .Z(n11) );
  XOR U19 ( .A(n415), .B(n413), .Z(n12) );
  NANDN U20 ( .A(n414), .B(n12), .Z(n13) );
  NAND U21 ( .A(n11), .B(n13), .Z(n422) );
  NAND U22 ( .A(n436), .B(n434), .Z(n14) );
  XOR U23 ( .A(n436), .B(n434), .Z(n15) );
  NANDN U24 ( .A(n435), .B(n15), .Z(n16) );
  NAND U25 ( .A(n14), .B(n16), .Z(n443) );
  NAND U26 ( .A(n457), .B(n455), .Z(n17) );
  XOR U27 ( .A(n457), .B(n455), .Z(n18) );
  NANDN U28 ( .A(n456), .B(n18), .Z(n19) );
  NAND U29 ( .A(n17), .B(n19), .Z(n464) );
  NAND U30 ( .A(n478), .B(n476), .Z(n20) );
  XOR U31 ( .A(n478), .B(n476), .Z(n21) );
  NANDN U32 ( .A(n477), .B(n21), .Z(n22) );
  NAND U33 ( .A(n20), .B(n22), .Z(n485) );
  NAND U34 ( .A(n499), .B(n497), .Z(n23) );
  XOR U35 ( .A(n499), .B(n497), .Z(n24) );
  NANDN U36 ( .A(n498), .B(n24), .Z(n25) );
  NAND U37 ( .A(n23), .B(n25), .Z(n506) );
  NAND U38 ( .A(n520), .B(n518), .Z(n26) );
  XOR U39 ( .A(n520), .B(n518), .Z(n27) );
  NANDN U40 ( .A(n519), .B(n27), .Z(n28) );
  NAND U41 ( .A(n26), .B(n28), .Z(n527) );
  NAND U42 ( .A(n541), .B(n539), .Z(n29) );
  XOR U43 ( .A(n541), .B(n539), .Z(n30) );
  NANDN U44 ( .A(n540), .B(n30), .Z(n31) );
  NAND U45 ( .A(n29), .B(n31), .Z(n548) );
  NAND U46 ( .A(n562), .B(n560), .Z(n32) );
  XOR U47 ( .A(n562), .B(n560), .Z(n33) );
  NANDN U48 ( .A(n561), .B(n33), .Z(n34) );
  NAND U49 ( .A(n32), .B(n34), .Z(n571) );
  NAND U50 ( .A(n583), .B(n581), .Z(n35) );
  XOR U51 ( .A(n583), .B(n581), .Z(n36) );
  NANDN U52 ( .A(n582), .B(n36), .Z(n37) );
  NAND U53 ( .A(n35), .B(n37), .Z(n590) );
  NAND U54 ( .A(n604), .B(n602), .Z(n38) );
  XOR U55 ( .A(n604), .B(n602), .Z(n39) );
  NANDN U56 ( .A(n603), .B(n39), .Z(n40) );
  NAND U57 ( .A(n38), .B(n40), .Z(n611) );
  NAND U58 ( .A(n625), .B(n623), .Z(n41) );
  XOR U59 ( .A(n625), .B(n623), .Z(n42) );
  NANDN U60 ( .A(n624), .B(n42), .Z(n43) );
  NAND U61 ( .A(n41), .B(n43), .Z(n632) );
  NAND U62 ( .A(n646), .B(n644), .Z(n44) );
  XOR U63 ( .A(n646), .B(n644), .Z(n45) );
  NANDN U64 ( .A(n645), .B(n45), .Z(n46) );
  NAND U65 ( .A(n44), .B(n46), .Z(n653) );
  NAND U66 ( .A(n667), .B(n665), .Z(n47) );
  XOR U67 ( .A(n667), .B(n665), .Z(n48) );
  NANDN U68 ( .A(n666), .B(n48), .Z(n49) );
  NAND U69 ( .A(n47), .B(n49), .Z(n674) );
  NAND U70 ( .A(n688), .B(n686), .Z(n50) );
  XOR U71 ( .A(n688), .B(n686), .Z(n51) );
  NANDN U72 ( .A(n687), .B(n51), .Z(n52) );
  NAND U73 ( .A(n50), .B(n52), .Z(n695) );
  NAND U74 ( .A(n709), .B(n707), .Z(n53) );
  XOR U75 ( .A(n709), .B(n707), .Z(n54) );
  NANDN U76 ( .A(n708), .B(n54), .Z(n55) );
  NAND U77 ( .A(n53), .B(n55), .Z(n716) );
  NAND U78 ( .A(n730), .B(n728), .Z(n56) );
  XOR U79 ( .A(n730), .B(n728), .Z(n57) );
  NANDN U80 ( .A(n729), .B(n57), .Z(n58) );
  NAND U81 ( .A(n56), .B(n58), .Z(n737) );
  NAND U82 ( .A(n751), .B(n749), .Z(n59) );
  XOR U83 ( .A(n751), .B(n749), .Z(n60) );
  NANDN U84 ( .A(n750), .B(n60), .Z(n61) );
  NAND U85 ( .A(n59), .B(n61), .Z(n758) );
  NAND U86 ( .A(n772), .B(n770), .Z(n62) );
  XOR U87 ( .A(n772), .B(n770), .Z(n63) );
  NANDN U88 ( .A(n771), .B(n63), .Z(n64) );
  NAND U89 ( .A(n62), .B(n64), .Z(n779) );
  NAND U90 ( .A(n793), .B(n791), .Z(n65) );
  XOR U91 ( .A(n793), .B(n791), .Z(n66) );
  NANDN U92 ( .A(n792), .B(n66), .Z(n67) );
  NAND U93 ( .A(n65), .B(n67), .Z(n800) );
  NAND U94 ( .A(n411), .B(n410), .Z(n68) );
  XOR U95 ( .A(n411), .B(n410), .Z(n69) );
  NANDN U96 ( .A(sreg[67]), .B(n69), .Z(n70) );
  NAND U97 ( .A(n68), .B(n70), .Z(n418) );
  NAND U98 ( .A(n432), .B(n431), .Z(n71) );
  XOR U99 ( .A(n432), .B(n431), .Z(n72) );
  NANDN U100 ( .A(sreg[70]), .B(n72), .Z(n73) );
  NAND U101 ( .A(n71), .B(n73), .Z(n439) );
  NAND U102 ( .A(n453), .B(n452), .Z(n74) );
  XOR U103 ( .A(n453), .B(n452), .Z(n75) );
  NANDN U104 ( .A(sreg[73]), .B(n75), .Z(n76) );
  NAND U105 ( .A(n74), .B(n76), .Z(n460) );
  NAND U106 ( .A(n474), .B(n473), .Z(n77) );
  XOR U107 ( .A(n474), .B(n473), .Z(n78) );
  NANDN U108 ( .A(sreg[76]), .B(n78), .Z(n79) );
  NAND U109 ( .A(n77), .B(n79), .Z(n481) );
  NAND U110 ( .A(n495), .B(n494), .Z(n80) );
  XOR U111 ( .A(n495), .B(n494), .Z(n81) );
  NANDN U112 ( .A(sreg[79]), .B(n81), .Z(n82) );
  NAND U113 ( .A(n80), .B(n82), .Z(n502) );
  NAND U114 ( .A(n516), .B(n515), .Z(n83) );
  XOR U115 ( .A(n516), .B(n515), .Z(n84) );
  NANDN U116 ( .A(sreg[82]), .B(n84), .Z(n85) );
  NAND U117 ( .A(n83), .B(n85), .Z(n523) );
  NAND U118 ( .A(n537), .B(n536), .Z(n86) );
  XOR U119 ( .A(n537), .B(n536), .Z(n87) );
  NANDN U120 ( .A(sreg[85]), .B(n87), .Z(n88) );
  NAND U121 ( .A(n86), .B(n88), .Z(n544) );
  NAND U122 ( .A(n558), .B(n557), .Z(n89) );
  XOR U123 ( .A(n558), .B(n557), .Z(n90) );
  NANDN U124 ( .A(sreg[88]), .B(n90), .Z(n91) );
  NAND U125 ( .A(n89), .B(n91), .Z(n565) );
  XOR U126 ( .A(n579), .B(sreg[91]), .Z(n92) );
  NANDN U127 ( .A(n578), .B(n92), .Z(n93) );
  NAND U128 ( .A(n579), .B(sreg[91]), .Z(n94) );
  AND U129 ( .A(n93), .B(n94), .Z(n586) );
  NAND U130 ( .A(n600), .B(n599), .Z(n95) );
  XOR U131 ( .A(n600), .B(n599), .Z(n96) );
  NANDN U132 ( .A(sreg[94]), .B(n96), .Z(n97) );
  NAND U133 ( .A(n95), .B(n97), .Z(n607) );
  NAND U134 ( .A(n621), .B(n620), .Z(n98) );
  XOR U135 ( .A(n621), .B(n620), .Z(n99) );
  NANDN U136 ( .A(sreg[97]), .B(n99), .Z(n100) );
  NAND U137 ( .A(n98), .B(n100), .Z(n628) );
  NAND U138 ( .A(n642), .B(n641), .Z(n101) );
  XOR U139 ( .A(n642), .B(n641), .Z(n102) );
  NANDN U140 ( .A(sreg[100]), .B(n102), .Z(n103) );
  NAND U141 ( .A(n101), .B(n103), .Z(n649) );
  NAND U142 ( .A(n663), .B(n662), .Z(n104) );
  XOR U143 ( .A(n663), .B(n662), .Z(n105) );
  NANDN U144 ( .A(sreg[103]), .B(n105), .Z(n106) );
  NAND U145 ( .A(n104), .B(n106), .Z(n670) );
  NAND U146 ( .A(n684), .B(n683), .Z(n107) );
  XOR U147 ( .A(n684), .B(n683), .Z(n108) );
  NANDN U148 ( .A(sreg[106]), .B(n108), .Z(n109) );
  NAND U149 ( .A(n107), .B(n109), .Z(n691) );
  NAND U150 ( .A(n705), .B(n704), .Z(n110) );
  XOR U151 ( .A(n705), .B(n704), .Z(n111) );
  NANDN U152 ( .A(sreg[109]), .B(n111), .Z(n112) );
  NAND U153 ( .A(n110), .B(n112), .Z(n712) );
  NAND U154 ( .A(n726), .B(n725), .Z(n113) );
  XOR U155 ( .A(n726), .B(n725), .Z(n114) );
  NANDN U156 ( .A(sreg[112]), .B(n114), .Z(n115) );
  NAND U157 ( .A(n113), .B(n115), .Z(n733) );
  NAND U158 ( .A(n747), .B(n746), .Z(n116) );
  XOR U159 ( .A(n747), .B(n746), .Z(n117) );
  NANDN U160 ( .A(sreg[115]), .B(n117), .Z(n118) );
  NAND U161 ( .A(n116), .B(n118), .Z(n754) );
  NAND U162 ( .A(n768), .B(n767), .Z(n119) );
  XOR U163 ( .A(n768), .B(n767), .Z(n120) );
  NANDN U164 ( .A(sreg[118]), .B(n120), .Z(n121) );
  NAND U165 ( .A(n119), .B(n121), .Z(n775) );
  NAND U166 ( .A(n789), .B(n788), .Z(n122) );
  XOR U167 ( .A(n789), .B(n788), .Z(n123) );
  NANDN U168 ( .A(sreg[121]), .B(n123), .Z(n124) );
  NAND U169 ( .A(n122), .B(n124), .Z(n796) );
  NAND U170 ( .A(n809), .B(n808), .Z(n125) );
  XOR U171 ( .A(n809), .B(n808), .Z(n126) );
  NANDN U172 ( .A(sreg[124]), .B(n126), .Z(n127) );
  NAND U173 ( .A(n125), .B(n127), .Z(n812) );
  NAND U174 ( .A(n401), .B(n399), .Z(n128) );
  XOR U175 ( .A(n401), .B(n399), .Z(n129) );
  NANDN U176 ( .A(n400), .B(n129), .Z(n130) );
  NAND U177 ( .A(n128), .B(n130), .Z(n408) );
  NAND U178 ( .A(n422), .B(n420), .Z(n131) );
  XOR U179 ( .A(n422), .B(n420), .Z(n132) );
  NANDN U180 ( .A(n421), .B(n132), .Z(n133) );
  NAND U181 ( .A(n131), .B(n133), .Z(n429) );
  NAND U182 ( .A(n443), .B(n441), .Z(n134) );
  XOR U183 ( .A(n443), .B(n441), .Z(n135) );
  NANDN U184 ( .A(n442), .B(n135), .Z(n136) );
  NAND U185 ( .A(n134), .B(n136), .Z(n450) );
  NAND U186 ( .A(n464), .B(n462), .Z(n137) );
  XOR U187 ( .A(n464), .B(n462), .Z(n138) );
  NANDN U188 ( .A(n463), .B(n138), .Z(n139) );
  NAND U189 ( .A(n137), .B(n139), .Z(n471) );
  NAND U190 ( .A(n485), .B(n483), .Z(n140) );
  XOR U191 ( .A(n485), .B(n483), .Z(n141) );
  NANDN U192 ( .A(n484), .B(n141), .Z(n142) );
  NAND U193 ( .A(n140), .B(n142), .Z(n492) );
  NAND U194 ( .A(n506), .B(n504), .Z(n143) );
  XOR U195 ( .A(n506), .B(n504), .Z(n144) );
  NANDN U196 ( .A(n505), .B(n144), .Z(n145) );
  NAND U197 ( .A(n143), .B(n145), .Z(n513) );
  NAND U198 ( .A(n527), .B(n525), .Z(n146) );
  XOR U199 ( .A(n527), .B(n525), .Z(n147) );
  NANDN U200 ( .A(n526), .B(n147), .Z(n148) );
  NAND U201 ( .A(n146), .B(n148), .Z(n534) );
  NAND U202 ( .A(n548), .B(n546), .Z(n149) );
  XOR U203 ( .A(n548), .B(n546), .Z(n150) );
  NANDN U204 ( .A(n547), .B(n150), .Z(n151) );
  NAND U205 ( .A(n149), .B(n151), .Z(n555) );
  NAND U206 ( .A(n571), .B(n569), .Z(n152) );
  XOR U207 ( .A(n571), .B(n569), .Z(n153) );
  NANDN U208 ( .A(n570), .B(n153), .Z(n154) );
  NAND U209 ( .A(n152), .B(n154), .Z(n576) );
  NAND U210 ( .A(n590), .B(n588), .Z(n155) );
  XOR U211 ( .A(n590), .B(n588), .Z(n156) );
  NANDN U212 ( .A(n589), .B(n156), .Z(n157) );
  NAND U213 ( .A(n155), .B(n157), .Z(n597) );
  NAND U214 ( .A(n611), .B(n609), .Z(n158) );
  XOR U215 ( .A(n611), .B(n609), .Z(n159) );
  NANDN U216 ( .A(n610), .B(n159), .Z(n160) );
  NAND U217 ( .A(n158), .B(n160), .Z(n618) );
  NAND U218 ( .A(n632), .B(n630), .Z(n161) );
  XOR U219 ( .A(n632), .B(n630), .Z(n162) );
  NANDN U220 ( .A(n631), .B(n162), .Z(n163) );
  NAND U221 ( .A(n161), .B(n163), .Z(n639) );
  NAND U222 ( .A(n653), .B(n651), .Z(n164) );
  XOR U223 ( .A(n653), .B(n651), .Z(n165) );
  NANDN U224 ( .A(n652), .B(n165), .Z(n166) );
  NAND U225 ( .A(n164), .B(n166), .Z(n660) );
  NAND U226 ( .A(n674), .B(n672), .Z(n167) );
  XOR U227 ( .A(n674), .B(n672), .Z(n168) );
  NANDN U228 ( .A(n673), .B(n168), .Z(n169) );
  NAND U229 ( .A(n167), .B(n169), .Z(n681) );
  NAND U230 ( .A(n695), .B(n693), .Z(n170) );
  XOR U231 ( .A(n695), .B(n693), .Z(n171) );
  NANDN U232 ( .A(n694), .B(n171), .Z(n172) );
  NAND U233 ( .A(n170), .B(n172), .Z(n702) );
  NAND U234 ( .A(n716), .B(n714), .Z(n173) );
  XOR U235 ( .A(n716), .B(n714), .Z(n174) );
  NANDN U236 ( .A(n715), .B(n174), .Z(n175) );
  NAND U237 ( .A(n173), .B(n175), .Z(n723) );
  NAND U238 ( .A(n737), .B(n735), .Z(n176) );
  XOR U239 ( .A(n737), .B(n735), .Z(n177) );
  NANDN U240 ( .A(n736), .B(n177), .Z(n178) );
  NAND U241 ( .A(n176), .B(n178), .Z(n744) );
  NAND U242 ( .A(n758), .B(n756), .Z(n179) );
  XOR U243 ( .A(n758), .B(n756), .Z(n180) );
  NANDN U244 ( .A(n757), .B(n180), .Z(n181) );
  NAND U245 ( .A(n179), .B(n181), .Z(n765) );
  NAND U246 ( .A(n779), .B(n777), .Z(n182) );
  XOR U247 ( .A(n779), .B(n777), .Z(n183) );
  NANDN U248 ( .A(n778), .B(n183), .Z(n184) );
  NAND U249 ( .A(n182), .B(n184), .Z(n786) );
  NAND U250 ( .A(n397), .B(n396), .Z(n185) );
  XOR U251 ( .A(n397), .B(n396), .Z(n186) );
  NANDN U252 ( .A(sreg[65]), .B(n186), .Z(n187) );
  NAND U253 ( .A(n185), .B(n187), .Z(n404) );
  NAND U254 ( .A(n418), .B(n417), .Z(n188) );
  XOR U255 ( .A(n418), .B(n417), .Z(n189) );
  NANDN U256 ( .A(sreg[68]), .B(n189), .Z(n190) );
  NAND U257 ( .A(n188), .B(n190), .Z(n425) );
  NAND U258 ( .A(n439), .B(n438), .Z(n191) );
  XOR U259 ( .A(n439), .B(n438), .Z(n192) );
  NANDN U260 ( .A(sreg[71]), .B(n192), .Z(n193) );
  NAND U261 ( .A(n191), .B(n193), .Z(n446) );
  NAND U262 ( .A(n460), .B(n459), .Z(n194) );
  XOR U263 ( .A(n460), .B(n459), .Z(n195) );
  NANDN U264 ( .A(sreg[74]), .B(n195), .Z(n196) );
  NAND U265 ( .A(n194), .B(n196), .Z(n467) );
  NAND U266 ( .A(n481), .B(n480), .Z(n197) );
  XOR U267 ( .A(n481), .B(n480), .Z(n198) );
  NANDN U268 ( .A(sreg[77]), .B(n198), .Z(n199) );
  NAND U269 ( .A(n197), .B(n199), .Z(n488) );
  NAND U270 ( .A(n502), .B(n501), .Z(n200) );
  XOR U271 ( .A(n502), .B(n501), .Z(n201) );
  NANDN U272 ( .A(sreg[80]), .B(n201), .Z(n202) );
  NAND U273 ( .A(n200), .B(n202), .Z(n509) );
  NAND U274 ( .A(n523), .B(n522), .Z(n203) );
  XOR U275 ( .A(n523), .B(n522), .Z(n204) );
  NANDN U276 ( .A(sreg[83]), .B(n204), .Z(n205) );
  NAND U277 ( .A(n203), .B(n205), .Z(n530) );
  NAND U278 ( .A(n544), .B(n543), .Z(n206) );
  XOR U279 ( .A(n544), .B(n543), .Z(n207) );
  NANDN U280 ( .A(sreg[86]), .B(n207), .Z(n208) );
  NAND U281 ( .A(n206), .B(n208), .Z(n551) );
  NAND U282 ( .A(n565), .B(n564), .Z(n209) );
  XOR U283 ( .A(n565), .B(n564), .Z(n210) );
  NANDN U284 ( .A(sreg[89]), .B(n210), .Z(n211) );
  NAND U285 ( .A(n209), .B(n211), .Z(n568) );
  NAND U286 ( .A(n586), .B(n585), .Z(n212) );
  XOR U287 ( .A(n586), .B(n585), .Z(n213) );
  NANDN U288 ( .A(sreg[92]), .B(n213), .Z(n214) );
  NAND U289 ( .A(n212), .B(n214), .Z(n593) );
  NAND U290 ( .A(n607), .B(n606), .Z(n215) );
  XOR U291 ( .A(n607), .B(n606), .Z(n216) );
  NANDN U292 ( .A(sreg[95]), .B(n216), .Z(n217) );
  NAND U293 ( .A(n215), .B(n217), .Z(n614) );
  NAND U294 ( .A(n628), .B(n627), .Z(n218) );
  XOR U295 ( .A(n628), .B(n627), .Z(n219) );
  NANDN U296 ( .A(sreg[98]), .B(n219), .Z(n220) );
  NAND U297 ( .A(n218), .B(n220), .Z(n635) );
  NAND U298 ( .A(n649), .B(n648), .Z(n221) );
  XOR U299 ( .A(n649), .B(n648), .Z(n222) );
  NANDN U300 ( .A(sreg[101]), .B(n222), .Z(n223) );
  NAND U301 ( .A(n221), .B(n223), .Z(n656) );
  NAND U302 ( .A(n670), .B(n669), .Z(n224) );
  XOR U303 ( .A(n670), .B(n669), .Z(n225) );
  NANDN U304 ( .A(sreg[104]), .B(n225), .Z(n226) );
  NAND U305 ( .A(n224), .B(n226), .Z(n677) );
  NAND U306 ( .A(n691), .B(n690), .Z(n227) );
  XOR U307 ( .A(n691), .B(n690), .Z(n228) );
  NANDN U308 ( .A(sreg[107]), .B(n228), .Z(n229) );
  NAND U309 ( .A(n227), .B(n229), .Z(n698) );
  NAND U310 ( .A(n712), .B(n711), .Z(n230) );
  XOR U311 ( .A(n712), .B(n711), .Z(n231) );
  NANDN U312 ( .A(sreg[110]), .B(n231), .Z(n232) );
  NAND U313 ( .A(n230), .B(n232), .Z(n719) );
  NAND U314 ( .A(n733), .B(n732), .Z(n233) );
  XOR U315 ( .A(n733), .B(n732), .Z(n234) );
  NANDN U316 ( .A(sreg[113]), .B(n234), .Z(n235) );
  NAND U317 ( .A(n233), .B(n235), .Z(n740) );
  NAND U318 ( .A(n754), .B(n753), .Z(n236) );
  XOR U319 ( .A(n754), .B(n753), .Z(n237) );
  NANDN U320 ( .A(sreg[116]), .B(n237), .Z(n238) );
  NAND U321 ( .A(n236), .B(n238), .Z(n761) );
  NAND U322 ( .A(n775), .B(n774), .Z(n239) );
  XOR U323 ( .A(n775), .B(n774), .Z(n240) );
  NANDN U324 ( .A(sreg[119]), .B(n240), .Z(n241) );
  NAND U325 ( .A(n239), .B(n241), .Z(n782) );
  NAND U326 ( .A(n796), .B(n795), .Z(n242) );
  XOR U327 ( .A(n796), .B(n795), .Z(n243) );
  NANDN U328 ( .A(sreg[122]), .B(n243), .Z(n244) );
  NAND U329 ( .A(n242), .B(n244), .Z(n803) );
  NAND U330 ( .A(n812), .B(n811), .Z(n245) );
  XOR U331 ( .A(n812), .B(n811), .Z(n246) );
  NANDN U332 ( .A(sreg[125]), .B(n246), .Z(n247) );
  NAND U333 ( .A(n245), .B(n247), .Z(n821) );
  NAND U334 ( .A(n408), .B(n406), .Z(n248) );
  XOR U335 ( .A(n408), .B(n406), .Z(n249) );
  NANDN U336 ( .A(n407), .B(n249), .Z(n250) );
  NAND U337 ( .A(n248), .B(n250), .Z(n415) );
  NAND U338 ( .A(n429), .B(n427), .Z(n251) );
  XOR U339 ( .A(n429), .B(n427), .Z(n252) );
  NANDN U340 ( .A(n428), .B(n252), .Z(n253) );
  NAND U341 ( .A(n251), .B(n253), .Z(n436) );
  NAND U342 ( .A(n450), .B(n448), .Z(n254) );
  XOR U343 ( .A(n450), .B(n448), .Z(n255) );
  NANDN U344 ( .A(n449), .B(n255), .Z(n256) );
  NAND U345 ( .A(n254), .B(n256), .Z(n457) );
  NAND U346 ( .A(n471), .B(n469), .Z(n257) );
  XOR U347 ( .A(n471), .B(n469), .Z(n258) );
  NANDN U348 ( .A(n470), .B(n258), .Z(n259) );
  NAND U349 ( .A(n257), .B(n259), .Z(n478) );
  NAND U350 ( .A(n492), .B(n490), .Z(n260) );
  XOR U351 ( .A(n492), .B(n490), .Z(n261) );
  NANDN U352 ( .A(n491), .B(n261), .Z(n262) );
  NAND U353 ( .A(n260), .B(n262), .Z(n499) );
  NAND U354 ( .A(n513), .B(n511), .Z(n263) );
  XOR U355 ( .A(n513), .B(n511), .Z(n264) );
  NANDN U356 ( .A(n512), .B(n264), .Z(n265) );
  NAND U357 ( .A(n263), .B(n265), .Z(n520) );
  NAND U358 ( .A(n534), .B(n532), .Z(n266) );
  XOR U359 ( .A(n534), .B(n532), .Z(n267) );
  NANDN U360 ( .A(n533), .B(n267), .Z(n268) );
  NAND U361 ( .A(n266), .B(n268), .Z(n541) );
  NAND U362 ( .A(n555), .B(n553), .Z(n269) );
  XOR U363 ( .A(n555), .B(n553), .Z(n270) );
  NANDN U364 ( .A(n554), .B(n270), .Z(n271) );
  NAND U365 ( .A(n269), .B(n271), .Z(n562) );
  NAND U366 ( .A(n576), .B(n574), .Z(n272) );
  XOR U367 ( .A(n576), .B(n574), .Z(n273) );
  NANDN U368 ( .A(n575), .B(n273), .Z(n274) );
  NAND U369 ( .A(n272), .B(n274), .Z(n583) );
  NAND U370 ( .A(n597), .B(n595), .Z(n275) );
  XOR U371 ( .A(n597), .B(n595), .Z(n276) );
  NANDN U372 ( .A(n596), .B(n276), .Z(n277) );
  NAND U373 ( .A(n275), .B(n277), .Z(n604) );
  NAND U374 ( .A(n618), .B(n616), .Z(n278) );
  XOR U375 ( .A(n618), .B(n616), .Z(n279) );
  NANDN U376 ( .A(n617), .B(n279), .Z(n280) );
  NAND U377 ( .A(n278), .B(n280), .Z(n625) );
  NAND U378 ( .A(n639), .B(n637), .Z(n281) );
  XOR U379 ( .A(n639), .B(n637), .Z(n282) );
  NANDN U380 ( .A(n638), .B(n282), .Z(n283) );
  NAND U381 ( .A(n281), .B(n283), .Z(n646) );
  NAND U382 ( .A(n660), .B(n658), .Z(n284) );
  XOR U383 ( .A(n660), .B(n658), .Z(n285) );
  NANDN U384 ( .A(n659), .B(n285), .Z(n286) );
  NAND U385 ( .A(n284), .B(n286), .Z(n667) );
  NAND U386 ( .A(n681), .B(n679), .Z(n287) );
  XOR U387 ( .A(n681), .B(n679), .Z(n288) );
  NANDN U388 ( .A(n680), .B(n288), .Z(n289) );
  NAND U389 ( .A(n287), .B(n289), .Z(n688) );
  NAND U390 ( .A(n702), .B(n700), .Z(n290) );
  XOR U391 ( .A(n702), .B(n700), .Z(n291) );
  NANDN U392 ( .A(n701), .B(n291), .Z(n292) );
  NAND U393 ( .A(n290), .B(n292), .Z(n709) );
  NAND U394 ( .A(n723), .B(n721), .Z(n293) );
  XOR U395 ( .A(n723), .B(n721), .Z(n294) );
  NANDN U396 ( .A(n722), .B(n294), .Z(n295) );
  NAND U397 ( .A(n293), .B(n295), .Z(n730) );
  NAND U398 ( .A(n744), .B(n742), .Z(n296) );
  XOR U399 ( .A(n744), .B(n742), .Z(n297) );
  NANDN U400 ( .A(n743), .B(n297), .Z(n298) );
  NAND U401 ( .A(n296), .B(n298), .Z(n751) );
  NAND U402 ( .A(n765), .B(n763), .Z(n299) );
  XOR U403 ( .A(n765), .B(n763), .Z(n300) );
  NANDN U404 ( .A(n764), .B(n300), .Z(n301) );
  NAND U405 ( .A(n299), .B(n301), .Z(n772) );
  NAND U406 ( .A(n786), .B(n784), .Z(n302) );
  XOR U407 ( .A(n786), .B(n784), .Z(n303) );
  NANDN U408 ( .A(n785), .B(n303), .Z(n304) );
  NAND U409 ( .A(n302), .B(n304), .Z(n793) );
  NAND U410 ( .A(n404), .B(n403), .Z(n305) );
  XOR U411 ( .A(n404), .B(n403), .Z(n306) );
  NANDN U412 ( .A(sreg[66]), .B(n306), .Z(n307) );
  NAND U413 ( .A(n305), .B(n307), .Z(n411) );
  NAND U414 ( .A(n425), .B(n424), .Z(n308) );
  XOR U415 ( .A(n425), .B(n424), .Z(n309) );
  NANDN U416 ( .A(sreg[69]), .B(n309), .Z(n310) );
  NAND U417 ( .A(n308), .B(n310), .Z(n432) );
  NAND U418 ( .A(n446), .B(n445), .Z(n311) );
  XOR U419 ( .A(n446), .B(n445), .Z(n312) );
  NANDN U420 ( .A(sreg[72]), .B(n312), .Z(n313) );
  NAND U421 ( .A(n311), .B(n313), .Z(n453) );
  NAND U422 ( .A(n467), .B(n466), .Z(n314) );
  XOR U423 ( .A(n467), .B(n466), .Z(n315) );
  NANDN U424 ( .A(sreg[75]), .B(n315), .Z(n316) );
  NAND U425 ( .A(n314), .B(n316), .Z(n474) );
  NAND U426 ( .A(n488), .B(n487), .Z(n317) );
  XOR U427 ( .A(n488), .B(n487), .Z(n318) );
  NANDN U428 ( .A(sreg[78]), .B(n318), .Z(n319) );
  NAND U429 ( .A(n317), .B(n319), .Z(n495) );
  NAND U430 ( .A(n509), .B(n508), .Z(n320) );
  XOR U431 ( .A(n509), .B(n508), .Z(n321) );
  NANDN U432 ( .A(sreg[81]), .B(n321), .Z(n322) );
  NAND U433 ( .A(n320), .B(n322), .Z(n516) );
  NAND U434 ( .A(n530), .B(n529), .Z(n323) );
  XOR U435 ( .A(n530), .B(n529), .Z(n324) );
  NANDN U436 ( .A(sreg[84]), .B(n324), .Z(n325) );
  NAND U437 ( .A(n323), .B(n325), .Z(n537) );
  NAND U438 ( .A(n551), .B(n550), .Z(n326) );
  XOR U439 ( .A(n551), .B(n550), .Z(n327) );
  NANDN U440 ( .A(sreg[87]), .B(n327), .Z(n328) );
  NAND U441 ( .A(n326), .B(n328), .Z(n558) );
  NAND U442 ( .A(n568), .B(n567), .Z(n329) );
  XOR U443 ( .A(n568), .B(n567), .Z(n330) );
  NANDN U444 ( .A(sreg[90]), .B(n330), .Z(n331) );
  NAND U445 ( .A(n329), .B(n331), .Z(n578) );
  NAND U446 ( .A(n593), .B(n592), .Z(n332) );
  XOR U447 ( .A(n593), .B(n592), .Z(n333) );
  NANDN U448 ( .A(sreg[93]), .B(n333), .Z(n334) );
  NAND U449 ( .A(n332), .B(n334), .Z(n600) );
  NAND U450 ( .A(n614), .B(n613), .Z(n335) );
  XOR U451 ( .A(n614), .B(n613), .Z(n336) );
  NANDN U452 ( .A(sreg[96]), .B(n336), .Z(n337) );
  NAND U453 ( .A(n335), .B(n337), .Z(n621) );
  NAND U454 ( .A(n635), .B(n634), .Z(n338) );
  XOR U455 ( .A(n635), .B(n634), .Z(n339) );
  NANDN U456 ( .A(sreg[99]), .B(n339), .Z(n340) );
  NAND U457 ( .A(n338), .B(n340), .Z(n642) );
  NAND U458 ( .A(n656), .B(n655), .Z(n341) );
  XOR U459 ( .A(n656), .B(n655), .Z(n342) );
  NANDN U460 ( .A(sreg[102]), .B(n342), .Z(n343) );
  NAND U461 ( .A(n341), .B(n343), .Z(n663) );
  NAND U462 ( .A(n677), .B(n676), .Z(n344) );
  XOR U463 ( .A(n677), .B(n676), .Z(n345) );
  NANDN U464 ( .A(sreg[105]), .B(n345), .Z(n346) );
  NAND U465 ( .A(n344), .B(n346), .Z(n684) );
  NAND U466 ( .A(n698), .B(n697), .Z(n347) );
  XOR U467 ( .A(n698), .B(n697), .Z(n348) );
  NANDN U468 ( .A(sreg[108]), .B(n348), .Z(n349) );
  NAND U469 ( .A(n347), .B(n349), .Z(n705) );
  NAND U470 ( .A(n719), .B(n718), .Z(n350) );
  XOR U471 ( .A(n719), .B(n718), .Z(n351) );
  NANDN U472 ( .A(sreg[111]), .B(n351), .Z(n352) );
  NAND U473 ( .A(n350), .B(n352), .Z(n726) );
  NAND U474 ( .A(n740), .B(n739), .Z(n353) );
  XOR U475 ( .A(n740), .B(n739), .Z(n354) );
  NANDN U476 ( .A(sreg[114]), .B(n354), .Z(n355) );
  NAND U477 ( .A(n353), .B(n355), .Z(n747) );
  NAND U478 ( .A(n761), .B(n760), .Z(n356) );
  XOR U479 ( .A(n761), .B(n760), .Z(n357) );
  NANDN U480 ( .A(sreg[117]), .B(n357), .Z(n358) );
  NAND U481 ( .A(n356), .B(n358), .Z(n768) );
  NAND U482 ( .A(n782), .B(n781), .Z(n359) );
  XOR U483 ( .A(n782), .B(n781), .Z(n360) );
  NANDN U484 ( .A(sreg[120]), .B(n360), .Z(n361) );
  NAND U485 ( .A(n359), .B(n361), .Z(n789) );
  NAND U486 ( .A(n803), .B(n802), .Z(n362) );
  XOR U487 ( .A(n803), .B(n802), .Z(n363) );
  NANDN U488 ( .A(sreg[123]), .B(n363), .Z(n364) );
  NAND U489 ( .A(n362), .B(n364), .Z(n809) );
  XOR U490 ( .A(n822), .B(n821), .Z(n365) );
  NANDN U491 ( .A(n820), .B(n365), .Z(n366) );
  NAND U492 ( .A(n821), .B(n822), .Z(n367) );
  AND U493 ( .A(n366), .B(n367), .Z(c[127]) );
  AND U494 ( .A(b[0]), .B(a[0]), .Z(n368) );
  XOR U495 ( .A(n368), .B(sreg[62]), .Z(c[62]) );
  AND U496 ( .A(b[0]), .B(a[1]), .Z(n392) );
  NAND U497 ( .A(b[1]), .B(a[0]), .Z(n380) );
  XOR U498 ( .A(n392), .B(n380), .Z(n375) );
  AND U499 ( .A(n368), .B(sreg[62]), .Z(n374) );
  IV U500 ( .A(n374), .Z(n373) );
  XNOR U501 ( .A(sreg[63]), .B(n373), .Z(n369) );
  XNOR U502 ( .A(n375), .B(n369), .Z(c[63]) );
  ANDN U503 ( .B(n392), .A(n380), .Z(n394) );
  AND U504 ( .A(a[2]), .B(b[0]), .Z(n371) );
  NAND U505 ( .A(a[1]), .B(b[1]), .Z(n370) );
  XNOR U506 ( .A(n371), .B(n370), .Z(n372) );
  XNOR U507 ( .A(n394), .B(n372), .Z(n386) );
  IV U508 ( .A(n386), .Z(n384) );
  NANDN U509 ( .A(sreg[63]), .B(n373), .Z(n378) );
  AND U510 ( .A(sreg[63]), .B(n374), .Z(n376) );
  NANDN U511 ( .A(n376), .B(n375), .Z(n377) );
  AND U512 ( .A(n378), .B(n377), .Z(n385) );
  XNOR U513 ( .A(n384), .B(n385), .Z(n379) );
  XNOR U514 ( .A(sreg[64]), .B(n379), .Z(c[64]) );
  AND U515 ( .A(b[0]), .B(a[3]), .Z(n391) );
  NAND U516 ( .A(b[1]), .B(a[2]), .Z(n393) );
  XNOR U517 ( .A(n392), .B(n393), .Z(n382) );
  NAND U518 ( .A(n392), .B(n380), .Z(n381) );
  NAND U519 ( .A(n382), .B(n381), .Z(n383) );
  XOR U520 ( .A(n391), .B(n383), .Z(n396) );
  NAND U521 ( .A(n384), .B(n385), .Z(n389) );
  ANDN U522 ( .B(n386), .A(n385), .Z(n387) );
  NANDN U523 ( .A(n387), .B(sreg[64]), .Z(n388) );
  AND U524 ( .A(n389), .B(n388), .Z(n397) );
  XNOR U525 ( .A(n397), .B(sreg[65]), .Z(n390) );
  XNOR U526 ( .A(n396), .B(n390), .Z(c[65]) );
  NAND U527 ( .A(b[0]), .B(a[4]), .Z(n400) );
  AND U528 ( .A(b[1]), .B(a[3]), .Z(n399) );
  XNOR U529 ( .A(n401), .B(n399), .Z(n395) );
  XNOR U530 ( .A(n400), .B(n395), .Z(n403) );
  XNOR U531 ( .A(n404), .B(sreg[66]), .Z(n398) );
  XNOR U532 ( .A(n403), .B(n398), .Z(c[66]) );
  NAND U533 ( .A(b[0]), .B(a[5]), .Z(n407) );
  AND U534 ( .A(b[1]), .B(a[4]), .Z(n406) );
  XNOR U535 ( .A(n408), .B(n406), .Z(n402) );
  XNOR U536 ( .A(n407), .B(n402), .Z(n410) );
  XNOR U537 ( .A(n411), .B(sreg[67]), .Z(n405) );
  XNOR U538 ( .A(n410), .B(n405), .Z(c[67]) );
  NAND U539 ( .A(b[0]), .B(a[6]), .Z(n414) );
  AND U540 ( .A(b[1]), .B(a[5]), .Z(n413) );
  XNOR U541 ( .A(n415), .B(n413), .Z(n409) );
  XNOR U542 ( .A(n414), .B(n409), .Z(n417) );
  XNOR U543 ( .A(n418), .B(sreg[68]), .Z(n412) );
  XNOR U544 ( .A(n417), .B(n412), .Z(c[68]) );
  NAND U545 ( .A(b[0]), .B(a[7]), .Z(n421) );
  AND U546 ( .A(b[1]), .B(a[6]), .Z(n420) );
  XNOR U547 ( .A(n422), .B(n420), .Z(n416) );
  XNOR U548 ( .A(n421), .B(n416), .Z(n424) );
  XNOR U549 ( .A(n425), .B(sreg[69]), .Z(n419) );
  XNOR U550 ( .A(n424), .B(n419), .Z(c[69]) );
  NAND U551 ( .A(b[0]), .B(a[8]), .Z(n428) );
  AND U552 ( .A(b[1]), .B(a[7]), .Z(n427) );
  XNOR U553 ( .A(n429), .B(n427), .Z(n423) );
  XNOR U554 ( .A(n428), .B(n423), .Z(n431) );
  XNOR U555 ( .A(n432), .B(sreg[70]), .Z(n426) );
  XNOR U556 ( .A(n431), .B(n426), .Z(c[70]) );
  NAND U557 ( .A(b[0]), .B(a[9]), .Z(n435) );
  AND U558 ( .A(b[1]), .B(a[8]), .Z(n434) );
  XNOR U559 ( .A(n436), .B(n434), .Z(n430) );
  XNOR U560 ( .A(n435), .B(n430), .Z(n438) );
  XNOR U561 ( .A(n439), .B(sreg[71]), .Z(n433) );
  XNOR U562 ( .A(n438), .B(n433), .Z(c[71]) );
  NAND U563 ( .A(b[0]), .B(a[10]), .Z(n442) );
  AND U564 ( .A(b[1]), .B(a[9]), .Z(n441) );
  XNOR U565 ( .A(n443), .B(n441), .Z(n437) );
  XNOR U566 ( .A(n442), .B(n437), .Z(n445) );
  XNOR U567 ( .A(n446), .B(sreg[72]), .Z(n440) );
  XNOR U568 ( .A(n445), .B(n440), .Z(c[72]) );
  NAND U569 ( .A(b[0]), .B(a[11]), .Z(n449) );
  AND U570 ( .A(b[1]), .B(a[10]), .Z(n448) );
  XNOR U571 ( .A(n450), .B(n448), .Z(n444) );
  XNOR U572 ( .A(n449), .B(n444), .Z(n452) );
  XNOR U573 ( .A(n453), .B(sreg[73]), .Z(n447) );
  XNOR U574 ( .A(n452), .B(n447), .Z(c[73]) );
  NAND U575 ( .A(b[0]), .B(a[12]), .Z(n456) );
  AND U576 ( .A(b[1]), .B(a[11]), .Z(n455) );
  XNOR U577 ( .A(n457), .B(n455), .Z(n451) );
  XNOR U578 ( .A(n456), .B(n451), .Z(n459) );
  XNOR U579 ( .A(n460), .B(sreg[74]), .Z(n454) );
  XNOR U580 ( .A(n459), .B(n454), .Z(c[74]) );
  NAND U581 ( .A(b[0]), .B(a[13]), .Z(n463) );
  AND U582 ( .A(b[1]), .B(a[12]), .Z(n462) );
  XNOR U583 ( .A(n464), .B(n462), .Z(n458) );
  XNOR U584 ( .A(n463), .B(n458), .Z(n466) );
  XNOR U585 ( .A(n467), .B(sreg[75]), .Z(n461) );
  XNOR U586 ( .A(n466), .B(n461), .Z(c[75]) );
  NAND U587 ( .A(b[0]), .B(a[14]), .Z(n470) );
  AND U588 ( .A(b[1]), .B(a[13]), .Z(n469) );
  XNOR U589 ( .A(n471), .B(n469), .Z(n465) );
  XNOR U590 ( .A(n470), .B(n465), .Z(n473) );
  XNOR U591 ( .A(n474), .B(sreg[76]), .Z(n468) );
  XNOR U592 ( .A(n473), .B(n468), .Z(c[76]) );
  NAND U593 ( .A(b[0]), .B(a[15]), .Z(n477) );
  AND U594 ( .A(b[1]), .B(a[14]), .Z(n476) );
  XNOR U595 ( .A(n478), .B(n476), .Z(n472) );
  XNOR U596 ( .A(n477), .B(n472), .Z(n480) );
  XNOR U597 ( .A(n481), .B(sreg[77]), .Z(n475) );
  XNOR U598 ( .A(n480), .B(n475), .Z(c[77]) );
  NAND U599 ( .A(b[0]), .B(a[16]), .Z(n484) );
  AND U600 ( .A(b[1]), .B(a[15]), .Z(n483) );
  XNOR U601 ( .A(n485), .B(n483), .Z(n479) );
  XNOR U602 ( .A(n484), .B(n479), .Z(n487) );
  XNOR U603 ( .A(n488), .B(sreg[78]), .Z(n482) );
  XNOR U604 ( .A(n487), .B(n482), .Z(c[78]) );
  NAND U605 ( .A(b[0]), .B(a[17]), .Z(n491) );
  AND U606 ( .A(b[1]), .B(a[16]), .Z(n490) );
  XNOR U607 ( .A(n492), .B(n490), .Z(n486) );
  XNOR U608 ( .A(n491), .B(n486), .Z(n494) );
  XNOR U609 ( .A(n495), .B(sreg[79]), .Z(n489) );
  XNOR U610 ( .A(n494), .B(n489), .Z(c[79]) );
  NAND U611 ( .A(b[0]), .B(a[18]), .Z(n498) );
  AND U612 ( .A(b[1]), .B(a[17]), .Z(n497) );
  XNOR U613 ( .A(n499), .B(n497), .Z(n493) );
  XNOR U614 ( .A(n498), .B(n493), .Z(n501) );
  XNOR U615 ( .A(n502), .B(sreg[80]), .Z(n496) );
  XNOR U616 ( .A(n501), .B(n496), .Z(c[80]) );
  NAND U617 ( .A(b[0]), .B(a[19]), .Z(n505) );
  AND U618 ( .A(b[1]), .B(a[18]), .Z(n504) );
  XNOR U619 ( .A(n506), .B(n504), .Z(n500) );
  XNOR U620 ( .A(n505), .B(n500), .Z(n508) );
  XNOR U621 ( .A(n509), .B(sreg[81]), .Z(n503) );
  XNOR U622 ( .A(n508), .B(n503), .Z(c[81]) );
  NAND U623 ( .A(b[0]), .B(a[20]), .Z(n512) );
  AND U624 ( .A(b[1]), .B(a[19]), .Z(n511) );
  XNOR U625 ( .A(n513), .B(n511), .Z(n507) );
  XNOR U626 ( .A(n512), .B(n507), .Z(n515) );
  XNOR U627 ( .A(n516), .B(sreg[82]), .Z(n510) );
  XNOR U628 ( .A(n515), .B(n510), .Z(c[82]) );
  NAND U629 ( .A(b[0]), .B(a[21]), .Z(n519) );
  AND U630 ( .A(b[1]), .B(a[20]), .Z(n518) );
  XNOR U631 ( .A(n520), .B(n518), .Z(n514) );
  XNOR U632 ( .A(n519), .B(n514), .Z(n522) );
  XNOR U633 ( .A(n523), .B(sreg[83]), .Z(n517) );
  XNOR U634 ( .A(n522), .B(n517), .Z(c[83]) );
  NAND U635 ( .A(b[0]), .B(a[22]), .Z(n526) );
  AND U636 ( .A(b[1]), .B(a[21]), .Z(n525) );
  XNOR U637 ( .A(n527), .B(n525), .Z(n521) );
  XNOR U638 ( .A(n526), .B(n521), .Z(n529) );
  XNOR U639 ( .A(n530), .B(sreg[84]), .Z(n524) );
  XNOR U640 ( .A(n529), .B(n524), .Z(c[84]) );
  NAND U641 ( .A(b[0]), .B(a[23]), .Z(n533) );
  AND U642 ( .A(b[1]), .B(a[22]), .Z(n532) );
  XNOR U643 ( .A(n534), .B(n532), .Z(n528) );
  XNOR U644 ( .A(n533), .B(n528), .Z(n536) );
  XNOR U645 ( .A(n537), .B(sreg[85]), .Z(n531) );
  XNOR U646 ( .A(n536), .B(n531), .Z(c[85]) );
  NAND U647 ( .A(b[0]), .B(a[24]), .Z(n540) );
  AND U648 ( .A(b[1]), .B(a[23]), .Z(n539) );
  XNOR U649 ( .A(n541), .B(n539), .Z(n535) );
  XNOR U650 ( .A(n540), .B(n535), .Z(n543) );
  XNOR U651 ( .A(n544), .B(sreg[86]), .Z(n538) );
  XNOR U652 ( .A(n543), .B(n538), .Z(c[86]) );
  NAND U653 ( .A(b[0]), .B(a[25]), .Z(n547) );
  AND U654 ( .A(b[1]), .B(a[24]), .Z(n546) );
  XNOR U655 ( .A(n548), .B(n546), .Z(n542) );
  XNOR U656 ( .A(n547), .B(n542), .Z(n550) );
  XNOR U657 ( .A(n551), .B(sreg[87]), .Z(n545) );
  XNOR U658 ( .A(n550), .B(n545), .Z(c[87]) );
  NAND U659 ( .A(b[0]), .B(a[26]), .Z(n554) );
  AND U660 ( .A(b[1]), .B(a[25]), .Z(n553) );
  XNOR U661 ( .A(n555), .B(n553), .Z(n549) );
  XNOR U662 ( .A(n554), .B(n549), .Z(n557) );
  XNOR U663 ( .A(n558), .B(sreg[88]), .Z(n552) );
  XNOR U664 ( .A(n557), .B(n552), .Z(c[88]) );
  NAND U665 ( .A(b[0]), .B(a[27]), .Z(n561) );
  AND U666 ( .A(b[1]), .B(a[26]), .Z(n560) );
  XNOR U667 ( .A(n562), .B(n560), .Z(n556) );
  XNOR U668 ( .A(n561), .B(n556), .Z(n564) );
  XNOR U669 ( .A(n565), .B(sreg[89]), .Z(n559) );
  XNOR U670 ( .A(n564), .B(n559), .Z(c[89]) );
  NAND U671 ( .A(b[0]), .B(a[28]), .Z(n570) );
  AND U672 ( .A(b[1]), .B(a[27]), .Z(n569) );
  XNOR U673 ( .A(n571), .B(n569), .Z(n563) );
  XNOR U674 ( .A(n570), .B(n563), .Z(n567) );
  XNOR U675 ( .A(n568), .B(sreg[90]), .Z(n566) );
  XNOR U676 ( .A(n567), .B(n566), .Z(c[90]) );
  NAND U677 ( .A(b[0]), .B(a[29]), .Z(n575) );
  AND U678 ( .A(b[1]), .B(a[28]), .Z(n574) );
  XNOR U679 ( .A(n576), .B(n574), .Z(n572) );
  XOR U680 ( .A(n575), .B(n572), .Z(n579) );
  XNOR U681 ( .A(n579), .B(sreg[91]), .Z(n573) );
  XOR U682 ( .A(n578), .B(n573), .Z(c[91]) );
  NAND U683 ( .A(b[0]), .B(a[30]), .Z(n582) );
  AND U684 ( .A(b[1]), .B(a[29]), .Z(n581) );
  XNOR U685 ( .A(n583), .B(n581), .Z(n577) );
  XNOR U686 ( .A(n582), .B(n577), .Z(n585) );
  XNOR U687 ( .A(n586), .B(sreg[92]), .Z(n580) );
  XNOR U688 ( .A(n585), .B(n580), .Z(c[92]) );
  NAND U689 ( .A(b[0]), .B(a[31]), .Z(n589) );
  AND U690 ( .A(b[1]), .B(a[30]), .Z(n588) );
  XNOR U691 ( .A(n590), .B(n588), .Z(n584) );
  XNOR U692 ( .A(n589), .B(n584), .Z(n592) );
  XNOR U693 ( .A(n593), .B(sreg[93]), .Z(n587) );
  XNOR U694 ( .A(n592), .B(n587), .Z(c[93]) );
  NAND U695 ( .A(b[0]), .B(a[32]), .Z(n596) );
  AND U696 ( .A(b[1]), .B(a[31]), .Z(n595) );
  XNOR U697 ( .A(n597), .B(n595), .Z(n591) );
  XNOR U698 ( .A(n596), .B(n591), .Z(n599) );
  XNOR U699 ( .A(n600), .B(sreg[94]), .Z(n594) );
  XNOR U700 ( .A(n599), .B(n594), .Z(c[94]) );
  NAND U701 ( .A(b[0]), .B(a[33]), .Z(n603) );
  AND U702 ( .A(b[1]), .B(a[32]), .Z(n602) );
  XNOR U703 ( .A(n604), .B(n602), .Z(n598) );
  XNOR U704 ( .A(n603), .B(n598), .Z(n606) );
  XNOR U705 ( .A(n607), .B(sreg[95]), .Z(n601) );
  XNOR U706 ( .A(n606), .B(n601), .Z(c[95]) );
  NAND U707 ( .A(b[0]), .B(a[34]), .Z(n610) );
  AND U708 ( .A(b[1]), .B(a[33]), .Z(n609) );
  XNOR U709 ( .A(n611), .B(n609), .Z(n605) );
  XNOR U710 ( .A(n610), .B(n605), .Z(n613) );
  XNOR U711 ( .A(n614), .B(sreg[96]), .Z(n608) );
  XNOR U712 ( .A(n613), .B(n608), .Z(c[96]) );
  NAND U713 ( .A(b[0]), .B(a[35]), .Z(n617) );
  AND U714 ( .A(b[1]), .B(a[34]), .Z(n616) );
  XNOR U715 ( .A(n618), .B(n616), .Z(n612) );
  XNOR U716 ( .A(n617), .B(n612), .Z(n620) );
  XNOR U717 ( .A(n621), .B(sreg[97]), .Z(n615) );
  XNOR U718 ( .A(n620), .B(n615), .Z(c[97]) );
  NAND U719 ( .A(b[0]), .B(a[36]), .Z(n624) );
  AND U720 ( .A(b[1]), .B(a[35]), .Z(n623) );
  XNOR U721 ( .A(n625), .B(n623), .Z(n619) );
  XNOR U722 ( .A(n624), .B(n619), .Z(n627) );
  XNOR U723 ( .A(n628), .B(sreg[98]), .Z(n622) );
  XNOR U724 ( .A(n627), .B(n622), .Z(c[98]) );
  NAND U725 ( .A(b[0]), .B(a[37]), .Z(n631) );
  AND U726 ( .A(b[1]), .B(a[36]), .Z(n630) );
  XNOR U727 ( .A(n632), .B(n630), .Z(n626) );
  XNOR U728 ( .A(n631), .B(n626), .Z(n634) );
  XNOR U729 ( .A(n635), .B(sreg[99]), .Z(n629) );
  XNOR U730 ( .A(n634), .B(n629), .Z(c[99]) );
  NAND U731 ( .A(b[0]), .B(a[38]), .Z(n638) );
  AND U732 ( .A(b[1]), .B(a[37]), .Z(n637) );
  XNOR U733 ( .A(n639), .B(n637), .Z(n633) );
  XNOR U734 ( .A(n638), .B(n633), .Z(n641) );
  XNOR U735 ( .A(n642), .B(sreg[100]), .Z(n636) );
  XNOR U736 ( .A(n641), .B(n636), .Z(c[100]) );
  NAND U737 ( .A(b[0]), .B(a[39]), .Z(n645) );
  AND U738 ( .A(b[1]), .B(a[38]), .Z(n644) );
  XNOR U739 ( .A(n646), .B(n644), .Z(n640) );
  XNOR U740 ( .A(n645), .B(n640), .Z(n648) );
  XNOR U741 ( .A(n649), .B(sreg[101]), .Z(n643) );
  XNOR U742 ( .A(n648), .B(n643), .Z(c[101]) );
  NAND U743 ( .A(b[0]), .B(a[40]), .Z(n652) );
  AND U744 ( .A(b[1]), .B(a[39]), .Z(n651) );
  XNOR U745 ( .A(n653), .B(n651), .Z(n647) );
  XNOR U746 ( .A(n652), .B(n647), .Z(n655) );
  XNOR U747 ( .A(n656), .B(sreg[102]), .Z(n650) );
  XNOR U748 ( .A(n655), .B(n650), .Z(c[102]) );
  NAND U749 ( .A(b[0]), .B(a[41]), .Z(n659) );
  AND U750 ( .A(b[1]), .B(a[40]), .Z(n658) );
  XNOR U751 ( .A(n660), .B(n658), .Z(n654) );
  XNOR U752 ( .A(n659), .B(n654), .Z(n662) );
  XNOR U753 ( .A(n663), .B(sreg[103]), .Z(n657) );
  XNOR U754 ( .A(n662), .B(n657), .Z(c[103]) );
  NAND U755 ( .A(b[0]), .B(a[42]), .Z(n666) );
  AND U756 ( .A(b[1]), .B(a[41]), .Z(n665) );
  XNOR U757 ( .A(n667), .B(n665), .Z(n661) );
  XNOR U758 ( .A(n666), .B(n661), .Z(n669) );
  XNOR U759 ( .A(n670), .B(sreg[104]), .Z(n664) );
  XNOR U760 ( .A(n669), .B(n664), .Z(c[104]) );
  NAND U761 ( .A(b[0]), .B(a[43]), .Z(n673) );
  AND U762 ( .A(b[1]), .B(a[42]), .Z(n672) );
  XNOR U763 ( .A(n674), .B(n672), .Z(n668) );
  XNOR U764 ( .A(n673), .B(n668), .Z(n676) );
  XNOR U765 ( .A(n677), .B(sreg[105]), .Z(n671) );
  XNOR U766 ( .A(n676), .B(n671), .Z(c[105]) );
  NAND U767 ( .A(b[0]), .B(a[44]), .Z(n680) );
  AND U768 ( .A(b[1]), .B(a[43]), .Z(n679) );
  XNOR U769 ( .A(n681), .B(n679), .Z(n675) );
  XNOR U770 ( .A(n680), .B(n675), .Z(n683) );
  XNOR U771 ( .A(n684), .B(sreg[106]), .Z(n678) );
  XNOR U772 ( .A(n683), .B(n678), .Z(c[106]) );
  NAND U773 ( .A(b[0]), .B(a[45]), .Z(n687) );
  AND U774 ( .A(b[1]), .B(a[44]), .Z(n686) );
  XNOR U775 ( .A(n688), .B(n686), .Z(n682) );
  XNOR U776 ( .A(n687), .B(n682), .Z(n690) );
  XNOR U777 ( .A(n691), .B(sreg[107]), .Z(n685) );
  XNOR U778 ( .A(n690), .B(n685), .Z(c[107]) );
  NAND U779 ( .A(b[0]), .B(a[46]), .Z(n694) );
  AND U780 ( .A(b[1]), .B(a[45]), .Z(n693) );
  XNOR U781 ( .A(n695), .B(n693), .Z(n689) );
  XNOR U782 ( .A(n694), .B(n689), .Z(n697) );
  XNOR U783 ( .A(n698), .B(sreg[108]), .Z(n692) );
  XNOR U784 ( .A(n697), .B(n692), .Z(c[108]) );
  NAND U785 ( .A(b[0]), .B(a[47]), .Z(n701) );
  AND U786 ( .A(b[1]), .B(a[46]), .Z(n700) );
  XNOR U787 ( .A(n702), .B(n700), .Z(n696) );
  XNOR U788 ( .A(n701), .B(n696), .Z(n704) );
  XNOR U789 ( .A(n705), .B(sreg[109]), .Z(n699) );
  XNOR U790 ( .A(n704), .B(n699), .Z(c[109]) );
  NAND U791 ( .A(b[0]), .B(a[48]), .Z(n708) );
  AND U792 ( .A(b[1]), .B(a[47]), .Z(n707) );
  XNOR U793 ( .A(n709), .B(n707), .Z(n703) );
  XNOR U794 ( .A(n708), .B(n703), .Z(n711) );
  XNOR U795 ( .A(n712), .B(sreg[110]), .Z(n706) );
  XNOR U796 ( .A(n711), .B(n706), .Z(c[110]) );
  NAND U797 ( .A(b[0]), .B(a[49]), .Z(n715) );
  AND U798 ( .A(b[1]), .B(a[48]), .Z(n714) );
  XNOR U799 ( .A(n716), .B(n714), .Z(n710) );
  XNOR U800 ( .A(n715), .B(n710), .Z(n718) );
  XNOR U801 ( .A(n719), .B(sreg[111]), .Z(n713) );
  XNOR U802 ( .A(n718), .B(n713), .Z(c[111]) );
  NAND U803 ( .A(b[0]), .B(a[50]), .Z(n722) );
  AND U804 ( .A(b[1]), .B(a[49]), .Z(n721) );
  XNOR U805 ( .A(n723), .B(n721), .Z(n717) );
  XNOR U806 ( .A(n722), .B(n717), .Z(n725) );
  XNOR U807 ( .A(n726), .B(sreg[112]), .Z(n720) );
  XNOR U808 ( .A(n725), .B(n720), .Z(c[112]) );
  NAND U809 ( .A(b[0]), .B(a[51]), .Z(n729) );
  AND U810 ( .A(b[1]), .B(a[50]), .Z(n728) );
  XNOR U811 ( .A(n730), .B(n728), .Z(n724) );
  XNOR U812 ( .A(n729), .B(n724), .Z(n732) );
  XNOR U813 ( .A(n733), .B(sreg[113]), .Z(n727) );
  XNOR U814 ( .A(n732), .B(n727), .Z(c[113]) );
  NAND U815 ( .A(b[0]), .B(a[52]), .Z(n736) );
  AND U816 ( .A(b[1]), .B(a[51]), .Z(n735) );
  XNOR U817 ( .A(n737), .B(n735), .Z(n731) );
  XNOR U818 ( .A(n736), .B(n731), .Z(n739) );
  XNOR U819 ( .A(n740), .B(sreg[114]), .Z(n734) );
  XNOR U820 ( .A(n739), .B(n734), .Z(c[114]) );
  NAND U821 ( .A(b[0]), .B(a[53]), .Z(n743) );
  AND U822 ( .A(b[1]), .B(a[52]), .Z(n742) );
  XNOR U823 ( .A(n744), .B(n742), .Z(n738) );
  XNOR U824 ( .A(n743), .B(n738), .Z(n746) );
  XNOR U825 ( .A(n747), .B(sreg[115]), .Z(n741) );
  XNOR U826 ( .A(n746), .B(n741), .Z(c[115]) );
  NAND U827 ( .A(b[0]), .B(a[54]), .Z(n750) );
  AND U828 ( .A(b[1]), .B(a[53]), .Z(n749) );
  XNOR U829 ( .A(n751), .B(n749), .Z(n745) );
  XNOR U830 ( .A(n750), .B(n745), .Z(n753) );
  XNOR U831 ( .A(n754), .B(sreg[116]), .Z(n748) );
  XNOR U832 ( .A(n753), .B(n748), .Z(c[116]) );
  NAND U833 ( .A(b[0]), .B(a[55]), .Z(n757) );
  AND U834 ( .A(b[1]), .B(a[54]), .Z(n756) );
  XNOR U835 ( .A(n758), .B(n756), .Z(n752) );
  XNOR U836 ( .A(n757), .B(n752), .Z(n760) );
  XNOR U837 ( .A(n761), .B(sreg[117]), .Z(n755) );
  XNOR U838 ( .A(n760), .B(n755), .Z(c[117]) );
  NAND U839 ( .A(b[0]), .B(a[56]), .Z(n764) );
  AND U840 ( .A(b[1]), .B(a[55]), .Z(n763) );
  XNOR U841 ( .A(n765), .B(n763), .Z(n759) );
  XNOR U842 ( .A(n764), .B(n759), .Z(n767) );
  XNOR U843 ( .A(n768), .B(sreg[118]), .Z(n762) );
  XNOR U844 ( .A(n767), .B(n762), .Z(c[118]) );
  NAND U845 ( .A(b[0]), .B(a[57]), .Z(n771) );
  AND U846 ( .A(b[1]), .B(a[56]), .Z(n770) );
  XNOR U847 ( .A(n772), .B(n770), .Z(n766) );
  XNOR U848 ( .A(n771), .B(n766), .Z(n774) );
  XNOR U849 ( .A(n775), .B(sreg[119]), .Z(n769) );
  XNOR U850 ( .A(n774), .B(n769), .Z(c[119]) );
  NAND U851 ( .A(b[0]), .B(a[58]), .Z(n778) );
  AND U852 ( .A(b[1]), .B(a[57]), .Z(n777) );
  XNOR U853 ( .A(n779), .B(n777), .Z(n773) );
  XNOR U854 ( .A(n778), .B(n773), .Z(n781) );
  XNOR U855 ( .A(n782), .B(sreg[120]), .Z(n776) );
  XNOR U856 ( .A(n781), .B(n776), .Z(c[120]) );
  NAND U857 ( .A(b[0]), .B(a[59]), .Z(n785) );
  AND U858 ( .A(b[1]), .B(a[58]), .Z(n784) );
  XNOR U859 ( .A(n786), .B(n784), .Z(n780) );
  XNOR U860 ( .A(n785), .B(n780), .Z(n788) );
  XNOR U861 ( .A(n789), .B(sreg[121]), .Z(n783) );
  XNOR U862 ( .A(n788), .B(n783), .Z(c[121]) );
  NAND U863 ( .A(b[0]), .B(a[60]), .Z(n792) );
  AND U864 ( .A(b[1]), .B(a[59]), .Z(n791) );
  XNOR U865 ( .A(n793), .B(n791), .Z(n787) );
  XNOR U866 ( .A(n792), .B(n787), .Z(n795) );
  XNOR U867 ( .A(n796), .B(sreg[122]), .Z(n790) );
  XNOR U868 ( .A(n795), .B(n790), .Z(c[122]) );
  NAND U869 ( .A(b[0]), .B(a[61]), .Z(n799) );
  AND U870 ( .A(b[1]), .B(a[60]), .Z(n798) );
  XNOR U871 ( .A(n800), .B(n798), .Z(n794) );
  XNOR U872 ( .A(n799), .B(n794), .Z(n802) );
  XNOR U873 ( .A(n803), .B(sreg[123]), .Z(n797) );
  XNOR U874 ( .A(n802), .B(n797), .Z(c[123]) );
  NAND U875 ( .A(a[62]), .B(b[0]), .Z(n806) );
  AND U876 ( .A(b[1]), .B(a[61]), .Z(n805) );
  XNOR U877 ( .A(n807), .B(n805), .Z(n801) );
  XNOR U878 ( .A(n806), .B(n801), .Z(n808) );
  XNOR U879 ( .A(n809), .B(sreg[124]), .Z(n804) );
  XNOR U880 ( .A(n808), .B(n804), .Z(c[124]) );
  AND U881 ( .A(b[1]), .B(a[62]), .Z(n813) );
  NAND U882 ( .A(b[0]), .B(a[63]), .Z(n814) );
  XNOR U883 ( .A(n813), .B(n814), .Z(n816) );
  XNOR U884 ( .A(n816), .B(n815), .Z(n811) );
  XNOR U885 ( .A(n812), .B(sreg[125]), .Z(n810) );
  XNOR U886 ( .A(n811), .B(n810), .Z(c[125]) );
  NANDN U887 ( .A(n814), .B(n813), .Z(n818) );
  NAND U888 ( .A(n816), .B(n815), .Z(n817) );
  AND U889 ( .A(n818), .B(n817), .Z(n822) );
  AND U890 ( .A(b[1]), .B(a[63]), .Z(n820) );
  XNOR U891 ( .A(n822), .B(n820), .Z(n819) );
  XNOR U892 ( .A(n821), .B(n819), .Z(c[126]) );
endmodule

