
module compare_N16384_CC8 ( clk, rst, x, y, g, e );
  input [2047:0] x;
  input [2047:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  NANDN U10 ( .A(n4419), .B(n4418), .Z(n8) );
  ANDN U11 ( .B(n8), .A(n5511), .Z(n9) );
  ANDN U12 ( .B(n8994), .A(n5507), .Z(n10) );
  NAND U13 ( .A(n5509), .B(n9), .Z(n11) );
  AND U14 ( .A(n10), .B(n11), .Z(n12) );
  ANDN U15 ( .B(n5510), .A(n12), .Z(n13) );
  NAND U16 ( .A(n12237), .B(n13), .Z(n14) );
  AND U17 ( .A(n5508), .B(n14), .Z(n15) );
  NAND U18 ( .A(n8995), .B(n15), .Z(n16) );
  NAND U19 ( .A(n12241), .B(n16), .Z(n17) );
  ANDN U20 ( .B(n17), .A(n12242), .Z(n18) );
  NANDN U21 ( .A(n18), .B(n12244), .Z(n19) );
  NAND U22 ( .A(n12247), .B(n19), .Z(n20) );
  NAND U23 ( .A(n12249), .B(n20), .Z(n4421) );
  AND U24 ( .A(n9121), .B(n12480), .Z(n21) );
  NANDN U25 ( .A(n4440), .B(n4439), .Z(n22) );
  AND U26 ( .A(n21), .B(n22), .Z(n23) );
  AND U27 ( .A(n5427), .B(n12485), .Z(n24) );
  OR U28 ( .A(n12483), .B(n23), .Z(n25) );
  AND U29 ( .A(n24), .B(n25), .Z(n26) );
  NOR U30 ( .A(n26), .B(n9125), .Z(n27) );
  NAND U31 ( .A(n12491), .B(n27), .Z(n28) );
  AND U32 ( .A(n5428), .B(n28), .Z(n29) );
  NAND U33 ( .A(n29), .B(n12493), .Z(n30) );
  NANDN U34 ( .A(n12495), .B(n30), .Z(n31) );
  AND U35 ( .A(n12497), .B(n31), .Z(n32) );
  OR U36 ( .A(n12499), .B(n32), .Z(n33) );
  NAND U37 ( .A(n12501), .B(n33), .Z(n34) );
  NANDN U38 ( .A(n12503), .B(n34), .Z(n35) );
  ANDN U39 ( .B(n35), .A(n12504), .Z(n4441) );
  NAND U40 ( .A(n5318), .B(n5322), .Z(n36) );
  ANDN U41 ( .B(n36), .A(n4478), .Z(n37) );
  NAND U42 ( .A(n4477), .B(n4476), .Z(n38) );
  AND U43 ( .A(n5329), .B(n38), .Z(n39) );
  NAND U44 ( .A(n39), .B(n5325), .Z(n40) );
  NOR U45 ( .A(n5327), .B(n12901), .Z(n41) );
  NAND U46 ( .A(n40), .B(n41), .Z(n42) );
  NAND U47 ( .A(n12903), .B(n42), .Z(n43) );
  OR U48 ( .A(n43), .B(n5324), .Z(n44) );
  NAND U49 ( .A(n12905), .B(n44), .Z(n45) );
  NANDN U50 ( .A(n12907), .B(n45), .Z(n46) );
  NANDN U51 ( .A(n12908), .B(n46), .Z(n47) );
  NAND U52 ( .A(n12910), .B(n47), .Z(n48) );
  AND U53 ( .A(n5317), .B(n48), .Z(n49) );
  NANDN U54 ( .A(n12913), .B(n49), .Z(n50) );
  NAND U55 ( .A(n12915), .B(n50), .Z(n51) );
  ANDN U56 ( .B(n51), .A(n37), .Z(n4480) );
  AND U57 ( .A(n5280), .B(n13010), .Z(n52) );
  NAND U58 ( .A(n4495), .B(n52), .Z(n53) );
  NANDN U59 ( .A(n5279), .B(n53), .Z(n54) );
  AND U60 ( .A(n5281), .B(n5276), .Z(n55) );
  OR U61 ( .A(n54), .B(n5283), .Z(n56) );
  AND U62 ( .A(n55), .B(n56), .Z(n57) );
  NOR U63 ( .A(n5274), .B(n57), .Z(n58) );
  NAND U64 ( .A(n5278), .B(n58), .Z(n59) );
  AND U65 ( .A(n13027), .B(n59), .Z(n60) );
  NAND U66 ( .A(n60), .B(n5277), .Z(n61) );
  AND U67 ( .A(n13028), .B(n61), .Z(n62) );
  NAND U68 ( .A(n62), .B(n5275), .Z(n63) );
  ANDN U69 ( .B(n5272), .A(n5273), .Z(n64) );
  NANDN U70 ( .A(n13031), .B(n63), .Z(n65) );
  NAND U71 ( .A(n64), .B(n65), .Z(n4496) );
  NANDN U72 ( .A(n4509), .B(n13207), .Z(n66) );
  NAND U73 ( .A(n13209), .B(n66), .Z(n67) );
  AND U74 ( .A(n13211), .B(n67), .Z(n68) );
  ANDN U75 ( .B(n9386), .A(n5222), .Z(n69) );
  NANDN U76 ( .A(n68), .B(n13213), .Z(n70) );
  AND U77 ( .A(n69), .B(n70), .Z(n71) );
  NOR U78 ( .A(n5224), .B(n71), .Z(n72) );
  NAND U79 ( .A(n9388), .B(n72), .Z(n73) );
  AND U80 ( .A(n5223), .B(n73), .Z(n74) );
  NANDN U81 ( .A(n74), .B(n9389), .Z(n75) );
  NANDN U82 ( .A(n13223), .B(n75), .Z(n76) );
  NAND U83 ( .A(n13225), .B(n76), .Z(n77) );
  NANDN U84 ( .A(n13227), .B(n77), .Z(n78) );
  NAND U85 ( .A(n13229), .B(n78), .Z(n79) );
  ANDN U86 ( .B(n79), .A(n13230), .Z(n80) );
  OR U87 ( .A(n13232), .B(n80), .Z(n81) );
  ANDN U88 ( .B(n81), .A(n13234), .Z(n4510) );
  NAND U89 ( .A(n13409), .B(n4525), .Z(n82) );
  NAND U90 ( .A(n13410), .B(n82), .Z(n83) );
  ANDN U91 ( .B(n83), .A(n13413), .Z(n84) );
  OR U92 ( .A(n13414), .B(n84), .Z(n85) );
  NAND U93 ( .A(n13416), .B(n85), .Z(n86) );
  NAND U94 ( .A(n13419), .B(n86), .Z(n87) );
  NANDN U95 ( .A(n13421), .B(n87), .Z(n88) );
  NAND U96 ( .A(n13423), .B(n88), .Z(n89) );
  ANDN U97 ( .B(n89), .A(n13425), .Z(n90) );
  AND U98 ( .A(n13428), .B(n5158), .Z(n91) );
  OR U99 ( .A(n13426), .B(n90), .Z(n92) );
  AND U100 ( .A(n91), .B(n92), .Z(n93) );
  NOR U101 ( .A(n13435), .B(n13431), .Z(n94) );
  NANDN U102 ( .A(n93), .B(n94), .Z(n95) );
  AND U103 ( .A(n5157), .B(n95), .Z(n96) );
  NANDN U104 ( .A(n13437), .B(n96), .Z(n4526) );
  NANDN U105 ( .A(n13483), .B(n4560), .Z(n97) );
  NAND U106 ( .A(n13485), .B(n97), .Z(n98) );
  ANDN U107 ( .B(n98), .A(n13487), .Z(n99) );
  NANDN U108 ( .A(n99), .B(n13489), .Z(n100) );
  NANDN U109 ( .A(n13491), .B(n100), .Z(n101) );
  NAND U110 ( .A(n13493), .B(n101), .Z(n102) );
  NOR U111 ( .A(n13495), .B(n5131), .Z(n103) );
  NANDN U112 ( .A(n102), .B(n5133), .Z(n104) );
  AND U113 ( .A(n103), .B(n104), .Z(n105) );
  NOR U114 ( .A(n5134), .B(n105), .Z(n106) );
  NAND U115 ( .A(n5129), .B(n106), .Z(n107) );
  AND U116 ( .A(n13503), .B(n107), .Z(n108) );
  NAND U117 ( .A(n5132), .B(n108), .Z(n109) );
  ANDN U118 ( .B(n109), .A(n5130), .Z(n110) );
  NANDN U119 ( .A(n13505), .B(n110), .Z(n4561) );
  NAND U120 ( .A(n4593), .B(n4592), .Z(n111) );
  AND U121 ( .A(n5076), .B(n111), .Z(n112) );
  NAND U122 ( .A(n112), .B(n9530), .Z(n113) );
  ANDN U123 ( .B(n5074), .A(n13651), .Z(n114) );
  NAND U124 ( .A(n113), .B(n114), .Z(n115) );
  NAND U125 ( .A(n5075), .B(n115), .Z(n116) );
  NOR U126 ( .A(n5073), .B(n5069), .Z(n117) );
  NANDN U127 ( .A(n116), .B(n5071), .Z(n118) );
  AND U128 ( .A(n117), .B(n118), .Z(n119) );
  ANDN U129 ( .B(n5072), .A(n119), .Z(n120) );
  NAND U130 ( .A(n9532), .B(n120), .Z(n121) );
  ANDN U131 ( .B(n121), .A(n13663), .Z(n122) );
  NAND U132 ( .A(n122), .B(n5070), .Z(n123) );
  AND U133 ( .A(n5067), .B(n123), .Z(n124) );
  NAND U134 ( .A(n124), .B(n9531), .Z(n125) );
  NANDN U135 ( .A(n13669), .B(n125), .Z(n4595) );
  OR U136 ( .A(n10157), .B(n10158), .Z(n126) );
  NAND U137 ( .A(n14667), .B(n126), .Z(n127) );
  NANDN U138 ( .A(n10159), .B(n127), .Z(n128) );
  NANDN U139 ( .A(n128), .B(n10160), .Z(n129) );
  AND U140 ( .A(n10161), .B(n129), .Z(n130) );
  ANDN U141 ( .B(n10162), .A(n130), .Z(n131) );
  NANDN U142 ( .A(y[2022]), .B(x[2022]), .Z(n132) );
  NAND U143 ( .A(n131), .B(n132), .Z(n133) );
  NAND U144 ( .A(n14678), .B(n133), .Z(n134) );
  NANDN U145 ( .A(n14681), .B(n134), .Z(n135) );
  AND U146 ( .A(n14683), .B(n135), .Z(n136) );
  OR U147 ( .A(n136), .B(n14685), .Z(n137) );
  NAND U148 ( .A(n14686), .B(n137), .Z(n138) );
  AND U149 ( .A(n14687), .B(n138), .Z(n139) );
  ANDN U150 ( .B(n14689), .A(n14691), .Z(n140) );
  OR U151 ( .A(n139), .B(n14688), .Z(n141) );
  NAND U152 ( .A(n140), .B(n141), .Z(n142) );
  ANDN U153 ( .B(n142), .A(n10165), .Z(n10166) );
  NAND U154 ( .A(n11867), .B(n4385), .Z(n143) );
  ANDN U155 ( .B(n143), .A(n5626), .Z(n144) );
  NANDN U156 ( .A(n11869), .B(n144), .Z(n145) );
  NAND U157 ( .A(n11871), .B(n145), .Z(n146) );
  NANDN U158 ( .A(n5628), .B(n146), .Z(n147) );
  AND U159 ( .A(n11875), .B(n147), .Z(n148) );
  NOR U160 ( .A(n11877), .B(n148), .Z(n149) );
  NAND U161 ( .A(n11878), .B(n149), .Z(n150) );
  AND U162 ( .A(n11881), .B(n150), .Z(n151) );
  ANDN U163 ( .B(n5621), .A(n151), .Z(n152) );
  NAND U164 ( .A(n11883), .B(n152), .Z(n153) );
  AND U165 ( .A(n11884), .B(n153), .Z(n154) );
  NAND U166 ( .A(n5619), .B(n154), .Z(n155) );
  ANDN U167 ( .B(n155), .A(n5622), .Z(n156) );
  NANDN U168 ( .A(n11891), .B(n156), .Z(n157) );
  AND U169 ( .A(n5620), .B(n11893), .Z(n158) );
  NAND U170 ( .A(n157), .B(n158), .Z(n159) );
  NANDN U171 ( .A(n11895), .B(n159), .Z(n4386) );
  AND U172 ( .A(n4392), .B(n4391), .Z(n160) );
  NAND U173 ( .A(n5584), .B(n160), .Z(n161) );
  NAND U174 ( .A(n5582), .B(n161), .Z(n162) );
  NANDN U175 ( .A(n162), .B(n5578), .Z(n163) );
  AND U176 ( .A(n5580), .B(n163), .Z(n164) );
  AND U177 ( .A(n5573), .B(n5577), .Z(n165) );
  NANDN U178 ( .A(n5575), .B(n164), .Z(n166) );
  NAND U179 ( .A(n165), .B(n166), .Z(n167) );
  ANDN U180 ( .B(n5576), .A(n11959), .Z(n168) );
  NAND U181 ( .A(n167), .B(n168), .Z(n169) );
  NAND U182 ( .A(n11961), .B(n169), .Z(n170) );
  NANDN U183 ( .A(n170), .B(n5574), .Z(n171) );
  NANDN U184 ( .A(n11963), .B(n171), .Z(n172) );
  NAND U185 ( .A(n11965), .B(n172), .Z(n173) );
  NAND U186 ( .A(n11967), .B(n173), .Z(n4393) );
  ANDN U187 ( .B(n12177), .A(n8970), .Z(n174) );
  NANDN U188 ( .A(n4414), .B(n12175), .Z(n175) );
  AND U189 ( .A(n174), .B(n175), .Z(n176) );
  NAND U190 ( .A(n4415), .B(n4416), .Z(n177) );
  NANDN U191 ( .A(n176), .B(n177), .Z(n178) );
  ANDN U192 ( .B(n178), .A(n8973), .Z(n179) );
  NANDN U193 ( .A(n179), .B(n12187), .Z(n180) );
  NAND U194 ( .A(n12188), .B(n180), .Z(n181) );
  NAND U195 ( .A(n12191), .B(n181), .Z(n182) );
  NAND U196 ( .A(n12193), .B(n182), .Z(n183) );
  AND U197 ( .A(n5521), .B(n183), .Z(n184) );
  NAND U198 ( .A(n184), .B(n8981), .Z(n185) );
  ANDN U199 ( .B(n8985), .A(n8983), .Z(n186) );
  NAND U200 ( .A(n185), .B(n186), .Z(n187) );
  NAND U201 ( .A(n8987), .B(n187), .Z(n188) );
  OR U202 ( .A(n5520), .B(n188), .Z(n189) );
  AND U203 ( .A(n8984), .B(n189), .Z(n4417) );
  OR U204 ( .A(n12275), .B(n4423), .Z(n190) );
  NAND U205 ( .A(n12277), .B(n190), .Z(n191) );
  NANDN U206 ( .A(n12279), .B(n191), .Z(n192) );
  NAND U207 ( .A(n12281), .B(n192), .Z(n193) );
  AND U208 ( .A(n12283), .B(n193), .Z(n194) );
  NANDN U209 ( .A(n9033), .B(n194), .Z(n195) );
  ANDN U210 ( .B(n12289), .A(n12284), .Z(n196) );
  NAND U211 ( .A(n195), .B(n196), .Z(n197) );
  NANDN U212 ( .A(n9034), .B(n197), .Z(n198) );
  OR U213 ( .A(n198), .B(n12290), .Z(n199) );
  NANDN U214 ( .A(n12293), .B(n199), .Z(n200) );
  NAND U215 ( .A(n12295), .B(n200), .Z(n201) );
  NANDN U216 ( .A(n201), .B(n5500), .Z(n202) );
  ANDN U217 ( .B(n202), .A(n5498), .Z(n203) );
  NAND U218 ( .A(n203), .B(n12296), .Z(n204) );
  AND U219 ( .A(n5496), .B(n204), .Z(n205) );
  NAND U220 ( .A(n205), .B(n5501), .Z(n4424) );
  NAND U221 ( .A(n4428), .B(n12355), .Z(n206) );
  NANDN U222 ( .A(n12356), .B(n206), .Z(n207) );
  AND U223 ( .A(n12358), .B(n207), .Z(n208) );
  NAND U224 ( .A(n5477), .B(n208), .Z(n209) );
  ANDN U225 ( .B(n209), .A(n5474), .Z(n210) );
  NANDN U226 ( .A(n12361), .B(n210), .Z(n211) );
  AND U227 ( .A(n5472), .B(n5476), .Z(n212) );
  NAND U228 ( .A(n211), .B(n212), .Z(n213) );
  NAND U229 ( .A(n5475), .B(n213), .Z(n214) );
  NANDN U230 ( .A(n214), .B(n5470), .Z(n215) );
  ANDN U231 ( .B(n215), .A(n5473), .Z(n216) );
  NAND U232 ( .A(n216), .B(n5468), .Z(n217) );
  AND U233 ( .A(n5471), .B(n217), .Z(n218) );
  NAND U234 ( .A(n218), .B(n12373), .Z(n4431) );
  NAND U235 ( .A(n4441), .B(n5426), .Z(n219) );
  AND U236 ( .A(n12511), .B(n219), .Z(n220) );
  NAND U237 ( .A(n220), .B(n12506), .Z(n221) );
  ANDN U238 ( .B(n5423), .A(n5425), .Z(n222) );
  NAND U239 ( .A(n221), .B(n222), .Z(n223) );
  NAND U240 ( .A(n12515), .B(n223), .Z(n224) );
  AND U241 ( .A(n5422), .B(n5424), .Z(n225) );
  NAND U242 ( .A(n224), .B(n225), .Z(n226) );
  NAND U243 ( .A(n12522), .B(n226), .Z(n227) );
  ANDN U244 ( .B(n5420), .A(n5421), .Z(n228) );
  OR U245 ( .A(n227), .B(n9140), .Z(n229) );
  AND U246 ( .A(n228), .B(n229), .Z(n230) );
  NANDN U247 ( .A(n230), .B(n12527), .Z(n231) );
  ANDN U248 ( .B(n231), .A(n5418), .Z(n4442) );
  ANDN U249 ( .B(n5452), .A(n12396), .Z(n232) );
  ANDN U250 ( .B(n9097), .A(n5453), .Z(n233) );
  NAND U251 ( .A(n12390), .B(n233), .Z(n234) );
  AND U252 ( .A(n232), .B(n234), .Z(n235) );
  NANDN U253 ( .A(n235), .B(n12398), .Z(n236) );
  ANDN U254 ( .B(n236), .A(n12401), .Z(n237) );
  NANDN U255 ( .A(n237), .B(n12403), .Z(n238) );
  NANDN U256 ( .A(n12404), .B(n238), .Z(n239) );
  NAND U257 ( .A(n9098), .B(n239), .Z(n240) );
  NANDN U258 ( .A(n240), .B(n12407), .Z(n241) );
  NAND U259 ( .A(n9099), .B(n241), .Z(n242) );
  NAND U260 ( .A(n9100), .B(n242), .Z(n243) );
  OR U261 ( .A(n9102), .B(n9101), .Z(n244) );
  NANDN U262 ( .A(n243), .B(n244), .Z(n245) );
  ANDN U263 ( .B(n245), .A(n12413), .Z(n246) );
  OR U264 ( .A(n12414), .B(n246), .Z(n247) );
  NANDN U265 ( .A(n9103), .B(n247), .Z(n248) );
  NANDN U266 ( .A(n12419), .B(n248), .Z(n9106) );
  NANDN U267 ( .A(n5374), .B(n4454), .Z(n249) );
  ANDN U268 ( .B(n5371), .A(n9206), .Z(n250) );
  OR U269 ( .A(n249), .B(n5372), .Z(n251) );
  AND U270 ( .A(n250), .B(n251), .Z(n252) );
  ANDN U271 ( .B(n5368), .A(n252), .Z(n253) );
  NAND U272 ( .A(n5373), .B(n253), .Z(n254) );
  ANDN U273 ( .B(n254), .A(n5370), .Z(n255) );
  NANDN U274 ( .A(n5364), .B(n255), .Z(n256) );
  NAND U275 ( .A(n5369), .B(n256), .Z(n257) );
  ANDN U276 ( .B(n257), .A(n5365), .Z(n258) );
  NANDN U277 ( .A(n12718), .B(n258), .Z(n259) );
  NANDN U278 ( .A(n12721), .B(n259), .Z(n260) );
  AND U279 ( .A(n5362), .B(n260), .Z(n261) );
  NOR U280 ( .A(n9209), .B(n261), .Z(n262) );
  NAND U281 ( .A(n12722), .B(n262), .Z(n263) );
  AND U282 ( .A(n5360), .B(n263), .Z(n4457) );
  AND U283 ( .A(n12876), .B(n5334), .Z(n264) );
  NAND U284 ( .A(n4474), .B(n4475), .Z(n265) );
  AND U285 ( .A(n264), .B(n265), .Z(n266) );
  NOR U286 ( .A(n12879), .B(n12883), .Z(n267) );
  NANDN U287 ( .A(n266), .B(n267), .Z(n268) );
  AND U288 ( .A(n5333), .B(n268), .Z(n269) );
  NAND U289 ( .A(n12885), .B(n269), .Z(n270) );
  NANDN U290 ( .A(n12886), .B(n270), .Z(n271) );
  AND U291 ( .A(n12888), .B(n271), .Z(n272) );
  NAND U292 ( .A(n272), .B(n5330), .Z(n273) );
  ANDN U293 ( .B(n273), .A(n5328), .Z(n274) );
  NANDN U294 ( .A(n12891), .B(n274), .Z(n4476) );
  ANDN U295 ( .B(n5304), .A(n5307), .Z(n275) );
  NANDN U296 ( .A(n4482), .B(n4481), .Z(n276) );
  AND U297 ( .A(n275), .B(n276), .Z(n277) );
  ANDN U298 ( .B(n5305), .A(n277), .Z(n278) );
  NAND U299 ( .A(n12943), .B(n278), .Z(n279) );
  ANDN U300 ( .B(n279), .A(n5303), .Z(n280) );
  NAND U301 ( .A(n280), .B(n12945), .Z(n281) );
  NAND U302 ( .A(n12947), .B(n281), .Z(n282) );
  AND U303 ( .A(n12949), .B(n282), .Z(n283) );
  OR U304 ( .A(n12951), .B(n283), .Z(n284) );
  AND U305 ( .A(n12953), .B(n284), .Z(n285) );
  OR U306 ( .A(n12955), .B(n285), .Z(n286) );
  NAND U307 ( .A(n12957), .B(n286), .Z(n287) );
  NANDN U308 ( .A(n12958), .B(n287), .Z(n4492) );
  ANDN U309 ( .B(n5271), .A(n9313), .Z(n288) );
  ANDN U310 ( .B(n4496), .A(n13038), .Z(n289) );
  NAND U311 ( .A(n13034), .B(n289), .Z(n290) );
  AND U312 ( .A(n288), .B(n290), .Z(n291) );
  NANDN U313 ( .A(n291), .B(n13043), .Z(n292) );
  NANDN U314 ( .A(n13044), .B(n292), .Z(n293) );
  NAND U315 ( .A(n13047), .B(n293), .Z(n294) );
  NANDN U316 ( .A(n13048), .B(n294), .Z(n295) );
  NANDN U317 ( .A(n13050), .B(n295), .Z(n296) );
  AND U318 ( .A(n13053), .B(n296), .Z(n297) );
  OR U319 ( .A(n13054), .B(n297), .Z(n298) );
  NAND U320 ( .A(n13057), .B(n298), .Z(n299) );
  NANDN U321 ( .A(n13058), .B(n299), .Z(n300) );
  NAND U322 ( .A(n13061), .B(n300), .Z(n301) );
  NANDN U323 ( .A(n13062), .B(n301), .Z(n302) );
  AND U324 ( .A(n5270), .B(n302), .Z(n4497) );
  NAND U325 ( .A(n9292), .B(n9293), .Z(n303) );
  ANDN U326 ( .B(n303), .A(n9294), .Z(n304) );
  AND U327 ( .A(n9296), .B(n9295), .Z(n305) );
  NANDN U328 ( .A(n12969), .B(n304), .Z(n306) );
  AND U329 ( .A(n305), .B(n306), .Z(n307) );
  NOR U330 ( .A(n12977), .B(n307), .Z(n308) );
  NANDN U331 ( .A(y[1302]), .B(x[1302]), .Z(n309) );
  NAND U332 ( .A(n308), .B(n309), .Z(n310) );
  AND U333 ( .A(n5294), .B(n310), .Z(n311) );
  AND U334 ( .A(n9297), .B(n311), .Z(n312) );
  ANDN U335 ( .B(n312), .A(n9299), .Z(n313) );
  NANDN U336 ( .A(n313), .B(n12981), .Z(n314) );
  NAND U337 ( .A(n12983), .B(n314), .Z(n315) );
  NANDN U338 ( .A(n12984), .B(n315), .Z(n316) );
  NAND U339 ( .A(n12986), .B(n316), .Z(n9302) );
  AND U340 ( .A(n4502), .B(n13135), .Z(n317) );
  NAND U341 ( .A(n5249), .B(n317), .Z(n318) );
  ANDN U342 ( .B(n318), .A(n5246), .Z(n319) );
  AND U343 ( .A(n5248), .B(n9362), .Z(n320) );
  NANDN U344 ( .A(n13137), .B(n319), .Z(n321) );
  NAND U345 ( .A(n320), .B(n321), .Z(n322) );
  ANDN U346 ( .B(n322), .A(n13144), .Z(n323) );
  NAND U347 ( .A(n323), .B(n5247), .Z(n324) );
  AND U348 ( .A(n13146), .B(n324), .Z(n325) );
  NAND U349 ( .A(n325), .B(n9363), .Z(n326) );
  ANDN U350 ( .B(n5242), .A(n5245), .Z(n327) );
  NANDN U351 ( .A(n13149), .B(n326), .Z(n328) );
  NAND U352 ( .A(n327), .B(n328), .Z(n4503) );
  NANDN U353 ( .A(n9407), .B(n9399), .Z(n329) );
  AND U354 ( .A(n4511), .B(n329), .Z(n4512) );
  NANDN U355 ( .A(n5224), .B(n5225), .Z(n330) );
  ANDN U356 ( .B(n9385), .A(n9387), .Z(n331) );
  NAND U357 ( .A(n9386), .B(n331), .Z(n332) );
  NANDN U358 ( .A(n330), .B(n332), .Z(n333) );
  NAND U359 ( .A(n13219), .B(n333), .Z(n334) );
  NAND U360 ( .A(n13220), .B(n334), .Z(n335) );
  ANDN U361 ( .B(n335), .A(n13223), .Z(n336) );
  NANDN U362 ( .A(n336), .B(n13225), .Z(n337) );
  ANDN U363 ( .B(n337), .A(n13227), .Z(n338) );
  ANDN U364 ( .B(n9390), .A(n338), .Z(n339) );
  NAND U365 ( .A(n13229), .B(n339), .Z(n340) );
  ANDN U366 ( .B(n340), .A(n13230), .Z(n341) );
  NANDN U367 ( .A(n13234), .B(n341), .Z(n9391) );
  NANDN U368 ( .A(n13313), .B(n4519), .Z(n342) );
  NAND U369 ( .A(n4520), .B(n342), .Z(n343) );
  NAND U370 ( .A(n13321), .B(n343), .Z(n344) );
  AND U371 ( .A(n9427), .B(n5195), .Z(n345) );
  NANDN U372 ( .A(n344), .B(n13317), .Z(n346) );
  AND U373 ( .A(n345), .B(n346), .Z(n347) );
  NOR U374 ( .A(n347), .B(n5193), .Z(n348) );
  NAND U375 ( .A(n13327), .B(n348), .Z(n349) );
  AND U376 ( .A(n9428), .B(n349), .Z(n350) );
  NAND U377 ( .A(n350), .B(n13329), .Z(n351) );
  NANDN U378 ( .A(n13331), .B(n351), .Z(n352) );
  AND U379 ( .A(n13333), .B(n352), .Z(n353) );
  NAND U380 ( .A(n5190), .B(n353), .Z(n354) );
  ANDN U381 ( .B(n354), .A(n5188), .Z(n355) );
  NANDN U382 ( .A(n13335), .B(n355), .Z(n4521) );
  AND U383 ( .A(n9446), .B(n9445), .Z(n356) );
  AND U384 ( .A(n13385), .B(n13389), .Z(n357) );
  NANDN U385 ( .A(n13383), .B(n356), .Z(n358) );
  NAND U386 ( .A(n357), .B(n358), .Z(n359) );
  AND U387 ( .A(n5169), .B(n13390), .Z(n360) );
  NAND U388 ( .A(n359), .B(n360), .Z(n361) );
  NAND U389 ( .A(n13393), .B(n361), .Z(n362) );
  NANDN U390 ( .A(n13395), .B(n362), .Z(n363) );
  NAND U391 ( .A(n13397), .B(n363), .Z(n364) );
  AND U392 ( .A(n13398), .B(n364), .Z(n365) );
  ANDN U393 ( .B(n13403), .A(n9447), .Z(n366) );
  NANDN U394 ( .A(n365), .B(n13401), .Z(n367) );
  AND U395 ( .A(n366), .B(n367), .Z(n368) );
  OR U396 ( .A(n13405), .B(n368), .Z(n369) );
  NANDN U397 ( .A(n9448), .B(n369), .Z(n370) );
  NAND U398 ( .A(n9449), .B(n370), .Z(n371) );
  AND U399 ( .A(n9450), .B(n9451), .Z(n372) );
  NAND U400 ( .A(n371), .B(n372), .Z(n373) );
  NAND U401 ( .A(n9452), .B(n373), .Z(n9453) );
  NAND U402 ( .A(n5139), .B(n5138), .Z(n374) );
  NAND U403 ( .A(n9463), .B(n9464), .Z(n375) );
  NAND U404 ( .A(n9465), .B(n375), .Z(n376) );
  AND U405 ( .A(n13468), .B(n376), .Z(n377) );
  NANDN U406 ( .A(n377), .B(n13471), .Z(n378) );
  AND U407 ( .A(n13473), .B(n378), .Z(n379) );
  NANDN U408 ( .A(n379), .B(n13475), .Z(n380) );
  NAND U409 ( .A(n13477), .B(n380), .Z(n381) );
  NANDN U410 ( .A(n9475), .B(n381), .Z(n382) );
  AND U411 ( .A(n13480), .B(n5140), .Z(n383) );
  OR U412 ( .A(n382), .B(n13479), .Z(n384) );
  AND U413 ( .A(n383), .B(n384), .Z(n385) );
  AND U414 ( .A(n5136), .B(n5137), .Z(n386) );
  OR U415 ( .A(n374), .B(n385), .Z(n387) );
  AND U416 ( .A(n386), .B(n387), .Z(n388) );
  ANDN U417 ( .B(n9477), .A(n388), .Z(n389) );
  NAND U418 ( .A(n9476), .B(n389), .Z(n390) );
  AND U419 ( .A(n13493), .B(n390), .Z(n391) );
  NANDN U420 ( .A(n9478), .B(n391), .Z(n9479) );
  NAND U421 ( .A(n4561), .B(n13507), .Z(n392) );
  AND U422 ( .A(n4562), .B(n392), .Z(n393) );
  ANDN U423 ( .B(n13515), .A(n393), .Z(n394) );
  NAND U424 ( .A(n13510), .B(n394), .Z(n395) );
  ANDN U425 ( .B(n395), .A(n5124), .Z(n396) );
  NAND U426 ( .A(n5126), .B(n396), .Z(n397) );
  NANDN U427 ( .A(n13519), .B(n397), .Z(n398) );
  NAND U428 ( .A(n13521), .B(n398), .Z(n399) );
  ANDN U429 ( .B(n13522), .A(n5119), .Z(n400) );
  NANDN U430 ( .A(n399), .B(n5122), .Z(n401) );
  AND U431 ( .A(n400), .B(n401), .Z(n402) );
  NOR U432 ( .A(n5121), .B(n402), .Z(n403) );
  NAND U433 ( .A(n5118), .B(n403), .Z(n404) );
  ANDN U434 ( .B(n404), .A(n5115), .Z(n405) );
  NAND U435 ( .A(n405), .B(n5120), .Z(n406) );
  AND U436 ( .A(n5114), .B(n406), .Z(n407) );
  NANDN U437 ( .A(n5117), .B(n407), .Z(n4563) );
  ANDN U438 ( .B(n5079), .A(n5078), .Z(n408) );
  NANDN U439 ( .A(n9521), .B(n9520), .Z(n409) );
  AND U440 ( .A(n408), .B(n409), .Z(n410) );
  NOR U441 ( .A(n13621), .B(n5077), .Z(n411) );
  NOR U442 ( .A(n13615), .B(n13619), .Z(n412) );
  NANDN U443 ( .A(n410), .B(n412), .Z(n413) );
  AND U444 ( .A(n411), .B(n413), .Z(n414) );
  AND U445 ( .A(n9524), .B(n13625), .Z(n415) );
  NANDN U446 ( .A(n414), .B(n13623), .Z(n416) );
  AND U447 ( .A(n415), .B(n416), .Z(n417) );
  NANDN U448 ( .A(n417), .B(n13626), .Z(n418) );
  NANDN U449 ( .A(n9525), .B(n418), .Z(n419) );
  NAND U450 ( .A(n13630), .B(n419), .Z(n420) );
  NANDN U451 ( .A(n13633), .B(n420), .Z(n9527) );
  NANDN U452 ( .A(n4596), .B(n13674), .Z(n421) );
  AND U453 ( .A(n4597), .B(n421), .Z(n422) );
  ANDN U454 ( .B(n4595), .A(n13672), .Z(n423) );
  NAND U455 ( .A(n13668), .B(n423), .Z(n424) );
  ANDN U456 ( .B(n424), .A(n422), .Z(n425) );
  OR U457 ( .A(n13677), .B(n425), .Z(n426) );
  NANDN U458 ( .A(n13679), .B(n426), .Z(n427) );
  NAND U459 ( .A(n5064), .B(n427), .Z(n428) );
  ANDN U460 ( .B(n13687), .A(n5065), .Z(n429) );
  OR U461 ( .A(n428), .B(n13680), .Z(n430) );
  AND U462 ( .A(n429), .B(n430), .Z(n431) );
  ANDN U463 ( .B(n5063), .A(n431), .Z(n432) );
  NAND U464 ( .A(n13688), .B(n432), .Z(n433) );
  ANDN U465 ( .B(n433), .A(n13690), .Z(n434) );
  ANDN U466 ( .B(n5061), .A(n434), .Z(n435) );
  NAND U467 ( .A(n13692), .B(n435), .Z(n436) );
  ANDN U468 ( .B(n436), .A(n9537), .Z(n4598) );
  NAND U469 ( .A(n5050), .B(n5051), .Z(n437) );
  NOR U470 ( .A(n13727), .B(n9546), .Z(n438) );
  NAND U471 ( .A(n9545), .B(n438), .Z(n439) );
  NANDN U472 ( .A(n437), .B(n439), .Z(n440) );
  ANDN U473 ( .B(n440), .A(n9547), .Z(n441) );
  NAND U474 ( .A(n441), .B(n13734), .Z(n442) );
  AND U475 ( .A(n5049), .B(n442), .Z(n443) );
  NANDN U476 ( .A(n13737), .B(n443), .Z(n444) );
  NANDN U477 ( .A(n13739), .B(n444), .Z(n445) );
  NAND U478 ( .A(n13741), .B(n445), .Z(n446) );
  ANDN U479 ( .B(n446), .A(n13742), .Z(n447) );
  ANDN U480 ( .B(n9548), .A(n447), .Z(n448) );
  NAND U481 ( .A(n13744), .B(n448), .Z(n449) );
  ANDN U482 ( .B(n449), .A(n13747), .Z(n450) );
  NANDN U483 ( .A(n13751), .B(n450), .Z(n9549) );
  NANDN U484 ( .A(n4604), .B(n4603), .Z(n451) );
  NAND U485 ( .A(n5032), .B(n451), .Z(n452) );
  NAND U486 ( .A(n9557), .B(n452), .Z(n453) );
  AND U487 ( .A(n5033), .B(n5028), .Z(n454) );
  OR U488 ( .A(n453), .B(n5030), .Z(n455) );
  AND U489 ( .A(n454), .B(n455), .Z(n456) );
  ANDN U490 ( .B(n5031), .A(n456), .Z(n457) );
  NAND U491 ( .A(n5027), .B(n457), .Z(n458) );
  AND U492 ( .A(n13780), .B(n458), .Z(n459) );
  NOR U493 ( .A(n13783), .B(n5026), .Z(n460) );
  NANDN U494 ( .A(n5029), .B(n459), .Z(n461) );
  NAND U495 ( .A(n460), .B(n461), .Z(n462) );
  NAND U496 ( .A(n13785), .B(n462), .Z(n463) );
  NAND U497 ( .A(n13787), .B(n463), .Z(n464) );
  AND U498 ( .A(n5025), .B(n464), .Z(n465) );
  NAND U499 ( .A(n13789), .B(n465), .Z(n4605) );
  NANDN U500 ( .A(n10184), .B(n10180), .Z(n466) );
  NAND U501 ( .A(n4628), .B(n466), .Z(n467) );
  NANDN U502 ( .A(n10182), .B(n467), .Z(n9635) );
  ANDN U503 ( .B(n4643), .A(n9679), .Z(n468) );
  NAND U504 ( .A(n14023), .B(n468), .Z(n469) );
  NANDN U505 ( .A(n14024), .B(n469), .Z(n470) );
  OR U506 ( .A(n470), .B(n9681), .Z(n471) );
  NAND U507 ( .A(n14026), .B(n471), .Z(n472) );
  NAND U508 ( .A(n14029), .B(n472), .Z(n473) );
  NAND U509 ( .A(n14031), .B(n473), .Z(n474) );
  NANDN U510 ( .A(n14033), .B(n474), .Z(n475) );
  AND U511 ( .A(n14035), .B(n475), .Z(n476) );
  NOR U512 ( .A(n9687), .B(n476), .Z(n477) );
  NAND U513 ( .A(n14036), .B(n477), .Z(n478) );
  ANDN U514 ( .B(n478), .A(n14039), .Z(n479) );
  NAND U515 ( .A(n479), .B(n4940), .Z(n480) );
  AND U516 ( .A(n9688), .B(n480), .Z(n481) );
  NAND U517 ( .A(n481), .B(n4938), .Z(n4644) );
  NANDN U518 ( .A(n14181), .B(n4656), .Z(n482) );
  NAND U519 ( .A(n14183), .B(n482), .Z(n483) );
  AND U520 ( .A(n9821), .B(n483), .Z(n484) );
  ANDN U521 ( .B(n9820), .A(n9823), .Z(n485) );
  NANDN U522 ( .A(n9818), .B(n484), .Z(n486) );
  NAND U523 ( .A(n485), .B(n486), .Z(n487) );
  NAND U524 ( .A(n9824), .B(n4891), .Z(n488) );
  ANDN U525 ( .B(n9822), .A(n4892), .Z(n489) );
  NAND U526 ( .A(n487), .B(n489), .Z(n490) );
  NANDN U527 ( .A(n488), .B(n490), .Z(n491) );
  ANDN U528 ( .B(n4893), .A(n9825), .Z(n492) );
  NAND U529 ( .A(n491), .B(n492), .Z(n493) );
  NAND U530 ( .A(n9828), .B(n493), .Z(n494) );
  OR U531 ( .A(n494), .B(n4890), .Z(n495) );
  NAND U532 ( .A(n14201), .B(n495), .Z(n496) );
  NAND U533 ( .A(n14203), .B(n496), .Z(n4657) );
  NANDN U534 ( .A(n4659), .B(n4660), .Z(n497) );
  NAND U535 ( .A(n14255), .B(n497), .Z(n498) );
  AND U536 ( .A(n14257), .B(n498), .Z(n499) );
  OR U537 ( .A(n499), .B(n14259), .Z(n500) );
  NANDN U538 ( .A(n14260), .B(n500), .Z(n501) );
  AND U539 ( .A(n14262), .B(n501), .Z(n502) );
  NANDN U540 ( .A(n502), .B(n14265), .Z(n503) );
  NAND U541 ( .A(n14267), .B(n503), .Z(n504) );
  NAND U542 ( .A(n9862), .B(n504), .Z(n505) );
  OR U543 ( .A(n14271), .B(n4662), .Z(n506) );
  OR U544 ( .A(n505), .B(n14275), .Z(n507) );
  AND U545 ( .A(n506), .B(n507), .Z(n508) );
  NANDN U546 ( .A(n508), .B(n9874), .Z(n509) );
  NAND U547 ( .A(n14278), .B(n509), .Z(n510) );
  NAND U548 ( .A(n14281), .B(n510), .Z(n4663) );
  ANDN U549 ( .B(n4837), .A(n14336), .Z(n511) );
  NANDN U550 ( .A(n14334), .B(n4666), .Z(n512) );
  AND U551 ( .A(n511), .B(n512), .Z(n513) );
  ANDN U552 ( .B(n9927), .A(n4836), .Z(n514) );
  OR U553 ( .A(n14340), .B(n513), .Z(n515) );
  AND U554 ( .A(n514), .B(n515), .Z(n516) );
  NOR U555 ( .A(n14342), .B(n4834), .Z(n517) );
  NANDN U556 ( .A(n516), .B(n517), .Z(n518) );
  AND U557 ( .A(n9926), .B(n518), .Z(n519) );
  NAND U558 ( .A(n4831), .B(n519), .Z(n520) );
  ANDN U559 ( .B(n520), .A(n4829), .Z(n521) );
  NANDN U560 ( .A(n4833), .B(n521), .Z(n522) );
  AND U561 ( .A(n4832), .B(n14355), .Z(n523) );
  NAND U562 ( .A(n522), .B(n523), .Z(n524) );
  NANDN U563 ( .A(n14356), .B(n524), .Z(n4667) );
  NAND U564 ( .A(n4675), .B(n4674), .Z(n525) );
  NANDN U565 ( .A(n4676), .B(n525), .Z(n526) );
  NANDN U566 ( .A(n14467), .B(n526), .Z(n527) );
  NAND U567 ( .A(n14469), .B(n527), .Z(n528) );
  NANDN U568 ( .A(n14471), .B(n528), .Z(n529) );
  AND U569 ( .A(n14473), .B(n529), .Z(n530) );
  ANDN U570 ( .B(n4783), .A(n14476), .Z(n531) );
  NANDN U571 ( .A(n530), .B(n14474), .Z(n532) );
  AND U572 ( .A(n531), .B(n532), .Z(n533) );
  ANDN U573 ( .B(n4781), .A(n533), .Z(n534) );
  NAND U574 ( .A(n14478), .B(n534), .Z(n535) );
  ANDN U575 ( .B(n535), .A(n14484), .Z(n536) );
  NANDN U576 ( .A(n4782), .B(n536), .Z(n4677) );
  NANDN U577 ( .A(n10130), .B(n4694), .Z(n537) );
  NAND U578 ( .A(n10131), .B(n537), .Z(n538) );
  AND U579 ( .A(n14576), .B(n538), .Z(n539) );
  ANDN U580 ( .B(n10133), .A(n539), .Z(n540) );
  NAND U581 ( .A(n10134), .B(n540), .Z(n541) );
  AND U582 ( .A(n14584), .B(n541), .Z(n542) );
  NAND U583 ( .A(n542), .B(n14580), .Z(n543) );
  AND U584 ( .A(n10135), .B(n543), .Z(n544) );
  NANDN U585 ( .A(n14586), .B(n544), .Z(n545) );
  NANDN U586 ( .A(n14588), .B(n545), .Z(n546) );
  NAND U587 ( .A(n14591), .B(n546), .Z(n547) );
  ANDN U588 ( .B(n547), .A(n14592), .Z(n548) );
  ANDN U589 ( .B(n4757), .A(n548), .Z(n549) );
  NAND U590 ( .A(n14595), .B(n549), .Z(n550) );
  AND U591 ( .A(n14601), .B(n550), .Z(n551) );
  ANDN U592 ( .B(n10139), .A(n4756), .Z(n552) );
  NANDN U593 ( .A(n4759), .B(n551), .Z(n553) );
  NAND U594 ( .A(n552), .B(n553), .Z(n4698) );
  OR U595 ( .A(n14685), .B(n14684), .Z(n554) );
  NAND U596 ( .A(n14686), .B(n554), .Z(n555) );
  AND U597 ( .A(n14687), .B(n555), .Z(n556) );
  OR U598 ( .A(n14688), .B(n556), .Z(n557) );
  AND U599 ( .A(n14689), .B(n557), .Z(n558) );
  ANDN U600 ( .B(n14690), .A(n558), .Z(n559) );
  NANDN U601 ( .A(x[2031]), .B(y[2031]), .Z(n560) );
  NAND U602 ( .A(n559), .B(n560), .Z(n561) );
  NANDN U603 ( .A(n14691), .B(n561), .Z(n562) );
  NAND U604 ( .A(n14692), .B(n562), .Z(n563) );
  AND U605 ( .A(n14693), .B(n563), .Z(n564) );
  NANDN U606 ( .A(n564), .B(n14694), .Z(n565) );
  NAND U607 ( .A(n14695), .B(n565), .Z(n566) );
  NAND U608 ( .A(n14696), .B(n566), .Z(n567) );
  NAND U609 ( .A(n14697), .B(n567), .Z(n568) );
  NANDN U610 ( .A(y[2039]), .B(n568), .Z(n569) );
  AND U611 ( .A(n14698), .B(n569), .Z(n570) );
  XNOR U612 ( .A(y[2039]), .B(n568), .Z(n571) );
  NAND U613 ( .A(n571), .B(x[2039]), .Z(n572) );
  NAND U614 ( .A(n570), .B(n572), .Z(n14699) );
  NAND U615 ( .A(n11603), .B(n4319), .Z(n573) );
  NANDN U616 ( .A(n11605), .B(n573), .Z(n574) );
  NAND U617 ( .A(n11607), .B(n574), .Z(n575) );
  NANDN U618 ( .A(n11609), .B(n575), .Z(n576) );
  NAND U619 ( .A(n11611), .B(n576), .Z(n577) );
  AND U620 ( .A(n11613), .B(n577), .Z(n578) );
  OR U621 ( .A(n11615), .B(n578), .Z(n579) );
  NAND U622 ( .A(n11617), .B(n579), .Z(n580) );
  NAND U623 ( .A(n11619), .B(n580), .Z(n581) );
  NAND U624 ( .A(n11620), .B(n581), .Z(n582) );
  NAND U625 ( .A(n11623), .B(n582), .Z(n583) );
  AND U626 ( .A(n11625), .B(n583), .Z(n584) );
  NANDN U627 ( .A(n584), .B(n11627), .Z(n585) );
  AND U628 ( .A(n11629), .B(n585), .Z(n4322) );
  NAND U629 ( .A(n4328), .B(n4327), .Z(n586) );
  NANDN U630 ( .A(n4329), .B(n586), .Z(n587) );
  NANDN U631 ( .A(n11678), .B(n587), .Z(n588) );
  NAND U632 ( .A(n11680), .B(n588), .Z(n589) );
  NANDN U633 ( .A(n11683), .B(n589), .Z(n590) );
  AND U634 ( .A(n11685), .B(n590), .Z(n591) );
  OR U635 ( .A(n11687), .B(n591), .Z(n592) );
  AND U636 ( .A(n11689), .B(n592), .Z(n593) );
  OR U637 ( .A(n593), .B(n11690), .Z(n594) );
  NAND U638 ( .A(n11692), .B(n594), .Z(n595) );
  NANDN U639 ( .A(n11695), .B(n595), .Z(n4330) );
  NAND U640 ( .A(n4386), .B(n11897), .Z(n596) );
  NANDN U641 ( .A(n11899), .B(n596), .Z(n597) );
  AND U642 ( .A(n11901), .B(n597), .Z(n598) );
  NANDN U643 ( .A(n598), .B(n11902), .Z(n599) );
  AND U644 ( .A(n11905), .B(n599), .Z(n600) );
  ANDN U645 ( .B(n5608), .A(n600), .Z(n601) );
  NAND U646 ( .A(n11907), .B(n601), .Z(n602) );
  AND U647 ( .A(n11908), .B(n602), .Z(n603) );
  NAND U648 ( .A(n5606), .B(n603), .Z(n604) );
  ANDN U649 ( .B(n604), .A(n5605), .Z(n605) );
  NANDN U650 ( .A(n5609), .B(n605), .Z(n606) );
  AND U651 ( .A(n5602), .B(n5607), .Z(n607) );
  NAND U652 ( .A(n606), .B(n607), .Z(n608) );
  NAND U653 ( .A(n5604), .B(n608), .Z(n609) );
  AND U654 ( .A(n5603), .B(n5598), .Z(n610) );
  OR U655 ( .A(n609), .B(n5601), .Z(n611) );
  AND U656 ( .A(n610), .B(n611), .Z(n4388) );
  NOR U657 ( .A(n11971), .B(n5570), .Z(n612) );
  NANDN U658 ( .A(n4394), .B(n4393), .Z(n613) );
  AND U659 ( .A(n612), .B(n613), .Z(n614) );
  NOR U660 ( .A(n8817), .B(n614), .Z(n615) );
  NAND U661 ( .A(n11977), .B(n615), .Z(n616) );
  AND U662 ( .A(n5571), .B(n616), .Z(n617) );
  NANDN U663 ( .A(n11978), .B(n617), .Z(n618) );
  NAND U664 ( .A(n11980), .B(n618), .Z(n619) );
  AND U665 ( .A(n5569), .B(n619), .Z(n620) );
  AND U666 ( .A(n11985), .B(n11989), .Z(n621) );
  NANDN U667 ( .A(n11983), .B(n620), .Z(n622) );
  NAND U668 ( .A(n621), .B(n622), .Z(n4395) );
  AND U669 ( .A(n8723), .B(n8724), .Z(n623) );
  NANDN U670 ( .A(n8722), .B(n8721), .Z(n624) );
  NAND U671 ( .A(n623), .B(n624), .Z(n625) );
  NOR U672 ( .A(n8726), .B(n8725), .Z(n626) );
  NAND U673 ( .A(n625), .B(n626), .Z(n627) );
  NAND U674 ( .A(n8727), .B(n627), .Z(n628) );
  ANDN U675 ( .B(n8728), .A(n8729), .Z(n629) );
  NANDN U676 ( .A(n628), .B(n11829), .Z(n630) );
  AND U677 ( .A(n629), .B(n630), .Z(n631) );
  NANDN U678 ( .A(n631), .B(n11833), .Z(n632) );
  ANDN U679 ( .B(n632), .A(n11834), .Z(n633) );
  ANDN U680 ( .B(n11836), .A(n11841), .Z(n634) );
  NANDN U681 ( .A(n8730), .B(n633), .Z(n635) );
  NAND U682 ( .A(n634), .B(n635), .Z(n636) );
  AND U683 ( .A(n8731), .B(n11842), .Z(n637) );
  NAND U684 ( .A(n636), .B(n637), .Z(n638) );
  NANDN U685 ( .A(n11845), .B(n638), .Z(n8732) );
  AND U686 ( .A(n5559), .B(n12037), .Z(n639) );
  NANDN U687 ( .A(n5557), .B(n4397), .Z(n640) );
  NAND U688 ( .A(n639), .B(n640), .Z(n641) );
  NAND U689 ( .A(n5556), .B(n12038), .Z(n642) );
  NAND U690 ( .A(n4398), .B(n642), .Z(n643) );
  AND U691 ( .A(n641), .B(n643), .Z(n644) );
  NANDN U692 ( .A(n644), .B(n12041), .Z(n645) );
  NANDN U693 ( .A(n12042), .B(n645), .Z(n646) );
  NAND U694 ( .A(n12044), .B(n646), .Z(n647) );
  NANDN U695 ( .A(n12047), .B(n647), .Z(n648) );
  NAND U696 ( .A(n12049), .B(n648), .Z(n649) );
  ANDN U697 ( .B(n649), .A(n12051), .Z(n650) );
  NAND U698 ( .A(n5549), .B(n650), .Z(n4406) );
  NANDN U699 ( .A(n12107), .B(n4412), .Z(n651) );
  NANDN U700 ( .A(n12109), .B(n651), .Z(n652) );
  AND U701 ( .A(n12111), .B(n652), .Z(n653) );
  OR U702 ( .A(n12113), .B(n653), .Z(n654) );
  NAND U703 ( .A(n12115), .B(n654), .Z(n655) );
  NANDN U704 ( .A(n12117), .B(n655), .Z(n656) );
  NAND U705 ( .A(n12119), .B(n656), .Z(n657) );
  NANDN U706 ( .A(n12121), .B(n657), .Z(n658) );
  AND U707 ( .A(n12123), .B(n658), .Z(n659) );
  OR U708 ( .A(n12125), .B(n659), .Z(n660) );
  NAND U709 ( .A(n12127), .B(n660), .Z(n661) );
  NANDN U710 ( .A(n12129), .B(n661), .Z(n662) );
  NAND U711 ( .A(n12131), .B(n662), .Z(n663) );
  NANDN U712 ( .A(n12133), .B(n663), .Z(n664) );
  ANDN U713 ( .B(n664), .A(n12135), .Z(n665) );
  NAND U714 ( .A(n5531), .B(n665), .Z(n666) );
  ANDN U715 ( .B(n666), .A(n5529), .Z(n667) );
  NANDN U716 ( .A(n12137), .B(n667), .Z(n668) );
  AND U717 ( .A(n5530), .B(n668), .Z(n4413) );
  NAND U718 ( .A(n5519), .B(n4417), .Z(n669) );
  ANDN U719 ( .B(n669), .A(n5516), .Z(n670) );
  NANDN U720 ( .A(n8986), .B(n670), .Z(n671) );
  ANDN U721 ( .B(n12209), .A(n5518), .Z(n672) );
  NAND U722 ( .A(n671), .B(n672), .Z(n673) );
  NAND U723 ( .A(n5515), .B(n673), .Z(n674) );
  NANDN U724 ( .A(n674), .B(n5517), .Z(n675) );
  ANDN U725 ( .B(n675), .A(n12212), .Z(n676) );
  AND U726 ( .A(n12221), .B(n12216), .Z(n677) );
  ANDN U727 ( .B(n5513), .A(n676), .Z(n678) );
  NAND U728 ( .A(n12213), .B(n678), .Z(n679) );
  AND U729 ( .A(n677), .B(n679), .Z(n680) );
  NOR U730 ( .A(n12222), .B(n5514), .Z(n681) );
  NANDN U731 ( .A(n680), .B(n681), .Z(n682) );
  AND U732 ( .A(n12225), .B(n682), .Z(n4419) );
  NAND U733 ( .A(n8886), .B(n12068), .Z(n683) );
  AND U734 ( .A(n12071), .B(n683), .Z(n684) );
  NOR U735 ( .A(n8887), .B(n12073), .Z(n685) );
  NANDN U736 ( .A(n684), .B(n685), .Z(n686) );
  NAND U737 ( .A(n8888), .B(n686), .Z(n687) );
  NOR U738 ( .A(n8890), .B(n8889), .Z(n688) );
  NANDN U739 ( .A(n687), .B(n12074), .Z(n689) );
  AND U740 ( .A(n688), .B(n689), .Z(n690) );
  ANDN U741 ( .B(n8891), .A(n690), .Z(n691) );
  NAND U742 ( .A(n8892), .B(n691), .Z(n692) );
  ANDN U743 ( .B(n692), .A(n8893), .Z(n693) );
  AND U744 ( .A(n12087), .B(n5541), .Z(n694) );
  NANDN U745 ( .A(n8894), .B(n693), .Z(n695) );
  NAND U746 ( .A(n694), .B(n695), .Z(n696) );
  AND U747 ( .A(n8895), .B(n12089), .Z(n697) );
  NAND U748 ( .A(n696), .B(n697), .Z(n698) );
  NAND U749 ( .A(n12091), .B(n698), .Z(n699) );
  NANDN U750 ( .A(n12093), .B(n699), .Z(n700) );
  NAND U751 ( .A(n12095), .B(n700), .Z(n8896) );
  NAND U752 ( .A(n5499), .B(n4424), .Z(n701) );
  AND U753 ( .A(n5497), .B(n5493), .Z(n702) );
  NANDN U754 ( .A(n701), .B(n4425), .Z(n703) );
  AND U755 ( .A(n702), .B(n703), .Z(n704) );
  NOR U756 ( .A(n12308), .B(n704), .Z(n705) );
  NAND U757 ( .A(n5495), .B(n705), .Z(n706) );
  AND U758 ( .A(n5492), .B(n706), .Z(n707) );
  NAND U759 ( .A(n12310), .B(n707), .Z(n708) );
  NANDN U760 ( .A(n12313), .B(n708), .Z(n709) );
  NAND U761 ( .A(n12315), .B(n709), .Z(n710) );
  AND U762 ( .A(n5489), .B(n12316), .Z(n711) );
  NANDN U763 ( .A(n710), .B(n5490), .Z(n712) );
  AND U764 ( .A(n711), .B(n712), .Z(n713) );
  ANDN U765 ( .B(n5486), .A(n713), .Z(n714) );
  NAND U766 ( .A(n5491), .B(n714), .Z(n715) );
  ANDN U767 ( .B(n715), .A(n5488), .Z(n716) );
  NANDN U768 ( .A(n5484), .B(n716), .Z(n4426) );
  AND U769 ( .A(n8961), .B(n8962), .Z(n717) );
  NAND U770 ( .A(n8963), .B(n717), .Z(n718) );
  NANDN U771 ( .A(n8964), .B(n718), .Z(n719) );
  OR U772 ( .A(n719), .B(n8965), .Z(n720) );
  NAND U773 ( .A(n8966), .B(n720), .Z(n721) );
  NANDN U774 ( .A(n8967), .B(n721), .Z(n722) );
  AND U775 ( .A(n12175), .B(n12170), .Z(n723) );
  OR U776 ( .A(n722), .B(n8968), .Z(n724) );
  AND U777 ( .A(n723), .B(n724), .Z(n725) );
  ANDN U778 ( .B(n8969), .A(n725), .Z(n726) );
  NAND U779 ( .A(n12177), .B(n726), .Z(n727) );
  AND U780 ( .A(n12179), .B(n727), .Z(n728) );
  AND U781 ( .A(n12183), .B(n8971), .Z(n729) );
  OR U782 ( .A(n8970), .B(n728), .Z(n730) );
  AND U783 ( .A(n729), .B(n730), .Z(n731) );
  NOR U784 ( .A(n731), .B(n8973), .Z(n732) );
  NAND U785 ( .A(n8972), .B(n732), .Z(n733) );
  ANDN U786 ( .B(n733), .A(n8974), .Z(n8975) );
  ANDN U787 ( .B(n4431), .A(n5469), .Z(n734) );
  NAND U788 ( .A(n12374), .B(n734), .Z(n735) );
  AND U789 ( .A(n12377), .B(n735), .Z(n736) );
  OR U790 ( .A(n5467), .B(n736), .Z(n737) );
  AND U791 ( .A(n12381), .B(n737), .Z(n738) );
  NANDN U792 ( .A(n5461), .B(n5466), .Z(n739) );
  NAND U793 ( .A(n4432), .B(n739), .Z(n740) );
  ANDN U794 ( .B(n740), .A(n738), .Z(n741) );
  NAND U795 ( .A(n741), .B(n5465), .Z(n742) );
  NANDN U796 ( .A(n5457), .B(n742), .Z(n743) );
  AND U797 ( .A(n5462), .B(n743), .Z(n744) );
  NAND U798 ( .A(n5456), .B(n744), .Z(n745) );
  ANDN U799 ( .B(n745), .A(n5458), .Z(n746) );
  NANDN U800 ( .A(n12388), .B(n746), .Z(n4433) );
  ANDN U801 ( .B(n12254), .A(n9007), .Z(n747) );
  NAND U802 ( .A(n9006), .B(n9005), .Z(n748) );
  AND U803 ( .A(n747), .B(n748), .Z(n749) );
  ANDN U804 ( .B(n9008), .A(n749), .Z(n750) );
  NAND U805 ( .A(n12257), .B(n750), .Z(n751) );
  ANDN U806 ( .B(n751), .A(n12259), .Z(n752) );
  NANDN U807 ( .A(n752), .B(n12261), .Z(n753) );
  NAND U808 ( .A(n12263), .B(n753), .Z(n754) );
  NAND U809 ( .A(n9013), .B(n754), .Z(n755) );
  ANDN U810 ( .B(n9016), .A(n9015), .Z(n756) );
  OR U811 ( .A(n755), .B(n9014), .Z(n757) );
  AND U812 ( .A(n756), .B(n757), .Z(n758) );
  ANDN U813 ( .B(n9017), .A(n758), .Z(n759) );
  NAND U814 ( .A(n9018), .B(n759), .Z(n760) );
  ANDN U815 ( .B(n760), .A(n9019), .Z(n761) );
  ANDN U816 ( .B(n9021), .A(n9022), .Z(n762) );
  NANDN U817 ( .A(n9020), .B(n761), .Z(n763) );
  NAND U818 ( .A(n762), .B(n763), .Z(n764) );
  NAND U819 ( .A(n9023), .B(n764), .Z(n9024) );
  NANDN U820 ( .A(n4438), .B(n4437), .Z(n765) );
  NAND U821 ( .A(n12445), .B(n765), .Z(n766) );
  NANDN U822 ( .A(n12447), .B(n766), .Z(n767) );
  ANDN U823 ( .B(n5438), .A(n12448), .Z(n768) );
  NAND U824 ( .A(n767), .B(n768), .Z(n769) );
  NANDN U825 ( .A(n12454), .B(n769), .Z(n770) );
  AND U826 ( .A(n12457), .B(n5437), .Z(n771) );
  NANDN U827 ( .A(n770), .B(n12450), .Z(n772) );
  AND U828 ( .A(n771), .B(n772), .Z(n773) );
  AND U829 ( .A(n9120), .B(n12461), .Z(n774) );
  OR U830 ( .A(n12459), .B(n773), .Z(n775) );
  AND U831 ( .A(n774), .B(n775), .Z(n776) );
  NOR U832 ( .A(n776), .B(n5434), .Z(n777) );
  NAND U833 ( .A(n12467), .B(n777), .Z(n778) );
  AND U834 ( .A(n12468), .B(n778), .Z(n779) );
  NAND U835 ( .A(n779), .B(n9119), .Z(n780) );
  NANDN U836 ( .A(n12471), .B(n780), .Z(n781) );
  AND U837 ( .A(n9122), .B(n781), .Z(n782) );
  NAND U838 ( .A(n12473), .B(n782), .Z(n4439) );
  NAND U839 ( .A(n4443), .B(n4442), .Z(n783) );
  AND U840 ( .A(n12530), .B(n783), .Z(n784) );
  NANDN U841 ( .A(n9145), .B(n784), .Z(n785) );
  AND U842 ( .A(n4444), .B(n5419), .Z(n786) );
  NAND U843 ( .A(n785), .B(n786), .Z(n787) );
  NANDN U844 ( .A(n12539), .B(n787), .Z(n788) );
  AND U845 ( .A(n5417), .B(n12541), .Z(n789) );
  NAND U846 ( .A(n788), .B(n789), .Z(n790) );
  NAND U847 ( .A(n12542), .B(n790), .Z(n791) );
  AND U848 ( .A(n5416), .B(n5413), .Z(n792) );
  NANDN U849 ( .A(n791), .B(n5414), .Z(n793) );
  AND U850 ( .A(n792), .B(n793), .Z(n794) );
  NOR U851 ( .A(n12551), .B(n5415), .Z(n795) );
  NANDN U852 ( .A(n794), .B(n795), .Z(n796) );
  AND U853 ( .A(n12553), .B(n796), .Z(n797) );
  NAND U854 ( .A(n5412), .B(n797), .Z(n798) );
  NANDN U855 ( .A(n12555), .B(n798), .Z(n799) );
  AND U856 ( .A(n12557), .B(n799), .Z(n800) );
  NAND U857 ( .A(n5411), .B(n800), .Z(n4445) );
  AND U858 ( .A(n12421), .B(n5443), .Z(n9107) );
  NANDN U859 ( .A(n9174), .B(n4447), .Z(n801) );
  ANDN U860 ( .B(n5405), .A(n12610), .Z(n802) );
  OR U861 ( .A(n801), .B(n5406), .Z(n803) );
  AND U862 ( .A(n802), .B(n803), .Z(n804) );
  OR U863 ( .A(n804), .B(n12613), .Z(n805) );
  AND U864 ( .A(n12615), .B(n805), .Z(n806) );
  NOR U865 ( .A(n806), .B(n12617), .Z(n807) );
  NANDN U866 ( .A(n5402), .B(n807), .Z(n808) );
  NAND U867 ( .A(n5400), .B(n808), .Z(n809) );
  AND U868 ( .A(n5398), .B(n5401), .Z(n810) );
  OR U869 ( .A(n809), .B(n12619), .Z(n811) );
  AND U870 ( .A(n810), .B(n811), .Z(n812) );
  NOR U871 ( .A(n12626), .B(n812), .Z(n813) );
  NAND U872 ( .A(n5399), .B(n813), .Z(n814) );
  AND U873 ( .A(n12628), .B(n814), .Z(n815) );
  NAND U874 ( .A(n5397), .B(n815), .Z(n4448) );
  ANDN U875 ( .B(n5430), .A(n5429), .Z(n816) );
  NANDN U876 ( .A(n9124), .B(n9123), .Z(n817) );
  NAND U877 ( .A(n816), .B(n817), .Z(n818) );
  NANDN U878 ( .A(n9125), .B(n9126), .Z(n819) );
  AND U879 ( .A(n12485), .B(n12480), .Z(n820) );
  NAND U880 ( .A(n818), .B(n820), .Z(n821) );
  NANDN U881 ( .A(n819), .B(n821), .Z(n822) );
  AND U882 ( .A(n12491), .B(n9127), .Z(n823) );
  NANDN U883 ( .A(n12489), .B(n822), .Z(n824) );
  NAND U884 ( .A(n823), .B(n824), .Z(n825) );
  ANDN U885 ( .B(n12493), .A(n9128), .Z(n826) );
  NAND U886 ( .A(n825), .B(n826), .Z(n827) );
  NAND U887 ( .A(n9129), .B(n827), .Z(n828) );
  NANDN U888 ( .A(n828), .B(n9130), .Z(n829) );
  ANDN U889 ( .B(n829), .A(n9131), .Z(n830) );
  AND U890 ( .A(n9134), .B(n9133), .Z(n831) );
  NANDN U891 ( .A(n9132), .B(n830), .Z(n832) );
  NAND U892 ( .A(n831), .B(n832), .Z(n9135) );
  AND U893 ( .A(n4453), .B(n5378), .Z(n833) );
  NAND U894 ( .A(n12686), .B(n833), .Z(n834) );
  NANDN U895 ( .A(n9201), .B(n834), .Z(n835) );
  AND U896 ( .A(n12695), .B(n5379), .Z(n836) );
  OR U897 ( .A(n835), .B(n5381), .Z(n837) );
  AND U898 ( .A(n836), .B(n837), .Z(n838) );
  NOR U899 ( .A(n12697), .B(n9202), .Z(n839) );
  NANDN U900 ( .A(n838), .B(n839), .Z(n840) );
  ANDN U901 ( .B(n840), .A(n12698), .Z(n841) );
  ANDN U902 ( .B(n5376), .A(n841), .Z(n842) );
  NAND U903 ( .A(n12700), .B(n842), .Z(n843) );
  AND U904 ( .A(n5375), .B(n843), .Z(n844) );
  AND U905 ( .A(n5377), .B(n9207), .Z(n845) );
  NANDN U906 ( .A(n12703), .B(n844), .Z(n846) );
  NAND U907 ( .A(n845), .B(n846), .Z(n4454) );
  NAND U908 ( .A(n12562), .B(n9152), .Z(n847) );
  NANDN U909 ( .A(n12564), .B(n847), .Z(n848) );
  NAND U910 ( .A(n9155), .B(n848), .Z(n849) );
  ANDN U911 ( .B(n12573), .A(n12569), .Z(n850) );
  NANDN U912 ( .A(n849), .B(n12566), .Z(n851) );
  AND U913 ( .A(n850), .B(n851), .Z(n852) );
  NOR U914 ( .A(n9156), .B(n852), .Z(n853) );
  NAND U915 ( .A(n12575), .B(n853), .Z(n854) );
  AND U916 ( .A(n12577), .B(n854), .Z(n855) );
  OR U917 ( .A(n12578), .B(n855), .Z(n856) );
  AND U918 ( .A(n9159), .B(n856), .Z(n857) );
  ANDN U919 ( .B(n12582), .A(n9160), .Z(n858) );
  NANDN U920 ( .A(n12580), .B(n857), .Z(n859) );
  NAND U921 ( .A(n858), .B(n859), .Z(n860) );
  AND U922 ( .A(n9162), .B(n9161), .Z(n861) );
  NAND U923 ( .A(n860), .B(n861), .Z(n862) );
  NANDN U924 ( .A(n9163), .B(n862), .Z(n9164) );
  ANDN U925 ( .B(n5349), .A(n12773), .Z(n863) );
  NAND U926 ( .A(n4462), .B(n12770), .Z(n864) );
  AND U927 ( .A(n863), .B(n864), .Z(n865) );
  ANDN U928 ( .B(n12779), .A(n865), .Z(n866) );
  NAND U929 ( .A(n12775), .B(n866), .Z(n867) );
  ANDN U930 ( .B(n867), .A(n12780), .Z(n868) );
  NAND U931 ( .A(n868), .B(n5348), .Z(n869) );
  NANDN U932 ( .A(n12783), .B(n869), .Z(n870) );
  AND U933 ( .A(n12785), .B(n870), .Z(n871) );
  ANDN U934 ( .B(n5347), .A(n12789), .Z(n872) );
  OR U935 ( .A(n12787), .B(n871), .Z(n873) );
  AND U936 ( .A(n872), .B(n873), .Z(n874) );
  ANDN U937 ( .B(n12791), .A(n874), .Z(n875) );
  NAND U938 ( .A(n12794), .B(n875), .Z(n876) );
  AND U939 ( .A(n5346), .B(n876), .Z(n877) );
  NANDN U940 ( .A(n12797), .B(n877), .Z(n878) );
  NANDN U941 ( .A(n12799), .B(n878), .Z(n879) );
  AND U942 ( .A(n9238), .B(n879), .Z(n880) );
  NAND U943 ( .A(n12801), .B(n880), .Z(n4465) );
  ANDN U944 ( .B(n5393), .A(n5392), .Z(n881) );
  OR U945 ( .A(n9186), .B(n9187), .Z(n882) );
  NAND U946 ( .A(n881), .B(n882), .Z(n883) );
  AND U947 ( .A(n12655), .B(n9188), .Z(n884) );
  NANDN U948 ( .A(n12653), .B(n883), .Z(n885) );
  NAND U949 ( .A(n884), .B(n885), .Z(n886) );
  ANDN U950 ( .B(n12657), .A(n9189), .Z(n887) );
  NAND U951 ( .A(n886), .B(n887), .Z(n888) );
  NAND U952 ( .A(n9190), .B(n888), .Z(n889) );
  AND U953 ( .A(n5388), .B(n5389), .Z(n890) );
  OR U954 ( .A(n889), .B(n9191), .Z(n891) );
  AND U955 ( .A(n890), .B(n891), .Z(n892) );
  NOR U956 ( .A(n9192), .B(n9193), .Z(n893) );
  NANDN U957 ( .A(n892), .B(n893), .Z(n894) );
  AND U958 ( .A(n9194), .B(n894), .Z(n895) );
  AND U959 ( .A(n5387), .B(n5386), .Z(n896) );
  NANDN U960 ( .A(n9195), .B(n895), .Z(n897) );
  NAND U961 ( .A(n896), .B(n897), .Z(n9196) );
  AND U962 ( .A(n4473), .B(n12854), .Z(n898) );
  NAND U963 ( .A(n12851), .B(n898), .Z(n899) );
  NAND U964 ( .A(n5340), .B(n899), .Z(n900) );
  OR U965 ( .A(n12857), .B(n900), .Z(n901) );
  ANDN U966 ( .B(n901), .A(n12859), .Z(n902) );
  ANDN U967 ( .B(n5338), .A(n902), .Z(n903) );
  NAND U968 ( .A(n12861), .B(n903), .Z(n904) );
  NANDN U969 ( .A(n12863), .B(n904), .Z(n905) );
  AND U970 ( .A(n5339), .B(n9261), .Z(n906) );
  OR U971 ( .A(n905), .B(n5336), .Z(n907) );
  AND U972 ( .A(n906), .B(n907), .Z(n908) );
  NOR U973 ( .A(n12870), .B(n908), .Z(n909) );
  NAND U974 ( .A(n5337), .B(n909), .Z(n910) );
  AND U975 ( .A(n12872), .B(n910), .Z(n911) );
  NAND U976 ( .A(n9262), .B(n911), .Z(n4474) );
  NANDN U977 ( .A(n9211), .B(n9210), .Z(n912) );
  NAND U978 ( .A(n12734), .B(n912), .Z(n913) );
  AND U979 ( .A(n12737), .B(n913), .Z(n914) );
  AND U980 ( .A(n12740), .B(n9212), .Z(n915) );
  OR U981 ( .A(n12739), .B(n914), .Z(n916) );
  AND U982 ( .A(n915), .B(n916), .Z(n917) );
  NOR U983 ( .A(n9213), .B(n917), .Z(n918) );
  NAND U984 ( .A(n12743), .B(n918), .Z(n919) );
  AND U985 ( .A(n9214), .B(n919), .Z(n920) );
  NAND U986 ( .A(n9215), .B(n920), .Z(n921) );
  ANDN U987 ( .B(n921), .A(n9216), .Z(n922) );
  NANDN U988 ( .A(n9217), .B(n922), .Z(n923) );
  ANDN U989 ( .B(n9218), .A(n12753), .Z(n924) );
  NAND U990 ( .A(n923), .B(n924), .Z(n925) );
  NANDN U991 ( .A(n9219), .B(n925), .Z(n926) );
  NANDN U992 ( .A(n926), .B(n12755), .Z(n927) );
  NAND U993 ( .A(n12757), .B(n927), .Z(n928) );
  NAND U994 ( .A(n12758), .B(n928), .Z(n929) );
  NAND U995 ( .A(n12761), .B(n929), .Z(n9224) );
  NANDN U996 ( .A(n12807), .B(n9244), .Z(n930) );
  NAND U997 ( .A(n12809), .B(n930), .Z(n931) );
  NANDN U998 ( .A(n12811), .B(n931), .Z(n932) );
  ANDN U999 ( .B(n12813), .A(n9245), .Z(n933) );
  NAND U1000 ( .A(n932), .B(n933), .Z(n934) );
  NAND U1001 ( .A(n9246), .B(n934), .Z(n935) );
  NOR U1002 ( .A(n9247), .B(n9248), .Z(n936) );
  OR U1003 ( .A(n935), .B(n12814), .Z(n937) );
  AND U1004 ( .A(n936), .B(n937), .Z(n938) );
  AND U1005 ( .A(n9250), .B(n9249), .Z(n939) );
  NANDN U1006 ( .A(y[1238]), .B(x[1238]), .Z(n940) );
  NANDN U1007 ( .A(n938), .B(n939), .Z(n941) );
  NAND U1008 ( .A(n940), .B(n941), .Z(n942) );
  AND U1009 ( .A(n12826), .B(n9251), .Z(n943) );
  OR U1010 ( .A(n942), .B(n12825), .Z(n944) );
  AND U1011 ( .A(n943), .B(n944), .Z(n945) );
  AND U1012 ( .A(n9252), .B(n12831), .Z(n946) );
  OR U1013 ( .A(n945), .B(n12829), .Z(n947) );
  NAND U1014 ( .A(n946), .B(n947), .Z(n9253) );
  AND U1015 ( .A(n4492), .B(n5295), .Z(n948) );
  NAND U1016 ( .A(n12960), .B(n948), .Z(n949) );
  AND U1017 ( .A(n12963), .B(n949), .Z(n950) );
  ANDN U1018 ( .B(n5300), .A(n950), .Z(n951) );
  OR U1019 ( .A(n3404), .B(n5296), .Z(n952) );
  NAND U1020 ( .A(n951), .B(n952), .Z(n953) );
  NAND U1021 ( .A(n12966), .B(n953), .Z(n954) );
  NANDN U1022 ( .A(n12969), .B(n954), .Z(n955) );
  ANDN U1023 ( .B(n955), .A(n12971), .Z(n956) );
  NANDN U1024 ( .A(n956), .B(n12973), .Z(n957) );
  NANDN U1025 ( .A(n12975), .B(n957), .Z(n958) );
  NAND U1026 ( .A(n5294), .B(n958), .Z(n959) );
  OR U1027 ( .A(n959), .B(n12977), .Z(n960) );
  NANDN U1028 ( .A(n12979), .B(n960), .Z(n961) );
  NAND U1029 ( .A(n9301), .B(n961), .Z(n962) );
  NAND U1030 ( .A(n12983), .B(n962), .Z(n963) );
  AND U1031 ( .A(n5293), .B(n963), .Z(n964) );
  NANDN U1032 ( .A(n12984), .B(n964), .Z(n4494) );
  ANDN U1033 ( .B(n12885), .A(n9264), .Z(n965) );
  NAND U1034 ( .A(n12888), .B(n965), .Z(n966) );
  AND U1035 ( .A(n9265), .B(n966), .Z(n967) );
  NANDN U1036 ( .A(n12891), .B(n967), .Z(n968) );
  NANDN U1037 ( .A(n12893), .B(n968), .Z(n969) );
  AND U1038 ( .A(n12895), .B(n969), .Z(n970) );
  OR U1039 ( .A(n970), .B(n12897), .Z(n971) );
  NAND U1040 ( .A(n12899), .B(n971), .Z(n972) );
  NANDN U1041 ( .A(n9266), .B(n972), .Z(n973) );
  AND U1042 ( .A(n12903), .B(n5323), .Z(n974) );
  OR U1043 ( .A(n973), .B(n12901), .Z(n975) );
  AND U1044 ( .A(n974), .B(n975), .Z(n976) );
  NOR U1045 ( .A(n976), .B(n9268), .Z(n977) );
  NAND U1046 ( .A(n9267), .B(n977), .Z(n978) );
  AND U1047 ( .A(n12910), .B(n978), .Z(n979) );
  OR U1048 ( .A(n9269), .B(n9270), .Z(n980) );
  NAND U1049 ( .A(n979), .B(n980), .Z(n981) );
  NANDN U1050 ( .A(n12913), .B(n981), .Z(n9271) );
  AND U1051 ( .A(n5259), .B(n5263), .Z(n982) );
  OR U1052 ( .A(n5260), .B(n4499), .Z(n983) );
  AND U1053 ( .A(n982), .B(n983), .Z(n984) );
  NOR U1054 ( .A(n5256), .B(n5261), .Z(n985) );
  NANDN U1055 ( .A(n984), .B(n985), .Z(n986) );
  AND U1056 ( .A(n5258), .B(n986), .Z(n987) );
  XNOR U1057 ( .A(y[1350]), .B(x[1350]), .Z(n988) );
  NAND U1058 ( .A(n987), .B(n988), .Z(n989) );
  NAND U1059 ( .A(n5257), .B(n989), .Z(n990) );
  NAND U1060 ( .A(n5255), .B(n990), .Z(n991) );
  NANDN U1061 ( .A(n13095), .B(n991), .Z(n992) );
  AND U1062 ( .A(n13097), .B(n992), .Z(n993) );
  OR U1063 ( .A(n13099), .B(n993), .Z(n994) );
  NAND U1064 ( .A(n13101), .B(n994), .Z(n995) );
  NANDN U1065 ( .A(n13102), .B(n995), .Z(n996) );
  NANDN U1066 ( .A(n9347), .B(n996), .Z(n4500) );
  NAND U1067 ( .A(n9303), .B(n9302), .Z(n997) );
  AND U1068 ( .A(n9304), .B(n997), .Z(n998) );
  NANDN U1069 ( .A(n12990), .B(n998), .Z(n999) );
  NANDN U1070 ( .A(n9305), .B(n9306), .Z(n1000) );
  AND U1071 ( .A(n12993), .B(n12997), .Z(n1001) );
  NAND U1072 ( .A(n999), .B(n1001), .Z(n1002) );
  NANDN U1073 ( .A(n1000), .B(n1002), .Z(n1003) );
  NAND U1074 ( .A(n13001), .B(n1003), .Z(n1004) );
  NANDN U1075 ( .A(n13003), .B(n1004), .Z(n1005) );
  AND U1076 ( .A(n13005), .B(n1005), .Z(n1006) );
  ANDN U1077 ( .B(n9307), .A(n1006), .Z(n1007) );
  NAND U1078 ( .A(n13007), .B(n1007), .Z(n1008) );
  ANDN U1079 ( .B(n1008), .A(n13009), .Z(n1009) );
  ANDN U1080 ( .B(n5284), .A(n1009), .Z(n1010) );
  NAND U1081 ( .A(n13010), .B(n1010), .Z(n1011) );
  ANDN U1082 ( .B(n1011), .A(n13017), .Z(n1012) );
  NANDN U1083 ( .A(n1012), .B(n13019), .Z(n1013) );
  NANDN U1084 ( .A(n13021), .B(n1013), .Z(n1014) );
  NAND U1085 ( .A(n13023), .B(n1014), .Z(n9308) );
  AND U1086 ( .A(n9372), .B(n4508), .Z(n1015) );
  NAND U1087 ( .A(n5233), .B(n4507), .Z(n1016) );
  AND U1088 ( .A(n1015), .B(n1016), .Z(n1017) );
  ANDN U1089 ( .B(n5229), .A(n1017), .Z(n1018) );
  NAND U1090 ( .A(n5232), .B(n1018), .Z(n1019) );
  ANDN U1091 ( .B(n1019), .A(n13189), .Z(n1020) );
  NAND U1092 ( .A(n1020), .B(n5230), .Z(n1021) );
  AND U1093 ( .A(n5228), .B(n1021), .Z(n1022) );
  NAND U1094 ( .A(n1022), .B(n13191), .Z(n1023) );
  AND U1095 ( .A(n13195), .B(n5227), .Z(n1024) );
  NANDN U1096 ( .A(n13193), .B(n1023), .Z(n1025) );
  NAND U1097 ( .A(n1024), .B(n1025), .Z(n1026) );
  NOR U1098 ( .A(n13197), .B(n9377), .Z(n1027) );
  NAND U1099 ( .A(n1026), .B(n1027), .Z(n1028) );
  NANDN U1100 ( .A(n13202), .B(n1028), .Z(n1029) );
  ANDN U1101 ( .B(n9376), .A(n9380), .Z(n1030) );
  OR U1102 ( .A(n1029), .B(n5226), .Z(n1031) );
  AND U1103 ( .A(n1030), .B(n1031), .Z(n4509) );
  NANDN U1104 ( .A(n9352), .B(n13119), .Z(n1032) );
  NAND U1105 ( .A(n13121), .B(n1032), .Z(n1033) );
  ANDN U1106 ( .B(n1033), .A(n9353), .Z(n1034) );
  ANDN U1107 ( .B(n9354), .A(n9355), .Z(n1035) );
  NANDN U1108 ( .A(n13123), .B(n1034), .Z(n1036) );
  NAND U1109 ( .A(n1035), .B(n1036), .Z(n1037) );
  NAND U1110 ( .A(n9358), .B(n9359), .Z(n1038) );
  NOR U1111 ( .A(n9357), .B(n9356), .Z(n1039) );
  NAND U1112 ( .A(n1037), .B(n1039), .Z(n1040) );
  NANDN U1113 ( .A(n1038), .B(n1040), .Z(n1041) );
  ANDN U1114 ( .B(n13135), .A(n9360), .Z(n1042) );
  NAND U1115 ( .A(n1041), .B(n1042), .Z(n1043) );
  NAND U1116 ( .A(n9361), .B(n1043), .Z(n1044) );
  OR U1117 ( .A(n1044), .B(n13137), .Z(n1045) );
  NANDN U1118 ( .A(n13139), .B(n1045), .Z(n1046) );
  NAND U1119 ( .A(n13141), .B(n1046), .Z(n1047) );
  ANDN U1120 ( .B(n9364), .A(n13144), .Z(n1048) );
  NANDN U1121 ( .A(n13143), .B(n1047), .Z(n1049) );
  NAND U1122 ( .A(n1048), .B(n1049), .Z(n9365) );
  NOR U1123 ( .A(n4513), .B(n4512), .Z(n1050) );
  NAND U1124 ( .A(n9404), .B(n1050), .Z(n1051) );
  ANDN U1125 ( .B(n1051), .A(n5214), .Z(n1052) );
  NOR U1126 ( .A(n9405), .B(n1052), .Z(n1053) );
  NAND U1127 ( .A(n5212), .B(n1053), .Z(n1054) );
  ANDN U1128 ( .B(n1054), .A(n5216), .Z(n1055) );
  AND U1129 ( .A(n5208), .B(n5213), .Z(n1056) );
  NANDN U1130 ( .A(n5210), .B(n1055), .Z(n1057) );
  NAND U1131 ( .A(n1056), .B(n1057), .Z(n1058) );
  NANDN U1132 ( .A(n5211), .B(n1058), .Z(n1059) );
  AND U1133 ( .A(n13274), .B(n5209), .Z(n1060) );
  NANDN U1134 ( .A(n1059), .B(n13273), .Z(n1061) );
  AND U1135 ( .A(n1060), .B(n1061), .Z(n1062) );
  OR U1136 ( .A(n13277), .B(n1062), .Z(n1063) );
  NAND U1137 ( .A(n13279), .B(n1063), .Z(n1064) );
  NANDN U1138 ( .A(n13281), .B(n1064), .Z(n1065) );
  NANDN U1139 ( .A(n13283), .B(n1065), .Z(n4515) );
  AND U1140 ( .A(n13236), .B(n5221), .Z(n9392) );
  NANDN U1141 ( .A(n13293), .B(n9416), .Z(n1066) );
  NAND U1142 ( .A(n13295), .B(n1066), .Z(n1067) );
  AND U1143 ( .A(n13296), .B(n1067), .Z(n1068) );
  AND U1144 ( .A(n13301), .B(n9417), .Z(n1069) );
  NANDN U1145 ( .A(n1068), .B(n13299), .Z(n1070) );
  AND U1146 ( .A(n1069), .B(n1070), .Z(n1071) );
  NOR U1147 ( .A(n13303), .B(n1071), .Z(n1072) );
  NAND U1148 ( .A(n9418), .B(n1072), .Z(n1073) );
  AND U1149 ( .A(n9419), .B(n1073), .Z(n1074) );
  NAND U1150 ( .A(n9420), .B(n9421), .Z(n1075) );
  NAND U1151 ( .A(n9422), .B(n1075), .Z(n1076) );
  AND U1152 ( .A(n1074), .B(n1076), .Z(n1077) );
  NAND U1153 ( .A(n1077), .B(n9423), .Z(n1078) );
  AND U1154 ( .A(n13311), .B(n1078), .Z(n1079) );
  NANDN U1155 ( .A(n5196), .B(n1079), .Z(n1080) );
  AND U1156 ( .A(n9424), .B(n13317), .Z(n1081) );
  NAND U1157 ( .A(n1080), .B(n1081), .Z(n1082) );
  NANDN U1158 ( .A(n13319), .B(n1082), .Z(n9425) );
  ANDN U1159 ( .B(n4522), .A(n13355), .Z(n1083) );
  NAND U1160 ( .A(n9433), .B(n1083), .Z(n1084) );
  NANDN U1161 ( .A(n13357), .B(n1084), .Z(n1085) );
  NAND U1162 ( .A(n13359), .B(n1085), .Z(n1086) );
  NAND U1163 ( .A(n13361), .B(n1086), .Z(n1087) );
  AND U1164 ( .A(n13363), .B(n1087), .Z(n1088) );
  NOR U1165 ( .A(n13365), .B(n1088), .Z(n1089) );
  NAND U1166 ( .A(n5172), .B(n1089), .Z(n1090) );
  AND U1167 ( .A(n13367), .B(n1090), .Z(n1091) );
  NANDN U1168 ( .A(n1091), .B(n5175), .Z(n1092) );
  NANDN U1169 ( .A(n13370), .B(n1092), .Z(n1093) );
  NAND U1170 ( .A(n13373), .B(n1093), .Z(n1094) );
  NOR U1171 ( .A(n13375), .B(n9442), .Z(n1095) );
  NANDN U1172 ( .A(n1094), .B(n5171), .Z(n1096) );
  AND U1173 ( .A(n1095), .B(n1096), .Z(n1097) );
  ANDN U1174 ( .B(n9444), .A(n1097), .Z(n1098) );
  NAND U1175 ( .A(n5170), .B(n1098), .Z(n1099) );
  ANDN U1176 ( .B(n1099), .A(n13383), .Z(n4524) );
  NAND U1177 ( .A(n9453), .B(n9454), .Z(n1100) );
  NANDN U1178 ( .A(n13413), .B(n1100), .Z(n1101) );
  AND U1179 ( .A(n9455), .B(n1101), .Z(n1102) );
  OR U1180 ( .A(n5160), .B(n5161), .Z(n1103) );
  AND U1181 ( .A(n5162), .B(n1103), .Z(n1104) );
  NANDN U1182 ( .A(n13414), .B(n1102), .Z(n1105) );
  NAND U1183 ( .A(n13416), .B(n1105), .Z(n1106) );
  AND U1184 ( .A(n1104), .B(n1106), .Z(n1107) );
  OR U1185 ( .A(n13421), .B(n1107), .Z(n1108) );
  NAND U1186 ( .A(n13423), .B(n1108), .Z(n1109) );
  NANDN U1187 ( .A(n13425), .B(n1109), .Z(n1110) );
  NAND U1188 ( .A(n9456), .B(n1110), .Z(n1111) );
  NAND U1189 ( .A(n13428), .B(n1111), .Z(n1112) );
  AND U1190 ( .A(n5159), .B(n1112), .Z(n1113) );
  NANDN U1191 ( .A(n13431), .B(n1113), .Z(n1114) );
  ANDN U1192 ( .B(n5156), .A(n13435), .Z(n1115) );
  NANDN U1193 ( .A(n13433), .B(n1114), .Z(n1116) );
  NAND U1194 ( .A(n1115), .B(n1116), .Z(n9457) );
  NAND U1195 ( .A(n9480), .B(n9479), .Z(n1117) );
  NANDN U1196 ( .A(n13497), .B(n1117), .Z(n1118) );
  NAND U1197 ( .A(n13499), .B(n1118), .Z(n1119) );
  AND U1198 ( .A(n13503), .B(n5128), .Z(n1120) );
  NANDN U1199 ( .A(n13501), .B(n1119), .Z(n1121) );
  NAND U1200 ( .A(n1120), .B(n1121), .Z(n1122) );
  ANDN U1201 ( .B(n9481), .A(n13505), .Z(n1123) );
  NAND U1202 ( .A(n1122), .B(n1123), .Z(n1124) );
  NAND U1203 ( .A(n13510), .B(n1124), .Z(n1125) );
  NANDN U1204 ( .A(n1125), .B(n9482), .Z(n1126) );
  ANDN U1205 ( .B(n1126), .A(n13513), .Z(n1127) );
  NANDN U1206 ( .A(n5124), .B(n13521), .Z(n1128) );
  ANDN U1207 ( .B(n5125), .A(n1127), .Z(n1129) );
  NAND U1208 ( .A(n13515), .B(n1129), .Z(n1130) );
  NANDN U1209 ( .A(n1128), .B(n1130), .Z(n1131) );
  AND U1210 ( .A(n5123), .B(n13522), .Z(n1132) );
  NAND U1211 ( .A(n1131), .B(n1132), .Z(n1133) );
  NAND U1212 ( .A(n13525), .B(n1133), .Z(n1134) );
  NAND U1213 ( .A(n13527), .B(n1134), .Z(n9483) );
  NAND U1214 ( .A(n4565), .B(n4564), .Z(n1135) );
  NANDN U1215 ( .A(n13558), .B(n1135), .Z(n1136) );
  AND U1216 ( .A(n13560), .B(n1136), .Z(n1137) );
  OR U1217 ( .A(n13563), .B(n1137), .Z(n1138) );
  NANDN U1218 ( .A(n13565), .B(n1138), .Z(n1139) );
  NAND U1219 ( .A(n13567), .B(n1139), .Z(n1140) );
  NANDN U1220 ( .A(n13569), .B(n1140), .Z(n1141) );
  NAND U1221 ( .A(n13571), .B(n1141), .Z(n1142) );
  ANDN U1222 ( .B(n1142), .A(n13573), .Z(n1143) );
  NANDN U1223 ( .A(n5094), .B(n1143), .Z(n1144) );
  NAND U1224 ( .A(n13575), .B(n1144), .Z(n1145) );
  ANDN U1225 ( .B(n1145), .A(n5096), .Z(n1146) );
  NAND U1226 ( .A(n1146), .B(n13578), .Z(n1147) );
  NANDN U1227 ( .A(n13581), .B(n1147), .Z(n1148) );
  ANDN U1228 ( .B(n1148), .A(n5092), .Z(n4566) );
  NANDN U1229 ( .A(n9526), .B(n9527), .Z(n1149) );
  NAND U1230 ( .A(n9528), .B(n1149), .Z(n1150) );
  AND U1231 ( .A(n13638), .B(n1150), .Z(n1151) );
  OR U1232 ( .A(n13641), .B(n1151), .Z(n1152) );
  NANDN U1233 ( .A(n9529), .B(n1152), .Z(n1153) );
  NANDN U1234 ( .A(n13647), .B(n1153), .Z(n1154) );
  NAND U1235 ( .A(n9530), .B(n1154), .Z(n1155) );
  NANDN U1236 ( .A(n13651), .B(n1155), .Z(n1156) );
  ANDN U1237 ( .B(n1156), .A(n13653), .Z(n1157) );
  NANDN U1238 ( .A(n1157), .B(n13655), .Z(n1158) );
  NANDN U1239 ( .A(n13657), .B(n1158), .Z(n1159) );
  NAND U1240 ( .A(n13659), .B(n1159), .Z(n1160) );
  NAND U1241 ( .A(n13661), .B(n1160), .Z(n1161) );
  AND U1242 ( .A(n5068), .B(n1161), .Z(n1162) );
  NANDN U1243 ( .A(n13663), .B(n1162), .Z(n1163) );
  NAND U1244 ( .A(n13665), .B(n1163), .Z(n1164) );
  NANDN U1245 ( .A(n9533), .B(n1164), .Z(n9534) );
  AND U1246 ( .A(n9540), .B(n5060), .Z(n1165) );
  NANDN U1247 ( .A(n13695), .B(n4598), .Z(n1166) );
  NAND U1248 ( .A(n1165), .B(n1166), .Z(n1167) );
  NANDN U1249 ( .A(n9538), .B(n1167), .Z(n1168) );
  AND U1250 ( .A(n5056), .B(n9541), .Z(n1169) );
  OR U1251 ( .A(n1168), .B(n5058), .Z(n1170) );
  AND U1252 ( .A(n1169), .B(n1170), .Z(n1171) );
  ANDN U1253 ( .B(n5059), .A(n1171), .Z(n1172) );
  NAND U1254 ( .A(n13707), .B(n1172), .Z(n1173) );
  AND U1255 ( .A(n5057), .B(n1173), .Z(n1174) );
  NAND U1256 ( .A(n1174), .B(n13709), .Z(n1175) );
  NANDN U1257 ( .A(n13711), .B(n1175), .Z(n1176) );
  AND U1258 ( .A(n5052), .B(n1176), .Z(n1177) );
  NAND U1259 ( .A(n1177), .B(n13713), .Z(n1178) );
  NAND U1260 ( .A(n13714), .B(n1178), .Z(n1179) );
  AND U1261 ( .A(n5053), .B(n1179), .Z(n1180) );
  OR U1262 ( .A(n13719), .B(n1180), .Z(n1181) );
  AND U1263 ( .A(n9543), .B(n1181), .Z(n4601) );
  AND U1264 ( .A(n13753), .B(n5042), .Z(n9550) );
  AND U1265 ( .A(n5024), .B(n13792), .Z(n1182) );
  NANDN U1266 ( .A(n13791), .B(n4605), .Z(n1183) );
  NAND U1267 ( .A(n1182), .B(n1183), .Z(n1184) );
  NANDN U1268 ( .A(n13799), .B(n1184), .Z(n1185) );
  NAND U1269 ( .A(n13801), .B(n1185), .Z(n1186) );
  ANDN U1270 ( .B(n1186), .A(n13803), .Z(n1187) );
  NANDN U1271 ( .A(n1187), .B(n13805), .Z(n1188) );
  NANDN U1272 ( .A(n13807), .B(n1188), .Z(n1189) );
  NAND U1273 ( .A(n13809), .B(n1189), .Z(n1190) );
  NANDN U1274 ( .A(n13810), .B(n1190), .Z(n1191) );
  AND U1275 ( .A(n5013), .B(n13813), .Z(n1192) );
  NANDN U1276 ( .A(n1191), .B(n5014), .Z(n1193) );
  AND U1277 ( .A(n1192), .B(n1193), .Z(n1194) );
  NOR U1278 ( .A(n5015), .B(n13819), .Z(n1195) );
  NANDN U1279 ( .A(n1194), .B(n1195), .Z(n1196) );
  AND U1280 ( .A(n13821), .B(n1196), .Z(n1197) );
  NAND U1281 ( .A(n1197), .B(n5012), .Z(n1198) );
  NANDN U1282 ( .A(n13823), .B(n1198), .Z(n1199) );
  AND U1283 ( .A(n13825), .B(n1199), .Z(n4607) );
  ANDN U1284 ( .B(n9641), .A(n4989), .Z(n1200) );
  NAND U1285 ( .A(n4990), .B(n1200), .Z(n1201) );
  ANDN U1286 ( .B(n1201), .A(n9642), .Z(n1202) );
  NAND U1287 ( .A(n1202), .B(n9643), .Z(n1203) );
  AND U1288 ( .A(n4987), .B(n1203), .Z(n1204) );
  NAND U1289 ( .A(n1204), .B(n4988), .Z(n1205) );
  AND U1290 ( .A(n4986), .B(n4985), .Z(n1206) );
  NAND U1291 ( .A(n1206), .B(n1205), .Z(n1207) );
  AND U1292 ( .A(n4984), .B(n1207), .Z(n1208) );
  NAND U1293 ( .A(n1208), .B(n4983), .Z(n1209) );
  AND U1294 ( .A(n9644), .B(n13932), .Z(n1210) );
  NAND U1295 ( .A(n1209), .B(n1210), .Z(n1211) );
  NANDN U1296 ( .A(n9645), .B(n1211), .Z(n1212) );
  OR U1297 ( .A(n1212), .B(n13935), .Z(n1213) );
  NAND U1298 ( .A(n13937), .B(n1213), .Z(n1214) );
  NANDN U1299 ( .A(n13939), .B(n1214), .Z(n1215) );
  NAND U1300 ( .A(n13941), .B(n1215), .Z(n9650) );
  AND U1301 ( .A(n13971), .B(n9662), .Z(n1216) );
  NANDN U1302 ( .A(n4641), .B(n4640), .Z(n1217) );
  NAND U1303 ( .A(n1216), .B(n1217), .Z(n1218) );
  ANDN U1304 ( .B(n9664), .A(n13973), .Z(n1219) );
  NAND U1305 ( .A(n1218), .B(n1219), .Z(n1220) );
  NANDN U1306 ( .A(n13975), .B(n1220), .Z(n1221) );
  NAND U1307 ( .A(n13977), .B(n1221), .Z(n1222) );
  NANDN U1308 ( .A(n13979), .B(n1222), .Z(n1223) );
  ANDN U1309 ( .B(n1223), .A(n13981), .Z(n1224) );
  ANDN U1310 ( .B(n4961), .A(n13985), .Z(n1225) );
  NANDN U1311 ( .A(n1224), .B(n13983), .Z(n1226) );
  AND U1312 ( .A(n1225), .B(n1226), .Z(n1227) );
  NOR U1313 ( .A(n13987), .B(n4960), .Z(n1228) );
  NANDN U1314 ( .A(n1227), .B(n1228), .Z(n1229) );
  AND U1315 ( .A(n4962), .B(n1229), .Z(n1230) );
  NAND U1316 ( .A(n4958), .B(n1230), .Z(n4642) );
  NAND U1317 ( .A(n9671), .B(n9670), .Z(n1231) );
  ANDN U1318 ( .B(n1231), .A(n9672), .Z(n1232) );
  ANDN U1319 ( .B(n9673), .A(n9674), .Z(n1233) );
  NANDN U1320 ( .A(n13999), .B(n1232), .Z(n1234) );
  NAND U1321 ( .A(n1233), .B(n1234), .Z(n1235) );
  AND U1322 ( .A(n4954), .B(n4953), .Z(n1236) );
  NAND U1323 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1324 ( .A(n4952), .B(n1237), .Z(n1238) );
  NAND U1325 ( .A(n1238), .B(n4951), .Z(n1239) );
  AND U1326 ( .A(n4950), .B(n4949), .Z(n1240) );
  NAND U1327 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U1328 ( .A(n9676), .B(n1241), .Z(n1242) );
  NAND U1329 ( .A(n1242), .B(n9675), .Z(n1243) );
  NOR U1330 ( .A(n9677), .B(n14014), .Z(n1244) );
  NAND U1331 ( .A(n1243), .B(n1244), .Z(n1245) );
  NAND U1332 ( .A(n9678), .B(n1245), .Z(n1246) );
  OR U1333 ( .A(n1246), .B(n14017), .Z(n1247) );
  NAND U1334 ( .A(n14019), .B(n1247), .Z(n1248) );
  NAND U1335 ( .A(n14021), .B(n1248), .Z(n9683) );
  NANDN U1336 ( .A(n4650), .B(n4649), .Z(n1249) );
  NAND U1337 ( .A(n14069), .B(n1249), .Z(n1250) );
  ANDN U1338 ( .B(n1250), .A(n14075), .Z(n1251) );
  NAND U1339 ( .A(n1251), .B(n9719), .Z(n1252) );
  NAND U1340 ( .A(n14077), .B(n1252), .Z(n1253) );
  ANDN U1341 ( .B(n1253), .A(n14079), .Z(n1254) );
  OR U1342 ( .A(n14081), .B(n1254), .Z(n1255) );
  AND U1343 ( .A(n14083), .B(n1255), .Z(n1256) );
  NOR U1344 ( .A(n14085), .B(n1256), .Z(n1257) );
  NAND U1345 ( .A(n4923), .B(n1257), .Z(n1258) );
  AND U1346 ( .A(n14087), .B(n1258), .Z(n1259) );
  NAND U1347 ( .A(n1259), .B(n4922), .Z(n1260) );
  AND U1348 ( .A(n4924), .B(n1260), .Z(n1261) );
  NANDN U1349 ( .A(n4919), .B(n1261), .Z(n4651) );
  ANDN U1350 ( .B(n9747), .A(n9748), .Z(n1262) );
  NAND U1351 ( .A(n14099), .B(n1262), .Z(n1263) );
  NAND U1352 ( .A(n9749), .B(n1263), .Z(n1264) );
  NOR U1353 ( .A(n9752), .B(n9751), .Z(n1265) );
  NANDN U1354 ( .A(n1264), .B(n9750), .Z(n1266) );
  AND U1355 ( .A(n1265), .B(n1266), .Z(n1267) );
  ANDN U1356 ( .B(n9753), .A(n1267), .Z(n1268) );
  NAND U1357 ( .A(n9754), .B(n1268), .Z(n1269) );
  ANDN U1358 ( .B(n1269), .A(n9755), .Z(n1270) );
  AND U1359 ( .A(n4916), .B(n4915), .Z(n1271) );
  NANDN U1360 ( .A(n9756), .B(n1270), .Z(n1272) );
  NAND U1361 ( .A(n1271), .B(n1272), .Z(n1273) );
  ANDN U1362 ( .B(n1273), .A(n9757), .Z(n1274) );
  NOR U1363 ( .A(n14116), .B(n4914), .Z(n1275) );
  NANDN U1364 ( .A(n14115), .B(n1274), .Z(n1276) );
  NAND U1365 ( .A(n1275), .B(n1276), .Z(n1277) );
  NAND U1366 ( .A(n14118), .B(n1277), .Z(n1278) );
  NANDN U1367 ( .A(n14121), .B(n1278), .Z(n9758) );
  NAND U1368 ( .A(n4653), .B(n14151), .Z(n1279) );
  ANDN U1369 ( .B(n1279), .A(n14152), .Z(n1280) );
  NANDN U1370 ( .A(n1280), .B(n14155), .Z(n1281) );
  NANDN U1371 ( .A(n14156), .B(n1281), .Z(n1282) );
  NAND U1372 ( .A(n14159), .B(n1282), .Z(n1283) );
  AND U1373 ( .A(n4900), .B(n14163), .Z(n1284) );
  NANDN U1374 ( .A(n14161), .B(n1283), .Z(n1285) );
  NAND U1375 ( .A(n1284), .B(n1285), .Z(n1286) );
  ANDN U1376 ( .B(n9805), .A(n14165), .Z(n1287) );
  NAND U1377 ( .A(n1286), .B(n1287), .Z(n1288) );
  NANDN U1378 ( .A(n4898), .B(n1288), .Z(n1289) );
  ANDN U1379 ( .B(n9811), .A(n9804), .Z(n1290) );
  NANDN U1380 ( .A(n1289), .B(n4901), .Z(n1291) );
  AND U1381 ( .A(n1290), .B(n1291), .Z(n1292) );
  NANDN U1382 ( .A(n1292), .B(n14174), .Z(n1293) );
  NAND U1383 ( .A(n14177), .B(n1293), .Z(n1294) );
  NAND U1384 ( .A(n14179), .B(n1294), .Z(n4656) );
  NANDN U1385 ( .A(y[1834]), .B(x[1834]), .Z(n1295) );
  AND U1386 ( .A(n4879), .B(n1295), .Z(n1296) );
  NAND U1387 ( .A(n9832), .B(n9831), .Z(n1297) );
  AND U1388 ( .A(n9833), .B(n1297), .Z(n1298) );
  NAND U1389 ( .A(n1298), .B(n9834), .Z(n1299) );
  NAND U1390 ( .A(n4885), .B(n4884), .Z(n1300) );
  AND U1391 ( .A(n4887), .B(n4886), .Z(n1301) );
  NAND U1392 ( .A(n1299), .B(n1301), .Z(n1302) );
  NANDN U1393 ( .A(n1300), .B(n1302), .Z(n1303) );
  AND U1394 ( .A(n4882), .B(n4883), .Z(n1304) );
  NAND U1395 ( .A(n1304), .B(n1303), .Z(n1305) );
  AND U1396 ( .A(n9835), .B(n1305), .Z(n1306) );
  NANDN U1397 ( .A(n14216), .B(n1306), .Z(n1307) );
  ANDN U1398 ( .B(n14218), .A(n9836), .Z(n1308) );
  NAND U1399 ( .A(n1307), .B(n1308), .Z(n1309) );
  NAND U1400 ( .A(n14221), .B(n1309), .Z(n1310) );
  AND U1401 ( .A(n14225), .B(n14222), .Z(n1311) );
  NAND U1402 ( .A(n1310), .B(n1311), .Z(n1312) );
  NAND U1403 ( .A(n1296), .B(n1312), .Z(n9837) );
  NANDN U1404 ( .A(n4664), .B(n14307), .Z(n1313) );
  NANDN U1405 ( .A(n4665), .B(n1313), .Z(n1314) );
  NANDN U1406 ( .A(n14311), .B(n1314), .Z(n1315) );
  NAND U1407 ( .A(n14313), .B(n1315), .Z(n1316) );
  NANDN U1408 ( .A(n14315), .B(n1316), .Z(n1317) );
  ANDN U1409 ( .B(n1317), .A(n14317), .Z(n1318) );
  ANDN U1410 ( .B(n14319), .A(n1318), .Z(n1319) );
  NAND U1411 ( .A(n4843), .B(n1319), .Z(n1320) );
  ANDN U1412 ( .B(n1320), .A(n4842), .Z(n1321) );
  NAND U1413 ( .A(n1321), .B(n9912), .Z(n1322) );
  AND U1414 ( .A(n14327), .B(n1322), .Z(n1323) );
  NAND U1415 ( .A(n1323), .B(n4844), .Z(n1324) );
  ANDN U1416 ( .B(n4841), .A(n14329), .Z(n1325) );
  NAND U1417 ( .A(n1324), .B(n1325), .Z(n1326) );
  NAND U1418 ( .A(n14331), .B(n1326), .Z(n1327) );
  NAND U1419 ( .A(n14333), .B(n1327), .Z(n4666) );
  NANDN U1420 ( .A(n4669), .B(n4670), .Z(n1328) );
  NAND U1421 ( .A(n14387), .B(n1328), .Z(n1329) );
  AND U1422 ( .A(n14389), .B(n1329), .Z(n1330) );
  OR U1423 ( .A(n14391), .B(n1330), .Z(n1331) );
  AND U1424 ( .A(n14393), .B(n1331), .Z(n1332) );
  ANDN U1425 ( .B(n9974), .A(n1332), .Z(n1333) );
  NAND U1426 ( .A(n14394), .B(n1333), .Z(n1334) );
  ANDN U1427 ( .B(n1334), .A(n14396), .Z(n1335) );
  NAND U1428 ( .A(n9975), .B(n1335), .Z(n1336) );
  ANDN U1429 ( .B(n1336), .A(n9973), .Z(n1337) );
  NANDN U1430 ( .A(n4819), .B(n1337), .Z(n1338) );
  AND U1431 ( .A(n4818), .B(n9976), .Z(n1339) );
  NAND U1432 ( .A(n1338), .B(n1339), .Z(n1340) );
  NAND U1433 ( .A(n14407), .B(n1340), .Z(n1341) );
  OR U1434 ( .A(n4820), .B(n1341), .Z(n1342) );
  ANDN U1435 ( .B(n1342), .A(n14409), .Z(n4672) );
  NAND U1436 ( .A(n4678), .B(n4677), .Z(n1343) );
  NAND U1437 ( .A(n4679), .B(n1343), .Z(n1344) );
  AND U1438 ( .A(n14490), .B(n1344), .Z(n1345) );
  OR U1439 ( .A(n14493), .B(n1345), .Z(n1346) );
  NANDN U1440 ( .A(n14495), .B(n1346), .Z(n1347) );
  NAND U1441 ( .A(n14497), .B(n1347), .Z(n1348) );
  NAND U1442 ( .A(n14499), .B(n1348), .Z(n1349) );
  NAND U1443 ( .A(n14500), .B(n1349), .Z(n1350) );
  AND U1444 ( .A(n14503), .B(n1350), .Z(n1351) );
  NOR U1445 ( .A(n10075), .B(n1351), .Z(n1352) );
  NANDN U1446 ( .A(n10083), .B(n1352), .Z(n1353) );
  AND U1447 ( .A(n14507), .B(n1353), .Z(n1354) );
  NANDN U1448 ( .A(n1354), .B(n14509), .Z(n1355) );
  NAND U1449 ( .A(n14515), .B(n1355), .Z(n1356) );
  NANDN U1450 ( .A(n10091), .B(n1356), .Z(n4682) );
  ANDN U1451 ( .B(n10120), .A(n10121), .Z(n1357) );
  NAND U1452 ( .A(n14546), .B(n1357), .Z(n1358) );
  NAND U1453 ( .A(n14549), .B(n1358), .Z(n1359) );
  NANDN U1454 ( .A(n14550), .B(n1359), .Z(n1360) );
  NAND U1455 ( .A(n14552), .B(n1360), .Z(n1361) );
  ANDN U1456 ( .B(n1361), .A(n14555), .Z(n1362) );
  NANDN U1457 ( .A(n1362), .B(n14557), .Z(n1363) );
  NAND U1458 ( .A(n10126), .B(n1363), .Z(n1364) );
  NAND U1459 ( .A(n14561), .B(n1364), .Z(n1365) );
  AND U1460 ( .A(n4767), .B(n14565), .Z(n1366) );
  NANDN U1461 ( .A(n14563), .B(n1365), .Z(n1367) );
  NAND U1462 ( .A(n1366), .B(n1367), .Z(n1368) );
  AND U1463 ( .A(n4766), .B(n14566), .Z(n1369) );
  NAND U1464 ( .A(n1368), .B(n1369), .Z(n1370) );
  NAND U1465 ( .A(n10127), .B(n1370), .Z(n1371) );
  NANDN U1466 ( .A(n10128), .B(n1371), .Z(n10129) );
  NOR U1467 ( .A(n4697), .B(n4754), .Z(n1372) );
  NAND U1468 ( .A(n4698), .B(n1372), .Z(n1373) );
  NANDN U1469 ( .A(n14608), .B(n1373), .Z(n1374) );
  NAND U1470 ( .A(n14610), .B(n1374), .Z(n1375) );
  NAND U1471 ( .A(n14613), .B(n1375), .Z(n1376) );
  AND U1472 ( .A(n10174), .B(n1376), .Z(n1377) );
  ANDN U1473 ( .B(n1377), .A(n4751), .Z(n1378) );
  AND U1474 ( .A(n14622), .B(n10175), .Z(n1379) );
  OR U1475 ( .A(n1378), .B(n4750), .Z(n1380) );
  AND U1476 ( .A(n1379), .B(n1380), .Z(n1381) );
  NANDN U1477 ( .A(n1381), .B(n14625), .Z(n1382) );
  NAND U1478 ( .A(n10143), .B(n1382), .Z(n1383) );
  NAND U1479 ( .A(n10145), .B(n1383), .Z(n1384) );
  ANDN U1480 ( .B(n10142), .A(n10146), .Z(n1385) );
  NAND U1481 ( .A(n1384), .B(n1385), .Z(n1386) );
  NANDN U1482 ( .A(n10144), .B(n1386), .Z(n4706) );
  ANDN U1483 ( .B(n4748), .A(n14641), .Z(n1387) );
  OR U1484 ( .A(n10148), .B(n10149), .Z(n1388) );
  NAND U1485 ( .A(n1387), .B(n1388), .Z(n1389) );
  NOR U1486 ( .A(n10150), .B(n14643), .Z(n1390) );
  NAND U1487 ( .A(n1389), .B(n1390), .Z(n1391) );
  NAND U1488 ( .A(n14645), .B(n1391), .Z(n1392) );
  AND U1489 ( .A(n4747), .B(n4746), .Z(n1393) );
  NAND U1490 ( .A(n1392), .B(n1393), .Z(n1394) );
  NAND U1491 ( .A(n10171), .B(n1394), .Z(n1395) );
  NANDN U1492 ( .A(n10153), .B(n1395), .Z(n1396) );
  NOR U1493 ( .A(n10172), .B(n4743), .Z(n1397) );
  OR U1494 ( .A(n1396), .B(n10170), .Z(n1398) );
  AND U1495 ( .A(n1397), .B(n1398), .Z(n1399) );
  NANDN U1496 ( .A(n1399), .B(n10154), .Z(n1400) );
  ANDN U1497 ( .B(n1400), .A(n10155), .Z(n1401) );
  ANDN U1498 ( .B(n4742), .A(n4741), .Z(n1402) );
  NANDN U1499 ( .A(n10156), .B(n1401), .Z(n1403) );
  AND U1500 ( .A(n1402), .B(n1403), .Z(n10157) );
  AND U1501 ( .A(n4729), .B(n3195), .Z(n1404) );
  NANDN U1502 ( .A(n4713), .B(n4712), .Z(n1405) );
  AND U1503 ( .A(n1404), .B(n1405), .Z(n1406) );
  ANDN U1504 ( .B(n4731), .A(n1406), .Z(n1407) );
  NAND U1505 ( .A(n10164), .B(n1407), .Z(n1408) );
  ANDN U1506 ( .B(n1408), .A(n4728), .Z(n1409) );
  AND U1507 ( .A(n10163), .B(n4724), .Z(n1410) );
  NANDN U1508 ( .A(n4727), .B(n1409), .Z(n1411) );
  NAND U1509 ( .A(n1410), .B(n1411), .Z(n1412) );
  AND U1510 ( .A(n4726), .B(n1412), .Z(n1413) );
  XNOR U1511 ( .A(y[2031]), .B(x[2031]), .Z(n1414) );
  AND U1512 ( .A(n1413), .B(n1414), .Z(n1415) );
  NANDN U1513 ( .A(n1415), .B(n4725), .Z(n1416) );
  AND U1514 ( .A(n14690), .B(n1416), .Z(n1417) );
  OR U1515 ( .A(n14691), .B(n1417), .Z(n1418) );
  NANDN U1516 ( .A(n10165), .B(n1418), .Z(n1419) );
  NAND U1517 ( .A(n14693), .B(n1419), .Z(n4720) );
  NANDN U1518 ( .A(y[2041]), .B(x[2041]), .Z(n1420) );
  AND U1519 ( .A(n14701), .B(n1420), .Z(n14700) );
  AND U1520 ( .A(n8214), .B(n8216), .Z(n1421) );
  NAND U1521 ( .A(n8215), .B(n1421), .Z(n1422) );
  ANDN U1522 ( .B(n1422), .A(n8217), .Z(n1423) );
  NANDN U1523 ( .A(n8218), .B(n1423), .Z(n1424) );
  NAND U1524 ( .A(n8219), .B(n1424), .Z(n1425) );
  NANDN U1525 ( .A(x[646]), .B(n1425), .Z(n1426) );
  ANDN U1526 ( .B(n1426), .A(n8220), .Z(n1427) );
  XNOR U1527 ( .A(n1425), .B(x[646]), .Z(n1428) );
  NAND U1528 ( .A(n1428), .B(y[646]), .Z(n1429) );
  AND U1529 ( .A(n1427), .B(n1429), .Z(n1430) );
  NANDN U1530 ( .A(n1430), .B(n11476), .Z(n1431) );
  ANDN U1531 ( .B(n1431), .A(n11479), .Z(n1432) );
  NANDN U1532 ( .A(n1432), .B(n11481), .Z(n1433) );
  NANDN U1533 ( .A(n11483), .B(n1433), .Z(n1434) );
  NAND U1534 ( .A(n11485), .B(n1434), .Z(n8221) );
  NANDN U1535 ( .A(n4322), .B(n11631), .Z(n1435) );
  NAND U1536 ( .A(n11632), .B(n1435), .Z(n1436) );
  NANDN U1537 ( .A(n11635), .B(n1436), .Z(n1437) );
  NAND U1538 ( .A(n11637), .B(n1437), .Z(n1438) );
  NANDN U1539 ( .A(n11639), .B(n1438), .Z(n1439) );
  AND U1540 ( .A(n11641), .B(n1439), .Z(n1440) );
  NANDN U1541 ( .A(n1440), .B(n11643), .Z(n1441) );
  AND U1542 ( .A(n11644), .B(n1441), .Z(n1442) );
  OR U1543 ( .A(n11647), .B(n1442), .Z(n1443) );
  NAND U1544 ( .A(n11649), .B(n1443), .Z(n1444) );
  NANDN U1545 ( .A(n11651), .B(n1444), .Z(n4325) );
  NAND U1546 ( .A(n4330), .B(n11697), .Z(n1445) );
  NAND U1547 ( .A(n11699), .B(n1445), .Z(n1446) );
  NAND U1548 ( .A(n11701), .B(n1446), .Z(n1447) );
  NAND U1549 ( .A(n11703), .B(n1447), .Z(n1448) );
  NAND U1550 ( .A(n11704), .B(n1448), .Z(n1449) );
  AND U1551 ( .A(n11707), .B(n1449), .Z(n1450) );
  OR U1552 ( .A(n1450), .B(n5664), .Z(n1451) );
  NAND U1553 ( .A(n8553), .B(n1451), .Z(n1452) );
  AND U1554 ( .A(n11713), .B(n1452), .Z(n1453) );
  NANDN U1555 ( .A(n1453), .B(n11715), .Z(n1454) );
  NAND U1556 ( .A(n11716), .B(n1454), .Z(n1455) );
  NANDN U1557 ( .A(n11719), .B(n1455), .Z(n1456) );
  NAND U1558 ( .A(n11721), .B(n1456), .Z(n4331) );
  NANDN U1559 ( .A(n4384), .B(n4383), .Z(n1457) );
  AND U1560 ( .A(n11839), .B(n1457), .Z(n1458) );
  NOR U1561 ( .A(n11841), .B(n1458), .Z(n1459) );
  NAND U1562 ( .A(n5635), .B(n1459), .Z(n1460) );
  NAND U1563 ( .A(n11842), .B(n1460), .Z(n1461) );
  ANDN U1564 ( .B(n5634), .A(n8734), .Z(n1462) );
  NANDN U1565 ( .A(n1461), .B(n5632), .Z(n1463) );
  AND U1566 ( .A(n1462), .B(n1463), .Z(n1464) );
  ANDN U1567 ( .B(n5633), .A(n1464), .Z(n1465) );
  NAND U1568 ( .A(n11851), .B(n1465), .Z(n1466) );
  ANDN U1569 ( .B(n1466), .A(n11853), .Z(n1467) );
  NAND U1570 ( .A(n1467), .B(n8733), .Z(n1468) );
  NAND U1571 ( .A(n11855), .B(n1468), .Z(n1469) );
  ANDN U1572 ( .B(n1469), .A(n11857), .Z(n1470) );
  NANDN U1573 ( .A(n1470), .B(n11859), .Z(n1471) );
  NANDN U1574 ( .A(n11861), .B(n1471), .Z(n1472) );
  NAND U1575 ( .A(n11863), .B(n1472), .Z(n1473) );
  NANDN U1576 ( .A(n11865), .B(n1473), .Z(n4385) );
  AND U1577 ( .A(n5599), .B(n11925), .Z(n1474) );
  NANDN U1578 ( .A(n4388), .B(n4387), .Z(n1475) );
  AND U1579 ( .A(n1474), .B(n1475), .Z(n1476) );
  OR U1580 ( .A(n1476), .B(n11927), .Z(n1477) );
  NAND U1581 ( .A(n11929), .B(n1477), .Z(n1478) );
  NANDN U1582 ( .A(n11931), .B(n1478), .Z(n1479) );
  NAND U1583 ( .A(n11933), .B(n1479), .Z(n1480) );
  NANDN U1584 ( .A(n11935), .B(n1480), .Z(n1481) );
  AND U1585 ( .A(n11937), .B(n1481), .Z(n1482) );
  NOR U1586 ( .A(n11939), .B(n5589), .Z(n1483) );
  NANDN U1587 ( .A(n1482), .B(n1483), .Z(n1484) );
  AND U1588 ( .A(n11941), .B(n1484), .Z(n1485) );
  OR U1589 ( .A(n5593), .B(n1485), .Z(n1486) );
  AND U1590 ( .A(n5585), .B(n1486), .Z(n1487) );
  NOR U1591 ( .A(n5590), .B(n5583), .Z(n1488) );
  NANDN U1592 ( .A(n1487), .B(n1488), .Z(n1489) );
  AND U1593 ( .A(n5587), .B(n1489), .Z(n1490) );
  NAND U1594 ( .A(n5581), .B(n1490), .Z(n4392) );
  NOR U1595 ( .A(n11990), .B(n5568), .Z(n1491) );
  NAND U1596 ( .A(n4395), .B(n1491), .Z(n1492) );
  AND U1597 ( .A(n11992), .B(n1492), .Z(n1493) );
  NOR U1598 ( .A(n11995), .B(n1493), .Z(n1494) );
  NAND U1599 ( .A(n5566), .B(n1494), .Z(n1495) );
  ANDN U1600 ( .B(n1495), .A(n11997), .Z(n1496) );
  ANDN U1601 ( .B(n5567), .A(n12002), .Z(n1497) );
  NANDN U1602 ( .A(n5565), .B(n1496), .Z(n1498) );
  NAND U1603 ( .A(n1497), .B(n1498), .Z(n1499) );
  AND U1604 ( .A(n5564), .B(n12004), .Z(n1500) );
  NAND U1605 ( .A(n1499), .B(n1500), .Z(n1501) );
  NANDN U1606 ( .A(n12007), .B(n1501), .Z(n4396) );
  NAND U1607 ( .A(n4407), .B(n4406), .Z(n1502) );
  NAND U1608 ( .A(n4408), .B(n1502), .Z(n1503) );
  AND U1609 ( .A(n12061), .B(n1503), .Z(n1504) );
  ANDN U1610 ( .B(n8885), .A(n1504), .Z(n1505) );
  NAND U1611 ( .A(n8883), .B(n1505), .Z(n1506) );
  ANDN U1612 ( .B(n1506), .A(n5546), .Z(n1507) );
  NAND U1613 ( .A(n5545), .B(n1507), .Z(n1508) );
  ANDN U1614 ( .B(n1508), .A(n8884), .Z(n1509) );
  NANDN U1615 ( .A(n5542), .B(n1509), .Z(n1510) );
  NOR U1616 ( .A(n5544), .B(n12073), .Z(n1511) );
  NAND U1617 ( .A(n1510), .B(n1511), .Z(n1512) );
  NAND U1618 ( .A(n12074), .B(n1512), .Z(n1513) );
  NANDN U1619 ( .A(n1513), .B(n5543), .Z(n1514) );
  NANDN U1620 ( .A(n12077), .B(n1514), .Z(n1515) );
  NAND U1621 ( .A(n12079), .B(n1515), .Z(n1516) );
  NANDN U1622 ( .A(n12081), .B(n1516), .Z(n4409) );
  NAND U1623 ( .A(n8766), .B(n11872), .Z(n1517) );
  NANDN U1624 ( .A(n8767), .B(n1517), .Z(n1518) );
  AND U1625 ( .A(n8768), .B(n1518), .Z(n1519) );
  AND U1626 ( .A(n11883), .B(n11878), .Z(n1520) );
  ANDN U1627 ( .B(n5624), .A(n1519), .Z(n1521) );
  NAND U1628 ( .A(n5625), .B(n1521), .Z(n1522) );
  AND U1629 ( .A(n1520), .B(n1522), .Z(n1523) );
  ANDN U1630 ( .B(n5623), .A(n1523), .Z(n1524) );
  NAND U1631 ( .A(n11884), .B(n1524), .Z(n1525) );
  ANDN U1632 ( .B(n1525), .A(n11887), .Z(n1526) );
  NOR U1633 ( .A(n11891), .B(n8769), .Z(n1527) );
  NANDN U1634 ( .A(n1526), .B(n11889), .Z(n1528) );
  AND U1635 ( .A(n1527), .B(n1528), .Z(n1529) );
  ANDN U1636 ( .B(n11893), .A(n1529), .Z(n1530) );
  NAND U1637 ( .A(n8770), .B(n1530), .Z(n1531) );
  ANDN U1638 ( .B(n1531), .A(n8771), .Z(n1532) );
  ANDN U1639 ( .B(n8773), .A(n8774), .Z(n1533) );
  NANDN U1640 ( .A(n8772), .B(n1532), .Z(n1534) );
  NAND U1641 ( .A(n1533), .B(n1534), .Z(n8775) );
  NAND U1642 ( .A(n4413), .B(n5526), .Z(n1535) );
  AND U1643 ( .A(n5528), .B(n1535), .Z(n1536) );
  NANDN U1644 ( .A(n12145), .B(n1536), .Z(n1537) );
  AND U1645 ( .A(n5527), .B(n12146), .Z(n1538) );
  NAND U1646 ( .A(n1537), .B(n1538), .Z(n1539) );
  NANDN U1647 ( .A(n12149), .B(n1539), .Z(n1540) );
  NAND U1648 ( .A(n12151), .B(n1540), .Z(n1541) );
  NANDN U1649 ( .A(n12153), .B(n1541), .Z(n1542) );
  AND U1650 ( .A(n12155), .B(n1542), .Z(n1543) );
  OR U1651 ( .A(n12157), .B(n1543), .Z(n1544) );
  NAND U1652 ( .A(n12159), .B(n1544), .Z(n1545) );
  NAND U1653 ( .A(n12161), .B(n1545), .Z(n1546) );
  NANDN U1654 ( .A(n12163), .B(n1546), .Z(n1547) );
  NAND U1655 ( .A(n12165), .B(n1547), .Z(n1548) );
  ANDN U1656 ( .B(n1548), .A(n12167), .Z(n1549) );
  NANDN U1657 ( .A(n1549), .B(n12169), .Z(n1550) );
  NAND U1658 ( .A(n12170), .B(n1550), .Z(n1551) );
  NAND U1659 ( .A(n12173), .B(n1551), .Z(n1552) );
  NANDN U1660 ( .A(n5522), .B(n1552), .Z(n4414) );
  NAND U1661 ( .A(n8863), .B(n8862), .Z(n1553) );
  NAND U1662 ( .A(n8866), .B(n1553), .Z(n1554) );
  ANDN U1663 ( .B(n1554), .A(n12023), .Z(n1555) );
  AND U1664 ( .A(n12025), .B(n8868), .Z(n1556) );
  NANDN U1665 ( .A(n8867), .B(n1555), .Z(n1557) );
  NAND U1666 ( .A(n1556), .B(n1557), .Z(n1558) );
  NANDN U1667 ( .A(n12026), .B(n1558), .Z(n1559) );
  NAND U1668 ( .A(n12028), .B(n1559), .Z(n1560) );
  ANDN U1669 ( .B(n1560), .A(n12031), .Z(n1561) );
  NANDN U1670 ( .A(n1561), .B(n12033), .Z(n1562) );
  NANDN U1671 ( .A(n12035), .B(n1562), .Z(n1563) );
  NAND U1672 ( .A(n12037), .B(n1563), .Z(n1564) );
  AND U1673 ( .A(n5555), .B(n12038), .Z(n1565) );
  NAND U1674 ( .A(n1564), .B(n1565), .Z(n1566) );
  NAND U1675 ( .A(n12041), .B(n1566), .Z(n8873) );
  NANDN U1676 ( .A(n4422), .B(n4421), .Z(n1567) );
  ANDN U1677 ( .B(n1567), .A(n12252), .Z(n1568) );
  ANDN U1678 ( .B(n5503), .A(n1568), .Z(n1569) );
  NAND U1679 ( .A(n12254), .B(n1569), .Z(n1570) );
  NAND U1680 ( .A(n12257), .B(n1570), .Z(n1571) );
  NOR U1681 ( .A(n5504), .B(n9011), .Z(n1572) );
  NANDN U1682 ( .A(n1571), .B(n9010), .Z(n1573) );
  AND U1683 ( .A(n1572), .B(n1573), .Z(n1574) );
  NOR U1684 ( .A(n9014), .B(n1574), .Z(n1575) );
  NAND U1685 ( .A(n9009), .B(n1575), .Z(n1576) );
  AND U1686 ( .A(n9016), .B(n1576), .Z(n1577) );
  NAND U1687 ( .A(n9012), .B(n1577), .Z(n1578) );
  NAND U1688 ( .A(n12269), .B(n1578), .Z(n1579) );
  NANDN U1689 ( .A(n12271), .B(n1579), .Z(n1580) );
  AND U1690 ( .A(n12273), .B(n1580), .Z(n4423) );
  ANDN U1691 ( .B(n8896), .A(n8897), .Z(n1581) );
  NAND U1692 ( .A(n1581), .B(n12097), .Z(n1582) );
  AND U1693 ( .A(n5534), .B(n1582), .Z(n1583) );
  NANDN U1694 ( .A(n12099), .B(n1583), .Z(n1584) );
  NOR U1695 ( .A(n8899), .B(n8898), .Z(n1585) );
  NAND U1696 ( .A(n1584), .B(n1585), .Z(n1586) );
  NAND U1697 ( .A(n8900), .B(n1586), .Z(n1587) );
  AND U1698 ( .A(n8901), .B(n8902), .Z(n1588) );
  NAND U1699 ( .A(n1587), .B(n1588), .Z(n1589) );
  NANDN U1700 ( .A(n8903), .B(n1589), .Z(n1590) );
  OR U1701 ( .A(n12107), .B(n1590), .Z(n1591) );
  AND U1702 ( .A(n8904), .B(n1591), .Z(n1592) );
  NOR U1703 ( .A(n8907), .B(n8906), .Z(n1593) );
  NAND U1704 ( .A(n1592), .B(n8905), .Z(n1594) );
  AND U1705 ( .A(n1593), .B(n1594), .Z(n1595) );
  ANDN U1706 ( .B(n8908), .A(n1595), .Z(n1596) );
  NAND U1707 ( .A(n8909), .B(n1596), .Z(n1597) );
  ANDN U1708 ( .B(n1597), .A(n8910), .Z(n1598) );
  NANDN U1709 ( .A(n8911), .B(n1598), .Z(n8912) );
  NAND U1710 ( .A(n4427), .B(n4426), .Z(n1599) );
  AND U1711 ( .A(n9039), .B(n1599), .Z(n1600) );
  NAND U1712 ( .A(n1600), .B(n5485), .Z(n1601) );
  ANDN U1713 ( .B(n5482), .A(n9042), .Z(n1602) );
  NAND U1714 ( .A(n1601), .B(n1602), .Z(n1603) );
  NAND U1715 ( .A(n12333), .B(n1603), .Z(n1604) );
  NAND U1716 ( .A(n12334), .B(n1604), .Z(n1605) );
  NAND U1717 ( .A(n12337), .B(n1605), .Z(n1606) );
  AND U1718 ( .A(n12339), .B(n1606), .Z(n1607) );
  NANDN U1719 ( .A(n1607), .B(n12341), .Z(n1608) );
  NANDN U1720 ( .A(n12343), .B(n1608), .Z(n1609) );
  NAND U1721 ( .A(n12345), .B(n1609), .Z(n1610) );
  NOR U1722 ( .A(n5480), .B(n12346), .Z(n1611) );
  NAND U1723 ( .A(n1610), .B(n1611), .Z(n1612) );
  NAND U1724 ( .A(n12352), .B(n1612), .Z(n1613) );
  NANDN U1725 ( .A(n1613), .B(n12349), .Z(n1614) );
  AND U1726 ( .A(n5479), .B(n1614), .Z(n4428) );
  NANDN U1727 ( .A(n8976), .B(n8975), .Z(n1615) );
  NAND U1728 ( .A(n8979), .B(n1615), .Z(n1616) );
  NANDN U1729 ( .A(n8980), .B(n1616), .Z(n1617) );
  ANDN U1730 ( .B(n8982), .A(n8983), .Z(n1618) );
  NANDN U1731 ( .A(n1617), .B(n8981), .Z(n1619) );
  AND U1732 ( .A(n1618), .B(n1619), .Z(n1620) );
  NANDN U1733 ( .A(n1620), .B(n12199), .Z(n1621) );
  NAND U1734 ( .A(n12200), .B(n1621), .Z(n1622) );
  NAND U1735 ( .A(n12203), .B(n1622), .Z(n1623) );
  NAND U1736 ( .A(n12205), .B(n1623), .Z(n1624) );
  NAND U1737 ( .A(n12207), .B(n1624), .Z(n1625) );
  AND U1738 ( .A(n8988), .B(n1625), .Z(n1626) );
  NAND U1739 ( .A(n1626), .B(n12209), .Z(n1627) );
  AND U1740 ( .A(n8989), .B(n12216), .Z(n1628) );
  NANDN U1741 ( .A(n12211), .B(n1627), .Z(n1629) );
  NAND U1742 ( .A(n1628), .B(n1629), .Z(n1630) );
  AND U1743 ( .A(n12221), .B(n8990), .Z(n1631) );
  NANDN U1744 ( .A(n12219), .B(n1630), .Z(n1632) );
  NAND U1745 ( .A(n1631), .B(n1632), .Z(n8991) );
  ANDN U1746 ( .B(n4433), .A(n3438), .Z(n1633) );
  NAND U1747 ( .A(n5455), .B(n1633), .Z(n1634) );
  NANDN U1748 ( .A(n12393), .B(n1634), .Z(n1635) );
  ANDN U1749 ( .B(n5450), .A(n5453), .Z(n1636) );
  NAND U1750 ( .A(n1635), .B(n1636), .Z(n1637) );
  NANDN U1751 ( .A(n12396), .B(n1637), .Z(n1638) );
  AND U1752 ( .A(n5451), .B(n5446), .Z(n1639) );
  NANDN U1753 ( .A(n1638), .B(n5448), .Z(n1640) );
  AND U1754 ( .A(n1639), .B(n1640), .Z(n1641) );
  NOR U1755 ( .A(n5445), .B(n5449), .Z(n1642) );
  NANDN U1756 ( .A(n1641), .B(n1642), .Z(n1643) );
  AND U1757 ( .A(n12407), .B(n1643), .Z(n1644) );
  NAND U1758 ( .A(n1644), .B(n5447), .Z(n1645) );
  AND U1759 ( .A(n9099), .B(n1645), .Z(n1646) );
  NAND U1760 ( .A(n1646), .B(n5444), .Z(n1647) );
  AND U1761 ( .A(n12411), .B(n1647), .Z(n4436) );
  AND U1762 ( .A(n12296), .B(n5502), .Z(n1648) );
  NOR U1763 ( .A(n9026), .B(n9025), .Z(n1649) );
  NAND U1764 ( .A(n9024), .B(n1649), .Z(n1650) );
  NAND U1765 ( .A(n9027), .B(n1650), .Z(n1651) );
  NOR U1766 ( .A(n9029), .B(n9030), .Z(n1652) );
  NANDN U1767 ( .A(n1651), .B(n9028), .Z(n1653) );
  AND U1768 ( .A(n1652), .B(n1653), .Z(n1654) );
  ANDN U1769 ( .B(n9031), .A(n1654), .Z(n1655) );
  NAND U1770 ( .A(n12283), .B(n1655), .Z(n1656) );
  ANDN U1771 ( .B(n1656), .A(n9032), .Z(n1657) );
  NANDN U1772 ( .A(n12284), .B(n1657), .Z(n1658) );
  NAND U1773 ( .A(n12286), .B(n1658), .Z(n1659) );
  AND U1774 ( .A(n9035), .B(n1659), .Z(n1660) );
  NAND U1775 ( .A(n1660), .B(n12289), .Z(n1661) );
  AND U1776 ( .A(n12295), .B(n1661), .Z(n1662) );
  NANDN U1777 ( .A(n12290), .B(n1662), .Z(n1663) );
  NAND U1778 ( .A(n1648), .B(n1663), .Z(n9036) );
  ANDN U1779 ( .B(n4445), .A(n9150), .Z(n1664) );
  NAND U1780 ( .A(n12558), .B(n1664), .Z(n1665) );
  NAND U1781 ( .A(n5410), .B(n1665), .Z(n1666) );
  ANDN U1782 ( .B(n12566), .A(n9151), .Z(n1667) );
  NANDN U1783 ( .A(n1666), .B(n9153), .Z(n1668) );
  AND U1784 ( .A(n1667), .B(n1668), .Z(n1669) );
  NOR U1785 ( .A(n12569), .B(n1669), .Z(n1670) );
  NAND U1786 ( .A(n9154), .B(n1670), .Z(n1671) );
  ANDN U1787 ( .B(n1671), .A(n12571), .Z(n1672) );
  ANDN U1788 ( .B(n5409), .A(n1672), .Z(n1673) );
  NAND U1789 ( .A(n12573), .B(n1673), .Z(n1674) );
  AND U1790 ( .A(n12575), .B(n1674), .Z(n1675) );
  NAND U1791 ( .A(n9157), .B(n1675), .Z(n1676) );
  ANDN U1792 ( .B(n1676), .A(n5408), .Z(n1677) );
  NANDN U1793 ( .A(n12580), .B(n1677), .Z(n1678) );
  AND U1794 ( .A(n9158), .B(n1678), .Z(n4446) );
  NAND U1795 ( .A(n9107), .B(n9106), .Z(n1679) );
  AND U1796 ( .A(n12427), .B(n1679), .Z(n1680) );
  NAND U1797 ( .A(n1680), .B(n12422), .Z(n1681) );
  AND U1798 ( .A(n9108), .B(n12428), .Z(n1682) );
  NAND U1799 ( .A(n1681), .B(n1682), .Z(n1683) );
  NANDN U1800 ( .A(n12430), .B(n1683), .Z(n1684) );
  NAND U1801 ( .A(n12432), .B(n1684), .Z(n1685) );
  NANDN U1802 ( .A(n12434), .B(n1685), .Z(n1686) );
  ANDN U1803 ( .B(n1686), .A(n9113), .Z(n1687) );
  NOR U1804 ( .A(n9114), .B(n12441), .Z(n1688) );
  NANDN U1805 ( .A(n12436), .B(n1687), .Z(n1689) );
  NAND U1806 ( .A(n1688), .B(n1689), .Z(n1690) );
  AND U1807 ( .A(n12443), .B(n9115), .Z(n1691) );
  NAND U1808 ( .A(n1690), .B(n1691), .Z(n1692) );
  NANDN U1809 ( .A(n9116), .B(n1692), .Z(n9118) );
  NAND U1810 ( .A(n4449), .B(n4448), .Z(n1693) );
  ANDN U1811 ( .B(n1693), .A(n4450), .Z(n1694) );
  NAND U1812 ( .A(n5396), .B(n1694), .Z(n1695) );
  ANDN U1813 ( .B(n1695), .A(n9183), .Z(n1696) );
  NANDN U1814 ( .A(n12635), .B(n1696), .Z(n1697) );
  AND U1815 ( .A(n9185), .B(n5395), .Z(n1698) );
  NAND U1816 ( .A(n1697), .B(n1698), .Z(n1699) );
  NANDN U1817 ( .A(n12642), .B(n1699), .Z(n1700) );
  AND U1818 ( .A(n9184), .B(n12645), .Z(n1701) );
  OR U1819 ( .A(n1700), .B(n9182), .Z(n1702) );
  AND U1820 ( .A(n1701), .B(n1702), .Z(n1703) );
  AND U1821 ( .A(n5391), .B(n12649), .Z(n1704) );
  OR U1822 ( .A(n12647), .B(n1703), .Z(n1705) );
  AND U1823 ( .A(n1704), .B(n1705), .Z(n1706) );
  NOR U1824 ( .A(n5392), .B(n1706), .Z(n1707) );
  NAND U1825 ( .A(n12655), .B(n1707), .Z(n1708) );
  AND U1826 ( .A(n5390), .B(n1708), .Z(n4451) );
  AND U1827 ( .A(n12530), .B(n9143), .Z(n1709) );
  ANDN U1828 ( .B(n9137), .A(n9136), .Z(n1710) );
  NAND U1829 ( .A(n9135), .B(n1710), .Z(n1711) );
  AND U1830 ( .A(n12506), .B(n1711), .Z(n1712) );
  NAND U1831 ( .A(n1712), .B(n9138), .Z(n1713) );
  NAND U1832 ( .A(n12509), .B(n1713), .Z(n1714) );
  AND U1833 ( .A(n9139), .B(n1714), .Z(n1715) );
  NAND U1834 ( .A(n1715), .B(n12511), .Z(n1716) );
  AND U1835 ( .A(n5424), .B(n1716), .Z(n1717) );
  NAND U1836 ( .A(n1717), .B(n5423), .Z(n1718) );
  ANDN U1837 ( .B(n9141), .A(n9140), .Z(n1719) );
  NAND U1838 ( .A(n1718), .B(n1719), .Z(n1720) );
  NAND U1839 ( .A(n12521), .B(n1720), .Z(n1721) );
  AND U1840 ( .A(n12522), .B(n9142), .Z(n1722) );
  NAND U1841 ( .A(n1722), .B(n1721), .Z(n1723) );
  AND U1842 ( .A(n5420), .B(n1723), .Z(n1724) );
  NANDN U1843 ( .A(n12528), .B(n1724), .Z(n1725) );
  NAND U1844 ( .A(n1709), .B(n1725), .Z(n9144) );
  NAND U1845 ( .A(n4458), .B(n4457), .Z(n1726) );
  ANDN U1846 ( .B(n1726), .A(n4459), .Z(n1727) );
  NAND U1847 ( .A(n1727), .B(n5358), .Z(n1728) );
  ANDN U1848 ( .B(n1728), .A(n5356), .Z(n1729) );
  NANDN U1849 ( .A(n12732), .B(n1729), .Z(n1730) );
  AND U1850 ( .A(n5355), .B(n5359), .Z(n1731) );
  NAND U1851 ( .A(n1730), .B(n1731), .Z(n1732) );
  NAND U1852 ( .A(n12740), .B(n1732), .Z(n1733) );
  AND U1853 ( .A(n5354), .B(n12743), .Z(n1734) );
  NANDN U1854 ( .A(n1733), .B(n5357), .Z(n1735) );
  AND U1855 ( .A(n1734), .B(n1735), .Z(n1736) );
  OR U1856 ( .A(n12744), .B(n1736), .Z(n1737) );
  NAND U1857 ( .A(n12746), .B(n1737), .Z(n1738) );
  NANDN U1858 ( .A(n12749), .B(n1738), .Z(n4460) );
  ANDN U1859 ( .B(n9166), .A(n12592), .Z(n1739) );
  OR U1860 ( .A(n9165), .B(n9164), .Z(n1740) );
  AND U1861 ( .A(n1739), .B(n1740), .Z(n1741) );
  ANDN U1862 ( .B(n9167), .A(n1741), .Z(n1742) );
  NAND U1863 ( .A(n9168), .B(n1742), .Z(n1743) );
  ANDN U1864 ( .B(n1743), .A(n10188), .Z(n1744) );
  ANDN U1865 ( .B(n9170), .A(n10189), .Z(n1745) );
  NANDN U1866 ( .A(n9169), .B(n1744), .Z(n1746) );
  NAND U1867 ( .A(n1745), .B(n1746), .Z(n1747) );
  NOR U1868 ( .A(n9171), .B(n12601), .Z(n1748) );
  NAND U1869 ( .A(n1747), .B(n1748), .Z(n1749) );
  NAND U1870 ( .A(n9172), .B(n1749), .Z(n1750) );
  NANDN U1871 ( .A(n1750), .B(n9173), .Z(n1751) );
  NAND U1872 ( .A(n12605), .B(n1751), .Z(n1752) );
  NAND U1873 ( .A(n12607), .B(n1752), .Z(n1753) );
  ANDN U1874 ( .B(n9175), .A(n9174), .Z(n1754) );
  NAND U1875 ( .A(n1753), .B(n1754), .Z(n1755) );
  NANDN U1876 ( .A(n9176), .B(n1755), .Z(n9178) );
  NAND U1877 ( .A(n4465), .B(n12803), .Z(n1756) );
  AND U1878 ( .A(n9243), .B(n1756), .Z(n1757) );
  OR U1879 ( .A(n4468), .B(n9239), .Z(n1758) );
  NAND U1880 ( .A(n1757), .B(n1758), .Z(n1759) );
  NANDN U1881 ( .A(n12807), .B(n1759), .Z(n1760) );
  NAND U1882 ( .A(n12809), .B(n1760), .Z(n1761) );
  NANDN U1883 ( .A(n12811), .B(n1761), .Z(n1762) );
  AND U1884 ( .A(n12813), .B(n1762), .Z(n1763) );
  OR U1885 ( .A(n12814), .B(n1763), .Z(n1764) );
  NAND U1886 ( .A(n12816), .B(n1764), .Z(n1765) );
  NANDN U1887 ( .A(n12819), .B(n1765), .Z(n4471) );
  ANDN U1888 ( .B(n9198), .A(n9197), .Z(n1766) );
  AND U1889 ( .A(n9196), .B(n5385), .Z(n1767) );
  NAND U1890 ( .A(n12673), .B(n1767), .Z(n1768) );
  AND U1891 ( .A(n1766), .B(n1768), .Z(n1769) );
  AND U1892 ( .A(n9199), .B(n12679), .Z(n1770) );
  OR U1893 ( .A(n12677), .B(n1769), .Z(n1771) );
  AND U1894 ( .A(n1770), .B(n1771), .Z(n1772) );
  AND U1895 ( .A(n12686), .B(n9200), .Z(n1773) );
  NOR U1896 ( .A(n5382), .B(n1772), .Z(n1774) );
  NAND U1897 ( .A(n12685), .B(n1774), .Z(n1775) );
  AND U1898 ( .A(n1773), .B(n1775), .Z(n1776) );
  OR U1899 ( .A(n12689), .B(n1776), .Z(n1777) );
  NANDN U1900 ( .A(n12690), .B(n1777), .Z(n1778) );
  NAND U1901 ( .A(n12692), .B(n1778), .Z(n1779) );
  AND U1902 ( .A(n9203), .B(n12695), .Z(n1780) );
  NAND U1903 ( .A(n1779), .B(n1780), .Z(n1781) );
  NANDN U1904 ( .A(n12697), .B(n1781), .Z(n9204) );
  ANDN U1905 ( .B(n5326), .A(n5331), .Z(n4477) );
  NAND U1906 ( .A(n9224), .B(n12763), .Z(n1782) );
  NAND U1907 ( .A(n9227), .B(n1782), .Z(n1783) );
  AND U1908 ( .A(n12767), .B(n1783), .Z(n1784) );
  OR U1909 ( .A(n12768), .B(n1784), .Z(n1785) );
  NAND U1910 ( .A(n12770), .B(n1785), .Z(n1786) );
  NANDN U1911 ( .A(n12773), .B(n1786), .Z(n1787) );
  NAND U1912 ( .A(n12775), .B(n1787), .Z(n1788) );
  NANDN U1913 ( .A(n12777), .B(n1788), .Z(n1789) );
  AND U1914 ( .A(n9228), .B(n1789), .Z(n1790) );
  NAND U1915 ( .A(n1790), .B(n12779), .Z(n1791) );
  NANDN U1916 ( .A(n12780), .B(n1791), .Z(n1792) );
  AND U1917 ( .A(n9229), .B(n1792), .Z(n9231) );
  ANDN U1918 ( .B(n9255), .A(n9254), .Z(n1793) );
  ANDN U1919 ( .B(n9253), .A(n12836), .Z(n1794) );
  NAND U1920 ( .A(n12832), .B(n1794), .Z(n1795) );
  AND U1921 ( .A(n1793), .B(n1795), .Z(n1796) );
  AND U1922 ( .A(n9256), .B(n12842), .Z(n1797) );
  OR U1923 ( .A(n12840), .B(n1796), .Z(n1798) );
  AND U1924 ( .A(n1797), .B(n1798), .Z(n1799) );
  NOR U1925 ( .A(n12849), .B(n12845), .Z(n1800) );
  NANDN U1926 ( .A(n1799), .B(n1800), .Z(n1801) );
  AND U1927 ( .A(n9257), .B(n1801), .Z(n1802) );
  NAND U1928 ( .A(n1802), .B(n12851), .Z(n1803) );
  NANDN U1929 ( .A(n12852), .B(n1803), .Z(n1804) );
  AND U1930 ( .A(n9258), .B(n1804), .Z(n9259) );
  AND U1931 ( .A(n4494), .B(n12986), .Z(n1805) );
  NAND U1932 ( .A(n4493), .B(n1805), .Z(n1806) );
  NAND U1933 ( .A(n12993), .B(n1806), .Z(n1807) );
  NANDN U1934 ( .A(n1807), .B(n5292), .Z(n1808) );
  ANDN U1935 ( .B(n1808), .A(n12995), .Z(n1809) );
  ANDN U1936 ( .B(n12997), .A(n1809), .Z(n1810) );
  NAND U1937 ( .A(n5291), .B(n1810), .Z(n1811) );
  NANDN U1938 ( .A(n9305), .B(n1811), .Z(n1812) );
  NOR U1939 ( .A(n5290), .B(n5286), .Z(n1813) );
  NANDN U1940 ( .A(n1812), .B(n5288), .Z(n1814) );
  AND U1941 ( .A(n1813), .B(n1814), .Z(n1815) );
  ANDN U1942 ( .B(n5289), .A(n1815), .Z(n1816) );
  NAND U1943 ( .A(n13007), .B(n1816), .Z(n1817) );
  AND U1944 ( .A(n5287), .B(n1817), .Z(n1818) );
  NAND U1945 ( .A(n1818), .B(n5285), .Z(n1819) );
  NAND U1946 ( .A(n13013), .B(n1819), .Z(n1820) );
  AND U1947 ( .A(n13012), .B(n1820), .Z(n1821) );
  NAND U1948 ( .A(n5282), .B(n1821), .Z(n4495) );
  NOR U1949 ( .A(n12917), .B(n9272), .Z(n1822) );
  NAND U1950 ( .A(n9271), .B(n12915), .Z(n1823) );
  AND U1951 ( .A(n1822), .B(n1823), .Z(n1824) );
  NOR U1952 ( .A(n12919), .B(n1824), .Z(n1825) );
  NAND U1953 ( .A(n9273), .B(n1825), .Z(n1826) );
  ANDN U1954 ( .B(n1826), .A(n9274), .Z(n1827) );
  NAND U1955 ( .A(n1827), .B(n12925), .Z(n1828) );
  AND U1956 ( .A(n9275), .B(n1828), .Z(n1829) );
  NAND U1957 ( .A(n1829), .B(n9276), .Z(n1830) );
  NANDN U1958 ( .A(n12929), .B(n1830), .Z(n1831) );
  NAND U1959 ( .A(n12931), .B(n1831), .Z(n1832) );
  ANDN U1960 ( .B(n1832), .A(n12933), .Z(n1833) );
  NANDN U1961 ( .A(n1833), .B(n12935), .Z(n1834) );
  NAND U1962 ( .A(n12937), .B(n1834), .Z(n1835) );
  NANDN U1963 ( .A(n12939), .B(n1835), .Z(n1836) );
  NAND U1964 ( .A(n12941), .B(n1836), .Z(n1837) );
  AND U1965 ( .A(n12943), .B(n1837), .Z(n1838) );
  NANDN U1966 ( .A(n9277), .B(n1838), .Z(n9278) );
  AND U1967 ( .A(n12966), .B(n9291), .Z(n9292) );
  NAND U1968 ( .A(n4501), .B(n4500), .Z(n1839) );
  NANDN U1969 ( .A(n5252), .B(n1839), .Z(n1840) );
  ANDN U1970 ( .B(n1840), .A(n9349), .Z(n1841) );
  NAND U1971 ( .A(n1841), .B(n13113), .Z(n1842) );
  AND U1972 ( .A(n9351), .B(n1842), .Z(n1843) );
  NAND U1973 ( .A(n1843), .B(n13115), .Z(n1844) );
  NOR U1974 ( .A(n9348), .B(n5250), .Z(n1845) );
  NAND U1975 ( .A(n1844), .B(n1845), .Z(n1846) );
  NANDN U1976 ( .A(n13123), .B(n1846), .Z(n1847) );
  ANDN U1977 ( .B(n5251), .A(n9355), .Z(n1848) );
  OR U1978 ( .A(n1847), .B(n9350), .Z(n1849) );
  AND U1979 ( .A(n1848), .B(n1849), .Z(n1850) );
  NANDN U1980 ( .A(n1850), .B(n13127), .Z(n1851) );
  NAND U1981 ( .A(n13128), .B(n1851), .Z(n1852) );
  NAND U1982 ( .A(n13131), .B(n1852), .Z(n1853) );
  NANDN U1983 ( .A(n13133), .B(n1853), .Z(n4502) );
  NAND U1984 ( .A(n9308), .B(n13025), .Z(n1854) );
  AND U1985 ( .A(n13027), .B(n1854), .Z(n1855) );
  NAND U1986 ( .A(n1855), .B(n9309), .Z(n1856) );
  NAND U1987 ( .A(n13034), .B(n9310), .Z(n1857) );
  ANDN U1988 ( .B(n13028), .A(n5273), .Z(n1858) );
  NAND U1989 ( .A(n1856), .B(n1858), .Z(n1859) );
  NANDN U1990 ( .A(n1857), .B(n1859), .Z(n1860) );
  NOR U1991 ( .A(n13038), .B(n9311), .Z(n1861) );
  NANDN U1992 ( .A(n13037), .B(n1860), .Z(n1862) );
  NAND U1993 ( .A(n1861), .B(n1862), .Z(n1863) );
  ANDN U1994 ( .B(n9312), .A(n9313), .Z(n1864) );
  NAND U1995 ( .A(n1863), .B(n1864), .Z(n1865) );
  NANDN U1996 ( .A(n9314), .B(n1865), .Z(n1866) );
  AND U1997 ( .A(n9317), .B(n9316), .Z(n1867) );
  OR U1998 ( .A(n1866), .B(n9315), .Z(n1868) );
  AND U1999 ( .A(n1867), .B(n1868), .Z(n1869) );
  NOR U2000 ( .A(n9318), .B(n1869), .Z(n1870) );
  NANDN U2001 ( .A(n9319), .B(n1870), .Z(n1871) );
  AND U2002 ( .A(n9320), .B(n1871), .Z(n9321) );
  ANDN U2003 ( .B(n9367), .A(n13153), .Z(n1872) );
  NANDN U2004 ( .A(n9366), .B(n9365), .Z(n1873) );
  AND U2005 ( .A(n1872), .B(n1873), .Z(n1874) );
  NANDN U2006 ( .A(n1874), .B(n13155), .Z(n1875) );
  NAND U2007 ( .A(n13157), .B(n1875), .Z(n1876) );
  NANDN U2008 ( .A(n13159), .B(n1876), .Z(n1877) );
  NAND U2009 ( .A(n13161), .B(n1877), .Z(n1878) );
  NANDN U2010 ( .A(n13163), .B(n1878), .Z(n1879) );
  ANDN U2011 ( .B(n1879), .A(n13165), .Z(n1880) );
  NANDN U2012 ( .A(n1880), .B(n13167), .Z(n1881) );
  ANDN U2013 ( .B(n1881), .A(n13169), .Z(n1882) );
  ANDN U2014 ( .B(n9370), .A(n9369), .Z(n1883) );
  OR U2015 ( .A(n9368), .B(n1882), .Z(n1884) );
  AND U2016 ( .A(n1883), .B(n1884), .Z(n1885) );
  NOR U2017 ( .A(n1885), .B(n5234), .Z(n1886) );
  NAND U2018 ( .A(n13179), .B(n1886), .Z(n1887) );
  ANDN U2019 ( .B(n1887), .A(n9371), .Z(n1888) );
  NAND U2020 ( .A(n9372), .B(n1888), .Z(n9373) );
  AND U2021 ( .A(n4516), .B(n13286), .Z(n1889) );
  NANDN U2022 ( .A(n4514), .B(n4515), .Z(n1890) );
  AND U2023 ( .A(n1889), .B(n1890), .Z(n1891) );
  NANDN U2024 ( .A(n1891), .B(n13288), .Z(n1892) );
  AND U2025 ( .A(n5200), .B(n1892), .Z(n1893) );
  AND U2026 ( .A(n13295), .B(n13299), .Z(n1894) );
  OR U2027 ( .A(n13293), .B(n1893), .Z(n1895) );
  NAND U2028 ( .A(n1894), .B(n1895), .Z(n1896) );
  NAND U2029 ( .A(n13301), .B(n13296), .Z(n1897) );
  NAND U2030 ( .A(n4518), .B(n1897), .Z(n1898) );
  AND U2031 ( .A(n1896), .B(n1898), .Z(n1899) );
  OR U2032 ( .A(n13303), .B(n1899), .Z(n1900) );
  AND U2033 ( .A(n13305), .B(n1900), .Z(n1901) );
  NANDN U2034 ( .A(n1901), .B(n9418), .Z(n1902) );
  NAND U2035 ( .A(n13308), .B(n1902), .Z(n1903) );
  NAND U2036 ( .A(n13311), .B(n1903), .Z(n4519) );
  NAND U2037 ( .A(n9392), .B(n9391), .Z(n1904) );
  AND U2038 ( .A(n9395), .B(n1904), .Z(n1905) );
  ANDN U2039 ( .B(n5220), .A(n1905), .Z(n1906) );
  NAND U2040 ( .A(n13240), .B(n1906), .Z(n1907) );
  NANDN U2041 ( .A(n13243), .B(n1907), .Z(n1908) );
  ANDN U2042 ( .B(n5219), .A(n13249), .Z(n1909) );
  NANDN U2043 ( .A(n1908), .B(n13247), .Z(n1910) );
  AND U2044 ( .A(n1909), .B(n1910), .Z(n1911) );
  OR U2045 ( .A(n13251), .B(n1911), .Z(n1912) );
  AND U2046 ( .A(n9398), .B(n1912), .Z(n1913) );
  AND U2047 ( .A(n13259), .B(n13255), .Z(n1914) );
  NANDN U2048 ( .A(n13253), .B(n1913), .Z(n1915) );
  NAND U2049 ( .A(n1914), .B(n1915), .Z(n1916) );
  AND U2050 ( .A(n5218), .B(n13260), .Z(n1917) );
  NAND U2051 ( .A(n1916), .B(n1917), .Z(n1918) );
  NANDN U2052 ( .A(n13262), .B(n1918), .Z(n1919) );
  NAND U2053 ( .A(n13264), .B(n1919), .Z(n9411) );
  NAND U2054 ( .A(n9426), .B(n9425), .Z(n1920) );
  NANDN U2055 ( .A(n13325), .B(n1920), .Z(n1921) );
  AND U2056 ( .A(n9429), .B(n1921), .Z(n1922) );
  NAND U2057 ( .A(n1922), .B(n13327), .Z(n1923) );
  AND U2058 ( .A(n13333), .B(n1923), .Z(n1924) );
  NAND U2059 ( .A(n1924), .B(n13329), .Z(n1925) );
  ANDN U2060 ( .B(n5192), .A(n13335), .Z(n1926) );
  NAND U2061 ( .A(n1925), .B(n1926), .Z(n1927) );
  NANDN U2062 ( .A(n13337), .B(n1927), .Z(n1928) );
  NAND U2063 ( .A(n13339), .B(n1928), .Z(n1929) );
  NANDN U2064 ( .A(n13341), .B(n1929), .Z(n1930) );
  AND U2065 ( .A(n13343), .B(n1930), .Z(n1931) );
  OR U2066 ( .A(n13345), .B(n1931), .Z(n1932) );
  NAND U2067 ( .A(n13347), .B(n1932), .Z(n1933) );
  NAND U2068 ( .A(n13349), .B(n1933), .Z(n1934) );
  NAND U2069 ( .A(n13351), .B(n1934), .Z(n1935) );
  AND U2070 ( .A(n5179), .B(n1935), .Z(n1936) );
  NANDN U2071 ( .A(n5178), .B(n1936), .Z(n9434) );
  AND U2072 ( .A(n9443), .B(n13385), .Z(n1937) );
  NANDN U2073 ( .A(n9441), .B(n4524), .Z(n1938) );
  AND U2074 ( .A(n1937), .B(n1938), .Z(n1939) );
  AND U2075 ( .A(n5165), .B(n13389), .Z(n1940) );
  OR U2076 ( .A(n13387), .B(n1939), .Z(n1941) );
  AND U2077 ( .A(n1940), .B(n1941), .Z(n1942) );
  NANDN U2078 ( .A(n1942), .B(n13390), .Z(n1943) );
  NAND U2079 ( .A(n5168), .B(n1943), .Z(n1944) );
  NANDN U2080 ( .A(n13395), .B(n1944), .Z(n1945) );
  NAND U2081 ( .A(n13403), .B(n13398), .Z(n1946) );
  AND U2082 ( .A(n5164), .B(n13397), .Z(n1947) );
  NAND U2083 ( .A(n1945), .B(n1947), .Z(n1948) );
  NANDN U2084 ( .A(n1946), .B(n1948), .Z(n1949) );
  NOR U2085 ( .A(n5163), .B(n13405), .Z(n1950) );
  NAND U2086 ( .A(n1949), .B(n1950), .Z(n1951) );
  NAND U2087 ( .A(n13407), .B(n1951), .Z(n4525) );
  NANDN U2088 ( .A(n4550), .B(n4551), .Z(n1952) );
  NAND U2089 ( .A(n13467), .B(n1952), .Z(n1953) );
  NAND U2090 ( .A(n5146), .B(n1953), .Z(n1954) );
  ANDN U2091 ( .B(n9467), .A(n5145), .Z(n1955) );
  NANDN U2092 ( .A(n5143), .B(n1954), .Z(n1956) );
  NAND U2093 ( .A(n1955), .B(n1956), .Z(n1957) );
  NANDN U2094 ( .A(n5144), .B(n1957), .Z(n1958) );
  NANDN U2095 ( .A(n9469), .B(n1958), .Z(n1959) );
  AND U2096 ( .A(n9471), .B(n1959), .Z(n1960) );
  NOR U2097 ( .A(n9472), .B(n5141), .Z(n1961) );
  NANDN U2098 ( .A(n1960), .B(n1961), .Z(n1962) );
  ANDN U2099 ( .B(n1962), .A(n13479), .Z(n1963) );
  AND U2100 ( .A(n5142), .B(n13480), .Z(n1964) );
  NANDN U2101 ( .A(n9473), .B(n1963), .Z(n1965) );
  NAND U2102 ( .A(n1964), .B(n1965), .Z(n4560) );
  AND U2103 ( .A(n5154), .B(n5155), .Z(n1966) );
  NOR U2104 ( .A(n13437), .B(n13441), .Z(n1967) );
  NAND U2105 ( .A(n9457), .B(n1967), .Z(n1968) );
  AND U2106 ( .A(n1966), .B(n1968), .Z(n1969) );
  ANDN U2107 ( .B(n13447), .A(n13451), .Z(n1970) );
  OR U2108 ( .A(n1969), .B(n13445), .Z(n1971) );
  AND U2109 ( .A(n1970), .B(n1971), .Z(n1972) );
  NOR U2110 ( .A(n5151), .B(n1972), .Z(n1973) );
  NAND U2111 ( .A(n13448), .B(n1973), .Z(n1974) );
  AND U2112 ( .A(n13455), .B(n1974), .Z(n1975) );
  NANDN U2113 ( .A(n1975), .B(n13457), .Z(n1976) );
  NANDN U2114 ( .A(n13458), .B(n1976), .Z(n1977) );
  NANDN U2115 ( .A(n9460), .B(n1977), .Z(n1978) );
  NANDN U2116 ( .A(n9461), .B(n1978), .Z(n1979) );
  NAND U2117 ( .A(n9462), .B(n1979), .Z(n1980) );
  AND U2118 ( .A(n5147), .B(n1980), .Z(n1981) );
  NAND U2119 ( .A(n1981), .B(n5148), .Z(n9463) );
  ANDN U2120 ( .B(n9481), .A(n5127), .Z(n4562) );
  ANDN U2121 ( .B(n5116), .A(n5115), .Z(n1982) );
  NAND U2122 ( .A(n13529), .B(n9483), .Z(n1983) );
  AND U2123 ( .A(n1982), .B(n1983), .Z(n1984) );
  AND U2124 ( .A(n13538), .B(n5113), .Z(n1985) );
  NOR U2125 ( .A(n13537), .B(n1984), .Z(n1986) );
  NAND U2126 ( .A(n5114), .B(n1986), .Z(n1987) );
  AND U2127 ( .A(n1985), .B(n1987), .Z(n1988) );
  ANDN U2128 ( .B(n9484), .A(n1988), .Z(n1989) );
  NAND U2129 ( .A(n13541), .B(n1989), .Z(n1990) );
  ANDN U2130 ( .B(n1990), .A(n9485), .Z(n1991) );
  NANDN U2131 ( .A(n13542), .B(n1991), .Z(n1992) );
  NAND U2132 ( .A(n9486), .B(n1992), .Z(n1993) );
  ANDN U2133 ( .B(n1993), .A(n10186), .Z(n1994) );
  NANDN U2134 ( .A(n1994), .B(n13548), .Z(n1995) );
  NANDN U2135 ( .A(n13551), .B(n1995), .Z(n1996) );
  NAND U2136 ( .A(n13553), .B(n1996), .Z(n9489) );
  NAND U2137 ( .A(n4566), .B(n5087), .Z(n1997) );
  NAND U2138 ( .A(n13585), .B(n1997), .Z(n1998) );
  AND U2139 ( .A(n5090), .B(n1998), .Z(n1999) );
  AND U2140 ( .A(n13591), .B(n5086), .Z(n2000) );
  OR U2141 ( .A(n13589), .B(n1999), .Z(n2001) );
  AND U2142 ( .A(n2000), .B(n2001), .Z(n2002) );
  NOR U2143 ( .A(n13593), .B(n2002), .Z(n2003) );
  NAND U2144 ( .A(n13597), .B(n2003), .Z(n2004) );
  AND U2145 ( .A(n5085), .B(n2004), .Z(n2005) );
  NAND U2146 ( .A(n2005), .B(n13598), .Z(n2006) );
  NANDN U2147 ( .A(n13600), .B(n2006), .Z(n2007) );
  AND U2148 ( .A(n5081), .B(n2007), .Z(n2008) );
  NAND U2149 ( .A(n2008), .B(n13602), .Z(n2009) );
  NANDN U2150 ( .A(n13605), .B(n2009), .Z(n2010) );
  AND U2151 ( .A(n5083), .B(n2010), .Z(n4568) );
  NANDN U2152 ( .A(n9534), .B(n13667), .Z(n2011) );
  NANDN U2153 ( .A(n13672), .B(n2011), .Z(n2012) );
  NAND U2154 ( .A(n9535), .B(n2012), .Z(n2013) );
  NOR U2155 ( .A(n13680), .B(n13677), .Z(n2014) );
  NANDN U2156 ( .A(n2013), .B(n13674), .Z(n2015) );
  AND U2157 ( .A(n2014), .B(n2015), .Z(n2016) );
  NOR U2158 ( .A(n2016), .B(n5065), .Z(n2017) );
  NAND U2159 ( .A(n5066), .B(n2017), .Z(n2018) );
  ANDN U2160 ( .B(n2018), .A(n13685), .Z(n2019) );
  ANDN U2161 ( .B(n9536), .A(n2019), .Z(n2020) );
  NAND U2162 ( .A(n13687), .B(n2020), .Z(n2021) );
  AND U2163 ( .A(n13688), .B(n2021), .Z(n2022) );
  NAND U2164 ( .A(n2022), .B(n13692), .Z(n2023) );
  AND U2165 ( .A(n5062), .B(n2023), .Z(n2024) );
  NANDN U2166 ( .A(n13695), .B(n2024), .Z(n2025) );
  NANDN U2167 ( .A(n13697), .B(n2025), .Z(n9539) );
  NANDN U2168 ( .A(n4601), .B(n13723), .Z(n2026) );
  NANDN U2169 ( .A(n13727), .B(n2026), .Z(n2027) );
  ANDN U2170 ( .B(n2027), .A(n13729), .Z(n2028) );
  NANDN U2171 ( .A(n2028), .B(n13731), .Z(n2029) );
  NANDN U2172 ( .A(n13732), .B(n2029), .Z(n2030) );
  NAND U2173 ( .A(n5048), .B(n2030), .Z(n2031) );
  NOR U2174 ( .A(n13737), .B(n5045), .Z(n2032) );
  NANDN U2175 ( .A(n2031), .B(n13734), .Z(n2033) );
  AND U2176 ( .A(n2032), .B(n2033), .Z(n2034) );
  ANDN U2177 ( .B(n5044), .A(n2034), .Z(n2035) );
  NAND U2178 ( .A(n5047), .B(n2035), .Z(n2036) );
  AND U2179 ( .A(n13744), .B(n2036), .Z(n2037) );
  ANDN U2180 ( .B(n5043), .A(n13747), .Z(n2038) );
  NANDN U2181 ( .A(n5046), .B(n2037), .Z(n2039) );
  NAND U2182 ( .A(n2038), .B(n2039), .Z(n4602) );
  NAND U2183 ( .A(n9550), .B(n9549), .Z(n2040) );
  NANDN U2184 ( .A(n13754), .B(n2040), .Z(n2041) );
  NAND U2185 ( .A(n13756), .B(n2041), .Z(n2042) );
  NANDN U2186 ( .A(n13759), .B(n2042), .Z(n2043) );
  NANDN U2187 ( .A(n13761), .B(n2043), .Z(n2044) );
  AND U2188 ( .A(n13763), .B(n2044), .Z(n2045) );
  NOR U2189 ( .A(n2045), .B(n9554), .Z(n2046) );
  NAND U2190 ( .A(n9553), .B(n2046), .Z(n2047) );
  NANDN U2191 ( .A(n9555), .B(n2047), .Z(n2048) );
  NAND U2192 ( .A(n13769), .B(n2048), .Z(n2049) );
  NAND U2193 ( .A(n13773), .B(n2049), .Z(n2050) );
  AND U2194 ( .A(n13775), .B(n2050), .Z(n2051) );
  OR U2195 ( .A(n2051), .B(n13777), .Z(n2052) );
  NAND U2196 ( .A(n13779), .B(n2052), .Z(n2053) );
  AND U2197 ( .A(n9558), .B(n2053), .Z(n2054) );
  NAND U2198 ( .A(n13780), .B(n2054), .Z(n9559) );
  OR U2199 ( .A(n13827), .B(n4607), .Z(n2055) );
  NAND U2200 ( .A(n13829), .B(n2055), .Z(n2056) );
  NAND U2201 ( .A(n13831), .B(n2056), .Z(n2057) );
  AND U2202 ( .A(n5008), .B(n13832), .Z(n2058) );
  NAND U2203 ( .A(n2057), .B(n2058), .Z(n2059) );
  NAND U2204 ( .A(n5007), .B(n2059), .Z(n2060) );
  OR U2205 ( .A(n13835), .B(n2060), .Z(n2061) );
  AND U2206 ( .A(n5009), .B(n2061), .Z(n2062) );
  NAND U2207 ( .A(n2062), .B(n5004), .Z(n2063) );
  AND U2208 ( .A(n5003), .B(n2063), .Z(n2064) );
  NANDN U2209 ( .A(n5006), .B(n2064), .Z(n2065) );
  AND U2210 ( .A(n5005), .B(n13844), .Z(n2066) );
  NAND U2211 ( .A(n2065), .B(n2066), .Z(n2067) );
  NANDN U2212 ( .A(n13847), .B(n2067), .Z(n4609) );
  NANDN U2213 ( .A(n9620), .B(n9621), .Z(n2068) );
  NANDN U2214 ( .A(n13865), .B(n2068), .Z(n2069) );
  NANDN U2215 ( .A(n13867), .B(n2069), .Z(n2070) );
  NAND U2216 ( .A(n13869), .B(n2070), .Z(n2071) );
  ANDN U2217 ( .B(n2071), .A(n13871), .Z(n2072) );
  NANDN U2218 ( .A(n9622), .B(n2072), .Z(n2073) );
  AND U2219 ( .A(n9623), .B(n13873), .Z(n2074) );
  NAND U2220 ( .A(n2073), .B(n2074), .Z(n2075) );
  NAND U2221 ( .A(n9624), .B(n2075), .Z(n2076) );
  OR U2222 ( .A(n9625), .B(n2076), .Z(n2077) );
  AND U2223 ( .A(n9626), .B(n2077), .Z(n2078) );
  NANDN U2224 ( .A(y[1682]), .B(x[1682]), .Z(n2079) );
  NAND U2225 ( .A(n2078), .B(n2079), .Z(n2080) );
  NANDN U2226 ( .A(n9627), .B(n2080), .Z(n2081) );
  OR U2227 ( .A(n9628), .B(n2081), .Z(n2082) );
  AND U2228 ( .A(n13885), .B(n2082), .Z(n2083) );
  NANDN U2229 ( .A(y[1684]), .B(x[1684]), .Z(n2084) );
  NAND U2230 ( .A(n2083), .B(n2084), .Z(n2085) );
  NANDN U2231 ( .A(n9629), .B(n2085), .Z(n9630) );
  NANDN U2232 ( .A(n4636), .B(n9637), .Z(n2086) );
  NANDN U2233 ( .A(n9638), .B(n2086), .Z(n2087) );
  ANDN U2234 ( .B(n2087), .A(n9639), .Z(n2088) );
  AND U2235 ( .A(n9643), .B(n9640), .Z(n2089) );
  OR U2236 ( .A(n4989), .B(n2088), .Z(n2090) );
  AND U2237 ( .A(n2089), .B(n2090), .Z(n2091) );
  NANDN U2238 ( .A(n2091), .B(n13922), .Z(n2092) );
  NAND U2239 ( .A(n13925), .B(n2092), .Z(n2093) );
  NAND U2240 ( .A(n13927), .B(n2093), .Z(n2094) );
  NANDN U2241 ( .A(n13929), .B(n2094), .Z(n2095) );
  NAND U2242 ( .A(n13931), .B(n2095), .Z(n2096) );
  ANDN U2243 ( .B(n2096), .A(n9646), .Z(n2097) );
  NAND U2244 ( .A(n2097), .B(n13932), .Z(n2098) );
  AND U2245 ( .A(n9649), .B(n2098), .Z(n2099) );
  NANDN U2246 ( .A(n13935), .B(n2099), .Z(n2100) );
  AND U2247 ( .A(n9647), .B(n2100), .Z(n4639) );
  NAND U2248 ( .A(n9651), .B(n9650), .Z(n2101) );
  NAND U2249 ( .A(n9654), .B(n2101), .Z(n2102) );
  ANDN U2250 ( .B(n2102), .A(n9655), .Z(n2103) );
  AND U2251 ( .A(n4978), .B(n4977), .Z(n2104) );
  NANDN U2252 ( .A(n13947), .B(n2103), .Z(n2105) );
  NAND U2253 ( .A(n2104), .B(n2105), .Z(n2106) );
  NAND U2254 ( .A(n4974), .B(n4973), .Z(n2107) );
  AND U2255 ( .A(n4975), .B(n4976), .Z(n2108) );
  NAND U2256 ( .A(n2106), .B(n2108), .Z(n2109) );
  NANDN U2257 ( .A(n2107), .B(n2109), .Z(n2110) );
  AND U2258 ( .A(n4972), .B(n4971), .Z(n2111) );
  NAND U2259 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2260 ( .A(n9657), .B(n2112), .Z(n2113) );
  NAND U2261 ( .A(n2113), .B(n9656), .Z(n2114) );
  NOR U2262 ( .A(n9658), .B(n13963), .Z(n2115) );
  NAND U2263 ( .A(n2114), .B(n2115), .Z(n2116) );
  NAND U2264 ( .A(n9659), .B(n2116), .Z(n2117) );
  NANDN U2265 ( .A(n2117), .B(n9660), .Z(n2118) );
  AND U2266 ( .A(n13966), .B(n2118), .Z(n9665) );
  AND U2267 ( .A(n4642), .B(n4959), .Z(n2119) );
  NAND U2268 ( .A(n4955), .B(n2119), .Z(n2120) );
  NAND U2269 ( .A(n13996), .B(n2120), .Z(n2121) );
  NOR U2270 ( .A(n13999), .B(n4956), .Z(n2122) );
  NANDN U2271 ( .A(n2121), .B(n4957), .Z(n2123) );
  AND U2272 ( .A(n2122), .B(n2123), .Z(n2124) );
  NANDN U2273 ( .A(n2124), .B(n14001), .Z(n2125) );
  NAND U2274 ( .A(n14002), .B(n2125), .Z(n2126) );
  NANDN U2275 ( .A(n14005), .B(n2126), .Z(n2127) );
  NANDN U2276 ( .A(n14007), .B(n2127), .Z(n2128) );
  NAND U2277 ( .A(n14009), .B(n2128), .Z(n2129) );
  ANDN U2278 ( .B(n2129), .A(n14011), .Z(n2130) );
  NANDN U2279 ( .A(n2130), .B(n14013), .Z(n2131) );
  ANDN U2280 ( .B(n2131), .A(n14014), .Z(n2132) );
  NAND U2281 ( .A(n2132), .B(n9680), .Z(n2133) );
  AND U2282 ( .A(n9682), .B(n2133), .Z(n2134) );
  NANDN U2283 ( .A(n14017), .B(n2134), .Z(n4643) );
  NAND U2284 ( .A(n4947), .B(n4946), .Z(n2135) );
  NOR U2285 ( .A(n14024), .B(n9685), .Z(n2136) );
  NAND U2286 ( .A(n9684), .B(n9683), .Z(n2137) );
  AND U2287 ( .A(n2136), .B(n2137), .Z(n2138) );
  AND U2288 ( .A(n4944), .B(n4945), .Z(n2139) );
  OR U2289 ( .A(n2135), .B(n2138), .Z(n2140) );
  AND U2290 ( .A(n2139), .B(n2140), .Z(n2141) );
  ANDN U2291 ( .B(n4943), .A(n2141), .Z(n2142) );
  NAND U2292 ( .A(n4942), .B(n2142), .Z(n2143) );
  AND U2293 ( .A(n14036), .B(n2143), .Z(n2144) );
  NANDN U2294 ( .A(y[1750]), .B(x[1750]), .Z(n2145) );
  NAND U2295 ( .A(n2144), .B(n2145), .Z(n2146) );
  NANDN U2296 ( .A(n9686), .B(n2146), .Z(n2147) );
  OR U2297 ( .A(n2147), .B(n14039), .Z(n2148) );
  NAND U2298 ( .A(n14041), .B(n2148), .Z(n2149) );
  NANDN U2299 ( .A(n14043), .B(n2149), .Z(n2150) );
  NAND U2300 ( .A(n14045), .B(n2150), .Z(n9689) );
  AND U2301 ( .A(n4651), .B(n4921), .Z(n2151) );
  NAND U2302 ( .A(n4917), .B(n2151), .Z(n2152) );
  NANDN U2303 ( .A(n14097), .B(n2152), .Z(n2153) );
  AND U2304 ( .A(n4918), .B(n14099), .Z(n2154) );
  NANDN U2305 ( .A(n2153), .B(n4920), .Z(n2155) );
  AND U2306 ( .A(n2154), .B(n2155), .Z(n2156) );
  NANDN U2307 ( .A(n2156), .B(n14101), .Z(n2157) );
  NANDN U2308 ( .A(n14103), .B(n2157), .Z(n2158) );
  NAND U2309 ( .A(n14105), .B(n2158), .Z(n2159) );
  NANDN U2310 ( .A(n14107), .B(n2159), .Z(n2160) );
  NAND U2311 ( .A(n14109), .B(n2160), .Z(n2161) );
  ANDN U2312 ( .B(n2161), .A(n14111), .Z(n2162) );
  NANDN U2313 ( .A(n2162), .B(n14113), .Z(n2163) );
  ANDN U2314 ( .B(n2163), .A(n4913), .Z(n2164) );
  ANDN U2315 ( .B(n4910), .A(n14116), .Z(n2165) );
  NANDN U2316 ( .A(n14115), .B(n2164), .Z(n2166) );
  NAND U2317 ( .A(n2165), .B(n2166), .Z(n4652) );
  AND U2318 ( .A(n14123), .B(n4909), .Z(n9759) );
  NAND U2319 ( .A(n4657), .B(n14204), .Z(n2167) );
  NANDN U2320 ( .A(n14207), .B(n2167), .Z(n2168) );
  ANDN U2321 ( .B(n2168), .A(n14209), .Z(n2169) );
  NANDN U2322 ( .A(n2169), .B(n14211), .Z(n2170) );
  ANDN U2323 ( .B(n2170), .A(n14212), .Z(n2171) );
  NOR U2324 ( .A(n14216), .B(n4880), .Z(n2172) );
  NANDN U2325 ( .A(n2171), .B(n14214), .Z(n2173) );
  AND U2326 ( .A(n2172), .B(n2173), .Z(n2174) );
  ANDN U2327 ( .B(n14222), .A(n2174), .Z(n2175) );
  NAND U2328 ( .A(n14218), .B(n2175), .Z(n2176) );
  AND U2329 ( .A(n14225), .B(n2176), .Z(n2177) );
  NAND U2330 ( .A(n4881), .B(n2177), .Z(n4658) );
  AND U2331 ( .A(n9837), .B(n9838), .Z(n2178) );
  ANDN U2332 ( .B(n9839), .A(n2178), .Z(n2179) );
  NANDN U2333 ( .A(y[1836]), .B(x[1836]), .Z(n2180) );
  NAND U2334 ( .A(n2179), .B(n2180), .Z(n2181) );
  AND U2335 ( .A(n4875), .B(n4876), .Z(n2182) );
  NAND U2336 ( .A(n2181), .B(n2182), .Z(n2183) );
  NANDN U2337 ( .A(n14236), .B(n2183), .Z(n2184) );
  NANDN U2338 ( .A(y[1838]), .B(x[1838]), .Z(n2185) );
  NANDN U2339 ( .A(n2184), .B(n2185), .Z(n2186) );
  AND U2340 ( .A(n9840), .B(n2186), .Z(n2187) );
  NANDN U2341 ( .A(n14239), .B(n2187), .Z(n2188) );
  NAND U2342 ( .A(n14241), .B(n2188), .Z(n2189) );
  ANDN U2343 ( .B(n2189), .A(n14243), .Z(n2190) );
  NANDN U2344 ( .A(n2190), .B(n14245), .Z(n2191) );
  AND U2345 ( .A(n14246), .B(n2191), .Z(n2192) );
  NOR U2346 ( .A(n9841), .B(n2192), .Z(n2193) );
  NAND U2347 ( .A(n9842), .B(n2193), .Z(n2194) );
  ANDN U2348 ( .B(n2194), .A(n9843), .Z(n2195) );
  NAND U2349 ( .A(n9844), .B(n2195), .Z(n9845) );
  NAND U2350 ( .A(n4663), .B(n14283), .Z(n2196) );
  NANDN U2351 ( .A(n14285), .B(n2196), .Z(n2197) );
  AND U2352 ( .A(n14287), .B(n2197), .Z(n2198) );
  NOR U2353 ( .A(n2198), .B(n9880), .Z(n2199) );
  NAND U2354 ( .A(n9884), .B(n2199), .Z(n2200) );
  NAND U2355 ( .A(n9887), .B(n2200), .Z(n2201) );
  AND U2356 ( .A(n4851), .B(n9885), .Z(n2202) );
  NANDN U2357 ( .A(n2201), .B(n9883), .Z(n2203) );
  AND U2358 ( .A(n2202), .B(n2203), .Z(n2204) );
  NOR U2359 ( .A(n9886), .B(n4849), .Z(n2205) );
  NANDN U2360 ( .A(n2204), .B(n2205), .Z(n2206) );
  ANDN U2361 ( .B(n2206), .A(n9888), .Z(n2207) );
  NAND U2362 ( .A(n2207), .B(n4852), .Z(n2208) );
  AND U2363 ( .A(n9891), .B(n2208), .Z(n2209) );
  NAND U2364 ( .A(n2209), .B(n4850), .Z(n2210) );
  AND U2365 ( .A(n14304), .B(n2210), .Z(n4664) );
  NOR U2366 ( .A(n9922), .B(n14336), .Z(n2211) );
  NANDN U2367 ( .A(n9923), .B(n2211), .Z(n2212) );
  NAND U2368 ( .A(n9924), .B(n2212), .Z(n2213) );
  NANDN U2369 ( .A(n2213), .B(n9925), .Z(n2214) );
  AND U2370 ( .A(n14339), .B(n2214), .Z(n2215) );
  NOR U2371 ( .A(n14342), .B(n2215), .Z(n2216) );
  NAND U2372 ( .A(n4835), .B(n2216), .Z(n2217) );
  ANDN U2373 ( .B(n2217), .A(n14347), .Z(n2218) );
  NANDN U2374 ( .A(n2218), .B(n14349), .Z(n2219) );
  NANDN U2375 ( .A(n14351), .B(n2219), .Z(n2220) );
  NAND U2376 ( .A(n14353), .B(n2220), .Z(n2221) );
  ANDN U2377 ( .B(n14355), .A(n9928), .Z(n2222) );
  NAND U2378 ( .A(n2221), .B(n2222), .Z(n2223) );
  NAND U2379 ( .A(n9929), .B(n2223), .Z(n2224) );
  AND U2380 ( .A(n9931), .B(n9930), .Z(n2225) );
  OR U2381 ( .A(n2224), .B(n14356), .Z(n2226) );
  AND U2382 ( .A(n2225), .B(n2226), .Z(n9935) );
  NAND U2383 ( .A(n4672), .B(n4817), .Z(n2227) );
  NANDN U2384 ( .A(n14411), .B(n2227), .Z(n2228) );
  AND U2385 ( .A(n14413), .B(n2228), .Z(n2229) );
  OR U2386 ( .A(n2229), .B(n14415), .Z(n2230) );
  NAND U2387 ( .A(n14417), .B(n2230), .Z(n2231) );
  ANDN U2388 ( .B(n2231), .A(n14419), .Z(n2232) );
  NANDN U2389 ( .A(n2232), .B(n14421), .Z(n2233) );
  AND U2390 ( .A(n14423), .B(n2233), .Z(n2234) );
  NOR U2391 ( .A(n4806), .B(n14425), .Z(n2235) );
  NANDN U2392 ( .A(n2234), .B(n2235), .Z(n2236) );
  AND U2393 ( .A(n14427), .B(n2236), .Z(n2237) );
  NAND U2394 ( .A(n2237), .B(n4803), .Z(n2238) );
  AND U2395 ( .A(n4805), .B(n2238), .Z(n2239) );
  NANDN U2396 ( .A(n14433), .B(n2239), .Z(n2240) );
  AND U2397 ( .A(n4804), .B(n14435), .Z(n2241) );
  NAND U2398 ( .A(n2240), .B(n2241), .Z(n2242) );
  NANDN U2399 ( .A(n14436), .B(n2242), .Z(n2243) );
  NAND U2400 ( .A(n14439), .B(n2243), .Z(n4673) );
  NAND U2401 ( .A(n4683), .B(n4682), .Z(n2244) );
  NANDN U2402 ( .A(n4685), .B(n2244), .Z(n2245) );
  AND U2403 ( .A(n14523), .B(n2245), .Z(n2246) );
  OR U2404 ( .A(n14524), .B(n2246), .Z(n2247) );
  NAND U2405 ( .A(n14527), .B(n2247), .Z(n2248) );
  NAND U2406 ( .A(n14528), .B(n2248), .Z(n2249) );
  NAND U2407 ( .A(n14537), .B(n14532), .Z(n2250) );
  AND U2408 ( .A(n10109), .B(n14531), .Z(n2251) );
  NAND U2409 ( .A(n2249), .B(n2251), .Z(n2252) );
  NANDN U2410 ( .A(n2250), .B(n2252), .Z(n2253) );
  NOR U2411 ( .A(n10110), .B(n14538), .Z(n2254) );
  NAND U2412 ( .A(n2253), .B(n2254), .Z(n2255) );
  NAND U2413 ( .A(n14541), .B(n2255), .Z(n2256) );
  NAND U2414 ( .A(n14543), .B(n2256), .Z(n2257) );
  AND U2415 ( .A(n10123), .B(n2257), .Z(n2258) );
  NANDN U2416 ( .A(n14544), .B(n2258), .Z(n4689) );
  NANDN U2417 ( .A(n10130), .B(n10129), .Z(n2259) );
  NAND U2418 ( .A(n10131), .B(n2259), .Z(n2260) );
  NAND U2419 ( .A(n10132), .B(n2260), .Z(n2261) );
  NAND U2420 ( .A(n10133), .B(n2261), .Z(n2262) );
  AND U2421 ( .A(n4765), .B(n2262), .Z(n2263) );
  NAND U2422 ( .A(n2263), .B(n14580), .Z(n2264) );
  NAND U2423 ( .A(n14583), .B(n2264), .Z(n2265) );
  AND U2424 ( .A(n14584), .B(n2265), .Z(n2266) );
  NAND U2425 ( .A(n2266), .B(n4764), .Z(n2267) );
  ANDN U2426 ( .B(n2267), .A(n10136), .Z(n2268) );
  AND U2427 ( .A(n4762), .B(n4763), .Z(n2269) );
  NANDN U2428 ( .A(n14586), .B(n2268), .Z(n2270) );
  NAND U2429 ( .A(n2269), .B(n2270), .Z(n2271) );
  NANDN U2430 ( .A(n4759), .B(n4760), .Z(n2272) );
  AND U2431 ( .A(n4761), .B(n14595), .Z(n2273) );
  NAND U2432 ( .A(n2271), .B(n2273), .Z(n2274) );
  NANDN U2433 ( .A(n2272), .B(n2274), .Z(n10137) );
  NANDN U2434 ( .A(n4706), .B(n4705), .Z(n2275) );
  NAND U2435 ( .A(n14634), .B(n2275), .Z(n2276) );
  AND U2436 ( .A(n4748), .B(n2276), .Z(n2277) );
  NANDN U2437 ( .A(n2277), .B(n14639), .Z(n2278) );
  ANDN U2438 ( .B(n2278), .A(n14641), .Z(n2279) );
  OR U2439 ( .A(n14643), .B(n2279), .Z(n2280) );
  NAND U2440 ( .A(n10152), .B(n2280), .Z(n2281) );
  NAND U2441 ( .A(n14647), .B(n2281), .Z(n2282) );
  ANDN U2442 ( .B(n4745), .A(n10151), .Z(n2283) );
  NAND U2443 ( .A(n2282), .B(n2283), .Z(n2284) );
  NANDN U2444 ( .A(n14651), .B(n2284), .Z(n2285) );
  NOR U2445 ( .A(n4744), .B(n10172), .Z(n2286) );
  NAND U2446 ( .A(n2285), .B(n2286), .Z(n2287) );
  NAND U2447 ( .A(n14654), .B(n2287), .Z(n2288) );
  NAND U2448 ( .A(n14657), .B(n2288), .Z(n4711) );
  NANDN U2449 ( .A(n10166), .B(n14693), .Z(n2289) );
  NAND U2450 ( .A(n14694), .B(n2289), .Z(n2290) );
  NAND U2451 ( .A(n14695), .B(n2290), .Z(n2291) );
  AND U2452 ( .A(n3192), .B(n3189), .Z(n2292) );
  AND U2453 ( .A(n14704), .B(n2292), .Z(n2293) );
  ANDN U2454 ( .B(n2293), .A(n3188), .Z(n2294) );
  AND U2455 ( .A(n3191), .B(n2294), .Z(n2295) );
  XNOR U2456 ( .A(y[2039]), .B(x[2039]), .Z(n2296) );
  NAND U2457 ( .A(n2295), .B(n2296), .Z(n2297) );
  NANDN U2458 ( .A(n4721), .B(n4720), .Z(n2298) );
  NANDN U2459 ( .A(n4722), .B(n2298), .Z(n2299) );
  NANDN U2460 ( .A(n2297), .B(n2299), .Z(n2300) );
  AND U2461 ( .A(n14705), .B(n14702), .Z(n2301) );
  AND U2462 ( .A(n14703), .B(n2301), .Z(n2302) );
  NANDN U2463 ( .A(n14706), .B(n2302), .Z(n2303) );
  NAND U2464 ( .A(n14696), .B(n2291), .Z(n2304) );
  ANDN U2465 ( .B(n2304), .A(n2303), .Z(n2305) );
  NANDN U2466 ( .A(n2300), .B(n2305), .Z(n10167) );
  AND U2467 ( .A(n6468), .B(n6467), .Z(n2306) );
  NAND U2468 ( .A(n6469), .B(n2306), .Z(n2307) );
  ANDN U2469 ( .B(n2307), .A(n6470), .Z(n2308) );
  NANDN U2470 ( .A(n2308), .B(n6471), .Z(n2309) );
  NAND U2471 ( .A(n10486), .B(n2309), .Z(n2310) );
  NANDN U2472 ( .A(n10489), .B(n2310), .Z(n2311) );
  NANDN U2473 ( .A(n6472), .B(n2311), .Z(n2312) );
  NAND U2474 ( .A(n6473), .B(n2312), .Z(n2313) );
  ANDN U2475 ( .B(n2313), .A(n6474), .Z(n2314) );
  AND U2476 ( .A(n6476), .B(n6477), .Z(n2315) );
  NANDN U2477 ( .A(n6475), .B(n2314), .Z(n2316) );
  NAND U2478 ( .A(n2315), .B(n2316), .Z(n2317) );
  ANDN U2479 ( .B(n2317), .A(n6478), .Z(n2318) );
  AND U2480 ( .A(n5877), .B(n5876), .Z(n2319) );
  NANDN U2481 ( .A(n6479), .B(n2318), .Z(n2320) );
  NAND U2482 ( .A(n2319), .B(n2320), .Z(n2321) );
  ANDN U2483 ( .B(n2321), .A(n6480), .Z(n2322) );
  NANDN U2484 ( .A(n6481), .B(n2322), .Z(n6482) );
  NAND U2485 ( .A(n6888), .B(n6889), .Z(n2323) );
  ANDN U2486 ( .B(n2323), .A(n6890), .Z(n2324) );
  AND U2487 ( .A(n5838), .B(n5839), .Z(n2325) );
  NANDN U2488 ( .A(n6891), .B(n2324), .Z(n2326) );
  AND U2489 ( .A(n2325), .B(n2326), .Z(n2327) );
  NOR U2490 ( .A(n6892), .B(n2327), .Z(n2328) );
  NANDN U2491 ( .A(n6893), .B(n2328), .Z(n2329) );
  NAND U2492 ( .A(n6894), .B(n2329), .Z(n2330) );
  NOR U2493 ( .A(n6896), .B(n6897), .Z(n2331) );
  NANDN U2494 ( .A(n2330), .B(n6895), .Z(n2332) );
  AND U2495 ( .A(n2331), .B(n2332), .Z(n2333) );
  ANDN U2496 ( .B(n6899), .A(n2333), .Z(n2334) );
  NAND U2497 ( .A(n6898), .B(n2334), .Z(n2335) );
  ANDN U2498 ( .B(n2335), .A(n10738), .Z(n2336) );
  AND U2499 ( .A(n10739), .B(n5837), .Z(n2337) );
  NANDN U2500 ( .A(n6900), .B(n2336), .Z(n2338) );
  NAND U2501 ( .A(n2337), .B(n2338), .Z(n2339) );
  ANDN U2502 ( .B(n2339), .A(n6901), .Z(n2340) );
  NANDN U2503 ( .A(n6902), .B(n2340), .Z(n6903) );
  NANDN U2504 ( .A(x[0]), .B(y[0]), .Z(n2341) );
  NAND U2505 ( .A(n5927), .B(n2341), .Z(n2342) );
  NANDN U2506 ( .A(n5929), .B(n2342), .Z(n2343) );
  NAND U2507 ( .A(n5931), .B(n2343), .Z(n2344) );
  NANDN U2508 ( .A(n5934), .B(n2344), .Z(n2345) );
  AND U2509 ( .A(n5936), .B(n2345), .Z(n2346) );
  OR U2510 ( .A(n2346), .B(n5938), .Z(n2347) );
  NAND U2511 ( .A(n10193), .B(n2347), .Z(n2348) );
  NANDN U2512 ( .A(n10195), .B(n2348), .Z(n2349) );
  NAND U2513 ( .A(n10197), .B(n2349), .Z(n2350) );
  NANDN U2514 ( .A(n10199), .B(n2350), .Z(n2351) );
  AND U2515 ( .A(n10201), .B(n2351), .Z(n3609) );
  NANDN U2516 ( .A(n11486), .B(n8221), .Z(n2352) );
  NAND U2517 ( .A(n11488), .B(n2352), .Z(n2353) );
  ANDN U2518 ( .B(n2353), .A(n11491), .Z(n2354) );
  NANDN U2519 ( .A(n2354), .B(n11493), .Z(n2355) );
  NANDN U2520 ( .A(n8222), .B(n2355), .Z(n2356) );
  NAND U2521 ( .A(n8223), .B(n2356), .Z(n2357) );
  NOR U2522 ( .A(n8225), .B(n8224), .Z(n2358) );
  NAND U2523 ( .A(n2357), .B(n2358), .Z(n2359) );
  NAND U2524 ( .A(n8226), .B(n2359), .Z(n2360) );
  NOR U2525 ( .A(n8229), .B(n8228), .Z(n2361) );
  NANDN U2526 ( .A(n2360), .B(n8227), .Z(n2362) );
  AND U2527 ( .A(n2361), .B(n2362), .Z(n2363) );
  ANDN U2528 ( .B(n8231), .A(n2363), .Z(n2364) );
  NAND U2529 ( .A(n8230), .B(n2364), .Z(n2365) );
  ANDN U2530 ( .B(n2365), .A(n8232), .Z(n2366) );
  NANDN U2531 ( .A(n8233), .B(n2366), .Z(n8234) );
  NANDN U2532 ( .A(n4324), .B(n4325), .Z(n2367) );
  NAND U2533 ( .A(n4326), .B(n2367), .Z(n2368) );
  NAND U2534 ( .A(n11656), .B(n2368), .Z(n2369) );
  NANDN U2535 ( .A(n11659), .B(n2369), .Z(n2370) );
  NAND U2536 ( .A(n11661), .B(n2370), .Z(n2371) );
  ANDN U2537 ( .B(n2371), .A(n11663), .Z(n2372) );
  NANDN U2538 ( .A(n2372), .B(n11665), .Z(n2373) );
  ANDN U2539 ( .B(n2373), .A(n11666), .Z(n2374) );
  NANDN U2540 ( .A(n2374), .B(n11668), .Z(n2375) );
  NANDN U2541 ( .A(n11671), .B(n2375), .Z(n2376) );
  NAND U2542 ( .A(n11673), .B(n2376), .Z(n4327) );
  NAND U2543 ( .A(n4332), .B(n4331), .Z(n2377) );
  NANDN U2544 ( .A(n4333), .B(n2377), .Z(n2378) );
  NANDN U2545 ( .A(n11726), .B(n2378), .Z(n2379) );
  NAND U2546 ( .A(n11728), .B(n2379), .Z(n2380) );
  NAND U2547 ( .A(n8587), .B(n2380), .Z(n2381) );
  ANDN U2548 ( .B(n2381), .A(n8589), .Z(n2382) );
  NANDN U2549 ( .A(n2382), .B(n8591), .Z(n2383) );
  NANDN U2550 ( .A(n8594), .B(n2383), .Z(n2384) );
  NAND U2551 ( .A(n8596), .B(n2384), .Z(n2385) );
  NANDN U2552 ( .A(n8598), .B(n2385), .Z(n2386) );
  NAND U2553 ( .A(n8600), .B(n2386), .Z(n2387) );
  ANDN U2554 ( .B(n2387), .A(n8601), .Z(n2388) );
  NANDN U2555 ( .A(n2388), .B(n8603), .Z(n2389) );
  ANDN U2556 ( .B(n2389), .A(n8606), .Z(n2390) );
  NANDN U2557 ( .A(n2390), .B(n8608), .Z(n2391) );
  NAND U2558 ( .A(n11752), .B(n2391), .Z(n2392) );
  NANDN U2559 ( .A(n11755), .B(n2392), .Z(n4342) );
  NAND U2560 ( .A(n4396), .B(n12009), .Z(n2393) );
  NAND U2561 ( .A(n12011), .B(n2393), .Z(n2394) );
  NAND U2562 ( .A(n12013), .B(n2394), .Z(n2395) );
  NAND U2563 ( .A(n12015), .B(n2395), .Z(n2396) );
  NANDN U2564 ( .A(n12017), .B(n2396), .Z(n2397) );
  AND U2565 ( .A(n12019), .B(n2397), .Z(n2398) );
  ANDN U2566 ( .B(n5560), .A(n12023), .Z(n2399) );
  OR U2567 ( .A(n12021), .B(n2398), .Z(n2400) );
  AND U2568 ( .A(n2399), .B(n2400), .Z(n2401) );
  NOR U2569 ( .A(n8870), .B(n2401), .Z(n2402) );
  NAND U2570 ( .A(n12025), .B(n2402), .Z(n2403) );
  AND U2571 ( .A(n5561), .B(n2403), .Z(n2404) );
  NAND U2572 ( .A(n8871), .B(n2404), .Z(n2405) );
  ANDN U2573 ( .B(n2405), .A(n5558), .Z(n2406) );
  NANDN U2574 ( .A(n8869), .B(n2406), .Z(n2407) );
  AND U2575 ( .A(n8872), .B(n2407), .Z(n4397) );
  NAND U2576 ( .A(n12083), .B(n4409), .Z(n2408) );
  NANDN U2577 ( .A(n12085), .B(n2408), .Z(n2409) );
  AND U2578 ( .A(n12087), .B(n2409), .Z(n2410) );
  NAND U2579 ( .A(n2410), .B(n5540), .Z(n2411) );
  AND U2580 ( .A(n12089), .B(n2411), .Z(n2412) );
  NANDN U2581 ( .A(n5538), .B(n2412), .Z(n2413) );
  ANDN U2582 ( .B(n5535), .A(n5539), .Z(n2414) );
  NAND U2583 ( .A(n2413), .B(n2414), .Z(n2415) );
  NAND U2584 ( .A(n12097), .B(n2415), .Z(n2416) );
  ANDN U2585 ( .B(n5536), .A(n12099), .Z(n2417) );
  NANDN U2586 ( .A(n2416), .B(n5537), .Z(n2418) );
  AND U2587 ( .A(n2417), .B(n2418), .Z(n2419) );
  NANDN U2588 ( .A(n2419), .B(n12101), .Z(n2420) );
  NAND U2589 ( .A(n12103), .B(n2420), .Z(n2421) );
  NANDN U2590 ( .A(n12105), .B(n2421), .Z(n4412) );
  NAND U2591 ( .A(n8798), .B(n8797), .Z(n2422) );
  AND U2592 ( .A(n8799), .B(n2422), .Z(n2423) );
  NAND U2593 ( .A(n2423), .B(n8800), .Z(n2424) );
  NANDN U2594 ( .A(n11939), .B(n5594), .Z(n2425) );
  ANDN U2595 ( .B(n2425), .A(n5595), .Z(n2426) );
  AND U2596 ( .A(n11937), .B(n8801), .Z(n2427) );
  NAND U2597 ( .A(n2424), .B(n2427), .Z(n2428) );
  NANDN U2598 ( .A(n2426), .B(n2428), .Z(n2429) );
  NAND U2599 ( .A(n11941), .B(n2429), .Z(n2430) );
  NANDN U2600 ( .A(n11943), .B(n2430), .Z(n2431) );
  AND U2601 ( .A(n11945), .B(n2431), .Z(n2432) );
  NANDN U2602 ( .A(n2432), .B(n11947), .Z(n2433) );
  AND U2603 ( .A(n11949), .B(n2433), .Z(n2434) );
  NANDN U2604 ( .A(n2434), .B(n11951), .Z(n2435) );
  NANDN U2605 ( .A(n11953), .B(n2435), .Z(n2436) );
  NAND U2606 ( .A(n11955), .B(n2436), .Z(n2437) );
  ANDN U2607 ( .B(n8802), .A(n11959), .Z(n2438) );
  NANDN U2608 ( .A(n11957), .B(n2437), .Z(n2439) );
  NAND U2609 ( .A(n2438), .B(n2439), .Z(n8804) );
  NAND U2610 ( .A(n8874), .B(n8873), .Z(n2440) );
  ANDN U2611 ( .B(n2440), .A(n8875), .Z(n2441) );
  ANDN U2612 ( .B(n8876), .A(n2441), .Z(n2442) );
  NANDN U2613 ( .A(y[918]), .B(x[918]), .Z(n2443) );
  NAND U2614 ( .A(n2442), .B(n2443), .Z(n2444) );
  NANDN U2615 ( .A(n8877), .B(n2444), .Z(n2445) );
  ANDN U2616 ( .B(n5550), .A(n12051), .Z(n2446) );
  OR U2617 ( .A(n2445), .B(n8878), .Z(n2447) );
  AND U2618 ( .A(n2446), .B(n2447), .Z(n2448) );
  NOR U2619 ( .A(n8880), .B(n2448), .Z(n2449) );
  NAND U2620 ( .A(n8879), .B(n2449), .Z(n2450) );
  AND U2621 ( .A(n12055), .B(n2450), .Z(n2451) );
  ANDN U2622 ( .B(n8881), .A(n2451), .Z(n2452) );
  NAND U2623 ( .A(n12056), .B(n2452), .Z(n2453) );
  AND U2624 ( .A(n8882), .B(n2453), .Z(n2454) );
  NAND U2625 ( .A(n2454), .B(n8883), .Z(n2455) );
  AND U2626 ( .A(n5547), .B(n2455), .Z(n2456) );
  NANDN U2627 ( .A(n5546), .B(n2456), .Z(n2457) );
  NAND U2628 ( .A(n12067), .B(n2457), .Z(n8886) );
  NOR U2629 ( .A(n5533), .B(n5532), .Z(n2458) );
  NAND U2630 ( .A(n2458), .B(n8912), .Z(n2459) );
  AND U2631 ( .A(n8914), .B(n2459), .Z(n2460) );
  NAND U2632 ( .A(n2460), .B(n8913), .Z(n2461) );
  NOR U2633 ( .A(n8916), .B(n8915), .Z(n2462) );
  NAND U2634 ( .A(n2461), .B(n2462), .Z(n2463) );
  NAND U2635 ( .A(n8917), .B(n2463), .Z(n2464) );
  OR U2636 ( .A(n8918), .B(n2464), .Z(n2465) );
  AND U2637 ( .A(n8919), .B(n2465), .Z(n2466) );
  NOR U2638 ( .A(n8922), .B(n8921), .Z(n2467) );
  NAND U2639 ( .A(n2466), .B(n8920), .Z(n2468) );
  AND U2640 ( .A(n2467), .B(n2468), .Z(n2469) );
  ANDN U2641 ( .B(n8923), .A(n2469), .Z(n2470) );
  NAND U2642 ( .A(n8924), .B(n2470), .Z(n2471) );
  ANDN U2643 ( .B(n2471), .A(n8925), .Z(n2472) );
  ANDN U2644 ( .B(n8926), .A(n12137), .Z(n2473) );
  NANDN U2645 ( .A(n12135), .B(n2472), .Z(n2474) );
  NAND U2646 ( .A(n2473), .B(n2474), .Z(n2475) );
  NAND U2647 ( .A(n12139), .B(n2475), .Z(n8927) );
  ANDN U2648 ( .B(n5512), .A(n5511), .Z(n2476) );
  ANDN U2649 ( .B(n8991), .A(n12222), .Z(n2477) );
  NAND U2650 ( .A(n8992), .B(n2477), .Z(n2478) );
  AND U2651 ( .A(n2476), .B(n2478), .Z(n2479) );
  NANDN U2652 ( .A(n2479), .B(n12231), .Z(n2480) );
  NAND U2653 ( .A(n12232), .B(n2480), .Z(n2481) );
  NAND U2654 ( .A(n12235), .B(n2481), .Z(n2482) );
  AND U2655 ( .A(n8995), .B(n12237), .Z(n2483) );
  NAND U2656 ( .A(n2482), .B(n2483), .Z(n2484) );
  NAND U2657 ( .A(n8996), .B(n2484), .Z(n2485) );
  NOR U2658 ( .A(n8998), .B(n8997), .Z(n2486) );
  NANDN U2659 ( .A(n2485), .B(n12238), .Z(n2487) );
  AND U2660 ( .A(n2486), .B(n2487), .Z(n2488) );
  ANDN U2661 ( .B(n8999), .A(n2488), .Z(n2489) );
  NAND U2662 ( .A(n9000), .B(n2489), .Z(n2490) );
  ANDN U2663 ( .B(n2490), .A(n9001), .Z(n2491) );
  NOR U2664 ( .A(n5506), .B(n5505), .Z(n2492) );
  NANDN U2665 ( .A(n9002), .B(n2491), .Z(n2493) );
  NAND U2666 ( .A(n2492), .B(n2493), .Z(n9006) );
  ANDN U2667 ( .B(n9105), .A(n12414), .Z(n2494) );
  OR U2668 ( .A(n12413), .B(n4436), .Z(n2495) );
  AND U2669 ( .A(n2494), .B(n2495), .Z(n2496) );
  NAND U2670 ( .A(n12422), .B(n9104), .Z(n2497) );
  NOR U2671 ( .A(n2496), .B(n9103), .Z(n2498) );
  NAND U2672 ( .A(n12421), .B(n2498), .Z(n2499) );
  NANDN U2673 ( .A(n2497), .B(n2499), .Z(n2500) );
  AND U2674 ( .A(n12427), .B(n5441), .Z(n2501) );
  NANDN U2675 ( .A(n12425), .B(n2500), .Z(n2502) );
  NAND U2676 ( .A(n2501), .B(n2502), .Z(n2503) );
  ANDN U2677 ( .B(n12428), .A(n9109), .Z(n2504) );
  NAND U2678 ( .A(n2503), .B(n2504), .Z(n2505) );
  NAND U2679 ( .A(n5442), .B(n2505), .Z(n2506) );
  NANDN U2680 ( .A(n2506), .B(n9111), .Z(n2507) );
  ANDN U2681 ( .B(n2507), .A(n12436), .Z(n2508) );
  ANDN U2682 ( .B(n9112), .A(n12441), .Z(n2509) );
  NANDN U2683 ( .A(n9110), .B(n2508), .Z(n2510) );
  NAND U2684 ( .A(n2509), .B(n2510), .Z(n4437) );
  NANDN U2685 ( .A(n12299), .B(n9036), .Z(n2511) );
  AND U2686 ( .A(n12301), .B(n2511), .Z(n2512) );
  OR U2687 ( .A(n2512), .B(n12303), .Z(n2513) );
  NAND U2688 ( .A(n12305), .B(n2513), .Z(n2514) );
  NANDN U2689 ( .A(n12307), .B(n2514), .Z(n2515) );
  NAND U2690 ( .A(n12310), .B(n12315), .Z(n2516) );
  ANDN U2691 ( .B(n9037), .A(n12308), .Z(n2517) );
  NAND U2692 ( .A(n2515), .B(n2517), .Z(n2518) );
  NANDN U2693 ( .A(n2516), .B(n2518), .Z(n2519) );
  AND U2694 ( .A(n9038), .B(n12316), .Z(n2520) );
  NAND U2695 ( .A(n2519), .B(n2520), .Z(n2521) );
  NANDN U2696 ( .A(n12319), .B(n2521), .Z(n2522) );
  NAND U2697 ( .A(n12321), .B(n2522), .Z(n2523) );
  NAND U2698 ( .A(n12322), .B(n2523), .Z(n2524) );
  AND U2699 ( .A(n12325), .B(n2524), .Z(n2525) );
  NANDN U2700 ( .A(n2525), .B(n12327), .Z(n2526) );
  AND U2701 ( .A(n9039), .B(n2526), .Z(n9040) );
  NAND U2702 ( .A(n4446), .B(n12582), .Z(n2527) );
  NANDN U2703 ( .A(n12585), .B(n2527), .Z(n2528) );
  AND U2704 ( .A(n12587), .B(n2528), .Z(n2529) );
  NANDN U2705 ( .A(n2529), .B(n12589), .Z(n2530) );
  NANDN U2706 ( .A(n12591), .B(n2530), .Z(n2531) );
  NANDN U2707 ( .A(n12592), .B(n2531), .Z(n2532) );
  OR U2708 ( .A(n2532), .B(n10188), .Z(n2533) );
  NANDN U2709 ( .A(n12595), .B(n2533), .Z(n2534) );
  NANDN U2710 ( .A(n10190), .B(n2534), .Z(n2535) );
  NAND U2711 ( .A(n12599), .B(n2535), .Z(n2536) );
  ANDN U2712 ( .B(n2536), .A(n12601), .Z(n2537) );
  NANDN U2713 ( .A(n5407), .B(n2537), .Z(n2538) );
  AND U2714 ( .A(n9173), .B(n2538), .Z(n2539) );
  NANDN U2715 ( .A(n5404), .B(n2539), .Z(n4447) );
  ANDN U2716 ( .B(n5440), .A(n5439), .Z(n2540) );
  NANDN U2717 ( .A(n9118), .B(n9117), .Z(n2541) );
  AND U2718 ( .A(n2540), .B(n2541), .Z(n2542) );
  ANDN U2719 ( .B(n5436), .A(n12454), .Z(n2543) );
  OR U2720 ( .A(n12452), .B(n2542), .Z(n2544) );
  AND U2721 ( .A(n2543), .B(n2544), .Z(n2545) );
  ANDN U2722 ( .B(n5435), .A(n5434), .Z(n2546) );
  ANDN U2723 ( .B(n12461), .A(n2545), .Z(n2547) );
  NAND U2724 ( .A(n12457), .B(n2547), .Z(n2548) );
  AND U2725 ( .A(n2546), .B(n2548), .Z(n2549) );
  AND U2726 ( .A(n5433), .B(n12467), .Z(n2550) );
  OR U2727 ( .A(n12465), .B(n2549), .Z(n2551) );
  AND U2728 ( .A(n2550), .B(n2551), .Z(n2552) );
  ANDN U2729 ( .B(n5432), .A(n5431), .Z(n2553) );
  ANDN U2730 ( .B(n12473), .A(n2552), .Z(n2554) );
  NAND U2731 ( .A(n12468), .B(n2554), .Z(n2555) );
  AND U2732 ( .A(n2553), .B(n2555), .Z(n9124) );
  AND U2733 ( .A(n12685), .B(n5380), .Z(n2556) );
  NANDN U2734 ( .A(n4452), .B(n4451), .Z(n2557) );
  NAND U2735 ( .A(n12659), .B(n2557), .Z(n2558) );
  AND U2736 ( .A(n12661), .B(n2558), .Z(n2559) );
  NANDN U2737 ( .A(n2559), .B(n12663), .Z(n2560) );
  NAND U2738 ( .A(n12665), .B(n2560), .Z(n2561) );
  NANDN U2739 ( .A(n12667), .B(n2561), .Z(n2562) );
  NAND U2740 ( .A(n12669), .B(n2562), .Z(n2563) );
  NANDN U2741 ( .A(n12671), .B(n2563), .Z(n2564) );
  AND U2742 ( .A(n5384), .B(n2564), .Z(n2565) );
  NAND U2743 ( .A(n2565), .B(n12673), .Z(n2566) );
  AND U2744 ( .A(n12679), .B(n2566), .Z(n2567) );
  NANDN U2745 ( .A(n9197), .B(n2567), .Z(n2568) );
  ANDN U2746 ( .B(n5383), .A(n5382), .Z(n2569) );
  NAND U2747 ( .A(n2568), .B(n2569), .Z(n2570) );
  NANDN U2748 ( .A(n12683), .B(n2570), .Z(n2571) );
  NAND U2749 ( .A(n2556), .B(n2571), .Z(n4453) );
  NANDN U2750 ( .A(n12537), .B(n12541), .Z(n2572) );
  ANDN U2751 ( .B(n9146), .A(n9145), .Z(n2573) );
  NAND U2752 ( .A(n9144), .B(n12533), .Z(n2574) );
  AND U2753 ( .A(n2573), .B(n2574), .Z(n2575) );
  ANDN U2754 ( .B(n12542), .A(n9147), .Z(n2576) );
  OR U2755 ( .A(n2572), .B(n2575), .Z(n2577) );
  AND U2756 ( .A(n2576), .B(n2577), .Z(n2578) );
  NANDN U2757 ( .A(n2578), .B(n12545), .Z(n2579) );
  NANDN U2758 ( .A(n12547), .B(n2579), .Z(n2580) );
  NAND U2759 ( .A(n12549), .B(n2580), .Z(n2581) );
  ANDN U2760 ( .B(n2581), .A(n9148), .Z(n2582) );
  AND U2761 ( .A(n12553), .B(n12557), .Z(n2583) );
  NANDN U2762 ( .A(n12551), .B(n2582), .Z(n2584) );
  NAND U2763 ( .A(n2583), .B(n2584), .Z(n2585) );
  AND U2764 ( .A(n12558), .B(n9149), .Z(n2586) );
  NAND U2765 ( .A(n2585), .B(n2586), .Z(n2587) );
  NANDN U2766 ( .A(n12560), .B(n2587), .Z(n9152) );
  ANDN U2767 ( .B(n5353), .A(n12753), .Z(n2588) );
  NANDN U2768 ( .A(n4461), .B(n4460), .Z(n2589) );
  NAND U2769 ( .A(n2588), .B(n2589), .Z(n2590) );
  AND U2770 ( .A(n9221), .B(n12755), .Z(n2591) );
  NAND U2771 ( .A(n2590), .B(n2591), .Z(n2592) );
  NANDN U2772 ( .A(n5352), .B(n2592), .Z(n2593) );
  ANDN U2773 ( .B(n9223), .A(n9220), .Z(n2594) );
  OR U2774 ( .A(n2593), .B(n5350), .Z(n2595) );
  AND U2775 ( .A(n2594), .B(n2595), .Z(n2596) );
  ANDN U2776 ( .B(n5351), .A(n2596), .Z(n2597) );
  NAND U2777 ( .A(n9226), .B(n2597), .Z(n2598) );
  ANDN U2778 ( .B(n2598), .A(n9222), .Z(n2599) );
  NAND U2779 ( .A(n2599), .B(n12767), .Z(n2600) );
  AND U2780 ( .A(n9225), .B(n2600), .Z(n2601) );
  NANDN U2781 ( .A(n12768), .B(n2601), .Z(n4462) );
  NANDN U2782 ( .A(n9178), .B(n9177), .Z(n2602) );
  AND U2783 ( .A(n9179), .B(n2602), .Z(n2603) );
  ANDN U2784 ( .B(n5403), .A(n12619), .Z(n2604) );
  NANDN U2785 ( .A(n12617), .B(n2603), .Z(n2605) );
  AND U2786 ( .A(n2604), .B(n2605), .Z(n2606) );
  OR U2787 ( .A(n12621), .B(n2606), .Z(n2607) );
  NAND U2788 ( .A(n12623), .B(n2607), .Z(n2608) );
  NANDN U2789 ( .A(n12624), .B(n2608), .Z(n2609) );
  ANDN U2790 ( .B(n9180), .A(n12626), .Z(n2610) );
  NAND U2791 ( .A(n2609), .B(n2610), .Z(n2611) );
  NAND U2792 ( .A(n12628), .B(n2611), .Z(n2612) );
  ANDN U2793 ( .B(n9181), .A(n12635), .Z(n2613) );
  NANDN U2794 ( .A(n2612), .B(n12632), .Z(n2614) );
  AND U2795 ( .A(n2613), .B(n2614), .Z(n2615) );
  OR U2796 ( .A(n2615), .B(n12637), .Z(n2616) );
  AND U2797 ( .A(n12639), .B(n2616), .Z(n2617) );
  ANDN U2798 ( .B(n5394), .A(n12642), .Z(n2618) );
  OR U2799 ( .A(n12640), .B(n2617), .Z(n2619) );
  AND U2800 ( .A(n2618), .B(n2619), .Z(n9186) );
  NANDN U2801 ( .A(n4472), .B(n4471), .Z(n2620) );
  NANDN U2802 ( .A(n12823), .B(n2620), .Z(n2621) );
  AND U2803 ( .A(n5344), .B(n2621), .Z(n2622) );
  AND U2804 ( .A(n12826), .B(n12831), .Z(n2623) );
  NANDN U2805 ( .A(n12825), .B(n2622), .Z(n2624) );
  NAND U2806 ( .A(n2623), .B(n2624), .Z(n2625) );
  AND U2807 ( .A(n5345), .B(n12832), .Z(n2626) );
  NAND U2808 ( .A(n2625), .B(n2626), .Z(n2627) );
  NANDN U2809 ( .A(n12835), .B(n2627), .Z(n2628) );
  ANDN U2810 ( .B(n5342), .A(n12836), .Z(n2629) );
  NAND U2811 ( .A(n2628), .B(n2629), .Z(n2630) );
  NAND U2812 ( .A(n12842), .B(n2630), .Z(n2631) );
  ANDN U2813 ( .B(n5343), .A(n12845), .Z(n2632) );
  NANDN U2814 ( .A(n2631), .B(n12838), .Z(n2633) );
  AND U2815 ( .A(n2632), .B(n2633), .Z(n2634) );
  ANDN U2816 ( .B(n5341), .A(n12849), .Z(n2635) );
  OR U2817 ( .A(n2634), .B(n12847), .Z(n2636) );
  NAND U2818 ( .A(n2635), .B(n2636), .Z(n4473) );
  NANDN U2819 ( .A(x[840]), .B(y[840]), .Z(n2637) );
  AND U2820 ( .A(n5627), .B(n2637), .Z(n11871) );
  ANDN U2821 ( .B(n9205), .A(n12703), .Z(n2638) );
  NANDN U2822 ( .A(n9204), .B(n12700), .Z(n2639) );
  NAND U2823 ( .A(n2638), .B(n2639), .Z(n2640) );
  NANDN U2824 ( .A(n12705), .B(n2640), .Z(n2641) );
  NAND U2825 ( .A(n12707), .B(n2641), .Z(n2642) );
  AND U2826 ( .A(n12709), .B(n2642), .Z(n2643) );
  NANDN U2827 ( .A(n2643), .B(n12711), .Z(n2644) );
  AND U2828 ( .A(n12713), .B(n2644), .Z(n2645) );
  NANDN U2829 ( .A(n2645), .B(n12715), .Z(n2646) );
  NANDN U2830 ( .A(n12716), .B(n2646), .Z(n2647) );
  NAND U2831 ( .A(n9208), .B(n2647), .Z(n2648) );
  AND U2832 ( .A(n5363), .B(n12722), .Z(n2649) );
  NANDN U2833 ( .A(n12718), .B(n2648), .Z(n2650) );
  NAND U2834 ( .A(n2649), .B(n2650), .Z(n2651) );
  NAND U2835 ( .A(n12725), .B(n2651), .Z(n2652) );
  AND U2836 ( .A(n12731), .B(n2652), .Z(n2653) );
  NANDN U2837 ( .A(n9209), .B(n2653), .Z(n9210) );
  OR U2838 ( .A(n9230), .B(n9231), .Z(n2654) );
  AND U2839 ( .A(n9232), .B(n2654), .Z(n2655) );
  NOR U2840 ( .A(n9234), .B(n12789), .Z(n2656) );
  NAND U2841 ( .A(n2655), .B(n9233), .Z(n2657) );
  AND U2842 ( .A(n2656), .B(n2657), .Z(n2658) );
  ANDN U2843 ( .B(n9235), .A(n2658), .Z(n2659) );
  NAND U2844 ( .A(n12791), .B(n2659), .Z(n2660) );
  ANDN U2845 ( .B(n2660), .A(n12792), .Z(n2661) );
  ANDN U2846 ( .B(n9236), .A(n2661), .Z(n2662) );
  NAND U2847 ( .A(n12794), .B(n2662), .Z(n2663) );
  ANDN U2848 ( .B(n2663), .A(n12797), .Z(n2664) );
  NAND U2849 ( .A(n2664), .B(n12801), .Z(n2665) );
  AND U2850 ( .A(n9237), .B(n2665), .Z(n2666) );
  NAND U2851 ( .A(n2666), .B(n12803), .Z(n2667) );
  NANDN U2852 ( .A(n12805), .B(n2667), .Z(n9244) );
  NANDN U2853 ( .A(n4480), .B(n4479), .Z(n2668) );
  NAND U2854 ( .A(n12921), .B(n2668), .Z(n2669) );
  NANDN U2855 ( .A(n12923), .B(n2669), .Z(n2670) );
  AND U2856 ( .A(n9275), .B(n12925), .Z(n2671) );
  NAND U2857 ( .A(n2670), .B(n2671), .Z(n2672) );
  NANDN U2858 ( .A(n12926), .B(n2672), .Z(n2673) );
  OR U2859 ( .A(n5313), .B(n2673), .Z(n2674) );
  AND U2860 ( .A(n5315), .B(n2674), .Z(n2675) );
  NAND U2861 ( .A(n2675), .B(n5312), .Z(n2676) );
  AND U2862 ( .A(n5314), .B(n2676), .Z(n2677) );
  NANDN U2863 ( .A(n5310), .B(n2677), .Z(n2678) );
  AND U2864 ( .A(n5308), .B(n5311), .Z(n2679) );
  NAND U2865 ( .A(n2678), .B(n2679), .Z(n2680) );
  NANDN U2866 ( .A(n5309), .B(n2680), .Z(n4482) );
  NAND U2867 ( .A(n9259), .B(n12854), .Z(n2681) );
  ANDN U2868 ( .B(n2681), .A(n12857), .Z(n2682) );
  ANDN U2869 ( .B(n9260), .A(n12863), .Z(n2683) );
  NAND U2870 ( .A(n2682), .B(n12861), .Z(n2684) );
  AND U2871 ( .A(n2683), .B(n2684), .Z(n2685) );
  OR U2872 ( .A(n12865), .B(n2685), .Z(n2686) );
  NAND U2873 ( .A(n12867), .B(n2686), .Z(n2687) );
  NAND U2874 ( .A(n12869), .B(n2687), .Z(n2688) );
  ANDN U2875 ( .B(n9263), .A(n12870), .Z(n2689) );
  NAND U2876 ( .A(n2688), .B(n2689), .Z(n2690) );
  NAND U2877 ( .A(n12872), .B(n2690), .Z(n2691) );
  ANDN U2878 ( .B(n5335), .A(n12879), .Z(n2692) );
  NANDN U2879 ( .A(n2691), .B(n12876), .Z(n2693) );
  AND U2880 ( .A(n2692), .B(n2693), .Z(n2694) );
  ANDN U2881 ( .B(n5332), .A(n12883), .Z(n2695) );
  OR U2882 ( .A(n12881), .B(n2694), .Z(n2696) );
  AND U2883 ( .A(n2695), .B(n2696), .Z(n9264) );
  NANDN U2884 ( .A(n3451), .B(n8964), .Z(n2697) );
  ANDN U2885 ( .B(n2697), .A(n8967), .Z(n12169) );
  NAND U2886 ( .A(n9278), .B(n12945), .Z(n2698) );
  NANDN U2887 ( .A(n9279), .B(n2698), .Z(n2699) );
  NAND U2888 ( .A(n9280), .B(n2699), .Z(n2700) );
  ANDN U2889 ( .B(n2700), .A(n9281), .Z(n2701) );
  AND U2890 ( .A(n5301), .B(n5302), .Z(n2702) );
  NANDN U2891 ( .A(n9282), .B(n2701), .Z(n2703) );
  NAND U2892 ( .A(n2702), .B(n2703), .Z(n2704) );
  AND U2893 ( .A(n9283), .B(n9284), .Z(n2705) );
  NAND U2894 ( .A(n2704), .B(n2705), .Z(n2706) );
  NANDN U2895 ( .A(n9285), .B(n2706), .Z(n2707) );
  OR U2896 ( .A(n9286), .B(n2707), .Z(n2708) );
  AND U2897 ( .A(n9287), .B(n2708), .Z(n2709) );
  NAND U2898 ( .A(n2709), .B(n9288), .Z(n2710) );
  AND U2899 ( .A(n12960), .B(n2710), .Z(n2711) );
  NANDN U2900 ( .A(n9289), .B(n2711), .Z(n2712) );
  AND U2901 ( .A(n12963), .B(n9290), .Z(n2713) );
  NAND U2902 ( .A(n2712), .B(n2713), .Z(n2714) );
  NANDN U2903 ( .A(n12964), .B(n2714), .Z(n9293) );
  NOR U2904 ( .A(n13066), .B(n5267), .Z(n2715) );
  NANDN U2905 ( .A(n4498), .B(n4497), .Z(n2716) );
  AND U2906 ( .A(n2715), .B(n2716), .Z(n2717) );
  ANDN U2907 ( .B(n5266), .A(n2717), .Z(n2718) );
  NAND U2908 ( .A(n5269), .B(n2718), .Z(n2719) );
  ANDN U2909 ( .B(n2719), .A(n13075), .Z(n2720) );
  NAND U2910 ( .A(n2720), .B(n5268), .Z(n2721) );
  AND U2911 ( .A(n13077), .B(n2721), .Z(n2722) );
  NAND U2912 ( .A(n2722), .B(n5265), .Z(n2723) );
  AND U2913 ( .A(n5262), .B(n13080), .Z(n2724) );
  NANDN U2914 ( .A(n13078), .B(n2723), .Z(n2725) );
  NAND U2915 ( .A(n2724), .B(n2725), .Z(n2726) );
  NANDN U2916 ( .A(n13083), .B(n2726), .Z(n4499) );
  NANDN U2917 ( .A(n9026), .B(n9021), .Z(n2727) );
  AND U2918 ( .A(n9028), .B(n2727), .Z(n2728) );
  NOR U2919 ( .A(n9025), .B(n9030), .Z(n2729) );
  NANDN U2920 ( .A(n3447), .B(n2728), .Z(n2730) );
  AND U2921 ( .A(n2729), .B(n2730), .Z(n12277) );
  OR U2922 ( .A(n4429), .B(n9085), .Z(n2731) );
  AND U2923 ( .A(n9089), .B(n2731), .Z(n12377) );
  NAND U2924 ( .A(n4504), .B(n4503), .Z(n2732) );
  NAND U2925 ( .A(n5244), .B(n2732), .Z(n2733) );
  NAND U2926 ( .A(n13157), .B(n2733), .Z(n2734) );
  NOR U2927 ( .A(n5240), .B(n13159), .Z(n2735) );
  NAND U2928 ( .A(n2734), .B(n2735), .Z(n2736) );
  NAND U2929 ( .A(n5238), .B(n2736), .Z(n2737) );
  NANDN U2930 ( .A(n2737), .B(n13161), .Z(n2738) );
  AND U2931 ( .A(n5239), .B(n2738), .Z(n2739) );
  XNOR U2932 ( .A(y[1380]), .B(x[1380]), .Z(n2740) );
  NAND U2933 ( .A(n2739), .B(n2740), .Z(n2741) );
  NAND U2934 ( .A(n5237), .B(n2741), .Z(n2742) );
  NAND U2935 ( .A(n5236), .B(n2742), .Z(n2743) );
  NANDN U2936 ( .A(n13169), .B(n2743), .Z(n2744) );
  ANDN U2937 ( .B(n2744), .A(n9368), .Z(n2745) );
  NANDN U2938 ( .A(n2745), .B(n9370), .Z(n2746) );
  NANDN U2939 ( .A(n5234), .B(n2746), .Z(n2747) );
  NAND U2940 ( .A(n13177), .B(n2747), .Z(n2748) );
  AND U2941 ( .A(n13179), .B(n2748), .Z(n4507) );
  NAND U2942 ( .A(n9345), .B(n13087), .Z(n2749) );
  NANDN U2943 ( .A(n13088), .B(n2749), .Z(n2750) );
  AND U2944 ( .A(n13090), .B(n2750), .Z(n2751) );
  NANDN U2945 ( .A(n2751), .B(n13093), .Z(n2752) );
  ANDN U2946 ( .B(n2752), .A(n13095), .Z(n2753) );
  ANDN U2947 ( .B(n5253), .A(n13099), .Z(n2754) );
  NANDN U2948 ( .A(n2753), .B(n13097), .Z(n2755) );
  AND U2949 ( .A(n2754), .B(n2755), .Z(n2756) );
  NOR U2950 ( .A(n9346), .B(n13105), .Z(n2757) );
  NANDN U2951 ( .A(n2756), .B(n13101), .Z(n2758) );
  AND U2952 ( .A(n2757), .B(n2758), .Z(n2759) );
  AND U2953 ( .A(n13109), .B(n13113), .Z(n2760) );
  OR U2954 ( .A(n9347), .B(n2759), .Z(n2761) );
  AND U2955 ( .A(n2760), .B(n2761), .Z(n2762) );
  NOR U2956 ( .A(n2762), .B(n5252), .Z(n2763) );
  NAND U2957 ( .A(n13115), .B(n2763), .Z(n2764) );
  AND U2958 ( .A(n13116), .B(n2764), .Z(n9352) );
  AND U2959 ( .A(n13236), .B(n13240), .Z(n2765) );
  NAND U2960 ( .A(n4510), .B(n9394), .Z(n2766) );
  AND U2961 ( .A(n2765), .B(n2766), .Z(n2767) );
  NOR U2962 ( .A(n13243), .B(n2767), .Z(n2768) );
  NAND U2963 ( .A(n9393), .B(n2768), .Z(n2769) );
  ANDN U2964 ( .B(n2769), .A(n13245), .Z(n2770) );
  ANDN U2965 ( .B(n9397), .A(n2770), .Z(n2771) );
  NAND U2966 ( .A(n13247), .B(n2771), .Z(n2772) );
  ANDN U2967 ( .B(n2772), .A(n13253), .Z(n2773) );
  AND U2968 ( .A(n9396), .B(n13255), .Z(n2774) );
  NANDN U2969 ( .A(n13249), .B(n2773), .Z(n2775) );
  NAND U2970 ( .A(n2774), .B(n2775), .Z(n2776) );
  ANDN U2971 ( .B(n13259), .A(n9400), .Z(n2777) );
  NANDN U2972 ( .A(n13257), .B(n2776), .Z(n2778) );
  NAND U2973 ( .A(n2777), .B(n2778), .Z(n2779) );
  AND U2974 ( .A(n13260), .B(n2779), .Z(n4513) );
  NAND U2975 ( .A(n9373), .B(n13182), .Z(n2780) );
  ANDN U2976 ( .B(n2780), .A(n13185), .Z(n2781) );
  NOR U2977 ( .A(n13189), .B(n9374), .Z(n2782) );
  NANDN U2978 ( .A(n2781), .B(n13187), .Z(n2783) );
  NAND U2979 ( .A(n2782), .B(n2783), .Z(n2784) );
  AND U2980 ( .A(n13191), .B(n13195), .Z(n2785) );
  NAND U2981 ( .A(n2784), .B(n2785), .Z(n2786) );
  NANDN U2982 ( .A(n9375), .B(n2786), .Z(n2787) );
  OR U2983 ( .A(n2787), .B(n13197), .Z(n2788) );
  NAND U2984 ( .A(n13199), .B(n2788), .Z(n2789) );
  NANDN U2985 ( .A(n13200), .B(n2789), .Z(n2790) );
  ANDN U2986 ( .B(n9378), .A(n13202), .Z(n2791) );
  NAND U2987 ( .A(n2790), .B(n2791), .Z(n2792) );
  NAND U2988 ( .A(n9379), .B(n2792), .Z(n2793) );
  OR U2989 ( .A(n9380), .B(n2793), .Z(n2794) );
  ANDN U2990 ( .B(n2794), .A(n9381), .Z(n2795) );
  AND U2991 ( .A(n9384), .B(n9383), .Z(n2796) );
  NANDN U2992 ( .A(n9382), .B(n2795), .Z(n2797) );
  NAND U2993 ( .A(n2796), .B(n2797), .Z(n9385) );
  NAND U2994 ( .A(n9411), .B(n9412), .Z(n2798) );
  NAND U2995 ( .A(n13268), .B(n2798), .Z(n2799) );
  NANDN U2996 ( .A(n13271), .B(n2799), .Z(n2800) );
  NAND U2997 ( .A(n13274), .B(n9413), .Z(n2801) );
  AND U2998 ( .A(n5207), .B(n13273), .Z(n2802) );
  NAND U2999 ( .A(n2800), .B(n2802), .Z(n2803) );
  NANDN U3000 ( .A(n2801), .B(n2803), .Z(n2804) );
  AND U3001 ( .A(n5205), .B(n5206), .Z(n2805) );
  NAND U3002 ( .A(n2805), .B(n2804), .Z(n2806) );
  AND U3003 ( .A(n5204), .B(n2806), .Z(n2807) );
  NAND U3004 ( .A(n2807), .B(n5203), .Z(n2808) );
  AND U3005 ( .A(n5202), .B(n5201), .Z(n2809) );
  NAND U3006 ( .A(n2809), .B(n2808), .Z(n2810) );
  AND U3007 ( .A(n13286), .B(n2810), .Z(n2811) );
  NAND U3008 ( .A(n2811), .B(n9414), .Z(n2812) );
  ANDN U3009 ( .B(n13288), .A(n9415), .Z(n2813) );
  NAND U3010 ( .A(n2812), .B(n2813), .Z(n2814) );
  NAND U3011 ( .A(n13291), .B(n2814), .Z(n9416) );
  AND U3012 ( .A(n3344), .B(n4521), .Z(n2815) );
  NAND U3013 ( .A(n5186), .B(n2815), .Z(n2816) );
  AND U3014 ( .A(n5189), .B(n2816), .Z(n2817) );
  NOR U3015 ( .A(n5187), .B(n5183), .Z(n2818) );
  NAND U3016 ( .A(n5185), .B(n2817), .Z(n2819) );
  AND U3017 ( .A(n2818), .B(n2819), .Z(n2820) );
  NOR U3018 ( .A(n2820), .B(n5184), .Z(n2821) );
  NAND U3019 ( .A(n5181), .B(n2821), .Z(n2822) );
  NAND U3020 ( .A(n5182), .B(n2822), .Z(n2823) );
  NANDN U3021 ( .A(n2823), .B(n9431), .Z(n2824) );
  ANDN U3022 ( .B(n2824), .A(n5180), .Z(n2825) );
  NOR U3023 ( .A(n9430), .B(n5178), .Z(n2826) );
  NANDN U3024 ( .A(n9432), .B(n2825), .Z(n2827) );
  NAND U3025 ( .A(n2826), .B(n2827), .Z(n4522) );
  ANDN U3026 ( .B(n9434), .A(n9435), .Z(n2828) );
  NAND U3027 ( .A(n9436), .B(n2828), .Z(n2829) );
  NAND U3028 ( .A(n9437), .B(n2829), .Z(n2830) );
  AND U3029 ( .A(n5177), .B(n5176), .Z(n2831) );
  OR U3030 ( .A(n2830), .B(n9438), .Z(n2832) );
  AND U3031 ( .A(n2831), .B(n2832), .Z(n2833) );
  NOR U3032 ( .A(n13365), .B(n9439), .Z(n2834) );
  NANDN U3033 ( .A(n2833), .B(n2834), .Z(n2835) );
  AND U3034 ( .A(n13367), .B(n2835), .Z(n2836) );
  NANDN U3035 ( .A(n9440), .B(n2836), .Z(n2837) );
  NAND U3036 ( .A(n13369), .B(n2837), .Z(n2838) );
  ANDN U3037 ( .B(n2838), .A(n13370), .Z(n2839) );
  NANDN U3038 ( .A(n2839), .B(n13373), .Z(n2840) );
  ANDN U3039 ( .B(n2840), .A(n13375), .Z(n2841) );
  OR U3040 ( .A(n13376), .B(n2841), .Z(n2842) );
  NAND U3041 ( .A(n13378), .B(n2842), .Z(n2843) );
  NANDN U3042 ( .A(n13381), .B(n2843), .Z(n9445) );
  NAND U3043 ( .A(n13012), .B(n5285), .Z(n13009) );
  ANDN U3044 ( .B(n13541), .A(n13537), .Z(n2844) );
  NAND U3045 ( .A(n13535), .B(n4563), .Z(n2845) );
  AND U3046 ( .A(n2844), .B(n2845), .Z(n2846) );
  NOR U3047 ( .A(n13542), .B(n2846), .Z(n2847) );
  NAND U3048 ( .A(n13538), .B(n2847), .Z(n2848) );
  ANDN U3049 ( .B(n2848), .A(n13544), .Z(n2849) );
  ANDN U3050 ( .B(n10187), .A(n2849), .Z(n2850) );
  NAND U3051 ( .A(n9487), .B(n2850), .Z(n2851) );
  ANDN U3052 ( .B(n2851), .A(n5111), .Z(n2852) );
  ANDN U3053 ( .B(n9488), .A(n2852), .Z(n2853) );
  NAND U3054 ( .A(n5109), .B(n2853), .Z(n2854) );
  ANDN U3055 ( .B(n2854), .A(n5112), .Z(n2855) );
  ANDN U3056 ( .B(n5110), .A(n13555), .Z(n2856) );
  NANDN U3057 ( .A(n5107), .B(n2855), .Z(n2857) );
  NAND U3058 ( .A(n2856), .B(n2857), .Z(n4564) );
  AND U3059 ( .A(n13585), .B(n5091), .Z(n2858) );
  NANDN U3060 ( .A(n9516), .B(n9515), .Z(n2859) );
  AND U3061 ( .A(n2858), .B(n2859), .Z(n2860) );
  NANDN U3062 ( .A(n2860), .B(n13587), .Z(n2861) );
  NANDN U3063 ( .A(n13589), .B(n2861), .Z(n2862) );
  NAND U3064 ( .A(n13591), .B(n2862), .Z(n2863) );
  NANDN U3065 ( .A(n13593), .B(n2863), .Z(n2864) );
  NANDN U3066 ( .A(n13595), .B(n2864), .Z(n2865) );
  AND U3067 ( .A(n9517), .B(n2865), .Z(n2866) );
  NAND U3068 ( .A(n2866), .B(n13597), .Z(n2867) );
  AND U3069 ( .A(n13602), .B(n2867), .Z(n2868) );
  NAND U3070 ( .A(n2868), .B(n13598), .Z(n2869) );
  ANDN U3071 ( .B(n5084), .A(n13605), .Z(n2870) );
  NAND U3072 ( .A(n2869), .B(n2870), .Z(n2871) );
  NAND U3073 ( .A(n13607), .B(n2871), .Z(n2872) );
  AND U3074 ( .A(n13609), .B(n2872), .Z(n9521) );
  NAND U3075 ( .A(n13643), .B(n4594), .Z(n2873) );
  AND U3076 ( .A(n13649), .B(n2873), .Z(n9530) );
  NAND U3077 ( .A(n13709), .B(n13713), .Z(n2874) );
  NAND U3078 ( .A(n9539), .B(n13699), .Z(n2875) );
  NAND U3079 ( .A(n9542), .B(n2875), .Z(n2876) );
  AND U3080 ( .A(n13702), .B(n2876), .Z(n2877) );
  AND U3081 ( .A(n13707), .B(n5055), .Z(n2878) );
  OR U3082 ( .A(n13705), .B(n2877), .Z(n2879) );
  AND U3083 ( .A(n2878), .B(n2879), .Z(n2880) );
  AND U3084 ( .A(n5054), .B(n13714), .Z(n2881) );
  OR U3085 ( .A(n2874), .B(n2880), .Z(n2882) );
  AND U3086 ( .A(n2881), .B(n2882), .Z(n2883) );
  OR U3087 ( .A(n13716), .B(n2883), .Z(n2884) );
  ANDN U3088 ( .B(n2884), .A(n13719), .Z(n2885) );
  AND U3089 ( .A(n9544), .B(n13723), .Z(n2886) );
  NANDN U3090 ( .A(n2885), .B(n9543), .Z(n2887) );
  NAND U3091 ( .A(n2886), .B(n2887), .Z(n9545) );
  ANDN U3092 ( .B(n9551), .A(n13751), .Z(n2888) );
  NANDN U3093 ( .A(n13749), .B(n4602), .Z(n2889) );
  AND U3094 ( .A(n2888), .B(n2889), .Z(n2890) );
  NOR U3095 ( .A(n5041), .B(n2890), .Z(n2891) );
  NAND U3096 ( .A(n13753), .B(n2891), .Z(n2892) );
  AND U3097 ( .A(n9552), .B(n2892), .Z(n2893) );
  NAND U3098 ( .A(n5038), .B(n2893), .Z(n2894) );
  ANDN U3099 ( .B(n2894), .A(n5037), .Z(n2895) );
  NANDN U3100 ( .A(n5040), .B(n2895), .Z(n2896) );
  AND U3101 ( .A(n5039), .B(n2896), .Z(n2897) );
  XNOR U3102 ( .A(x[1634]), .B(y[1634]), .Z(n2898) );
  AND U3103 ( .A(n2897), .B(n2898), .Z(n2899) );
  NANDN U3104 ( .A(n2899), .B(n5036), .Z(n2900) );
  AND U3105 ( .A(n5035), .B(n2900), .Z(n2901) );
  NANDN U3106 ( .A(n2901), .B(n9553), .Z(n2902) );
  NANDN U3107 ( .A(n9555), .B(n2902), .Z(n2903) );
  NANDN U3108 ( .A(n13771), .B(n2903), .Z(n4604) );
  OR U3109 ( .A(n3324), .B(n9450), .Z(n2904) );
  AND U3110 ( .A(n9454), .B(n2904), .Z(n13410) );
  NOR U3111 ( .A(n13783), .B(n9560), .Z(n2905) );
  NAND U3112 ( .A(n9559), .B(n2905), .Z(n2906) );
  AND U3113 ( .A(n9561), .B(n2906), .Z(n2907) );
  NAND U3114 ( .A(n13789), .B(n2907), .Z(n2908) );
  ANDN U3115 ( .B(n2908), .A(n9562), .Z(n2909) );
  NANDN U3116 ( .A(n9563), .B(n2909), .Z(n2910) );
  NAND U3117 ( .A(n13795), .B(n2910), .Z(n2911) );
  AND U3118 ( .A(n13794), .B(n2911), .Z(n2912) );
  NAND U3119 ( .A(n2912), .B(n5023), .Z(n2913) );
  AND U3120 ( .A(n5022), .B(n13792), .Z(n2914) );
  NAND U3121 ( .A(n2913), .B(n2914), .Z(n2915) );
  NANDN U3122 ( .A(n9564), .B(n2915), .Z(n2916) );
  AND U3123 ( .A(n5020), .B(n5021), .Z(n2917) );
  OR U3124 ( .A(n2916), .B(n9565), .Z(n2918) );
  AND U3125 ( .A(n2917), .B(n2918), .Z(n2919) );
  ANDN U3126 ( .B(n5019), .A(n2919), .Z(n2920) );
  NAND U3127 ( .A(n5018), .B(n2920), .Z(n2921) );
  AND U3128 ( .A(n9566), .B(n2921), .Z(n9567) );
  NANDN U3129 ( .A(n5145), .B(n5143), .Z(n2922) );
  ANDN U3130 ( .B(n2922), .A(n5144), .Z(n13471) );
  NANDN U3131 ( .A(n4609), .B(n4608), .Z(n2923) );
  NAND U3132 ( .A(n13849), .B(n2923), .Z(n2924) );
  ANDN U3133 ( .B(n2924), .A(n13850), .Z(n2925) );
  NANDN U3134 ( .A(n2925), .B(n13852), .Z(n2926) );
  AND U3135 ( .A(n13855), .B(n2926), .Z(n2927) );
  OR U3136 ( .A(n9613), .B(n2927), .Z(n2928) );
  NAND U3137 ( .A(n13859), .B(n2928), .Z(n2929) );
  NAND U3138 ( .A(n9619), .B(n2929), .Z(n2930) );
  ANDN U3139 ( .B(n4996), .A(n9620), .Z(n2931) );
  NAND U3140 ( .A(n2930), .B(n2931), .Z(n2932) );
  NANDN U3141 ( .A(n13865), .B(n2932), .Z(n2933) );
  NANDN U3142 ( .A(n2933), .B(n4995), .Z(n2934) );
  ANDN U3143 ( .B(n2934), .A(n13871), .Z(n2935) );
  AND U3144 ( .A(n13873), .B(n4994), .Z(n2936) );
  NANDN U3145 ( .A(n4997), .B(n2935), .Z(n2937) );
  NAND U3146 ( .A(n2936), .B(n2937), .Z(n4610) );
  OR U3147 ( .A(n13887), .B(n9630), .Z(n2938) );
  NAND U3148 ( .A(n13889), .B(n2938), .Z(n2939) );
  ANDN U3149 ( .B(n2939), .A(n13891), .Z(n2940) );
  NANDN U3150 ( .A(n2940), .B(n13893), .Z(n2941) );
  NANDN U3151 ( .A(n13895), .B(n2941), .Z(n2942) );
  NAND U3152 ( .A(n9631), .B(n2942), .Z(n2943) );
  AND U3153 ( .A(n13898), .B(n4991), .Z(n2944) );
  OR U3154 ( .A(n2943), .B(n13896), .Z(n2945) );
  AND U3155 ( .A(n2944), .B(n2945), .Z(n2946) );
  NOR U3156 ( .A(n9632), .B(n2946), .Z(n2947) );
  NAND U3157 ( .A(n10185), .B(n2947), .Z(n2948) );
  AND U3158 ( .A(n9633), .B(n2948), .Z(n2949) );
  NANDN U3159 ( .A(n9634), .B(n2949), .Z(n2950) );
  NANDN U3160 ( .A(n9635), .B(n2950), .Z(n2951) );
  ANDN U3161 ( .B(n2951), .A(n9636), .Z(n2952) );
  NANDN U3162 ( .A(n2952), .B(n9637), .Z(n2953) );
  NANDN U3163 ( .A(n9638), .B(n2953), .Z(n2954) );
  NAND U3164 ( .A(n13917), .B(n2954), .Z(n9641) );
  AND U3165 ( .A(n9648), .B(n4980), .Z(n2955) );
  NANDN U3166 ( .A(n4981), .B(n4639), .Z(n2956) );
  AND U3167 ( .A(n2955), .B(n2956), .Z(n2957) );
  NOR U3168 ( .A(n9652), .B(n2957), .Z(n2958) );
  NAND U3169 ( .A(n4982), .B(n2958), .Z(n2959) );
  ANDN U3170 ( .B(n2959), .A(n13947), .Z(n2960) );
  NAND U3171 ( .A(n2960), .B(n4979), .Z(n2961) );
  NANDN U3172 ( .A(n13949), .B(n2961), .Z(n2962) );
  AND U3173 ( .A(n13951), .B(n2962), .Z(n2963) );
  OR U3174 ( .A(n13953), .B(n2963), .Z(n2964) );
  AND U3175 ( .A(n13955), .B(n2964), .Z(n2965) );
  OR U3176 ( .A(n13957), .B(n2965), .Z(n2966) );
  NAND U3177 ( .A(n13959), .B(n2966), .Z(n2967) );
  NAND U3178 ( .A(n13961), .B(n2967), .Z(n2968) );
  NOR U3179 ( .A(n9661), .B(n13963), .Z(n2969) );
  NAND U3180 ( .A(n2968), .B(n2969), .Z(n2970) );
  NAND U3181 ( .A(n9660), .B(n2970), .Z(n4641) );
  OR U3182 ( .A(n3281), .B(n9524), .Z(n2971) );
  ANDN U3183 ( .B(n2971), .A(n9525), .Z(n13629) );
  ANDN U3184 ( .B(n4970), .A(n4969), .Z(n2972) );
  NANDN U3185 ( .A(n9665), .B(n13969), .Z(n2973) );
  NAND U3186 ( .A(n2972), .B(n2973), .Z(n2974) );
  ANDN U3187 ( .B(n2974), .A(n9666), .Z(n2975) );
  AND U3188 ( .A(n4968), .B(n4967), .Z(n2976) );
  NANDN U3189 ( .A(n13973), .B(n2975), .Z(n2977) );
  NAND U3190 ( .A(n2976), .B(n2977), .Z(n2978) );
  NAND U3191 ( .A(n4964), .B(n4963), .Z(n2979) );
  AND U3192 ( .A(n4966), .B(n4965), .Z(n2980) );
  NAND U3193 ( .A(n2978), .B(n2980), .Z(n2981) );
  NANDN U3194 ( .A(n2979), .B(n2981), .Z(n2982) );
  ANDN U3195 ( .B(n9667), .A(n13985), .Z(n2983) );
  NAND U3196 ( .A(n2982), .B(n2983), .Z(n2984) );
  NANDN U3197 ( .A(n9668), .B(n2984), .Z(n2985) );
  OR U3198 ( .A(n13987), .B(n2985), .Z(n2986) );
  AND U3199 ( .A(n13989), .B(n2986), .Z(n2987) );
  OR U3200 ( .A(n13991), .B(n2987), .Z(n2988) );
  NAND U3201 ( .A(n13993), .B(n2988), .Z(n2989) );
  NANDN U3202 ( .A(n13995), .B(n2989), .Z(n9671) );
  AND U3203 ( .A(n14023), .B(n4948), .Z(n9684) );
  ANDN U3204 ( .B(n4936), .A(n4941), .Z(n2990) );
  NAND U3205 ( .A(n4644), .B(n2990), .Z(n2991) );
  AND U3206 ( .A(n14049), .B(n2991), .Z(n2992) );
  NAND U3207 ( .A(n4939), .B(n2992), .Z(n2993) );
  ANDN U3208 ( .B(n2993), .A(n4937), .Z(n2994) );
  NANDN U3209 ( .A(n14051), .B(n2994), .Z(n2995) );
  NAND U3210 ( .A(n14053), .B(n2995), .Z(n2996) );
  NANDN U3211 ( .A(n14055), .B(n2996), .Z(n2997) );
  AND U3212 ( .A(n14057), .B(n2997), .Z(n2998) );
  OR U3213 ( .A(n14059), .B(n2998), .Z(n2999) );
  NAND U3214 ( .A(n14061), .B(n2999), .Z(n3000) );
  NANDN U3215 ( .A(n14062), .B(n3000), .Z(n3001) );
  NAND U3216 ( .A(n14064), .B(n3001), .Z(n3002) );
  NAND U3217 ( .A(n14067), .B(n3002), .Z(n3003) );
  ANDN U3218 ( .B(n3003), .A(n4926), .Z(n4650) );
  ANDN U3219 ( .B(n4652), .A(n4912), .Z(n3004) );
  NAND U3220 ( .A(n14123), .B(n3004), .Z(n3005) );
  AND U3221 ( .A(n4911), .B(n3005), .Z(n3006) );
  NANDN U3222 ( .A(n14124), .B(n3006), .Z(n3007) );
  NANDN U3223 ( .A(n14127), .B(n3007), .Z(n3008) );
  AND U3224 ( .A(n14129), .B(n3008), .Z(n3009) );
  OR U3225 ( .A(n14131), .B(n3009), .Z(n3010) );
  NAND U3226 ( .A(n14133), .B(n3010), .Z(n3011) );
  NANDN U3227 ( .A(n14135), .B(n3011), .Z(n3012) );
  NAND U3228 ( .A(n10177), .B(n3012), .Z(n3013) );
  NANDN U3229 ( .A(n4903), .B(n3013), .Z(n3014) );
  ANDN U3230 ( .B(n3014), .A(n9781), .Z(n3015) );
  NANDN U3231 ( .A(n3015), .B(n14143), .Z(n3016) );
  NANDN U3232 ( .A(n14144), .B(n3016), .Z(n3017) );
  NAND U3233 ( .A(n14146), .B(n3017), .Z(n3018) );
  NANDN U3234 ( .A(n14149), .B(n3018), .Z(n4653) );
  AND U3235 ( .A(n9816), .B(n9815), .Z(n3019) );
  NAND U3236 ( .A(n9814), .B(n9813), .Z(n3020) );
  AND U3237 ( .A(n3019), .B(n3020), .Z(n3021) );
  ANDN U3238 ( .B(n4895), .A(n3021), .Z(n3022) );
  NAND U3239 ( .A(n4894), .B(n3022), .Z(n3023) );
  AND U3240 ( .A(n9817), .B(n3023), .Z(n3024) );
  ANDN U3241 ( .B(n9820), .A(n9819), .Z(n3025) );
  NANDN U3242 ( .A(n9818), .B(n3024), .Z(n3026) );
  NAND U3243 ( .A(n3025), .B(n3026), .Z(n3027) );
  NAND U3244 ( .A(n14188), .B(n3027), .Z(n3028) );
  NAND U3245 ( .A(n14191), .B(n3028), .Z(n3029) );
  AND U3246 ( .A(n14192), .B(n3029), .Z(n3030) );
  ANDN U3247 ( .B(n9826), .A(n9825), .Z(n3031) );
  NANDN U3248 ( .A(n3030), .B(n14195), .Z(n3032) );
  AND U3249 ( .A(n3031), .B(n3032), .Z(n3033) );
  NOR U3250 ( .A(n3033), .B(n9827), .Z(n3034) );
  NAND U3251 ( .A(n9828), .B(n3034), .Z(n3035) );
  AND U3252 ( .A(n9829), .B(n3035), .Z(n3036) );
  NANDN U3253 ( .A(n9830), .B(n3036), .Z(n9831) );
  NANDN U3254 ( .A(n14226), .B(n4658), .Z(n3037) );
  NAND U3255 ( .A(n14229), .B(n3037), .Z(n3038) );
  NANDN U3256 ( .A(n14230), .B(n3038), .Z(n3039) );
  NAND U3257 ( .A(n14233), .B(n3039), .Z(n3040) );
  NANDN U3258 ( .A(n14234), .B(n3040), .Z(n3041) );
  ANDN U3259 ( .B(n3041), .A(n14236), .Z(n3042) );
  NAND U3260 ( .A(n3042), .B(n4874), .Z(n3043) );
  AND U3261 ( .A(n4871), .B(n3043), .Z(n3044) );
  NANDN U3262 ( .A(n14239), .B(n3044), .Z(n3045) );
  AND U3263 ( .A(n4870), .B(n4873), .Z(n3046) );
  NAND U3264 ( .A(n3045), .B(n3046), .Z(n3047) );
  NANDN U3265 ( .A(n4867), .B(n3047), .Z(n3048) );
  OR U3266 ( .A(n4872), .B(n3048), .Z(n3049) );
  ANDN U3267 ( .B(n3049), .A(n9841), .Z(n3050) );
  NAND U3268 ( .A(n3050), .B(n4869), .Z(n3051) );
  AND U3269 ( .A(n4868), .B(n3051), .Z(n3052) );
  NAND U3270 ( .A(n3052), .B(n9844), .Z(n4660) );
  NAND U3271 ( .A(n9877), .B(n9876), .Z(n3053) );
  ANDN U3272 ( .B(n3053), .A(n9878), .Z(n3054) );
  NOR U3273 ( .A(n4853), .B(n4854), .Z(n3055) );
  NANDN U3274 ( .A(n9879), .B(n3054), .Z(n3056) );
  AND U3275 ( .A(n3055), .B(n3056), .Z(n3057) );
  NOR U3276 ( .A(n9880), .B(n3057), .Z(n3058) );
  NAND U3277 ( .A(n9881), .B(n3058), .Z(n3059) );
  ANDN U3278 ( .B(n3059), .A(n9882), .Z(n3060) );
  NAND U3279 ( .A(n3060), .B(n9883), .Z(n3061) );
  NAND U3280 ( .A(n14292), .B(n3061), .Z(n3062) );
  AND U3281 ( .A(n14295), .B(n3062), .Z(n3063) );
  NANDN U3282 ( .A(n3063), .B(n14296), .Z(n3064) );
  AND U3283 ( .A(n14299), .B(n3064), .Z(n3065) );
  NOR U3284 ( .A(n9888), .B(n3065), .Z(n3066) );
  NAND U3285 ( .A(n9889), .B(n3066), .Z(n3067) );
  ANDN U3286 ( .B(n3067), .A(n9890), .Z(n3068) );
  NAND U3287 ( .A(n9891), .B(n3068), .Z(n3069) );
  AND U3288 ( .A(n9892), .B(n3069), .Z(n3070) );
  NANDN U3289 ( .A(n9893), .B(n3070), .Z(n9894) );
  NANDN U3290 ( .A(n4667), .B(n4830), .Z(n3071) );
  NAND U3291 ( .A(n14358), .B(n3071), .Z(n3072) );
  AND U3292 ( .A(n14361), .B(n3072), .Z(n3073) );
  OR U3293 ( .A(n3073), .B(n14363), .Z(n3074) );
  AND U3294 ( .A(n14365), .B(n3074), .Z(n3075) );
  OR U3295 ( .A(n3075), .B(n14366), .Z(n3076) );
  NAND U3296 ( .A(n14368), .B(n3076), .Z(n3077) );
  NAND U3297 ( .A(n14371), .B(n3077), .Z(n3078) );
  NAND U3298 ( .A(n14373), .B(n3078), .Z(n3079) );
  AND U3299 ( .A(n9949), .B(n3079), .Z(n3080) );
  NAND U3300 ( .A(n3080), .B(n4822), .Z(n3081) );
  NAND U3301 ( .A(n14377), .B(n3081), .Z(n3082) );
  AND U3302 ( .A(n9956), .B(n3082), .Z(n3083) );
  NANDN U3303 ( .A(n4821), .B(n3083), .Z(n4670) );
  NAND U3304 ( .A(n9965), .B(n9966), .Z(n3084) );
  NAND U3305 ( .A(n9967), .B(n3084), .Z(n3085) );
  AND U3306 ( .A(n9968), .B(n3085), .Z(n3086) );
  OR U3307 ( .A(n9969), .B(n3086), .Z(n3087) );
  NAND U3308 ( .A(n9970), .B(n3087), .Z(n3088) );
  NANDN U3309 ( .A(n9971), .B(n3088), .Z(n3089) );
  ANDN U3310 ( .B(n9972), .A(n14396), .Z(n3090) );
  NANDN U3311 ( .A(n3089), .B(n14394), .Z(n3091) );
  AND U3312 ( .A(n3090), .B(n3091), .Z(n3092) );
  NANDN U3313 ( .A(n3092), .B(n14398), .Z(n3093) );
  NANDN U3314 ( .A(n14400), .B(n3093), .Z(n3094) );
  NAND U3315 ( .A(n14402), .B(n3094), .Z(n3095) );
  AND U3316 ( .A(n14407), .B(n9977), .Z(n3096) );
  NANDN U3317 ( .A(n14405), .B(n3095), .Z(n3097) );
  NAND U3318 ( .A(n3096), .B(n3097), .Z(n3098) );
  NANDN U3319 ( .A(n9978), .B(n3098), .Z(n9980) );
  NANDN U3320 ( .A(n14441), .B(n4673), .Z(n3099) );
  NAND U3321 ( .A(n14443), .B(n3099), .Z(n3100) );
  NAND U3322 ( .A(n14445), .B(n3100), .Z(n3101) );
  AND U3323 ( .A(n4798), .B(n10016), .Z(n3102) );
  NAND U3324 ( .A(n3101), .B(n3102), .Z(n3103) );
  NAND U3325 ( .A(n14449), .B(n3103), .Z(n3104) );
  ANDN U3326 ( .B(n4799), .A(n4794), .Z(n3105) );
  NANDN U3327 ( .A(n3104), .B(n4796), .Z(n3106) );
  AND U3328 ( .A(n3105), .B(n3106), .Z(n3107) );
  ANDN U3329 ( .B(n4797), .A(n3107), .Z(n3108) );
  NAND U3330 ( .A(n4793), .B(n3108), .Z(n3109) );
  ANDN U3331 ( .B(n3109), .A(n14459), .Z(n3110) );
  NAND U3332 ( .A(n3110), .B(n4795), .Z(n3111) );
  AND U3333 ( .A(n4792), .B(n3111), .Z(n3112) );
  NAND U3334 ( .A(n3112), .B(n14461), .Z(n4674) );
  AND U3335 ( .A(n14486), .B(n4780), .Z(n4678) );
  ANDN U3336 ( .B(n4689), .A(n4688), .Z(n3113) );
  NAND U3337 ( .A(n10124), .B(n3113), .Z(n3114) );
  ANDN U3338 ( .B(n3114), .A(n10122), .Z(n3115) );
  AND U3339 ( .A(n10125), .B(n4771), .Z(n3116) );
  NANDN U3340 ( .A(n4772), .B(n3115), .Z(n3117) );
  NAND U3341 ( .A(n3116), .B(n3117), .Z(n3118) );
  AND U3342 ( .A(n4773), .B(n3118), .Z(n3119) );
  XNOR U3343 ( .A(y[1973]), .B(x[1973]), .Z(n3120) );
  AND U3344 ( .A(n3119), .B(n3120), .Z(n3121) );
  NANDN U3345 ( .A(n3121), .B(n4770), .Z(n3122) );
  NAND U3346 ( .A(n4769), .B(n3122), .Z(n3123) );
  NAND U3347 ( .A(n10126), .B(n3123), .Z(n3124) );
  NAND U3348 ( .A(n14561), .B(n3124), .Z(n3125) );
  NANDN U3349 ( .A(n14563), .B(n3125), .Z(n3126) );
  AND U3350 ( .A(n14565), .B(n3126), .Z(n3127) );
  NANDN U3351 ( .A(n3127), .B(n14566), .Z(n3128) );
  NAND U3352 ( .A(n14569), .B(n3128), .Z(n3129) );
  NAND U3353 ( .A(n14571), .B(n3129), .Z(n4694) );
  ANDN U3354 ( .B(n10137), .A(n10138), .Z(n3130) );
  NAND U3355 ( .A(n3130), .B(n10139), .Z(n3131) );
  AND U3356 ( .A(n4755), .B(n3131), .Z(n3132) );
  NANDN U3357 ( .A(n4754), .B(n3132), .Z(n3133) );
  NANDN U3358 ( .A(y[1994]), .B(x[1994]), .Z(n3134) );
  AND U3359 ( .A(n4753), .B(n3134), .Z(n3135) );
  NAND U3360 ( .A(n3135), .B(n3133), .Z(n3136) );
  AND U3361 ( .A(n4752), .B(n3136), .Z(n3137) );
  NANDN U3362 ( .A(n4751), .B(n3137), .Z(n3138) );
  AND U3363 ( .A(n4749), .B(n3138), .Z(n3139) );
  ANDN U3364 ( .B(n3139), .A(n10140), .Z(n3140) );
  ANDN U3365 ( .B(n3140), .A(n4750), .Z(n3141) );
  NANDN U3366 ( .A(n3141), .B(n14622), .Z(n3142) );
  NANDN U3367 ( .A(n10141), .B(n3142), .Z(n3143) );
  NAND U3368 ( .A(n14627), .B(n3143), .Z(n3144) );
  NAND U3369 ( .A(n14629), .B(n3144), .Z(n3145) );
  ANDN U3370 ( .B(n3145), .A(n10147), .Z(n3146) );
  NANDN U3371 ( .A(n10146), .B(n3146), .Z(n3147) );
  ANDN U3372 ( .B(n3147), .A(n14632), .Z(n10148) );
  NAND U3373 ( .A(n14659), .B(n4711), .Z(n3148) );
  NAND U3374 ( .A(n14661), .B(n3148), .Z(n3149) );
  ANDN U3375 ( .B(n3149), .A(n4741), .Z(n3150) );
  NAND U3376 ( .A(n4738), .B(n3150), .Z(n3151) );
  AND U3377 ( .A(n10160), .B(n3151), .Z(n3152) );
  NANDN U3378 ( .A(n14665), .B(n3152), .Z(n3153) );
  AND U3379 ( .A(n14670), .B(n4739), .Z(n3154) );
  NAND U3380 ( .A(n3153), .B(n3154), .Z(n3155) );
  NAND U3381 ( .A(n14673), .B(n3155), .Z(n3156) );
  AND U3382 ( .A(n14675), .B(n4736), .Z(n3157) );
  NAND U3383 ( .A(n3156), .B(n3157), .Z(n3158) );
  NANDN U3384 ( .A(n4735), .B(n3158), .Z(n3159) );
  AND U3385 ( .A(n4733), .B(n4737), .Z(n3160) );
  NANDN U3386 ( .A(n3159), .B(n10162), .Z(n3161) );
  AND U3387 ( .A(n3160), .B(n3161), .Z(n4713) );
  ANDN U3388 ( .B(n10167), .A(ebreg), .Z(n3162) );
  NANDN U3389 ( .A(y[2046]), .B(x[2046]), .Z(n3163) );
  AND U3390 ( .A(n10168), .B(n3163), .Z(n3164) );
  NANDN U3391 ( .A(x[2040]), .B(y[2040]), .Z(n3165) );
  NAND U3392 ( .A(n14699), .B(n3165), .Z(n3166) );
  NAND U3393 ( .A(n14700), .B(n3166), .Z(n3167) );
  AND U3394 ( .A(n3167), .B(n14703), .Z(n3168) );
  NANDN U3395 ( .A(n14702), .B(n14701), .Z(n3169) );
  AND U3396 ( .A(n3168), .B(n3169), .Z(n3170) );
  NANDN U3397 ( .A(n3170), .B(n14704), .Z(n3171) );
  AND U3398 ( .A(n14705), .B(n3171), .Z(n3172) );
  NANDN U3399 ( .A(x[2046]), .B(y[2046]), .Z(n3173) );
  NANDN U3400 ( .A(n3172), .B(n3164), .Z(n3174) );
  NAND U3401 ( .A(n3173), .B(n3174), .Z(n3175) );
  NAND U3402 ( .A(n10169), .B(n3175), .Z(n3176) );
  NANDN U3403 ( .A(n3162), .B(g), .Z(n3177) );
  ANDN U3404 ( .B(n3176), .A(n14706), .Z(n3178) );
  NAND U3405 ( .A(n3162), .B(n3178), .Z(n3179) );
  NAND U3406 ( .A(n3177), .B(n3179), .Z(n4) );
  IV U3407 ( .A(ebreg), .Z(e) );
  NANDN U3408 ( .A(x[2042]), .B(y[2042]), .Z(n3181) );
  NANDN U3409 ( .A(x[2041]), .B(y[2041]), .Z(n3180) );
  AND U3410 ( .A(n3181), .B(n3180), .Z(n14702) );
  NANDN U3411 ( .A(x[2043]), .B(y[2043]), .Z(n14703) );
  NANDN U3412 ( .A(x[2044]), .B(y[2044]), .Z(n3183) );
  NANDN U3413 ( .A(x[2045]), .B(y[2045]), .Z(n3182) );
  AND U3414 ( .A(n3183), .B(n3182), .Z(n14705) );
  ANDN U3415 ( .B(y[2047]), .A(x[2047]), .Z(n14706) );
  NANDN U3416 ( .A(y[2044]), .B(x[2044]), .Z(n3185) );
  NANDN U3417 ( .A(y[2043]), .B(x[2043]), .Z(n3184) );
  AND U3418 ( .A(n3185), .B(n3184), .Z(n14704) );
  NANDN U3419 ( .A(x[2037]), .B(y[2037]), .Z(n3187) );
  NANDN U3420 ( .A(x[2038]), .B(y[2038]), .Z(n3186) );
  AND U3421 ( .A(n3187), .B(n3186), .Z(n14696) );
  IV U3422 ( .A(n14696), .Z(n3188) );
  NANDN U3423 ( .A(y[2042]), .B(x[2042]), .Z(n14701) );
  XNOR U3424 ( .A(x[2040]), .B(y[2040]), .Z(n14698) );
  AND U3425 ( .A(n14700), .B(n14698), .Z(n3189) );
  NANDN U3426 ( .A(y[2047]), .B(x[2047]), .Z(n10169) );
  NANDN U3427 ( .A(y[2045]), .B(x[2045]), .Z(n10168) );
  AND U3428 ( .A(n10169), .B(n10168), .Z(n3190) );
  NANDN U3429 ( .A(y[2038]), .B(x[2038]), .Z(n14697) );
  AND U3430 ( .A(n3190), .B(n14697), .Z(n3192) );
  XNOR U3431 ( .A(y[2046]), .B(x[2046]), .Z(n3191) );
  ANDN U3432 ( .B(x[2036]), .A(y[2036]), .Z(n4722) );
  NANDN U3433 ( .A(x[2035]), .B(y[2035]), .Z(n3194) );
  NANDN U3434 ( .A(x[2036]), .B(y[2036]), .Z(n3193) );
  AND U3435 ( .A(n3194), .B(n3193), .Z(n14694) );
  IV U3436 ( .A(n14694), .Z(n4721) );
  NANDN U3437 ( .A(x[2032]), .B(y[2032]), .Z(n14690) );
  NANDN U3438 ( .A(y[2031]), .B(x[2031]), .Z(n4725) );
  NANDN U3439 ( .A(x[2030]), .B(y[2030]), .Z(n4726) );
  NANDN U3440 ( .A(y[2030]), .B(x[2030]), .Z(n4724) );
  ANDN U3441 ( .B(y[2028]), .A(x[2028]), .Z(n4728) );
  NANDN U3442 ( .A(y[2028]), .B(x[2028]), .Z(n10164) );
  NANDN U3443 ( .A(x[2027]), .B(y[2027]), .Z(n4729) );
  ANDN U3444 ( .B(y[2026]), .A(x[2026]), .Z(n4732) );
  IV U3445 ( .A(n4732), .Z(n3195) );
  NANDN U3446 ( .A(x[2024]), .B(y[2024]), .Z(n4737) );
  ANDN U3447 ( .B(x[2023]), .A(y[2023]), .Z(n14676) );
  IV U3448 ( .A(n14676), .Z(n10162) );
  NANDN U3449 ( .A(x[2020]), .B(y[2020]), .Z(n4739) );
  NANDN U3450 ( .A(x[2021]), .B(y[2021]), .Z(n14670) );
  ANDN U3451 ( .B(x[2020]), .A(y[2020]), .Z(n14668) );
  IV U3452 ( .A(n14668), .Z(n10160) );
  NANDN U3453 ( .A(x[2019]), .B(y[2019]), .Z(n4738) );
  NANDN U3454 ( .A(y[2018]), .B(x[2018]), .Z(n4740) );
  ANDN U3455 ( .B(x[2017]), .A(y[2017]), .Z(n10155) );
  ANDN U3456 ( .B(n4740), .A(n10155), .Z(n14661) );
  NANDN U3457 ( .A(x[2017]), .B(y[2017]), .Z(n4742) );
  NANDN U3458 ( .A(x[2016]), .B(y[2016]), .Z(n3196) );
  AND U3459 ( .A(n4742), .B(n3196), .Z(n14659) );
  ANDN U3460 ( .B(x[2013]), .A(y[2013]), .Z(n4744) );
  NANDN U3461 ( .A(y[2012]), .B(x[2012]), .Z(n4745) );
  NANDN U3462 ( .A(y[2011]), .B(x[2011]), .Z(n14646) );
  IV U3463 ( .A(n14646), .Z(n10151) );
  NANDN U3464 ( .A(y[2010]), .B(x[2010]), .Z(n10152) );
  NANDN U3465 ( .A(y[2007]), .B(x[2007]), .Z(n3198) );
  NANDN U3466 ( .A(y[2006]), .B(x[2006]), .Z(n3197) );
  NAND U3467 ( .A(n3198), .B(n3197), .Z(n14637) );
  IV U3468 ( .A(n14637), .Z(n4748) );
  ANDN U3469 ( .B(y[2004]), .A(x[2004]), .Z(n10147) );
  NANDN U3470 ( .A(y[2005]), .B(x[2005]), .Z(n4704) );
  NAND U3471 ( .A(n10147), .B(n4704), .Z(n3201) );
  NANDN U3472 ( .A(x[2006]), .B(y[2006]), .Z(n3200) );
  NANDN U3473 ( .A(x[2005]), .B(y[2005]), .Z(n3199) );
  NAND U3474 ( .A(n3200), .B(n3199), .Z(n10149) );
  ANDN U3475 ( .B(n3201), .A(n10149), .Z(n14634) );
  ANDN U3476 ( .B(x[2003]), .A(y[2003]), .Z(n10144) );
  NANDN U3477 ( .A(x[2002]), .B(y[2002]), .Z(n10142) );
  NANDN U3478 ( .A(y[2002]), .B(x[2002]), .Z(n10145) );
  NANDN U3479 ( .A(x[2001]), .B(y[2001]), .Z(n10143) );
  NANDN U3480 ( .A(x[1998]), .B(y[1998]), .Z(n10175) );
  NANDN U3481 ( .A(x[1999]), .B(y[1999]), .Z(n3202) );
  NANDN U3482 ( .A(x[2000]), .B(y[2000]), .Z(n4699) );
  AND U3483 ( .A(n3202), .B(n4699), .Z(n14622) );
  NANDN U3484 ( .A(x[1997]), .B(y[1997]), .Z(n10174) );
  NANDN U3485 ( .A(y[1993]), .B(x[1993]), .Z(n4758) );
  XNOR U3486 ( .A(y[1994]), .B(x[1994]), .Z(n3203) );
  NAND U3487 ( .A(n4758), .B(n3203), .Z(n14608) );
  NANDN U3488 ( .A(x[1993]), .B(y[1993]), .Z(n14606) );
  IV U3489 ( .A(n14606), .Z(n4754) );
  ANDN U3490 ( .B(x[1991]), .A(y[1991]), .Z(n4756) );
  NANDN U3491 ( .A(x[1990]), .B(y[1990]), .Z(n14596) );
  IV U3492 ( .A(n14596), .Z(n4759) );
  NANDN U3493 ( .A(x[1988]), .B(y[1988]), .Z(n4763) );
  NANDN U3494 ( .A(x[1989]), .B(y[1989]), .Z(n4760) );
  NAND U3495 ( .A(n4763), .B(n4760), .Z(n14592) );
  NANDN U3496 ( .A(y[1988]), .B(x[1988]), .Z(n4761) );
  ANDN U3497 ( .B(x[1987]), .A(y[1987]), .Z(n10136) );
  ANDN U3498 ( .B(n4761), .A(n10136), .Z(n14591) );
  NANDN U3499 ( .A(x[1986]), .B(y[1986]), .Z(n4764) );
  NANDN U3500 ( .A(x[1987]), .B(y[1987]), .Z(n4762) );
  NAND U3501 ( .A(n4764), .B(n4762), .Z(n14588) );
  NANDN U3502 ( .A(y[1985]), .B(x[1985]), .Z(n10135) );
  ANDN U3503 ( .B(x[1986]), .A(y[1986]), .Z(n14586) );
  NANDN U3504 ( .A(x[1985]), .B(y[1985]), .Z(n14584) );
  NANDN U3505 ( .A(y[1978]), .B(x[1978]), .Z(n14566) );
  NANDN U3506 ( .A(x[1977]), .B(y[1977]), .Z(n14565) );
  NANDN U3507 ( .A(y[1976]), .B(x[1976]), .Z(n3205) );
  NANDN U3508 ( .A(y[1977]), .B(x[1977]), .Z(n3204) );
  NAND U3509 ( .A(n3205), .B(n3204), .Z(n14563) );
  NANDN U3510 ( .A(x[1976]), .B(y[1976]), .Z(n3207) );
  NANDN U3511 ( .A(x[1975]), .B(y[1975]), .Z(n3206) );
  AND U3512 ( .A(n3207), .B(n3206), .Z(n14561) );
  NANDN U3513 ( .A(x[1974]), .B(y[1974]), .Z(n4769) );
  NANDN U3514 ( .A(y[1973]), .B(x[1973]), .Z(n4770) );
  NANDN U3515 ( .A(x[1972]), .B(y[1972]), .Z(n4773) );
  NANDN U3516 ( .A(y[1971]), .B(x[1971]), .Z(n10125) );
  ANDN U3517 ( .B(y[1970]), .A(x[1970]), .Z(n10122) );
  NANDN U3518 ( .A(y[1970]), .B(x[1970]), .Z(n10124) );
  NANDN U3519 ( .A(x[1969]), .B(y[1969]), .Z(n10123) );
  ANDN U3520 ( .B(y[1968]), .A(x[1968]), .Z(n14544) );
  NANDN U3521 ( .A(x[1966]), .B(y[1966]), .Z(n3209) );
  NANDN U3522 ( .A(x[1967]), .B(y[1967]), .Z(n3208) );
  AND U3523 ( .A(n3209), .B(n3208), .Z(n14541) );
  ANDN U3524 ( .B(x[1965]), .A(y[1965]), .Z(n10110) );
  XOR U3525 ( .A(x[1966]), .B(y[1966]), .Z(n14538) );
  NANDN U3526 ( .A(y[1962]), .B(x[1962]), .Z(n3211) );
  NANDN U3527 ( .A(y[1961]), .B(x[1961]), .Z(n3210) );
  AND U3528 ( .A(n3211), .B(n3210), .Z(n14527) );
  NANDN U3529 ( .A(x[1960]), .B(y[1960]), .Z(n3213) );
  NANDN U3530 ( .A(x[1961]), .B(y[1961]), .Z(n3212) );
  NAND U3531 ( .A(n3213), .B(n3212), .Z(n14524) );
  NANDN U3532 ( .A(y[1958]), .B(x[1958]), .Z(n3215) );
  NANDN U3533 ( .A(y[1957]), .B(x[1957]), .Z(n3214) );
  NAND U3534 ( .A(n3215), .B(n3214), .Z(n14518) );
  IV U3535 ( .A(n14518), .Z(n4683) );
  NANDN U3536 ( .A(x[1956]), .B(y[1956]), .Z(n3217) );
  NANDN U3537 ( .A(x[1957]), .B(y[1957]), .Z(n3216) );
  AND U3538 ( .A(n3217), .B(n3216), .Z(n14516) );
  IV U3539 ( .A(n14516), .Z(n10091) );
  NANDN U3540 ( .A(y[1954]), .B(x[1954]), .Z(n14510) );
  ANDN U3541 ( .B(x[1953]), .A(y[1953]), .Z(n10080) );
  ANDN U3542 ( .B(n14510), .A(n10080), .Z(n14507) );
  NANDN U3543 ( .A(x[1953]), .B(y[1953]), .Z(n14511) );
  IV U3544 ( .A(n14511), .Z(n10083) );
  ANDN U3545 ( .B(x[1951]), .A(y[1951]), .Z(n10071) );
  ANDN U3546 ( .B(x[1952]), .A(y[1952]), .Z(n10082) );
  NOR U3547 ( .A(n10071), .B(n10082), .Z(n14503) );
  NANDN U3548 ( .A(x[1950]), .B(y[1950]), .Z(n10068) );
  NANDN U3549 ( .A(x[1951]), .B(y[1951]), .Z(n10076) );
  AND U3550 ( .A(n10068), .B(n10076), .Z(n14500) );
  ANDN U3551 ( .B(x[1948]), .A(y[1948]), .Z(n10066) );
  NANDN U3552 ( .A(y[1947]), .B(x[1947]), .Z(n4775) );
  NANDN U3553 ( .A(n10066), .B(n4775), .Z(n14495) );
  NANDN U3554 ( .A(x[1947]), .B(y[1947]), .Z(n10062) );
  NANDN U3555 ( .A(x[1946]), .B(y[1946]), .Z(n4778) );
  NAND U3556 ( .A(n10062), .B(n4778), .Z(n14493) );
  NANDN U3557 ( .A(y[1946]), .B(x[1946]), .Z(n4776) );
  ANDN U3558 ( .B(x[1945]), .A(y[1945]), .Z(n10055) );
  ANDN U3559 ( .B(n4776), .A(n10055), .Z(n14490) );
  NANDN U3560 ( .A(y[1943]), .B(x[1943]), .Z(n4780) );
  NANDN U3561 ( .A(y[1944]), .B(x[1944]), .Z(n14486) );
  ANDN U3562 ( .B(y[1943]), .A(x[1943]), .Z(n14484) );
  NANDN U3563 ( .A(y[1942]), .B(x[1942]), .Z(n4781) );
  NANDN U3564 ( .A(x[1941]), .B(y[1941]), .Z(n4783) );
  ANDN U3565 ( .B(y[1940]), .A(x[1940]), .Z(n14476) );
  NANDN U3566 ( .A(x[1938]), .B(y[1938]), .Z(n4786) );
  NANDN U3567 ( .A(x[1939]), .B(y[1939]), .Z(n10044) );
  AND U3568 ( .A(n4786), .B(n10044), .Z(n14473) );
  NANDN U3569 ( .A(y[1937]), .B(x[1937]), .Z(n4788) );
  NANDN U3570 ( .A(y[1938]), .B(x[1938]), .Z(n4784) );
  NAND U3571 ( .A(n4788), .B(n4784), .Z(n14471) );
  NANDN U3572 ( .A(x[1936]), .B(y[1936]), .Z(n10034) );
  NANDN U3573 ( .A(x[1937]), .B(y[1937]), .Z(n4787) );
  AND U3574 ( .A(n10034), .B(n4787), .Z(n14469) );
  NANDN U3575 ( .A(y[1933]), .B(x[1933]), .Z(n10026) );
  NANDN U3576 ( .A(y[1934]), .B(x[1934]), .Z(n4790) );
  NAND U3577 ( .A(n10026), .B(n4790), .Z(n14462) );
  IV U3578 ( .A(n14462), .Z(n4675) );
  NANDN U3579 ( .A(y[1931]), .B(x[1931]), .Z(n4795) );
  NANDN U3580 ( .A(x[1930]), .B(y[1930]), .Z(n4797) );
  NANDN U3581 ( .A(y[1929]), .B(x[1929]), .Z(n4799) );
  NANDN U3582 ( .A(x[1929]), .B(y[1929]), .Z(n4796) );
  NANDN U3583 ( .A(y[1928]), .B(x[1928]), .Z(n4798) );
  ANDN U3584 ( .B(x[1927]), .A(y[1927]), .Z(n14447) );
  IV U3585 ( .A(n14447), .Z(n10016) );
  ANDN U3586 ( .B(x[1925]), .A(y[1925]), .Z(n4801) );
  ANDN U3587 ( .B(x[1926]), .A(y[1926]), .Z(n10018) );
  NOR U3588 ( .A(n4801), .B(n10018), .Z(n14443) );
  ANDN U3589 ( .B(y[1924]), .A(x[1924]), .Z(n10006) );
  NANDN U3590 ( .A(x[1925]), .B(y[1925]), .Z(n10011) );
  NANDN U3591 ( .A(n10006), .B(n10011), .Z(n14441) );
  NANDN U3592 ( .A(y[1923]), .B(x[1923]), .Z(n4802) );
  ANDN U3593 ( .B(x[1924]), .A(y[1924]), .Z(n4800) );
  ANDN U3594 ( .B(n4802), .A(n4800), .Z(n14439) );
  ANDN U3595 ( .B(y[1922]), .A(x[1922]), .Z(n10001) );
  ANDN U3596 ( .B(y[1923]), .A(x[1923]), .Z(n10007) );
  OR U3597 ( .A(n10001), .B(n10007), .Z(n14436) );
  NANDN U3598 ( .A(y[1921]), .B(x[1921]), .Z(n4804) );
  NANDN U3599 ( .A(y[1922]), .B(x[1922]), .Z(n14435) );
  ANDN U3600 ( .B(y[1921]), .A(x[1921]), .Z(n14433) );
  NANDN U3601 ( .A(y[1920]), .B(x[1920]), .Z(n4803) );
  ANDN U3602 ( .B(y[1919]), .A(x[1919]), .Z(n4806) );
  ANDN U3603 ( .B(y[1918]), .A(x[1918]), .Z(n14425) );
  NANDN U3604 ( .A(y[1915]), .B(x[1915]), .Z(n4811) );
  NANDN U3605 ( .A(y[1916]), .B(x[1916]), .Z(n4808) );
  NAND U3606 ( .A(n4811), .B(n4808), .Z(n14419) );
  NANDN U3607 ( .A(x[1914]), .B(y[1914]), .Z(n4813) );
  NANDN U3608 ( .A(x[1915]), .B(y[1915]), .Z(n4810) );
  AND U3609 ( .A(n4813), .B(n4810), .Z(n14417) );
  NANDN U3610 ( .A(y[1913]), .B(x[1913]), .Z(n4815) );
  NANDN U3611 ( .A(y[1914]), .B(x[1914]), .Z(n4812) );
  NAND U3612 ( .A(n4815), .B(n4812), .Z(n14415) );
  NANDN U3613 ( .A(x[1913]), .B(y[1913]), .Z(n4814) );
  ANDN U3614 ( .B(y[1912]), .A(x[1912]), .Z(n9978) );
  ANDN U3615 ( .B(n4814), .A(n9978), .Z(n14413) );
  NANDN U3616 ( .A(y[1911]), .B(x[1911]), .Z(n9977) );
  NANDN U3617 ( .A(y[1912]), .B(x[1912]), .Z(n4816) );
  NAND U3618 ( .A(n9977), .B(n4816), .Z(n14411) );
  ANDN U3619 ( .B(x[1909]), .A(y[1909]), .Z(n4820) );
  NANDN U3620 ( .A(x[1908]), .B(y[1908]), .Z(n9976) );
  ANDN U3621 ( .B(x[1907]), .A(y[1907]), .Z(n9973) );
  NANDN U3622 ( .A(x[1907]), .B(y[1907]), .Z(n9975) );
  NANDN U3623 ( .A(y[1905]), .B(x[1905]), .Z(n14394) );
  NANDN U3624 ( .A(y[1906]), .B(x[1906]), .Z(n9974) );
  NANDN U3625 ( .A(x[1904]), .B(y[1904]), .Z(n9970) );
  NANDN U3626 ( .A(x[1905]), .B(y[1905]), .Z(n9972) );
  AND U3627 ( .A(n9970), .B(n9972), .Z(n14393) );
  ANDN U3628 ( .B(x[1903]), .A(y[1903]), .Z(n9969) );
  ANDN U3629 ( .B(x[1904]), .A(y[1904]), .Z(n9971) );
  OR U3630 ( .A(n9969), .B(n9971), .Z(n14391) );
  XOR U3631 ( .A(x[1900]), .B(y[1900]), .Z(n14378) );
  IV U3632 ( .A(n14378), .Z(n9956) );
  NANDN U3633 ( .A(x[1898]), .B(y[1898]), .Z(n4823) );
  NANDN U3634 ( .A(x[1899]), .B(y[1899]), .Z(n14380) );
  IV U3635 ( .A(n14380), .Z(n9955) );
  ANDN U3636 ( .B(n4823), .A(n9955), .Z(n14377) );
  ANDN U3637 ( .B(x[1897]), .A(y[1897]), .Z(n14375) );
  IV U3638 ( .A(n14375), .Z(n9949) );
  NANDN U3639 ( .A(x[1896]), .B(y[1896]), .Z(n9945) );
  NANDN U3640 ( .A(x[1897]), .B(y[1897]), .Z(n4824) );
  AND U3641 ( .A(n9945), .B(n4824), .Z(n14373) );
  NANDN U3642 ( .A(y[1891]), .B(x[1891]), .Z(n9930) );
  NANDN U3643 ( .A(y[1892]), .B(x[1892]), .Z(n4828) );
  NAND U3644 ( .A(n9930), .B(n4828), .Z(n14363) );
  ANDN U3645 ( .B(y[1889]), .A(x[1889]), .Z(n14356) );
  NANDN U3646 ( .A(y[1887]), .B(x[1887]), .Z(n4832) );
  ANDN U3647 ( .B(y[1886]), .A(x[1886]), .Z(n4833) );
  NANDN U3648 ( .A(y[1885]), .B(x[1885]), .Z(n9926) );
  ANDN U3649 ( .B(y[1884]), .A(x[1884]), .Z(n14342) );
  NANDN U3650 ( .A(x[1882]), .B(y[1882]), .Z(n9924) );
  NANDN U3651 ( .A(x[1883]), .B(y[1883]), .Z(n4835) );
  NAND U3652 ( .A(n9924), .B(n4835), .Z(n14340) );
  NANDN U3653 ( .A(x[1880]), .B(y[1880]), .Z(n4839) );
  NANDN U3654 ( .A(x[1881]), .B(y[1881]), .Z(n9925) );
  NAND U3655 ( .A(n4839), .B(n9925), .Z(n14334) );
  ANDN U3656 ( .B(x[1878]), .A(y[1878]), .Z(n14329) );
  NANDN U3657 ( .A(x[1876]), .B(y[1876]), .Z(n4844) );
  ANDN U3658 ( .B(x[1875]), .A(y[1875]), .Z(n14321) );
  IV U3659 ( .A(n14321), .Z(n9912) );
  NANDN U3660 ( .A(x[1874]), .B(y[1874]), .Z(n14319) );
  NANDN U3661 ( .A(x[1875]), .B(y[1875]), .Z(n4843) );
  NANDN U3662 ( .A(y[1873]), .B(x[1873]), .Z(n9903) );
  NANDN U3663 ( .A(y[1874]), .B(x[1874]), .Z(n9910) );
  NAND U3664 ( .A(n9903), .B(n9910), .Z(n14317) );
  ANDN U3665 ( .B(y[1873]), .A(x[1873]), .Z(n9908) );
  NANDN U3666 ( .A(x[1872]), .B(y[1872]), .Z(n4845) );
  NANDN U3667 ( .A(n9908), .B(n4845), .Z(n14315) );
  NANDN U3668 ( .A(y[1871]), .B(x[1871]), .Z(n9896) );
  NANDN U3669 ( .A(y[1872]), .B(x[1872]), .Z(n9905) );
  AND U3670 ( .A(n9896), .B(n9905), .Z(n14313) );
  NANDN U3671 ( .A(x[1870]), .B(y[1870]), .Z(n4848) );
  NANDN U3672 ( .A(x[1871]), .B(y[1871]), .Z(n4846) );
  NAND U3673 ( .A(n4848), .B(n4846), .Z(n14311) );
  ANDN U3674 ( .B(y[1867]), .A(x[1867]), .Z(n14302) );
  IV U3675 ( .A(n14302), .Z(n9891) );
  NANDN U3676 ( .A(y[1865]), .B(x[1865]), .Z(n4852) );
  ANDN U3677 ( .B(y[1864]), .A(x[1864]), .Z(n9886) );
  NANDN U3678 ( .A(y[1863]), .B(x[1863]), .Z(n9885) );
  ANDN U3679 ( .B(y[1862]), .A(x[1862]), .Z(n14290) );
  IV U3680 ( .A(n14290), .Z(n9883) );
  NANDN U3681 ( .A(y[1861]), .B(x[1861]), .Z(n14288) );
  IV U3682 ( .A(n14288), .Z(n9880) );
  NANDN U3683 ( .A(y[1862]), .B(x[1862]), .Z(n9884) );
  ANDN U3684 ( .B(y[1860]), .A(x[1860]), .Z(n4854) );
  ANDN U3685 ( .B(y[1861]), .A(x[1861]), .Z(n9882) );
  NOR U3686 ( .A(n4854), .B(n9882), .Z(n14287) );
  ANDN U3687 ( .B(x[1859]), .A(y[1859]), .Z(n9878) );
  NANDN U3688 ( .A(y[1860]), .B(x[1860]), .Z(n9881) );
  NANDN U3689 ( .A(n9878), .B(n9881), .Z(n14285) );
  NANDN U3690 ( .A(x[1858]), .B(y[1858]), .Z(n4855) );
  ANDN U3691 ( .B(y[1859]), .A(x[1859]), .Z(n4853) );
  ANDN U3692 ( .B(n4855), .A(n4853), .Z(n14283) );
  ANDN U3693 ( .B(x[1853]), .A(y[1853]), .Z(n14269) );
  IV U3694 ( .A(n14269), .Z(n9862) );
  NANDN U3695 ( .A(x[1852]), .B(y[1852]), .Z(n9858) );
  NANDN U3696 ( .A(x[1853]), .B(y[1853]), .Z(n4858) );
  AND U3697 ( .A(n9858), .B(n4858), .Z(n14267) );
  NANDN U3698 ( .A(y[1849]), .B(x[1849]), .Z(n4864) );
  NANDN U3699 ( .A(y[1850]), .B(x[1850]), .Z(n4859) );
  NAND U3700 ( .A(n4864), .B(n4859), .Z(n14260) );
  ANDN U3701 ( .B(y[1848]), .A(x[1848]), .Z(n9848) );
  NANDN U3702 ( .A(x[1849]), .B(y[1849]), .Z(n4862) );
  NANDN U3703 ( .A(n9848), .B(n4862), .Z(n14259) );
  NANDN U3704 ( .A(y[1847]), .B(x[1847]), .Z(n4865) );
  NANDN U3705 ( .A(y[1848]), .B(x[1848]), .Z(n4863) );
  AND U3706 ( .A(n4865), .B(n4863), .Z(n14257) );
  ANDN U3707 ( .B(y[1845]), .A(x[1845]), .Z(n14250) );
  IV U3708 ( .A(n14250), .Z(n9844) );
  NANDN U3709 ( .A(y[1843]), .B(x[1843]), .Z(n4869) );
  ANDN U3710 ( .B(y[1842]), .A(x[1842]), .Z(n4872) );
  NANDN U3711 ( .A(y[1842]), .B(x[1842]), .Z(n4870) );
  ANDN U3712 ( .B(y[1840]), .A(x[1840]), .Z(n14239) );
  NANDN U3713 ( .A(y[1840]), .B(x[1840]), .Z(n4874) );
  NANDN U3714 ( .A(x[1838]), .B(y[1838]), .Z(n3218) );
  NANDN U3715 ( .A(x[1839]), .B(y[1839]), .Z(n9840) );
  NAND U3716 ( .A(n3218), .B(n9840), .Z(n14234) );
  XNOR U3717 ( .A(x[1838]), .B(y[1838]), .Z(n4876) );
  NANDN U3718 ( .A(y[1837]), .B(x[1837]), .Z(n9839) );
  AND U3719 ( .A(n4876), .B(n9839), .Z(n14233) );
  NANDN U3720 ( .A(x[1836]), .B(y[1836]), .Z(n3219) );
  NANDN U3721 ( .A(x[1837]), .B(y[1837]), .Z(n4875) );
  NAND U3722 ( .A(n3219), .B(n4875), .Z(n14230) );
  XNOR U3723 ( .A(x[1836]), .B(y[1836]), .Z(n4878) );
  NANDN U3724 ( .A(y[1835]), .B(x[1835]), .Z(n4879) );
  AND U3725 ( .A(n4878), .B(n4879), .Z(n14229) );
  NANDN U3726 ( .A(x[1834]), .B(y[1834]), .Z(n3220) );
  NANDN U3727 ( .A(x[1835]), .B(y[1835]), .Z(n4877) );
  NAND U3728 ( .A(n3220), .B(n4877), .Z(n14226) );
  XNOR U3729 ( .A(x[1834]), .B(y[1834]), .Z(n14225) );
  NANDN U3730 ( .A(x[1833]), .B(y[1833]), .Z(n14222) );
  NANDN U3731 ( .A(x[1832]), .B(y[1832]), .Z(n14218) );
  ANDN U3732 ( .B(x[1831]), .A(y[1831]), .Z(n14216) );
  NANDN U3733 ( .A(x[1830]), .B(y[1830]), .Z(n4883) );
  ANDN U3734 ( .B(y[1831]), .A(x[1831]), .Z(n9836) );
  ANDN U3735 ( .B(n4883), .A(n9836), .Z(n14214) );
  NANDN U3736 ( .A(y[1827]), .B(x[1827]), .Z(n9833) );
  NANDN U3737 ( .A(y[1828]), .B(x[1828]), .Z(n4885) );
  NAND U3738 ( .A(n9833), .B(n4885), .Z(n14209) );
  NANDN U3739 ( .A(x[1826]), .B(y[1826]), .Z(n4889) );
  NANDN U3740 ( .A(x[1827]), .B(y[1827]), .Z(n4887) );
  NAND U3741 ( .A(n4889), .B(n4887), .Z(n14207) );
  NANDN U3742 ( .A(y[1825]), .B(x[1825]), .Z(n9829) );
  NANDN U3743 ( .A(y[1826]), .B(x[1826]), .Z(n9834) );
  AND U3744 ( .A(n9829), .B(n9834), .Z(n14204) );
  ANDN U3745 ( .B(y[1823]), .A(x[1823]), .Z(n14199) );
  IV U3746 ( .A(n14199), .Z(n9828) );
  NANDN U3747 ( .A(y[1821]), .B(x[1821]), .Z(n4893) );
  NANDN U3748 ( .A(x[1821]), .B(y[1821]), .Z(n4891) );
  NANDN U3749 ( .A(x[1820]), .B(y[1820]), .Z(n9824) );
  ANDN U3750 ( .B(x[1820]), .A(y[1820]), .Z(n4892) );
  NANDN U3751 ( .A(y[1819]), .B(x[1819]), .Z(n9822) );
  ANDN U3752 ( .B(y[1818]), .A(x[1818]), .Z(n14186) );
  IV U3753 ( .A(n14186), .Z(n9820) );
  NANDN U3754 ( .A(y[1817]), .B(x[1817]), .Z(n14184) );
  IV U3755 ( .A(n14184), .Z(n9818) );
  NANDN U3756 ( .A(y[1818]), .B(x[1818]), .Z(n9821) );
  NANDN U3757 ( .A(x[1816]), .B(y[1816]), .Z(n4894) );
  ANDN U3758 ( .B(y[1817]), .A(x[1817]), .Z(n9819) );
  ANDN U3759 ( .B(n4894), .A(n9819), .Z(n14183) );
  NANDN U3760 ( .A(y[1815]), .B(x[1815]), .Z(n9815) );
  NANDN U3761 ( .A(y[1816]), .B(x[1816]), .Z(n9817) );
  NAND U3762 ( .A(n9815), .B(n9817), .Z(n14181) );
  NANDN U3763 ( .A(x[1814]), .B(y[1814]), .Z(n4897) );
  NANDN U3764 ( .A(x[1815]), .B(y[1815]), .Z(n4895) );
  AND U3765 ( .A(n4897), .B(n4895), .Z(n14179) );
  ANDN U3766 ( .B(x[1812]), .A(y[1812]), .Z(n14172) );
  IV U3767 ( .A(n14172), .Z(n9811) );
  NANDN U3768 ( .A(x[1810]), .B(y[1810]), .Z(n4901) );
  ANDN U3769 ( .B(x[1809]), .A(y[1809]), .Z(n14165) );
  NANDN U3770 ( .A(x[1809]), .B(y[1809]), .Z(n4900) );
  NANDN U3771 ( .A(x[1807]), .B(y[1807]), .Z(n3222) );
  NANDN U3772 ( .A(x[1806]), .B(y[1806]), .Z(n3221) );
  AND U3773 ( .A(n3222), .B(n3221), .Z(n14159) );
  NANDN U3774 ( .A(y[1805]), .B(x[1805]), .Z(n3224) );
  NANDN U3775 ( .A(y[1806]), .B(x[1806]), .Z(n3223) );
  NAND U3776 ( .A(n3224), .B(n3223), .Z(n14156) );
  NANDN U3777 ( .A(x[1805]), .B(y[1805]), .Z(n3226) );
  NANDN U3778 ( .A(x[1804]), .B(y[1804]), .Z(n3225) );
  AND U3779 ( .A(n3226), .B(n3225), .Z(n14155) );
  ANDN U3780 ( .B(x[1804]), .A(y[1804]), .Z(n9791) );
  NANDN U3781 ( .A(y[1803]), .B(x[1803]), .Z(n3227) );
  NANDN U3782 ( .A(n9791), .B(n3227), .Z(n14152) );
  NANDN U3783 ( .A(x[1803]), .B(y[1803]), .Z(n3228) );
  ANDN U3784 ( .B(y[1802]), .A(x[1802]), .Z(n9788) );
  ANDN U3785 ( .B(n3228), .A(n9788), .Z(n14151) );
  NANDN U3786 ( .A(y[1801]), .B(x[1801]), .Z(n9783) );
  NANDN U3787 ( .A(y[1802]), .B(x[1802]), .Z(n9790) );
  NAND U3788 ( .A(n9783), .B(n9790), .Z(n14149) );
  ANDN U3789 ( .B(x[1800]), .A(y[1800]), .Z(n14144) );
  NANDN U3790 ( .A(x[1800]), .B(y[1800]), .Z(n3230) );
  NANDN U3791 ( .A(x[1799]), .B(y[1799]), .Z(n3229) );
  AND U3792 ( .A(n3230), .B(n3229), .Z(n14143) );
  NANDN U3793 ( .A(y[1799]), .B(x[1799]), .Z(n14141) );
  NANDN U3794 ( .A(y[1798]), .B(x[1798]), .Z(n10176) );
  NAND U3795 ( .A(n14141), .B(n10176), .Z(n9781) );
  NANDN U3796 ( .A(x[1798]), .B(y[1798]), .Z(n14138) );
  IV U3797 ( .A(n14138), .Z(n4903) );
  NANDN U3798 ( .A(y[1797]), .B(x[1797]), .Z(n10177) );
  NANDN U3799 ( .A(x[1796]), .B(y[1796]), .Z(n9773) );
  NANDN U3800 ( .A(x[1797]), .B(y[1797]), .Z(n4902) );
  NAND U3801 ( .A(n9773), .B(n4902), .Z(n14135) );
  NANDN U3802 ( .A(y[1796]), .B(x[1796]), .Z(n4904) );
  ANDN U3803 ( .B(x[1795]), .A(y[1795]), .Z(n9769) );
  ANDN U3804 ( .B(n4904), .A(n9769), .Z(n14133) );
  ANDN U3805 ( .B(y[1795]), .A(x[1795]), .Z(n9775) );
  NANDN U3806 ( .A(x[1794]), .B(y[1794]), .Z(n9767) );
  NANDN U3807 ( .A(n9775), .B(n9767), .Z(n14131) );
  XNOR U3808 ( .A(x[1794]), .B(y[1794]), .Z(n3231) );
  ANDN U3809 ( .B(x[1793]), .A(y[1793]), .Z(n9765) );
  ANDN U3810 ( .B(n3231), .A(n9765), .Z(n14129) );
  NANDN U3811 ( .A(x[1792]), .B(y[1792]), .Z(n3233) );
  NANDN U3812 ( .A(x[1793]), .B(y[1793]), .Z(n3232) );
  AND U3813 ( .A(n3233), .B(n3232), .Z(n4908) );
  NANDN U3814 ( .A(y[1791]), .B(x[1791]), .Z(n3234) );
  ANDN U3815 ( .B(x[1792]), .A(y[1792]), .Z(n4906) );
  ANDN U3816 ( .B(n3234), .A(n4906), .Z(n3238) );
  NANDN U3817 ( .A(x[1790]), .B(y[1790]), .Z(n4909) );
  NANDN U3818 ( .A(x[1791]), .B(y[1791]), .Z(n4905) );
  NAND U3819 ( .A(n4909), .B(n4905), .Z(n3235) );
  NAND U3820 ( .A(n3238), .B(n3235), .Z(n3236) );
  NAND U3821 ( .A(n4908), .B(n3236), .Z(n14127) );
  NANDN U3822 ( .A(y[1790]), .B(x[1790]), .Z(n3237) );
  NAND U3823 ( .A(n3238), .B(n3237), .Z(n14124) );
  NANDN U3824 ( .A(y[1789]), .B(x[1789]), .Z(n4911) );
  NANDN U3825 ( .A(x[1789]), .B(y[1789]), .Z(n14123) );
  NANDN U3826 ( .A(y[1788]), .B(x[1788]), .Z(n4910) );
  ANDN U3827 ( .B(y[1786]), .A(x[1786]), .Z(n14115) );
  NANDN U3828 ( .A(y[1785]), .B(x[1785]), .Z(n4915) );
  ANDN U3829 ( .B(x[1786]), .A(y[1786]), .Z(n4914) );
  ANDN U3830 ( .B(n4915), .A(n4914), .Z(n14113) );
  ANDN U3831 ( .B(y[1784]), .A(x[1784]), .Z(n9755) );
  ANDN U3832 ( .B(y[1785]), .A(x[1785]), .Z(n9757) );
  OR U3833 ( .A(n9755), .B(n9757), .Z(n14111) );
  NANDN U3834 ( .A(y[1783]), .B(x[1783]), .Z(n9754) );
  NANDN U3835 ( .A(y[1784]), .B(x[1784]), .Z(n4916) );
  AND U3836 ( .A(n9754), .B(n4916), .Z(n14109) );
  ANDN U3837 ( .B(y[1782]), .A(x[1782]), .Z(n9751) );
  ANDN U3838 ( .B(y[1783]), .A(x[1783]), .Z(n9756) );
  OR U3839 ( .A(n9751), .B(n9756), .Z(n14107) );
  NANDN U3840 ( .A(y[1781]), .B(x[1781]), .Z(n9749) );
  NANDN U3841 ( .A(y[1782]), .B(x[1782]), .Z(n9753) );
  AND U3842 ( .A(n9749), .B(n9753), .Z(n14105) );
  ANDN U3843 ( .B(y[1780]), .A(x[1780]), .Z(n9748) );
  ANDN U3844 ( .B(y[1781]), .A(x[1781]), .Z(n9752) );
  OR U3845 ( .A(n9748), .B(n9752), .Z(n14103) );
  NANDN U3846 ( .A(y[1777]), .B(x[1777]), .Z(n4920) );
  NANDN U3847 ( .A(x[1776]), .B(y[1776]), .Z(n4921) );
  NANDN U3848 ( .A(y[1771]), .B(x[1771]), .Z(n9727) );
  NANDN U3849 ( .A(y[1772]), .B(x[1772]), .Z(n9734) );
  NAND U3850 ( .A(n9727), .B(n9734), .Z(n14081) );
  ANDN U3851 ( .B(y[1770]), .A(x[1770]), .Z(n9724) );
  ANDN U3852 ( .B(y[1771]), .A(x[1771]), .Z(n9733) );
  OR U3853 ( .A(n9724), .B(n9733), .Z(n14079) );
  NANDN U3854 ( .A(y[1769]), .B(x[1769]), .Z(n4925) );
  NANDN U3855 ( .A(y[1770]), .B(x[1770]), .Z(n9728) );
  AND U3856 ( .A(n4925), .B(n9728), .Z(n14077) );
  ANDN U3857 ( .B(y[1769]), .A(x[1769]), .Z(n14075) );
  NANDN U3858 ( .A(y[1767]), .B(x[1767]), .Z(n4927) );
  ANDN U3859 ( .B(x[1768]), .A(y[1768]), .Z(n10178) );
  ANDN U3860 ( .B(n4927), .A(n10178), .Z(n14069) );
  NANDN U3861 ( .A(x[1766]), .B(y[1766]), .Z(n3240) );
  NANDN U3862 ( .A(x[1765]), .B(y[1765]), .Z(n3239) );
  AND U3863 ( .A(n3240), .B(n3239), .Z(n9715) );
  NANDN U3864 ( .A(x[1764]), .B(y[1764]), .Z(n3241) );
  AND U3865 ( .A(n9715), .B(n3241), .Z(n14067) );
  NANDN U3866 ( .A(y[1764]), .B(x[1764]), .Z(n9713) );
  NANDN U3867 ( .A(y[1763]), .B(x[1763]), .Z(n4928) );
  AND U3868 ( .A(n9713), .B(n4928), .Z(n14064) );
  NANDN U3869 ( .A(x[1760]), .B(y[1760]), .Z(n4935) );
  NANDN U3870 ( .A(x[1761]), .B(y[1761]), .Z(n4930) );
  NAND U3871 ( .A(n4935), .B(n4930), .Z(n14059) );
  NANDN U3872 ( .A(y[1759]), .B(x[1759]), .Z(n9697) );
  NANDN U3873 ( .A(y[1760]), .B(x[1760]), .Z(n4933) );
  AND U3874 ( .A(n9697), .B(n4933), .Z(n14057) );
  ANDN U3875 ( .B(y[1758]), .A(x[1758]), .Z(n9694) );
  NANDN U3876 ( .A(x[1759]), .B(y[1759]), .Z(n4934) );
  NANDN U3877 ( .A(n9694), .B(n4934), .Z(n14055) );
  NANDN U3878 ( .A(y[1757]), .B(x[1757]), .Z(n9690) );
  ANDN U3879 ( .B(x[1758]), .A(y[1758]), .Z(n9699) );
  ANDN U3880 ( .B(n9690), .A(n9699), .Z(n14053) );
  ANDN U3881 ( .B(y[1757]), .A(x[1757]), .Z(n14051) );
  NANDN U3882 ( .A(y[1755]), .B(x[1755]), .Z(n4939) );
  ANDN U3883 ( .B(y[1754]), .A(x[1754]), .Z(n4941) );
  NANDN U3884 ( .A(y[1753]), .B(x[1753]), .Z(n9688) );
  NANDN U3885 ( .A(y[1751]), .B(x[1751]), .Z(n14036) );
  NANDN U3886 ( .A(x[1750]), .B(y[1750]), .Z(n3242) );
  ANDN U3887 ( .B(y[1751]), .A(x[1751]), .Z(n9686) );
  ANDN U3888 ( .B(n3242), .A(n9686), .Z(n14035) );
  XNOR U3889 ( .A(x[1750]), .B(y[1750]), .Z(n4942) );
  NANDN U3890 ( .A(y[1749]), .B(x[1749]), .Z(n4944) );
  NAND U3891 ( .A(n4942), .B(n4944), .Z(n14033) );
  NANDN U3892 ( .A(x[1748]), .B(y[1748]), .Z(n4947) );
  NANDN U3893 ( .A(x[1749]), .B(y[1749]), .Z(n4943) );
  AND U3894 ( .A(n4947), .B(n4943), .Z(n14031) );
  ANDN U3895 ( .B(x[1745]), .A(y[1745]), .Z(n9681) );
  NANDN U3896 ( .A(x[1745]), .B(y[1745]), .Z(n14023) );
  NANDN U3897 ( .A(y[1744]), .B(x[1744]), .Z(n9682) );
  ANDN U3898 ( .B(y[1742]), .A(x[1742]), .Z(n14014) );
  NANDN U3899 ( .A(y[1741]), .B(x[1741]), .Z(n9676) );
  NANDN U3900 ( .A(y[1742]), .B(x[1742]), .Z(n9678) );
  AND U3901 ( .A(n9676), .B(n9678), .Z(n14013) );
  ANDN U3902 ( .B(y[1741]), .A(x[1741]), .Z(n9677) );
  NANDN U3903 ( .A(x[1740]), .B(y[1740]), .Z(n4950) );
  NANDN U3904 ( .A(n9677), .B(n4950), .Z(n14011) );
  NANDN U3905 ( .A(y[1739]), .B(x[1739]), .Z(n4951) );
  NANDN U3906 ( .A(y[1740]), .B(x[1740]), .Z(n9675) );
  AND U3907 ( .A(n4951), .B(n9675), .Z(n14009) );
  NANDN U3908 ( .A(x[1738]), .B(y[1738]), .Z(n4954) );
  NANDN U3909 ( .A(x[1739]), .B(y[1739]), .Z(n4949) );
  NAND U3910 ( .A(n4954), .B(n4949), .Z(n14007) );
  NANDN U3911 ( .A(y[1737]), .B(x[1737]), .Z(n9673) );
  NANDN U3912 ( .A(y[1738]), .B(x[1738]), .Z(n4952) );
  NAND U3913 ( .A(n9673), .B(n4952), .Z(n14005) );
  NANDN U3914 ( .A(x[1737]), .B(y[1737]), .Z(n4953) );
  ANDN U3915 ( .B(y[1736]), .A(x[1736]), .Z(n9672) );
  ANDN U3916 ( .B(n4953), .A(n9672), .Z(n14002) );
  NANDN U3917 ( .A(y[1734]), .B(x[1734]), .Z(n13996) );
  NANDN U3918 ( .A(x[1732]), .B(y[1732]), .Z(n4959) );
  NANDN U3919 ( .A(y[1731]), .B(x[1731]), .Z(n4962) );
  ANDN U3920 ( .B(y[1730]), .A(x[1730]), .Z(n13987) );
  NANDN U3921 ( .A(y[1727]), .B(x[1727]), .Z(n4965) );
  NANDN U3922 ( .A(y[1728]), .B(x[1728]), .Z(n9667) );
  NAND U3923 ( .A(n4965), .B(n9667), .Z(n13981) );
  NANDN U3924 ( .A(x[1726]), .B(y[1726]), .Z(n4968) );
  NANDN U3925 ( .A(x[1727]), .B(y[1727]), .Z(n4963) );
  NAND U3926 ( .A(n4968), .B(n4963), .Z(n13979) );
  NANDN U3927 ( .A(y[1726]), .B(x[1726]), .Z(n4966) );
  ANDN U3928 ( .B(x[1725]), .A(y[1725]), .Z(n9666) );
  ANDN U3929 ( .B(n4966), .A(n9666), .Z(n13977) );
  NANDN U3930 ( .A(x[1724]), .B(y[1724]), .Z(n4970) );
  NANDN U3931 ( .A(x[1725]), .B(y[1725]), .Z(n4967) );
  NAND U3932 ( .A(n4970), .B(n4967), .Z(n13975) );
  NANDN U3933 ( .A(y[1723]), .B(x[1723]), .Z(n9664) );
  ANDN U3934 ( .B(x[1724]), .A(y[1724]), .Z(n13973) );
  NANDN U3935 ( .A(x[1723]), .B(y[1723]), .Z(n13971) );
  NANDN U3936 ( .A(x[1722]), .B(y[1722]), .Z(n9662) );
  ANDN U3937 ( .B(x[1721]), .A(y[1721]), .Z(n13964) );
  IV U3938 ( .A(n13964), .Z(n9660) );
  NANDN U3939 ( .A(x[1718]), .B(y[1718]), .Z(n4971) );
  ANDN U3940 ( .B(y[1719]), .A(x[1719]), .Z(n9658) );
  ANDN U3941 ( .B(n4971), .A(n9658), .Z(n13959) );
  NANDN U3942 ( .A(y[1717]), .B(x[1717]), .Z(n4973) );
  NANDN U3943 ( .A(y[1718]), .B(x[1718]), .Z(n9656) );
  NAND U3944 ( .A(n4973), .B(n9656), .Z(n13957) );
  NANDN U3945 ( .A(x[1716]), .B(y[1716]), .Z(n4975) );
  NANDN U3946 ( .A(x[1717]), .B(y[1717]), .Z(n4972) );
  AND U3947 ( .A(n4975), .B(n4972), .Z(n13955) );
  NANDN U3948 ( .A(y[1715]), .B(x[1715]), .Z(n4978) );
  NANDN U3949 ( .A(y[1716]), .B(x[1716]), .Z(n4974) );
  NAND U3950 ( .A(n4978), .B(n4974), .Z(n13953) );
  NANDN U3951 ( .A(x[1715]), .B(y[1715]), .Z(n4976) );
  ANDN U3952 ( .B(y[1714]), .A(x[1714]), .Z(n9655) );
  ANDN U3953 ( .B(n4976), .A(n9655), .Z(n13951) );
  NANDN U3954 ( .A(y[1713]), .B(x[1713]), .Z(n9653) );
  NANDN U3955 ( .A(y[1714]), .B(x[1714]), .Z(n4977) );
  NAND U3956 ( .A(n9653), .B(n4977), .Z(n13949) );
  NANDN U3957 ( .A(y[1712]), .B(x[1712]), .Z(n13944) );
  IV U3958 ( .A(n13944), .Z(n9652) );
  NANDN U3959 ( .A(y[1711]), .B(x[1711]), .Z(n4982) );
  NANDN U3960 ( .A(x[1711]), .B(y[1711]), .Z(n4980) );
  NANDN U3961 ( .A(x[1710]), .B(y[1710]), .Z(n9648) );
  ANDN U3962 ( .B(x[1710]), .A(y[1710]), .Z(n4981) );
  NANDN U3963 ( .A(y[1709]), .B(x[1709]), .Z(n9647) );
  NANDN U3964 ( .A(y[1707]), .B(x[1707]), .Z(n13932) );
  NANDN U3965 ( .A(x[1706]), .B(y[1706]), .Z(n4984) );
  ANDN U3966 ( .B(y[1707]), .A(x[1707]), .Z(n9645) );
  ANDN U3967 ( .B(n4984), .A(n9645), .Z(n13931) );
  NANDN U3968 ( .A(y[1705]), .B(x[1705]), .Z(n4985) );
  NANDN U3969 ( .A(y[1706]), .B(x[1706]), .Z(n9644) );
  NAND U3970 ( .A(n4985), .B(n9644), .Z(n13929) );
  NANDN U3971 ( .A(x[1704]), .B(y[1704]), .Z(n4988) );
  NANDN U3972 ( .A(x[1705]), .B(y[1705]), .Z(n4983) );
  AND U3973 ( .A(n4988), .B(n4983), .Z(n13927) );
  ANDN U3974 ( .B(x[1702]), .A(y[1702]), .Z(n13920) );
  IV U3975 ( .A(n13920), .Z(n9643) );
  NANDN U3976 ( .A(x[1701]), .B(y[1701]), .Z(n13919) );
  IV U3977 ( .A(n13919), .Z(n4989) );
  NANDN U3978 ( .A(y[1697]), .B(x[1697]), .Z(n3244) );
  NANDN U3979 ( .A(y[1696]), .B(x[1696]), .Z(n3243) );
  NAND U3980 ( .A(n3244), .B(n3243), .Z(n10182) );
  NANDN U3981 ( .A(x[1695]), .B(y[1695]), .Z(n3245) );
  ANDN U3982 ( .B(y[1696]), .A(x[1696]), .Z(n10181) );
  ANDN U3983 ( .B(n3245), .A(n10181), .Z(n4628) );
  ANDN U3984 ( .B(x[1694]), .A(y[1694]), .Z(n10184) );
  NANDN U3985 ( .A(y[1695]), .B(x[1695]), .Z(n10180) );
  NANDN U3986 ( .A(y[1691]), .B(x[1691]), .Z(n9631) );
  ANDN U3987 ( .B(x[1692]), .A(y[1692]), .Z(n9632) );
  ANDN U3988 ( .B(n9631), .A(n9632), .Z(n13901) );
  NANDN U3989 ( .A(x[1691]), .B(y[1691]), .Z(n13898) );
  ANDN U3990 ( .B(x[1690]), .A(y[1690]), .Z(n13896) );
  NANDN U3991 ( .A(x[1689]), .B(y[1689]), .Z(n3247) );
  NANDN U3992 ( .A(x[1690]), .B(y[1690]), .Z(n3246) );
  NAND U3993 ( .A(n3247), .B(n3246), .Z(n13895) );
  NANDN U3994 ( .A(y[1689]), .B(x[1689]), .Z(n3249) );
  NANDN U3995 ( .A(y[1688]), .B(x[1688]), .Z(n3248) );
  AND U3996 ( .A(n3249), .B(n3248), .Z(n13893) );
  NANDN U3997 ( .A(x[1687]), .B(y[1687]), .Z(n3251) );
  NANDN U3998 ( .A(x[1688]), .B(y[1688]), .Z(n3250) );
  NAND U3999 ( .A(n3251), .B(n3250), .Z(n13891) );
  NANDN U4000 ( .A(y[1687]), .B(x[1687]), .Z(n4993) );
  ANDN U4001 ( .B(y[1686]), .A(x[1686]), .Z(n13887) );
  NANDN U4002 ( .A(y[1686]), .B(x[1686]), .Z(n4992) );
  ANDN U4003 ( .B(y[1685]), .A(x[1685]), .Z(n9629) );
  NANDN U4004 ( .A(x[1684]), .B(y[1684]), .Z(n3252) );
  NANDN U4005 ( .A(n9629), .B(n3252), .Z(n13882) );
  NANDN U4006 ( .A(y[1683]), .B(x[1683]), .Z(n9626) );
  XOR U4007 ( .A(x[1684]), .B(y[1684]), .Z(n9628) );
  ANDN U4008 ( .B(n9626), .A(n9628), .Z(n13881) );
  ANDN U4009 ( .B(y[1683]), .A(x[1683]), .Z(n9627) );
  NANDN U4010 ( .A(x[1682]), .B(y[1682]), .Z(n3253) );
  NANDN U4011 ( .A(n9627), .B(n3253), .Z(n13879) );
  XNOR U4012 ( .A(x[1682]), .B(y[1682]), .Z(n9624) );
  NANDN U4013 ( .A(y[1681]), .B(x[1681]), .Z(n9623) );
  AND U4014 ( .A(n9624), .B(n9623), .Z(n13877) );
  ANDN U4015 ( .B(y[1680]), .A(x[1680]), .Z(n9622) );
  ANDN U4016 ( .B(y[1681]), .A(x[1681]), .Z(n9625) );
  OR U4017 ( .A(n9622), .B(n9625), .Z(n13875) );
  NANDN U4018 ( .A(y[1680]), .B(x[1680]), .Z(n13873) );
  ANDN U4019 ( .B(y[1678]), .A(x[1678]), .Z(n4997) );
  NANDN U4020 ( .A(y[1675]), .B(x[1675]), .Z(n3255) );
  NANDN U4021 ( .A(y[1676]), .B(x[1676]), .Z(n3254) );
  NAND U4022 ( .A(n3255), .B(n3254), .Z(n13861) );
  IV U4023 ( .A(n13861), .Z(n9619) );
  NANDN U4024 ( .A(x[1675]), .B(y[1675]), .Z(n3257) );
  NANDN U4025 ( .A(x[1674]), .B(y[1674]), .Z(n3256) );
  AND U4026 ( .A(n3257), .B(n3256), .Z(n13859) );
  NANDN U4027 ( .A(y[1673]), .B(x[1673]), .Z(n3259) );
  NANDN U4028 ( .A(y[1674]), .B(x[1674]), .Z(n3258) );
  AND U4029 ( .A(n3259), .B(n3258), .Z(n13857) );
  IV U4030 ( .A(n13857), .Z(n9613) );
  NANDN U4031 ( .A(x[1672]), .B(y[1672]), .Z(n3260) );
  ANDN U4032 ( .B(y[1673]), .A(x[1673]), .Z(n9612) );
  ANDN U4033 ( .B(n3260), .A(n9612), .Z(n13855) );
  NANDN U4034 ( .A(y[1671]), .B(x[1671]), .Z(n4999) );
  NANDN U4035 ( .A(y[1672]), .B(x[1672]), .Z(n9611) );
  AND U4036 ( .A(n4999), .B(n9611), .Z(n13852) );
  ANDN U4037 ( .B(y[1669]), .A(x[1669]), .Z(n13847) );
  NANDN U4038 ( .A(y[1667]), .B(x[1667]), .Z(n5005) );
  ANDN U4039 ( .B(y[1666]), .A(x[1666]), .Z(n5006) );
  NANDN U4040 ( .A(y[1665]), .B(x[1665]), .Z(n5009) );
  ANDN U4041 ( .B(y[1664]), .A(x[1664]), .Z(n13835) );
  XNOR U4042 ( .A(x[1660]), .B(y[1660]), .Z(n9583) );
  NANDN U4043 ( .A(y[1659]), .B(x[1659]), .Z(n5011) );
  AND U4044 ( .A(n9583), .B(n5011), .Z(n13825) );
  ANDN U4045 ( .B(y[1658]), .A(x[1658]), .Z(n9577) );
  ANDN U4046 ( .B(y[1659]), .A(x[1659]), .Z(n9582) );
  OR U4047 ( .A(n9577), .B(n9582), .Z(n13823) );
  NANDN U4048 ( .A(y[1658]), .B(x[1658]), .Z(n13821) );
  NANDN U4049 ( .A(y[1656]), .B(x[1656]), .Z(n5013) );
  NANDN U4050 ( .A(y[1655]), .B(x[1655]), .Z(n13813) );
  ANDN U4051 ( .B(y[1654]), .A(x[1654]), .Z(n13810) );
  XNOR U4052 ( .A(x[1654]), .B(y[1654]), .Z(n5017) );
  NANDN U4053 ( .A(y[1653]), .B(x[1653]), .Z(n9566) );
  AND U4054 ( .A(n5017), .B(n9566), .Z(n13809) );
  NANDN U4055 ( .A(x[1652]), .B(y[1652]), .Z(n5018) );
  NANDN U4056 ( .A(x[1653]), .B(y[1653]), .Z(n5016) );
  NAND U4057 ( .A(n5018), .B(n5016), .Z(n13807) );
  NANDN U4058 ( .A(y[1651]), .B(x[1651]), .Z(n5020) );
  NANDN U4059 ( .A(y[1652]), .B(x[1652]), .Z(n9568) );
  AND U4060 ( .A(n5020), .B(n9568), .Z(n13805) );
  ANDN U4061 ( .B(y[1650]), .A(x[1650]), .Z(n9564) );
  NANDN U4062 ( .A(x[1651]), .B(y[1651]), .Z(n5019) );
  NANDN U4063 ( .A(n9564), .B(n5019), .Z(n13803) );
  NANDN U4064 ( .A(y[1649]), .B(x[1649]), .Z(n5022) );
  NANDN U4065 ( .A(y[1650]), .B(x[1650]), .Z(n5021) );
  AND U4066 ( .A(n5022), .B(n5021), .Z(n13801) );
  ANDN U4067 ( .B(y[1649]), .A(x[1649]), .Z(n9565) );
  NANDN U4068 ( .A(x[1648]), .B(y[1648]), .Z(n5023) );
  NANDN U4069 ( .A(n9565), .B(n5023), .Z(n13799) );
  NANDN U4070 ( .A(y[1648]), .B(x[1648]), .Z(n13792) );
  ANDN U4071 ( .B(y[1646]), .A(x[1646]), .Z(n9562) );
  NANDN U4072 ( .A(x[1647]), .B(y[1647]), .Z(n13794) );
  NANDN U4073 ( .A(n9562), .B(n13794), .Z(n13791) );
  NANDN U4074 ( .A(y[1645]), .B(x[1645]), .Z(n13789) );
  ANDN U4075 ( .B(y[1644]), .A(x[1644]), .Z(n9560) );
  ANDN U4076 ( .B(y[1645]), .A(x[1645]), .Z(n9563) );
  NOR U4077 ( .A(n9560), .B(n9563), .Z(n13787) );
  NANDN U4078 ( .A(y[1643]), .B(x[1643]), .Z(n9558) );
  NANDN U4079 ( .A(y[1644]), .B(x[1644]), .Z(n9561) );
  AND U4080 ( .A(n9558), .B(n9561), .Z(n13785) );
  ANDN U4081 ( .B(y[1642]), .A(x[1642]), .Z(n5026) );
  NANDN U4082 ( .A(y[1642]), .B(x[1642]), .Z(n13780) );
  NANDN U4083 ( .A(x[1641]), .B(y[1641]), .Z(n5027) );
  NANDN U4084 ( .A(y[1639]), .B(x[1639]), .Z(n5033) );
  NANDN U4085 ( .A(x[1638]), .B(y[1638]), .Z(n9557) );
  NANDN U4086 ( .A(y[1638]), .B(x[1638]), .Z(n5032) );
  ANDN U4087 ( .B(y[1636]), .A(x[1636]), .Z(n9554) );
  NANDN U4088 ( .A(y[1637]), .B(x[1637]), .Z(n3262) );
  AND U4089 ( .A(n9554), .B(n3262), .Z(n13771) );
  NANDN U4090 ( .A(y[1636]), .B(x[1636]), .Z(n3261) );
  AND U4091 ( .A(n3262), .B(n3261), .Z(n13767) );
  IV U4092 ( .A(n13767), .Z(n9555) );
  NANDN U4093 ( .A(y[1635]), .B(x[1635]), .Z(n5035) );
  NANDN U4094 ( .A(x[1634]), .B(y[1634]), .Z(n5036) );
  NANDN U4095 ( .A(y[1633]), .B(x[1633]), .Z(n5039) );
  ANDN U4096 ( .B(y[1632]), .A(x[1632]), .Z(n5040) );
  NANDN U4097 ( .A(y[1631]), .B(x[1631]), .Z(n9552) );
  NANDN U4098 ( .A(x[1630]), .B(y[1630]), .Z(n13753) );
  NANDN U4099 ( .A(y[1630]), .B(x[1630]), .Z(n9551) );
  NANDN U4100 ( .A(x[1628]), .B(y[1628]), .Z(n9548) );
  NANDN U4101 ( .A(x[1629]), .B(y[1629]), .Z(n5042) );
  NAND U4102 ( .A(n9548), .B(n5042), .Z(n13749) );
  NANDN U4103 ( .A(y[1627]), .B(x[1627]), .Z(n5043) );
  ANDN U4104 ( .B(x[1628]), .A(y[1628]), .Z(n13747) );
  NANDN U4105 ( .A(x[1627]), .B(y[1627]), .Z(n13744) );
  NANDN U4106 ( .A(y[1626]), .B(x[1626]), .Z(n5044) );
  ANDN U4107 ( .B(y[1624]), .A(x[1624]), .Z(n13737) );
  NANDN U4108 ( .A(y[1623]), .B(x[1623]), .Z(n13734) );
  NANDN U4109 ( .A(y[1624]), .B(x[1624]), .Z(n5048) );
  NANDN U4110 ( .A(x[1622]), .B(y[1622]), .Z(n5050) );
  NANDN U4111 ( .A(x[1623]), .B(y[1623]), .Z(n5049) );
  NAND U4112 ( .A(n5050), .B(n5049), .Z(n13732) );
  ANDN U4113 ( .B(x[1621]), .A(y[1621]), .Z(n9546) );
  ANDN U4114 ( .B(x[1622]), .A(y[1622]), .Z(n9547) );
  NOR U4115 ( .A(n9546), .B(n9547), .Z(n13731) );
  NANDN U4116 ( .A(x[1620]), .B(y[1620]), .Z(n9544) );
  NANDN U4117 ( .A(x[1621]), .B(y[1621]), .Z(n5051) );
  NAND U4118 ( .A(n9544), .B(n5051), .Z(n13729) );
  ANDN U4119 ( .B(x[1620]), .A(y[1620]), .Z(n13727) );
  NANDN U4120 ( .A(y[1618]), .B(x[1618]), .Z(n13721) );
  NANDN U4121 ( .A(y[1619]), .B(x[1619]), .Z(n13724) );
  AND U4122 ( .A(n13721), .B(n13724), .Z(n9543) );
  NANDN U4123 ( .A(y[1617]), .B(x[1617]), .Z(n5053) );
  NANDN U4124 ( .A(x[1616]), .B(y[1616]), .Z(n13714) );
  NANDN U4125 ( .A(y[1616]), .B(x[1616]), .Z(n5052) );
  NANDN U4126 ( .A(x[1614]), .B(y[1614]), .Z(n5055) );
  NANDN U4127 ( .A(x[1615]), .B(y[1615]), .Z(n5054) );
  NAND U4128 ( .A(n5055), .B(n5054), .Z(n13711) );
  NANDN U4129 ( .A(y[1613]), .B(x[1613]), .Z(n5057) );
  NANDN U4130 ( .A(y[1612]), .B(x[1612]), .Z(n5056) );
  NANDN U4131 ( .A(y[1611]), .B(x[1611]), .Z(n9541) );
  ANDN U4132 ( .B(y[1610]), .A(x[1610]), .Z(n9538) );
  NANDN U4133 ( .A(y[1610]), .B(x[1610]), .Z(n9540) );
  ANDN U4134 ( .B(y[1608]), .A(x[1608]), .Z(n13695) );
  NANDN U4135 ( .A(x[1606]), .B(y[1606]), .Z(n9536) );
  NANDN U4136 ( .A(x[1607]), .B(y[1607]), .Z(n5062) );
  NAND U4137 ( .A(n9536), .B(n5062), .Z(n13690) );
  NANDN U4138 ( .A(x[1604]), .B(y[1604]), .Z(n13682) );
  IV U4139 ( .A(n13682), .Z(n5065) );
  NANDN U4140 ( .A(x[1605]), .B(y[1605]), .Z(n13687) );
  ANDN U4141 ( .B(x[1603]), .A(y[1603]), .Z(n13680) );
  NANDN U4142 ( .A(y[1604]), .B(x[1604]), .Z(n5064) );
  NANDN U4143 ( .A(x[1602]), .B(y[1602]), .Z(n9535) );
  NANDN U4144 ( .A(x[1603]), .B(y[1603]), .Z(n5066) );
  NAND U4145 ( .A(n9535), .B(n5066), .Z(n13679) );
  ANDN U4146 ( .B(x[1602]), .A(y[1602]), .Z(n13677) );
  NANDN U4147 ( .A(y[1601]), .B(x[1601]), .Z(n4597) );
  NANDN U4148 ( .A(y[1600]), .B(x[1600]), .Z(n3263) );
  NAND U4149 ( .A(n4597), .B(n3263), .Z(n13672) );
  NANDN U4150 ( .A(y[1599]), .B(x[1599]), .Z(n13668) );
  NANDN U4151 ( .A(y[1598]), .B(x[1598]), .Z(n5067) );
  NANDN U4152 ( .A(y[1597]), .B(x[1597]), .Z(n9531) );
  ANDN U4153 ( .B(y[1597]), .A(x[1597]), .Z(n13663) );
  NANDN U4154 ( .A(y[1596]), .B(x[1596]), .Z(n9532) );
  ANDN U4155 ( .B(y[1594]), .A(x[1594]), .Z(n5073) );
  NANDN U4156 ( .A(y[1593]), .B(x[1593]), .Z(n5075) );
  ANDN U4157 ( .B(y[1592]), .A(x[1592]), .Z(n13651) );
  NANDN U4158 ( .A(y[1592]), .B(x[1592]), .Z(n5076) );
  NANDN U4159 ( .A(x[1591]), .B(y[1591]), .Z(n4594) );
  NANDN U4160 ( .A(x[1590]), .B(y[1590]), .Z(n3264) );
  NAND U4161 ( .A(n4594), .B(n3264), .Z(n13647) );
  IV U4162 ( .A(n13647), .Z(n4593) );
  NANDN U4163 ( .A(y[1589]), .B(x[1589]), .Z(n13644) );
  IV U4164 ( .A(n13644), .Z(n9529) );
  NANDN U4165 ( .A(x[1589]), .B(y[1589]), .Z(n3266) );
  NANDN U4166 ( .A(x[1588]), .B(y[1588]), .Z(n3265) );
  NAND U4167 ( .A(n3266), .B(n3265), .Z(n13641) );
  NANDN U4168 ( .A(y[1587]), .B(x[1587]), .Z(n3268) );
  NANDN U4169 ( .A(y[1588]), .B(x[1588]), .Z(n3267) );
  AND U4170 ( .A(n3268), .B(n3267), .Z(n13638) );
  NANDN U4171 ( .A(x[1587]), .B(y[1587]), .Z(n3270) );
  NANDN U4172 ( .A(x[1586]), .B(y[1586]), .Z(n3269) );
  NAND U4173 ( .A(n3270), .B(n3269), .Z(n13636) );
  NANDN U4174 ( .A(y[1583]), .B(x[1583]), .Z(n3272) );
  ANDN U4175 ( .B(x[1584]), .A(y[1584]), .Z(n3271) );
  ANDN U4176 ( .B(n3272), .A(n3271), .Z(n3276) );
  XNOR U4177 ( .A(x[1583]), .B(y[1583]), .Z(n3274) );
  ANDN U4178 ( .B(x[1582]), .A(y[1582]), .Z(n3273) );
  NAND U4179 ( .A(n3274), .B(n3273), .Z(n3275) );
  AND U4180 ( .A(n3276), .B(n3275), .Z(n13630) );
  NANDN U4181 ( .A(x[1580]), .B(y[1580]), .Z(n9524) );
  ANDN U4182 ( .B(x[1581]), .A(y[1581]), .Z(n3281) );
  NANDN U4183 ( .A(x[1582]), .B(y[1582]), .Z(n3278) );
  NANDN U4184 ( .A(x[1581]), .B(y[1581]), .Z(n3277) );
  AND U4185 ( .A(n3278), .B(n3277), .Z(n3280) );
  NANDN U4186 ( .A(x[1583]), .B(y[1583]), .Z(n3279) );
  NAND U4187 ( .A(n3280), .B(n3279), .Z(n9525) );
  NANDN U4188 ( .A(y[1580]), .B(x[1580]), .Z(n3282) );
  ANDN U4189 ( .B(n3282), .A(n3281), .Z(n13626) );
  NANDN U4190 ( .A(y[1579]), .B(x[1579]), .Z(n9522) );
  ANDN U4191 ( .B(y[1578]), .A(x[1578]), .Z(n13621) );
  NANDN U4192 ( .A(x[1579]), .B(y[1579]), .Z(n13625) );
  NANDN U4193 ( .A(n13621), .B(n13625), .Z(n4577) );
  NANDN U4194 ( .A(y[1575]), .B(x[1575]), .Z(n9519) );
  ANDN U4195 ( .B(x[1576]), .A(y[1576]), .Z(n13615) );
  ANDN U4196 ( .B(n9519), .A(n13615), .Z(n4572) );
  NANDN U4197 ( .A(x[1575]), .B(y[1575]), .Z(n13612) );
  NANDN U4198 ( .A(y[1574]), .B(x[1574]), .Z(n9518) );
  NANDN U4199 ( .A(x[1573]), .B(y[1573]), .Z(n5080) );
  NANDN U4200 ( .A(x[1572]), .B(y[1572]), .Z(n3283) );
  NAND U4201 ( .A(n5080), .B(n3283), .Z(n13605) );
  NANDN U4202 ( .A(y[1571]), .B(x[1571]), .Z(n13602) );
  NANDN U4203 ( .A(x[1570]), .B(y[1570]), .Z(n9517) );
  NANDN U4204 ( .A(x[1571]), .B(y[1571]), .Z(n5084) );
  NAND U4205 ( .A(n9517), .B(n5084), .Z(n13600) );
  NANDN U4206 ( .A(y[1570]), .B(x[1570]), .Z(n13598) );
  ANDN U4207 ( .B(y[1568]), .A(x[1568]), .Z(n13593) );
  NANDN U4208 ( .A(x[1569]), .B(y[1569]), .Z(n13597) );
  NANDN U4209 ( .A(y[1567]), .B(x[1567]), .Z(n13591) );
  NANDN U4210 ( .A(x[1567]), .B(y[1567]), .Z(n3285) );
  NANDN U4211 ( .A(x[1566]), .B(y[1566]), .Z(n3284) );
  NAND U4212 ( .A(n3285), .B(n3284), .Z(n13589) );
  NANDN U4213 ( .A(y[1566]), .B(x[1566]), .Z(n3287) );
  NANDN U4214 ( .A(y[1565]), .B(x[1565]), .Z(n3286) );
  AND U4215 ( .A(n3287), .B(n3286), .Z(n5090) );
  NANDN U4216 ( .A(x[1562]), .B(y[1562]), .Z(n9514) );
  NANDN U4217 ( .A(x[1563]), .B(y[1563]), .Z(n5091) );
  NAND U4218 ( .A(n9514), .B(n5091), .Z(n13581) );
  ANDN U4219 ( .B(x[1561]), .A(y[1561]), .Z(n5096) );
  NANDN U4220 ( .A(x[1561]), .B(y[1561]), .Z(n5093) );
  NANDN U4221 ( .A(x[1560]), .B(y[1560]), .Z(n3288) );
  AND U4222 ( .A(n5093), .B(n3288), .Z(n13575) );
  ANDN U4223 ( .B(x[1559]), .A(y[1559]), .Z(n13573) );
  NANDN U4224 ( .A(x[1558]), .B(y[1558]), .Z(n5098) );
  NANDN U4225 ( .A(x[1559]), .B(y[1559]), .Z(n5097) );
  AND U4226 ( .A(n5098), .B(n5097), .Z(n13571) );
  ANDN U4227 ( .B(x[1557]), .A(y[1557]), .Z(n9502) );
  ANDN U4228 ( .B(x[1558]), .A(y[1558]), .Z(n9508) );
  OR U4229 ( .A(n9502), .B(n9508), .Z(n13569) );
  NANDN U4230 ( .A(x[1556]), .B(y[1556]), .Z(n9498) );
  NANDN U4231 ( .A(x[1557]), .B(y[1557]), .Z(n5099) );
  AND U4232 ( .A(n9498), .B(n5099), .Z(n13567) );
  ANDN U4233 ( .B(x[1556]), .A(y[1556]), .Z(n9503) );
  NANDN U4234 ( .A(y[1555]), .B(x[1555]), .Z(n5100) );
  NANDN U4235 ( .A(n9503), .B(n5100), .Z(n13565) );
  NANDN U4236 ( .A(x[1554]), .B(y[1554]), .Z(n5102) );
  NANDN U4237 ( .A(x[1555]), .B(y[1555]), .Z(n9497) );
  NAND U4238 ( .A(n5102), .B(n9497), .Z(n13563) );
  NANDN U4239 ( .A(y[1553]), .B(x[1553]), .Z(n5104) );
  NANDN U4240 ( .A(y[1554]), .B(x[1554]), .Z(n5101) );
  AND U4241 ( .A(n5104), .B(n5101), .Z(n13560) );
  NANDN U4242 ( .A(y[1551]), .B(x[1551]), .Z(n5108) );
  NANDN U4243 ( .A(y[1552]), .B(x[1552]), .Z(n13557) );
  IV U4244 ( .A(n13557), .Z(n5105) );
  ANDN U4245 ( .B(n5108), .A(n5105), .Z(n4565) );
  ANDN U4246 ( .B(y[1551]), .A(x[1551]), .Z(n13555) );
  NANDN U4247 ( .A(x[1550]), .B(y[1550]), .Z(n5110) );
  ANDN U4248 ( .B(x[1549]), .A(y[1549]), .Z(n5112) );
  NANDN U4249 ( .A(x[1549]), .B(y[1549]), .Z(n5109) );
  ANDN U4250 ( .B(x[1548]), .A(y[1548]), .Z(n5111) );
  NANDN U4251 ( .A(x[1547]), .B(y[1547]), .Z(n9487) );
  ANDN U4252 ( .B(y[1546]), .A(x[1546]), .Z(n9485) );
  NANDN U4253 ( .A(y[1547]), .B(x[1547]), .Z(n3290) );
  NAND U4254 ( .A(n9485), .B(n3290), .Z(n10187) );
  NANDN U4255 ( .A(y[1546]), .B(x[1546]), .Z(n3289) );
  AND U4256 ( .A(n3290), .B(n3289), .Z(n9486) );
  NANDN U4257 ( .A(y[1545]), .B(x[1545]), .Z(n9484) );
  NAND U4258 ( .A(n9486), .B(n9484), .Z(n13544) );
  NANDN U4259 ( .A(x[1544]), .B(y[1544]), .Z(n13538) );
  ANDN U4260 ( .B(y[1545]), .A(x[1545]), .Z(n13542) );
  NANDN U4261 ( .A(y[1544]), .B(x[1544]), .Z(n13541) );
  NANDN U4262 ( .A(x[1542]), .B(y[1542]), .Z(n5116) );
  NANDN U4263 ( .A(x[1543]), .B(y[1543]), .Z(n5113) );
  AND U4264 ( .A(n5116), .B(n5113), .Z(n13535) );
  ANDN U4265 ( .B(x[1542]), .A(y[1542]), .Z(n13533) );
  IV U4266 ( .A(n13533), .Z(n5114) );
  NANDN U4267 ( .A(x[1540]), .B(y[1540]), .Z(n5120) );
  NANDN U4268 ( .A(y[1540]), .B(x[1540]), .Z(n5118) );
  ANDN U4269 ( .B(x[1539]), .A(y[1539]), .Z(n5121) );
  NANDN U4270 ( .A(x[1538]), .B(y[1538]), .Z(n13522) );
  NANDN U4271 ( .A(y[1538]), .B(x[1538]), .Z(n5122) );
  NANDN U4272 ( .A(x[1536]), .B(y[1536]), .Z(n5125) );
  NANDN U4273 ( .A(x[1537]), .B(y[1537]), .Z(n5123) );
  NAND U4274 ( .A(n5125), .B(n5123), .Z(n13519) );
  NANDN U4275 ( .A(y[1535]), .B(x[1535]), .Z(n5126) );
  NANDN U4276 ( .A(x[1534]), .B(y[1534]), .Z(n13510) );
  NANDN U4277 ( .A(x[1535]), .B(y[1535]), .Z(n13515) );
  NANDN U4278 ( .A(x[1532]), .B(y[1532]), .Z(n5128) );
  NANDN U4279 ( .A(x[1533]), .B(y[1533]), .Z(n9482) );
  AND U4280 ( .A(n5128), .B(n9482), .Z(n13507) );
  ANDN U4281 ( .B(x[1532]), .A(y[1532]), .Z(n13505) );
  NANDN U4282 ( .A(x[1530]), .B(y[1530]), .Z(n5132) );
  NANDN U4283 ( .A(y[1530]), .B(x[1530]), .Z(n5129) );
  ANDN U4284 ( .B(x[1529]), .A(y[1529]), .Z(n5134) );
  ANDN U4285 ( .B(y[1528]), .A(x[1528]), .Z(n13495) );
  NANDN U4286 ( .A(y[1528]), .B(x[1528]), .Z(n5133) );
  NANDN U4287 ( .A(x[1526]), .B(y[1526]), .Z(n9477) );
  NANDN U4288 ( .A(x[1527]), .B(y[1527]), .Z(n5135) );
  NAND U4289 ( .A(n9477), .B(n5135), .Z(n13491) );
  NANDN U4290 ( .A(y[1525]), .B(x[1525]), .Z(n5137) );
  ANDN U4291 ( .B(x[1526]), .A(y[1526]), .Z(n9478) );
  ANDN U4292 ( .B(n5137), .A(n9478), .Z(n13489) );
  NANDN U4293 ( .A(x[1524]), .B(y[1524]), .Z(n5138) );
  NANDN U4294 ( .A(x[1525]), .B(y[1525]), .Z(n9476) );
  NAND U4295 ( .A(n5138), .B(n9476), .Z(n13487) );
  NANDN U4296 ( .A(y[1523]), .B(x[1523]), .Z(n5140) );
  NANDN U4297 ( .A(y[1524]), .B(x[1524]), .Z(n5136) );
  AND U4298 ( .A(n5140), .B(n5136), .Z(n13485) );
  ANDN U4299 ( .B(y[1522]), .A(x[1522]), .Z(n9475) );
  NANDN U4300 ( .A(x[1523]), .B(y[1523]), .Z(n5139) );
  NANDN U4301 ( .A(n9475), .B(n5139), .Z(n13483) );
  NANDN U4302 ( .A(y[1522]), .B(x[1522]), .Z(n13480) );
  ANDN U4303 ( .B(y[1521]), .A(x[1521]), .Z(n13479) );
  NANDN U4304 ( .A(y[1517]), .B(x[1517]), .Z(n3292) );
  NANDN U4305 ( .A(y[1518]), .B(x[1518]), .Z(n3291) );
  NAND U4306 ( .A(n3292), .B(n3291), .Z(n9469) );
  NANDN U4307 ( .A(x[1517]), .B(y[1517]), .Z(n9466) );
  NANDN U4308 ( .A(x[1516]), .B(y[1516]), .Z(n3293) );
  NAND U4309 ( .A(n9466), .B(n3293), .Z(n5144) );
  ANDN U4310 ( .B(x[1515]), .A(y[1515]), .Z(n5145) );
  NANDN U4311 ( .A(x[1515]), .B(y[1515]), .Z(n3295) );
  NANDN U4312 ( .A(x[1514]), .B(y[1514]), .Z(n3294) );
  NAND U4313 ( .A(n3295), .B(n3294), .Z(n5143) );
  NANDN U4314 ( .A(x[1513]), .B(y[1513]), .Z(n4554) );
  XNOR U4315 ( .A(x[1513]), .B(y[1513]), .Z(n3297) );
  NANDN U4316 ( .A(y[1512]), .B(x[1512]), .Z(n3296) );
  NAND U4317 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U4318 ( .A(n4554), .B(n3298), .Z(n3300) );
  NANDN U4319 ( .A(y[1514]), .B(x[1514]), .Z(n3299) );
  AND U4320 ( .A(n3300), .B(n3299), .Z(n5146) );
  NANDN U4321 ( .A(x[1509]), .B(y[1509]), .Z(n5148) );
  NANDN U4322 ( .A(x[1508]), .B(y[1508]), .Z(n3302) );
  NANDN U4323 ( .A(x[1507]), .B(y[1507]), .Z(n3301) );
  NAND U4324 ( .A(n3302), .B(n3301), .Z(n9461) );
  ANDN U4325 ( .B(n5148), .A(n9461), .Z(n13463) );
  NANDN U4326 ( .A(y[1506]), .B(x[1506]), .Z(n3304) );
  NANDN U4327 ( .A(y[1507]), .B(x[1507]), .Z(n3303) );
  AND U4328 ( .A(n3304), .B(n3303), .Z(n13460) );
  IV U4329 ( .A(n13460), .Z(n9460) );
  NANDN U4330 ( .A(x[1506]), .B(y[1506]), .Z(n3306) );
  NANDN U4331 ( .A(x[1505]), .B(y[1505]), .Z(n3305) );
  NAND U4332 ( .A(n3306), .B(n3305), .Z(n13458) );
  ANDN U4333 ( .B(x[1505]), .A(y[1505]), .Z(n9458) );
  NANDN U4334 ( .A(x[1504]), .B(y[1504]), .Z(n5150) );
  ANDN U4335 ( .B(x[1504]), .A(y[1504]), .Z(n9459) );
  IV U4336 ( .A(n9459), .Z(n4540) );
  ANDN U4337 ( .B(y[1502]), .A(x[1502]), .Z(n13451) );
  IV U4338 ( .A(n13451), .Z(n4535) );
  NANDN U4339 ( .A(y[1502]), .B(x[1502]), .Z(n13448) );
  IV U4340 ( .A(n13448), .Z(n4533) );
  NANDN U4341 ( .A(x[1500]), .B(y[1500]), .Z(n13442) );
  NANDN U4342 ( .A(x[1501]), .B(y[1501]), .Z(n13447) );
  NAND U4343 ( .A(n13442), .B(n13447), .Z(n4530) );
  ANDN U4344 ( .B(x[1499]), .A(y[1499]), .Z(n13441) );
  XNOR U4345 ( .A(x[1500]), .B(y[1500]), .Z(n5154) );
  NANDN U4346 ( .A(x[1498]), .B(y[1498]), .Z(n5156) );
  NANDN U4347 ( .A(x[1499]), .B(y[1499]), .Z(n5155) );
  NAND U4348 ( .A(n5156), .B(n5155), .Z(n13439) );
  ANDN U4349 ( .B(x[1498]), .A(y[1498]), .Z(n13437) );
  ANDN U4350 ( .B(y[1496]), .A(x[1496]), .Z(n13431) );
  NANDN U4351 ( .A(y[1495]), .B(x[1495]), .Z(n13428) );
  NANDN U4352 ( .A(y[1496]), .B(x[1496]), .Z(n5158) );
  NANDN U4353 ( .A(x[1494]), .B(y[1494]), .Z(n9456) );
  NANDN U4354 ( .A(x[1495]), .B(y[1495]), .Z(n5159) );
  NAND U4355 ( .A(n9456), .B(n5159), .Z(n13426) );
  NANDN U4356 ( .A(y[1493]), .B(x[1493]), .Z(n3308) );
  NANDN U4357 ( .A(y[1494]), .B(x[1494]), .Z(n3307) );
  NAND U4358 ( .A(n3308), .B(n3307), .Z(n13425) );
  NANDN U4359 ( .A(x[1493]), .B(y[1493]), .Z(n3310) );
  NANDN U4360 ( .A(x[1492]), .B(y[1492]), .Z(n3309) );
  AND U4361 ( .A(n3310), .B(n3309), .Z(n13423) );
  NANDN U4362 ( .A(y[1491]), .B(x[1491]), .Z(n3312) );
  NANDN U4363 ( .A(y[1492]), .B(x[1492]), .Z(n3311) );
  NAND U4364 ( .A(n3312), .B(n3311), .Z(n13421) );
  NANDN U4365 ( .A(x[1491]), .B(y[1491]), .Z(n3314) );
  NANDN U4366 ( .A(x[1490]), .B(y[1490]), .Z(n3313) );
  AND U4367 ( .A(n3314), .B(n3313), .Z(n5162) );
  NANDN U4368 ( .A(y[1489]), .B(x[1489]), .Z(n3315) );
  ANDN U4369 ( .B(x[1490]), .A(y[1490]), .Z(n5161) );
  ANDN U4370 ( .B(n3315), .A(n5161), .Z(n3319) );
  NANDN U4371 ( .A(x[1489]), .B(y[1489]), .Z(n5160) );
  NANDN U4372 ( .A(x[1488]), .B(y[1488]), .Z(n9455) );
  NAND U4373 ( .A(n5160), .B(n9455), .Z(n3316) );
  NAND U4374 ( .A(n3319), .B(n3316), .Z(n3317) );
  AND U4375 ( .A(n5162), .B(n3317), .Z(n13419) );
  NANDN U4376 ( .A(y[1488]), .B(x[1488]), .Z(n3318) );
  AND U4377 ( .A(n3319), .B(n3318), .Z(n13416) );
  ANDN U4378 ( .B(y[1487]), .A(x[1487]), .Z(n13414) );
  NANDN U4379 ( .A(y[1487]), .B(x[1487]), .Z(n3321) );
  NANDN U4380 ( .A(y[1486]), .B(x[1486]), .Z(n3320) );
  NAND U4381 ( .A(n3321), .B(n3320), .Z(n13413) );
  NANDN U4382 ( .A(x[1486]), .B(y[1486]), .Z(n3323) );
  NANDN U4383 ( .A(x[1485]), .B(y[1485]), .Z(n3322) );
  AND U4384 ( .A(n3323), .B(n3322), .Z(n9454) );
  NANDN U4385 ( .A(x[1484]), .B(y[1484]), .Z(n9450) );
  ANDN U4386 ( .B(x[1485]), .A(y[1485]), .Z(n3324) );
  NANDN U4387 ( .A(y[1484]), .B(x[1484]), .Z(n3325) );
  ANDN U4388 ( .B(n3325), .A(n3324), .Z(n9452) );
  NANDN U4389 ( .A(y[1482]), .B(x[1482]), .Z(n3327) );
  NANDN U4390 ( .A(y[1483]), .B(x[1483]), .Z(n3326) );
  AND U4391 ( .A(n3327), .B(n3326), .Z(n9449) );
  NANDN U4392 ( .A(x[1483]), .B(y[1483]), .Z(n9451) );
  NANDN U4393 ( .A(n9449), .B(n9451), .Z(n3328) );
  AND U4394 ( .A(n9452), .B(n3328), .Z(n13409) );
  ANDN U4395 ( .B(y[1480]), .A(x[1480]), .Z(n9447) );
  NANDN U4396 ( .A(y[1481]), .B(x[1481]), .Z(n3334) );
  NAND U4397 ( .A(n9447), .B(n3334), .Z(n3329) );
  AND U4398 ( .A(n3329), .B(n9451), .Z(n3332) );
  NANDN U4399 ( .A(x[1481]), .B(y[1481]), .Z(n3331) );
  NANDN U4400 ( .A(x[1482]), .B(y[1482]), .Z(n3330) );
  NAND U4401 ( .A(n3331), .B(n3330), .Z(n9448) );
  ANDN U4402 ( .B(n3332), .A(n9448), .Z(n13407) );
  NANDN U4403 ( .A(y[1480]), .B(x[1480]), .Z(n3333) );
  NAND U4404 ( .A(n3334), .B(n3333), .Z(n13405) );
  NANDN U4405 ( .A(x[1478]), .B(y[1478]), .Z(n13398) );
  NANDN U4406 ( .A(x[1479]), .B(y[1479]), .Z(n13403) );
  NANDN U4407 ( .A(y[1477]), .B(x[1477]), .Z(n13397) );
  NANDN U4408 ( .A(x[1477]), .B(y[1477]), .Z(n3336) );
  NANDN U4409 ( .A(x[1476]), .B(y[1476]), .Z(n3335) );
  NAND U4410 ( .A(n3336), .B(n3335), .Z(n13395) );
  NANDN U4411 ( .A(y[1476]), .B(x[1476]), .Z(n3338) );
  NANDN U4412 ( .A(y[1475]), .B(x[1475]), .Z(n3337) );
  AND U4413 ( .A(n3338), .B(n3337), .Z(n5168) );
  NANDN U4414 ( .A(x[1474]), .B(y[1474]), .Z(n3339) );
  ANDN U4415 ( .B(y[1475]), .A(x[1475]), .Z(n5166) );
  ANDN U4416 ( .B(n3339), .A(n5166), .Z(n13390) );
  NANDN U4417 ( .A(y[1473]), .B(x[1473]), .Z(n13389) );
  NANDN U4418 ( .A(x[1472]), .B(y[1472]), .Z(n9446) );
  NANDN U4419 ( .A(x[1473]), .B(y[1473]), .Z(n5169) );
  NAND U4420 ( .A(n9446), .B(n5169), .Z(n13387) );
  NANDN U4421 ( .A(y[1471]), .B(x[1471]), .Z(n9443) );
  ANDN U4422 ( .B(y[1470]), .A(x[1470]), .Z(n9441) );
  NANDN U4423 ( .A(y[1469]), .B(x[1469]), .Z(n5170) );
  ANDN U4424 ( .B(y[1468]), .A(x[1468]), .Z(n13375) );
  NANDN U4425 ( .A(y[1468]), .B(x[1468]), .Z(n5171) );
  NANDN U4426 ( .A(x[1467]), .B(y[1467]), .Z(n3341) );
  NANDN U4427 ( .A(x[1466]), .B(y[1466]), .Z(n3340) );
  NAND U4428 ( .A(n3341), .B(n3340), .Z(n13370) );
  NANDN U4429 ( .A(y[1466]), .B(x[1466]), .Z(n3343) );
  NANDN U4430 ( .A(y[1465]), .B(x[1465]), .Z(n3342) );
  AND U4431 ( .A(n3343), .B(n3342), .Z(n5175) );
  NANDN U4432 ( .A(y[1464]), .B(x[1464]), .Z(n5172) );
  ANDN U4433 ( .B(x[1463]), .A(y[1463]), .Z(n13365) );
  NANDN U4434 ( .A(x[1462]), .B(y[1462]), .Z(n5177) );
  ANDN U4435 ( .B(y[1463]), .A(x[1463]), .Z(n9440) );
  ANDN U4436 ( .B(n5177), .A(n9440), .Z(n13363) );
  NANDN U4437 ( .A(y[1461]), .B(x[1461]), .Z(n9437) );
  ANDN U4438 ( .B(x[1462]), .A(y[1462]), .Z(n9439) );
  ANDN U4439 ( .B(n9437), .A(n9439), .Z(n13361) );
  NANDN U4440 ( .A(x[1461]), .B(y[1461]), .Z(n5176) );
  ANDN U4441 ( .B(y[1460]), .A(x[1460]), .Z(n9435) );
  ANDN U4442 ( .B(n5176), .A(n9435), .Z(n13359) );
  ANDN U4443 ( .B(x[1460]), .A(y[1460]), .Z(n9438) );
  NANDN U4444 ( .A(y[1459]), .B(x[1459]), .Z(n5179) );
  NANDN U4445 ( .A(n9438), .B(n5179), .Z(n13357) );
  NANDN U4446 ( .A(x[1458]), .B(y[1458]), .Z(n9433) );
  ANDN U4447 ( .B(y[1459]), .A(x[1459]), .Z(n13355) );
  ANDN U4448 ( .B(x[1457]), .A(y[1457]), .Z(n9430) );
  ANDN U4449 ( .B(y[1456]), .A(x[1456]), .Z(n5180) );
  NANDN U4450 ( .A(y[1456]), .B(x[1456]), .Z(n9431) );
  NANDN U4451 ( .A(x[1455]), .B(y[1455]), .Z(n5181) );
  ANDN U4452 ( .B(y[1454]), .A(x[1454]), .Z(n5184) );
  ANDN U4453 ( .B(x[1453]), .A(y[1453]), .Z(n5187) );
  NANDN U4454 ( .A(x[1453]), .B(y[1453]), .Z(n5185) );
  NANDN U4455 ( .A(y[1452]), .B(x[1452]), .Z(n5186) );
  ANDN U4456 ( .B(x[1451]), .A(y[1451]), .Z(n5191) );
  IV U4457 ( .A(n5191), .Z(n3344) );
  ANDN U4458 ( .B(y[1450]), .A(x[1450]), .Z(n13335) );
  NANDN U4459 ( .A(y[1450]), .B(x[1450]), .Z(n5190) );
  NANDN U4460 ( .A(x[1448]), .B(y[1448]), .Z(n9429) );
  NANDN U4461 ( .A(x[1449]), .B(y[1449]), .Z(n5192) );
  NAND U4462 ( .A(n9429), .B(n5192), .Z(n13331) );
  NANDN U4463 ( .A(y[1448]), .B(x[1448]), .Z(n13329) );
  NANDN U4464 ( .A(x[1446]), .B(y[1446]), .Z(n13322) );
  IV U4465 ( .A(n13322), .Z(n5193) );
  NANDN U4466 ( .A(x[1447]), .B(y[1447]), .Z(n13327) );
  NANDN U4467 ( .A(y[1445]), .B(x[1445]), .Z(n5195) );
  NANDN U4468 ( .A(x[1445]), .B(y[1445]), .Z(n13321) );
  NANDN U4469 ( .A(x[1442]), .B(y[1442]), .Z(n9423) );
  NANDN U4470 ( .A(x[1443]), .B(y[1443]), .Z(n9424) );
  NAND U4471 ( .A(n9423), .B(n9424), .Z(n13313) );
  NANDN U4472 ( .A(y[1442]), .B(x[1442]), .Z(n13311) );
  NANDN U4473 ( .A(y[1441]), .B(x[1441]), .Z(n3347) );
  NANDN U4474 ( .A(x[1441]), .B(y[1441]), .Z(n9419) );
  NANDN U4475 ( .A(x[1440]), .B(y[1440]), .Z(n9420) );
  NAND U4476 ( .A(n9419), .B(n9420), .Z(n3345) );
  NAND U4477 ( .A(n3347), .B(n3345), .Z(n13308) );
  NANDN U4478 ( .A(y[1440]), .B(x[1440]), .Z(n3346) );
  AND U4479 ( .A(n3347), .B(n3346), .Z(n9422) );
  NANDN U4480 ( .A(y[1439]), .B(x[1439]), .Z(n3348) );
  NAND U4481 ( .A(n9422), .B(n3348), .Z(n13306) );
  IV U4482 ( .A(n13306), .Z(n9418) );
  NANDN U4483 ( .A(x[1438]), .B(y[1438]), .Z(n9417) );
  NANDN U4484 ( .A(x[1439]), .B(y[1439]), .Z(n9421) );
  AND U4485 ( .A(n9417), .B(n9421), .Z(n13305) );
  ANDN U4486 ( .B(x[1438]), .A(y[1438]), .Z(n13303) );
  NANDN U4487 ( .A(y[1435]), .B(x[1435]), .Z(n13295) );
  NANDN U4488 ( .A(x[1435]), .B(y[1435]), .Z(n3350) );
  NANDN U4489 ( .A(x[1434]), .B(y[1434]), .Z(n3349) );
  NAND U4490 ( .A(n3350), .B(n3349), .Z(n13293) );
  NANDN U4491 ( .A(y[1434]), .B(x[1434]), .Z(n3352) );
  NANDN U4492 ( .A(y[1433]), .B(x[1433]), .Z(n3351) );
  AND U4493 ( .A(n3352), .B(n3351), .Z(n5200) );
  NANDN U4494 ( .A(x[1432]), .B(y[1432]), .Z(n3353) );
  ANDN U4495 ( .B(y[1433]), .A(x[1433]), .Z(n5198) );
  ANDN U4496 ( .B(n3353), .A(n5198), .Z(n13288) );
  NANDN U4497 ( .A(y[1429]), .B(x[1429]), .Z(n5203) );
  NANDN U4498 ( .A(y[1430]), .B(x[1430]), .Z(n9414) );
  NAND U4499 ( .A(n5203), .B(n9414), .Z(n13283) );
  NANDN U4500 ( .A(x[1428]), .B(y[1428]), .Z(n5205) );
  NANDN U4501 ( .A(x[1429]), .B(y[1429]), .Z(n5201) );
  NAND U4502 ( .A(n5205), .B(n5201), .Z(n13281) );
  NANDN U4503 ( .A(y[1427]), .B(x[1427]), .Z(n9413) );
  NANDN U4504 ( .A(y[1428]), .B(x[1428]), .Z(n5204) );
  AND U4505 ( .A(n9413), .B(n5204), .Z(n13279) );
  NANDN U4506 ( .A(x[1426]), .B(y[1426]), .Z(n5207) );
  NANDN U4507 ( .A(x[1427]), .B(y[1427]), .Z(n5206) );
  NAND U4508 ( .A(n5207), .B(n5206), .Z(n13277) );
  NANDN U4509 ( .A(y[1425]), .B(x[1425]), .Z(n5209) );
  NANDN U4510 ( .A(y[1426]), .B(x[1426]), .Z(n13274) );
  ANDN U4511 ( .B(y[1424]), .A(x[1424]), .Z(n5211) );
  NANDN U4512 ( .A(y[1424]), .B(x[1424]), .Z(n5208) );
  NANDN U4513 ( .A(y[1423]), .B(x[1423]), .Z(n5213) );
  ANDN U4514 ( .B(y[1422]), .A(x[1422]), .Z(n5216) );
  NANDN U4515 ( .A(y[1422]), .B(x[1422]), .Z(n5212) );
  NANDN U4516 ( .A(x[1421]), .B(y[1421]), .Z(n3355) );
  NANDN U4517 ( .A(x[1420]), .B(y[1420]), .Z(n3354) );
  NAND U4518 ( .A(n3355), .B(n3354), .Z(n5214) );
  NANDN U4519 ( .A(y[1420]), .B(x[1420]), .Z(n3357) );
  NANDN U4520 ( .A(y[1419]), .B(x[1419]), .Z(n3356) );
  AND U4521 ( .A(n3357), .B(n3356), .Z(n9404) );
  NANDN U4522 ( .A(x[1418]), .B(y[1418]), .Z(n3358) );
  ANDN U4523 ( .B(y[1419]), .A(x[1419]), .Z(n9408) );
  ANDN U4524 ( .B(n3358), .A(n9408), .Z(n4511) );
  NANDN U4525 ( .A(x[1417]), .B(y[1417]), .Z(n3359) );
  AND U4526 ( .A(n4511), .B(n3359), .Z(n9402) );
  NANDN U4527 ( .A(x[1416]), .B(y[1416]), .Z(n3360) );
  AND U4528 ( .A(n9402), .B(n3360), .Z(n13260) );
  ANDN U4529 ( .B(x[1416]), .A(y[1416]), .Z(n9400) );
  NANDN U4530 ( .A(y[1415]), .B(x[1415]), .Z(n13259) );
  NANDN U4531 ( .A(y[1414]), .B(x[1414]), .Z(n13255) );
  NANDN U4532 ( .A(y[1413]), .B(x[1413]), .Z(n9396) );
  ANDN U4533 ( .B(y[1413]), .A(x[1413]), .Z(n13253) );
  NANDN U4534 ( .A(y[1412]), .B(x[1412]), .Z(n9397) );
  NANDN U4535 ( .A(x[1410]), .B(y[1410]), .Z(n5220) );
  NANDN U4536 ( .A(x[1411]), .B(y[1411]), .Z(n5219) );
  NAND U4537 ( .A(n5220), .B(n5219), .Z(n13245) );
  ANDN U4538 ( .B(x[1410]), .A(y[1410]), .Z(n13243) );
  NANDN U4539 ( .A(x[1408]), .B(y[1408]), .Z(n13236) );
  NANDN U4540 ( .A(x[1405]), .B(y[1405]), .Z(n13229) );
  NANDN U4541 ( .A(y[1404]), .B(x[1404]), .Z(n3362) );
  NANDN U4542 ( .A(y[1405]), .B(x[1405]), .Z(n3361) );
  NAND U4543 ( .A(n3362), .B(n3361), .Z(n13227) );
  NANDN U4544 ( .A(x[1403]), .B(y[1403]), .Z(n3364) );
  NANDN U4545 ( .A(x[1404]), .B(y[1404]), .Z(n3363) );
  AND U4546 ( .A(n3364), .B(n3363), .Z(n13225) );
  NANDN U4547 ( .A(y[1403]), .B(x[1403]), .Z(n3366) );
  NANDN U4548 ( .A(y[1402]), .B(x[1402]), .Z(n3365) );
  NAND U4549 ( .A(n3366), .B(n3365), .Z(n13223) );
  NANDN U4550 ( .A(x[1402]), .B(y[1402]), .Z(n9389) );
  NANDN U4551 ( .A(y[1401]), .B(x[1401]), .Z(n5223) );
  NANDN U4552 ( .A(x[1401]), .B(y[1401]), .Z(n9388) );
  ANDN U4553 ( .B(x[1399]), .A(y[1399]), .Z(n13214) );
  IV U4554 ( .A(n13214), .Z(n9386) );
  NANDN U4555 ( .A(x[1398]), .B(y[1398]), .Z(n9384) );
  NANDN U4556 ( .A(x[1399]), .B(y[1399]), .Z(n5225) );
  AND U4557 ( .A(n9384), .B(n5225), .Z(n13213) );
  XNOR U4558 ( .A(y[1398]), .B(x[1398]), .Z(n3367) );
  ANDN U4559 ( .B(x[1397]), .A(y[1397]), .Z(n9381) );
  ANDN U4560 ( .B(n3367), .A(n9381), .Z(n13211) );
  NANDN U4561 ( .A(x[1396]), .B(y[1396]), .Z(n9379) );
  NANDN U4562 ( .A(x[1397]), .B(y[1397]), .Z(n9383) );
  AND U4563 ( .A(n9379), .B(n9383), .Z(n13209) );
  NANDN U4564 ( .A(x[1394]), .B(y[1394]), .Z(n9376) );
  NANDN U4565 ( .A(x[1395]), .B(y[1395]), .Z(n13204) );
  IV U4566 ( .A(n13204), .Z(n9380) );
  ANDN U4567 ( .B(x[1393]), .A(y[1393]), .Z(n5226) );
  ANDN U4568 ( .B(y[1392]), .A(x[1392]), .Z(n13197) );
  NANDN U4569 ( .A(y[1392]), .B(x[1392]), .Z(n5227) );
  ANDN U4570 ( .B(y[1390]), .A(x[1390]), .Z(n9374) );
  ANDN U4571 ( .B(y[1391]), .A(x[1391]), .Z(n9375) );
  OR U4572 ( .A(n9374), .B(n9375), .Z(n13193) );
  NANDN U4573 ( .A(y[1389]), .B(x[1389]), .Z(n5228) );
  NANDN U4574 ( .A(y[1390]), .B(x[1390]), .Z(n13191) );
  ANDN U4575 ( .B(y[1389]), .A(x[1389]), .Z(n13189) );
  NANDN U4576 ( .A(y[1388]), .B(x[1388]), .Z(n5229) );
  ANDN U4577 ( .B(y[1386]), .A(x[1386]), .Z(n13180) );
  IV U4578 ( .A(n13180), .Z(n9372) );
  ANDN U4579 ( .B(y[1384]), .A(x[1384]), .Z(n9369) );
  ANDN U4580 ( .B(y[1385]), .A(x[1385]), .Z(n9371) );
  NOR U4581 ( .A(n9369), .B(n9371), .Z(n13177) );
  NANDN U4582 ( .A(y[1384]), .B(x[1384]), .Z(n13174) );
  IV U4583 ( .A(n13174), .Z(n5234) );
  ANDN U4584 ( .B(y[1383]), .A(x[1383]), .Z(n13172) );
  IV U4585 ( .A(n13172), .Z(n9370) );
  NANDN U4586 ( .A(y[1383]), .B(x[1383]), .Z(n3369) );
  NANDN U4587 ( .A(y[1382]), .B(x[1382]), .Z(n3368) );
  AND U4588 ( .A(n3369), .B(n3368), .Z(n13171) );
  IV U4589 ( .A(n13171), .Z(n9368) );
  NANDN U4590 ( .A(y[1381]), .B(x[1381]), .Z(n5236) );
  NANDN U4591 ( .A(x[1380]), .B(y[1380]), .Z(n5237) );
  NANDN U4592 ( .A(y[1379]), .B(x[1379]), .Z(n5239) );
  NANDN U4593 ( .A(x[1379]), .B(y[1379]), .Z(n5238) );
  ANDN U4594 ( .B(x[1377]), .A(y[1377]), .Z(n13159) );
  NANDN U4595 ( .A(x[1376]), .B(y[1376]), .Z(n3371) );
  NANDN U4596 ( .A(x[1377]), .B(y[1377]), .Z(n3370) );
  AND U4597 ( .A(n3371), .B(n3370), .Z(n13157) );
  NANDN U4598 ( .A(y[1376]), .B(x[1376]), .Z(n3373) );
  NANDN U4599 ( .A(y[1375]), .B(x[1375]), .Z(n3372) );
  AND U4600 ( .A(n3373), .B(n3372), .Z(n5244) );
  NANDN U4601 ( .A(x[1375]), .B(y[1375]), .Z(n5241) );
  NANDN U4602 ( .A(x[1374]), .B(y[1374]), .Z(n3374) );
  NAND U4603 ( .A(n5241), .B(n3374), .Z(n13153) );
  IV U4604 ( .A(n13153), .Z(n4504) );
  NANDN U4605 ( .A(y[1373]), .B(x[1373]), .Z(n13151) );
  IV U4606 ( .A(n13151), .Z(n5245) );
  NANDN U4607 ( .A(x[1372]), .B(y[1372]), .Z(n9364) );
  NANDN U4608 ( .A(x[1373]), .B(y[1373]), .Z(n9367) );
  NAND U4609 ( .A(n9364), .B(n9367), .Z(n13149) );
  NANDN U4610 ( .A(y[1371]), .B(x[1371]), .Z(n9363) );
  NANDN U4611 ( .A(y[1372]), .B(x[1372]), .Z(n13146) );
  ANDN U4612 ( .B(y[1371]), .A(x[1371]), .Z(n13144) );
  NANDN U4613 ( .A(y[1370]), .B(x[1370]), .Z(n9362) );
  ANDN U4614 ( .B(y[1368]), .A(x[1368]), .Z(n13137) );
  NANDN U4615 ( .A(y[1367]), .B(x[1367]), .Z(n13135) );
  NANDN U4616 ( .A(y[1368]), .B(x[1368]), .Z(n5249) );
  NANDN U4617 ( .A(x[1366]), .B(y[1366]), .Z(n9359) );
  NANDN U4618 ( .A(x[1367]), .B(y[1367]), .Z(n9361) );
  NAND U4619 ( .A(n9359), .B(n9361), .Z(n13133) );
  ANDN U4620 ( .B(x[1365]), .A(y[1365]), .Z(n9356) );
  ANDN U4621 ( .B(x[1366]), .A(y[1366]), .Z(n9360) );
  NOR U4622 ( .A(n9356), .B(n9360), .Z(n13131) );
  NANDN U4623 ( .A(x[1364]), .B(y[1364]), .Z(n9354) );
  NANDN U4624 ( .A(x[1365]), .B(y[1365]), .Z(n9358) );
  AND U4625 ( .A(n9354), .B(n9358), .Z(n13128) );
  NANDN U4626 ( .A(x[1362]), .B(y[1362]), .Z(n5251) );
  NANDN U4627 ( .A(x[1363]), .B(y[1363]), .Z(n13125) );
  IV U4628 ( .A(n13125), .Z(n9355) );
  ANDN U4629 ( .B(x[1361]), .A(y[1361]), .Z(n9350) );
  ANDN U4630 ( .B(y[1360]), .A(x[1360]), .Z(n9348) );
  NANDN U4631 ( .A(y[1360]), .B(x[1360]), .Z(n9351) );
  NANDN U4632 ( .A(x[1358]), .B(y[1358]), .Z(n13113) );
  NANDN U4633 ( .A(y[1358]), .B(x[1358]), .Z(n13110) );
  IV U4634 ( .A(n13110), .Z(n5252) );
  ANDN U4635 ( .B(y[1356]), .A(x[1356]), .Z(n13105) );
  NANDN U4636 ( .A(x[1357]), .B(y[1357]), .Z(n13109) );
  NANDN U4637 ( .A(n13105), .B(n13109), .Z(n3375) );
  NANDN U4638 ( .A(y[1357]), .B(x[1357]), .Z(n3376) );
  NAND U4639 ( .A(n3375), .B(n3376), .Z(n4501) );
  NANDN U4640 ( .A(y[1356]), .B(x[1356]), .Z(n3377) );
  AND U4641 ( .A(n3377), .B(n3376), .Z(n13107) );
  IV U4642 ( .A(n13107), .Z(n9347) );
  NANDN U4643 ( .A(y[1355]), .B(x[1355]), .Z(n3380) );
  ANDN U4644 ( .B(y[1355]), .A(x[1355]), .Z(n9346) );
  NANDN U4645 ( .A(x[1354]), .B(y[1354]), .Z(n5253) );
  NANDN U4646 ( .A(n9346), .B(n5253), .Z(n3378) );
  AND U4647 ( .A(n3380), .B(n3378), .Z(n13102) );
  NANDN U4648 ( .A(y[1354]), .B(x[1354]), .Z(n3379) );
  AND U4649 ( .A(n3380), .B(n3379), .Z(n13101) );
  NANDN U4650 ( .A(y[1353]), .B(x[1353]), .Z(n3382) );
  NANDN U4651 ( .A(y[1352]), .B(x[1352]), .Z(n3381) );
  AND U4652 ( .A(n3382), .B(n3381), .Z(n13097) );
  NANDN U4653 ( .A(x[1351]), .B(y[1351]), .Z(n3384) );
  NANDN U4654 ( .A(x[1352]), .B(y[1352]), .Z(n3383) );
  NAND U4655 ( .A(n3384), .B(n3383), .Z(n13095) );
  NANDN U4656 ( .A(y[1351]), .B(x[1351]), .Z(n5255) );
  NANDN U4657 ( .A(x[1350]), .B(y[1350]), .Z(n5257) );
  NANDN U4658 ( .A(y[1349]), .B(x[1349]), .Z(n5258) );
  ANDN U4659 ( .B(y[1348]), .A(x[1348]), .Z(n5261) );
  NANDN U4660 ( .A(y[1347]), .B(x[1347]), .Z(n5263) );
  ANDN U4661 ( .B(y[1346]), .A(x[1346]), .Z(n13083) );
  NANDN U4662 ( .A(y[1346]), .B(x[1346]), .Z(n5262) );
  NANDN U4663 ( .A(x[1344]), .B(y[1344]), .Z(n9337) );
  NANDN U4664 ( .A(x[1345]), .B(y[1345]), .Z(n5264) );
  NAND U4665 ( .A(n9337), .B(n5264), .Z(n13078) );
  NANDN U4666 ( .A(y[1343]), .B(x[1343]), .Z(n5265) );
  NANDN U4667 ( .A(y[1344]), .B(x[1344]), .Z(n13077) );
  ANDN U4668 ( .B(y[1343]), .A(x[1343]), .Z(n13075) );
  NANDN U4669 ( .A(y[1342]), .B(x[1342]), .Z(n5266) );
  ANDN U4670 ( .B(y[1340]), .A(x[1340]), .Z(n13066) );
  NANDN U4671 ( .A(y[1339]), .B(x[1339]), .Z(n13065) );
  IV U4672 ( .A(n13065), .Z(n4498) );
  NANDN U4673 ( .A(y[1340]), .B(x[1340]), .Z(n5270) );
  NANDN U4674 ( .A(x[1338]), .B(y[1338]), .Z(n3386) );
  NANDN U4675 ( .A(x[1339]), .B(y[1339]), .Z(n3385) );
  NAND U4676 ( .A(n3386), .B(n3385), .Z(n13062) );
  NANDN U4677 ( .A(y[1338]), .B(x[1338]), .Z(n3388) );
  NANDN U4678 ( .A(y[1337]), .B(x[1337]), .Z(n3387) );
  AND U4679 ( .A(n3388), .B(n3387), .Z(n13061) );
  NANDN U4680 ( .A(x[1336]), .B(y[1336]), .Z(n3390) );
  NANDN U4681 ( .A(x[1337]), .B(y[1337]), .Z(n3389) );
  NAND U4682 ( .A(n3390), .B(n3389), .Z(n13058) );
  NANDN U4683 ( .A(y[1336]), .B(x[1336]), .Z(n3392) );
  NANDN U4684 ( .A(y[1335]), .B(x[1335]), .Z(n3391) );
  AND U4685 ( .A(n3392), .B(n3391), .Z(n13057) );
  NANDN U4686 ( .A(x[1334]), .B(y[1334]), .Z(n3394) );
  NANDN U4687 ( .A(x[1335]), .B(y[1335]), .Z(n3393) );
  NAND U4688 ( .A(n3394), .B(n3393), .Z(n13054) );
  NANDN U4689 ( .A(y[1334]), .B(x[1334]), .Z(n9326) );
  NANDN U4690 ( .A(y[1333]), .B(x[1333]), .Z(n3395) );
  AND U4691 ( .A(n9326), .B(n3395), .Z(n13053) );
  ANDN U4692 ( .B(y[1332]), .A(x[1332]), .Z(n9318) );
  NANDN U4693 ( .A(x[1333]), .B(y[1333]), .Z(n9324) );
  NANDN U4694 ( .A(n9318), .B(n9324), .Z(n13050) );
  NANDN U4695 ( .A(y[1331]), .B(x[1331]), .Z(n9317) );
  NANDN U4696 ( .A(y[1332]), .B(x[1332]), .Z(n9320) );
  NAND U4697 ( .A(n9317), .B(n9320), .Z(n13048) );
  ANDN U4698 ( .B(y[1330]), .A(x[1330]), .Z(n9314) );
  ANDN U4699 ( .B(y[1331]), .A(x[1331]), .Z(n9319) );
  NOR U4700 ( .A(n9314), .B(n9319), .Z(n13047) );
  ANDN U4701 ( .B(y[1328]), .A(x[1328]), .Z(n9311) );
  ANDN U4702 ( .B(y[1329]), .A(x[1329]), .Z(n9315) );
  NOR U4703 ( .A(n9311), .B(n9315), .Z(n13043) );
  ANDN U4704 ( .B(y[1327]), .A(x[1327]), .Z(n13038) );
  NANDN U4705 ( .A(x[1326]), .B(y[1326]), .Z(n13034) );
  NANDN U4706 ( .A(y[1325]), .B(x[1325]), .Z(n13033) );
  IV U4707 ( .A(n13033), .Z(n5273) );
  NANDN U4708 ( .A(x[1324]), .B(y[1324]), .Z(n9309) );
  NANDN U4709 ( .A(x[1325]), .B(y[1325]), .Z(n9310) );
  NAND U4710 ( .A(n9309), .B(n9310), .Z(n13031) );
  NANDN U4711 ( .A(y[1323]), .B(x[1323]), .Z(n5275) );
  NANDN U4712 ( .A(x[1323]), .B(y[1323]), .Z(n13027) );
  NANDN U4713 ( .A(y[1321]), .B(x[1321]), .Z(n5278) );
  NANDN U4714 ( .A(x[1321]), .B(y[1321]), .Z(n5276) );
  ANDN U4715 ( .B(x[1319]), .A(y[1319]), .Z(n5283) );
  NANDN U4716 ( .A(x[1319]), .B(y[1319]), .Z(n5280) );
  NANDN U4717 ( .A(y[1317]), .B(x[1317]), .Z(n13012) );
  NANDN U4718 ( .A(x[1316]), .B(y[1316]), .Z(n9307) );
  NANDN U4719 ( .A(x[1317]), .B(y[1317]), .Z(n5284) );
  AND U4720 ( .A(n9307), .B(n5284), .Z(n13013) );
  NANDN U4721 ( .A(y[1315]), .B(x[1315]), .Z(n5287) );
  NANDN U4722 ( .A(x[1314]), .B(y[1314]), .Z(n5289) );
  ANDN U4723 ( .B(x[1313]), .A(y[1313]), .Z(n5290) );
  NANDN U4724 ( .A(x[1310]), .B(y[1310]), .Z(n9304) );
  NANDN U4725 ( .A(x[1311]), .B(y[1311]), .Z(n9306) );
  NAND U4726 ( .A(n9304), .B(n9306), .Z(n12995) );
  NANDN U4727 ( .A(y[1309]), .B(x[1309]), .Z(n5292) );
  NANDN U4728 ( .A(x[1308]), .B(y[1308]), .Z(n12986) );
  NANDN U4729 ( .A(x[1307]), .B(y[1307]), .Z(n3397) );
  NANDN U4730 ( .A(x[1306]), .B(y[1306]), .Z(n3396) );
  AND U4731 ( .A(n3397), .B(n3396), .Z(n12983) );
  NANDN U4732 ( .A(y[1306]), .B(x[1306]), .Z(n3399) );
  NANDN U4733 ( .A(y[1305]), .B(x[1305]), .Z(n3398) );
  AND U4734 ( .A(n3399), .B(n3398), .Z(n9301) );
  ANDN U4735 ( .B(y[1305]), .A(x[1305]), .Z(n9299) );
  NANDN U4736 ( .A(x[1304]), .B(y[1304]), .Z(n3400) );
  NANDN U4737 ( .A(n9299), .B(n3400), .Z(n12979) );
  ANDN U4738 ( .B(x[1303]), .A(y[1303]), .Z(n12977) );
  XNOR U4739 ( .A(x[1304]), .B(y[1304]), .Z(n5294) );
  NANDN U4740 ( .A(x[1302]), .B(y[1302]), .Z(n3401) );
  NANDN U4741 ( .A(x[1303]), .B(y[1303]), .Z(n9297) );
  NAND U4742 ( .A(n3401), .B(n9297), .Z(n12975) );
  XNOR U4743 ( .A(x[1302]), .B(y[1302]), .Z(n9295) );
  ANDN U4744 ( .B(x[1301]), .A(y[1301]), .Z(n9294) );
  ANDN U4745 ( .B(n9295), .A(n9294), .Z(n12973) );
  NANDN U4746 ( .A(x[1300]), .B(y[1300]), .Z(n9291) );
  NANDN U4747 ( .A(x[1301]), .B(y[1301]), .Z(n9296) );
  NAND U4748 ( .A(n9291), .B(n9296), .Z(n12971) );
  NANDN U4749 ( .A(x[1299]), .B(y[1299]), .Z(n12966) );
  NANDN U4750 ( .A(y[1299]), .B(x[1299]), .Z(n3403) );
  NANDN U4751 ( .A(y[1298]), .B(x[1298]), .Z(n3402) );
  AND U4752 ( .A(n3403), .B(n3402), .Z(n5300) );
  NANDN U4753 ( .A(y[1297]), .B(x[1297]), .Z(n5296) );
  ANDN U4754 ( .B(y[1298]), .A(x[1298]), .Z(n3404) );
  NANDN U4755 ( .A(x[1297]), .B(y[1297]), .Z(n3405) );
  ANDN U4756 ( .B(n3405), .A(n3404), .Z(n5298) );
  NANDN U4757 ( .A(x[1296]), .B(y[1296]), .Z(n3406) );
  AND U4758 ( .A(n5298), .B(n3406), .Z(n12963) );
  NANDN U4759 ( .A(y[1295]), .B(x[1295]), .Z(n12960) );
  NANDN U4760 ( .A(x[1294]), .B(y[1294]), .Z(n9287) );
  NANDN U4761 ( .A(x[1295]), .B(y[1295]), .Z(n9290) );
  NAND U4762 ( .A(n9287), .B(n9290), .Z(n12958) );
  ANDN U4763 ( .B(x[1293]), .A(y[1293]), .Z(n9285) );
  ANDN U4764 ( .B(x[1294]), .A(y[1294]), .Z(n9289) );
  NOR U4765 ( .A(n9285), .B(n9289), .Z(n12957) );
  NANDN U4766 ( .A(x[1292]), .B(y[1292]), .Z(n9284) );
  NANDN U4767 ( .A(x[1293]), .B(y[1293]), .Z(n9288) );
  NAND U4768 ( .A(n9284), .B(n9288), .Z(n12955) );
  NANDN U4769 ( .A(y[1291]), .B(x[1291]), .Z(n5302) );
  ANDN U4770 ( .B(x[1292]), .A(y[1292]), .Z(n9286) );
  ANDN U4771 ( .B(n5302), .A(n9286), .Z(n12953) );
  ANDN U4772 ( .B(y[1290]), .A(x[1290]), .Z(n9281) );
  NANDN U4773 ( .A(x[1291]), .B(y[1291]), .Z(n9283) );
  NANDN U4774 ( .A(n9281), .B(n9283), .Z(n12951) );
  ANDN U4775 ( .B(x[1285]), .A(y[1285]), .Z(n5303) );
  NANDN U4776 ( .A(x[1284]), .B(y[1284]), .Z(n5305) );
  NANDN U4777 ( .A(y[1284]), .B(x[1284]), .Z(n5304) );
  ANDN U4778 ( .B(x[1283]), .A(y[1283]), .Z(n5307) );
  ANDN U4779 ( .B(y[1282]), .A(x[1282]), .Z(n5309) );
  NANDN U4780 ( .A(y[1282]), .B(x[1282]), .Z(n5308) );
  NANDN U4781 ( .A(x[1280]), .B(y[1280]), .Z(n5314) );
  NANDN U4782 ( .A(y[1279]), .B(x[1279]), .Z(n5315) );
  ANDN U4783 ( .B(y[1278]), .A(x[1278]), .Z(n12926) );
  NANDN U4784 ( .A(y[1277]), .B(x[1277]), .Z(n12925) );
  XNOR U4785 ( .A(x[1278]), .B(y[1278]), .Z(n9275) );
  NANDN U4786 ( .A(x[1276]), .B(y[1276]), .Z(n9273) );
  NANDN U4787 ( .A(x[1277]), .B(y[1277]), .Z(n9276) );
  NAND U4788 ( .A(n9273), .B(n9276), .Z(n12923) );
  ANDN U4789 ( .B(x[1275]), .A(y[1275]), .Z(n9272) );
  ANDN U4790 ( .B(x[1276]), .A(y[1276]), .Z(n9274) );
  NOR U4791 ( .A(n9272), .B(n9274), .Z(n12921) );
  NANDN U4792 ( .A(x[1273]), .B(y[1273]), .Z(n3407) );
  ANDN U4793 ( .B(y[1274]), .A(x[1274]), .Z(n4478) );
  ANDN U4794 ( .B(n3407), .A(n4478), .Z(n5320) );
  NANDN U4795 ( .A(x[1272]), .B(y[1272]), .Z(n3408) );
  AND U4796 ( .A(n5320), .B(n3408), .Z(n12915) );
  ANDN U4797 ( .B(x[1271]), .A(y[1271]), .Z(n12913) );
  NANDN U4798 ( .A(x[1270]), .B(y[1270]), .Z(n3410) );
  NANDN U4799 ( .A(x[1271]), .B(y[1271]), .Z(n3409) );
  AND U4800 ( .A(n3410), .B(n3409), .Z(n12910) );
  NANDN U4801 ( .A(y[1269]), .B(x[1269]), .Z(n3411) );
  XOR U4802 ( .A(x[1270]), .B(y[1270]), .Z(n9269) );
  ANDN U4803 ( .B(n3411), .A(n9269), .Z(n9267) );
  IV U4804 ( .A(n9267), .Z(n12908) );
  NANDN U4805 ( .A(x[1268]), .B(y[1268]), .Z(n5323) );
  NANDN U4806 ( .A(x[1269]), .B(y[1269]), .Z(n9270) );
  NAND U4807 ( .A(n5323), .B(n9270), .Z(n12907) );
  ANDN U4808 ( .B(y[1266]), .A(x[1266]), .Z(n5324) );
  NANDN U4809 ( .A(x[1267]), .B(y[1267]), .Z(n12903) );
  ANDN U4810 ( .B(x[1266]), .A(y[1266]), .Z(n12901) );
  NANDN U4811 ( .A(x[1265]), .B(y[1265]), .Z(n5325) );
  NANDN U4812 ( .A(y[1264]), .B(x[1264]), .Z(n5326) );
  ANDN U4813 ( .B(x[1263]), .A(y[1263]), .Z(n5331) );
  ANDN U4814 ( .B(y[1262]), .A(x[1262]), .Z(n12891) );
  NANDN U4815 ( .A(y[1262]), .B(x[1262]), .Z(n5330) );
  NANDN U4816 ( .A(x[1260]), .B(y[1260]), .Z(n5332) );
  NANDN U4817 ( .A(x[1261]), .B(y[1261]), .Z(n9265) );
  NAND U4818 ( .A(n5332), .B(n9265), .Z(n12886) );
  NANDN U4819 ( .A(y[1260]), .B(x[1260]), .Z(n12885) );
  ANDN U4820 ( .B(y[1258]), .A(x[1258]), .Z(n12879) );
  NANDN U4821 ( .A(y[1257]), .B(x[1257]), .Z(n12876) );
  NANDN U4822 ( .A(y[1258]), .B(x[1258]), .Z(n5334) );
  NANDN U4823 ( .A(x[1256]), .B(y[1256]), .Z(n9263) );
  NANDN U4824 ( .A(x[1257]), .B(y[1257]), .Z(n5335) );
  NAND U4825 ( .A(n9263), .B(n5335), .Z(n12874) );
  IV U4826 ( .A(n12874), .Z(n4475) );
  NANDN U4827 ( .A(y[1254]), .B(x[1254]), .Z(n9261) );
  NANDN U4828 ( .A(y[1253]), .B(x[1253]), .Z(n5339) );
  ANDN U4829 ( .B(y[1252]), .A(x[1252]), .Z(n12863) );
  NANDN U4830 ( .A(y[1252]), .B(x[1252]), .Z(n5338) );
  NANDN U4831 ( .A(x[1250]), .B(y[1250]), .Z(n9258) );
  NANDN U4832 ( .A(x[1251]), .B(y[1251]), .Z(n9260) );
  NAND U4833 ( .A(n9258), .B(n9260), .Z(n12859) );
  ANDN U4834 ( .B(x[1250]), .A(y[1250]), .Z(n12857) );
  NANDN U4835 ( .A(x[1248]), .B(y[1248]), .Z(n12851) );
  ANDN U4836 ( .B(x[1247]), .A(y[1247]), .Z(n12849) );
  NANDN U4837 ( .A(y[1248]), .B(x[1248]), .Z(n5341) );
  NANDN U4838 ( .A(x[1246]), .B(y[1246]), .Z(n9256) );
  NANDN U4839 ( .A(x[1247]), .B(y[1247]), .Z(n9257) );
  NAND U4840 ( .A(n9256), .B(n9257), .Z(n12847) );
  NANDN U4841 ( .A(x[1245]), .B(y[1245]), .Z(n12842) );
  NANDN U4842 ( .A(y[1244]), .B(x[1244]), .Z(n5342) );
  NANDN U4843 ( .A(x[1242]), .B(y[1242]), .Z(n9252) );
  NANDN U4844 ( .A(x[1243]), .B(y[1243]), .Z(n9255) );
  NAND U4845 ( .A(n9252), .B(n9255), .Z(n12835) );
  NANDN U4846 ( .A(y[1242]), .B(x[1242]), .Z(n12832) );
  NANDN U4847 ( .A(x[1240]), .B(y[1240]), .Z(n12826) );
  NANDN U4848 ( .A(x[1241]), .B(y[1241]), .Z(n12831) );
  ANDN U4849 ( .B(x[1239]), .A(y[1239]), .Z(n12825) );
  NANDN U4850 ( .A(x[1238]), .B(y[1238]), .Z(n9250) );
  NANDN U4851 ( .A(x[1239]), .B(y[1239]), .Z(n9251) );
  NAND U4852 ( .A(n9250), .B(n9251), .Z(n12823) );
  XNOR U4853 ( .A(y[1238]), .B(x[1238]), .Z(n3412) );
  ANDN U4854 ( .B(x[1237]), .A(y[1237]), .Z(n9247) );
  ANDN U4855 ( .B(n3412), .A(n9247), .Z(n12821) );
  IV U4856 ( .A(n12821), .Z(n4472) );
  ANDN U4857 ( .B(y[1235]), .A(x[1235]), .Z(n12814) );
  NANDN U4858 ( .A(y[1234]), .B(x[1234]), .Z(n12813) );
  NANDN U4859 ( .A(x[1233]), .B(y[1233]), .Z(n3414) );
  NANDN U4860 ( .A(x[1234]), .B(y[1234]), .Z(n3413) );
  NAND U4861 ( .A(n3414), .B(n3413), .Z(n12811) );
  NANDN U4862 ( .A(y[1232]), .B(x[1232]), .Z(n3416) );
  NANDN U4863 ( .A(y[1233]), .B(x[1233]), .Z(n3415) );
  AND U4864 ( .A(n3416), .B(n3415), .Z(n12809) );
  NANDN U4865 ( .A(x[1229]), .B(y[1229]), .Z(n3417) );
  ANDN U4866 ( .B(y[1230]), .A(x[1230]), .Z(n4468) );
  ANDN U4867 ( .B(n3417), .A(n4468), .Z(n9241) );
  NANDN U4868 ( .A(x[1228]), .B(y[1228]), .Z(n3418) );
  AND U4869 ( .A(n9241), .B(n3418), .Z(n12803) );
  NANDN U4870 ( .A(y[1227]), .B(x[1227]), .Z(n12801) );
  NANDN U4871 ( .A(x[1226]), .B(y[1226]), .Z(n9236) );
  NANDN U4872 ( .A(x[1227]), .B(y[1227]), .Z(n9237) );
  NAND U4873 ( .A(n9236), .B(n9237), .Z(n12799) );
  ANDN U4874 ( .B(x[1226]), .A(y[1226]), .Z(n12797) );
  NANDN U4875 ( .A(x[1224]), .B(y[1224]), .Z(n12791) );
  NANDN U4876 ( .A(x[1222]), .B(y[1222]), .Z(n9232) );
  NANDN U4877 ( .A(x[1223]), .B(y[1223]), .Z(n9235) );
  NAND U4878 ( .A(n9232), .B(n9235), .Z(n12787) );
  NANDN U4879 ( .A(y[1220]), .B(x[1220]), .Z(n3420) );
  NANDN U4880 ( .A(y[1221]), .B(x[1221]), .Z(n3419) );
  NAND U4881 ( .A(n3420), .B(n3419), .Z(n9230) );
  NANDN U4882 ( .A(x[1221]), .B(y[1221]), .Z(n9233) );
  NAND U4883 ( .A(n9230), .B(n9233), .Z(n3421) );
  ANDN U4884 ( .B(x[1222]), .A(y[1222]), .Z(n9234) );
  ANDN U4885 ( .B(n3421), .A(n9234), .Z(n12785) );
  NANDN U4886 ( .A(x[1219]), .B(y[1219]), .Z(n3423) );
  NANDN U4887 ( .A(x[1220]), .B(y[1220]), .Z(n3422) );
  AND U4888 ( .A(n3423), .B(n3422), .Z(n9229) );
  NANDN U4889 ( .A(x[1218]), .B(y[1218]), .Z(n9228) );
  NANDN U4890 ( .A(y[1219]), .B(x[1219]), .Z(n4464) );
  NANDN U4891 ( .A(n9228), .B(n4464), .Z(n3424) );
  AND U4892 ( .A(n3424), .B(n9233), .Z(n3425) );
  NAND U4893 ( .A(n9229), .B(n3425), .Z(n12783) );
  NANDN U4894 ( .A(y[1217]), .B(x[1217]), .Z(n5348) );
  NANDN U4895 ( .A(x[1216]), .B(y[1216]), .Z(n12775) );
  NANDN U4896 ( .A(x[1215]), .B(y[1215]), .Z(n3427) );
  NANDN U4897 ( .A(x[1214]), .B(y[1214]), .Z(n3426) );
  AND U4898 ( .A(n3427), .B(n3426), .Z(n12770) );
  ANDN U4899 ( .B(x[1214]), .A(y[1214]), .Z(n12768) );
  NANDN U4900 ( .A(y[1213]), .B(x[1213]), .Z(n9225) );
  ANDN U4901 ( .B(y[1212]), .A(x[1212]), .Z(n9222) );
  NANDN U4902 ( .A(y[1212]), .B(x[1212]), .Z(n9226) );
  NANDN U4903 ( .A(x[1211]), .B(y[1211]), .Z(n9223) );
  ANDN U4904 ( .B(y[1210]), .A(x[1210]), .Z(n9220) );
  ANDN U4905 ( .B(x[1209]), .A(y[1209]), .Z(n5352) );
  NANDN U4906 ( .A(x[1209]), .B(y[1209]), .Z(n9221) );
  ANDN U4907 ( .B(x[1207]), .A(y[1207]), .Z(n12753) );
  ANDN U4908 ( .B(y[1206]), .A(x[1206]), .Z(n9216) );
  ANDN U4909 ( .B(y[1207]), .A(x[1207]), .Z(n9219) );
  NOR U4910 ( .A(n9216), .B(n9219), .Z(n12751) );
  IV U4911 ( .A(n12751), .Z(n4461) );
  NANDN U4912 ( .A(y[1205]), .B(x[1205]), .Z(n9214) );
  NANDN U4913 ( .A(y[1206]), .B(x[1206]), .Z(n9218) );
  NAND U4914 ( .A(n9214), .B(n9218), .Z(n12749) );
  ANDN U4915 ( .B(y[1204]), .A(x[1204]), .Z(n9213) );
  ANDN U4916 ( .B(y[1205]), .A(x[1205]), .Z(n9217) );
  NOR U4917 ( .A(n9213), .B(n9217), .Z(n12746) );
  NANDN U4918 ( .A(x[1202]), .B(y[1202]), .Z(n5354) );
  NANDN U4919 ( .A(x[1203]), .B(y[1203]), .Z(n12743) );
  NANDN U4920 ( .A(y[1202]), .B(x[1202]), .Z(n12740) );
  NANDN U4921 ( .A(x[1201]), .B(y[1201]), .Z(n5355) );
  NANDN U4922 ( .A(x[1200]), .B(y[1200]), .Z(n5359) );
  ANDN U4923 ( .B(x[1199]), .A(y[1199]), .Z(n12732) );
  NANDN U4924 ( .A(x[1199]), .B(y[1199]), .Z(n5358) );
  ANDN U4925 ( .B(x[1197]), .A(y[1197]), .Z(n5361) );
  IV U4926 ( .A(n5361), .Z(n4458) );
  NANDN U4927 ( .A(x[1196]), .B(y[1196]), .Z(n12722) );
  NANDN U4928 ( .A(x[1197]), .B(y[1197]), .Z(n12727) );
  IV U4929 ( .A(n12727), .Z(n9209) );
  NANDN U4930 ( .A(y[1196]), .B(x[1196]), .Z(n5362) );
  NANDN U4931 ( .A(y[1195]), .B(x[1195]), .Z(n4456) );
  NANDN U4932 ( .A(x[1194]), .B(y[1194]), .Z(n9208) );
  NANDN U4933 ( .A(x[1195]), .B(y[1195]), .Z(n5363) );
  NAND U4934 ( .A(n9208), .B(n5363), .Z(n3428) );
  AND U4935 ( .A(n4456), .B(n3428), .Z(n12721) );
  ANDN U4936 ( .B(x[1193]), .A(y[1193]), .Z(n5365) );
  NANDN U4937 ( .A(x[1193]), .B(y[1193]), .Z(n5367) );
  NANDN U4938 ( .A(x[1192]), .B(y[1192]), .Z(n3429) );
  AND U4939 ( .A(n5367), .B(n3429), .Z(n5369) );
  ANDN U4940 ( .B(x[1191]), .A(y[1191]), .Z(n5370) );
  NANDN U4941 ( .A(x[1191]), .B(y[1191]), .Z(n5368) );
  NANDN U4942 ( .A(y[1190]), .B(x[1190]), .Z(n5371) );
  ANDN U4943 ( .B(x[1189]), .A(y[1189]), .Z(n9206) );
  ANDN U4944 ( .B(y[1188]), .A(x[1188]), .Z(n5374) );
  NANDN U4945 ( .A(y[1188]), .B(x[1188]), .Z(n9207) );
  ANDN U4946 ( .B(y[1186]), .A(x[1186]), .Z(n12703) );
  NANDN U4947 ( .A(x[1184]), .B(y[1184]), .Z(n9203) );
  NANDN U4948 ( .A(x[1185]), .B(y[1185]), .Z(n9205) );
  NAND U4949 ( .A(n9203), .B(n9205), .Z(n12698) );
  ANDN U4950 ( .B(x[1184]), .A(y[1184]), .Z(n12697) );
  NANDN U4951 ( .A(x[1182]), .B(y[1182]), .Z(n5379) );
  ANDN U4952 ( .B(x[1181]), .A(y[1181]), .Z(n5381) );
  NANDN U4953 ( .A(x[1180]), .B(y[1180]), .Z(n12686) );
  NANDN U4954 ( .A(x[1178]), .B(y[1178]), .Z(n9199) );
  NANDN U4955 ( .A(x[1179]), .B(y[1179]), .Z(n9200) );
  NAND U4956 ( .A(n9199), .B(n9200), .Z(n12683) );
  NANDN U4957 ( .A(y[1177]), .B(x[1177]), .Z(n5383) );
  NANDN U4958 ( .A(x[1176]), .B(y[1176]), .Z(n12674) );
  IV U4959 ( .A(n12674), .Z(n9197) );
  NANDN U4960 ( .A(x[1177]), .B(y[1177]), .Z(n12679) );
  NANDN U4961 ( .A(y[1175]), .B(x[1175]), .Z(n12673) );
  NANDN U4962 ( .A(x[1174]), .B(y[1174]), .Z(n5386) );
  NANDN U4963 ( .A(x[1175]), .B(y[1175]), .Z(n9198) );
  NAND U4964 ( .A(n5386), .B(n9198), .Z(n12671) );
  NANDN U4965 ( .A(y[1173]), .B(x[1173]), .Z(n9194) );
  NANDN U4966 ( .A(y[1174]), .B(x[1174]), .Z(n5385) );
  AND U4967 ( .A(n9194), .B(n5385), .Z(n12669) );
  ANDN U4968 ( .B(y[1172]), .A(x[1172]), .Z(n9193) );
  NANDN U4969 ( .A(x[1173]), .B(y[1173]), .Z(n5387) );
  NANDN U4970 ( .A(n9193), .B(n5387), .Z(n12667) );
  NANDN U4971 ( .A(y[1171]), .B(x[1171]), .Z(n5388) );
  ANDN U4972 ( .B(x[1172]), .A(y[1172]), .Z(n9195) );
  ANDN U4973 ( .B(n5388), .A(n9195), .Z(n12665) );
  NANDN U4974 ( .A(x[1170]), .B(y[1170]), .Z(n9190) );
  ANDN U4975 ( .B(y[1171]), .A(x[1171]), .Z(n9192) );
  ANDN U4976 ( .B(n9190), .A(n9192), .Z(n12663) );
  NANDN U4977 ( .A(y[1170]), .B(x[1170]), .Z(n5389) );
  ANDN U4978 ( .B(x[1169]), .A(y[1169]), .Z(n9189) );
  ANDN U4979 ( .B(n5389), .A(n9189), .Z(n12661) );
  NANDN U4980 ( .A(x[1168]), .B(y[1168]), .Z(n9188) );
  ANDN U4981 ( .B(y[1169]), .A(x[1169]), .Z(n9191) );
  ANDN U4982 ( .B(n9188), .A(n9191), .Z(n12659) );
  NANDN U4983 ( .A(y[1168]), .B(x[1168]), .Z(n12657) );
  IV U4984 ( .A(n12657), .Z(n4452) );
  NANDN U4985 ( .A(x[1166]), .B(y[1166]), .Z(n12650) );
  IV U4986 ( .A(n12650), .Z(n5392) );
  NANDN U4987 ( .A(x[1167]), .B(y[1167]), .Z(n12655) );
  NANDN U4988 ( .A(y[1165]), .B(x[1165]), .Z(n12649) );
  NANDN U4989 ( .A(x[1164]), .B(y[1164]), .Z(n5394) );
  NANDN U4990 ( .A(x[1165]), .B(y[1165]), .Z(n5393) );
  NAND U4991 ( .A(n5394), .B(n5393), .Z(n12647) );
  NANDN U4992 ( .A(y[1164]), .B(x[1164]), .Z(n12645) );
  NANDN U4993 ( .A(y[1163]), .B(x[1163]), .Z(n9184) );
  ANDN U4994 ( .B(y[1163]), .A(x[1163]), .Z(n12642) );
  NANDN U4995 ( .A(y[1162]), .B(x[1162]), .Z(n9185) );
  ANDN U4996 ( .B(y[1160]), .A(x[1160]), .Z(n12635) );
  NANDN U4997 ( .A(x[1158]), .B(y[1158]), .Z(n9180) );
  NANDN U4998 ( .A(x[1159]), .B(y[1159]), .Z(n9181) );
  NAND U4999 ( .A(n9180), .B(n9181), .Z(n12630) );
  IV U5000 ( .A(n12630), .Z(n4449) );
  NANDN U5001 ( .A(y[1156]), .B(x[1156]), .Z(n5398) );
  NANDN U5002 ( .A(y[1155]), .B(x[1155]), .Z(n5401) );
  ANDN U5003 ( .B(y[1154]), .A(x[1154]), .Z(n12619) );
  NANDN U5004 ( .A(x[1155]), .B(y[1155]), .Z(n5400) );
  ANDN U5005 ( .B(x[1153]), .A(y[1153]), .Z(n12617) );
  NANDN U5006 ( .A(x[1153]), .B(y[1153]), .Z(n5403) );
  ANDN U5007 ( .B(y[1152]), .A(x[1152]), .Z(n9176) );
  ANDN U5008 ( .B(n5403), .A(n9176), .Z(n12615) );
  NANDN U5009 ( .A(y[1151]), .B(x[1151]), .Z(n9175) );
  NANDN U5010 ( .A(y[1152]), .B(x[1152]), .Z(n9179) );
  NAND U5011 ( .A(n9175), .B(n9179), .Z(n12613) );
  NANDN U5012 ( .A(x[1150]), .B(y[1150]), .Z(n5405) );
  ANDN U5013 ( .B(y[1151]), .A(x[1151]), .Z(n12610) );
  ANDN U5014 ( .B(x[1149]), .A(y[1149]), .Z(n5406) );
  ANDN U5015 ( .B(y[1148]), .A(x[1148]), .Z(n12603) );
  IV U5016 ( .A(n12603), .Z(n9173) );
  ANDN U5017 ( .B(x[1145]), .A(y[1145]), .Z(n9169) );
  ANDN U5018 ( .B(x[1146]), .A(y[1146]), .Z(n9171) );
  OR U5019 ( .A(n9169), .B(n9171), .Z(n10190) );
  ANDN U5020 ( .B(y[1145]), .A(x[1145]), .Z(n10189) );
  NANDN U5021 ( .A(x[1144]), .B(y[1144]), .Z(n9167) );
  NANDN U5022 ( .A(n10189), .B(n9167), .Z(n12595) );
  ANDN U5023 ( .B(x[1144]), .A(y[1144]), .Z(n10188) );
  ANDN U5024 ( .B(y[1142]), .A(x[1142]), .Z(n9163) );
  NANDN U5025 ( .A(x[1143]), .B(y[1143]), .Z(n9168) );
  NANDN U5026 ( .A(n9163), .B(n9168), .Z(n12591) );
  NANDN U5027 ( .A(y[1141]), .B(x[1141]), .Z(n9162) );
  NANDN U5028 ( .A(y[1142]), .B(x[1142]), .Z(n9166) );
  AND U5029 ( .A(n9162), .B(n9166), .Z(n12589) );
  ANDN U5030 ( .B(y[1140]), .A(x[1140]), .Z(n9160) );
  ANDN U5031 ( .B(y[1141]), .A(x[1141]), .Z(n9165) );
  NOR U5032 ( .A(n9160), .B(n9165), .Z(n12587) );
  NANDN U5033 ( .A(y[1139]), .B(x[1139]), .Z(n9159) );
  NANDN U5034 ( .A(y[1140]), .B(x[1140]), .Z(n9161) );
  NAND U5035 ( .A(n9159), .B(n9161), .Z(n12585) );
  NANDN U5036 ( .A(x[1139]), .B(y[1139]), .Z(n12582) );
  ANDN U5037 ( .B(x[1137]), .A(y[1137]), .Z(n5408) );
  ANDN U5038 ( .B(y[1135]), .A(x[1135]), .Z(n9156) );
  NANDN U5039 ( .A(x[1134]), .B(y[1134]), .Z(n9155) );
  NANDN U5040 ( .A(n9156), .B(n9155), .Z(n12571) );
  ANDN U5041 ( .B(x[1134]), .A(y[1134]), .Z(n12569) );
  ANDN U5042 ( .B(y[1132]), .A(x[1132]), .Z(n9151) );
  NANDN U5043 ( .A(y[1131]), .B(x[1131]), .Z(n5410) );
  NANDN U5044 ( .A(x[1130]), .B(y[1130]), .Z(n12558) );
  NANDN U5045 ( .A(y[1130]), .B(x[1130]), .Z(n5411) );
  ANDN U5046 ( .B(y[1128]), .A(x[1128]), .Z(n9148) );
  NANDN U5047 ( .A(x[1129]), .B(y[1129]), .Z(n9149) );
  NANDN U5048 ( .A(n9148), .B(n9149), .Z(n12555) );
  NANDN U5049 ( .A(y[1127]), .B(x[1127]), .Z(n5412) );
  ANDN U5050 ( .B(y[1126]), .A(x[1126]), .Z(n5415) );
  NANDN U5051 ( .A(y[1125]), .B(x[1125]), .Z(n5416) );
  NANDN U5052 ( .A(x[1124]), .B(y[1124]), .Z(n12542) );
  NANDN U5053 ( .A(y[1124]), .B(x[1124]), .Z(n5417) );
  ANDN U5054 ( .B(y[1123]), .A(x[1123]), .Z(n9147) );
  NANDN U5055 ( .A(x[1122]), .B(y[1122]), .Z(n9146) );
  NANDN U5056 ( .A(n9147), .B(n9146), .Z(n12539) );
  NANDN U5057 ( .A(x[1120]), .B(y[1120]), .Z(n12530) );
  NANDN U5058 ( .A(x[1121]), .B(y[1121]), .Z(n12535) );
  IV U5059 ( .A(n12535), .Z(n9145) );
  ANDN U5060 ( .B(x[1119]), .A(y[1119]), .Z(n12528) );
  IV U5061 ( .A(n12528), .Z(n4443) );
  NANDN U5062 ( .A(x[1118]), .B(y[1118]), .Z(n9142) );
  NANDN U5063 ( .A(x[1119]), .B(y[1119]), .Z(n9143) );
  AND U5064 ( .A(n9142), .B(n9143), .Z(n12527) );
  ANDN U5065 ( .B(x[1117]), .A(y[1117]), .Z(n5421) );
  NANDN U5066 ( .A(x[1116]), .B(y[1116]), .Z(n12518) );
  IV U5067 ( .A(n12518), .Z(n9140) );
  NANDN U5068 ( .A(x[1117]), .B(y[1117]), .Z(n12522) );
  ANDN U5069 ( .B(x[1113]), .A(y[1113]), .Z(n5425) );
  NANDN U5070 ( .A(x[1112]), .B(y[1112]), .Z(n12506) );
  NANDN U5071 ( .A(x[1113]), .B(y[1113]), .Z(n12511) );
  NANDN U5072 ( .A(y[1112]), .B(x[1112]), .Z(n5426) );
  XNOR U5073 ( .A(y[1110]), .B(x[1110]), .Z(n3430) );
  ANDN U5074 ( .B(x[1109]), .A(y[1109]), .Z(n9131) );
  ANDN U5075 ( .B(n3430), .A(n9131), .Z(n12501) );
  NANDN U5076 ( .A(x[1108]), .B(y[1108]), .Z(n9129) );
  NANDN U5077 ( .A(x[1109]), .B(y[1109]), .Z(n9133) );
  NAND U5078 ( .A(n9129), .B(n9133), .Z(n12499) );
  ANDN U5079 ( .B(x[1107]), .A(y[1107]), .Z(n9128) );
  ANDN U5080 ( .B(x[1108]), .A(y[1108]), .Z(n9132) );
  NOR U5081 ( .A(n9128), .B(n9132), .Z(n12497) );
  NANDN U5082 ( .A(x[1106]), .B(y[1106]), .Z(n9127) );
  NANDN U5083 ( .A(x[1107]), .B(y[1107]), .Z(n9130) );
  NAND U5084 ( .A(n9127), .B(n9130), .Z(n12495) );
  NANDN U5085 ( .A(y[1106]), .B(x[1106]), .Z(n12493) );
  NANDN U5086 ( .A(x[1104]), .B(y[1104]), .Z(n12486) );
  IV U5087 ( .A(n12486), .Z(n9125) );
  NANDN U5088 ( .A(x[1105]), .B(y[1105]), .Z(n12491) );
  NANDN U5089 ( .A(y[1103]), .B(x[1103]), .Z(n12485) );
  NANDN U5090 ( .A(x[1102]), .B(y[1102]), .Z(n5430) );
  NANDN U5091 ( .A(x[1103]), .B(y[1103]), .Z(n9126) );
  NAND U5092 ( .A(n5430), .B(n9126), .Z(n12483) );
  NANDN U5093 ( .A(y[1101]), .B(x[1101]), .Z(n9121) );
  NANDN U5094 ( .A(x[1100]), .B(y[1100]), .Z(n12474) );
  IV U5095 ( .A(n12474), .Z(n5431) );
  NANDN U5096 ( .A(x[1101]), .B(y[1101]), .Z(n12479) );
  NANDN U5097 ( .A(n5431), .B(n12479), .Z(n4440) );
  NANDN U5098 ( .A(y[1099]), .B(x[1099]), .Z(n12473) );
  NANDN U5099 ( .A(x[1098]), .B(y[1098]), .Z(n5433) );
  NANDN U5100 ( .A(x[1099]), .B(y[1099]), .Z(n5432) );
  NAND U5101 ( .A(n5433), .B(n5432), .Z(n12471) );
  NANDN U5102 ( .A(y[1097]), .B(x[1097]), .Z(n9119) );
  NANDN U5103 ( .A(x[1096]), .B(y[1096]), .Z(n12462) );
  IV U5104 ( .A(n12462), .Z(n5434) );
  NANDN U5105 ( .A(x[1097]), .B(y[1097]), .Z(n12467) );
  NANDN U5106 ( .A(y[1095]), .B(x[1095]), .Z(n12461) );
  NANDN U5107 ( .A(x[1094]), .B(y[1094]), .Z(n5436) );
  NANDN U5108 ( .A(x[1095]), .B(y[1095]), .Z(n5435) );
  NAND U5109 ( .A(n5436), .B(n5435), .Z(n12459) );
  NANDN U5110 ( .A(y[1093]), .B(x[1093]), .Z(n5437) );
  NANDN U5111 ( .A(x[1092]), .B(y[1092]), .Z(n12450) );
  ANDN U5112 ( .B(x[1089]), .A(y[1089]), .Z(n9114) );
  ANDN U5113 ( .B(x[1090]), .A(y[1090]), .Z(n9116) );
  NOR U5114 ( .A(n9114), .B(n9116), .Z(n12445) );
  NANDN U5115 ( .A(x[1088]), .B(y[1088]), .Z(n12438) );
  IV U5116 ( .A(n12438), .Z(n9113) );
  NANDN U5117 ( .A(x[1089]), .B(y[1089]), .Z(n12443) );
  NANDN U5118 ( .A(n9113), .B(n12443), .Z(n4438) );
  ANDN U5119 ( .B(y[1087]), .A(x[1087]), .Z(n12436) );
  NANDN U5120 ( .A(y[1086]), .B(x[1086]), .Z(n9111) );
  NANDN U5121 ( .A(x[1084]), .B(y[1084]), .Z(n12428) );
  NANDN U5122 ( .A(y[1083]), .B(x[1083]), .Z(n12427) );
  NANDN U5123 ( .A(y[1082]), .B(x[1082]), .Z(n12422) );
  NANDN U5124 ( .A(y[1081]), .B(x[1081]), .Z(n9104) );
  NANDN U5125 ( .A(x[1080]), .B(y[1080]), .Z(n12416) );
  IV U5126 ( .A(n12416), .Z(n9103) );
  NANDN U5127 ( .A(x[1081]), .B(y[1081]), .Z(n12421) );
  NANDN U5128 ( .A(y[1080]), .B(x[1080]), .Z(n9105) );
  ANDN U5129 ( .B(x[1079]), .A(y[1079]), .Z(n12414) );
  NANDN U5130 ( .A(x[1079]), .B(y[1079]), .Z(n3432) );
  NANDN U5131 ( .A(x[1078]), .B(y[1078]), .Z(n3431) );
  NAND U5132 ( .A(n3432), .B(n3431), .Z(n12413) );
  NANDN U5133 ( .A(y[1078]), .B(x[1078]), .Z(n3434) );
  NANDN U5134 ( .A(y[1077]), .B(x[1077]), .Z(n3433) );
  AND U5135 ( .A(n3434), .B(n3433), .Z(n9100) );
  NANDN U5136 ( .A(x[1076]), .B(y[1076]), .Z(n3435) );
  ANDN U5137 ( .B(y[1077]), .A(x[1077]), .Z(n9101) );
  ANDN U5138 ( .B(n3435), .A(n9101), .Z(n4435) );
  NANDN U5139 ( .A(y[1076]), .B(x[1076]), .Z(n9102) );
  NANDN U5140 ( .A(y[1075]), .B(x[1075]), .Z(n9098) );
  NAND U5141 ( .A(n9102), .B(n9098), .Z(n3436) );
  NAND U5142 ( .A(n4435), .B(n3436), .Z(n3437) );
  AND U5143 ( .A(n9100), .B(n3437), .Z(n12411) );
  NANDN U5144 ( .A(x[1074]), .B(y[1074]), .Z(n5444) );
  NANDN U5145 ( .A(y[1073]), .B(x[1073]), .Z(n5447) );
  ANDN U5146 ( .B(y[1072]), .A(x[1072]), .Z(n5449) );
  NANDN U5147 ( .A(y[1071]), .B(x[1071]), .Z(n5451) );
  ANDN U5148 ( .B(y[1070]), .A(x[1070]), .Z(n12396) );
  NANDN U5149 ( .A(y[1070]), .B(x[1070]), .Z(n5450) );
  NANDN U5150 ( .A(x[1068]), .B(y[1068]), .Z(n5454) );
  NANDN U5151 ( .A(x[1069]), .B(y[1069]), .Z(n5452) );
  NAND U5152 ( .A(n5454), .B(n5452), .Z(n12393) );
  NANDN U5153 ( .A(y[1067]), .B(x[1067]), .Z(n5455) );
  NANDN U5154 ( .A(y[1068]), .B(x[1068]), .Z(n12390) );
  IV U5155 ( .A(n12390), .Z(n3438) );
  ANDN U5156 ( .B(y[1067]), .A(x[1067]), .Z(n12388) );
  NANDN U5157 ( .A(y[1066]), .B(x[1066]), .Z(n5456) );
  NANDN U5158 ( .A(x[1065]), .B(y[1065]), .Z(n3440) );
  NANDN U5159 ( .A(x[1064]), .B(y[1064]), .Z(n3439) );
  NAND U5160 ( .A(n3440), .B(n3439), .Z(n5457) );
  NANDN U5161 ( .A(y[1063]), .B(x[1063]), .Z(n3442) );
  NANDN U5162 ( .A(y[1064]), .B(x[1064]), .Z(n3441) );
  AND U5163 ( .A(n3442), .B(n3441), .Z(n5465) );
  NANDN U5164 ( .A(x[1063]), .B(y[1063]), .Z(n5460) );
  NANDN U5165 ( .A(x[1062]), .B(y[1062]), .Z(n3443) );
  AND U5166 ( .A(n5460), .B(n3443), .Z(n4432) );
  NANDN U5167 ( .A(x[1061]), .B(y[1061]), .Z(n3444) );
  AND U5168 ( .A(n4432), .B(n3444), .Z(n12381) );
  NANDN U5169 ( .A(x[1060]), .B(y[1060]), .Z(n3446) );
  NANDN U5170 ( .A(x[1059]), .B(y[1059]), .Z(n3445) );
  AND U5171 ( .A(n3446), .B(n3445), .Z(n9089) );
  NANDN U5172 ( .A(x[1058]), .B(y[1058]), .Z(n9085) );
  ANDN U5173 ( .B(x[1059]), .A(y[1059]), .Z(n4429) );
  ANDN U5174 ( .B(x[1057]), .A(y[1057]), .Z(n5469) );
  NANDN U5175 ( .A(x[1057]), .B(y[1057]), .Z(n12373) );
  ANDN U5176 ( .B(x[1055]), .A(y[1055]), .Z(n5473) );
  NANDN U5177 ( .A(x[1055]), .B(y[1055]), .Z(n5470) );
  NANDN U5178 ( .A(y[1054]), .B(x[1054]), .Z(n5472) );
  NANDN U5179 ( .A(y[1053]), .B(x[1053]), .Z(n5476) );
  ANDN U5180 ( .B(y[1052]), .A(x[1052]), .Z(n12361) );
  NANDN U5181 ( .A(y[1052]), .B(x[1052]), .Z(n5477) );
  NANDN U5182 ( .A(x[1050]), .B(y[1050]), .Z(n9072) );
  NANDN U5183 ( .A(x[1051]), .B(y[1051]), .Z(n5478) );
  NAND U5184 ( .A(n9072), .B(n5478), .Z(n12356) );
  NANDN U5185 ( .A(y[1050]), .B(x[1050]), .Z(n12355) );
  NANDN U5186 ( .A(x[1049]), .B(y[1049]), .Z(n12352) );
  NANDN U5187 ( .A(x[1047]), .B(y[1047]), .Z(n5481) );
  ANDN U5188 ( .B(y[1046]), .A(x[1046]), .Z(n9063) );
  ANDN U5189 ( .B(n5481), .A(n9063), .Z(n12345) );
  NANDN U5190 ( .A(y[1045]), .B(x[1045]), .Z(n9059) );
  NANDN U5191 ( .A(y[1046]), .B(x[1046]), .Z(n9067) );
  NAND U5192 ( .A(n9059), .B(n9067), .Z(n12343) );
  ANDN U5193 ( .B(y[1044]), .A(x[1044]), .Z(n9054) );
  ANDN U5194 ( .B(y[1045]), .A(x[1045]), .Z(n9065) );
  NOR U5195 ( .A(n9054), .B(n9065), .Z(n12341) );
  NANDN U5196 ( .A(y[1043]), .B(x[1043]), .Z(n9051) );
  NANDN U5197 ( .A(y[1044]), .B(x[1044]), .Z(n9058) );
  AND U5198 ( .A(n9051), .B(n9058), .Z(n12339) );
  ANDN U5199 ( .B(y[1040]), .A(x[1040]), .Z(n9041) );
  ANDN U5200 ( .B(y[1041]), .A(x[1041]), .Z(n9049) );
  NOR U5201 ( .A(n9041), .B(n9049), .Z(n12333) );
  NANDN U5202 ( .A(y[1038]), .B(x[1038]), .Z(n5483) );
  NANDN U5203 ( .A(y[1037]), .B(x[1037]), .Z(n5487) );
  AND U5204 ( .A(n5483), .B(n5487), .Z(n4427) );
  ANDN U5205 ( .B(y[1036]), .A(x[1036]), .Z(n5488) );
  NANDN U5206 ( .A(y[1036]), .B(x[1036]), .Z(n5486) );
  NANDN U5207 ( .A(x[1034]), .B(y[1034]), .Z(n12316) );
  NANDN U5208 ( .A(y[1033]), .B(x[1033]), .Z(n12315) );
  NANDN U5209 ( .A(x[1032]), .B(y[1032]), .Z(n9037) );
  NANDN U5210 ( .A(x[1033]), .B(y[1033]), .Z(n9038) );
  NAND U5211 ( .A(n9037), .B(n9038), .Z(n12313) );
  NANDN U5212 ( .A(y[1031]), .B(x[1031]), .Z(n5492) );
  NANDN U5213 ( .A(y[1030]), .B(x[1030]), .Z(n5493) );
  NANDN U5214 ( .A(y[1029]), .B(x[1029]), .Z(n5497) );
  NANDN U5215 ( .A(x[1028]), .B(y[1028]), .Z(n5499) );
  NANDN U5216 ( .A(y[1028]), .B(x[1028]), .Z(n5496) );
  NANDN U5217 ( .A(x[1026]), .B(y[1026]), .Z(n12296) );
  NANDN U5218 ( .A(y[1025]), .B(x[1025]), .Z(n12295) );
  NANDN U5219 ( .A(x[1024]), .B(y[1024]), .Z(n9035) );
  NANDN U5220 ( .A(x[1025]), .B(y[1025]), .Z(n5502) );
  NAND U5221 ( .A(n9035), .B(n5502), .Z(n12293) );
  ANDN U5222 ( .B(x[1023]), .A(y[1023]), .Z(n9034) );
  ANDN U5223 ( .B(y[1022]), .A(x[1022]), .Z(n12284) );
  NANDN U5224 ( .A(y[1021]), .B(x[1021]), .Z(n12283) );
  ANDN U5225 ( .B(y[1020]), .A(x[1020]), .Z(n9029) );
  ANDN U5226 ( .B(y[1021]), .A(x[1021]), .Z(n9032) );
  NOR U5227 ( .A(n9029), .B(n9032), .Z(n12281) );
  NANDN U5228 ( .A(y[1019]), .B(x[1019]), .Z(n9027) );
  NANDN U5229 ( .A(y[1020]), .B(x[1020]), .Z(n9031) );
  NAND U5230 ( .A(n9027), .B(n9031), .Z(n12279) );
  ANDN U5231 ( .B(y[1019]), .A(x[1019]), .Z(n9030) );
  ANDN U5232 ( .B(y[1018]), .A(x[1018]), .Z(n9025) );
  ANDN U5233 ( .B(x[1017]), .A(y[1017]), .Z(n3447) );
  NANDN U5234 ( .A(y[1018]), .B(x[1018]), .Z(n9028) );
  ANDN U5235 ( .B(y[1017]), .A(x[1017]), .Z(n9026) );
  NANDN U5236 ( .A(x[1016]), .B(y[1016]), .Z(n9021) );
  NANDN U5237 ( .A(y[1016]), .B(x[1016]), .Z(n3448) );
  ANDN U5238 ( .B(n3448), .A(n3447), .Z(n9023) );
  ANDN U5239 ( .B(x[1015]), .A(y[1015]), .Z(n9019) );
  ANDN U5240 ( .B(n9028), .A(n9019), .Z(n3449) );
  NAND U5241 ( .A(n9023), .B(n3449), .Z(n12275) );
  NANDN U5242 ( .A(x[1014]), .B(y[1014]), .Z(n9018) );
  ANDN U5243 ( .B(y[1015]), .A(x[1015]), .Z(n9022) );
  ANDN U5244 ( .B(n9018), .A(n9022), .Z(n12273) );
  ANDN U5245 ( .B(x[1012]), .A(y[1012]), .Z(n12267) );
  IV U5246 ( .A(n12267), .Z(n9016) );
  NANDN U5247 ( .A(x[1010]), .B(y[1010]), .Z(n9009) );
  ANDN U5248 ( .B(x[1009]), .A(y[1009]), .Z(n5504) );
  NANDN U5249 ( .A(x[1008]), .B(y[1008]), .Z(n12257) );
  NANDN U5250 ( .A(x[1006]), .B(y[1006]), .Z(n9004) );
  NANDN U5251 ( .A(x[1007]), .B(y[1007]), .Z(n9008) );
  NAND U5252 ( .A(n9004), .B(n9008), .Z(n12252) );
  ANDN U5253 ( .B(x[1005]), .A(y[1005]), .Z(n5506) );
  ANDN U5254 ( .B(x[1006]), .A(y[1006]), .Z(n9007) );
  NOR U5255 ( .A(n5506), .B(n9007), .Z(n12251) );
  IV U5256 ( .A(n12251), .Z(n4422) );
  NANDN U5257 ( .A(x[1005]), .B(y[1005]), .Z(n9003) );
  ANDN U5258 ( .B(y[1004]), .A(x[1004]), .Z(n9001) );
  ANDN U5259 ( .B(n9003), .A(n9001), .Z(n12249) );
  NANDN U5260 ( .A(y[1003]), .B(x[1003]), .Z(n9000) );
  ANDN U5261 ( .B(x[1004]), .A(y[1004]), .Z(n5505) );
  ANDN U5262 ( .B(n9000), .A(n5505), .Z(n12247) );
  ANDN U5263 ( .B(y[1002]), .A(x[1002]), .Z(n8997) );
  ANDN U5264 ( .B(y[1003]), .A(x[1003]), .Z(n9002) );
  NOR U5265 ( .A(n8997), .B(n9002), .Z(n12244) );
  NANDN U5266 ( .A(y[999]), .B(x[999]), .Z(n5508) );
  NANDN U5267 ( .A(x[998]), .B(y[998]), .Z(n5510) );
  NANDN U5268 ( .A(x[999]), .B(y[999]), .Z(n12237) );
  NANDN U5269 ( .A(y[997]), .B(x[997]), .Z(n8994) );
  NANDN U5270 ( .A(x[992]), .B(y[992]), .Z(n12216) );
  NANDN U5271 ( .A(x[993]), .B(y[993]), .Z(n12221) );
  NANDN U5272 ( .A(x[990]), .B(y[990]), .Z(n8988) );
  NANDN U5273 ( .A(x[991]), .B(y[991]), .Z(n8989) );
  NAND U5274 ( .A(n8988), .B(n8989), .Z(n12212) );
  NANDN U5275 ( .A(y[989]), .B(x[989]), .Z(n5517) );
  NANDN U5276 ( .A(x[989]), .B(y[989]), .Z(n12209) );
  ANDN U5277 ( .B(y[988]), .A(x[988]), .Z(n5518) );
  ANDN U5278 ( .B(x[987]), .A(y[987]), .Z(n8986) );
  NANDN U5279 ( .A(x[987]), .B(y[987]), .Z(n5519) );
  ANDN U5280 ( .B(x[985]), .A(y[985]), .Z(n5520) );
  ANDN U5281 ( .B(x[983]), .A(y[983]), .Z(n12195) );
  IV U5282 ( .A(n12195), .Z(n8981) );
  NANDN U5283 ( .A(x[982]), .B(y[982]), .Z(n8978) );
  NANDN U5284 ( .A(x[983]), .B(y[983]), .Z(n8982) );
  AND U5285 ( .A(n8978), .B(n8982), .Z(n12193) );
  NANDN U5286 ( .A(y[979]), .B(x[979]), .Z(n8971) );
  ANDN U5287 ( .B(x[980]), .A(y[980]), .Z(n8976) );
  ANDN U5288 ( .B(n8971), .A(n8976), .Z(n12187) );
  NANDN U5289 ( .A(x[979]), .B(y[979]), .Z(n12185) );
  IV U5290 ( .A(n12185), .Z(n8973) );
  NANDN U5291 ( .A(x[976]), .B(y[976]), .Z(n12177) );
  NANDN U5292 ( .A(x[978]), .B(y[978]), .Z(n4416) );
  NANDN U5293 ( .A(x[977]), .B(y[977]), .Z(n3450) );
  AND U5294 ( .A(n4416), .B(n3450), .Z(n12181) );
  IV U5295 ( .A(n12181), .Z(n8970) );
  ANDN U5296 ( .B(x[976]), .A(y[976]), .Z(n5522) );
  NANDN U5297 ( .A(x[975]), .B(y[975]), .Z(n8969) );
  ANDN U5298 ( .B(y[974]), .A(x[974]), .Z(n8968) );
  ANDN U5299 ( .B(n8969), .A(n8968), .Z(n12173) );
  ANDN U5300 ( .B(x[973]), .A(y[973]), .Z(n3451) );
  ANDN U5301 ( .B(y[972]), .A(x[972]), .Z(n8964) );
  ANDN U5302 ( .B(y[973]), .A(x[973]), .Z(n8967) );
  NANDN U5303 ( .A(y[972]), .B(x[972]), .Z(n3452) );
  ANDN U5304 ( .B(n3452), .A(n3451), .Z(n8966) );
  NANDN U5305 ( .A(y[971]), .B(x[971]), .Z(n8962) );
  NAND U5306 ( .A(n8966), .B(n8962), .Z(n12167) );
  NANDN U5307 ( .A(x[970]), .B(y[970]), .Z(n8957) );
  ANDN U5308 ( .B(y[971]), .A(x[971]), .Z(n8965) );
  ANDN U5309 ( .B(n8957), .A(n8965), .Z(n12165) );
  NANDN U5310 ( .A(y[969]), .B(x[969]), .Z(n5525) );
  NANDN U5311 ( .A(y[970]), .B(x[970]), .Z(n8963) );
  NAND U5312 ( .A(n5525), .B(n8963), .Z(n12163) );
  NANDN U5313 ( .A(x[969]), .B(y[969]), .Z(n8958) );
  ANDN U5314 ( .B(y[968]), .A(x[968]), .Z(n8952) );
  ANDN U5315 ( .B(n8958), .A(n8952), .Z(n12161) );
  NANDN U5316 ( .A(y[967]), .B(x[967]), .Z(n8948) );
  NANDN U5317 ( .A(y[968]), .B(x[968]), .Z(n5524) );
  AND U5318 ( .A(n8948), .B(n5524), .Z(n12159) );
  ANDN U5319 ( .B(y[966]), .A(x[966]), .Z(n8943) );
  ANDN U5320 ( .B(y[967]), .A(x[967]), .Z(n8953) );
  OR U5321 ( .A(n8943), .B(n8953), .Z(n12157) );
  NANDN U5322 ( .A(y[965]), .B(x[965]), .Z(n8940) );
  NANDN U5323 ( .A(y[966]), .B(x[966]), .Z(n8947) );
  AND U5324 ( .A(n8940), .B(n8947), .Z(n12155) );
  ANDN U5325 ( .B(y[964]), .A(x[964]), .Z(n8936) );
  ANDN U5326 ( .B(y[965]), .A(x[965]), .Z(n8946) );
  OR U5327 ( .A(n8936), .B(n8946), .Z(n12153) );
  NANDN U5328 ( .A(y[963]), .B(x[963]), .Z(n8932) );
  NANDN U5329 ( .A(y[964]), .B(x[964]), .Z(n8941) );
  AND U5330 ( .A(n8932), .B(n8941), .Z(n12151) );
  ANDN U5331 ( .B(y[962]), .A(x[962]), .Z(n8931) );
  ANDN U5332 ( .B(y[963]), .A(x[963]), .Z(n8938) );
  OR U5333 ( .A(n8931), .B(n8938), .Z(n12149) );
  NANDN U5334 ( .A(y[962]), .B(x[962]), .Z(n12146) );
  ANDN U5335 ( .B(y[961]), .A(x[961]), .Z(n12145) );
  NANDN U5336 ( .A(y[960]), .B(x[960]), .Z(n5526) );
  ANDN U5337 ( .B(y[958]), .A(x[958]), .Z(n12137) );
  ANDN U5338 ( .B(x[955]), .A(y[955]), .Z(n8921) );
  ANDN U5339 ( .B(x[956]), .A(y[956]), .Z(n8925) );
  NOR U5340 ( .A(n8921), .B(n8925), .Z(n12131) );
  NANDN U5341 ( .A(x[954]), .B(y[954]), .Z(n8919) );
  NANDN U5342 ( .A(x[955]), .B(y[955]), .Z(n8923) );
  NAND U5343 ( .A(n8919), .B(n8923), .Z(n12129) );
  NANDN U5344 ( .A(y[953]), .B(x[953]), .Z(n8917) );
  ANDN U5345 ( .B(x[954]), .A(y[954]), .Z(n8922) );
  ANDN U5346 ( .B(n8917), .A(n8922), .Z(n12127) );
  ANDN U5347 ( .B(y[952]), .A(x[952]), .Z(n8915) );
  NANDN U5348 ( .A(x[953]), .B(y[953]), .Z(n8920) );
  NANDN U5349 ( .A(n8915), .B(n8920), .Z(n12125) );
  NANDN U5350 ( .A(y[951]), .B(x[951]), .Z(n8914) );
  ANDN U5351 ( .B(x[952]), .A(y[952]), .Z(n8918) );
  ANDN U5352 ( .B(n8914), .A(n8918), .Z(n12123) );
  ANDN U5353 ( .B(y[950]), .A(x[950]), .Z(n5533) );
  ANDN U5354 ( .B(y[951]), .A(x[951]), .Z(n8916) );
  OR U5355 ( .A(n5533), .B(n8916), .Z(n12121) );
  NANDN U5356 ( .A(y[950]), .B(x[950]), .Z(n8913) );
  ANDN U5357 ( .B(x[949]), .A(y[949]), .Z(n8910) );
  ANDN U5358 ( .B(n8913), .A(n8910), .Z(n12119) );
  ANDN U5359 ( .B(y[949]), .A(x[949]), .Z(n5532) );
  NANDN U5360 ( .A(x[948]), .B(y[948]), .Z(n8909) );
  NANDN U5361 ( .A(n5532), .B(n8909), .Z(n12117) );
  ANDN U5362 ( .B(x[947]), .A(y[947]), .Z(n8906) );
  ANDN U5363 ( .B(x[948]), .A(y[948]), .Z(n8911) );
  NOR U5364 ( .A(n8906), .B(n8911), .Z(n12115) );
  NANDN U5365 ( .A(x[946]), .B(y[946]), .Z(n8904) );
  NANDN U5366 ( .A(x[947]), .B(y[947]), .Z(n8908) );
  NAND U5367 ( .A(n8904), .B(n8908), .Z(n12113) );
  ANDN U5368 ( .B(x[945]), .A(y[945]), .Z(n8903) );
  ANDN U5369 ( .B(x[946]), .A(y[946]), .Z(n8907) );
  NOR U5370 ( .A(n8903), .B(n8907), .Z(n12111) );
  NANDN U5371 ( .A(x[944]), .B(y[944]), .Z(n8901) );
  NANDN U5372 ( .A(x[945]), .B(y[945]), .Z(n8905) );
  NAND U5373 ( .A(n8901), .B(n8905), .Z(n12109) );
  NANDN U5374 ( .A(y[943]), .B(x[943]), .Z(n4411) );
  ANDN U5375 ( .B(y[942]), .A(x[942]), .Z(n8898) );
  NANDN U5376 ( .A(x[943]), .B(y[943]), .Z(n8902) );
  NANDN U5377 ( .A(n8898), .B(n8902), .Z(n3453) );
  AND U5378 ( .A(n4411), .B(n3453), .Z(n12105) );
  ANDN U5379 ( .B(x[940]), .A(y[940]), .Z(n12099) );
  NANDN U5380 ( .A(x[938]), .B(y[938]), .Z(n5537) );
  NANDN U5381 ( .A(y[938]), .B(x[938]), .Z(n5535) );
  ANDN U5382 ( .B(x[937]), .A(y[937]), .Z(n5539) );
  NANDN U5383 ( .A(x[936]), .B(y[936]), .Z(n12089) );
  NANDN U5384 ( .A(y[936]), .B(x[936]), .Z(n5540) );
  ANDN U5385 ( .B(y[934]), .A(x[934]), .Z(n8893) );
  NANDN U5386 ( .A(x[935]), .B(y[935]), .Z(n8895) );
  NANDN U5387 ( .A(n8893), .B(n8895), .Z(n12085) );
  NANDN U5388 ( .A(y[933]), .B(x[933]), .Z(n8892) );
  NANDN U5389 ( .A(y[934]), .B(x[934]), .Z(n5541) );
  AND U5390 ( .A(n8892), .B(n5541), .Z(n12083) );
  ANDN U5391 ( .B(y[932]), .A(x[932]), .Z(n8889) );
  ANDN U5392 ( .B(y[933]), .A(x[933]), .Z(n8894) );
  OR U5393 ( .A(n8889), .B(n8894), .Z(n12081) );
  NANDN U5394 ( .A(y[931]), .B(x[931]), .Z(n8888) );
  NANDN U5395 ( .A(y[932]), .B(x[932]), .Z(n8891) );
  AND U5396 ( .A(n8888), .B(n8891), .Z(n12079) );
  ANDN U5397 ( .B(y[930]), .A(x[930]), .Z(n8887) );
  ANDN U5398 ( .B(y[931]), .A(x[931]), .Z(n8890) );
  OR U5399 ( .A(n8887), .B(n8890), .Z(n12077) );
  NANDN U5400 ( .A(y[930]), .B(x[930]), .Z(n12074) );
  NANDN U5401 ( .A(x[923]), .B(y[923]), .Z(n12056) );
  NANDN U5402 ( .A(x[922]), .B(y[922]), .Z(n12053) );
  IV U5403 ( .A(n12053), .Z(n8880) );
  ANDN U5404 ( .B(n12056), .A(n8880), .Z(n4407) );
  ANDN U5405 ( .B(x[921]), .A(y[921]), .Z(n12051) );
  NANDN U5406 ( .A(x[921]), .B(y[921]), .Z(n8879) );
  ANDN U5407 ( .B(y[920]), .A(x[920]), .Z(n8877) );
  ANDN U5408 ( .B(n8879), .A(n8877), .Z(n12049) );
  NANDN U5409 ( .A(x[912]), .B(y[912]), .Z(n5559) );
  NANDN U5410 ( .A(x[914]), .B(y[914]), .Z(n4398) );
  NANDN U5411 ( .A(x[913]), .B(y[913]), .Z(n3454) );
  AND U5412 ( .A(n4398), .B(n3454), .Z(n12037) );
  ANDN U5413 ( .B(x[912]), .A(y[912]), .Z(n5557) );
  NANDN U5414 ( .A(y[911]), .B(x[911]), .Z(n8872) );
  ANDN U5415 ( .B(y[910]), .A(x[910]), .Z(n8869) );
  NANDN U5416 ( .A(y[910]), .B(x[910]), .Z(n8871) );
  NANDN U5417 ( .A(x[908]), .B(y[908]), .Z(n12025) );
  NANDN U5418 ( .A(x[906]), .B(y[906]), .Z(n8865) );
  NANDN U5419 ( .A(x[907]), .B(y[907]), .Z(n8868) );
  NAND U5420 ( .A(n8865), .B(n8868), .Z(n12021) );
  ANDN U5421 ( .B(x[905]), .A(y[905]), .Z(n5563) );
  ANDN U5422 ( .B(x[906]), .A(y[906]), .Z(n8867) );
  NOR U5423 ( .A(n5563), .B(n8867), .Z(n12019) );
  ANDN U5424 ( .B(y[904]), .A(x[904]), .Z(n8859) );
  NANDN U5425 ( .A(x[905]), .B(y[905]), .Z(n8864) );
  NANDN U5426 ( .A(n8859), .B(n8864), .Z(n12017) );
  NANDN U5427 ( .A(y[903]), .B(x[903]), .Z(n8855) );
  ANDN U5428 ( .B(x[904]), .A(y[904]), .Z(n5562) );
  ANDN U5429 ( .B(n8855), .A(n5562), .Z(n12015) );
  NANDN U5430 ( .A(x[902]), .B(y[902]), .Z(n3455) );
  ANDN U5431 ( .B(y[903]), .A(x[903]), .Z(n8860) );
  ANDN U5432 ( .B(n3455), .A(n8860), .Z(n12013) );
  NANDN U5433 ( .A(y[901]), .B(x[901]), .Z(n8847) );
  XOR U5434 ( .A(x[902]), .B(y[902]), .Z(n8853) );
  ANDN U5435 ( .B(n8847), .A(n8853), .Z(n12011) );
  ANDN U5436 ( .B(y[900]), .A(x[900]), .Z(n8844) );
  ANDN U5437 ( .B(y[901]), .A(x[901]), .Z(n8850) );
  NOR U5438 ( .A(n8844), .B(n8850), .Z(n12009) );
  NANDN U5439 ( .A(x[898]), .B(y[898]), .Z(n5564) );
  NANDN U5440 ( .A(x[899]), .B(y[899]), .Z(n12004) );
  ANDN U5441 ( .B(x[898]), .A(y[898]), .Z(n12002) );
  NANDN U5442 ( .A(y[897]), .B(x[897]), .Z(n5567) );
  ANDN U5443 ( .B(y[896]), .A(x[896]), .Z(n11997) );
  ANDN U5444 ( .B(x[894]), .A(y[894]), .Z(n11990) );
  NANDN U5445 ( .A(x[892]), .B(y[892]), .Z(n11985) );
  ANDN U5446 ( .B(x[891]), .A(y[891]), .Z(n11983) );
  ANDN U5447 ( .B(y[890]), .A(x[890]), .Z(n8823) );
  ANDN U5448 ( .B(y[891]), .A(x[891]), .Z(n8826) );
  NOR U5449 ( .A(n8823), .B(n8826), .Z(n11980) );
  ANDN U5450 ( .B(x[890]), .A(y[890]), .Z(n11978) );
  NANDN U5451 ( .A(x[888]), .B(y[888]), .Z(n11973) );
  IV U5452 ( .A(n11973), .Z(n8817) );
  ANDN U5453 ( .B(x[887]), .A(y[887]), .Z(n11971) );
  NANDN U5454 ( .A(x[886]), .B(y[886]), .Z(n3456) );
  NANDN U5455 ( .A(x[887]), .B(y[887]), .Z(n8816) );
  AND U5456 ( .A(n3456), .B(n8816), .Z(n11968) );
  IV U5457 ( .A(n11968), .Z(n4394) );
  NANDN U5458 ( .A(y[883]), .B(x[883]), .Z(n8802) );
  NANDN U5459 ( .A(y[884]), .B(x[884]), .Z(n8809) );
  NAND U5460 ( .A(n8802), .B(n8809), .Z(n11963) );
  NANDN U5461 ( .A(x[881]), .B(y[881]), .Z(n5573) );
  NANDN U5462 ( .A(x[880]), .B(y[880]), .Z(n5577) );
  NANDN U5463 ( .A(y[879]), .B(x[879]), .Z(n5580) );
  NANDN U5464 ( .A(x[879]), .B(y[879]), .Z(n5578) );
  NANDN U5465 ( .A(y[877]), .B(x[877]), .Z(n5584) );
  NANDN U5466 ( .A(x[876]), .B(y[876]), .Z(n5587) );
  NANDN U5467 ( .A(y[873]), .B(x[873]), .Z(n3458) );
  NANDN U5468 ( .A(y[874]), .B(x[874]), .Z(n3457) );
  NAND U5469 ( .A(n3458), .B(n3457), .Z(n5593) );
  NANDN U5470 ( .A(x[873]), .B(y[873]), .Z(n5588) );
  NANDN U5471 ( .A(x[872]), .B(y[872]), .Z(n3459) );
  AND U5472 ( .A(n5588), .B(n3459), .Z(n11941) );
  ANDN U5473 ( .B(x[871]), .A(y[871]), .Z(n11939) );
  NANDN U5474 ( .A(x[870]), .B(y[870]), .Z(n3460) );
  ANDN U5475 ( .B(y[871]), .A(x[871]), .Z(n5595) );
  ANDN U5476 ( .B(n3460), .A(n5595), .Z(n11937) );
  NANDN U5477 ( .A(y[869]), .B(x[869]), .Z(n8799) );
  NANDN U5478 ( .A(y[870]), .B(x[870]), .Z(n5594) );
  NAND U5479 ( .A(n8799), .B(n5594), .Z(n11935) );
  NANDN U5480 ( .A(x[868]), .B(y[868]), .Z(n5597) );
  NANDN U5481 ( .A(x[869]), .B(y[869]), .Z(n8801) );
  AND U5482 ( .A(n5597), .B(n8801), .Z(n11933) );
  ANDN U5483 ( .B(x[867]), .A(y[867]), .Z(n8794) );
  NANDN U5484 ( .A(y[868]), .B(x[868]), .Z(n8800) );
  NANDN U5485 ( .A(n8794), .B(n8800), .Z(n11931) );
  NANDN U5486 ( .A(x[866]), .B(y[866]), .Z(n8790) );
  NANDN U5487 ( .A(x[867]), .B(y[867]), .Z(n5596) );
  AND U5488 ( .A(n8790), .B(n5596), .Z(n11929) );
  ANDN U5489 ( .B(x[865]), .A(y[865]), .Z(n8789) );
  ANDN U5490 ( .B(x[866]), .A(y[866]), .Z(n8795) );
  OR U5491 ( .A(n8789), .B(n8795), .Z(n11927) );
  NANDN U5492 ( .A(x[865]), .B(y[865]), .Z(n11925) );
  NANDN U5493 ( .A(x[863]), .B(y[863]), .Z(n5598) );
  NANDN U5494 ( .A(x[862]), .B(y[862]), .Z(n5603) );
  NANDN U5495 ( .A(y[861]), .B(x[861]), .Z(n5604) );
  NANDN U5496 ( .A(x[861]), .B(y[861]), .Z(n5602) );
  ANDN U5497 ( .B(x[859]), .A(y[859]), .Z(n5609) );
  NANDN U5498 ( .A(x[858]), .B(y[858]), .Z(n11908) );
  NANDN U5499 ( .A(x[857]), .B(y[857]), .Z(n5610) );
  ANDN U5500 ( .B(y[856]), .A(x[856]), .Z(n5611) );
  ANDN U5501 ( .B(n5610), .A(n5611), .Z(n11905) );
  NANDN U5502 ( .A(y[856]), .B(x[856]), .Z(n5614) );
  NANDN U5503 ( .A(y[855]), .B(x[855]), .Z(n3461) );
  AND U5504 ( .A(n5614), .B(n3461), .Z(n11902) );
  NANDN U5505 ( .A(x[854]), .B(y[854]), .Z(n8773) );
  ANDN U5506 ( .B(y[855]), .A(x[855]), .Z(n5612) );
  ANDN U5507 ( .B(n8773), .A(n5612), .Z(n11901) );
  ANDN U5508 ( .B(x[853]), .A(y[853]), .Z(n8771) );
  NANDN U5509 ( .A(y[854]), .B(x[854]), .Z(n8777) );
  NANDN U5510 ( .A(n8771), .B(n8777), .Z(n11899) );
  NANDN U5511 ( .A(x[852]), .B(y[852]), .Z(n8770) );
  ANDN U5512 ( .B(y[853]), .A(x[853]), .Z(n8774) );
  ANDN U5513 ( .B(n8770), .A(n8774), .Z(n11897) );
  ANDN U5514 ( .B(x[851]), .A(y[851]), .Z(n8769) );
  ANDN U5515 ( .B(x[852]), .A(y[852]), .Z(n8772) );
  OR U5516 ( .A(n8769), .B(n8772), .Z(n11895) );
  NANDN U5517 ( .A(x[850]), .B(y[850]), .Z(n5620) );
  NANDN U5518 ( .A(x[851]), .B(y[851]), .Z(n11893) );
  ANDN U5519 ( .B(x[850]), .A(y[850]), .Z(n11891) );
  NANDN U5520 ( .A(x[849]), .B(y[849]), .Z(n5619) );
  NANDN U5521 ( .A(y[847]), .B(x[847]), .Z(n11883) );
  NANDN U5522 ( .A(x[846]), .B(y[846]), .Z(n5624) );
  NANDN U5523 ( .A(x[847]), .B(y[847]), .Z(n5623) );
  AND U5524 ( .A(n5624), .B(n5623), .Z(n11881) );
  NANDN U5525 ( .A(x[845]), .B(y[845]), .Z(n5625) );
  NANDN U5526 ( .A(y[845]), .B(x[845]), .Z(n3463) );
  NANDN U5527 ( .A(y[844]), .B(x[844]), .Z(n3462) );
  AND U5528 ( .A(n3463), .B(n3462), .Z(n8768) );
  ANDN U5529 ( .B(n5625), .A(n8768), .Z(n11877) );
  NANDN U5530 ( .A(y[843]), .B(x[843]), .Z(n3471) );
  XNOR U5531 ( .A(y[843]), .B(x[843]), .Z(n3465) );
  NANDN U5532 ( .A(x[842]), .B(y[842]), .Z(n3464) );
  NAND U5533 ( .A(n3465), .B(n3464), .Z(n3466) );
  NAND U5534 ( .A(n3471), .B(n3466), .Z(n3468) );
  NANDN U5535 ( .A(x[844]), .B(y[844]), .Z(n3467) );
  NAND U5536 ( .A(n3468), .B(n3467), .Z(n8767) );
  ANDN U5537 ( .B(n5625), .A(n8767), .Z(n11875) );
  NANDN U5538 ( .A(y[842]), .B(x[842]), .Z(n3470) );
  NANDN U5539 ( .A(y[841]), .B(x[841]), .Z(n3469) );
  AND U5540 ( .A(n3470), .B(n3469), .Z(n3472) );
  NAND U5541 ( .A(n3472), .B(n3471), .Z(n5628) );
  NANDN U5542 ( .A(x[841]), .B(y[841]), .Z(n5627) );
  ANDN U5543 ( .B(x[839]), .A(y[839]), .Z(n11869) );
  NANDN U5544 ( .A(x[838]), .B(y[838]), .Z(n8757) );
  NANDN U5545 ( .A(x[839]), .B(y[839]), .Z(n8763) );
  AND U5546 ( .A(n8757), .B(n8763), .Z(n11867) );
  ANDN U5547 ( .B(x[838]), .A(y[838]), .Z(n8760) );
  NANDN U5548 ( .A(y[837]), .B(x[837]), .Z(n8752) );
  NANDN U5549 ( .A(n8760), .B(n8752), .Z(n11865) );
  NANDN U5550 ( .A(x[836]), .B(y[836]), .Z(n5631) );
  NANDN U5551 ( .A(x[837]), .B(y[837]), .Z(n8758) );
  AND U5552 ( .A(n5631), .B(n8758), .Z(n11863) );
  ANDN U5553 ( .B(x[835]), .A(y[835]), .Z(n8747) );
  NANDN U5554 ( .A(y[836]), .B(x[836]), .Z(n8753) );
  NANDN U5555 ( .A(n8747), .B(n8753), .Z(n11861) );
  NANDN U5556 ( .A(x[834]), .B(y[834]), .Z(n8743) );
  NANDN U5557 ( .A(x[835]), .B(y[835]), .Z(n5630) );
  AND U5558 ( .A(n8743), .B(n5630), .Z(n11859) );
  ANDN U5559 ( .B(x[833]), .A(y[833]), .Z(n8739) );
  ANDN U5560 ( .B(x[834]), .A(y[834]), .Z(n8748) );
  OR U5561 ( .A(n8739), .B(n8748), .Z(n11857) );
  NANDN U5562 ( .A(x[832]), .B(y[832]), .Z(n8737) );
  NANDN U5563 ( .A(x[833]), .B(y[833]), .Z(n8742) );
  AND U5564 ( .A(n8737), .B(n8742), .Z(n11855) );
  ANDN U5565 ( .B(x[832]), .A(y[832]), .Z(n11853) );
  NANDN U5566 ( .A(x[830]), .B(y[830]), .Z(n5633) );
  NANDN U5567 ( .A(y[829]), .B(x[829]), .Z(n5634) );
  NANDN U5568 ( .A(x[828]), .B(y[828]), .Z(n11842) );
  NANDN U5569 ( .A(x[827]), .B(y[827]), .Z(n8731) );
  ANDN U5570 ( .B(y[826]), .A(x[826]), .Z(n8730) );
  ANDN U5571 ( .B(n8731), .A(n8730), .Z(n11839) );
  ANDN U5572 ( .B(y[824]), .A(x[824]), .Z(n11831) );
  IV U5573 ( .A(n11831), .Z(n8728) );
  ANDN U5574 ( .B(y[825]), .A(x[825]), .Z(n11834) );
  ANDN U5575 ( .B(n8728), .A(n11834), .Z(n4382) );
  ANDN U5576 ( .B(y[822]), .A(x[822]), .Z(n8725) );
  ANDN U5577 ( .B(y[823]), .A(x[823]), .Z(n8729) );
  NOR U5578 ( .A(n8725), .B(n8729), .Z(n11827) );
  NANDN U5579 ( .A(y[821]), .B(x[821]), .Z(n8724) );
  NANDN U5580 ( .A(y[822]), .B(x[822]), .Z(n8727) );
  NAND U5581 ( .A(n8724), .B(n8727), .Z(n11825) );
  NANDN U5582 ( .A(x[820]), .B(y[820]), .Z(n5638) );
  ANDN U5583 ( .B(y[821]), .A(x[821]), .Z(n8726) );
  ANDN U5584 ( .B(n5638), .A(n8726), .Z(n11823) );
  NANDN U5585 ( .A(y[819]), .B(x[819]), .Z(n5640) );
  NANDN U5586 ( .A(y[820]), .B(x[820]), .Z(n8723) );
  NAND U5587 ( .A(n5640), .B(n8723), .Z(n11821) );
  NANDN U5588 ( .A(x[819]), .B(y[819]), .Z(n5639) );
  ANDN U5589 ( .B(y[818]), .A(x[818]), .Z(n8716) );
  ANDN U5590 ( .B(n5639), .A(n8716), .Z(n11819) );
  NANDN U5591 ( .A(y[817]), .B(x[817]), .Z(n8712) );
  NANDN U5592 ( .A(y[818]), .B(x[818]), .Z(n5641) );
  NAND U5593 ( .A(n8712), .B(n5641), .Z(n11817) );
  NANDN U5594 ( .A(x[816]), .B(y[816]), .Z(n5642) );
  ANDN U5595 ( .B(y[817]), .A(x[817]), .Z(n8717) );
  ANDN U5596 ( .B(n5642), .A(n8717), .Z(n11815) );
  NANDN U5597 ( .A(y[815]), .B(x[815]), .Z(n5644) );
  NANDN U5598 ( .A(y[816]), .B(x[816]), .Z(n8711) );
  NAND U5599 ( .A(n5644), .B(n8711), .Z(n11813) );
  NANDN U5600 ( .A(x[815]), .B(y[815]), .Z(n5643) );
  ANDN U5601 ( .B(y[814]), .A(x[814]), .Z(n8704) );
  ANDN U5602 ( .B(n5643), .A(n8704), .Z(n11811) );
  NANDN U5603 ( .A(y[813]), .B(x[813]), .Z(n8700) );
  NANDN U5604 ( .A(y[814]), .B(x[814]), .Z(n5645) );
  NAND U5605 ( .A(n8700), .B(n5645), .Z(n11809) );
  ANDN U5606 ( .B(y[812]), .A(x[812]), .Z(n5647) );
  ANDN U5607 ( .B(y[813]), .A(x[813]), .Z(n8705) );
  NOR U5608 ( .A(n5647), .B(n8705), .Z(n11807) );
  ANDN U5609 ( .B(x[811]), .A(y[811]), .Z(n8694) );
  XNOR U5610 ( .A(y[812]), .B(x[812]), .Z(n3473) );
  NANDN U5611 ( .A(n8694), .B(n3473), .Z(n11805) );
  NANDN U5612 ( .A(x[810]), .B(y[810]), .Z(n8690) );
  ANDN U5613 ( .B(y[811]), .A(x[811]), .Z(n5646) );
  ANDN U5614 ( .B(n8690), .A(n5646), .Z(n11803) );
  ANDN U5615 ( .B(x[809]), .A(y[809]), .Z(n8688) );
  ANDN U5616 ( .B(x[810]), .A(y[810]), .Z(n8695) );
  OR U5617 ( .A(n8688), .B(n8695), .Z(n11801) );
  NANDN U5618 ( .A(x[808]), .B(y[808]), .Z(n3474) );
  NANDN U5619 ( .A(x[809]), .B(y[809]), .Z(n8689) );
  AND U5620 ( .A(n3474), .B(n8689), .Z(n11799) );
  XNOR U5621 ( .A(x[808]), .B(y[808]), .Z(n8682) );
  NANDN U5622 ( .A(y[807]), .B(x[807]), .Z(n8677) );
  NAND U5623 ( .A(n8682), .B(n8677), .Z(n11797) );
  NANDN U5624 ( .A(x[806]), .B(y[806]), .Z(n5649) );
  NANDN U5625 ( .A(x[807]), .B(y[807]), .Z(n8683) );
  AND U5626 ( .A(n5649), .B(n8683), .Z(n11795) );
  ANDN U5627 ( .B(x[805]), .A(y[805]), .Z(n8672) );
  NANDN U5628 ( .A(y[806]), .B(x[806]), .Z(n8678) );
  NANDN U5629 ( .A(n8672), .B(n8678), .Z(n11793) );
  NANDN U5630 ( .A(x[804]), .B(y[804]), .Z(n8668) );
  NANDN U5631 ( .A(x[805]), .B(y[805]), .Z(n5648) );
  AND U5632 ( .A(n8668), .B(n5648), .Z(n11791) );
  ANDN U5633 ( .B(x[803]), .A(y[803]), .Z(n8663) );
  ANDN U5634 ( .B(x[804]), .A(y[804]), .Z(n8673) );
  OR U5635 ( .A(n8663), .B(n8673), .Z(n11789) );
  NANDN U5636 ( .A(x[802]), .B(y[802]), .Z(n8660) );
  NANDN U5637 ( .A(x[803]), .B(y[803]), .Z(n8667) );
  AND U5638 ( .A(n8660), .B(n8667), .Z(n11787) );
  ANDN U5639 ( .B(x[801]), .A(y[801]), .Z(n8656) );
  XNOR U5640 ( .A(y[802]), .B(x[802]), .Z(n3475) );
  NANDN U5641 ( .A(n8656), .B(n3475), .Z(n11785) );
  NANDN U5642 ( .A(x[800]), .B(y[800]), .Z(n8652) );
  NANDN U5643 ( .A(x[801]), .B(y[801]), .Z(n8661) );
  AND U5644 ( .A(n8652), .B(n8661), .Z(n11783) );
  ANDN U5645 ( .B(x[799]), .A(y[799]), .Z(n5651) );
  ANDN U5646 ( .B(x[800]), .A(y[800]), .Z(n8658) );
  OR U5647 ( .A(n5651), .B(n8658), .Z(n11781) );
  NANDN U5648 ( .A(x[799]), .B(y[799]), .Z(n8651) );
  ANDN U5649 ( .B(y[798]), .A(x[798]), .Z(n8646) );
  ANDN U5650 ( .B(n8651), .A(n8646), .Z(n11779) );
  ANDN U5651 ( .B(x[798]), .A(y[798]), .Z(n5650) );
  NANDN U5652 ( .A(y[797]), .B(x[797]), .Z(n8642) );
  NANDN U5653 ( .A(n5650), .B(n8642), .Z(n11777) );
  ANDN U5654 ( .B(y[796]), .A(x[796]), .Z(n5653) );
  ANDN U5655 ( .B(y[797]), .A(x[797]), .Z(n8647) );
  NOR U5656 ( .A(n5653), .B(n8647), .Z(n11775) );
  ANDN U5657 ( .B(x[795]), .A(y[795]), .Z(n8636) );
  NANDN U5658 ( .A(y[796]), .B(x[796]), .Z(n8641) );
  NANDN U5659 ( .A(n8636), .B(n8641), .Z(n11773) );
  NANDN U5660 ( .A(x[794]), .B(y[794]), .Z(n5654) );
  ANDN U5661 ( .B(y[795]), .A(x[795]), .Z(n5652) );
  ANDN U5662 ( .B(n5654), .A(n5652), .Z(n11771) );
  ANDN U5663 ( .B(x[794]), .A(y[794]), .Z(n8637) );
  NANDN U5664 ( .A(y[793]), .B(x[793]), .Z(n8630) );
  NANDN U5665 ( .A(n8637), .B(n8630), .Z(n11769) );
  NANDN U5666 ( .A(x[793]), .B(y[793]), .Z(n5655) );
  ANDN U5667 ( .B(y[792]), .A(x[792]), .Z(n8628) );
  ANDN U5668 ( .B(n5655), .A(n8628), .Z(n11767) );
  ANDN U5669 ( .B(x[792]), .A(y[792]), .Z(n8632) );
  NANDN U5670 ( .A(y[791]), .B(x[791]), .Z(n5656) );
  NANDN U5671 ( .A(n8632), .B(n5656), .Z(n11765) );
  NANDN U5672 ( .A(x[790]), .B(y[790]), .Z(n8620) );
  ANDN U5673 ( .B(y[791]), .A(x[791]), .Z(n8625) );
  ANDN U5674 ( .B(n8620), .A(n8625), .Z(n11763) );
  ANDN U5675 ( .B(x[789]), .A(y[789]), .Z(n8616) );
  XNOR U5676 ( .A(y[790]), .B(x[790]), .Z(n3476) );
  NANDN U5677 ( .A(n8616), .B(n3476), .Z(n11761) );
  NANDN U5678 ( .A(x[788]), .B(y[788]), .Z(n8614) );
  ANDN U5679 ( .B(y[789]), .A(x[789]), .Z(n8622) );
  ANDN U5680 ( .B(n8614), .A(n8622), .Z(n11759) );
  XNOR U5681 ( .A(x[788]), .B(y[788]), .Z(n3477) );
  ANDN U5682 ( .B(x[787]), .A(y[787]), .Z(n8612) );
  ANDN U5683 ( .B(n3477), .A(n8612), .Z(n11757) );
  IV U5684 ( .A(n11757), .Z(n4343) );
  NANDN U5685 ( .A(x[787]), .B(y[787]), .Z(n3479) );
  NANDN U5686 ( .A(x[786]), .B(y[786]), .Z(n3478) );
  NAND U5687 ( .A(n3479), .B(n3478), .Z(n11755) );
  NANDN U5688 ( .A(y[785]), .B(x[785]), .Z(n3481) );
  NANDN U5689 ( .A(y[786]), .B(x[786]), .Z(n3480) );
  AND U5690 ( .A(n3481), .B(n3480), .Z(n11752) );
  NANDN U5691 ( .A(x[783]), .B(y[783]), .Z(n3483) );
  NANDN U5692 ( .A(x[782]), .B(y[782]), .Z(n3482) );
  NAND U5693 ( .A(n3483), .B(n3482), .Z(n11747) );
  IV U5694 ( .A(n11747), .Z(n8603) );
  NANDN U5695 ( .A(y[781]), .B(x[781]), .Z(n3485) );
  NANDN U5696 ( .A(y[782]), .B(x[782]), .Z(n3484) );
  AND U5697 ( .A(n3485), .B(n3484), .Z(n11745) );
  IV U5698 ( .A(n11745), .Z(n8601) );
  NANDN U5699 ( .A(x[781]), .B(y[781]), .Z(n3487) );
  NANDN U5700 ( .A(x[780]), .B(y[780]), .Z(n3486) );
  NAND U5701 ( .A(n3487), .B(n3486), .Z(n11743) );
  IV U5702 ( .A(n11743), .Z(n8600) );
  NANDN U5703 ( .A(y[779]), .B(x[779]), .Z(n3489) );
  NANDN U5704 ( .A(y[780]), .B(x[780]), .Z(n3488) );
  AND U5705 ( .A(n3489), .B(n3488), .Z(n11740) );
  IV U5706 ( .A(n11740), .Z(n8598) );
  NANDN U5707 ( .A(x[777]), .B(y[777]), .Z(n3491) );
  NANDN U5708 ( .A(x[776]), .B(y[776]), .Z(n3490) );
  NAND U5709 ( .A(n3491), .B(n3490), .Z(n11735) );
  IV U5710 ( .A(n11735), .Z(n8591) );
  NANDN U5711 ( .A(y[775]), .B(x[775]), .Z(n3493) );
  NANDN U5712 ( .A(y[776]), .B(x[776]), .Z(n3492) );
  AND U5713 ( .A(n3493), .B(n3492), .Z(n11733) );
  IV U5714 ( .A(n11733), .Z(n8589) );
  NANDN U5715 ( .A(x[775]), .B(y[775]), .Z(n3495) );
  NANDN U5716 ( .A(x[774]), .B(y[774]), .Z(n3494) );
  NAND U5717 ( .A(n3495), .B(n3494), .Z(n11731) );
  IV U5718 ( .A(n11731), .Z(n8587) );
  NANDN U5719 ( .A(y[774]), .B(x[774]), .Z(n8586) );
  NANDN U5720 ( .A(y[773]), .B(x[773]), .Z(n3496) );
  AND U5721 ( .A(n8586), .B(n3496), .Z(n11728) );
  NANDN U5722 ( .A(x[770]), .B(y[770]), .Z(n5659) );
  NANDN U5723 ( .A(x[771]), .B(y[771]), .Z(n8577) );
  NAND U5724 ( .A(n5659), .B(n8577), .Z(n11723) );
  IV U5725 ( .A(n11723), .Z(n4332) );
  NANDN U5726 ( .A(y[770]), .B(x[770]), .Z(n8572) );
  ANDN U5727 ( .B(x[769]), .A(y[769]), .Z(n8566) );
  ANDN U5728 ( .B(n8572), .A(n8566), .Z(n11721) );
  NANDN U5729 ( .A(x[768]), .B(y[768]), .Z(n8562) );
  NANDN U5730 ( .A(x[769]), .B(y[769]), .Z(n5658) );
  NAND U5731 ( .A(n8562), .B(n5658), .Z(n11719) );
  ANDN U5732 ( .B(x[767]), .A(y[767]), .Z(n5661) );
  ANDN U5733 ( .B(x[768]), .A(y[768]), .Z(n8567) );
  NOR U5734 ( .A(n5661), .B(n8567), .Z(n11716) );
  NANDN U5735 ( .A(x[765]), .B(y[765]), .Z(n3498) );
  NANDN U5736 ( .A(x[764]), .B(y[764]), .Z(n3497) );
  NAND U5737 ( .A(n3498), .B(n3497), .Z(n11711) );
  IV U5738 ( .A(n11711), .Z(n8553) );
  NANDN U5739 ( .A(y[763]), .B(x[763]), .Z(n3500) );
  NANDN U5740 ( .A(y[764]), .B(x[764]), .Z(n3499) );
  AND U5741 ( .A(n3500), .B(n3499), .Z(n11709) );
  IV U5742 ( .A(n11709), .Z(n5664) );
  NANDN U5743 ( .A(x[762]), .B(y[762]), .Z(n3501) );
  ANDN U5744 ( .B(y[763]), .A(x[763]), .Z(n5663) );
  ANDN U5745 ( .B(n3501), .A(n5663), .Z(n11707) );
  NANDN U5746 ( .A(y[761]), .B(x[761]), .Z(n5666) );
  XNOR U5747 ( .A(y[762]), .B(x[762]), .Z(n3502) );
  AND U5748 ( .A(n5666), .B(n3502), .Z(n11704) );
  NANDN U5749 ( .A(x[758]), .B(y[758]), .Z(n8535) );
  ANDN U5750 ( .B(y[759]), .A(x[759]), .Z(n8545) );
  ANDN U5751 ( .B(n8535), .A(n8545), .Z(n11699) );
  NANDN U5752 ( .A(y[757]), .B(x[757]), .Z(n5668) );
  ANDN U5753 ( .B(x[758]), .A(y[758]), .Z(n8541) );
  ANDN U5754 ( .B(n5668), .A(n8541), .Z(n11697) );
  NANDN U5755 ( .A(x[756]), .B(y[756]), .Z(n5670) );
  NANDN U5756 ( .A(x[757]), .B(y[757]), .Z(n8534) );
  NAND U5757 ( .A(n5670), .B(n8534), .Z(n11695) );
  NANDN U5758 ( .A(y[756]), .B(x[756]), .Z(n5669) );
  ANDN U5759 ( .B(x[755]), .A(y[755]), .Z(n8527) );
  ANDN U5760 ( .B(n5669), .A(n8527), .Z(n11692) );
  NANDN U5761 ( .A(x[752]), .B(y[752]), .Z(n5674) );
  NANDN U5762 ( .A(x[753]), .B(y[753]), .Z(n8522) );
  NAND U5763 ( .A(n5674), .B(n8522), .Z(n11687) );
  NANDN U5764 ( .A(y[752]), .B(x[752]), .Z(n5673) );
  ANDN U5765 ( .B(x[751]), .A(y[751]), .Z(n8515) );
  ANDN U5766 ( .B(n5673), .A(n8515), .Z(n11685) );
  NANDN U5767 ( .A(x[750]), .B(y[750]), .Z(n8511) );
  NANDN U5768 ( .A(x[751]), .B(y[751]), .Z(n5675) );
  NAND U5769 ( .A(n8511), .B(n5675), .Z(n11683) );
  NANDN U5770 ( .A(y[749]), .B(x[749]), .Z(n5676) );
  ANDN U5771 ( .B(x[750]), .A(y[750]), .Z(n8516) );
  ANDN U5772 ( .B(n5676), .A(n8516), .Z(n11680) );
  NANDN U5773 ( .A(x[746]), .B(y[746]), .Z(n8499) );
  NANDN U5774 ( .A(x[747]), .B(y[747]), .Z(n5679) );
  NAND U5775 ( .A(n8499), .B(n5679), .Z(n11675) );
  IV U5776 ( .A(n11675), .Z(n4328) );
  NANDN U5777 ( .A(y[745]), .B(x[745]), .Z(n5680) );
  ANDN U5778 ( .B(x[746]), .A(y[746]), .Z(n8504) );
  ANDN U5779 ( .B(n5680), .A(n8504), .Z(n11673) );
  NANDN U5780 ( .A(x[744]), .B(y[744]), .Z(n5682) );
  NANDN U5781 ( .A(x[745]), .B(y[745]), .Z(n8498) );
  NAND U5782 ( .A(n5682), .B(n8498), .Z(n11671) );
  NANDN U5783 ( .A(y[744]), .B(x[744]), .Z(n5681) );
  ANDN U5784 ( .B(x[743]), .A(y[743]), .Z(n8491) );
  ANDN U5785 ( .B(n5681), .A(n8491), .Z(n11668) );
  NANDN U5786 ( .A(x[740]), .B(y[740]), .Z(n5686) );
  NANDN U5787 ( .A(x[741]), .B(y[741]), .Z(n8486) );
  NAND U5788 ( .A(n5686), .B(n8486), .Z(n11663) );
  NANDN U5789 ( .A(y[740]), .B(x[740]), .Z(n5685) );
  ANDN U5790 ( .B(x[739]), .A(y[739]), .Z(n8479) );
  ANDN U5791 ( .B(n5685), .A(n8479), .Z(n11661) );
  NANDN U5792 ( .A(x[738]), .B(y[738]), .Z(n8475) );
  NANDN U5793 ( .A(x[739]), .B(y[739]), .Z(n5687) );
  NAND U5794 ( .A(n8475), .B(n5687), .Z(n11659) );
  NANDN U5795 ( .A(y[737]), .B(x[737]), .Z(n5688) );
  ANDN U5796 ( .B(x[738]), .A(y[738]), .Z(n8480) );
  ANDN U5797 ( .B(n5688), .A(n8480), .Z(n11656) );
  NANDN U5798 ( .A(x[734]), .B(y[734]), .Z(n3503) );
  NANDN U5799 ( .A(x[735]), .B(y[735]), .Z(n5691) );
  NAND U5800 ( .A(n3503), .B(n5691), .Z(n11651) );
  XNOR U5801 ( .A(x[734]), .B(y[734]), .Z(n8463) );
  NANDN U5802 ( .A(y[733]), .B(x[733]), .Z(n5693) );
  AND U5803 ( .A(n8463), .B(n5693), .Z(n11649) );
  NANDN U5804 ( .A(x[732]), .B(y[732]), .Z(n8457) );
  NANDN U5805 ( .A(x[733]), .B(y[733]), .Z(n8462) );
  NAND U5806 ( .A(n8457), .B(n8462), .Z(n11647) );
  XNOR U5807 ( .A(y[732]), .B(x[732]), .Z(n3504) );
  ANDN U5808 ( .B(x[731]), .A(y[731]), .Z(n8453) );
  ANDN U5809 ( .B(n3504), .A(n8453), .Z(n11644) );
  NANDN U5810 ( .A(x[729]), .B(y[729]), .Z(n3506) );
  NANDN U5811 ( .A(x[728]), .B(y[728]), .Z(n3505) );
  NAND U5812 ( .A(n3506), .B(n3505), .Z(n11639) );
  NANDN U5813 ( .A(y[727]), .B(x[727]), .Z(n3508) );
  NANDN U5814 ( .A(y[728]), .B(x[728]), .Z(n3507) );
  AND U5815 ( .A(n3508), .B(n3507), .Z(n11637) );
  NANDN U5816 ( .A(x[726]), .B(y[726]), .Z(n3509) );
  NANDN U5817 ( .A(x[727]), .B(y[727]), .Z(n5694) );
  NAND U5818 ( .A(n3509), .B(n5694), .Z(n11635) );
  NANDN U5819 ( .A(y[725]), .B(x[725]), .Z(n8438) );
  XNOR U5820 ( .A(y[726]), .B(x[726]), .Z(n3510) );
  AND U5821 ( .A(n8438), .B(n3510), .Z(n11632) );
  NANDN U5822 ( .A(x[722]), .B(y[722]), .Z(n5696) );
  ANDN U5823 ( .B(y[723]), .A(x[723]), .Z(n8436) );
  ANDN U5824 ( .B(n5696), .A(n8436), .Z(n11627) );
  NANDN U5825 ( .A(y[721]), .B(x[721]), .Z(n5698) );
  NANDN U5826 ( .A(y[722]), .B(x[722]), .Z(n8429) );
  AND U5827 ( .A(n5698), .B(n8429), .Z(n11625) );
  NANDN U5828 ( .A(x[721]), .B(y[721]), .Z(n5697) );
  ANDN U5829 ( .B(y[720]), .A(x[720]), .Z(n8422) );
  ANDN U5830 ( .B(n5697), .A(n8422), .Z(n11623) );
  NANDN U5831 ( .A(y[719]), .B(x[719]), .Z(n8418) );
  NANDN U5832 ( .A(y[720]), .B(x[720]), .Z(n5699) );
  AND U5833 ( .A(n8418), .B(n5699), .Z(n11620) );
  NANDN U5834 ( .A(x[717]), .B(y[717]), .Z(n3512) );
  NANDN U5835 ( .A(x[716]), .B(y[716]), .Z(n3511) );
  NAND U5836 ( .A(n3512), .B(n3511), .Z(n11615) );
  NANDN U5837 ( .A(x[715]), .B(y[715]), .Z(n3514) );
  NANDN U5838 ( .A(x[714]), .B(y[714]), .Z(n3513) );
  AND U5839 ( .A(n3514), .B(n3513), .Z(n11611) );
  NANDN U5840 ( .A(y[713]), .B(x[713]), .Z(n3516) );
  NANDN U5841 ( .A(y[714]), .B(x[714]), .Z(n3515) );
  NAND U5842 ( .A(n3516), .B(n3515), .Z(n11609) );
  NANDN U5843 ( .A(x[713]), .B(y[713]), .Z(n8408) );
  NANDN U5844 ( .A(x[712]), .B(y[712]), .Z(n3517) );
  AND U5845 ( .A(n8408), .B(n3517), .Z(n11607) );
  ANDN U5846 ( .B(x[711]), .A(y[711]), .Z(n5701) );
  NANDN U5847 ( .A(y[712]), .B(x[712]), .Z(n8406) );
  NANDN U5848 ( .A(n5701), .B(n8406), .Z(n11605) );
  NANDN U5849 ( .A(x[711]), .B(y[711]), .Z(n8401) );
  ANDN U5850 ( .B(y[710]), .A(x[710]), .Z(n8396) );
  ANDN U5851 ( .B(n8401), .A(n8396), .Z(n11603) );
  ANDN U5852 ( .B(x[710]), .A(y[710]), .Z(n5700) );
  NANDN U5853 ( .A(y[709]), .B(x[709]), .Z(n8392) );
  NANDN U5854 ( .A(n5700), .B(n8392), .Z(n11601) );
  ANDN U5855 ( .B(y[708]), .A(x[708]), .Z(n8387) );
  ANDN U5856 ( .B(y[709]), .A(x[709]), .Z(n8397) );
  NOR U5857 ( .A(n8387), .B(n8397), .Z(n11599) );
  NANDN U5858 ( .A(y[707]), .B(x[707]), .Z(n8384) );
  NANDN U5859 ( .A(y[708]), .B(x[708]), .Z(n8391) );
  NAND U5860 ( .A(n8384), .B(n8391), .Z(n11597) );
  ANDN U5861 ( .B(y[706]), .A(x[706]), .Z(n8380) );
  ANDN U5862 ( .B(y[707]), .A(x[707]), .Z(n8390) );
  NOR U5863 ( .A(n8380), .B(n8390), .Z(n11595) );
  NANDN U5864 ( .A(y[705]), .B(x[705]), .Z(n8376) );
  XNOR U5865 ( .A(y[706]), .B(x[706]), .Z(n3518) );
  NAND U5866 ( .A(n8376), .B(n3518), .Z(n11593) );
  NANDN U5867 ( .A(x[704]), .B(y[704]), .Z(n8374) );
  ANDN U5868 ( .B(y[705]), .A(x[705]), .Z(n8382) );
  ANDN U5869 ( .B(n8374), .A(n8382), .Z(n11591) );
  ANDN U5870 ( .B(x[703]), .A(y[703]), .Z(n8372) );
  NANDN U5871 ( .A(y[704]), .B(x[704]), .Z(n8378) );
  NANDN U5872 ( .A(n8372), .B(n8378), .Z(n11589) );
  NANDN U5873 ( .A(x[703]), .B(y[703]), .Z(n3520) );
  NANDN U5874 ( .A(x[702]), .B(y[702]), .Z(n3519) );
  AND U5875 ( .A(n3520), .B(n3519), .Z(n11587) );
  NANDN U5876 ( .A(y[701]), .B(x[701]), .Z(n3522) );
  NANDN U5877 ( .A(y[702]), .B(x[702]), .Z(n3521) );
  NAND U5878 ( .A(n3522), .B(n3521), .Z(n11585) );
  NANDN U5879 ( .A(x[701]), .B(y[701]), .Z(n5702) );
  NANDN U5880 ( .A(x[700]), .B(y[700]), .Z(n3523) );
  AND U5881 ( .A(n5702), .B(n3523), .Z(n11583) );
  ANDN U5882 ( .B(x[699]), .A(y[699]), .Z(n8361) );
  ANDN U5883 ( .B(x[700]), .A(y[700]), .Z(n5703) );
  OR U5884 ( .A(n8361), .B(n5703), .Z(n11581) );
  NANDN U5885 ( .A(x[698]), .B(y[698]), .Z(n8359) );
  NANDN U5886 ( .A(x[699]), .B(y[699]), .Z(n8365) );
  AND U5887 ( .A(n8359), .B(n8365), .Z(n11579) );
  ANDN U5888 ( .B(x[697]), .A(y[697]), .Z(n5704) );
  ANDN U5889 ( .B(x[698]), .A(y[698]), .Z(n8363) );
  OR U5890 ( .A(n5704), .B(n8363), .Z(n11577) );
  NANDN U5891 ( .A(x[697]), .B(y[697]), .Z(n5707) );
  NANDN U5892 ( .A(x[696]), .B(y[696]), .Z(n3524) );
  AND U5893 ( .A(n5707), .B(n3524), .Z(n11575) );
  ANDN U5894 ( .B(x[695]), .A(y[695]), .Z(n8351) );
  XNOR U5895 ( .A(y[696]), .B(x[696]), .Z(n3525) );
  NANDN U5896 ( .A(n8351), .B(n3525), .Z(n11573) );
  NANDN U5897 ( .A(x[694]), .B(y[694]), .Z(n5709) );
  NANDN U5898 ( .A(x[695]), .B(y[695]), .Z(n5708) );
  AND U5899 ( .A(n5709), .B(n5708), .Z(n11571) );
  ANDN U5900 ( .B(x[694]), .A(y[694]), .Z(n8353) );
  NANDN U5901 ( .A(y[693]), .B(x[693]), .Z(n8345) );
  NANDN U5902 ( .A(n8353), .B(n8345), .Z(n11569) );
  NANDN U5903 ( .A(x[693]), .B(y[693]), .Z(n5710) );
  ANDN U5904 ( .B(y[692]), .A(x[692]), .Z(n8341) );
  ANDN U5905 ( .B(n5710), .A(n8341), .Z(n11567) );
  ANDN U5906 ( .B(x[692]), .A(y[692]), .Z(n8347) );
  NANDN U5907 ( .A(y[691]), .B(x[691]), .Z(n8337) );
  NANDN U5908 ( .A(n8347), .B(n8337), .Z(n11565) );
  ANDN U5909 ( .B(y[690]), .A(x[690]), .Z(n8332) );
  ANDN U5910 ( .B(y[691]), .A(x[691]), .Z(n8343) );
  NOR U5911 ( .A(n8332), .B(n8343), .Z(n11563) );
  NANDN U5912 ( .A(y[689]), .B(x[689]), .Z(n8329) );
  NANDN U5913 ( .A(y[690]), .B(x[690]), .Z(n8336) );
  NAND U5914 ( .A(n8329), .B(n8336), .Z(n11561) );
  NANDN U5915 ( .A(x[688]), .B(y[688]), .Z(n8324) );
  ANDN U5916 ( .B(y[689]), .A(x[689]), .Z(n8335) );
  ANDN U5917 ( .B(n8324), .A(n8335), .Z(n11559) );
  NANDN U5918 ( .A(y[687]), .B(x[687]), .Z(n5712) );
  NANDN U5919 ( .A(y[688]), .B(x[688]), .Z(n8330) );
  NAND U5920 ( .A(n5712), .B(n8330), .Z(n11557) );
  NANDN U5921 ( .A(x[687]), .B(y[687]), .Z(n8325) );
  ANDN U5922 ( .B(y[686]), .A(x[686]), .Z(n8319) );
  ANDN U5923 ( .B(n8325), .A(n8319), .Z(n11555) );
  NANDN U5924 ( .A(y[685]), .B(x[685]), .Z(n8315) );
  NANDN U5925 ( .A(y[686]), .B(x[686]), .Z(n5711) );
  NAND U5926 ( .A(n8315), .B(n5711), .Z(n11553) );
  ANDN U5927 ( .B(y[684]), .A(x[684]), .Z(n8310) );
  ANDN U5928 ( .B(y[685]), .A(x[685]), .Z(n8320) );
  NOR U5929 ( .A(n8310), .B(n8320), .Z(n11551) );
  NANDN U5930 ( .A(y[683]), .B(x[683]), .Z(n8307) );
  NANDN U5931 ( .A(y[684]), .B(x[684]), .Z(n8314) );
  NAND U5932 ( .A(n8307), .B(n8314), .Z(n11549) );
  NANDN U5933 ( .A(x[682]), .B(y[682]), .Z(n8302) );
  ANDN U5934 ( .B(y[683]), .A(x[683]), .Z(n8313) );
  ANDN U5935 ( .B(n8302), .A(n8313), .Z(n11547) );
  NANDN U5936 ( .A(y[681]), .B(x[681]), .Z(n5714) );
  NANDN U5937 ( .A(y[682]), .B(x[682]), .Z(n8308) );
  NAND U5938 ( .A(n5714), .B(n8308), .Z(n11545) );
  NANDN U5939 ( .A(x[681]), .B(y[681]), .Z(n8303) );
  ANDN U5940 ( .B(y[680]), .A(x[680]), .Z(n8297) );
  ANDN U5941 ( .B(n8303), .A(n8297), .Z(n11543) );
  NANDN U5942 ( .A(y[679]), .B(x[679]), .Z(n8293) );
  NANDN U5943 ( .A(y[680]), .B(x[680]), .Z(n5713) );
  NAND U5944 ( .A(n8293), .B(n5713), .Z(n11541) );
  ANDN U5945 ( .B(y[678]), .A(x[678]), .Z(n8288) );
  ANDN U5946 ( .B(y[679]), .A(x[679]), .Z(n8298) );
  NOR U5947 ( .A(n8288), .B(n8298), .Z(n11539) );
  NANDN U5948 ( .A(y[677]), .B(x[677]), .Z(n8285) );
  NANDN U5949 ( .A(y[678]), .B(x[678]), .Z(n8292) );
  NAND U5950 ( .A(n8285), .B(n8292), .Z(n11537) );
  NANDN U5951 ( .A(x[676]), .B(y[676]), .Z(n8280) );
  ANDN U5952 ( .B(y[677]), .A(x[677]), .Z(n8291) );
  ANDN U5953 ( .B(n8280), .A(n8291), .Z(n11535) );
  NANDN U5954 ( .A(y[675]), .B(x[675]), .Z(n5716) );
  NANDN U5955 ( .A(y[676]), .B(x[676]), .Z(n8286) );
  NAND U5956 ( .A(n5716), .B(n8286), .Z(n11533) );
  NANDN U5957 ( .A(x[675]), .B(y[675]), .Z(n8281) );
  ANDN U5958 ( .B(y[674]), .A(x[674]), .Z(n8275) );
  ANDN U5959 ( .B(n8281), .A(n8275), .Z(n11531) );
  NANDN U5960 ( .A(y[673]), .B(x[673]), .Z(n8271) );
  NANDN U5961 ( .A(y[674]), .B(x[674]), .Z(n5715) );
  NAND U5962 ( .A(n8271), .B(n5715), .Z(n11529) );
  ANDN U5963 ( .B(y[672]), .A(x[672]), .Z(n8266) );
  ANDN U5964 ( .B(y[673]), .A(x[673]), .Z(n8276) );
  NOR U5965 ( .A(n8266), .B(n8276), .Z(n11527) );
  NANDN U5966 ( .A(y[671]), .B(x[671]), .Z(n8263) );
  NANDN U5967 ( .A(y[672]), .B(x[672]), .Z(n8270) );
  NAND U5968 ( .A(n8263), .B(n8270), .Z(n11525) );
  NANDN U5969 ( .A(x[670]), .B(y[670]), .Z(n8258) );
  ANDN U5970 ( .B(y[671]), .A(x[671]), .Z(n8269) );
  ANDN U5971 ( .B(n8258), .A(n8269), .Z(n11523) );
  NANDN U5972 ( .A(y[669]), .B(x[669]), .Z(n5718) );
  NANDN U5973 ( .A(y[670]), .B(x[670]), .Z(n8264) );
  NAND U5974 ( .A(n5718), .B(n8264), .Z(n11521) );
  NANDN U5975 ( .A(x[669]), .B(y[669]), .Z(n8259) );
  ANDN U5976 ( .B(y[668]), .A(x[668]), .Z(n8253) );
  ANDN U5977 ( .B(n8259), .A(n8253), .Z(n11519) );
  NANDN U5978 ( .A(y[667]), .B(x[667]), .Z(n8249) );
  NANDN U5979 ( .A(y[668]), .B(x[668]), .Z(n5717) );
  NAND U5980 ( .A(n8249), .B(n5717), .Z(n11517) );
  ANDN U5981 ( .B(y[666]), .A(x[666]), .Z(n8244) );
  ANDN U5982 ( .B(y[667]), .A(x[667]), .Z(n8254) );
  NOR U5983 ( .A(n8244), .B(n8254), .Z(n11515) );
  NANDN U5984 ( .A(y[665]), .B(x[665]), .Z(n8241) );
  NANDN U5985 ( .A(y[666]), .B(x[666]), .Z(n8248) );
  NAND U5986 ( .A(n8241), .B(n8248), .Z(n11513) );
  NANDN U5987 ( .A(x[664]), .B(y[664]), .Z(n8236) );
  ANDN U5988 ( .B(y[665]), .A(x[665]), .Z(n8247) );
  ANDN U5989 ( .B(n8236), .A(n8247), .Z(n11511) );
  NANDN U5990 ( .A(y[663]), .B(x[663]), .Z(n5720) );
  NANDN U5991 ( .A(y[664]), .B(x[664]), .Z(n8242) );
  NAND U5992 ( .A(n5720), .B(n8242), .Z(n11509) );
  NANDN U5993 ( .A(x[663]), .B(y[663]), .Z(n8237) );
  ANDN U5994 ( .B(y[662]), .A(x[662]), .Z(n8232) );
  ANDN U5995 ( .B(n8237), .A(n8232), .Z(n11507) );
  NANDN U5996 ( .A(y[661]), .B(x[661]), .Z(n8231) );
  NANDN U5997 ( .A(y[662]), .B(x[662]), .Z(n5719) );
  NAND U5998 ( .A(n8231), .B(n5719), .Z(n11505) );
  ANDN U5999 ( .B(y[660]), .A(x[660]), .Z(n8228) );
  ANDN U6000 ( .B(y[661]), .A(x[661]), .Z(n8233) );
  NOR U6001 ( .A(n8228), .B(n8233), .Z(n11503) );
  NANDN U6002 ( .A(y[659]), .B(x[659]), .Z(n8226) );
  NANDN U6003 ( .A(y[660]), .B(x[660]), .Z(n8230) );
  NAND U6004 ( .A(n8226), .B(n8230), .Z(n11501) );
  ANDN U6005 ( .B(y[658]), .A(x[658]), .Z(n8224) );
  ANDN U6006 ( .B(y[659]), .A(x[659]), .Z(n8229) );
  NOR U6007 ( .A(n8224), .B(n8229), .Z(n11499) );
  NANDN U6008 ( .A(y[657]), .B(x[657]), .Z(n8223) );
  NANDN U6009 ( .A(y[658]), .B(x[658]), .Z(n8227) );
  NAND U6010 ( .A(n8223), .B(n8227), .Z(n11497) );
  ANDN U6011 ( .B(y[656]), .A(x[656]), .Z(n8222) );
  ANDN U6012 ( .B(y[657]), .A(x[657]), .Z(n8225) );
  NOR U6013 ( .A(n8222), .B(n8225), .Z(n11495) );
  NANDN U6014 ( .A(y[653]), .B(x[653]), .Z(n3527) );
  NANDN U6015 ( .A(y[654]), .B(x[654]), .Z(n3526) );
  AND U6016 ( .A(n3527), .B(n3526), .Z(n11488) );
  NANDN U6017 ( .A(x[653]), .B(y[653]), .Z(n3529) );
  NANDN U6018 ( .A(x[652]), .B(y[652]), .Z(n3528) );
  NAND U6019 ( .A(n3529), .B(n3528), .Z(n11486) );
  NANDN U6020 ( .A(y[651]), .B(x[651]), .Z(n3531) );
  NANDN U6021 ( .A(y[652]), .B(x[652]), .Z(n3530) );
  AND U6022 ( .A(n3531), .B(n3530), .Z(n11485) );
  NANDN U6023 ( .A(x[651]), .B(y[651]), .Z(n3533) );
  NANDN U6024 ( .A(x[650]), .B(y[650]), .Z(n3532) );
  NAND U6025 ( .A(n3533), .B(n3532), .Z(n11483) );
  NANDN U6026 ( .A(y[647]), .B(x[647]), .Z(n3535) );
  NANDN U6027 ( .A(y[648]), .B(x[648]), .Z(n3534) );
  AND U6028 ( .A(n3535), .B(n3534), .Z(n11476) );
  NANDN U6029 ( .A(x[646]), .B(y[646]), .Z(n3536) );
  ANDN U6030 ( .B(y[647]), .A(x[647]), .Z(n8220) );
  ANDN U6031 ( .B(n3536), .A(n8220), .Z(n11475) );
  ANDN U6032 ( .B(x[645]), .A(y[645]), .Z(n8217) );
  NANDN U6033 ( .A(y[646]), .B(x[646]), .Z(n3537) );
  NANDN U6034 ( .A(n8217), .B(n3537), .Z(n11473) );
  NANDN U6035 ( .A(x[644]), .B(y[644]), .Z(n8215) );
  NANDN U6036 ( .A(x[645]), .B(y[645]), .Z(n8219) );
  AND U6037 ( .A(n8215), .B(n8219), .Z(n11471) );
  ANDN U6038 ( .B(x[643]), .A(y[643]), .Z(n8213) );
  ANDN U6039 ( .B(x[644]), .A(y[644]), .Z(n8218) );
  OR U6040 ( .A(n8213), .B(n8218), .Z(n11469) );
  NANDN U6041 ( .A(x[642]), .B(y[642]), .Z(n5722) );
  NANDN U6042 ( .A(x[643]), .B(y[643]), .Z(n8216) );
  AND U6043 ( .A(n5722), .B(n8216), .Z(n11467) );
  ANDN U6044 ( .B(x[641]), .A(y[641]), .Z(n8205) );
  XNOR U6045 ( .A(y[642]), .B(x[642]), .Z(n3538) );
  NANDN U6046 ( .A(n8205), .B(n3538), .Z(n11465) );
  NANDN U6047 ( .A(x[640]), .B(y[640]), .Z(n8201) );
  NANDN U6048 ( .A(x[641]), .B(y[641]), .Z(n5721) );
  AND U6049 ( .A(n8201), .B(n5721), .Z(n11463) );
  ANDN U6050 ( .B(x[639]), .A(y[639]), .Z(n8196) );
  ANDN U6051 ( .B(x[640]), .A(y[640]), .Z(n8206) );
  OR U6052 ( .A(n8196), .B(n8206), .Z(n11461) );
  NANDN U6053 ( .A(x[638]), .B(y[638]), .Z(n8193) );
  NANDN U6054 ( .A(x[639]), .B(y[639]), .Z(n8200) );
  AND U6055 ( .A(n8193), .B(n8200), .Z(n11459) );
  ANDN U6056 ( .B(x[637]), .A(y[637]), .Z(n8191) );
  ANDN U6057 ( .B(x[638]), .A(y[638]), .Z(n8199) );
  OR U6058 ( .A(n8191), .B(n8199), .Z(n11457) );
  NANDN U6059 ( .A(x[636]), .B(y[636]), .Z(n5724) );
  NANDN U6060 ( .A(x[637]), .B(y[637]), .Z(n8194) );
  AND U6061 ( .A(n5724), .B(n8194), .Z(n11455) );
  ANDN U6062 ( .B(x[635]), .A(y[635]), .Z(n8183) );
  ANDN U6063 ( .B(x[636]), .A(y[636]), .Z(n8188) );
  OR U6064 ( .A(n8183), .B(n8188), .Z(n11453) );
  NANDN U6065 ( .A(x[634]), .B(y[634]), .Z(n8179) );
  NANDN U6066 ( .A(x[635]), .B(y[635]), .Z(n5723) );
  AND U6067 ( .A(n8179), .B(n5723), .Z(n11451) );
  ANDN U6068 ( .B(x[633]), .A(y[633]), .Z(n8174) );
  ANDN U6069 ( .B(x[634]), .A(y[634]), .Z(n8184) );
  OR U6070 ( .A(n8174), .B(n8184), .Z(n11449) );
  NANDN U6071 ( .A(x[632]), .B(y[632]), .Z(n8171) );
  NANDN U6072 ( .A(x[633]), .B(y[633]), .Z(n8178) );
  AND U6073 ( .A(n8171), .B(n8178), .Z(n11447) );
  ANDN U6074 ( .B(x[631]), .A(y[631]), .Z(n8169) );
  XNOR U6075 ( .A(y[632]), .B(x[632]), .Z(n3539) );
  NANDN U6076 ( .A(n8169), .B(n3539), .Z(n11445) );
  NANDN U6077 ( .A(x[630]), .B(y[630]), .Z(n5726) );
  NANDN U6078 ( .A(x[631]), .B(y[631]), .Z(n8172) );
  AND U6079 ( .A(n5726), .B(n8172), .Z(n11443) );
  ANDN U6080 ( .B(x[629]), .A(y[629]), .Z(n8161) );
  ANDN U6081 ( .B(x[630]), .A(y[630]), .Z(n8166) );
  OR U6082 ( .A(n8161), .B(n8166), .Z(n11441) );
  NANDN U6083 ( .A(x[628]), .B(y[628]), .Z(n8157) );
  NANDN U6084 ( .A(x[629]), .B(y[629]), .Z(n5725) );
  AND U6085 ( .A(n8157), .B(n5725), .Z(n11439) );
  ANDN U6086 ( .B(x[627]), .A(y[627]), .Z(n8152) );
  ANDN U6087 ( .B(x[628]), .A(y[628]), .Z(n8162) );
  OR U6088 ( .A(n8152), .B(n8162), .Z(n11437) );
  NANDN U6089 ( .A(x[626]), .B(y[626]), .Z(n8149) );
  NANDN U6090 ( .A(x[627]), .B(y[627]), .Z(n8156) );
  AND U6091 ( .A(n8149), .B(n8156), .Z(n11435) );
  ANDN U6092 ( .B(x[625]), .A(y[625]), .Z(n8147) );
  ANDN U6093 ( .B(x[626]), .A(y[626]), .Z(n8155) );
  OR U6094 ( .A(n8147), .B(n8155), .Z(n11433) );
  NANDN U6095 ( .A(x[624]), .B(y[624]), .Z(n5728) );
  NANDN U6096 ( .A(x[625]), .B(y[625]), .Z(n8150) );
  AND U6097 ( .A(n5728), .B(n8150), .Z(n11431) );
  ANDN U6098 ( .B(x[623]), .A(y[623]), .Z(n8139) );
  XNOR U6099 ( .A(y[624]), .B(x[624]), .Z(n3540) );
  NANDN U6100 ( .A(n8139), .B(n3540), .Z(n11429) );
  NANDN U6101 ( .A(x[622]), .B(y[622]), .Z(n8135) );
  NANDN U6102 ( .A(x[623]), .B(y[623]), .Z(n5727) );
  AND U6103 ( .A(n8135), .B(n5727), .Z(n11427) );
  ANDN U6104 ( .B(x[621]), .A(y[621]), .Z(n8130) );
  ANDN U6105 ( .B(x[622]), .A(y[622]), .Z(n8140) );
  OR U6106 ( .A(n8130), .B(n8140), .Z(n11425) );
  NANDN U6107 ( .A(x[620]), .B(y[620]), .Z(n8127) );
  NANDN U6108 ( .A(x[621]), .B(y[621]), .Z(n8134) );
  AND U6109 ( .A(n8127), .B(n8134), .Z(n11423) );
  ANDN U6110 ( .B(x[619]), .A(y[619]), .Z(n8125) );
  ANDN U6111 ( .B(x[620]), .A(y[620]), .Z(n8133) );
  OR U6112 ( .A(n8125), .B(n8133), .Z(n11421) );
  NANDN U6113 ( .A(x[618]), .B(y[618]), .Z(n5730) );
  NANDN U6114 ( .A(x[619]), .B(y[619]), .Z(n8128) );
  AND U6115 ( .A(n5730), .B(n8128), .Z(n11419) );
  ANDN U6116 ( .B(x[617]), .A(y[617]), .Z(n8117) );
  ANDN U6117 ( .B(x[618]), .A(y[618]), .Z(n8122) );
  OR U6118 ( .A(n8117), .B(n8122), .Z(n11417) );
  NANDN U6119 ( .A(x[616]), .B(y[616]), .Z(n8113) );
  NANDN U6120 ( .A(x[617]), .B(y[617]), .Z(n5729) );
  AND U6121 ( .A(n8113), .B(n5729), .Z(n11415) );
  ANDN U6122 ( .B(x[615]), .A(y[615]), .Z(n8108) );
  ANDN U6123 ( .B(x[616]), .A(y[616]), .Z(n8118) );
  OR U6124 ( .A(n8108), .B(n8118), .Z(n11413) );
  NANDN U6125 ( .A(x[614]), .B(y[614]), .Z(n8105) );
  NANDN U6126 ( .A(x[615]), .B(y[615]), .Z(n8112) );
  AND U6127 ( .A(n8105), .B(n8112), .Z(n11411) );
  ANDN U6128 ( .B(x[613]), .A(y[613]), .Z(n8103) );
  ANDN U6129 ( .B(x[614]), .A(y[614]), .Z(n8111) );
  OR U6130 ( .A(n8103), .B(n8111), .Z(n11409) );
  NANDN U6131 ( .A(x[612]), .B(y[612]), .Z(n5732) );
  NANDN U6132 ( .A(x[613]), .B(y[613]), .Z(n8106) );
  AND U6133 ( .A(n5732), .B(n8106), .Z(n11407) );
  ANDN U6134 ( .B(x[611]), .A(y[611]), .Z(n8095) );
  ANDN U6135 ( .B(x[612]), .A(y[612]), .Z(n8100) );
  OR U6136 ( .A(n8095), .B(n8100), .Z(n11405) );
  NANDN U6137 ( .A(x[610]), .B(y[610]), .Z(n8091) );
  NANDN U6138 ( .A(x[611]), .B(y[611]), .Z(n5731) );
  AND U6139 ( .A(n8091), .B(n5731), .Z(n11403) );
  ANDN U6140 ( .B(x[609]), .A(y[609]), .Z(n8086) );
  ANDN U6141 ( .B(x[610]), .A(y[610]), .Z(n8096) );
  OR U6142 ( .A(n8086), .B(n8096), .Z(n11401) );
  NANDN U6143 ( .A(x[608]), .B(y[608]), .Z(n8083) );
  NANDN U6144 ( .A(x[609]), .B(y[609]), .Z(n8090) );
  AND U6145 ( .A(n8083), .B(n8090), .Z(n11399) );
  ANDN U6146 ( .B(x[607]), .A(y[607]), .Z(n8081) );
  ANDN U6147 ( .B(x[608]), .A(y[608]), .Z(n8089) );
  OR U6148 ( .A(n8081), .B(n8089), .Z(n11397) );
  NANDN U6149 ( .A(x[606]), .B(y[606]), .Z(n5734) );
  NANDN U6150 ( .A(x[607]), .B(y[607]), .Z(n8084) );
  AND U6151 ( .A(n5734), .B(n8084), .Z(n11395) );
  ANDN U6152 ( .B(x[605]), .A(y[605]), .Z(n8073) );
  ANDN U6153 ( .B(x[606]), .A(y[606]), .Z(n8078) );
  OR U6154 ( .A(n8073), .B(n8078), .Z(n11393) );
  NANDN U6155 ( .A(x[604]), .B(y[604]), .Z(n8069) );
  NANDN U6156 ( .A(x[605]), .B(y[605]), .Z(n5733) );
  AND U6157 ( .A(n8069), .B(n5733), .Z(n11391) );
  ANDN U6158 ( .B(x[603]), .A(y[603]), .Z(n8064) );
  ANDN U6159 ( .B(x[604]), .A(y[604]), .Z(n8074) );
  OR U6160 ( .A(n8064), .B(n8074), .Z(n11389) );
  NANDN U6161 ( .A(x[602]), .B(y[602]), .Z(n8061) );
  NANDN U6162 ( .A(x[603]), .B(y[603]), .Z(n8068) );
  AND U6163 ( .A(n8061), .B(n8068), .Z(n11387) );
  ANDN U6164 ( .B(x[601]), .A(y[601]), .Z(n8059) );
  XNOR U6165 ( .A(y[602]), .B(x[602]), .Z(n3541) );
  NANDN U6166 ( .A(n8059), .B(n3541), .Z(n11385) );
  NANDN U6167 ( .A(x[600]), .B(y[600]), .Z(n5736) );
  NANDN U6168 ( .A(x[601]), .B(y[601]), .Z(n8062) );
  AND U6169 ( .A(n5736), .B(n8062), .Z(n11383) );
  ANDN U6170 ( .B(x[599]), .A(y[599]), .Z(n8051) );
  XNOR U6171 ( .A(y[600]), .B(x[600]), .Z(n3542) );
  NANDN U6172 ( .A(n8051), .B(n3542), .Z(n11381) );
  NANDN U6173 ( .A(x[598]), .B(y[598]), .Z(n8047) );
  NANDN U6174 ( .A(x[599]), .B(y[599]), .Z(n5735) );
  AND U6175 ( .A(n8047), .B(n5735), .Z(n11379) );
  ANDN U6176 ( .B(x[597]), .A(y[597]), .Z(n8042) );
  ANDN U6177 ( .B(x[598]), .A(y[598]), .Z(n8052) );
  OR U6178 ( .A(n8042), .B(n8052), .Z(n11377) );
  NANDN U6179 ( .A(x[596]), .B(y[596]), .Z(n8039) );
  NANDN U6180 ( .A(x[597]), .B(y[597]), .Z(n8046) );
  AND U6181 ( .A(n8039), .B(n8046), .Z(n11375) );
  ANDN U6182 ( .B(x[595]), .A(y[595]), .Z(n8037) );
  XNOR U6183 ( .A(y[596]), .B(x[596]), .Z(n3543) );
  NANDN U6184 ( .A(n8037), .B(n3543), .Z(n11373) );
  NANDN U6185 ( .A(x[594]), .B(y[594]), .Z(n5738) );
  NANDN U6186 ( .A(x[595]), .B(y[595]), .Z(n8040) );
  AND U6187 ( .A(n5738), .B(n8040), .Z(n11371) );
  ANDN U6188 ( .B(x[593]), .A(y[593]), .Z(n8029) );
  XNOR U6189 ( .A(y[594]), .B(x[594]), .Z(n3544) );
  NANDN U6190 ( .A(n8029), .B(n3544), .Z(n11369) );
  NANDN U6191 ( .A(x[592]), .B(y[592]), .Z(n8025) );
  NANDN U6192 ( .A(x[593]), .B(y[593]), .Z(n5737) );
  AND U6193 ( .A(n8025), .B(n5737), .Z(n11367) );
  ANDN U6194 ( .B(x[591]), .A(y[591]), .Z(n8020) );
  ANDN U6195 ( .B(x[592]), .A(y[592]), .Z(n8030) );
  OR U6196 ( .A(n8020), .B(n8030), .Z(n11365) );
  NANDN U6197 ( .A(x[590]), .B(y[590]), .Z(n8017) );
  NANDN U6198 ( .A(x[591]), .B(y[591]), .Z(n8024) );
  AND U6199 ( .A(n8017), .B(n8024), .Z(n11363) );
  ANDN U6200 ( .B(x[589]), .A(y[589]), .Z(n8015) );
  ANDN U6201 ( .B(x[590]), .A(y[590]), .Z(n8023) );
  OR U6202 ( .A(n8015), .B(n8023), .Z(n11361) );
  NANDN U6203 ( .A(x[588]), .B(y[588]), .Z(n5740) );
  NANDN U6204 ( .A(x[589]), .B(y[589]), .Z(n8018) );
  AND U6205 ( .A(n5740), .B(n8018), .Z(n11359) );
  ANDN U6206 ( .B(x[587]), .A(y[587]), .Z(n8007) );
  ANDN U6207 ( .B(x[588]), .A(y[588]), .Z(n8012) );
  OR U6208 ( .A(n8007), .B(n8012), .Z(n11357) );
  NANDN U6209 ( .A(x[586]), .B(y[586]), .Z(n8003) );
  NANDN U6210 ( .A(x[587]), .B(y[587]), .Z(n5739) );
  AND U6211 ( .A(n8003), .B(n5739), .Z(n11355) );
  ANDN U6212 ( .B(x[585]), .A(y[585]), .Z(n7998) );
  ANDN U6213 ( .B(x[586]), .A(y[586]), .Z(n8008) );
  OR U6214 ( .A(n7998), .B(n8008), .Z(n11353) );
  NANDN U6215 ( .A(x[584]), .B(y[584]), .Z(n7995) );
  NANDN U6216 ( .A(x[585]), .B(y[585]), .Z(n8002) );
  AND U6217 ( .A(n7995), .B(n8002), .Z(n11351) );
  ANDN U6218 ( .B(x[583]), .A(y[583]), .Z(n7993) );
  ANDN U6219 ( .B(x[584]), .A(y[584]), .Z(n8001) );
  OR U6220 ( .A(n7993), .B(n8001), .Z(n11349) );
  NANDN U6221 ( .A(x[582]), .B(y[582]), .Z(n5742) );
  NANDN U6222 ( .A(x[583]), .B(y[583]), .Z(n7996) );
  AND U6223 ( .A(n5742), .B(n7996), .Z(n11347) );
  ANDN U6224 ( .B(x[581]), .A(y[581]), .Z(n7985) );
  ANDN U6225 ( .B(x[582]), .A(y[582]), .Z(n7990) );
  OR U6226 ( .A(n7985), .B(n7990), .Z(n11345) );
  NANDN U6227 ( .A(x[580]), .B(y[580]), .Z(n7981) );
  NANDN U6228 ( .A(x[581]), .B(y[581]), .Z(n5741) );
  AND U6229 ( .A(n7981), .B(n5741), .Z(n11343) );
  ANDN U6230 ( .B(x[579]), .A(y[579]), .Z(n7976) );
  ANDN U6231 ( .B(x[580]), .A(y[580]), .Z(n7986) );
  OR U6232 ( .A(n7976), .B(n7986), .Z(n11341) );
  NANDN U6233 ( .A(x[578]), .B(y[578]), .Z(n7973) );
  NANDN U6234 ( .A(x[579]), .B(y[579]), .Z(n7980) );
  AND U6235 ( .A(n7973), .B(n7980), .Z(n11339) );
  ANDN U6236 ( .B(x[577]), .A(y[577]), .Z(n7971) );
  ANDN U6237 ( .B(x[578]), .A(y[578]), .Z(n7979) );
  OR U6238 ( .A(n7971), .B(n7979), .Z(n11337) );
  NANDN U6239 ( .A(x[576]), .B(y[576]), .Z(n5744) );
  NANDN U6240 ( .A(x[577]), .B(y[577]), .Z(n7974) );
  AND U6241 ( .A(n5744), .B(n7974), .Z(n11335) );
  ANDN U6242 ( .B(x[575]), .A(y[575]), .Z(n7963) );
  XNOR U6243 ( .A(y[576]), .B(x[576]), .Z(n3545) );
  NANDN U6244 ( .A(n7963), .B(n3545), .Z(n11333) );
  NANDN U6245 ( .A(x[574]), .B(y[574]), .Z(n7959) );
  NANDN U6246 ( .A(x[575]), .B(y[575]), .Z(n5743) );
  AND U6247 ( .A(n7959), .B(n5743), .Z(n11331) );
  ANDN U6248 ( .B(x[573]), .A(y[573]), .Z(n7954) );
  ANDN U6249 ( .B(x[574]), .A(y[574]), .Z(n7964) );
  OR U6250 ( .A(n7954), .B(n7964), .Z(n11329) );
  NANDN U6251 ( .A(x[572]), .B(y[572]), .Z(n7951) );
  NANDN U6252 ( .A(x[573]), .B(y[573]), .Z(n7958) );
  AND U6253 ( .A(n7951), .B(n7958), .Z(n11327) );
  ANDN U6254 ( .B(x[571]), .A(y[571]), .Z(n7949) );
  XNOR U6255 ( .A(y[572]), .B(x[572]), .Z(n3546) );
  NANDN U6256 ( .A(n7949), .B(n3546), .Z(n11325) );
  NANDN U6257 ( .A(x[570]), .B(y[570]), .Z(n5746) );
  NANDN U6258 ( .A(x[571]), .B(y[571]), .Z(n7952) );
  AND U6259 ( .A(n5746), .B(n7952), .Z(n11323) );
  ANDN U6260 ( .B(x[569]), .A(y[569]), .Z(n7941) );
  XNOR U6261 ( .A(y[570]), .B(x[570]), .Z(n3547) );
  NANDN U6262 ( .A(n7941), .B(n3547), .Z(n11321) );
  NANDN U6263 ( .A(x[568]), .B(y[568]), .Z(n7937) );
  NANDN U6264 ( .A(x[569]), .B(y[569]), .Z(n5745) );
  AND U6265 ( .A(n7937), .B(n5745), .Z(n11319) );
  ANDN U6266 ( .B(x[567]), .A(y[567]), .Z(n7932) );
  ANDN U6267 ( .B(x[568]), .A(y[568]), .Z(n7942) );
  OR U6268 ( .A(n7932), .B(n7942), .Z(n11317) );
  NANDN U6269 ( .A(x[566]), .B(y[566]), .Z(n7929) );
  NANDN U6270 ( .A(x[567]), .B(y[567]), .Z(n7936) );
  AND U6271 ( .A(n7929), .B(n7936), .Z(n11315) );
  ANDN U6272 ( .B(x[565]), .A(y[565]), .Z(n7927) );
  XNOR U6273 ( .A(y[566]), .B(x[566]), .Z(n3548) );
  NANDN U6274 ( .A(n7927), .B(n3548), .Z(n11313) );
  NANDN U6275 ( .A(x[564]), .B(y[564]), .Z(n5748) );
  NANDN U6276 ( .A(x[565]), .B(y[565]), .Z(n7930) );
  AND U6277 ( .A(n5748), .B(n7930), .Z(n11311) );
  ANDN U6278 ( .B(x[563]), .A(y[563]), .Z(n7919) );
  ANDN U6279 ( .B(x[564]), .A(y[564]), .Z(n7924) );
  OR U6280 ( .A(n7919), .B(n7924), .Z(n11309) );
  NANDN U6281 ( .A(x[562]), .B(y[562]), .Z(n7915) );
  NANDN U6282 ( .A(x[563]), .B(y[563]), .Z(n5747) );
  AND U6283 ( .A(n7915), .B(n5747), .Z(n11307) );
  ANDN U6284 ( .B(x[561]), .A(y[561]), .Z(n7910) );
  ANDN U6285 ( .B(x[562]), .A(y[562]), .Z(n7920) );
  OR U6286 ( .A(n7910), .B(n7920), .Z(n11305) );
  NANDN U6287 ( .A(x[560]), .B(y[560]), .Z(n7907) );
  NANDN U6288 ( .A(x[561]), .B(y[561]), .Z(n7914) );
  AND U6289 ( .A(n7907), .B(n7914), .Z(n11303) );
  ANDN U6290 ( .B(x[559]), .A(y[559]), .Z(n7905) );
  ANDN U6291 ( .B(x[560]), .A(y[560]), .Z(n7913) );
  OR U6292 ( .A(n7905), .B(n7913), .Z(n11301) );
  NANDN U6293 ( .A(x[558]), .B(y[558]), .Z(n5750) );
  NANDN U6294 ( .A(x[559]), .B(y[559]), .Z(n7908) );
  AND U6295 ( .A(n5750), .B(n7908), .Z(n11299) );
  ANDN U6296 ( .B(x[557]), .A(y[557]), .Z(n7897) );
  ANDN U6297 ( .B(x[558]), .A(y[558]), .Z(n7902) );
  OR U6298 ( .A(n7897), .B(n7902), .Z(n11297) );
  NANDN U6299 ( .A(x[556]), .B(y[556]), .Z(n7893) );
  NANDN U6300 ( .A(x[557]), .B(y[557]), .Z(n5749) );
  AND U6301 ( .A(n7893), .B(n5749), .Z(n11295) );
  ANDN U6302 ( .B(x[555]), .A(y[555]), .Z(n7888) );
  ANDN U6303 ( .B(x[556]), .A(y[556]), .Z(n7898) );
  OR U6304 ( .A(n7888), .B(n7898), .Z(n11293) );
  NANDN U6305 ( .A(x[554]), .B(y[554]), .Z(n7885) );
  NANDN U6306 ( .A(x[555]), .B(y[555]), .Z(n7892) );
  AND U6307 ( .A(n7885), .B(n7892), .Z(n11291) );
  ANDN U6308 ( .B(x[553]), .A(y[553]), .Z(n7883) );
  ANDN U6309 ( .B(x[554]), .A(y[554]), .Z(n7891) );
  OR U6310 ( .A(n7883), .B(n7891), .Z(n11289) );
  NANDN U6311 ( .A(x[552]), .B(y[552]), .Z(n5752) );
  NANDN U6312 ( .A(x[553]), .B(y[553]), .Z(n7886) );
  AND U6313 ( .A(n5752), .B(n7886), .Z(n11287) );
  ANDN U6314 ( .B(x[551]), .A(y[551]), .Z(n7875) );
  ANDN U6315 ( .B(x[552]), .A(y[552]), .Z(n7880) );
  OR U6316 ( .A(n7875), .B(n7880), .Z(n11285) );
  NANDN U6317 ( .A(x[550]), .B(y[550]), .Z(n7871) );
  NANDN U6318 ( .A(x[551]), .B(y[551]), .Z(n5751) );
  AND U6319 ( .A(n7871), .B(n5751), .Z(n11283) );
  ANDN U6320 ( .B(x[549]), .A(y[549]), .Z(n7866) );
  ANDN U6321 ( .B(x[550]), .A(y[550]), .Z(n7876) );
  OR U6322 ( .A(n7866), .B(n7876), .Z(n11281) );
  NANDN U6323 ( .A(x[548]), .B(y[548]), .Z(n7863) );
  NANDN U6324 ( .A(x[549]), .B(y[549]), .Z(n7870) );
  AND U6325 ( .A(n7863), .B(n7870), .Z(n11279) );
  ANDN U6326 ( .B(x[547]), .A(y[547]), .Z(n7861) );
  XNOR U6327 ( .A(y[548]), .B(x[548]), .Z(n3549) );
  NANDN U6328 ( .A(n7861), .B(n3549), .Z(n11277) );
  NANDN U6329 ( .A(x[546]), .B(y[546]), .Z(n5754) );
  NANDN U6330 ( .A(x[547]), .B(y[547]), .Z(n7864) );
  AND U6331 ( .A(n5754), .B(n7864), .Z(n11275) );
  ANDN U6332 ( .B(x[545]), .A(y[545]), .Z(n7853) );
  ANDN U6333 ( .B(x[546]), .A(y[546]), .Z(n7858) );
  OR U6334 ( .A(n7853), .B(n7858), .Z(n11273) );
  NANDN U6335 ( .A(x[544]), .B(y[544]), .Z(n7849) );
  NANDN U6336 ( .A(x[545]), .B(y[545]), .Z(n5753) );
  AND U6337 ( .A(n7849), .B(n5753), .Z(n11271) );
  ANDN U6338 ( .B(x[543]), .A(y[543]), .Z(n7844) );
  ANDN U6339 ( .B(x[544]), .A(y[544]), .Z(n7854) );
  OR U6340 ( .A(n7844), .B(n7854), .Z(n11269) );
  NANDN U6341 ( .A(x[542]), .B(y[542]), .Z(n7841) );
  NANDN U6342 ( .A(x[543]), .B(y[543]), .Z(n7848) );
  AND U6343 ( .A(n7841), .B(n7848), .Z(n11267) );
  ANDN U6344 ( .B(x[541]), .A(y[541]), .Z(n7839) );
  XNOR U6345 ( .A(y[542]), .B(x[542]), .Z(n3550) );
  NANDN U6346 ( .A(n7839), .B(n3550), .Z(n11265) );
  NANDN U6347 ( .A(x[540]), .B(y[540]), .Z(n5756) );
  NANDN U6348 ( .A(x[541]), .B(y[541]), .Z(n7842) );
  AND U6349 ( .A(n5756), .B(n7842), .Z(n11263) );
  ANDN U6350 ( .B(x[539]), .A(y[539]), .Z(n7831) );
  ANDN U6351 ( .B(x[540]), .A(y[540]), .Z(n7836) );
  OR U6352 ( .A(n7831), .B(n7836), .Z(n11261) );
  NANDN U6353 ( .A(x[538]), .B(y[538]), .Z(n7827) );
  NANDN U6354 ( .A(x[539]), .B(y[539]), .Z(n5755) );
  AND U6355 ( .A(n7827), .B(n5755), .Z(n11259) );
  ANDN U6356 ( .B(x[537]), .A(y[537]), .Z(n7822) );
  ANDN U6357 ( .B(x[538]), .A(y[538]), .Z(n7832) );
  OR U6358 ( .A(n7822), .B(n7832), .Z(n11257) );
  NANDN U6359 ( .A(x[536]), .B(y[536]), .Z(n7819) );
  NANDN U6360 ( .A(x[537]), .B(y[537]), .Z(n7826) );
  AND U6361 ( .A(n7819), .B(n7826), .Z(n11255) );
  ANDN U6362 ( .B(x[535]), .A(y[535]), .Z(n7817) );
  XNOR U6363 ( .A(y[536]), .B(x[536]), .Z(n3551) );
  NANDN U6364 ( .A(n7817), .B(n3551), .Z(n11253) );
  NANDN U6365 ( .A(x[534]), .B(y[534]), .Z(n3552) );
  NANDN U6366 ( .A(x[535]), .B(y[535]), .Z(n7820) );
  AND U6367 ( .A(n3552), .B(n7820), .Z(n11251) );
  ANDN U6368 ( .B(x[533]), .A(y[533]), .Z(n7809) );
  XNOR U6369 ( .A(x[534]), .B(y[534]), .Z(n5757) );
  NANDN U6370 ( .A(n7809), .B(n5757), .Z(n11249) );
  NANDN U6371 ( .A(x[532]), .B(y[532]), .Z(n7805) );
  NANDN U6372 ( .A(x[533]), .B(y[533]), .Z(n5758) );
  AND U6373 ( .A(n7805), .B(n5758), .Z(n11247) );
  ANDN U6374 ( .B(x[531]), .A(y[531]), .Z(n7800) );
  ANDN U6375 ( .B(x[532]), .A(y[532]), .Z(n7810) );
  OR U6376 ( .A(n7800), .B(n7810), .Z(n11245) );
  NANDN U6377 ( .A(x[530]), .B(y[530]), .Z(n7797) );
  NANDN U6378 ( .A(x[531]), .B(y[531]), .Z(n7804) );
  AND U6379 ( .A(n7797), .B(n7804), .Z(n11243) );
  ANDN U6380 ( .B(x[529]), .A(y[529]), .Z(n7795) );
  ANDN U6381 ( .B(x[530]), .A(y[530]), .Z(n7803) );
  OR U6382 ( .A(n7795), .B(n7803), .Z(n11241) );
  NANDN U6383 ( .A(x[528]), .B(y[528]), .Z(n5760) );
  NANDN U6384 ( .A(x[529]), .B(y[529]), .Z(n7798) );
  AND U6385 ( .A(n5760), .B(n7798), .Z(n11239) );
  ANDN U6386 ( .B(x[527]), .A(y[527]), .Z(n7787) );
  ANDN U6387 ( .B(x[528]), .A(y[528]), .Z(n7792) );
  OR U6388 ( .A(n7787), .B(n7792), .Z(n11237) );
  NANDN U6389 ( .A(x[526]), .B(y[526]), .Z(n7783) );
  NANDN U6390 ( .A(x[527]), .B(y[527]), .Z(n5759) );
  AND U6391 ( .A(n7783), .B(n5759), .Z(n11235) );
  ANDN U6392 ( .B(x[525]), .A(y[525]), .Z(n7778) );
  ANDN U6393 ( .B(x[526]), .A(y[526]), .Z(n7788) );
  OR U6394 ( .A(n7778), .B(n7788), .Z(n11233) );
  NANDN U6395 ( .A(x[524]), .B(y[524]), .Z(n7775) );
  NANDN U6396 ( .A(x[525]), .B(y[525]), .Z(n7782) );
  AND U6397 ( .A(n7775), .B(n7782), .Z(n11231) );
  ANDN U6398 ( .B(x[523]), .A(y[523]), .Z(n7773) );
  ANDN U6399 ( .B(x[524]), .A(y[524]), .Z(n7781) );
  OR U6400 ( .A(n7773), .B(n7781), .Z(n11229) );
  NANDN U6401 ( .A(x[522]), .B(y[522]), .Z(n5762) );
  NANDN U6402 ( .A(x[523]), .B(y[523]), .Z(n7776) );
  AND U6403 ( .A(n5762), .B(n7776), .Z(n11227) );
  ANDN U6404 ( .B(x[521]), .A(y[521]), .Z(n7765) );
  ANDN U6405 ( .B(x[522]), .A(y[522]), .Z(n7770) );
  OR U6406 ( .A(n7765), .B(n7770), .Z(n11225) );
  NANDN U6407 ( .A(x[520]), .B(y[520]), .Z(n7761) );
  NANDN U6408 ( .A(x[521]), .B(y[521]), .Z(n5761) );
  AND U6409 ( .A(n7761), .B(n5761), .Z(n11223) );
  ANDN U6410 ( .B(x[519]), .A(y[519]), .Z(n7756) );
  ANDN U6411 ( .B(x[520]), .A(y[520]), .Z(n7766) );
  OR U6412 ( .A(n7756), .B(n7766), .Z(n11221) );
  NANDN U6413 ( .A(x[518]), .B(y[518]), .Z(n7753) );
  NANDN U6414 ( .A(x[519]), .B(y[519]), .Z(n7760) );
  AND U6415 ( .A(n7753), .B(n7760), .Z(n11219) );
  ANDN U6416 ( .B(x[517]), .A(y[517]), .Z(n7751) );
  ANDN U6417 ( .B(x[518]), .A(y[518]), .Z(n7759) );
  OR U6418 ( .A(n7751), .B(n7759), .Z(n11217) );
  NANDN U6419 ( .A(x[516]), .B(y[516]), .Z(n5764) );
  NANDN U6420 ( .A(x[517]), .B(y[517]), .Z(n7754) );
  AND U6421 ( .A(n5764), .B(n7754), .Z(n11215) );
  ANDN U6422 ( .B(x[515]), .A(y[515]), .Z(n7743) );
  ANDN U6423 ( .B(x[516]), .A(y[516]), .Z(n7748) );
  OR U6424 ( .A(n7743), .B(n7748), .Z(n11213) );
  NANDN U6425 ( .A(x[514]), .B(y[514]), .Z(n7739) );
  NANDN U6426 ( .A(x[515]), .B(y[515]), .Z(n5763) );
  AND U6427 ( .A(n7739), .B(n5763), .Z(n11211) );
  ANDN U6428 ( .B(x[513]), .A(y[513]), .Z(n7734) );
  ANDN U6429 ( .B(x[514]), .A(y[514]), .Z(n7744) );
  OR U6430 ( .A(n7734), .B(n7744), .Z(n11209) );
  NANDN U6431 ( .A(x[512]), .B(y[512]), .Z(n7731) );
  NANDN U6432 ( .A(x[513]), .B(y[513]), .Z(n7738) );
  AND U6433 ( .A(n7731), .B(n7738), .Z(n11207) );
  ANDN U6434 ( .B(x[511]), .A(y[511]), .Z(n7729) );
  ANDN U6435 ( .B(x[512]), .A(y[512]), .Z(n7737) );
  OR U6436 ( .A(n7729), .B(n7737), .Z(n11205) );
  NANDN U6437 ( .A(x[510]), .B(y[510]), .Z(n5766) );
  NANDN U6438 ( .A(x[511]), .B(y[511]), .Z(n7732) );
  AND U6439 ( .A(n5766), .B(n7732), .Z(n11203) );
  ANDN U6440 ( .B(x[509]), .A(y[509]), .Z(n7721) );
  ANDN U6441 ( .B(x[510]), .A(y[510]), .Z(n7726) );
  OR U6442 ( .A(n7721), .B(n7726), .Z(n11201) );
  NANDN U6443 ( .A(x[508]), .B(y[508]), .Z(n7717) );
  NANDN U6444 ( .A(x[509]), .B(y[509]), .Z(n5765) );
  AND U6445 ( .A(n7717), .B(n5765), .Z(n11199) );
  ANDN U6446 ( .B(x[507]), .A(y[507]), .Z(n7712) );
  ANDN U6447 ( .B(x[508]), .A(y[508]), .Z(n7722) );
  OR U6448 ( .A(n7712), .B(n7722), .Z(n11197) );
  NANDN U6449 ( .A(x[506]), .B(y[506]), .Z(n7709) );
  NANDN U6450 ( .A(x[507]), .B(y[507]), .Z(n7716) );
  AND U6451 ( .A(n7709), .B(n7716), .Z(n11195) );
  ANDN U6452 ( .B(x[505]), .A(y[505]), .Z(n7707) );
  ANDN U6453 ( .B(x[506]), .A(y[506]), .Z(n7715) );
  OR U6454 ( .A(n7707), .B(n7715), .Z(n11193) );
  NANDN U6455 ( .A(x[504]), .B(y[504]), .Z(n5768) );
  NANDN U6456 ( .A(x[505]), .B(y[505]), .Z(n7710) );
  AND U6457 ( .A(n5768), .B(n7710), .Z(n11191) );
  ANDN U6458 ( .B(x[503]), .A(y[503]), .Z(n7699) );
  ANDN U6459 ( .B(x[504]), .A(y[504]), .Z(n7704) );
  OR U6460 ( .A(n7699), .B(n7704), .Z(n11189) );
  NANDN U6461 ( .A(x[502]), .B(y[502]), .Z(n7695) );
  NANDN U6462 ( .A(x[503]), .B(y[503]), .Z(n5767) );
  AND U6463 ( .A(n7695), .B(n5767), .Z(n11187) );
  ANDN U6464 ( .B(x[501]), .A(y[501]), .Z(n7690) );
  ANDN U6465 ( .B(x[502]), .A(y[502]), .Z(n7700) );
  OR U6466 ( .A(n7690), .B(n7700), .Z(n11185) );
  NANDN U6467 ( .A(x[500]), .B(y[500]), .Z(n7687) );
  NANDN U6468 ( .A(x[501]), .B(y[501]), .Z(n7694) );
  AND U6469 ( .A(n7687), .B(n7694), .Z(n11183) );
  ANDN U6470 ( .B(x[499]), .A(y[499]), .Z(n7685) );
  ANDN U6471 ( .B(x[500]), .A(y[500]), .Z(n7693) );
  OR U6472 ( .A(n7685), .B(n7693), .Z(n11181) );
  NANDN U6473 ( .A(x[498]), .B(y[498]), .Z(n5770) );
  NANDN U6474 ( .A(x[499]), .B(y[499]), .Z(n7688) );
  AND U6475 ( .A(n5770), .B(n7688), .Z(n11179) );
  ANDN U6476 ( .B(x[497]), .A(y[497]), .Z(n7677) );
  ANDN U6477 ( .B(x[498]), .A(y[498]), .Z(n7682) );
  OR U6478 ( .A(n7677), .B(n7682), .Z(n11177) );
  NANDN U6479 ( .A(x[496]), .B(y[496]), .Z(n7673) );
  NANDN U6480 ( .A(x[497]), .B(y[497]), .Z(n5769) );
  AND U6481 ( .A(n7673), .B(n5769), .Z(n11175) );
  ANDN U6482 ( .B(x[495]), .A(y[495]), .Z(n7668) );
  ANDN U6483 ( .B(x[496]), .A(y[496]), .Z(n7678) );
  OR U6484 ( .A(n7668), .B(n7678), .Z(n11173) );
  NANDN U6485 ( .A(x[494]), .B(y[494]), .Z(n7665) );
  NANDN U6486 ( .A(x[495]), .B(y[495]), .Z(n7672) );
  AND U6487 ( .A(n7665), .B(n7672), .Z(n11171) );
  ANDN U6488 ( .B(x[493]), .A(y[493]), .Z(n7663) );
  XNOR U6489 ( .A(y[494]), .B(x[494]), .Z(n3553) );
  NANDN U6490 ( .A(n7663), .B(n3553), .Z(n11169) );
  NANDN U6491 ( .A(x[492]), .B(y[492]), .Z(n5772) );
  NANDN U6492 ( .A(x[493]), .B(y[493]), .Z(n7666) );
  AND U6493 ( .A(n5772), .B(n7666), .Z(n11167) );
  ANDN U6494 ( .B(x[491]), .A(y[491]), .Z(n7655) );
  ANDN U6495 ( .B(x[492]), .A(y[492]), .Z(n7660) );
  OR U6496 ( .A(n7655), .B(n7660), .Z(n11165) );
  NANDN U6497 ( .A(x[490]), .B(y[490]), .Z(n7651) );
  NANDN U6498 ( .A(x[491]), .B(y[491]), .Z(n5771) );
  AND U6499 ( .A(n7651), .B(n5771), .Z(n11163) );
  ANDN U6500 ( .B(x[489]), .A(y[489]), .Z(n7646) );
  ANDN U6501 ( .B(x[490]), .A(y[490]), .Z(n7656) );
  OR U6502 ( .A(n7646), .B(n7656), .Z(n11161) );
  NANDN U6503 ( .A(x[488]), .B(y[488]), .Z(n7643) );
  NANDN U6504 ( .A(x[489]), .B(y[489]), .Z(n7650) );
  AND U6505 ( .A(n7643), .B(n7650), .Z(n11159) );
  ANDN U6506 ( .B(x[487]), .A(y[487]), .Z(n7641) );
  XNOR U6507 ( .A(y[488]), .B(x[488]), .Z(n3554) );
  NANDN U6508 ( .A(n7641), .B(n3554), .Z(n11157) );
  NANDN U6509 ( .A(x[486]), .B(y[486]), .Z(n5774) );
  NANDN U6510 ( .A(x[487]), .B(y[487]), .Z(n7644) );
  AND U6511 ( .A(n5774), .B(n7644), .Z(n11155) );
  ANDN U6512 ( .B(x[485]), .A(y[485]), .Z(n7633) );
  ANDN U6513 ( .B(x[486]), .A(y[486]), .Z(n7638) );
  OR U6514 ( .A(n7633), .B(n7638), .Z(n11153) );
  NANDN U6515 ( .A(x[484]), .B(y[484]), .Z(n7629) );
  NANDN U6516 ( .A(x[485]), .B(y[485]), .Z(n5773) );
  AND U6517 ( .A(n7629), .B(n5773), .Z(n11151) );
  ANDN U6518 ( .B(x[483]), .A(y[483]), .Z(n7624) );
  ANDN U6519 ( .B(x[484]), .A(y[484]), .Z(n7634) );
  OR U6520 ( .A(n7624), .B(n7634), .Z(n11149) );
  NANDN U6521 ( .A(x[482]), .B(y[482]), .Z(n7621) );
  NANDN U6522 ( .A(x[483]), .B(y[483]), .Z(n7628) );
  AND U6523 ( .A(n7621), .B(n7628), .Z(n11147) );
  ANDN U6524 ( .B(x[481]), .A(y[481]), .Z(n7619) );
  XNOR U6525 ( .A(y[482]), .B(x[482]), .Z(n3555) );
  NANDN U6526 ( .A(n7619), .B(n3555), .Z(n11145) );
  NANDN U6527 ( .A(x[480]), .B(y[480]), .Z(n5776) );
  NANDN U6528 ( .A(x[481]), .B(y[481]), .Z(n7622) );
  AND U6529 ( .A(n5776), .B(n7622), .Z(n11143) );
  ANDN U6530 ( .B(x[479]), .A(y[479]), .Z(n7611) );
  XNOR U6531 ( .A(y[480]), .B(x[480]), .Z(n3556) );
  NANDN U6532 ( .A(n7611), .B(n3556), .Z(n11141) );
  NANDN U6533 ( .A(x[478]), .B(y[478]), .Z(n7607) );
  NANDN U6534 ( .A(x[479]), .B(y[479]), .Z(n5775) );
  AND U6535 ( .A(n7607), .B(n5775), .Z(n11139) );
  ANDN U6536 ( .B(x[477]), .A(y[477]), .Z(n7602) );
  ANDN U6537 ( .B(x[478]), .A(y[478]), .Z(n7612) );
  OR U6538 ( .A(n7602), .B(n7612), .Z(n11137) );
  NANDN U6539 ( .A(x[476]), .B(y[476]), .Z(n7599) );
  NANDN U6540 ( .A(x[477]), .B(y[477]), .Z(n7606) );
  AND U6541 ( .A(n7599), .B(n7606), .Z(n11135) );
  ANDN U6542 ( .B(x[475]), .A(y[475]), .Z(n7597) );
  ANDN U6543 ( .B(x[476]), .A(y[476]), .Z(n7605) );
  OR U6544 ( .A(n7597), .B(n7605), .Z(n11133) );
  NANDN U6545 ( .A(x[474]), .B(y[474]), .Z(n5778) );
  NANDN U6546 ( .A(x[475]), .B(y[475]), .Z(n7600) );
  AND U6547 ( .A(n5778), .B(n7600), .Z(n11131) );
  ANDN U6548 ( .B(x[473]), .A(y[473]), .Z(n7589) );
  ANDN U6549 ( .B(x[474]), .A(y[474]), .Z(n7594) );
  OR U6550 ( .A(n7589), .B(n7594), .Z(n11129) );
  NANDN U6551 ( .A(x[472]), .B(y[472]), .Z(n7585) );
  NANDN U6552 ( .A(x[473]), .B(y[473]), .Z(n5777) );
  AND U6553 ( .A(n7585), .B(n5777), .Z(n11127) );
  ANDN U6554 ( .B(x[471]), .A(y[471]), .Z(n7580) );
  ANDN U6555 ( .B(x[472]), .A(y[472]), .Z(n7590) );
  OR U6556 ( .A(n7580), .B(n7590), .Z(n11125) );
  NANDN U6557 ( .A(x[470]), .B(y[470]), .Z(n7577) );
  NANDN U6558 ( .A(x[471]), .B(y[471]), .Z(n7584) );
  AND U6559 ( .A(n7577), .B(n7584), .Z(n11123) );
  ANDN U6560 ( .B(x[469]), .A(y[469]), .Z(n7575) );
  ANDN U6561 ( .B(x[470]), .A(y[470]), .Z(n7583) );
  OR U6562 ( .A(n7575), .B(n7583), .Z(n11121) );
  NANDN U6563 ( .A(x[468]), .B(y[468]), .Z(n5780) );
  NANDN U6564 ( .A(x[469]), .B(y[469]), .Z(n7578) );
  AND U6565 ( .A(n5780), .B(n7578), .Z(n11119) );
  ANDN U6566 ( .B(x[467]), .A(y[467]), .Z(n7567) );
  XNOR U6567 ( .A(y[468]), .B(x[468]), .Z(n3557) );
  NANDN U6568 ( .A(n7567), .B(n3557), .Z(n11117) );
  NANDN U6569 ( .A(x[466]), .B(y[466]), .Z(n7563) );
  NANDN U6570 ( .A(x[467]), .B(y[467]), .Z(n5779) );
  AND U6571 ( .A(n7563), .B(n5779), .Z(n11115) );
  ANDN U6572 ( .B(x[465]), .A(y[465]), .Z(n7558) );
  ANDN U6573 ( .B(x[466]), .A(y[466]), .Z(n7568) );
  OR U6574 ( .A(n7558), .B(n7568), .Z(n11113) );
  NANDN U6575 ( .A(x[464]), .B(y[464]), .Z(n7555) );
  NANDN U6576 ( .A(x[465]), .B(y[465]), .Z(n7562) );
  AND U6577 ( .A(n7555), .B(n7562), .Z(n11111) );
  ANDN U6578 ( .B(x[463]), .A(y[463]), .Z(n7553) );
  XNOR U6579 ( .A(y[464]), .B(x[464]), .Z(n3558) );
  NANDN U6580 ( .A(n7553), .B(n3558), .Z(n11109) );
  NANDN U6581 ( .A(x[462]), .B(y[462]), .Z(n5782) );
  NANDN U6582 ( .A(x[463]), .B(y[463]), .Z(n7556) );
  AND U6583 ( .A(n5782), .B(n7556), .Z(n11107) );
  ANDN U6584 ( .B(x[461]), .A(y[461]), .Z(n7545) );
  XNOR U6585 ( .A(y[462]), .B(x[462]), .Z(n3559) );
  NANDN U6586 ( .A(n7545), .B(n3559), .Z(n11105) );
  NANDN U6587 ( .A(x[460]), .B(y[460]), .Z(n7541) );
  NANDN U6588 ( .A(x[461]), .B(y[461]), .Z(n5781) );
  AND U6589 ( .A(n7541), .B(n5781), .Z(n11103) );
  ANDN U6590 ( .B(x[459]), .A(y[459]), .Z(n7536) );
  ANDN U6591 ( .B(x[460]), .A(y[460]), .Z(n7546) );
  OR U6592 ( .A(n7536), .B(n7546), .Z(n11101) );
  NANDN U6593 ( .A(x[458]), .B(y[458]), .Z(n7533) );
  NANDN U6594 ( .A(x[459]), .B(y[459]), .Z(n7540) );
  AND U6595 ( .A(n7533), .B(n7540), .Z(n11099) );
  ANDN U6596 ( .B(x[457]), .A(y[457]), .Z(n7531) );
  ANDN U6597 ( .B(x[458]), .A(y[458]), .Z(n7539) );
  OR U6598 ( .A(n7531), .B(n7539), .Z(n11097) );
  NANDN U6599 ( .A(x[456]), .B(y[456]), .Z(n5784) );
  NANDN U6600 ( .A(x[457]), .B(y[457]), .Z(n7534) );
  AND U6601 ( .A(n5784), .B(n7534), .Z(n11095) );
  ANDN U6602 ( .B(x[455]), .A(y[455]), .Z(n7523) );
  XNOR U6603 ( .A(y[456]), .B(x[456]), .Z(n3560) );
  NANDN U6604 ( .A(n7523), .B(n3560), .Z(n11093) );
  NANDN U6605 ( .A(x[454]), .B(y[454]), .Z(n7519) );
  NANDN U6606 ( .A(x[455]), .B(y[455]), .Z(n5783) );
  AND U6607 ( .A(n7519), .B(n5783), .Z(n11091) );
  ANDN U6608 ( .B(x[453]), .A(y[453]), .Z(n7514) );
  ANDN U6609 ( .B(x[454]), .A(y[454]), .Z(n7524) );
  OR U6610 ( .A(n7514), .B(n7524), .Z(n11089) );
  NANDN U6611 ( .A(x[452]), .B(y[452]), .Z(n7511) );
  NANDN U6612 ( .A(x[453]), .B(y[453]), .Z(n7518) );
  AND U6613 ( .A(n7511), .B(n7518), .Z(n11087) );
  ANDN U6614 ( .B(x[451]), .A(y[451]), .Z(n7509) );
  ANDN U6615 ( .B(x[452]), .A(y[452]), .Z(n7517) );
  OR U6616 ( .A(n7509), .B(n7517), .Z(n11085) );
  NANDN U6617 ( .A(x[450]), .B(y[450]), .Z(n5786) );
  NANDN U6618 ( .A(x[451]), .B(y[451]), .Z(n7512) );
  AND U6619 ( .A(n5786), .B(n7512), .Z(n11083) );
  ANDN U6620 ( .B(x[449]), .A(y[449]), .Z(n7501) );
  ANDN U6621 ( .B(x[450]), .A(y[450]), .Z(n7506) );
  OR U6622 ( .A(n7501), .B(n7506), .Z(n11081) );
  NANDN U6623 ( .A(x[448]), .B(y[448]), .Z(n7497) );
  NANDN U6624 ( .A(x[449]), .B(y[449]), .Z(n5785) );
  AND U6625 ( .A(n7497), .B(n5785), .Z(n11079) );
  ANDN U6626 ( .B(x[447]), .A(y[447]), .Z(n7492) );
  ANDN U6627 ( .B(x[448]), .A(y[448]), .Z(n7502) );
  OR U6628 ( .A(n7492), .B(n7502), .Z(n11077) );
  NANDN U6629 ( .A(x[446]), .B(y[446]), .Z(n7489) );
  NANDN U6630 ( .A(x[447]), .B(y[447]), .Z(n7496) );
  AND U6631 ( .A(n7489), .B(n7496), .Z(n11075) );
  ANDN U6632 ( .B(x[445]), .A(y[445]), .Z(n7487) );
  ANDN U6633 ( .B(x[446]), .A(y[446]), .Z(n7495) );
  OR U6634 ( .A(n7487), .B(n7495), .Z(n11073) );
  NANDN U6635 ( .A(x[444]), .B(y[444]), .Z(n5788) );
  NANDN U6636 ( .A(x[445]), .B(y[445]), .Z(n7490) );
  AND U6637 ( .A(n5788), .B(n7490), .Z(n11071) );
  ANDN U6638 ( .B(x[443]), .A(y[443]), .Z(n7479) );
  ANDN U6639 ( .B(x[444]), .A(y[444]), .Z(n7484) );
  OR U6640 ( .A(n7479), .B(n7484), .Z(n11069) );
  NANDN U6641 ( .A(x[442]), .B(y[442]), .Z(n7475) );
  NANDN U6642 ( .A(x[443]), .B(y[443]), .Z(n5787) );
  AND U6643 ( .A(n7475), .B(n5787), .Z(n11067) );
  ANDN U6644 ( .B(x[441]), .A(y[441]), .Z(n7470) );
  ANDN U6645 ( .B(x[442]), .A(y[442]), .Z(n7480) );
  OR U6646 ( .A(n7470), .B(n7480), .Z(n11065) );
  NANDN U6647 ( .A(x[440]), .B(y[440]), .Z(n7467) );
  NANDN U6648 ( .A(x[441]), .B(y[441]), .Z(n7474) );
  AND U6649 ( .A(n7467), .B(n7474), .Z(n11063) );
  ANDN U6650 ( .B(x[439]), .A(y[439]), .Z(n7465) );
  XNOR U6651 ( .A(y[440]), .B(x[440]), .Z(n3561) );
  NANDN U6652 ( .A(n7465), .B(n3561), .Z(n11061) );
  NANDN U6653 ( .A(x[438]), .B(y[438]), .Z(n5790) );
  NANDN U6654 ( .A(x[439]), .B(y[439]), .Z(n7468) );
  AND U6655 ( .A(n5790), .B(n7468), .Z(n11059) );
  ANDN U6656 ( .B(x[437]), .A(y[437]), .Z(n7457) );
  ANDN U6657 ( .B(x[438]), .A(y[438]), .Z(n7462) );
  OR U6658 ( .A(n7457), .B(n7462), .Z(n11057) );
  NANDN U6659 ( .A(x[436]), .B(y[436]), .Z(n7453) );
  NANDN U6660 ( .A(x[437]), .B(y[437]), .Z(n5789) );
  AND U6661 ( .A(n7453), .B(n5789), .Z(n11055) );
  ANDN U6662 ( .B(x[435]), .A(y[435]), .Z(n7451) );
  ANDN U6663 ( .B(x[436]), .A(y[436]), .Z(n7458) );
  OR U6664 ( .A(n7451), .B(n7458), .Z(n11053) );
  NANDN U6665 ( .A(x[434]), .B(y[434]), .Z(n3562) );
  NANDN U6666 ( .A(x[435]), .B(y[435]), .Z(n7452) );
  AND U6667 ( .A(n3562), .B(n7452), .Z(n11051) );
  ANDN U6668 ( .B(x[433]), .A(y[433]), .Z(n7443) );
  XNOR U6669 ( .A(x[434]), .B(y[434]), .Z(n7445) );
  NANDN U6670 ( .A(n7443), .B(n7445), .Z(n11049) );
  NANDN U6671 ( .A(x[432]), .B(y[432]), .Z(n5792) );
  NANDN U6672 ( .A(x[433]), .B(y[433]), .Z(n7446) );
  AND U6673 ( .A(n5792), .B(n7446), .Z(n11047) );
  ANDN U6674 ( .B(x[431]), .A(y[431]), .Z(n7435) );
  ANDN U6675 ( .B(x[432]), .A(y[432]), .Z(n7440) );
  OR U6676 ( .A(n7435), .B(n7440), .Z(n11045) );
  NANDN U6677 ( .A(x[430]), .B(y[430]), .Z(n7431) );
  NANDN U6678 ( .A(x[431]), .B(y[431]), .Z(n5791) );
  AND U6679 ( .A(n7431), .B(n5791), .Z(n11043) );
  ANDN U6680 ( .B(x[429]), .A(y[429]), .Z(n7426) );
  ANDN U6681 ( .B(x[430]), .A(y[430]), .Z(n7436) );
  OR U6682 ( .A(n7426), .B(n7436), .Z(n11041) );
  NANDN U6683 ( .A(x[428]), .B(y[428]), .Z(n7423) );
  NANDN U6684 ( .A(x[429]), .B(y[429]), .Z(n7430) );
  AND U6685 ( .A(n7423), .B(n7430), .Z(n11039) );
  ANDN U6686 ( .B(x[427]), .A(y[427]), .Z(n7421) );
  ANDN U6687 ( .B(x[428]), .A(y[428]), .Z(n7429) );
  OR U6688 ( .A(n7421), .B(n7429), .Z(n11037) );
  NANDN U6689 ( .A(x[426]), .B(y[426]), .Z(n5794) );
  NANDN U6690 ( .A(x[427]), .B(y[427]), .Z(n7424) );
  AND U6691 ( .A(n5794), .B(n7424), .Z(n11035) );
  ANDN U6692 ( .B(x[425]), .A(y[425]), .Z(n7413) );
  ANDN U6693 ( .B(x[426]), .A(y[426]), .Z(n7418) );
  OR U6694 ( .A(n7413), .B(n7418), .Z(n11033) );
  NANDN U6695 ( .A(x[424]), .B(y[424]), .Z(n7409) );
  NANDN U6696 ( .A(x[425]), .B(y[425]), .Z(n5793) );
  AND U6697 ( .A(n7409), .B(n5793), .Z(n11031) );
  ANDN U6698 ( .B(x[423]), .A(y[423]), .Z(n7404) );
  ANDN U6699 ( .B(x[424]), .A(y[424]), .Z(n7414) );
  OR U6700 ( .A(n7404), .B(n7414), .Z(n11029) );
  NANDN U6701 ( .A(x[422]), .B(y[422]), .Z(n7401) );
  NANDN U6702 ( .A(x[423]), .B(y[423]), .Z(n7408) );
  AND U6703 ( .A(n7401), .B(n7408), .Z(n11027) );
  ANDN U6704 ( .B(x[421]), .A(y[421]), .Z(n7399) );
  XNOR U6705 ( .A(y[422]), .B(x[422]), .Z(n3563) );
  NANDN U6706 ( .A(n7399), .B(n3563), .Z(n11025) );
  NANDN U6707 ( .A(x[420]), .B(y[420]), .Z(n5796) );
  NANDN U6708 ( .A(x[421]), .B(y[421]), .Z(n7402) );
  AND U6709 ( .A(n5796), .B(n7402), .Z(n11023) );
  ANDN U6710 ( .B(x[419]), .A(y[419]), .Z(n7391) );
  ANDN U6711 ( .B(x[420]), .A(y[420]), .Z(n7396) );
  OR U6712 ( .A(n7391), .B(n7396), .Z(n11021) );
  NANDN U6713 ( .A(x[418]), .B(y[418]), .Z(n7387) );
  NANDN U6714 ( .A(x[419]), .B(y[419]), .Z(n5795) );
  AND U6715 ( .A(n7387), .B(n5795), .Z(n11019) );
  ANDN U6716 ( .B(x[417]), .A(y[417]), .Z(n7385) );
  ANDN U6717 ( .B(x[418]), .A(y[418]), .Z(n7392) );
  OR U6718 ( .A(n7385), .B(n7392), .Z(n11017) );
  NANDN U6719 ( .A(x[416]), .B(y[416]), .Z(n7383) );
  NANDN U6720 ( .A(x[417]), .B(y[417]), .Z(n7386) );
  AND U6721 ( .A(n7383), .B(n7386), .Z(n11015) );
  ANDN U6722 ( .B(x[416]), .A(y[416]), .Z(n7381) );
  ANDN U6723 ( .B(x[415]), .A(y[415]), .Z(n7377) );
  OR U6724 ( .A(n7381), .B(n7377), .Z(n11013) );
  NANDN U6725 ( .A(x[415]), .B(y[415]), .Z(n7379) );
  NANDN U6726 ( .A(x[414]), .B(y[414]), .Z(n5798) );
  AND U6727 ( .A(n7379), .B(n5798), .Z(n11011) );
  ANDN U6728 ( .B(x[413]), .A(y[413]), .Z(n7369) );
  ANDN U6729 ( .B(x[414]), .A(y[414]), .Z(n7374) );
  OR U6730 ( .A(n7369), .B(n7374), .Z(n11009) );
  NANDN U6731 ( .A(x[412]), .B(y[412]), .Z(n7365) );
  NANDN U6732 ( .A(x[413]), .B(y[413]), .Z(n5797) );
  AND U6733 ( .A(n7365), .B(n5797), .Z(n11007) );
  ANDN U6734 ( .B(x[411]), .A(y[411]), .Z(n7360) );
  ANDN U6735 ( .B(x[412]), .A(y[412]), .Z(n7370) );
  OR U6736 ( .A(n7360), .B(n7370), .Z(n11005) );
  NANDN U6737 ( .A(x[410]), .B(y[410]), .Z(n7357) );
  NANDN U6738 ( .A(x[411]), .B(y[411]), .Z(n7364) );
  AND U6739 ( .A(n7357), .B(n7364), .Z(n11003) );
  ANDN U6740 ( .B(x[409]), .A(y[409]), .Z(n7355) );
  ANDN U6741 ( .B(x[410]), .A(y[410]), .Z(n7363) );
  OR U6742 ( .A(n7355), .B(n7363), .Z(n11001) );
  NANDN U6743 ( .A(x[408]), .B(y[408]), .Z(n5800) );
  NANDN U6744 ( .A(x[409]), .B(y[409]), .Z(n7358) );
  AND U6745 ( .A(n5800), .B(n7358), .Z(n10999) );
  ANDN U6746 ( .B(x[407]), .A(y[407]), .Z(n7347) );
  ANDN U6747 ( .B(x[408]), .A(y[408]), .Z(n7352) );
  OR U6748 ( .A(n7347), .B(n7352), .Z(n10997) );
  NANDN U6749 ( .A(x[406]), .B(y[406]), .Z(n7343) );
  NANDN U6750 ( .A(x[407]), .B(y[407]), .Z(n5799) );
  AND U6751 ( .A(n7343), .B(n5799), .Z(n10995) );
  ANDN U6752 ( .B(x[405]), .A(y[405]), .Z(n7338) );
  ANDN U6753 ( .B(x[406]), .A(y[406]), .Z(n7348) );
  OR U6754 ( .A(n7338), .B(n7348), .Z(n10993) );
  NANDN U6755 ( .A(x[404]), .B(y[404]), .Z(n7335) );
  NANDN U6756 ( .A(x[405]), .B(y[405]), .Z(n7342) );
  AND U6757 ( .A(n7335), .B(n7342), .Z(n10991) );
  ANDN U6758 ( .B(x[403]), .A(y[403]), .Z(n7333) );
  ANDN U6759 ( .B(x[404]), .A(y[404]), .Z(n7341) );
  OR U6760 ( .A(n7333), .B(n7341), .Z(n10989) );
  NANDN U6761 ( .A(x[402]), .B(y[402]), .Z(n5802) );
  NANDN U6762 ( .A(x[403]), .B(y[403]), .Z(n7336) );
  AND U6763 ( .A(n5802), .B(n7336), .Z(n10987) );
  ANDN U6764 ( .B(x[401]), .A(y[401]), .Z(n7325) );
  ANDN U6765 ( .B(x[402]), .A(y[402]), .Z(n7330) );
  OR U6766 ( .A(n7325), .B(n7330), .Z(n10985) );
  NANDN U6767 ( .A(x[400]), .B(y[400]), .Z(n7321) );
  NANDN U6768 ( .A(x[401]), .B(y[401]), .Z(n5801) );
  AND U6769 ( .A(n7321), .B(n5801), .Z(n10983) );
  ANDN U6770 ( .B(x[399]), .A(y[399]), .Z(n7316) );
  ANDN U6771 ( .B(x[400]), .A(y[400]), .Z(n7326) );
  OR U6772 ( .A(n7316), .B(n7326), .Z(n10981) );
  NANDN U6773 ( .A(x[398]), .B(y[398]), .Z(n7313) );
  NANDN U6774 ( .A(x[399]), .B(y[399]), .Z(n7320) );
  AND U6775 ( .A(n7313), .B(n7320), .Z(n10979) );
  ANDN U6776 ( .B(x[397]), .A(y[397]), .Z(n7311) );
  XNOR U6777 ( .A(y[398]), .B(x[398]), .Z(n3564) );
  NANDN U6778 ( .A(n7311), .B(n3564), .Z(n10977) );
  NANDN U6779 ( .A(x[396]), .B(y[396]), .Z(n5804) );
  NANDN U6780 ( .A(x[397]), .B(y[397]), .Z(n7314) );
  AND U6781 ( .A(n5804), .B(n7314), .Z(n10975) );
  ANDN U6782 ( .B(x[395]), .A(y[395]), .Z(n7303) );
  ANDN U6783 ( .B(x[396]), .A(y[396]), .Z(n7308) );
  OR U6784 ( .A(n7303), .B(n7308), .Z(n10973) );
  NANDN U6785 ( .A(x[394]), .B(y[394]), .Z(n7299) );
  NANDN U6786 ( .A(x[395]), .B(y[395]), .Z(n5803) );
  AND U6787 ( .A(n7299), .B(n5803), .Z(n10971) );
  ANDN U6788 ( .B(x[393]), .A(y[393]), .Z(n7294) );
  ANDN U6789 ( .B(x[394]), .A(y[394]), .Z(n7304) );
  OR U6790 ( .A(n7294), .B(n7304), .Z(n10969) );
  NANDN U6791 ( .A(x[392]), .B(y[392]), .Z(n7291) );
  NANDN U6792 ( .A(x[393]), .B(y[393]), .Z(n7298) );
  AND U6793 ( .A(n7291), .B(n7298), .Z(n10967) );
  ANDN U6794 ( .B(x[391]), .A(y[391]), .Z(n7289) );
  ANDN U6795 ( .B(x[392]), .A(y[392]), .Z(n7297) );
  OR U6796 ( .A(n7289), .B(n7297), .Z(n10965) );
  NANDN U6797 ( .A(x[390]), .B(y[390]), .Z(n7285) );
  NANDN U6798 ( .A(x[391]), .B(y[391]), .Z(n7292) );
  AND U6799 ( .A(n7285), .B(n7292), .Z(n10963) );
  ANDN U6800 ( .B(x[389]), .A(y[389]), .Z(n7283) );
  ANDN U6801 ( .B(x[390]), .A(y[390]), .Z(n7286) );
  OR U6802 ( .A(n7283), .B(n7286), .Z(n10961) );
  NANDN U6803 ( .A(x[389]), .B(y[389]), .Z(n3566) );
  NANDN U6804 ( .A(x[388]), .B(y[388]), .Z(n3565) );
  AND U6805 ( .A(n3566), .B(n3565), .Z(n10959) );
  NANDN U6806 ( .A(y[387]), .B(x[387]), .Z(n3568) );
  NANDN U6807 ( .A(y[388]), .B(x[388]), .Z(n3567) );
  NAND U6808 ( .A(n3568), .B(n3567), .Z(n10957) );
  NANDN U6809 ( .A(x[387]), .B(y[387]), .Z(n3570) );
  NANDN U6810 ( .A(x[386]), .B(y[386]), .Z(n3569) );
  AND U6811 ( .A(n3570), .B(n3569), .Z(n10955) );
  NANDN U6812 ( .A(y[385]), .B(x[385]), .Z(n3572) );
  NANDN U6813 ( .A(y[386]), .B(x[386]), .Z(n3571) );
  NAND U6814 ( .A(n3572), .B(n3571), .Z(n10953) );
  NANDN U6815 ( .A(x[384]), .B(y[384]), .Z(n3574) );
  NANDN U6816 ( .A(x[385]), .B(y[385]), .Z(n3573) );
  AND U6817 ( .A(n3574), .B(n3573), .Z(n10951) );
  ANDN U6818 ( .B(x[383]), .A(y[383]), .Z(n7269) );
  XNOR U6819 ( .A(y[384]), .B(x[384]), .Z(n3575) );
  NANDN U6820 ( .A(n7269), .B(n3575), .Z(n10949) );
  NANDN U6821 ( .A(x[383]), .B(y[383]), .Z(n7273) );
  NANDN U6822 ( .A(x[382]), .B(y[382]), .Z(n7267) );
  AND U6823 ( .A(n7273), .B(n7267), .Z(n10947) );
  ANDN U6824 ( .B(x[381]), .A(y[381]), .Z(n7266) );
  ANDN U6825 ( .B(x[382]), .A(y[382]), .Z(n7272) );
  OR U6826 ( .A(n7266), .B(n7272), .Z(n10945) );
  NANDN U6827 ( .A(x[381]), .B(y[381]), .Z(n3577) );
  NANDN U6828 ( .A(x[380]), .B(y[380]), .Z(n3576) );
  AND U6829 ( .A(n3577), .B(n3576), .Z(n10943) );
  NANDN U6830 ( .A(y[379]), .B(x[379]), .Z(n3579) );
  NANDN U6831 ( .A(y[380]), .B(x[380]), .Z(n3578) );
  NAND U6832 ( .A(n3579), .B(n3578), .Z(n10941) );
  NANDN U6833 ( .A(x[379]), .B(y[379]), .Z(n7262) );
  NANDN U6834 ( .A(x[378]), .B(y[378]), .Z(n3580) );
  AND U6835 ( .A(n7262), .B(n3580), .Z(n10939) );
  ANDN U6836 ( .B(x[377]), .A(y[377]), .Z(n7254) );
  NANDN U6837 ( .A(y[378]), .B(x[378]), .Z(n7260) );
  NANDN U6838 ( .A(n7254), .B(n7260), .Z(n10937) );
  NANDN U6839 ( .A(x[376]), .B(y[376]), .Z(n5806) );
  NANDN U6840 ( .A(x[377]), .B(y[377]), .Z(n7256) );
  AND U6841 ( .A(n5806), .B(n7256), .Z(n10935) );
  ANDN U6842 ( .B(x[375]), .A(y[375]), .Z(n7246) );
  ANDN U6843 ( .B(x[376]), .A(y[376]), .Z(n7251) );
  OR U6844 ( .A(n7246), .B(n7251), .Z(n10933) );
  NANDN U6845 ( .A(x[374]), .B(y[374]), .Z(n7242) );
  NANDN U6846 ( .A(x[375]), .B(y[375]), .Z(n5805) );
  AND U6847 ( .A(n7242), .B(n5805), .Z(n10931) );
  ANDN U6848 ( .B(x[373]), .A(y[373]), .Z(n7237) );
  ANDN U6849 ( .B(x[374]), .A(y[374]), .Z(n7247) );
  OR U6850 ( .A(n7237), .B(n7247), .Z(n10929) );
  NANDN U6851 ( .A(x[372]), .B(y[372]), .Z(n7234) );
  NANDN U6852 ( .A(x[373]), .B(y[373]), .Z(n7241) );
  AND U6853 ( .A(n7234), .B(n7241), .Z(n10927) );
  ANDN U6854 ( .B(x[371]), .A(y[371]), .Z(n7232) );
  ANDN U6855 ( .B(x[372]), .A(y[372]), .Z(n7240) );
  OR U6856 ( .A(n7232), .B(n7240), .Z(n10925) );
  NANDN U6857 ( .A(x[370]), .B(y[370]), .Z(n5808) );
  NANDN U6858 ( .A(x[371]), .B(y[371]), .Z(n7235) );
  AND U6859 ( .A(n5808), .B(n7235), .Z(n10923) );
  ANDN U6860 ( .B(x[369]), .A(y[369]), .Z(n7224) );
  ANDN U6861 ( .B(x[370]), .A(y[370]), .Z(n7229) );
  OR U6862 ( .A(n7224), .B(n7229), .Z(n10921) );
  NANDN U6863 ( .A(x[368]), .B(y[368]), .Z(n7220) );
  NANDN U6864 ( .A(x[369]), .B(y[369]), .Z(n5807) );
  AND U6865 ( .A(n7220), .B(n5807), .Z(n10919) );
  ANDN U6866 ( .B(x[367]), .A(y[367]), .Z(n7215) );
  XNOR U6867 ( .A(y[368]), .B(x[368]), .Z(n3581) );
  NANDN U6868 ( .A(n7215), .B(n3581), .Z(n10917) );
  NANDN U6869 ( .A(x[366]), .B(y[366]), .Z(n7212) );
  NANDN U6870 ( .A(x[367]), .B(y[367]), .Z(n7219) );
  AND U6871 ( .A(n7212), .B(n7219), .Z(n10915) );
  ANDN U6872 ( .B(x[365]), .A(y[365]), .Z(n7210) );
  ANDN U6873 ( .B(x[366]), .A(y[366]), .Z(n7218) );
  OR U6874 ( .A(n7210), .B(n7218), .Z(n10913) );
  NANDN U6875 ( .A(x[364]), .B(y[364]), .Z(n5810) );
  NANDN U6876 ( .A(x[365]), .B(y[365]), .Z(n7213) );
  AND U6877 ( .A(n5810), .B(n7213), .Z(n10911) );
  ANDN U6878 ( .B(x[363]), .A(y[363]), .Z(n7202) );
  ANDN U6879 ( .B(x[364]), .A(y[364]), .Z(n7207) );
  OR U6880 ( .A(n7202), .B(n7207), .Z(n10909) );
  NANDN U6881 ( .A(x[362]), .B(y[362]), .Z(n7198) );
  NANDN U6882 ( .A(x[363]), .B(y[363]), .Z(n5809) );
  AND U6883 ( .A(n7198), .B(n5809), .Z(n10907) );
  ANDN U6884 ( .B(x[361]), .A(y[361]), .Z(n7193) );
  ANDN U6885 ( .B(x[362]), .A(y[362]), .Z(n7203) );
  OR U6886 ( .A(n7193), .B(n7203), .Z(n10905) );
  NANDN U6887 ( .A(x[360]), .B(y[360]), .Z(n7190) );
  NANDN U6888 ( .A(x[361]), .B(y[361]), .Z(n7197) );
  AND U6889 ( .A(n7190), .B(n7197), .Z(n10903) );
  ANDN U6890 ( .B(x[359]), .A(y[359]), .Z(n7188) );
  ANDN U6891 ( .B(x[360]), .A(y[360]), .Z(n7196) );
  OR U6892 ( .A(n7188), .B(n7196), .Z(n10901) );
  NANDN U6893 ( .A(x[358]), .B(y[358]), .Z(n5812) );
  NANDN U6894 ( .A(x[359]), .B(y[359]), .Z(n7191) );
  AND U6895 ( .A(n5812), .B(n7191), .Z(n10899) );
  ANDN U6896 ( .B(x[357]), .A(y[357]), .Z(n7180) );
  ANDN U6897 ( .B(x[358]), .A(y[358]), .Z(n7185) );
  OR U6898 ( .A(n7180), .B(n7185), .Z(n10897) );
  NANDN U6899 ( .A(x[356]), .B(y[356]), .Z(n7176) );
  NANDN U6900 ( .A(x[357]), .B(y[357]), .Z(n5811) );
  AND U6901 ( .A(n7176), .B(n5811), .Z(n10895) );
  ANDN U6902 ( .B(x[355]), .A(y[355]), .Z(n7171) );
  ANDN U6903 ( .B(x[356]), .A(y[356]), .Z(n7181) );
  OR U6904 ( .A(n7171), .B(n7181), .Z(n10893) );
  NANDN U6905 ( .A(x[354]), .B(y[354]), .Z(n7168) );
  NANDN U6906 ( .A(x[355]), .B(y[355]), .Z(n7175) );
  AND U6907 ( .A(n7168), .B(n7175), .Z(n10891) );
  ANDN U6908 ( .B(x[353]), .A(y[353]), .Z(n7166) );
  ANDN U6909 ( .B(x[354]), .A(y[354]), .Z(n7174) );
  OR U6910 ( .A(n7166), .B(n7174), .Z(n10889) );
  NANDN U6911 ( .A(x[352]), .B(y[352]), .Z(n5814) );
  NANDN U6912 ( .A(x[353]), .B(y[353]), .Z(n7169) );
  AND U6913 ( .A(n5814), .B(n7169), .Z(n10887) );
  ANDN U6914 ( .B(x[351]), .A(y[351]), .Z(n7158) );
  ANDN U6915 ( .B(x[352]), .A(y[352]), .Z(n7163) );
  OR U6916 ( .A(n7158), .B(n7163), .Z(n10885) );
  NANDN U6917 ( .A(x[350]), .B(y[350]), .Z(n7154) );
  NANDN U6918 ( .A(x[351]), .B(y[351]), .Z(n5813) );
  AND U6919 ( .A(n7154), .B(n5813), .Z(n10883) );
  ANDN U6920 ( .B(x[349]), .A(y[349]), .Z(n7149) );
  ANDN U6921 ( .B(x[350]), .A(y[350]), .Z(n7159) );
  OR U6922 ( .A(n7149), .B(n7159), .Z(n10881) );
  NANDN U6923 ( .A(x[348]), .B(y[348]), .Z(n7146) );
  NANDN U6924 ( .A(x[349]), .B(y[349]), .Z(n7153) );
  AND U6925 ( .A(n7146), .B(n7153), .Z(n10879) );
  ANDN U6926 ( .B(x[347]), .A(y[347]), .Z(n7144) );
  XNOR U6927 ( .A(y[348]), .B(x[348]), .Z(n3582) );
  NANDN U6928 ( .A(n7144), .B(n3582), .Z(n10877) );
  NANDN U6929 ( .A(x[346]), .B(y[346]), .Z(n5816) );
  NANDN U6930 ( .A(x[347]), .B(y[347]), .Z(n7147) );
  AND U6931 ( .A(n5816), .B(n7147), .Z(n10875) );
  ANDN U6932 ( .B(x[345]), .A(y[345]), .Z(n7136) );
  ANDN U6933 ( .B(x[346]), .A(y[346]), .Z(n7141) );
  OR U6934 ( .A(n7136), .B(n7141), .Z(n10873) );
  NANDN U6935 ( .A(x[344]), .B(y[344]), .Z(n7132) );
  NANDN U6936 ( .A(x[345]), .B(y[345]), .Z(n5815) );
  AND U6937 ( .A(n7132), .B(n5815), .Z(n10871) );
  ANDN U6938 ( .B(x[343]), .A(y[343]), .Z(n7127) );
  ANDN U6939 ( .B(x[344]), .A(y[344]), .Z(n7137) );
  OR U6940 ( .A(n7127), .B(n7137), .Z(n10869) );
  NANDN U6941 ( .A(x[342]), .B(y[342]), .Z(n7124) );
  NANDN U6942 ( .A(x[343]), .B(y[343]), .Z(n7131) );
  AND U6943 ( .A(n7124), .B(n7131), .Z(n10867) );
  ANDN U6944 ( .B(x[341]), .A(y[341]), .Z(n7122) );
  ANDN U6945 ( .B(x[342]), .A(y[342]), .Z(n7130) );
  OR U6946 ( .A(n7122), .B(n7130), .Z(n10865) );
  NANDN U6947 ( .A(x[340]), .B(y[340]), .Z(n5818) );
  NANDN U6948 ( .A(x[341]), .B(y[341]), .Z(n7125) );
  AND U6949 ( .A(n5818), .B(n7125), .Z(n10863) );
  ANDN U6950 ( .B(x[339]), .A(y[339]), .Z(n7114) );
  ANDN U6951 ( .B(x[340]), .A(y[340]), .Z(n7119) );
  OR U6952 ( .A(n7114), .B(n7119), .Z(n10861) );
  NANDN U6953 ( .A(x[338]), .B(y[338]), .Z(n7110) );
  NANDN U6954 ( .A(x[339]), .B(y[339]), .Z(n5817) );
  AND U6955 ( .A(n7110), .B(n5817), .Z(n10859) );
  ANDN U6956 ( .B(x[337]), .A(y[337]), .Z(n7105) );
  ANDN U6957 ( .B(x[338]), .A(y[338]), .Z(n7115) );
  OR U6958 ( .A(n7105), .B(n7115), .Z(n10857) );
  NANDN U6959 ( .A(x[336]), .B(y[336]), .Z(n7102) );
  NANDN U6960 ( .A(x[337]), .B(y[337]), .Z(n7109) );
  AND U6961 ( .A(n7102), .B(n7109), .Z(n10855) );
  ANDN U6962 ( .B(x[335]), .A(y[335]), .Z(n7100) );
  ANDN U6963 ( .B(x[336]), .A(y[336]), .Z(n7108) );
  OR U6964 ( .A(n7100), .B(n7108), .Z(n10853) );
  NANDN U6965 ( .A(x[334]), .B(y[334]), .Z(n5820) );
  NANDN U6966 ( .A(x[335]), .B(y[335]), .Z(n7103) );
  AND U6967 ( .A(n5820), .B(n7103), .Z(n10851) );
  ANDN U6968 ( .B(x[333]), .A(y[333]), .Z(n7092) );
  ANDN U6969 ( .B(x[334]), .A(y[334]), .Z(n7097) );
  OR U6970 ( .A(n7092), .B(n7097), .Z(n10849) );
  NANDN U6971 ( .A(x[332]), .B(y[332]), .Z(n7088) );
  NANDN U6972 ( .A(x[333]), .B(y[333]), .Z(n5819) );
  AND U6973 ( .A(n7088), .B(n5819), .Z(n10847) );
  ANDN U6974 ( .B(x[331]), .A(y[331]), .Z(n7083) );
  XNOR U6975 ( .A(y[332]), .B(x[332]), .Z(n3583) );
  NANDN U6976 ( .A(n7083), .B(n3583), .Z(n10845) );
  NANDN U6977 ( .A(x[330]), .B(y[330]), .Z(n7080) );
  NANDN U6978 ( .A(x[331]), .B(y[331]), .Z(n7087) );
  AND U6979 ( .A(n7080), .B(n7087), .Z(n10843) );
  ANDN U6980 ( .B(x[329]), .A(y[329]), .Z(n7078) );
  ANDN U6981 ( .B(x[330]), .A(y[330]), .Z(n7086) );
  OR U6982 ( .A(n7078), .B(n7086), .Z(n10841) );
  NANDN U6983 ( .A(x[328]), .B(y[328]), .Z(n5822) );
  NANDN U6984 ( .A(x[329]), .B(y[329]), .Z(n7081) );
  AND U6985 ( .A(n5822), .B(n7081), .Z(n10839) );
  ANDN U6986 ( .B(x[327]), .A(y[327]), .Z(n7070) );
  ANDN U6987 ( .B(x[328]), .A(y[328]), .Z(n7075) );
  OR U6988 ( .A(n7070), .B(n7075), .Z(n10837) );
  NANDN U6989 ( .A(x[326]), .B(y[326]), .Z(n7066) );
  NANDN U6990 ( .A(x[327]), .B(y[327]), .Z(n5821) );
  AND U6991 ( .A(n7066), .B(n5821), .Z(n10835) );
  ANDN U6992 ( .B(x[325]), .A(y[325]), .Z(n7061) );
  ANDN U6993 ( .B(x[326]), .A(y[326]), .Z(n7071) );
  OR U6994 ( .A(n7061), .B(n7071), .Z(n10833) );
  NANDN U6995 ( .A(x[324]), .B(y[324]), .Z(n7058) );
  NANDN U6996 ( .A(x[325]), .B(y[325]), .Z(n7065) );
  AND U6997 ( .A(n7058), .B(n7065), .Z(n10831) );
  ANDN U6998 ( .B(x[323]), .A(y[323]), .Z(n7056) );
  XNOR U6999 ( .A(y[324]), .B(x[324]), .Z(n3584) );
  NANDN U7000 ( .A(n7056), .B(n3584), .Z(n10829) );
  NANDN U7001 ( .A(x[322]), .B(y[322]), .Z(n5824) );
  NANDN U7002 ( .A(x[323]), .B(y[323]), .Z(n7059) );
  AND U7003 ( .A(n5824), .B(n7059), .Z(n10827) );
  ANDN U7004 ( .B(x[321]), .A(y[321]), .Z(n7048) );
  ANDN U7005 ( .B(x[322]), .A(y[322]), .Z(n7053) );
  OR U7006 ( .A(n7048), .B(n7053), .Z(n10825) );
  NANDN U7007 ( .A(x[320]), .B(y[320]), .Z(n7044) );
  NANDN U7008 ( .A(x[321]), .B(y[321]), .Z(n5823) );
  AND U7009 ( .A(n7044), .B(n5823), .Z(n10823) );
  ANDN U7010 ( .B(x[319]), .A(y[319]), .Z(n7042) );
  ANDN U7011 ( .B(x[320]), .A(y[320]), .Z(n7049) );
  OR U7012 ( .A(n7042), .B(n7049), .Z(n10821) );
  NANDN U7013 ( .A(x[318]), .B(y[318]), .Z(n3585) );
  NANDN U7014 ( .A(x[319]), .B(y[319]), .Z(n7043) );
  AND U7015 ( .A(n3585), .B(n7043), .Z(n10819) );
  ANDN U7016 ( .B(x[317]), .A(y[317]), .Z(n7034) );
  XNOR U7017 ( .A(x[318]), .B(y[318]), .Z(n7036) );
  NANDN U7018 ( .A(n7034), .B(n7036), .Z(n10817) );
  NANDN U7019 ( .A(x[316]), .B(y[316]), .Z(n5826) );
  NANDN U7020 ( .A(x[317]), .B(y[317]), .Z(n7037) );
  AND U7021 ( .A(n5826), .B(n7037), .Z(n10815) );
  ANDN U7022 ( .B(x[315]), .A(y[315]), .Z(n7026) );
  ANDN U7023 ( .B(x[316]), .A(y[316]), .Z(n7031) );
  OR U7024 ( .A(n7026), .B(n7031), .Z(n10813) );
  NANDN U7025 ( .A(x[314]), .B(y[314]), .Z(n7022) );
  NANDN U7026 ( .A(x[315]), .B(y[315]), .Z(n5825) );
  AND U7027 ( .A(n7022), .B(n5825), .Z(n10811) );
  ANDN U7028 ( .B(x[313]), .A(y[313]), .Z(n7017) );
  ANDN U7029 ( .B(x[314]), .A(y[314]), .Z(n7027) );
  OR U7030 ( .A(n7017), .B(n7027), .Z(n10809) );
  NANDN U7031 ( .A(x[312]), .B(y[312]), .Z(n7014) );
  NANDN U7032 ( .A(x[313]), .B(y[313]), .Z(n7021) );
  AND U7033 ( .A(n7014), .B(n7021), .Z(n10807) );
  ANDN U7034 ( .B(x[311]), .A(y[311]), .Z(n7012) );
  ANDN U7035 ( .B(x[312]), .A(y[312]), .Z(n7020) );
  OR U7036 ( .A(n7012), .B(n7020), .Z(n10805) );
  NANDN U7037 ( .A(x[310]), .B(y[310]), .Z(n5828) );
  NANDN U7038 ( .A(x[311]), .B(y[311]), .Z(n7015) );
  AND U7039 ( .A(n5828), .B(n7015), .Z(n10803) );
  ANDN U7040 ( .B(x[309]), .A(y[309]), .Z(n7004) );
  ANDN U7041 ( .B(x[310]), .A(y[310]), .Z(n7009) );
  OR U7042 ( .A(n7004), .B(n7009), .Z(n10801) );
  NANDN U7043 ( .A(x[308]), .B(y[308]), .Z(n7000) );
  NANDN U7044 ( .A(x[309]), .B(y[309]), .Z(n5827) );
  AND U7045 ( .A(n7000), .B(n5827), .Z(n10799) );
  ANDN U7046 ( .B(x[307]), .A(y[307]), .Z(n6995) );
  XNOR U7047 ( .A(y[308]), .B(x[308]), .Z(n3586) );
  NANDN U7048 ( .A(n6995), .B(n3586), .Z(n10797) );
  NANDN U7049 ( .A(x[306]), .B(y[306]), .Z(n6992) );
  NANDN U7050 ( .A(x[307]), .B(y[307]), .Z(n6999) );
  AND U7051 ( .A(n6992), .B(n6999), .Z(n10795) );
  ANDN U7052 ( .B(x[305]), .A(y[305]), .Z(n6990) );
  XNOR U7053 ( .A(y[306]), .B(x[306]), .Z(n3587) );
  NANDN U7054 ( .A(n6990), .B(n3587), .Z(n10793) );
  NANDN U7055 ( .A(x[304]), .B(y[304]), .Z(n5830) );
  NANDN U7056 ( .A(x[305]), .B(y[305]), .Z(n6993) );
  AND U7057 ( .A(n5830), .B(n6993), .Z(n10791) );
  ANDN U7058 ( .B(x[303]), .A(y[303]), .Z(n6982) );
  ANDN U7059 ( .B(x[304]), .A(y[304]), .Z(n6987) );
  OR U7060 ( .A(n6982), .B(n6987), .Z(n10789) );
  NANDN U7061 ( .A(x[302]), .B(y[302]), .Z(n6978) );
  NANDN U7062 ( .A(x[303]), .B(y[303]), .Z(n5829) );
  AND U7063 ( .A(n6978), .B(n5829), .Z(n10787) );
  ANDN U7064 ( .B(x[301]), .A(y[301]), .Z(n6973) );
  ANDN U7065 ( .B(x[302]), .A(y[302]), .Z(n6983) );
  OR U7066 ( .A(n6973), .B(n6983), .Z(n10785) );
  NANDN U7067 ( .A(x[300]), .B(y[300]), .Z(n6970) );
  NANDN U7068 ( .A(x[301]), .B(y[301]), .Z(n6977) );
  AND U7069 ( .A(n6970), .B(n6977), .Z(n10783) );
  ANDN U7070 ( .B(x[299]), .A(y[299]), .Z(n6968) );
  ANDN U7071 ( .B(x[300]), .A(y[300]), .Z(n6976) );
  OR U7072 ( .A(n6968), .B(n6976), .Z(n10781) );
  NANDN U7073 ( .A(x[298]), .B(y[298]), .Z(n5832) );
  NANDN U7074 ( .A(x[299]), .B(y[299]), .Z(n6971) );
  AND U7075 ( .A(n5832), .B(n6971), .Z(n10779) );
  ANDN U7076 ( .B(x[297]), .A(y[297]), .Z(n6960) );
  ANDN U7077 ( .B(x[298]), .A(y[298]), .Z(n6965) );
  OR U7078 ( .A(n6960), .B(n6965), .Z(n10777) );
  NANDN U7079 ( .A(x[296]), .B(y[296]), .Z(n6956) );
  NANDN U7080 ( .A(x[297]), .B(y[297]), .Z(n5831) );
  AND U7081 ( .A(n6956), .B(n5831), .Z(n10775) );
  ANDN U7082 ( .B(x[295]), .A(y[295]), .Z(n6951) );
  ANDN U7083 ( .B(x[296]), .A(y[296]), .Z(n6961) );
  OR U7084 ( .A(n6951), .B(n6961), .Z(n10773) );
  NANDN U7085 ( .A(x[294]), .B(y[294]), .Z(n6948) );
  NANDN U7086 ( .A(x[295]), .B(y[295]), .Z(n6955) );
  AND U7087 ( .A(n6948), .B(n6955), .Z(n10771) );
  ANDN U7088 ( .B(x[293]), .A(y[293]), .Z(n6946) );
  ANDN U7089 ( .B(x[294]), .A(y[294]), .Z(n6954) );
  OR U7090 ( .A(n6946), .B(n6954), .Z(n10769) );
  NANDN U7091 ( .A(x[292]), .B(y[292]), .Z(n5834) );
  NANDN U7092 ( .A(x[293]), .B(y[293]), .Z(n6949) );
  AND U7093 ( .A(n5834), .B(n6949), .Z(n10767) );
  ANDN U7094 ( .B(x[291]), .A(y[291]), .Z(n6938) );
  ANDN U7095 ( .B(x[292]), .A(y[292]), .Z(n6943) );
  OR U7096 ( .A(n6938), .B(n6943), .Z(n10765) );
  NANDN U7097 ( .A(x[290]), .B(y[290]), .Z(n6934) );
  NANDN U7098 ( .A(x[291]), .B(y[291]), .Z(n5833) );
  AND U7099 ( .A(n6934), .B(n5833), .Z(n10763) );
  ANDN U7100 ( .B(x[289]), .A(y[289]), .Z(n6929) );
  ANDN U7101 ( .B(x[290]), .A(y[290]), .Z(n6939) );
  OR U7102 ( .A(n6929), .B(n6939), .Z(n10761) );
  NANDN U7103 ( .A(x[288]), .B(y[288]), .Z(n6926) );
  NANDN U7104 ( .A(x[289]), .B(y[289]), .Z(n6933) );
  AND U7105 ( .A(n6926), .B(n6933), .Z(n10759) );
  ANDN U7106 ( .B(x[287]), .A(y[287]), .Z(n6924) );
  ANDN U7107 ( .B(x[288]), .A(y[288]), .Z(n6932) );
  OR U7108 ( .A(n6924), .B(n6932), .Z(n10757) );
  NANDN U7109 ( .A(x[286]), .B(y[286]), .Z(n5836) );
  NANDN U7110 ( .A(x[287]), .B(y[287]), .Z(n6927) );
  AND U7111 ( .A(n5836), .B(n6927), .Z(n10755) );
  ANDN U7112 ( .B(x[285]), .A(y[285]), .Z(n6916) );
  ANDN U7113 ( .B(x[286]), .A(y[286]), .Z(n6921) );
  OR U7114 ( .A(n6916), .B(n6921), .Z(n10753) );
  NANDN U7115 ( .A(x[284]), .B(y[284]), .Z(n6912) );
  NANDN U7116 ( .A(x[285]), .B(y[285]), .Z(n5835) );
  AND U7117 ( .A(n6912), .B(n5835), .Z(n10751) );
  ANDN U7118 ( .B(x[283]), .A(y[283]), .Z(n6907) );
  ANDN U7119 ( .B(x[284]), .A(y[284]), .Z(n6917) );
  OR U7120 ( .A(n6907), .B(n6917), .Z(n10749) );
  NANDN U7121 ( .A(x[282]), .B(y[282]), .Z(n6904) );
  NANDN U7122 ( .A(x[283]), .B(y[283]), .Z(n6911) );
  AND U7123 ( .A(n6904), .B(n6911), .Z(n10747) );
  ANDN U7124 ( .B(x[281]), .A(y[281]), .Z(n6902) );
  ANDN U7125 ( .B(x[282]), .A(y[282]), .Z(n6910) );
  OR U7126 ( .A(n6902), .B(n6910), .Z(n10745) );
  NANDN U7127 ( .A(x[280]), .B(y[280]), .Z(n3588) );
  NANDN U7128 ( .A(x[281]), .B(y[281]), .Z(n6905) );
  AND U7129 ( .A(n3588), .B(n6905), .Z(n10743) );
  ANDN U7130 ( .B(x[279]), .A(y[279]), .Z(n10738) );
  NANDN U7131 ( .A(x[278]), .B(y[278]), .Z(n6899) );
  NANDN U7132 ( .A(x[279]), .B(y[279]), .Z(n5837) );
  AND U7133 ( .A(n6899), .B(n5837), .Z(n10737) );
  ANDN U7134 ( .B(x[277]), .A(y[277]), .Z(n6896) );
  ANDN U7135 ( .B(x[278]), .A(y[278]), .Z(n6900) );
  OR U7136 ( .A(n6896), .B(n6900), .Z(n10735) );
  NANDN U7137 ( .A(x[276]), .B(y[276]), .Z(n6894) );
  NANDN U7138 ( .A(x[277]), .B(y[277]), .Z(n6898) );
  AND U7139 ( .A(n6894), .B(n6898), .Z(n10733) );
  ANDN U7140 ( .B(x[275]), .A(y[275]), .Z(n6893) );
  ANDN U7141 ( .B(x[276]), .A(y[276]), .Z(n6897) );
  OR U7142 ( .A(n6893), .B(n6897), .Z(n10731) );
  NANDN U7143 ( .A(x[274]), .B(y[274]), .Z(n5839) );
  NANDN U7144 ( .A(x[275]), .B(y[275]), .Z(n6895) );
  AND U7145 ( .A(n5839), .B(n6895), .Z(n10729) );
  ANDN U7146 ( .B(x[273]), .A(y[273]), .Z(n6890) );
  ANDN U7147 ( .B(x[274]), .A(y[274]), .Z(n6892) );
  OR U7148 ( .A(n6890), .B(n6892), .Z(n10727) );
  NANDN U7149 ( .A(x[272]), .B(y[272]), .Z(n6887) );
  NANDN U7150 ( .A(x[273]), .B(y[273]), .Z(n5838) );
  AND U7151 ( .A(n6887), .B(n5838), .Z(n10725) );
  ANDN U7152 ( .B(x[271]), .A(y[271]), .Z(n6882) );
  ANDN U7153 ( .B(x[272]), .A(y[272]), .Z(n6891) );
  OR U7154 ( .A(n6882), .B(n6891), .Z(n10723) );
  NANDN U7155 ( .A(x[270]), .B(y[270]), .Z(n6879) );
  NANDN U7156 ( .A(x[271]), .B(y[271]), .Z(n6886) );
  AND U7157 ( .A(n6879), .B(n6886), .Z(n10721) );
  ANDN U7158 ( .B(x[269]), .A(y[269]), .Z(n6877) );
  ANDN U7159 ( .B(x[270]), .A(y[270]), .Z(n6885) );
  OR U7160 ( .A(n6877), .B(n6885), .Z(n10719) );
  NANDN U7161 ( .A(x[268]), .B(y[268]), .Z(n5841) );
  NANDN U7162 ( .A(x[269]), .B(y[269]), .Z(n6880) );
  AND U7163 ( .A(n5841), .B(n6880), .Z(n10717) );
  ANDN U7164 ( .B(x[267]), .A(y[267]), .Z(n6869) );
  ANDN U7165 ( .B(x[268]), .A(y[268]), .Z(n6874) );
  OR U7166 ( .A(n6869), .B(n6874), .Z(n10715) );
  NANDN U7167 ( .A(x[266]), .B(y[266]), .Z(n6865) );
  NANDN U7168 ( .A(x[267]), .B(y[267]), .Z(n5840) );
  AND U7169 ( .A(n6865), .B(n5840), .Z(n10713) );
  ANDN U7170 ( .B(x[265]), .A(y[265]), .Z(n6860) );
  ANDN U7171 ( .B(x[266]), .A(y[266]), .Z(n6870) );
  OR U7172 ( .A(n6860), .B(n6870), .Z(n10711) );
  NANDN U7173 ( .A(x[264]), .B(y[264]), .Z(n6857) );
  NANDN U7174 ( .A(x[265]), .B(y[265]), .Z(n6864) );
  AND U7175 ( .A(n6857), .B(n6864), .Z(n10709) );
  ANDN U7176 ( .B(x[263]), .A(y[263]), .Z(n6855) );
  ANDN U7177 ( .B(x[264]), .A(y[264]), .Z(n6863) );
  OR U7178 ( .A(n6855), .B(n6863), .Z(n10707) );
  NANDN U7179 ( .A(x[262]), .B(y[262]), .Z(n5843) );
  NANDN U7180 ( .A(x[263]), .B(y[263]), .Z(n6858) );
  AND U7181 ( .A(n5843), .B(n6858), .Z(n10705) );
  ANDN U7182 ( .B(x[261]), .A(y[261]), .Z(n6847) );
  ANDN U7183 ( .B(x[262]), .A(y[262]), .Z(n6852) );
  OR U7184 ( .A(n6847), .B(n6852), .Z(n10703) );
  NANDN U7185 ( .A(x[260]), .B(y[260]), .Z(n6843) );
  NANDN U7186 ( .A(x[261]), .B(y[261]), .Z(n5842) );
  AND U7187 ( .A(n6843), .B(n5842), .Z(n10701) );
  ANDN U7188 ( .B(x[259]), .A(y[259]), .Z(n6838) );
  ANDN U7189 ( .B(x[260]), .A(y[260]), .Z(n6848) );
  OR U7190 ( .A(n6838), .B(n6848), .Z(n10699) );
  NANDN U7191 ( .A(x[258]), .B(y[258]), .Z(n6835) );
  NANDN U7192 ( .A(x[259]), .B(y[259]), .Z(n6842) );
  AND U7193 ( .A(n6835), .B(n6842), .Z(n10697) );
  ANDN U7194 ( .B(x[257]), .A(y[257]), .Z(n6833) );
  ANDN U7195 ( .B(x[258]), .A(y[258]), .Z(n6841) );
  OR U7196 ( .A(n6833), .B(n6841), .Z(n10695) );
  NANDN U7197 ( .A(x[256]), .B(y[256]), .Z(n5845) );
  NANDN U7198 ( .A(x[257]), .B(y[257]), .Z(n6836) );
  AND U7199 ( .A(n5845), .B(n6836), .Z(n10693) );
  ANDN U7200 ( .B(x[255]), .A(y[255]), .Z(n6825) );
  ANDN U7201 ( .B(x[256]), .A(y[256]), .Z(n6830) );
  OR U7202 ( .A(n6825), .B(n6830), .Z(n10691) );
  NANDN U7203 ( .A(x[254]), .B(y[254]), .Z(n6821) );
  NANDN U7204 ( .A(x[255]), .B(y[255]), .Z(n5844) );
  AND U7205 ( .A(n6821), .B(n5844), .Z(n10689) );
  ANDN U7206 ( .B(x[253]), .A(y[253]), .Z(n6816) );
  ANDN U7207 ( .B(x[254]), .A(y[254]), .Z(n6826) );
  OR U7208 ( .A(n6816), .B(n6826), .Z(n10687) );
  NANDN U7209 ( .A(x[252]), .B(y[252]), .Z(n6813) );
  NANDN U7210 ( .A(x[253]), .B(y[253]), .Z(n6820) );
  AND U7211 ( .A(n6813), .B(n6820), .Z(n10685) );
  ANDN U7212 ( .B(x[251]), .A(y[251]), .Z(n6811) );
  ANDN U7213 ( .B(x[252]), .A(y[252]), .Z(n6819) );
  OR U7214 ( .A(n6811), .B(n6819), .Z(n10683) );
  NANDN U7215 ( .A(x[250]), .B(y[250]), .Z(n5847) );
  NANDN U7216 ( .A(x[251]), .B(y[251]), .Z(n6814) );
  AND U7217 ( .A(n5847), .B(n6814), .Z(n10681) );
  ANDN U7218 ( .B(x[249]), .A(y[249]), .Z(n6803) );
  ANDN U7219 ( .B(x[250]), .A(y[250]), .Z(n6808) );
  OR U7220 ( .A(n6803), .B(n6808), .Z(n10679) );
  NANDN U7221 ( .A(x[248]), .B(y[248]), .Z(n6799) );
  NANDN U7222 ( .A(x[249]), .B(y[249]), .Z(n5846) );
  AND U7223 ( .A(n6799), .B(n5846), .Z(n10677) );
  ANDN U7224 ( .B(x[247]), .A(y[247]), .Z(n6794) );
  ANDN U7225 ( .B(x[248]), .A(y[248]), .Z(n6804) );
  OR U7226 ( .A(n6794), .B(n6804), .Z(n10675) );
  NANDN U7227 ( .A(x[246]), .B(y[246]), .Z(n6791) );
  NANDN U7228 ( .A(x[247]), .B(y[247]), .Z(n6798) );
  AND U7229 ( .A(n6791), .B(n6798), .Z(n10673) );
  ANDN U7230 ( .B(x[245]), .A(y[245]), .Z(n6789) );
  ANDN U7231 ( .B(x[246]), .A(y[246]), .Z(n6797) );
  OR U7232 ( .A(n6789), .B(n6797), .Z(n10671) );
  NANDN U7233 ( .A(x[244]), .B(y[244]), .Z(n5849) );
  NANDN U7234 ( .A(x[245]), .B(y[245]), .Z(n6792) );
  AND U7235 ( .A(n5849), .B(n6792), .Z(n10669) );
  ANDN U7236 ( .B(x[243]), .A(y[243]), .Z(n6781) );
  ANDN U7237 ( .B(x[244]), .A(y[244]), .Z(n6786) );
  OR U7238 ( .A(n6781), .B(n6786), .Z(n10667) );
  NANDN U7239 ( .A(x[242]), .B(y[242]), .Z(n6777) );
  NANDN U7240 ( .A(x[243]), .B(y[243]), .Z(n5848) );
  AND U7241 ( .A(n6777), .B(n5848), .Z(n10665) );
  ANDN U7242 ( .B(x[241]), .A(y[241]), .Z(n6772) );
  ANDN U7243 ( .B(x[242]), .A(y[242]), .Z(n6782) );
  OR U7244 ( .A(n6772), .B(n6782), .Z(n10663) );
  NANDN U7245 ( .A(x[240]), .B(y[240]), .Z(n6769) );
  NANDN U7246 ( .A(x[241]), .B(y[241]), .Z(n6776) );
  AND U7247 ( .A(n6769), .B(n6776), .Z(n10661) );
  ANDN U7248 ( .B(x[239]), .A(y[239]), .Z(n6767) );
  ANDN U7249 ( .B(x[240]), .A(y[240]), .Z(n6775) );
  OR U7250 ( .A(n6767), .B(n6775), .Z(n10659) );
  NANDN U7251 ( .A(x[238]), .B(y[238]), .Z(n5851) );
  NANDN U7252 ( .A(x[239]), .B(y[239]), .Z(n6770) );
  AND U7253 ( .A(n5851), .B(n6770), .Z(n10657) );
  ANDN U7254 ( .B(x[237]), .A(y[237]), .Z(n6759) );
  ANDN U7255 ( .B(x[238]), .A(y[238]), .Z(n6764) );
  OR U7256 ( .A(n6759), .B(n6764), .Z(n10655) );
  NANDN U7257 ( .A(x[236]), .B(y[236]), .Z(n6755) );
  NANDN U7258 ( .A(x[237]), .B(y[237]), .Z(n5850) );
  AND U7259 ( .A(n6755), .B(n5850), .Z(n10653) );
  ANDN U7260 ( .B(x[235]), .A(y[235]), .Z(n6750) );
  ANDN U7261 ( .B(x[236]), .A(y[236]), .Z(n6760) );
  OR U7262 ( .A(n6750), .B(n6760), .Z(n10651) );
  NANDN U7263 ( .A(x[234]), .B(y[234]), .Z(n6747) );
  NANDN U7264 ( .A(x[235]), .B(y[235]), .Z(n6754) );
  AND U7265 ( .A(n6747), .B(n6754), .Z(n10649) );
  ANDN U7266 ( .B(x[233]), .A(y[233]), .Z(n6745) );
  ANDN U7267 ( .B(x[234]), .A(y[234]), .Z(n6753) );
  OR U7268 ( .A(n6745), .B(n6753), .Z(n10647) );
  NANDN U7269 ( .A(x[232]), .B(y[232]), .Z(n5853) );
  NANDN U7270 ( .A(x[233]), .B(y[233]), .Z(n6748) );
  AND U7271 ( .A(n5853), .B(n6748), .Z(n10645) );
  ANDN U7272 ( .B(x[231]), .A(y[231]), .Z(n6737) );
  ANDN U7273 ( .B(x[232]), .A(y[232]), .Z(n6742) );
  OR U7274 ( .A(n6737), .B(n6742), .Z(n10643) );
  NANDN U7275 ( .A(x[230]), .B(y[230]), .Z(n6733) );
  NANDN U7276 ( .A(x[231]), .B(y[231]), .Z(n5852) );
  AND U7277 ( .A(n6733), .B(n5852), .Z(n10641) );
  ANDN U7278 ( .B(x[229]), .A(y[229]), .Z(n6728) );
  ANDN U7279 ( .B(x[230]), .A(y[230]), .Z(n6738) );
  OR U7280 ( .A(n6728), .B(n6738), .Z(n10639) );
  NANDN U7281 ( .A(x[228]), .B(y[228]), .Z(n6725) );
  NANDN U7282 ( .A(x[229]), .B(y[229]), .Z(n6732) );
  AND U7283 ( .A(n6725), .B(n6732), .Z(n10637) );
  ANDN U7284 ( .B(x[227]), .A(y[227]), .Z(n6723) );
  ANDN U7285 ( .B(x[228]), .A(y[228]), .Z(n6731) );
  OR U7286 ( .A(n6723), .B(n6731), .Z(n10635) );
  NANDN U7287 ( .A(x[226]), .B(y[226]), .Z(n5855) );
  NANDN U7288 ( .A(x[227]), .B(y[227]), .Z(n6726) );
  AND U7289 ( .A(n5855), .B(n6726), .Z(n10633) );
  ANDN U7290 ( .B(x[225]), .A(y[225]), .Z(n6715) );
  ANDN U7291 ( .B(x[226]), .A(y[226]), .Z(n6720) );
  OR U7292 ( .A(n6715), .B(n6720), .Z(n10631) );
  NANDN U7293 ( .A(x[224]), .B(y[224]), .Z(n6711) );
  NANDN U7294 ( .A(x[225]), .B(y[225]), .Z(n5854) );
  AND U7295 ( .A(n6711), .B(n5854), .Z(n10629) );
  ANDN U7296 ( .B(x[223]), .A(y[223]), .Z(n6706) );
  ANDN U7297 ( .B(x[224]), .A(y[224]), .Z(n6716) );
  OR U7298 ( .A(n6706), .B(n6716), .Z(n10627) );
  NANDN U7299 ( .A(x[222]), .B(y[222]), .Z(n6703) );
  NANDN U7300 ( .A(x[223]), .B(y[223]), .Z(n6710) );
  AND U7301 ( .A(n6703), .B(n6710), .Z(n10625) );
  ANDN U7302 ( .B(x[221]), .A(y[221]), .Z(n6701) );
  ANDN U7303 ( .B(x[222]), .A(y[222]), .Z(n6709) );
  OR U7304 ( .A(n6701), .B(n6709), .Z(n10623) );
  NANDN U7305 ( .A(x[220]), .B(y[220]), .Z(n5857) );
  NANDN U7306 ( .A(x[221]), .B(y[221]), .Z(n6704) );
  AND U7307 ( .A(n5857), .B(n6704), .Z(n10621) );
  ANDN U7308 ( .B(x[219]), .A(y[219]), .Z(n6693) );
  ANDN U7309 ( .B(x[220]), .A(y[220]), .Z(n6698) );
  OR U7310 ( .A(n6693), .B(n6698), .Z(n10619) );
  NANDN U7311 ( .A(x[218]), .B(y[218]), .Z(n6689) );
  NANDN U7312 ( .A(x[219]), .B(y[219]), .Z(n5856) );
  AND U7313 ( .A(n6689), .B(n5856), .Z(n10617) );
  ANDN U7314 ( .B(x[217]), .A(y[217]), .Z(n6687) );
  ANDN U7315 ( .B(x[218]), .A(y[218]), .Z(n6694) );
  OR U7316 ( .A(n6687), .B(n6694), .Z(n10615) );
  NANDN U7317 ( .A(x[216]), .B(y[216]), .Z(n3589) );
  NANDN U7318 ( .A(x[217]), .B(y[217]), .Z(n6688) );
  AND U7319 ( .A(n3589), .B(n6688), .Z(n10613) );
  ANDN U7320 ( .B(x[215]), .A(y[215]), .Z(n6679) );
  XNOR U7321 ( .A(x[216]), .B(y[216]), .Z(n6681) );
  NANDN U7322 ( .A(n6679), .B(n6681), .Z(n10611) );
  NANDN U7323 ( .A(x[214]), .B(y[214]), .Z(n5859) );
  NANDN U7324 ( .A(x[215]), .B(y[215]), .Z(n6682) );
  AND U7325 ( .A(n5859), .B(n6682), .Z(n10609) );
  ANDN U7326 ( .B(x[213]), .A(y[213]), .Z(n6671) );
  ANDN U7327 ( .B(x[214]), .A(y[214]), .Z(n6676) );
  OR U7328 ( .A(n6671), .B(n6676), .Z(n10607) );
  NANDN U7329 ( .A(x[212]), .B(y[212]), .Z(n6667) );
  NANDN U7330 ( .A(x[213]), .B(y[213]), .Z(n5858) );
  AND U7331 ( .A(n6667), .B(n5858), .Z(n10605) );
  ANDN U7332 ( .B(x[211]), .A(y[211]), .Z(n6662) );
  ANDN U7333 ( .B(x[212]), .A(y[212]), .Z(n6672) );
  OR U7334 ( .A(n6662), .B(n6672), .Z(n10603) );
  NANDN U7335 ( .A(x[210]), .B(y[210]), .Z(n6659) );
  NANDN U7336 ( .A(x[211]), .B(y[211]), .Z(n6666) );
  AND U7337 ( .A(n6659), .B(n6666), .Z(n10601) );
  ANDN U7338 ( .B(x[209]), .A(y[209]), .Z(n6657) );
  ANDN U7339 ( .B(x[210]), .A(y[210]), .Z(n6665) );
  OR U7340 ( .A(n6657), .B(n6665), .Z(n10599) );
  NANDN U7341 ( .A(x[208]), .B(y[208]), .Z(n5861) );
  NANDN U7342 ( .A(x[209]), .B(y[209]), .Z(n6660) );
  AND U7343 ( .A(n5861), .B(n6660), .Z(n10597) );
  ANDN U7344 ( .B(x[207]), .A(y[207]), .Z(n6649) );
  ANDN U7345 ( .B(x[208]), .A(y[208]), .Z(n6654) );
  OR U7346 ( .A(n6649), .B(n6654), .Z(n10595) );
  NANDN U7347 ( .A(x[206]), .B(y[206]), .Z(n6645) );
  NANDN U7348 ( .A(x[207]), .B(y[207]), .Z(n5860) );
  AND U7349 ( .A(n6645), .B(n5860), .Z(n10593) );
  ANDN U7350 ( .B(x[205]), .A(y[205]), .Z(n6643) );
  ANDN U7351 ( .B(x[206]), .A(y[206]), .Z(n6650) );
  OR U7352 ( .A(n6643), .B(n6650), .Z(n10591) );
  NANDN U7353 ( .A(x[204]), .B(y[204]), .Z(n3590) );
  NANDN U7354 ( .A(x[205]), .B(y[205]), .Z(n6644) );
  AND U7355 ( .A(n3590), .B(n6644), .Z(n10589) );
  ANDN U7356 ( .B(x[203]), .A(y[203]), .Z(n6635) );
  XNOR U7357 ( .A(x[204]), .B(y[204]), .Z(n6637) );
  NANDN U7358 ( .A(n6635), .B(n6637), .Z(n10587) );
  NANDN U7359 ( .A(x[202]), .B(y[202]), .Z(n5863) );
  NANDN U7360 ( .A(x[203]), .B(y[203]), .Z(n6638) );
  AND U7361 ( .A(n5863), .B(n6638), .Z(n10585) );
  ANDN U7362 ( .B(x[201]), .A(y[201]), .Z(n6627) );
  ANDN U7363 ( .B(x[202]), .A(y[202]), .Z(n6632) );
  OR U7364 ( .A(n6627), .B(n6632), .Z(n10583) );
  NANDN U7365 ( .A(x[200]), .B(y[200]), .Z(n6623) );
  NANDN U7366 ( .A(x[201]), .B(y[201]), .Z(n5862) );
  AND U7367 ( .A(n6623), .B(n5862), .Z(n10581) );
  ANDN U7368 ( .B(x[199]), .A(y[199]), .Z(n6618) );
  ANDN U7369 ( .B(x[200]), .A(y[200]), .Z(n6628) );
  OR U7370 ( .A(n6618), .B(n6628), .Z(n10579) );
  NANDN U7371 ( .A(x[198]), .B(y[198]), .Z(n6615) );
  NANDN U7372 ( .A(x[199]), .B(y[199]), .Z(n6622) );
  AND U7373 ( .A(n6615), .B(n6622), .Z(n10577) );
  ANDN U7374 ( .B(x[197]), .A(y[197]), .Z(n6613) );
  ANDN U7375 ( .B(x[198]), .A(y[198]), .Z(n6621) );
  OR U7376 ( .A(n6613), .B(n6621), .Z(n10575) );
  NANDN U7377 ( .A(x[196]), .B(y[196]), .Z(n5865) );
  NANDN U7378 ( .A(x[197]), .B(y[197]), .Z(n6616) );
  AND U7379 ( .A(n5865), .B(n6616), .Z(n10573) );
  ANDN U7380 ( .B(x[195]), .A(y[195]), .Z(n6605) );
  ANDN U7381 ( .B(x[196]), .A(y[196]), .Z(n6610) );
  OR U7382 ( .A(n6605), .B(n6610), .Z(n10571) );
  NANDN U7383 ( .A(x[194]), .B(y[194]), .Z(n6601) );
  NANDN U7384 ( .A(x[195]), .B(y[195]), .Z(n5864) );
  AND U7385 ( .A(n6601), .B(n5864), .Z(n10569) );
  ANDN U7386 ( .B(x[193]), .A(y[193]), .Z(n6596) );
  ANDN U7387 ( .B(x[194]), .A(y[194]), .Z(n6606) );
  OR U7388 ( .A(n6596), .B(n6606), .Z(n10567) );
  NANDN U7389 ( .A(x[192]), .B(y[192]), .Z(n6593) );
  NANDN U7390 ( .A(x[193]), .B(y[193]), .Z(n6600) );
  AND U7391 ( .A(n6593), .B(n6600), .Z(n10565) );
  ANDN U7392 ( .B(x[191]), .A(y[191]), .Z(n6591) );
  ANDN U7393 ( .B(x[192]), .A(y[192]), .Z(n6599) );
  OR U7394 ( .A(n6591), .B(n6599), .Z(n10563) );
  NANDN U7395 ( .A(x[190]), .B(y[190]), .Z(n5867) );
  NANDN U7396 ( .A(x[191]), .B(y[191]), .Z(n6594) );
  AND U7397 ( .A(n5867), .B(n6594), .Z(n10561) );
  ANDN U7398 ( .B(x[189]), .A(y[189]), .Z(n6583) );
  ANDN U7399 ( .B(x[190]), .A(y[190]), .Z(n6588) );
  OR U7400 ( .A(n6583), .B(n6588), .Z(n10559) );
  NANDN U7401 ( .A(x[188]), .B(y[188]), .Z(n6579) );
  NANDN U7402 ( .A(x[189]), .B(y[189]), .Z(n5866) );
  AND U7403 ( .A(n6579), .B(n5866), .Z(n10557) );
  ANDN U7404 ( .B(x[187]), .A(y[187]), .Z(n6574) );
  ANDN U7405 ( .B(x[188]), .A(y[188]), .Z(n6584) );
  OR U7406 ( .A(n6574), .B(n6584), .Z(n10555) );
  NANDN U7407 ( .A(x[186]), .B(y[186]), .Z(n6571) );
  NANDN U7408 ( .A(x[187]), .B(y[187]), .Z(n6578) );
  AND U7409 ( .A(n6571), .B(n6578), .Z(n10553) );
  ANDN U7410 ( .B(x[185]), .A(y[185]), .Z(n6569) );
  ANDN U7411 ( .B(x[186]), .A(y[186]), .Z(n6577) );
  OR U7412 ( .A(n6569), .B(n6577), .Z(n10551) );
  NANDN U7413 ( .A(x[184]), .B(y[184]), .Z(n5869) );
  NANDN U7414 ( .A(x[185]), .B(y[185]), .Z(n6572) );
  AND U7415 ( .A(n5869), .B(n6572), .Z(n10549) );
  ANDN U7416 ( .B(x[183]), .A(y[183]), .Z(n6561) );
  ANDN U7417 ( .B(x[184]), .A(y[184]), .Z(n6566) );
  OR U7418 ( .A(n6561), .B(n6566), .Z(n10547) );
  NANDN U7419 ( .A(x[182]), .B(y[182]), .Z(n6557) );
  NANDN U7420 ( .A(x[183]), .B(y[183]), .Z(n5868) );
  AND U7421 ( .A(n6557), .B(n5868), .Z(n10545) );
  ANDN U7422 ( .B(x[181]), .A(y[181]), .Z(n6555) );
  ANDN U7423 ( .B(x[182]), .A(y[182]), .Z(n6562) );
  OR U7424 ( .A(n6555), .B(n6562), .Z(n10543) );
  NANDN U7425 ( .A(x[180]), .B(y[180]), .Z(n3591) );
  NANDN U7426 ( .A(x[181]), .B(y[181]), .Z(n6556) );
  AND U7427 ( .A(n3591), .B(n6556), .Z(n10541) );
  ANDN U7428 ( .B(x[179]), .A(y[179]), .Z(n6547) );
  XNOR U7429 ( .A(x[180]), .B(y[180]), .Z(n6549) );
  NANDN U7430 ( .A(n6547), .B(n6549), .Z(n10539) );
  NANDN U7431 ( .A(x[178]), .B(y[178]), .Z(n5871) );
  NANDN U7432 ( .A(x[179]), .B(y[179]), .Z(n6550) );
  AND U7433 ( .A(n5871), .B(n6550), .Z(n10537) );
  ANDN U7434 ( .B(x[177]), .A(y[177]), .Z(n6539) );
  ANDN U7435 ( .B(x[178]), .A(y[178]), .Z(n6544) );
  OR U7436 ( .A(n6539), .B(n6544), .Z(n10535) );
  NANDN U7437 ( .A(x[176]), .B(y[176]), .Z(n6535) );
  NANDN U7438 ( .A(x[177]), .B(y[177]), .Z(n5870) );
  AND U7439 ( .A(n6535), .B(n5870), .Z(n10533) );
  ANDN U7440 ( .B(x[175]), .A(y[175]), .Z(n6530) );
  ANDN U7441 ( .B(x[176]), .A(y[176]), .Z(n6540) );
  OR U7442 ( .A(n6530), .B(n6540), .Z(n10531) );
  NANDN U7443 ( .A(x[174]), .B(y[174]), .Z(n6527) );
  NANDN U7444 ( .A(x[175]), .B(y[175]), .Z(n6534) );
  AND U7445 ( .A(n6527), .B(n6534), .Z(n10529) );
  ANDN U7446 ( .B(x[173]), .A(y[173]), .Z(n6525) );
  ANDN U7447 ( .B(x[174]), .A(y[174]), .Z(n6533) );
  OR U7448 ( .A(n6525), .B(n6533), .Z(n10527) );
  NANDN U7449 ( .A(x[172]), .B(y[172]), .Z(n5873) );
  NANDN U7450 ( .A(x[173]), .B(y[173]), .Z(n6528) );
  AND U7451 ( .A(n5873), .B(n6528), .Z(n10525) );
  ANDN U7452 ( .B(x[171]), .A(y[171]), .Z(n6517) );
  ANDN U7453 ( .B(x[172]), .A(y[172]), .Z(n6522) );
  OR U7454 ( .A(n6517), .B(n6522), .Z(n10523) );
  NANDN U7455 ( .A(x[170]), .B(y[170]), .Z(n6513) );
  NANDN U7456 ( .A(x[171]), .B(y[171]), .Z(n5872) );
  AND U7457 ( .A(n6513), .B(n5872), .Z(n10521) );
  ANDN U7458 ( .B(x[169]), .A(y[169]), .Z(n6508) );
  ANDN U7459 ( .B(x[170]), .A(y[170]), .Z(n6518) );
  OR U7460 ( .A(n6508), .B(n6518), .Z(n10519) );
  NANDN U7461 ( .A(x[168]), .B(y[168]), .Z(n6505) );
  NANDN U7462 ( .A(x[169]), .B(y[169]), .Z(n6512) );
  AND U7463 ( .A(n6505), .B(n6512), .Z(n10517) );
  ANDN U7464 ( .B(x[167]), .A(y[167]), .Z(n6503) );
  ANDN U7465 ( .B(x[168]), .A(y[168]), .Z(n6511) );
  OR U7466 ( .A(n6503), .B(n6511), .Z(n10515) );
  NANDN U7467 ( .A(x[166]), .B(y[166]), .Z(n5875) );
  NANDN U7468 ( .A(x[167]), .B(y[167]), .Z(n6506) );
  AND U7469 ( .A(n5875), .B(n6506), .Z(n10513) );
  ANDN U7470 ( .B(x[165]), .A(y[165]), .Z(n6495) );
  ANDN U7471 ( .B(x[166]), .A(y[166]), .Z(n6500) );
  OR U7472 ( .A(n6495), .B(n6500), .Z(n10511) );
  NANDN U7473 ( .A(x[164]), .B(y[164]), .Z(n6491) );
  NANDN U7474 ( .A(x[165]), .B(y[165]), .Z(n5874) );
  AND U7475 ( .A(n6491), .B(n5874), .Z(n10509) );
  ANDN U7476 ( .B(x[163]), .A(y[163]), .Z(n6486) );
  ANDN U7477 ( .B(x[164]), .A(y[164]), .Z(n6496) );
  OR U7478 ( .A(n6486), .B(n6496), .Z(n10507) );
  NANDN U7479 ( .A(x[162]), .B(y[162]), .Z(n6483) );
  NANDN U7480 ( .A(x[163]), .B(y[163]), .Z(n6490) );
  AND U7481 ( .A(n6483), .B(n6490), .Z(n10505) );
  ANDN U7482 ( .B(x[161]), .A(y[161]), .Z(n6481) );
  ANDN U7483 ( .B(x[162]), .A(y[162]), .Z(n6489) );
  OR U7484 ( .A(n6481), .B(n6489), .Z(n10503) );
  NANDN U7485 ( .A(x[160]), .B(y[160]), .Z(n5877) );
  NANDN U7486 ( .A(x[161]), .B(y[161]), .Z(n6484) );
  AND U7487 ( .A(n5877), .B(n6484), .Z(n10501) );
  ANDN U7488 ( .B(x[159]), .A(y[159]), .Z(n6478) );
  ANDN U7489 ( .B(x[160]), .A(y[160]), .Z(n6480) );
  OR U7490 ( .A(n6478), .B(n6480), .Z(n10499) );
  NANDN U7491 ( .A(x[158]), .B(y[158]), .Z(n6477) );
  NANDN U7492 ( .A(x[159]), .B(y[159]), .Z(n5876) );
  AND U7493 ( .A(n6477), .B(n5876), .Z(n10497) );
  ANDN U7494 ( .B(x[157]), .A(y[157]), .Z(n6474) );
  ANDN U7495 ( .B(x[158]), .A(y[158]), .Z(n6479) );
  OR U7496 ( .A(n6474), .B(n6479), .Z(n10495) );
  NANDN U7497 ( .A(x[156]), .B(y[156]), .Z(n6473) );
  NANDN U7498 ( .A(x[157]), .B(y[157]), .Z(n6476) );
  AND U7499 ( .A(n6473), .B(n6476), .Z(n10493) );
  ANDN U7500 ( .B(x[155]), .A(y[155]), .Z(n6472) );
  ANDN U7501 ( .B(x[156]), .A(y[156]), .Z(n6475) );
  OR U7502 ( .A(n6472), .B(n6475), .Z(n10491) );
  NANDN U7503 ( .A(y[153]), .B(x[153]), .Z(n3593) );
  NANDN U7504 ( .A(y[154]), .B(x[154]), .Z(n3592) );
  AND U7505 ( .A(n3593), .B(n3592), .Z(n10486) );
  NANDN U7506 ( .A(x[153]), .B(y[153]), .Z(n6471) );
  NANDN U7507 ( .A(x[152]), .B(y[152]), .Z(n6468) );
  AND U7508 ( .A(n6471), .B(n6468), .Z(n10485) );
  ANDN U7509 ( .B(x[152]), .A(y[152]), .Z(n6470) );
  ANDN U7510 ( .B(x[151]), .A(y[151]), .Z(n6466) );
  OR U7511 ( .A(n6470), .B(n6466), .Z(n10483) );
  NANDN U7512 ( .A(x[150]), .B(y[150]), .Z(n5879) );
  NANDN U7513 ( .A(x[151]), .B(y[151]), .Z(n6469) );
  AND U7514 ( .A(n5879), .B(n6469), .Z(n10481) );
  ANDN U7515 ( .B(x[149]), .A(y[149]), .Z(n6458) );
  ANDN U7516 ( .B(x[150]), .A(y[150]), .Z(n6463) );
  OR U7517 ( .A(n6458), .B(n6463), .Z(n10479) );
  NANDN U7518 ( .A(x[148]), .B(y[148]), .Z(n6454) );
  NANDN U7519 ( .A(x[149]), .B(y[149]), .Z(n5878) );
  AND U7520 ( .A(n6454), .B(n5878), .Z(n10477) );
  ANDN U7521 ( .B(x[147]), .A(y[147]), .Z(n6449) );
  ANDN U7522 ( .B(x[148]), .A(y[148]), .Z(n6459) );
  OR U7523 ( .A(n6449), .B(n6459), .Z(n10475) );
  NANDN U7524 ( .A(x[146]), .B(y[146]), .Z(n6447) );
  NANDN U7525 ( .A(x[147]), .B(y[147]), .Z(n6453) );
  AND U7526 ( .A(n6447), .B(n6453), .Z(n10473) );
  ANDN U7527 ( .B(x[145]), .A(y[145]), .Z(n6441) );
  ANDN U7528 ( .B(x[146]), .A(y[146]), .Z(n6452) );
  OR U7529 ( .A(n6441), .B(n6452), .Z(n10471) );
  NANDN U7530 ( .A(x[145]), .B(y[145]), .Z(n6444) );
  NANDN U7531 ( .A(x[144]), .B(y[144]), .Z(n3594) );
  AND U7532 ( .A(n6444), .B(n3594), .Z(n10469) );
  ANDN U7533 ( .B(x[143]), .A(y[143]), .Z(n6436) );
  ANDN U7534 ( .B(x[144]), .A(y[144]), .Z(n6442) );
  OR U7535 ( .A(n6436), .B(n6442), .Z(n10467) );
  NANDN U7536 ( .A(x[142]), .B(y[142]), .Z(n6432) );
  NANDN U7537 ( .A(x[143]), .B(y[143]), .Z(n5880) );
  AND U7538 ( .A(n6432), .B(n5880), .Z(n10465) );
  ANDN U7539 ( .B(x[141]), .A(y[141]), .Z(n6427) );
  ANDN U7540 ( .B(x[142]), .A(y[142]), .Z(n6437) );
  OR U7541 ( .A(n6427), .B(n6437), .Z(n10463) );
  NANDN U7542 ( .A(x[140]), .B(y[140]), .Z(n6424) );
  NANDN U7543 ( .A(x[141]), .B(y[141]), .Z(n6431) );
  AND U7544 ( .A(n6424), .B(n6431), .Z(n10461) );
  ANDN U7545 ( .B(x[139]), .A(y[139]), .Z(n6422) );
  ANDN U7546 ( .B(x[140]), .A(y[140]), .Z(n6430) );
  OR U7547 ( .A(n6422), .B(n6430), .Z(n10459) );
  NANDN U7548 ( .A(x[138]), .B(y[138]), .Z(n5882) );
  NANDN U7549 ( .A(x[139]), .B(y[139]), .Z(n6425) );
  AND U7550 ( .A(n5882), .B(n6425), .Z(n10457) );
  ANDN U7551 ( .B(x[137]), .A(y[137]), .Z(n6414) );
  ANDN U7552 ( .B(x[138]), .A(y[138]), .Z(n6419) );
  OR U7553 ( .A(n6414), .B(n6419), .Z(n10455) );
  NANDN U7554 ( .A(x[136]), .B(y[136]), .Z(n6410) );
  NANDN U7555 ( .A(x[137]), .B(y[137]), .Z(n5881) );
  AND U7556 ( .A(n6410), .B(n5881), .Z(n10453) );
  ANDN U7557 ( .B(x[135]), .A(y[135]), .Z(n6405) );
  ANDN U7558 ( .B(x[136]), .A(y[136]), .Z(n6415) );
  OR U7559 ( .A(n6405), .B(n6415), .Z(n10451) );
  NANDN U7560 ( .A(x[134]), .B(y[134]), .Z(n6402) );
  NANDN U7561 ( .A(x[135]), .B(y[135]), .Z(n6409) );
  AND U7562 ( .A(n6402), .B(n6409), .Z(n10449) );
  ANDN U7563 ( .B(x[133]), .A(y[133]), .Z(n6400) );
  ANDN U7564 ( .B(x[134]), .A(y[134]), .Z(n6408) );
  OR U7565 ( .A(n6400), .B(n6408), .Z(n10447) );
  NANDN U7566 ( .A(x[132]), .B(y[132]), .Z(n5884) );
  NANDN U7567 ( .A(x[133]), .B(y[133]), .Z(n6403) );
  AND U7568 ( .A(n5884), .B(n6403), .Z(n10445) );
  ANDN U7569 ( .B(x[131]), .A(y[131]), .Z(n6392) );
  ANDN U7570 ( .B(x[132]), .A(y[132]), .Z(n6397) );
  OR U7571 ( .A(n6392), .B(n6397), .Z(n10443) );
  NANDN U7572 ( .A(x[130]), .B(y[130]), .Z(n6388) );
  NANDN U7573 ( .A(x[131]), .B(y[131]), .Z(n5883) );
  AND U7574 ( .A(n6388), .B(n5883), .Z(n10441) );
  ANDN U7575 ( .B(x[129]), .A(y[129]), .Z(n6383) );
  ANDN U7576 ( .B(x[130]), .A(y[130]), .Z(n6393) );
  OR U7577 ( .A(n6383), .B(n6393), .Z(n10439) );
  NANDN U7578 ( .A(x[128]), .B(y[128]), .Z(n6381) );
  NANDN U7579 ( .A(x[129]), .B(y[129]), .Z(n6387) );
  AND U7580 ( .A(n6381), .B(n6387), .Z(n10437) );
  ANDN U7581 ( .B(x[127]), .A(y[127]), .Z(n5885) );
  ANDN U7582 ( .B(x[128]), .A(y[128]), .Z(n6386) );
  OR U7583 ( .A(n5885), .B(n6386), .Z(n10435) );
  NANDN U7584 ( .A(x[127]), .B(y[127]), .Z(n5888) );
  NANDN U7585 ( .A(x[126]), .B(y[126]), .Z(n3595) );
  AND U7586 ( .A(n5888), .B(n3595), .Z(n10433) );
  ANDN U7587 ( .B(x[125]), .A(y[125]), .Z(n6372) );
  ANDN U7588 ( .B(x[126]), .A(y[126]), .Z(n5886) );
  OR U7589 ( .A(n6372), .B(n5886), .Z(n10431) );
  NANDN U7590 ( .A(x[124]), .B(y[124]), .Z(n6369) );
  NANDN U7591 ( .A(x[125]), .B(y[125]), .Z(n6376) );
  AND U7592 ( .A(n6369), .B(n6376), .Z(n10429) );
  ANDN U7593 ( .B(x[123]), .A(y[123]), .Z(n6367) );
  ANDN U7594 ( .B(x[124]), .A(y[124]), .Z(n6375) );
  OR U7595 ( .A(n6367), .B(n6375), .Z(n10427) );
  NANDN U7596 ( .A(x[122]), .B(y[122]), .Z(n5890) );
  NANDN U7597 ( .A(x[123]), .B(y[123]), .Z(n6370) );
  AND U7598 ( .A(n5890), .B(n6370), .Z(n10425) );
  ANDN U7599 ( .B(x[121]), .A(y[121]), .Z(n6359) );
  ANDN U7600 ( .B(x[122]), .A(y[122]), .Z(n6364) );
  OR U7601 ( .A(n6359), .B(n6364), .Z(n10423) );
  NANDN U7602 ( .A(x[120]), .B(y[120]), .Z(n6355) );
  NANDN U7603 ( .A(x[121]), .B(y[121]), .Z(n5889) );
  AND U7604 ( .A(n6355), .B(n5889), .Z(n10421) );
  ANDN U7605 ( .B(x[119]), .A(y[119]), .Z(n6350) );
  ANDN U7606 ( .B(x[120]), .A(y[120]), .Z(n6360) );
  OR U7607 ( .A(n6350), .B(n6360), .Z(n10419) );
  NANDN U7608 ( .A(x[118]), .B(y[118]), .Z(n6347) );
  NANDN U7609 ( .A(x[119]), .B(y[119]), .Z(n6354) );
  AND U7610 ( .A(n6347), .B(n6354), .Z(n10417) );
  ANDN U7611 ( .B(x[117]), .A(y[117]), .Z(n6345) );
  ANDN U7612 ( .B(x[118]), .A(y[118]), .Z(n6353) );
  OR U7613 ( .A(n6345), .B(n6353), .Z(n10415) );
  NANDN U7614 ( .A(x[116]), .B(y[116]), .Z(n5892) );
  NANDN U7615 ( .A(x[117]), .B(y[117]), .Z(n6348) );
  AND U7616 ( .A(n5892), .B(n6348), .Z(n10413) );
  ANDN U7617 ( .B(x[115]), .A(y[115]), .Z(n6337) );
  ANDN U7618 ( .B(x[116]), .A(y[116]), .Z(n6342) );
  OR U7619 ( .A(n6337), .B(n6342), .Z(n10411) );
  NANDN U7620 ( .A(x[114]), .B(y[114]), .Z(n6333) );
  NANDN U7621 ( .A(x[115]), .B(y[115]), .Z(n5891) );
  AND U7622 ( .A(n6333), .B(n5891), .Z(n10409) );
  ANDN U7623 ( .B(x[113]), .A(y[113]), .Z(n6328) );
  ANDN U7624 ( .B(x[114]), .A(y[114]), .Z(n6338) );
  OR U7625 ( .A(n6328), .B(n6338), .Z(n10407) );
  NANDN U7626 ( .A(x[112]), .B(y[112]), .Z(n6325) );
  NANDN U7627 ( .A(x[113]), .B(y[113]), .Z(n6332) );
  AND U7628 ( .A(n6325), .B(n6332), .Z(n10405) );
  ANDN U7629 ( .B(x[111]), .A(y[111]), .Z(n6323) );
  ANDN U7630 ( .B(x[112]), .A(y[112]), .Z(n6331) );
  OR U7631 ( .A(n6323), .B(n6331), .Z(n10403) );
  NANDN U7632 ( .A(x[110]), .B(y[110]), .Z(n5894) );
  NANDN U7633 ( .A(x[111]), .B(y[111]), .Z(n6326) );
  AND U7634 ( .A(n5894), .B(n6326), .Z(n10401) );
  ANDN U7635 ( .B(x[109]), .A(y[109]), .Z(n6315) );
  ANDN U7636 ( .B(x[110]), .A(y[110]), .Z(n6320) );
  OR U7637 ( .A(n6315), .B(n6320), .Z(n10399) );
  NANDN U7638 ( .A(x[108]), .B(y[108]), .Z(n6311) );
  NANDN U7639 ( .A(x[109]), .B(y[109]), .Z(n5893) );
  AND U7640 ( .A(n6311), .B(n5893), .Z(n10397) );
  ANDN U7641 ( .B(x[107]), .A(y[107]), .Z(n6306) );
  ANDN U7642 ( .B(x[108]), .A(y[108]), .Z(n6316) );
  OR U7643 ( .A(n6306), .B(n6316), .Z(n10395) );
  NANDN U7644 ( .A(x[106]), .B(y[106]), .Z(n6303) );
  NANDN U7645 ( .A(x[107]), .B(y[107]), .Z(n6310) );
  AND U7646 ( .A(n6303), .B(n6310), .Z(n10393) );
  ANDN U7647 ( .B(x[105]), .A(y[105]), .Z(n6301) );
  ANDN U7648 ( .B(x[106]), .A(y[106]), .Z(n6309) );
  OR U7649 ( .A(n6301), .B(n6309), .Z(n10391) );
  NANDN U7650 ( .A(x[104]), .B(y[104]), .Z(n5896) );
  NANDN U7651 ( .A(x[105]), .B(y[105]), .Z(n6304) );
  AND U7652 ( .A(n5896), .B(n6304), .Z(n10389) );
  ANDN U7653 ( .B(x[103]), .A(y[103]), .Z(n6293) );
  ANDN U7654 ( .B(x[104]), .A(y[104]), .Z(n6298) );
  OR U7655 ( .A(n6293), .B(n6298), .Z(n10387) );
  NANDN U7656 ( .A(x[102]), .B(y[102]), .Z(n6289) );
  NANDN U7657 ( .A(x[103]), .B(y[103]), .Z(n5895) );
  AND U7658 ( .A(n6289), .B(n5895), .Z(n10385) );
  ANDN U7659 ( .B(x[101]), .A(y[101]), .Z(n6284) );
  ANDN U7660 ( .B(x[102]), .A(y[102]), .Z(n6294) );
  OR U7661 ( .A(n6284), .B(n6294), .Z(n10383) );
  NANDN U7662 ( .A(x[100]), .B(y[100]), .Z(n6281) );
  NANDN U7663 ( .A(x[101]), .B(y[101]), .Z(n6288) );
  AND U7664 ( .A(n6281), .B(n6288), .Z(n10381) );
  ANDN U7665 ( .B(x[99]), .A(y[99]), .Z(n6279) );
  ANDN U7666 ( .B(x[100]), .A(y[100]), .Z(n6287) );
  OR U7667 ( .A(n6279), .B(n6287), .Z(n10379) );
  NANDN U7668 ( .A(x[98]), .B(y[98]), .Z(n5898) );
  NANDN U7669 ( .A(x[99]), .B(y[99]), .Z(n6282) );
  AND U7670 ( .A(n5898), .B(n6282), .Z(n10377) );
  ANDN U7671 ( .B(x[97]), .A(y[97]), .Z(n6271) );
  ANDN U7672 ( .B(x[98]), .A(y[98]), .Z(n6276) );
  OR U7673 ( .A(n6271), .B(n6276), .Z(n10375) );
  NANDN U7674 ( .A(x[96]), .B(y[96]), .Z(n6267) );
  NANDN U7675 ( .A(x[97]), .B(y[97]), .Z(n5897) );
  AND U7676 ( .A(n6267), .B(n5897), .Z(n10373) );
  ANDN U7677 ( .B(x[95]), .A(y[95]), .Z(n6262) );
  ANDN U7678 ( .B(x[96]), .A(y[96]), .Z(n6272) );
  OR U7679 ( .A(n6262), .B(n6272), .Z(n10371) );
  NANDN U7680 ( .A(x[94]), .B(y[94]), .Z(n6259) );
  NANDN U7681 ( .A(x[95]), .B(y[95]), .Z(n6266) );
  AND U7682 ( .A(n6259), .B(n6266), .Z(n10369) );
  ANDN U7683 ( .B(x[93]), .A(y[93]), .Z(n6257) );
  ANDN U7684 ( .B(x[94]), .A(y[94]), .Z(n6265) );
  OR U7685 ( .A(n6257), .B(n6265), .Z(n10367) );
  NANDN U7686 ( .A(x[92]), .B(y[92]), .Z(n5900) );
  NANDN U7687 ( .A(x[93]), .B(y[93]), .Z(n6260) );
  AND U7688 ( .A(n5900), .B(n6260), .Z(n10365) );
  ANDN U7689 ( .B(x[91]), .A(y[91]), .Z(n6249) );
  ANDN U7690 ( .B(x[92]), .A(y[92]), .Z(n6254) );
  OR U7691 ( .A(n6249), .B(n6254), .Z(n10363) );
  NANDN U7692 ( .A(x[90]), .B(y[90]), .Z(n6245) );
  NANDN U7693 ( .A(x[91]), .B(y[91]), .Z(n5899) );
  AND U7694 ( .A(n6245), .B(n5899), .Z(n10361) );
  ANDN U7695 ( .B(x[89]), .A(y[89]), .Z(n6240) );
  ANDN U7696 ( .B(x[90]), .A(y[90]), .Z(n6250) );
  OR U7697 ( .A(n6240), .B(n6250), .Z(n10359) );
  NANDN U7698 ( .A(x[88]), .B(y[88]), .Z(n6237) );
  NANDN U7699 ( .A(x[89]), .B(y[89]), .Z(n6244) );
  AND U7700 ( .A(n6237), .B(n6244), .Z(n10357) );
  ANDN U7701 ( .B(x[87]), .A(y[87]), .Z(n6235) );
  ANDN U7702 ( .B(x[88]), .A(y[88]), .Z(n6243) );
  OR U7703 ( .A(n6235), .B(n6243), .Z(n10355) );
  NANDN U7704 ( .A(x[86]), .B(y[86]), .Z(n5902) );
  NANDN U7705 ( .A(x[87]), .B(y[87]), .Z(n6238) );
  AND U7706 ( .A(n5902), .B(n6238), .Z(n10353) );
  ANDN U7707 ( .B(x[85]), .A(y[85]), .Z(n6227) );
  ANDN U7708 ( .B(x[86]), .A(y[86]), .Z(n6232) );
  OR U7709 ( .A(n6227), .B(n6232), .Z(n10351) );
  NANDN U7710 ( .A(x[84]), .B(y[84]), .Z(n6223) );
  NANDN U7711 ( .A(x[85]), .B(y[85]), .Z(n5901) );
  AND U7712 ( .A(n6223), .B(n5901), .Z(n10349) );
  ANDN U7713 ( .B(x[83]), .A(y[83]), .Z(n6218) );
  ANDN U7714 ( .B(x[84]), .A(y[84]), .Z(n6228) );
  OR U7715 ( .A(n6218), .B(n6228), .Z(n10347) );
  NANDN U7716 ( .A(x[82]), .B(y[82]), .Z(n6215) );
  NANDN U7717 ( .A(x[83]), .B(y[83]), .Z(n6222) );
  AND U7718 ( .A(n6215), .B(n6222), .Z(n10345) );
  ANDN U7719 ( .B(x[81]), .A(y[81]), .Z(n6213) );
  ANDN U7720 ( .B(x[82]), .A(y[82]), .Z(n6221) );
  OR U7721 ( .A(n6213), .B(n6221), .Z(n10343) );
  NANDN U7722 ( .A(x[80]), .B(y[80]), .Z(n5904) );
  NANDN U7723 ( .A(x[81]), .B(y[81]), .Z(n6216) );
  AND U7724 ( .A(n5904), .B(n6216), .Z(n10341) );
  ANDN U7725 ( .B(x[79]), .A(y[79]), .Z(n6205) );
  ANDN U7726 ( .B(x[80]), .A(y[80]), .Z(n6210) );
  OR U7727 ( .A(n6205), .B(n6210), .Z(n10339) );
  NANDN U7728 ( .A(x[78]), .B(y[78]), .Z(n6203) );
  NANDN U7729 ( .A(x[79]), .B(y[79]), .Z(n5903) );
  AND U7730 ( .A(n6203), .B(n5903), .Z(n10337) );
  ANDN U7731 ( .B(x[77]), .A(y[77]), .Z(n6200) );
  ANDN U7732 ( .B(x[78]), .A(y[78]), .Z(n6206) );
  OR U7733 ( .A(n6200), .B(n6206), .Z(n10335) );
  NANDN U7734 ( .A(x[77]), .B(y[77]), .Z(n6199) );
  NANDN U7735 ( .A(x[76]), .B(y[76]), .Z(n3596) );
  AND U7736 ( .A(n6199), .B(n3596), .Z(n10333) );
  ANDN U7737 ( .B(x[75]), .A(y[75]), .Z(n6188) );
  NANDN U7738 ( .A(y[76]), .B(x[76]), .Z(n6197) );
  NANDN U7739 ( .A(n6188), .B(n6197), .Z(n10331) );
  NANDN U7740 ( .A(x[74]), .B(y[74]), .Z(n6185) );
  NANDN U7741 ( .A(x[75]), .B(y[75]), .Z(n6192) );
  AND U7742 ( .A(n6185), .B(n6192), .Z(n10329) );
  ANDN U7743 ( .B(x[73]), .A(y[73]), .Z(n6183) );
  ANDN U7744 ( .B(x[74]), .A(y[74]), .Z(n6191) );
  OR U7745 ( .A(n6183), .B(n6191), .Z(n10327) );
  NANDN U7746 ( .A(x[72]), .B(y[72]), .Z(n5906) );
  NANDN U7747 ( .A(x[73]), .B(y[73]), .Z(n6186) );
  AND U7748 ( .A(n5906), .B(n6186), .Z(n10325) );
  ANDN U7749 ( .B(x[71]), .A(y[71]), .Z(n6175) );
  ANDN U7750 ( .B(x[72]), .A(y[72]), .Z(n6180) );
  OR U7751 ( .A(n6175), .B(n6180), .Z(n10323) );
  NANDN U7752 ( .A(x[70]), .B(y[70]), .Z(n6171) );
  NANDN U7753 ( .A(x[71]), .B(y[71]), .Z(n5905) );
  AND U7754 ( .A(n6171), .B(n5905), .Z(n10321) );
  ANDN U7755 ( .B(x[69]), .A(y[69]), .Z(n6166) );
  ANDN U7756 ( .B(x[70]), .A(y[70]), .Z(n6176) );
  OR U7757 ( .A(n6166), .B(n6176), .Z(n10319) );
  NANDN U7758 ( .A(x[68]), .B(y[68]), .Z(n6163) );
  NANDN U7759 ( .A(x[69]), .B(y[69]), .Z(n6170) );
  AND U7760 ( .A(n6163), .B(n6170), .Z(n10317) );
  ANDN U7761 ( .B(x[67]), .A(y[67]), .Z(n6161) );
  ANDN U7762 ( .B(x[68]), .A(y[68]), .Z(n6169) );
  OR U7763 ( .A(n6161), .B(n6169), .Z(n10315) );
  NANDN U7764 ( .A(x[66]), .B(y[66]), .Z(n5908) );
  NANDN U7765 ( .A(x[67]), .B(y[67]), .Z(n6164) );
  AND U7766 ( .A(n5908), .B(n6164), .Z(n10313) );
  ANDN U7767 ( .B(x[65]), .A(y[65]), .Z(n6153) );
  ANDN U7768 ( .B(x[66]), .A(y[66]), .Z(n6158) );
  OR U7769 ( .A(n6153), .B(n6158), .Z(n10311) );
  NANDN U7770 ( .A(x[64]), .B(y[64]), .Z(n6149) );
  NANDN U7771 ( .A(x[65]), .B(y[65]), .Z(n5907) );
  AND U7772 ( .A(n6149), .B(n5907), .Z(n10309) );
  ANDN U7773 ( .B(x[63]), .A(y[63]), .Z(n6144) );
  ANDN U7774 ( .B(x[64]), .A(y[64]), .Z(n6154) );
  OR U7775 ( .A(n6144), .B(n6154), .Z(n10307) );
  NANDN U7776 ( .A(x[62]), .B(y[62]), .Z(n6141) );
  NANDN U7777 ( .A(x[63]), .B(y[63]), .Z(n6148) );
  AND U7778 ( .A(n6141), .B(n6148), .Z(n10305) );
  ANDN U7779 ( .B(x[61]), .A(y[61]), .Z(n6139) );
  ANDN U7780 ( .B(x[62]), .A(y[62]), .Z(n6147) );
  OR U7781 ( .A(n6139), .B(n6147), .Z(n10303) );
  NANDN U7782 ( .A(x[60]), .B(y[60]), .Z(n5910) );
  NANDN U7783 ( .A(x[61]), .B(y[61]), .Z(n6142) );
  AND U7784 ( .A(n5910), .B(n6142), .Z(n10301) );
  ANDN U7785 ( .B(x[59]), .A(y[59]), .Z(n6131) );
  ANDN U7786 ( .B(x[60]), .A(y[60]), .Z(n6136) );
  OR U7787 ( .A(n6131), .B(n6136), .Z(n10299) );
  NANDN U7788 ( .A(x[58]), .B(y[58]), .Z(n6127) );
  NANDN U7789 ( .A(x[59]), .B(y[59]), .Z(n5909) );
  AND U7790 ( .A(n6127), .B(n5909), .Z(n10297) );
  ANDN U7791 ( .B(x[57]), .A(y[57]), .Z(n6122) );
  ANDN U7792 ( .B(x[58]), .A(y[58]), .Z(n6132) );
  OR U7793 ( .A(n6122), .B(n6132), .Z(n10295) );
  NANDN U7794 ( .A(x[56]), .B(y[56]), .Z(n6119) );
  NANDN U7795 ( .A(x[57]), .B(y[57]), .Z(n6126) );
  AND U7796 ( .A(n6119), .B(n6126), .Z(n10293) );
  ANDN U7797 ( .B(x[55]), .A(y[55]), .Z(n6117) );
  ANDN U7798 ( .B(x[56]), .A(y[56]), .Z(n6125) );
  OR U7799 ( .A(n6117), .B(n6125), .Z(n10291) );
  NANDN U7800 ( .A(x[54]), .B(y[54]), .Z(n5912) );
  NANDN U7801 ( .A(x[55]), .B(y[55]), .Z(n6120) );
  AND U7802 ( .A(n5912), .B(n6120), .Z(n10289) );
  ANDN U7803 ( .B(x[53]), .A(y[53]), .Z(n6109) );
  ANDN U7804 ( .B(x[54]), .A(y[54]), .Z(n6114) );
  OR U7805 ( .A(n6109), .B(n6114), .Z(n10287) );
  NANDN U7806 ( .A(x[52]), .B(y[52]), .Z(n6105) );
  NANDN U7807 ( .A(x[53]), .B(y[53]), .Z(n5911) );
  AND U7808 ( .A(n6105), .B(n5911), .Z(n10285) );
  ANDN U7809 ( .B(x[51]), .A(y[51]), .Z(n6100) );
  ANDN U7810 ( .B(x[52]), .A(y[52]), .Z(n6110) );
  OR U7811 ( .A(n6100), .B(n6110), .Z(n10283) );
  NANDN U7812 ( .A(x[50]), .B(y[50]), .Z(n6097) );
  NANDN U7813 ( .A(x[51]), .B(y[51]), .Z(n6104) );
  AND U7814 ( .A(n6097), .B(n6104), .Z(n10281) );
  ANDN U7815 ( .B(x[49]), .A(y[49]), .Z(n6095) );
  ANDN U7816 ( .B(x[50]), .A(y[50]), .Z(n6103) );
  OR U7817 ( .A(n6095), .B(n6103), .Z(n10279) );
  NANDN U7818 ( .A(x[48]), .B(y[48]), .Z(n5914) );
  NANDN U7819 ( .A(x[49]), .B(y[49]), .Z(n6098) );
  AND U7820 ( .A(n5914), .B(n6098), .Z(n10277) );
  ANDN U7821 ( .B(x[47]), .A(y[47]), .Z(n6087) );
  ANDN U7822 ( .B(x[48]), .A(y[48]), .Z(n6092) );
  OR U7823 ( .A(n6087), .B(n6092), .Z(n10275) );
  NANDN U7824 ( .A(x[46]), .B(y[46]), .Z(n6083) );
  NANDN U7825 ( .A(x[47]), .B(y[47]), .Z(n5913) );
  AND U7826 ( .A(n6083), .B(n5913), .Z(n10273) );
  ANDN U7827 ( .B(x[45]), .A(y[45]), .Z(n6078) );
  ANDN U7828 ( .B(x[46]), .A(y[46]), .Z(n6088) );
  OR U7829 ( .A(n6078), .B(n6088), .Z(n10271) );
  NANDN U7830 ( .A(x[44]), .B(y[44]), .Z(n6075) );
  NANDN U7831 ( .A(x[45]), .B(y[45]), .Z(n6082) );
  AND U7832 ( .A(n6075), .B(n6082), .Z(n10269) );
  ANDN U7833 ( .B(x[43]), .A(y[43]), .Z(n6073) );
  ANDN U7834 ( .B(x[44]), .A(y[44]), .Z(n6081) );
  OR U7835 ( .A(n6073), .B(n6081), .Z(n10267) );
  NANDN U7836 ( .A(x[42]), .B(y[42]), .Z(n5916) );
  NANDN U7837 ( .A(x[43]), .B(y[43]), .Z(n6076) );
  AND U7838 ( .A(n5916), .B(n6076), .Z(n10265) );
  ANDN U7839 ( .B(x[41]), .A(y[41]), .Z(n6065) );
  ANDN U7840 ( .B(x[42]), .A(y[42]), .Z(n6070) );
  OR U7841 ( .A(n6065), .B(n6070), .Z(n10263) );
  NANDN U7842 ( .A(x[40]), .B(y[40]), .Z(n6061) );
  NANDN U7843 ( .A(x[41]), .B(y[41]), .Z(n5915) );
  AND U7844 ( .A(n6061), .B(n5915), .Z(n10261) );
  ANDN U7845 ( .B(x[39]), .A(y[39]), .Z(n6056) );
  ANDN U7846 ( .B(x[40]), .A(y[40]), .Z(n6066) );
  OR U7847 ( .A(n6056), .B(n6066), .Z(n10259) );
  NANDN U7848 ( .A(x[38]), .B(y[38]), .Z(n6053) );
  NANDN U7849 ( .A(x[39]), .B(y[39]), .Z(n6060) );
  AND U7850 ( .A(n6053), .B(n6060), .Z(n10257) );
  ANDN U7851 ( .B(x[37]), .A(y[37]), .Z(n6051) );
  ANDN U7852 ( .B(x[38]), .A(y[38]), .Z(n6059) );
  OR U7853 ( .A(n6051), .B(n6059), .Z(n10255) );
  NANDN U7854 ( .A(x[36]), .B(y[36]), .Z(n5918) );
  NANDN U7855 ( .A(x[37]), .B(y[37]), .Z(n6054) );
  AND U7856 ( .A(n5918), .B(n6054), .Z(n10253) );
  ANDN U7857 ( .B(x[35]), .A(y[35]), .Z(n6043) );
  ANDN U7858 ( .B(x[36]), .A(y[36]), .Z(n6048) );
  OR U7859 ( .A(n6043), .B(n6048), .Z(n10251) );
  NANDN U7860 ( .A(x[34]), .B(y[34]), .Z(n6039) );
  NANDN U7861 ( .A(x[35]), .B(y[35]), .Z(n5917) );
  AND U7862 ( .A(n6039), .B(n5917), .Z(n10249) );
  ANDN U7863 ( .B(x[33]), .A(y[33]), .Z(n6034) );
  ANDN U7864 ( .B(x[34]), .A(y[34]), .Z(n6044) );
  OR U7865 ( .A(n6034), .B(n6044), .Z(n10247) );
  NANDN U7866 ( .A(x[32]), .B(y[32]), .Z(n6031) );
  NANDN U7867 ( .A(x[33]), .B(y[33]), .Z(n6038) );
  AND U7868 ( .A(n6031), .B(n6038), .Z(n10245) );
  ANDN U7869 ( .B(x[31]), .A(y[31]), .Z(n6029) );
  ANDN U7870 ( .B(x[32]), .A(y[32]), .Z(n6037) );
  OR U7871 ( .A(n6029), .B(n6037), .Z(n10243) );
  NANDN U7872 ( .A(x[30]), .B(y[30]), .Z(n3597) );
  NANDN U7873 ( .A(x[31]), .B(y[31]), .Z(n6032) );
  AND U7874 ( .A(n3597), .B(n6032), .Z(n10241) );
  ANDN U7875 ( .B(x[29]), .A(y[29]), .Z(n6021) );
  XNOR U7876 ( .A(x[30]), .B(y[30]), .Z(n5919) );
  NANDN U7877 ( .A(n6021), .B(n5919), .Z(n10239) );
  NANDN U7878 ( .A(x[28]), .B(y[28]), .Z(n6017) );
  NANDN U7879 ( .A(x[29]), .B(y[29]), .Z(n5920) );
  AND U7880 ( .A(n6017), .B(n5920), .Z(n10237) );
  ANDN U7881 ( .B(x[27]), .A(y[27]), .Z(n6012) );
  ANDN U7882 ( .B(x[28]), .A(y[28]), .Z(n6022) );
  OR U7883 ( .A(n6012), .B(n6022), .Z(n10235) );
  NANDN U7884 ( .A(x[26]), .B(y[26]), .Z(n6009) );
  NANDN U7885 ( .A(x[27]), .B(y[27]), .Z(n6016) );
  AND U7886 ( .A(n6009), .B(n6016), .Z(n10233) );
  ANDN U7887 ( .B(x[25]), .A(y[25]), .Z(n6007) );
  ANDN U7888 ( .B(x[26]), .A(y[26]), .Z(n6015) );
  OR U7889 ( .A(n6007), .B(n6015), .Z(n10231) );
  NANDN U7890 ( .A(x[24]), .B(y[24]), .Z(n5922) );
  NANDN U7891 ( .A(x[25]), .B(y[25]), .Z(n6010) );
  AND U7892 ( .A(n5922), .B(n6010), .Z(n10229) );
  ANDN U7893 ( .B(x[23]), .A(y[23]), .Z(n5999) );
  ANDN U7894 ( .B(x[24]), .A(y[24]), .Z(n6004) );
  OR U7895 ( .A(n5999), .B(n6004), .Z(n10227) );
  NANDN U7896 ( .A(x[22]), .B(y[22]), .Z(n5995) );
  NANDN U7897 ( .A(x[23]), .B(y[23]), .Z(n5921) );
  AND U7898 ( .A(n5995), .B(n5921), .Z(n10225) );
  ANDN U7899 ( .B(x[21]), .A(y[21]), .Z(n5990) );
  ANDN U7900 ( .B(x[22]), .A(y[22]), .Z(n6000) );
  OR U7901 ( .A(n5990), .B(n6000), .Z(n10223) );
  NANDN U7902 ( .A(x[20]), .B(y[20]), .Z(n5987) );
  NANDN U7903 ( .A(x[21]), .B(y[21]), .Z(n5994) );
  AND U7904 ( .A(n5987), .B(n5994), .Z(n10221) );
  ANDN U7905 ( .B(x[19]), .A(y[19]), .Z(n5985) );
  ANDN U7906 ( .B(x[20]), .A(y[20]), .Z(n5993) );
  OR U7907 ( .A(n5985), .B(n5993), .Z(n10219) );
  NANDN U7908 ( .A(x[18]), .B(y[18]), .Z(n5924) );
  NANDN U7909 ( .A(x[19]), .B(y[19]), .Z(n5988) );
  AND U7910 ( .A(n5924), .B(n5988), .Z(n10217) );
  ANDN U7911 ( .B(x[17]), .A(y[17]), .Z(n5977) );
  ANDN U7912 ( .B(x[18]), .A(y[18]), .Z(n5982) );
  OR U7913 ( .A(n5977), .B(n5982), .Z(n10215) );
  NANDN U7914 ( .A(x[16]), .B(y[16]), .Z(n5973) );
  NANDN U7915 ( .A(x[17]), .B(y[17]), .Z(n5923) );
  AND U7916 ( .A(n5973), .B(n5923), .Z(n10213) );
  ANDN U7917 ( .B(x[15]), .A(y[15]), .Z(n5968) );
  ANDN U7918 ( .B(x[16]), .A(y[16]), .Z(n5978) );
  OR U7919 ( .A(n5968), .B(n5978), .Z(n10211) );
  NANDN U7920 ( .A(x[14]), .B(y[14]), .Z(n5965) );
  NANDN U7921 ( .A(x[15]), .B(y[15]), .Z(n5972) );
  AND U7922 ( .A(n5965), .B(n5972), .Z(n10209) );
  ANDN U7923 ( .B(x[13]), .A(y[13]), .Z(n5963) );
  ANDN U7924 ( .B(x[14]), .A(y[14]), .Z(n5971) );
  OR U7925 ( .A(n5963), .B(n5971), .Z(n10207) );
  NANDN U7926 ( .A(x[12]), .B(y[12]), .Z(n5926) );
  NANDN U7927 ( .A(x[13]), .B(y[13]), .Z(n5966) );
  AND U7928 ( .A(n5926), .B(n5966), .Z(n10205) );
  ANDN U7929 ( .B(x[11]), .A(y[11]), .Z(n5955) );
  ANDN U7930 ( .B(x[12]), .A(y[12]), .Z(n5960) );
  OR U7931 ( .A(n5955), .B(n5960), .Z(n10203) );
  NANDN U7932 ( .A(x[10]), .B(y[10]), .Z(n5951) );
  NANDN U7933 ( .A(x[11]), .B(y[11]), .Z(n5925) );
  AND U7934 ( .A(n5951), .B(n5925), .Z(n10201) );
  ANDN U7935 ( .B(x[9]), .A(y[9]), .Z(n5949) );
  ANDN U7936 ( .B(x[10]), .A(y[10]), .Z(n5956) );
  OR U7937 ( .A(n5949), .B(n5956), .Z(n10199) );
  NANDN U7938 ( .A(x[8]), .B(y[8]), .Z(n3598) );
  NANDN U7939 ( .A(x[9]), .B(y[9]), .Z(n5950) );
  AND U7940 ( .A(n3598), .B(n5950), .Z(n10197) );
  ANDN U7941 ( .B(x[7]), .A(y[7]), .Z(n5941) );
  XNOR U7942 ( .A(x[8]), .B(y[8]), .Z(n5943) );
  NANDN U7943 ( .A(n5941), .B(n5943), .Z(n10195) );
  NANDN U7944 ( .A(x[6]), .B(y[6]), .Z(n5939) );
  NANDN U7945 ( .A(x[7]), .B(y[7]), .Z(n5944) );
  AND U7946 ( .A(n5939), .B(n5944), .Z(n10193) );
  NANDN U7947 ( .A(y[4]), .B(x[4]), .Z(n3600) );
  NANDN U7948 ( .A(y[3]), .B(x[3]), .Z(n3599) );
  NAND U7949 ( .A(n3600), .B(n3599), .Z(n5934) );
  NANDN U7950 ( .A(x[2]), .B(y[2]), .Z(n3602) );
  NANDN U7951 ( .A(x[3]), .B(y[3]), .Z(n3601) );
  AND U7952 ( .A(n3602), .B(n3601), .Z(n5931) );
  NANDN U7953 ( .A(y[2]), .B(x[2]), .Z(n3604) );
  NANDN U7954 ( .A(y[1]), .B(x[1]), .Z(n3603) );
  NAND U7955 ( .A(n3604), .B(n3603), .Z(n5929) );
  NANDN U7956 ( .A(x[1]), .B(y[1]), .Z(n5927) );
  NANDN U7957 ( .A(x[4]), .B(y[4]), .Z(n3606) );
  NANDN U7958 ( .A(x[5]), .B(y[5]), .Z(n3605) );
  AND U7959 ( .A(n3606), .B(n3605), .Z(n5936) );
  NANDN U7960 ( .A(y[6]), .B(x[6]), .Z(n3608) );
  NANDN U7961 ( .A(y[5]), .B(x[5]), .Z(n3607) );
  NAND U7962 ( .A(n3608), .B(n3607), .Z(n5938) );
  OR U7963 ( .A(n10203), .B(n3609), .Z(n3610) );
  NAND U7964 ( .A(n10205), .B(n3610), .Z(n3611) );
  NANDN U7965 ( .A(n10207), .B(n3611), .Z(n3612) );
  NAND U7966 ( .A(n10209), .B(n3612), .Z(n3613) );
  NANDN U7967 ( .A(n10211), .B(n3613), .Z(n3614) );
  AND U7968 ( .A(n10213), .B(n3614), .Z(n3615) );
  OR U7969 ( .A(n10215), .B(n3615), .Z(n3616) );
  NAND U7970 ( .A(n10217), .B(n3616), .Z(n3617) );
  NANDN U7971 ( .A(n10219), .B(n3617), .Z(n3618) );
  NAND U7972 ( .A(n10221), .B(n3618), .Z(n3619) );
  NANDN U7973 ( .A(n10223), .B(n3619), .Z(n3620) );
  AND U7974 ( .A(n10225), .B(n3620), .Z(n3621) );
  OR U7975 ( .A(n10227), .B(n3621), .Z(n3622) );
  NAND U7976 ( .A(n10229), .B(n3622), .Z(n3623) );
  NANDN U7977 ( .A(n10231), .B(n3623), .Z(n3624) );
  NAND U7978 ( .A(n10233), .B(n3624), .Z(n3625) );
  NANDN U7979 ( .A(n10235), .B(n3625), .Z(n3626) );
  AND U7980 ( .A(n10237), .B(n3626), .Z(n3627) );
  OR U7981 ( .A(n10239), .B(n3627), .Z(n3628) );
  NAND U7982 ( .A(n10241), .B(n3628), .Z(n3629) );
  NANDN U7983 ( .A(n10243), .B(n3629), .Z(n3630) );
  NAND U7984 ( .A(n10245), .B(n3630), .Z(n3631) );
  NANDN U7985 ( .A(n10247), .B(n3631), .Z(n3632) );
  AND U7986 ( .A(n10249), .B(n3632), .Z(n3633) );
  OR U7987 ( .A(n10251), .B(n3633), .Z(n3634) );
  NAND U7988 ( .A(n10253), .B(n3634), .Z(n3635) );
  NANDN U7989 ( .A(n10255), .B(n3635), .Z(n3636) );
  NAND U7990 ( .A(n10257), .B(n3636), .Z(n3637) );
  NANDN U7991 ( .A(n10259), .B(n3637), .Z(n3638) );
  AND U7992 ( .A(n10261), .B(n3638), .Z(n3639) );
  OR U7993 ( .A(n10263), .B(n3639), .Z(n3640) );
  NAND U7994 ( .A(n10265), .B(n3640), .Z(n3641) );
  NANDN U7995 ( .A(n10267), .B(n3641), .Z(n3642) );
  NAND U7996 ( .A(n10269), .B(n3642), .Z(n3643) );
  NANDN U7997 ( .A(n10271), .B(n3643), .Z(n3644) );
  AND U7998 ( .A(n10273), .B(n3644), .Z(n3645) );
  OR U7999 ( .A(n10275), .B(n3645), .Z(n3646) );
  NAND U8000 ( .A(n10277), .B(n3646), .Z(n3647) );
  NANDN U8001 ( .A(n10279), .B(n3647), .Z(n3648) );
  NAND U8002 ( .A(n10281), .B(n3648), .Z(n3649) );
  NANDN U8003 ( .A(n10283), .B(n3649), .Z(n3650) );
  AND U8004 ( .A(n10285), .B(n3650), .Z(n3651) );
  OR U8005 ( .A(n10287), .B(n3651), .Z(n3652) );
  NAND U8006 ( .A(n10289), .B(n3652), .Z(n3653) );
  NANDN U8007 ( .A(n10291), .B(n3653), .Z(n3654) );
  NAND U8008 ( .A(n10293), .B(n3654), .Z(n3655) );
  NANDN U8009 ( .A(n10295), .B(n3655), .Z(n3656) );
  AND U8010 ( .A(n10297), .B(n3656), .Z(n3657) );
  OR U8011 ( .A(n10299), .B(n3657), .Z(n3658) );
  NAND U8012 ( .A(n10301), .B(n3658), .Z(n3659) );
  NANDN U8013 ( .A(n10303), .B(n3659), .Z(n3660) );
  NAND U8014 ( .A(n10305), .B(n3660), .Z(n3661) );
  NANDN U8015 ( .A(n10307), .B(n3661), .Z(n3662) );
  AND U8016 ( .A(n10309), .B(n3662), .Z(n3663) );
  OR U8017 ( .A(n10311), .B(n3663), .Z(n3664) );
  NAND U8018 ( .A(n10313), .B(n3664), .Z(n3665) );
  NANDN U8019 ( .A(n10315), .B(n3665), .Z(n3666) );
  NAND U8020 ( .A(n10317), .B(n3666), .Z(n3667) );
  NANDN U8021 ( .A(n10319), .B(n3667), .Z(n3668) );
  AND U8022 ( .A(n10321), .B(n3668), .Z(n3669) );
  OR U8023 ( .A(n10323), .B(n3669), .Z(n3670) );
  NAND U8024 ( .A(n10325), .B(n3670), .Z(n3671) );
  NANDN U8025 ( .A(n10327), .B(n3671), .Z(n3672) );
  NAND U8026 ( .A(n10329), .B(n3672), .Z(n3673) );
  NANDN U8027 ( .A(n10331), .B(n3673), .Z(n3674) );
  AND U8028 ( .A(n10333), .B(n3674), .Z(n3675) );
  OR U8029 ( .A(n10335), .B(n3675), .Z(n3676) );
  NAND U8030 ( .A(n10337), .B(n3676), .Z(n3677) );
  NANDN U8031 ( .A(n10339), .B(n3677), .Z(n3678) );
  NAND U8032 ( .A(n10341), .B(n3678), .Z(n3679) );
  NANDN U8033 ( .A(n10343), .B(n3679), .Z(n3680) );
  AND U8034 ( .A(n10345), .B(n3680), .Z(n3681) );
  OR U8035 ( .A(n10347), .B(n3681), .Z(n3682) );
  NAND U8036 ( .A(n10349), .B(n3682), .Z(n3683) );
  NANDN U8037 ( .A(n10351), .B(n3683), .Z(n3684) );
  NAND U8038 ( .A(n10353), .B(n3684), .Z(n3685) );
  NANDN U8039 ( .A(n10355), .B(n3685), .Z(n3686) );
  AND U8040 ( .A(n10357), .B(n3686), .Z(n3687) );
  OR U8041 ( .A(n10359), .B(n3687), .Z(n3688) );
  NAND U8042 ( .A(n10361), .B(n3688), .Z(n3689) );
  NANDN U8043 ( .A(n10363), .B(n3689), .Z(n3690) );
  NAND U8044 ( .A(n10365), .B(n3690), .Z(n3691) );
  NANDN U8045 ( .A(n10367), .B(n3691), .Z(n3692) );
  AND U8046 ( .A(n10369), .B(n3692), .Z(n3693) );
  OR U8047 ( .A(n10371), .B(n3693), .Z(n3694) );
  NAND U8048 ( .A(n10373), .B(n3694), .Z(n3695) );
  NANDN U8049 ( .A(n10375), .B(n3695), .Z(n3696) );
  NAND U8050 ( .A(n10377), .B(n3696), .Z(n3697) );
  NANDN U8051 ( .A(n10379), .B(n3697), .Z(n3698) );
  AND U8052 ( .A(n10381), .B(n3698), .Z(n3699) );
  OR U8053 ( .A(n10383), .B(n3699), .Z(n3700) );
  NAND U8054 ( .A(n10385), .B(n3700), .Z(n3701) );
  NANDN U8055 ( .A(n10387), .B(n3701), .Z(n3702) );
  NAND U8056 ( .A(n10389), .B(n3702), .Z(n3703) );
  NANDN U8057 ( .A(n10391), .B(n3703), .Z(n3704) );
  AND U8058 ( .A(n10393), .B(n3704), .Z(n3705) );
  OR U8059 ( .A(n10395), .B(n3705), .Z(n3706) );
  NAND U8060 ( .A(n10397), .B(n3706), .Z(n3707) );
  NANDN U8061 ( .A(n10399), .B(n3707), .Z(n3708) );
  NAND U8062 ( .A(n10401), .B(n3708), .Z(n3709) );
  NANDN U8063 ( .A(n10403), .B(n3709), .Z(n3710) );
  AND U8064 ( .A(n10405), .B(n3710), .Z(n3711) );
  OR U8065 ( .A(n10407), .B(n3711), .Z(n3712) );
  NAND U8066 ( .A(n10409), .B(n3712), .Z(n3713) );
  NANDN U8067 ( .A(n10411), .B(n3713), .Z(n3714) );
  NAND U8068 ( .A(n10413), .B(n3714), .Z(n3715) );
  NANDN U8069 ( .A(n10415), .B(n3715), .Z(n3716) );
  AND U8070 ( .A(n10417), .B(n3716), .Z(n3717) );
  OR U8071 ( .A(n10419), .B(n3717), .Z(n3718) );
  NAND U8072 ( .A(n10421), .B(n3718), .Z(n3719) );
  NANDN U8073 ( .A(n10423), .B(n3719), .Z(n3720) );
  NAND U8074 ( .A(n10425), .B(n3720), .Z(n3721) );
  NANDN U8075 ( .A(n10427), .B(n3721), .Z(n3722) );
  AND U8076 ( .A(n10429), .B(n3722), .Z(n3723) );
  OR U8077 ( .A(n10431), .B(n3723), .Z(n3724) );
  NAND U8078 ( .A(n10433), .B(n3724), .Z(n3725) );
  NANDN U8079 ( .A(n10435), .B(n3725), .Z(n3726) );
  NAND U8080 ( .A(n10437), .B(n3726), .Z(n3727) );
  NANDN U8081 ( .A(n10439), .B(n3727), .Z(n3728) );
  AND U8082 ( .A(n10441), .B(n3728), .Z(n3729) );
  OR U8083 ( .A(n10443), .B(n3729), .Z(n3730) );
  NAND U8084 ( .A(n10445), .B(n3730), .Z(n3731) );
  NANDN U8085 ( .A(n10447), .B(n3731), .Z(n3732) );
  NAND U8086 ( .A(n10449), .B(n3732), .Z(n3733) );
  NANDN U8087 ( .A(n10451), .B(n3733), .Z(n3734) );
  AND U8088 ( .A(n10453), .B(n3734), .Z(n3735) );
  OR U8089 ( .A(n10455), .B(n3735), .Z(n3736) );
  NAND U8090 ( .A(n10457), .B(n3736), .Z(n3737) );
  NANDN U8091 ( .A(n10459), .B(n3737), .Z(n3738) );
  NAND U8092 ( .A(n10461), .B(n3738), .Z(n3739) );
  NANDN U8093 ( .A(n10463), .B(n3739), .Z(n3740) );
  AND U8094 ( .A(n10465), .B(n3740), .Z(n3741) );
  OR U8095 ( .A(n10467), .B(n3741), .Z(n3742) );
  NAND U8096 ( .A(n10469), .B(n3742), .Z(n3743) );
  NANDN U8097 ( .A(n10471), .B(n3743), .Z(n3744) );
  NAND U8098 ( .A(n10473), .B(n3744), .Z(n3745) );
  NANDN U8099 ( .A(n10475), .B(n3745), .Z(n3746) );
  AND U8100 ( .A(n10477), .B(n3746), .Z(n3747) );
  OR U8101 ( .A(n10479), .B(n3747), .Z(n3748) );
  NAND U8102 ( .A(n10481), .B(n3748), .Z(n3749) );
  NANDN U8103 ( .A(n10483), .B(n3749), .Z(n3750) );
  NAND U8104 ( .A(n10485), .B(n3750), .Z(n3751) );
  NAND U8105 ( .A(n10486), .B(n3751), .Z(n3754) );
  NANDN U8106 ( .A(x[155]), .B(y[155]), .Z(n3753) );
  NANDN U8107 ( .A(x[154]), .B(y[154]), .Z(n3752) );
  NAND U8108 ( .A(n3753), .B(n3752), .Z(n10489) );
  ANDN U8109 ( .B(n3754), .A(n10489), .Z(n3755) );
  OR U8110 ( .A(n10491), .B(n3755), .Z(n3756) );
  NAND U8111 ( .A(n10493), .B(n3756), .Z(n3757) );
  NANDN U8112 ( .A(n10495), .B(n3757), .Z(n3758) );
  NAND U8113 ( .A(n10497), .B(n3758), .Z(n3759) );
  NANDN U8114 ( .A(n10499), .B(n3759), .Z(n3760) );
  AND U8115 ( .A(n10501), .B(n3760), .Z(n3761) );
  OR U8116 ( .A(n10503), .B(n3761), .Z(n3762) );
  NAND U8117 ( .A(n10505), .B(n3762), .Z(n3763) );
  NANDN U8118 ( .A(n10507), .B(n3763), .Z(n3764) );
  NAND U8119 ( .A(n10509), .B(n3764), .Z(n3765) );
  NANDN U8120 ( .A(n10511), .B(n3765), .Z(n3766) );
  AND U8121 ( .A(n10513), .B(n3766), .Z(n3767) );
  OR U8122 ( .A(n10515), .B(n3767), .Z(n3768) );
  NAND U8123 ( .A(n10517), .B(n3768), .Z(n3769) );
  NANDN U8124 ( .A(n10519), .B(n3769), .Z(n3770) );
  NAND U8125 ( .A(n10521), .B(n3770), .Z(n3771) );
  NANDN U8126 ( .A(n10523), .B(n3771), .Z(n3772) );
  AND U8127 ( .A(n10525), .B(n3772), .Z(n3773) );
  OR U8128 ( .A(n10527), .B(n3773), .Z(n3774) );
  NAND U8129 ( .A(n10529), .B(n3774), .Z(n3775) );
  NANDN U8130 ( .A(n10531), .B(n3775), .Z(n3776) );
  NAND U8131 ( .A(n10533), .B(n3776), .Z(n3777) );
  NANDN U8132 ( .A(n10535), .B(n3777), .Z(n3778) );
  AND U8133 ( .A(n10537), .B(n3778), .Z(n3779) );
  OR U8134 ( .A(n10539), .B(n3779), .Z(n3780) );
  NAND U8135 ( .A(n10541), .B(n3780), .Z(n3781) );
  NANDN U8136 ( .A(n10543), .B(n3781), .Z(n3782) );
  NAND U8137 ( .A(n10545), .B(n3782), .Z(n3783) );
  NANDN U8138 ( .A(n10547), .B(n3783), .Z(n3784) );
  AND U8139 ( .A(n10549), .B(n3784), .Z(n3785) );
  OR U8140 ( .A(n10551), .B(n3785), .Z(n3786) );
  NAND U8141 ( .A(n10553), .B(n3786), .Z(n3787) );
  NANDN U8142 ( .A(n10555), .B(n3787), .Z(n3788) );
  NAND U8143 ( .A(n10557), .B(n3788), .Z(n3789) );
  NANDN U8144 ( .A(n10559), .B(n3789), .Z(n3790) );
  AND U8145 ( .A(n10561), .B(n3790), .Z(n3791) );
  OR U8146 ( .A(n10563), .B(n3791), .Z(n3792) );
  NAND U8147 ( .A(n10565), .B(n3792), .Z(n3793) );
  NANDN U8148 ( .A(n10567), .B(n3793), .Z(n3794) );
  NAND U8149 ( .A(n10569), .B(n3794), .Z(n3795) );
  NANDN U8150 ( .A(n10571), .B(n3795), .Z(n3796) );
  AND U8151 ( .A(n10573), .B(n3796), .Z(n3797) );
  OR U8152 ( .A(n10575), .B(n3797), .Z(n3798) );
  NAND U8153 ( .A(n10577), .B(n3798), .Z(n3799) );
  NANDN U8154 ( .A(n10579), .B(n3799), .Z(n3800) );
  NAND U8155 ( .A(n10581), .B(n3800), .Z(n3801) );
  NANDN U8156 ( .A(n10583), .B(n3801), .Z(n3802) );
  AND U8157 ( .A(n10585), .B(n3802), .Z(n3803) );
  OR U8158 ( .A(n10587), .B(n3803), .Z(n3804) );
  NAND U8159 ( .A(n10589), .B(n3804), .Z(n3805) );
  NANDN U8160 ( .A(n10591), .B(n3805), .Z(n3806) );
  NAND U8161 ( .A(n10593), .B(n3806), .Z(n3807) );
  NANDN U8162 ( .A(n10595), .B(n3807), .Z(n3808) );
  AND U8163 ( .A(n10597), .B(n3808), .Z(n3809) );
  OR U8164 ( .A(n10599), .B(n3809), .Z(n3810) );
  NAND U8165 ( .A(n10601), .B(n3810), .Z(n3811) );
  NANDN U8166 ( .A(n10603), .B(n3811), .Z(n3812) );
  NAND U8167 ( .A(n10605), .B(n3812), .Z(n3813) );
  NANDN U8168 ( .A(n10607), .B(n3813), .Z(n3814) );
  AND U8169 ( .A(n10609), .B(n3814), .Z(n3815) );
  OR U8170 ( .A(n10611), .B(n3815), .Z(n3816) );
  NAND U8171 ( .A(n10613), .B(n3816), .Z(n3817) );
  NANDN U8172 ( .A(n10615), .B(n3817), .Z(n3818) );
  NAND U8173 ( .A(n10617), .B(n3818), .Z(n3819) );
  NANDN U8174 ( .A(n10619), .B(n3819), .Z(n3820) );
  AND U8175 ( .A(n10621), .B(n3820), .Z(n3821) );
  OR U8176 ( .A(n10623), .B(n3821), .Z(n3822) );
  NAND U8177 ( .A(n10625), .B(n3822), .Z(n3823) );
  NANDN U8178 ( .A(n10627), .B(n3823), .Z(n3824) );
  NAND U8179 ( .A(n10629), .B(n3824), .Z(n3825) );
  NANDN U8180 ( .A(n10631), .B(n3825), .Z(n3826) );
  AND U8181 ( .A(n10633), .B(n3826), .Z(n3827) );
  OR U8182 ( .A(n10635), .B(n3827), .Z(n3828) );
  NAND U8183 ( .A(n10637), .B(n3828), .Z(n3829) );
  NANDN U8184 ( .A(n10639), .B(n3829), .Z(n3830) );
  NAND U8185 ( .A(n10641), .B(n3830), .Z(n3831) );
  NANDN U8186 ( .A(n10643), .B(n3831), .Z(n3832) );
  AND U8187 ( .A(n10645), .B(n3832), .Z(n3833) );
  OR U8188 ( .A(n10647), .B(n3833), .Z(n3834) );
  NAND U8189 ( .A(n10649), .B(n3834), .Z(n3835) );
  NANDN U8190 ( .A(n10651), .B(n3835), .Z(n3836) );
  NAND U8191 ( .A(n10653), .B(n3836), .Z(n3837) );
  NANDN U8192 ( .A(n10655), .B(n3837), .Z(n3838) );
  AND U8193 ( .A(n10657), .B(n3838), .Z(n3839) );
  OR U8194 ( .A(n10659), .B(n3839), .Z(n3840) );
  NAND U8195 ( .A(n10661), .B(n3840), .Z(n3841) );
  NANDN U8196 ( .A(n10663), .B(n3841), .Z(n3842) );
  NAND U8197 ( .A(n10665), .B(n3842), .Z(n3843) );
  NANDN U8198 ( .A(n10667), .B(n3843), .Z(n3844) );
  AND U8199 ( .A(n10669), .B(n3844), .Z(n3845) );
  OR U8200 ( .A(n10671), .B(n3845), .Z(n3846) );
  NAND U8201 ( .A(n10673), .B(n3846), .Z(n3847) );
  NANDN U8202 ( .A(n10675), .B(n3847), .Z(n3848) );
  NAND U8203 ( .A(n10677), .B(n3848), .Z(n3849) );
  NANDN U8204 ( .A(n10679), .B(n3849), .Z(n3850) );
  AND U8205 ( .A(n10681), .B(n3850), .Z(n3851) );
  OR U8206 ( .A(n10683), .B(n3851), .Z(n3852) );
  NAND U8207 ( .A(n10685), .B(n3852), .Z(n3853) );
  NANDN U8208 ( .A(n10687), .B(n3853), .Z(n3854) );
  NAND U8209 ( .A(n10689), .B(n3854), .Z(n3855) );
  NANDN U8210 ( .A(n10691), .B(n3855), .Z(n3856) );
  AND U8211 ( .A(n10693), .B(n3856), .Z(n3857) );
  OR U8212 ( .A(n10695), .B(n3857), .Z(n3858) );
  NAND U8213 ( .A(n10697), .B(n3858), .Z(n3859) );
  NANDN U8214 ( .A(n10699), .B(n3859), .Z(n3860) );
  NAND U8215 ( .A(n10701), .B(n3860), .Z(n3861) );
  NANDN U8216 ( .A(n10703), .B(n3861), .Z(n3862) );
  AND U8217 ( .A(n10705), .B(n3862), .Z(n3863) );
  OR U8218 ( .A(n10707), .B(n3863), .Z(n3864) );
  NAND U8219 ( .A(n10709), .B(n3864), .Z(n3865) );
  NANDN U8220 ( .A(n10711), .B(n3865), .Z(n3866) );
  NAND U8221 ( .A(n10713), .B(n3866), .Z(n3867) );
  NANDN U8222 ( .A(n10715), .B(n3867), .Z(n3868) );
  AND U8223 ( .A(n10717), .B(n3868), .Z(n3869) );
  OR U8224 ( .A(n10719), .B(n3869), .Z(n3870) );
  NAND U8225 ( .A(n10721), .B(n3870), .Z(n3871) );
  NANDN U8226 ( .A(n10723), .B(n3871), .Z(n3872) );
  NAND U8227 ( .A(n10725), .B(n3872), .Z(n3873) );
  NANDN U8228 ( .A(n10727), .B(n3873), .Z(n3874) );
  AND U8229 ( .A(n10729), .B(n3874), .Z(n3875) );
  OR U8230 ( .A(n10731), .B(n3875), .Z(n3876) );
  NAND U8231 ( .A(n10733), .B(n3876), .Z(n3877) );
  NANDN U8232 ( .A(n10735), .B(n3877), .Z(n3878) );
  NAND U8233 ( .A(n10737), .B(n3878), .Z(n3879) );
  ANDN U8234 ( .B(x[280]), .A(y[280]), .Z(n6901) );
  ANDN U8235 ( .B(n3879), .A(n6901), .Z(n3880) );
  NANDN U8236 ( .A(n10738), .B(n3880), .Z(n3881) );
  NAND U8237 ( .A(n10743), .B(n3881), .Z(n3882) );
  NANDN U8238 ( .A(n10745), .B(n3882), .Z(n3883) );
  AND U8239 ( .A(n10747), .B(n3883), .Z(n3884) );
  OR U8240 ( .A(n10749), .B(n3884), .Z(n3885) );
  NAND U8241 ( .A(n10751), .B(n3885), .Z(n3886) );
  NANDN U8242 ( .A(n10753), .B(n3886), .Z(n3887) );
  NAND U8243 ( .A(n10755), .B(n3887), .Z(n3888) );
  NANDN U8244 ( .A(n10757), .B(n3888), .Z(n3889) );
  AND U8245 ( .A(n10759), .B(n3889), .Z(n3890) );
  OR U8246 ( .A(n10761), .B(n3890), .Z(n3891) );
  NAND U8247 ( .A(n10763), .B(n3891), .Z(n3892) );
  NANDN U8248 ( .A(n10765), .B(n3892), .Z(n3893) );
  NAND U8249 ( .A(n10767), .B(n3893), .Z(n3894) );
  NANDN U8250 ( .A(n10769), .B(n3894), .Z(n3895) );
  AND U8251 ( .A(n10771), .B(n3895), .Z(n3896) );
  OR U8252 ( .A(n10773), .B(n3896), .Z(n3897) );
  NAND U8253 ( .A(n10775), .B(n3897), .Z(n3898) );
  NANDN U8254 ( .A(n10777), .B(n3898), .Z(n3899) );
  NAND U8255 ( .A(n10779), .B(n3899), .Z(n3900) );
  NANDN U8256 ( .A(n10781), .B(n3900), .Z(n3901) );
  AND U8257 ( .A(n10783), .B(n3901), .Z(n3902) );
  OR U8258 ( .A(n10785), .B(n3902), .Z(n3903) );
  NAND U8259 ( .A(n10787), .B(n3903), .Z(n3904) );
  NANDN U8260 ( .A(n10789), .B(n3904), .Z(n3905) );
  NAND U8261 ( .A(n10791), .B(n3905), .Z(n3906) );
  NANDN U8262 ( .A(n10793), .B(n3906), .Z(n3907) );
  AND U8263 ( .A(n10795), .B(n3907), .Z(n3908) );
  OR U8264 ( .A(n10797), .B(n3908), .Z(n3909) );
  NAND U8265 ( .A(n10799), .B(n3909), .Z(n3910) );
  NANDN U8266 ( .A(n10801), .B(n3910), .Z(n3911) );
  NAND U8267 ( .A(n10803), .B(n3911), .Z(n3912) );
  NANDN U8268 ( .A(n10805), .B(n3912), .Z(n3913) );
  AND U8269 ( .A(n10807), .B(n3913), .Z(n3914) );
  OR U8270 ( .A(n10809), .B(n3914), .Z(n3915) );
  NAND U8271 ( .A(n10811), .B(n3915), .Z(n3916) );
  NANDN U8272 ( .A(n10813), .B(n3916), .Z(n3917) );
  NAND U8273 ( .A(n10815), .B(n3917), .Z(n3918) );
  NANDN U8274 ( .A(n10817), .B(n3918), .Z(n3919) );
  AND U8275 ( .A(n10819), .B(n3919), .Z(n3920) );
  OR U8276 ( .A(n10821), .B(n3920), .Z(n3921) );
  NAND U8277 ( .A(n10823), .B(n3921), .Z(n3922) );
  NANDN U8278 ( .A(n10825), .B(n3922), .Z(n3923) );
  NAND U8279 ( .A(n10827), .B(n3923), .Z(n3924) );
  NANDN U8280 ( .A(n10829), .B(n3924), .Z(n3925) );
  AND U8281 ( .A(n10831), .B(n3925), .Z(n3926) );
  OR U8282 ( .A(n10833), .B(n3926), .Z(n3927) );
  NAND U8283 ( .A(n10835), .B(n3927), .Z(n3928) );
  NANDN U8284 ( .A(n10837), .B(n3928), .Z(n3929) );
  NAND U8285 ( .A(n10839), .B(n3929), .Z(n3930) );
  NANDN U8286 ( .A(n10841), .B(n3930), .Z(n3931) );
  AND U8287 ( .A(n10843), .B(n3931), .Z(n3932) );
  OR U8288 ( .A(n10845), .B(n3932), .Z(n3933) );
  NAND U8289 ( .A(n10847), .B(n3933), .Z(n3934) );
  NANDN U8290 ( .A(n10849), .B(n3934), .Z(n3935) );
  NAND U8291 ( .A(n10851), .B(n3935), .Z(n3936) );
  NANDN U8292 ( .A(n10853), .B(n3936), .Z(n3937) );
  AND U8293 ( .A(n10855), .B(n3937), .Z(n3938) );
  OR U8294 ( .A(n10857), .B(n3938), .Z(n3939) );
  NAND U8295 ( .A(n10859), .B(n3939), .Z(n3940) );
  NANDN U8296 ( .A(n10861), .B(n3940), .Z(n3941) );
  NAND U8297 ( .A(n10863), .B(n3941), .Z(n3942) );
  NANDN U8298 ( .A(n10865), .B(n3942), .Z(n3943) );
  AND U8299 ( .A(n10867), .B(n3943), .Z(n3944) );
  OR U8300 ( .A(n10869), .B(n3944), .Z(n3945) );
  NAND U8301 ( .A(n10871), .B(n3945), .Z(n3946) );
  NANDN U8302 ( .A(n10873), .B(n3946), .Z(n3947) );
  NAND U8303 ( .A(n10875), .B(n3947), .Z(n3948) );
  NANDN U8304 ( .A(n10877), .B(n3948), .Z(n3949) );
  AND U8305 ( .A(n10879), .B(n3949), .Z(n3950) );
  OR U8306 ( .A(n10881), .B(n3950), .Z(n3951) );
  NAND U8307 ( .A(n10883), .B(n3951), .Z(n3952) );
  NANDN U8308 ( .A(n10885), .B(n3952), .Z(n3953) );
  NAND U8309 ( .A(n10887), .B(n3953), .Z(n3954) );
  NANDN U8310 ( .A(n10889), .B(n3954), .Z(n3955) );
  AND U8311 ( .A(n10891), .B(n3955), .Z(n3956) );
  OR U8312 ( .A(n10893), .B(n3956), .Z(n3957) );
  NAND U8313 ( .A(n10895), .B(n3957), .Z(n3958) );
  NANDN U8314 ( .A(n10897), .B(n3958), .Z(n3959) );
  NAND U8315 ( .A(n10899), .B(n3959), .Z(n3960) );
  NANDN U8316 ( .A(n10901), .B(n3960), .Z(n3961) );
  AND U8317 ( .A(n10903), .B(n3961), .Z(n3962) );
  OR U8318 ( .A(n10905), .B(n3962), .Z(n3963) );
  NAND U8319 ( .A(n10907), .B(n3963), .Z(n3964) );
  NANDN U8320 ( .A(n10909), .B(n3964), .Z(n3965) );
  NAND U8321 ( .A(n10911), .B(n3965), .Z(n3966) );
  NANDN U8322 ( .A(n10913), .B(n3966), .Z(n3967) );
  AND U8323 ( .A(n10915), .B(n3967), .Z(n3968) );
  OR U8324 ( .A(n10917), .B(n3968), .Z(n3969) );
  NAND U8325 ( .A(n10919), .B(n3969), .Z(n3970) );
  NANDN U8326 ( .A(n10921), .B(n3970), .Z(n3971) );
  NAND U8327 ( .A(n10923), .B(n3971), .Z(n3972) );
  NANDN U8328 ( .A(n10925), .B(n3972), .Z(n3973) );
  AND U8329 ( .A(n10927), .B(n3973), .Z(n3974) );
  OR U8330 ( .A(n10929), .B(n3974), .Z(n3975) );
  NAND U8331 ( .A(n10931), .B(n3975), .Z(n3976) );
  NANDN U8332 ( .A(n10933), .B(n3976), .Z(n3977) );
  NAND U8333 ( .A(n10935), .B(n3977), .Z(n3978) );
  NANDN U8334 ( .A(n10937), .B(n3978), .Z(n3979) );
  AND U8335 ( .A(n10939), .B(n3979), .Z(n3980) );
  OR U8336 ( .A(n10941), .B(n3980), .Z(n3981) );
  NAND U8337 ( .A(n10943), .B(n3981), .Z(n3982) );
  NANDN U8338 ( .A(n10945), .B(n3982), .Z(n3983) );
  NAND U8339 ( .A(n10947), .B(n3983), .Z(n3984) );
  NANDN U8340 ( .A(n10949), .B(n3984), .Z(n3985) );
  AND U8341 ( .A(n10951), .B(n3985), .Z(n3986) );
  OR U8342 ( .A(n10953), .B(n3986), .Z(n3987) );
  NAND U8343 ( .A(n10955), .B(n3987), .Z(n3988) );
  NANDN U8344 ( .A(n10957), .B(n3988), .Z(n3989) );
  NAND U8345 ( .A(n10959), .B(n3989), .Z(n3990) );
  NANDN U8346 ( .A(n10961), .B(n3990), .Z(n3991) );
  AND U8347 ( .A(n10963), .B(n3991), .Z(n3992) );
  OR U8348 ( .A(n10965), .B(n3992), .Z(n3993) );
  NAND U8349 ( .A(n10967), .B(n3993), .Z(n3994) );
  NANDN U8350 ( .A(n10969), .B(n3994), .Z(n3995) );
  NAND U8351 ( .A(n10971), .B(n3995), .Z(n3996) );
  NANDN U8352 ( .A(n10973), .B(n3996), .Z(n3997) );
  AND U8353 ( .A(n10975), .B(n3997), .Z(n3998) );
  OR U8354 ( .A(n10977), .B(n3998), .Z(n3999) );
  NAND U8355 ( .A(n10979), .B(n3999), .Z(n4000) );
  NANDN U8356 ( .A(n10981), .B(n4000), .Z(n4001) );
  NAND U8357 ( .A(n10983), .B(n4001), .Z(n4002) );
  NANDN U8358 ( .A(n10985), .B(n4002), .Z(n4003) );
  AND U8359 ( .A(n10987), .B(n4003), .Z(n4004) );
  OR U8360 ( .A(n10989), .B(n4004), .Z(n4005) );
  NAND U8361 ( .A(n10991), .B(n4005), .Z(n4006) );
  NANDN U8362 ( .A(n10993), .B(n4006), .Z(n4007) );
  NAND U8363 ( .A(n10995), .B(n4007), .Z(n4008) );
  NANDN U8364 ( .A(n10997), .B(n4008), .Z(n4009) );
  AND U8365 ( .A(n10999), .B(n4009), .Z(n4010) );
  OR U8366 ( .A(n11001), .B(n4010), .Z(n4011) );
  NAND U8367 ( .A(n11003), .B(n4011), .Z(n4012) );
  NANDN U8368 ( .A(n11005), .B(n4012), .Z(n4013) );
  NAND U8369 ( .A(n11007), .B(n4013), .Z(n4014) );
  NANDN U8370 ( .A(n11009), .B(n4014), .Z(n4015) );
  AND U8371 ( .A(n11011), .B(n4015), .Z(n4016) );
  OR U8372 ( .A(n11013), .B(n4016), .Z(n4017) );
  NAND U8373 ( .A(n11015), .B(n4017), .Z(n4018) );
  NANDN U8374 ( .A(n11017), .B(n4018), .Z(n4019) );
  NAND U8375 ( .A(n11019), .B(n4019), .Z(n4020) );
  NANDN U8376 ( .A(n11021), .B(n4020), .Z(n4021) );
  AND U8377 ( .A(n11023), .B(n4021), .Z(n4022) );
  OR U8378 ( .A(n11025), .B(n4022), .Z(n4023) );
  NAND U8379 ( .A(n11027), .B(n4023), .Z(n4024) );
  NANDN U8380 ( .A(n11029), .B(n4024), .Z(n4025) );
  NAND U8381 ( .A(n11031), .B(n4025), .Z(n4026) );
  NANDN U8382 ( .A(n11033), .B(n4026), .Z(n4027) );
  AND U8383 ( .A(n11035), .B(n4027), .Z(n4028) );
  OR U8384 ( .A(n11037), .B(n4028), .Z(n4029) );
  NAND U8385 ( .A(n11039), .B(n4029), .Z(n4030) );
  NANDN U8386 ( .A(n11041), .B(n4030), .Z(n4031) );
  NAND U8387 ( .A(n11043), .B(n4031), .Z(n4032) );
  NANDN U8388 ( .A(n11045), .B(n4032), .Z(n4033) );
  AND U8389 ( .A(n11047), .B(n4033), .Z(n4034) );
  OR U8390 ( .A(n11049), .B(n4034), .Z(n4035) );
  NAND U8391 ( .A(n11051), .B(n4035), .Z(n4036) );
  NANDN U8392 ( .A(n11053), .B(n4036), .Z(n4037) );
  NAND U8393 ( .A(n11055), .B(n4037), .Z(n4038) );
  NANDN U8394 ( .A(n11057), .B(n4038), .Z(n4039) );
  AND U8395 ( .A(n11059), .B(n4039), .Z(n4040) );
  OR U8396 ( .A(n11061), .B(n4040), .Z(n4041) );
  NAND U8397 ( .A(n11063), .B(n4041), .Z(n4042) );
  NANDN U8398 ( .A(n11065), .B(n4042), .Z(n4043) );
  NAND U8399 ( .A(n11067), .B(n4043), .Z(n4044) );
  NANDN U8400 ( .A(n11069), .B(n4044), .Z(n4045) );
  AND U8401 ( .A(n11071), .B(n4045), .Z(n4046) );
  OR U8402 ( .A(n11073), .B(n4046), .Z(n4047) );
  NAND U8403 ( .A(n11075), .B(n4047), .Z(n4048) );
  NANDN U8404 ( .A(n11077), .B(n4048), .Z(n4049) );
  NAND U8405 ( .A(n11079), .B(n4049), .Z(n4050) );
  NANDN U8406 ( .A(n11081), .B(n4050), .Z(n4051) );
  AND U8407 ( .A(n11083), .B(n4051), .Z(n4052) );
  OR U8408 ( .A(n11085), .B(n4052), .Z(n4053) );
  NAND U8409 ( .A(n11087), .B(n4053), .Z(n4054) );
  NANDN U8410 ( .A(n11089), .B(n4054), .Z(n4055) );
  NAND U8411 ( .A(n11091), .B(n4055), .Z(n4056) );
  NANDN U8412 ( .A(n11093), .B(n4056), .Z(n4057) );
  AND U8413 ( .A(n11095), .B(n4057), .Z(n4058) );
  OR U8414 ( .A(n11097), .B(n4058), .Z(n4059) );
  NAND U8415 ( .A(n11099), .B(n4059), .Z(n4060) );
  NANDN U8416 ( .A(n11101), .B(n4060), .Z(n4061) );
  NAND U8417 ( .A(n11103), .B(n4061), .Z(n4062) );
  NANDN U8418 ( .A(n11105), .B(n4062), .Z(n4063) );
  AND U8419 ( .A(n11107), .B(n4063), .Z(n4064) );
  OR U8420 ( .A(n11109), .B(n4064), .Z(n4065) );
  NAND U8421 ( .A(n11111), .B(n4065), .Z(n4066) );
  NANDN U8422 ( .A(n11113), .B(n4066), .Z(n4067) );
  NAND U8423 ( .A(n11115), .B(n4067), .Z(n4068) );
  NANDN U8424 ( .A(n11117), .B(n4068), .Z(n4069) );
  AND U8425 ( .A(n11119), .B(n4069), .Z(n4070) );
  OR U8426 ( .A(n11121), .B(n4070), .Z(n4071) );
  NAND U8427 ( .A(n11123), .B(n4071), .Z(n4072) );
  NANDN U8428 ( .A(n11125), .B(n4072), .Z(n4073) );
  NAND U8429 ( .A(n11127), .B(n4073), .Z(n4074) );
  NANDN U8430 ( .A(n11129), .B(n4074), .Z(n4075) );
  AND U8431 ( .A(n11131), .B(n4075), .Z(n4076) );
  OR U8432 ( .A(n11133), .B(n4076), .Z(n4077) );
  NAND U8433 ( .A(n11135), .B(n4077), .Z(n4078) );
  NANDN U8434 ( .A(n11137), .B(n4078), .Z(n4079) );
  NAND U8435 ( .A(n11139), .B(n4079), .Z(n4080) );
  NANDN U8436 ( .A(n11141), .B(n4080), .Z(n4081) );
  AND U8437 ( .A(n11143), .B(n4081), .Z(n4082) );
  OR U8438 ( .A(n11145), .B(n4082), .Z(n4083) );
  NAND U8439 ( .A(n11147), .B(n4083), .Z(n4084) );
  NANDN U8440 ( .A(n11149), .B(n4084), .Z(n4085) );
  NAND U8441 ( .A(n11151), .B(n4085), .Z(n4086) );
  NANDN U8442 ( .A(n11153), .B(n4086), .Z(n4087) );
  AND U8443 ( .A(n11155), .B(n4087), .Z(n4088) );
  OR U8444 ( .A(n11157), .B(n4088), .Z(n4089) );
  NAND U8445 ( .A(n11159), .B(n4089), .Z(n4090) );
  NANDN U8446 ( .A(n11161), .B(n4090), .Z(n4091) );
  NAND U8447 ( .A(n11163), .B(n4091), .Z(n4092) );
  NANDN U8448 ( .A(n11165), .B(n4092), .Z(n4093) );
  AND U8449 ( .A(n11167), .B(n4093), .Z(n4094) );
  OR U8450 ( .A(n11169), .B(n4094), .Z(n4095) );
  NAND U8451 ( .A(n11171), .B(n4095), .Z(n4096) );
  NANDN U8452 ( .A(n11173), .B(n4096), .Z(n4097) );
  NAND U8453 ( .A(n11175), .B(n4097), .Z(n4098) );
  NANDN U8454 ( .A(n11177), .B(n4098), .Z(n4099) );
  AND U8455 ( .A(n11179), .B(n4099), .Z(n4100) );
  OR U8456 ( .A(n11181), .B(n4100), .Z(n4101) );
  NAND U8457 ( .A(n11183), .B(n4101), .Z(n4102) );
  NANDN U8458 ( .A(n11185), .B(n4102), .Z(n4103) );
  NAND U8459 ( .A(n11187), .B(n4103), .Z(n4104) );
  NANDN U8460 ( .A(n11189), .B(n4104), .Z(n4105) );
  AND U8461 ( .A(n11191), .B(n4105), .Z(n4106) );
  OR U8462 ( .A(n11193), .B(n4106), .Z(n4107) );
  NAND U8463 ( .A(n11195), .B(n4107), .Z(n4108) );
  NANDN U8464 ( .A(n11197), .B(n4108), .Z(n4109) );
  NAND U8465 ( .A(n11199), .B(n4109), .Z(n4110) );
  NANDN U8466 ( .A(n11201), .B(n4110), .Z(n4111) );
  AND U8467 ( .A(n11203), .B(n4111), .Z(n4112) );
  OR U8468 ( .A(n11205), .B(n4112), .Z(n4113) );
  NAND U8469 ( .A(n11207), .B(n4113), .Z(n4114) );
  NANDN U8470 ( .A(n11209), .B(n4114), .Z(n4115) );
  NAND U8471 ( .A(n11211), .B(n4115), .Z(n4116) );
  NANDN U8472 ( .A(n11213), .B(n4116), .Z(n4117) );
  AND U8473 ( .A(n11215), .B(n4117), .Z(n4118) );
  OR U8474 ( .A(n11217), .B(n4118), .Z(n4119) );
  NAND U8475 ( .A(n11219), .B(n4119), .Z(n4120) );
  NANDN U8476 ( .A(n11221), .B(n4120), .Z(n4121) );
  NAND U8477 ( .A(n11223), .B(n4121), .Z(n4122) );
  NANDN U8478 ( .A(n11225), .B(n4122), .Z(n4123) );
  AND U8479 ( .A(n11227), .B(n4123), .Z(n4124) );
  OR U8480 ( .A(n11229), .B(n4124), .Z(n4125) );
  NAND U8481 ( .A(n11231), .B(n4125), .Z(n4126) );
  NANDN U8482 ( .A(n11233), .B(n4126), .Z(n4127) );
  NAND U8483 ( .A(n11235), .B(n4127), .Z(n4128) );
  NANDN U8484 ( .A(n11237), .B(n4128), .Z(n4129) );
  AND U8485 ( .A(n11239), .B(n4129), .Z(n4130) );
  OR U8486 ( .A(n11241), .B(n4130), .Z(n4131) );
  NAND U8487 ( .A(n11243), .B(n4131), .Z(n4132) );
  NANDN U8488 ( .A(n11245), .B(n4132), .Z(n4133) );
  NAND U8489 ( .A(n11247), .B(n4133), .Z(n4134) );
  NANDN U8490 ( .A(n11249), .B(n4134), .Z(n4135) );
  AND U8491 ( .A(n11251), .B(n4135), .Z(n4136) );
  OR U8492 ( .A(n11253), .B(n4136), .Z(n4137) );
  NAND U8493 ( .A(n11255), .B(n4137), .Z(n4138) );
  NANDN U8494 ( .A(n11257), .B(n4138), .Z(n4139) );
  NAND U8495 ( .A(n11259), .B(n4139), .Z(n4140) );
  NANDN U8496 ( .A(n11261), .B(n4140), .Z(n4141) );
  AND U8497 ( .A(n11263), .B(n4141), .Z(n4142) );
  OR U8498 ( .A(n11265), .B(n4142), .Z(n4143) );
  NAND U8499 ( .A(n11267), .B(n4143), .Z(n4144) );
  NANDN U8500 ( .A(n11269), .B(n4144), .Z(n4145) );
  NAND U8501 ( .A(n11271), .B(n4145), .Z(n4146) );
  NANDN U8502 ( .A(n11273), .B(n4146), .Z(n4147) );
  AND U8503 ( .A(n11275), .B(n4147), .Z(n4148) );
  OR U8504 ( .A(n11277), .B(n4148), .Z(n4149) );
  NAND U8505 ( .A(n11279), .B(n4149), .Z(n4150) );
  NANDN U8506 ( .A(n11281), .B(n4150), .Z(n4151) );
  NAND U8507 ( .A(n11283), .B(n4151), .Z(n4152) );
  NANDN U8508 ( .A(n11285), .B(n4152), .Z(n4153) );
  AND U8509 ( .A(n11287), .B(n4153), .Z(n4154) );
  OR U8510 ( .A(n11289), .B(n4154), .Z(n4155) );
  NAND U8511 ( .A(n11291), .B(n4155), .Z(n4156) );
  NANDN U8512 ( .A(n11293), .B(n4156), .Z(n4157) );
  NAND U8513 ( .A(n11295), .B(n4157), .Z(n4158) );
  NANDN U8514 ( .A(n11297), .B(n4158), .Z(n4159) );
  AND U8515 ( .A(n11299), .B(n4159), .Z(n4160) );
  OR U8516 ( .A(n11301), .B(n4160), .Z(n4161) );
  NAND U8517 ( .A(n11303), .B(n4161), .Z(n4162) );
  NANDN U8518 ( .A(n11305), .B(n4162), .Z(n4163) );
  NAND U8519 ( .A(n11307), .B(n4163), .Z(n4164) );
  NANDN U8520 ( .A(n11309), .B(n4164), .Z(n4165) );
  AND U8521 ( .A(n11311), .B(n4165), .Z(n4166) );
  OR U8522 ( .A(n11313), .B(n4166), .Z(n4167) );
  NAND U8523 ( .A(n11315), .B(n4167), .Z(n4168) );
  NANDN U8524 ( .A(n11317), .B(n4168), .Z(n4169) );
  NAND U8525 ( .A(n11319), .B(n4169), .Z(n4170) );
  NANDN U8526 ( .A(n11321), .B(n4170), .Z(n4171) );
  AND U8527 ( .A(n11323), .B(n4171), .Z(n4172) );
  OR U8528 ( .A(n11325), .B(n4172), .Z(n4173) );
  NAND U8529 ( .A(n11327), .B(n4173), .Z(n4174) );
  NANDN U8530 ( .A(n11329), .B(n4174), .Z(n4175) );
  NAND U8531 ( .A(n11331), .B(n4175), .Z(n4176) );
  NANDN U8532 ( .A(n11333), .B(n4176), .Z(n4177) );
  AND U8533 ( .A(n11335), .B(n4177), .Z(n4178) );
  OR U8534 ( .A(n11337), .B(n4178), .Z(n4179) );
  NAND U8535 ( .A(n11339), .B(n4179), .Z(n4180) );
  NANDN U8536 ( .A(n11341), .B(n4180), .Z(n4181) );
  NAND U8537 ( .A(n11343), .B(n4181), .Z(n4182) );
  NANDN U8538 ( .A(n11345), .B(n4182), .Z(n4183) );
  AND U8539 ( .A(n11347), .B(n4183), .Z(n4184) );
  OR U8540 ( .A(n11349), .B(n4184), .Z(n4185) );
  NAND U8541 ( .A(n11351), .B(n4185), .Z(n4186) );
  NANDN U8542 ( .A(n11353), .B(n4186), .Z(n4187) );
  NAND U8543 ( .A(n11355), .B(n4187), .Z(n4188) );
  NANDN U8544 ( .A(n11357), .B(n4188), .Z(n4189) );
  AND U8545 ( .A(n11359), .B(n4189), .Z(n4190) );
  OR U8546 ( .A(n11361), .B(n4190), .Z(n4191) );
  NAND U8547 ( .A(n11363), .B(n4191), .Z(n4192) );
  NANDN U8548 ( .A(n11365), .B(n4192), .Z(n4193) );
  NAND U8549 ( .A(n11367), .B(n4193), .Z(n4194) );
  NANDN U8550 ( .A(n11369), .B(n4194), .Z(n4195) );
  AND U8551 ( .A(n11371), .B(n4195), .Z(n4196) );
  OR U8552 ( .A(n11373), .B(n4196), .Z(n4197) );
  NAND U8553 ( .A(n11375), .B(n4197), .Z(n4198) );
  NANDN U8554 ( .A(n11377), .B(n4198), .Z(n4199) );
  NAND U8555 ( .A(n11379), .B(n4199), .Z(n4200) );
  NANDN U8556 ( .A(n11381), .B(n4200), .Z(n4201) );
  AND U8557 ( .A(n11383), .B(n4201), .Z(n4202) );
  OR U8558 ( .A(n11385), .B(n4202), .Z(n4203) );
  NAND U8559 ( .A(n11387), .B(n4203), .Z(n4204) );
  NANDN U8560 ( .A(n11389), .B(n4204), .Z(n4205) );
  NAND U8561 ( .A(n11391), .B(n4205), .Z(n4206) );
  NANDN U8562 ( .A(n11393), .B(n4206), .Z(n4207) );
  AND U8563 ( .A(n11395), .B(n4207), .Z(n4208) );
  OR U8564 ( .A(n11397), .B(n4208), .Z(n4209) );
  NAND U8565 ( .A(n11399), .B(n4209), .Z(n4210) );
  NANDN U8566 ( .A(n11401), .B(n4210), .Z(n4211) );
  NAND U8567 ( .A(n11403), .B(n4211), .Z(n4212) );
  NANDN U8568 ( .A(n11405), .B(n4212), .Z(n4213) );
  AND U8569 ( .A(n11407), .B(n4213), .Z(n4214) );
  OR U8570 ( .A(n11409), .B(n4214), .Z(n4215) );
  NAND U8571 ( .A(n11411), .B(n4215), .Z(n4216) );
  NANDN U8572 ( .A(n11413), .B(n4216), .Z(n4217) );
  NAND U8573 ( .A(n11415), .B(n4217), .Z(n4218) );
  NANDN U8574 ( .A(n11417), .B(n4218), .Z(n4219) );
  AND U8575 ( .A(n11419), .B(n4219), .Z(n4220) );
  OR U8576 ( .A(n11421), .B(n4220), .Z(n4221) );
  NAND U8577 ( .A(n11423), .B(n4221), .Z(n4222) );
  NANDN U8578 ( .A(n11425), .B(n4222), .Z(n4223) );
  NAND U8579 ( .A(n11427), .B(n4223), .Z(n4224) );
  NANDN U8580 ( .A(n11429), .B(n4224), .Z(n4225) );
  AND U8581 ( .A(n11431), .B(n4225), .Z(n4226) );
  OR U8582 ( .A(n11433), .B(n4226), .Z(n4227) );
  NAND U8583 ( .A(n11435), .B(n4227), .Z(n4228) );
  NANDN U8584 ( .A(n11437), .B(n4228), .Z(n4229) );
  NAND U8585 ( .A(n11439), .B(n4229), .Z(n4230) );
  NANDN U8586 ( .A(n11441), .B(n4230), .Z(n4231) );
  AND U8587 ( .A(n11443), .B(n4231), .Z(n4232) );
  OR U8588 ( .A(n11445), .B(n4232), .Z(n4233) );
  NAND U8589 ( .A(n11447), .B(n4233), .Z(n4234) );
  NANDN U8590 ( .A(n11449), .B(n4234), .Z(n4235) );
  NAND U8591 ( .A(n11451), .B(n4235), .Z(n4236) );
  NANDN U8592 ( .A(n11453), .B(n4236), .Z(n4237) );
  AND U8593 ( .A(n11455), .B(n4237), .Z(n4238) );
  OR U8594 ( .A(n11457), .B(n4238), .Z(n4239) );
  NAND U8595 ( .A(n11459), .B(n4239), .Z(n4240) );
  NANDN U8596 ( .A(n11461), .B(n4240), .Z(n4241) );
  NAND U8597 ( .A(n11463), .B(n4241), .Z(n4242) );
  NANDN U8598 ( .A(n11465), .B(n4242), .Z(n4243) );
  AND U8599 ( .A(n11467), .B(n4243), .Z(n4244) );
  OR U8600 ( .A(n11469), .B(n4244), .Z(n4245) );
  NAND U8601 ( .A(n11471), .B(n4245), .Z(n4246) );
  NANDN U8602 ( .A(n11473), .B(n4246), .Z(n4247) );
  NAND U8603 ( .A(n11475), .B(n4247), .Z(n4248) );
  NAND U8604 ( .A(n11476), .B(n4248), .Z(n4251) );
  NANDN U8605 ( .A(x[649]), .B(y[649]), .Z(n4250) );
  NANDN U8606 ( .A(x[648]), .B(y[648]), .Z(n4249) );
  NAND U8607 ( .A(n4250), .B(n4249), .Z(n11479) );
  ANDN U8608 ( .B(n4251), .A(n11479), .Z(n4254) );
  NANDN U8609 ( .A(y[649]), .B(x[649]), .Z(n4253) );
  NANDN U8610 ( .A(y[650]), .B(x[650]), .Z(n4252) );
  AND U8611 ( .A(n4253), .B(n4252), .Z(n11481) );
  NANDN U8612 ( .A(n4254), .B(n11481), .Z(n4255) );
  NANDN U8613 ( .A(n11483), .B(n4255), .Z(n4256) );
  NAND U8614 ( .A(n11485), .B(n4256), .Z(n4257) );
  NANDN U8615 ( .A(n11486), .B(n4257), .Z(n4258) );
  NAND U8616 ( .A(n11488), .B(n4258), .Z(n4261) );
  NANDN U8617 ( .A(x[655]), .B(y[655]), .Z(n4260) );
  NANDN U8618 ( .A(x[654]), .B(y[654]), .Z(n4259) );
  NAND U8619 ( .A(n4260), .B(n4259), .Z(n11491) );
  ANDN U8620 ( .B(n4261), .A(n11491), .Z(n4264) );
  NANDN U8621 ( .A(y[655]), .B(x[655]), .Z(n4263) );
  NANDN U8622 ( .A(y[656]), .B(x[656]), .Z(n4262) );
  AND U8623 ( .A(n4263), .B(n4262), .Z(n11493) );
  NANDN U8624 ( .A(n4264), .B(n11493), .Z(n4265) );
  NAND U8625 ( .A(n11495), .B(n4265), .Z(n4266) );
  NANDN U8626 ( .A(n11497), .B(n4266), .Z(n4267) );
  NAND U8627 ( .A(n11499), .B(n4267), .Z(n4268) );
  NANDN U8628 ( .A(n11501), .B(n4268), .Z(n4269) );
  AND U8629 ( .A(n11503), .B(n4269), .Z(n4270) );
  OR U8630 ( .A(n11505), .B(n4270), .Z(n4271) );
  NAND U8631 ( .A(n11507), .B(n4271), .Z(n4272) );
  NANDN U8632 ( .A(n11509), .B(n4272), .Z(n4273) );
  NAND U8633 ( .A(n11511), .B(n4273), .Z(n4274) );
  NANDN U8634 ( .A(n11513), .B(n4274), .Z(n4275) );
  AND U8635 ( .A(n11515), .B(n4275), .Z(n4276) );
  OR U8636 ( .A(n11517), .B(n4276), .Z(n4277) );
  NAND U8637 ( .A(n11519), .B(n4277), .Z(n4278) );
  NANDN U8638 ( .A(n11521), .B(n4278), .Z(n4279) );
  NAND U8639 ( .A(n11523), .B(n4279), .Z(n4280) );
  NANDN U8640 ( .A(n11525), .B(n4280), .Z(n4281) );
  AND U8641 ( .A(n11527), .B(n4281), .Z(n4282) );
  OR U8642 ( .A(n11529), .B(n4282), .Z(n4283) );
  NAND U8643 ( .A(n11531), .B(n4283), .Z(n4284) );
  NANDN U8644 ( .A(n11533), .B(n4284), .Z(n4285) );
  NAND U8645 ( .A(n11535), .B(n4285), .Z(n4286) );
  NANDN U8646 ( .A(n11537), .B(n4286), .Z(n4287) );
  AND U8647 ( .A(n11539), .B(n4287), .Z(n4288) );
  OR U8648 ( .A(n11541), .B(n4288), .Z(n4289) );
  NAND U8649 ( .A(n11543), .B(n4289), .Z(n4290) );
  NANDN U8650 ( .A(n11545), .B(n4290), .Z(n4291) );
  NAND U8651 ( .A(n11547), .B(n4291), .Z(n4292) );
  NANDN U8652 ( .A(n11549), .B(n4292), .Z(n4293) );
  AND U8653 ( .A(n11551), .B(n4293), .Z(n4294) );
  OR U8654 ( .A(n11553), .B(n4294), .Z(n4295) );
  NAND U8655 ( .A(n11555), .B(n4295), .Z(n4296) );
  NANDN U8656 ( .A(n11557), .B(n4296), .Z(n4297) );
  NAND U8657 ( .A(n11559), .B(n4297), .Z(n4298) );
  NANDN U8658 ( .A(n11561), .B(n4298), .Z(n4299) );
  AND U8659 ( .A(n11563), .B(n4299), .Z(n4300) );
  OR U8660 ( .A(n11565), .B(n4300), .Z(n4301) );
  NAND U8661 ( .A(n11567), .B(n4301), .Z(n4302) );
  NANDN U8662 ( .A(n11569), .B(n4302), .Z(n4303) );
  NAND U8663 ( .A(n11571), .B(n4303), .Z(n4304) );
  NANDN U8664 ( .A(n11573), .B(n4304), .Z(n4305) );
  AND U8665 ( .A(n11575), .B(n4305), .Z(n4306) );
  OR U8666 ( .A(n11577), .B(n4306), .Z(n4307) );
  NAND U8667 ( .A(n11579), .B(n4307), .Z(n4308) );
  NANDN U8668 ( .A(n11581), .B(n4308), .Z(n4309) );
  NAND U8669 ( .A(n11583), .B(n4309), .Z(n4310) );
  NANDN U8670 ( .A(n11585), .B(n4310), .Z(n4311) );
  AND U8671 ( .A(n11587), .B(n4311), .Z(n4312) );
  OR U8672 ( .A(n11589), .B(n4312), .Z(n4313) );
  NAND U8673 ( .A(n11591), .B(n4313), .Z(n4314) );
  NANDN U8674 ( .A(n11593), .B(n4314), .Z(n4315) );
  NAND U8675 ( .A(n11595), .B(n4315), .Z(n4316) );
  NANDN U8676 ( .A(n11597), .B(n4316), .Z(n4317) );
  AND U8677 ( .A(n11599), .B(n4317), .Z(n4318) );
  OR U8678 ( .A(n11601), .B(n4318), .Z(n4319) );
  NANDN U8679 ( .A(y[715]), .B(x[715]), .Z(n4321) );
  NANDN U8680 ( .A(y[716]), .B(x[716]), .Z(n4320) );
  AND U8681 ( .A(n4321), .B(n4320), .Z(n11613) );
  NANDN U8682 ( .A(y[717]), .B(x[717]), .Z(n8414) );
  NANDN U8683 ( .A(y[718]), .B(x[718]), .Z(n8417) );
  AND U8684 ( .A(n8414), .B(n8417), .Z(n11617) );
  ANDN U8685 ( .B(y[718]), .A(x[718]), .Z(n8416) );
  ANDN U8686 ( .B(y[719]), .A(x[719]), .Z(n8423) );
  NOR U8687 ( .A(n8416), .B(n8423), .Z(n11619) );
  NANDN U8688 ( .A(y[723]), .B(x[723]), .Z(n8430) );
  ANDN U8689 ( .B(x[724]), .A(y[724]), .Z(n8440) );
  ANDN U8690 ( .B(n8430), .A(n8440), .Z(n11629) );
  NANDN U8691 ( .A(x[725]), .B(y[725]), .Z(n8442) );
  ANDN U8692 ( .B(y[724]), .A(x[724]), .Z(n8434) );
  ANDN U8693 ( .B(n8442), .A(n8434), .Z(n11631) );
  XNOR U8694 ( .A(x[730]), .B(y[730]), .Z(n4323) );
  ANDN U8695 ( .B(x[729]), .A(y[729]), .Z(n8449) );
  ANDN U8696 ( .B(n4323), .A(n8449), .Z(n11641) );
  NANDN U8697 ( .A(x[730]), .B(y[730]), .Z(n8451) );
  ANDN U8698 ( .B(y[731]), .A(x[731]), .Z(n8459) );
  ANDN U8699 ( .B(n8451), .A(n8459), .Z(n11643) );
  NANDN U8700 ( .A(y[736]), .B(x[736]), .Z(n5689) );
  ANDN U8701 ( .B(x[735]), .A(y[735]), .Z(n8467) );
  ANDN U8702 ( .B(n5689), .A(n8467), .Z(n11653) );
  IV U8703 ( .A(n11653), .Z(n4324) );
  NANDN U8704 ( .A(x[736]), .B(y[736]), .Z(n5690) );
  NANDN U8705 ( .A(x[737]), .B(y[737]), .Z(n8474) );
  NAND U8706 ( .A(n5690), .B(n8474), .Z(n11654) );
  IV U8707 ( .A(n11654), .Z(n4326) );
  NANDN U8708 ( .A(y[741]), .B(x[741]), .Z(n5684) );
  ANDN U8709 ( .B(x[742]), .A(y[742]), .Z(n8492) );
  ANDN U8710 ( .B(n5684), .A(n8492), .Z(n11665) );
  NANDN U8711 ( .A(x[742]), .B(y[742]), .Z(n8487) );
  NANDN U8712 ( .A(x[743]), .B(y[743]), .Z(n5683) );
  NAND U8713 ( .A(n8487), .B(n5683), .Z(n11666) );
  NANDN U8714 ( .A(y[748]), .B(x[748]), .Z(n5677) );
  ANDN U8715 ( .B(x[747]), .A(y[747]), .Z(n8503) );
  ANDN U8716 ( .B(n5677), .A(n8503), .Z(n11677) );
  IV U8717 ( .A(n11677), .Z(n4329) );
  NANDN U8718 ( .A(x[748]), .B(y[748]), .Z(n5678) );
  NANDN U8719 ( .A(x[749]), .B(y[749]), .Z(n8510) );
  NAND U8720 ( .A(n5678), .B(n8510), .Z(n11678) );
  NANDN U8721 ( .A(y[753]), .B(x[753]), .Z(n5672) );
  ANDN U8722 ( .B(x[754]), .A(y[754]), .Z(n8528) );
  ANDN U8723 ( .B(n5672), .A(n8528), .Z(n11689) );
  NANDN U8724 ( .A(x[754]), .B(y[754]), .Z(n8523) );
  NANDN U8725 ( .A(x[755]), .B(y[755]), .Z(n5671) );
  NAND U8726 ( .A(n8523), .B(n5671), .Z(n11690) );
  NANDN U8727 ( .A(y[760]), .B(x[760]), .Z(n5667) );
  ANDN U8728 ( .B(x[759]), .A(y[759]), .Z(n8539) );
  ANDN U8729 ( .B(n5667), .A(n8539), .Z(n11701) );
  NANDN U8730 ( .A(x[760]), .B(y[760]), .Z(n8543) );
  ANDN U8731 ( .B(y[761]), .A(x[761]), .Z(n8550) );
  ANDN U8732 ( .B(n8543), .A(n8550), .Z(n11703) );
  NANDN U8733 ( .A(y[765]), .B(x[765]), .Z(n8556) );
  ANDN U8734 ( .B(x[766]), .A(y[766]), .Z(n5660) );
  ANDN U8735 ( .B(n8556), .A(n5660), .Z(n11713) );
  NANDN U8736 ( .A(x[767]), .B(y[767]), .Z(n8561) );
  ANDN U8737 ( .B(y[766]), .A(x[766]), .Z(n8558) );
  ANDN U8738 ( .B(n8561), .A(n8558), .Z(n11715) );
  NANDN U8739 ( .A(y[771]), .B(x[771]), .Z(n8571) );
  NANDN U8740 ( .A(y[772]), .B(x[772]), .Z(n8579) );
  AND U8741 ( .A(n8571), .B(n8579), .Z(n11725) );
  IV U8742 ( .A(n11725), .Z(n4333) );
  NANDN U8743 ( .A(x[772]), .B(y[772]), .Z(n8576) );
  NANDN U8744 ( .A(x[773]), .B(y[773]), .Z(n8584) );
  NAND U8745 ( .A(n8576), .B(n8584), .Z(n11726) );
  NANDN U8746 ( .A(y[777]), .B(x[777]), .Z(n4335) );
  NANDN U8747 ( .A(y[778]), .B(x[778]), .Z(n4334) );
  AND U8748 ( .A(n4335), .B(n4334), .Z(n11737) );
  IV U8749 ( .A(n11737), .Z(n8594) );
  NANDN U8750 ( .A(x[779]), .B(y[779]), .Z(n4337) );
  NANDN U8751 ( .A(x[778]), .B(y[778]), .Z(n4336) );
  NAND U8752 ( .A(n4337), .B(n4336), .Z(n11738) );
  IV U8753 ( .A(n11738), .Z(n8596) );
  NANDN U8754 ( .A(y[783]), .B(x[783]), .Z(n4339) );
  NANDN U8755 ( .A(y[784]), .B(x[784]), .Z(n4338) );
  AND U8756 ( .A(n4339), .B(n4338), .Z(n11749) );
  IV U8757 ( .A(n11749), .Z(n8606) );
  NANDN U8758 ( .A(x[785]), .B(y[785]), .Z(n4341) );
  NANDN U8759 ( .A(x[784]), .B(y[784]), .Z(n4340) );
  NAND U8760 ( .A(n4341), .B(n4340), .Z(n11750) );
  IV U8761 ( .A(n11750), .Z(n8608) );
  NANDN U8762 ( .A(n4343), .B(n4342), .Z(n4344) );
  NAND U8763 ( .A(n11759), .B(n4344), .Z(n4345) );
  NANDN U8764 ( .A(n11761), .B(n4345), .Z(n4346) );
  NAND U8765 ( .A(n11763), .B(n4346), .Z(n4347) );
  NANDN U8766 ( .A(n11765), .B(n4347), .Z(n4348) );
  AND U8767 ( .A(n11767), .B(n4348), .Z(n4349) );
  OR U8768 ( .A(n11769), .B(n4349), .Z(n4350) );
  NAND U8769 ( .A(n11771), .B(n4350), .Z(n4351) );
  NANDN U8770 ( .A(n11773), .B(n4351), .Z(n4352) );
  NAND U8771 ( .A(n11775), .B(n4352), .Z(n4353) );
  NANDN U8772 ( .A(n11777), .B(n4353), .Z(n4354) );
  AND U8773 ( .A(n11779), .B(n4354), .Z(n4355) );
  OR U8774 ( .A(n11781), .B(n4355), .Z(n4356) );
  NAND U8775 ( .A(n11783), .B(n4356), .Z(n4357) );
  NANDN U8776 ( .A(n11785), .B(n4357), .Z(n4358) );
  NAND U8777 ( .A(n11787), .B(n4358), .Z(n4359) );
  NANDN U8778 ( .A(n11789), .B(n4359), .Z(n4360) );
  AND U8779 ( .A(n11791), .B(n4360), .Z(n4361) );
  OR U8780 ( .A(n11793), .B(n4361), .Z(n4362) );
  NAND U8781 ( .A(n11795), .B(n4362), .Z(n4363) );
  NANDN U8782 ( .A(n11797), .B(n4363), .Z(n4364) );
  NAND U8783 ( .A(n11799), .B(n4364), .Z(n4365) );
  NANDN U8784 ( .A(n11801), .B(n4365), .Z(n4366) );
  AND U8785 ( .A(n11803), .B(n4366), .Z(n4367) );
  OR U8786 ( .A(n11805), .B(n4367), .Z(n4368) );
  NAND U8787 ( .A(n11807), .B(n4368), .Z(n4369) );
  NANDN U8788 ( .A(n11809), .B(n4369), .Z(n4370) );
  NAND U8789 ( .A(n11811), .B(n4370), .Z(n4371) );
  NANDN U8790 ( .A(n11813), .B(n4371), .Z(n4372) );
  AND U8791 ( .A(n11815), .B(n4372), .Z(n4373) );
  OR U8792 ( .A(n11817), .B(n4373), .Z(n4374) );
  NAND U8793 ( .A(n11819), .B(n4374), .Z(n4375) );
  NANDN U8794 ( .A(n11821), .B(n4375), .Z(n4376) );
  NAND U8795 ( .A(n11823), .B(n4376), .Z(n4377) );
  NANDN U8796 ( .A(n11825), .B(n4377), .Z(n4378) );
  AND U8797 ( .A(n11827), .B(n4378), .Z(n4380) );
  NANDN U8798 ( .A(y[824]), .B(x[824]), .Z(n5637) );
  NANDN U8799 ( .A(y[823]), .B(x[823]), .Z(n11829) );
  AND U8800 ( .A(n5637), .B(n11829), .Z(n4379) );
  NANDN U8801 ( .A(n4380), .B(n4379), .Z(n4381) );
  AND U8802 ( .A(n4382), .B(n4381), .Z(n4384) );
  NANDN U8803 ( .A(y[825]), .B(x[825]), .Z(n5636) );
  NANDN U8804 ( .A(y[826]), .B(x[826]), .Z(n11836) );
  AND U8805 ( .A(n5636), .B(n11836), .Z(n4383) );
  NANDN U8806 ( .A(y[828]), .B(x[828]), .Z(n5635) );
  ANDN U8807 ( .B(x[827]), .A(y[827]), .Z(n11841) );
  NANDN U8808 ( .A(x[829]), .B(y[829]), .Z(n5632) );
  ANDN U8809 ( .B(x[830]), .A(y[830]), .Z(n8734) );
  NANDN U8810 ( .A(x[831]), .B(y[831]), .Z(n11851) );
  NANDN U8811 ( .A(y[831]), .B(x[831]), .Z(n8733) );
  ANDN U8812 ( .B(x[840]), .A(y[840]), .Z(n5626) );
  NANDN U8813 ( .A(y[846]), .B(x[846]), .Z(n11878) );
  NANDN U8814 ( .A(y[848]), .B(x[848]), .Z(n5621) );
  NANDN U8815 ( .A(x[848]), .B(y[848]), .Z(n11884) );
  ANDN U8816 ( .B(x[849]), .A(y[849]), .Z(n5622) );
  NANDN U8817 ( .A(y[858]), .B(x[858]), .Z(n5608) );
  NANDN U8818 ( .A(y[857]), .B(x[857]), .Z(n11907) );
  NANDN U8819 ( .A(x[859]), .B(y[859]), .Z(n5606) );
  ANDN U8820 ( .B(x[860]), .A(y[860]), .Z(n5605) );
  NANDN U8821 ( .A(x[860]), .B(y[860]), .Z(n5607) );
  ANDN U8822 ( .B(x[862]), .A(y[862]), .Z(n5601) );
  NANDN U8823 ( .A(y[863]), .B(x[863]), .Z(n5600) );
  ANDN U8824 ( .B(x[864]), .A(y[864]), .Z(n11923) );
  ANDN U8825 ( .B(n5600), .A(n11923), .Z(n4387) );
  NANDN U8826 ( .A(x[864]), .B(y[864]), .Z(n5599) );
  ANDN U8827 ( .B(x[872]), .A(y[872]), .Z(n5589) );
  NANDN U8828 ( .A(x[875]), .B(y[875]), .Z(n4390) );
  NANDN U8829 ( .A(x[874]), .B(y[874]), .Z(n4389) );
  AND U8830 ( .A(n4390), .B(n4389), .Z(n5585) );
  ANDN U8831 ( .B(x[876]), .A(y[876]), .Z(n5583) );
  ANDN U8832 ( .B(x[875]), .A(y[875]), .Z(n5590) );
  NANDN U8833 ( .A(x[877]), .B(y[877]), .Z(n5581) );
  ANDN U8834 ( .B(x[878]), .A(y[878]), .Z(n5579) );
  IV U8835 ( .A(n5579), .Z(n4391) );
  NANDN U8836 ( .A(x[878]), .B(y[878]), .Z(n5582) );
  ANDN U8837 ( .B(x[880]), .A(y[880]), .Z(n5575) );
  NANDN U8838 ( .A(y[881]), .B(x[881]), .Z(n5576) );
  ANDN U8839 ( .B(x[882]), .A(y[882]), .Z(n11959) );
  NANDN U8840 ( .A(x[883]), .B(y[883]), .Z(n11961) );
  NANDN U8841 ( .A(x[882]), .B(y[882]), .Z(n5574) );
  ANDN U8842 ( .B(y[884]), .A(x[884]), .Z(n8803) );
  ANDN U8843 ( .B(y[885]), .A(x[885]), .Z(n8812) );
  NOR U8844 ( .A(n8803), .B(n8812), .Z(n11965) );
  NANDN U8845 ( .A(y[885]), .B(x[885]), .Z(n8807) );
  XOR U8846 ( .A(x[886]), .B(y[886]), .Z(n8811) );
  ANDN U8847 ( .B(n8807), .A(n8811), .Z(n11967) );
  ANDN U8848 ( .B(x[888]), .A(y[888]), .Z(n5570) );
  NANDN U8849 ( .A(x[889]), .B(y[889]), .Z(n11977) );
  NANDN U8850 ( .A(y[889]), .B(x[889]), .Z(n5571) );
  NANDN U8851 ( .A(y[892]), .B(x[892]), .Z(n5569) );
  NANDN U8852 ( .A(x[893]), .B(y[893]), .Z(n11989) );
  ANDN U8853 ( .B(x[893]), .A(y[893]), .Z(n5568) );
  NANDN U8854 ( .A(x[895]), .B(y[895]), .Z(n8836) );
  ANDN U8855 ( .B(y[894]), .A(x[894]), .Z(n8832) );
  ANDN U8856 ( .B(n8836), .A(n8832), .Z(n11992) );
  NANDN U8857 ( .A(y[896]), .B(x[896]), .Z(n5566) );
  ANDN U8858 ( .B(x[895]), .A(y[895]), .Z(n11995) );
  ANDN U8859 ( .B(y[897]), .A(x[897]), .Z(n5565) );
  NANDN U8860 ( .A(y[899]), .B(x[899]), .Z(n8840) );
  NANDN U8861 ( .A(y[900]), .B(x[900]), .Z(n8848) );
  NAND U8862 ( .A(n8840), .B(n8848), .Z(n12007) );
  ANDN U8863 ( .B(x[907]), .A(y[907]), .Z(n12023) );
  NANDN U8864 ( .A(y[908]), .B(x[908]), .Z(n5560) );
  ANDN U8865 ( .B(y[909]), .A(x[909]), .Z(n8870) );
  NANDN U8866 ( .A(y[909]), .B(x[909]), .Z(n5561) );
  ANDN U8867 ( .B(y[911]), .A(x[911]), .Z(n5558) );
  NANDN U8868 ( .A(y[914]), .B(x[914]), .Z(n12038) );
  NANDN U8869 ( .A(y[913]), .B(x[913]), .Z(n5556) );
  NANDN U8870 ( .A(x[916]), .B(y[916]), .Z(n4399) );
  ANDN U8871 ( .B(y[917]), .A(x[917]), .Z(n5552) );
  ANDN U8872 ( .B(n4399), .A(n5552), .Z(n4402) );
  NANDN U8873 ( .A(x[915]), .B(y[915]), .Z(n4400) );
  AND U8874 ( .A(n4402), .B(n4400), .Z(n12041) );
  NANDN U8875 ( .A(y[917]), .B(x[917]), .Z(n5554) );
  NANDN U8876 ( .A(y[916]), .B(x[916]), .Z(n5551) );
  NANDN U8877 ( .A(y[915]), .B(x[915]), .Z(n5555) );
  NAND U8878 ( .A(n5551), .B(n5555), .Z(n4401) );
  NAND U8879 ( .A(n4402), .B(n4401), .Z(n4403) );
  AND U8880 ( .A(n5554), .B(n4403), .Z(n4405) );
  XNOR U8881 ( .A(y[918]), .B(x[918]), .Z(n4404) );
  NAND U8882 ( .A(n4405), .B(n4404), .Z(n12042) );
  ANDN U8883 ( .B(y[918]), .A(x[918]), .Z(n8875) );
  ANDN U8884 ( .B(y[919]), .A(x[919]), .Z(n8878) );
  NOR U8885 ( .A(n8875), .B(n8878), .Z(n12044) );
  NANDN U8886 ( .A(y[919]), .B(x[919]), .Z(n8876) );
  NANDN U8887 ( .A(y[920]), .B(x[920]), .Z(n5550) );
  NAND U8888 ( .A(n8876), .B(n5550), .Z(n12047) );
  NANDN U8889 ( .A(y[922]), .B(x[922]), .Z(n5549) );
  NANDN U8890 ( .A(y[923]), .B(x[923]), .Z(n5548) );
  ANDN U8891 ( .B(x[924]), .A(y[924]), .Z(n12059) );
  IV U8892 ( .A(n12059), .Z(n8882) );
  AND U8893 ( .A(n5548), .B(n8882), .Z(n4408) );
  NANDN U8894 ( .A(x[924]), .B(y[924]), .Z(n8881) );
  NANDN U8895 ( .A(x[925]), .B(y[925]), .Z(n5547) );
  AND U8896 ( .A(n8881), .B(n5547), .Z(n12061) );
  NANDN U8897 ( .A(y[926]), .B(x[926]), .Z(n8885) );
  ANDN U8898 ( .B(x[925]), .A(y[925]), .Z(n12063) );
  IV U8899 ( .A(n12063), .Z(n8883) );
  NANDN U8900 ( .A(x[926]), .B(y[926]), .Z(n12065) );
  IV U8901 ( .A(n12065), .Z(n5546) );
  NANDN U8902 ( .A(x[927]), .B(y[927]), .Z(n5545) );
  ANDN U8903 ( .B(x[928]), .A(y[928]), .Z(n5542) );
  ANDN U8904 ( .B(x[927]), .A(y[927]), .Z(n8884) );
  ANDN U8905 ( .B(y[928]), .A(x[928]), .Z(n5544) );
  ANDN U8906 ( .B(y[929]), .A(x[929]), .Z(n12073) );
  NANDN U8907 ( .A(y[929]), .B(x[929]), .Z(n5543) );
  NANDN U8908 ( .A(y[935]), .B(x[935]), .Z(n12087) );
  ANDN U8909 ( .B(y[937]), .A(x[937]), .Z(n5538) );
  NANDN U8910 ( .A(x[939]), .B(y[939]), .Z(n12097) );
  NANDN U8911 ( .A(y[939]), .B(x[939]), .Z(n5536) );
  ANDN U8912 ( .B(y[940]), .A(x[940]), .Z(n8897) );
  ANDN U8913 ( .B(y[941]), .A(x[941]), .Z(n8899) );
  NOR U8914 ( .A(n8897), .B(n8899), .Z(n12101) );
  NANDN U8915 ( .A(y[942]), .B(x[942]), .Z(n4410) );
  AND U8916 ( .A(n4411), .B(n4410), .Z(n8900) );
  NANDN U8917 ( .A(y[941]), .B(x[941]), .Z(n5534) );
  AND U8918 ( .A(n8900), .B(n5534), .Z(n12103) );
  ANDN U8919 ( .B(x[944]), .A(y[944]), .Z(n12107) );
  NANDN U8920 ( .A(x[956]), .B(y[956]), .Z(n8924) );
  NANDN U8921 ( .A(x[957]), .B(y[957]), .Z(n8926) );
  NAND U8922 ( .A(n8924), .B(n8926), .Z(n12133) );
  ANDN U8923 ( .B(x[957]), .A(y[957]), .Z(n12135) );
  NANDN U8924 ( .A(y[958]), .B(x[958]), .Z(n5531) );
  ANDN U8925 ( .B(y[959]), .A(x[959]), .Z(n5529) );
  NANDN U8926 ( .A(y[959]), .B(x[959]), .Z(n5530) );
  NANDN U8927 ( .A(x[960]), .B(y[960]), .Z(n5528) );
  NANDN U8928 ( .A(y[961]), .B(x[961]), .Z(n5527) );
  NANDN U8929 ( .A(y[974]), .B(x[974]), .Z(n12170) );
  NANDN U8930 ( .A(y[975]), .B(x[975]), .Z(n12175) );
  NANDN U8931 ( .A(y[977]), .B(x[977]), .Z(n5523) );
  NANDN U8932 ( .A(y[978]), .B(x[978]), .Z(n12183) );
  NAND U8933 ( .A(n5523), .B(n12183), .Z(n4415) );
  NANDN U8934 ( .A(x[980]), .B(y[980]), .Z(n8972) );
  NANDN U8935 ( .A(x[981]), .B(y[981]), .Z(n8977) );
  AND U8936 ( .A(n8972), .B(n8977), .Z(n12188) );
  ANDN U8937 ( .B(x[981]), .A(y[981]), .Z(n8974) );
  ANDN U8938 ( .B(x[982]), .A(y[982]), .Z(n8980) );
  NOR U8939 ( .A(n8974), .B(n8980), .Z(n12191) );
  NANDN U8940 ( .A(y[984]), .B(x[984]), .Z(n5521) );
  NANDN U8941 ( .A(x[984]), .B(y[984]), .Z(n12197) );
  IV U8942 ( .A(n12197), .Z(n8983) );
  NANDN U8943 ( .A(x[985]), .B(y[985]), .Z(n8985) );
  NANDN U8944 ( .A(y[986]), .B(x[986]), .Z(n8987) );
  NANDN U8945 ( .A(x[986]), .B(y[986]), .Z(n8984) );
  ANDN U8946 ( .B(x[988]), .A(y[988]), .Z(n5516) );
  NANDN U8947 ( .A(y[990]), .B(x[990]), .Z(n5515) );
  NANDN U8948 ( .A(y[992]), .B(x[992]), .Z(n5513) );
  NANDN U8949 ( .A(y[991]), .B(x[991]), .Z(n12213) );
  ANDN U8950 ( .B(x[993]), .A(y[993]), .Z(n5514) );
  ANDN U8951 ( .B(x[994]), .A(y[994]), .Z(n12222) );
  NANDN U8952 ( .A(x[994]), .B(y[994]), .Z(n8990) );
  NANDN U8953 ( .A(x[995]), .B(y[995]), .Z(n5512) );
  AND U8954 ( .A(n8990), .B(n5512), .Z(n12225) );
  NANDN U8955 ( .A(y[996]), .B(x[996]), .Z(n8993) );
  ANDN U8956 ( .B(x[995]), .A(y[995]), .Z(n12226) );
  IV U8957 ( .A(n12226), .Z(n8992) );
  AND U8958 ( .A(n8993), .B(n8992), .Z(n4418) );
  NANDN U8959 ( .A(x[996]), .B(y[996]), .Z(n12228) );
  IV U8960 ( .A(n12228), .Z(n5511) );
  NANDN U8961 ( .A(x[997]), .B(y[997]), .Z(n5509) );
  ANDN U8962 ( .B(x[998]), .A(y[998]), .Z(n5507) );
  XNOR U8963 ( .A(y[1000]), .B(x[1000]), .Z(n8995) );
  NANDN U8964 ( .A(x[1000]), .B(y[1000]), .Z(n4420) );
  ANDN U8965 ( .B(y[1001]), .A(x[1001]), .Z(n8998) );
  ANDN U8966 ( .B(n4420), .A(n8998), .Z(n12241) );
  NANDN U8967 ( .A(y[1001]), .B(x[1001]), .Z(n8996) );
  NANDN U8968 ( .A(y[1002]), .B(x[1002]), .Z(n8999) );
  NAND U8969 ( .A(n8996), .B(n8999), .Z(n12242) );
  NANDN U8970 ( .A(y[1008]), .B(x[1008]), .Z(n5503) );
  NANDN U8971 ( .A(y[1007]), .B(x[1007]), .Z(n12254) );
  NANDN U8972 ( .A(x[1009]), .B(y[1009]), .Z(n9010) );
  ANDN U8973 ( .B(x[1010]), .A(y[1010]), .Z(n9011) );
  NANDN U8974 ( .A(x[1011]), .B(y[1011]), .Z(n12264) );
  IV U8975 ( .A(n12264), .Z(n9014) );
  NANDN U8976 ( .A(y[1011]), .B(x[1011]), .Z(n9012) );
  NANDN U8977 ( .A(x[1012]), .B(y[1012]), .Z(n9013) );
  NANDN U8978 ( .A(x[1013]), .B(y[1013]), .Z(n9017) );
  AND U8979 ( .A(n9013), .B(n9017), .Z(n12269) );
  ANDN U8980 ( .B(x[1013]), .A(y[1013]), .Z(n9015) );
  ANDN U8981 ( .B(x[1014]), .A(y[1014]), .Z(n9020) );
  OR U8982 ( .A(n9015), .B(n9020), .Z(n12271) );
  ANDN U8983 ( .B(x[1022]), .A(y[1022]), .Z(n9033) );
  NANDN U8984 ( .A(x[1023]), .B(y[1023]), .Z(n12289) );
  ANDN U8985 ( .B(x[1024]), .A(y[1024]), .Z(n12290) );
  NANDN U8986 ( .A(y[1026]), .B(x[1026]), .Z(n5500) );
  ANDN U8987 ( .B(y[1027]), .A(x[1027]), .Z(n5498) );
  NANDN U8988 ( .A(y[1027]), .B(x[1027]), .Z(n5501) );
  ANDN U8989 ( .B(y[1029]), .A(x[1029]), .Z(n5494) );
  IV U8990 ( .A(n5494), .Z(n4425) );
  NANDN U8991 ( .A(x[1030]), .B(y[1030]), .Z(n5495) );
  ANDN U8992 ( .B(y[1031]), .A(x[1031]), .Z(n12308) );
  NANDN U8993 ( .A(y[1032]), .B(x[1032]), .Z(n12310) );
  NANDN U8994 ( .A(y[1034]), .B(x[1034]), .Z(n5490) );
  NANDN U8995 ( .A(x[1035]), .B(y[1035]), .Z(n5489) );
  NANDN U8996 ( .A(y[1035]), .B(x[1035]), .Z(n5491) );
  ANDN U8997 ( .B(y[1037]), .A(x[1037]), .Z(n5484) );
  NANDN U8998 ( .A(x[1038]), .B(y[1038]), .Z(n5485) );
  ANDN U8999 ( .B(y[1039]), .A(x[1039]), .Z(n12329) );
  IV U9000 ( .A(n12329), .Z(n9039) );
  NANDN U9001 ( .A(y[1040]), .B(x[1040]), .Z(n12331) );
  IV U9002 ( .A(n12331), .Z(n9042) );
  NANDN U9003 ( .A(y[1039]), .B(x[1039]), .Z(n5482) );
  NANDN U9004 ( .A(y[1041]), .B(x[1041]), .Z(n9043) );
  NANDN U9005 ( .A(y[1042]), .B(x[1042]), .Z(n9052) );
  AND U9006 ( .A(n9043), .B(n9052), .Z(n12334) );
  ANDN U9007 ( .B(y[1042]), .A(x[1042]), .Z(n9047) );
  ANDN U9008 ( .B(y[1043]), .A(x[1043]), .Z(n9057) );
  NOR U9009 ( .A(n9047), .B(n9057), .Z(n12337) );
  ANDN U9010 ( .B(x[1048]), .A(y[1048]), .Z(n5480) );
  ANDN U9011 ( .B(x[1047]), .A(y[1047]), .Z(n12346) );
  NANDN U9012 ( .A(x[1048]), .B(y[1048]), .Z(n12349) );
  NANDN U9013 ( .A(y[1049]), .B(x[1049]), .Z(n5479) );
  NANDN U9014 ( .A(y[1051]), .B(x[1051]), .Z(n12358) );
  ANDN U9015 ( .B(y[1053]), .A(x[1053]), .Z(n5474) );
  NANDN U9016 ( .A(x[1054]), .B(y[1054]), .Z(n5475) );
  NANDN U9017 ( .A(y[1056]), .B(x[1056]), .Z(n5468) );
  NANDN U9018 ( .A(x[1056]), .B(y[1056]), .Z(n5471) );
  NANDN U9019 ( .A(y[1058]), .B(x[1058]), .Z(n4430) );
  ANDN U9020 ( .B(n4430), .A(n4429), .Z(n12374) );
  ANDN U9021 ( .B(x[1060]), .A(y[1060]), .Z(n5467) );
  ANDN U9022 ( .B(x[1062]), .A(y[1062]), .Z(n5461) );
  NANDN U9023 ( .A(y[1061]), .B(x[1061]), .Z(n5466) );
  NANDN U9024 ( .A(y[1065]), .B(x[1065]), .Z(n5462) );
  ANDN U9025 ( .B(y[1066]), .A(x[1066]), .Z(n5458) );
  NANDN U9026 ( .A(y[1069]), .B(x[1069]), .Z(n12395) );
  IV U9027 ( .A(n12395), .Z(n5453) );
  NANDN U9028 ( .A(x[1071]), .B(y[1071]), .Z(n5448) );
  NANDN U9029 ( .A(y[1072]), .B(x[1072]), .Z(n5446) );
  ANDN U9030 ( .B(y[1073]), .A(x[1073]), .Z(n5445) );
  NANDN U9031 ( .A(y[1074]), .B(x[1074]), .Z(n12407) );
  NANDN U9032 ( .A(x[1075]), .B(y[1075]), .Z(n4434) );
  NAND U9033 ( .A(n4435), .B(n4434), .Z(n12408) );
  IV U9034 ( .A(n12408), .Z(n9099) );
  NANDN U9035 ( .A(x[1082]), .B(y[1082]), .Z(n5443) );
  NANDN U9036 ( .A(x[1083]), .B(y[1083]), .Z(n9108) );
  NAND U9037 ( .A(n5443), .B(n9108), .Z(n12425) );
  NANDN U9038 ( .A(y[1084]), .B(x[1084]), .Z(n5441) );
  ANDN U9039 ( .B(y[1085]), .A(x[1085]), .Z(n9109) );
  NANDN U9040 ( .A(y[1085]), .B(x[1085]), .Z(n5442) );
  ANDN U9041 ( .B(y[1086]), .A(x[1086]), .Z(n9110) );
  ANDN U9042 ( .B(x[1088]), .A(y[1088]), .Z(n12441) );
  NANDN U9043 ( .A(y[1087]), .B(x[1087]), .Z(n9112) );
  NANDN U9044 ( .A(x[1090]), .B(y[1090]), .Z(n9115) );
  NANDN U9045 ( .A(x[1091]), .B(y[1091]), .Z(n5440) );
  NAND U9046 ( .A(n9115), .B(n5440), .Z(n12447) );
  ANDN U9047 ( .B(x[1091]), .A(y[1091]), .Z(n12448) );
  NANDN U9048 ( .A(y[1092]), .B(x[1092]), .Z(n5438) );
  ANDN U9049 ( .B(y[1093]), .A(x[1093]), .Z(n12454) );
  NANDN U9050 ( .A(y[1094]), .B(x[1094]), .Z(n12457) );
  NANDN U9051 ( .A(y[1096]), .B(x[1096]), .Z(n9120) );
  NANDN U9052 ( .A(y[1098]), .B(x[1098]), .Z(n12468) );
  NANDN U9053 ( .A(y[1100]), .B(x[1100]), .Z(n9122) );
  NANDN U9054 ( .A(y[1102]), .B(x[1102]), .Z(n12480) );
  NANDN U9055 ( .A(y[1104]), .B(x[1104]), .Z(n5427) );
  NANDN U9056 ( .A(y[1105]), .B(x[1105]), .Z(n5428) );
  NANDN U9057 ( .A(x[1110]), .B(y[1110]), .Z(n9134) );
  NANDN U9058 ( .A(x[1111]), .B(y[1111]), .Z(n9138) );
  NAND U9059 ( .A(n9134), .B(n9138), .Z(n12503) );
  ANDN U9060 ( .B(x[1111]), .A(y[1111]), .Z(n12504) );
  ANDN U9061 ( .B(x[1114]), .A(y[1114]), .Z(n12513) );
  IV U9062 ( .A(n12513), .Z(n5423) );
  NANDN U9063 ( .A(x[1114]), .B(y[1114]), .Z(n9139) );
  NANDN U9064 ( .A(x[1115]), .B(y[1115]), .Z(n9141) );
  AND U9065 ( .A(n9139), .B(n9141), .Z(n12515) );
  NANDN U9066 ( .A(y[1116]), .B(x[1116]), .Z(n5422) );
  ANDN U9067 ( .B(x[1115]), .A(y[1115]), .Z(n12516) );
  IV U9068 ( .A(n12516), .Z(n5424) );
  ANDN U9069 ( .B(x[1118]), .A(y[1118]), .Z(n12525) );
  IV U9070 ( .A(n12525), .Z(n5420) );
  ANDN U9071 ( .B(x[1120]), .A(y[1120]), .Z(n5418) );
  NANDN U9072 ( .A(y[1121]), .B(x[1121]), .Z(n5419) );
  ANDN U9073 ( .B(x[1122]), .A(y[1122]), .Z(n12537) );
  IV U9074 ( .A(n12537), .Z(n4444) );
  NANDN U9075 ( .A(y[1123]), .B(x[1123]), .Z(n12541) );
  NANDN U9076 ( .A(x[1125]), .B(y[1125]), .Z(n5414) );
  NANDN U9077 ( .A(y[1126]), .B(x[1126]), .Z(n5413) );
  ANDN U9078 ( .B(y[1127]), .A(x[1127]), .Z(n12551) );
  NANDN U9079 ( .A(y[1128]), .B(x[1128]), .Z(n12553) );
  NANDN U9080 ( .A(y[1129]), .B(x[1129]), .Z(n12557) );
  ANDN U9081 ( .B(y[1131]), .A(x[1131]), .Z(n9150) );
  NANDN U9082 ( .A(y[1132]), .B(x[1132]), .Z(n9153) );
  NANDN U9083 ( .A(x[1133]), .B(y[1133]), .Z(n12566) );
  NANDN U9084 ( .A(y[1133]), .B(x[1133]), .Z(n9154) );
  NANDN U9085 ( .A(y[1136]), .B(x[1136]), .Z(n5409) );
  NANDN U9086 ( .A(y[1135]), .B(x[1135]), .Z(n12573) );
  NANDN U9087 ( .A(x[1136]), .B(y[1136]), .Z(n12575) );
  NANDN U9088 ( .A(x[1137]), .B(y[1137]), .Z(n9157) );
  ANDN U9089 ( .B(x[1138]), .A(y[1138]), .Z(n12580) );
  NANDN U9090 ( .A(x[1138]), .B(y[1138]), .Z(n9158) );
  ANDN U9091 ( .B(x[1143]), .A(y[1143]), .Z(n12592) );
  NANDN U9092 ( .A(x[1146]), .B(y[1146]), .Z(n9170) );
  NANDN U9093 ( .A(x[1147]), .B(y[1147]), .Z(n9172) );
  AND U9094 ( .A(n9170), .B(n9172), .Z(n12599) );
  ANDN U9095 ( .B(x[1148]), .A(y[1148]), .Z(n5407) );
  ANDN U9096 ( .B(x[1147]), .A(y[1147]), .Z(n12601) );
  ANDN U9097 ( .B(y[1149]), .A(x[1149]), .Z(n5404) );
  NANDN U9098 ( .A(y[1150]), .B(x[1150]), .Z(n12609) );
  IV U9099 ( .A(n12609), .Z(n9174) );
  ANDN U9100 ( .B(x[1154]), .A(y[1154]), .Z(n5402) );
  NANDN U9101 ( .A(x[1156]), .B(y[1156]), .Z(n5399) );
  ANDN U9102 ( .B(y[1157]), .A(x[1157]), .Z(n12626) );
  NANDN U9103 ( .A(y[1158]), .B(x[1158]), .Z(n12628) );
  NANDN U9104 ( .A(y[1157]), .B(x[1157]), .Z(n5397) );
  NANDN U9105 ( .A(y[1159]), .B(x[1159]), .Z(n12632) );
  IV U9106 ( .A(n12632), .Z(n4450) );
  NANDN U9107 ( .A(y[1160]), .B(x[1160]), .Z(n5396) );
  ANDN U9108 ( .B(y[1161]), .A(x[1161]), .Z(n9183) );
  NANDN U9109 ( .A(y[1161]), .B(x[1161]), .Z(n5395) );
  ANDN U9110 ( .B(y[1162]), .A(x[1162]), .Z(n9182) );
  NANDN U9111 ( .A(y[1166]), .B(x[1166]), .Z(n5391) );
  NANDN U9112 ( .A(y[1167]), .B(x[1167]), .Z(n5390) );
  NANDN U9113 ( .A(y[1176]), .B(x[1176]), .Z(n5384) );
  NANDN U9114 ( .A(y[1178]), .B(x[1178]), .Z(n12681) );
  IV U9115 ( .A(n12681), .Z(n5382) );
  NANDN U9116 ( .A(y[1180]), .B(x[1180]), .Z(n5380) );
  NANDN U9117 ( .A(y[1179]), .B(x[1179]), .Z(n12685) );
  NANDN U9118 ( .A(x[1181]), .B(y[1181]), .Z(n5378) );
  ANDN U9119 ( .B(x[1182]), .A(y[1182]), .Z(n9201) );
  NANDN U9120 ( .A(x[1183]), .B(y[1183]), .Z(n12695) );
  ANDN U9121 ( .B(x[1183]), .A(y[1183]), .Z(n9202) );
  NANDN U9122 ( .A(y[1185]), .B(x[1185]), .Z(n12700) );
  NANDN U9123 ( .A(y[1186]), .B(x[1186]), .Z(n5376) );
  NANDN U9124 ( .A(x[1187]), .B(y[1187]), .Z(n5375) );
  NANDN U9125 ( .A(y[1187]), .B(x[1187]), .Z(n5377) );
  ANDN U9126 ( .B(y[1189]), .A(x[1189]), .Z(n5372) );
  NANDN U9127 ( .A(x[1190]), .B(y[1190]), .Z(n5373) );
  ANDN U9128 ( .B(x[1192]), .A(y[1192]), .Z(n5364) );
  NANDN U9129 ( .A(y[1194]), .B(x[1194]), .Z(n4455) );
  NAND U9130 ( .A(n4456), .B(n4455), .Z(n12718) );
  ANDN U9131 ( .B(x[1198]), .A(y[1198]), .Z(n12729) );
  IV U9132 ( .A(n12729), .Z(n5360) );
  NANDN U9133 ( .A(x[1198]), .B(y[1198]), .Z(n12731) );
  IV U9134 ( .A(n12731), .Z(n4459) );
  ANDN U9135 ( .B(x[1200]), .A(y[1200]), .Z(n5356) );
  NANDN U9136 ( .A(y[1201]), .B(x[1201]), .Z(n5357) );
  NANDN U9137 ( .A(y[1203]), .B(x[1203]), .Z(n9212) );
  NANDN U9138 ( .A(y[1204]), .B(x[1204]), .Z(n9215) );
  NAND U9139 ( .A(n9212), .B(n9215), .Z(n12744) );
  NANDN U9140 ( .A(y[1208]), .B(x[1208]), .Z(n5353) );
  NANDN U9141 ( .A(x[1208]), .B(y[1208]), .Z(n12755) );
  ANDN U9142 ( .B(x[1210]), .A(y[1210]), .Z(n5350) );
  NANDN U9143 ( .A(y[1211]), .B(x[1211]), .Z(n5351) );
  NANDN U9144 ( .A(x[1213]), .B(y[1213]), .Z(n12767) );
  ANDN U9145 ( .B(x[1215]), .A(y[1215]), .Z(n12773) );
  NANDN U9146 ( .A(y[1216]), .B(x[1216]), .Z(n5349) );
  NANDN U9147 ( .A(x[1217]), .B(y[1217]), .Z(n12779) );
  NANDN U9148 ( .A(y[1218]), .B(x[1218]), .Z(n4463) );
  NAND U9149 ( .A(n4464), .B(n4463), .Z(n12780) );
  ANDN U9150 ( .B(x[1223]), .A(y[1223]), .Z(n12789) );
  NANDN U9151 ( .A(y[1224]), .B(x[1224]), .Z(n5347) );
  NANDN U9152 ( .A(x[1225]), .B(y[1225]), .Z(n12794) );
  NANDN U9153 ( .A(y[1225]), .B(x[1225]), .Z(n5346) );
  NANDN U9154 ( .A(y[1228]), .B(x[1228]), .Z(n9238) );
  NANDN U9155 ( .A(y[1230]), .B(x[1230]), .Z(n4467) );
  NANDN U9156 ( .A(y[1231]), .B(x[1231]), .Z(n4466) );
  AND U9157 ( .A(n4467), .B(n4466), .Z(n9243) );
  NANDN U9158 ( .A(y[1229]), .B(x[1229]), .Z(n9239) );
  NANDN U9159 ( .A(x[1232]), .B(y[1232]), .Z(n4470) );
  NANDN U9160 ( .A(x[1231]), .B(y[1231]), .Z(n4469) );
  NAND U9161 ( .A(n4470), .B(n4469), .Z(n12807) );
  ANDN U9162 ( .B(x[1235]), .A(y[1235]), .Z(n9245) );
  ANDN U9163 ( .B(x[1236]), .A(y[1236]), .Z(n9248) );
  NOR U9164 ( .A(n9245), .B(n9248), .Z(n12816) );
  NANDN U9165 ( .A(x[1236]), .B(y[1236]), .Z(n9246) );
  NANDN U9166 ( .A(x[1237]), .B(y[1237]), .Z(n9249) );
  NAND U9167 ( .A(n9246), .B(n9249), .Z(n12819) );
  NANDN U9168 ( .A(y[1240]), .B(x[1240]), .Z(n5344) );
  NANDN U9169 ( .A(y[1241]), .B(x[1241]), .Z(n5345) );
  ANDN U9170 ( .B(x[1243]), .A(y[1243]), .Z(n12836) );
  NANDN U9171 ( .A(x[1244]), .B(y[1244]), .Z(n12838) );
  ANDN U9172 ( .B(x[1246]), .A(y[1246]), .Z(n12845) );
  NANDN U9173 ( .A(y[1245]), .B(x[1245]), .Z(n5343) );
  NANDN U9174 ( .A(x[1249]), .B(y[1249]), .Z(n12854) );
  NANDN U9175 ( .A(y[1249]), .B(x[1249]), .Z(n5340) );
  NANDN U9176 ( .A(y[1251]), .B(x[1251]), .Z(n12861) );
  ANDN U9177 ( .B(y[1253]), .A(x[1253]), .Z(n5336) );
  NANDN U9178 ( .A(x[1254]), .B(y[1254]), .Z(n5337) );
  ANDN U9179 ( .B(y[1255]), .A(x[1255]), .Z(n12870) );
  NANDN U9180 ( .A(y[1256]), .B(x[1256]), .Z(n12872) );
  NANDN U9181 ( .A(y[1255]), .B(x[1255]), .Z(n9262) );
  ANDN U9182 ( .B(y[1259]), .A(x[1259]), .Z(n12883) );
  NANDN U9183 ( .A(y[1259]), .B(x[1259]), .Z(n5333) );
  NANDN U9184 ( .A(y[1261]), .B(x[1261]), .Z(n12888) );
  ANDN U9185 ( .B(y[1263]), .A(x[1263]), .Z(n5328) );
  NANDN U9186 ( .A(x[1264]), .B(y[1264]), .Z(n5329) );
  ANDN U9187 ( .B(x[1265]), .A(y[1265]), .Z(n5327) );
  ANDN U9188 ( .B(x[1267]), .A(y[1267]), .Z(n9266) );
  ANDN U9189 ( .B(x[1268]), .A(y[1268]), .Z(n9268) );
  NOR U9190 ( .A(n9266), .B(n9268), .Z(n12905) );
  NANDN U9191 ( .A(y[1272]), .B(x[1272]), .Z(n5317) );
  NANDN U9192 ( .A(y[1273]), .B(x[1273]), .Z(n5318) );
  NANDN U9193 ( .A(y[1274]), .B(x[1274]), .Z(n5322) );
  ANDN U9194 ( .B(y[1275]), .A(x[1275]), .Z(n12919) );
  IV U9195 ( .A(n12919), .Z(n4479) );
  ANDN U9196 ( .B(y[1279]), .A(x[1279]), .Z(n5313) );
  NANDN U9197 ( .A(y[1280]), .B(x[1280]), .Z(n5312) );
  ANDN U9198 ( .B(y[1281]), .A(x[1281]), .Z(n5310) );
  NANDN U9199 ( .A(y[1281]), .B(x[1281]), .Z(n5311) );
  ANDN U9200 ( .B(y[1283]), .A(x[1283]), .Z(n5306) );
  IV U9201 ( .A(n5306), .Z(n4481) );
  NANDN U9202 ( .A(x[1285]), .B(y[1285]), .Z(n12943) );
  NANDN U9203 ( .A(y[1287]), .B(x[1287]), .Z(n4484) );
  NANDN U9204 ( .A(y[1286]), .B(x[1286]), .Z(n4483) );
  AND U9205 ( .A(n4484), .B(n4483), .Z(n12945) );
  ANDN U9206 ( .B(y[1286]), .A(x[1286]), .Z(n9277) );
  NAND U9207 ( .A(n9277), .B(n4484), .Z(n4485) );
  ANDN U9208 ( .B(y[1289]), .A(x[1289]), .Z(n9282) );
  ANDN U9209 ( .B(n4485), .A(n9282), .Z(n4488) );
  NANDN U9210 ( .A(x[1287]), .B(y[1287]), .Z(n4487) );
  NANDN U9211 ( .A(x[1288]), .B(y[1288]), .Z(n4486) );
  NAND U9212 ( .A(n4487), .B(n4486), .Z(n9279) );
  ANDN U9213 ( .B(n4488), .A(n9279), .Z(n12947) );
  NANDN U9214 ( .A(y[1290]), .B(x[1290]), .Z(n5301) );
  NANDN U9215 ( .A(y[1288]), .B(x[1288]), .Z(n4490) );
  NANDN U9216 ( .A(y[1289]), .B(x[1289]), .Z(n4489) );
  AND U9217 ( .A(n4490), .B(n4489), .Z(n9280) );
  OR U9218 ( .A(n9280), .B(n9282), .Z(n4491) );
  AND U9219 ( .A(n5301), .B(n4491), .Z(n12949) );
  NANDN U9220 ( .A(y[1296]), .B(x[1296]), .Z(n5295) );
  ANDN U9221 ( .B(x[1300]), .A(y[1300]), .Z(n12969) );
  ANDN U9222 ( .B(x[1307]), .A(y[1307]), .Z(n12984) );
  NANDN U9223 ( .A(y[1308]), .B(x[1308]), .Z(n5293) );
  ANDN U9224 ( .B(y[1309]), .A(x[1309]), .Z(n12990) );
  IV U9225 ( .A(n12990), .Z(n4493) );
  NANDN U9226 ( .A(y[1310]), .B(x[1310]), .Z(n12993) );
  NANDN U9227 ( .A(y[1312]), .B(x[1312]), .Z(n5291) );
  NANDN U9228 ( .A(y[1311]), .B(x[1311]), .Z(n12997) );
  NANDN U9229 ( .A(x[1312]), .B(y[1312]), .Z(n12998) );
  IV U9230 ( .A(n12998), .Z(n9305) );
  NANDN U9231 ( .A(x[1313]), .B(y[1313]), .Z(n5288) );
  ANDN U9232 ( .B(x[1314]), .A(y[1314]), .Z(n5286) );
  NANDN U9233 ( .A(x[1315]), .B(y[1315]), .Z(n13007) );
  NANDN U9234 ( .A(y[1316]), .B(x[1316]), .Z(n5285) );
  NANDN U9235 ( .A(y[1318]), .B(x[1318]), .Z(n5282) );
  NANDN U9236 ( .A(x[1318]), .B(y[1318]), .Z(n13010) );
  ANDN U9237 ( .B(x[1320]), .A(y[1320]), .Z(n5279) );
  NANDN U9238 ( .A(x[1320]), .B(y[1320]), .Z(n5281) );
  ANDN U9239 ( .B(x[1322]), .A(y[1322]), .Z(n5274) );
  NANDN U9240 ( .A(x[1322]), .B(y[1322]), .Z(n5277) );
  NANDN U9241 ( .A(y[1324]), .B(x[1324]), .Z(n13028) );
  NANDN U9242 ( .A(y[1326]), .B(x[1326]), .Z(n5272) );
  NANDN U9243 ( .A(y[1327]), .B(x[1327]), .Z(n5271) );
  NANDN U9244 ( .A(y[1328]), .B(x[1328]), .Z(n13040) );
  IV U9245 ( .A(n13040), .Z(n9313) );
  NANDN U9246 ( .A(y[1329]), .B(x[1329]), .Z(n9312) );
  NANDN U9247 ( .A(y[1330]), .B(x[1330]), .Z(n9316) );
  NAND U9248 ( .A(n9312), .B(n9316), .Z(n13044) );
  ANDN U9249 ( .B(y[1341]), .A(x[1341]), .Z(n5267) );
  NANDN U9250 ( .A(y[1341]), .B(x[1341]), .Z(n5269) );
  NANDN U9251 ( .A(x[1342]), .B(y[1342]), .Z(n5268) );
  NANDN U9252 ( .A(y[1345]), .B(x[1345]), .Z(n13080) );
  ANDN U9253 ( .B(y[1347]), .A(x[1347]), .Z(n5260) );
  NANDN U9254 ( .A(y[1348]), .B(x[1348]), .Z(n5259) );
  ANDN U9255 ( .B(y[1349]), .A(x[1349]), .Z(n5256) );
  ANDN U9256 ( .B(y[1353]), .A(x[1353]), .Z(n13099) );
  ANDN U9257 ( .B(y[1359]), .A(x[1359]), .Z(n9349) );
  NANDN U9258 ( .A(y[1359]), .B(x[1359]), .Z(n13115) );
  ANDN U9259 ( .B(y[1361]), .A(x[1361]), .Z(n5250) );
  ANDN U9260 ( .B(x[1362]), .A(y[1362]), .Z(n13123) );
  ANDN U9261 ( .B(x[1363]), .A(y[1363]), .Z(n9353) );
  ANDN U9262 ( .B(x[1364]), .A(y[1364]), .Z(n9357) );
  NOR U9263 ( .A(n9353), .B(n9357), .Z(n13127) );
  ANDN U9264 ( .B(y[1369]), .A(x[1369]), .Z(n5246) );
  NANDN U9265 ( .A(y[1369]), .B(x[1369]), .Z(n5248) );
  NANDN U9266 ( .A(x[1370]), .B(y[1370]), .Z(n5247) );
  NANDN U9267 ( .A(y[1374]), .B(x[1374]), .Z(n5242) );
  ANDN U9268 ( .B(x[1378]), .A(y[1378]), .Z(n5240) );
  NANDN U9269 ( .A(x[1378]), .B(y[1378]), .Z(n13161) );
  NANDN U9270 ( .A(x[1381]), .B(y[1381]), .Z(n4506) );
  NANDN U9271 ( .A(x[1382]), .B(y[1382]), .Z(n4505) );
  NAND U9272 ( .A(n4506), .B(n4505), .Z(n13169) );
  NANDN U9273 ( .A(y[1385]), .B(x[1385]), .Z(n13179) );
  NANDN U9274 ( .A(y[1386]), .B(x[1386]), .Z(n5233) );
  ANDN U9275 ( .B(y[1387]), .A(x[1387]), .Z(n5231) );
  IV U9276 ( .A(n5231), .Z(n4508) );
  NANDN U9277 ( .A(y[1387]), .B(x[1387]), .Z(n5232) );
  NANDN U9278 ( .A(x[1388]), .B(y[1388]), .Z(n5230) );
  NANDN U9279 ( .A(y[1391]), .B(x[1391]), .Z(n13195) );
  ANDN U9280 ( .B(y[1393]), .A(x[1393]), .Z(n9377) );
  ANDN U9281 ( .B(x[1394]), .A(y[1394]), .Z(n13202) );
  NANDN U9282 ( .A(y[1395]), .B(x[1395]), .Z(n9378) );
  ANDN U9283 ( .B(x[1396]), .A(y[1396]), .Z(n9382) );
  ANDN U9284 ( .B(n9378), .A(n9382), .Z(n13207) );
  ANDN U9285 ( .B(x[1400]), .A(y[1400]), .Z(n5222) );
  NANDN U9286 ( .A(x[1400]), .B(y[1400]), .Z(n13216) );
  IV U9287 ( .A(n13216), .Z(n5224) );
  ANDN U9288 ( .B(x[1406]), .A(y[1406]), .Z(n13230) );
  NANDN U9289 ( .A(x[1406]), .B(y[1406]), .Z(n9390) );
  NANDN U9290 ( .A(x[1407]), .B(y[1407]), .Z(n5221) );
  NAND U9291 ( .A(n9390), .B(n5221), .Z(n13232) );
  ANDN U9292 ( .B(x[1407]), .A(y[1407]), .Z(n13234) );
  NANDN U9293 ( .A(y[1408]), .B(x[1408]), .Z(n9394) );
  NANDN U9294 ( .A(x[1409]), .B(y[1409]), .Z(n13240) );
  NANDN U9295 ( .A(y[1409]), .B(x[1409]), .Z(n9393) );
  NANDN U9296 ( .A(y[1411]), .B(x[1411]), .Z(n13247) );
  ANDN U9297 ( .B(y[1412]), .A(x[1412]), .Z(n13249) );
  NANDN U9298 ( .A(x[1414]), .B(y[1414]), .Z(n9398) );
  NANDN U9299 ( .A(x[1415]), .B(y[1415]), .Z(n5218) );
  NAND U9300 ( .A(n9398), .B(n5218), .Z(n13257) );
  ANDN U9301 ( .B(x[1418]), .A(y[1418]), .Z(n9407) );
  NANDN U9302 ( .A(y[1417]), .B(x[1417]), .Z(n9399) );
  NANDN U9303 ( .A(y[1421]), .B(x[1421]), .Z(n5215) );
  IV U9304 ( .A(n5215), .Z(n9405) );
  ANDN U9305 ( .B(y[1423]), .A(x[1423]), .Z(n5210) );
  NANDN U9306 ( .A(x[1425]), .B(y[1425]), .Z(n13273) );
  NANDN U9307 ( .A(x[1430]), .B(y[1430]), .Z(n5202) );
  ANDN U9308 ( .B(y[1431]), .A(x[1431]), .Z(n9415) );
  ANDN U9309 ( .B(n5202), .A(n9415), .Z(n13285) );
  IV U9310 ( .A(n13285), .Z(n4514) );
  NANDN U9311 ( .A(y[1431]), .B(x[1431]), .Z(n13286) );
  ANDN U9312 ( .B(x[1432]), .A(y[1432]), .Z(n5197) );
  IV U9313 ( .A(n5197), .Z(n4516) );
  NANDN U9314 ( .A(y[1437]), .B(x[1437]), .Z(n4518) );
  NANDN U9315 ( .A(y[1436]), .B(x[1436]), .Z(n4517) );
  AND U9316 ( .A(n4518), .B(n4517), .Z(n13299) );
  NANDN U9317 ( .A(x[1436]), .B(y[1436]), .Z(n13296) );
  NANDN U9318 ( .A(x[1437]), .B(y[1437]), .Z(n13301) );
  NANDN U9319 ( .A(y[1444]), .B(x[1444]), .Z(n5194) );
  NANDN U9320 ( .A(y[1443]), .B(x[1443]), .Z(n13315) );
  IV U9321 ( .A(n13315), .Z(n5196) );
  ANDN U9322 ( .B(n5194), .A(n5196), .Z(n4520) );
  NANDN U9323 ( .A(x[1444]), .B(y[1444]), .Z(n13317) );
  NANDN U9324 ( .A(y[1446]), .B(x[1446]), .Z(n9427) );
  NANDN U9325 ( .A(y[1447]), .B(x[1447]), .Z(n9428) );
  NANDN U9326 ( .A(y[1449]), .B(x[1449]), .Z(n13333) );
  ANDN U9327 ( .B(y[1451]), .A(x[1451]), .Z(n5188) );
  NANDN U9328 ( .A(x[1452]), .B(y[1452]), .Z(n5189) );
  ANDN U9329 ( .B(x[1454]), .A(y[1454]), .Z(n5183) );
  NANDN U9330 ( .A(y[1455]), .B(x[1455]), .Z(n5182) );
  ANDN U9331 ( .B(y[1457]), .A(x[1457]), .Z(n9432) );
  NANDN U9332 ( .A(y[1458]), .B(x[1458]), .Z(n13352) );
  IV U9333 ( .A(n13352), .Z(n5178) );
  NANDN U9334 ( .A(x[1464]), .B(y[1464]), .Z(n4523) );
  ANDN U9335 ( .B(y[1465]), .A(x[1465]), .Z(n5173) );
  ANDN U9336 ( .B(n4523), .A(n5173), .Z(n13367) );
  NANDN U9337 ( .A(y[1467]), .B(x[1467]), .Z(n13373) );
  ANDN U9338 ( .B(y[1469]), .A(x[1469]), .Z(n9442) );
  NANDN U9339 ( .A(y[1470]), .B(x[1470]), .Z(n9444) );
  ANDN U9340 ( .B(y[1471]), .A(x[1471]), .Z(n13383) );
  NANDN U9341 ( .A(y[1472]), .B(x[1472]), .Z(n13385) );
  NANDN U9342 ( .A(y[1474]), .B(x[1474]), .Z(n5165) );
  NANDN U9343 ( .A(y[1478]), .B(x[1478]), .Z(n5164) );
  ANDN U9344 ( .B(x[1479]), .A(y[1479]), .Z(n5163) );
  ANDN U9345 ( .B(y[1497]), .A(x[1497]), .Z(n13435) );
  NANDN U9346 ( .A(y[1497]), .B(x[1497]), .Z(n5157) );
  NANDN U9347 ( .A(n13439), .B(n4526), .Z(n4527) );
  AND U9348 ( .A(n5154), .B(n4527), .Z(n4528) );
  NANDN U9349 ( .A(n13441), .B(n4528), .Z(n4529) );
  NANDN U9350 ( .A(n4530), .B(n4529), .Z(n4531) );
  NANDN U9351 ( .A(y[1501]), .B(x[1501]), .Z(n5153) );
  AND U9352 ( .A(n4531), .B(n5153), .Z(n4532) );
  NANDN U9353 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U9354 ( .A(n4535), .B(n4534), .Z(n4537) );
  ANDN U9355 ( .B(y[1503]), .A(x[1503]), .Z(n5149) );
  IV U9356 ( .A(n5149), .Z(n4536) );
  NANDN U9357 ( .A(n4537), .B(n4536), .Z(n4538) );
  NANDN U9358 ( .A(y[1503]), .B(x[1503]), .Z(n13453) );
  IV U9359 ( .A(n13453), .Z(n5151) );
  ANDN U9360 ( .B(n4538), .A(n5151), .Z(n4539) );
  NAND U9361 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U9362 ( .A(n5150), .B(n4541), .Z(n4542) );
  NANDN U9363 ( .A(n9458), .B(n4542), .Z(n4543) );
  NANDN U9364 ( .A(n13458), .B(n4543), .Z(n4544) );
  NANDN U9365 ( .A(n9460), .B(n4544), .Z(n4545) );
  NAND U9366 ( .A(n13463), .B(n4545), .Z(n4551) );
  NANDN U9367 ( .A(y[1510]), .B(x[1510]), .Z(n4546) );
  ANDN U9368 ( .B(x[1511]), .A(y[1511]), .Z(n4556) );
  ANDN U9369 ( .B(n4546), .A(n4556), .Z(n9464) );
  NANDN U9370 ( .A(y[1509]), .B(x[1509]), .Z(n4548) );
  NANDN U9371 ( .A(y[1508]), .B(x[1508]), .Z(n4547) );
  AND U9372 ( .A(n4548), .B(n4547), .Z(n9462) );
  NANDN U9373 ( .A(n9462), .B(n5148), .Z(n4549) );
  AND U9374 ( .A(n9464), .B(n4549), .Z(n13464) );
  IV U9375 ( .A(n13464), .Z(n4550) );
  NANDN U9376 ( .A(x[1512]), .B(y[1512]), .Z(n4553) );
  NANDN U9377 ( .A(x[1511]), .B(y[1511]), .Z(n4552) );
  AND U9378 ( .A(n4553), .B(n4552), .Z(n4555) );
  AND U9379 ( .A(n4555), .B(n4554), .Z(n9465) );
  NANDN U9380 ( .A(x[1510]), .B(y[1510]), .Z(n5147) );
  OR U9381 ( .A(n4556), .B(n5147), .Z(n4557) );
  AND U9382 ( .A(n9465), .B(n4557), .Z(n13467) );
  NANDN U9383 ( .A(y[1516]), .B(x[1516]), .Z(n9467) );
  NANDN U9384 ( .A(x[1519]), .B(y[1519]), .Z(n4559) );
  NANDN U9385 ( .A(x[1518]), .B(y[1518]), .Z(n4558) );
  AND U9386 ( .A(n4559), .B(n4558), .Z(n9471) );
  ANDN U9387 ( .B(x[1520]), .A(y[1520]), .Z(n5141) );
  ANDN U9388 ( .B(x[1519]), .A(y[1519]), .Z(n9472) );
  ANDN U9389 ( .B(y[1520]), .A(x[1520]), .Z(n9473) );
  NANDN U9390 ( .A(y[1521]), .B(x[1521]), .Z(n5142) );
  NANDN U9391 ( .A(y[1527]), .B(x[1527]), .Z(n13493) );
  ANDN U9392 ( .B(y[1529]), .A(x[1529]), .Z(n5131) );
  NANDN U9393 ( .A(x[1531]), .B(y[1531]), .Z(n13503) );
  ANDN U9394 ( .B(x[1531]), .A(y[1531]), .Z(n5130) );
  ANDN U9395 ( .B(x[1533]), .A(y[1533]), .Z(n13508) );
  IV U9396 ( .A(n13508), .Z(n9481) );
  ANDN U9397 ( .B(x[1534]), .A(y[1534]), .Z(n5127) );
  NANDN U9398 ( .A(y[1536]), .B(x[1536]), .Z(n13516) );
  IV U9399 ( .A(n13516), .Z(n5124) );
  NANDN U9400 ( .A(y[1537]), .B(x[1537]), .Z(n13521) );
  ANDN U9401 ( .B(y[1539]), .A(x[1539]), .Z(n5119) );
  NANDN U9402 ( .A(x[1541]), .B(y[1541]), .Z(n13530) );
  IV U9403 ( .A(n13530), .Z(n5115) );
  ANDN U9404 ( .B(x[1541]), .A(y[1541]), .Z(n5117) );
  ANDN U9405 ( .B(x[1543]), .A(y[1543]), .Z(n13537) );
  NANDN U9406 ( .A(x[1548]), .B(y[1548]), .Z(n9488) );
  ANDN U9407 ( .B(x[1550]), .A(y[1550]), .Z(n5107) );
  NANDN U9408 ( .A(x[1552]), .B(y[1552]), .Z(n5106) );
  NANDN U9409 ( .A(x[1553]), .B(y[1553]), .Z(n5103) );
  NAND U9410 ( .A(n5106), .B(n5103), .Z(n13558) );
  ANDN U9411 ( .B(x[1560]), .A(y[1560]), .Z(n5094) );
  NANDN U9412 ( .A(y[1562]), .B(x[1562]), .Z(n13578) );
  NANDN U9413 ( .A(y[1563]), .B(x[1563]), .Z(n13583) );
  IV U9414 ( .A(n13583), .Z(n5092) );
  NANDN U9415 ( .A(y[1564]), .B(x[1564]), .Z(n5087) );
  NANDN U9416 ( .A(x[1564]), .B(y[1564]), .Z(n4567) );
  ANDN U9417 ( .B(y[1565]), .A(x[1565]), .Z(n5088) );
  ANDN U9418 ( .B(n4567), .A(n5088), .Z(n13585) );
  NANDN U9419 ( .A(y[1568]), .B(x[1568]), .Z(n5086) );
  NANDN U9420 ( .A(y[1569]), .B(x[1569]), .Z(n5085) );
  NANDN U9421 ( .A(y[1572]), .B(x[1572]), .Z(n5081) );
  NANDN U9422 ( .A(y[1573]), .B(x[1573]), .Z(n5083) );
  NAND U9423 ( .A(n9518), .B(n4568), .Z(n4569) );
  NAND U9424 ( .A(n13612), .B(n4569), .Z(n4570) );
  NANDN U9425 ( .A(x[1574]), .B(y[1574]), .Z(n13609) );
  NANDN U9426 ( .A(n4570), .B(n13609), .Z(n4571) );
  AND U9427 ( .A(n4572), .B(n4571), .Z(n4573) );
  ANDN U9428 ( .B(y[1577]), .A(x[1577]), .Z(n5077) );
  NANDN U9429 ( .A(x[1576]), .B(y[1576]), .Z(n5079) );
  NANDN U9430 ( .A(n5077), .B(n5079), .Z(n13617) );
  OR U9431 ( .A(n4573), .B(n13617), .Z(n4574) );
  ANDN U9432 ( .B(x[1577]), .A(y[1577]), .Z(n13619) );
  ANDN U9433 ( .B(n4574), .A(n13619), .Z(n4575) );
  NANDN U9434 ( .A(y[1578]), .B(x[1578]), .Z(n9523) );
  NAND U9435 ( .A(n4575), .B(n9523), .Z(n4576) );
  NANDN U9436 ( .A(n4577), .B(n4576), .Z(n4578) );
  AND U9437 ( .A(n9522), .B(n4578), .Z(n4579) );
  NAND U9438 ( .A(n13626), .B(n4579), .Z(n4580) );
  NAND U9439 ( .A(n13629), .B(n4580), .Z(n4581) );
  NAND U9440 ( .A(n13630), .B(n4581), .Z(n4584) );
  NANDN U9441 ( .A(x[1585]), .B(y[1585]), .Z(n4583) );
  NANDN U9442 ( .A(x[1584]), .B(y[1584]), .Z(n4582) );
  NAND U9443 ( .A(n4583), .B(n4582), .Z(n13633) );
  ANDN U9444 ( .B(n4584), .A(n13633), .Z(n4587) );
  NANDN U9445 ( .A(y[1585]), .B(x[1585]), .Z(n4586) );
  NANDN U9446 ( .A(y[1586]), .B(x[1586]), .Z(n4585) );
  AND U9447 ( .A(n4586), .B(n4585), .Z(n13635) );
  NANDN U9448 ( .A(n4587), .B(n13635), .Z(n4588) );
  NANDN U9449 ( .A(n13636), .B(n4588), .Z(n4589) );
  NAND U9450 ( .A(n13638), .B(n4589), .Z(n4590) );
  NANDN U9451 ( .A(n13641), .B(n4590), .Z(n4591) );
  NANDN U9452 ( .A(n9529), .B(n4591), .Z(n4592) );
  ANDN U9453 ( .B(x[1590]), .A(y[1590]), .Z(n13643) );
  NANDN U9454 ( .A(y[1591]), .B(x[1591]), .Z(n13649) );
  NANDN U9455 ( .A(x[1593]), .B(y[1593]), .Z(n5074) );
  NANDN U9456 ( .A(y[1594]), .B(x[1594]), .Z(n5071) );
  ANDN U9457 ( .B(y[1595]), .A(x[1595]), .Z(n5069) );
  NANDN U9458 ( .A(y[1595]), .B(x[1595]), .Z(n5072) );
  NANDN U9459 ( .A(x[1596]), .B(y[1596]), .Z(n5070) );
  ANDN U9460 ( .B(y[1599]), .A(x[1599]), .Z(n9533) );
  NANDN U9461 ( .A(x[1598]), .B(y[1598]), .Z(n5068) );
  NANDN U9462 ( .A(n9533), .B(n5068), .Z(n13669) );
  NANDN U9463 ( .A(x[1600]), .B(y[1600]), .Z(n13667) );
  IV U9464 ( .A(n13667), .Z(n4596) );
  NANDN U9465 ( .A(x[1601]), .B(y[1601]), .Z(n13674) );
  NANDN U9466 ( .A(y[1606]), .B(x[1606]), .Z(n13688) );
  NANDN U9467 ( .A(y[1605]), .B(x[1605]), .Z(n5063) );
  NANDN U9468 ( .A(y[1607]), .B(x[1607]), .Z(n13692) );
  NANDN U9469 ( .A(y[1608]), .B(x[1608]), .Z(n5061) );
  ANDN U9470 ( .B(y[1609]), .A(x[1609]), .Z(n9537) );
  NANDN U9471 ( .A(y[1609]), .B(x[1609]), .Z(n5060) );
  ANDN U9472 ( .B(y[1611]), .A(x[1611]), .Z(n5058) );
  NANDN U9473 ( .A(x[1612]), .B(y[1612]), .Z(n5059) );
  NANDN U9474 ( .A(x[1613]), .B(y[1613]), .Z(n13707) );
  NANDN U9475 ( .A(y[1614]), .B(x[1614]), .Z(n13709) );
  NANDN U9476 ( .A(y[1615]), .B(x[1615]), .Z(n13713) );
  NANDN U9477 ( .A(x[1618]), .B(y[1618]), .Z(n4600) );
  NANDN U9478 ( .A(x[1617]), .B(y[1617]), .Z(n4599) );
  NAND U9479 ( .A(n4600), .B(n4599), .Z(n13719) );
  NANDN U9480 ( .A(x[1619]), .B(y[1619]), .Z(n13723) );
  ANDN U9481 ( .B(y[1625]), .A(x[1625]), .Z(n5045) );
  NANDN U9482 ( .A(y[1625]), .B(x[1625]), .Z(n5047) );
  ANDN U9483 ( .B(y[1626]), .A(x[1626]), .Z(n5046) );
  ANDN U9484 ( .B(x[1629]), .A(y[1629]), .Z(n13751) );
  ANDN U9485 ( .B(y[1631]), .A(x[1631]), .Z(n5041) );
  NANDN U9486 ( .A(y[1632]), .B(x[1632]), .Z(n5038) );
  ANDN U9487 ( .B(y[1633]), .A(x[1633]), .Z(n5037) );
  ANDN U9488 ( .B(y[1635]), .A(x[1635]), .Z(n13765) );
  IV U9489 ( .A(n13765), .Z(n9553) );
  ANDN U9490 ( .B(y[1637]), .A(x[1637]), .Z(n9556) );
  IV U9491 ( .A(n9556), .Z(n4603) );
  ANDN U9492 ( .B(y[1639]), .A(x[1639]), .Z(n5030) );
  NANDN U9493 ( .A(y[1640]), .B(x[1640]), .Z(n5028) );
  NANDN U9494 ( .A(x[1640]), .B(y[1640]), .Z(n5031) );
  ANDN U9495 ( .B(x[1641]), .A(y[1641]), .Z(n5029) );
  ANDN U9496 ( .B(y[1643]), .A(x[1643]), .Z(n13783) );
  NANDN U9497 ( .A(y[1646]), .B(x[1646]), .Z(n5025) );
  NANDN U9498 ( .A(y[1647]), .B(x[1647]), .Z(n5024) );
  NANDN U9499 ( .A(x[1655]), .B(y[1655]), .Z(n5014) );
  ANDN U9500 ( .B(y[1656]), .A(x[1656]), .Z(n5015) );
  ANDN U9501 ( .B(y[1657]), .A(x[1657]), .Z(n13819) );
  NANDN U9502 ( .A(y[1657]), .B(x[1657]), .Z(n5012) );
  ANDN U9503 ( .B(y[1661]), .A(x[1661]), .Z(n9592) );
  NANDN U9504 ( .A(x[1660]), .B(y[1660]), .Z(n4606) );
  NANDN U9505 ( .A(n9592), .B(n4606), .Z(n13827) );
  NANDN U9506 ( .A(y[1661]), .B(x[1661]), .Z(n9586) );
  NANDN U9507 ( .A(y[1662]), .B(x[1662]), .Z(n9594) );
  AND U9508 ( .A(n9586), .B(n9594), .Z(n13829) );
  NANDN U9509 ( .A(x[1663]), .B(y[1663]), .Z(n5010) );
  ANDN U9510 ( .B(y[1662]), .A(x[1662]), .Z(n9590) );
  ANDN U9511 ( .B(n5010), .A(n9590), .Z(n13831) );
  NANDN U9512 ( .A(y[1663]), .B(x[1663]), .Z(n13832) );
  NANDN U9513 ( .A(y[1664]), .B(x[1664]), .Z(n5008) );
  NANDN U9514 ( .A(x[1665]), .B(y[1665]), .Z(n5007) );
  NANDN U9515 ( .A(y[1666]), .B(x[1666]), .Z(n5004) );
  NANDN U9516 ( .A(x[1667]), .B(y[1667]), .Z(n5003) );
  NANDN U9517 ( .A(y[1668]), .B(x[1668]), .Z(n13844) );
  ANDN U9518 ( .B(y[1668]), .A(x[1668]), .Z(n5002) );
  IV U9519 ( .A(n5002), .Z(n4608) );
  NANDN U9520 ( .A(y[1670]), .B(x[1670]), .Z(n5000) );
  ANDN U9521 ( .B(x[1669]), .A(y[1669]), .Z(n9604) );
  ANDN U9522 ( .B(n5000), .A(n9604), .Z(n13849) );
  NANDN U9523 ( .A(x[1670]), .B(y[1670]), .Z(n5001) );
  NANDN U9524 ( .A(x[1671]), .B(y[1671]), .Z(n4998) );
  NAND U9525 ( .A(n5001), .B(n4998), .Z(n13850) );
  NANDN U9526 ( .A(x[1677]), .B(y[1677]), .Z(n4996) );
  NANDN U9527 ( .A(x[1676]), .B(y[1676]), .Z(n13863) );
  IV U9528 ( .A(n13863), .Z(n9620) );
  ANDN U9529 ( .B(x[1677]), .A(y[1677]), .Z(n13865) );
  NANDN U9530 ( .A(y[1678]), .B(x[1678]), .Z(n4995) );
  ANDN U9531 ( .B(y[1679]), .A(x[1679]), .Z(n13871) );
  NANDN U9532 ( .A(y[1679]), .B(x[1679]), .Z(n4994) );
  NANDN U9533 ( .A(n13875), .B(n4610), .Z(n4611) );
  AND U9534 ( .A(n13877), .B(n4611), .Z(n4612) );
  OR U9535 ( .A(n13879), .B(n4612), .Z(n4613) );
  NAND U9536 ( .A(n13881), .B(n4613), .Z(n4614) );
  NANDN U9537 ( .A(n13882), .B(n4614), .Z(n4615) );
  NANDN U9538 ( .A(y[1685]), .B(x[1685]), .Z(n13885) );
  AND U9539 ( .A(n4615), .B(n13885), .Z(n4616) );
  NAND U9540 ( .A(n4992), .B(n4616), .Z(n4617) );
  NANDN U9541 ( .A(n13887), .B(n4617), .Z(n4618) );
  AND U9542 ( .A(n4993), .B(n4618), .Z(n4619) );
  OR U9543 ( .A(n13891), .B(n4619), .Z(n4620) );
  NAND U9544 ( .A(n13893), .B(n4620), .Z(n4621) );
  NANDN U9545 ( .A(n13895), .B(n4621), .Z(n4622) );
  NANDN U9546 ( .A(n13896), .B(n4622), .Z(n4623) );
  NAND U9547 ( .A(n13898), .B(n4623), .Z(n4624) );
  AND U9548 ( .A(n13901), .B(n4624), .Z(n4625) );
  NANDN U9549 ( .A(x[1692]), .B(y[1692]), .Z(n4991) );
  NANDN U9550 ( .A(x[1693]), .B(y[1693]), .Z(n9633) );
  NAND U9551 ( .A(n4991), .B(n9633), .Z(n13903) );
  OR U9552 ( .A(n4625), .B(n13903), .Z(n4626) );
  NANDN U9553 ( .A(y[1693]), .B(x[1693]), .Z(n10185) );
  AND U9554 ( .A(n4626), .B(n10185), .Z(n4629) );
  NANDN U9555 ( .A(x[1694]), .B(y[1694]), .Z(n4627) );
  AND U9556 ( .A(n4628), .B(n4627), .Z(n13906) );
  IV U9557 ( .A(n13906), .Z(n9634) );
  OR U9558 ( .A(n4629), .B(n9634), .Z(n4630) );
  NANDN U9559 ( .A(n9635), .B(n4630), .Z(n4633) );
  NANDN U9560 ( .A(x[1697]), .B(y[1697]), .Z(n4632) );
  NANDN U9561 ( .A(x[1698]), .B(y[1698]), .Z(n4631) );
  AND U9562 ( .A(n4632), .B(n4631), .Z(n13910) );
  IV U9563 ( .A(n13910), .Z(n9636) );
  ANDN U9564 ( .B(n4633), .A(n9636), .Z(n4636) );
  NANDN U9565 ( .A(y[1699]), .B(x[1699]), .Z(n4635) );
  NANDN U9566 ( .A(y[1698]), .B(x[1698]), .Z(n4634) );
  NAND U9567 ( .A(n4635), .B(n4634), .Z(n13913) );
  IV U9568 ( .A(n13913), .Z(n9637) );
  NANDN U9569 ( .A(x[1699]), .B(y[1699]), .Z(n4638) );
  NANDN U9570 ( .A(x[1700]), .B(y[1700]), .Z(n4637) );
  AND U9571 ( .A(n4638), .B(n4637), .Z(n13915) );
  IV U9572 ( .A(n13915), .Z(n9638) );
  ANDN U9573 ( .B(x[1700]), .A(y[1700]), .Z(n9639) );
  NANDN U9574 ( .A(y[1701]), .B(x[1701]), .Z(n9640) );
  NANDN U9575 ( .A(x[1702]), .B(y[1702]), .Z(n4990) );
  NANDN U9576 ( .A(x[1703]), .B(y[1703]), .Z(n4987) );
  AND U9577 ( .A(n4990), .B(n4987), .Z(n13922) );
  NANDN U9578 ( .A(y[1704]), .B(x[1704]), .Z(n4986) );
  ANDN U9579 ( .B(x[1703]), .A(y[1703]), .Z(n9642) );
  ANDN U9580 ( .B(n4986), .A(n9642), .Z(n13925) );
  ANDN U9581 ( .B(x[1708]), .A(y[1708]), .Z(n9646) );
  ANDN U9582 ( .B(y[1708]), .A(x[1708]), .Z(n13935) );
  NANDN U9583 ( .A(x[1709]), .B(y[1709]), .Z(n9649) );
  ANDN U9584 ( .B(y[1713]), .A(x[1713]), .Z(n13947) );
  NANDN U9585 ( .A(x[1712]), .B(y[1712]), .Z(n4979) );
  NANDN U9586 ( .A(y[1719]), .B(x[1719]), .Z(n9657) );
  NANDN U9587 ( .A(y[1720]), .B(x[1720]), .Z(n9659) );
  AND U9588 ( .A(n9657), .B(n9659), .Z(n13961) );
  ANDN U9589 ( .B(y[1721]), .A(x[1721]), .Z(n9661) );
  ANDN U9590 ( .B(y[1720]), .A(x[1720]), .Z(n13963) );
  ANDN U9591 ( .B(x[1722]), .A(y[1722]), .Z(n9663) );
  IV U9592 ( .A(n9663), .Z(n4640) );
  NANDN U9593 ( .A(x[1728]), .B(y[1728]), .Z(n4964) );
  ANDN U9594 ( .B(y[1729]), .A(x[1729]), .Z(n9668) );
  ANDN U9595 ( .B(n4964), .A(n9668), .Z(n13983) );
  NANDN U9596 ( .A(y[1730]), .B(x[1730]), .Z(n4961) );
  ANDN U9597 ( .B(x[1729]), .A(y[1729]), .Z(n13985) );
  ANDN U9598 ( .B(y[1731]), .A(x[1731]), .Z(n4960) );
  NANDN U9599 ( .A(y[1732]), .B(x[1732]), .Z(n4958) );
  NANDN U9600 ( .A(x[1733]), .B(y[1733]), .Z(n4955) );
  NANDN U9601 ( .A(y[1733]), .B(x[1733]), .Z(n4957) );
  ANDN U9602 ( .B(y[1734]), .A(x[1734]), .Z(n4956) );
  ANDN U9603 ( .B(y[1735]), .A(x[1735]), .Z(n13999) );
  NANDN U9604 ( .A(y[1735]), .B(x[1735]), .Z(n9669) );
  ANDN U9605 ( .B(x[1736]), .A(y[1736]), .Z(n9674) );
  ANDN U9606 ( .B(n9669), .A(n9674), .Z(n14001) );
  NANDN U9607 ( .A(x[1743]), .B(y[1743]), .Z(n9680) );
  ANDN U9608 ( .B(x[1743]), .A(y[1743]), .Z(n14017) );
  ANDN U9609 ( .B(y[1744]), .A(x[1744]), .Z(n9679) );
  ANDN U9610 ( .B(x[1746]), .A(y[1746]), .Z(n14024) );
  NANDN U9611 ( .A(x[1746]), .B(y[1746]), .Z(n4948) );
  NANDN U9612 ( .A(x[1747]), .B(y[1747]), .Z(n4946) );
  AND U9613 ( .A(n4948), .B(n4946), .Z(n14026) );
  NANDN U9614 ( .A(y[1748]), .B(x[1748]), .Z(n4945) );
  ANDN U9615 ( .B(x[1747]), .A(y[1747]), .Z(n9685) );
  ANDN U9616 ( .B(n4945), .A(n9685), .Z(n14029) );
  ANDN U9617 ( .B(x[1752]), .A(y[1752]), .Z(n9687) );
  ANDN U9618 ( .B(y[1752]), .A(x[1752]), .Z(n14039) );
  NANDN U9619 ( .A(x[1753]), .B(y[1753]), .Z(n4940) );
  NANDN U9620 ( .A(y[1754]), .B(x[1754]), .Z(n4938) );
  NANDN U9621 ( .A(x[1755]), .B(y[1755]), .Z(n4936) );
  NANDN U9622 ( .A(y[1756]), .B(x[1756]), .Z(n14049) );
  ANDN U9623 ( .B(y[1756]), .A(x[1756]), .Z(n4937) );
  NANDN U9624 ( .A(y[1761]), .B(x[1761]), .Z(n4932) );
  NANDN U9625 ( .A(y[1762]), .B(x[1762]), .Z(n4929) );
  AND U9626 ( .A(n4932), .B(n4929), .Z(n14061) );
  NANDN U9627 ( .A(x[1762]), .B(y[1762]), .Z(n4931) );
  NANDN U9628 ( .A(x[1763]), .B(y[1763]), .Z(n9708) );
  NAND U9629 ( .A(n4931), .B(n9708), .Z(n14062) );
  ANDN U9630 ( .B(x[1765]), .A(y[1765]), .Z(n4645) );
  NAND U9631 ( .A(n4645), .B(x[1766]), .Z(n4648) );
  XOR U9632 ( .A(n4645), .B(x[1766]), .Z(n4646) );
  NANDN U9633 ( .A(y[1766]), .B(n4646), .Z(n4647) );
  AND U9634 ( .A(n4648), .B(n4647), .Z(n14070) );
  IV U9635 ( .A(n14070), .Z(n4926) );
  ANDN U9636 ( .B(y[1767]), .A(x[1767]), .Z(n9718) );
  IV U9637 ( .A(n9718), .Z(n4649) );
  NANDN U9638 ( .A(x[1768]), .B(y[1768]), .Z(n9719) );
  ANDN U9639 ( .B(y[1772]), .A(x[1772]), .Z(n9730) );
  ANDN U9640 ( .B(y[1773]), .A(x[1773]), .Z(n9738) );
  NOR U9641 ( .A(n9730), .B(n9738), .Z(n14083) );
  NANDN U9642 ( .A(y[1774]), .B(x[1774]), .Z(n4923) );
  ANDN U9643 ( .B(x[1773]), .A(y[1773]), .Z(n14085) );
  NANDN U9644 ( .A(x[1774]), .B(y[1774]), .Z(n14087) );
  NANDN U9645 ( .A(x[1775]), .B(y[1775]), .Z(n4922) );
  NANDN U9646 ( .A(y[1775]), .B(x[1775]), .Z(n4924) );
  ANDN U9647 ( .B(x[1776]), .A(y[1776]), .Z(n4919) );
  NANDN U9648 ( .A(x[1777]), .B(y[1777]), .Z(n4917) );
  ANDN U9649 ( .B(x[1778]), .A(y[1778]), .Z(n14097) );
  NANDN U9650 ( .A(x[1779]), .B(y[1779]), .Z(n14099) );
  NANDN U9651 ( .A(x[1778]), .B(y[1778]), .Z(n4918) );
  NANDN U9652 ( .A(y[1779]), .B(x[1779]), .Z(n9744) );
  NANDN U9653 ( .A(y[1780]), .B(x[1780]), .Z(n9750) );
  AND U9654 ( .A(n9744), .B(n9750), .Z(n14101) );
  ANDN U9655 ( .B(y[1787]), .A(x[1787]), .Z(n4913) );
  ANDN U9656 ( .B(x[1787]), .A(y[1787]), .Z(n14116) );
  ANDN U9657 ( .B(y[1788]), .A(x[1788]), .Z(n4912) );
  NANDN U9658 ( .A(x[1801]), .B(y[1801]), .Z(n14146) );
  NANDN U9659 ( .A(y[1808]), .B(x[1808]), .Z(n4655) );
  NANDN U9660 ( .A(y[1807]), .B(x[1807]), .Z(n4654) );
  NAND U9661 ( .A(n4655), .B(n4654), .Z(n14161) );
  NANDN U9662 ( .A(x[1808]), .B(y[1808]), .Z(n14163) );
  NANDN U9663 ( .A(y[1810]), .B(x[1810]), .Z(n9805) );
  NANDN U9664 ( .A(x[1811]), .B(y[1811]), .Z(n14171) );
  IV U9665 ( .A(n14171), .Z(n4898) );
  ANDN U9666 ( .B(x[1811]), .A(y[1811]), .Z(n9804) );
  NANDN U9667 ( .A(x[1812]), .B(y[1812]), .Z(n4899) );
  NANDN U9668 ( .A(x[1813]), .B(y[1813]), .Z(n4896) );
  AND U9669 ( .A(n4899), .B(n4896), .Z(n14174) );
  NANDN U9670 ( .A(y[1814]), .B(x[1814]), .Z(n9816) );
  ANDN U9671 ( .B(x[1813]), .A(y[1813]), .Z(n9810) );
  ANDN U9672 ( .B(n9816), .A(n9810), .Z(n14177) );
  ANDN U9673 ( .B(y[1819]), .A(x[1819]), .Z(n9823) );
  NANDN U9674 ( .A(y[1822]), .B(x[1822]), .Z(n14197) );
  IV U9675 ( .A(n14197), .Z(n9825) );
  ANDN U9676 ( .B(y[1822]), .A(x[1822]), .Z(n4890) );
  NANDN U9677 ( .A(y[1823]), .B(x[1823]), .Z(n9826) );
  ANDN U9678 ( .B(x[1824]), .A(y[1824]), .Z(n9830) );
  ANDN U9679 ( .B(n9826), .A(n9830), .Z(n14201) );
  NANDN U9680 ( .A(x[1825]), .B(y[1825]), .Z(n4888) );
  ANDN U9681 ( .B(y[1824]), .A(x[1824]), .Z(n9827) );
  ANDN U9682 ( .B(n4888), .A(n9827), .Z(n14203) );
  NANDN U9683 ( .A(x[1828]), .B(y[1828]), .Z(n4886) );
  NANDN U9684 ( .A(x[1829]), .B(y[1829]), .Z(n4882) );
  AND U9685 ( .A(n4886), .B(n4882), .Z(n14211) );
  NANDN U9686 ( .A(y[1829]), .B(x[1829]), .Z(n4884) );
  NANDN U9687 ( .A(y[1830]), .B(x[1830]), .Z(n9835) );
  NAND U9688 ( .A(n4884), .B(n9835), .Z(n14212) );
  ANDN U9689 ( .B(x[1832]), .A(y[1832]), .Z(n4880) );
  NANDN U9690 ( .A(y[1833]), .B(x[1833]), .Z(n4881) );
  ANDN U9691 ( .B(x[1839]), .A(y[1839]), .Z(n14236) );
  NANDN U9692 ( .A(x[1841]), .B(y[1841]), .Z(n4871) );
  NANDN U9693 ( .A(y[1841]), .B(x[1841]), .Z(n4873) );
  ANDN U9694 ( .B(y[1843]), .A(x[1843]), .Z(n4867) );
  NANDN U9695 ( .A(y[1844]), .B(x[1844]), .Z(n14249) );
  IV U9696 ( .A(n14249), .Z(n9841) );
  NANDN U9697 ( .A(x[1844]), .B(y[1844]), .Z(n4868) );
  NANDN U9698 ( .A(y[1845]), .B(x[1845]), .Z(n9842) );
  NANDN U9699 ( .A(y[1846]), .B(x[1846]), .Z(n4866) );
  AND U9700 ( .A(n9842), .B(n4866), .Z(n14252) );
  IV U9701 ( .A(n14252), .Z(n4659) );
  ANDN U9702 ( .B(y[1846]), .A(x[1846]), .Z(n9843) );
  ANDN U9703 ( .B(y[1847]), .A(x[1847]), .Z(n9849) );
  NOR U9704 ( .A(n9843), .B(n9849), .Z(n14255) );
  NANDN U9705 ( .A(x[1850]), .B(y[1850]), .Z(n4861) );
  NANDN U9706 ( .A(x[1851]), .B(y[1851]), .Z(n9857) );
  AND U9707 ( .A(n4861), .B(n9857), .Z(n14262) );
  NANDN U9708 ( .A(y[1851]), .B(x[1851]), .Z(n4860) );
  ANDN U9709 ( .B(x[1852]), .A(y[1852]), .Z(n9863) );
  ANDN U9710 ( .B(n4860), .A(n9863), .Z(n14265) );
  NANDN U9711 ( .A(y[1854]), .B(x[1854]), .Z(n4661) );
  ANDN U9712 ( .B(x[1855]), .A(y[1855]), .Z(n4662) );
  ANDN U9713 ( .B(n4661), .A(n4662), .Z(n9868) );
  IV U9714 ( .A(n9868), .Z(n14275) );
  NANDN U9715 ( .A(x[1854]), .B(y[1854]), .Z(n4857) );
  NANDN U9716 ( .A(x[1855]), .B(y[1855]), .Z(n14274) );
  AND U9717 ( .A(n4857), .B(n14274), .Z(n14271) );
  ANDN U9718 ( .B(x[1856]), .A(y[1856]), .Z(n14272) );
  IV U9719 ( .A(n14272), .Z(n9874) );
  NANDN U9720 ( .A(x[1856]), .B(y[1856]), .Z(n9869) );
  NANDN U9721 ( .A(x[1857]), .B(y[1857]), .Z(n4856) );
  AND U9722 ( .A(n9869), .B(n4856), .Z(n14278) );
  ANDN U9723 ( .B(x[1857]), .A(y[1857]), .Z(n9873) );
  ANDN U9724 ( .B(x[1858]), .A(y[1858]), .Z(n9879) );
  NOR U9725 ( .A(n9873), .B(n9879), .Z(n14281) );
  NANDN U9726 ( .A(x[1863]), .B(y[1863]), .Z(n9887) );
  NANDN U9727 ( .A(y[1864]), .B(x[1864]), .Z(n4851) );
  ANDN U9728 ( .B(y[1865]), .A(x[1865]), .Z(n4849) );
  NANDN U9729 ( .A(y[1866]), .B(x[1866]), .Z(n14301) );
  IV U9730 ( .A(n14301), .Z(n9888) );
  NANDN U9731 ( .A(x[1866]), .B(y[1866]), .Z(n4850) );
  NANDN U9732 ( .A(y[1867]), .B(x[1867]), .Z(n9889) );
  ANDN U9733 ( .B(x[1868]), .A(y[1868]), .Z(n9893) );
  ANDN U9734 ( .B(n9889), .A(n9893), .Z(n14304) );
  NANDN U9735 ( .A(x[1869]), .B(y[1869]), .Z(n4847) );
  ANDN U9736 ( .B(y[1868]), .A(x[1868]), .Z(n9890) );
  ANDN U9737 ( .B(n4847), .A(n9890), .Z(n14307) );
  NANDN U9738 ( .A(y[1869]), .B(x[1869]), .Z(n9892) );
  NANDN U9739 ( .A(y[1870]), .B(x[1870]), .Z(n9897) );
  AND U9740 ( .A(n9892), .B(n9897), .Z(n14309) );
  IV U9741 ( .A(n14309), .Z(n4665) );
  ANDN U9742 ( .B(x[1876]), .A(y[1876]), .Z(n4842) );
  NANDN U9743 ( .A(x[1877]), .B(y[1877]), .Z(n14327) );
  NANDN U9744 ( .A(y[1877]), .B(x[1877]), .Z(n4841) );
  NANDN U9745 ( .A(x[1878]), .B(y[1878]), .Z(n4840) );
  NANDN U9746 ( .A(x[1879]), .B(y[1879]), .Z(n4838) );
  AND U9747 ( .A(n4840), .B(n4838), .Z(n14331) );
  ANDN U9748 ( .B(x[1879]), .A(y[1879]), .Z(n9918) );
  ANDN U9749 ( .B(x[1880]), .A(y[1880]), .Z(n9922) );
  NOR U9750 ( .A(n9918), .B(n9922), .Z(n14333) );
  ANDN U9751 ( .B(x[1881]), .A(y[1881]), .Z(n14336) );
  NANDN U9752 ( .A(y[1882]), .B(x[1882]), .Z(n4837) );
  NANDN U9753 ( .A(y[1883]), .B(x[1883]), .Z(n14341) );
  IV U9754 ( .A(n14341), .Z(n4836) );
  NANDN U9755 ( .A(y[1884]), .B(x[1884]), .Z(n9927) );
  ANDN U9756 ( .B(y[1885]), .A(x[1885]), .Z(n4834) );
  NANDN U9757 ( .A(y[1886]), .B(x[1886]), .Z(n4831) );
  ANDN U9758 ( .B(y[1887]), .A(x[1887]), .Z(n4829) );
  NANDN U9759 ( .A(y[1888]), .B(x[1888]), .Z(n14355) );
  NANDN U9760 ( .A(x[1888]), .B(y[1888]), .Z(n4830) );
  NANDN U9761 ( .A(y[1890]), .B(x[1890]), .Z(n9931) );
  ANDN U9762 ( .B(x[1889]), .A(y[1889]), .Z(n9928) );
  ANDN U9763 ( .B(n9931), .A(n9928), .Z(n14358) );
  NANDN U9764 ( .A(x[1890]), .B(y[1890]), .Z(n9929) );
  NANDN U9765 ( .A(x[1891]), .B(y[1891]), .Z(n9933) );
  AND U9766 ( .A(n9929), .B(n9933), .Z(n14361) );
  NANDN U9767 ( .A(x[1892]), .B(y[1892]), .Z(n9932) );
  NANDN U9768 ( .A(x[1893]), .B(y[1893]), .Z(n9939) );
  AND U9769 ( .A(n9932), .B(n9939), .Z(n14365) );
  NANDN U9770 ( .A(y[1893]), .B(x[1893]), .Z(n4827) );
  NANDN U9771 ( .A(y[1894]), .B(x[1894]), .Z(n4826) );
  NAND U9772 ( .A(n4827), .B(n4826), .Z(n14366) );
  NANDN U9773 ( .A(x[1894]), .B(y[1894]), .Z(n9938) );
  NANDN U9774 ( .A(x[1895]), .B(y[1895]), .Z(n9947) );
  AND U9775 ( .A(n9938), .B(n9947), .Z(n14368) );
  NANDN U9776 ( .A(y[1895]), .B(x[1895]), .Z(n4825) );
  ANDN U9777 ( .B(x[1896]), .A(y[1896]), .Z(n9950) );
  ANDN U9778 ( .B(n4825), .A(n9950), .Z(n14371) );
  NANDN U9779 ( .A(y[1898]), .B(x[1898]), .Z(n4822) );
  ANDN U9780 ( .B(x[1899]), .A(y[1899]), .Z(n4821) );
  NANDN U9781 ( .A(x[1900]), .B(y[1900]), .Z(n4668) );
  NANDN U9782 ( .A(x[1901]), .B(y[1901]), .Z(n9964) );
  AND U9783 ( .A(n4668), .B(n9964), .Z(n14384) );
  IV U9784 ( .A(n14384), .Z(n4669) );
  NANDN U9785 ( .A(y[1902]), .B(x[1902]), .Z(n9967) );
  ANDN U9786 ( .B(x[1901]), .A(y[1901]), .Z(n9960) );
  ANDN U9787 ( .B(n9967), .A(n9960), .Z(n14387) );
  NANDN U9788 ( .A(x[1903]), .B(y[1903]), .Z(n9968) );
  NANDN U9789 ( .A(x[1902]), .B(y[1902]), .Z(n4671) );
  AND U9790 ( .A(n9968), .B(n4671), .Z(n14389) );
  ANDN U9791 ( .B(y[1906]), .A(x[1906]), .Z(n14396) );
  ANDN U9792 ( .B(x[1908]), .A(y[1908]), .Z(n4819) );
  NANDN U9793 ( .A(x[1909]), .B(y[1909]), .Z(n4818) );
  NANDN U9794 ( .A(y[1910]), .B(x[1910]), .Z(n14407) );
  ANDN U9795 ( .B(y[1911]), .A(x[1911]), .Z(n14409) );
  NANDN U9796 ( .A(x[1910]), .B(y[1910]), .Z(n4817) );
  NANDN U9797 ( .A(x[1916]), .B(y[1916]), .Z(n4809) );
  ANDN U9798 ( .B(y[1917]), .A(x[1917]), .Z(n9994) );
  ANDN U9799 ( .B(n4809), .A(n9994), .Z(n14421) );
  NANDN U9800 ( .A(y[1917]), .B(x[1917]), .Z(n4807) );
  XOR U9801 ( .A(x[1918]), .B(y[1918]), .Z(n9992) );
  ANDN U9802 ( .B(n4807), .A(n9992), .Z(n14423) );
  NANDN U9803 ( .A(y[1919]), .B(x[1919]), .Z(n14427) );
  NANDN U9804 ( .A(x[1920]), .B(y[1920]), .Z(n4805) );
  NANDN U9805 ( .A(x[1926]), .B(y[1926]), .Z(n10012) );
  NANDN U9806 ( .A(x[1927]), .B(y[1927]), .Z(n10020) );
  AND U9807 ( .A(n10012), .B(n10020), .Z(n14445) );
  NANDN U9808 ( .A(x[1928]), .B(y[1928]), .Z(n14449) );
  ANDN U9809 ( .B(x[1930]), .A(y[1930]), .Z(n4794) );
  NANDN U9810 ( .A(x[1931]), .B(y[1931]), .Z(n4793) );
  ANDN U9811 ( .B(x[1932]), .A(y[1932]), .Z(n14459) );
  NANDN U9812 ( .A(x[1933]), .B(y[1933]), .Z(n14461) );
  NANDN U9813 ( .A(x[1932]), .B(y[1932]), .Z(n4792) );
  NANDN U9814 ( .A(x[1935]), .B(y[1935]), .Z(n10035) );
  ANDN U9815 ( .B(y[1934]), .A(x[1934]), .Z(n10030) );
  ANDN U9816 ( .B(n10035), .A(n10030), .Z(n14464) );
  IV U9817 ( .A(n14464), .Z(n4676) );
  NANDN U9818 ( .A(y[1935]), .B(x[1935]), .Z(n4791) );
  NANDN U9819 ( .A(y[1936]), .B(x[1936]), .Z(n4789) );
  NAND U9820 ( .A(n4791), .B(n4789), .Z(n14467) );
  NANDN U9821 ( .A(y[1939]), .B(x[1939]), .Z(n4785) );
  ANDN U9822 ( .B(x[1940]), .A(y[1940]), .Z(n10048) );
  ANDN U9823 ( .B(n4785), .A(n10048), .Z(n14474) );
  NANDN U9824 ( .A(y[1941]), .B(x[1941]), .Z(n14478) );
  ANDN U9825 ( .B(y[1942]), .A(x[1942]), .Z(n4782) );
  NANDN U9826 ( .A(x[1944]), .B(y[1944]), .Z(n4779) );
  NANDN U9827 ( .A(x[1945]), .B(y[1945]), .Z(n4777) );
  NAND U9828 ( .A(n4779), .B(n4777), .Z(n14488) );
  IV U9829 ( .A(n14488), .Z(n4679) );
  NANDN U9830 ( .A(x[1949]), .B(y[1949]), .Z(n10069) );
  NANDN U9831 ( .A(x[1948]), .B(y[1948]), .Z(n4680) );
  AND U9832 ( .A(n10069), .B(n4680), .Z(n14497) );
  ANDN U9833 ( .B(x[1949]), .A(y[1949]), .Z(n10064) );
  ANDN U9834 ( .B(x[1950]), .A(y[1950]), .Z(n10074) );
  NOR U9835 ( .A(n10064), .B(n10074), .Z(n14499) );
  NANDN U9836 ( .A(x[1952]), .B(y[1952]), .Z(n14504) );
  IV U9837 ( .A(n14504), .Z(n10075) );
  NANDN U9838 ( .A(x[1955]), .B(y[1955]), .Z(n10089) );
  ANDN U9839 ( .B(y[1954]), .A(x[1954]), .Z(n10086) );
  ANDN U9840 ( .B(n10089), .A(n10086), .Z(n14509) );
  NANDN U9841 ( .A(y[1955]), .B(x[1955]), .Z(n4681) );
  ANDN U9842 ( .B(x[1956]), .A(y[1956]), .Z(n10090) );
  ANDN U9843 ( .B(n4681), .A(n10090), .Z(n14515) );
  NANDN U9844 ( .A(x[1959]), .B(y[1959]), .Z(n4684) );
  ANDN U9845 ( .B(y[1958]), .A(x[1958]), .Z(n10097) );
  ANDN U9846 ( .B(n4684), .A(n10097), .Z(n14520) );
  IV U9847 ( .A(n14520), .Z(n4685) );
  NANDN U9848 ( .A(y[1960]), .B(x[1960]), .Z(n10103) );
  NANDN U9849 ( .A(y[1959]), .B(x[1959]), .Z(n4686) );
  AND U9850 ( .A(n10103), .B(n4686), .Z(n14523) );
  NANDN U9851 ( .A(x[1963]), .B(y[1963]), .Z(n4774) );
  NANDN U9852 ( .A(x[1962]), .B(y[1962]), .Z(n4687) );
  AND U9853 ( .A(n4774), .B(n4687), .Z(n14528) );
  NANDN U9854 ( .A(y[1963]), .B(x[1963]), .Z(n14531) );
  NANDN U9855 ( .A(y[1964]), .B(x[1964]), .Z(n10109) );
  NANDN U9856 ( .A(x[1964]), .B(y[1964]), .Z(n14532) );
  NANDN U9857 ( .A(x[1965]), .B(y[1965]), .Z(n14537) );
  ANDN U9858 ( .B(x[1967]), .A(y[1967]), .Z(n10116) );
  ANDN U9859 ( .B(x[1968]), .A(y[1968]), .Z(n10121) );
  NOR U9860 ( .A(n10116), .B(n10121), .Z(n14543) );
  NANDN U9861 ( .A(y[1969]), .B(x[1969]), .Z(n14546) );
  IV U9862 ( .A(n14546), .Z(n4688) );
  ANDN U9863 ( .B(y[1971]), .A(x[1971]), .Z(n4772) );
  NANDN U9864 ( .A(y[1972]), .B(x[1972]), .Z(n4771) );
  NANDN U9865 ( .A(y[1975]), .B(x[1975]), .Z(n4691) );
  NANDN U9866 ( .A(y[1974]), .B(x[1974]), .Z(n4690) );
  NAND U9867 ( .A(n4691), .B(n4690), .Z(n14559) );
  IV U9868 ( .A(n14559), .Z(n10126) );
  NANDN U9869 ( .A(x[1979]), .B(y[1979]), .Z(n10127) );
  NANDN U9870 ( .A(x[1978]), .B(y[1978]), .Z(n4767) );
  AND U9871 ( .A(n10127), .B(n4767), .Z(n14569) );
  NANDN U9872 ( .A(y[1979]), .B(x[1979]), .Z(n4766) );
  ANDN U9873 ( .B(x[1980]), .A(y[1980]), .Z(n10128) );
  ANDN U9874 ( .B(n4766), .A(n10128), .Z(n14571) );
  NANDN U9875 ( .A(x[1980]), .B(y[1980]), .Z(n4693) );
  NANDN U9876 ( .A(x[1981]), .B(y[1981]), .Z(n4692) );
  AND U9877 ( .A(n4693), .B(n4692), .Z(n14572) );
  IV U9878 ( .A(n14572), .Z(n10130) );
  NANDN U9879 ( .A(y[1982]), .B(x[1982]), .Z(n4696) );
  NANDN U9880 ( .A(y[1981]), .B(x[1981]), .Z(n4695) );
  NAND U9881 ( .A(n4696), .B(n4695), .Z(n14574) );
  IV U9882 ( .A(n14574), .Z(n10131) );
  NANDN U9883 ( .A(x[1982]), .B(y[1982]), .Z(n10132) );
  NANDN U9884 ( .A(x[1983]), .B(y[1983]), .Z(n4765) );
  AND U9885 ( .A(n10132), .B(n4765), .Z(n14576) );
  NANDN U9886 ( .A(y[1984]), .B(x[1984]), .Z(n10134) );
  ANDN U9887 ( .B(x[1983]), .A(y[1983]), .Z(n14578) );
  IV U9888 ( .A(n14578), .Z(n10133) );
  NANDN U9889 ( .A(x[1984]), .B(y[1984]), .Z(n14580) );
  NANDN U9890 ( .A(y[1989]), .B(x[1989]), .Z(n14595) );
  NANDN U9891 ( .A(y[1990]), .B(x[1990]), .Z(n4757) );
  NANDN U9892 ( .A(x[1991]), .B(y[1991]), .Z(n14601) );
  ANDN U9893 ( .B(x[1992]), .A(y[1992]), .Z(n14604) );
  IV U9894 ( .A(n14604), .Z(n10139) );
  NANDN U9895 ( .A(x[1992]), .B(y[1992]), .Z(n14600) );
  IV U9896 ( .A(n14600), .Z(n4697) );
  NANDN U9897 ( .A(x[1994]), .B(y[1994]), .Z(n4755) );
  NANDN U9898 ( .A(x[1995]), .B(y[1995]), .Z(n4752) );
  AND U9899 ( .A(n4755), .B(n4752), .Z(n14610) );
  NANDN U9900 ( .A(y[1995]), .B(x[1995]), .Z(n4753) );
  ANDN U9901 ( .B(x[1996]), .A(y[1996]), .Z(n10140) );
  ANDN U9902 ( .B(n4753), .A(n10140), .Z(n14613) );
  NANDN U9903 ( .A(x[1996]), .B(y[1996]), .Z(n14615) );
  IV U9904 ( .A(n14615), .Z(n4751) );
  NANDN U9905 ( .A(y[1998]), .B(x[1998]), .Z(n14621) );
  NANDN U9906 ( .A(y[1997]), .B(x[1997]), .Z(n14617) );
  NAND U9907 ( .A(n14621), .B(n14617), .Z(n4750) );
  NANDN U9908 ( .A(y[1999]), .B(x[1999]), .Z(n4749) );
  NANDN U9909 ( .A(n4749), .B(n4699), .Z(n4702) );
  NANDN U9910 ( .A(y[2001]), .B(x[2001]), .Z(n4701) );
  NANDN U9911 ( .A(y[2000]), .B(x[2000]), .Z(n4700) );
  NAND U9912 ( .A(n4701), .B(n4700), .Z(n10141) );
  ANDN U9913 ( .B(n4702), .A(n10141), .Z(n14625) );
  NANDN U9914 ( .A(x[2003]), .B(y[2003]), .Z(n14630) );
  IV U9915 ( .A(n14630), .Z(n10146) );
  NANDN U9916 ( .A(y[2004]), .B(x[2004]), .Z(n4703) );
  NAND U9917 ( .A(n4704), .B(n4703), .Z(n14632) );
  IV U9918 ( .A(n14632), .Z(n4705) );
  NANDN U9919 ( .A(x[2007]), .B(y[2007]), .Z(n4708) );
  NANDN U9920 ( .A(x[2008]), .B(y[2008]), .Z(n4707) );
  AND U9921 ( .A(n4708), .B(n4707), .Z(n14639) );
  NANDN U9922 ( .A(y[2009]), .B(x[2009]), .Z(n4710) );
  NANDN U9923 ( .A(y[2008]), .B(x[2008]), .Z(n4709) );
  NAND U9924 ( .A(n4710), .B(n4709), .Z(n14641) );
  ANDN U9925 ( .B(y[2009]), .A(x[2009]), .Z(n14643) );
  NANDN U9926 ( .A(x[2011]), .B(y[2011]), .Z(n4746) );
  ANDN U9927 ( .B(y[2010]), .A(x[2010]), .Z(n10150) );
  ANDN U9928 ( .B(n4746), .A(n10150), .Z(n14647) );
  ANDN U9929 ( .B(y[2013]), .A(x[2013]), .Z(n10170) );
  NANDN U9930 ( .A(x[2012]), .B(y[2012]), .Z(n4747) );
  NANDN U9931 ( .A(n10170), .B(n4747), .Z(n14651) );
  ANDN U9932 ( .B(x[2014]), .A(y[2014]), .Z(n10172) );
  NANDN U9933 ( .A(x[2015]), .B(y[2015]), .Z(n10154) );
  ANDN U9934 ( .B(y[2014]), .A(x[2014]), .Z(n10153) );
  ANDN U9935 ( .B(n10154), .A(n10153), .Z(n14654) );
  ANDN U9936 ( .B(x[2015]), .A(y[2015]), .Z(n4743) );
  ANDN U9937 ( .B(x[2016]), .A(y[2016]), .Z(n10156) );
  NOR U9938 ( .A(n4743), .B(n10156), .Z(n14657) );
  NANDN U9939 ( .A(x[2018]), .B(y[2018]), .Z(n14662) );
  IV U9940 ( .A(n14662), .Z(n4741) );
  ANDN U9941 ( .B(x[2019]), .A(y[2019]), .Z(n14665) );
  XNOR U9942 ( .A(y[2022]), .B(x[2022]), .Z(n10161) );
  ANDN U9943 ( .B(x[2021]), .A(y[2021]), .Z(n10159) );
  ANDN U9944 ( .B(n10161), .A(n10159), .Z(n14673) );
  NANDN U9945 ( .A(x[2022]), .B(y[2022]), .Z(n14675) );
  NANDN U9946 ( .A(x[2023]), .B(y[2023]), .Z(n4736) );
  ANDN U9947 ( .B(x[2024]), .A(y[2024]), .Z(n4735) );
  NANDN U9948 ( .A(x[2025]), .B(y[2025]), .Z(n4733) );
  NANDN U9949 ( .A(y[2026]), .B(x[2026]), .Z(n4730) );
  NANDN U9950 ( .A(y[2025]), .B(x[2025]), .Z(n4734) );
  AND U9951 ( .A(n4730), .B(n4734), .Z(n4712) );
  NANDN U9952 ( .A(y[2027]), .B(x[2027]), .Z(n4731) );
  ANDN U9953 ( .B(y[2029]), .A(x[2029]), .Z(n4727) );
  NANDN U9954 ( .A(y[2029]), .B(x[2029]), .Z(n10163) );
  NANDN U9955 ( .A(y[2033]), .B(x[2033]), .Z(n4715) );
  NANDN U9956 ( .A(y[2032]), .B(x[2032]), .Z(n4714) );
  NAND U9957 ( .A(n4715), .B(n4714), .Z(n14691) );
  NANDN U9958 ( .A(x[2033]), .B(y[2033]), .Z(n4717) );
  NANDN U9959 ( .A(x[2034]), .B(y[2034]), .Z(n4716) );
  AND U9960 ( .A(n4717), .B(n4716), .Z(n14692) );
  IV U9961 ( .A(n14692), .Z(n10165) );
  NANDN U9962 ( .A(y[2035]), .B(x[2035]), .Z(n4719) );
  NANDN U9963 ( .A(y[2034]), .B(x[2034]), .Z(n4718) );
  AND U9964 ( .A(n4719), .B(n4718), .Z(n14693) );
  NANDN U9965 ( .A(y[2037]), .B(x[2037]), .Z(n4723) );
  ANDN U9966 ( .B(n4723), .A(n4722), .Z(n14695) );
  AND U9967 ( .A(n4725), .B(n4724), .Z(n14689) );
  NANDN U9968 ( .A(n4727), .B(n4726), .Z(n14688) );
  ANDN U9969 ( .B(n4729), .A(n4728), .Z(n14686) );
  NAND U9970 ( .A(n4731), .B(n4730), .Z(n14685) );
  ANDN U9971 ( .B(n4733), .A(n4732), .Z(n14683) );
  NANDN U9972 ( .A(n4735), .B(n4734), .Z(n14681) );
  AND U9973 ( .A(n4737), .B(n4736), .Z(n14678) );
  AND U9974 ( .A(n4739), .B(n4738), .Z(n14667) );
  NANDN U9975 ( .A(n14665), .B(n4740), .Z(n10158) );
  ANDN U9976 ( .B(n4745), .A(n4744), .Z(n10171) );
  ANDN U9977 ( .B(n4757), .A(n4756), .Z(n14599) );
  NAND U9978 ( .A(n14599), .B(n4758), .Z(n10138) );
  NANDN U9979 ( .A(x[1973]), .B(y[1973]), .Z(n4768) );
  AND U9980 ( .A(n4769), .B(n4768), .Z(n14557) );
  NAND U9981 ( .A(n4771), .B(n4770), .Z(n14555) );
  ANDN U9982 ( .B(n4773), .A(n4772), .Z(n14552) );
  AND U9983 ( .A(n14532), .B(n4774), .Z(n10108) );
  AND U9984 ( .A(n14515), .B(n14510), .Z(n10088) );
  NAND U9985 ( .A(n4776), .B(n4775), .Z(n10060) );
  AND U9986 ( .A(n4778), .B(n4777), .Z(n10058) );
  ANDN U9987 ( .B(n4779), .A(n14484), .Z(n10053) );
  NAND U9988 ( .A(n4781), .B(n4780), .Z(n14482) );
  ANDN U9989 ( .B(n4783), .A(n4782), .Z(n14481) );
  AND U9990 ( .A(n4785), .B(n4784), .Z(n10043) );
  NAND U9991 ( .A(n4787), .B(n4786), .Z(n10041) );
  AND U9992 ( .A(n4789), .B(n4788), .Z(n10039) );
  AND U9993 ( .A(n4791), .B(n4790), .Z(n10033) );
  NAND U9994 ( .A(n4793), .B(n4792), .Z(n14457) );
  ANDN U9995 ( .B(n4795), .A(n4794), .Z(n14455) );
  NAND U9996 ( .A(n4797), .B(n4796), .Z(n14453) );
  AND U9997 ( .A(n4799), .B(n4798), .Z(n14451) );
  NOR U9998 ( .A(n4801), .B(n4800), .Z(n10010) );
  AND U9999 ( .A(n14435), .B(n4802), .Z(n10004) );
  AND U10000 ( .A(n4804), .B(n4803), .Z(n14431) );
  NANDN U10001 ( .A(n4806), .B(n4805), .Z(n14428) );
  AND U10002 ( .A(n4808), .B(n4807), .Z(n9990) );
  NAND U10003 ( .A(n4810), .B(n4809), .Z(n9988) );
  AND U10004 ( .A(n4812), .B(n4811), .Z(n9986) );
  NAND U10005 ( .A(n4814), .B(n4813), .Z(n9984) );
  AND U10006 ( .A(n4816), .B(n4815), .Z(n9982) );
  NAND U10007 ( .A(n4818), .B(n4817), .Z(n14405) );
  NOR U10008 ( .A(n4820), .B(n4819), .Z(n14402) );
  XNOR U10009 ( .A(x[1902]), .B(y[1902]), .Z(n9966) );
  ANDN U10010 ( .B(x[1900]), .A(y[1900]), .Z(n9962) );
  ANDN U10011 ( .B(n4822), .A(n4821), .Z(n14381) );
  AND U10012 ( .A(n4824), .B(n4823), .Z(n9953) );
  AND U10013 ( .A(n4826), .B(n4825), .Z(n9943) );
  AND U10014 ( .A(n4828), .B(n4827), .Z(n9937) );
  ANDN U10015 ( .B(n4830), .A(n4829), .Z(n14353) );
  NAND U10016 ( .A(n4832), .B(n4831), .Z(n14351) );
  NOR U10017 ( .A(n4834), .B(n4833), .Z(n14349) );
  ANDN U10018 ( .B(n4837), .A(n4836), .Z(n14339) );
  AND U10019 ( .A(n4839), .B(n4838), .Z(n9921) );
  AND U10020 ( .A(n14327), .B(n4840), .Z(n9916) );
  NANDN U10021 ( .A(n4842), .B(n4841), .Z(n14325) );
  AND U10022 ( .A(n4844), .B(n4843), .Z(n14323) );
  AND U10023 ( .A(n4846), .B(n4845), .Z(n9901) );
  AND U10024 ( .A(n4848), .B(n4847), .Z(n9895) );
  ANDN U10025 ( .B(n4850), .A(n4849), .Z(n14299) );
  AND U10026 ( .A(n4852), .B(n4851), .Z(n14296) );
  AND U10027 ( .A(n4856), .B(n4855), .Z(n9877) );
  AND U10028 ( .A(n4858), .B(n4857), .Z(n9866) );
  AND U10029 ( .A(n4860), .B(n4859), .Z(n9856) );
  NAND U10030 ( .A(n4862), .B(n4861), .Z(n9854) );
  AND U10031 ( .A(n4864), .B(n4863), .Z(n9852) );
  AND U10032 ( .A(n4866), .B(n4865), .Z(n9846) );
  ANDN U10033 ( .B(n4868), .A(n4867), .Z(n14246) );
  AND U10034 ( .A(n4870), .B(n4869), .Z(n14245) );
  NANDN U10035 ( .A(n4872), .B(n4871), .Z(n14243) );
  AND U10036 ( .A(n4874), .B(n4873), .Z(n14241) );
  AND U10037 ( .A(n4878), .B(n4877), .Z(n9838) );
  ANDN U10038 ( .B(n4881), .A(n4880), .Z(n14221) );
  AND U10039 ( .A(n4889), .B(n4888), .Z(n9832) );
  ANDN U10040 ( .B(n4891), .A(n4890), .Z(n14195) );
  ANDN U10041 ( .B(n4893), .A(n4892), .Z(n14192) );
  AND U10042 ( .A(n4897), .B(n4896), .Z(n9814) );
  ANDN U10043 ( .B(n4899), .A(n4898), .Z(n9808) );
  AND U10044 ( .A(n4901), .B(n4900), .Z(n14167) );
  NANDN U10045 ( .A(n4903), .B(n4902), .Z(n9779) );
  AND U10046 ( .A(n10177), .B(n4904), .Z(n9777) );
  ANDN U10047 ( .B(x[1794]), .A(y[1794]), .Z(n9771) );
  OR U10048 ( .A(n4906), .B(n4905), .Z(n4907) );
  AND U10049 ( .A(n4908), .B(n4907), .Z(n9763) );
  NAND U10050 ( .A(n4911), .B(n4910), .Z(n14121) );
  NOR U10051 ( .A(n4913), .B(n4912), .Z(n14118) );
  NAND U10052 ( .A(n4918), .B(n4917), .Z(n14095) );
  ANDN U10053 ( .B(n4920), .A(n4919), .Z(n14093) );
  NAND U10054 ( .A(n4922), .B(n4921), .Z(n14091) );
  AND U10055 ( .A(n4924), .B(n4923), .Z(n14089) );
  ANDN U10056 ( .B(n4925), .A(n10178), .Z(n9722) );
  ANDN U10057 ( .B(n4927), .A(n4926), .Z(n9717) );
  XNOR U10058 ( .A(x[1764]), .B(y[1764]), .Z(n9711) );
  AND U10059 ( .A(n4929), .B(n4928), .Z(n9707) );
  AND U10060 ( .A(n4931), .B(n4930), .Z(n9705) );
  NAND U10061 ( .A(n4933), .B(n4932), .Z(n9703) );
  AND U10062 ( .A(n4935), .B(n4934), .Z(n9701) );
  NANDN U10063 ( .A(n4937), .B(n4936), .Z(n14046) );
  AND U10064 ( .A(n4939), .B(n4938), .Z(n14045) );
  NANDN U10065 ( .A(n4941), .B(n4940), .Z(n14043) );
  NANDN U10066 ( .A(n4956), .B(n4955), .Z(n13995) );
  AND U10067 ( .A(n4958), .B(n4957), .Z(n13993) );
  NANDN U10068 ( .A(n4960), .B(n4959), .Z(n13991) );
  AND U10069 ( .A(n4962), .B(n4961), .Z(n13989) );
  IV U10070 ( .A(n13971), .Z(n4969) );
  NAND U10071 ( .A(n4980), .B(n4979), .Z(n13942) );
  IV U10072 ( .A(n13942), .Z(n9651) );
  ANDN U10073 ( .B(n4982), .A(n4981), .Z(n13941) );
  AND U10074 ( .A(n4993), .B(n4992), .Z(n13889) );
  AND U10075 ( .A(n4995), .B(n4994), .Z(n13869) );
  NANDN U10076 ( .A(n4997), .B(n4996), .Z(n13867) );
  AND U10077 ( .A(n13855), .B(n4998), .Z(n9610) );
  NAND U10078 ( .A(n5000), .B(n4999), .Z(n9608) );
  ANDN U10079 ( .B(n5001), .A(n13847), .Z(n9606) );
  ANDN U10080 ( .B(n5003), .A(n5002), .Z(n13843) );
  NAND U10081 ( .A(n5005), .B(n5004), .Z(n13841) );
  ANDN U10082 ( .B(n5007), .A(n5006), .Z(n13839) );
  NAND U10083 ( .A(n5009), .B(n5008), .Z(n13837) );
  ANDN U10084 ( .B(n5010), .A(n13835), .Z(n9597) );
  NANDN U10085 ( .A(y[1660]), .B(x[1660]), .Z(n9588) );
  AND U10086 ( .A(n13821), .B(n5011), .Z(n9580) );
  AND U10087 ( .A(n5013), .B(n5012), .Z(n13817) );
  NANDN U10088 ( .A(n5015), .B(n5014), .Z(n13815) );
  NAND U10089 ( .A(n5017), .B(n5016), .Z(n9570) );
  AND U10090 ( .A(n5025), .B(n5024), .Z(n13795) );
  ANDN U10091 ( .B(n5027), .A(n5026), .Z(n13779) );
  NANDN U10092 ( .A(n5029), .B(n5028), .Z(n13777) );
  ANDN U10093 ( .B(n5031), .A(n5030), .Z(n13775) );
  AND U10094 ( .A(n5033), .B(n5032), .Z(n13773) );
  NANDN U10095 ( .A(y[1634]), .B(x[1634]), .Z(n5034) );
  AND U10096 ( .A(n5035), .B(n5034), .Z(n13763) );
  NANDN U10097 ( .A(n5037), .B(n5036), .Z(n13761) );
  NAND U10098 ( .A(n5039), .B(n5038), .Z(n13759) );
  NOR U10099 ( .A(n5041), .B(n5040), .Z(n13756) );
  NAND U10100 ( .A(n5044), .B(n5043), .Z(n13742) );
  NOR U10101 ( .A(n5046), .B(n5045), .Z(n13741) );
  NAND U10102 ( .A(n5048), .B(n5047), .Z(n13739) );
  NAND U10103 ( .A(n5053), .B(n5052), .Z(n13716) );
  NAND U10104 ( .A(n5057), .B(n5056), .Z(n13705) );
  ANDN U10105 ( .B(n5059), .A(n5058), .Z(n13702) );
  NAND U10106 ( .A(n5061), .B(n5060), .Z(n13697) );
  NAND U10107 ( .A(n5064), .B(n5063), .Z(n13685) );
  AND U10108 ( .A(n13668), .B(n5067), .Z(n13665) );
  ANDN U10109 ( .B(n5070), .A(n5069), .Z(n13659) );
  NAND U10110 ( .A(n5072), .B(n5071), .Z(n13657) );
  ANDN U10111 ( .B(n5074), .A(n5073), .Z(n13655) );
  NAND U10112 ( .A(n5076), .B(n5075), .Z(n13653) );
  IV U10113 ( .A(n13612), .Z(n5078) );
  NANDN U10114 ( .A(n5081), .B(n5080), .Z(n5082) );
  AND U10115 ( .A(n5083), .B(n5082), .Z(n13607) );
  NAND U10116 ( .A(n5086), .B(n5085), .Z(n13595) );
  OR U10117 ( .A(n5088), .B(n5087), .Z(n5089) );
  AND U10118 ( .A(n5090), .B(n5089), .Z(n13587) );
  NANDN U10119 ( .A(n5092), .B(n13578), .Z(n9516) );
  NAND U10120 ( .A(n5094), .B(n5093), .Z(n5095) );
  NANDN U10121 ( .A(n5096), .B(n5095), .Z(n13577) );
  AND U10122 ( .A(n5097), .B(n13575), .Z(n9511) );
  AND U10123 ( .A(n5099), .B(n5098), .Z(n9506) );
  NAND U10124 ( .A(n5101), .B(n5100), .Z(n9496) );
  AND U10125 ( .A(n5103), .B(n5102), .Z(n9494) );
  NANDN U10126 ( .A(n5105), .B(n5104), .Z(n9492) );
  ANDN U10127 ( .B(n5106), .A(n13555), .Z(n9490) );
  ANDN U10128 ( .B(n5108), .A(n5107), .Z(n13553) );
  NAND U10129 ( .A(n5110), .B(n5109), .Z(n13551) );
  NOR U10130 ( .A(n5112), .B(n5111), .Z(n13548) );
  ANDN U10131 ( .B(n5118), .A(n5117), .Z(n13529) );
  ANDN U10132 ( .B(n5120), .A(n5119), .Z(n13527) );
  ANDN U10133 ( .B(n5122), .A(n5121), .Z(n13525) );
  NANDN U10134 ( .A(n5127), .B(n5126), .Z(n13513) );
  NANDN U10135 ( .A(n5130), .B(n5129), .Z(n13501) );
  ANDN U10136 ( .B(n5132), .A(n5131), .Z(n13499) );
  NANDN U10137 ( .A(n5134), .B(n5133), .Z(n13497) );
  ANDN U10138 ( .B(n5135), .A(n13495), .Z(n9480) );
  ANDN U10139 ( .B(n5142), .A(n5141), .Z(n13477) );
  ANDN U10140 ( .B(n5146), .A(n5145), .Z(n13468) );
  ANDN U10141 ( .B(n5150), .A(n5149), .Z(n13455) );
  NANDN U10142 ( .A(y[1500]), .B(x[1500]), .Z(n5152) );
  NAND U10143 ( .A(n5153), .B(n5152), .Z(n13445) );
  NAND U10144 ( .A(n5158), .B(n5157), .Z(n13433) );
  ANDN U10145 ( .B(n5164), .A(n5163), .Z(n13401) );
  OR U10146 ( .A(n5166), .B(n5165), .Z(n5167) );
  AND U10147 ( .A(n5168), .B(n5167), .Z(n13393) );
  NAND U10148 ( .A(n5171), .B(n5170), .Z(n13376) );
  OR U10149 ( .A(n5173), .B(n5172), .Z(n5174) );
  AND U10150 ( .A(n5175), .B(n5174), .Z(n13369) );
  ANDN U10151 ( .B(n5181), .A(n5180), .Z(n13347) );
  NANDN U10152 ( .A(n5183), .B(n5182), .Z(n13345) );
  ANDN U10153 ( .B(n5185), .A(n5184), .Z(n13343) );
  NANDN U10154 ( .A(n5187), .B(n5186), .Z(n13341) );
  ANDN U10155 ( .B(n5189), .A(n5188), .Z(n13339) );
  NANDN U10156 ( .A(n5191), .B(n5190), .Z(n13337) );
  ANDN U10157 ( .B(n13321), .A(n5193), .Z(n9426) );
  NAND U10158 ( .A(n5195), .B(n5194), .Z(n13319) );
  NANDN U10159 ( .A(n5198), .B(n5197), .Z(n5199) );
  AND U10160 ( .A(n5200), .B(n5199), .Z(n13291) );
  NAND U10161 ( .A(n5209), .B(n5208), .Z(n13271) );
  NOR U10162 ( .A(n5211), .B(n5210), .Z(n13268) );
  NAND U10163 ( .A(n5213), .B(n5212), .Z(n13266) );
  IV U10164 ( .A(n13266), .Z(n9412) );
  NAND U10165 ( .A(n5215), .B(n5214), .Z(n5217) );
  ANDN U10166 ( .B(n5217), .A(n5216), .Z(n13264) );
  ANDN U10167 ( .B(n5223), .A(n5222), .Z(n13219) );
  ANDN U10168 ( .B(n5227), .A(n5226), .Z(n13199) );
  AND U10169 ( .A(n5229), .B(n5228), .Z(n13187) );
  NANDN U10170 ( .A(n5231), .B(n5230), .Z(n13185) );
  AND U10171 ( .A(n5233), .B(n5232), .Z(n13182) );
  NANDN U10172 ( .A(y[1380]), .B(x[1380]), .Z(n5235) );
  AND U10173 ( .A(n5236), .B(n5235), .Z(n13167) );
  NAND U10174 ( .A(n5238), .B(n5237), .Z(n13165) );
  NANDN U10175 ( .A(n5240), .B(n5239), .Z(n13163) );
  NANDN U10176 ( .A(n5242), .B(n5241), .Z(n5243) );
  AND U10177 ( .A(n5244), .B(n5243), .Z(n13155) );
  NANDN U10178 ( .A(n5245), .B(n13146), .Z(n9366) );
  ANDN U10179 ( .B(n5247), .A(n5246), .Z(n13141) );
  NAND U10180 ( .A(n5249), .B(n5248), .Z(n13139) );
  ANDN U10181 ( .B(n5251), .A(n5250), .Z(n13121) );
  NANDN U10182 ( .A(y[1350]), .B(x[1350]), .Z(n5254) );
  AND U10183 ( .A(n5255), .B(n5254), .Z(n13093) );
  ANDN U10184 ( .B(n5257), .A(n5256), .Z(n13090) );
  NAND U10185 ( .A(n5259), .B(n5258), .Z(n13088) );
  NOR U10186 ( .A(n5261), .B(n5260), .Z(n13087) );
  NAND U10187 ( .A(n5263), .B(n5262), .Z(n13085) );
  ANDN U10188 ( .B(n5264), .A(n13083), .Z(n9343) );
  NAND U10189 ( .A(n5266), .B(n5265), .Z(n13073) );
  ANDN U10190 ( .B(n5268), .A(n5267), .Z(n13071) );
  NAND U10191 ( .A(n5270), .B(n5269), .Z(n13069) );
  XNOR U10192 ( .A(y[1333]), .B(x[1333]), .Z(n9322) );
  NAND U10193 ( .A(n5272), .B(n5271), .Z(n13037) );
  ANDN U10194 ( .B(n5275), .A(n5274), .Z(n13025) );
  AND U10195 ( .A(n5277), .B(n5276), .Z(n13023) );
  NANDN U10196 ( .A(n5279), .B(n5278), .Z(n13021) );
  AND U10197 ( .A(n5281), .B(n5280), .Z(n13019) );
  NANDN U10198 ( .A(n5283), .B(n5282), .Z(n13017) );
  ANDN U10199 ( .B(n5287), .A(n5286), .Z(n13005) );
  NAND U10200 ( .A(n5289), .B(n5288), .Z(n13003) );
  ANDN U10201 ( .B(n5291), .A(n5290), .Z(n13001) );
  NAND U10202 ( .A(n5293), .B(n5292), .Z(n12988) );
  IV U10203 ( .A(n12988), .Z(n9303) );
  NAND U10204 ( .A(n5296), .B(n5295), .Z(n5297) );
  NAND U10205 ( .A(n5298), .B(n5297), .Z(n5299) );
  NAND U10206 ( .A(n5300), .B(n5299), .Z(n12964) );
  ANDN U10207 ( .B(n5304), .A(n5303), .Z(n12941) );
  NANDN U10208 ( .A(n5306), .B(n5305), .Z(n12939) );
  ANDN U10209 ( .B(n5308), .A(n5307), .Z(n12937) );
  NOR U10210 ( .A(n5310), .B(n5309), .Z(n12935) );
  NAND U10211 ( .A(n5312), .B(n5311), .Z(n12933) );
  ANDN U10212 ( .B(n5314), .A(n5313), .Z(n12931) );
  NANDN U10213 ( .A(y[1278]), .B(x[1278]), .Z(n5316) );
  NAND U10214 ( .A(n5316), .B(n5315), .Z(n12929) );
  NAND U10215 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U10216 ( .A(n5320), .B(n5319), .Z(n5321) );
  NAND U10217 ( .A(n5322), .B(n5321), .Z(n12917) );
  ANDN U10218 ( .B(n5325), .A(n5324), .Z(n12899) );
  NANDN U10219 ( .A(n5327), .B(n5326), .Z(n12897) );
  ANDN U10220 ( .B(n5329), .A(n5328), .Z(n12895) );
  NANDN U10221 ( .A(n5331), .B(n5330), .Z(n12893) );
  NAND U10222 ( .A(n5334), .B(n5333), .Z(n12881) );
  ANDN U10223 ( .B(n5337), .A(n5336), .Z(n12867) );
  NAND U10224 ( .A(n5339), .B(n5338), .Z(n12865) );
  NAND U10225 ( .A(n5341), .B(n5340), .Z(n12852) );
  NAND U10226 ( .A(n5343), .B(n5342), .Z(n12840) );
  NAND U10227 ( .A(n5345), .B(n5344), .Z(n12829) );
  NAND U10228 ( .A(n5347), .B(n5346), .Z(n12792) );
  NAND U10229 ( .A(n5349), .B(n5348), .Z(n12777) );
  ANDN U10230 ( .B(n5351), .A(n5350), .Z(n12761) );
  ANDN U10231 ( .B(n5353), .A(n5352), .Z(n12757) );
  NAND U10232 ( .A(n5355), .B(n5354), .Z(n12739) );
  ANDN U10233 ( .B(n5357), .A(n5356), .Z(n12737) );
  AND U10234 ( .A(n5359), .B(n5358), .Z(n12734) );
  NANDN U10235 ( .A(n12732), .B(n5360), .Z(n9211) );
  ANDN U10236 ( .B(n5362), .A(n5361), .Z(n12725) );
  OR U10237 ( .A(n5365), .B(n5364), .Z(n5366) );
  AND U10238 ( .A(n5367), .B(n5366), .Z(n12716) );
  AND U10239 ( .A(n5369), .B(n5368), .Z(n12715) );
  ANDN U10240 ( .B(n5371), .A(n5370), .Z(n12713) );
  ANDN U10241 ( .B(n5373), .A(n5372), .Z(n12711) );
  ANDN U10242 ( .B(n5375), .A(n5374), .Z(n12707) );
  NAND U10243 ( .A(n5377), .B(n5376), .Z(n12705) );
  NAND U10244 ( .A(n5379), .B(n5378), .Z(n12690) );
  NANDN U10245 ( .A(n5381), .B(n5380), .Z(n12689) );
  NAND U10246 ( .A(n5384), .B(n5383), .Z(n12677) );
  NAND U10247 ( .A(n5391), .B(n5390), .Z(n12653) );
  NAND U10248 ( .A(n12649), .B(n12645), .Z(n9187) );
  NAND U10249 ( .A(n5396), .B(n5395), .Z(n12637) );
  NAND U10250 ( .A(n5398), .B(n5397), .Z(n12624) );
  AND U10251 ( .A(n5400), .B(n5399), .Z(n12623) );
  NANDN U10252 ( .A(n5402), .B(n5401), .Z(n12621) );
  ANDN U10253 ( .B(n5405), .A(n5404), .Z(n12607) );
  NOR U10254 ( .A(n5407), .B(n5406), .Z(n12605) );
  ANDN U10255 ( .B(n5409), .A(n5408), .Z(n12577) );
  NAND U10256 ( .A(n5411), .B(n5410), .Z(n12560) );
  AND U10257 ( .A(n5413), .B(n5412), .Z(n12549) );
  NANDN U10258 ( .A(n5415), .B(n5414), .Z(n12547) );
  AND U10259 ( .A(n5417), .B(n5416), .Z(n12545) );
  ANDN U10260 ( .B(n5419), .A(n5418), .Z(n12533) );
  ANDN U10261 ( .B(n5422), .A(n5421), .Z(n12521) );
  ANDN U10262 ( .B(n5426), .A(n5425), .Z(n12509) );
  ANDN U10263 ( .B(x[1110]), .A(y[1110]), .Z(n9136) );
  NAND U10264 ( .A(n5428), .B(n5427), .Z(n12489) );
  IV U10265 ( .A(n12479), .Z(n5429) );
  NAND U10266 ( .A(n5438), .B(n5437), .Z(n12452) );
  IV U10267 ( .A(n12450), .Z(n5439) );
  NAND U10268 ( .A(n5442), .B(n5441), .Z(n12430) );
  NANDN U10269 ( .A(n5445), .B(n5444), .Z(n12404) );
  AND U10270 ( .A(n5447), .B(n5446), .Z(n12403) );
  NANDN U10271 ( .A(n5449), .B(n5448), .Z(n12401) );
  AND U10272 ( .A(n5451), .B(n5450), .Z(n12398) );
  ANDN U10273 ( .B(n5454), .A(n12388), .Z(n9096) );
  NAND U10274 ( .A(n5456), .B(n5455), .Z(n12386) );
  NAND U10275 ( .A(n5462), .B(n5457), .Z(n5459) );
  ANDN U10276 ( .B(n5459), .A(n5458), .Z(n12385) );
  NAND U10277 ( .A(n5461), .B(n5460), .Z(n5463) );
  AND U10278 ( .A(n5463), .B(n5462), .Z(n5464) );
  NAND U10279 ( .A(n5465), .B(n5464), .Z(n12383) );
  NANDN U10280 ( .A(n5467), .B(n5466), .Z(n12379) );
  NANDN U10281 ( .A(n5469), .B(n5468), .Z(n12370) );
  AND U10282 ( .A(n5471), .B(n5470), .Z(n12369) );
  NANDN U10283 ( .A(n5473), .B(n5472), .Z(n12367) );
  ANDN U10284 ( .B(n5475), .A(n5474), .Z(n12365) );
  NAND U10285 ( .A(n5477), .B(n5476), .Z(n12363) );
  ANDN U10286 ( .B(n5478), .A(n12361), .Z(n9078) );
  NANDN U10287 ( .A(n5480), .B(n5479), .Z(n12351) );
  AND U10288 ( .A(n12349), .B(n5481), .Z(n9070) );
  AND U10289 ( .A(n5483), .B(n5482), .Z(n12327) );
  ANDN U10290 ( .B(n5485), .A(n5484), .Z(n12325) );
  AND U10291 ( .A(n5487), .B(n5486), .Z(n12322) );
  ANDN U10292 ( .B(n5489), .A(n5488), .Z(n12321) );
  NAND U10293 ( .A(n5491), .B(n5490), .Z(n12319) );
  NAND U10294 ( .A(n5493), .B(n5492), .Z(n12307) );
  ANDN U10295 ( .B(n5495), .A(n5494), .Z(n12305) );
  NAND U10296 ( .A(n5497), .B(n5496), .Z(n12303) );
  ANDN U10297 ( .B(n5499), .A(n5498), .Z(n12301) );
  NAND U10298 ( .A(n5501), .B(n5500), .Z(n12299) );
  NANDN U10299 ( .A(n5504), .B(n5503), .Z(n12259) );
  ANDN U10300 ( .B(n5508), .A(n5507), .Z(n12235) );
  AND U10301 ( .A(n5510), .B(n5509), .Z(n12232) );
  NANDN U10302 ( .A(n5514), .B(n5513), .Z(n12219) );
  NAND U10303 ( .A(n12213), .B(n5515), .Z(n12211) );
  ANDN U10304 ( .B(n5517), .A(n5516), .Z(n12207) );
  ANDN U10305 ( .B(n5519), .A(n5518), .Z(n12205) );
  ANDN U10306 ( .B(n5521), .A(n5520), .Z(n12199) );
  ANDN U10307 ( .B(n5523), .A(n5522), .Z(n12179) );
  AND U10308 ( .A(n5525), .B(n5524), .Z(n8956) );
  AND U10309 ( .A(n5527), .B(n5526), .Z(n12143) );
  NANDN U10310 ( .A(n5529), .B(n5528), .Z(n12141) );
  AND U10311 ( .A(n5531), .B(n5530), .Z(n12139) );
  AND U10312 ( .A(n5536), .B(n5535), .Z(n12095) );
  NANDN U10313 ( .A(n5538), .B(n5537), .Z(n12093) );
  ANDN U10314 ( .B(n5540), .A(n5539), .Z(n12091) );
  ANDN U10315 ( .B(n5543), .A(n5542), .Z(n12071) );
  ANDN U10316 ( .B(n5545), .A(n5544), .Z(n12068) );
  AND U10317 ( .A(n5549), .B(n5548), .Z(n12055) );
  OR U10318 ( .A(n5552), .B(n5551), .Z(n5553) );
  AND U10319 ( .A(n5554), .B(n5553), .Z(n8874) );
  NANDN U10320 ( .A(n5557), .B(n5556), .Z(n12035) );
  ANDN U10321 ( .B(n5559), .A(n5558), .Z(n12033) );
  NAND U10322 ( .A(n5561), .B(n5560), .Z(n12026) );
  NOR U10323 ( .A(n5563), .B(n5562), .Z(n8863) );
  NANDN U10324 ( .A(y[902]), .B(x[902]), .Z(n8857) );
  NANDN U10325 ( .A(n5565), .B(n5564), .Z(n12001) );
  AND U10326 ( .A(n5567), .B(n5566), .Z(n11999) );
  ANDN U10327 ( .B(n5569), .A(n5568), .Z(n11987) );
  ANDN U10328 ( .B(n5571), .A(n5570), .Z(n11975) );
  NANDN U10329 ( .A(y[886]), .B(x[886]), .Z(n5572) );
  ANDN U10330 ( .B(n5572), .A(n11971), .Z(n8815) );
  NAND U10331 ( .A(n5574), .B(n5573), .Z(n11957) );
  ANDN U10332 ( .B(n5576), .A(n5575), .Z(n11955) );
  NAND U10333 ( .A(n5578), .B(n5577), .Z(n11953) );
  ANDN U10334 ( .B(n5580), .A(n5579), .Z(n11951) );
  AND U10335 ( .A(n5582), .B(n5581), .Z(n11949) );
  ANDN U10336 ( .B(n5584), .A(n5583), .Z(n11947) );
  OR U10337 ( .A(n5590), .B(n5585), .Z(n5586) );
  AND U10338 ( .A(n5587), .B(n5586), .Z(n11945) );
  NAND U10339 ( .A(n5589), .B(n5588), .Z(n5591) );
  ANDN U10340 ( .B(n5591), .A(n5590), .Z(n5592) );
  NANDN U10341 ( .A(n5593), .B(n5592), .Z(n11943) );
  AND U10342 ( .A(n5597), .B(n5596), .Z(n8798) );
  AND U10343 ( .A(n5599), .B(n5598), .Z(n11921) );
  NANDN U10344 ( .A(n5601), .B(n5600), .Z(n11919) );
  AND U10345 ( .A(n5603), .B(n5602), .Z(n11917) );
  NANDN U10346 ( .A(n5605), .B(n5604), .Z(n11915) );
  AND U10347 ( .A(n5607), .B(n5606), .Z(n11913) );
  NANDN U10348 ( .A(n5609), .B(n5608), .Z(n11911) );
  AND U10349 ( .A(n5610), .B(n11908), .Z(n5617) );
  OR U10350 ( .A(n5612), .B(n5611), .Z(n5613) );
  AND U10351 ( .A(n5614), .B(n5613), .Z(n5615) );
  NAND U10352 ( .A(n11907), .B(n5615), .Z(n5616) );
  AND U10353 ( .A(n5617), .B(n5616), .Z(n8780) );
  IV U10354 ( .A(n11907), .Z(n5618) );
  ANDN U10355 ( .B(n11902), .A(n5618), .Z(n8776) );
  AND U10356 ( .A(n5620), .B(n5619), .Z(n11889) );
  NANDN U10357 ( .A(n5622), .B(n5621), .Z(n11887) );
  NAND U10358 ( .A(n5627), .B(n5626), .Z(n5629) );
  ANDN U10359 ( .B(n5629), .A(n5628), .Z(n11872) );
  AND U10360 ( .A(n5631), .B(n5630), .Z(n8751) );
  AND U10361 ( .A(n5633), .B(n5632), .Z(n11847) );
  NAND U10362 ( .A(n5635), .B(n5634), .Z(n11845) );
  AND U10363 ( .A(n5637), .B(n5636), .Z(n11833) );
  NAND U10364 ( .A(n5639), .B(n5638), .Z(n8722) );
  AND U10365 ( .A(n5641), .B(n5640), .Z(n8720) );
  NAND U10366 ( .A(n5643), .B(n5642), .Z(n8710) );
  AND U10367 ( .A(n5645), .B(n5644), .Z(n8708) );
  NOR U10368 ( .A(n5647), .B(n5646), .Z(n8698) );
  AND U10369 ( .A(n5649), .B(n5648), .Z(n8676) );
  ANDN U10370 ( .B(x[802]), .A(y[802]), .Z(n8666) );
  NOR U10371 ( .A(n5651), .B(n5650), .Z(n8650) );
  NOR U10372 ( .A(n5653), .B(n5652), .Z(n8640) );
  AND U10373 ( .A(n5655), .B(n5654), .Z(n8634) );
  NANDN U10374 ( .A(y[790]), .B(x[790]), .Z(n5657) );
  AND U10375 ( .A(n5657), .B(n5656), .Z(n8624) );
  ANDN U10376 ( .B(x[788]), .A(y[788]), .Z(n8618) );
  XNOR U10377 ( .A(y[773]), .B(x[773]), .Z(n8582) );
  AND U10378 ( .A(n5659), .B(n5658), .Z(n8570) );
  NOR U10379 ( .A(n5661), .B(n5660), .Z(n8560) );
  NANDN U10380 ( .A(y[762]), .B(x[762]), .Z(n5662) );
  OR U10381 ( .A(n5663), .B(n5662), .Z(n5665) );
  ANDN U10382 ( .B(n5665), .A(n5664), .Z(n8552) );
  AND U10383 ( .A(n5667), .B(n5666), .Z(n8547) );
  NAND U10384 ( .A(n5669), .B(n5668), .Z(n8533) );
  AND U10385 ( .A(n5671), .B(n5670), .Z(n8531) );
  NAND U10386 ( .A(n5673), .B(n5672), .Z(n8521) );
  AND U10387 ( .A(n5675), .B(n5674), .Z(n8519) );
  NAND U10388 ( .A(n5677), .B(n5676), .Z(n8509) );
  AND U10389 ( .A(n5679), .B(n5678), .Z(n8507) );
  NAND U10390 ( .A(n5681), .B(n5680), .Z(n8497) );
  AND U10391 ( .A(n5683), .B(n5682), .Z(n8495) );
  NAND U10392 ( .A(n5685), .B(n5684), .Z(n8485) );
  AND U10393 ( .A(n5687), .B(n5686), .Z(n8483) );
  NAND U10394 ( .A(n5689), .B(n5688), .Z(n8473) );
  AND U10395 ( .A(n5691), .B(n5690), .Z(n8471) );
  NANDN U10396 ( .A(y[732]), .B(x[732]), .Z(n5692) );
  AND U10397 ( .A(n5693), .B(n5692), .Z(n8461) );
  ANDN U10398 ( .B(x[730]), .A(y[730]), .Z(n8455) );
  ANDN U10399 ( .B(x[726]), .A(y[726]), .Z(n5695) );
  NAND U10400 ( .A(n5695), .B(n5694), .Z(n8445) );
  NAND U10401 ( .A(n5697), .B(n5696), .Z(n8428) );
  AND U10402 ( .A(n5699), .B(n5698), .Z(n8426) );
  XNOR U10403 ( .A(x[712]), .B(y[712]), .Z(n8404) );
  NOR U10404 ( .A(n5701), .B(n5700), .Z(n8400) );
  NAND U10405 ( .A(n5703), .B(n5702), .Z(n8368) );
  ANDN U10406 ( .B(x[696]), .A(y[696]), .Z(n5705) );
  OR U10407 ( .A(n5705), .B(n5704), .Z(n5706) );
  AND U10408 ( .A(n5707), .B(n5706), .Z(n8357) );
  AND U10409 ( .A(n11575), .B(n5708), .Z(n8355) );
  AND U10410 ( .A(n5710), .B(n5709), .Z(n8349) );
  AND U10411 ( .A(n5712), .B(n5711), .Z(n8323) );
  AND U10412 ( .A(n5714), .B(n5713), .Z(n8301) );
  AND U10413 ( .A(n5716), .B(n5715), .Z(n8279) );
  AND U10414 ( .A(n5718), .B(n5717), .Z(n8257) );
  AND U10415 ( .A(n5720), .B(n5719), .Z(n8235) );
  AND U10416 ( .A(n5722), .B(n5721), .Z(n8209) );
  AND U10417 ( .A(n5724), .B(n5723), .Z(n8187) );
  ANDN U10418 ( .B(x[632]), .A(y[632]), .Z(n8177) );
  AND U10419 ( .A(n5726), .B(n5725), .Z(n8165) );
  AND U10420 ( .A(n5728), .B(n5727), .Z(n8143) );
  AND U10421 ( .A(n5730), .B(n5729), .Z(n8121) );
  AND U10422 ( .A(n5732), .B(n5731), .Z(n8099) );
  AND U10423 ( .A(n5734), .B(n5733), .Z(n8077) );
  ANDN U10424 ( .B(x[602]), .A(y[602]), .Z(n8067) );
  AND U10425 ( .A(n5736), .B(n5735), .Z(n8055) );
  ANDN U10426 ( .B(x[596]), .A(y[596]), .Z(n8045) );
  AND U10427 ( .A(n5738), .B(n5737), .Z(n8033) );
  AND U10428 ( .A(n5740), .B(n5739), .Z(n8011) );
  AND U10429 ( .A(n5742), .B(n5741), .Z(n7989) );
  AND U10430 ( .A(n5744), .B(n5743), .Z(n7967) );
  ANDN U10431 ( .B(x[572]), .A(y[572]), .Z(n7957) );
  AND U10432 ( .A(n5746), .B(n5745), .Z(n7945) );
  ANDN U10433 ( .B(x[566]), .A(y[566]), .Z(n7935) );
  AND U10434 ( .A(n5748), .B(n5747), .Z(n7923) );
  AND U10435 ( .A(n5750), .B(n5749), .Z(n7901) );
  AND U10436 ( .A(n5752), .B(n5751), .Z(n7879) );
  ANDN U10437 ( .B(x[548]), .A(y[548]), .Z(n7869) );
  AND U10438 ( .A(n5754), .B(n5753), .Z(n7857) );
  ANDN U10439 ( .B(x[542]), .A(y[542]), .Z(n7847) );
  AND U10440 ( .A(n5756), .B(n5755), .Z(n7835) );
  ANDN U10441 ( .B(x[536]), .A(y[536]), .Z(n7825) );
  ANDN U10442 ( .B(x[534]), .A(y[534]), .Z(n7815) );
  AND U10443 ( .A(n5758), .B(n5757), .Z(n7813) );
  AND U10444 ( .A(n5760), .B(n5759), .Z(n7791) );
  AND U10445 ( .A(n5762), .B(n5761), .Z(n7769) );
  AND U10446 ( .A(n5764), .B(n5763), .Z(n7747) );
  AND U10447 ( .A(n5766), .B(n5765), .Z(n7725) );
  AND U10448 ( .A(n5768), .B(n5767), .Z(n7703) );
  AND U10449 ( .A(n5770), .B(n5769), .Z(n7681) );
  ANDN U10450 ( .B(x[494]), .A(y[494]), .Z(n7671) );
  AND U10451 ( .A(n5772), .B(n5771), .Z(n7659) );
  ANDN U10452 ( .B(x[488]), .A(y[488]), .Z(n7649) );
  AND U10453 ( .A(n5774), .B(n5773), .Z(n7637) );
  ANDN U10454 ( .B(x[482]), .A(y[482]), .Z(n7627) );
  AND U10455 ( .A(n5776), .B(n5775), .Z(n7615) );
  AND U10456 ( .A(n5778), .B(n5777), .Z(n7593) );
  AND U10457 ( .A(n5780), .B(n5779), .Z(n7571) );
  ANDN U10458 ( .B(x[464]), .A(y[464]), .Z(n7561) );
  AND U10459 ( .A(n5782), .B(n5781), .Z(n7549) );
  AND U10460 ( .A(n5784), .B(n5783), .Z(n7527) );
  AND U10461 ( .A(n5786), .B(n5785), .Z(n7505) );
  AND U10462 ( .A(n5788), .B(n5787), .Z(n7483) );
  ANDN U10463 ( .B(x[440]), .A(y[440]), .Z(n7473) );
  AND U10464 ( .A(n5790), .B(n5789), .Z(n7461) );
  AND U10465 ( .A(n5792), .B(n5791), .Z(n7439) );
  AND U10466 ( .A(n5794), .B(n5793), .Z(n7417) );
  ANDN U10467 ( .B(x[422]), .A(y[422]), .Z(n7407) );
  AND U10468 ( .A(n5796), .B(n5795), .Z(n7395) );
  AND U10469 ( .A(n5798), .B(n5797), .Z(n7373) );
  AND U10470 ( .A(n5800), .B(n5799), .Z(n7351) );
  AND U10471 ( .A(n5802), .B(n5801), .Z(n7329) );
  ANDN U10472 ( .B(x[398]), .A(y[398]), .Z(n7319) );
  AND U10473 ( .A(n5804), .B(n5803), .Z(n7307) );
  ANDN U10474 ( .B(x[384]), .A(y[384]), .Z(n7276) );
  XNOR U10475 ( .A(x[378]), .B(y[378]), .Z(n7258) );
  AND U10476 ( .A(n5806), .B(n5805), .Z(n7250) );
  AND U10477 ( .A(n5808), .B(n5807), .Z(n7228) );
  AND U10478 ( .A(n5810), .B(n5809), .Z(n7206) );
  AND U10479 ( .A(n5812), .B(n5811), .Z(n7184) );
  AND U10480 ( .A(n5814), .B(n5813), .Z(n7162) );
  ANDN U10481 ( .B(x[348]), .A(y[348]), .Z(n7152) );
  AND U10482 ( .A(n5816), .B(n5815), .Z(n7140) );
  AND U10483 ( .A(n5818), .B(n5817), .Z(n7118) );
  AND U10484 ( .A(n5820), .B(n5819), .Z(n7096) );
  AND U10485 ( .A(n5822), .B(n5821), .Z(n7074) );
  ANDN U10486 ( .B(x[324]), .A(y[324]), .Z(n7064) );
  AND U10487 ( .A(n5824), .B(n5823), .Z(n7052) );
  AND U10488 ( .A(n5826), .B(n5825), .Z(n7030) );
  AND U10489 ( .A(n5828), .B(n5827), .Z(n7008) );
  ANDN U10490 ( .B(x[306]), .A(y[306]), .Z(n6998) );
  AND U10491 ( .A(n5830), .B(n5829), .Z(n6986) );
  AND U10492 ( .A(n5832), .B(n5831), .Z(n6964) );
  AND U10493 ( .A(n5834), .B(n5833), .Z(n6942) );
  AND U10494 ( .A(n5836), .B(n5835), .Z(n6920) );
  XNOR U10495 ( .A(x[280]), .B(y[280]), .Z(n10739) );
  AND U10496 ( .A(n5841), .B(n5840), .Z(n6873) );
  AND U10497 ( .A(n5843), .B(n5842), .Z(n6851) );
  AND U10498 ( .A(n5845), .B(n5844), .Z(n6829) );
  AND U10499 ( .A(n5847), .B(n5846), .Z(n6807) );
  AND U10500 ( .A(n5849), .B(n5848), .Z(n6785) );
  AND U10501 ( .A(n5851), .B(n5850), .Z(n6763) );
  AND U10502 ( .A(n5853), .B(n5852), .Z(n6741) );
  AND U10503 ( .A(n5855), .B(n5854), .Z(n6719) );
  AND U10504 ( .A(n5857), .B(n5856), .Z(n6697) );
  AND U10505 ( .A(n5859), .B(n5858), .Z(n6675) );
  AND U10506 ( .A(n5861), .B(n5860), .Z(n6653) );
  AND U10507 ( .A(n5863), .B(n5862), .Z(n6631) );
  AND U10508 ( .A(n5865), .B(n5864), .Z(n6609) );
  AND U10509 ( .A(n5867), .B(n5866), .Z(n6587) );
  AND U10510 ( .A(n5869), .B(n5868), .Z(n6565) );
  AND U10511 ( .A(n5871), .B(n5870), .Z(n6543) );
  AND U10512 ( .A(n5873), .B(n5872), .Z(n6521) );
  AND U10513 ( .A(n5875), .B(n5874), .Z(n6499) );
  AND U10514 ( .A(n5879), .B(n5878), .Z(n6462) );
  AND U10515 ( .A(n5880), .B(n10469), .Z(n6440) );
  AND U10516 ( .A(n5882), .B(n5881), .Z(n6418) );
  AND U10517 ( .A(n5884), .B(n5883), .Z(n6396) );
  OR U10518 ( .A(n5886), .B(n5885), .Z(n5887) );
  AND U10519 ( .A(n5888), .B(n5887), .Z(n6380) );
  AND U10520 ( .A(n5890), .B(n5889), .Z(n6363) );
  AND U10521 ( .A(n5892), .B(n5891), .Z(n6341) );
  AND U10522 ( .A(n5894), .B(n5893), .Z(n6319) );
  AND U10523 ( .A(n5896), .B(n5895), .Z(n6297) );
  AND U10524 ( .A(n5898), .B(n5897), .Z(n6275) );
  AND U10525 ( .A(n5900), .B(n5899), .Z(n6253) );
  AND U10526 ( .A(n5902), .B(n5901), .Z(n6231) );
  AND U10527 ( .A(n5904), .B(n5903), .Z(n6209) );
  XNOR U10528 ( .A(x[76]), .B(y[76]), .Z(n6195) );
  AND U10529 ( .A(n5906), .B(n5905), .Z(n6179) );
  AND U10530 ( .A(n5908), .B(n5907), .Z(n6157) );
  AND U10531 ( .A(n5910), .B(n5909), .Z(n6135) );
  AND U10532 ( .A(n5912), .B(n5911), .Z(n6113) );
  AND U10533 ( .A(n5914), .B(n5913), .Z(n6091) );
  AND U10534 ( .A(n5916), .B(n5915), .Z(n6069) );
  AND U10535 ( .A(n5918), .B(n5917), .Z(n6047) );
  ANDN U10536 ( .B(x[30]), .A(y[30]), .Z(n6027) );
  AND U10537 ( .A(n5920), .B(n5919), .Z(n6025) );
  AND U10538 ( .A(n5922), .B(n5921), .Z(n6003) );
  AND U10539 ( .A(n5924), .B(n5923), .Z(n5981) );
  AND U10540 ( .A(n5926), .B(n5925), .Z(n5959) );
  ANDN U10541 ( .B(n5927), .A(y[0]), .Z(n5928) );
  NAND U10542 ( .A(x[0]), .B(n5928), .Z(n5930) );
  ANDN U10543 ( .B(n5930), .A(n5929), .Z(n5932) );
  NANDN U10544 ( .A(n5932), .B(n5931), .Z(n5933) );
  NANDN U10545 ( .A(n5934), .B(n5933), .Z(n5935) );
  NAND U10546 ( .A(n5936), .B(n5935), .Z(n5937) );
  NANDN U10547 ( .A(n5938), .B(n5937), .Z(n10192) );
  NAND U10548 ( .A(n5939), .B(n10192), .Z(n5940) );
  NANDN U10549 ( .A(n5941), .B(n5940), .Z(n5942) );
  AND U10550 ( .A(n5943), .B(n5942), .Z(n5945) );
  NAND U10551 ( .A(n5945), .B(n5944), .Z(n5947) );
  ANDN U10552 ( .B(x[8]), .A(y[8]), .Z(n5946) );
  ANDN U10553 ( .B(n5947), .A(n5946), .Z(n5948) );
  NANDN U10554 ( .A(n5949), .B(n5948), .Z(n5953) );
  AND U10555 ( .A(n5951), .B(n5950), .Z(n5952) );
  NAND U10556 ( .A(n5953), .B(n5952), .Z(n5954) );
  NANDN U10557 ( .A(n5955), .B(n5954), .Z(n5957) );
  OR U10558 ( .A(n5957), .B(n5956), .Z(n5958) );
  AND U10559 ( .A(n5959), .B(n5958), .Z(n5961) );
  NOR U10560 ( .A(n5961), .B(n5960), .Z(n5962) );
  NANDN U10561 ( .A(n5963), .B(n5962), .Z(n5964) );
  AND U10562 ( .A(n5965), .B(n5964), .Z(n5967) );
  NAND U10563 ( .A(n5967), .B(n5966), .Z(n5969) );
  ANDN U10564 ( .B(n5969), .A(n5968), .Z(n5970) );
  NANDN U10565 ( .A(n5971), .B(n5970), .Z(n5975) );
  AND U10566 ( .A(n5973), .B(n5972), .Z(n5974) );
  NAND U10567 ( .A(n5975), .B(n5974), .Z(n5976) );
  NANDN U10568 ( .A(n5977), .B(n5976), .Z(n5979) );
  OR U10569 ( .A(n5979), .B(n5978), .Z(n5980) );
  AND U10570 ( .A(n5981), .B(n5980), .Z(n5983) );
  NOR U10571 ( .A(n5983), .B(n5982), .Z(n5984) );
  NANDN U10572 ( .A(n5985), .B(n5984), .Z(n5986) );
  AND U10573 ( .A(n5987), .B(n5986), .Z(n5989) );
  NAND U10574 ( .A(n5989), .B(n5988), .Z(n5991) );
  ANDN U10575 ( .B(n5991), .A(n5990), .Z(n5992) );
  NANDN U10576 ( .A(n5993), .B(n5992), .Z(n5997) );
  AND U10577 ( .A(n5995), .B(n5994), .Z(n5996) );
  NAND U10578 ( .A(n5997), .B(n5996), .Z(n5998) );
  NANDN U10579 ( .A(n5999), .B(n5998), .Z(n6001) );
  OR U10580 ( .A(n6001), .B(n6000), .Z(n6002) );
  AND U10581 ( .A(n6003), .B(n6002), .Z(n6005) );
  NOR U10582 ( .A(n6005), .B(n6004), .Z(n6006) );
  NANDN U10583 ( .A(n6007), .B(n6006), .Z(n6008) );
  AND U10584 ( .A(n6009), .B(n6008), .Z(n6011) );
  NAND U10585 ( .A(n6011), .B(n6010), .Z(n6013) );
  ANDN U10586 ( .B(n6013), .A(n6012), .Z(n6014) );
  NANDN U10587 ( .A(n6015), .B(n6014), .Z(n6019) );
  AND U10588 ( .A(n6017), .B(n6016), .Z(n6018) );
  NAND U10589 ( .A(n6019), .B(n6018), .Z(n6020) );
  NANDN U10590 ( .A(n6021), .B(n6020), .Z(n6023) );
  OR U10591 ( .A(n6023), .B(n6022), .Z(n6024) );
  AND U10592 ( .A(n6025), .B(n6024), .Z(n6026) );
  NOR U10593 ( .A(n6027), .B(n6026), .Z(n6028) );
  NANDN U10594 ( .A(n6029), .B(n6028), .Z(n6030) );
  AND U10595 ( .A(n6031), .B(n6030), .Z(n6033) );
  NAND U10596 ( .A(n6033), .B(n6032), .Z(n6035) );
  ANDN U10597 ( .B(n6035), .A(n6034), .Z(n6036) );
  NANDN U10598 ( .A(n6037), .B(n6036), .Z(n6041) );
  AND U10599 ( .A(n6039), .B(n6038), .Z(n6040) );
  NAND U10600 ( .A(n6041), .B(n6040), .Z(n6042) );
  NANDN U10601 ( .A(n6043), .B(n6042), .Z(n6045) );
  OR U10602 ( .A(n6045), .B(n6044), .Z(n6046) );
  AND U10603 ( .A(n6047), .B(n6046), .Z(n6049) );
  NOR U10604 ( .A(n6049), .B(n6048), .Z(n6050) );
  NANDN U10605 ( .A(n6051), .B(n6050), .Z(n6052) );
  AND U10606 ( .A(n6053), .B(n6052), .Z(n6055) );
  NAND U10607 ( .A(n6055), .B(n6054), .Z(n6057) );
  ANDN U10608 ( .B(n6057), .A(n6056), .Z(n6058) );
  NANDN U10609 ( .A(n6059), .B(n6058), .Z(n6063) );
  AND U10610 ( .A(n6061), .B(n6060), .Z(n6062) );
  NAND U10611 ( .A(n6063), .B(n6062), .Z(n6064) );
  NANDN U10612 ( .A(n6065), .B(n6064), .Z(n6067) );
  OR U10613 ( .A(n6067), .B(n6066), .Z(n6068) );
  AND U10614 ( .A(n6069), .B(n6068), .Z(n6071) );
  NOR U10615 ( .A(n6071), .B(n6070), .Z(n6072) );
  NANDN U10616 ( .A(n6073), .B(n6072), .Z(n6074) );
  AND U10617 ( .A(n6075), .B(n6074), .Z(n6077) );
  NAND U10618 ( .A(n6077), .B(n6076), .Z(n6079) );
  ANDN U10619 ( .B(n6079), .A(n6078), .Z(n6080) );
  NANDN U10620 ( .A(n6081), .B(n6080), .Z(n6085) );
  AND U10621 ( .A(n6083), .B(n6082), .Z(n6084) );
  NAND U10622 ( .A(n6085), .B(n6084), .Z(n6086) );
  NANDN U10623 ( .A(n6087), .B(n6086), .Z(n6089) );
  OR U10624 ( .A(n6089), .B(n6088), .Z(n6090) );
  AND U10625 ( .A(n6091), .B(n6090), .Z(n6093) );
  NOR U10626 ( .A(n6093), .B(n6092), .Z(n6094) );
  NANDN U10627 ( .A(n6095), .B(n6094), .Z(n6096) );
  AND U10628 ( .A(n6097), .B(n6096), .Z(n6099) );
  NAND U10629 ( .A(n6099), .B(n6098), .Z(n6101) );
  ANDN U10630 ( .B(n6101), .A(n6100), .Z(n6102) );
  NANDN U10631 ( .A(n6103), .B(n6102), .Z(n6107) );
  AND U10632 ( .A(n6105), .B(n6104), .Z(n6106) );
  NAND U10633 ( .A(n6107), .B(n6106), .Z(n6108) );
  NANDN U10634 ( .A(n6109), .B(n6108), .Z(n6111) );
  OR U10635 ( .A(n6111), .B(n6110), .Z(n6112) );
  AND U10636 ( .A(n6113), .B(n6112), .Z(n6115) );
  NOR U10637 ( .A(n6115), .B(n6114), .Z(n6116) );
  NANDN U10638 ( .A(n6117), .B(n6116), .Z(n6118) );
  AND U10639 ( .A(n6119), .B(n6118), .Z(n6121) );
  NAND U10640 ( .A(n6121), .B(n6120), .Z(n6123) );
  ANDN U10641 ( .B(n6123), .A(n6122), .Z(n6124) );
  NANDN U10642 ( .A(n6125), .B(n6124), .Z(n6129) );
  AND U10643 ( .A(n6127), .B(n6126), .Z(n6128) );
  NAND U10644 ( .A(n6129), .B(n6128), .Z(n6130) );
  NANDN U10645 ( .A(n6131), .B(n6130), .Z(n6133) );
  OR U10646 ( .A(n6133), .B(n6132), .Z(n6134) );
  AND U10647 ( .A(n6135), .B(n6134), .Z(n6137) );
  NOR U10648 ( .A(n6137), .B(n6136), .Z(n6138) );
  NANDN U10649 ( .A(n6139), .B(n6138), .Z(n6140) );
  AND U10650 ( .A(n6141), .B(n6140), .Z(n6143) );
  NAND U10651 ( .A(n6143), .B(n6142), .Z(n6145) );
  ANDN U10652 ( .B(n6145), .A(n6144), .Z(n6146) );
  NANDN U10653 ( .A(n6147), .B(n6146), .Z(n6151) );
  AND U10654 ( .A(n6149), .B(n6148), .Z(n6150) );
  NAND U10655 ( .A(n6151), .B(n6150), .Z(n6152) );
  NANDN U10656 ( .A(n6153), .B(n6152), .Z(n6155) );
  OR U10657 ( .A(n6155), .B(n6154), .Z(n6156) );
  AND U10658 ( .A(n6157), .B(n6156), .Z(n6159) );
  NOR U10659 ( .A(n6159), .B(n6158), .Z(n6160) );
  NANDN U10660 ( .A(n6161), .B(n6160), .Z(n6162) );
  AND U10661 ( .A(n6163), .B(n6162), .Z(n6165) );
  NAND U10662 ( .A(n6165), .B(n6164), .Z(n6167) );
  ANDN U10663 ( .B(n6167), .A(n6166), .Z(n6168) );
  NANDN U10664 ( .A(n6169), .B(n6168), .Z(n6173) );
  AND U10665 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U10666 ( .A(n6173), .B(n6172), .Z(n6174) );
  NANDN U10667 ( .A(n6175), .B(n6174), .Z(n6177) );
  OR U10668 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U10669 ( .A(n6179), .B(n6178), .Z(n6181) );
  NOR U10670 ( .A(n6181), .B(n6180), .Z(n6182) );
  NANDN U10671 ( .A(n6183), .B(n6182), .Z(n6184) );
  AND U10672 ( .A(n6185), .B(n6184), .Z(n6187) );
  NAND U10673 ( .A(n6187), .B(n6186), .Z(n6189) );
  ANDN U10674 ( .B(n6189), .A(n6188), .Z(n6190) );
  NANDN U10675 ( .A(n6191), .B(n6190), .Z(n6193) );
  AND U10676 ( .A(n6193), .B(n6192), .Z(n6194) );
  NAND U10677 ( .A(n6195), .B(n6194), .Z(n6196) );
  NAND U10678 ( .A(n6197), .B(n6196), .Z(n6198) );
  AND U10679 ( .A(n6199), .B(n6198), .Z(n6201) );
  OR U10680 ( .A(n6201), .B(n6200), .Z(n6202) );
  NAND U10681 ( .A(n6203), .B(n6202), .Z(n6204) );
  NANDN U10682 ( .A(n6205), .B(n6204), .Z(n6207) );
  OR U10683 ( .A(n6207), .B(n6206), .Z(n6208) );
  AND U10684 ( .A(n6209), .B(n6208), .Z(n6211) );
  NOR U10685 ( .A(n6211), .B(n6210), .Z(n6212) );
  NANDN U10686 ( .A(n6213), .B(n6212), .Z(n6214) );
  AND U10687 ( .A(n6215), .B(n6214), .Z(n6217) );
  NAND U10688 ( .A(n6217), .B(n6216), .Z(n6219) );
  ANDN U10689 ( .B(n6219), .A(n6218), .Z(n6220) );
  NANDN U10690 ( .A(n6221), .B(n6220), .Z(n6225) );
  AND U10691 ( .A(n6223), .B(n6222), .Z(n6224) );
  NAND U10692 ( .A(n6225), .B(n6224), .Z(n6226) );
  NANDN U10693 ( .A(n6227), .B(n6226), .Z(n6229) );
  OR U10694 ( .A(n6229), .B(n6228), .Z(n6230) );
  AND U10695 ( .A(n6231), .B(n6230), .Z(n6233) );
  NOR U10696 ( .A(n6233), .B(n6232), .Z(n6234) );
  NANDN U10697 ( .A(n6235), .B(n6234), .Z(n6236) );
  AND U10698 ( .A(n6237), .B(n6236), .Z(n6239) );
  NAND U10699 ( .A(n6239), .B(n6238), .Z(n6241) );
  ANDN U10700 ( .B(n6241), .A(n6240), .Z(n6242) );
  NANDN U10701 ( .A(n6243), .B(n6242), .Z(n6247) );
  AND U10702 ( .A(n6245), .B(n6244), .Z(n6246) );
  NAND U10703 ( .A(n6247), .B(n6246), .Z(n6248) );
  NANDN U10704 ( .A(n6249), .B(n6248), .Z(n6251) );
  OR U10705 ( .A(n6251), .B(n6250), .Z(n6252) );
  AND U10706 ( .A(n6253), .B(n6252), .Z(n6255) );
  NOR U10707 ( .A(n6255), .B(n6254), .Z(n6256) );
  NANDN U10708 ( .A(n6257), .B(n6256), .Z(n6258) );
  AND U10709 ( .A(n6259), .B(n6258), .Z(n6261) );
  NAND U10710 ( .A(n6261), .B(n6260), .Z(n6263) );
  ANDN U10711 ( .B(n6263), .A(n6262), .Z(n6264) );
  NANDN U10712 ( .A(n6265), .B(n6264), .Z(n6269) );
  AND U10713 ( .A(n6267), .B(n6266), .Z(n6268) );
  NAND U10714 ( .A(n6269), .B(n6268), .Z(n6270) );
  NANDN U10715 ( .A(n6271), .B(n6270), .Z(n6273) );
  OR U10716 ( .A(n6273), .B(n6272), .Z(n6274) );
  AND U10717 ( .A(n6275), .B(n6274), .Z(n6277) );
  NOR U10718 ( .A(n6277), .B(n6276), .Z(n6278) );
  NANDN U10719 ( .A(n6279), .B(n6278), .Z(n6280) );
  AND U10720 ( .A(n6281), .B(n6280), .Z(n6283) );
  NAND U10721 ( .A(n6283), .B(n6282), .Z(n6285) );
  ANDN U10722 ( .B(n6285), .A(n6284), .Z(n6286) );
  NANDN U10723 ( .A(n6287), .B(n6286), .Z(n6291) );
  AND U10724 ( .A(n6289), .B(n6288), .Z(n6290) );
  NAND U10725 ( .A(n6291), .B(n6290), .Z(n6292) );
  NANDN U10726 ( .A(n6293), .B(n6292), .Z(n6295) );
  OR U10727 ( .A(n6295), .B(n6294), .Z(n6296) );
  AND U10728 ( .A(n6297), .B(n6296), .Z(n6299) );
  NOR U10729 ( .A(n6299), .B(n6298), .Z(n6300) );
  NANDN U10730 ( .A(n6301), .B(n6300), .Z(n6302) );
  AND U10731 ( .A(n6303), .B(n6302), .Z(n6305) );
  NAND U10732 ( .A(n6305), .B(n6304), .Z(n6307) );
  ANDN U10733 ( .B(n6307), .A(n6306), .Z(n6308) );
  NANDN U10734 ( .A(n6309), .B(n6308), .Z(n6313) );
  AND U10735 ( .A(n6311), .B(n6310), .Z(n6312) );
  NAND U10736 ( .A(n6313), .B(n6312), .Z(n6314) );
  NANDN U10737 ( .A(n6315), .B(n6314), .Z(n6317) );
  OR U10738 ( .A(n6317), .B(n6316), .Z(n6318) );
  AND U10739 ( .A(n6319), .B(n6318), .Z(n6321) );
  NOR U10740 ( .A(n6321), .B(n6320), .Z(n6322) );
  NANDN U10741 ( .A(n6323), .B(n6322), .Z(n6324) );
  AND U10742 ( .A(n6325), .B(n6324), .Z(n6327) );
  NAND U10743 ( .A(n6327), .B(n6326), .Z(n6329) );
  ANDN U10744 ( .B(n6329), .A(n6328), .Z(n6330) );
  NANDN U10745 ( .A(n6331), .B(n6330), .Z(n6335) );
  AND U10746 ( .A(n6333), .B(n6332), .Z(n6334) );
  NAND U10747 ( .A(n6335), .B(n6334), .Z(n6336) );
  NANDN U10748 ( .A(n6337), .B(n6336), .Z(n6339) );
  OR U10749 ( .A(n6339), .B(n6338), .Z(n6340) );
  AND U10750 ( .A(n6341), .B(n6340), .Z(n6343) );
  NOR U10751 ( .A(n6343), .B(n6342), .Z(n6344) );
  NANDN U10752 ( .A(n6345), .B(n6344), .Z(n6346) );
  AND U10753 ( .A(n6347), .B(n6346), .Z(n6349) );
  NAND U10754 ( .A(n6349), .B(n6348), .Z(n6351) );
  ANDN U10755 ( .B(n6351), .A(n6350), .Z(n6352) );
  NANDN U10756 ( .A(n6353), .B(n6352), .Z(n6357) );
  AND U10757 ( .A(n6355), .B(n6354), .Z(n6356) );
  NAND U10758 ( .A(n6357), .B(n6356), .Z(n6358) );
  NANDN U10759 ( .A(n6359), .B(n6358), .Z(n6361) );
  OR U10760 ( .A(n6361), .B(n6360), .Z(n6362) );
  AND U10761 ( .A(n6363), .B(n6362), .Z(n6365) );
  NOR U10762 ( .A(n6365), .B(n6364), .Z(n6366) );
  NANDN U10763 ( .A(n6367), .B(n6366), .Z(n6368) );
  AND U10764 ( .A(n6369), .B(n6368), .Z(n6371) );
  NAND U10765 ( .A(n6371), .B(n6370), .Z(n6373) );
  ANDN U10766 ( .B(n6373), .A(n6372), .Z(n6374) );
  NANDN U10767 ( .A(n6375), .B(n6374), .Z(n6378) );
  AND U10768 ( .A(n10433), .B(n6376), .Z(n6377) );
  NAND U10769 ( .A(n6378), .B(n6377), .Z(n6379) );
  NANDN U10770 ( .A(n6380), .B(n6379), .Z(n6382) );
  NAND U10771 ( .A(n6382), .B(n6381), .Z(n6384) );
  ANDN U10772 ( .B(n6384), .A(n6383), .Z(n6385) );
  NANDN U10773 ( .A(n6386), .B(n6385), .Z(n6390) );
  AND U10774 ( .A(n6388), .B(n6387), .Z(n6389) );
  NAND U10775 ( .A(n6390), .B(n6389), .Z(n6391) );
  NANDN U10776 ( .A(n6392), .B(n6391), .Z(n6394) );
  OR U10777 ( .A(n6394), .B(n6393), .Z(n6395) );
  AND U10778 ( .A(n6396), .B(n6395), .Z(n6398) );
  NOR U10779 ( .A(n6398), .B(n6397), .Z(n6399) );
  NANDN U10780 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U10781 ( .A(n6402), .B(n6401), .Z(n6404) );
  NAND U10782 ( .A(n6404), .B(n6403), .Z(n6406) );
  ANDN U10783 ( .B(n6406), .A(n6405), .Z(n6407) );
  NANDN U10784 ( .A(n6408), .B(n6407), .Z(n6412) );
  AND U10785 ( .A(n6410), .B(n6409), .Z(n6411) );
  NAND U10786 ( .A(n6412), .B(n6411), .Z(n6413) );
  NANDN U10787 ( .A(n6414), .B(n6413), .Z(n6416) );
  OR U10788 ( .A(n6416), .B(n6415), .Z(n6417) );
  AND U10789 ( .A(n6418), .B(n6417), .Z(n6420) );
  NOR U10790 ( .A(n6420), .B(n6419), .Z(n6421) );
  NANDN U10791 ( .A(n6422), .B(n6421), .Z(n6423) );
  AND U10792 ( .A(n6424), .B(n6423), .Z(n6426) );
  NAND U10793 ( .A(n6426), .B(n6425), .Z(n6428) );
  ANDN U10794 ( .B(n6428), .A(n6427), .Z(n6429) );
  NANDN U10795 ( .A(n6430), .B(n6429), .Z(n6434) );
  AND U10796 ( .A(n6432), .B(n6431), .Z(n6433) );
  NAND U10797 ( .A(n6434), .B(n6433), .Z(n6435) );
  NANDN U10798 ( .A(n6436), .B(n6435), .Z(n6438) );
  OR U10799 ( .A(n6438), .B(n6437), .Z(n6439) );
  AND U10800 ( .A(n6440), .B(n6439), .Z(n6446) );
  OR U10801 ( .A(n6442), .B(n6441), .Z(n6443) );
  NAND U10802 ( .A(n6444), .B(n6443), .Z(n6445) );
  NANDN U10803 ( .A(n6446), .B(n6445), .Z(n6448) );
  NAND U10804 ( .A(n6448), .B(n6447), .Z(n6450) );
  ANDN U10805 ( .B(n6450), .A(n6449), .Z(n6451) );
  NANDN U10806 ( .A(n6452), .B(n6451), .Z(n6456) );
  AND U10807 ( .A(n6454), .B(n6453), .Z(n6455) );
  NAND U10808 ( .A(n6456), .B(n6455), .Z(n6457) );
  NANDN U10809 ( .A(n6458), .B(n6457), .Z(n6460) );
  OR U10810 ( .A(n6460), .B(n6459), .Z(n6461) );
  AND U10811 ( .A(n6462), .B(n6461), .Z(n6464) );
  NOR U10812 ( .A(n6464), .B(n6463), .Z(n6465) );
  NANDN U10813 ( .A(n6466), .B(n6465), .Z(n6467) );
  AND U10814 ( .A(n6483), .B(n6482), .Z(n6485) );
  NAND U10815 ( .A(n6485), .B(n6484), .Z(n6487) );
  ANDN U10816 ( .B(n6487), .A(n6486), .Z(n6488) );
  NANDN U10817 ( .A(n6489), .B(n6488), .Z(n6493) );
  AND U10818 ( .A(n6491), .B(n6490), .Z(n6492) );
  NAND U10819 ( .A(n6493), .B(n6492), .Z(n6494) );
  NANDN U10820 ( .A(n6495), .B(n6494), .Z(n6497) );
  OR U10821 ( .A(n6497), .B(n6496), .Z(n6498) );
  AND U10822 ( .A(n6499), .B(n6498), .Z(n6501) );
  NOR U10823 ( .A(n6501), .B(n6500), .Z(n6502) );
  NANDN U10824 ( .A(n6503), .B(n6502), .Z(n6504) );
  AND U10825 ( .A(n6505), .B(n6504), .Z(n6507) );
  NAND U10826 ( .A(n6507), .B(n6506), .Z(n6509) );
  ANDN U10827 ( .B(n6509), .A(n6508), .Z(n6510) );
  NANDN U10828 ( .A(n6511), .B(n6510), .Z(n6515) );
  AND U10829 ( .A(n6513), .B(n6512), .Z(n6514) );
  NAND U10830 ( .A(n6515), .B(n6514), .Z(n6516) );
  NANDN U10831 ( .A(n6517), .B(n6516), .Z(n6519) );
  OR U10832 ( .A(n6519), .B(n6518), .Z(n6520) );
  AND U10833 ( .A(n6521), .B(n6520), .Z(n6523) );
  NOR U10834 ( .A(n6523), .B(n6522), .Z(n6524) );
  NANDN U10835 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U10836 ( .A(n6527), .B(n6526), .Z(n6529) );
  NAND U10837 ( .A(n6529), .B(n6528), .Z(n6531) );
  ANDN U10838 ( .B(n6531), .A(n6530), .Z(n6532) );
  NANDN U10839 ( .A(n6533), .B(n6532), .Z(n6537) );
  AND U10840 ( .A(n6535), .B(n6534), .Z(n6536) );
  NAND U10841 ( .A(n6537), .B(n6536), .Z(n6538) );
  NANDN U10842 ( .A(n6539), .B(n6538), .Z(n6541) );
  OR U10843 ( .A(n6541), .B(n6540), .Z(n6542) );
  AND U10844 ( .A(n6543), .B(n6542), .Z(n6545) );
  NOR U10845 ( .A(n6545), .B(n6544), .Z(n6546) );
  NANDN U10846 ( .A(n6547), .B(n6546), .Z(n6548) );
  AND U10847 ( .A(n6549), .B(n6548), .Z(n6551) );
  NAND U10848 ( .A(n6551), .B(n6550), .Z(n6553) );
  ANDN U10849 ( .B(x[180]), .A(y[180]), .Z(n6552) );
  ANDN U10850 ( .B(n6553), .A(n6552), .Z(n6554) );
  NANDN U10851 ( .A(n6555), .B(n6554), .Z(n6559) );
  AND U10852 ( .A(n6557), .B(n6556), .Z(n6558) );
  NAND U10853 ( .A(n6559), .B(n6558), .Z(n6560) );
  NANDN U10854 ( .A(n6561), .B(n6560), .Z(n6563) );
  OR U10855 ( .A(n6563), .B(n6562), .Z(n6564) );
  AND U10856 ( .A(n6565), .B(n6564), .Z(n6567) );
  NOR U10857 ( .A(n6567), .B(n6566), .Z(n6568) );
  NANDN U10858 ( .A(n6569), .B(n6568), .Z(n6570) );
  AND U10859 ( .A(n6571), .B(n6570), .Z(n6573) );
  NAND U10860 ( .A(n6573), .B(n6572), .Z(n6575) );
  ANDN U10861 ( .B(n6575), .A(n6574), .Z(n6576) );
  NANDN U10862 ( .A(n6577), .B(n6576), .Z(n6581) );
  AND U10863 ( .A(n6579), .B(n6578), .Z(n6580) );
  NAND U10864 ( .A(n6581), .B(n6580), .Z(n6582) );
  NANDN U10865 ( .A(n6583), .B(n6582), .Z(n6585) );
  OR U10866 ( .A(n6585), .B(n6584), .Z(n6586) );
  AND U10867 ( .A(n6587), .B(n6586), .Z(n6589) );
  NOR U10868 ( .A(n6589), .B(n6588), .Z(n6590) );
  NANDN U10869 ( .A(n6591), .B(n6590), .Z(n6592) );
  AND U10870 ( .A(n6593), .B(n6592), .Z(n6595) );
  NAND U10871 ( .A(n6595), .B(n6594), .Z(n6597) );
  ANDN U10872 ( .B(n6597), .A(n6596), .Z(n6598) );
  NANDN U10873 ( .A(n6599), .B(n6598), .Z(n6603) );
  AND U10874 ( .A(n6601), .B(n6600), .Z(n6602) );
  NAND U10875 ( .A(n6603), .B(n6602), .Z(n6604) );
  NANDN U10876 ( .A(n6605), .B(n6604), .Z(n6607) );
  OR U10877 ( .A(n6607), .B(n6606), .Z(n6608) );
  AND U10878 ( .A(n6609), .B(n6608), .Z(n6611) );
  NOR U10879 ( .A(n6611), .B(n6610), .Z(n6612) );
  NANDN U10880 ( .A(n6613), .B(n6612), .Z(n6614) );
  AND U10881 ( .A(n6615), .B(n6614), .Z(n6617) );
  NAND U10882 ( .A(n6617), .B(n6616), .Z(n6619) );
  ANDN U10883 ( .B(n6619), .A(n6618), .Z(n6620) );
  NANDN U10884 ( .A(n6621), .B(n6620), .Z(n6625) );
  AND U10885 ( .A(n6623), .B(n6622), .Z(n6624) );
  NAND U10886 ( .A(n6625), .B(n6624), .Z(n6626) );
  NANDN U10887 ( .A(n6627), .B(n6626), .Z(n6629) );
  OR U10888 ( .A(n6629), .B(n6628), .Z(n6630) );
  AND U10889 ( .A(n6631), .B(n6630), .Z(n6633) );
  NOR U10890 ( .A(n6633), .B(n6632), .Z(n6634) );
  NANDN U10891 ( .A(n6635), .B(n6634), .Z(n6636) );
  AND U10892 ( .A(n6637), .B(n6636), .Z(n6639) );
  NAND U10893 ( .A(n6639), .B(n6638), .Z(n6641) );
  ANDN U10894 ( .B(x[204]), .A(y[204]), .Z(n6640) );
  ANDN U10895 ( .B(n6641), .A(n6640), .Z(n6642) );
  NANDN U10896 ( .A(n6643), .B(n6642), .Z(n6647) );
  AND U10897 ( .A(n6645), .B(n6644), .Z(n6646) );
  NAND U10898 ( .A(n6647), .B(n6646), .Z(n6648) );
  NANDN U10899 ( .A(n6649), .B(n6648), .Z(n6651) );
  OR U10900 ( .A(n6651), .B(n6650), .Z(n6652) );
  AND U10901 ( .A(n6653), .B(n6652), .Z(n6655) );
  NOR U10902 ( .A(n6655), .B(n6654), .Z(n6656) );
  NANDN U10903 ( .A(n6657), .B(n6656), .Z(n6658) );
  AND U10904 ( .A(n6659), .B(n6658), .Z(n6661) );
  NAND U10905 ( .A(n6661), .B(n6660), .Z(n6663) );
  ANDN U10906 ( .B(n6663), .A(n6662), .Z(n6664) );
  NANDN U10907 ( .A(n6665), .B(n6664), .Z(n6669) );
  AND U10908 ( .A(n6667), .B(n6666), .Z(n6668) );
  NAND U10909 ( .A(n6669), .B(n6668), .Z(n6670) );
  NANDN U10910 ( .A(n6671), .B(n6670), .Z(n6673) );
  OR U10911 ( .A(n6673), .B(n6672), .Z(n6674) );
  AND U10912 ( .A(n6675), .B(n6674), .Z(n6677) );
  NOR U10913 ( .A(n6677), .B(n6676), .Z(n6678) );
  NANDN U10914 ( .A(n6679), .B(n6678), .Z(n6680) );
  AND U10915 ( .A(n6681), .B(n6680), .Z(n6683) );
  NAND U10916 ( .A(n6683), .B(n6682), .Z(n6685) );
  ANDN U10917 ( .B(x[216]), .A(y[216]), .Z(n6684) );
  ANDN U10918 ( .B(n6685), .A(n6684), .Z(n6686) );
  NANDN U10919 ( .A(n6687), .B(n6686), .Z(n6691) );
  AND U10920 ( .A(n6689), .B(n6688), .Z(n6690) );
  NAND U10921 ( .A(n6691), .B(n6690), .Z(n6692) );
  NANDN U10922 ( .A(n6693), .B(n6692), .Z(n6695) );
  OR U10923 ( .A(n6695), .B(n6694), .Z(n6696) );
  AND U10924 ( .A(n6697), .B(n6696), .Z(n6699) );
  NOR U10925 ( .A(n6699), .B(n6698), .Z(n6700) );
  NANDN U10926 ( .A(n6701), .B(n6700), .Z(n6702) );
  AND U10927 ( .A(n6703), .B(n6702), .Z(n6705) );
  NAND U10928 ( .A(n6705), .B(n6704), .Z(n6707) );
  ANDN U10929 ( .B(n6707), .A(n6706), .Z(n6708) );
  NANDN U10930 ( .A(n6709), .B(n6708), .Z(n6713) );
  AND U10931 ( .A(n6711), .B(n6710), .Z(n6712) );
  NAND U10932 ( .A(n6713), .B(n6712), .Z(n6714) );
  NANDN U10933 ( .A(n6715), .B(n6714), .Z(n6717) );
  OR U10934 ( .A(n6717), .B(n6716), .Z(n6718) );
  AND U10935 ( .A(n6719), .B(n6718), .Z(n6721) );
  NOR U10936 ( .A(n6721), .B(n6720), .Z(n6722) );
  NANDN U10937 ( .A(n6723), .B(n6722), .Z(n6724) );
  AND U10938 ( .A(n6725), .B(n6724), .Z(n6727) );
  NAND U10939 ( .A(n6727), .B(n6726), .Z(n6729) );
  ANDN U10940 ( .B(n6729), .A(n6728), .Z(n6730) );
  NANDN U10941 ( .A(n6731), .B(n6730), .Z(n6735) );
  AND U10942 ( .A(n6733), .B(n6732), .Z(n6734) );
  NAND U10943 ( .A(n6735), .B(n6734), .Z(n6736) );
  NANDN U10944 ( .A(n6737), .B(n6736), .Z(n6739) );
  OR U10945 ( .A(n6739), .B(n6738), .Z(n6740) );
  AND U10946 ( .A(n6741), .B(n6740), .Z(n6743) );
  NOR U10947 ( .A(n6743), .B(n6742), .Z(n6744) );
  NANDN U10948 ( .A(n6745), .B(n6744), .Z(n6746) );
  AND U10949 ( .A(n6747), .B(n6746), .Z(n6749) );
  NAND U10950 ( .A(n6749), .B(n6748), .Z(n6751) );
  ANDN U10951 ( .B(n6751), .A(n6750), .Z(n6752) );
  NANDN U10952 ( .A(n6753), .B(n6752), .Z(n6757) );
  AND U10953 ( .A(n6755), .B(n6754), .Z(n6756) );
  NAND U10954 ( .A(n6757), .B(n6756), .Z(n6758) );
  NANDN U10955 ( .A(n6759), .B(n6758), .Z(n6761) );
  OR U10956 ( .A(n6761), .B(n6760), .Z(n6762) );
  AND U10957 ( .A(n6763), .B(n6762), .Z(n6765) );
  NOR U10958 ( .A(n6765), .B(n6764), .Z(n6766) );
  NANDN U10959 ( .A(n6767), .B(n6766), .Z(n6768) );
  AND U10960 ( .A(n6769), .B(n6768), .Z(n6771) );
  NAND U10961 ( .A(n6771), .B(n6770), .Z(n6773) );
  ANDN U10962 ( .B(n6773), .A(n6772), .Z(n6774) );
  NANDN U10963 ( .A(n6775), .B(n6774), .Z(n6779) );
  AND U10964 ( .A(n6777), .B(n6776), .Z(n6778) );
  NAND U10965 ( .A(n6779), .B(n6778), .Z(n6780) );
  NANDN U10966 ( .A(n6781), .B(n6780), .Z(n6783) );
  OR U10967 ( .A(n6783), .B(n6782), .Z(n6784) );
  AND U10968 ( .A(n6785), .B(n6784), .Z(n6787) );
  NOR U10969 ( .A(n6787), .B(n6786), .Z(n6788) );
  NANDN U10970 ( .A(n6789), .B(n6788), .Z(n6790) );
  AND U10971 ( .A(n6791), .B(n6790), .Z(n6793) );
  NAND U10972 ( .A(n6793), .B(n6792), .Z(n6795) );
  ANDN U10973 ( .B(n6795), .A(n6794), .Z(n6796) );
  NANDN U10974 ( .A(n6797), .B(n6796), .Z(n6801) );
  AND U10975 ( .A(n6799), .B(n6798), .Z(n6800) );
  NAND U10976 ( .A(n6801), .B(n6800), .Z(n6802) );
  NANDN U10977 ( .A(n6803), .B(n6802), .Z(n6805) );
  OR U10978 ( .A(n6805), .B(n6804), .Z(n6806) );
  AND U10979 ( .A(n6807), .B(n6806), .Z(n6809) );
  NOR U10980 ( .A(n6809), .B(n6808), .Z(n6810) );
  NANDN U10981 ( .A(n6811), .B(n6810), .Z(n6812) );
  AND U10982 ( .A(n6813), .B(n6812), .Z(n6815) );
  NAND U10983 ( .A(n6815), .B(n6814), .Z(n6817) );
  ANDN U10984 ( .B(n6817), .A(n6816), .Z(n6818) );
  NANDN U10985 ( .A(n6819), .B(n6818), .Z(n6823) );
  AND U10986 ( .A(n6821), .B(n6820), .Z(n6822) );
  NAND U10987 ( .A(n6823), .B(n6822), .Z(n6824) );
  NANDN U10988 ( .A(n6825), .B(n6824), .Z(n6827) );
  OR U10989 ( .A(n6827), .B(n6826), .Z(n6828) );
  AND U10990 ( .A(n6829), .B(n6828), .Z(n6831) );
  NOR U10991 ( .A(n6831), .B(n6830), .Z(n6832) );
  NANDN U10992 ( .A(n6833), .B(n6832), .Z(n6834) );
  AND U10993 ( .A(n6835), .B(n6834), .Z(n6837) );
  NAND U10994 ( .A(n6837), .B(n6836), .Z(n6839) );
  ANDN U10995 ( .B(n6839), .A(n6838), .Z(n6840) );
  NANDN U10996 ( .A(n6841), .B(n6840), .Z(n6845) );
  AND U10997 ( .A(n6843), .B(n6842), .Z(n6844) );
  NAND U10998 ( .A(n6845), .B(n6844), .Z(n6846) );
  NANDN U10999 ( .A(n6847), .B(n6846), .Z(n6849) );
  OR U11000 ( .A(n6849), .B(n6848), .Z(n6850) );
  AND U11001 ( .A(n6851), .B(n6850), .Z(n6853) );
  NOR U11002 ( .A(n6853), .B(n6852), .Z(n6854) );
  NANDN U11003 ( .A(n6855), .B(n6854), .Z(n6856) );
  AND U11004 ( .A(n6857), .B(n6856), .Z(n6859) );
  NAND U11005 ( .A(n6859), .B(n6858), .Z(n6861) );
  ANDN U11006 ( .B(n6861), .A(n6860), .Z(n6862) );
  NANDN U11007 ( .A(n6863), .B(n6862), .Z(n6867) );
  AND U11008 ( .A(n6865), .B(n6864), .Z(n6866) );
  NAND U11009 ( .A(n6867), .B(n6866), .Z(n6868) );
  NANDN U11010 ( .A(n6869), .B(n6868), .Z(n6871) );
  OR U11011 ( .A(n6871), .B(n6870), .Z(n6872) );
  AND U11012 ( .A(n6873), .B(n6872), .Z(n6875) );
  NOR U11013 ( .A(n6875), .B(n6874), .Z(n6876) );
  NANDN U11014 ( .A(n6877), .B(n6876), .Z(n6878) );
  AND U11015 ( .A(n6879), .B(n6878), .Z(n6881) );
  NAND U11016 ( .A(n6881), .B(n6880), .Z(n6883) );
  ANDN U11017 ( .B(n6883), .A(n6882), .Z(n6884) );
  NANDN U11018 ( .A(n6885), .B(n6884), .Z(n6889) );
  AND U11019 ( .A(n6887), .B(n6886), .Z(n6888) );
  AND U11020 ( .A(n6904), .B(n6903), .Z(n6906) );
  NAND U11021 ( .A(n6906), .B(n6905), .Z(n6908) );
  ANDN U11022 ( .B(n6908), .A(n6907), .Z(n6909) );
  NANDN U11023 ( .A(n6910), .B(n6909), .Z(n6914) );
  AND U11024 ( .A(n6912), .B(n6911), .Z(n6913) );
  NAND U11025 ( .A(n6914), .B(n6913), .Z(n6915) );
  NANDN U11026 ( .A(n6916), .B(n6915), .Z(n6918) );
  OR U11027 ( .A(n6918), .B(n6917), .Z(n6919) );
  AND U11028 ( .A(n6920), .B(n6919), .Z(n6922) );
  NOR U11029 ( .A(n6922), .B(n6921), .Z(n6923) );
  NANDN U11030 ( .A(n6924), .B(n6923), .Z(n6925) );
  AND U11031 ( .A(n6926), .B(n6925), .Z(n6928) );
  NAND U11032 ( .A(n6928), .B(n6927), .Z(n6930) );
  ANDN U11033 ( .B(n6930), .A(n6929), .Z(n6931) );
  NANDN U11034 ( .A(n6932), .B(n6931), .Z(n6936) );
  AND U11035 ( .A(n6934), .B(n6933), .Z(n6935) );
  NAND U11036 ( .A(n6936), .B(n6935), .Z(n6937) );
  NANDN U11037 ( .A(n6938), .B(n6937), .Z(n6940) );
  OR U11038 ( .A(n6940), .B(n6939), .Z(n6941) );
  AND U11039 ( .A(n6942), .B(n6941), .Z(n6944) );
  NOR U11040 ( .A(n6944), .B(n6943), .Z(n6945) );
  NANDN U11041 ( .A(n6946), .B(n6945), .Z(n6947) );
  AND U11042 ( .A(n6948), .B(n6947), .Z(n6950) );
  NAND U11043 ( .A(n6950), .B(n6949), .Z(n6952) );
  ANDN U11044 ( .B(n6952), .A(n6951), .Z(n6953) );
  NANDN U11045 ( .A(n6954), .B(n6953), .Z(n6958) );
  AND U11046 ( .A(n6956), .B(n6955), .Z(n6957) );
  NAND U11047 ( .A(n6958), .B(n6957), .Z(n6959) );
  NANDN U11048 ( .A(n6960), .B(n6959), .Z(n6962) );
  OR U11049 ( .A(n6962), .B(n6961), .Z(n6963) );
  AND U11050 ( .A(n6964), .B(n6963), .Z(n6966) );
  NOR U11051 ( .A(n6966), .B(n6965), .Z(n6967) );
  NANDN U11052 ( .A(n6968), .B(n6967), .Z(n6969) );
  AND U11053 ( .A(n6970), .B(n6969), .Z(n6972) );
  NAND U11054 ( .A(n6972), .B(n6971), .Z(n6974) );
  ANDN U11055 ( .B(n6974), .A(n6973), .Z(n6975) );
  NANDN U11056 ( .A(n6976), .B(n6975), .Z(n6980) );
  AND U11057 ( .A(n6978), .B(n6977), .Z(n6979) );
  NAND U11058 ( .A(n6980), .B(n6979), .Z(n6981) );
  NANDN U11059 ( .A(n6982), .B(n6981), .Z(n6984) );
  OR U11060 ( .A(n6984), .B(n6983), .Z(n6985) );
  AND U11061 ( .A(n6986), .B(n6985), .Z(n6988) );
  NOR U11062 ( .A(n6988), .B(n6987), .Z(n6989) );
  NANDN U11063 ( .A(n6990), .B(n6989), .Z(n6991) );
  AND U11064 ( .A(n6992), .B(n6991), .Z(n6994) );
  NAND U11065 ( .A(n6994), .B(n6993), .Z(n6996) );
  ANDN U11066 ( .B(n6996), .A(n6995), .Z(n6997) );
  NANDN U11067 ( .A(n6998), .B(n6997), .Z(n7002) );
  AND U11068 ( .A(n7000), .B(n6999), .Z(n7001) );
  NAND U11069 ( .A(n7002), .B(n7001), .Z(n7003) );
  NANDN U11070 ( .A(n7004), .B(n7003), .Z(n7006) );
  ANDN U11071 ( .B(x[308]), .A(y[308]), .Z(n7005) );
  OR U11072 ( .A(n7006), .B(n7005), .Z(n7007) );
  AND U11073 ( .A(n7008), .B(n7007), .Z(n7010) );
  NOR U11074 ( .A(n7010), .B(n7009), .Z(n7011) );
  NANDN U11075 ( .A(n7012), .B(n7011), .Z(n7013) );
  AND U11076 ( .A(n7014), .B(n7013), .Z(n7016) );
  NAND U11077 ( .A(n7016), .B(n7015), .Z(n7018) );
  ANDN U11078 ( .B(n7018), .A(n7017), .Z(n7019) );
  NANDN U11079 ( .A(n7020), .B(n7019), .Z(n7024) );
  AND U11080 ( .A(n7022), .B(n7021), .Z(n7023) );
  NAND U11081 ( .A(n7024), .B(n7023), .Z(n7025) );
  NANDN U11082 ( .A(n7026), .B(n7025), .Z(n7028) );
  OR U11083 ( .A(n7028), .B(n7027), .Z(n7029) );
  AND U11084 ( .A(n7030), .B(n7029), .Z(n7032) );
  NOR U11085 ( .A(n7032), .B(n7031), .Z(n7033) );
  NANDN U11086 ( .A(n7034), .B(n7033), .Z(n7035) );
  AND U11087 ( .A(n7036), .B(n7035), .Z(n7038) );
  NAND U11088 ( .A(n7038), .B(n7037), .Z(n7040) );
  ANDN U11089 ( .B(x[318]), .A(y[318]), .Z(n7039) );
  ANDN U11090 ( .B(n7040), .A(n7039), .Z(n7041) );
  NANDN U11091 ( .A(n7042), .B(n7041), .Z(n7046) );
  AND U11092 ( .A(n7044), .B(n7043), .Z(n7045) );
  NAND U11093 ( .A(n7046), .B(n7045), .Z(n7047) );
  NANDN U11094 ( .A(n7048), .B(n7047), .Z(n7050) );
  OR U11095 ( .A(n7050), .B(n7049), .Z(n7051) );
  AND U11096 ( .A(n7052), .B(n7051), .Z(n7054) );
  NOR U11097 ( .A(n7054), .B(n7053), .Z(n7055) );
  NANDN U11098 ( .A(n7056), .B(n7055), .Z(n7057) );
  AND U11099 ( .A(n7058), .B(n7057), .Z(n7060) );
  NAND U11100 ( .A(n7060), .B(n7059), .Z(n7062) );
  ANDN U11101 ( .B(n7062), .A(n7061), .Z(n7063) );
  NANDN U11102 ( .A(n7064), .B(n7063), .Z(n7068) );
  AND U11103 ( .A(n7066), .B(n7065), .Z(n7067) );
  NAND U11104 ( .A(n7068), .B(n7067), .Z(n7069) );
  NANDN U11105 ( .A(n7070), .B(n7069), .Z(n7072) );
  OR U11106 ( .A(n7072), .B(n7071), .Z(n7073) );
  AND U11107 ( .A(n7074), .B(n7073), .Z(n7076) );
  NOR U11108 ( .A(n7076), .B(n7075), .Z(n7077) );
  NANDN U11109 ( .A(n7078), .B(n7077), .Z(n7079) );
  AND U11110 ( .A(n7080), .B(n7079), .Z(n7082) );
  NAND U11111 ( .A(n7082), .B(n7081), .Z(n7084) );
  ANDN U11112 ( .B(n7084), .A(n7083), .Z(n7085) );
  NANDN U11113 ( .A(n7086), .B(n7085), .Z(n7090) );
  AND U11114 ( .A(n7088), .B(n7087), .Z(n7089) );
  NAND U11115 ( .A(n7090), .B(n7089), .Z(n7091) );
  NANDN U11116 ( .A(n7092), .B(n7091), .Z(n7094) );
  ANDN U11117 ( .B(x[332]), .A(y[332]), .Z(n7093) );
  OR U11118 ( .A(n7094), .B(n7093), .Z(n7095) );
  AND U11119 ( .A(n7096), .B(n7095), .Z(n7098) );
  NOR U11120 ( .A(n7098), .B(n7097), .Z(n7099) );
  NANDN U11121 ( .A(n7100), .B(n7099), .Z(n7101) );
  AND U11122 ( .A(n7102), .B(n7101), .Z(n7104) );
  NAND U11123 ( .A(n7104), .B(n7103), .Z(n7106) );
  ANDN U11124 ( .B(n7106), .A(n7105), .Z(n7107) );
  NANDN U11125 ( .A(n7108), .B(n7107), .Z(n7112) );
  AND U11126 ( .A(n7110), .B(n7109), .Z(n7111) );
  NAND U11127 ( .A(n7112), .B(n7111), .Z(n7113) );
  NANDN U11128 ( .A(n7114), .B(n7113), .Z(n7116) );
  OR U11129 ( .A(n7116), .B(n7115), .Z(n7117) );
  AND U11130 ( .A(n7118), .B(n7117), .Z(n7120) );
  NOR U11131 ( .A(n7120), .B(n7119), .Z(n7121) );
  NANDN U11132 ( .A(n7122), .B(n7121), .Z(n7123) );
  AND U11133 ( .A(n7124), .B(n7123), .Z(n7126) );
  NAND U11134 ( .A(n7126), .B(n7125), .Z(n7128) );
  ANDN U11135 ( .B(n7128), .A(n7127), .Z(n7129) );
  NANDN U11136 ( .A(n7130), .B(n7129), .Z(n7134) );
  AND U11137 ( .A(n7132), .B(n7131), .Z(n7133) );
  NAND U11138 ( .A(n7134), .B(n7133), .Z(n7135) );
  NANDN U11139 ( .A(n7136), .B(n7135), .Z(n7138) );
  OR U11140 ( .A(n7138), .B(n7137), .Z(n7139) );
  AND U11141 ( .A(n7140), .B(n7139), .Z(n7142) );
  NOR U11142 ( .A(n7142), .B(n7141), .Z(n7143) );
  NANDN U11143 ( .A(n7144), .B(n7143), .Z(n7145) );
  AND U11144 ( .A(n7146), .B(n7145), .Z(n7148) );
  NAND U11145 ( .A(n7148), .B(n7147), .Z(n7150) );
  ANDN U11146 ( .B(n7150), .A(n7149), .Z(n7151) );
  NANDN U11147 ( .A(n7152), .B(n7151), .Z(n7156) );
  AND U11148 ( .A(n7154), .B(n7153), .Z(n7155) );
  NAND U11149 ( .A(n7156), .B(n7155), .Z(n7157) );
  NANDN U11150 ( .A(n7158), .B(n7157), .Z(n7160) );
  OR U11151 ( .A(n7160), .B(n7159), .Z(n7161) );
  AND U11152 ( .A(n7162), .B(n7161), .Z(n7164) );
  NOR U11153 ( .A(n7164), .B(n7163), .Z(n7165) );
  NANDN U11154 ( .A(n7166), .B(n7165), .Z(n7167) );
  AND U11155 ( .A(n7168), .B(n7167), .Z(n7170) );
  NAND U11156 ( .A(n7170), .B(n7169), .Z(n7172) );
  ANDN U11157 ( .B(n7172), .A(n7171), .Z(n7173) );
  NANDN U11158 ( .A(n7174), .B(n7173), .Z(n7178) );
  AND U11159 ( .A(n7176), .B(n7175), .Z(n7177) );
  NAND U11160 ( .A(n7178), .B(n7177), .Z(n7179) );
  NANDN U11161 ( .A(n7180), .B(n7179), .Z(n7182) );
  OR U11162 ( .A(n7182), .B(n7181), .Z(n7183) );
  AND U11163 ( .A(n7184), .B(n7183), .Z(n7186) );
  NOR U11164 ( .A(n7186), .B(n7185), .Z(n7187) );
  NANDN U11165 ( .A(n7188), .B(n7187), .Z(n7189) );
  AND U11166 ( .A(n7190), .B(n7189), .Z(n7192) );
  NAND U11167 ( .A(n7192), .B(n7191), .Z(n7194) );
  ANDN U11168 ( .B(n7194), .A(n7193), .Z(n7195) );
  NANDN U11169 ( .A(n7196), .B(n7195), .Z(n7200) );
  AND U11170 ( .A(n7198), .B(n7197), .Z(n7199) );
  NAND U11171 ( .A(n7200), .B(n7199), .Z(n7201) );
  NANDN U11172 ( .A(n7202), .B(n7201), .Z(n7204) );
  OR U11173 ( .A(n7204), .B(n7203), .Z(n7205) );
  AND U11174 ( .A(n7206), .B(n7205), .Z(n7208) );
  NOR U11175 ( .A(n7208), .B(n7207), .Z(n7209) );
  NANDN U11176 ( .A(n7210), .B(n7209), .Z(n7211) );
  AND U11177 ( .A(n7212), .B(n7211), .Z(n7214) );
  NAND U11178 ( .A(n7214), .B(n7213), .Z(n7216) );
  ANDN U11179 ( .B(n7216), .A(n7215), .Z(n7217) );
  NANDN U11180 ( .A(n7218), .B(n7217), .Z(n7222) );
  AND U11181 ( .A(n7220), .B(n7219), .Z(n7221) );
  NAND U11182 ( .A(n7222), .B(n7221), .Z(n7223) );
  NANDN U11183 ( .A(n7224), .B(n7223), .Z(n7226) );
  ANDN U11184 ( .B(x[368]), .A(y[368]), .Z(n7225) );
  OR U11185 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U11186 ( .A(n7228), .B(n7227), .Z(n7230) );
  NOR U11187 ( .A(n7230), .B(n7229), .Z(n7231) );
  NANDN U11188 ( .A(n7232), .B(n7231), .Z(n7233) );
  AND U11189 ( .A(n7234), .B(n7233), .Z(n7236) );
  NAND U11190 ( .A(n7236), .B(n7235), .Z(n7238) );
  ANDN U11191 ( .B(n7238), .A(n7237), .Z(n7239) );
  NANDN U11192 ( .A(n7240), .B(n7239), .Z(n7244) );
  AND U11193 ( .A(n7242), .B(n7241), .Z(n7243) );
  NAND U11194 ( .A(n7244), .B(n7243), .Z(n7245) );
  NANDN U11195 ( .A(n7246), .B(n7245), .Z(n7248) );
  OR U11196 ( .A(n7248), .B(n7247), .Z(n7249) );
  AND U11197 ( .A(n7250), .B(n7249), .Z(n7252) );
  NOR U11198 ( .A(n7252), .B(n7251), .Z(n7253) );
  NANDN U11199 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U11200 ( .A(n7256), .B(n7255), .Z(n7257) );
  NAND U11201 ( .A(n7258), .B(n7257), .Z(n7259) );
  NAND U11202 ( .A(n7260), .B(n7259), .Z(n7261) );
  AND U11203 ( .A(n7262), .B(n7261), .Z(n7263) );
  OR U11204 ( .A(n7263), .B(n10941), .Z(n7264) );
  NAND U11205 ( .A(n10943), .B(n7264), .Z(n7265) );
  NANDN U11206 ( .A(n7266), .B(n7265), .Z(n7268) );
  NAND U11207 ( .A(n7268), .B(n7267), .Z(n7270) );
  ANDN U11208 ( .B(n7270), .A(n7269), .Z(n7271) );
  NANDN U11209 ( .A(n7272), .B(n7271), .Z(n7274) );
  NAND U11210 ( .A(n7274), .B(n7273), .Z(n7275) );
  NANDN U11211 ( .A(n7276), .B(n7275), .Z(n7277) );
  AND U11212 ( .A(n10951), .B(n7277), .Z(n7278) );
  OR U11213 ( .A(n10953), .B(n7278), .Z(n7279) );
  NAND U11214 ( .A(n10955), .B(n7279), .Z(n7280) );
  NANDN U11215 ( .A(n10957), .B(n7280), .Z(n7281) );
  NAND U11216 ( .A(n10959), .B(n7281), .Z(n7282) );
  NANDN U11217 ( .A(n7283), .B(n7282), .Z(n7284) );
  AND U11218 ( .A(n7285), .B(n7284), .Z(n7287) );
  NOR U11219 ( .A(n7287), .B(n7286), .Z(n7288) );
  NANDN U11220 ( .A(n7289), .B(n7288), .Z(n7290) );
  AND U11221 ( .A(n7291), .B(n7290), .Z(n7293) );
  NAND U11222 ( .A(n7293), .B(n7292), .Z(n7295) );
  ANDN U11223 ( .B(n7295), .A(n7294), .Z(n7296) );
  NANDN U11224 ( .A(n7297), .B(n7296), .Z(n7301) );
  AND U11225 ( .A(n7299), .B(n7298), .Z(n7300) );
  NAND U11226 ( .A(n7301), .B(n7300), .Z(n7302) );
  NANDN U11227 ( .A(n7303), .B(n7302), .Z(n7305) );
  OR U11228 ( .A(n7305), .B(n7304), .Z(n7306) );
  AND U11229 ( .A(n7307), .B(n7306), .Z(n7309) );
  NOR U11230 ( .A(n7309), .B(n7308), .Z(n7310) );
  NANDN U11231 ( .A(n7311), .B(n7310), .Z(n7312) );
  AND U11232 ( .A(n7313), .B(n7312), .Z(n7315) );
  NAND U11233 ( .A(n7315), .B(n7314), .Z(n7317) );
  ANDN U11234 ( .B(n7317), .A(n7316), .Z(n7318) );
  NANDN U11235 ( .A(n7319), .B(n7318), .Z(n7323) );
  AND U11236 ( .A(n7321), .B(n7320), .Z(n7322) );
  NAND U11237 ( .A(n7323), .B(n7322), .Z(n7324) );
  NANDN U11238 ( .A(n7325), .B(n7324), .Z(n7327) );
  OR U11239 ( .A(n7327), .B(n7326), .Z(n7328) );
  AND U11240 ( .A(n7329), .B(n7328), .Z(n7331) );
  NOR U11241 ( .A(n7331), .B(n7330), .Z(n7332) );
  NANDN U11242 ( .A(n7333), .B(n7332), .Z(n7334) );
  AND U11243 ( .A(n7335), .B(n7334), .Z(n7337) );
  NAND U11244 ( .A(n7337), .B(n7336), .Z(n7339) );
  ANDN U11245 ( .B(n7339), .A(n7338), .Z(n7340) );
  NANDN U11246 ( .A(n7341), .B(n7340), .Z(n7345) );
  AND U11247 ( .A(n7343), .B(n7342), .Z(n7344) );
  NAND U11248 ( .A(n7345), .B(n7344), .Z(n7346) );
  NANDN U11249 ( .A(n7347), .B(n7346), .Z(n7349) );
  OR U11250 ( .A(n7349), .B(n7348), .Z(n7350) );
  AND U11251 ( .A(n7351), .B(n7350), .Z(n7353) );
  NOR U11252 ( .A(n7353), .B(n7352), .Z(n7354) );
  NANDN U11253 ( .A(n7355), .B(n7354), .Z(n7356) );
  AND U11254 ( .A(n7357), .B(n7356), .Z(n7359) );
  NAND U11255 ( .A(n7359), .B(n7358), .Z(n7361) );
  ANDN U11256 ( .B(n7361), .A(n7360), .Z(n7362) );
  NANDN U11257 ( .A(n7363), .B(n7362), .Z(n7367) );
  AND U11258 ( .A(n7365), .B(n7364), .Z(n7366) );
  NAND U11259 ( .A(n7367), .B(n7366), .Z(n7368) );
  NANDN U11260 ( .A(n7369), .B(n7368), .Z(n7371) );
  OR U11261 ( .A(n7371), .B(n7370), .Z(n7372) );
  AND U11262 ( .A(n7373), .B(n7372), .Z(n7375) );
  NOR U11263 ( .A(n7375), .B(n7374), .Z(n7376) );
  NANDN U11264 ( .A(n7377), .B(n7376), .Z(n7378) );
  AND U11265 ( .A(n7379), .B(n7378), .Z(n7380) );
  OR U11266 ( .A(n7381), .B(n7380), .Z(n7382) );
  NAND U11267 ( .A(n7383), .B(n7382), .Z(n7384) );
  NANDN U11268 ( .A(n7385), .B(n7384), .Z(n7389) );
  AND U11269 ( .A(n7387), .B(n7386), .Z(n7388) );
  NAND U11270 ( .A(n7389), .B(n7388), .Z(n7390) );
  NANDN U11271 ( .A(n7391), .B(n7390), .Z(n7393) );
  OR U11272 ( .A(n7393), .B(n7392), .Z(n7394) );
  AND U11273 ( .A(n7395), .B(n7394), .Z(n7397) );
  NOR U11274 ( .A(n7397), .B(n7396), .Z(n7398) );
  NANDN U11275 ( .A(n7399), .B(n7398), .Z(n7400) );
  AND U11276 ( .A(n7401), .B(n7400), .Z(n7403) );
  NAND U11277 ( .A(n7403), .B(n7402), .Z(n7405) );
  ANDN U11278 ( .B(n7405), .A(n7404), .Z(n7406) );
  NANDN U11279 ( .A(n7407), .B(n7406), .Z(n7411) );
  AND U11280 ( .A(n7409), .B(n7408), .Z(n7410) );
  NAND U11281 ( .A(n7411), .B(n7410), .Z(n7412) );
  NANDN U11282 ( .A(n7413), .B(n7412), .Z(n7415) );
  OR U11283 ( .A(n7415), .B(n7414), .Z(n7416) );
  AND U11284 ( .A(n7417), .B(n7416), .Z(n7419) );
  NOR U11285 ( .A(n7419), .B(n7418), .Z(n7420) );
  NANDN U11286 ( .A(n7421), .B(n7420), .Z(n7422) );
  AND U11287 ( .A(n7423), .B(n7422), .Z(n7425) );
  NAND U11288 ( .A(n7425), .B(n7424), .Z(n7427) );
  ANDN U11289 ( .B(n7427), .A(n7426), .Z(n7428) );
  NANDN U11290 ( .A(n7429), .B(n7428), .Z(n7433) );
  AND U11291 ( .A(n7431), .B(n7430), .Z(n7432) );
  NAND U11292 ( .A(n7433), .B(n7432), .Z(n7434) );
  NANDN U11293 ( .A(n7435), .B(n7434), .Z(n7437) );
  OR U11294 ( .A(n7437), .B(n7436), .Z(n7438) );
  AND U11295 ( .A(n7439), .B(n7438), .Z(n7441) );
  NOR U11296 ( .A(n7441), .B(n7440), .Z(n7442) );
  NANDN U11297 ( .A(n7443), .B(n7442), .Z(n7444) );
  AND U11298 ( .A(n7445), .B(n7444), .Z(n7447) );
  NAND U11299 ( .A(n7447), .B(n7446), .Z(n7449) );
  ANDN U11300 ( .B(x[434]), .A(y[434]), .Z(n7448) );
  ANDN U11301 ( .B(n7449), .A(n7448), .Z(n7450) );
  NANDN U11302 ( .A(n7451), .B(n7450), .Z(n7455) );
  AND U11303 ( .A(n7453), .B(n7452), .Z(n7454) );
  NAND U11304 ( .A(n7455), .B(n7454), .Z(n7456) );
  NANDN U11305 ( .A(n7457), .B(n7456), .Z(n7459) );
  OR U11306 ( .A(n7459), .B(n7458), .Z(n7460) );
  AND U11307 ( .A(n7461), .B(n7460), .Z(n7463) );
  NOR U11308 ( .A(n7463), .B(n7462), .Z(n7464) );
  NANDN U11309 ( .A(n7465), .B(n7464), .Z(n7466) );
  AND U11310 ( .A(n7467), .B(n7466), .Z(n7469) );
  NAND U11311 ( .A(n7469), .B(n7468), .Z(n7471) );
  ANDN U11312 ( .B(n7471), .A(n7470), .Z(n7472) );
  NANDN U11313 ( .A(n7473), .B(n7472), .Z(n7477) );
  AND U11314 ( .A(n7475), .B(n7474), .Z(n7476) );
  NAND U11315 ( .A(n7477), .B(n7476), .Z(n7478) );
  NANDN U11316 ( .A(n7479), .B(n7478), .Z(n7481) );
  OR U11317 ( .A(n7481), .B(n7480), .Z(n7482) );
  AND U11318 ( .A(n7483), .B(n7482), .Z(n7485) );
  NOR U11319 ( .A(n7485), .B(n7484), .Z(n7486) );
  NANDN U11320 ( .A(n7487), .B(n7486), .Z(n7488) );
  AND U11321 ( .A(n7489), .B(n7488), .Z(n7491) );
  NAND U11322 ( .A(n7491), .B(n7490), .Z(n7493) );
  ANDN U11323 ( .B(n7493), .A(n7492), .Z(n7494) );
  NANDN U11324 ( .A(n7495), .B(n7494), .Z(n7499) );
  AND U11325 ( .A(n7497), .B(n7496), .Z(n7498) );
  NAND U11326 ( .A(n7499), .B(n7498), .Z(n7500) );
  NANDN U11327 ( .A(n7501), .B(n7500), .Z(n7503) );
  OR U11328 ( .A(n7503), .B(n7502), .Z(n7504) );
  AND U11329 ( .A(n7505), .B(n7504), .Z(n7507) );
  NOR U11330 ( .A(n7507), .B(n7506), .Z(n7508) );
  NANDN U11331 ( .A(n7509), .B(n7508), .Z(n7510) );
  AND U11332 ( .A(n7511), .B(n7510), .Z(n7513) );
  NAND U11333 ( .A(n7513), .B(n7512), .Z(n7515) );
  ANDN U11334 ( .B(n7515), .A(n7514), .Z(n7516) );
  NANDN U11335 ( .A(n7517), .B(n7516), .Z(n7521) );
  AND U11336 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U11337 ( .A(n7521), .B(n7520), .Z(n7522) );
  NANDN U11338 ( .A(n7523), .B(n7522), .Z(n7525) );
  OR U11339 ( .A(n7525), .B(n7524), .Z(n7526) );
  AND U11340 ( .A(n7527), .B(n7526), .Z(n7529) );
  ANDN U11341 ( .B(x[456]), .A(y[456]), .Z(n7528) );
  NOR U11342 ( .A(n7529), .B(n7528), .Z(n7530) );
  NANDN U11343 ( .A(n7531), .B(n7530), .Z(n7532) );
  AND U11344 ( .A(n7533), .B(n7532), .Z(n7535) );
  NAND U11345 ( .A(n7535), .B(n7534), .Z(n7537) );
  ANDN U11346 ( .B(n7537), .A(n7536), .Z(n7538) );
  NANDN U11347 ( .A(n7539), .B(n7538), .Z(n7543) );
  AND U11348 ( .A(n7541), .B(n7540), .Z(n7542) );
  NAND U11349 ( .A(n7543), .B(n7542), .Z(n7544) );
  NANDN U11350 ( .A(n7545), .B(n7544), .Z(n7547) );
  OR U11351 ( .A(n7547), .B(n7546), .Z(n7548) );
  AND U11352 ( .A(n7549), .B(n7548), .Z(n7551) );
  ANDN U11353 ( .B(x[462]), .A(y[462]), .Z(n7550) );
  NOR U11354 ( .A(n7551), .B(n7550), .Z(n7552) );
  NANDN U11355 ( .A(n7553), .B(n7552), .Z(n7554) );
  AND U11356 ( .A(n7555), .B(n7554), .Z(n7557) );
  NAND U11357 ( .A(n7557), .B(n7556), .Z(n7559) );
  ANDN U11358 ( .B(n7559), .A(n7558), .Z(n7560) );
  NANDN U11359 ( .A(n7561), .B(n7560), .Z(n7565) );
  AND U11360 ( .A(n7563), .B(n7562), .Z(n7564) );
  NAND U11361 ( .A(n7565), .B(n7564), .Z(n7566) );
  NANDN U11362 ( .A(n7567), .B(n7566), .Z(n7569) );
  OR U11363 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U11364 ( .A(n7571), .B(n7570), .Z(n7573) );
  ANDN U11365 ( .B(x[468]), .A(y[468]), .Z(n7572) );
  NOR U11366 ( .A(n7573), .B(n7572), .Z(n7574) );
  NANDN U11367 ( .A(n7575), .B(n7574), .Z(n7576) );
  AND U11368 ( .A(n7577), .B(n7576), .Z(n7579) );
  NAND U11369 ( .A(n7579), .B(n7578), .Z(n7581) );
  ANDN U11370 ( .B(n7581), .A(n7580), .Z(n7582) );
  NANDN U11371 ( .A(n7583), .B(n7582), .Z(n7587) );
  AND U11372 ( .A(n7585), .B(n7584), .Z(n7586) );
  NAND U11373 ( .A(n7587), .B(n7586), .Z(n7588) );
  NANDN U11374 ( .A(n7589), .B(n7588), .Z(n7591) );
  OR U11375 ( .A(n7591), .B(n7590), .Z(n7592) );
  AND U11376 ( .A(n7593), .B(n7592), .Z(n7595) );
  NOR U11377 ( .A(n7595), .B(n7594), .Z(n7596) );
  NANDN U11378 ( .A(n7597), .B(n7596), .Z(n7598) );
  AND U11379 ( .A(n7599), .B(n7598), .Z(n7601) );
  NAND U11380 ( .A(n7601), .B(n7600), .Z(n7603) );
  ANDN U11381 ( .B(n7603), .A(n7602), .Z(n7604) );
  NANDN U11382 ( .A(n7605), .B(n7604), .Z(n7609) );
  AND U11383 ( .A(n7607), .B(n7606), .Z(n7608) );
  NAND U11384 ( .A(n7609), .B(n7608), .Z(n7610) );
  NANDN U11385 ( .A(n7611), .B(n7610), .Z(n7613) );
  OR U11386 ( .A(n7613), .B(n7612), .Z(n7614) );
  AND U11387 ( .A(n7615), .B(n7614), .Z(n7617) );
  ANDN U11388 ( .B(x[480]), .A(y[480]), .Z(n7616) );
  NOR U11389 ( .A(n7617), .B(n7616), .Z(n7618) );
  NANDN U11390 ( .A(n7619), .B(n7618), .Z(n7620) );
  AND U11391 ( .A(n7621), .B(n7620), .Z(n7623) );
  NAND U11392 ( .A(n7623), .B(n7622), .Z(n7625) );
  ANDN U11393 ( .B(n7625), .A(n7624), .Z(n7626) );
  NANDN U11394 ( .A(n7627), .B(n7626), .Z(n7631) );
  AND U11395 ( .A(n7629), .B(n7628), .Z(n7630) );
  NAND U11396 ( .A(n7631), .B(n7630), .Z(n7632) );
  NANDN U11397 ( .A(n7633), .B(n7632), .Z(n7635) );
  OR U11398 ( .A(n7635), .B(n7634), .Z(n7636) );
  AND U11399 ( .A(n7637), .B(n7636), .Z(n7639) );
  NOR U11400 ( .A(n7639), .B(n7638), .Z(n7640) );
  NANDN U11401 ( .A(n7641), .B(n7640), .Z(n7642) );
  AND U11402 ( .A(n7643), .B(n7642), .Z(n7645) );
  NAND U11403 ( .A(n7645), .B(n7644), .Z(n7647) );
  ANDN U11404 ( .B(n7647), .A(n7646), .Z(n7648) );
  NANDN U11405 ( .A(n7649), .B(n7648), .Z(n7653) );
  AND U11406 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U11407 ( .A(n7653), .B(n7652), .Z(n7654) );
  NANDN U11408 ( .A(n7655), .B(n7654), .Z(n7657) );
  OR U11409 ( .A(n7657), .B(n7656), .Z(n7658) );
  AND U11410 ( .A(n7659), .B(n7658), .Z(n7661) );
  NOR U11411 ( .A(n7661), .B(n7660), .Z(n7662) );
  NANDN U11412 ( .A(n7663), .B(n7662), .Z(n7664) );
  AND U11413 ( .A(n7665), .B(n7664), .Z(n7667) );
  NAND U11414 ( .A(n7667), .B(n7666), .Z(n7669) );
  ANDN U11415 ( .B(n7669), .A(n7668), .Z(n7670) );
  NANDN U11416 ( .A(n7671), .B(n7670), .Z(n7675) );
  AND U11417 ( .A(n7673), .B(n7672), .Z(n7674) );
  NAND U11418 ( .A(n7675), .B(n7674), .Z(n7676) );
  NANDN U11419 ( .A(n7677), .B(n7676), .Z(n7679) );
  OR U11420 ( .A(n7679), .B(n7678), .Z(n7680) );
  AND U11421 ( .A(n7681), .B(n7680), .Z(n7683) );
  NOR U11422 ( .A(n7683), .B(n7682), .Z(n7684) );
  NANDN U11423 ( .A(n7685), .B(n7684), .Z(n7686) );
  AND U11424 ( .A(n7687), .B(n7686), .Z(n7689) );
  NAND U11425 ( .A(n7689), .B(n7688), .Z(n7691) );
  ANDN U11426 ( .B(n7691), .A(n7690), .Z(n7692) );
  NANDN U11427 ( .A(n7693), .B(n7692), .Z(n7697) );
  AND U11428 ( .A(n7695), .B(n7694), .Z(n7696) );
  NAND U11429 ( .A(n7697), .B(n7696), .Z(n7698) );
  NANDN U11430 ( .A(n7699), .B(n7698), .Z(n7701) );
  OR U11431 ( .A(n7701), .B(n7700), .Z(n7702) );
  AND U11432 ( .A(n7703), .B(n7702), .Z(n7705) );
  NOR U11433 ( .A(n7705), .B(n7704), .Z(n7706) );
  NANDN U11434 ( .A(n7707), .B(n7706), .Z(n7708) );
  AND U11435 ( .A(n7709), .B(n7708), .Z(n7711) );
  NAND U11436 ( .A(n7711), .B(n7710), .Z(n7713) );
  ANDN U11437 ( .B(n7713), .A(n7712), .Z(n7714) );
  NANDN U11438 ( .A(n7715), .B(n7714), .Z(n7719) );
  AND U11439 ( .A(n7717), .B(n7716), .Z(n7718) );
  NAND U11440 ( .A(n7719), .B(n7718), .Z(n7720) );
  NANDN U11441 ( .A(n7721), .B(n7720), .Z(n7723) );
  OR U11442 ( .A(n7723), .B(n7722), .Z(n7724) );
  AND U11443 ( .A(n7725), .B(n7724), .Z(n7727) );
  NOR U11444 ( .A(n7727), .B(n7726), .Z(n7728) );
  NANDN U11445 ( .A(n7729), .B(n7728), .Z(n7730) );
  AND U11446 ( .A(n7731), .B(n7730), .Z(n7733) );
  NAND U11447 ( .A(n7733), .B(n7732), .Z(n7735) );
  ANDN U11448 ( .B(n7735), .A(n7734), .Z(n7736) );
  NANDN U11449 ( .A(n7737), .B(n7736), .Z(n7741) );
  AND U11450 ( .A(n7739), .B(n7738), .Z(n7740) );
  NAND U11451 ( .A(n7741), .B(n7740), .Z(n7742) );
  NANDN U11452 ( .A(n7743), .B(n7742), .Z(n7745) );
  OR U11453 ( .A(n7745), .B(n7744), .Z(n7746) );
  AND U11454 ( .A(n7747), .B(n7746), .Z(n7749) );
  NOR U11455 ( .A(n7749), .B(n7748), .Z(n7750) );
  NANDN U11456 ( .A(n7751), .B(n7750), .Z(n7752) );
  AND U11457 ( .A(n7753), .B(n7752), .Z(n7755) );
  NAND U11458 ( .A(n7755), .B(n7754), .Z(n7757) );
  ANDN U11459 ( .B(n7757), .A(n7756), .Z(n7758) );
  NANDN U11460 ( .A(n7759), .B(n7758), .Z(n7763) );
  AND U11461 ( .A(n7761), .B(n7760), .Z(n7762) );
  NAND U11462 ( .A(n7763), .B(n7762), .Z(n7764) );
  NANDN U11463 ( .A(n7765), .B(n7764), .Z(n7767) );
  OR U11464 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U11465 ( .A(n7769), .B(n7768), .Z(n7771) );
  NOR U11466 ( .A(n7771), .B(n7770), .Z(n7772) );
  NANDN U11467 ( .A(n7773), .B(n7772), .Z(n7774) );
  AND U11468 ( .A(n7775), .B(n7774), .Z(n7777) );
  NAND U11469 ( .A(n7777), .B(n7776), .Z(n7779) );
  ANDN U11470 ( .B(n7779), .A(n7778), .Z(n7780) );
  NANDN U11471 ( .A(n7781), .B(n7780), .Z(n7785) );
  AND U11472 ( .A(n7783), .B(n7782), .Z(n7784) );
  NAND U11473 ( .A(n7785), .B(n7784), .Z(n7786) );
  NANDN U11474 ( .A(n7787), .B(n7786), .Z(n7789) );
  OR U11475 ( .A(n7789), .B(n7788), .Z(n7790) );
  AND U11476 ( .A(n7791), .B(n7790), .Z(n7793) );
  NOR U11477 ( .A(n7793), .B(n7792), .Z(n7794) );
  NANDN U11478 ( .A(n7795), .B(n7794), .Z(n7796) );
  AND U11479 ( .A(n7797), .B(n7796), .Z(n7799) );
  NAND U11480 ( .A(n7799), .B(n7798), .Z(n7801) );
  ANDN U11481 ( .B(n7801), .A(n7800), .Z(n7802) );
  NANDN U11482 ( .A(n7803), .B(n7802), .Z(n7807) );
  AND U11483 ( .A(n7805), .B(n7804), .Z(n7806) );
  NAND U11484 ( .A(n7807), .B(n7806), .Z(n7808) );
  NANDN U11485 ( .A(n7809), .B(n7808), .Z(n7811) );
  OR U11486 ( .A(n7811), .B(n7810), .Z(n7812) );
  AND U11487 ( .A(n7813), .B(n7812), .Z(n7814) );
  NOR U11488 ( .A(n7815), .B(n7814), .Z(n7816) );
  NANDN U11489 ( .A(n7817), .B(n7816), .Z(n7818) );
  AND U11490 ( .A(n7819), .B(n7818), .Z(n7821) );
  NAND U11491 ( .A(n7821), .B(n7820), .Z(n7823) );
  ANDN U11492 ( .B(n7823), .A(n7822), .Z(n7824) );
  NANDN U11493 ( .A(n7825), .B(n7824), .Z(n7829) );
  AND U11494 ( .A(n7827), .B(n7826), .Z(n7828) );
  NAND U11495 ( .A(n7829), .B(n7828), .Z(n7830) );
  NANDN U11496 ( .A(n7831), .B(n7830), .Z(n7833) );
  OR U11497 ( .A(n7833), .B(n7832), .Z(n7834) );
  AND U11498 ( .A(n7835), .B(n7834), .Z(n7837) );
  NOR U11499 ( .A(n7837), .B(n7836), .Z(n7838) );
  NANDN U11500 ( .A(n7839), .B(n7838), .Z(n7840) );
  AND U11501 ( .A(n7841), .B(n7840), .Z(n7843) );
  NAND U11502 ( .A(n7843), .B(n7842), .Z(n7845) );
  ANDN U11503 ( .B(n7845), .A(n7844), .Z(n7846) );
  NANDN U11504 ( .A(n7847), .B(n7846), .Z(n7851) );
  AND U11505 ( .A(n7849), .B(n7848), .Z(n7850) );
  NAND U11506 ( .A(n7851), .B(n7850), .Z(n7852) );
  NANDN U11507 ( .A(n7853), .B(n7852), .Z(n7855) );
  OR U11508 ( .A(n7855), .B(n7854), .Z(n7856) );
  AND U11509 ( .A(n7857), .B(n7856), .Z(n7859) );
  NOR U11510 ( .A(n7859), .B(n7858), .Z(n7860) );
  NANDN U11511 ( .A(n7861), .B(n7860), .Z(n7862) );
  AND U11512 ( .A(n7863), .B(n7862), .Z(n7865) );
  NAND U11513 ( .A(n7865), .B(n7864), .Z(n7867) );
  ANDN U11514 ( .B(n7867), .A(n7866), .Z(n7868) );
  NANDN U11515 ( .A(n7869), .B(n7868), .Z(n7873) );
  AND U11516 ( .A(n7871), .B(n7870), .Z(n7872) );
  NAND U11517 ( .A(n7873), .B(n7872), .Z(n7874) );
  NANDN U11518 ( .A(n7875), .B(n7874), .Z(n7877) );
  OR U11519 ( .A(n7877), .B(n7876), .Z(n7878) );
  AND U11520 ( .A(n7879), .B(n7878), .Z(n7881) );
  NOR U11521 ( .A(n7881), .B(n7880), .Z(n7882) );
  NANDN U11522 ( .A(n7883), .B(n7882), .Z(n7884) );
  AND U11523 ( .A(n7885), .B(n7884), .Z(n7887) );
  NAND U11524 ( .A(n7887), .B(n7886), .Z(n7889) );
  ANDN U11525 ( .B(n7889), .A(n7888), .Z(n7890) );
  NANDN U11526 ( .A(n7891), .B(n7890), .Z(n7895) );
  AND U11527 ( .A(n7893), .B(n7892), .Z(n7894) );
  NAND U11528 ( .A(n7895), .B(n7894), .Z(n7896) );
  NANDN U11529 ( .A(n7897), .B(n7896), .Z(n7899) );
  OR U11530 ( .A(n7899), .B(n7898), .Z(n7900) );
  AND U11531 ( .A(n7901), .B(n7900), .Z(n7903) );
  NOR U11532 ( .A(n7903), .B(n7902), .Z(n7904) );
  NANDN U11533 ( .A(n7905), .B(n7904), .Z(n7906) );
  AND U11534 ( .A(n7907), .B(n7906), .Z(n7909) );
  NAND U11535 ( .A(n7909), .B(n7908), .Z(n7911) );
  ANDN U11536 ( .B(n7911), .A(n7910), .Z(n7912) );
  NANDN U11537 ( .A(n7913), .B(n7912), .Z(n7917) );
  AND U11538 ( .A(n7915), .B(n7914), .Z(n7916) );
  NAND U11539 ( .A(n7917), .B(n7916), .Z(n7918) );
  NANDN U11540 ( .A(n7919), .B(n7918), .Z(n7921) );
  OR U11541 ( .A(n7921), .B(n7920), .Z(n7922) );
  AND U11542 ( .A(n7923), .B(n7922), .Z(n7925) );
  NOR U11543 ( .A(n7925), .B(n7924), .Z(n7926) );
  NANDN U11544 ( .A(n7927), .B(n7926), .Z(n7928) );
  AND U11545 ( .A(n7929), .B(n7928), .Z(n7931) );
  NAND U11546 ( .A(n7931), .B(n7930), .Z(n7933) );
  ANDN U11547 ( .B(n7933), .A(n7932), .Z(n7934) );
  NANDN U11548 ( .A(n7935), .B(n7934), .Z(n7939) );
  AND U11549 ( .A(n7937), .B(n7936), .Z(n7938) );
  NAND U11550 ( .A(n7939), .B(n7938), .Z(n7940) );
  NANDN U11551 ( .A(n7941), .B(n7940), .Z(n7943) );
  OR U11552 ( .A(n7943), .B(n7942), .Z(n7944) );
  AND U11553 ( .A(n7945), .B(n7944), .Z(n7947) );
  ANDN U11554 ( .B(x[570]), .A(y[570]), .Z(n7946) );
  NOR U11555 ( .A(n7947), .B(n7946), .Z(n7948) );
  NANDN U11556 ( .A(n7949), .B(n7948), .Z(n7950) );
  AND U11557 ( .A(n7951), .B(n7950), .Z(n7953) );
  NAND U11558 ( .A(n7953), .B(n7952), .Z(n7955) );
  ANDN U11559 ( .B(n7955), .A(n7954), .Z(n7956) );
  NANDN U11560 ( .A(n7957), .B(n7956), .Z(n7961) );
  AND U11561 ( .A(n7959), .B(n7958), .Z(n7960) );
  NAND U11562 ( .A(n7961), .B(n7960), .Z(n7962) );
  NANDN U11563 ( .A(n7963), .B(n7962), .Z(n7965) );
  OR U11564 ( .A(n7965), .B(n7964), .Z(n7966) );
  AND U11565 ( .A(n7967), .B(n7966), .Z(n7969) );
  ANDN U11566 ( .B(x[576]), .A(y[576]), .Z(n7968) );
  NOR U11567 ( .A(n7969), .B(n7968), .Z(n7970) );
  NANDN U11568 ( .A(n7971), .B(n7970), .Z(n7972) );
  AND U11569 ( .A(n7973), .B(n7972), .Z(n7975) );
  NAND U11570 ( .A(n7975), .B(n7974), .Z(n7977) );
  ANDN U11571 ( .B(n7977), .A(n7976), .Z(n7978) );
  NANDN U11572 ( .A(n7979), .B(n7978), .Z(n7983) );
  AND U11573 ( .A(n7981), .B(n7980), .Z(n7982) );
  NAND U11574 ( .A(n7983), .B(n7982), .Z(n7984) );
  NANDN U11575 ( .A(n7985), .B(n7984), .Z(n7987) );
  OR U11576 ( .A(n7987), .B(n7986), .Z(n7988) );
  AND U11577 ( .A(n7989), .B(n7988), .Z(n7991) );
  NOR U11578 ( .A(n7991), .B(n7990), .Z(n7992) );
  NANDN U11579 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U11580 ( .A(n7995), .B(n7994), .Z(n7997) );
  NAND U11581 ( .A(n7997), .B(n7996), .Z(n7999) );
  ANDN U11582 ( .B(n7999), .A(n7998), .Z(n8000) );
  NANDN U11583 ( .A(n8001), .B(n8000), .Z(n8005) );
  AND U11584 ( .A(n8003), .B(n8002), .Z(n8004) );
  NAND U11585 ( .A(n8005), .B(n8004), .Z(n8006) );
  NANDN U11586 ( .A(n8007), .B(n8006), .Z(n8009) );
  OR U11587 ( .A(n8009), .B(n8008), .Z(n8010) );
  AND U11588 ( .A(n8011), .B(n8010), .Z(n8013) );
  NOR U11589 ( .A(n8013), .B(n8012), .Z(n8014) );
  NANDN U11590 ( .A(n8015), .B(n8014), .Z(n8016) );
  AND U11591 ( .A(n8017), .B(n8016), .Z(n8019) );
  NAND U11592 ( .A(n8019), .B(n8018), .Z(n8021) );
  ANDN U11593 ( .B(n8021), .A(n8020), .Z(n8022) );
  NANDN U11594 ( .A(n8023), .B(n8022), .Z(n8027) );
  AND U11595 ( .A(n8025), .B(n8024), .Z(n8026) );
  NAND U11596 ( .A(n8027), .B(n8026), .Z(n8028) );
  NANDN U11597 ( .A(n8029), .B(n8028), .Z(n8031) );
  OR U11598 ( .A(n8031), .B(n8030), .Z(n8032) );
  AND U11599 ( .A(n8033), .B(n8032), .Z(n8035) );
  ANDN U11600 ( .B(x[594]), .A(y[594]), .Z(n8034) );
  NOR U11601 ( .A(n8035), .B(n8034), .Z(n8036) );
  NANDN U11602 ( .A(n8037), .B(n8036), .Z(n8038) );
  AND U11603 ( .A(n8039), .B(n8038), .Z(n8041) );
  NAND U11604 ( .A(n8041), .B(n8040), .Z(n8043) );
  ANDN U11605 ( .B(n8043), .A(n8042), .Z(n8044) );
  NANDN U11606 ( .A(n8045), .B(n8044), .Z(n8049) );
  AND U11607 ( .A(n8047), .B(n8046), .Z(n8048) );
  NAND U11608 ( .A(n8049), .B(n8048), .Z(n8050) );
  NANDN U11609 ( .A(n8051), .B(n8050), .Z(n8053) );
  OR U11610 ( .A(n8053), .B(n8052), .Z(n8054) );
  AND U11611 ( .A(n8055), .B(n8054), .Z(n8057) );
  ANDN U11612 ( .B(x[600]), .A(y[600]), .Z(n8056) );
  NOR U11613 ( .A(n8057), .B(n8056), .Z(n8058) );
  NANDN U11614 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U11615 ( .A(n8061), .B(n8060), .Z(n8063) );
  NAND U11616 ( .A(n8063), .B(n8062), .Z(n8065) );
  ANDN U11617 ( .B(n8065), .A(n8064), .Z(n8066) );
  NANDN U11618 ( .A(n8067), .B(n8066), .Z(n8071) );
  AND U11619 ( .A(n8069), .B(n8068), .Z(n8070) );
  NAND U11620 ( .A(n8071), .B(n8070), .Z(n8072) );
  NANDN U11621 ( .A(n8073), .B(n8072), .Z(n8075) );
  OR U11622 ( .A(n8075), .B(n8074), .Z(n8076) );
  AND U11623 ( .A(n8077), .B(n8076), .Z(n8079) );
  NOR U11624 ( .A(n8079), .B(n8078), .Z(n8080) );
  NANDN U11625 ( .A(n8081), .B(n8080), .Z(n8082) );
  AND U11626 ( .A(n8083), .B(n8082), .Z(n8085) );
  NAND U11627 ( .A(n8085), .B(n8084), .Z(n8087) );
  ANDN U11628 ( .B(n8087), .A(n8086), .Z(n8088) );
  NANDN U11629 ( .A(n8089), .B(n8088), .Z(n8093) );
  AND U11630 ( .A(n8091), .B(n8090), .Z(n8092) );
  NAND U11631 ( .A(n8093), .B(n8092), .Z(n8094) );
  NANDN U11632 ( .A(n8095), .B(n8094), .Z(n8097) );
  OR U11633 ( .A(n8097), .B(n8096), .Z(n8098) );
  AND U11634 ( .A(n8099), .B(n8098), .Z(n8101) );
  NOR U11635 ( .A(n8101), .B(n8100), .Z(n8102) );
  NANDN U11636 ( .A(n8103), .B(n8102), .Z(n8104) );
  AND U11637 ( .A(n8105), .B(n8104), .Z(n8107) );
  NAND U11638 ( .A(n8107), .B(n8106), .Z(n8109) );
  ANDN U11639 ( .B(n8109), .A(n8108), .Z(n8110) );
  NANDN U11640 ( .A(n8111), .B(n8110), .Z(n8115) );
  AND U11641 ( .A(n8113), .B(n8112), .Z(n8114) );
  NAND U11642 ( .A(n8115), .B(n8114), .Z(n8116) );
  NANDN U11643 ( .A(n8117), .B(n8116), .Z(n8119) );
  OR U11644 ( .A(n8119), .B(n8118), .Z(n8120) );
  AND U11645 ( .A(n8121), .B(n8120), .Z(n8123) );
  NOR U11646 ( .A(n8123), .B(n8122), .Z(n8124) );
  NANDN U11647 ( .A(n8125), .B(n8124), .Z(n8126) );
  AND U11648 ( .A(n8127), .B(n8126), .Z(n8129) );
  NAND U11649 ( .A(n8129), .B(n8128), .Z(n8131) );
  ANDN U11650 ( .B(n8131), .A(n8130), .Z(n8132) );
  NANDN U11651 ( .A(n8133), .B(n8132), .Z(n8137) );
  AND U11652 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND U11653 ( .A(n8137), .B(n8136), .Z(n8138) );
  NANDN U11654 ( .A(n8139), .B(n8138), .Z(n8141) );
  OR U11655 ( .A(n8141), .B(n8140), .Z(n8142) );
  AND U11656 ( .A(n8143), .B(n8142), .Z(n8145) );
  ANDN U11657 ( .B(x[624]), .A(y[624]), .Z(n8144) );
  NOR U11658 ( .A(n8145), .B(n8144), .Z(n8146) );
  NANDN U11659 ( .A(n8147), .B(n8146), .Z(n8148) );
  AND U11660 ( .A(n8149), .B(n8148), .Z(n8151) );
  NAND U11661 ( .A(n8151), .B(n8150), .Z(n8153) );
  ANDN U11662 ( .B(n8153), .A(n8152), .Z(n8154) );
  NANDN U11663 ( .A(n8155), .B(n8154), .Z(n8159) );
  AND U11664 ( .A(n8157), .B(n8156), .Z(n8158) );
  NAND U11665 ( .A(n8159), .B(n8158), .Z(n8160) );
  NANDN U11666 ( .A(n8161), .B(n8160), .Z(n8163) );
  OR U11667 ( .A(n8163), .B(n8162), .Z(n8164) );
  AND U11668 ( .A(n8165), .B(n8164), .Z(n8167) );
  NOR U11669 ( .A(n8167), .B(n8166), .Z(n8168) );
  NANDN U11670 ( .A(n8169), .B(n8168), .Z(n8170) );
  AND U11671 ( .A(n8171), .B(n8170), .Z(n8173) );
  NAND U11672 ( .A(n8173), .B(n8172), .Z(n8175) );
  ANDN U11673 ( .B(n8175), .A(n8174), .Z(n8176) );
  NANDN U11674 ( .A(n8177), .B(n8176), .Z(n8181) );
  AND U11675 ( .A(n8179), .B(n8178), .Z(n8180) );
  NAND U11676 ( .A(n8181), .B(n8180), .Z(n8182) );
  NANDN U11677 ( .A(n8183), .B(n8182), .Z(n8185) );
  OR U11678 ( .A(n8185), .B(n8184), .Z(n8186) );
  AND U11679 ( .A(n8187), .B(n8186), .Z(n8189) );
  NOR U11680 ( .A(n8189), .B(n8188), .Z(n8190) );
  NANDN U11681 ( .A(n8191), .B(n8190), .Z(n8192) );
  AND U11682 ( .A(n8193), .B(n8192), .Z(n8195) );
  NAND U11683 ( .A(n8195), .B(n8194), .Z(n8197) );
  ANDN U11684 ( .B(n8197), .A(n8196), .Z(n8198) );
  NANDN U11685 ( .A(n8199), .B(n8198), .Z(n8203) );
  AND U11686 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND U11687 ( .A(n8203), .B(n8202), .Z(n8204) );
  NANDN U11688 ( .A(n8205), .B(n8204), .Z(n8207) );
  OR U11689 ( .A(n8207), .B(n8206), .Z(n8208) );
  AND U11690 ( .A(n8209), .B(n8208), .Z(n8211) );
  ANDN U11691 ( .B(x[642]), .A(y[642]), .Z(n8210) );
  NOR U11692 ( .A(n8211), .B(n8210), .Z(n8212) );
  NANDN U11693 ( .A(n8213), .B(n8212), .Z(n8214) );
  AND U11694 ( .A(n8235), .B(n8234), .Z(n8239) );
  NAND U11695 ( .A(n8237), .B(n8236), .Z(n8238) );
  OR U11696 ( .A(n8239), .B(n8238), .Z(n8240) );
  AND U11697 ( .A(n8241), .B(n8240), .Z(n8243) );
  NAND U11698 ( .A(n8243), .B(n8242), .Z(n8245) );
  ANDN U11699 ( .B(n8245), .A(n8244), .Z(n8246) );
  NANDN U11700 ( .A(n8247), .B(n8246), .Z(n8251) );
  AND U11701 ( .A(n8249), .B(n8248), .Z(n8250) );
  NAND U11702 ( .A(n8251), .B(n8250), .Z(n8252) );
  NANDN U11703 ( .A(n8253), .B(n8252), .Z(n8255) );
  OR U11704 ( .A(n8255), .B(n8254), .Z(n8256) );
  AND U11705 ( .A(n8257), .B(n8256), .Z(n8261) );
  NAND U11706 ( .A(n8259), .B(n8258), .Z(n8260) );
  OR U11707 ( .A(n8261), .B(n8260), .Z(n8262) );
  AND U11708 ( .A(n8263), .B(n8262), .Z(n8265) );
  NAND U11709 ( .A(n8265), .B(n8264), .Z(n8267) );
  ANDN U11710 ( .B(n8267), .A(n8266), .Z(n8268) );
  NANDN U11711 ( .A(n8269), .B(n8268), .Z(n8273) );
  AND U11712 ( .A(n8271), .B(n8270), .Z(n8272) );
  NAND U11713 ( .A(n8273), .B(n8272), .Z(n8274) );
  NANDN U11714 ( .A(n8275), .B(n8274), .Z(n8277) );
  OR U11715 ( .A(n8277), .B(n8276), .Z(n8278) );
  AND U11716 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U11717 ( .A(n8281), .B(n8280), .Z(n8282) );
  OR U11718 ( .A(n8283), .B(n8282), .Z(n8284) );
  AND U11719 ( .A(n8285), .B(n8284), .Z(n8287) );
  NAND U11720 ( .A(n8287), .B(n8286), .Z(n8289) );
  ANDN U11721 ( .B(n8289), .A(n8288), .Z(n8290) );
  NANDN U11722 ( .A(n8291), .B(n8290), .Z(n8295) );
  AND U11723 ( .A(n8293), .B(n8292), .Z(n8294) );
  NAND U11724 ( .A(n8295), .B(n8294), .Z(n8296) );
  NANDN U11725 ( .A(n8297), .B(n8296), .Z(n8299) );
  OR U11726 ( .A(n8299), .B(n8298), .Z(n8300) );
  AND U11727 ( .A(n8301), .B(n8300), .Z(n8305) );
  NAND U11728 ( .A(n8303), .B(n8302), .Z(n8304) );
  OR U11729 ( .A(n8305), .B(n8304), .Z(n8306) );
  AND U11730 ( .A(n8307), .B(n8306), .Z(n8309) );
  NAND U11731 ( .A(n8309), .B(n8308), .Z(n8311) );
  ANDN U11732 ( .B(n8311), .A(n8310), .Z(n8312) );
  NANDN U11733 ( .A(n8313), .B(n8312), .Z(n8317) );
  AND U11734 ( .A(n8315), .B(n8314), .Z(n8316) );
  NAND U11735 ( .A(n8317), .B(n8316), .Z(n8318) );
  NANDN U11736 ( .A(n8319), .B(n8318), .Z(n8321) );
  OR U11737 ( .A(n8321), .B(n8320), .Z(n8322) );
  AND U11738 ( .A(n8323), .B(n8322), .Z(n8327) );
  NAND U11739 ( .A(n8325), .B(n8324), .Z(n8326) );
  OR U11740 ( .A(n8327), .B(n8326), .Z(n8328) );
  AND U11741 ( .A(n8329), .B(n8328), .Z(n8331) );
  NAND U11742 ( .A(n8331), .B(n8330), .Z(n8333) );
  ANDN U11743 ( .B(n8333), .A(n8332), .Z(n8334) );
  NANDN U11744 ( .A(n8335), .B(n8334), .Z(n8339) );
  AND U11745 ( .A(n8337), .B(n8336), .Z(n8338) );
  NAND U11746 ( .A(n8339), .B(n8338), .Z(n8340) );
  NANDN U11747 ( .A(n8341), .B(n8340), .Z(n8342) );
  OR U11748 ( .A(n8343), .B(n8342), .Z(n8344) );
  AND U11749 ( .A(n8345), .B(n8344), .Z(n8346) );
  NANDN U11750 ( .A(n8347), .B(n8346), .Z(n8348) );
  NAND U11751 ( .A(n8349), .B(n8348), .Z(n8350) );
  NANDN U11752 ( .A(n8351), .B(n8350), .Z(n8352) );
  OR U11753 ( .A(n8353), .B(n8352), .Z(n8354) );
  AND U11754 ( .A(n8355), .B(n8354), .Z(n8356) );
  OR U11755 ( .A(n8357), .B(n8356), .Z(n8358) );
  NAND U11756 ( .A(n8359), .B(n8358), .Z(n8360) );
  NANDN U11757 ( .A(n8361), .B(n8360), .Z(n8362) );
  OR U11758 ( .A(n8363), .B(n8362), .Z(n8364) );
  AND U11759 ( .A(n11583), .B(n8364), .Z(n8366) );
  NAND U11760 ( .A(n8366), .B(n8365), .Z(n8367) );
  NAND U11761 ( .A(n8368), .B(n8367), .Z(n8369) );
  OR U11762 ( .A(n11585), .B(n8369), .Z(n8370) );
  AND U11763 ( .A(n11587), .B(n8370), .Z(n8371) );
  OR U11764 ( .A(n8372), .B(n8371), .Z(n8373) );
  AND U11765 ( .A(n8374), .B(n8373), .Z(n8375) );
  ANDN U11766 ( .B(n8376), .A(n8375), .Z(n8377) );
  NAND U11767 ( .A(n8378), .B(n8377), .Z(n8379) );
  NANDN U11768 ( .A(n8380), .B(n8379), .Z(n8381) );
  OR U11769 ( .A(n8382), .B(n8381), .Z(n8383) );
  AND U11770 ( .A(n8384), .B(n8383), .Z(n8386) );
  NANDN U11771 ( .A(y[706]), .B(x[706]), .Z(n8385) );
  NAND U11772 ( .A(n8386), .B(n8385), .Z(n8388) );
  ANDN U11773 ( .B(n8388), .A(n8387), .Z(n8389) );
  NANDN U11774 ( .A(n8390), .B(n8389), .Z(n8394) );
  AND U11775 ( .A(n8392), .B(n8391), .Z(n8393) );
  NAND U11776 ( .A(n8394), .B(n8393), .Z(n8395) );
  NANDN U11777 ( .A(n8396), .B(n8395), .Z(n8398) );
  OR U11778 ( .A(n8398), .B(n8397), .Z(n8399) );
  NAND U11779 ( .A(n8400), .B(n8399), .Z(n8402) );
  AND U11780 ( .A(n8402), .B(n8401), .Z(n8403) );
  NAND U11781 ( .A(n8404), .B(n8403), .Z(n8405) );
  NAND U11782 ( .A(n8406), .B(n8405), .Z(n8407) );
  AND U11783 ( .A(n8408), .B(n8407), .Z(n8409) );
  OR U11784 ( .A(n8409), .B(n11609), .Z(n8410) );
  NAND U11785 ( .A(n11611), .B(n8410), .Z(n8411) );
  NAND U11786 ( .A(n11613), .B(n8411), .Z(n8412) );
  NANDN U11787 ( .A(n11615), .B(n8412), .Z(n8413) );
  NAND U11788 ( .A(n8414), .B(n8413), .Z(n8415) );
  NANDN U11789 ( .A(n8416), .B(n8415), .Z(n8420) );
  AND U11790 ( .A(n8418), .B(n8417), .Z(n8419) );
  NAND U11791 ( .A(n8420), .B(n8419), .Z(n8421) );
  NANDN U11792 ( .A(n8422), .B(n8421), .Z(n8424) );
  OR U11793 ( .A(n8424), .B(n8423), .Z(n8425) );
  NAND U11794 ( .A(n8426), .B(n8425), .Z(n8427) );
  NANDN U11795 ( .A(n8428), .B(n8427), .Z(n8432) );
  AND U11796 ( .A(n8430), .B(n8429), .Z(n8431) );
  NAND U11797 ( .A(n8432), .B(n8431), .Z(n8433) );
  NANDN U11798 ( .A(n8434), .B(n8433), .Z(n8435) );
  OR U11799 ( .A(n8436), .B(n8435), .Z(n8437) );
  AND U11800 ( .A(n8438), .B(n8437), .Z(n8439) );
  NANDN U11801 ( .A(n8440), .B(n8439), .Z(n8441) );
  ANDN U11802 ( .B(n8441), .A(n11635), .Z(n8443) );
  NAND U11803 ( .A(n8443), .B(n8442), .Z(n8444) );
  NAND U11804 ( .A(n8445), .B(n8444), .Z(n8446) );
  NANDN U11805 ( .A(n8446), .B(n11637), .Z(n8447) );
  ANDN U11806 ( .B(n8447), .A(n11639), .Z(n8448) );
  OR U11807 ( .A(n8449), .B(n8448), .Z(n8450) );
  NAND U11808 ( .A(n8451), .B(n8450), .Z(n8452) );
  NANDN U11809 ( .A(n8453), .B(n8452), .Z(n8454) );
  OR U11810 ( .A(n8455), .B(n8454), .Z(n8456) );
  AND U11811 ( .A(n8457), .B(n8456), .Z(n8458) );
  NANDN U11812 ( .A(n8459), .B(n8458), .Z(n8460) );
  NAND U11813 ( .A(n8461), .B(n8460), .Z(n8465) );
  AND U11814 ( .A(n8463), .B(n8462), .Z(n8464) );
  NAND U11815 ( .A(n8465), .B(n8464), .Z(n8466) );
  NANDN U11816 ( .A(n8467), .B(n8466), .Z(n8469) );
  ANDN U11817 ( .B(x[734]), .A(y[734]), .Z(n8468) );
  OR U11818 ( .A(n8469), .B(n8468), .Z(n8470) );
  NAND U11819 ( .A(n8471), .B(n8470), .Z(n8472) );
  NANDN U11820 ( .A(n8473), .B(n8472), .Z(n8477) );
  AND U11821 ( .A(n8475), .B(n8474), .Z(n8476) );
  NAND U11822 ( .A(n8477), .B(n8476), .Z(n8478) );
  NANDN U11823 ( .A(n8479), .B(n8478), .Z(n8481) );
  OR U11824 ( .A(n8481), .B(n8480), .Z(n8482) );
  NAND U11825 ( .A(n8483), .B(n8482), .Z(n8484) );
  NANDN U11826 ( .A(n8485), .B(n8484), .Z(n8489) );
  AND U11827 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U11828 ( .A(n8489), .B(n8488), .Z(n8490) );
  NANDN U11829 ( .A(n8491), .B(n8490), .Z(n8493) );
  OR U11830 ( .A(n8493), .B(n8492), .Z(n8494) );
  NAND U11831 ( .A(n8495), .B(n8494), .Z(n8496) );
  NANDN U11832 ( .A(n8497), .B(n8496), .Z(n8501) );
  AND U11833 ( .A(n8499), .B(n8498), .Z(n8500) );
  NAND U11834 ( .A(n8501), .B(n8500), .Z(n8502) );
  NANDN U11835 ( .A(n8503), .B(n8502), .Z(n8505) );
  OR U11836 ( .A(n8505), .B(n8504), .Z(n8506) );
  NAND U11837 ( .A(n8507), .B(n8506), .Z(n8508) );
  NANDN U11838 ( .A(n8509), .B(n8508), .Z(n8513) );
  AND U11839 ( .A(n8511), .B(n8510), .Z(n8512) );
  NAND U11840 ( .A(n8513), .B(n8512), .Z(n8514) );
  NANDN U11841 ( .A(n8515), .B(n8514), .Z(n8517) );
  OR U11842 ( .A(n8517), .B(n8516), .Z(n8518) );
  NAND U11843 ( .A(n8519), .B(n8518), .Z(n8520) );
  NANDN U11844 ( .A(n8521), .B(n8520), .Z(n8525) );
  AND U11845 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U11846 ( .A(n8525), .B(n8524), .Z(n8526) );
  NANDN U11847 ( .A(n8527), .B(n8526), .Z(n8529) );
  OR U11848 ( .A(n8529), .B(n8528), .Z(n8530) );
  NAND U11849 ( .A(n8531), .B(n8530), .Z(n8532) );
  NANDN U11850 ( .A(n8533), .B(n8532), .Z(n8537) );
  AND U11851 ( .A(n8535), .B(n8534), .Z(n8536) );
  NAND U11852 ( .A(n8537), .B(n8536), .Z(n8538) );
  NANDN U11853 ( .A(n8539), .B(n8538), .Z(n8540) );
  OR U11854 ( .A(n8541), .B(n8540), .Z(n8542) );
  AND U11855 ( .A(n8543), .B(n8542), .Z(n8544) );
  NANDN U11856 ( .A(n8545), .B(n8544), .Z(n8546) );
  AND U11857 ( .A(n8547), .B(n8546), .Z(n8548) );
  ANDN U11858 ( .B(n11707), .A(n8548), .Z(n8549) );
  NANDN U11859 ( .A(n8550), .B(n8549), .Z(n8551) );
  AND U11860 ( .A(n8552), .B(n8551), .Z(n8554) );
  NANDN U11861 ( .A(n8554), .B(n8553), .Z(n8555) );
  AND U11862 ( .A(n8556), .B(n8555), .Z(n8557) );
  OR U11863 ( .A(n8558), .B(n8557), .Z(n8559) );
  NAND U11864 ( .A(n8560), .B(n8559), .Z(n8564) );
  AND U11865 ( .A(n8562), .B(n8561), .Z(n8563) );
  NAND U11866 ( .A(n8564), .B(n8563), .Z(n8565) );
  NANDN U11867 ( .A(n8566), .B(n8565), .Z(n8568) );
  OR U11868 ( .A(n8568), .B(n8567), .Z(n8569) );
  AND U11869 ( .A(n8570), .B(n8569), .Z(n8574) );
  NAND U11870 ( .A(n8572), .B(n8571), .Z(n8573) );
  OR U11871 ( .A(n8574), .B(n8573), .Z(n8575) );
  AND U11872 ( .A(n8576), .B(n8575), .Z(n8578) );
  NAND U11873 ( .A(n8578), .B(n8577), .Z(n8580) );
  AND U11874 ( .A(n8580), .B(n8579), .Z(n8581) );
  NAND U11875 ( .A(n8582), .B(n8581), .Z(n8583) );
  NAND U11876 ( .A(n8584), .B(n8583), .Z(n8585) );
  AND U11877 ( .A(n8586), .B(n8585), .Z(n8588) );
  NANDN U11878 ( .A(n8588), .B(n8587), .Z(n8590) );
  ANDN U11879 ( .B(n8590), .A(n8589), .Z(n8592) );
  NANDN U11880 ( .A(n8592), .B(n8591), .Z(n8593) );
  NANDN U11881 ( .A(n8594), .B(n8593), .Z(n8595) );
  NAND U11882 ( .A(n8596), .B(n8595), .Z(n8597) );
  NANDN U11883 ( .A(n8598), .B(n8597), .Z(n8599) );
  NAND U11884 ( .A(n8600), .B(n8599), .Z(n8602) );
  ANDN U11885 ( .B(n8602), .A(n8601), .Z(n8604) );
  NANDN U11886 ( .A(n8604), .B(n8603), .Z(n8605) );
  NANDN U11887 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U11888 ( .A(n8608), .B(n8607), .Z(n8609) );
  NAND U11889 ( .A(n11752), .B(n8609), .Z(n8610) );
  ANDN U11890 ( .B(n8610), .A(n11755), .Z(n8611) );
  OR U11891 ( .A(n8612), .B(n8611), .Z(n8613) );
  NAND U11892 ( .A(n8614), .B(n8613), .Z(n8615) );
  NANDN U11893 ( .A(n8616), .B(n8615), .Z(n8617) );
  OR U11894 ( .A(n8618), .B(n8617), .Z(n8619) );
  AND U11895 ( .A(n8620), .B(n8619), .Z(n8621) );
  NANDN U11896 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U11897 ( .A(n8624), .B(n8623), .Z(n8626) );
  NOR U11898 ( .A(n8626), .B(n8625), .Z(n8627) );
  NANDN U11899 ( .A(n8628), .B(n8627), .Z(n8629) );
  AND U11900 ( .A(n8630), .B(n8629), .Z(n8631) );
  NANDN U11901 ( .A(n8632), .B(n8631), .Z(n8633) );
  NAND U11902 ( .A(n8634), .B(n8633), .Z(n8635) );
  NANDN U11903 ( .A(n8636), .B(n8635), .Z(n8638) );
  OR U11904 ( .A(n8638), .B(n8637), .Z(n8639) );
  NAND U11905 ( .A(n8640), .B(n8639), .Z(n8644) );
  AND U11906 ( .A(n8642), .B(n8641), .Z(n8643) );
  NAND U11907 ( .A(n8644), .B(n8643), .Z(n8645) );
  NANDN U11908 ( .A(n8646), .B(n8645), .Z(n8648) );
  OR U11909 ( .A(n8648), .B(n8647), .Z(n8649) );
  NAND U11910 ( .A(n8650), .B(n8649), .Z(n8654) );
  AND U11911 ( .A(n8652), .B(n8651), .Z(n8653) );
  NAND U11912 ( .A(n8654), .B(n8653), .Z(n8655) );
  NANDN U11913 ( .A(n8656), .B(n8655), .Z(n8657) );
  OR U11914 ( .A(n8658), .B(n8657), .Z(n8659) );
  AND U11915 ( .A(n8660), .B(n8659), .Z(n8662) );
  NAND U11916 ( .A(n8662), .B(n8661), .Z(n8664) );
  ANDN U11917 ( .B(n8664), .A(n8663), .Z(n8665) );
  NANDN U11918 ( .A(n8666), .B(n8665), .Z(n8670) );
  AND U11919 ( .A(n8668), .B(n8667), .Z(n8669) );
  NAND U11920 ( .A(n8670), .B(n8669), .Z(n8671) );
  NANDN U11921 ( .A(n8672), .B(n8671), .Z(n8674) );
  OR U11922 ( .A(n8674), .B(n8673), .Z(n8675) );
  AND U11923 ( .A(n8676), .B(n8675), .Z(n8680) );
  NAND U11924 ( .A(n8678), .B(n8677), .Z(n8679) );
  OR U11925 ( .A(n8680), .B(n8679), .Z(n8681) );
  AND U11926 ( .A(n8682), .B(n8681), .Z(n8684) );
  NAND U11927 ( .A(n8684), .B(n8683), .Z(n8686) );
  ANDN U11928 ( .B(x[808]), .A(y[808]), .Z(n8685) );
  ANDN U11929 ( .B(n8686), .A(n8685), .Z(n8687) );
  NANDN U11930 ( .A(n8688), .B(n8687), .Z(n8692) );
  AND U11931 ( .A(n8690), .B(n8689), .Z(n8691) );
  NAND U11932 ( .A(n8692), .B(n8691), .Z(n8693) );
  NANDN U11933 ( .A(n8694), .B(n8693), .Z(n8696) );
  OR U11934 ( .A(n8696), .B(n8695), .Z(n8697) );
  NAND U11935 ( .A(n8698), .B(n8697), .Z(n8702) );
  NANDN U11936 ( .A(y[812]), .B(x[812]), .Z(n8699) );
  AND U11937 ( .A(n8700), .B(n8699), .Z(n8701) );
  NAND U11938 ( .A(n8702), .B(n8701), .Z(n8703) );
  NANDN U11939 ( .A(n8704), .B(n8703), .Z(n8706) );
  OR U11940 ( .A(n8706), .B(n8705), .Z(n8707) );
  NAND U11941 ( .A(n8708), .B(n8707), .Z(n8709) );
  NANDN U11942 ( .A(n8710), .B(n8709), .Z(n8714) );
  AND U11943 ( .A(n8712), .B(n8711), .Z(n8713) );
  NAND U11944 ( .A(n8714), .B(n8713), .Z(n8715) );
  NANDN U11945 ( .A(n8716), .B(n8715), .Z(n8718) );
  OR U11946 ( .A(n8718), .B(n8717), .Z(n8719) );
  NAND U11947 ( .A(n8720), .B(n8719), .Z(n8721) );
  AND U11948 ( .A(n11847), .B(n8732), .Z(n8735) );
  NANDN U11949 ( .A(n8734), .B(n8733), .Z(n11849) );
  OR U11950 ( .A(n8735), .B(n11849), .Z(n8736) );
  AND U11951 ( .A(n8737), .B(n8736), .Z(n8738) );
  NAND U11952 ( .A(n8738), .B(n11851), .Z(n8740) );
  ANDN U11953 ( .B(n8740), .A(n8739), .Z(n8741) );
  NANDN U11954 ( .A(n11853), .B(n8741), .Z(n8745) );
  AND U11955 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U11956 ( .A(n8745), .B(n8744), .Z(n8746) );
  NANDN U11957 ( .A(n8747), .B(n8746), .Z(n8749) );
  OR U11958 ( .A(n8749), .B(n8748), .Z(n8750) );
  AND U11959 ( .A(n8751), .B(n8750), .Z(n8755) );
  NAND U11960 ( .A(n8753), .B(n8752), .Z(n8754) );
  OR U11961 ( .A(n8755), .B(n8754), .Z(n8756) );
  AND U11962 ( .A(n8757), .B(n8756), .Z(n8759) );
  NAND U11963 ( .A(n8759), .B(n8758), .Z(n8761) );
  ANDN U11964 ( .B(n8761), .A(n8760), .Z(n8762) );
  NANDN U11965 ( .A(n11869), .B(n8762), .Z(n8765) );
  AND U11966 ( .A(n11871), .B(n8763), .Z(n8764) );
  NAND U11967 ( .A(n8765), .B(n8764), .Z(n8766) );
  AND U11968 ( .A(n8776), .B(n8775), .Z(n8778) );
  NAND U11969 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U11970 ( .A(n8780), .B(n8779), .Z(n8781) );
  NANDN U11971 ( .A(n11911), .B(n8781), .Z(n8782) );
  AND U11972 ( .A(n11913), .B(n8782), .Z(n8783) );
  OR U11973 ( .A(n11915), .B(n8783), .Z(n8784) );
  NAND U11974 ( .A(n11917), .B(n8784), .Z(n8785) );
  NANDN U11975 ( .A(n11919), .B(n8785), .Z(n8786) );
  NAND U11976 ( .A(n11921), .B(n8786), .Z(n8787) );
  ANDN U11977 ( .B(n8787), .A(n11923), .Z(n8788) );
  NANDN U11978 ( .A(n8789), .B(n8788), .Z(n8792) );
  AND U11979 ( .A(n8790), .B(n11925), .Z(n8791) );
  NAND U11980 ( .A(n8792), .B(n8791), .Z(n8793) );
  NANDN U11981 ( .A(n8794), .B(n8793), .Z(n8796) );
  OR U11982 ( .A(n8796), .B(n8795), .Z(n8797) );
  ANDN U11983 ( .B(n8804), .A(n8803), .Z(n8805) );
  NAND U11984 ( .A(n11961), .B(n8805), .Z(n8806) );
  AND U11985 ( .A(n8807), .B(n8806), .Z(n8808) );
  NAND U11986 ( .A(n8809), .B(n8808), .Z(n8810) );
  NANDN U11987 ( .A(n8811), .B(n8810), .Z(n8813) );
  OR U11988 ( .A(n8813), .B(n8812), .Z(n8814) );
  AND U11989 ( .A(n8815), .B(n8814), .Z(n8819) );
  NANDN U11990 ( .A(n8817), .B(n8816), .Z(n8818) );
  OR U11991 ( .A(n8819), .B(n8818), .Z(n8820) );
  AND U11992 ( .A(n11975), .B(n8820), .Z(n8821) );
  ANDN U11993 ( .B(n11977), .A(n8821), .Z(n8822) );
  NANDN U11994 ( .A(n8823), .B(n8822), .Z(n8824) );
  ANDN U11995 ( .B(n8824), .A(n11978), .Z(n8825) );
  NANDN U11996 ( .A(n11983), .B(n8825), .Z(n8827) );
  ANDN U11997 ( .B(n8827), .A(n8826), .Z(n8828) );
  NAND U11998 ( .A(n11985), .B(n8828), .Z(n8829) );
  NAND U11999 ( .A(n11987), .B(n8829), .Z(n8830) );
  AND U12000 ( .A(n8830), .B(n11989), .Z(n8831) );
  NANDN U12001 ( .A(n8832), .B(n8831), .Z(n8833) );
  ANDN U12002 ( .B(n8833), .A(n11995), .Z(n8834) );
  NANDN U12003 ( .A(n11990), .B(n8834), .Z(n8835) );
  AND U12004 ( .A(n8836), .B(n8835), .Z(n8837) );
  NANDN U12005 ( .A(n11997), .B(n8837), .Z(n8838) );
  NAND U12006 ( .A(n11999), .B(n8838), .Z(n8839) );
  NANDN U12007 ( .A(n12001), .B(n8839), .Z(n8842) );
  ANDN U12008 ( .B(n8840), .A(n12002), .Z(n8841) );
  NAND U12009 ( .A(n8842), .B(n8841), .Z(n8843) );
  NANDN U12010 ( .A(n8844), .B(n8843), .Z(n8845) );
  NANDN U12011 ( .A(n8845), .B(n12004), .Z(n8846) );
  AND U12012 ( .A(n8847), .B(n8846), .Z(n8849) );
  NAND U12013 ( .A(n8849), .B(n8848), .Z(n8851) );
  ANDN U12014 ( .B(n8851), .A(n8850), .Z(n8852) );
  NANDN U12015 ( .A(n8853), .B(n8852), .Z(n8854) );
  AND U12016 ( .A(n8855), .B(n8854), .Z(n8856) );
  NAND U12017 ( .A(n8857), .B(n8856), .Z(n8858) );
  NANDN U12018 ( .A(n8859), .B(n8858), .Z(n8861) );
  OR U12019 ( .A(n8861), .B(n8860), .Z(n8862) );
  AND U12020 ( .A(n8865), .B(n8864), .Z(n8866) );
  NOR U12021 ( .A(n8870), .B(n8869), .Z(n12028) );
  NAND U12022 ( .A(n8872), .B(n8871), .Z(n12031) );
  ANDN U12023 ( .B(n8885), .A(n8884), .Z(n12067) );
  NANDN U12024 ( .A(n12141), .B(n8927), .Z(n8928) );
  NAND U12025 ( .A(n12143), .B(n8928), .Z(n8929) );
  ANDN U12026 ( .B(n8929), .A(n12145), .Z(n8930) );
  NANDN U12027 ( .A(n8931), .B(n8930), .Z(n8934) );
  AND U12028 ( .A(n8932), .B(n12146), .Z(n8933) );
  NAND U12029 ( .A(n8934), .B(n8933), .Z(n8935) );
  NANDN U12030 ( .A(n8936), .B(n8935), .Z(n8937) );
  OR U12031 ( .A(n8938), .B(n8937), .Z(n8939) );
  AND U12032 ( .A(n8940), .B(n8939), .Z(n8942) );
  NAND U12033 ( .A(n8942), .B(n8941), .Z(n8944) );
  ANDN U12034 ( .B(n8944), .A(n8943), .Z(n8945) );
  NANDN U12035 ( .A(n8946), .B(n8945), .Z(n8950) );
  AND U12036 ( .A(n8948), .B(n8947), .Z(n8949) );
  NAND U12037 ( .A(n8950), .B(n8949), .Z(n8951) );
  NANDN U12038 ( .A(n8952), .B(n8951), .Z(n8954) );
  OR U12039 ( .A(n8954), .B(n8953), .Z(n8955) );
  AND U12040 ( .A(n8956), .B(n8955), .Z(n8960) );
  NAND U12041 ( .A(n8958), .B(n8957), .Z(n8959) );
  OR U12042 ( .A(n8960), .B(n8959), .Z(n8961) );
  AND U12043 ( .A(n8978), .B(n8977), .Z(n8979) );
  AND U12044 ( .A(n8985), .B(n8984), .Z(n12200) );
  ANDN U12045 ( .B(n8987), .A(n8986), .Z(n12203) );
  AND U12046 ( .A(n8994), .B(n8993), .Z(n12231) );
  NANDN U12047 ( .A(y[1000]), .B(x[1000]), .Z(n12238) );
  AND U12048 ( .A(n9004), .B(n9003), .Z(n9005) );
  AND U12049 ( .A(n9010), .B(n9009), .Z(n12261) );
  ANDN U12050 ( .B(n9012), .A(n9011), .Z(n12263) );
  NOR U12051 ( .A(n9034), .B(n9033), .Z(n12286) );
  NANDN U12052 ( .A(n9041), .B(n9040), .Z(n9045) );
  ANDN U12053 ( .B(n9043), .A(n9042), .Z(n9044) );
  NAND U12054 ( .A(n9045), .B(n9044), .Z(n9046) );
  NANDN U12055 ( .A(n9047), .B(n9046), .Z(n9048) );
  OR U12056 ( .A(n9049), .B(n9048), .Z(n9050) );
  AND U12057 ( .A(n9051), .B(n9050), .Z(n9053) );
  NAND U12058 ( .A(n9053), .B(n9052), .Z(n9055) );
  ANDN U12059 ( .B(n9055), .A(n9054), .Z(n9056) );
  NANDN U12060 ( .A(n9057), .B(n9056), .Z(n9061) );
  AND U12061 ( .A(n9059), .B(n9058), .Z(n9060) );
  NAND U12062 ( .A(n9061), .B(n9060), .Z(n9062) );
  NANDN U12063 ( .A(n9063), .B(n9062), .Z(n9064) );
  OR U12064 ( .A(n9065), .B(n9064), .Z(n9066) );
  AND U12065 ( .A(n9067), .B(n9066), .Z(n9068) );
  NANDN U12066 ( .A(n12346), .B(n9068), .Z(n9069) );
  NAND U12067 ( .A(n9070), .B(n9069), .Z(n9071) );
  NANDN U12068 ( .A(n12351), .B(n9071), .Z(n9074) );
  AND U12069 ( .A(n9072), .B(n12352), .Z(n9073) );
  NAND U12070 ( .A(n9074), .B(n9073), .Z(n9075) );
  NAND U12071 ( .A(n12355), .B(n9075), .Z(n9076) );
  NANDN U12072 ( .A(n9076), .B(n12358), .Z(n9077) );
  AND U12073 ( .A(n9078), .B(n9077), .Z(n9079) );
  OR U12074 ( .A(n12363), .B(n9079), .Z(n9080) );
  NAND U12075 ( .A(n12365), .B(n9080), .Z(n9081) );
  NANDN U12076 ( .A(n12367), .B(n9081), .Z(n9082) );
  NAND U12077 ( .A(n12369), .B(n9082), .Z(n9083) );
  NANDN U12078 ( .A(n12370), .B(n9083), .Z(n9084) );
  AND U12079 ( .A(n9085), .B(n9084), .Z(n9086) );
  AND U12080 ( .A(n9086), .B(n12373), .Z(n9087) );
  NANDN U12081 ( .A(n9087), .B(n12374), .Z(n9088) );
  AND U12082 ( .A(n9089), .B(n9088), .Z(n9090) );
  OR U12083 ( .A(n12379), .B(n9090), .Z(n9091) );
  NAND U12084 ( .A(n12381), .B(n9091), .Z(n9092) );
  NANDN U12085 ( .A(n12383), .B(n9092), .Z(n9093) );
  AND U12086 ( .A(n12385), .B(n9093), .Z(n9094) );
  OR U12087 ( .A(n12386), .B(n9094), .Z(n9095) );
  NAND U12088 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U12089 ( .A(n9105), .B(n9104), .Z(n12419) );
  NOR U12090 ( .A(n9110), .B(n9109), .Z(n12432) );
  NAND U12091 ( .A(n9112), .B(n9111), .Z(n12434) );
  IV U12092 ( .A(n12448), .Z(n9117) );
  NAND U12093 ( .A(n9120), .B(n9119), .Z(n12465) );
  NAND U12094 ( .A(n9122), .B(n9121), .Z(n12477) );
  IV U12095 ( .A(n12477), .Z(n9123) );
  IV U12096 ( .A(n12504), .Z(n9137) );
  NOR U12097 ( .A(n9151), .B(n9150), .Z(n12562) );
  NAND U12098 ( .A(n9154), .B(n9153), .Z(n12564) );
  NAND U12099 ( .A(n9158), .B(n9157), .Z(n12578) );
  IV U12100 ( .A(n12610), .Z(n9177) );
  NOR U12101 ( .A(n9183), .B(n9182), .Z(n12639) );
  NAND U12102 ( .A(n9185), .B(n9184), .Z(n12640) );
  NOR U12103 ( .A(n9202), .B(n9201), .Z(n12692) );
  ANDN U12104 ( .B(n9207), .A(n9206), .Z(n12709) );
  ANDN U12105 ( .B(n9221), .A(n9220), .Z(n12758) );
  ANDN U12106 ( .B(n9223), .A(n9222), .Z(n12763) );
  NAND U12107 ( .A(n9226), .B(n9225), .Z(n12765) );
  IV U12108 ( .A(n12765), .Z(n9227) );
  NAND U12109 ( .A(n9239), .B(n9238), .Z(n9240) );
  NAND U12110 ( .A(n9241), .B(n9240), .Z(n9242) );
  NAND U12111 ( .A(n9243), .B(n9242), .Z(n12805) );
  IV U12112 ( .A(n12838), .Z(n9254) );
  AND U12113 ( .A(n9262), .B(n9261), .Z(n12869) );
  NANDN U12114 ( .A(y[1304]), .B(x[1304]), .Z(n9298) );
  OR U12115 ( .A(n9299), .B(n9298), .Z(n9300) );
  AND U12116 ( .A(n9301), .B(n9300), .Z(n12981) );
  NAND U12117 ( .A(n9322), .B(n9321), .Z(n9323) );
  NAND U12118 ( .A(n9324), .B(n9323), .Z(n9325) );
  AND U12119 ( .A(n9326), .B(n9325), .Z(n9327) );
  OR U12120 ( .A(n13054), .B(n9327), .Z(n9328) );
  AND U12121 ( .A(n13057), .B(n9328), .Z(n9329) );
  OR U12122 ( .A(n9329), .B(n13058), .Z(n9330) );
  AND U12123 ( .A(n13061), .B(n9330), .Z(n9331) );
  OR U12124 ( .A(n9331), .B(n13062), .Z(n9332) );
  NAND U12125 ( .A(n13065), .B(n9332), .Z(n9333) );
  ANDN U12126 ( .B(n9333), .A(n13066), .Z(n9334) );
  OR U12127 ( .A(n13069), .B(n9334), .Z(n9335) );
  NAND U12128 ( .A(n13071), .B(n9335), .Z(n9336) );
  NANDN U12129 ( .A(n13073), .B(n9336), .Z(n9339) );
  ANDN U12130 ( .B(n9337), .A(n13075), .Z(n9338) );
  NAND U12131 ( .A(n9339), .B(n9338), .Z(n9340) );
  NAND U12132 ( .A(n13077), .B(n9340), .Z(n9341) );
  NANDN U12133 ( .A(n9341), .B(n13080), .Z(n9342) );
  AND U12134 ( .A(n9343), .B(n9342), .Z(n9344) );
  OR U12135 ( .A(n13085), .B(n9344), .Z(n9345) );
  NOR U12136 ( .A(n9349), .B(n9348), .Z(n13116) );
  ANDN U12137 ( .B(n9351), .A(n9350), .Z(n13119) );
  NAND U12138 ( .A(n9363), .B(n9362), .Z(n13143) );
  NANDN U12139 ( .A(n9377), .B(n9376), .Z(n13200) );
  ANDN U12140 ( .B(x[1398]), .A(y[1398]), .Z(n9387) );
  AND U12141 ( .A(n9389), .B(n9388), .Z(n13220) );
  NAND U12142 ( .A(n9394), .B(n9393), .Z(n13238) );
  IV U12143 ( .A(n13238), .Z(n9395) );
  NAND U12144 ( .A(n9397), .B(n9396), .Z(n13251) );
  NANDN U12145 ( .A(n9400), .B(n9399), .Z(n9401) );
  NAND U12146 ( .A(n9402), .B(n9401), .Z(n9403) );
  AND U12147 ( .A(n9404), .B(n9403), .Z(n9406) );
  ANDN U12148 ( .B(n9406), .A(n9405), .Z(n9410) );
  NANDN U12149 ( .A(n9408), .B(n9407), .Z(n9409) );
  NAND U12150 ( .A(n9410), .B(n9409), .Z(n13262) );
  NAND U12151 ( .A(n9428), .B(n9427), .Z(n13325) );
  ANDN U12152 ( .B(n9431), .A(n9430), .Z(n13349) );
  ANDN U12153 ( .B(n9433), .A(n9432), .Z(n13351) );
  IV U12154 ( .A(n13355), .Z(n9436) );
  NOR U12155 ( .A(n9442), .B(n9441), .Z(n13378) );
  NAND U12156 ( .A(n9444), .B(n9443), .Z(n13381) );
  NOR U12157 ( .A(n9459), .B(n9458), .Z(n13457) );
  NANDN U12158 ( .A(n9467), .B(n9466), .Z(n9468) );
  ANDN U12159 ( .B(n9468), .A(n9472), .Z(n9470) );
  ANDN U12160 ( .B(n9470), .A(n9469), .Z(n13473) );
  OR U12161 ( .A(n9472), .B(n9471), .Z(n9474) );
  ANDN U12162 ( .B(n9474), .A(n9473), .Z(n13475) );
  NAND U12163 ( .A(n9488), .B(n9487), .Z(n10186) );
  AND U12164 ( .A(n9490), .B(n9489), .Z(n9491) );
  OR U12165 ( .A(n9492), .B(n9491), .Z(n9493) );
  NAND U12166 ( .A(n9494), .B(n9493), .Z(n9495) );
  NANDN U12167 ( .A(n9496), .B(n9495), .Z(n9500) );
  AND U12168 ( .A(n9498), .B(n9497), .Z(n9499) );
  NAND U12169 ( .A(n9500), .B(n9499), .Z(n9501) );
  NANDN U12170 ( .A(n9502), .B(n9501), .Z(n9504) );
  OR U12171 ( .A(n9504), .B(n9503), .Z(n9505) );
  NAND U12172 ( .A(n9506), .B(n9505), .Z(n9507) );
  NANDN U12173 ( .A(n9508), .B(n9507), .Z(n9509) );
  OR U12174 ( .A(n9509), .B(n13573), .Z(n9510) );
  AND U12175 ( .A(n9511), .B(n9510), .Z(n9512) );
  OR U12176 ( .A(n13577), .B(n9512), .Z(n9513) );
  NAND U12177 ( .A(n9514), .B(n9513), .Z(n9515) );
  NAND U12178 ( .A(n9519), .B(n9518), .Z(n13610) );
  IV U12179 ( .A(n13610), .Z(n9520) );
  AND U12180 ( .A(n9523), .B(n9522), .Z(n13623) );
  IV U12181 ( .A(n13635), .Z(n9526) );
  IV U12182 ( .A(n13636), .Z(n9528) );
  AND U12183 ( .A(n9532), .B(n9531), .Z(n13661) );
  NOR U12184 ( .A(n9538), .B(n9537), .Z(n13699) );
  NAND U12185 ( .A(n9541), .B(n9540), .Z(n13700) );
  IV U12186 ( .A(n13700), .Z(n9542) );
  NAND U12187 ( .A(n9552), .B(n9551), .Z(n13754) );
  ANDN U12188 ( .B(n9557), .A(n9556), .Z(n13769) );
  NAND U12189 ( .A(n9568), .B(n9567), .Z(n9569) );
  NANDN U12190 ( .A(n9570), .B(n9569), .Z(n9571) );
  AND U12191 ( .A(n9571), .B(n13813), .Z(n9573) );
  NANDN U12192 ( .A(y[1654]), .B(x[1654]), .Z(n9572) );
  AND U12193 ( .A(n9573), .B(n9572), .Z(n9574) );
  OR U12194 ( .A(n13815), .B(n9574), .Z(n9575) );
  NAND U12195 ( .A(n13817), .B(n9575), .Z(n9576) );
  NANDN U12196 ( .A(n9577), .B(n9576), .Z(n9578) );
  OR U12197 ( .A(n13819), .B(n9578), .Z(n9579) );
  AND U12198 ( .A(n9580), .B(n9579), .Z(n9581) );
  NOR U12199 ( .A(n9582), .B(n9581), .Z(n9584) );
  NAND U12200 ( .A(n9584), .B(n9583), .Z(n9585) );
  AND U12201 ( .A(n9586), .B(n9585), .Z(n9587) );
  NAND U12202 ( .A(n9588), .B(n9587), .Z(n9589) );
  NANDN U12203 ( .A(n9590), .B(n9589), .Z(n9591) );
  OR U12204 ( .A(n9592), .B(n9591), .Z(n9593) );
  AND U12205 ( .A(n9594), .B(n9593), .Z(n9595) );
  NAND U12206 ( .A(n13832), .B(n9595), .Z(n9596) );
  AND U12207 ( .A(n9597), .B(n9596), .Z(n9598) );
  OR U12208 ( .A(n13837), .B(n9598), .Z(n9599) );
  NAND U12209 ( .A(n13839), .B(n9599), .Z(n9600) );
  NANDN U12210 ( .A(n13841), .B(n9600), .Z(n9601) );
  NAND U12211 ( .A(n13843), .B(n9601), .Z(n9602) );
  AND U12212 ( .A(n9602), .B(n13844), .Z(n9603) );
  NANDN U12213 ( .A(n9604), .B(n9603), .Z(n9605) );
  NAND U12214 ( .A(n9606), .B(n9605), .Z(n9607) );
  NANDN U12215 ( .A(n9608), .B(n9607), .Z(n9609) );
  AND U12216 ( .A(n9610), .B(n9609), .Z(n9616) );
  OR U12217 ( .A(n9612), .B(n9611), .Z(n9614) );
  ANDN U12218 ( .B(n9614), .A(n9613), .Z(n9615) );
  NANDN U12219 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U12220 ( .A(n13859), .B(n9617), .Z(n9618) );
  NAND U12221 ( .A(n9619), .B(n9618), .Z(n9621) );
  ANDN U12222 ( .B(n9640), .A(n9639), .Z(n13917) );
  ANDN U12223 ( .B(n9647), .A(n9646), .Z(n13937) );
  NAND U12224 ( .A(n9649), .B(n9648), .Z(n13939) );
  ANDN U12225 ( .B(n9653), .A(n9652), .Z(n9654) );
  ANDN U12226 ( .B(n9662), .A(n9661), .Z(n13966) );
  ANDN U12227 ( .B(n9664), .A(n9663), .Z(n13969) );
  AND U12228 ( .A(n9669), .B(n13996), .Z(n9670) );
  ANDN U12229 ( .B(n9680), .A(n9679), .Z(n14019) );
  ANDN U12230 ( .B(n9682), .A(n9681), .Z(n14021) );
  ANDN U12231 ( .B(n9688), .A(n9687), .Z(n14041) );
  NANDN U12232 ( .A(n14046), .B(n9689), .Z(n9692) );
  AND U12233 ( .A(n9690), .B(n14049), .Z(n9691) );
  NAND U12234 ( .A(n9692), .B(n9691), .Z(n9693) );
  NANDN U12235 ( .A(n9694), .B(n9693), .Z(n9695) );
  OR U12236 ( .A(n14051), .B(n9695), .Z(n9696) );
  AND U12237 ( .A(n9697), .B(n9696), .Z(n9698) );
  NANDN U12238 ( .A(n9699), .B(n9698), .Z(n9700) );
  AND U12239 ( .A(n9701), .B(n9700), .Z(n9702) );
  OR U12240 ( .A(n9703), .B(n9702), .Z(n9704) );
  NAND U12241 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND U12242 ( .A(n9707), .B(n9706), .Z(n9709) );
  AND U12243 ( .A(n9709), .B(n9708), .Z(n9710) );
  NAND U12244 ( .A(n9711), .B(n9710), .Z(n9712) );
  NAND U12245 ( .A(n9713), .B(n9712), .Z(n9714) );
  AND U12246 ( .A(n9715), .B(n9714), .Z(n9716) );
  ANDN U12247 ( .B(n9717), .A(n9716), .Z(n9720) );
  ANDN U12248 ( .B(n9719), .A(n9718), .Z(n10179) );
  NANDN U12249 ( .A(n9720), .B(n10179), .Z(n9721) );
  NAND U12250 ( .A(n9722), .B(n9721), .Z(n9723) );
  NANDN U12251 ( .A(n9724), .B(n9723), .Z(n9725) );
  OR U12252 ( .A(n14075), .B(n9725), .Z(n9726) );
  AND U12253 ( .A(n9727), .B(n9726), .Z(n9729) );
  NAND U12254 ( .A(n9729), .B(n9728), .Z(n9731) );
  ANDN U12255 ( .B(n9731), .A(n9730), .Z(n9732) );
  NANDN U12256 ( .A(n9733), .B(n9732), .Z(n9736) );
  ANDN U12257 ( .B(n9734), .A(n14085), .Z(n9735) );
  NAND U12258 ( .A(n9736), .B(n9735), .Z(n9737) );
  NANDN U12259 ( .A(n9738), .B(n9737), .Z(n9739) );
  NANDN U12260 ( .A(n9739), .B(n14087), .Z(n9740) );
  AND U12261 ( .A(n14089), .B(n9740), .Z(n9741) );
  OR U12262 ( .A(n14091), .B(n9741), .Z(n9742) );
  NAND U12263 ( .A(n14093), .B(n9742), .Z(n9743) );
  NANDN U12264 ( .A(n14095), .B(n9743), .Z(n9746) );
  ANDN U12265 ( .B(n9744), .A(n14097), .Z(n9745) );
  NAND U12266 ( .A(n9746), .B(n9745), .Z(n9747) );
  AND U12267 ( .A(n9759), .B(n9758), .Z(n9761) );
  IV U12268 ( .A(n14124), .Z(n9760) );
  NANDN U12269 ( .A(n9761), .B(n9760), .Z(n9762) );
  AND U12270 ( .A(n9763), .B(n9762), .Z(n9764) );
  OR U12271 ( .A(n9765), .B(n9764), .Z(n9766) );
  NAND U12272 ( .A(n9767), .B(n9766), .Z(n9768) );
  NANDN U12273 ( .A(n9769), .B(n9768), .Z(n9770) );
  OR U12274 ( .A(n9771), .B(n9770), .Z(n9772) );
  AND U12275 ( .A(n9773), .B(n9772), .Z(n9774) );
  NANDN U12276 ( .A(n9775), .B(n9774), .Z(n9776) );
  AND U12277 ( .A(n9777), .B(n9776), .Z(n9778) );
  OR U12278 ( .A(n9779), .B(n9778), .Z(n9780) );
  NANDN U12279 ( .A(n9781), .B(n9780), .Z(n9782) );
  NAND U12280 ( .A(n14143), .B(n9782), .Z(n9785) );
  ANDN U12281 ( .B(n9783), .A(n14144), .Z(n9784) );
  NAND U12282 ( .A(n9785), .B(n9784), .Z(n9786) );
  NAND U12283 ( .A(n14146), .B(n9786), .Z(n9787) );
  OR U12284 ( .A(n9788), .B(n9787), .Z(n9789) );
  AND U12285 ( .A(n9790), .B(n9789), .Z(n9793) );
  NANDN U12286 ( .A(n9793), .B(x[1803]), .Z(n9792) );
  ANDN U12287 ( .B(n9792), .A(n9791), .Z(n9796) );
  XNOR U12288 ( .A(x[1803]), .B(n9793), .Z(n9794) );
  NANDN U12289 ( .A(y[1803]), .B(n9794), .Z(n9795) );
  NAND U12290 ( .A(n9796), .B(n9795), .Z(n9797) );
  AND U12291 ( .A(n14155), .B(n9797), .Z(n9798) );
  OR U12292 ( .A(n14156), .B(n9798), .Z(n9799) );
  NAND U12293 ( .A(n14159), .B(n9799), .Z(n9800) );
  NANDN U12294 ( .A(n14161), .B(n9800), .Z(n9801) );
  NAND U12295 ( .A(n9801), .B(n14163), .Z(n9802) );
  NANDN U12296 ( .A(n14165), .B(n9802), .Z(n9803) );
  AND U12297 ( .A(n14167), .B(n9803), .Z(n9806) );
  ANDN U12298 ( .B(n9805), .A(n9804), .Z(n14168) );
  NANDN U12299 ( .A(n9806), .B(n14168), .Z(n9807) );
  NAND U12300 ( .A(n9808), .B(n9807), .Z(n9809) );
  NANDN U12301 ( .A(n9810), .B(n9809), .Z(n9812) );
  NANDN U12302 ( .A(n9812), .B(n9811), .Z(n9813) );
  AND U12303 ( .A(n9822), .B(n9821), .Z(n14188) );
  ANDN U12304 ( .B(n9824), .A(n9823), .Z(n14191) );
  NAND U12305 ( .A(n9846), .B(n9845), .Z(n9847) );
  NANDN U12306 ( .A(n9848), .B(n9847), .Z(n9850) );
  OR U12307 ( .A(n9850), .B(n9849), .Z(n9851) );
  AND U12308 ( .A(n9852), .B(n9851), .Z(n9853) );
  OR U12309 ( .A(n9854), .B(n9853), .Z(n9855) );
  NAND U12310 ( .A(n9856), .B(n9855), .Z(n9860) );
  AND U12311 ( .A(n9858), .B(n9857), .Z(n9859) );
  NAND U12312 ( .A(n9860), .B(n9859), .Z(n9861) );
  NAND U12313 ( .A(n9862), .B(n9861), .Z(n9864) );
  OR U12314 ( .A(n9864), .B(n9863), .Z(n9865) );
  NAND U12315 ( .A(n9866), .B(n9865), .Z(n9867) );
  NAND U12316 ( .A(n9868), .B(n9867), .Z(n9871) );
  AND U12317 ( .A(n9869), .B(n14274), .Z(n9870) );
  NAND U12318 ( .A(n9871), .B(n9870), .Z(n9872) );
  NANDN U12319 ( .A(n9873), .B(n9872), .Z(n9875) );
  NANDN U12320 ( .A(n9875), .B(n9874), .Z(n9876) );
  AND U12321 ( .A(n9885), .B(n9884), .Z(n14292) );
  ANDN U12322 ( .B(n9887), .A(n9886), .Z(n14295) );
  AND U12323 ( .A(n9895), .B(n9894), .Z(n9899) );
  NAND U12324 ( .A(n9897), .B(n9896), .Z(n9898) );
  OR U12325 ( .A(n9899), .B(n9898), .Z(n9900) );
  AND U12326 ( .A(n9901), .B(n9900), .Z(n9902) );
  ANDN U12327 ( .B(n9903), .A(n9902), .Z(n9904) );
  NAND U12328 ( .A(n9905), .B(n9904), .Z(n9906) );
  NAND U12329 ( .A(n14319), .B(n9906), .Z(n9907) );
  OR U12330 ( .A(n9908), .B(n9907), .Z(n9909) );
  AND U12331 ( .A(n9910), .B(n9909), .Z(n9911) );
  NAND U12332 ( .A(n9912), .B(n9911), .Z(n9913) );
  AND U12333 ( .A(n14323), .B(n9913), .Z(n9914) );
  OR U12334 ( .A(n14325), .B(n9914), .Z(n9915) );
  NAND U12335 ( .A(n9916), .B(n9915), .Z(n9917) );
  NANDN U12336 ( .A(n9918), .B(n9917), .Z(n9919) );
  OR U12337 ( .A(n9919), .B(n14329), .Z(n9920) );
  AND U12338 ( .A(n9921), .B(n9920), .Z(n9923) );
  NAND U12339 ( .A(n9927), .B(n9926), .Z(n14347) );
  NAND U12340 ( .A(n9933), .B(n9932), .Z(n9934) );
  OR U12341 ( .A(n9935), .B(n9934), .Z(n9936) );
  AND U12342 ( .A(n9937), .B(n9936), .Z(n9941) );
  NAND U12343 ( .A(n9939), .B(n9938), .Z(n9940) );
  OR U12344 ( .A(n9941), .B(n9940), .Z(n9942) );
  AND U12345 ( .A(n9943), .B(n9942), .Z(n9944) );
  ANDN U12346 ( .B(n9945), .A(n9944), .Z(n9946) );
  NAND U12347 ( .A(n9947), .B(n9946), .Z(n9948) );
  NAND U12348 ( .A(n9949), .B(n9948), .Z(n9951) );
  OR U12349 ( .A(n9951), .B(n9950), .Z(n9952) );
  NAND U12350 ( .A(n9953), .B(n9952), .Z(n9954) );
  NAND U12351 ( .A(n14381), .B(n9954), .Z(n9958) );
  ANDN U12352 ( .B(n9956), .A(n9955), .Z(n9957) );
  NAND U12353 ( .A(n9958), .B(n9957), .Z(n9959) );
  NANDN U12354 ( .A(n9960), .B(n9959), .Z(n9961) );
  OR U12355 ( .A(n9962), .B(n9961), .Z(n9963) );
  AND U12356 ( .A(n9964), .B(n9963), .Z(n9965) );
  ANDN U12357 ( .B(n9974), .A(n9973), .Z(n14398) );
  NAND U12358 ( .A(n9976), .B(n9975), .Z(n14400) );
  IV U12359 ( .A(n14409), .Z(n9979) );
  NANDN U12360 ( .A(n9980), .B(n9979), .Z(n9981) );
  NAND U12361 ( .A(n9982), .B(n9981), .Z(n9983) );
  NANDN U12362 ( .A(n9984), .B(n9983), .Z(n9985) );
  NAND U12363 ( .A(n9986), .B(n9985), .Z(n9987) );
  NANDN U12364 ( .A(n9988), .B(n9987), .Z(n9989) );
  AND U12365 ( .A(n9990), .B(n9989), .Z(n9991) );
  NOR U12366 ( .A(n9992), .B(n9991), .Z(n9993) );
  NANDN U12367 ( .A(n9994), .B(n9993), .Z(n9995) );
  AND U12368 ( .A(n14427), .B(n9995), .Z(n9997) );
  NANDN U12369 ( .A(y[1918]), .B(x[1918]), .Z(n9996) );
  AND U12370 ( .A(n9997), .B(n9996), .Z(n9998) );
  OR U12371 ( .A(n14428), .B(n9998), .Z(n9999) );
  NAND U12372 ( .A(n14431), .B(n9999), .Z(n10000) );
  NANDN U12373 ( .A(n14433), .B(n10000), .Z(n10002) );
  OR U12374 ( .A(n10002), .B(n10001), .Z(n10003) );
  NAND U12375 ( .A(n10004), .B(n10003), .Z(n10005) );
  NANDN U12376 ( .A(n10006), .B(n10005), .Z(n10008) );
  OR U12377 ( .A(n10008), .B(n10007), .Z(n10009) );
  NAND U12378 ( .A(n10010), .B(n10009), .Z(n10014) );
  AND U12379 ( .A(n10012), .B(n10011), .Z(n10013) );
  NAND U12380 ( .A(n10014), .B(n10013), .Z(n10015) );
  NAND U12381 ( .A(n10016), .B(n10015), .Z(n10017) );
  OR U12382 ( .A(n10018), .B(n10017), .Z(n10019) );
  AND U12383 ( .A(n10020), .B(n10019), .Z(n10021) );
  NAND U12384 ( .A(n14449), .B(n10021), .Z(n10022) );
  AND U12385 ( .A(n14451), .B(n10022), .Z(n10023) );
  OR U12386 ( .A(n14453), .B(n10023), .Z(n10024) );
  NAND U12387 ( .A(n14455), .B(n10024), .Z(n10025) );
  NANDN U12388 ( .A(n14457), .B(n10025), .Z(n10028) );
  ANDN U12389 ( .B(n10026), .A(n14459), .Z(n10027) );
  NAND U12390 ( .A(n10028), .B(n10027), .Z(n10029) );
  NANDN U12391 ( .A(n10030), .B(n10029), .Z(n10031) );
  NANDN U12392 ( .A(n10031), .B(n14461), .Z(n10032) );
  AND U12393 ( .A(n10033), .B(n10032), .Z(n10037) );
  NAND U12394 ( .A(n10035), .B(n10034), .Z(n10036) );
  OR U12395 ( .A(n10037), .B(n10036), .Z(n10038) );
  AND U12396 ( .A(n10039), .B(n10038), .Z(n10040) );
  OR U12397 ( .A(n10041), .B(n10040), .Z(n10042) );
  NAND U12398 ( .A(n10043), .B(n10042), .Z(n10046) );
  ANDN U12399 ( .B(n10044), .A(n14476), .Z(n10045) );
  NAND U12400 ( .A(n10046), .B(n10045), .Z(n10047) );
  NANDN U12401 ( .A(n10048), .B(n10047), .Z(n10049) );
  NANDN U12402 ( .A(n10049), .B(n14478), .Z(n10050) );
  AND U12403 ( .A(n14481), .B(n10050), .Z(n10051) );
  OR U12404 ( .A(n14482), .B(n10051), .Z(n10052) );
  NAND U12405 ( .A(n10053), .B(n10052), .Z(n10054) );
  NANDN U12406 ( .A(n10055), .B(n10054), .Z(n10056) );
  NANDN U12407 ( .A(n10056), .B(n14486), .Z(n10057) );
  AND U12408 ( .A(n10058), .B(n10057), .Z(n10059) );
  OR U12409 ( .A(n10060), .B(n10059), .Z(n10061) );
  NAND U12410 ( .A(n10062), .B(n10061), .Z(n10063) );
  NANDN U12411 ( .A(n10064), .B(n10063), .Z(n10065) );
  OR U12412 ( .A(n10066), .B(n10065), .Z(n10067) );
  AND U12413 ( .A(n10068), .B(n10067), .Z(n10070) );
  NAND U12414 ( .A(n10070), .B(n10069), .Z(n10072) );
  ANDN U12415 ( .B(n10072), .A(n10071), .Z(n10073) );
  NANDN U12416 ( .A(n10074), .B(n10073), .Z(n10078) );
  ANDN U12417 ( .B(n10076), .A(n10075), .Z(n10077) );
  NAND U12418 ( .A(n10078), .B(n10077), .Z(n10079) );
  NANDN U12419 ( .A(n10080), .B(n10079), .Z(n10081) );
  OR U12420 ( .A(n10082), .B(n10081), .Z(n10084) );
  ANDN U12421 ( .B(n10084), .A(n10083), .Z(n10085) );
  NANDN U12422 ( .A(n10086), .B(n10085), .Z(n10087) );
  AND U12423 ( .A(n10088), .B(n10087), .Z(n10094) );
  OR U12424 ( .A(n10090), .B(n10089), .Z(n10092) );
  ANDN U12425 ( .B(n10092), .A(n10091), .Z(n10093) );
  NANDN U12426 ( .A(n10094), .B(n10093), .Z(n10095) );
  NANDN U12427 ( .A(n14518), .B(n10095), .Z(n10096) );
  NANDN U12428 ( .A(n10097), .B(n10096), .Z(n10098) );
  NANDN U12429 ( .A(x[1959]), .B(n10098), .Z(n10101) );
  XNOR U12430 ( .A(x[1959]), .B(n10098), .Z(n10099) );
  NAND U12431 ( .A(n10099), .B(y[1959]), .Z(n10100) );
  NAND U12432 ( .A(n10101), .B(n10100), .Z(n10102) );
  AND U12433 ( .A(n10103), .B(n10102), .Z(n10104) );
  OR U12434 ( .A(n14524), .B(n10104), .Z(n10105) );
  AND U12435 ( .A(n14527), .B(n10105), .Z(n10106) );
  NAND U12436 ( .A(n14531), .B(n10106), .Z(n10107) );
  AND U12437 ( .A(n10108), .B(n10107), .Z(n10111) );
  NANDN U12438 ( .A(n10110), .B(n10109), .Z(n14535) );
  OR U12439 ( .A(n10111), .B(n14535), .Z(n10112) );
  AND U12440 ( .A(n14537), .B(n10112), .Z(n10114) );
  XNOR U12441 ( .A(x[1966]), .B(y[1966]), .Z(n10113) );
  NAND U12442 ( .A(n10114), .B(n10113), .Z(n10115) );
  NANDN U12443 ( .A(n10116), .B(n10115), .Z(n10118) );
  ANDN U12444 ( .B(x[1966]), .A(y[1966]), .Z(n10117) );
  OR U12445 ( .A(n10118), .B(n10117), .Z(n10119) );
  NANDN U12446 ( .A(n14544), .B(n10119), .Z(n10120) );
  ANDN U12447 ( .B(n10123), .A(n10122), .Z(n14549) );
  NAND U12448 ( .A(n10125), .B(n10124), .Z(n14550) );
  AND U12449 ( .A(n10135), .B(n10134), .Z(n14583) );
  AND U12450 ( .A(n10143), .B(n10142), .Z(n14627) );
  ANDN U12451 ( .B(n10145), .A(n10144), .Z(n14629) );
  ANDN U12452 ( .B(n10152), .A(n10151), .Z(n14645) );
  AND U12453 ( .A(n10164), .B(n10163), .Z(n14687) );
  OR U12454 ( .A(n10167), .B(ebreg), .Z(n5) );
  OR U12455 ( .A(n10171), .B(n10170), .Z(n10173) );
  ANDN U12456 ( .B(n10173), .A(n10172), .Z(n14653) );
  AND U12457 ( .A(n10175), .B(n10174), .Z(n14619) );
  AND U12458 ( .A(n10177), .B(n10176), .Z(n14137) );
  OR U12459 ( .A(n10179), .B(n10178), .Z(n14073) );
  OR U12460 ( .A(n10181), .B(n10180), .Z(n10183) );
  ANDN U12461 ( .B(n10183), .A(n10182), .Z(n13909) );
  ANDN U12462 ( .B(n10185), .A(n10184), .Z(n13905) );
  ANDN U12463 ( .B(n10187), .A(n10186), .Z(n13547) );
  NANDN U12464 ( .A(n10189), .B(n10188), .Z(n10191) );
  ANDN U12465 ( .B(n10191), .A(n10190), .Z(n12597) );
  NAND U12466 ( .A(n10193), .B(n10192), .Z(n10194) );
  NANDN U12467 ( .A(n10195), .B(n10194), .Z(n10196) );
  AND U12468 ( .A(n10197), .B(n10196), .Z(n10198) );
  OR U12469 ( .A(n10199), .B(n10198), .Z(n10200) );
  NAND U12470 ( .A(n10201), .B(n10200), .Z(n10202) );
  NANDN U12471 ( .A(n10203), .B(n10202), .Z(n10204) );
  NAND U12472 ( .A(n10205), .B(n10204), .Z(n10206) );
  NANDN U12473 ( .A(n10207), .B(n10206), .Z(n10208) );
  AND U12474 ( .A(n10209), .B(n10208), .Z(n10210) );
  OR U12475 ( .A(n10211), .B(n10210), .Z(n10212) );
  NAND U12476 ( .A(n10213), .B(n10212), .Z(n10214) );
  NANDN U12477 ( .A(n10215), .B(n10214), .Z(n10216) );
  NAND U12478 ( .A(n10217), .B(n10216), .Z(n10218) );
  NANDN U12479 ( .A(n10219), .B(n10218), .Z(n10220) );
  AND U12480 ( .A(n10221), .B(n10220), .Z(n10222) );
  OR U12481 ( .A(n10223), .B(n10222), .Z(n10224) );
  NAND U12482 ( .A(n10225), .B(n10224), .Z(n10226) );
  NANDN U12483 ( .A(n10227), .B(n10226), .Z(n10228) );
  NAND U12484 ( .A(n10229), .B(n10228), .Z(n10230) );
  NANDN U12485 ( .A(n10231), .B(n10230), .Z(n10232) );
  AND U12486 ( .A(n10233), .B(n10232), .Z(n10234) );
  OR U12487 ( .A(n10235), .B(n10234), .Z(n10236) );
  NAND U12488 ( .A(n10237), .B(n10236), .Z(n10238) );
  NANDN U12489 ( .A(n10239), .B(n10238), .Z(n10240) );
  NAND U12490 ( .A(n10241), .B(n10240), .Z(n10242) );
  NANDN U12491 ( .A(n10243), .B(n10242), .Z(n10244) );
  AND U12492 ( .A(n10245), .B(n10244), .Z(n10246) );
  OR U12493 ( .A(n10247), .B(n10246), .Z(n10248) );
  NAND U12494 ( .A(n10249), .B(n10248), .Z(n10250) );
  NANDN U12495 ( .A(n10251), .B(n10250), .Z(n10252) );
  NAND U12496 ( .A(n10253), .B(n10252), .Z(n10254) );
  NANDN U12497 ( .A(n10255), .B(n10254), .Z(n10256) );
  AND U12498 ( .A(n10257), .B(n10256), .Z(n10258) );
  OR U12499 ( .A(n10259), .B(n10258), .Z(n10260) );
  NAND U12500 ( .A(n10261), .B(n10260), .Z(n10262) );
  NANDN U12501 ( .A(n10263), .B(n10262), .Z(n10264) );
  NAND U12502 ( .A(n10265), .B(n10264), .Z(n10266) );
  NANDN U12503 ( .A(n10267), .B(n10266), .Z(n10268) );
  AND U12504 ( .A(n10269), .B(n10268), .Z(n10270) );
  OR U12505 ( .A(n10271), .B(n10270), .Z(n10272) );
  NAND U12506 ( .A(n10273), .B(n10272), .Z(n10274) );
  NANDN U12507 ( .A(n10275), .B(n10274), .Z(n10276) );
  NAND U12508 ( .A(n10277), .B(n10276), .Z(n10278) );
  NANDN U12509 ( .A(n10279), .B(n10278), .Z(n10280) );
  AND U12510 ( .A(n10281), .B(n10280), .Z(n10282) );
  OR U12511 ( .A(n10283), .B(n10282), .Z(n10284) );
  NAND U12512 ( .A(n10285), .B(n10284), .Z(n10286) );
  NANDN U12513 ( .A(n10287), .B(n10286), .Z(n10288) );
  NAND U12514 ( .A(n10289), .B(n10288), .Z(n10290) );
  NANDN U12515 ( .A(n10291), .B(n10290), .Z(n10292) );
  AND U12516 ( .A(n10293), .B(n10292), .Z(n10294) );
  OR U12517 ( .A(n10295), .B(n10294), .Z(n10296) );
  NAND U12518 ( .A(n10297), .B(n10296), .Z(n10298) );
  NANDN U12519 ( .A(n10299), .B(n10298), .Z(n10300) );
  NAND U12520 ( .A(n10301), .B(n10300), .Z(n10302) );
  NANDN U12521 ( .A(n10303), .B(n10302), .Z(n10304) );
  AND U12522 ( .A(n10305), .B(n10304), .Z(n10306) );
  OR U12523 ( .A(n10307), .B(n10306), .Z(n10308) );
  NAND U12524 ( .A(n10309), .B(n10308), .Z(n10310) );
  NANDN U12525 ( .A(n10311), .B(n10310), .Z(n10312) );
  NAND U12526 ( .A(n10313), .B(n10312), .Z(n10314) );
  NANDN U12527 ( .A(n10315), .B(n10314), .Z(n10316) );
  AND U12528 ( .A(n10317), .B(n10316), .Z(n10318) );
  OR U12529 ( .A(n10319), .B(n10318), .Z(n10320) );
  NAND U12530 ( .A(n10321), .B(n10320), .Z(n10322) );
  NANDN U12531 ( .A(n10323), .B(n10322), .Z(n10324) );
  NAND U12532 ( .A(n10325), .B(n10324), .Z(n10326) );
  NANDN U12533 ( .A(n10327), .B(n10326), .Z(n10328) );
  AND U12534 ( .A(n10329), .B(n10328), .Z(n10330) );
  OR U12535 ( .A(n10331), .B(n10330), .Z(n10332) );
  NAND U12536 ( .A(n10333), .B(n10332), .Z(n10334) );
  NANDN U12537 ( .A(n10335), .B(n10334), .Z(n10336) );
  NAND U12538 ( .A(n10337), .B(n10336), .Z(n10338) );
  NANDN U12539 ( .A(n10339), .B(n10338), .Z(n10340) );
  AND U12540 ( .A(n10341), .B(n10340), .Z(n10342) );
  OR U12541 ( .A(n10343), .B(n10342), .Z(n10344) );
  NAND U12542 ( .A(n10345), .B(n10344), .Z(n10346) );
  NANDN U12543 ( .A(n10347), .B(n10346), .Z(n10348) );
  NAND U12544 ( .A(n10349), .B(n10348), .Z(n10350) );
  NANDN U12545 ( .A(n10351), .B(n10350), .Z(n10352) );
  AND U12546 ( .A(n10353), .B(n10352), .Z(n10354) );
  OR U12547 ( .A(n10355), .B(n10354), .Z(n10356) );
  NAND U12548 ( .A(n10357), .B(n10356), .Z(n10358) );
  NANDN U12549 ( .A(n10359), .B(n10358), .Z(n10360) );
  NAND U12550 ( .A(n10361), .B(n10360), .Z(n10362) );
  NANDN U12551 ( .A(n10363), .B(n10362), .Z(n10364) );
  AND U12552 ( .A(n10365), .B(n10364), .Z(n10366) );
  OR U12553 ( .A(n10367), .B(n10366), .Z(n10368) );
  NAND U12554 ( .A(n10369), .B(n10368), .Z(n10370) );
  NANDN U12555 ( .A(n10371), .B(n10370), .Z(n10372) );
  NAND U12556 ( .A(n10373), .B(n10372), .Z(n10374) );
  NANDN U12557 ( .A(n10375), .B(n10374), .Z(n10376) );
  AND U12558 ( .A(n10377), .B(n10376), .Z(n10378) );
  OR U12559 ( .A(n10379), .B(n10378), .Z(n10380) );
  NAND U12560 ( .A(n10381), .B(n10380), .Z(n10382) );
  NANDN U12561 ( .A(n10383), .B(n10382), .Z(n10384) );
  NAND U12562 ( .A(n10385), .B(n10384), .Z(n10386) );
  NANDN U12563 ( .A(n10387), .B(n10386), .Z(n10388) );
  AND U12564 ( .A(n10389), .B(n10388), .Z(n10390) );
  OR U12565 ( .A(n10391), .B(n10390), .Z(n10392) );
  NAND U12566 ( .A(n10393), .B(n10392), .Z(n10394) );
  NANDN U12567 ( .A(n10395), .B(n10394), .Z(n10396) );
  NAND U12568 ( .A(n10397), .B(n10396), .Z(n10398) );
  NANDN U12569 ( .A(n10399), .B(n10398), .Z(n10400) );
  AND U12570 ( .A(n10401), .B(n10400), .Z(n10402) );
  OR U12571 ( .A(n10403), .B(n10402), .Z(n10404) );
  NAND U12572 ( .A(n10405), .B(n10404), .Z(n10406) );
  NANDN U12573 ( .A(n10407), .B(n10406), .Z(n10408) );
  NAND U12574 ( .A(n10409), .B(n10408), .Z(n10410) );
  NANDN U12575 ( .A(n10411), .B(n10410), .Z(n10412) );
  AND U12576 ( .A(n10413), .B(n10412), .Z(n10414) );
  OR U12577 ( .A(n10415), .B(n10414), .Z(n10416) );
  NAND U12578 ( .A(n10417), .B(n10416), .Z(n10418) );
  NANDN U12579 ( .A(n10419), .B(n10418), .Z(n10420) );
  NAND U12580 ( .A(n10421), .B(n10420), .Z(n10422) );
  NANDN U12581 ( .A(n10423), .B(n10422), .Z(n10424) );
  AND U12582 ( .A(n10425), .B(n10424), .Z(n10426) );
  OR U12583 ( .A(n10427), .B(n10426), .Z(n10428) );
  NAND U12584 ( .A(n10429), .B(n10428), .Z(n10430) );
  NANDN U12585 ( .A(n10431), .B(n10430), .Z(n10432) );
  NAND U12586 ( .A(n10433), .B(n10432), .Z(n10434) );
  NANDN U12587 ( .A(n10435), .B(n10434), .Z(n10436) );
  AND U12588 ( .A(n10437), .B(n10436), .Z(n10438) );
  OR U12589 ( .A(n10439), .B(n10438), .Z(n10440) );
  NAND U12590 ( .A(n10441), .B(n10440), .Z(n10442) );
  NANDN U12591 ( .A(n10443), .B(n10442), .Z(n10444) );
  NAND U12592 ( .A(n10445), .B(n10444), .Z(n10446) );
  NANDN U12593 ( .A(n10447), .B(n10446), .Z(n10448) );
  AND U12594 ( .A(n10449), .B(n10448), .Z(n10450) );
  OR U12595 ( .A(n10451), .B(n10450), .Z(n10452) );
  NAND U12596 ( .A(n10453), .B(n10452), .Z(n10454) );
  NANDN U12597 ( .A(n10455), .B(n10454), .Z(n10456) );
  NAND U12598 ( .A(n10457), .B(n10456), .Z(n10458) );
  NANDN U12599 ( .A(n10459), .B(n10458), .Z(n10460) );
  AND U12600 ( .A(n10461), .B(n10460), .Z(n10462) );
  OR U12601 ( .A(n10463), .B(n10462), .Z(n10464) );
  NAND U12602 ( .A(n10465), .B(n10464), .Z(n10466) );
  NANDN U12603 ( .A(n10467), .B(n10466), .Z(n10468) );
  NAND U12604 ( .A(n10469), .B(n10468), .Z(n10470) );
  NANDN U12605 ( .A(n10471), .B(n10470), .Z(n10472) );
  AND U12606 ( .A(n10473), .B(n10472), .Z(n10474) );
  OR U12607 ( .A(n10475), .B(n10474), .Z(n10476) );
  NAND U12608 ( .A(n10477), .B(n10476), .Z(n10478) );
  NANDN U12609 ( .A(n10479), .B(n10478), .Z(n10480) );
  NAND U12610 ( .A(n10481), .B(n10480), .Z(n10482) );
  NANDN U12611 ( .A(n10483), .B(n10482), .Z(n10484) );
  AND U12612 ( .A(n10485), .B(n10484), .Z(n10487) );
  NANDN U12613 ( .A(n10487), .B(n10486), .Z(n10488) );
  NANDN U12614 ( .A(n10489), .B(n10488), .Z(n10490) );
  NANDN U12615 ( .A(n10491), .B(n10490), .Z(n10492) );
  NAND U12616 ( .A(n10493), .B(n10492), .Z(n10494) );
  NANDN U12617 ( .A(n10495), .B(n10494), .Z(n10496) );
  AND U12618 ( .A(n10497), .B(n10496), .Z(n10498) );
  OR U12619 ( .A(n10499), .B(n10498), .Z(n10500) );
  NAND U12620 ( .A(n10501), .B(n10500), .Z(n10502) );
  NANDN U12621 ( .A(n10503), .B(n10502), .Z(n10504) );
  NAND U12622 ( .A(n10505), .B(n10504), .Z(n10506) );
  NANDN U12623 ( .A(n10507), .B(n10506), .Z(n10508) );
  AND U12624 ( .A(n10509), .B(n10508), .Z(n10510) );
  OR U12625 ( .A(n10511), .B(n10510), .Z(n10512) );
  NAND U12626 ( .A(n10513), .B(n10512), .Z(n10514) );
  NANDN U12627 ( .A(n10515), .B(n10514), .Z(n10516) );
  NAND U12628 ( .A(n10517), .B(n10516), .Z(n10518) );
  NANDN U12629 ( .A(n10519), .B(n10518), .Z(n10520) );
  AND U12630 ( .A(n10521), .B(n10520), .Z(n10522) );
  OR U12631 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U12632 ( .A(n10525), .B(n10524), .Z(n10526) );
  NANDN U12633 ( .A(n10527), .B(n10526), .Z(n10528) );
  NAND U12634 ( .A(n10529), .B(n10528), .Z(n10530) );
  NANDN U12635 ( .A(n10531), .B(n10530), .Z(n10532) );
  AND U12636 ( .A(n10533), .B(n10532), .Z(n10534) );
  OR U12637 ( .A(n10535), .B(n10534), .Z(n10536) );
  NAND U12638 ( .A(n10537), .B(n10536), .Z(n10538) );
  NANDN U12639 ( .A(n10539), .B(n10538), .Z(n10540) );
  NAND U12640 ( .A(n10541), .B(n10540), .Z(n10542) );
  NANDN U12641 ( .A(n10543), .B(n10542), .Z(n10544) );
  AND U12642 ( .A(n10545), .B(n10544), .Z(n10546) );
  OR U12643 ( .A(n10547), .B(n10546), .Z(n10548) );
  NAND U12644 ( .A(n10549), .B(n10548), .Z(n10550) );
  NANDN U12645 ( .A(n10551), .B(n10550), .Z(n10552) );
  NAND U12646 ( .A(n10553), .B(n10552), .Z(n10554) );
  NANDN U12647 ( .A(n10555), .B(n10554), .Z(n10556) );
  AND U12648 ( .A(n10557), .B(n10556), .Z(n10558) );
  OR U12649 ( .A(n10559), .B(n10558), .Z(n10560) );
  NAND U12650 ( .A(n10561), .B(n10560), .Z(n10562) );
  NANDN U12651 ( .A(n10563), .B(n10562), .Z(n10564) );
  NAND U12652 ( .A(n10565), .B(n10564), .Z(n10566) );
  NANDN U12653 ( .A(n10567), .B(n10566), .Z(n10568) );
  AND U12654 ( .A(n10569), .B(n10568), .Z(n10570) );
  OR U12655 ( .A(n10571), .B(n10570), .Z(n10572) );
  NAND U12656 ( .A(n10573), .B(n10572), .Z(n10574) );
  NANDN U12657 ( .A(n10575), .B(n10574), .Z(n10576) );
  NAND U12658 ( .A(n10577), .B(n10576), .Z(n10578) );
  NANDN U12659 ( .A(n10579), .B(n10578), .Z(n10580) );
  AND U12660 ( .A(n10581), .B(n10580), .Z(n10582) );
  OR U12661 ( .A(n10583), .B(n10582), .Z(n10584) );
  NAND U12662 ( .A(n10585), .B(n10584), .Z(n10586) );
  NANDN U12663 ( .A(n10587), .B(n10586), .Z(n10588) );
  NAND U12664 ( .A(n10589), .B(n10588), .Z(n10590) );
  NANDN U12665 ( .A(n10591), .B(n10590), .Z(n10592) );
  AND U12666 ( .A(n10593), .B(n10592), .Z(n10594) );
  OR U12667 ( .A(n10595), .B(n10594), .Z(n10596) );
  NAND U12668 ( .A(n10597), .B(n10596), .Z(n10598) );
  NANDN U12669 ( .A(n10599), .B(n10598), .Z(n10600) );
  NAND U12670 ( .A(n10601), .B(n10600), .Z(n10602) );
  NANDN U12671 ( .A(n10603), .B(n10602), .Z(n10604) );
  AND U12672 ( .A(n10605), .B(n10604), .Z(n10606) );
  OR U12673 ( .A(n10607), .B(n10606), .Z(n10608) );
  NAND U12674 ( .A(n10609), .B(n10608), .Z(n10610) );
  NANDN U12675 ( .A(n10611), .B(n10610), .Z(n10612) );
  NAND U12676 ( .A(n10613), .B(n10612), .Z(n10614) );
  NANDN U12677 ( .A(n10615), .B(n10614), .Z(n10616) );
  AND U12678 ( .A(n10617), .B(n10616), .Z(n10618) );
  OR U12679 ( .A(n10619), .B(n10618), .Z(n10620) );
  NAND U12680 ( .A(n10621), .B(n10620), .Z(n10622) );
  NANDN U12681 ( .A(n10623), .B(n10622), .Z(n10624) );
  NAND U12682 ( .A(n10625), .B(n10624), .Z(n10626) );
  NANDN U12683 ( .A(n10627), .B(n10626), .Z(n10628) );
  AND U12684 ( .A(n10629), .B(n10628), .Z(n10630) );
  OR U12685 ( .A(n10631), .B(n10630), .Z(n10632) );
  NAND U12686 ( .A(n10633), .B(n10632), .Z(n10634) );
  NANDN U12687 ( .A(n10635), .B(n10634), .Z(n10636) );
  NAND U12688 ( .A(n10637), .B(n10636), .Z(n10638) );
  NANDN U12689 ( .A(n10639), .B(n10638), .Z(n10640) );
  AND U12690 ( .A(n10641), .B(n10640), .Z(n10642) );
  OR U12691 ( .A(n10643), .B(n10642), .Z(n10644) );
  NAND U12692 ( .A(n10645), .B(n10644), .Z(n10646) );
  NANDN U12693 ( .A(n10647), .B(n10646), .Z(n10648) );
  NAND U12694 ( .A(n10649), .B(n10648), .Z(n10650) );
  NANDN U12695 ( .A(n10651), .B(n10650), .Z(n10652) );
  AND U12696 ( .A(n10653), .B(n10652), .Z(n10654) );
  OR U12697 ( .A(n10655), .B(n10654), .Z(n10656) );
  NAND U12698 ( .A(n10657), .B(n10656), .Z(n10658) );
  NANDN U12699 ( .A(n10659), .B(n10658), .Z(n10660) );
  NAND U12700 ( .A(n10661), .B(n10660), .Z(n10662) );
  NANDN U12701 ( .A(n10663), .B(n10662), .Z(n10664) );
  AND U12702 ( .A(n10665), .B(n10664), .Z(n10666) );
  OR U12703 ( .A(n10667), .B(n10666), .Z(n10668) );
  NAND U12704 ( .A(n10669), .B(n10668), .Z(n10670) );
  NANDN U12705 ( .A(n10671), .B(n10670), .Z(n10672) );
  NAND U12706 ( .A(n10673), .B(n10672), .Z(n10674) );
  NANDN U12707 ( .A(n10675), .B(n10674), .Z(n10676) );
  AND U12708 ( .A(n10677), .B(n10676), .Z(n10678) );
  OR U12709 ( .A(n10679), .B(n10678), .Z(n10680) );
  NAND U12710 ( .A(n10681), .B(n10680), .Z(n10682) );
  NANDN U12711 ( .A(n10683), .B(n10682), .Z(n10684) );
  NAND U12712 ( .A(n10685), .B(n10684), .Z(n10686) );
  NANDN U12713 ( .A(n10687), .B(n10686), .Z(n10688) );
  AND U12714 ( .A(n10689), .B(n10688), .Z(n10690) );
  OR U12715 ( .A(n10691), .B(n10690), .Z(n10692) );
  NAND U12716 ( .A(n10693), .B(n10692), .Z(n10694) );
  NANDN U12717 ( .A(n10695), .B(n10694), .Z(n10696) );
  NAND U12718 ( .A(n10697), .B(n10696), .Z(n10698) );
  NANDN U12719 ( .A(n10699), .B(n10698), .Z(n10700) );
  AND U12720 ( .A(n10701), .B(n10700), .Z(n10702) );
  OR U12721 ( .A(n10703), .B(n10702), .Z(n10704) );
  NAND U12722 ( .A(n10705), .B(n10704), .Z(n10706) );
  NANDN U12723 ( .A(n10707), .B(n10706), .Z(n10708) );
  NAND U12724 ( .A(n10709), .B(n10708), .Z(n10710) );
  NANDN U12725 ( .A(n10711), .B(n10710), .Z(n10712) );
  AND U12726 ( .A(n10713), .B(n10712), .Z(n10714) );
  OR U12727 ( .A(n10715), .B(n10714), .Z(n10716) );
  NAND U12728 ( .A(n10717), .B(n10716), .Z(n10718) );
  NANDN U12729 ( .A(n10719), .B(n10718), .Z(n10720) );
  NAND U12730 ( .A(n10721), .B(n10720), .Z(n10722) );
  NANDN U12731 ( .A(n10723), .B(n10722), .Z(n10724) );
  AND U12732 ( .A(n10725), .B(n10724), .Z(n10726) );
  OR U12733 ( .A(n10727), .B(n10726), .Z(n10728) );
  NAND U12734 ( .A(n10729), .B(n10728), .Z(n10730) );
  NANDN U12735 ( .A(n10731), .B(n10730), .Z(n10732) );
  NAND U12736 ( .A(n10733), .B(n10732), .Z(n10734) );
  NANDN U12737 ( .A(n10735), .B(n10734), .Z(n10736) );
  AND U12738 ( .A(n10737), .B(n10736), .Z(n10741) );
  ANDN U12739 ( .B(n10739), .A(n10738), .Z(n10740) );
  NANDN U12740 ( .A(n10741), .B(n10740), .Z(n10742) );
  AND U12741 ( .A(n10743), .B(n10742), .Z(n10744) );
  OR U12742 ( .A(n10745), .B(n10744), .Z(n10746) );
  NAND U12743 ( .A(n10747), .B(n10746), .Z(n10748) );
  NANDN U12744 ( .A(n10749), .B(n10748), .Z(n10750) );
  NAND U12745 ( .A(n10751), .B(n10750), .Z(n10752) );
  NANDN U12746 ( .A(n10753), .B(n10752), .Z(n10754) );
  AND U12747 ( .A(n10755), .B(n10754), .Z(n10756) );
  OR U12748 ( .A(n10757), .B(n10756), .Z(n10758) );
  NAND U12749 ( .A(n10759), .B(n10758), .Z(n10760) );
  NANDN U12750 ( .A(n10761), .B(n10760), .Z(n10762) );
  NAND U12751 ( .A(n10763), .B(n10762), .Z(n10764) );
  NANDN U12752 ( .A(n10765), .B(n10764), .Z(n10766) );
  AND U12753 ( .A(n10767), .B(n10766), .Z(n10768) );
  OR U12754 ( .A(n10769), .B(n10768), .Z(n10770) );
  NAND U12755 ( .A(n10771), .B(n10770), .Z(n10772) );
  NANDN U12756 ( .A(n10773), .B(n10772), .Z(n10774) );
  NAND U12757 ( .A(n10775), .B(n10774), .Z(n10776) );
  NANDN U12758 ( .A(n10777), .B(n10776), .Z(n10778) );
  AND U12759 ( .A(n10779), .B(n10778), .Z(n10780) );
  OR U12760 ( .A(n10781), .B(n10780), .Z(n10782) );
  NAND U12761 ( .A(n10783), .B(n10782), .Z(n10784) );
  NANDN U12762 ( .A(n10785), .B(n10784), .Z(n10786) );
  NAND U12763 ( .A(n10787), .B(n10786), .Z(n10788) );
  NANDN U12764 ( .A(n10789), .B(n10788), .Z(n10790) );
  AND U12765 ( .A(n10791), .B(n10790), .Z(n10792) );
  OR U12766 ( .A(n10793), .B(n10792), .Z(n10794) );
  NAND U12767 ( .A(n10795), .B(n10794), .Z(n10796) );
  NANDN U12768 ( .A(n10797), .B(n10796), .Z(n10798) );
  NAND U12769 ( .A(n10799), .B(n10798), .Z(n10800) );
  NANDN U12770 ( .A(n10801), .B(n10800), .Z(n10802) );
  AND U12771 ( .A(n10803), .B(n10802), .Z(n10804) );
  OR U12772 ( .A(n10805), .B(n10804), .Z(n10806) );
  NAND U12773 ( .A(n10807), .B(n10806), .Z(n10808) );
  NANDN U12774 ( .A(n10809), .B(n10808), .Z(n10810) );
  NAND U12775 ( .A(n10811), .B(n10810), .Z(n10812) );
  NANDN U12776 ( .A(n10813), .B(n10812), .Z(n10814) );
  AND U12777 ( .A(n10815), .B(n10814), .Z(n10816) );
  OR U12778 ( .A(n10817), .B(n10816), .Z(n10818) );
  NAND U12779 ( .A(n10819), .B(n10818), .Z(n10820) );
  NANDN U12780 ( .A(n10821), .B(n10820), .Z(n10822) );
  NAND U12781 ( .A(n10823), .B(n10822), .Z(n10824) );
  NANDN U12782 ( .A(n10825), .B(n10824), .Z(n10826) );
  AND U12783 ( .A(n10827), .B(n10826), .Z(n10828) );
  OR U12784 ( .A(n10829), .B(n10828), .Z(n10830) );
  NAND U12785 ( .A(n10831), .B(n10830), .Z(n10832) );
  NANDN U12786 ( .A(n10833), .B(n10832), .Z(n10834) );
  NAND U12787 ( .A(n10835), .B(n10834), .Z(n10836) );
  NANDN U12788 ( .A(n10837), .B(n10836), .Z(n10838) );
  AND U12789 ( .A(n10839), .B(n10838), .Z(n10840) );
  OR U12790 ( .A(n10841), .B(n10840), .Z(n10842) );
  NAND U12791 ( .A(n10843), .B(n10842), .Z(n10844) );
  NANDN U12792 ( .A(n10845), .B(n10844), .Z(n10846) );
  NAND U12793 ( .A(n10847), .B(n10846), .Z(n10848) );
  NANDN U12794 ( .A(n10849), .B(n10848), .Z(n10850) );
  AND U12795 ( .A(n10851), .B(n10850), .Z(n10852) );
  OR U12796 ( .A(n10853), .B(n10852), .Z(n10854) );
  NAND U12797 ( .A(n10855), .B(n10854), .Z(n10856) );
  NANDN U12798 ( .A(n10857), .B(n10856), .Z(n10858) );
  NAND U12799 ( .A(n10859), .B(n10858), .Z(n10860) );
  NANDN U12800 ( .A(n10861), .B(n10860), .Z(n10862) );
  AND U12801 ( .A(n10863), .B(n10862), .Z(n10864) );
  OR U12802 ( .A(n10865), .B(n10864), .Z(n10866) );
  NAND U12803 ( .A(n10867), .B(n10866), .Z(n10868) );
  NANDN U12804 ( .A(n10869), .B(n10868), .Z(n10870) );
  NAND U12805 ( .A(n10871), .B(n10870), .Z(n10872) );
  NANDN U12806 ( .A(n10873), .B(n10872), .Z(n10874) );
  AND U12807 ( .A(n10875), .B(n10874), .Z(n10876) );
  OR U12808 ( .A(n10877), .B(n10876), .Z(n10878) );
  NAND U12809 ( .A(n10879), .B(n10878), .Z(n10880) );
  NANDN U12810 ( .A(n10881), .B(n10880), .Z(n10882) );
  NAND U12811 ( .A(n10883), .B(n10882), .Z(n10884) );
  NANDN U12812 ( .A(n10885), .B(n10884), .Z(n10886) );
  AND U12813 ( .A(n10887), .B(n10886), .Z(n10888) );
  OR U12814 ( .A(n10889), .B(n10888), .Z(n10890) );
  NAND U12815 ( .A(n10891), .B(n10890), .Z(n10892) );
  NANDN U12816 ( .A(n10893), .B(n10892), .Z(n10894) );
  NAND U12817 ( .A(n10895), .B(n10894), .Z(n10896) );
  NANDN U12818 ( .A(n10897), .B(n10896), .Z(n10898) );
  AND U12819 ( .A(n10899), .B(n10898), .Z(n10900) );
  OR U12820 ( .A(n10901), .B(n10900), .Z(n10902) );
  NAND U12821 ( .A(n10903), .B(n10902), .Z(n10904) );
  NANDN U12822 ( .A(n10905), .B(n10904), .Z(n10906) );
  NAND U12823 ( .A(n10907), .B(n10906), .Z(n10908) );
  NANDN U12824 ( .A(n10909), .B(n10908), .Z(n10910) );
  AND U12825 ( .A(n10911), .B(n10910), .Z(n10912) );
  OR U12826 ( .A(n10913), .B(n10912), .Z(n10914) );
  NAND U12827 ( .A(n10915), .B(n10914), .Z(n10916) );
  NANDN U12828 ( .A(n10917), .B(n10916), .Z(n10918) );
  NAND U12829 ( .A(n10919), .B(n10918), .Z(n10920) );
  NANDN U12830 ( .A(n10921), .B(n10920), .Z(n10922) );
  AND U12831 ( .A(n10923), .B(n10922), .Z(n10924) );
  OR U12832 ( .A(n10925), .B(n10924), .Z(n10926) );
  NAND U12833 ( .A(n10927), .B(n10926), .Z(n10928) );
  NANDN U12834 ( .A(n10929), .B(n10928), .Z(n10930) );
  NAND U12835 ( .A(n10931), .B(n10930), .Z(n10932) );
  NANDN U12836 ( .A(n10933), .B(n10932), .Z(n10934) );
  AND U12837 ( .A(n10935), .B(n10934), .Z(n10936) );
  OR U12838 ( .A(n10937), .B(n10936), .Z(n10938) );
  NAND U12839 ( .A(n10939), .B(n10938), .Z(n10940) );
  NANDN U12840 ( .A(n10941), .B(n10940), .Z(n10942) );
  NAND U12841 ( .A(n10943), .B(n10942), .Z(n10944) );
  NANDN U12842 ( .A(n10945), .B(n10944), .Z(n10946) );
  AND U12843 ( .A(n10947), .B(n10946), .Z(n10948) );
  OR U12844 ( .A(n10949), .B(n10948), .Z(n10950) );
  NAND U12845 ( .A(n10951), .B(n10950), .Z(n10952) );
  NANDN U12846 ( .A(n10953), .B(n10952), .Z(n10954) );
  NAND U12847 ( .A(n10955), .B(n10954), .Z(n10956) );
  NANDN U12848 ( .A(n10957), .B(n10956), .Z(n10958) );
  AND U12849 ( .A(n10959), .B(n10958), .Z(n10960) );
  OR U12850 ( .A(n10961), .B(n10960), .Z(n10962) );
  NAND U12851 ( .A(n10963), .B(n10962), .Z(n10964) );
  NANDN U12852 ( .A(n10965), .B(n10964), .Z(n10966) );
  NAND U12853 ( .A(n10967), .B(n10966), .Z(n10968) );
  NANDN U12854 ( .A(n10969), .B(n10968), .Z(n10970) );
  AND U12855 ( .A(n10971), .B(n10970), .Z(n10972) );
  OR U12856 ( .A(n10973), .B(n10972), .Z(n10974) );
  NAND U12857 ( .A(n10975), .B(n10974), .Z(n10976) );
  NANDN U12858 ( .A(n10977), .B(n10976), .Z(n10978) );
  NAND U12859 ( .A(n10979), .B(n10978), .Z(n10980) );
  NANDN U12860 ( .A(n10981), .B(n10980), .Z(n10982) );
  AND U12861 ( .A(n10983), .B(n10982), .Z(n10984) );
  OR U12862 ( .A(n10985), .B(n10984), .Z(n10986) );
  NAND U12863 ( .A(n10987), .B(n10986), .Z(n10988) );
  NANDN U12864 ( .A(n10989), .B(n10988), .Z(n10990) );
  NAND U12865 ( .A(n10991), .B(n10990), .Z(n10992) );
  NANDN U12866 ( .A(n10993), .B(n10992), .Z(n10994) );
  AND U12867 ( .A(n10995), .B(n10994), .Z(n10996) );
  OR U12868 ( .A(n10997), .B(n10996), .Z(n10998) );
  NAND U12869 ( .A(n10999), .B(n10998), .Z(n11000) );
  NANDN U12870 ( .A(n11001), .B(n11000), .Z(n11002) );
  NAND U12871 ( .A(n11003), .B(n11002), .Z(n11004) );
  NANDN U12872 ( .A(n11005), .B(n11004), .Z(n11006) );
  AND U12873 ( .A(n11007), .B(n11006), .Z(n11008) );
  OR U12874 ( .A(n11009), .B(n11008), .Z(n11010) );
  NAND U12875 ( .A(n11011), .B(n11010), .Z(n11012) );
  NANDN U12876 ( .A(n11013), .B(n11012), .Z(n11014) );
  NAND U12877 ( .A(n11015), .B(n11014), .Z(n11016) );
  NANDN U12878 ( .A(n11017), .B(n11016), .Z(n11018) );
  AND U12879 ( .A(n11019), .B(n11018), .Z(n11020) );
  OR U12880 ( .A(n11021), .B(n11020), .Z(n11022) );
  NAND U12881 ( .A(n11023), .B(n11022), .Z(n11024) );
  NANDN U12882 ( .A(n11025), .B(n11024), .Z(n11026) );
  NAND U12883 ( .A(n11027), .B(n11026), .Z(n11028) );
  NANDN U12884 ( .A(n11029), .B(n11028), .Z(n11030) );
  AND U12885 ( .A(n11031), .B(n11030), .Z(n11032) );
  OR U12886 ( .A(n11033), .B(n11032), .Z(n11034) );
  NAND U12887 ( .A(n11035), .B(n11034), .Z(n11036) );
  NANDN U12888 ( .A(n11037), .B(n11036), .Z(n11038) );
  NAND U12889 ( .A(n11039), .B(n11038), .Z(n11040) );
  NANDN U12890 ( .A(n11041), .B(n11040), .Z(n11042) );
  AND U12891 ( .A(n11043), .B(n11042), .Z(n11044) );
  OR U12892 ( .A(n11045), .B(n11044), .Z(n11046) );
  NAND U12893 ( .A(n11047), .B(n11046), .Z(n11048) );
  NANDN U12894 ( .A(n11049), .B(n11048), .Z(n11050) );
  NAND U12895 ( .A(n11051), .B(n11050), .Z(n11052) );
  NANDN U12896 ( .A(n11053), .B(n11052), .Z(n11054) );
  AND U12897 ( .A(n11055), .B(n11054), .Z(n11056) );
  OR U12898 ( .A(n11057), .B(n11056), .Z(n11058) );
  NAND U12899 ( .A(n11059), .B(n11058), .Z(n11060) );
  NANDN U12900 ( .A(n11061), .B(n11060), .Z(n11062) );
  NAND U12901 ( .A(n11063), .B(n11062), .Z(n11064) );
  NANDN U12902 ( .A(n11065), .B(n11064), .Z(n11066) );
  AND U12903 ( .A(n11067), .B(n11066), .Z(n11068) );
  OR U12904 ( .A(n11069), .B(n11068), .Z(n11070) );
  NAND U12905 ( .A(n11071), .B(n11070), .Z(n11072) );
  NANDN U12906 ( .A(n11073), .B(n11072), .Z(n11074) );
  NAND U12907 ( .A(n11075), .B(n11074), .Z(n11076) );
  NANDN U12908 ( .A(n11077), .B(n11076), .Z(n11078) );
  AND U12909 ( .A(n11079), .B(n11078), .Z(n11080) );
  OR U12910 ( .A(n11081), .B(n11080), .Z(n11082) );
  NAND U12911 ( .A(n11083), .B(n11082), .Z(n11084) );
  NANDN U12912 ( .A(n11085), .B(n11084), .Z(n11086) );
  NAND U12913 ( .A(n11087), .B(n11086), .Z(n11088) );
  NANDN U12914 ( .A(n11089), .B(n11088), .Z(n11090) );
  AND U12915 ( .A(n11091), .B(n11090), .Z(n11092) );
  OR U12916 ( .A(n11093), .B(n11092), .Z(n11094) );
  NAND U12917 ( .A(n11095), .B(n11094), .Z(n11096) );
  NANDN U12918 ( .A(n11097), .B(n11096), .Z(n11098) );
  NAND U12919 ( .A(n11099), .B(n11098), .Z(n11100) );
  NANDN U12920 ( .A(n11101), .B(n11100), .Z(n11102) );
  AND U12921 ( .A(n11103), .B(n11102), .Z(n11104) );
  OR U12922 ( .A(n11105), .B(n11104), .Z(n11106) );
  NAND U12923 ( .A(n11107), .B(n11106), .Z(n11108) );
  NANDN U12924 ( .A(n11109), .B(n11108), .Z(n11110) );
  NAND U12925 ( .A(n11111), .B(n11110), .Z(n11112) );
  NANDN U12926 ( .A(n11113), .B(n11112), .Z(n11114) );
  AND U12927 ( .A(n11115), .B(n11114), .Z(n11116) );
  OR U12928 ( .A(n11117), .B(n11116), .Z(n11118) );
  NAND U12929 ( .A(n11119), .B(n11118), .Z(n11120) );
  NANDN U12930 ( .A(n11121), .B(n11120), .Z(n11122) );
  NAND U12931 ( .A(n11123), .B(n11122), .Z(n11124) );
  NANDN U12932 ( .A(n11125), .B(n11124), .Z(n11126) );
  AND U12933 ( .A(n11127), .B(n11126), .Z(n11128) );
  OR U12934 ( .A(n11129), .B(n11128), .Z(n11130) );
  NAND U12935 ( .A(n11131), .B(n11130), .Z(n11132) );
  NANDN U12936 ( .A(n11133), .B(n11132), .Z(n11134) );
  NAND U12937 ( .A(n11135), .B(n11134), .Z(n11136) );
  NANDN U12938 ( .A(n11137), .B(n11136), .Z(n11138) );
  AND U12939 ( .A(n11139), .B(n11138), .Z(n11140) );
  OR U12940 ( .A(n11141), .B(n11140), .Z(n11142) );
  NAND U12941 ( .A(n11143), .B(n11142), .Z(n11144) );
  NANDN U12942 ( .A(n11145), .B(n11144), .Z(n11146) );
  NAND U12943 ( .A(n11147), .B(n11146), .Z(n11148) );
  NANDN U12944 ( .A(n11149), .B(n11148), .Z(n11150) );
  AND U12945 ( .A(n11151), .B(n11150), .Z(n11152) );
  OR U12946 ( .A(n11153), .B(n11152), .Z(n11154) );
  NAND U12947 ( .A(n11155), .B(n11154), .Z(n11156) );
  NANDN U12948 ( .A(n11157), .B(n11156), .Z(n11158) );
  NAND U12949 ( .A(n11159), .B(n11158), .Z(n11160) );
  NANDN U12950 ( .A(n11161), .B(n11160), .Z(n11162) );
  AND U12951 ( .A(n11163), .B(n11162), .Z(n11164) );
  OR U12952 ( .A(n11165), .B(n11164), .Z(n11166) );
  NAND U12953 ( .A(n11167), .B(n11166), .Z(n11168) );
  NANDN U12954 ( .A(n11169), .B(n11168), .Z(n11170) );
  NAND U12955 ( .A(n11171), .B(n11170), .Z(n11172) );
  NANDN U12956 ( .A(n11173), .B(n11172), .Z(n11174) );
  AND U12957 ( .A(n11175), .B(n11174), .Z(n11176) );
  OR U12958 ( .A(n11177), .B(n11176), .Z(n11178) );
  NAND U12959 ( .A(n11179), .B(n11178), .Z(n11180) );
  NANDN U12960 ( .A(n11181), .B(n11180), .Z(n11182) );
  NAND U12961 ( .A(n11183), .B(n11182), .Z(n11184) );
  NANDN U12962 ( .A(n11185), .B(n11184), .Z(n11186) );
  AND U12963 ( .A(n11187), .B(n11186), .Z(n11188) );
  OR U12964 ( .A(n11189), .B(n11188), .Z(n11190) );
  NAND U12965 ( .A(n11191), .B(n11190), .Z(n11192) );
  NANDN U12966 ( .A(n11193), .B(n11192), .Z(n11194) );
  NAND U12967 ( .A(n11195), .B(n11194), .Z(n11196) );
  NANDN U12968 ( .A(n11197), .B(n11196), .Z(n11198) );
  AND U12969 ( .A(n11199), .B(n11198), .Z(n11200) );
  OR U12970 ( .A(n11201), .B(n11200), .Z(n11202) );
  NAND U12971 ( .A(n11203), .B(n11202), .Z(n11204) );
  NANDN U12972 ( .A(n11205), .B(n11204), .Z(n11206) );
  NAND U12973 ( .A(n11207), .B(n11206), .Z(n11208) );
  NANDN U12974 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U12975 ( .A(n11211), .B(n11210), .Z(n11212) );
  OR U12976 ( .A(n11213), .B(n11212), .Z(n11214) );
  NAND U12977 ( .A(n11215), .B(n11214), .Z(n11216) );
  NANDN U12978 ( .A(n11217), .B(n11216), .Z(n11218) );
  NAND U12979 ( .A(n11219), .B(n11218), .Z(n11220) );
  NANDN U12980 ( .A(n11221), .B(n11220), .Z(n11222) );
  AND U12981 ( .A(n11223), .B(n11222), .Z(n11224) );
  OR U12982 ( .A(n11225), .B(n11224), .Z(n11226) );
  NAND U12983 ( .A(n11227), .B(n11226), .Z(n11228) );
  NANDN U12984 ( .A(n11229), .B(n11228), .Z(n11230) );
  NAND U12985 ( .A(n11231), .B(n11230), .Z(n11232) );
  NANDN U12986 ( .A(n11233), .B(n11232), .Z(n11234) );
  AND U12987 ( .A(n11235), .B(n11234), .Z(n11236) );
  OR U12988 ( .A(n11237), .B(n11236), .Z(n11238) );
  NAND U12989 ( .A(n11239), .B(n11238), .Z(n11240) );
  NANDN U12990 ( .A(n11241), .B(n11240), .Z(n11242) );
  NAND U12991 ( .A(n11243), .B(n11242), .Z(n11244) );
  NANDN U12992 ( .A(n11245), .B(n11244), .Z(n11246) );
  AND U12993 ( .A(n11247), .B(n11246), .Z(n11248) );
  OR U12994 ( .A(n11249), .B(n11248), .Z(n11250) );
  NAND U12995 ( .A(n11251), .B(n11250), .Z(n11252) );
  NANDN U12996 ( .A(n11253), .B(n11252), .Z(n11254) );
  NAND U12997 ( .A(n11255), .B(n11254), .Z(n11256) );
  NANDN U12998 ( .A(n11257), .B(n11256), .Z(n11258) );
  AND U12999 ( .A(n11259), .B(n11258), .Z(n11260) );
  OR U13000 ( .A(n11261), .B(n11260), .Z(n11262) );
  NAND U13001 ( .A(n11263), .B(n11262), .Z(n11264) );
  NANDN U13002 ( .A(n11265), .B(n11264), .Z(n11266) );
  NAND U13003 ( .A(n11267), .B(n11266), .Z(n11268) );
  NANDN U13004 ( .A(n11269), .B(n11268), .Z(n11270) );
  AND U13005 ( .A(n11271), .B(n11270), .Z(n11272) );
  OR U13006 ( .A(n11273), .B(n11272), .Z(n11274) );
  NAND U13007 ( .A(n11275), .B(n11274), .Z(n11276) );
  NANDN U13008 ( .A(n11277), .B(n11276), .Z(n11278) );
  NAND U13009 ( .A(n11279), .B(n11278), .Z(n11280) );
  NANDN U13010 ( .A(n11281), .B(n11280), .Z(n11282) );
  AND U13011 ( .A(n11283), .B(n11282), .Z(n11284) );
  OR U13012 ( .A(n11285), .B(n11284), .Z(n11286) );
  NAND U13013 ( .A(n11287), .B(n11286), .Z(n11288) );
  NANDN U13014 ( .A(n11289), .B(n11288), .Z(n11290) );
  NAND U13015 ( .A(n11291), .B(n11290), .Z(n11292) );
  NANDN U13016 ( .A(n11293), .B(n11292), .Z(n11294) );
  AND U13017 ( .A(n11295), .B(n11294), .Z(n11296) );
  OR U13018 ( .A(n11297), .B(n11296), .Z(n11298) );
  NAND U13019 ( .A(n11299), .B(n11298), .Z(n11300) );
  NANDN U13020 ( .A(n11301), .B(n11300), .Z(n11302) );
  NAND U13021 ( .A(n11303), .B(n11302), .Z(n11304) );
  NANDN U13022 ( .A(n11305), .B(n11304), .Z(n11306) );
  AND U13023 ( .A(n11307), .B(n11306), .Z(n11308) );
  OR U13024 ( .A(n11309), .B(n11308), .Z(n11310) );
  NAND U13025 ( .A(n11311), .B(n11310), .Z(n11312) );
  NANDN U13026 ( .A(n11313), .B(n11312), .Z(n11314) );
  NAND U13027 ( .A(n11315), .B(n11314), .Z(n11316) );
  NANDN U13028 ( .A(n11317), .B(n11316), .Z(n11318) );
  AND U13029 ( .A(n11319), .B(n11318), .Z(n11320) );
  OR U13030 ( .A(n11321), .B(n11320), .Z(n11322) );
  NAND U13031 ( .A(n11323), .B(n11322), .Z(n11324) );
  NANDN U13032 ( .A(n11325), .B(n11324), .Z(n11326) );
  NAND U13033 ( .A(n11327), .B(n11326), .Z(n11328) );
  NANDN U13034 ( .A(n11329), .B(n11328), .Z(n11330) );
  AND U13035 ( .A(n11331), .B(n11330), .Z(n11332) );
  OR U13036 ( .A(n11333), .B(n11332), .Z(n11334) );
  NAND U13037 ( .A(n11335), .B(n11334), .Z(n11336) );
  NANDN U13038 ( .A(n11337), .B(n11336), .Z(n11338) );
  NAND U13039 ( .A(n11339), .B(n11338), .Z(n11340) );
  NANDN U13040 ( .A(n11341), .B(n11340), .Z(n11342) );
  AND U13041 ( .A(n11343), .B(n11342), .Z(n11344) );
  OR U13042 ( .A(n11345), .B(n11344), .Z(n11346) );
  NAND U13043 ( .A(n11347), .B(n11346), .Z(n11348) );
  NANDN U13044 ( .A(n11349), .B(n11348), .Z(n11350) );
  NAND U13045 ( .A(n11351), .B(n11350), .Z(n11352) );
  NANDN U13046 ( .A(n11353), .B(n11352), .Z(n11354) );
  AND U13047 ( .A(n11355), .B(n11354), .Z(n11356) );
  OR U13048 ( .A(n11357), .B(n11356), .Z(n11358) );
  NAND U13049 ( .A(n11359), .B(n11358), .Z(n11360) );
  NANDN U13050 ( .A(n11361), .B(n11360), .Z(n11362) );
  NAND U13051 ( .A(n11363), .B(n11362), .Z(n11364) );
  NANDN U13052 ( .A(n11365), .B(n11364), .Z(n11366) );
  AND U13053 ( .A(n11367), .B(n11366), .Z(n11368) );
  OR U13054 ( .A(n11369), .B(n11368), .Z(n11370) );
  NAND U13055 ( .A(n11371), .B(n11370), .Z(n11372) );
  NANDN U13056 ( .A(n11373), .B(n11372), .Z(n11374) );
  NAND U13057 ( .A(n11375), .B(n11374), .Z(n11376) );
  NANDN U13058 ( .A(n11377), .B(n11376), .Z(n11378) );
  AND U13059 ( .A(n11379), .B(n11378), .Z(n11380) );
  OR U13060 ( .A(n11381), .B(n11380), .Z(n11382) );
  NAND U13061 ( .A(n11383), .B(n11382), .Z(n11384) );
  NANDN U13062 ( .A(n11385), .B(n11384), .Z(n11386) );
  NAND U13063 ( .A(n11387), .B(n11386), .Z(n11388) );
  NANDN U13064 ( .A(n11389), .B(n11388), .Z(n11390) );
  AND U13065 ( .A(n11391), .B(n11390), .Z(n11392) );
  OR U13066 ( .A(n11393), .B(n11392), .Z(n11394) );
  NAND U13067 ( .A(n11395), .B(n11394), .Z(n11396) );
  NANDN U13068 ( .A(n11397), .B(n11396), .Z(n11398) );
  NAND U13069 ( .A(n11399), .B(n11398), .Z(n11400) );
  NANDN U13070 ( .A(n11401), .B(n11400), .Z(n11402) );
  AND U13071 ( .A(n11403), .B(n11402), .Z(n11404) );
  OR U13072 ( .A(n11405), .B(n11404), .Z(n11406) );
  NAND U13073 ( .A(n11407), .B(n11406), .Z(n11408) );
  NANDN U13074 ( .A(n11409), .B(n11408), .Z(n11410) );
  NAND U13075 ( .A(n11411), .B(n11410), .Z(n11412) );
  NANDN U13076 ( .A(n11413), .B(n11412), .Z(n11414) );
  AND U13077 ( .A(n11415), .B(n11414), .Z(n11416) );
  OR U13078 ( .A(n11417), .B(n11416), .Z(n11418) );
  NAND U13079 ( .A(n11419), .B(n11418), .Z(n11420) );
  NANDN U13080 ( .A(n11421), .B(n11420), .Z(n11422) );
  NAND U13081 ( .A(n11423), .B(n11422), .Z(n11424) );
  NANDN U13082 ( .A(n11425), .B(n11424), .Z(n11426) );
  AND U13083 ( .A(n11427), .B(n11426), .Z(n11428) );
  OR U13084 ( .A(n11429), .B(n11428), .Z(n11430) );
  NAND U13085 ( .A(n11431), .B(n11430), .Z(n11432) );
  NANDN U13086 ( .A(n11433), .B(n11432), .Z(n11434) );
  NAND U13087 ( .A(n11435), .B(n11434), .Z(n11436) );
  NANDN U13088 ( .A(n11437), .B(n11436), .Z(n11438) );
  AND U13089 ( .A(n11439), .B(n11438), .Z(n11440) );
  OR U13090 ( .A(n11441), .B(n11440), .Z(n11442) );
  NAND U13091 ( .A(n11443), .B(n11442), .Z(n11444) );
  NANDN U13092 ( .A(n11445), .B(n11444), .Z(n11446) );
  NAND U13093 ( .A(n11447), .B(n11446), .Z(n11448) );
  NANDN U13094 ( .A(n11449), .B(n11448), .Z(n11450) );
  AND U13095 ( .A(n11451), .B(n11450), .Z(n11452) );
  OR U13096 ( .A(n11453), .B(n11452), .Z(n11454) );
  NAND U13097 ( .A(n11455), .B(n11454), .Z(n11456) );
  NANDN U13098 ( .A(n11457), .B(n11456), .Z(n11458) );
  NAND U13099 ( .A(n11459), .B(n11458), .Z(n11460) );
  NANDN U13100 ( .A(n11461), .B(n11460), .Z(n11462) );
  AND U13101 ( .A(n11463), .B(n11462), .Z(n11464) );
  OR U13102 ( .A(n11465), .B(n11464), .Z(n11466) );
  NAND U13103 ( .A(n11467), .B(n11466), .Z(n11468) );
  NANDN U13104 ( .A(n11469), .B(n11468), .Z(n11470) );
  NAND U13105 ( .A(n11471), .B(n11470), .Z(n11472) );
  NANDN U13106 ( .A(n11473), .B(n11472), .Z(n11474) );
  AND U13107 ( .A(n11475), .B(n11474), .Z(n11477) );
  NANDN U13108 ( .A(n11477), .B(n11476), .Z(n11478) );
  NANDN U13109 ( .A(n11479), .B(n11478), .Z(n11480) );
  NAND U13110 ( .A(n11481), .B(n11480), .Z(n11482) );
  NANDN U13111 ( .A(n11483), .B(n11482), .Z(n11484) );
  NAND U13112 ( .A(n11485), .B(n11484), .Z(n11487) );
  ANDN U13113 ( .B(n11487), .A(n11486), .Z(n11489) );
  NANDN U13114 ( .A(n11489), .B(n11488), .Z(n11490) );
  NANDN U13115 ( .A(n11491), .B(n11490), .Z(n11492) );
  NAND U13116 ( .A(n11493), .B(n11492), .Z(n11494) );
  NAND U13117 ( .A(n11495), .B(n11494), .Z(n11496) );
  NANDN U13118 ( .A(n11497), .B(n11496), .Z(n11498) );
  AND U13119 ( .A(n11499), .B(n11498), .Z(n11500) );
  OR U13120 ( .A(n11501), .B(n11500), .Z(n11502) );
  NAND U13121 ( .A(n11503), .B(n11502), .Z(n11504) );
  NANDN U13122 ( .A(n11505), .B(n11504), .Z(n11506) );
  NAND U13123 ( .A(n11507), .B(n11506), .Z(n11508) );
  NANDN U13124 ( .A(n11509), .B(n11508), .Z(n11510) );
  AND U13125 ( .A(n11511), .B(n11510), .Z(n11512) );
  OR U13126 ( .A(n11513), .B(n11512), .Z(n11514) );
  NAND U13127 ( .A(n11515), .B(n11514), .Z(n11516) );
  NANDN U13128 ( .A(n11517), .B(n11516), .Z(n11518) );
  NAND U13129 ( .A(n11519), .B(n11518), .Z(n11520) );
  NANDN U13130 ( .A(n11521), .B(n11520), .Z(n11522) );
  AND U13131 ( .A(n11523), .B(n11522), .Z(n11524) );
  OR U13132 ( .A(n11525), .B(n11524), .Z(n11526) );
  NAND U13133 ( .A(n11527), .B(n11526), .Z(n11528) );
  NANDN U13134 ( .A(n11529), .B(n11528), .Z(n11530) );
  NAND U13135 ( .A(n11531), .B(n11530), .Z(n11532) );
  NANDN U13136 ( .A(n11533), .B(n11532), .Z(n11534) );
  AND U13137 ( .A(n11535), .B(n11534), .Z(n11536) );
  OR U13138 ( .A(n11537), .B(n11536), .Z(n11538) );
  NAND U13139 ( .A(n11539), .B(n11538), .Z(n11540) );
  NANDN U13140 ( .A(n11541), .B(n11540), .Z(n11542) );
  NAND U13141 ( .A(n11543), .B(n11542), .Z(n11544) );
  NANDN U13142 ( .A(n11545), .B(n11544), .Z(n11546) );
  AND U13143 ( .A(n11547), .B(n11546), .Z(n11548) );
  OR U13144 ( .A(n11549), .B(n11548), .Z(n11550) );
  NAND U13145 ( .A(n11551), .B(n11550), .Z(n11552) );
  NANDN U13146 ( .A(n11553), .B(n11552), .Z(n11554) );
  NAND U13147 ( .A(n11555), .B(n11554), .Z(n11556) );
  NANDN U13148 ( .A(n11557), .B(n11556), .Z(n11558) );
  AND U13149 ( .A(n11559), .B(n11558), .Z(n11560) );
  OR U13150 ( .A(n11561), .B(n11560), .Z(n11562) );
  NAND U13151 ( .A(n11563), .B(n11562), .Z(n11564) );
  NANDN U13152 ( .A(n11565), .B(n11564), .Z(n11566) );
  NAND U13153 ( .A(n11567), .B(n11566), .Z(n11568) );
  NANDN U13154 ( .A(n11569), .B(n11568), .Z(n11570) );
  AND U13155 ( .A(n11571), .B(n11570), .Z(n11572) );
  OR U13156 ( .A(n11573), .B(n11572), .Z(n11574) );
  NAND U13157 ( .A(n11575), .B(n11574), .Z(n11576) );
  NANDN U13158 ( .A(n11577), .B(n11576), .Z(n11578) );
  NAND U13159 ( .A(n11579), .B(n11578), .Z(n11580) );
  NANDN U13160 ( .A(n11581), .B(n11580), .Z(n11582) );
  AND U13161 ( .A(n11583), .B(n11582), .Z(n11584) );
  OR U13162 ( .A(n11585), .B(n11584), .Z(n11586) );
  NAND U13163 ( .A(n11587), .B(n11586), .Z(n11588) );
  NANDN U13164 ( .A(n11589), .B(n11588), .Z(n11590) );
  NAND U13165 ( .A(n11591), .B(n11590), .Z(n11592) );
  NANDN U13166 ( .A(n11593), .B(n11592), .Z(n11594) );
  AND U13167 ( .A(n11595), .B(n11594), .Z(n11596) );
  OR U13168 ( .A(n11597), .B(n11596), .Z(n11598) );
  NAND U13169 ( .A(n11599), .B(n11598), .Z(n11600) );
  NANDN U13170 ( .A(n11601), .B(n11600), .Z(n11602) );
  NAND U13171 ( .A(n11603), .B(n11602), .Z(n11604) );
  NANDN U13172 ( .A(n11605), .B(n11604), .Z(n11606) );
  AND U13173 ( .A(n11607), .B(n11606), .Z(n11608) );
  OR U13174 ( .A(n11609), .B(n11608), .Z(n11610) );
  NAND U13175 ( .A(n11611), .B(n11610), .Z(n11612) );
  NAND U13176 ( .A(n11613), .B(n11612), .Z(n11614) );
  NANDN U13177 ( .A(n11615), .B(n11614), .Z(n11616) );
  NAND U13178 ( .A(n11617), .B(n11616), .Z(n11618) );
  AND U13179 ( .A(n11619), .B(n11618), .Z(n11621) );
  NANDN U13180 ( .A(n11621), .B(n11620), .Z(n11622) );
  NAND U13181 ( .A(n11623), .B(n11622), .Z(n11624) );
  NAND U13182 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U13183 ( .A(n11627), .B(n11626), .Z(n11628) );
  NAND U13184 ( .A(n11629), .B(n11628), .Z(n11630) );
  AND U13185 ( .A(n11631), .B(n11630), .Z(n11633) );
  NANDN U13186 ( .A(n11633), .B(n11632), .Z(n11634) );
  NANDN U13187 ( .A(n11635), .B(n11634), .Z(n11636) );
  NAND U13188 ( .A(n11637), .B(n11636), .Z(n11638) );
  NANDN U13189 ( .A(n11639), .B(n11638), .Z(n11640) );
  NAND U13190 ( .A(n11641), .B(n11640), .Z(n11642) );
  AND U13191 ( .A(n11643), .B(n11642), .Z(n11645) );
  NANDN U13192 ( .A(n11645), .B(n11644), .Z(n11646) );
  NANDN U13193 ( .A(n11647), .B(n11646), .Z(n11648) );
  NAND U13194 ( .A(n11649), .B(n11648), .Z(n11650) );
  NANDN U13195 ( .A(n11651), .B(n11650), .Z(n11652) );
  NAND U13196 ( .A(n11653), .B(n11652), .Z(n11655) );
  ANDN U13197 ( .B(n11655), .A(n11654), .Z(n11657) );
  NANDN U13198 ( .A(n11657), .B(n11656), .Z(n11658) );
  NANDN U13199 ( .A(n11659), .B(n11658), .Z(n11660) );
  NAND U13200 ( .A(n11661), .B(n11660), .Z(n11662) );
  NANDN U13201 ( .A(n11663), .B(n11662), .Z(n11664) );
  NAND U13202 ( .A(n11665), .B(n11664), .Z(n11667) );
  ANDN U13203 ( .B(n11667), .A(n11666), .Z(n11669) );
  NANDN U13204 ( .A(n11669), .B(n11668), .Z(n11670) );
  NANDN U13205 ( .A(n11671), .B(n11670), .Z(n11672) );
  NAND U13206 ( .A(n11673), .B(n11672), .Z(n11674) );
  NANDN U13207 ( .A(n11675), .B(n11674), .Z(n11676) );
  NAND U13208 ( .A(n11677), .B(n11676), .Z(n11679) );
  ANDN U13209 ( .B(n11679), .A(n11678), .Z(n11681) );
  NANDN U13210 ( .A(n11681), .B(n11680), .Z(n11682) );
  NANDN U13211 ( .A(n11683), .B(n11682), .Z(n11684) );
  NAND U13212 ( .A(n11685), .B(n11684), .Z(n11686) );
  NANDN U13213 ( .A(n11687), .B(n11686), .Z(n11688) );
  NAND U13214 ( .A(n11689), .B(n11688), .Z(n11691) );
  ANDN U13215 ( .B(n11691), .A(n11690), .Z(n11693) );
  NANDN U13216 ( .A(n11693), .B(n11692), .Z(n11694) );
  NANDN U13217 ( .A(n11695), .B(n11694), .Z(n11696) );
  NAND U13218 ( .A(n11697), .B(n11696), .Z(n11698) );
  NAND U13219 ( .A(n11699), .B(n11698), .Z(n11700) );
  NAND U13220 ( .A(n11701), .B(n11700), .Z(n11702) );
  AND U13221 ( .A(n11703), .B(n11702), .Z(n11705) );
  NANDN U13222 ( .A(n11705), .B(n11704), .Z(n11706) );
  NAND U13223 ( .A(n11707), .B(n11706), .Z(n11708) );
  NAND U13224 ( .A(n11709), .B(n11708), .Z(n11710) );
  NANDN U13225 ( .A(n11711), .B(n11710), .Z(n11712) );
  NAND U13226 ( .A(n11713), .B(n11712), .Z(n11714) );
  AND U13227 ( .A(n11715), .B(n11714), .Z(n11717) );
  NANDN U13228 ( .A(n11717), .B(n11716), .Z(n11718) );
  NANDN U13229 ( .A(n11719), .B(n11718), .Z(n11720) );
  NAND U13230 ( .A(n11721), .B(n11720), .Z(n11722) );
  NANDN U13231 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U13232 ( .A(n11725), .B(n11724), .Z(n11727) );
  ANDN U13233 ( .B(n11727), .A(n11726), .Z(n11729) );
  NANDN U13234 ( .A(n11729), .B(n11728), .Z(n11730) );
  NANDN U13235 ( .A(n11731), .B(n11730), .Z(n11732) );
  NAND U13236 ( .A(n11733), .B(n11732), .Z(n11734) );
  NANDN U13237 ( .A(n11735), .B(n11734), .Z(n11736) );
  NAND U13238 ( .A(n11737), .B(n11736), .Z(n11739) );
  ANDN U13239 ( .B(n11739), .A(n11738), .Z(n11741) );
  NANDN U13240 ( .A(n11741), .B(n11740), .Z(n11742) );
  NANDN U13241 ( .A(n11743), .B(n11742), .Z(n11744) );
  NAND U13242 ( .A(n11745), .B(n11744), .Z(n11746) );
  NANDN U13243 ( .A(n11747), .B(n11746), .Z(n11748) );
  NAND U13244 ( .A(n11749), .B(n11748), .Z(n11751) );
  ANDN U13245 ( .B(n11751), .A(n11750), .Z(n11753) );
  NANDN U13246 ( .A(n11753), .B(n11752), .Z(n11754) );
  NANDN U13247 ( .A(n11755), .B(n11754), .Z(n11756) );
  NAND U13248 ( .A(n11757), .B(n11756), .Z(n11758) );
  NAND U13249 ( .A(n11759), .B(n11758), .Z(n11760) );
  NANDN U13250 ( .A(n11761), .B(n11760), .Z(n11762) );
  AND U13251 ( .A(n11763), .B(n11762), .Z(n11764) );
  OR U13252 ( .A(n11765), .B(n11764), .Z(n11766) );
  NAND U13253 ( .A(n11767), .B(n11766), .Z(n11768) );
  NANDN U13254 ( .A(n11769), .B(n11768), .Z(n11770) );
  NAND U13255 ( .A(n11771), .B(n11770), .Z(n11772) );
  NANDN U13256 ( .A(n11773), .B(n11772), .Z(n11774) );
  AND U13257 ( .A(n11775), .B(n11774), .Z(n11776) );
  OR U13258 ( .A(n11777), .B(n11776), .Z(n11778) );
  NAND U13259 ( .A(n11779), .B(n11778), .Z(n11780) );
  NANDN U13260 ( .A(n11781), .B(n11780), .Z(n11782) );
  NAND U13261 ( .A(n11783), .B(n11782), .Z(n11784) );
  NANDN U13262 ( .A(n11785), .B(n11784), .Z(n11786) );
  AND U13263 ( .A(n11787), .B(n11786), .Z(n11788) );
  OR U13264 ( .A(n11789), .B(n11788), .Z(n11790) );
  NAND U13265 ( .A(n11791), .B(n11790), .Z(n11792) );
  NANDN U13266 ( .A(n11793), .B(n11792), .Z(n11794) );
  NAND U13267 ( .A(n11795), .B(n11794), .Z(n11796) );
  NANDN U13268 ( .A(n11797), .B(n11796), .Z(n11798) );
  AND U13269 ( .A(n11799), .B(n11798), .Z(n11800) );
  OR U13270 ( .A(n11801), .B(n11800), .Z(n11802) );
  NAND U13271 ( .A(n11803), .B(n11802), .Z(n11804) );
  NANDN U13272 ( .A(n11805), .B(n11804), .Z(n11806) );
  NAND U13273 ( .A(n11807), .B(n11806), .Z(n11808) );
  NANDN U13274 ( .A(n11809), .B(n11808), .Z(n11810) );
  AND U13275 ( .A(n11811), .B(n11810), .Z(n11812) );
  OR U13276 ( .A(n11813), .B(n11812), .Z(n11814) );
  NAND U13277 ( .A(n11815), .B(n11814), .Z(n11816) );
  NANDN U13278 ( .A(n11817), .B(n11816), .Z(n11818) );
  NAND U13279 ( .A(n11819), .B(n11818), .Z(n11820) );
  NANDN U13280 ( .A(n11821), .B(n11820), .Z(n11822) );
  AND U13281 ( .A(n11823), .B(n11822), .Z(n11824) );
  OR U13282 ( .A(n11825), .B(n11824), .Z(n11826) );
  NAND U13283 ( .A(n11827), .B(n11826), .Z(n11828) );
  NAND U13284 ( .A(n11829), .B(n11828), .Z(n11830) );
  NANDN U13285 ( .A(n11831), .B(n11830), .Z(n11832) );
  NAND U13286 ( .A(n11833), .B(n11832), .Z(n11835) );
  ANDN U13287 ( .B(n11835), .A(n11834), .Z(n11837) );
  NANDN U13288 ( .A(n11837), .B(n11836), .Z(n11838) );
  NAND U13289 ( .A(n11839), .B(n11838), .Z(n11840) );
  NANDN U13290 ( .A(n11841), .B(n11840), .Z(n11843) );
  NAND U13291 ( .A(n11843), .B(n11842), .Z(n11844) );
  NANDN U13292 ( .A(n11845), .B(n11844), .Z(n11846) );
  AND U13293 ( .A(n11847), .B(n11846), .Z(n11848) );
  OR U13294 ( .A(n11849), .B(n11848), .Z(n11850) );
  NAND U13295 ( .A(n11851), .B(n11850), .Z(n11852) );
  NANDN U13296 ( .A(n11853), .B(n11852), .Z(n11854) );
  NAND U13297 ( .A(n11855), .B(n11854), .Z(n11856) );
  NANDN U13298 ( .A(n11857), .B(n11856), .Z(n11858) );
  AND U13299 ( .A(n11859), .B(n11858), .Z(n11860) );
  OR U13300 ( .A(n11861), .B(n11860), .Z(n11862) );
  NAND U13301 ( .A(n11863), .B(n11862), .Z(n11864) );
  NANDN U13302 ( .A(n11865), .B(n11864), .Z(n11866) );
  NAND U13303 ( .A(n11867), .B(n11866), .Z(n11868) );
  NANDN U13304 ( .A(n11869), .B(n11868), .Z(n11870) );
  AND U13305 ( .A(n11871), .B(n11870), .Z(n11873) );
  NANDN U13306 ( .A(n11873), .B(n11872), .Z(n11874) );
  NAND U13307 ( .A(n11875), .B(n11874), .Z(n11876) );
  NANDN U13308 ( .A(n11877), .B(n11876), .Z(n11879) );
  NANDN U13309 ( .A(n11879), .B(n11878), .Z(n11880) );
  NAND U13310 ( .A(n11881), .B(n11880), .Z(n11882) );
  NAND U13311 ( .A(n11883), .B(n11882), .Z(n11885) );
  NAND U13312 ( .A(n11885), .B(n11884), .Z(n11886) );
  NANDN U13313 ( .A(n11887), .B(n11886), .Z(n11888) );
  AND U13314 ( .A(n11889), .B(n11888), .Z(n11890) );
  OR U13315 ( .A(n11891), .B(n11890), .Z(n11892) );
  NAND U13316 ( .A(n11893), .B(n11892), .Z(n11894) );
  NANDN U13317 ( .A(n11895), .B(n11894), .Z(n11896) );
  NAND U13318 ( .A(n11897), .B(n11896), .Z(n11898) );
  NANDN U13319 ( .A(n11899), .B(n11898), .Z(n11900) );
  AND U13320 ( .A(n11901), .B(n11900), .Z(n11903) );
  NANDN U13321 ( .A(n11903), .B(n11902), .Z(n11904) );
  NAND U13322 ( .A(n11905), .B(n11904), .Z(n11906) );
  NAND U13323 ( .A(n11907), .B(n11906), .Z(n11909) );
  NAND U13324 ( .A(n11909), .B(n11908), .Z(n11910) );
  NANDN U13325 ( .A(n11911), .B(n11910), .Z(n11912) );
  AND U13326 ( .A(n11913), .B(n11912), .Z(n11914) );
  OR U13327 ( .A(n11915), .B(n11914), .Z(n11916) );
  NAND U13328 ( .A(n11917), .B(n11916), .Z(n11918) );
  NANDN U13329 ( .A(n11919), .B(n11918), .Z(n11920) );
  NAND U13330 ( .A(n11921), .B(n11920), .Z(n11922) );
  NANDN U13331 ( .A(n11923), .B(n11922), .Z(n11924) );
  AND U13332 ( .A(n11925), .B(n11924), .Z(n11926) );
  OR U13333 ( .A(n11927), .B(n11926), .Z(n11928) );
  NAND U13334 ( .A(n11929), .B(n11928), .Z(n11930) );
  NANDN U13335 ( .A(n11931), .B(n11930), .Z(n11932) );
  NAND U13336 ( .A(n11933), .B(n11932), .Z(n11934) );
  NANDN U13337 ( .A(n11935), .B(n11934), .Z(n11936) );
  AND U13338 ( .A(n11937), .B(n11936), .Z(n11938) );
  OR U13339 ( .A(n11939), .B(n11938), .Z(n11940) );
  NAND U13340 ( .A(n11941), .B(n11940), .Z(n11942) );
  NANDN U13341 ( .A(n11943), .B(n11942), .Z(n11944) );
  NAND U13342 ( .A(n11945), .B(n11944), .Z(n11946) );
  NAND U13343 ( .A(n11947), .B(n11946), .Z(n11948) );
  NAND U13344 ( .A(n11949), .B(n11948), .Z(n11950) );
  NAND U13345 ( .A(n11951), .B(n11950), .Z(n11952) );
  NANDN U13346 ( .A(n11953), .B(n11952), .Z(n11954) );
  AND U13347 ( .A(n11955), .B(n11954), .Z(n11956) );
  OR U13348 ( .A(n11957), .B(n11956), .Z(n11958) );
  NANDN U13349 ( .A(n11959), .B(n11958), .Z(n11960) );
  NAND U13350 ( .A(n11961), .B(n11960), .Z(n11962) );
  NANDN U13351 ( .A(n11963), .B(n11962), .Z(n11964) );
  NAND U13352 ( .A(n11965), .B(n11964), .Z(n11966) );
  AND U13353 ( .A(n11967), .B(n11966), .Z(n11969) );
  NANDN U13354 ( .A(n11969), .B(n11968), .Z(n11970) );
  NANDN U13355 ( .A(n11971), .B(n11970), .Z(n11972) );
  NAND U13356 ( .A(n11973), .B(n11972), .Z(n11974) );
  NAND U13357 ( .A(n11975), .B(n11974), .Z(n11976) );
  NAND U13358 ( .A(n11977), .B(n11976), .Z(n11979) );
  ANDN U13359 ( .B(n11979), .A(n11978), .Z(n11981) );
  NANDN U13360 ( .A(n11981), .B(n11980), .Z(n11982) );
  NANDN U13361 ( .A(n11983), .B(n11982), .Z(n11984) );
  NAND U13362 ( .A(n11985), .B(n11984), .Z(n11986) );
  NAND U13363 ( .A(n11987), .B(n11986), .Z(n11988) );
  NAND U13364 ( .A(n11989), .B(n11988), .Z(n11991) );
  ANDN U13365 ( .B(n11991), .A(n11990), .Z(n11993) );
  NANDN U13366 ( .A(n11993), .B(n11992), .Z(n11994) );
  NANDN U13367 ( .A(n11995), .B(n11994), .Z(n11996) );
  NANDN U13368 ( .A(n11997), .B(n11996), .Z(n11998) );
  NAND U13369 ( .A(n11999), .B(n11998), .Z(n12000) );
  NANDN U13370 ( .A(n12001), .B(n12000), .Z(n12003) );
  ANDN U13371 ( .B(n12003), .A(n12002), .Z(n12005) );
  NANDN U13372 ( .A(n12005), .B(n12004), .Z(n12006) );
  NANDN U13373 ( .A(n12007), .B(n12006), .Z(n12008) );
  NAND U13374 ( .A(n12009), .B(n12008), .Z(n12010) );
  NAND U13375 ( .A(n12011), .B(n12010), .Z(n12012) );
  NAND U13376 ( .A(n12013), .B(n12012), .Z(n12014) );
  AND U13377 ( .A(n12015), .B(n12014), .Z(n12016) );
  OR U13378 ( .A(n12017), .B(n12016), .Z(n12018) );
  NAND U13379 ( .A(n12019), .B(n12018), .Z(n12020) );
  NANDN U13380 ( .A(n12021), .B(n12020), .Z(n12022) );
  NANDN U13381 ( .A(n12023), .B(n12022), .Z(n12024) );
  NAND U13382 ( .A(n12025), .B(n12024), .Z(n12027) );
  ANDN U13383 ( .B(n12027), .A(n12026), .Z(n12029) );
  NANDN U13384 ( .A(n12029), .B(n12028), .Z(n12030) );
  NANDN U13385 ( .A(n12031), .B(n12030), .Z(n12032) );
  NAND U13386 ( .A(n12033), .B(n12032), .Z(n12034) );
  NANDN U13387 ( .A(n12035), .B(n12034), .Z(n12036) );
  AND U13388 ( .A(n12037), .B(n12036), .Z(n12039) );
  NANDN U13389 ( .A(n12039), .B(n12038), .Z(n12040) );
  NAND U13390 ( .A(n12041), .B(n12040), .Z(n12043) );
  ANDN U13391 ( .B(n12043), .A(n12042), .Z(n12045) );
  NANDN U13392 ( .A(n12045), .B(n12044), .Z(n12046) );
  NANDN U13393 ( .A(n12047), .B(n12046), .Z(n12048) );
  NAND U13394 ( .A(n12049), .B(n12048), .Z(n12050) );
  NANDN U13395 ( .A(n12051), .B(n12050), .Z(n12052) );
  NAND U13396 ( .A(n12053), .B(n12052), .Z(n12054) );
  AND U13397 ( .A(n12055), .B(n12054), .Z(n12057) );
  NANDN U13398 ( .A(n12057), .B(n12056), .Z(n12058) );
  NANDN U13399 ( .A(n12059), .B(n12058), .Z(n12060) );
  NAND U13400 ( .A(n12061), .B(n12060), .Z(n12062) );
  NANDN U13401 ( .A(n12063), .B(n12062), .Z(n12064) );
  NAND U13402 ( .A(n12065), .B(n12064), .Z(n12066) );
  AND U13403 ( .A(n12067), .B(n12066), .Z(n12069) );
  NANDN U13404 ( .A(n12069), .B(n12068), .Z(n12070) );
  NAND U13405 ( .A(n12071), .B(n12070), .Z(n12072) );
  NANDN U13406 ( .A(n12073), .B(n12072), .Z(n12075) );
  NAND U13407 ( .A(n12075), .B(n12074), .Z(n12076) );
  NANDN U13408 ( .A(n12077), .B(n12076), .Z(n12078) );
  AND U13409 ( .A(n12079), .B(n12078), .Z(n12080) );
  OR U13410 ( .A(n12081), .B(n12080), .Z(n12082) );
  NAND U13411 ( .A(n12083), .B(n12082), .Z(n12084) );
  NANDN U13412 ( .A(n12085), .B(n12084), .Z(n12086) );
  NAND U13413 ( .A(n12087), .B(n12086), .Z(n12088) );
  NAND U13414 ( .A(n12089), .B(n12088), .Z(n12090) );
  AND U13415 ( .A(n12091), .B(n12090), .Z(n12092) );
  OR U13416 ( .A(n12093), .B(n12092), .Z(n12094) );
  NAND U13417 ( .A(n12095), .B(n12094), .Z(n12096) );
  NAND U13418 ( .A(n12097), .B(n12096), .Z(n12098) );
  NANDN U13419 ( .A(n12099), .B(n12098), .Z(n12100) );
  NAND U13420 ( .A(n12101), .B(n12100), .Z(n12102) );
  AND U13421 ( .A(n12103), .B(n12102), .Z(n12104) );
  OR U13422 ( .A(n12105), .B(n12104), .Z(n12106) );
  NANDN U13423 ( .A(n12107), .B(n12106), .Z(n12108) );
  NANDN U13424 ( .A(n12109), .B(n12108), .Z(n12110) );
  NAND U13425 ( .A(n12111), .B(n12110), .Z(n12112) );
  NANDN U13426 ( .A(n12113), .B(n12112), .Z(n12114) );
  AND U13427 ( .A(n12115), .B(n12114), .Z(n12116) );
  OR U13428 ( .A(n12117), .B(n12116), .Z(n12118) );
  NAND U13429 ( .A(n12119), .B(n12118), .Z(n12120) );
  NANDN U13430 ( .A(n12121), .B(n12120), .Z(n12122) );
  NAND U13431 ( .A(n12123), .B(n12122), .Z(n12124) );
  NANDN U13432 ( .A(n12125), .B(n12124), .Z(n12126) );
  AND U13433 ( .A(n12127), .B(n12126), .Z(n12128) );
  OR U13434 ( .A(n12129), .B(n12128), .Z(n12130) );
  NAND U13435 ( .A(n12131), .B(n12130), .Z(n12132) );
  NANDN U13436 ( .A(n12133), .B(n12132), .Z(n12134) );
  NANDN U13437 ( .A(n12135), .B(n12134), .Z(n12136) );
  NANDN U13438 ( .A(n12137), .B(n12136), .Z(n12138) );
  AND U13439 ( .A(n12139), .B(n12138), .Z(n12140) );
  OR U13440 ( .A(n12141), .B(n12140), .Z(n12142) );
  NAND U13441 ( .A(n12143), .B(n12142), .Z(n12144) );
  NANDN U13442 ( .A(n12145), .B(n12144), .Z(n12147) );
  NAND U13443 ( .A(n12147), .B(n12146), .Z(n12148) );
  NANDN U13444 ( .A(n12149), .B(n12148), .Z(n12150) );
  AND U13445 ( .A(n12151), .B(n12150), .Z(n12152) );
  OR U13446 ( .A(n12153), .B(n12152), .Z(n12154) );
  NAND U13447 ( .A(n12155), .B(n12154), .Z(n12156) );
  NANDN U13448 ( .A(n12157), .B(n12156), .Z(n12158) );
  NAND U13449 ( .A(n12159), .B(n12158), .Z(n12160) );
  NAND U13450 ( .A(n12161), .B(n12160), .Z(n12162) );
  NANDN U13451 ( .A(n12163), .B(n12162), .Z(n12164) );
  NAND U13452 ( .A(n12165), .B(n12164), .Z(n12166) );
  NANDN U13453 ( .A(n12167), .B(n12166), .Z(n12168) );
  AND U13454 ( .A(n12169), .B(n12168), .Z(n12171) );
  NANDN U13455 ( .A(n12171), .B(n12170), .Z(n12172) );
  NAND U13456 ( .A(n12173), .B(n12172), .Z(n12174) );
  NAND U13457 ( .A(n12175), .B(n12174), .Z(n12176) );
  NAND U13458 ( .A(n12177), .B(n12176), .Z(n12178) );
  NAND U13459 ( .A(n12179), .B(n12178), .Z(n12180) );
  NAND U13460 ( .A(n12181), .B(n12180), .Z(n12182) );
  NAND U13461 ( .A(n12183), .B(n12182), .Z(n12184) );
  NAND U13462 ( .A(n12185), .B(n12184), .Z(n12186) );
  AND U13463 ( .A(n12187), .B(n12186), .Z(n12189) );
  NANDN U13464 ( .A(n12189), .B(n12188), .Z(n12190) );
  NAND U13465 ( .A(n12191), .B(n12190), .Z(n12192) );
  NAND U13466 ( .A(n12193), .B(n12192), .Z(n12194) );
  NANDN U13467 ( .A(n12195), .B(n12194), .Z(n12196) );
  NAND U13468 ( .A(n12197), .B(n12196), .Z(n12198) );
  AND U13469 ( .A(n12199), .B(n12198), .Z(n12201) );
  NANDN U13470 ( .A(n12201), .B(n12200), .Z(n12202) );
  NAND U13471 ( .A(n12203), .B(n12202), .Z(n12204) );
  NAND U13472 ( .A(n12205), .B(n12204), .Z(n12206) );
  NAND U13473 ( .A(n12207), .B(n12206), .Z(n12208) );
  NAND U13474 ( .A(n12209), .B(n12208), .Z(n12210) );
  NANDN U13475 ( .A(n12211), .B(n12210), .Z(n12215) );
  NAND U13476 ( .A(n12213), .B(n12212), .Z(n12214) );
  AND U13477 ( .A(n12215), .B(n12214), .Z(n12217) );
  NAND U13478 ( .A(n12217), .B(n12216), .Z(n12218) );
  NANDN U13479 ( .A(n12219), .B(n12218), .Z(n12220) );
  AND U13480 ( .A(n12221), .B(n12220), .Z(n12223) );
  OR U13481 ( .A(n12223), .B(n12222), .Z(n12224) );
  NAND U13482 ( .A(n12225), .B(n12224), .Z(n12227) );
  ANDN U13483 ( .B(n12227), .A(n12226), .Z(n12229) );
  NANDN U13484 ( .A(n12229), .B(n12228), .Z(n12230) );
  AND U13485 ( .A(n12231), .B(n12230), .Z(n12233) );
  NANDN U13486 ( .A(n12233), .B(n12232), .Z(n12234) );
  NAND U13487 ( .A(n12235), .B(n12234), .Z(n12236) );
  NAND U13488 ( .A(n12237), .B(n12236), .Z(n12239) );
  NAND U13489 ( .A(n12239), .B(n12238), .Z(n12240) );
  NAND U13490 ( .A(n12241), .B(n12240), .Z(n12243) );
  ANDN U13491 ( .B(n12243), .A(n12242), .Z(n12245) );
  NANDN U13492 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND U13493 ( .A(n12247), .B(n12246), .Z(n12248) );
  NAND U13494 ( .A(n12249), .B(n12248), .Z(n12250) );
  NAND U13495 ( .A(n12251), .B(n12250), .Z(n12253) );
  ANDN U13496 ( .B(n12253), .A(n12252), .Z(n12255) );
  NANDN U13497 ( .A(n12255), .B(n12254), .Z(n12256) );
  NAND U13498 ( .A(n12257), .B(n12256), .Z(n12258) );
  NANDN U13499 ( .A(n12259), .B(n12258), .Z(n12260) );
  NAND U13500 ( .A(n12261), .B(n12260), .Z(n12262) );
  AND U13501 ( .A(n12263), .B(n12262), .Z(n12265) );
  NANDN U13502 ( .A(n12265), .B(n12264), .Z(n12266) );
  NANDN U13503 ( .A(n12267), .B(n12266), .Z(n12268) );
  NAND U13504 ( .A(n12269), .B(n12268), .Z(n12270) );
  NANDN U13505 ( .A(n12271), .B(n12270), .Z(n12272) );
  AND U13506 ( .A(n12273), .B(n12272), .Z(n12274) );
  OR U13507 ( .A(n12275), .B(n12274), .Z(n12276) );
  NAND U13508 ( .A(n12277), .B(n12276), .Z(n12278) );
  NANDN U13509 ( .A(n12279), .B(n12278), .Z(n12280) );
  NAND U13510 ( .A(n12281), .B(n12280), .Z(n12282) );
  NAND U13511 ( .A(n12283), .B(n12282), .Z(n12285) );
  ANDN U13512 ( .B(n12285), .A(n12284), .Z(n12287) );
  NANDN U13513 ( .A(n12287), .B(n12286), .Z(n12288) );
  AND U13514 ( .A(n12289), .B(n12288), .Z(n12291) );
  OR U13515 ( .A(n12291), .B(n12290), .Z(n12292) );
  NANDN U13516 ( .A(n12293), .B(n12292), .Z(n12294) );
  AND U13517 ( .A(n12295), .B(n12294), .Z(n12297) );
  NANDN U13518 ( .A(n12297), .B(n12296), .Z(n12298) );
  NANDN U13519 ( .A(n12299), .B(n12298), .Z(n12300) );
  AND U13520 ( .A(n12301), .B(n12300), .Z(n12302) );
  OR U13521 ( .A(n12303), .B(n12302), .Z(n12304) );
  NAND U13522 ( .A(n12305), .B(n12304), .Z(n12306) );
  NANDN U13523 ( .A(n12307), .B(n12306), .Z(n12309) );
  ANDN U13524 ( .B(n12309), .A(n12308), .Z(n12311) );
  NANDN U13525 ( .A(n12311), .B(n12310), .Z(n12312) );
  NANDN U13526 ( .A(n12313), .B(n12312), .Z(n12314) );
  AND U13527 ( .A(n12315), .B(n12314), .Z(n12317) );
  NANDN U13528 ( .A(n12317), .B(n12316), .Z(n12318) );
  NANDN U13529 ( .A(n12319), .B(n12318), .Z(n12320) );
  AND U13530 ( .A(n12321), .B(n12320), .Z(n12323) );
  NANDN U13531 ( .A(n12323), .B(n12322), .Z(n12324) );
  NAND U13532 ( .A(n12325), .B(n12324), .Z(n12326) );
  NAND U13533 ( .A(n12327), .B(n12326), .Z(n12328) );
  NANDN U13534 ( .A(n12329), .B(n12328), .Z(n12330) );
  NAND U13535 ( .A(n12331), .B(n12330), .Z(n12332) );
  AND U13536 ( .A(n12333), .B(n12332), .Z(n12335) );
  NANDN U13537 ( .A(n12335), .B(n12334), .Z(n12336) );
  NAND U13538 ( .A(n12337), .B(n12336), .Z(n12338) );
  NAND U13539 ( .A(n12339), .B(n12338), .Z(n12340) );
  NAND U13540 ( .A(n12341), .B(n12340), .Z(n12342) );
  NANDN U13541 ( .A(n12343), .B(n12342), .Z(n12344) );
  AND U13542 ( .A(n12345), .B(n12344), .Z(n12347) );
  OR U13543 ( .A(n12347), .B(n12346), .Z(n12348) );
  NAND U13544 ( .A(n12349), .B(n12348), .Z(n12350) );
  NANDN U13545 ( .A(n12351), .B(n12350), .Z(n12353) );
  NAND U13546 ( .A(n12353), .B(n12352), .Z(n12354) );
  NAND U13547 ( .A(n12355), .B(n12354), .Z(n12357) );
  ANDN U13548 ( .B(n12357), .A(n12356), .Z(n12359) );
  NANDN U13549 ( .A(n12359), .B(n12358), .Z(n12360) );
  NANDN U13550 ( .A(n12361), .B(n12360), .Z(n12362) );
  NANDN U13551 ( .A(n12363), .B(n12362), .Z(n12364) );
  NAND U13552 ( .A(n12365), .B(n12364), .Z(n12366) );
  NANDN U13553 ( .A(n12367), .B(n12366), .Z(n12368) );
  AND U13554 ( .A(n12369), .B(n12368), .Z(n12371) );
  OR U13555 ( .A(n12371), .B(n12370), .Z(n12372) );
  AND U13556 ( .A(n12373), .B(n12372), .Z(n12375) );
  NANDN U13557 ( .A(n12375), .B(n12374), .Z(n12376) );
  NAND U13558 ( .A(n12377), .B(n12376), .Z(n12378) );
  NANDN U13559 ( .A(n12379), .B(n12378), .Z(n12380) );
  NAND U13560 ( .A(n12381), .B(n12380), .Z(n12382) );
  NANDN U13561 ( .A(n12383), .B(n12382), .Z(n12384) );
  AND U13562 ( .A(n12385), .B(n12384), .Z(n12387) );
  OR U13563 ( .A(n12387), .B(n12386), .Z(n12389) );
  ANDN U13564 ( .B(n12389), .A(n12388), .Z(n12391) );
  NANDN U13565 ( .A(n12391), .B(n12390), .Z(n12392) );
  NANDN U13566 ( .A(n12393), .B(n12392), .Z(n12394) );
  NAND U13567 ( .A(n12395), .B(n12394), .Z(n12397) );
  ANDN U13568 ( .B(n12397), .A(n12396), .Z(n12399) );
  NANDN U13569 ( .A(n12399), .B(n12398), .Z(n12400) );
  NANDN U13570 ( .A(n12401), .B(n12400), .Z(n12402) );
  AND U13571 ( .A(n12403), .B(n12402), .Z(n12405) );
  OR U13572 ( .A(n12405), .B(n12404), .Z(n12406) );
  AND U13573 ( .A(n12407), .B(n12406), .Z(n12409) );
  OR U13574 ( .A(n12409), .B(n12408), .Z(n12410) );
  NAND U13575 ( .A(n12411), .B(n12410), .Z(n12412) );
  NANDN U13576 ( .A(n12413), .B(n12412), .Z(n12415) );
  ANDN U13577 ( .B(n12415), .A(n12414), .Z(n12417) );
  NANDN U13578 ( .A(n12417), .B(n12416), .Z(n12418) );
  NANDN U13579 ( .A(n12419), .B(n12418), .Z(n12420) );
  NAND U13580 ( .A(n12421), .B(n12420), .Z(n12423) );
  NAND U13581 ( .A(n12423), .B(n12422), .Z(n12424) );
  NANDN U13582 ( .A(n12425), .B(n12424), .Z(n12426) );
  AND U13583 ( .A(n12427), .B(n12426), .Z(n12429) );
  NANDN U13584 ( .A(n12429), .B(n12428), .Z(n12431) );
  ANDN U13585 ( .B(n12431), .A(n12430), .Z(n12433) );
  NANDN U13586 ( .A(n12433), .B(n12432), .Z(n12435) );
  ANDN U13587 ( .B(n12435), .A(n12434), .Z(n12437) );
  OR U13588 ( .A(n12437), .B(n12436), .Z(n12439) );
  NANDN U13589 ( .A(n12439), .B(n12438), .Z(n12440) );
  NANDN U13590 ( .A(n12441), .B(n12440), .Z(n12442) );
  NAND U13591 ( .A(n12443), .B(n12442), .Z(n12444) );
  NAND U13592 ( .A(n12445), .B(n12444), .Z(n12446) );
  NANDN U13593 ( .A(n12447), .B(n12446), .Z(n12449) );
  ANDN U13594 ( .B(n12449), .A(n12448), .Z(n12451) );
  NANDN U13595 ( .A(n12451), .B(n12450), .Z(n12453) );
  ANDN U13596 ( .B(n12453), .A(n12452), .Z(n12455) );
  OR U13597 ( .A(n12455), .B(n12454), .Z(n12456) );
  NAND U13598 ( .A(n12457), .B(n12456), .Z(n12458) );
  NANDN U13599 ( .A(n12459), .B(n12458), .Z(n12460) );
  AND U13600 ( .A(n12461), .B(n12460), .Z(n12463) );
  NANDN U13601 ( .A(n12463), .B(n12462), .Z(n12464) );
  NANDN U13602 ( .A(n12465), .B(n12464), .Z(n12466) );
  NAND U13603 ( .A(n12467), .B(n12466), .Z(n12469) );
  NAND U13604 ( .A(n12469), .B(n12468), .Z(n12470) );
  NANDN U13605 ( .A(n12471), .B(n12470), .Z(n12472) );
  AND U13606 ( .A(n12473), .B(n12472), .Z(n12475) );
  NANDN U13607 ( .A(n12475), .B(n12474), .Z(n12476) );
  NANDN U13608 ( .A(n12477), .B(n12476), .Z(n12478) );
  NAND U13609 ( .A(n12479), .B(n12478), .Z(n12481) );
  NAND U13610 ( .A(n12481), .B(n12480), .Z(n12482) );
  NANDN U13611 ( .A(n12483), .B(n12482), .Z(n12484) );
  AND U13612 ( .A(n12485), .B(n12484), .Z(n12487) );
  NANDN U13613 ( .A(n12487), .B(n12486), .Z(n12488) );
  NANDN U13614 ( .A(n12489), .B(n12488), .Z(n12490) );
  NAND U13615 ( .A(n12491), .B(n12490), .Z(n12492) );
  NAND U13616 ( .A(n12493), .B(n12492), .Z(n12494) );
  NANDN U13617 ( .A(n12495), .B(n12494), .Z(n12496) );
  NAND U13618 ( .A(n12497), .B(n12496), .Z(n12498) );
  NANDN U13619 ( .A(n12499), .B(n12498), .Z(n12500) );
  NAND U13620 ( .A(n12501), .B(n12500), .Z(n12502) );
  NANDN U13621 ( .A(n12503), .B(n12502), .Z(n12505) );
  ANDN U13622 ( .B(n12505), .A(n12504), .Z(n12507) );
  NANDN U13623 ( .A(n12507), .B(n12506), .Z(n12508) );
  NAND U13624 ( .A(n12509), .B(n12508), .Z(n12510) );
  NAND U13625 ( .A(n12511), .B(n12510), .Z(n12512) );
  NANDN U13626 ( .A(n12513), .B(n12512), .Z(n12514) );
  NAND U13627 ( .A(n12515), .B(n12514), .Z(n12517) );
  ANDN U13628 ( .B(n12517), .A(n12516), .Z(n12519) );
  NANDN U13629 ( .A(n12519), .B(n12518), .Z(n12520) );
  AND U13630 ( .A(n12521), .B(n12520), .Z(n12523) );
  NANDN U13631 ( .A(n12523), .B(n12522), .Z(n12524) );
  NANDN U13632 ( .A(n12525), .B(n12524), .Z(n12526) );
  NAND U13633 ( .A(n12527), .B(n12526), .Z(n12529) );
  ANDN U13634 ( .B(n12529), .A(n12528), .Z(n12531) );
  NANDN U13635 ( .A(n12531), .B(n12530), .Z(n12532) );
  NAND U13636 ( .A(n12533), .B(n12532), .Z(n12534) );
  NAND U13637 ( .A(n12535), .B(n12534), .Z(n12536) );
  NANDN U13638 ( .A(n12537), .B(n12536), .Z(n12538) );
  NANDN U13639 ( .A(n12539), .B(n12538), .Z(n12540) );
  AND U13640 ( .A(n12541), .B(n12540), .Z(n12543) );
  NANDN U13641 ( .A(n12543), .B(n12542), .Z(n12544) );
  AND U13642 ( .A(n12545), .B(n12544), .Z(n12546) );
  OR U13643 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND U13644 ( .A(n12549), .B(n12548), .Z(n12550) );
  NANDN U13645 ( .A(n12551), .B(n12550), .Z(n12552) );
  NAND U13646 ( .A(n12553), .B(n12552), .Z(n12554) );
  NANDN U13647 ( .A(n12555), .B(n12554), .Z(n12556) );
  AND U13648 ( .A(n12557), .B(n12556), .Z(n12559) );
  NANDN U13649 ( .A(n12559), .B(n12558), .Z(n12561) );
  ANDN U13650 ( .B(n12561), .A(n12560), .Z(n12563) );
  NANDN U13651 ( .A(n12563), .B(n12562), .Z(n12565) );
  ANDN U13652 ( .B(n12565), .A(n12564), .Z(n12567) );
  NANDN U13653 ( .A(n12567), .B(n12566), .Z(n12568) );
  NANDN U13654 ( .A(n12569), .B(n12568), .Z(n12570) );
  NANDN U13655 ( .A(n12571), .B(n12570), .Z(n12572) );
  NAND U13656 ( .A(n12573), .B(n12572), .Z(n12574) );
  NAND U13657 ( .A(n12575), .B(n12574), .Z(n12576) );
  AND U13658 ( .A(n12577), .B(n12576), .Z(n12579) );
  OR U13659 ( .A(n12579), .B(n12578), .Z(n12581) );
  ANDN U13660 ( .B(n12581), .A(n12580), .Z(n12583) );
  NANDN U13661 ( .A(n12583), .B(n12582), .Z(n12584) );
  NANDN U13662 ( .A(n12585), .B(n12584), .Z(n12586) );
  NAND U13663 ( .A(n12587), .B(n12586), .Z(n12588) );
  NAND U13664 ( .A(n12589), .B(n12588), .Z(n12590) );
  NANDN U13665 ( .A(n12591), .B(n12590), .Z(n12593) );
  ANDN U13666 ( .B(n12593), .A(n12592), .Z(n12594) );
  OR U13667 ( .A(n12595), .B(n12594), .Z(n12596) );
  NAND U13668 ( .A(n12597), .B(n12596), .Z(n12598) );
  NAND U13669 ( .A(n12599), .B(n12598), .Z(n12600) );
  NANDN U13670 ( .A(n12601), .B(n12600), .Z(n12602) );
  NANDN U13671 ( .A(n12603), .B(n12602), .Z(n12604) );
  NAND U13672 ( .A(n12605), .B(n12604), .Z(n12606) );
  NAND U13673 ( .A(n12607), .B(n12606), .Z(n12608) );
  NAND U13674 ( .A(n12609), .B(n12608), .Z(n12611) );
  ANDN U13675 ( .B(n12611), .A(n12610), .Z(n12612) );
  OR U13676 ( .A(n12613), .B(n12612), .Z(n12614) );
  NAND U13677 ( .A(n12615), .B(n12614), .Z(n12616) );
  NANDN U13678 ( .A(n12617), .B(n12616), .Z(n12618) );
  NANDN U13679 ( .A(n12619), .B(n12618), .Z(n12620) );
  NANDN U13680 ( .A(n12621), .B(n12620), .Z(n12622) );
  AND U13681 ( .A(n12623), .B(n12622), .Z(n12625) );
  OR U13682 ( .A(n12625), .B(n12624), .Z(n12627) );
  ANDN U13683 ( .B(n12627), .A(n12626), .Z(n12629) );
  NANDN U13684 ( .A(n12629), .B(n12628), .Z(n12631) );
  ANDN U13685 ( .B(n12631), .A(n12630), .Z(n12633) );
  NANDN U13686 ( .A(n12633), .B(n12632), .Z(n12634) );
  NANDN U13687 ( .A(n12635), .B(n12634), .Z(n12636) );
  NANDN U13688 ( .A(n12637), .B(n12636), .Z(n12638) );
  NAND U13689 ( .A(n12639), .B(n12638), .Z(n12641) );
  ANDN U13690 ( .B(n12641), .A(n12640), .Z(n12643) );
  OR U13691 ( .A(n12643), .B(n12642), .Z(n12644) );
  NAND U13692 ( .A(n12645), .B(n12644), .Z(n12646) );
  NANDN U13693 ( .A(n12647), .B(n12646), .Z(n12648) );
  AND U13694 ( .A(n12649), .B(n12648), .Z(n12651) );
  NANDN U13695 ( .A(n12651), .B(n12650), .Z(n12652) );
  NANDN U13696 ( .A(n12653), .B(n12652), .Z(n12654) );
  NAND U13697 ( .A(n12655), .B(n12654), .Z(n12656) );
  NAND U13698 ( .A(n12657), .B(n12656), .Z(n12658) );
  NAND U13699 ( .A(n12659), .B(n12658), .Z(n12660) );
  NAND U13700 ( .A(n12661), .B(n12660), .Z(n12662) );
  NAND U13701 ( .A(n12663), .B(n12662), .Z(n12664) );
  NAND U13702 ( .A(n12665), .B(n12664), .Z(n12666) );
  NANDN U13703 ( .A(n12667), .B(n12666), .Z(n12668) );
  NAND U13704 ( .A(n12669), .B(n12668), .Z(n12670) );
  NANDN U13705 ( .A(n12671), .B(n12670), .Z(n12672) );
  AND U13706 ( .A(n12673), .B(n12672), .Z(n12675) );
  NANDN U13707 ( .A(n12675), .B(n12674), .Z(n12676) );
  NANDN U13708 ( .A(n12677), .B(n12676), .Z(n12678) );
  NAND U13709 ( .A(n12679), .B(n12678), .Z(n12680) );
  NAND U13710 ( .A(n12681), .B(n12680), .Z(n12682) );
  NANDN U13711 ( .A(n12683), .B(n12682), .Z(n12684) );
  NAND U13712 ( .A(n12685), .B(n12684), .Z(n12687) );
  NAND U13713 ( .A(n12687), .B(n12686), .Z(n12688) );
  NANDN U13714 ( .A(n12689), .B(n12688), .Z(n12691) );
  ANDN U13715 ( .B(n12691), .A(n12690), .Z(n12693) );
  NANDN U13716 ( .A(n12693), .B(n12692), .Z(n12694) );
  AND U13717 ( .A(n12695), .B(n12694), .Z(n12696) );
  OR U13718 ( .A(n12697), .B(n12696), .Z(n12699) );
  ANDN U13719 ( .B(n12699), .A(n12698), .Z(n12701) );
  NANDN U13720 ( .A(n12701), .B(n12700), .Z(n12702) );
  NANDN U13721 ( .A(n12703), .B(n12702), .Z(n12704) );
  NANDN U13722 ( .A(n12705), .B(n12704), .Z(n12706) );
  NAND U13723 ( .A(n12707), .B(n12706), .Z(n12708) );
  NAND U13724 ( .A(n12709), .B(n12708), .Z(n12710) );
  NAND U13725 ( .A(n12711), .B(n12710), .Z(n12712) );
  NAND U13726 ( .A(n12713), .B(n12712), .Z(n12714) );
  NAND U13727 ( .A(n12715), .B(n12714), .Z(n12717) );
  ANDN U13728 ( .B(n12717), .A(n12716), .Z(n12719) );
  ANDN U13729 ( .B(n12719), .A(n12718), .Z(n12720) );
  OR U13730 ( .A(n12721), .B(n12720), .Z(n12723) );
  NANDN U13731 ( .A(n12723), .B(n12722), .Z(n12724) );
  NAND U13732 ( .A(n12725), .B(n12724), .Z(n12726) );
  NAND U13733 ( .A(n12727), .B(n12726), .Z(n12728) );
  NANDN U13734 ( .A(n12729), .B(n12728), .Z(n12730) );
  NAND U13735 ( .A(n12731), .B(n12730), .Z(n12733) );
  ANDN U13736 ( .B(n12733), .A(n12732), .Z(n12735) );
  NANDN U13737 ( .A(n12735), .B(n12734), .Z(n12736) );
  NAND U13738 ( .A(n12737), .B(n12736), .Z(n12738) );
  NANDN U13739 ( .A(n12739), .B(n12738), .Z(n12741) );
  NAND U13740 ( .A(n12741), .B(n12740), .Z(n12742) );
  NAND U13741 ( .A(n12743), .B(n12742), .Z(n12745) );
  ANDN U13742 ( .B(n12745), .A(n12744), .Z(n12747) );
  NANDN U13743 ( .A(n12747), .B(n12746), .Z(n12748) );
  NANDN U13744 ( .A(n12749), .B(n12748), .Z(n12750) );
  NAND U13745 ( .A(n12751), .B(n12750), .Z(n12752) );
  NANDN U13746 ( .A(n12753), .B(n12752), .Z(n12754) );
  NAND U13747 ( .A(n12755), .B(n12754), .Z(n12756) );
  AND U13748 ( .A(n12757), .B(n12756), .Z(n12759) );
  NANDN U13749 ( .A(n12759), .B(n12758), .Z(n12760) );
  NAND U13750 ( .A(n12761), .B(n12760), .Z(n12762) );
  NAND U13751 ( .A(n12763), .B(n12762), .Z(n12764) );
  NANDN U13752 ( .A(n12765), .B(n12764), .Z(n12766) );
  NAND U13753 ( .A(n12767), .B(n12766), .Z(n12769) );
  ANDN U13754 ( .B(n12769), .A(n12768), .Z(n12771) );
  NANDN U13755 ( .A(n12771), .B(n12770), .Z(n12772) );
  NANDN U13756 ( .A(n12773), .B(n12772), .Z(n12774) );
  NAND U13757 ( .A(n12775), .B(n12774), .Z(n12776) );
  NANDN U13758 ( .A(n12777), .B(n12776), .Z(n12778) );
  NAND U13759 ( .A(n12779), .B(n12778), .Z(n12781) );
  ANDN U13760 ( .B(n12781), .A(n12780), .Z(n12782) );
  OR U13761 ( .A(n12783), .B(n12782), .Z(n12784) );
  NAND U13762 ( .A(n12785), .B(n12784), .Z(n12786) );
  NANDN U13763 ( .A(n12787), .B(n12786), .Z(n12788) );
  NANDN U13764 ( .A(n12789), .B(n12788), .Z(n12790) );
  NAND U13765 ( .A(n12791), .B(n12790), .Z(n12793) );
  ANDN U13766 ( .B(n12793), .A(n12792), .Z(n12795) );
  NANDN U13767 ( .A(n12795), .B(n12794), .Z(n12796) );
  NANDN U13768 ( .A(n12797), .B(n12796), .Z(n12798) );
  NANDN U13769 ( .A(n12799), .B(n12798), .Z(n12800) );
  NAND U13770 ( .A(n12801), .B(n12800), .Z(n12802) );
  AND U13771 ( .A(n12803), .B(n12802), .Z(n12804) );
  OR U13772 ( .A(n12805), .B(n12804), .Z(n12806) );
  NANDN U13773 ( .A(n12807), .B(n12806), .Z(n12808) );
  NAND U13774 ( .A(n12809), .B(n12808), .Z(n12810) );
  NANDN U13775 ( .A(n12811), .B(n12810), .Z(n12812) );
  NAND U13776 ( .A(n12813), .B(n12812), .Z(n12815) );
  ANDN U13777 ( .B(n12815), .A(n12814), .Z(n12817) );
  NANDN U13778 ( .A(n12817), .B(n12816), .Z(n12818) );
  NANDN U13779 ( .A(n12819), .B(n12818), .Z(n12820) );
  NAND U13780 ( .A(n12821), .B(n12820), .Z(n12822) );
  NANDN U13781 ( .A(n12823), .B(n12822), .Z(n12824) );
  NANDN U13782 ( .A(n12825), .B(n12824), .Z(n12827) );
  NAND U13783 ( .A(n12827), .B(n12826), .Z(n12828) );
  NANDN U13784 ( .A(n12829), .B(n12828), .Z(n12830) );
  AND U13785 ( .A(n12831), .B(n12830), .Z(n12833) );
  NANDN U13786 ( .A(n12833), .B(n12832), .Z(n12834) );
  NANDN U13787 ( .A(n12835), .B(n12834), .Z(n12837) );
  ANDN U13788 ( .B(n12837), .A(n12836), .Z(n12839) );
  NANDN U13789 ( .A(n12839), .B(n12838), .Z(n12841) );
  ANDN U13790 ( .B(n12841), .A(n12840), .Z(n12843) );
  NANDN U13791 ( .A(n12843), .B(n12842), .Z(n12844) );
  NANDN U13792 ( .A(n12845), .B(n12844), .Z(n12846) );
  NANDN U13793 ( .A(n12847), .B(n12846), .Z(n12848) );
  NANDN U13794 ( .A(n12849), .B(n12848), .Z(n12850) );
  NAND U13795 ( .A(n12851), .B(n12850), .Z(n12853) );
  ANDN U13796 ( .B(n12853), .A(n12852), .Z(n12855) );
  NANDN U13797 ( .A(n12855), .B(n12854), .Z(n12856) );
  NANDN U13798 ( .A(n12857), .B(n12856), .Z(n12858) );
  NANDN U13799 ( .A(n12859), .B(n12858), .Z(n12860) );
  NAND U13800 ( .A(n12861), .B(n12860), .Z(n12862) );
  NANDN U13801 ( .A(n12863), .B(n12862), .Z(n12864) );
  NANDN U13802 ( .A(n12865), .B(n12864), .Z(n12866) );
  NAND U13803 ( .A(n12867), .B(n12866), .Z(n12868) );
  NAND U13804 ( .A(n12869), .B(n12868), .Z(n12871) );
  ANDN U13805 ( .B(n12871), .A(n12870), .Z(n12873) );
  NANDN U13806 ( .A(n12873), .B(n12872), .Z(n12875) );
  ANDN U13807 ( .B(n12875), .A(n12874), .Z(n12877) );
  NANDN U13808 ( .A(n12877), .B(n12876), .Z(n12878) );
  NANDN U13809 ( .A(n12879), .B(n12878), .Z(n12880) );
  NANDN U13810 ( .A(n12881), .B(n12880), .Z(n12882) );
  NANDN U13811 ( .A(n12883), .B(n12882), .Z(n12884) );
  NAND U13812 ( .A(n12885), .B(n12884), .Z(n12887) );
  ANDN U13813 ( .B(n12887), .A(n12886), .Z(n12889) );
  NANDN U13814 ( .A(n12889), .B(n12888), .Z(n12890) );
  NANDN U13815 ( .A(n12891), .B(n12890), .Z(n12892) );
  NANDN U13816 ( .A(n12893), .B(n12892), .Z(n12894) );
  NAND U13817 ( .A(n12895), .B(n12894), .Z(n12896) );
  NANDN U13818 ( .A(n12897), .B(n12896), .Z(n12898) );
  AND U13819 ( .A(n12899), .B(n12898), .Z(n12900) );
  OR U13820 ( .A(n12901), .B(n12900), .Z(n12902) );
  NAND U13821 ( .A(n12903), .B(n12902), .Z(n12904) );
  NAND U13822 ( .A(n12905), .B(n12904), .Z(n12906) );
  NANDN U13823 ( .A(n12907), .B(n12906), .Z(n12909) );
  ANDN U13824 ( .B(n12909), .A(n12908), .Z(n12911) );
  NANDN U13825 ( .A(n12911), .B(n12910), .Z(n12912) );
  NANDN U13826 ( .A(n12913), .B(n12912), .Z(n12914) );
  NAND U13827 ( .A(n12915), .B(n12914), .Z(n12916) );
  NANDN U13828 ( .A(n12917), .B(n12916), .Z(n12918) );
  NANDN U13829 ( .A(n12919), .B(n12918), .Z(n12920) );
  NAND U13830 ( .A(n12921), .B(n12920), .Z(n12922) );
  NANDN U13831 ( .A(n12923), .B(n12922), .Z(n12924) );
  NAND U13832 ( .A(n12925), .B(n12924), .Z(n12927) );
  ANDN U13833 ( .B(n12927), .A(n12926), .Z(n12928) );
  OR U13834 ( .A(n12929), .B(n12928), .Z(n12930) );
  NAND U13835 ( .A(n12931), .B(n12930), .Z(n12932) );
  NANDN U13836 ( .A(n12933), .B(n12932), .Z(n12934) );
  NAND U13837 ( .A(n12935), .B(n12934), .Z(n12936) );
  AND U13838 ( .A(n12937), .B(n12936), .Z(n12938) );
  OR U13839 ( .A(n12939), .B(n12938), .Z(n12940) );
  NAND U13840 ( .A(n12941), .B(n12940), .Z(n12942) );
  NAND U13841 ( .A(n12943), .B(n12942), .Z(n12944) );
  NAND U13842 ( .A(n12945), .B(n12944), .Z(n12946) );
  NAND U13843 ( .A(n12947), .B(n12946), .Z(n12948) );
  AND U13844 ( .A(n12949), .B(n12948), .Z(n12950) );
  OR U13845 ( .A(n12951), .B(n12950), .Z(n12952) );
  NAND U13846 ( .A(n12953), .B(n12952), .Z(n12954) );
  NANDN U13847 ( .A(n12955), .B(n12954), .Z(n12956) );
  NAND U13848 ( .A(n12957), .B(n12956), .Z(n12959) );
  ANDN U13849 ( .B(n12959), .A(n12958), .Z(n12961) );
  NANDN U13850 ( .A(n12961), .B(n12960), .Z(n12962) );
  NAND U13851 ( .A(n12963), .B(n12962), .Z(n12965) );
  ANDN U13852 ( .B(n12965), .A(n12964), .Z(n12967) );
  NANDN U13853 ( .A(n12967), .B(n12966), .Z(n12968) );
  NANDN U13854 ( .A(n12969), .B(n12968), .Z(n12970) );
  NANDN U13855 ( .A(n12971), .B(n12970), .Z(n12972) );
  AND U13856 ( .A(n12973), .B(n12972), .Z(n12974) );
  OR U13857 ( .A(n12975), .B(n12974), .Z(n12976) );
  NANDN U13858 ( .A(n12977), .B(n12976), .Z(n12978) );
  NANDN U13859 ( .A(n12979), .B(n12978), .Z(n12980) );
  NAND U13860 ( .A(n12981), .B(n12980), .Z(n12982) );
  NAND U13861 ( .A(n12983), .B(n12982), .Z(n12985) );
  ANDN U13862 ( .B(n12985), .A(n12984), .Z(n12987) );
  NANDN U13863 ( .A(n12987), .B(n12986), .Z(n12989) );
  ANDN U13864 ( .B(n12989), .A(n12988), .Z(n12991) );
  OR U13865 ( .A(n12991), .B(n12990), .Z(n12992) );
  NAND U13866 ( .A(n12993), .B(n12992), .Z(n12994) );
  NANDN U13867 ( .A(n12995), .B(n12994), .Z(n12996) );
  AND U13868 ( .A(n12997), .B(n12996), .Z(n12999) );
  NANDN U13869 ( .A(n12999), .B(n12998), .Z(n13000) );
  NAND U13870 ( .A(n13001), .B(n13000), .Z(n13002) );
  NANDN U13871 ( .A(n13003), .B(n13002), .Z(n13004) );
  NAND U13872 ( .A(n13005), .B(n13004), .Z(n13006) );
  NAND U13873 ( .A(n13007), .B(n13006), .Z(n13008) );
  NANDN U13874 ( .A(n13009), .B(n13008), .Z(n13011) );
  AND U13875 ( .A(n13011), .B(n13010), .Z(n13015) );
  NANDN U13876 ( .A(n13013), .B(n13012), .Z(n13014) );
  AND U13877 ( .A(n13015), .B(n13014), .Z(n13016) );
  OR U13878 ( .A(n13017), .B(n13016), .Z(n13018) );
  NAND U13879 ( .A(n13019), .B(n13018), .Z(n13020) );
  NANDN U13880 ( .A(n13021), .B(n13020), .Z(n13022) );
  NAND U13881 ( .A(n13023), .B(n13022), .Z(n13024) );
  AND U13882 ( .A(n13025), .B(n13024), .Z(n13026) );
  ANDN U13883 ( .B(n13027), .A(n13026), .Z(n13029) );
  NANDN U13884 ( .A(n13029), .B(n13028), .Z(n13030) );
  NANDN U13885 ( .A(n13031), .B(n13030), .Z(n13032) );
  NAND U13886 ( .A(n13033), .B(n13032), .Z(n13035) );
  NAND U13887 ( .A(n13035), .B(n13034), .Z(n13036) );
  NANDN U13888 ( .A(n13037), .B(n13036), .Z(n13039) );
  ANDN U13889 ( .B(n13039), .A(n13038), .Z(n13041) );
  NANDN U13890 ( .A(n13041), .B(n13040), .Z(n13042) );
  AND U13891 ( .A(n13043), .B(n13042), .Z(n13045) );
  OR U13892 ( .A(n13045), .B(n13044), .Z(n13046) );
  NAND U13893 ( .A(n13047), .B(n13046), .Z(n13049) );
  ANDN U13894 ( .B(n13049), .A(n13048), .Z(n13051) );
  OR U13895 ( .A(n13051), .B(n13050), .Z(n13052) );
  AND U13896 ( .A(n13053), .B(n13052), .Z(n13055) );
  OR U13897 ( .A(n13055), .B(n13054), .Z(n13056) );
  AND U13898 ( .A(n13057), .B(n13056), .Z(n13059) );
  OR U13899 ( .A(n13059), .B(n13058), .Z(n13060) );
  AND U13900 ( .A(n13061), .B(n13060), .Z(n13063) );
  OR U13901 ( .A(n13063), .B(n13062), .Z(n13064) );
  NAND U13902 ( .A(n13065), .B(n13064), .Z(n13067) );
  ANDN U13903 ( .B(n13067), .A(n13066), .Z(n13068) );
  OR U13904 ( .A(n13069), .B(n13068), .Z(n13070) );
  NAND U13905 ( .A(n13071), .B(n13070), .Z(n13072) );
  NANDN U13906 ( .A(n13073), .B(n13072), .Z(n13074) );
  NANDN U13907 ( .A(n13075), .B(n13074), .Z(n13076) );
  NAND U13908 ( .A(n13077), .B(n13076), .Z(n13079) );
  ANDN U13909 ( .B(n13079), .A(n13078), .Z(n13081) );
  NANDN U13910 ( .A(n13081), .B(n13080), .Z(n13082) );
  NANDN U13911 ( .A(n13083), .B(n13082), .Z(n13084) );
  NANDN U13912 ( .A(n13085), .B(n13084), .Z(n13086) );
  NAND U13913 ( .A(n13087), .B(n13086), .Z(n13089) );
  ANDN U13914 ( .B(n13089), .A(n13088), .Z(n13091) );
  NANDN U13915 ( .A(n13091), .B(n13090), .Z(n13092) );
  NAND U13916 ( .A(n13093), .B(n13092), .Z(n13094) );
  NANDN U13917 ( .A(n13095), .B(n13094), .Z(n13096) );
  NAND U13918 ( .A(n13097), .B(n13096), .Z(n13098) );
  NANDN U13919 ( .A(n13099), .B(n13098), .Z(n13100) );
  NAND U13920 ( .A(n13101), .B(n13100), .Z(n13103) );
  ANDN U13921 ( .B(n13103), .A(n13102), .Z(n13104) );
  NANDN U13922 ( .A(n13105), .B(n13104), .Z(n13106) );
  NAND U13923 ( .A(n13107), .B(n13106), .Z(n13108) );
  AND U13924 ( .A(n13109), .B(n13108), .Z(n13111) );
  NANDN U13925 ( .A(n13111), .B(n13110), .Z(n13112) );
  NAND U13926 ( .A(n13113), .B(n13112), .Z(n13114) );
  AND U13927 ( .A(n13115), .B(n13114), .Z(n13117) );
  NANDN U13928 ( .A(n13117), .B(n13116), .Z(n13118) );
  NAND U13929 ( .A(n13119), .B(n13118), .Z(n13120) );
  NAND U13930 ( .A(n13121), .B(n13120), .Z(n13122) );
  NANDN U13931 ( .A(n13123), .B(n13122), .Z(n13124) );
  NAND U13932 ( .A(n13125), .B(n13124), .Z(n13126) );
  AND U13933 ( .A(n13127), .B(n13126), .Z(n13129) );
  NANDN U13934 ( .A(n13129), .B(n13128), .Z(n13130) );
  NAND U13935 ( .A(n13131), .B(n13130), .Z(n13132) );
  NANDN U13936 ( .A(n13133), .B(n13132), .Z(n13134) );
  NAND U13937 ( .A(n13135), .B(n13134), .Z(n13136) );
  NANDN U13938 ( .A(n13137), .B(n13136), .Z(n13138) );
  NANDN U13939 ( .A(n13139), .B(n13138), .Z(n13140) );
  NAND U13940 ( .A(n13141), .B(n13140), .Z(n13142) );
  NANDN U13941 ( .A(n13143), .B(n13142), .Z(n13145) );
  ANDN U13942 ( .B(n13145), .A(n13144), .Z(n13147) );
  NANDN U13943 ( .A(n13147), .B(n13146), .Z(n13148) );
  NANDN U13944 ( .A(n13149), .B(n13148), .Z(n13150) );
  NAND U13945 ( .A(n13151), .B(n13150), .Z(n13152) );
  NANDN U13946 ( .A(n13153), .B(n13152), .Z(n13154) );
  NAND U13947 ( .A(n13155), .B(n13154), .Z(n13156) );
  AND U13948 ( .A(n13157), .B(n13156), .Z(n13158) );
  OR U13949 ( .A(n13159), .B(n13158), .Z(n13160) );
  NAND U13950 ( .A(n13161), .B(n13160), .Z(n13162) );
  NANDN U13951 ( .A(n13163), .B(n13162), .Z(n13164) );
  NANDN U13952 ( .A(n13165), .B(n13164), .Z(n13166) );
  NAND U13953 ( .A(n13167), .B(n13166), .Z(n13168) );
  NANDN U13954 ( .A(n13169), .B(n13168), .Z(n13170) );
  NAND U13955 ( .A(n13171), .B(n13170), .Z(n13173) );
  ANDN U13956 ( .B(n13173), .A(n13172), .Z(n13175) );
  NANDN U13957 ( .A(n13175), .B(n13174), .Z(n13176) );
  NAND U13958 ( .A(n13177), .B(n13176), .Z(n13178) );
  NAND U13959 ( .A(n13179), .B(n13178), .Z(n13181) );
  ANDN U13960 ( .B(n13181), .A(n13180), .Z(n13183) );
  NANDN U13961 ( .A(n13183), .B(n13182), .Z(n13184) );
  NANDN U13962 ( .A(n13185), .B(n13184), .Z(n13186) );
  AND U13963 ( .A(n13187), .B(n13186), .Z(n13188) );
  OR U13964 ( .A(n13189), .B(n13188), .Z(n13190) );
  NAND U13965 ( .A(n13191), .B(n13190), .Z(n13192) );
  NANDN U13966 ( .A(n13193), .B(n13192), .Z(n13194) );
  NAND U13967 ( .A(n13195), .B(n13194), .Z(n13196) );
  NANDN U13968 ( .A(n13197), .B(n13196), .Z(n13198) );
  AND U13969 ( .A(n13199), .B(n13198), .Z(n13201) );
  OR U13970 ( .A(n13201), .B(n13200), .Z(n13203) );
  ANDN U13971 ( .B(n13203), .A(n13202), .Z(n13205) );
  NANDN U13972 ( .A(n13205), .B(n13204), .Z(n13206) );
  NAND U13973 ( .A(n13207), .B(n13206), .Z(n13208) );
  NAND U13974 ( .A(n13209), .B(n13208), .Z(n13210) );
  NAND U13975 ( .A(n13211), .B(n13210), .Z(n13212) );
  NAND U13976 ( .A(n13213), .B(n13212), .Z(n13215) );
  ANDN U13977 ( .B(n13215), .A(n13214), .Z(n13217) );
  NANDN U13978 ( .A(n13217), .B(n13216), .Z(n13218) );
  AND U13979 ( .A(n13219), .B(n13218), .Z(n13221) );
  NANDN U13980 ( .A(n13221), .B(n13220), .Z(n13222) );
  NANDN U13981 ( .A(n13223), .B(n13222), .Z(n13224) );
  NAND U13982 ( .A(n13225), .B(n13224), .Z(n13226) );
  NANDN U13983 ( .A(n13227), .B(n13226), .Z(n13228) );
  NAND U13984 ( .A(n13229), .B(n13228), .Z(n13231) );
  ANDN U13985 ( .B(n13231), .A(n13230), .Z(n13233) );
  OR U13986 ( .A(n13233), .B(n13232), .Z(n13235) );
  ANDN U13987 ( .B(n13235), .A(n13234), .Z(n13237) );
  NANDN U13988 ( .A(n13237), .B(n13236), .Z(n13239) );
  ANDN U13989 ( .B(n13239), .A(n13238), .Z(n13241) );
  NANDN U13990 ( .A(n13241), .B(n13240), .Z(n13242) );
  NANDN U13991 ( .A(n13243), .B(n13242), .Z(n13244) );
  NANDN U13992 ( .A(n13245), .B(n13244), .Z(n13246) );
  NAND U13993 ( .A(n13247), .B(n13246), .Z(n13248) );
  NANDN U13994 ( .A(n13249), .B(n13248), .Z(n13250) );
  NANDN U13995 ( .A(n13251), .B(n13250), .Z(n13252) );
  NANDN U13996 ( .A(n13253), .B(n13252), .Z(n13254) );
  NAND U13997 ( .A(n13255), .B(n13254), .Z(n13256) );
  NANDN U13998 ( .A(n13257), .B(n13256), .Z(n13258) );
  AND U13999 ( .A(n13259), .B(n13258), .Z(n13261) );
  NANDN U14000 ( .A(n13261), .B(n13260), .Z(n13263) );
  ANDN U14001 ( .B(n13263), .A(n13262), .Z(n13265) );
  NANDN U14002 ( .A(n13265), .B(n13264), .Z(n13267) );
  ANDN U14003 ( .B(n13267), .A(n13266), .Z(n13269) );
  NANDN U14004 ( .A(n13269), .B(n13268), .Z(n13270) );
  NANDN U14005 ( .A(n13271), .B(n13270), .Z(n13272) );
  NAND U14006 ( .A(n13273), .B(n13272), .Z(n13275) );
  NAND U14007 ( .A(n13275), .B(n13274), .Z(n13276) );
  NANDN U14008 ( .A(n13277), .B(n13276), .Z(n13278) );
  AND U14009 ( .A(n13279), .B(n13278), .Z(n13280) );
  OR U14010 ( .A(n13281), .B(n13280), .Z(n13282) );
  NANDN U14011 ( .A(n13283), .B(n13282), .Z(n13284) );
  NAND U14012 ( .A(n13285), .B(n13284), .Z(n13287) );
  AND U14013 ( .A(n13287), .B(n13286), .Z(n13289) );
  NANDN U14014 ( .A(n13289), .B(n13288), .Z(n13290) );
  NAND U14015 ( .A(n13291), .B(n13290), .Z(n13292) );
  NANDN U14016 ( .A(n13293), .B(n13292), .Z(n13294) );
  AND U14017 ( .A(n13295), .B(n13294), .Z(n13297) );
  NANDN U14018 ( .A(n13297), .B(n13296), .Z(n13298) );
  NAND U14019 ( .A(n13299), .B(n13298), .Z(n13300) );
  NAND U14020 ( .A(n13301), .B(n13300), .Z(n13302) );
  NANDN U14021 ( .A(n13303), .B(n13302), .Z(n13304) );
  NAND U14022 ( .A(n13305), .B(n13304), .Z(n13307) );
  ANDN U14023 ( .B(n13307), .A(n13306), .Z(n13309) );
  NANDN U14024 ( .A(n13309), .B(n13308), .Z(n13310) );
  NAND U14025 ( .A(n13311), .B(n13310), .Z(n13312) );
  NANDN U14026 ( .A(n13313), .B(n13312), .Z(n13314) );
  NAND U14027 ( .A(n13315), .B(n13314), .Z(n13316) );
  NAND U14028 ( .A(n13317), .B(n13316), .Z(n13318) );
  NANDN U14029 ( .A(n13319), .B(n13318), .Z(n13320) );
  NAND U14030 ( .A(n13321), .B(n13320), .Z(n13323) );
  NANDN U14031 ( .A(n13323), .B(n13322), .Z(n13324) );
  NANDN U14032 ( .A(n13325), .B(n13324), .Z(n13326) );
  NAND U14033 ( .A(n13327), .B(n13326), .Z(n13328) );
  NAND U14034 ( .A(n13329), .B(n13328), .Z(n13330) );
  NANDN U14035 ( .A(n13331), .B(n13330), .Z(n13332) );
  NAND U14036 ( .A(n13333), .B(n13332), .Z(n13334) );
  NANDN U14037 ( .A(n13335), .B(n13334), .Z(n13336) );
  NANDN U14038 ( .A(n13337), .B(n13336), .Z(n13338) );
  AND U14039 ( .A(n13339), .B(n13338), .Z(n13340) );
  OR U14040 ( .A(n13341), .B(n13340), .Z(n13342) );
  NAND U14041 ( .A(n13343), .B(n13342), .Z(n13344) );
  NANDN U14042 ( .A(n13345), .B(n13344), .Z(n13346) );
  NAND U14043 ( .A(n13347), .B(n13346), .Z(n13348) );
  NAND U14044 ( .A(n13349), .B(n13348), .Z(n13350) );
  AND U14045 ( .A(n13351), .B(n13350), .Z(n13353) );
  NANDN U14046 ( .A(n13353), .B(n13352), .Z(n13354) );
  NANDN U14047 ( .A(n13355), .B(n13354), .Z(n13356) );
  NANDN U14048 ( .A(n13357), .B(n13356), .Z(n13358) );
  NAND U14049 ( .A(n13359), .B(n13358), .Z(n13360) );
  NAND U14050 ( .A(n13361), .B(n13360), .Z(n13362) );
  NAND U14051 ( .A(n13363), .B(n13362), .Z(n13364) );
  NANDN U14052 ( .A(n13365), .B(n13364), .Z(n13366) );
  NAND U14053 ( .A(n13367), .B(n13366), .Z(n13368) );
  AND U14054 ( .A(n13369), .B(n13368), .Z(n13371) );
  OR U14055 ( .A(n13371), .B(n13370), .Z(n13372) );
  AND U14056 ( .A(n13373), .B(n13372), .Z(n13374) );
  OR U14057 ( .A(n13375), .B(n13374), .Z(n13377) );
  ANDN U14058 ( .B(n13377), .A(n13376), .Z(n13379) );
  NANDN U14059 ( .A(n13379), .B(n13378), .Z(n13380) );
  NANDN U14060 ( .A(n13381), .B(n13380), .Z(n13382) );
  NANDN U14061 ( .A(n13383), .B(n13382), .Z(n13384) );
  NAND U14062 ( .A(n13385), .B(n13384), .Z(n13386) );
  NANDN U14063 ( .A(n13387), .B(n13386), .Z(n13388) );
  AND U14064 ( .A(n13389), .B(n13388), .Z(n13391) );
  NANDN U14065 ( .A(n13391), .B(n13390), .Z(n13392) );
  NAND U14066 ( .A(n13393), .B(n13392), .Z(n13394) );
  NANDN U14067 ( .A(n13395), .B(n13394), .Z(n13396) );
  AND U14068 ( .A(n13397), .B(n13396), .Z(n13399) );
  NANDN U14069 ( .A(n13399), .B(n13398), .Z(n13400) );
  NAND U14070 ( .A(n13401), .B(n13400), .Z(n13402) );
  NAND U14071 ( .A(n13403), .B(n13402), .Z(n13404) );
  NANDN U14072 ( .A(n13405), .B(n13404), .Z(n13406) );
  NAND U14073 ( .A(n13407), .B(n13406), .Z(n13408) );
  AND U14074 ( .A(n13409), .B(n13408), .Z(n13411) );
  NANDN U14075 ( .A(n13411), .B(n13410), .Z(n13412) );
  NANDN U14076 ( .A(n13413), .B(n13412), .Z(n13415) );
  ANDN U14077 ( .B(n13415), .A(n13414), .Z(n13417) );
  NANDN U14078 ( .A(n13417), .B(n13416), .Z(n13418) );
  NAND U14079 ( .A(n13419), .B(n13418), .Z(n13420) );
  NANDN U14080 ( .A(n13421), .B(n13420), .Z(n13422) );
  NAND U14081 ( .A(n13423), .B(n13422), .Z(n13424) );
  NANDN U14082 ( .A(n13425), .B(n13424), .Z(n13427) );
  ANDN U14083 ( .B(n13427), .A(n13426), .Z(n13429) );
  NANDN U14084 ( .A(n13429), .B(n13428), .Z(n13430) );
  NANDN U14085 ( .A(n13431), .B(n13430), .Z(n13432) );
  NANDN U14086 ( .A(n13433), .B(n13432), .Z(n13434) );
  NANDN U14087 ( .A(n13435), .B(n13434), .Z(n13436) );
  NANDN U14088 ( .A(n13437), .B(n13436), .Z(n13438) );
  NANDN U14089 ( .A(n13439), .B(n13438), .Z(n13440) );
  NANDN U14090 ( .A(n13441), .B(n13440), .Z(n13443) );
  NAND U14091 ( .A(n13443), .B(n13442), .Z(n13444) );
  NANDN U14092 ( .A(n13445), .B(n13444), .Z(n13446) );
  AND U14093 ( .A(n13447), .B(n13446), .Z(n13449) );
  NANDN U14094 ( .A(n13449), .B(n13448), .Z(n13450) );
  NANDN U14095 ( .A(n13451), .B(n13450), .Z(n13452) );
  NAND U14096 ( .A(n13453), .B(n13452), .Z(n13454) );
  NAND U14097 ( .A(n13455), .B(n13454), .Z(n13456) );
  NAND U14098 ( .A(n13457), .B(n13456), .Z(n13459) );
  ANDN U14099 ( .B(n13459), .A(n13458), .Z(n13461) );
  NANDN U14100 ( .A(n13461), .B(n13460), .Z(n13462) );
  AND U14101 ( .A(n13463), .B(n13462), .Z(n13465) );
  NANDN U14102 ( .A(n13465), .B(n13464), .Z(n13466) );
  AND U14103 ( .A(n13467), .B(n13466), .Z(n13469) );
  NANDN U14104 ( .A(n13469), .B(n13468), .Z(n13470) );
  NAND U14105 ( .A(n13471), .B(n13470), .Z(n13472) );
  NAND U14106 ( .A(n13473), .B(n13472), .Z(n13474) );
  NAND U14107 ( .A(n13475), .B(n13474), .Z(n13476) );
  NAND U14108 ( .A(n13477), .B(n13476), .Z(n13478) );
  NANDN U14109 ( .A(n13479), .B(n13478), .Z(n13481) );
  NAND U14110 ( .A(n13481), .B(n13480), .Z(n13482) );
  NANDN U14111 ( .A(n13483), .B(n13482), .Z(n13484) );
  AND U14112 ( .A(n13485), .B(n13484), .Z(n13486) );
  OR U14113 ( .A(n13487), .B(n13486), .Z(n13488) );
  NAND U14114 ( .A(n13489), .B(n13488), .Z(n13490) );
  NANDN U14115 ( .A(n13491), .B(n13490), .Z(n13492) );
  NAND U14116 ( .A(n13493), .B(n13492), .Z(n13494) );
  NANDN U14117 ( .A(n13495), .B(n13494), .Z(n13496) );
  NANDN U14118 ( .A(n13497), .B(n13496), .Z(n13498) );
  NAND U14119 ( .A(n13499), .B(n13498), .Z(n13500) );
  NANDN U14120 ( .A(n13501), .B(n13500), .Z(n13502) );
  AND U14121 ( .A(n13503), .B(n13502), .Z(n13504) );
  OR U14122 ( .A(n13505), .B(n13504), .Z(n13506) );
  AND U14123 ( .A(n13507), .B(n13506), .Z(n13509) );
  OR U14124 ( .A(n13509), .B(n13508), .Z(n13511) );
  NAND U14125 ( .A(n13511), .B(n13510), .Z(n13512) );
  NANDN U14126 ( .A(n13513), .B(n13512), .Z(n13514) );
  AND U14127 ( .A(n13515), .B(n13514), .Z(n13517) );
  NANDN U14128 ( .A(n13517), .B(n13516), .Z(n13518) );
  NANDN U14129 ( .A(n13519), .B(n13518), .Z(n13520) );
  AND U14130 ( .A(n13521), .B(n13520), .Z(n13523) );
  NANDN U14131 ( .A(n13523), .B(n13522), .Z(n13524) );
  NAND U14132 ( .A(n13525), .B(n13524), .Z(n13526) );
  NAND U14133 ( .A(n13527), .B(n13526), .Z(n13528) );
  AND U14134 ( .A(n13529), .B(n13528), .Z(n13531) );
  NANDN U14135 ( .A(n13531), .B(n13530), .Z(n13532) );
  NANDN U14136 ( .A(n13533), .B(n13532), .Z(n13534) );
  NAND U14137 ( .A(n13535), .B(n13534), .Z(n13536) );
  NANDN U14138 ( .A(n13537), .B(n13536), .Z(n13539) );
  NAND U14139 ( .A(n13539), .B(n13538), .Z(n13540) );
  NAND U14140 ( .A(n13541), .B(n13540), .Z(n13543) );
  ANDN U14141 ( .B(n13543), .A(n13542), .Z(n13545) );
  OR U14142 ( .A(n13545), .B(n13544), .Z(n13546) );
  AND U14143 ( .A(n13547), .B(n13546), .Z(n13549) );
  NANDN U14144 ( .A(n13549), .B(n13548), .Z(n13550) );
  NANDN U14145 ( .A(n13551), .B(n13550), .Z(n13552) );
  NAND U14146 ( .A(n13553), .B(n13552), .Z(n13554) );
  NANDN U14147 ( .A(n13555), .B(n13554), .Z(n13556) );
  NAND U14148 ( .A(n13557), .B(n13556), .Z(n13559) );
  ANDN U14149 ( .B(n13559), .A(n13558), .Z(n13561) );
  NANDN U14150 ( .A(n13561), .B(n13560), .Z(n13562) );
  NANDN U14151 ( .A(n13563), .B(n13562), .Z(n13564) );
  NANDN U14152 ( .A(n13565), .B(n13564), .Z(n13566) );
  NAND U14153 ( .A(n13567), .B(n13566), .Z(n13568) );
  NANDN U14154 ( .A(n13569), .B(n13568), .Z(n13570) );
  AND U14155 ( .A(n13571), .B(n13570), .Z(n13572) );
  OR U14156 ( .A(n13573), .B(n13572), .Z(n13574) );
  NAND U14157 ( .A(n13575), .B(n13574), .Z(n13576) );
  NANDN U14158 ( .A(n13577), .B(n13576), .Z(n13579) );
  NANDN U14159 ( .A(n13579), .B(n13578), .Z(n13580) );
  NANDN U14160 ( .A(n13581), .B(n13580), .Z(n13582) );
  NAND U14161 ( .A(n13583), .B(n13582), .Z(n13584) );
  NAND U14162 ( .A(n13585), .B(n13584), .Z(n13586) );
  NAND U14163 ( .A(n13587), .B(n13586), .Z(n13588) );
  NANDN U14164 ( .A(n13589), .B(n13588), .Z(n13590) );
  NAND U14165 ( .A(n13591), .B(n13590), .Z(n13592) );
  NANDN U14166 ( .A(n13593), .B(n13592), .Z(n13594) );
  NANDN U14167 ( .A(n13595), .B(n13594), .Z(n13596) );
  AND U14168 ( .A(n13597), .B(n13596), .Z(n13599) );
  NANDN U14169 ( .A(n13599), .B(n13598), .Z(n13601) );
  ANDN U14170 ( .B(n13601), .A(n13600), .Z(n13603) );
  NANDN U14171 ( .A(n13603), .B(n13602), .Z(n13604) );
  NANDN U14172 ( .A(n13605), .B(n13604), .Z(n13606) );
  NAND U14173 ( .A(n13607), .B(n13606), .Z(n13608) );
  NAND U14174 ( .A(n13609), .B(n13608), .Z(n13611) );
  ANDN U14175 ( .B(n13611), .A(n13610), .Z(n13613) );
  NANDN U14176 ( .A(n13613), .B(n13612), .Z(n13614) );
  NANDN U14177 ( .A(n13615), .B(n13614), .Z(n13616) );
  NANDN U14178 ( .A(n13617), .B(n13616), .Z(n13618) );
  NANDN U14179 ( .A(n13619), .B(n13618), .Z(n13620) );
  NANDN U14180 ( .A(n13621), .B(n13620), .Z(n13622) );
  NAND U14181 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U14182 ( .A(n13625), .B(n13624), .Z(n13627) );
  NANDN U14183 ( .A(n13627), .B(n13626), .Z(n13628) );
  AND U14184 ( .A(n13629), .B(n13628), .Z(n13631) );
  NANDN U14185 ( .A(n13631), .B(n13630), .Z(n13632) );
  NANDN U14186 ( .A(n13633), .B(n13632), .Z(n13634) );
  NAND U14187 ( .A(n13635), .B(n13634), .Z(n13637) );
  ANDN U14188 ( .B(n13637), .A(n13636), .Z(n13639) );
  NANDN U14189 ( .A(n13639), .B(n13638), .Z(n13640) );
  NANDN U14190 ( .A(n13641), .B(n13640), .Z(n13642) );
  NANDN U14191 ( .A(n13643), .B(n13642), .Z(n13645) );
  NANDN U14192 ( .A(n13645), .B(n13644), .Z(n13646) );
  NANDN U14193 ( .A(n13647), .B(n13646), .Z(n13648) );
  NAND U14194 ( .A(n13649), .B(n13648), .Z(n13650) );
  NANDN U14195 ( .A(n13651), .B(n13650), .Z(n13652) );
  NANDN U14196 ( .A(n13653), .B(n13652), .Z(n13654) );
  AND U14197 ( .A(n13655), .B(n13654), .Z(n13656) );
  OR U14198 ( .A(n13657), .B(n13656), .Z(n13658) );
  NAND U14199 ( .A(n13659), .B(n13658), .Z(n13660) );
  NAND U14200 ( .A(n13661), .B(n13660), .Z(n13662) );
  NANDN U14201 ( .A(n13663), .B(n13662), .Z(n13664) );
  NAND U14202 ( .A(n13665), .B(n13664), .Z(n13666) );
  NAND U14203 ( .A(n13667), .B(n13666), .Z(n13671) );
  NAND U14204 ( .A(n13669), .B(n13668), .Z(n13670) );
  NANDN U14205 ( .A(n13671), .B(n13670), .Z(n13673) );
  ANDN U14206 ( .B(n13673), .A(n13672), .Z(n13675) );
  NANDN U14207 ( .A(n13675), .B(n13674), .Z(n13676) );
  NANDN U14208 ( .A(n13677), .B(n13676), .Z(n13678) );
  NANDN U14209 ( .A(n13679), .B(n13678), .Z(n13681) );
  ANDN U14210 ( .B(n13681), .A(n13680), .Z(n13683) );
  NANDN U14211 ( .A(n13683), .B(n13682), .Z(n13684) );
  NANDN U14212 ( .A(n13685), .B(n13684), .Z(n13686) );
  AND U14213 ( .A(n13687), .B(n13686), .Z(n13689) );
  NANDN U14214 ( .A(n13689), .B(n13688), .Z(n13691) );
  ANDN U14215 ( .B(n13691), .A(n13690), .Z(n13693) );
  NANDN U14216 ( .A(n13693), .B(n13692), .Z(n13694) );
  NANDN U14217 ( .A(n13695), .B(n13694), .Z(n13696) );
  NANDN U14218 ( .A(n13697), .B(n13696), .Z(n13698) );
  NAND U14219 ( .A(n13699), .B(n13698), .Z(n13701) );
  ANDN U14220 ( .B(n13701), .A(n13700), .Z(n13703) );
  NANDN U14221 ( .A(n13703), .B(n13702), .Z(n13704) );
  NANDN U14222 ( .A(n13705), .B(n13704), .Z(n13706) );
  NAND U14223 ( .A(n13707), .B(n13706), .Z(n13708) );
  NAND U14224 ( .A(n13709), .B(n13708), .Z(n13710) );
  NANDN U14225 ( .A(n13711), .B(n13710), .Z(n13712) );
  AND U14226 ( .A(n13713), .B(n13712), .Z(n13715) );
  NANDN U14227 ( .A(n13715), .B(n13714), .Z(n13717) );
  ANDN U14228 ( .B(n13717), .A(n13716), .Z(n13718) );
  OR U14229 ( .A(n13719), .B(n13718), .Z(n13720) );
  NAND U14230 ( .A(n13721), .B(n13720), .Z(n13722) );
  NAND U14231 ( .A(n13723), .B(n13722), .Z(n13725) );
  AND U14232 ( .A(n13725), .B(n13724), .Z(n13726) );
  NANDN U14233 ( .A(n13727), .B(n13726), .Z(n13728) );
  NANDN U14234 ( .A(n13729), .B(n13728), .Z(n13730) );
  NAND U14235 ( .A(n13731), .B(n13730), .Z(n13733) );
  ANDN U14236 ( .B(n13733), .A(n13732), .Z(n13735) );
  NANDN U14237 ( .A(n13735), .B(n13734), .Z(n13736) );
  NANDN U14238 ( .A(n13737), .B(n13736), .Z(n13738) );
  NANDN U14239 ( .A(n13739), .B(n13738), .Z(n13740) );
  NAND U14240 ( .A(n13741), .B(n13740), .Z(n13743) );
  ANDN U14241 ( .B(n13743), .A(n13742), .Z(n13745) );
  NANDN U14242 ( .A(n13745), .B(n13744), .Z(n13746) );
  NANDN U14243 ( .A(n13747), .B(n13746), .Z(n13748) );
  NANDN U14244 ( .A(n13749), .B(n13748), .Z(n13750) );
  NANDN U14245 ( .A(n13751), .B(n13750), .Z(n13752) );
  NAND U14246 ( .A(n13753), .B(n13752), .Z(n13755) );
  ANDN U14247 ( .B(n13755), .A(n13754), .Z(n13757) );
  NANDN U14248 ( .A(n13757), .B(n13756), .Z(n13758) );
  NANDN U14249 ( .A(n13759), .B(n13758), .Z(n13760) );
  NANDN U14250 ( .A(n13761), .B(n13760), .Z(n13762) );
  NAND U14251 ( .A(n13763), .B(n13762), .Z(n13764) );
  NANDN U14252 ( .A(n13765), .B(n13764), .Z(n13766) );
  NAND U14253 ( .A(n13767), .B(n13766), .Z(n13768) );
  AND U14254 ( .A(n13769), .B(n13768), .Z(n13770) );
  NANDN U14255 ( .A(n13771), .B(n13770), .Z(n13772) );
  NAND U14256 ( .A(n13773), .B(n13772), .Z(n13774) );
  NAND U14257 ( .A(n13775), .B(n13774), .Z(n13776) );
  NANDN U14258 ( .A(n13777), .B(n13776), .Z(n13778) );
  AND U14259 ( .A(n13779), .B(n13778), .Z(n13781) );
  NANDN U14260 ( .A(n13781), .B(n13780), .Z(n13782) );
  NANDN U14261 ( .A(n13783), .B(n13782), .Z(n13784) );
  NAND U14262 ( .A(n13785), .B(n13784), .Z(n13786) );
  NAND U14263 ( .A(n13787), .B(n13786), .Z(n13788) );
  NAND U14264 ( .A(n13789), .B(n13788), .Z(n13790) );
  NANDN U14265 ( .A(n13791), .B(n13790), .Z(n13793) );
  AND U14266 ( .A(n13793), .B(n13792), .Z(n13797) );
  NANDN U14267 ( .A(n13795), .B(n13794), .Z(n13796) );
  AND U14268 ( .A(n13797), .B(n13796), .Z(n13798) );
  OR U14269 ( .A(n13799), .B(n13798), .Z(n13800) );
  NAND U14270 ( .A(n13801), .B(n13800), .Z(n13802) );
  NANDN U14271 ( .A(n13803), .B(n13802), .Z(n13804) );
  NAND U14272 ( .A(n13805), .B(n13804), .Z(n13806) );
  NANDN U14273 ( .A(n13807), .B(n13806), .Z(n13808) );
  AND U14274 ( .A(n13809), .B(n13808), .Z(n13811) );
  OR U14275 ( .A(n13811), .B(n13810), .Z(n13812) );
  NAND U14276 ( .A(n13813), .B(n13812), .Z(n13814) );
  NANDN U14277 ( .A(n13815), .B(n13814), .Z(n13816) );
  NAND U14278 ( .A(n13817), .B(n13816), .Z(n13818) );
  NANDN U14279 ( .A(n13819), .B(n13818), .Z(n13820) );
  AND U14280 ( .A(n13821), .B(n13820), .Z(n13822) );
  OR U14281 ( .A(n13823), .B(n13822), .Z(n13824) );
  NAND U14282 ( .A(n13825), .B(n13824), .Z(n13826) );
  NANDN U14283 ( .A(n13827), .B(n13826), .Z(n13828) );
  NAND U14284 ( .A(n13829), .B(n13828), .Z(n13830) );
  AND U14285 ( .A(n13831), .B(n13830), .Z(n13833) );
  NANDN U14286 ( .A(n13833), .B(n13832), .Z(n13834) );
  NANDN U14287 ( .A(n13835), .B(n13834), .Z(n13836) );
  NANDN U14288 ( .A(n13837), .B(n13836), .Z(n13838) );
  NAND U14289 ( .A(n13839), .B(n13838), .Z(n13840) );
  NANDN U14290 ( .A(n13841), .B(n13840), .Z(n13842) );
  AND U14291 ( .A(n13843), .B(n13842), .Z(n13845) );
  NANDN U14292 ( .A(n13845), .B(n13844), .Z(n13846) );
  NANDN U14293 ( .A(n13847), .B(n13846), .Z(n13848) );
  NAND U14294 ( .A(n13849), .B(n13848), .Z(n13851) );
  ANDN U14295 ( .B(n13851), .A(n13850), .Z(n13853) );
  NANDN U14296 ( .A(n13853), .B(n13852), .Z(n13854) );
  NAND U14297 ( .A(n13855), .B(n13854), .Z(n13856) );
  NAND U14298 ( .A(n13857), .B(n13856), .Z(n13858) );
  NAND U14299 ( .A(n13859), .B(n13858), .Z(n13860) );
  NANDN U14300 ( .A(n13861), .B(n13860), .Z(n13862) );
  NAND U14301 ( .A(n13863), .B(n13862), .Z(n13864) );
  NANDN U14302 ( .A(n13865), .B(n13864), .Z(n13866) );
  NANDN U14303 ( .A(n13867), .B(n13866), .Z(n13868) );
  AND U14304 ( .A(n13869), .B(n13868), .Z(n13870) );
  OR U14305 ( .A(n13871), .B(n13870), .Z(n13872) );
  NAND U14306 ( .A(n13873), .B(n13872), .Z(n13874) );
  NANDN U14307 ( .A(n13875), .B(n13874), .Z(n13876) );
  NAND U14308 ( .A(n13877), .B(n13876), .Z(n13878) );
  NANDN U14309 ( .A(n13879), .B(n13878), .Z(n13880) );
  AND U14310 ( .A(n13881), .B(n13880), .Z(n13883) );
  OR U14311 ( .A(n13883), .B(n13882), .Z(n13884) );
  AND U14312 ( .A(n13885), .B(n13884), .Z(n13886) );
  OR U14313 ( .A(n13887), .B(n13886), .Z(n13888) );
  NAND U14314 ( .A(n13889), .B(n13888), .Z(n13890) );
  NANDN U14315 ( .A(n13891), .B(n13890), .Z(n13892) );
  NAND U14316 ( .A(n13893), .B(n13892), .Z(n13894) );
  NANDN U14317 ( .A(n13895), .B(n13894), .Z(n13897) );
  ANDN U14318 ( .B(n13897), .A(n13896), .Z(n13899) );
  NANDN U14319 ( .A(n13899), .B(n13898), .Z(n13900) );
  AND U14320 ( .A(n13901), .B(n13900), .Z(n13902) );
  OR U14321 ( .A(n13903), .B(n13902), .Z(n13904) );
  AND U14322 ( .A(n13905), .B(n13904), .Z(n13907) );
  NANDN U14323 ( .A(n13907), .B(n13906), .Z(n13908) );
  AND U14324 ( .A(n13909), .B(n13908), .Z(n13911) );
  NANDN U14325 ( .A(n13911), .B(n13910), .Z(n13912) );
  NANDN U14326 ( .A(n13913), .B(n13912), .Z(n13914) );
  NAND U14327 ( .A(n13915), .B(n13914), .Z(n13916) );
  NAND U14328 ( .A(n13917), .B(n13916), .Z(n13918) );
  NAND U14329 ( .A(n13919), .B(n13918), .Z(n13921) );
  ANDN U14330 ( .B(n13921), .A(n13920), .Z(n13923) );
  NANDN U14331 ( .A(n13923), .B(n13922), .Z(n13924) );
  NAND U14332 ( .A(n13925), .B(n13924), .Z(n13926) );
  NAND U14333 ( .A(n13927), .B(n13926), .Z(n13928) );
  NANDN U14334 ( .A(n13929), .B(n13928), .Z(n13930) );
  AND U14335 ( .A(n13931), .B(n13930), .Z(n13933) );
  NANDN U14336 ( .A(n13933), .B(n13932), .Z(n13934) );
  NANDN U14337 ( .A(n13935), .B(n13934), .Z(n13936) );
  NAND U14338 ( .A(n13937), .B(n13936), .Z(n13938) );
  NANDN U14339 ( .A(n13939), .B(n13938), .Z(n13940) );
  NAND U14340 ( .A(n13941), .B(n13940), .Z(n13943) );
  ANDN U14341 ( .B(n13943), .A(n13942), .Z(n13945) );
  NANDN U14342 ( .A(n13945), .B(n13944), .Z(n13946) );
  NANDN U14343 ( .A(n13947), .B(n13946), .Z(n13948) );
  NANDN U14344 ( .A(n13949), .B(n13948), .Z(n13950) );
  NAND U14345 ( .A(n13951), .B(n13950), .Z(n13952) );
  NANDN U14346 ( .A(n13953), .B(n13952), .Z(n13954) );
  AND U14347 ( .A(n13955), .B(n13954), .Z(n13956) );
  OR U14348 ( .A(n13957), .B(n13956), .Z(n13958) );
  NAND U14349 ( .A(n13959), .B(n13958), .Z(n13960) );
  NAND U14350 ( .A(n13961), .B(n13960), .Z(n13962) );
  NANDN U14351 ( .A(n13963), .B(n13962), .Z(n13965) );
  ANDN U14352 ( .B(n13965), .A(n13964), .Z(n13967) );
  NANDN U14353 ( .A(n13967), .B(n13966), .Z(n13968) );
  NAND U14354 ( .A(n13969), .B(n13968), .Z(n13970) );
  NAND U14355 ( .A(n13971), .B(n13970), .Z(n13972) );
  NANDN U14356 ( .A(n13973), .B(n13972), .Z(n13974) );
  NANDN U14357 ( .A(n13975), .B(n13974), .Z(n13976) );
  AND U14358 ( .A(n13977), .B(n13976), .Z(n13978) );
  OR U14359 ( .A(n13979), .B(n13978), .Z(n13980) );
  NANDN U14360 ( .A(n13981), .B(n13980), .Z(n13982) );
  NAND U14361 ( .A(n13983), .B(n13982), .Z(n13984) );
  NANDN U14362 ( .A(n13985), .B(n13984), .Z(n13986) );
  NANDN U14363 ( .A(n13987), .B(n13986), .Z(n13988) );
  AND U14364 ( .A(n13989), .B(n13988), .Z(n13990) );
  OR U14365 ( .A(n13991), .B(n13990), .Z(n13992) );
  NAND U14366 ( .A(n13993), .B(n13992), .Z(n13994) );
  NANDN U14367 ( .A(n13995), .B(n13994), .Z(n13997) );
  NAND U14368 ( .A(n13997), .B(n13996), .Z(n13998) );
  NANDN U14369 ( .A(n13999), .B(n13998), .Z(n14000) );
  AND U14370 ( .A(n14001), .B(n14000), .Z(n14003) );
  NANDN U14371 ( .A(n14003), .B(n14002), .Z(n14004) );
  NANDN U14372 ( .A(n14005), .B(n14004), .Z(n14006) );
  NANDN U14373 ( .A(n14007), .B(n14006), .Z(n14008) );
  NAND U14374 ( .A(n14009), .B(n14008), .Z(n14010) );
  NANDN U14375 ( .A(n14011), .B(n14010), .Z(n14012) );
  AND U14376 ( .A(n14013), .B(n14012), .Z(n14015) );
  OR U14377 ( .A(n14015), .B(n14014), .Z(n14016) );
  NANDN U14378 ( .A(n14017), .B(n14016), .Z(n14018) );
  NAND U14379 ( .A(n14019), .B(n14018), .Z(n14020) );
  NAND U14380 ( .A(n14021), .B(n14020), .Z(n14022) );
  NAND U14381 ( .A(n14023), .B(n14022), .Z(n14025) );
  ANDN U14382 ( .B(n14025), .A(n14024), .Z(n14027) );
  NANDN U14383 ( .A(n14027), .B(n14026), .Z(n14028) );
  NAND U14384 ( .A(n14029), .B(n14028), .Z(n14030) );
  NAND U14385 ( .A(n14031), .B(n14030), .Z(n14032) );
  NANDN U14386 ( .A(n14033), .B(n14032), .Z(n14034) );
  AND U14387 ( .A(n14035), .B(n14034), .Z(n14037) );
  NANDN U14388 ( .A(n14037), .B(n14036), .Z(n14038) );
  NANDN U14389 ( .A(n14039), .B(n14038), .Z(n14040) );
  NAND U14390 ( .A(n14041), .B(n14040), .Z(n14042) );
  NANDN U14391 ( .A(n14043), .B(n14042), .Z(n14044) );
  AND U14392 ( .A(n14045), .B(n14044), .Z(n14047) );
  OR U14393 ( .A(n14047), .B(n14046), .Z(n14048) );
  AND U14394 ( .A(n14049), .B(n14048), .Z(n14050) );
  OR U14395 ( .A(n14051), .B(n14050), .Z(n14052) );
  AND U14396 ( .A(n14053), .B(n14052), .Z(n14054) );
  OR U14397 ( .A(n14055), .B(n14054), .Z(n14056) );
  NAND U14398 ( .A(n14057), .B(n14056), .Z(n14058) );
  NANDN U14399 ( .A(n14059), .B(n14058), .Z(n14060) );
  NAND U14400 ( .A(n14061), .B(n14060), .Z(n14063) );
  ANDN U14401 ( .B(n14063), .A(n14062), .Z(n14065) );
  NANDN U14402 ( .A(n14065), .B(n14064), .Z(n14066) );
  NAND U14403 ( .A(n14067), .B(n14066), .Z(n14068) );
  NAND U14404 ( .A(n14069), .B(n14068), .Z(n14071) );
  NANDN U14405 ( .A(n14071), .B(n14070), .Z(n14072) );
  NAND U14406 ( .A(n14073), .B(n14072), .Z(n14074) );
  OR U14407 ( .A(n14075), .B(n14074), .Z(n14076) );
  AND U14408 ( .A(n14077), .B(n14076), .Z(n14078) );
  OR U14409 ( .A(n14079), .B(n14078), .Z(n14080) );
  NANDN U14410 ( .A(n14081), .B(n14080), .Z(n14082) );
  NAND U14411 ( .A(n14083), .B(n14082), .Z(n14084) );
  NANDN U14412 ( .A(n14085), .B(n14084), .Z(n14086) );
  NAND U14413 ( .A(n14087), .B(n14086), .Z(n14088) );
  AND U14414 ( .A(n14089), .B(n14088), .Z(n14090) );
  OR U14415 ( .A(n14091), .B(n14090), .Z(n14092) );
  NAND U14416 ( .A(n14093), .B(n14092), .Z(n14094) );
  NANDN U14417 ( .A(n14095), .B(n14094), .Z(n14096) );
  NANDN U14418 ( .A(n14097), .B(n14096), .Z(n14098) );
  NAND U14419 ( .A(n14099), .B(n14098), .Z(n14100) );
  AND U14420 ( .A(n14101), .B(n14100), .Z(n14102) );
  OR U14421 ( .A(n14103), .B(n14102), .Z(n14104) );
  NAND U14422 ( .A(n14105), .B(n14104), .Z(n14106) );
  NANDN U14423 ( .A(n14107), .B(n14106), .Z(n14108) );
  AND U14424 ( .A(n14109), .B(n14108), .Z(n14110) );
  OR U14425 ( .A(n14111), .B(n14110), .Z(n14112) );
  NAND U14426 ( .A(n14113), .B(n14112), .Z(n14114) );
  NANDN U14427 ( .A(n14115), .B(n14114), .Z(n14117) );
  ANDN U14428 ( .B(n14117), .A(n14116), .Z(n14119) );
  NANDN U14429 ( .A(n14119), .B(n14118), .Z(n14120) );
  NANDN U14430 ( .A(n14121), .B(n14120), .Z(n14122) );
  NAND U14431 ( .A(n14123), .B(n14122), .Z(n14125) );
  ANDN U14432 ( .B(n14125), .A(n14124), .Z(n14126) );
  OR U14433 ( .A(n14127), .B(n14126), .Z(n14128) );
  NAND U14434 ( .A(n14129), .B(n14128), .Z(n14130) );
  NANDN U14435 ( .A(n14131), .B(n14130), .Z(n14132) );
  AND U14436 ( .A(n14133), .B(n14132), .Z(n14134) );
  OR U14437 ( .A(n14135), .B(n14134), .Z(n14136) );
  AND U14438 ( .A(n14137), .B(n14136), .Z(n14139) );
  NANDN U14439 ( .A(n14139), .B(n14138), .Z(n14140) );
  NAND U14440 ( .A(n14141), .B(n14140), .Z(n14142) );
  NAND U14441 ( .A(n14143), .B(n14142), .Z(n14145) );
  ANDN U14442 ( .B(n14145), .A(n14144), .Z(n14147) );
  NANDN U14443 ( .A(n14147), .B(n14146), .Z(n14148) );
  NANDN U14444 ( .A(n14149), .B(n14148), .Z(n14150) );
  AND U14445 ( .A(n14151), .B(n14150), .Z(n14153) );
  OR U14446 ( .A(n14153), .B(n14152), .Z(n14154) );
  AND U14447 ( .A(n14155), .B(n14154), .Z(n14157) );
  OR U14448 ( .A(n14157), .B(n14156), .Z(n14158) );
  AND U14449 ( .A(n14159), .B(n14158), .Z(n14160) );
  OR U14450 ( .A(n14161), .B(n14160), .Z(n14162) );
  NAND U14451 ( .A(n14163), .B(n14162), .Z(n14164) );
  NANDN U14452 ( .A(n14165), .B(n14164), .Z(n14166) );
  AND U14453 ( .A(n14167), .B(n14166), .Z(n14169) );
  NANDN U14454 ( .A(n14169), .B(n14168), .Z(n14170) );
  NAND U14455 ( .A(n14171), .B(n14170), .Z(n14173) );
  ANDN U14456 ( .B(n14173), .A(n14172), .Z(n14175) );
  NANDN U14457 ( .A(n14175), .B(n14174), .Z(n14176) );
  NAND U14458 ( .A(n14177), .B(n14176), .Z(n14178) );
  NAND U14459 ( .A(n14179), .B(n14178), .Z(n14180) );
  NANDN U14460 ( .A(n14181), .B(n14180), .Z(n14182) );
  AND U14461 ( .A(n14183), .B(n14182), .Z(n14185) );
  NANDN U14462 ( .A(n14185), .B(n14184), .Z(n14187) );
  ANDN U14463 ( .B(n14187), .A(n14186), .Z(n14189) );
  NANDN U14464 ( .A(n14189), .B(n14188), .Z(n14190) );
  AND U14465 ( .A(n14191), .B(n14190), .Z(n14193) );
  NANDN U14466 ( .A(n14193), .B(n14192), .Z(n14194) );
  NAND U14467 ( .A(n14195), .B(n14194), .Z(n14196) );
  NAND U14468 ( .A(n14197), .B(n14196), .Z(n14198) );
  NANDN U14469 ( .A(n14199), .B(n14198), .Z(n14200) );
  NAND U14470 ( .A(n14201), .B(n14200), .Z(n14202) );
  AND U14471 ( .A(n14203), .B(n14202), .Z(n14205) );
  NANDN U14472 ( .A(n14205), .B(n14204), .Z(n14206) );
  NANDN U14473 ( .A(n14207), .B(n14206), .Z(n14208) );
  NANDN U14474 ( .A(n14209), .B(n14208), .Z(n14210) );
  NAND U14475 ( .A(n14211), .B(n14210), .Z(n14213) );
  ANDN U14476 ( .B(n14213), .A(n14212), .Z(n14215) );
  NANDN U14477 ( .A(n14215), .B(n14214), .Z(n14217) );
  ANDN U14478 ( .B(n14217), .A(n14216), .Z(n14219) );
  NANDN U14479 ( .A(n14219), .B(n14218), .Z(n14220) );
  AND U14480 ( .A(n14221), .B(n14220), .Z(n14223) );
  NANDN U14481 ( .A(n14223), .B(n14222), .Z(n14224) );
  AND U14482 ( .A(n14225), .B(n14224), .Z(n14227) );
  OR U14483 ( .A(n14227), .B(n14226), .Z(n14228) );
  AND U14484 ( .A(n14229), .B(n14228), .Z(n14231) );
  OR U14485 ( .A(n14231), .B(n14230), .Z(n14232) );
  AND U14486 ( .A(n14233), .B(n14232), .Z(n14235) );
  OR U14487 ( .A(n14235), .B(n14234), .Z(n14237) );
  ANDN U14488 ( .B(n14237), .A(n14236), .Z(n14238) );
  OR U14489 ( .A(n14239), .B(n14238), .Z(n14240) );
  NAND U14490 ( .A(n14241), .B(n14240), .Z(n14242) );
  NANDN U14491 ( .A(n14243), .B(n14242), .Z(n14244) );
  AND U14492 ( .A(n14245), .B(n14244), .Z(n14247) );
  NANDN U14493 ( .A(n14247), .B(n14246), .Z(n14248) );
  NAND U14494 ( .A(n14249), .B(n14248), .Z(n14251) );
  ANDN U14495 ( .B(n14251), .A(n14250), .Z(n14253) );
  NANDN U14496 ( .A(n14253), .B(n14252), .Z(n14254) );
  NAND U14497 ( .A(n14255), .B(n14254), .Z(n14256) );
  NAND U14498 ( .A(n14257), .B(n14256), .Z(n14258) );
  NANDN U14499 ( .A(n14259), .B(n14258), .Z(n14261) );
  ANDN U14500 ( .B(n14261), .A(n14260), .Z(n14263) );
  NANDN U14501 ( .A(n14263), .B(n14262), .Z(n14264) );
  NAND U14502 ( .A(n14265), .B(n14264), .Z(n14266) );
  NAND U14503 ( .A(n14267), .B(n14266), .Z(n14268) );
  NANDN U14504 ( .A(n14269), .B(n14268), .Z(n14270) );
  NAND U14505 ( .A(n14271), .B(n14270), .Z(n14273) );
  ANDN U14506 ( .B(n14273), .A(n14272), .Z(n14277) );
  NAND U14507 ( .A(n14275), .B(n14274), .Z(n14276) );
  AND U14508 ( .A(n14277), .B(n14276), .Z(n14279) );
  NANDN U14509 ( .A(n14279), .B(n14278), .Z(n14280) );
  NAND U14510 ( .A(n14281), .B(n14280), .Z(n14282) );
  NAND U14511 ( .A(n14283), .B(n14282), .Z(n14284) );
  NANDN U14512 ( .A(n14285), .B(n14284), .Z(n14286) );
  AND U14513 ( .A(n14287), .B(n14286), .Z(n14289) );
  NANDN U14514 ( .A(n14289), .B(n14288), .Z(n14291) );
  ANDN U14515 ( .B(n14291), .A(n14290), .Z(n14293) );
  NANDN U14516 ( .A(n14293), .B(n14292), .Z(n14294) );
  AND U14517 ( .A(n14295), .B(n14294), .Z(n14297) );
  NANDN U14518 ( .A(n14297), .B(n14296), .Z(n14298) );
  NAND U14519 ( .A(n14299), .B(n14298), .Z(n14300) );
  NAND U14520 ( .A(n14301), .B(n14300), .Z(n14303) );
  ANDN U14521 ( .B(n14303), .A(n14302), .Z(n14305) );
  NANDN U14522 ( .A(n14305), .B(n14304), .Z(n14306) );
  NAND U14523 ( .A(n14307), .B(n14306), .Z(n14308) );
  NAND U14524 ( .A(n14309), .B(n14308), .Z(n14310) );
  NANDN U14525 ( .A(n14311), .B(n14310), .Z(n14312) );
  AND U14526 ( .A(n14313), .B(n14312), .Z(n14314) );
  OR U14527 ( .A(n14315), .B(n14314), .Z(n14316) );
  NANDN U14528 ( .A(n14317), .B(n14316), .Z(n14318) );
  NAND U14529 ( .A(n14319), .B(n14318), .Z(n14320) );
  NANDN U14530 ( .A(n14321), .B(n14320), .Z(n14322) );
  NAND U14531 ( .A(n14323), .B(n14322), .Z(n14324) );
  NANDN U14532 ( .A(n14325), .B(n14324), .Z(n14326) );
  AND U14533 ( .A(n14327), .B(n14326), .Z(n14328) );
  OR U14534 ( .A(n14329), .B(n14328), .Z(n14330) );
  NAND U14535 ( .A(n14331), .B(n14330), .Z(n14332) );
  AND U14536 ( .A(n14333), .B(n14332), .Z(n14335) );
  OR U14537 ( .A(n14335), .B(n14334), .Z(n14337) );
  ANDN U14538 ( .B(n14337), .A(n14336), .Z(n14338) );
  AND U14539 ( .A(n14339), .B(n14338), .Z(n14345) );
  NAND U14540 ( .A(n14341), .B(n14340), .Z(n14343) );
  ANDN U14541 ( .B(n14343), .A(n14342), .Z(n14344) );
  NANDN U14542 ( .A(n14345), .B(n14344), .Z(n14346) );
  NANDN U14543 ( .A(n14347), .B(n14346), .Z(n14348) );
  NAND U14544 ( .A(n14349), .B(n14348), .Z(n14350) );
  NANDN U14545 ( .A(n14351), .B(n14350), .Z(n14352) );
  NAND U14546 ( .A(n14353), .B(n14352), .Z(n14354) );
  NAND U14547 ( .A(n14355), .B(n14354), .Z(n14357) );
  ANDN U14548 ( .B(n14357), .A(n14356), .Z(n14359) );
  NANDN U14549 ( .A(n14359), .B(n14358), .Z(n14360) );
  NAND U14550 ( .A(n14361), .B(n14360), .Z(n14362) );
  NANDN U14551 ( .A(n14363), .B(n14362), .Z(n14364) );
  NAND U14552 ( .A(n14365), .B(n14364), .Z(n14367) );
  ANDN U14553 ( .B(n14367), .A(n14366), .Z(n14369) );
  NANDN U14554 ( .A(n14369), .B(n14368), .Z(n14370) );
  NAND U14555 ( .A(n14371), .B(n14370), .Z(n14372) );
  NAND U14556 ( .A(n14373), .B(n14372), .Z(n14374) );
  NANDN U14557 ( .A(n14375), .B(n14374), .Z(n14376) );
  NAND U14558 ( .A(n14377), .B(n14376), .Z(n14379) );
  ANDN U14559 ( .B(n14379), .A(n14378), .Z(n14383) );
  NANDN U14560 ( .A(n14381), .B(n14380), .Z(n14382) );
  AND U14561 ( .A(n14383), .B(n14382), .Z(n14385) );
  NANDN U14562 ( .A(n14385), .B(n14384), .Z(n14386) );
  NAND U14563 ( .A(n14387), .B(n14386), .Z(n14388) );
  NAND U14564 ( .A(n14389), .B(n14388), .Z(n14390) );
  NANDN U14565 ( .A(n14391), .B(n14390), .Z(n14392) );
  AND U14566 ( .A(n14393), .B(n14392), .Z(n14395) );
  NANDN U14567 ( .A(n14395), .B(n14394), .Z(n14397) );
  ANDN U14568 ( .B(n14397), .A(n14396), .Z(n14399) );
  NANDN U14569 ( .A(n14399), .B(n14398), .Z(n14401) );
  ANDN U14570 ( .B(n14401), .A(n14400), .Z(n14403) );
  NANDN U14571 ( .A(n14403), .B(n14402), .Z(n14404) );
  NANDN U14572 ( .A(n14405), .B(n14404), .Z(n14406) );
  NAND U14573 ( .A(n14407), .B(n14406), .Z(n14408) );
  NANDN U14574 ( .A(n14409), .B(n14408), .Z(n14410) );
  NANDN U14575 ( .A(n14411), .B(n14410), .Z(n14412) );
  AND U14576 ( .A(n14413), .B(n14412), .Z(n14414) );
  OR U14577 ( .A(n14415), .B(n14414), .Z(n14416) );
  NAND U14578 ( .A(n14417), .B(n14416), .Z(n14418) );
  NANDN U14579 ( .A(n14419), .B(n14418), .Z(n14420) );
  NAND U14580 ( .A(n14421), .B(n14420), .Z(n14422) );
  AND U14581 ( .A(n14423), .B(n14422), .Z(n14424) );
  OR U14582 ( .A(n14425), .B(n14424), .Z(n14426) );
  AND U14583 ( .A(n14427), .B(n14426), .Z(n14429) );
  OR U14584 ( .A(n14429), .B(n14428), .Z(n14430) );
  AND U14585 ( .A(n14431), .B(n14430), .Z(n14432) );
  OR U14586 ( .A(n14433), .B(n14432), .Z(n14434) );
  AND U14587 ( .A(n14435), .B(n14434), .Z(n14437) );
  OR U14588 ( .A(n14437), .B(n14436), .Z(n14438) );
  AND U14589 ( .A(n14439), .B(n14438), .Z(n14440) );
  OR U14590 ( .A(n14441), .B(n14440), .Z(n14442) );
  NAND U14591 ( .A(n14443), .B(n14442), .Z(n14444) );
  NAND U14592 ( .A(n14445), .B(n14444), .Z(n14446) );
  NANDN U14593 ( .A(n14447), .B(n14446), .Z(n14448) );
  NAND U14594 ( .A(n14449), .B(n14448), .Z(n14450) );
  AND U14595 ( .A(n14451), .B(n14450), .Z(n14452) );
  OR U14596 ( .A(n14453), .B(n14452), .Z(n14454) );
  NAND U14597 ( .A(n14455), .B(n14454), .Z(n14456) );
  NANDN U14598 ( .A(n14457), .B(n14456), .Z(n14458) );
  NANDN U14599 ( .A(n14459), .B(n14458), .Z(n14460) );
  NAND U14600 ( .A(n14461), .B(n14460), .Z(n14463) );
  ANDN U14601 ( .B(n14463), .A(n14462), .Z(n14465) );
  NANDN U14602 ( .A(n14465), .B(n14464), .Z(n14466) );
  NANDN U14603 ( .A(n14467), .B(n14466), .Z(n14468) );
  NAND U14604 ( .A(n14469), .B(n14468), .Z(n14470) );
  NANDN U14605 ( .A(n14471), .B(n14470), .Z(n14472) );
  AND U14606 ( .A(n14473), .B(n14472), .Z(n14475) );
  NANDN U14607 ( .A(n14475), .B(n14474), .Z(n14477) );
  ANDN U14608 ( .B(n14477), .A(n14476), .Z(n14479) );
  NANDN U14609 ( .A(n14479), .B(n14478), .Z(n14480) );
  AND U14610 ( .A(n14481), .B(n14480), .Z(n14483) );
  OR U14611 ( .A(n14483), .B(n14482), .Z(n14485) );
  ANDN U14612 ( .B(n14485), .A(n14484), .Z(n14487) );
  NANDN U14613 ( .A(n14487), .B(n14486), .Z(n14489) );
  ANDN U14614 ( .B(n14489), .A(n14488), .Z(n14491) );
  NANDN U14615 ( .A(n14491), .B(n14490), .Z(n14492) );
  NANDN U14616 ( .A(n14493), .B(n14492), .Z(n14494) );
  NANDN U14617 ( .A(n14495), .B(n14494), .Z(n14496) );
  NAND U14618 ( .A(n14497), .B(n14496), .Z(n14498) );
  AND U14619 ( .A(n14499), .B(n14498), .Z(n14501) );
  NANDN U14620 ( .A(n14501), .B(n14500), .Z(n14502) );
  AND U14621 ( .A(n14503), .B(n14502), .Z(n14505) );
  NANDN U14622 ( .A(n14505), .B(n14504), .Z(n14506) );
  NAND U14623 ( .A(n14507), .B(n14506), .Z(n14508) );
  NAND U14624 ( .A(n14509), .B(n14508), .Z(n14513) );
  NANDN U14625 ( .A(n14511), .B(n14510), .Z(n14512) );
  NANDN U14626 ( .A(n14513), .B(n14512), .Z(n14514) );
  AND U14627 ( .A(n14515), .B(n14514), .Z(n14517) );
  NANDN U14628 ( .A(n14517), .B(n14516), .Z(n14519) );
  ANDN U14629 ( .B(n14519), .A(n14518), .Z(n14521) );
  NANDN U14630 ( .A(n14521), .B(n14520), .Z(n14522) );
  AND U14631 ( .A(n14523), .B(n14522), .Z(n14525) );
  OR U14632 ( .A(n14525), .B(n14524), .Z(n14526) );
  AND U14633 ( .A(n14527), .B(n14526), .Z(n14529) );
  NANDN U14634 ( .A(n14529), .B(n14528), .Z(n14530) );
  NAND U14635 ( .A(n14531), .B(n14530), .Z(n14533) );
  NAND U14636 ( .A(n14533), .B(n14532), .Z(n14534) );
  NANDN U14637 ( .A(n14535), .B(n14534), .Z(n14536) );
  AND U14638 ( .A(n14537), .B(n14536), .Z(n14539) );
  OR U14639 ( .A(n14539), .B(n14538), .Z(n14540) );
  NAND U14640 ( .A(n14541), .B(n14540), .Z(n14542) );
  NAND U14641 ( .A(n14543), .B(n14542), .Z(n14545) );
  ANDN U14642 ( .B(n14545), .A(n14544), .Z(n14547) );
  NANDN U14643 ( .A(n14547), .B(n14546), .Z(n14548) );
  NAND U14644 ( .A(n14549), .B(n14548), .Z(n14551) );
  ANDN U14645 ( .B(n14551), .A(n14550), .Z(n14553) );
  NANDN U14646 ( .A(n14553), .B(n14552), .Z(n14554) );
  NANDN U14647 ( .A(n14555), .B(n14554), .Z(n14556) );
  NAND U14648 ( .A(n14557), .B(n14556), .Z(n14558) );
  NANDN U14649 ( .A(n14559), .B(n14558), .Z(n14560) );
  NAND U14650 ( .A(n14561), .B(n14560), .Z(n14562) );
  NANDN U14651 ( .A(n14563), .B(n14562), .Z(n14564) );
  AND U14652 ( .A(n14565), .B(n14564), .Z(n14567) );
  NANDN U14653 ( .A(n14567), .B(n14566), .Z(n14568) );
  NAND U14654 ( .A(n14569), .B(n14568), .Z(n14570) );
  AND U14655 ( .A(n14571), .B(n14570), .Z(n14573) );
  NANDN U14656 ( .A(n14573), .B(n14572), .Z(n14575) );
  ANDN U14657 ( .B(n14575), .A(n14574), .Z(n14577) );
  NANDN U14658 ( .A(n14577), .B(n14576), .Z(n14579) );
  ANDN U14659 ( .B(n14579), .A(n14578), .Z(n14581) );
  NANDN U14660 ( .A(n14581), .B(n14580), .Z(n14582) );
  AND U14661 ( .A(n14583), .B(n14582), .Z(n14585) );
  NANDN U14662 ( .A(n14585), .B(n14584), .Z(n14587) );
  ANDN U14663 ( .B(n14587), .A(n14586), .Z(n14589) );
  OR U14664 ( .A(n14589), .B(n14588), .Z(n14590) );
  AND U14665 ( .A(n14591), .B(n14590), .Z(n14593) );
  OR U14666 ( .A(n14593), .B(n14592), .Z(n14594) );
  AND U14667 ( .A(n14595), .B(n14594), .Z(n14597) );
  NANDN U14668 ( .A(n14597), .B(n14596), .Z(n14598) );
  AND U14669 ( .A(n14599), .B(n14598), .Z(n14603) );
  AND U14670 ( .A(n14601), .B(n14600), .Z(n14602) );
  NANDN U14671 ( .A(n14603), .B(n14602), .Z(n14605) );
  ANDN U14672 ( .B(n14605), .A(n14604), .Z(n14607) );
  NANDN U14673 ( .A(n14607), .B(n14606), .Z(n14609) );
  ANDN U14674 ( .B(n14609), .A(n14608), .Z(n14611) );
  NANDN U14675 ( .A(n14611), .B(n14610), .Z(n14612) );
  NAND U14676 ( .A(n14613), .B(n14612), .Z(n14614) );
  NAND U14677 ( .A(n14615), .B(n14614), .Z(n14616) );
  NAND U14678 ( .A(n14617), .B(n14616), .Z(n14618) );
  NAND U14679 ( .A(n14619), .B(n14618), .Z(n14620) );
  AND U14680 ( .A(n14621), .B(n14620), .Z(n14623) );
  NANDN U14681 ( .A(n14623), .B(n14622), .Z(n14624) );
  NAND U14682 ( .A(n14625), .B(n14624), .Z(n14626) );
  NAND U14683 ( .A(n14627), .B(n14626), .Z(n14628) );
  AND U14684 ( .A(n14629), .B(n14628), .Z(n14631) );
  NANDN U14685 ( .A(n14631), .B(n14630), .Z(n14633) );
  ANDN U14686 ( .B(n14633), .A(n14632), .Z(n14635) );
  NANDN U14687 ( .A(n14635), .B(n14634), .Z(n14636) );
  NANDN U14688 ( .A(n14637), .B(n14636), .Z(n14638) );
  NAND U14689 ( .A(n14639), .B(n14638), .Z(n14640) );
  NANDN U14690 ( .A(n14641), .B(n14640), .Z(n14642) );
  NANDN U14691 ( .A(n14643), .B(n14642), .Z(n14644) );
  NAND U14692 ( .A(n14645), .B(n14644), .Z(n14649) );
  NANDN U14693 ( .A(n14647), .B(n14646), .Z(n14648) );
  AND U14694 ( .A(n14649), .B(n14648), .Z(n14650) );
  NANDN U14695 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U14696 ( .A(n14653), .B(n14652), .Z(n14655) );
  NANDN U14697 ( .A(n14655), .B(n14654), .Z(n14656) );
  NAND U14698 ( .A(n14657), .B(n14656), .Z(n14658) );
  NAND U14699 ( .A(n14659), .B(n14658), .Z(n14660) );
  AND U14700 ( .A(n14661), .B(n14660), .Z(n14663) );
  NANDN U14701 ( .A(n14663), .B(n14662), .Z(n14664) );
  NANDN U14702 ( .A(n14665), .B(n14664), .Z(n14666) );
  NAND U14703 ( .A(n14667), .B(n14666), .Z(n14669) );
  ANDN U14704 ( .B(n14669), .A(n14668), .Z(n14671) );
  NANDN U14705 ( .A(n14671), .B(n14670), .Z(n14672) );
  NAND U14706 ( .A(n14673), .B(n14672), .Z(n14674) );
  NAND U14707 ( .A(n14675), .B(n14674), .Z(n14677) );
  ANDN U14708 ( .B(n14677), .A(n14676), .Z(n14679) );
  NANDN U14709 ( .A(n14679), .B(n14678), .Z(n14680) );
  NANDN U14710 ( .A(n14681), .B(n14680), .Z(n14682) );
  AND U14711 ( .A(n14683), .B(n14682), .Z(n14684) );
endmodule

