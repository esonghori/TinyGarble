
module alu ( x, y, c, o );
  input [3:0] x;
  input [3:0] y;
  input [2:0] c;
  output [7:0] o;
  wire   n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382;

  IV U123 ( .A(c[2]), .Z(n123) );
  NOR U124 ( .A(c[0]), .B(c[1]), .Z(n121) );
  IV U125 ( .A(n121), .Z(n122) );
  NOR U126 ( .A(n123), .B(n122), .Z(n124) );
  IV U127 ( .A(n124), .Z(n367) );
  IV U128 ( .A(x[0]), .Z(n224) );
  IV U129 ( .A(y[0]), .Z(n249) );
  NOR U130 ( .A(n224), .B(n249), .Z(n146) );
  IV U131 ( .A(n146), .Z(n172) );
  NOR U132 ( .A(n367), .B(n172), .Z(n128) );
  NOR U133 ( .A(c[1]), .B(y[0]), .Z(n125) );
  XOR U134 ( .A(x[0]), .B(n125), .Z(n126) );
  NOR U135 ( .A(c[2]), .B(n126), .Z(n127) );
  NOR U136 ( .A(n128), .B(n127), .Z(n129) );
  IV U137 ( .A(n129), .Z(o[0]) );
  IV U138 ( .A(c[1]), .Z(n195) );
  IV U139 ( .A(c[0]), .Z(n193) );
  XOR U140 ( .A(x[1]), .B(n193), .Z(n130) );
  NOR U141 ( .A(n195), .B(n130), .Z(n131) );
  IV U142 ( .A(n131), .Z(n132) );
  NOR U143 ( .A(c[2]), .B(n132), .Z(n206) );
  IV U144 ( .A(n206), .Z(n133) );
  NOR U145 ( .A(n224), .B(n133), .Z(n164) );
  NOR U146 ( .A(c[2]), .B(n193), .Z(n134) );
  IV U147 ( .A(n134), .Z(n148) );
  NOR U148 ( .A(n195), .B(n148), .Z(n135) );
  IV U149 ( .A(n135), .Z(n338) );
  NOR U150 ( .A(x[0]), .B(n338), .Z(n136) );
  IV U151 ( .A(n136), .Z(n137) );
  IV U152 ( .A(x[1]), .Z(n235) );
  NOR U153 ( .A(n137), .B(n235), .Z(n161) );
  NOR U154 ( .A(n235), .B(n249), .Z(n250) );
  IV U155 ( .A(y[1]), .Z(n228) );
  NOR U156 ( .A(n224), .B(n228), .Z(n138) );
  IV U157 ( .A(n138), .Z(n251) );
  XOR U158 ( .A(n250), .B(n251), .Z(n139) );
  NOR U159 ( .A(n367), .B(n139), .Z(n158) );
  NOR U160 ( .A(c[2]), .B(c[0]), .Z(n140) );
  IV U161 ( .A(n140), .Z(n144) );
  NOR U162 ( .A(n144), .B(n195), .Z(n141) );
  IV U163 ( .A(n141), .Z(n350) );
  NOR U164 ( .A(x[0]), .B(n350), .Z(n142) );
  IV U165 ( .A(n142), .Z(n143) );
  NOR U166 ( .A(n143), .B(x[1]), .Z(n155) );
  NOR U167 ( .A(c[1]), .B(n144), .Z(n145) );
  IV U168 ( .A(n145), .Z(n372) );
  XOR U169 ( .A(n235), .B(y[1]), .Z(n173) );
  XOR U170 ( .A(n173), .B(n146), .Z(n147) );
  NOR U171 ( .A(n372), .B(n147), .Z(n152) );
  NOR U172 ( .A(c[1]), .B(n148), .Z(n149) );
  IV U173 ( .A(n149), .Z(n324) );
  NOR U174 ( .A(x[0]), .B(n249), .Z(n168) );
  XOR U175 ( .A(n168), .B(n173), .Z(n150) );
  NOR U176 ( .A(n324), .B(n150), .Z(n151) );
  NOR U177 ( .A(n152), .B(n151), .Z(n153) );
  IV U178 ( .A(n153), .Z(n154) );
  NOR U179 ( .A(n155), .B(n154), .Z(n156) );
  IV U180 ( .A(n156), .Z(n157) );
  NOR U181 ( .A(n158), .B(n157), .Z(n159) );
  IV U182 ( .A(n159), .Z(n160) );
  NOR U183 ( .A(n161), .B(n160), .Z(n162) );
  IV U184 ( .A(n162), .Z(n163) );
  NOR U185 ( .A(n164), .B(n163), .Z(n165) );
  IV U186 ( .A(n165), .Z(o[1]) );
  NOR U187 ( .A(n235), .B(n224), .Z(n166) );
  IV U188 ( .A(n166), .Z(n314) );
  NOR U189 ( .A(n314), .B(n338), .Z(n184) );
  NOR U190 ( .A(y[1]), .B(n235), .Z(n170) );
  NOR U191 ( .A(x[1]), .B(n228), .Z(n167) );
  NOR U192 ( .A(n168), .B(n167), .Z(n169) );
  NOR U193 ( .A(n170), .B(n169), .Z(n291) );
  IV U194 ( .A(n291), .Z(n171) );
  NOR U195 ( .A(n324), .B(n171), .Z(n176) );
  NOR U196 ( .A(n235), .B(n228), .Z(n217) );
  NOR U197 ( .A(n173), .B(n172), .Z(n174) );
  NOR U198 ( .A(n217), .B(n174), .Z(n177) );
  NOR U199 ( .A(n372), .B(n177), .Z(n175) );
  NOR U200 ( .A(n176), .B(n175), .Z(n199) );
  NOR U201 ( .A(n199), .B(y[2]), .Z(n181) );
  IV U202 ( .A(n177), .Z(n318) );
  NOR U203 ( .A(n372), .B(n318), .Z(n179) );
  NOR U204 ( .A(n291), .B(n324), .Z(n178) );
  NOR U205 ( .A(n179), .B(n178), .Z(n198) );
  IV U206 ( .A(y[2]), .Z(n289) );
  NOR U207 ( .A(n198), .B(n289), .Z(n180) );
  NOR U208 ( .A(n181), .B(n180), .Z(n182) );
  IV U209 ( .A(n182), .Z(n183) );
  NOR U210 ( .A(n184), .B(n183), .Z(n185) );
  NOR U211 ( .A(x[2]), .B(n185), .Z(n215) );
  NOR U212 ( .A(x[2]), .B(x[0]), .Z(n186) );
  IV U213 ( .A(n186), .Z(n187) );
  NOR U214 ( .A(x[1]), .B(n187), .Z(n188) );
  IV U215 ( .A(n188), .Z(n348) );
  NOR U216 ( .A(n348), .B(n350), .Z(n287) );
  IV U217 ( .A(x[2]), .Z(n315) );
  NOR U218 ( .A(n251), .B(n235), .Z(n189) );
  XOR U219 ( .A(n315), .B(n189), .Z(n190) );
  NOR U220 ( .A(n249), .B(n190), .Z(n255) );
  NOR U221 ( .A(n224), .B(n289), .Z(n191) );
  IV U222 ( .A(n191), .Z(n218) );
  XOR U223 ( .A(n218), .B(n217), .Z(n256) );
  XOR U224 ( .A(n255), .B(n256), .Z(n192) );
  NOR U225 ( .A(n367), .B(n192), .Z(n210) );
  XOR U226 ( .A(x[0]), .B(n193), .Z(n194) );
  NOR U227 ( .A(n195), .B(n194), .Z(n196) );
  IV U228 ( .A(n196), .Z(n197) );
  NOR U229 ( .A(c[2]), .B(n197), .Z(n204) );
  NOR U230 ( .A(n198), .B(y[2]), .Z(n201) );
  NOR U231 ( .A(n199), .B(n289), .Z(n200) );
  NOR U232 ( .A(n201), .B(n200), .Z(n202) );
  IV U233 ( .A(n202), .Z(n203) );
  NOR U234 ( .A(n204), .B(n203), .Z(n205) );
  IV U235 ( .A(n205), .Z(n207) );
  NOR U236 ( .A(n207), .B(n206), .Z(n208) );
  NOR U237 ( .A(n315), .B(n208), .Z(n209) );
  NOR U238 ( .A(n210), .B(n209), .Z(n211) );
  IV U239 ( .A(n211), .Z(n212) );
  NOR U240 ( .A(n287), .B(n212), .Z(n213) );
  IV U241 ( .A(n213), .Z(n214) );
  NOR U242 ( .A(n215), .B(n214), .Z(n216) );
  IV U243 ( .A(n216), .Z(o[2]) );
  NOR U244 ( .A(n315), .B(n228), .Z(n223) );
  IV U245 ( .A(n223), .Z(n221) );
  IV U246 ( .A(n217), .Z(n219) );
  NOR U247 ( .A(n219), .B(n218), .Z(n220) );
  IV U248 ( .A(n220), .Z(n222) );
  NOR U249 ( .A(n221), .B(n222), .Z(n227) );
  XOR U250 ( .A(n223), .B(n222), .Z(n261) );
  IV U251 ( .A(y[3]), .Z(n373) );
  NOR U252 ( .A(n224), .B(n373), .Z(n232) );
  NOR U253 ( .A(n235), .B(n289), .Z(n225) );
  IV U254 ( .A(n225), .Z(n233) );
  XOR U255 ( .A(n232), .B(n233), .Z(n260) );
  NOR U256 ( .A(n261), .B(n260), .Z(n226) );
  NOR U257 ( .A(n227), .B(n226), .Z(n229) );
  IV U258 ( .A(x[3]), .Z(n362) );
  NOR U259 ( .A(n229), .B(n362), .Z(n246) );
  NOR U260 ( .A(n362), .B(n228), .Z(n231) );
  IV U261 ( .A(n229), .Z(n230) );
  NOR U262 ( .A(n231), .B(n230), .Z(n245) );
  NOR U263 ( .A(n315), .B(n289), .Z(n317) );
  IV U264 ( .A(n232), .Z(n234) );
  NOR U265 ( .A(n234), .B(n233), .Z(n240) );
  NOR U266 ( .A(n235), .B(n373), .Z(n241) );
  XOR U267 ( .A(n240), .B(n241), .Z(n236) );
  XOR U268 ( .A(n317), .B(n236), .Z(n237) );
  IV U269 ( .A(n237), .Z(n247) );
  NOR U270 ( .A(n245), .B(n247), .Z(n238) );
  NOR U271 ( .A(n246), .B(n238), .Z(n269) );
  NOR U272 ( .A(n362), .B(n289), .Z(n276) );
  IV U273 ( .A(n276), .Z(n274) );
  NOR U274 ( .A(n315), .B(n373), .Z(n239) );
  IV U275 ( .A(n239), .Z(n278) );
  NOR U276 ( .A(n240), .B(n317), .Z(n243) );
  IV U277 ( .A(n241), .Z(n242) );
  NOR U278 ( .A(n243), .B(n242), .Z(n277) );
  IV U279 ( .A(n277), .Z(n275) );
  XOR U280 ( .A(n278), .B(n275), .Z(n244) );
  XOR U281 ( .A(n274), .B(n244), .Z(n268) );
  NOR U282 ( .A(n269), .B(n268), .Z(n273) );
  NOR U283 ( .A(n246), .B(n245), .Z(n248) );
  XOR U284 ( .A(n248), .B(n247), .Z(n365) );
  NOR U285 ( .A(n362), .B(n249), .Z(n262) );
  IV U286 ( .A(n250), .Z(n252) );
  NOR U287 ( .A(n252), .B(n251), .Z(n253) );
  IV U288 ( .A(n253), .Z(n254) );
  NOR U289 ( .A(n315), .B(n254), .Z(n259) );
  IV U290 ( .A(n255), .Z(n257) );
  NOR U291 ( .A(n257), .B(n256), .Z(n258) );
  NOR U292 ( .A(n259), .B(n258), .Z(n263) );
  IV U293 ( .A(n263), .Z(n333) );
  NOR U294 ( .A(n262), .B(n333), .Z(n266) );
  XOR U295 ( .A(n261), .B(n260), .Z(n336) );
  IV U296 ( .A(n262), .Z(n334) );
  NOR U297 ( .A(n263), .B(n334), .Z(n264) );
  NOR U298 ( .A(n336), .B(n264), .Z(n265) );
  NOR U299 ( .A(n266), .B(n265), .Z(n364) );
  IV U300 ( .A(n364), .Z(n267) );
  NOR U301 ( .A(n365), .B(n267), .Z(n309) );
  IV U302 ( .A(n309), .Z(n271) );
  XOR U303 ( .A(n269), .B(n268), .Z(n270) );
  IV U304 ( .A(n270), .Z(n310) );
  NOR U305 ( .A(n271), .B(n310), .Z(n272) );
  NOR U306 ( .A(n273), .B(n272), .Z(n303) );
  NOR U307 ( .A(n275), .B(n274), .Z(n281) );
  NOR U308 ( .A(n277), .B(n276), .Z(n279) );
  NOR U309 ( .A(n279), .B(n278), .Z(n280) );
  NOR U310 ( .A(n281), .B(n280), .Z(n283) );
  NOR U311 ( .A(n373), .B(n362), .Z(n282) );
  XOR U312 ( .A(n283), .B(n282), .Z(n304) );
  NOR U313 ( .A(n303), .B(n304), .Z(n285) );
  NOR U314 ( .A(n283), .B(n362), .Z(n284) );
  NOR U315 ( .A(n285), .B(n284), .Z(n286) );
  NOR U316 ( .A(n286), .B(n367), .Z(n301) );
  IV U317 ( .A(n287), .Z(n288) );
  NOR U318 ( .A(x[3]), .B(n288), .Z(n299) );
  NOR U319 ( .A(y[2]), .B(n315), .Z(n293) );
  NOR U320 ( .A(x[2]), .B(n289), .Z(n290) );
  NOR U321 ( .A(n291), .B(n290), .Z(n292) );
  NOR U322 ( .A(n293), .B(n292), .Z(n325) );
  IV U323 ( .A(n325), .Z(n322) );
  NOR U324 ( .A(y[3]), .B(n362), .Z(n294) );
  NOR U325 ( .A(n322), .B(n294), .Z(n296) );
  NOR U326 ( .A(x[3]), .B(n373), .Z(n295) );
  NOR U327 ( .A(n296), .B(n295), .Z(n297) );
  NOR U328 ( .A(n324), .B(n297), .Z(n298) );
  NOR U329 ( .A(n299), .B(n298), .Z(n300) );
  IV U330 ( .A(n300), .Z(n377) );
  NOR U331 ( .A(n301), .B(n377), .Z(n302) );
  IV U332 ( .A(n302), .Z(o[7]) );
  XOR U333 ( .A(n304), .B(n303), .Z(n305) );
  IV U334 ( .A(n305), .Z(n306) );
  NOR U335 ( .A(n367), .B(n306), .Z(n307) );
  NOR U336 ( .A(n307), .B(n377), .Z(n308) );
  IV U337 ( .A(n308), .Z(o[6]) );
  XOR U338 ( .A(n310), .B(n309), .Z(n311) );
  NOR U339 ( .A(n367), .B(n311), .Z(n312) );
  NOR U340 ( .A(n312), .B(n377), .Z(n313) );
  IV U341 ( .A(n313), .Z(o[5]) );
  NOR U342 ( .A(n315), .B(n314), .Z(n339) );
  IV U343 ( .A(n339), .Z(n316) );
  NOR U344 ( .A(n316), .B(n338), .Z(n360) );
  NOR U345 ( .A(x[2]), .B(y[2]), .Z(n320) );
  NOR U346 ( .A(n318), .B(n317), .Z(n319) );
  NOR U347 ( .A(n320), .B(n319), .Z(n371) );
  IV U348 ( .A(n371), .Z(n321) );
  NOR U349 ( .A(n372), .B(n321), .Z(n361) );
  NOR U350 ( .A(n322), .B(n324), .Z(n323) );
  NOR U351 ( .A(n361), .B(n323), .Z(n341) );
  NOR U352 ( .A(n341), .B(y[3]), .Z(n329) );
  NOR U353 ( .A(n372), .B(n371), .Z(n327) );
  NOR U354 ( .A(n325), .B(n324), .Z(n326) );
  NOR U355 ( .A(n327), .B(n326), .Z(n340) );
  NOR U356 ( .A(n340), .B(n373), .Z(n328) );
  NOR U357 ( .A(n329), .B(n328), .Z(n330) );
  IV U358 ( .A(n330), .Z(n331) );
  NOR U359 ( .A(n360), .B(n331), .Z(n332) );
  NOR U360 ( .A(x[3]), .B(n332), .Z(n358) );
  XOR U361 ( .A(n334), .B(n333), .Z(n335) );
  XOR U362 ( .A(n336), .B(n335), .Z(n337) );
  NOR U363 ( .A(n367), .B(n337), .Z(n355) );
  NOR U364 ( .A(n339), .B(n338), .Z(n346) );
  NOR U365 ( .A(n340), .B(y[3]), .Z(n343) );
  NOR U366 ( .A(n341), .B(n373), .Z(n342) );
  NOR U367 ( .A(n343), .B(n342), .Z(n344) );
  IV U368 ( .A(n344), .Z(n345) );
  NOR U369 ( .A(n346), .B(n345), .Z(n347) );
  NOR U370 ( .A(n347), .B(n362), .Z(n352) );
  XOR U371 ( .A(x[3]), .B(n348), .Z(n349) );
  NOR U372 ( .A(n350), .B(n349), .Z(n351) );
  NOR U373 ( .A(n352), .B(n351), .Z(n353) );
  IV U374 ( .A(n353), .Z(n354) );
  NOR U375 ( .A(n355), .B(n354), .Z(n356) );
  IV U376 ( .A(n356), .Z(n357) );
  NOR U377 ( .A(n358), .B(n357), .Z(n359) );
  IV U378 ( .A(n359), .Z(o[3]) );
  NOR U379 ( .A(n361), .B(n360), .Z(n363) );
  NOR U380 ( .A(n363), .B(n362), .Z(n369) );
  XOR U381 ( .A(n365), .B(n364), .Z(n366) );
  NOR U382 ( .A(n367), .B(n366), .Z(n368) );
  NOR U383 ( .A(n369), .B(n368), .Z(n370) );
  IV U384 ( .A(n370), .Z(n381) );
  NOR U385 ( .A(x[3]), .B(n371), .Z(n376) );
  NOR U386 ( .A(n373), .B(n372), .Z(n374) );
  IV U387 ( .A(n374), .Z(n375) );
  NOR U388 ( .A(n376), .B(n375), .Z(n378) );
  NOR U389 ( .A(n378), .B(n377), .Z(n379) );
  IV U390 ( .A(n379), .Z(n380) );
  NOR U391 ( .A(n381), .B(n380), .Z(n382) );
  IV U392 ( .A(n382), .Z(o[4]) );
endmodule

