
module FA_2016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_2048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_2976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_97 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_2976 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_2944 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_2912 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_2880 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_2848 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_2816 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_2784 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_2752 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_2720 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_2688 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_2656 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_2624 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_2592 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_2560 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_2528 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_2496 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_2464 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_2432 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_2400 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_2368 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_2336 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_2304 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_2272 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_2240 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_2208 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_2176 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_2144 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_2112 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_2080 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_2048 \FAINST[30].FA_  ( .A(1'b0), .B(B[30]), .CI(1'b0), .S(S[30]) );
  FA_2016 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(1'b0), .S(S[31]) );
endmodule


module FA_3009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_98 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;
  wire   \C[31] ;

  FA_3039 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3038 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3037 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3036 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3035 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3034 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3033 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3032 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3031 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3030 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3029 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3028 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3027 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3026 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3025 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3024 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3023 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3022 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3021 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3020 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3019 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3018 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3017 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3016 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3015 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3014 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3013 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_3012 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_3011 \FAINST[29].FA_  ( .A(1'b0), .B(B[29]), .CI(1'b0), .S(S[29]) );
  FA_3010 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(1'b0), .S(S[30]), .CO(
        \C[31] ) );
  FA_3009 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(\C[31] ), .S(S[31]) );
endmodule


module FA_3041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_99 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3071 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3070 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3069 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3068 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3067 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3066 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3065 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3064 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3063 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3062 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3061 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3060 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3059 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3058 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3057 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3056 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3055 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3054 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3053 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3052 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3051 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3050 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3049 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3048 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3047 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3046 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3045 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_3044 \FAINST[28].FA_  ( .A(1'b0), .B(B[28]), .CI(1'b0), .S(S[28]) );
  FA_3043 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(1'b0), .S(S[29]), .CO(
        C[30]) );
  FA_3042 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3041 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_100 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3103 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3102 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3101 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3100 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3099 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3098 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3097 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3096 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3095 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3094 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3093 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3092 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3091 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3090 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3089 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3088 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3087 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3086 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3085 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3084 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3083 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3082 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3081 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3080 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3079 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3078 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3077 \FAINST[27].FA_  ( .A(1'b0), .B(B[27]), .CI(1'b0), .S(S[27]) );
  FA_3076 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(1'b0), .S(S[28]), .CO(
        C[29]) );
  FA_3075 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3074 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3073 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_101 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3135 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3134 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3133 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3132 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3131 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3130 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3129 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3128 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3127 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3126 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3125 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3124 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3123 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3122 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3121 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3120 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3119 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3118 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3117 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3116 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3115 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3114 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3113 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3112 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3111 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3110 \FAINST[26].FA_  ( .A(1'b0), .B(B[26]), .CI(1'b0), .S(S[26]) );
  FA_3109 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(1'b0), .S(S[27]), .CO(
        C[28]) );
  FA_3108 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3107 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3106 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3105 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_102 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3167 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3166 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3165 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3164 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3163 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3162 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3161 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3160 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3159 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3158 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3157 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3156 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3155 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3154 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3153 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3152 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3151 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3150 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3149 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3148 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3147 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3146 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3145 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3144 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3143 \FAINST[25].FA_  ( .A(1'b0), .B(B[25]), .CI(1'b0), .S(S[25]) );
  FA_3142 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(1'b0), .S(S[26]), .CO(
        C[27]) );
  FA_3141 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3140 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3139 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3138 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3137 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_103 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3199 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3198 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3197 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3196 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3195 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3194 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3193 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3192 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3191 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3190 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3189 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3188 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3187 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3186 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3185 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3184 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3183 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3182 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3181 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3180 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3179 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3178 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3177 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3176 \FAINST[24].FA_  ( .A(1'b0), .B(B[24]), .CI(1'b0), .S(S[24]) );
  FA_3175 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(1'b0), .S(S[25]), .CO(
        C[26]) );
  FA_3174 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3173 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3172 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3171 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3170 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3169 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_104 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3231 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3230 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3229 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3228 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3227 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3226 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3225 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3224 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3223 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3222 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3221 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3220 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3219 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3218 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3217 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3216 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3215 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3214 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3213 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3212 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3211 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3210 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3209 \FAINST[23].FA_  ( .A(1'b0), .B(B[23]), .CI(1'b0), .S(S[23]) );
  FA_3208 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(1'b0), .S(S[24]), .CO(
        C[25]) );
  FA_3207 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3206 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3205 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3204 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3203 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3202 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3201 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_105 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3263 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3262 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3261 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3260 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3259 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3258 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3257 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3256 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3255 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3254 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3253 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3252 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3251 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3250 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3249 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3248 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3247 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3246 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3245 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3244 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3243 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3242 \FAINST[22].FA_  ( .A(1'b0), .B(B[22]), .CI(1'b0), .S(S[22]) );
  FA_3241 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(1'b0), .S(S[23]), .CO(
        C[24]) );
  FA_3240 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3239 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3238 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3237 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3236 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3235 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3234 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3233 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_106 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3295 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3294 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3293 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3292 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3291 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3290 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3289 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3288 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3287 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3286 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3285 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3284 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3283 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3282 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3281 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3280 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3279 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3278 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3277 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3276 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3275 \FAINST[21].FA_  ( .A(1'b0), .B(B[21]), .CI(1'b0), .S(S[21]) );
  FA_3274 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(1'b0), .S(S[22]), .CO(
        C[23]) );
  FA_3273 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3272 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3271 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3270 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3269 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3268 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3267 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3266 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3265 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_107 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3327 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3326 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3325 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3324 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3323 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3322 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3321 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3320 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3319 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3318 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3317 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3316 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3315 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3314 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3313 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3312 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3311 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3310 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3309 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3308 \FAINST[20].FA_  ( .A(1'b0), .B(B[20]), .CI(1'b0), .S(S[20]) );
  FA_3307 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(1'b0), .S(S[21]), .CO(
        C[22]) );
  FA_3306 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3305 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3304 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3303 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3302 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3301 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3300 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3299 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3298 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3297 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_108 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3359 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3358 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3357 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3356 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3355 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3354 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3353 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3352 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3351 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3350 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3349 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3348 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3347 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3346 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3345 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3344 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3343 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3342 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3341 \FAINST[19].FA_  ( .A(1'b0), .B(B[19]), .CI(1'b0), .S(S[19]) );
  FA_3340 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(1'b0), .S(S[20]), .CO(
        C[21]) );
  FA_3339 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3338 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3337 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3336 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3335 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3334 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3333 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3332 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3331 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3330 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3329 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_109 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3391 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3390 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3389 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3388 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3387 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3386 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3385 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3384 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3383 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3382 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3381 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3380 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3379 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3378 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3377 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3376 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3375 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3374 \FAINST[18].FA_  ( .A(1'b0), .B(B[18]), .CI(1'b0), .S(S[18]) );
  FA_3373 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(1'b0), .S(S[19]), .CO(
        C[20]) );
  FA_3372 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3371 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3370 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3369 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3368 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3367 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3366 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3365 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3364 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3363 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3362 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3361 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_110 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3423 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3422 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3421 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3420 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3419 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3418 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3417 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3416 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3415 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3414 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3413 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3412 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3411 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3410 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3409 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3408 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3407 \FAINST[17].FA_  ( .A(1'b0), .B(B[17]), .CI(1'b0), .S(S[17]) );
  FA_3406 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(1'b0), .S(S[18]), .CO(
        C[19]) );
  FA_3405 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3404 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3403 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3402 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3401 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3400 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3399 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3398 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3397 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3396 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3395 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3394 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3393 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_111 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3455 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3454 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3453 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3452 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3451 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3450 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3449 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3448 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3447 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3446 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3445 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3444 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3443 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3442 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3441 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3440 \FAINST[16].FA_  ( .A(1'b0), .B(B[16]), .CI(1'b0), .S(S[16]) );
  FA_3439 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(1'b0), .S(S[17]), .CO(
        C[18]) );
  FA_3438 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3437 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3436 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3435 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3434 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3433 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3432 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3431 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3430 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3429 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3428 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3427 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3426 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3425 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_112 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3487 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3486 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3485 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3484 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3483 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3482 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3481 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3480 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3479 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3478 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3477 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3476 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3475 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3474 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3473 \FAINST[15].FA_  ( .A(1'b0), .B(B[15]), .CI(1'b0), .S(S[15]) );
  FA_3472 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(1'b0), .S(S[16]), .CO(
        C[17]) );
  FA_3471 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3470 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3469 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3468 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3467 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3466 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3465 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3464 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3463 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3462 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3461 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3460 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3459 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3458 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3457 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_113 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3519 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3518 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3517 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3516 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3515 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3514 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3513 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3512 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3511 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3510 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3509 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3508 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3507 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3506 \FAINST[14].FA_  ( .A(1'b0), .B(B[14]), .CI(1'b0), .S(S[14]) );
  FA_3505 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(1'b0), .S(S[15]), .CO(
        C[16]) );
  FA_3504 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3503 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3502 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3501 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3500 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3499 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3498 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3497 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3496 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3495 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3494 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3493 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3492 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3491 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3490 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3489 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_114 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3551 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3550 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3549 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3548 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3547 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3546 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3545 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3544 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3543 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3542 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3541 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3540 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3539 \FAINST[13].FA_  ( .A(1'b0), .B(B[13]), .CI(1'b0), .S(S[13]) );
  FA_3538 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(1'b0), .S(S[14]), .CO(
        C[15]) );
  FA_3537 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3536 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3535 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3534 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3533 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3532 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3531 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3530 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3529 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3528 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3527 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3526 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3525 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3524 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3523 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3522 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3521 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_115 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3583 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3582 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3581 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3580 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3579 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3578 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3577 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3576 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3575 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3574 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3573 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3572 \FAINST[12].FA_  ( .A(1'b0), .B(B[12]), .CI(1'b0), .S(S[12]) );
  FA_3571 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(1'b0), .S(S[13]), .CO(
        C[14]) );
  FA_3570 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3569 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3568 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3567 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3566 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3565 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3564 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3563 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3562 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3561 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3560 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3559 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3558 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3557 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3556 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3555 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3554 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3553 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_116 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3615 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3614 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3613 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3612 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3611 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3610 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3609 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3608 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3607 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3606 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3605 \FAINST[11].FA_  ( .A(1'b0), .B(B[11]), .CI(1'b0), .S(S[11]) );
  FA_3604 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(1'b0), .S(S[12]), .CO(
        C[13]) );
  FA_3603 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3602 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3601 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3600 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3599 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3598 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3597 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3596 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3595 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3594 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3593 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3592 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3591 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3590 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3589 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3588 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3587 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3586 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3585 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_117 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3647 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3646 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3645 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3644 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3643 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3642 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3641 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3640 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3639 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3638 \FAINST[10].FA_  ( .A(1'b0), .B(B[10]), .CI(1'b0), .S(S[10]) );
  FA_3637 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(1'b0), .S(S[11]), .CO(
        C[12]) );
  FA_3636 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3635 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3634 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3633 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3632 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3631 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3630 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3629 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3628 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3627 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3626 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3625 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3624 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3623 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3622 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3621 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3620 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3619 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3618 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3617 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_118 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3679 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3678 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3677 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3676 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3675 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3674 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3673 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3672 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3671 \FAINST[9].FA_  ( .A(1'b0), .B(B[9]), .CI(1'b0), .S(S[9]) );
  FA_3670 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(1'b0), .S(S[10]), .CO(
        C[11]) );
  FA_3669 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3668 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3667 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3666 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3665 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3664 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3663 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3662 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3661 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3660 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3659 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3658 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3657 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3656 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3655 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3654 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3653 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3652 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3651 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3650 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3649 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_119 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3711 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3710 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3709 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3708 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3707 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3706 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3705 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3704 \FAINST[8].FA_  ( .A(1'b0), .B(B[8]), .CI(1'b0), .S(S[8]) );
  FA_3703 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(1'b0), .S(S[9]), .CO(C[10]) );
  FA_3702 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3701 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3700 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3699 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3698 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3697 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3696 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3695 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3694 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3693 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3692 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3691 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3690 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3689 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3688 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3687 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3686 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3685 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3684 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3683 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3682 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3681 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_120 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3743 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3742 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3741 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3740 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3739 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3738 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3737 \FAINST[7].FA_  ( .A(1'b0), .B(B[7]), .CI(1'b0), .S(S[7]) );
  FA_3736 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(1'b0), .S(S[8]), .CO(C[9])
         );
  FA_3735 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3734 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3733 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3732 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3731 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3730 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3729 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3728 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3727 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3726 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3725 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3724 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3723 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3722 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3721 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3720 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3719 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3718 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3717 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3716 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3715 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3714 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3713 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_121 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3775 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3774 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3773 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3772 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3771 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3770 \FAINST[6].FA_  ( .A(1'b0), .B(B[6]), .CI(1'b0), .S(S[6]) );
  FA_3769 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(1'b0), .S(S[7]), .CO(C[8])
         );
  FA_3768 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3767 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3766 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3765 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3764 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3763 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3762 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3761 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3760 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3759 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3758 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3757 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3756 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3755 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3754 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3753 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3752 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3751 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3750 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3749 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3748 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3747 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3746 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3745 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_122 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3807 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3806 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3805 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3804 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3803 \FAINST[5].FA_  ( .A(1'b0), .B(B[5]), .CI(1'b0), .S(S[5]) );
  FA_3802 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(1'b0), .S(S[6]), .CO(C[7])
         );
  FA_3801 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3800 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3799 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3798 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3797 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3796 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3795 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3794 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3793 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3792 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3791 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3790 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3789 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3788 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3787 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3786 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3785 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3784 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3783 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3782 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3781 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3780 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3779 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3778 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3777 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_123 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3839 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3838 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3837 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3836 \FAINST[4].FA_  ( .A(1'b0), .B(B[4]), .CI(1'b0), .S(S[4]) );
  FA_3835 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(1'b0), .S(S[5]), .CO(C[6])
         );
  FA_3834 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3833 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3832 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3831 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3830 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3829 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3828 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3827 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3826 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3825 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3824 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3823 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3822 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3821 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3820 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3819 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3818 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3817 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3816 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3815 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3814 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3813 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3812 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3811 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3810 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3809 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_124 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3871 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3870 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3869 \FAINST[3].FA_  ( .A(1'b0), .B(B[3]), .CI(1'b0), .S(S[3]) );
  FA_3868 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(1'b0), .S(S[4]), .CO(C[5])
         );
  FA_3867 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3866 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3865 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3864 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3863 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3862 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3861 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3860 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3859 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3858 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3857 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3856 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3855 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3854 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3853 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3852 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3851 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3850 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3849 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3848 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3847 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3846 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3845 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3844 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3843 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3842 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3841 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_3903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_125 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3903 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3902 \FAINST[2].FA_  ( .A(1'b0), .B(B[2]), .CI(1'b0), .S(S[2]) );
  FA_3901 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(1'b0), .S(S[3]), .CO(C[4])
         );
  FA_3900 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3899 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3898 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3897 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3896 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3895 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3894 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3893 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3892 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3891 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3890 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3889 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3888 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3887 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3886 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3885 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3884 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3883 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3882 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3881 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3880 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3879 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3878 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3877 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3876 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3875 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3874 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3873 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_3935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N32_126 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3935 \FAINST[1].FA_  ( .A(1'b0), .B(B[1]), .CI(1'b0), .S(S[1]) );
  FA_3934 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(1'b0), .S(S[2]), .CO(C[3])
         );
  FA_3933 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3932 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3931 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3930 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3929 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3928 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3927 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3926 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3925 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3924 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3923 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3922 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3921 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3920 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3919 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3918 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3917 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3916 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3915 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3914 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3913 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3912 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3911 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3910 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3909 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3908 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3907 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3906 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3905 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module FA_3937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module FA_3967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   A;
  assign S = A;

endmodule


module ADD_N32_127 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;


  FA_3967 \FAINST[1].FA_  ( .A(A[1]), .B(1'b0), .CI(1'b0), .S(S[1]) );
  FA_3966 \FAINST[2].FA_  ( .A(A[2]), .B(1'b0), .CI(1'b0), .S(S[2]) );
  FA_3965 \FAINST[3].FA_  ( .A(A[3]), .B(1'b0), .CI(1'b0), .S(S[3]) );
  FA_3964 \FAINST[4].FA_  ( .A(A[4]), .B(1'b0), .CI(1'b0), .S(S[4]) );
  FA_3963 \FAINST[5].FA_  ( .A(A[5]), .B(1'b0), .CI(1'b0), .S(S[5]) );
  FA_3962 \FAINST[6].FA_  ( .A(A[6]), .B(1'b0), .CI(1'b0), .S(S[6]) );
  FA_3961 \FAINST[7].FA_  ( .A(A[7]), .B(1'b0), .CI(1'b0), .S(S[7]) );
  FA_3960 \FAINST[8].FA_  ( .A(A[8]), .B(1'b0), .CI(1'b0), .S(S[8]) );
  FA_3959 \FAINST[9].FA_  ( .A(A[9]), .B(1'b0), .CI(1'b0), .S(S[9]) );
  FA_3958 \FAINST[10].FA_  ( .A(A[10]), .B(1'b0), .CI(1'b0), .S(S[10]) );
  FA_3957 \FAINST[11].FA_  ( .A(A[11]), .B(1'b0), .CI(1'b0), .S(S[11]) );
  FA_3956 \FAINST[12].FA_  ( .A(A[12]), .B(1'b0), .CI(1'b0), .S(S[12]) );
  FA_3955 \FAINST[13].FA_  ( .A(A[13]), .B(1'b0), .CI(1'b0), .S(S[13]) );
  FA_3954 \FAINST[14].FA_  ( .A(A[14]), .B(1'b0), .CI(1'b0), .S(S[14]) );
  FA_3953 \FAINST[15].FA_  ( .A(A[15]), .B(1'b0), .CI(1'b0), .S(S[15]) );
  FA_3952 \FAINST[16].FA_  ( .A(A[16]), .B(1'b0), .CI(1'b0), .S(S[16]) );
  FA_3951 \FAINST[17].FA_  ( .A(A[17]), .B(1'b0), .CI(1'b0), .S(S[17]) );
  FA_3950 \FAINST[18].FA_  ( .A(A[18]), .B(1'b0), .CI(1'b0), .S(S[18]) );
  FA_3949 \FAINST[19].FA_  ( .A(A[19]), .B(1'b0), .CI(1'b0), .S(S[19]) );
  FA_3948 \FAINST[20].FA_  ( .A(A[20]), .B(1'b0), .CI(1'b0), .S(S[20]) );
  FA_3947 \FAINST[21].FA_  ( .A(A[21]), .B(1'b0), .CI(1'b0), .S(S[21]) );
  FA_3946 \FAINST[22].FA_  ( .A(A[22]), .B(1'b0), .CI(1'b0), .S(S[22]) );
  FA_3945 \FAINST[23].FA_  ( .A(A[23]), .B(1'b0), .CI(1'b0), .S(S[23]) );
  FA_3944 \FAINST[24].FA_  ( .A(A[24]), .B(1'b0), .CI(1'b0), .S(S[24]) );
  FA_3943 \FAINST[25].FA_  ( .A(A[25]), .B(1'b0), .CI(1'b0), .S(S[25]) );
  FA_3942 \FAINST[26].FA_  ( .A(A[26]), .B(1'b0), .CI(1'b0), .S(S[26]) );
  FA_3941 \FAINST[27].FA_  ( .A(A[27]), .B(1'b0), .CI(1'b0), .S(S[27]) );
  FA_3940 \FAINST[28].FA_  ( .A(A[28]), .B(1'b0), .CI(1'b0), .S(S[28]) );
  FA_3939 \FAINST[29].FA_  ( .A(A[29]), .B(1'b0), .CI(1'b0), .S(S[29]) );
  FA_3938 \FAINST[30].FA_  ( .A(A[30]), .B(1'b0), .CI(1'b0), .S(S[30]) );
  FA_3937 \FAINST[31].FA_  ( .A(A[31]), .B(1'b0), .CI(1'b0), .S(S[31]) );
endmodule


module MULT_N32_3 ( A, B, O );
  input [31:0] A;
  input [31:0] B;
  output [31:0] O;
  wire   \w[31][31] , \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] ,
         \w[31][26] , \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] ,
         \w[31][21] , \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] ,
         \w[31][16] , \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] ,
         \w[31][11] , \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] ,
         \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] ,
         \w[31][1] , \w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] ,
         \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] ,
         \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] ,
         \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] ,
         \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] ,
         \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] ,
         \w[30][2] , \w[30][1] , \w[29][31] , \w[29][30] , \w[29][29] ,
         \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] ,
         \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] ,
         \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] ,
         \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] ,
         \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] ,
         \w[29][3] , \w[29][2] , \w[29][1] , \w[28][31] , \w[28][30] ,
         \w[28][29] , \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] ,
         \w[28][24] , \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] ,
         \w[28][19] , \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] ,
         \w[28][14] , \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] ,
         \w[28][9] , \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] ,
         \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , \w[27][31] ,
         \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] ,
         \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] ,
         \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] ,
         \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] ,
         \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] ,
         \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] ,
         \w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] ,
         \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] ,
         \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] ,
         \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] ,
         \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] ,
         \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] ,
         \w[26][1] , \w[25][31] , \w[25][30] , \w[25][29] , \w[25][28] ,
         \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , \w[25][23] ,
         \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , \w[25][18] ,
         \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , \w[25][13] ,
         \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , \w[25][8] ,
         \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] ,
         \w[25][2] , \w[25][1] , \w[24][31] , \w[24][30] , \w[24][29] ,
         \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] ,
         \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] ,
         \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] ,
         \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] ,
         \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] ,
         \w[24][3] , \w[24][2] , \w[24][1] , \w[23][31] , \w[23][30] ,
         \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] ,
         \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] ,
         \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] ,
         \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] ,
         \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] ,
         \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , \w[22][31] ,
         \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , \w[22][26] ,
         \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , \w[22][21] ,
         \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , \w[22][16] ,
         \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , \w[22][11] ,
         \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , \w[22][6] ,
         \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] ,
         \w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] ,
         \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] ,
         \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] ,
         \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] ,
         \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] ,
         \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] ,
         \w[21][1] , \w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] ,
         \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] ,
         \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] ,
         \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] ,
         \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] ,
         \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] ,
         \w[20][2] , \w[20][1] , \w[19][31] , \w[19][30] , \w[19][29] ,
         \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] ,
         \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] ,
         \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] ,
         \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] ,
         \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] ,
         \w[19][3] , \w[19][2] , \w[19][1] , \w[18][31] , \w[18][30] ,
         \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] ,
         \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] ,
         \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] ,
         \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] ,
         \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] ,
         \w[18][4] , \w[18][3] , \w[18][2] , \w[18][1] , \w[17][31] ,
         \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] ,
         \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] ,
         \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] ,
         \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] ,
         \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] ,
         \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] ,
         \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] ,
         \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] ,
         \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] ,
         \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] ,
         \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] ,
         \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] ,
         \w[16][1] , \w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] ,
         \w[15][27] , \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] ,
         \w[15][22] , \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] ,
         \w[15][17] , \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] ,
         \w[15][12] , \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] ,
         \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] ,
         \w[15][2] , \w[15][1] , \w[14][31] , \w[14][30] , \w[14][29] ,
         \w[14][28] , \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] ,
         \w[14][23] , \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] ,
         \w[14][18] , \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] ,
         \w[14][13] , \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] ,
         \w[14][8] , \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] ,
         \w[14][3] , \w[14][2] , \w[14][1] , \w[13][31] , \w[13][30] ,
         \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] ,
         \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] ,
         \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] ,
         \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] ,
         \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] ,
         \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , \w[12][31] ,
         \w[12][30] , \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] ,
         \w[12][25] , \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] ,
         \w[12][20] , \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] ,
         \w[12][15] , \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] ,
         \w[12][10] , \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] ,
         \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , \w[12][1] ,
         \w[11][31] , \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] ,
         \w[11][26] , \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] ,
         \w[11][21] , \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] ,
         \w[11][16] , \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] ,
         \w[11][11] , \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] ,
         \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] ,
         \w[11][1] , \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] ,
         \w[10][27] , \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] ,
         \w[10][22] , \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] ,
         \w[10][17] , \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] ,
         \w[10][12] , \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] ,
         \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] ,
         \w[10][2] , \w[10][1] , \w[9][31] , \w[9][30] , \w[9][29] ,
         \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] ,
         \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] ,
         \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] ,
         \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] ,
         \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] ,
         \w[9][1] , \w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] ,
         \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] ,
         \w[8][21] , \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] ,
         \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , \w[8][12] ,
         \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , \w[8][6] ,
         \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , \w[7][31] ,
         \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] ,
         \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] ,
         \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] ,
         \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] ,
         \w[7][10] , \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] ,
         \w[7][4] , \w[7][3] , \w[7][2] , \w[7][1] , \w[6][31] , \w[6][30] ,
         \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] ,
         \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] ,
         \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] ,
         \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] ,
         \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] ,
         \w[6][2] , \w[6][1] , \w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] ,
         \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] ,
         \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] ,
         \w[5][17] , \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] ,
         \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] ,
         \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] ,
         \w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] ,
         \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] ,
         \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] ,
         \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] ,
         \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] ,
         \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , \w[3][31] ,
         \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] ,
         \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] ,
         \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] ,
         \w[3][15] , \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] ,
         \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] ,
         \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , \w[2][31] , \w[2][30] ,
         \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] ,
         \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] ,
         \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] ,
         \w[2][14] , \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] ,
         \w[2][8] , \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] ,
         \w[2][2] , \w[2][1] , \_0_net_[31] , \_0_net_[30] , \_0_net_[29] ,
         \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , \_0_net_[25] ,
         \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , \_0_net_[21] ,
         \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , \_0_net_[17] ,
         \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , \_0_net_[13] ,
         \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , \_0_net_[9] ,
         \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , \_0_net_[4] ,
         \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , \_2_net_[31] ,
         \_2_net_[30] , \_2_net_[29] , \_2_net_[28] , \_2_net_[27] ,
         \_2_net_[26] , \_2_net_[25] , \_2_net_[24] , \_2_net_[23] ,
         \_2_net_[22] , \_2_net_[21] , \_2_net_[20] , \_2_net_[19] ,
         \_2_net_[18] , \_2_net_[17] , \_2_net_[16] , \_2_net_[15] ,
         \_2_net_[14] , \_2_net_[13] , \_2_net_[12] , \_2_net_[11] ,
         \_2_net_[10] , \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] ,
         \_2_net_[5] , \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , \_4_net_[31] ,
         \_4_net_[30] , \_4_net_[29] , \_4_net_[28] , \_4_net_[27] ,
         \_4_net_[26] , \_4_net_[25] , \_4_net_[24] , \_4_net_[23] ,
         \_4_net_[22] , \_4_net_[21] , \_4_net_[20] , \_4_net_[19] ,
         \_4_net_[18] , \_4_net_[17] , \_4_net_[16] , \_4_net_[15] ,
         \_4_net_[14] , \_4_net_[13] , \_4_net_[12] , \_4_net_[11] ,
         \_4_net_[10] , \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] ,
         \_4_net_[5] , \_4_net_[4] , \_4_net_[3] , \_6_net_[31] ,
         \_6_net_[30] , \_6_net_[29] , \_6_net_[28] , \_6_net_[27] ,
         \_6_net_[26] , \_6_net_[25] , \_6_net_[24] , \_6_net_[23] ,
         \_6_net_[22] , \_6_net_[21] , \_6_net_[20] , \_6_net_[19] ,
         \_6_net_[18] , \_6_net_[17] , \_6_net_[16] , \_6_net_[15] ,
         \_6_net_[14] , \_6_net_[13] , \_6_net_[12] , \_6_net_[11] ,
         \_6_net_[10] , \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] ,
         \_6_net_[5] , \_6_net_[4] , \_8_net_[31] , \_8_net_[30] ,
         \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] ,
         \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] ,
         \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] ,
         \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] ,
         \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] ,
         \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] ,
         \_10_net_[31] , \_10_net_[30] , \_10_net_[29] , \_10_net_[28] ,
         \_10_net_[27] , \_10_net_[26] , \_10_net_[25] , \_10_net_[24] ,
         \_10_net_[23] , \_10_net_[22] , \_10_net_[21] , \_10_net_[20] ,
         \_10_net_[19] , \_10_net_[18] , \_10_net_[17] , \_10_net_[16] ,
         \_10_net_[15] , \_10_net_[14] , \_10_net_[13] , \_10_net_[12] ,
         \_10_net_[11] , \_10_net_[10] , \_10_net_[9] , \_10_net_[8] ,
         \_10_net_[7] , \_10_net_[6] , \_12_net_[31] , \_12_net_[30] ,
         \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] ,
         \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] ,
         \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] ,
         \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] ,
         \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] ,
         \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , \_14_net_[31] ,
         \_14_net_[30] , \_14_net_[29] , \_14_net_[28] , \_14_net_[27] ,
         \_14_net_[26] , \_14_net_[25] , \_14_net_[24] , \_14_net_[23] ,
         \_14_net_[22] , \_14_net_[21] , \_14_net_[20] , \_14_net_[19] ,
         \_14_net_[18] , \_14_net_[17] , \_14_net_[16] , \_14_net_[15] ,
         \_14_net_[14] , \_14_net_[13] , \_14_net_[12] , \_14_net_[11] ,
         \_14_net_[10] , \_14_net_[9] , \_14_net_[8] , \_16_net_[31] ,
         \_16_net_[30] , \_16_net_[29] , \_16_net_[28] , \_16_net_[27] ,
         \_16_net_[26] , \_16_net_[25] , \_16_net_[24] , \_16_net_[23] ,
         \_16_net_[22] , \_16_net_[21] , \_16_net_[20] , \_16_net_[19] ,
         \_16_net_[18] , \_16_net_[17] , \_16_net_[16] , \_16_net_[15] ,
         \_16_net_[14] , \_16_net_[13] , \_16_net_[12] , \_16_net_[11] ,
         \_16_net_[10] , \_16_net_[9] , \_18_net_[31] , \_18_net_[30] ,
         \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] ,
         \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] ,
         \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] ,
         \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] ,
         \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] ,
         \_20_net_[31] , \_20_net_[30] , \_20_net_[29] , \_20_net_[28] ,
         \_20_net_[27] , \_20_net_[26] , \_20_net_[25] , \_20_net_[24] ,
         \_20_net_[23] , \_20_net_[22] , \_20_net_[21] , \_20_net_[20] ,
         \_20_net_[19] , \_20_net_[18] , \_20_net_[17] , \_20_net_[16] ,
         \_20_net_[15] , \_20_net_[14] , \_20_net_[13] , \_20_net_[12] ,
         \_20_net_[11] , \_22_net_[31] , \_22_net_[30] , \_22_net_[29] ,
         \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , \_22_net_[25] ,
         \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , \_22_net_[21] ,
         \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , \_22_net_[17] ,
         \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , \_22_net_[13] ,
         \_22_net_[12] , \_24_net_[31] , \_24_net_[30] , \_24_net_[29] ,
         \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , \_24_net_[25] ,
         \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , \_24_net_[21] ,
         \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , \_24_net_[17] ,
         \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , \_24_net_[13] ,
         \_26_net_[31] , \_26_net_[30] , \_26_net_[29] , \_26_net_[28] ,
         \_26_net_[27] , \_26_net_[26] , \_26_net_[25] , \_26_net_[24] ,
         \_26_net_[23] , \_26_net_[22] , \_26_net_[21] , \_26_net_[20] ,
         \_26_net_[19] , \_26_net_[18] , \_26_net_[17] , \_26_net_[16] ,
         \_26_net_[15] , \_26_net_[14] , \_28_net_[31] , \_28_net_[30] ,
         \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] ,
         \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] ,
         \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] ,
         \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , \_30_net_[31] ,
         \_30_net_[30] , \_30_net_[29] , \_30_net_[28] , \_30_net_[27] ,
         \_30_net_[26] , \_30_net_[25] , \_30_net_[24] , \_30_net_[23] ,
         \_30_net_[22] , \_30_net_[21] , \_30_net_[20] , \_30_net_[19] ,
         \_30_net_[18] , \_30_net_[17] , \_30_net_[16] , \_32_net_[31] ,
         \_32_net_[30] , \_32_net_[29] , \_32_net_[28] , \_32_net_[27] ,
         \_32_net_[26] , \_32_net_[25] , \_32_net_[24] , \_32_net_[23] ,
         \_32_net_[22] , \_32_net_[21] , \_32_net_[20] , \_32_net_[19] ,
         \_32_net_[18] , \_32_net_[17] , \_34_net_[31] , \_34_net_[30] ,
         \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] ,
         \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] ,
         \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] ,
         \_36_net_[31] , \_36_net_[30] , \_36_net_[29] , \_36_net_[28] ,
         \_36_net_[27] , \_36_net_[26] , \_36_net_[25] , \_36_net_[24] ,
         \_36_net_[23] , \_36_net_[22] , \_36_net_[21] , \_36_net_[20] ,
         \_36_net_[19] , \_38_net_[31] , \_38_net_[30] , \_38_net_[29] ,
         \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , \_38_net_[25] ,
         \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , \_38_net_[21] ,
         \_38_net_[20] , \_40_net_[31] , \_40_net_[30] , \_40_net_[29] ,
         \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , \_40_net_[25] ,
         \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , \_40_net_[21] ,
         \_42_net_[31] , \_42_net_[30] , \_42_net_[29] , \_42_net_[28] ,
         \_42_net_[27] , \_42_net_[26] , \_42_net_[25] , \_42_net_[24] ,
         \_42_net_[23] , \_42_net_[22] , \_44_net_[31] , \_44_net_[30] ,
         \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] ,
         \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , \_46_net_[31] ,
         \_46_net_[30] , \_46_net_[29] , \_46_net_[28] , \_46_net_[27] ,
         \_46_net_[26] , \_46_net_[25] , \_46_net_[24] , \_48_net_[31] ,
         \_48_net_[30] , \_48_net_[29] , \_48_net_[28] , \_48_net_[27] ,
         \_48_net_[26] , \_48_net_[25] , \_50_net_[31] , \_50_net_[30] ,
         \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] ,
         \_52_net_[31] , \_52_net_[30] , \_52_net_[29] , \_52_net_[28] ,
         \_52_net_[27] , \_54_net_[31] , \_54_net_[30] , \_54_net_[29] ,
         \_54_net_[28] , \_56_net_[31] , \_56_net_[30] , \_56_net_[29] ,
         \_58_net_[31] , \_58_net_[30] , \_60_net_[31] ;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  ADD_N32_127 \FAINST[1].ADD_  ( .A({\_0_net_[31] , \_0_net_[30] , 
        \_0_net_[29] , \_0_net_[28] , \_0_net_[27] , \_0_net_[26] , 
        \_0_net_[25] , \_0_net_[24] , \_0_net_[23] , \_0_net_[22] , 
        \_0_net_[21] , \_0_net_[20] , \_0_net_[19] , \_0_net_[18] , 
        \_0_net_[17] , \_0_net_[16] , \_0_net_[15] , \_0_net_[14] , 
        \_0_net_[13] , \_0_net_[12] , \_0_net_[11] , \_0_net_[10] , 
        \_0_net_[9] , \_0_net_[8] , \_0_net_[7] , \_0_net_[6] , \_0_net_[5] , 
        \_0_net_[4] , \_0_net_[3] , \_0_net_[2] , \_0_net_[1] , 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .S({
        \w[2][31] , \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , 
        \w[2][25] , \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , 
        \w[2][19] , \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , 
        \w[2][13] , \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , 
        \w[2][7] , \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , 
        \w[2][1] , SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_126 \FAINST[2].ADD_  ( .A({\_2_net_[31] , \_2_net_[30] , 
        \_2_net_[29] , \_2_net_[28] , \_2_net_[27] , \_2_net_[26] , 
        \_2_net_[25] , \_2_net_[24] , \_2_net_[23] , \_2_net_[22] , 
        \_2_net_[21] , \_2_net_[20] , \_2_net_[19] , \_2_net_[18] , 
        \_2_net_[17] , \_2_net_[16] , \_2_net_[15] , \_2_net_[14] , 
        \_2_net_[13] , \_2_net_[12] , \_2_net_[11] , \_2_net_[10] , 
        \_2_net_[9] , \_2_net_[8] , \_2_net_[7] , \_2_net_[6] , \_2_net_[5] , 
        \_2_net_[4] , \_2_net_[3] , \_2_net_[2] , 1'b0, 1'b0}), .B({\w[2][31] , 
        \w[2][30] , \w[2][29] , \w[2][28] , \w[2][27] , \w[2][26] , \w[2][25] , 
        \w[2][24] , \w[2][23] , \w[2][22] , \w[2][21] , \w[2][20] , \w[2][19] , 
        \w[2][18] , \w[2][17] , \w[2][16] , \w[2][15] , \w[2][14] , \w[2][13] , 
        \w[2][12] , \w[2][11] , \w[2][10] , \w[2][9] , \w[2][8] , \w[2][7] , 
        \w[2][6] , \w[2][5] , \w[2][4] , \w[2][3] , \w[2][2] , \w[2][1] , 1'b0}), .CI(1'b0), .S({\w[3][31] , \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , 
        \w[3][26] , \w[3][25] , \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , 
        \w[3][20] , \w[3][19] , \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , 
        \w[3][14] , \w[3][13] , \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , 
        \w[3][8] , \w[3][7] , \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , 
        \w[3][2] , \w[3][1] , SYNOPSYS_UNCONNECTED__1}) );
  ADD_N32_125 \FAINST[3].ADD_  ( .A({\_4_net_[31] , \_4_net_[30] , 
        \_4_net_[29] , \_4_net_[28] , \_4_net_[27] , \_4_net_[26] , 
        \_4_net_[25] , \_4_net_[24] , \_4_net_[23] , \_4_net_[22] , 
        \_4_net_[21] , \_4_net_[20] , \_4_net_[19] , \_4_net_[18] , 
        \_4_net_[17] , \_4_net_[16] , \_4_net_[15] , \_4_net_[14] , 
        \_4_net_[13] , \_4_net_[12] , \_4_net_[11] , \_4_net_[10] , 
        \_4_net_[9] , \_4_net_[8] , \_4_net_[7] , \_4_net_[6] , \_4_net_[5] , 
        \_4_net_[4] , \_4_net_[3] , 1'b0, 1'b0, 1'b0}), .B({\w[3][31] , 
        \w[3][30] , \w[3][29] , \w[3][28] , \w[3][27] , \w[3][26] , \w[3][25] , 
        \w[3][24] , \w[3][23] , \w[3][22] , \w[3][21] , \w[3][20] , \w[3][19] , 
        \w[3][18] , \w[3][17] , \w[3][16] , \w[3][15] , \w[3][14] , \w[3][13] , 
        \w[3][12] , \w[3][11] , \w[3][10] , \w[3][9] , \w[3][8] , \w[3][7] , 
        \w[3][6] , \w[3][5] , \w[3][4] , \w[3][3] , \w[3][2] , \w[3][1] , 1'b0}), .CI(1'b0), .S({\w[4][31] , \w[4][30] , \w[4][29] , \w[4][28] , \w[4][27] , 
        \w[4][26] , \w[4][25] , \w[4][24] , \w[4][23] , \w[4][22] , \w[4][21] , 
        \w[4][20] , \w[4][19] , \w[4][18] , \w[4][17] , \w[4][16] , \w[4][15] , 
        \w[4][14] , \w[4][13] , \w[4][12] , \w[4][11] , \w[4][10] , \w[4][9] , 
        \w[4][8] , \w[4][7] , \w[4][6] , \w[4][5] , \w[4][4] , \w[4][3] , 
        \w[4][2] , \w[4][1] , SYNOPSYS_UNCONNECTED__2}) );
  ADD_N32_124 \FAINST[4].ADD_  ( .A({\_6_net_[31] , \_6_net_[30] , 
        \_6_net_[29] , \_6_net_[28] , \_6_net_[27] , \_6_net_[26] , 
        \_6_net_[25] , \_6_net_[24] , \_6_net_[23] , \_6_net_[22] , 
        \_6_net_[21] , \_6_net_[20] , \_6_net_[19] , \_6_net_[18] , 
        \_6_net_[17] , \_6_net_[16] , \_6_net_[15] , \_6_net_[14] , 
        \_6_net_[13] , \_6_net_[12] , \_6_net_[11] , \_6_net_[10] , 
        \_6_net_[9] , \_6_net_[8] , \_6_net_[7] , \_6_net_[6] , \_6_net_[5] , 
        \_6_net_[4] , 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[4][31] , \w[4][30] , 
        \w[4][29] , \w[4][28] , \w[4][27] , \w[4][26] , \w[4][25] , \w[4][24] , 
        \w[4][23] , \w[4][22] , \w[4][21] , \w[4][20] , \w[4][19] , \w[4][18] , 
        \w[4][17] , \w[4][16] , \w[4][15] , \w[4][14] , \w[4][13] , \w[4][12] , 
        \w[4][11] , \w[4][10] , \w[4][9] , \w[4][8] , \w[4][7] , \w[4][6] , 
        \w[4][5] , \w[4][4] , \w[4][3] , \w[4][2] , \w[4][1] , 1'b0}), .CI(
        1'b0), .S({\w[5][31] , \w[5][30] , \w[5][29] , \w[5][28] , \w[5][27] , 
        \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , \w[5][22] , \w[5][21] , 
        \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , \w[5][16] , \w[5][15] , 
        \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , \w[5][10] , \w[5][9] , 
        \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , \w[5][4] , \w[5][3] , 
        \w[5][2] , \w[5][1] , SYNOPSYS_UNCONNECTED__3}) );
  ADD_N32_123 \FAINST[5].ADD_  ( .A({\_8_net_[31] , \_8_net_[30] , 
        \_8_net_[29] , \_8_net_[28] , \_8_net_[27] , \_8_net_[26] , 
        \_8_net_[25] , \_8_net_[24] , \_8_net_[23] , \_8_net_[22] , 
        \_8_net_[21] , \_8_net_[20] , \_8_net_[19] , \_8_net_[18] , 
        \_8_net_[17] , \_8_net_[16] , \_8_net_[15] , \_8_net_[14] , 
        \_8_net_[13] , \_8_net_[12] , \_8_net_[11] , \_8_net_[10] , 
        \_8_net_[9] , \_8_net_[8] , \_8_net_[7] , \_8_net_[6] , \_8_net_[5] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[5][31] , \w[5][30] , \w[5][29] , 
        \w[5][28] , \w[5][27] , \w[5][26] , \w[5][25] , \w[5][24] , \w[5][23] , 
        \w[5][22] , \w[5][21] , \w[5][20] , \w[5][19] , \w[5][18] , \w[5][17] , 
        \w[5][16] , \w[5][15] , \w[5][14] , \w[5][13] , \w[5][12] , \w[5][11] , 
        \w[5][10] , \w[5][9] , \w[5][8] , \w[5][7] , \w[5][6] , \w[5][5] , 
        \w[5][4] , \w[5][3] , \w[5][2] , \w[5][1] , 1'b0}), .CI(1'b0), .S({
        \w[6][31] , \w[6][30] , \w[6][29] , \w[6][28] , \w[6][27] , \w[6][26] , 
        \w[6][25] , \w[6][24] , \w[6][23] , \w[6][22] , \w[6][21] , \w[6][20] , 
        \w[6][19] , \w[6][18] , \w[6][17] , \w[6][16] , \w[6][15] , \w[6][14] , 
        \w[6][13] , \w[6][12] , \w[6][11] , \w[6][10] , \w[6][9] , \w[6][8] , 
        \w[6][7] , \w[6][6] , \w[6][5] , \w[6][4] , \w[6][3] , \w[6][2] , 
        \w[6][1] , SYNOPSYS_UNCONNECTED__4}) );
  ADD_N32_122 \FAINST[6].ADD_  ( .A({\_10_net_[31] , \_10_net_[30] , 
        \_10_net_[29] , \_10_net_[28] , \_10_net_[27] , \_10_net_[26] , 
        \_10_net_[25] , \_10_net_[24] , \_10_net_[23] , \_10_net_[22] , 
        \_10_net_[21] , \_10_net_[20] , \_10_net_[19] , \_10_net_[18] , 
        \_10_net_[17] , \_10_net_[16] , \_10_net_[15] , \_10_net_[14] , 
        \_10_net_[13] , \_10_net_[12] , \_10_net_[11] , \_10_net_[10] , 
        \_10_net_[9] , \_10_net_[8] , \_10_net_[7] , \_10_net_[6] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[6][31] , \w[6][30] , \w[6][29] , 
        \w[6][28] , \w[6][27] , \w[6][26] , \w[6][25] , \w[6][24] , \w[6][23] , 
        \w[6][22] , \w[6][21] , \w[6][20] , \w[6][19] , \w[6][18] , \w[6][17] , 
        \w[6][16] , \w[6][15] , \w[6][14] , \w[6][13] , \w[6][12] , \w[6][11] , 
        \w[6][10] , \w[6][9] , \w[6][8] , \w[6][7] , \w[6][6] , \w[6][5] , 
        \w[6][4] , \w[6][3] , \w[6][2] , \w[6][1] , 1'b0}), .CI(1'b0), .S({
        \w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , \w[7][27] , \w[7][26] , 
        \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , \w[7][21] , \w[7][20] , 
        \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , \w[7][15] , \w[7][14] , 
        \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , \w[7][9] , \w[7][8] , 
        \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , \w[7][3] , \w[7][2] , 
        \w[7][1] , SYNOPSYS_UNCONNECTED__5}) );
  ADD_N32_121 \FAINST[7].ADD_  ( .A({\_12_net_[31] , \_12_net_[30] , 
        \_12_net_[29] , \_12_net_[28] , \_12_net_[27] , \_12_net_[26] , 
        \_12_net_[25] , \_12_net_[24] , \_12_net_[23] , \_12_net_[22] , 
        \_12_net_[21] , \_12_net_[20] , \_12_net_[19] , \_12_net_[18] , 
        \_12_net_[17] , \_12_net_[16] , \_12_net_[15] , \_12_net_[14] , 
        \_12_net_[13] , \_12_net_[12] , \_12_net_[11] , \_12_net_[10] , 
        \_12_net_[9] , \_12_net_[8] , \_12_net_[7] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[7][31] , \w[7][30] , \w[7][29] , \w[7][28] , 
        \w[7][27] , \w[7][26] , \w[7][25] , \w[7][24] , \w[7][23] , \w[7][22] , 
        \w[7][21] , \w[7][20] , \w[7][19] , \w[7][18] , \w[7][17] , \w[7][16] , 
        \w[7][15] , \w[7][14] , \w[7][13] , \w[7][12] , \w[7][11] , \w[7][10] , 
        \w[7][9] , \w[7][8] , \w[7][7] , \w[7][6] , \w[7][5] , \w[7][4] , 
        \w[7][3] , \w[7][2] , \w[7][1] , 1'b0}), .CI(1'b0), .S({\w[8][31] , 
        \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , \w[8][26] , \w[8][25] , 
        \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , \w[8][20] , \w[8][19] , 
        \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , \w[8][14] , \w[8][13] , 
        \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , \w[8][8] , \w[8][7] , 
        \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , \w[8][2] , \w[8][1] , 
        SYNOPSYS_UNCONNECTED__6}) );
  ADD_N32_120 \FAINST[8].ADD_  ( .A({\_14_net_[31] , \_14_net_[30] , 
        \_14_net_[29] , \_14_net_[28] , \_14_net_[27] , \_14_net_[26] , 
        \_14_net_[25] , \_14_net_[24] , \_14_net_[23] , \_14_net_[22] , 
        \_14_net_[21] , \_14_net_[20] , \_14_net_[19] , \_14_net_[18] , 
        \_14_net_[17] , \_14_net_[16] , \_14_net_[15] , \_14_net_[14] , 
        \_14_net_[13] , \_14_net_[12] , \_14_net_[11] , \_14_net_[10] , 
        \_14_net_[9] , \_14_net_[8] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[8][31] , \w[8][30] , \w[8][29] , \w[8][28] , \w[8][27] , 
        \w[8][26] , \w[8][25] , \w[8][24] , \w[8][23] , \w[8][22] , \w[8][21] , 
        \w[8][20] , \w[8][19] , \w[8][18] , \w[8][17] , \w[8][16] , \w[8][15] , 
        \w[8][14] , \w[8][13] , \w[8][12] , \w[8][11] , \w[8][10] , \w[8][9] , 
        \w[8][8] , \w[8][7] , \w[8][6] , \w[8][5] , \w[8][4] , \w[8][3] , 
        \w[8][2] , \w[8][1] , 1'b0}), .CI(1'b0), .S({\w[9][31] , \w[9][30] , 
        \w[9][29] , \w[9][28] , \w[9][27] , \w[9][26] , \w[9][25] , \w[9][24] , 
        \w[9][23] , \w[9][22] , \w[9][21] , \w[9][20] , \w[9][19] , \w[9][18] , 
        \w[9][17] , \w[9][16] , \w[9][15] , \w[9][14] , \w[9][13] , \w[9][12] , 
        \w[9][11] , \w[9][10] , \w[9][9] , \w[9][8] , \w[9][7] , \w[9][6] , 
        \w[9][5] , \w[9][4] , \w[9][3] , \w[9][2] , \w[9][1] , 
        SYNOPSYS_UNCONNECTED__7}) );
  ADD_N32_119 \FAINST[9].ADD_  ( .A({\_16_net_[31] , \_16_net_[30] , 
        \_16_net_[29] , \_16_net_[28] , \_16_net_[27] , \_16_net_[26] , 
        \_16_net_[25] , \_16_net_[24] , \_16_net_[23] , \_16_net_[22] , 
        \_16_net_[21] , \_16_net_[20] , \_16_net_[19] , \_16_net_[18] , 
        \_16_net_[17] , \_16_net_[16] , \_16_net_[15] , \_16_net_[14] , 
        \_16_net_[13] , \_16_net_[12] , \_16_net_[11] , \_16_net_[10] , 
        \_16_net_[9] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[9][31] , \w[9][30] , \w[9][29] , \w[9][28] , \w[9][27] , 
        \w[9][26] , \w[9][25] , \w[9][24] , \w[9][23] , \w[9][22] , \w[9][21] , 
        \w[9][20] , \w[9][19] , \w[9][18] , \w[9][17] , \w[9][16] , \w[9][15] , 
        \w[9][14] , \w[9][13] , \w[9][12] , \w[9][11] , \w[9][10] , \w[9][9] , 
        \w[9][8] , \w[9][7] , \w[9][6] , \w[9][5] , \w[9][4] , \w[9][3] , 
        \w[9][2] , \w[9][1] , 1'b0}), .CI(1'b0), .S({\w[10][31] , \w[10][30] , 
        \w[10][29] , \w[10][28] , \w[10][27] , \w[10][26] , \w[10][25] , 
        \w[10][24] , \w[10][23] , \w[10][22] , \w[10][21] , \w[10][20] , 
        \w[10][19] , \w[10][18] , \w[10][17] , \w[10][16] , \w[10][15] , 
        \w[10][14] , \w[10][13] , \w[10][12] , \w[10][11] , \w[10][10] , 
        \w[10][9] , \w[10][8] , \w[10][7] , \w[10][6] , \w[10][5] , \w[10][4] , 
        \w[10][3] , \w[10][2] , \w[10][1] , SYNOPSYS_UNCONNECTED__8}) );
  ADD_N32_118 \FAINST[10].ADD_  ( .A({\_18_net_[31] , \_18_net_[30] , 
        \_18_net_[29] , \_18_net_[28] , \_18_net_[27] , \_18_net_[26] , 
        \_18_net_[25] , \_18_net_[24] , \_18_net_[23] , \_18_net_[22] , 
        \_18_net_[21] , \_18_net_[20] , \_18_net_[19] , \_18_net_[18] , 
        \_18_net_[17] , \_18_net_[16] , \_18_net_[15] , \_18_net_[14] , 
        \_18_net_[13] , \_18_net_[12] , \_18_net_[11] , \_18_net_[10] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[10][31] , \w[10][30] , \w[10][29] , \w[10][28] , \w[10][27] , 
        \w[10][26] , \w[10][25] , \w[10][24] , \w[10][23] , \w[10][22] , 
        \w[10][21] , \w[10][20] , \w[10][19] , \w[10][18] , \w[10][17] , 
        \w[10][16] , \w[10][15] , \w[10][14] , \w[10][13] , \w[10][12] , 
        \w[10][11] , \w[10][10] , \w[10][9] , \w[10][8] , \w[10][7] , 
        \w[10][6] , \w[10][5] , \w[10][4] , \w[10][3] , \w[10][2] , \w[10][1] , 
        1'b0}), .CI(1'b0), .S({\w[11][31] , \w[11][30] , \w[11][29] , 
        \w[11][28] , \w[11][27] , \w[11][26] , \w[11][25] , \w[11][24] , 
        \w[11][23] , \w[11][22] , \w[11][21] , \w[11][20] , \w[11][19] , 
        \w[11][18] , \w[11][17] , \w[11][16] , \w[11][15] , \w[11][14] , 
        \w[11][13] , \w[11][12] , \w[11][11] , \w[11][10] , \w[11][9] , 
        \w[11][8] , \w[11][7] , \w[11][6] , \w[11][5] , \w[11][4] , \w[11][3] , 
        \w[11][2] , \w[11][1] , SYNOPSYS_UNCONNECTED__9}) );
  ADD_N32_117 \FAINST[11].ADD_  ( .A({\_20_net_[31] , \_20_net_[30] , 
        \_20_net_[29] , \_20_net_[28] , \_20_net_[27] , \_20_net_[26] , 
        \_20_net_[25] , \_20_net_[24] , \_20_net_[23] , \_20_net_[22] , 
        \_20_net_[21] , \_20_net_[20] , \_20_net_[19] , \_20_net_[18] , 
        \_20_net_[17] , \_20_net_[16] , \_20_net_[15] , \_20_net_[14] , 
        \_20_net_[13] , \_20_net_[12] , \_20_net_[11] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[11][31] , 
        \w[11][30] , \w[11][29] , \w[11][28] , \w[11][27] , \w[11][26] , 
        \w[11][25] , \w[11][24] , \w[11][23] , \w[11][22] , \w[11][21] , 
        \w[11][20] , \w[11][19] , \w[11][18] , \w[11][17] , \w[11][16] , 
        \w[11][15] , \w[11][14] , \w[11][13] , \w[11][12] , \w[11][11] , 
        \w[11][10] , \w[11][9] , \w[11][8] , \w[11][7] , \w[11][6] , 
        \w[11][5] , \w[11][4] , \w[11][3] , \w[11][2] , \w[11][1] , 1'b0}), 
        .CI(1'b0), .S({\w[12][31] , \w[12][30] , \w[12][29] , \w[12][28] , 
        \w[12][27] , \w[12][26] , \w[12][25] , \w[12][24] , \w[12][23] , 
        \w[12][22] , \w[12][21] , \w[12][20] , \w[12][19] , \w[12][18] , 
        \w[12][17] , \w[12][16] , \w[12][15] , \w[12][14] , \w[12][13] , 
        \w[12][12] , \w[12][11] , \w[12][10] , \w[12][9] , \w[12][8] , 
        \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , \w[12][3] , \w[12][2] , 
        \w[12][1] , SYNOPSYS_UNCONNECTED__10}) );
  ADD_N32_116 \FAINST[12].ADD_  ( .A({\_22_net_[31] , \_22_net_[30] , 
        \_22_net_[29] , \_22_net_[28] , \_22_net_[27] , \_22_net_[26] , 
        \_22_net_[25] , \_22_net_[24] , \_22_net_[23] , \_22_net_[22] , 
        \_22_net_[21] , \_22_net_[20] , \_22_net_[19] , \_22_net_[18] , 
        \_22_net_[17] , \_22_net_[16] , \_22_net_[15] , \_22_net_[14] , 
        \_22_net_[13] , \_22_net_[12] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[12][31] , \w[12][30] , 
        \w[12][29] , \w[12][28] , \w[12][27] , \w[12][26] , \w[12][25] , 
        \w[12][24] , \w[12][23] , \w[12][22] , \w[12][21] , \w[12][20] , 
        \w[12][19] , \w[12][18] , \w[12][17] , \w[12][16] , \w[12][15] , 
        \w[12][14] , \w[12][13] , \w[12][12] , \w[12][11] , \w[12][10] , 
        \w[12][9] , \w[12][8] , \w[12][7] , \w[12][6] , \w[12][5] , \w[12][4] , 
        \w[12][3] , \w[12][2] , \w[12][1] , 1'b0}), .CI(1'b0), .S({\w[13][31] , 
        \w[13][30] , \w[13][29] , \w[13][28] , \w[13][27] , \w[13][26] , 
        \w[13][25] , \w[13][24] , \w[13][23] , \w[13][22] , \w[13][21] , 
        \w[13][20] , \w[13][19] , \w[13][18] , \w[13][17] , \w[13][16] , 
        \w[13][15] , \w[13][14] , \w[13][13] , \w[13][12] , \w[13][11] , 
        \w[13][10] , \w[13][9] , \w[13][8] , \w[13][7] , \w[13][6] , 
        \w[13][5] , \w[13][4] , \w[13][3] , \w[13][2] , \w[13][1] , 
        SYNOPSYS_UNCONNECTED__11}) );
  ADD_N32_115 \FAINST[13].ADD_  ( .A({\_24_net_[31] , \_24_net_[30] , 
        \_24_net_[29] , \_24_net_[28] , \_24_net_[27] , \_24_net_[26] , 
        \_24_net_[25] , \_24_net_[24] , \_24_net_[23] , \_24_net_[22] , 
        \_24_net_[21] , \_24_net_[20] , \_24_net_[19] , \_24_net_[18] , 
        \_24_net_[17] , \_24_net_[16] , \_24_net_[15] , \_24_net_[14] , 
        \_24_net_[13] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[13][31] , \w[13][30] , \w[13][29] , 
        \w[13][28] , \w[13][27] , \w[13][26] , \w[13][25] , \w[13][24] , 
        \w[13][23] , \w[13][22] , \w[13][21] , \w[13][20] , \w[13][19] , 
        \w[13][18] , \w[13][17] , \w[13][16] , \w[13][15] , \w[13][14] , 
        \w[13][13] , \w[13][12] , \w[13][11] , \w[13][10] , \w[13][9] , 
        \w[13][8] , \w[13][7] , \w[13][6] , \w[13][5] , \w[13][4] , \w[13][3] , 
        \w[13][2] , \w[13][1] , 1'b0}), .CI(1'b0), .S({\w[14][31] , 
        \w[14][30] , \w[14][29] , \w[14][28] , \w[14][27] , \w[14][26] , 
        \w[14][25] , \w[14][24] , \w[14][23] , \w[14][22] , \w[14][21] , 
        \w[14][20] , \w[14][19] , \w[14][18] , \w[14][17] , \w[14][16] , 
        \w[14][15] , \w[14][14] , \w[14][13] , \w[14][12] , \w[14][11] , 
        \w[14][10] , \w[14][9] , \w[14][8] , \w[14][7] , \w[14][6] , 
        \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , \w[14][1] , 
        SYNOPSYS_UNCONNECTED__12}) );
  ADD_N32_114 \FAINST[14].ADD_  ( .A({\_26_net_[31] , \_26_net_[30] , 
        \_26_net_[29] , \_26_net_[28] , \_26_net_[27] , \_26_net_[26] , 
        \_26_net_[25] , \_26_net_[24] , \_26_net_[23] , \_26_net_[22] , 
        \_26_net_[21] , \_26_net_[20] , \_26_net_[19] , \_26_net_[18] , 
        \_26_net_[17] , \_26_net_[16] , \_26_net_[15] , \_26_net_[14] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[14][31] , \w[14][30] , \w[14][29] , \w[14][28] , 
        \w[14][27] , \w[14][26] , \w[14][25] , \w[14][24] , \w[14][23] , 
        \w[14][22] , \w[14][21] , \w[14][20] , \w[14][19] , \w[14][18] , 
        \w[14][17] , \w[14][16] , \w[14][15] , \w[14][14] , \w[14][13] , 
        \w[14][12] , \w[14][11] , \w[14][10] , \w[14][9] , \w[14][8] , 
        \w[14][7] , \w[14][6] , \w[14][5] , \w[14][4] , \w[14][3] , \w[14][2] , 
        \w[14][1] , 1'b0}), .CI(1'b0), .S({\w[15][31] , \w[15][30] , 
        \w[15][29] , \w[15][28] , \w[15][27] , \w[15][26] , \w[15][25] , 
        \w[15][24] , \w[15][23] , \w[15][22] , \w[15][21] , \w[15][20] , 
        \w[15][19] , \w[15][18] , \w[15][17] , \w[15][16] , \w[15][15] , 
        \w[15][14] , \w[15][13] , \w[15][12] , \w[15][11] , \w[15][10] , 
        \w[15][9] , \w[15][8] , \w[15][7] , \w[15][6] , \w[15][5] , \w[15][4] , 
        \w[15][3] , \w[15][2] , \w[15][1] , SYNOPSYS_UNCONNECTED__13}) );
  ADD_N32_113 \FAINST[15].ADD_  ( .A({\_28_net_[31] , \_28_net_[30] , 
        \_28_net_[29] , \_28_net_[28] , \_28_net_[27] , \_28_net_[26] , 
        \_28_net_[25] , \_28_net_[24] , \_28_net_[23] , \_28_net_[22] , 
        \_28_net_[21] , \_28_net_[20] , \_28_net_[19] , \_28_net_[18] , 
        \_28_net_[17] , \_28_net_[16] , \_28_net_[15] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[15][31] , \w[15][30] , \w[15][29] , \w[15][28] , \w[15][27] , 
        \w[15][26] , \w[15][25] , \w[15][24] , \w[15][23] , \w[15][22] , 
        \w[15][21] , \w[15][20] , \w[15][19] , \w[15][18] , \w[15][17] , 
        \w[15][16] , \w[15][15] , \w[15][14] , \w[15][13] , \w[15][12] , 
        \w[15][11] , \w[15][10] , \w[15][9] , \w[15][8] , \w[15][7] , 
        \w[15][6] , \w[15][5] , \w[15][4] , \w[15][3] , \w[15][2] , \w[15][1] , 
        1'b0}), .CI(1'b0), .S({\w[16][31] , \w[16][30] , \w[16][29] , 
        \w[16][28] , \w[16][27] , \w[16][26] , \w[16][25] , \w[16][24] , 
        \w[16][23] , \w[16][22] , \w[16][21] , \w[16][20] , \w[16][19] , 
        \w[16][18] , \w[16][17] , \w[16][16] , \w[16][15] , \w[16][14] , 
        \w[16][13] , \w[16][12] , \w[16][11] , \w[16][10] , \w[16][9] , 
        \w[16][8] , \w[16][7] , \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , 
        \w[16][2] , \w[16][1] , SYNOPSYS_UNCONNECTED__14}) );
  ADD_N32_112 \FAINST[16].ADD_  ( .A({\_30_net_[31] , \_30_net_[30] , 
        \_30_net_[29] , \_30_net_[28] , \_30_net_[27] , \_30_net_[26] , 
        \_30_net_[25] , \_30_net_[24] , \_30_net_[23] , \_30_net_[22] , 
        \_30_net_[21] , \_30_net_[20] , \_30_net_[19] , \_30_net_[18] , 
        \_30_net_[17] , \_30_net_[16] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[16][31] , \w[16][30] , \w[16][29] , \w[16][28] , \w[16][27] , 
        \w[16][26] , \w[16][25] , \w[16][24] , \w[16][23] , \w[16][22] , 
        \w[16][21] , \w[16][20] , \w[16][19] , \w[16][18] , \w[16][17] , 
        \w[16][16] , \w[16][15] , \w[16][14] , \w[16][13] , \w[16][12] , 
        \w[16][11] , \w[16][10] , \w[16][9] , \w[16][8] , \w[16][7] , 
        \w[16][6] , \w[16][5] , \w[16][4] , \w[16][3] , \w[16][2] , \w[16][1] , 
        1'b0}), .CI(1'b0), .S({\w[17][31] , \w[17][30] , \w[17][29] , 
        \w[17][28] , \w[17][27] , \w[17][26] , \w[17][25] , \w[17][24] , 
        \w[17][23] , \w[17][22] , \w[17][21] , \w[17][20] , \w[17][19] , 
        \w[17][18] , \w[17][17] , \w[17][16] , \w[17][15] , \w[17][14] , 
        \w[17][13] , \w[17][12] , \w[17][11] , \w[17][10] , \w[17][9] , 
        \w[17][8] , \w[17][7] , \w[17][6] , \w[17][5] , \w[17][4] , \w[17][3] , 
        \w[17][2] , \w[17][1] , SYNOPSYS_UNCONNECTED__15}) );
  ADD_N32_111 \FAINST[17].ADD_  ( .A({\_32_net_[31] , \_32_net_[30] , 
        \_32_net_[29] , \_32_net_[28] , \_32_net_[27] , \_32_net_[26] , 
        \_32_net_[25] , \_32_net_[24] , \_32_net_[23] , \_32_net_[22] , 
        \_32_net_[21] , \_32_net_[20] , \_32_net_[19] , \_32_net_[18] , 
        \_32_net_[17] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[17][31] , 
        \w[17][30] , \w[17][29] , \w[17][28] , \w[17][27] , \w[17][26] , 
        \w[17][25] , \w[17][24] , \w[17][23] , \w[17][22] , \w[17][21] , 
        \w[17][20] , \w[17][19] , \w[17][18] , \w[17][17] , \w[17][16] , 
        \w[17][15] , \w[17][14] , \w[17][13] , \w[17][12] , \w[17][11] , 
        \w[17][10] , \w[17][9] , \w[17][8] , \w[17][7] , \w[17][6] , 
        \w[17][5] , \w[17][4] , \w[17][3] , \w[17][2] , \w[17][1] , 1'b0}), 
        .CI(1'b0), .S({\w[18][31] , \w[18][30] , \w[18][29] , \w[18][28] , 
        \w[18][27] , \w[18][26] , \w[18][25] , \w[18][24] , \w[18][23] , 
        \w[18][22] , \w[18][21] , \w[18][20] , \w[18][19] , \w[18][18] , 
        \w[18][17] , \w[18][16] , \w[18][15] , \w[18][14] , \w[18][13] , 
        \w[18][12] , \w[18][11] , \w[18][10] , \w[18][9] , \w[18][8] , 
        \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , \w[18][3] , \w[18][2] , 
        \w[18][1] , SYNOPSYS_UNCONNECTED__16}) );
  ADD_N32_110 \FAINST[18].ADD_  ( .A({\_34_net_[31] , \_34_net_[30] , 
        \_34_net_[29] , \_34_net_[28] , \_34_net_[27] , \_34_net_[26] , 
        \_34_net_[25] , \_34_net_[24] , \_34_net_[23] , \_34_net_[22] , 
        \_34_net_[21] , \_34_net_[20] , \_34_net_[19] , \_34_net_[18] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[18][31] , \w[18][30] , 
        \w[18][29] , \w[18][28] , \w[18][27] , \w[18][26] , \w[18][25] , 
        \w[18][24] , \w[18][23] , \w[18][22] , \w[18][21] , \w[18][20] , 
        \w[18][19] , \w[18][18] , \w[18][17] , \w[18][16] , \w[18][15] , 
        \w[18][14] , \w[18][13] , \w[18][12] , \w[18][11] , \w[18][10] , 
        \w[18][9] , \w[18][8] , \w[18][7] , \w[18][6] , \w[18][5] , \w[18][4] , 
        \w[18][3] , \w[18][2] , \w[18][1] , 1'b0}), .CI(1'b0), .S({\w[19][31] , 
        \w[19][30] , \w[19][29] , \w[19][28] , \w[19][27] , \w[19][26] , 
        \w[19][25] , \w[19][24] , \w[19][23] , \w[19][22] , \w[19][21] , 
        \w[19][20] , \w[19][19] , \w[19][18] , \w[19][17] , \w[19][16] , 
        \w[19][15] , \w[19][14] , \w[19][13] , \w[19][12] , \w[19][11] , 
        \w[19][10] , \w[19][9] , \w[19][8] , \w[19][7] , \w[19][6] , 
        \w[19][5] , \w[19][4] , \w[19][3] , \w[19][2] , \w[19][1] , 
        SYNOPSYS_UNCONNECTED__17}) );
  ADD_N32_109 \FAINST[19].ADD_  ( .A({\_36_net_[31] , \_36_net_[30] , 
        \_36_net_[29] , \_36_net_[28] , \_36_net_[27] , \_36_net_[26] , 
        \_36_net_[25] , \_36_net_[24] , \_36_net_[23] , \_36_net_[22] , 
        \_36_net_[21] , \_36_net_[20] , \_36_net_[19] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[19][31] , \w[19][30] , \w[19][29] , 
        \w[19][28] , \w[19][27] , \w[19][26] , \w[19][25] , \w[19][24] , 
        \w[19][23] , \w[19][22] , \w[19][21] , \w[19][20] , \w[19][19] , 
        \w[19][18] , \w[19][17] , \w[19][16] , \w[19][15] , \w[19][14] , 
        \w[19][13] , \w[19][12] , \w[19][11] , \w[19][10] , \w[19][9] , 
        \w[19][8] , \w[19][7] , \w[19][6] , \w[19][5] , \w[19][4] , \w[19][3] , 
        \w[19][2] , \w[19][1] , 1'b0}), .CI(1'b0), .S({\w[20][31] , 
        \w[20][30] , \w[20][29] , \w[20][28] , \w[20][27] , \w[20][26] , 
        \w[20][25] , \w[20][24] , \w[20][23] , \w[20][22] , \w[20][21] , 
        \w[20][20] , \w[20][19] , \w[20][18] , \w[20][17] , \w[20][16] , 
        \w[20][15] , \w[20][14] , \w[20][13] , \w[20][12] , \w[20][11] , 
        \w[20][10] , \w[20][9] , \w[20][8] , \w[20][7] , \w[20][6] , 
        \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , \w[20][1] , 
        SYNOPSYS_UNCONNECTED__18}) );
  ADD_N32_108 \FAINST[20].ADD_  ( .A({\_38_net_[31] , \_38_net_[30] , 
        \_38_net_[29] , \_38_net_[28] , \_38_net_[27] , \_38_net_[26] , 
        \_38_net_[25] , \_38_net_[24] , \_38_net_[23] , \_38_net_[22] , 
        \_38_net_[21] , \_38_net_[20] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({\w[20][31] , \w[20][30] , \w[20][29] , \w[20][28] , 
        \w[20][27] , \w[20][26] , \w[20][25] , \w[20][24] , \w[20][23] , 
        \w[20][22] , \w[20][21] , \w[20][20] , \w[20][19] , \w[20][18] , 
        \w[20][17] , \w[20][16] , \w[20][15] , \w[20][14] , \w[20][13] , 
        \w[20][12] , \w[20][11] , \w[20][10] , \w[20][9] , \w[20][8] , 
        \w[20][7] , \w[20][6] , \w[20][5] , \w[20][4] , \w[20][3] , \w[20][2] , 
        \w[20][1] , 1'b0}), .CI(1'b0), .S({\w[21][31] , \w[21][30] , 
        \w[21][29] , \w[21][28] , \w[21][27] , \w[21][26] , \w[21][25] , 
        \w[21][24] , \w[21][23] , \w[21][22] , \w[21][21] , \w[21][20] , 
        \w[21][19] , \w[21][18] , \w[21][17] , \w[21][16] , \w[21][15] , 
        \w[21][14] , \w[21][13] , \w[21][12] , \w[21][11] , \w[21][10] , 
        \w[21][9] , \w[21][8] , \w[21][7] , \w[21][6] , \w[21][5] , \w[21][4] , 
        \w[21][3] , \w[21][2] , \w[21][1] , SYNOPSYS_UNCONNECTED__19}) );
  ADD_N32_107 \FAINST[21].ADD_  ( .A({\_40_net_[31] , \_40_net_[30] , 
        \_40_net_[29] , \_40_net_[28] , \_40_net_[27] , \_40_net_[26] , 
        \_40_net_[25] , \_40_net_[24] , \_40_net_[23] , \_40_net_[22] , 
        \_40_net_[21] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[21][31] , \w[21][30] , \w[21][29] , \w[21][28] , \w[21][27] , 
        \w[21][26] , \w[21][25] , \w[21][24] , \w[21][23] , \w[21][22] , 
        \w[21][21] , \w[21][20] , \w[21][19] , \w[21][18] , \w[21][17] , 
        \w[21][16] , \w[21][15] , \w[21][14] , \w[21][13] , \w[21][12] , 
        \w[21][11] , \w[21][10] , \w[21][9] , \w[21][8] , \w[21][7] , 
        \w[21][6] , \w[21][5] , \w[21][4] , \w[21][3] , \w[21][2] , \w[21][1] , 
        1'b0}), .CI(1'b0), .S({\w[22][31] , \w[22][30] , \w[22][29] , 
        \w[22][28] , \w[22][27] , \w[22][26] , \w[22][25] , \w[22][24] , 
        \w[22][23] , \w[22][22] , \w[22][21] , \w[22][20] , \w[22][19] , 
        \w[22][18] , \w[22][17] , \w[22][16] , \w[22][15] , \w[22][14] , 
        \w[22][13] , \w[22][12] , \w[22][11] , \w[22][10] , \w[22][9] , 
        \w[22][8] , \w[22][7] , \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , 
        \w[22][2] , \w[22][1] , SYNOPSYS_UNCONNECTED__20}) );
  ADD_N32_106 \FAINST[22].ADD_  ( .A({\_42_net_[31] , \_42_net_[30] , 
        \_42_net_[29] , \_42_net_[28] , \_42_net_[27] , \_42_net_[26] , 
        \_42_net_[25] , \_42_net_[24] , \_42_net_[23] , \_42_net_[22] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[22][31] , \w[22][30] , \w[22][29] , \w[22][28] , \w[22][27] , 
        \w[22][26] , \w[22][25] , \w[22][24] , \w[22][23] , \w[22][22] , 
        \w[22][21] , \w[22][20] , \w[22][19] , \w[22][18] , \w[22][17] , 
        \w[22][16] , \w[22][15] , \w[22][14] , \w[22][13] , \w[22][12] , 
        \w[22][11] , \w[22][10] , \w[22][9] , \w[22][8] , \w[22][7] , 
        \w[22][6] , \w[22][5] , \w[22][4] , \w[22][3] , \w[22][2] , \w[22][1] , 
        1'b0}), .CI(1'b0), .S({\w[23][31] , \w[23][30] , \w[23][29] , 
        \w[23][28] , \w[23][27] , \w[23][26] , \w[23][25] , \w[23][24] , 
        \w[23][23] , \w[23][22] , \w[23][21] , \w[23][20] , \w[23][19] , 
        \w[23][18] , \w[23][17] , \w[23][16] , \w[23][15] , \w[23][14] , 
        \w[23][13] , \w[23][12] , \w[23][11] , \w[23][10] , \w[23][9] , 
        \w[23][8] , \w[23][7] , \w[23][6] , \w[23][5] , \w[23][4] , \w[23][3] , 
        \w[23][2] , \w[23][1] , SYNOPSYS_UNCONNECTED__21}) );
  ADD_N32_105 \FAINST[23].ADD_  ( .A({\_44_net_[31] , \_44_net_[30] , 
        \_44_net_[29] , \_44_net_[28] , \_44_net_[27] , \_44_net_[26] , 
        \_44_net_[25] , \_44_net_[24] , \_44_net_[23] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[23][31] , 
        \w[23][30] , \w[23][29] , \w[23][28] , \w[23][27] , \w[23][26] , 
        \w[23][25] , \w[23][24] , \w[23][23] , \w[23][22] , \w[23][21] , 
        \w[23][20] , \w[23][19] , \w[23][18] , \w[23][17] , \w[23][16] , 
        \w[23][15] , \w[23][14] , \w[23][13] , \w[23][12] , \w[23][11] , 
        \w[23][10] , \w[23][9] , \w[23][8] , \w[23][7] , \w[23][6] , 
        \w[23][5] , \w[23][4] , \w[23][3] , \w[23][2] , \w[23][1] , 1'b0}), 
        .CI(1'b0), .S({\w[24][31] , \w[24][30] , \w[24][29] , \w[24][28] , 
        \w[24][27] , \w[24][26] , \w[24][25] , \w[24][24] , \w[24][23] , 
        \w[24][22] , \w[24][21] , \w[24][20] , \w[24][19] , \w[24][18] , 
        \w[24][17] , \w[24][16] , \w[24][15] , \w[24][14] , \w[24][13] , 
        \w[24][12] , \w[24][11] , \w[24][10] , \w[24][9] , \w[24][8] , 
        \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , \w[24][3] , \w[24][2] , 
        \w[24][1] , SYNOPSYS_UNCONNECTED__22}) );
  ADD_N32_104 \FAINST[24].ADD_  ( .A({\_46_net_[31] , \_46_net_[30] , 
        \_46_net_[29] , \_46_net_[28] , \_46_net_[27] , \_46_net_[26] , 
        \_46_net_[25] , \_46_net_[24] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[24][31] , \w[24][30] , 
        \w[24][29] , \w[24][28] , \w[24][27] , \w[24][26] , \w[24][25] , 
        \w[24][24] , \w[24][23] , \w[24][22] , \w[24][21] , \w[24][20] , 
        \w[24][19] , \w[24][18] , \w[24][17] , \w[24][16] , \w[24][15] , 
        \w[24][14] , \w[24][13] , \w[24][12] , \w[24][11] , \w[24][10] , 
        \w[24][9] , \w[24][8] , \w[24][7] , \w[24][6] , \w[24][5] , \w[24][4] , 
        \w[24][3] , \w[24][2] , \w[24][1] , 1'b0}), .CI(1'b0), .S({\w[25][31] , 
        \w[25][30] , \w[25][29] , \w[25][28] , \w[25][27] , \w[25][26] , 
        \w[25][25] , \w[25][24] , \w[25][23] , \w[25][22] , \w[25][21] , 
        \w[25][20] , \w[25][19] , \w[25][18] , \w[25][17] , \w[25][16] , 
        \w[25][15] , \w[25][14] , \w[25][13] , \w[25][12] , \w[25][11] , 
        \w[25][10] , \w[25][9] , \w[25][8] , \w[25][7] , \w[25][6] , 
        \w[25][5] , \w[25][4] , \w[25][3] , \w[25][2] , \w[25][1] , 
        SYNOPSYS_UNCONNECTED__23}) );
  ADD_N32_103 \FAINST[25].ADD_  ( .A({\_48_net_[31] , \_48_net_[30] , 
        \_48_net_[29] , \_48_net_[28] , \_48_net_[27] , \_48_net_[26] , 
        \_48_net_[25] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[25][31] , \w[25][30] , \w[25][29] , 
        \w[25][28] , \w[25][27] , \w[25][26] , \w[25][25] , \w[25][24] , 
        \w[25][23] , \w[25][22] , \w[25][21] , \w[25][20] , \w[25][19] , 
        \w[25][18] , \w[25][17] , \w[25][16] , \w[25][15] , \w[25][14] , 
        \w[25][13] , \w[25][12] , \w[25][11] , \w[25][10] , \w[25][9] , 
        \w[25][8] , \w[25][7] , \w[25][6] , \w[25][5] , \w[25][4] , \w[25][3] , 
        \w[25][2] , \w[25][1] , 1'b0}), .CI(1'b0), .S({\w[26][31] , 
        \w[26][30] , \w[26][29] , \w[26][28] , \w[26][27] , \w[26][26] , 
        \w[26][25] , \w[26][24] , \w[26][23] , \w[26][22] , \w[26][21] , 
        \w[26][20] , \w[26][19] , \w[26][18] , \w[26][17] , \w[26][16] , 
        \w[26][15] , \w[26][14] , \w[26][13] , \w[26][12] , \w[26][11] , 
        \w[26][10] , \w[26][9] , \w[26][8] , \w[26][7] , \w[26][6] , 
        \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , \w[26][1] , 
        SYNOPSYS_UNCONNECTED__24}) );
  ADD_N32_102 \FAINST[26].ADD_  ( .A({\_50_net_[31] , \_50_net_[30] , 
        \_50_net_[29] , \_50_net_[28] , \_50_net_[27] , \_50_net_[26] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({\w[26][31] , \w[26][30] , \w[26][29] , \w[26][28] , 
        \w[26][27] , \w[26][26] , \w[26][25] , \w[26][24] , \w[26][23] , 
        \w[26][22] , \w[26][21] , \w[26][20] , \w[26][19] , \w[26][18] , 
        \w[26][17] , \w[26][16] , \w[26][15] , \w[26][14] , \w[26][13] , 
        \w[26][12] , \w[26][11] , \w[26][10] , \w[26][9] , \w[26][8] , 
        \w[26][7] , \w[26][6] , \w[26][5] , \w[26][4] , \w[26][3] , \w[26][2] , 
        \w[26][1] , 1'b0}), .CI(1'b0), .S({\w[27][31] , \w[27][30] , 
        \w[27][29] , \w[27][28] , \w[27][27] , \w[27][26] , \w[27][25] , 
        \w[27][24] , \w[27][23] , \w[27][22] , \w[27][21] , \w[27][20] , 
        \w[27][19] , \w[27][18] , \w[27][17] , \w[27][16] , \w[27][15] , 
        \w[27][14] , \w[27][13] , \w[27][12] , \w[27][11] , \w[27][10] , 
        \w[27][9] , \w[27][8] , \w[27][7] , \w[27][6] , \w[27][5] , \w[27][4] , 
        \w[27][3] , \w[27][2] , \w[27][1] , SYNOPSYS_UNCONNECTED__25}) );
  ADD_N32_101 \FAINST[27].ADD_  ( .A({\_52_net_[31] , \_52_net_[30] , 
        \_52_net_[29] , \_52_net_[28] , \_52_net_[27] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .B({\w[27][31] , \w[27][30] , \w[27][29] , \w[27][28] , \w[27][27] , 
        \w[27][26] , \w[27][25] , \w[27][24] , \w[27][23] , \w[27][22] , 
        \w[27][21] , \w[27][20] , \w[27][19] , \w[27][18] , \w[27][17] , 
        \w[27][16] , \w[27][15] , \w[27][14] , \w[27][13] , \w[27][12] , 
        \w[27][11] , \w[27][10] , \w[27][9] , \w[27][8] , \w[27][7] , 
        \w[27][6] , \w[27][5] , \w[27][4] , \w[27][3] , \w[27][2] , \w[27][1] , 
        1'b0}), .CI(1'b0), .S({\w[28][31] , \w[28][30] , \w[28][29] , 
        \w[28][28] , \w[28][27] , \w[28][26] , \w[28][25] , \w[28][24] , 
        \w[28][23] , \w[28][22] , \w[28][21] , \w[28][20] , \w[28][19] , 
        \w[28][18] , \w[28][17] , \w[28][16] , \w[28][15] , \w[28][14] , 
        \w[28][13] , \w[28][12] , \w[28][11] , \w[28][10] , \w[28][9] , 
        \w[28][8] , \w[28][7] , \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , 
        \w[28][2] , \w[28][1] , SYNOPSYS_UNCONNECTED__26}) );
  ADD_N32_100 \FAINST[28].ADD_  ( .A({\_54_net_[31] , \_54_net_[30] , 
        \_54_net_[29] , \_54_net_[28] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({
        \w[28][31] , \w[28][30] , \w[28][29] , \w[28][28] , \w[28][27] , 
        \w[28][26] , \w[28][25] , \w[28][24] , \w[28][23] , \w[28][22] , 
        \w[28][21] , \w[28][20] , \w[28][19] , \w[28][18] , \w[28][17] , 
        \w[28][16] , \w[28][15] , \w[28][14] , \w[28][13] , \w[28][12] , 
        \w[28][11] , \w[28][10] , \w[28][9] , \w[28][8] , \w[28][7] , 
        \w[28][6] , \w[28][5] , \w[28][4] , \w[28][3] , \w[28][2] , \w[28][1] , 
        1'b0}), .CI(1'b0), .S({\w[29][31] , \w[29][30] , \w[29][29] , 
        \w[29][28] , \w[29][27] , \w[29][26] , \w[29][25] , \w[29][24] , 
        \w[29][23] , \w[29][22] , \w[29][21] , \w[29][20] , \w[29][19] , 
        \w[29][18] , \w[29][17] , \w[29][16] , \w[29][15] , \w[29][14] , 
        \w[29][13] , \w[29][12] , \w[29][11] , \w[29][10] , \w[29][9] , 
        \w[29][8] , \w[29][7] , \w[29][6] , \w[29][5] , \w[29][4] , \w[29][3] , 
        \w[29][2] , \w[29][1] , SYNOPSYS_UNCONNECTED__27}) );
  ADD_N32_99 \FAINST[29].ADD_  ( .A({\_56_net_[31] , \_56_net_[30] , 
        \_56_net_[29] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[29][31] , 
        \w[29][30] , \w[29][29] , \w[29][28] , \w[29][27] , \w[29][26] , 
        \w[29][25] , \w[29][24] , \w[29][23] , \w[29][22] , \w[29][21] , 
        \w[29][20] , \w[29][19] , \w[29][18] , \w[29][17] , \w[29][16] , 
        \w[29][15] , \w[29][14] , \w[29][13] , \w[29][12] , \w[29][11] , 
        \w[29][10] , \w[29][9] , \w[29][8] , \w[29][7] , \w[29][6] , 
        \w[29][5] , \w[29][4] , \w[29][3] , \w[29][2] , \w[29][1] , 1'b0}), 
        .CI(1'b0), .S({\w[30][31] , \w[30][30] , \w[30][29] , \w[30][28] , 
        \w[30][27] , \w[30][26] , \w[30][25] , \w[30][24] , \w[30][23] , 
        \w[30][22] , \w[30][21] , \w[30][20] , \w[30][19] , \w[30][18] , 
        \w[30][17] , \w[30][16] , \w[30][15] , \w[30][14] , \w[30][13] , 
        \w[30][12] , \w[30][11] , \w[30][10] , \w[30][9] , \w[30][8] , 
        \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , \w[30][3] , \w[30][2] , 
        \w[30][1] , SYNOPSYS_UNCONNECTED__28}) );
  ADD_N32_98 \FAINST[30].ADD_  ( .A({\_58_net_[31] , \_58_net_[30] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({\w[30][31] , \w[30][30] , 
        \w[30][29] , \w[30][28] , \w[30][27] , \w[30][26] , \w[30][25] , 
        \w[30][24] , \w[30][23] , \w[30][22] , \w[30][21] , \w[30][20] , 
        \w[30][19] , \w[30][18] , \w[30][17] , \w[30][16] , \w[30][15] , 
        \w[30][14] , \w[30][13] , \w[30][12] , \w[30][11] , \w[30][10] , 
        \w[30][9] , \w[30][8] , \w[30][7] , \w[30][6] , \w[30][5] , \w[30][4] , 
        \w[30][3] , \w[30][2] , \w[30][1] , 1'b0}), .CI(1'b0), .S({\w[31][31] , 
        \w[31][30] , \w[31][29] , \w[31][28] , \w[31][27] , \w[31][26] , 
        \w[31][25] , \w[31][24] , \w[31][23] , \w[31][22] , \w[31][21] , 
        \w[31][20] , \w[31][19] , \w[31][18] , \w[31][17] , \w[31][16] , 
        \w[31][15] , \w[31][14] , \w[31][13] , \w[31][12] , \w[31][11] , 
        \w[31][10] , \w[31][9] , \w[31][8] , \w[31][7] , \w[31][6] , 
        \w[31][5] , \w[31][4] , \w[31][3] , \w[31][2] , \w[31][1] , 
        SYNOPSYS_UNCONNECTED__29}) );
  ADD_N32_97 \FAINST[31].ADD_  ( .A({\_60_net_[31] , 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({\w[31][31] , \w[31][30] , \w[31][29] , 
        \w[31][28] , \w[31][27] , \w[31][26] , \w[31][25] , \w[31][24] , 
        \w[31][23] , \w[31][22] , \w[31][21] , \w[31][20] , \w[31][19] , 
        \w[31][18] , \w[31][17] , \w[31][16] , \w[31][15] , \w[31][14] , 
        \w[31][13] , \w[31][12] , \w[31][11] , \w[31][10] , \w[31][9] , 
        \w[31][8] , \w[31][7] , \w[31][6] , \w[31][5] , \w[31][4] , \w[31][3] , 
        \w[31][2] , \w[31][1] , 1'b0}), .CI(1'b0), .S({O[31:1], 
        SYNOPSYS_UNCONNECTED__30}) );
  AND U2 ( .A(A[5]), .B(B[4]), .Z(\_8_net_[9] ) );
  AND U3 ( .A(A[5]), .B(B[3]), .Z(\_8_net_[8] ) );
  AND U4 ( .A(A[5]), .B(B[2]), .Z(\_8_net_[7] ) );
  AND U5 ( .A(A[5]), .B(B[1]), .Z(\_8_net_[6] ) );
  AND U6 ( .A(A[5]), .B(B[0]), .Z(\_8_net_[5] ) );
  AND U7 ( .A(A[5]), .B(B[26]), .Z(\_8_net_[31] ) );
  AND U8 ( .A(A[5]), .B(B[25]), .Z(\_8_net_[30] ) );
  AND U9 ( .A(A[5]), .B(B[24]), .Z(\_8_net_[29] ) );
  AND U10 ( .A(A[5]), .B(B[23]), .Z(\_8_net_[28] ) );
  AND U11 ( .A(A[5]), .B(B[22]), .Z(\_8_net_[27] ) );
  AND U12 ( .A(A[5]), .B(B[21]), .Z(\_8_net_[26] ) );
  AND U13 ( .A(A[5]), .B(B[20]), .Z(\_8_net_[25] ) );
  AND U14 ( .A(A[5]), .B(B[19]), .Z(\_8_net_[24] ) );
  AND U15 ( .A(A[5]), .B(B[18]), .Z(\_8_net_[23] ) );
  AND U16 ( .A(A[5]), .B(B[17]), .Z(\_8_net_[22] ) );
  AND U17 ( .A(A[5]), .B(B[16]), .Z(\_8_net_[21] ) );
  AND U18 ( .A(A[5]), .B(B[15]), .Z(\_8_net_[20] ) );
  AND U19 ( .A(A[5]), .B(B[14]), .Z(\_8_net_[19] ) );
  AND U20 ( .A(A[5]), .B(B[13]), .Z(\_8_net_[18] ) );
  AND U21 ( .A(A[5]), .B(B[12]), .Z(\_8_net_[17] ) );
  AND U22 ( .A(A[5]), .B(B[11]), .Z(\_8_net_[16] ) );
  AND U23 ( .A(A[5]), .B(B[10]), .Z(\_8_net_[15] ) );
  AND U24 ( .A(A[5]), .B(B[9]), .Z(\_8_net_[14] ) );
  AND U25 ( .A(A[5]), .B(B[8]), .Z(\_8_net_[13] ) );
  AND U26 ( .A(A[5]), .B(B[7]), .Z(\_8_net_[12] ) );
  AND U27 ( .A(A[5]), .B(B[6]), .Z(\_8_net_[11] ) );
  AND U28 ( .A(A[5]), .B(B[5]), .Z(\_8_net_[10] ) );
  AND U29 ( .A(B[5]), .B(A[4]), .Z(\_6_net_[9] ) );
  AND U30 ( .A(B[4]), .B(A[4]), .Z(\_6_net_[8] ) );
  AND U31 ( .A(B[3]), .B(A[4]), .Z(\_6_net_[7] ) );
  AND U32 ( .A(B[2]), .B(A[4]), .Z(\_6_net_[6] ) );
  AND U33 ( .A(B[1]), .B(A[4]), .Z(\_6_net_[5] ) );
  AND U34 ( .A(B[0]), .B(A[4]), .Z(\_6_net_[4] ) );
  AND U35 ( .A(A[4]), .B(B[27]), .Z(\_6_net_[31] ) );
  AND U36 ( .A(B[26]), .B(A[4]), .Z(\_6_net_[30] ) );
  AND U37 ( .A(B[25]), .B(A[4]), .Z(\_6_net_[29] ) );
  AND U38 ( .A(B[24]), .B(A[4]), .Z(\_6_net_[28] ) );
  AND U39 ( .A(B[23]), .B(A[4]), .Z(\_6_net_[27] ) );
  AND U40 ( .A(B[22]), .B(A[4]), .Z(\_6_net_[26] ) );
  AND U41 ( .A(B[21]), .B(A[4]), .Z(\_6_net_[25] ) );
  AND U42 ( .A(B[20]), .B(A[4]), .Z(\_6_net_[24] ) );
  AND U43 ( .A(B[19]), .B(A[4]), .Z(\_6_net_[23] ) );
  AND U44 ( .A(B[18]), .B(A[4]), .Z(\_6_net_[22] ) );
  AND U45 ( .A(B[17]), .B(A[4]), .Z(\_6_net_[21] ) );
  AND U46 ( .A(B[16]), .B(A[4]), .Z(\_6_net_[20] ) );
  AND U47 ( .A(B[15]), .B(A[4]), .Z(\_6_net_[19] ) );
  AND U48 ( .A(B[14]), .B(A[4]), .Z(\_6_net_[18] ) );
  AND U49 ( .A(B[13]), .B(A[4]), .Z(\_6_net_[17] ) );
  AND U50 ( .A(B[12]), .B(A[4]), .Z(\_6_net_[16] ) );
  AND U51 ( .A(B[11]), .B(A[4]), .Z(\_6_net_[15] ) );
  AND U52 ( .A(B[10]), .B(A[4]), .Z(\_6_net_[14] ) );
  AND U53 ( .A(B[9]), .B(A[4]), .Z(\_6_net_[13] ) );
  AND U54 ( .A(B[8]), .B(A[4]), .Z(\_6_net_[12] ) );
  AND U55 ( .A(B[7]), .B(A[4]), .Z(\_6_net_[11] ) );
  AND U56 ( .A(B[6]), .B(A[4]), .Z(\_6_net_[10] ) );
  AND U57 ( .A(A[31]), .B(B[0]), .Z(\_60_net_[31] ) );
  AND U58 ( .A(B[1]), .B(A[30]), .Z(\_58_net_[31] ) );
  AND U59 ( .A(A[30]), .B(B[0]), .Z(\_58_net_[30] ) );
  AND U60 ( .A(B[2]), .B(A[29]), .Z(\_56_net_[31] ) );
  AND U61 ( .A(B[1]), .B(A[29]), .Z(\_56_net_[30] ) );
  AND U62 ( .A(A[29]), .B(B[0]), .Z(\_56_net_[29] ) );
  AND U63 ( .A(B[3]), .B(A[28]), .Z(\_54_net_[31] ) );
  AND U64 ( .A(B[2]), .B(A[28]), .Z(\_54_net_[30] ) );
  AND U65 ( .A(B[1]), .B(A[28]), .Z(\_54_net_[29] ) );
  AND U66 ( .A(A[28]), .B(B[0]), .Z(\_54_net_[28] ) );
  AND U67 ( .A(B[4]), .B(A[27]), .Z(\_52_net_[31] ) );
  AND U68 ( .A(B[3]), .B(A[27]), .Z(\_52_net_[30] ) );
  AND U69 ( .A(B[2]), .B(A[27]), .Z(\_52_net_[29] ) );
  AND U70 ( .A(B[1]), .B(A[27]), .Z(\_52_net_[28] ) );
  AND U71 ( .A(A[27]), .B(B[0]), .Z(\_52_net_[27] ) );
  AND U72 ( .A(B[5]), .B(A[26]), .Z(\_50_net_[31] ) );
  AND U73 ( .A(B[4]), .B(A[26]), .Z(\_50_net_[30] ) );
  AND U74 ( .A(B[3]), .B(A[26]), .Z(\_50_net_[29] ) );
  AND U75 ( .A(B[2]), .B(A[26]), .Z(\_50_net_[28] ) );
  AND U76 ( .A(B[1]), .B(A[26]), .Z(\_50_net_[27] ) );
  AND U77 ( .A(A[26]), .B(B[0]), .Z(\_50_net_[26] ) );
  AND U78 ( .A(B[6]), .B(A[3]), .Z(\_4_net_[9] ) );
  AND U79 ( .A(B[5]), .B(A[3]), .Z(\_4_net_[8] ) );
  AND U80 ( .A(B[4]), .B(A[3]), .Z(\_4_net_[7] ) );
  AND U81 ( .A(B[3]), .B(A[3]), .Z(\_4_net_[6] ) );
  AND U82 ( .A(B[2]), .B(A[3]), .Z(\_4_net_[5] ) );
  AND U83 ( .A(B[1]), .B(A[3]), .Z(\_4_net_[4] ) );
  AND U84 ( .A(B[0]), .B(A[3]), .Z(\_4_net_[3] ) );
  AND U85 ( .A(A[3]), .B(B[28]), .Z(\_4_net_[31] ) );
  AND U86 ( .A(B[27]), .B(A[3]), .Z(\_4_net_[30] ) );
  AND U87 ( .A(B[26]), .B(A[3]), .Z(\_4_net_[29] ) );
  AND U88 ( .A(B[25]), .B(A[3]), .Z(\_4_net_[28] ) );
  AND U89 ( .A(B[24]), .B(A[3]), .Z(\_4_net_[27] ) );
  AND U90 ( .A(B[23]), .B(A[3]), .Z(\_4_net_[26] ) );
  AND U91 ( .A(B[22]), .B(A[3]), .Z(\_4_net_[25] ) );
  AND U92 ( .A(B[21]), .B(A[3]), .Z(\_4_net_[24] ) );
  AND U93 ( .A(B[20]), .B(A[3]), .Z(\_4_net_[23] ) );
  AND U94 ( .A(B[19]), .B(A[3]), .Z(\_4_net_[22] ) );
  AND U95 ( .A(B[18]), .B(A[3]), .Z(\_4_net_[21] ) );
  AND U96 ( .A(B[17]), .B(A[3]), .Z(\_4_net_[20] ) );
  AND U97 ( .A(B[16]), .B(A[3]), .Z(\_4_net_[19] ) );
  AND U98 ( .A(B[15]), .B(A[3]), .Z(\_4_net_[18] ) );
  AND U99 ( .A(B[14]), .B(A[3]), .Z(\_4_net_[17] ) );
  AND U100 ( .A(B[13]), .B(A[3]), .Z(\_4_net_[16] ) );
  AND U101 ( .A(B[12]), .B(A[3]), .Z(\_4_net_[15] ) );
  AND U102 ( .A(B[11]), .B(A[3]), .Z(\_4_net_[14] ) );
  AND U103 ( .A(B[10]), .B(A[3]), .Z(\_4_net_[13] ) );
  AND U104 ( .A(B[9]), .B(A[3]), .Z(\_4_net_[12] ) );
  AND U105 ( .A(B[8]), .B(A[3]), .Z(\_4_net_[11] ) );
  AND U106 ( .A(B[7]), .B(A[3]), .Z(\_4_net_[10] ) );
  AND U107 ( .A(B[6]), .B(A[25]), .Z(\_48_net_[31] ) );
  AND U108 ( .A(B[5]), .B(A[25]), .Z(\_48_net_[30] ) );
  AND U109 ( .A(B[4]), .B(A[25]), .Z(\_48_net_[29] ) );
  AND U110 ( .A(B[3]), .B(A[25]), .Z(\_48_net_[28] ) );
  AND U111 ( .A(B[2]), .B(A[25]), .Z(\_48_net_[27] ) );
  AND U112 ( .A(B[1]), .B(A[25]), .Z(\_48_net_[26] ) );
  AND U113 ( .A(A[25]), .B(B[0]), .Z(\_48_net_[25] ) );
  AND U114 ( .A(B[7]), .B(A[24]), .Z(\_46_net_[31] ) );
  AND U115 ( .A(B[6]), .B(A[24]), .Z(\_46_net_[30] ) );
  AND U116 ( .A(B[5]), .B(A[24]), .Z(\_46_net_[29] ) );
  AND U117 ( .A(B[4]), .B(A[24]), .Z(\_46_net_[28] ) );
  AND U118 ( .A(B[3]), .B(A[24]), .Z(\_46_net_[27] ) );
  AND U119 ( .A(B[2]), .B(A[24]), .Z(\_46_net_[26] ) );
  AND U120 ( .A(B[1]), .B(A[24]), .Z(\_46_net_[25] ) );
  AND U121 ( .A(A[24]), .B(B[0]), .Z(\_46_net_[24] ) );
  AND U122 ( .A(B[8]), .B(A[23]), .Z(\_44_net_[31] ) );
  AND U123 ( .A(B[7]), .B(A[23]), .Z(\_44_net_[30] ) );
  AND U124 ( .A(B[6]), .B(A[23]), .Z(\_44_net_[29] ) );
  AND U125 ( .A(B[5]), .B(A[23]), .Z(\_44_net_[28] ) );
  AND U126 ( .A(B[4]), .B(A[23]), .Z(\_44_net_[27] ) );
  AND U127 ( .A(B[3]), .B(A[23]), .Z(\_44_net_[26] ) );
  AND U128 ( .A(B[2]), .B(A[23]), .Z(\_44_net_[25] ) );
  AND U129 ( .A(B[1]), .B(A[23]), .Z(\_44_net_[24] ) );
  AND U130 ( .A(A[23]), .B(B[0]), .Z(\_44_net_[23] ) );
  AND U131 ( .A(B[9]), .B(A[22]), .Z(\_42_net_[31] ) );
  AND U132 ( .A(B[8]), .B(A[22]), .Z(\_42_net_[30] ) );
  AND U133 ( .A(B[7]), .B(A[22]), .Z(\_42_net_[29] ) );
  AND U134 ( .A(B[6]), .B(A[22]), .Z(\_42_net_[28] ) );
  AND U135 ( .A(B[5]), .B(A[22]), .Z(\_42_net_[27] ) );
  AND U136 ( .A(B[4]), .B(A[22]), .Z(\_42_net_[26] ) );
  AND U137 ( .A(B[3]), .B(A[22]), .Z(\_42_net_[25] ) );
  AND U138 ( .A(B[2]), .B(A[22]), .Z(\_42_net_[24] ) );
  AND U139 ( .A(B[1]), .B(A[22]), .Z(\_42_net_[23] ) );
  AND U140 ( .A(A[22]), .B(B[0]), .Z(\_42_net_[22] ) );
  AND U141 ( .A(B[10]), .B(A[21]), .Z(\_40_net_[31] ) );
  AND U142 ( .A(B[9]), .B(A[21]), .Z(\_40_net_[30] ) );
  AND U143 ( .A(B[8]), .B(A[21]), .Z(\_40_net_[29] ) );
  AND U144 ( .A(B[7]), .B(A[21]), .Z(\_40_net_[28] ) );
  AND U145 ( .A(B[6]), .B(A[21]), .Z(\_40_net_[27] ) );
  AND U146 ( .A(B[5]), .B(A[21]), .Z(\_40_net_[26] ) );
  AND U147 ( .A(B[4]), .B(A[21]), .Z(\_40_net_[25] ) );
  AND U148 ( .A(B[3]), .B(A[21]), .Z(\_40_net_[24] ) );
  AND U149 ( .A(B[2]), .B(A[21]), .Z(\_40_net_[23] ) );
  AND U150 ( .A(B[1]), .B(A[21]), .Z(\_40_net_[22] ) );
  AND U151 ( .A(A[21]), .B(B[0]), .Z(\_40_net_[21] ) );
  AND U152 ( .A(B[11]), .B(A[20]), .Z(\_38_net_[31] ) );
  AND U153 ( .A(B[10]), .B(A[20]), .Z(\_38_net_[30] ) );
  AND U154 ( .A(B[9]), .B(A[20]), .Z(\_38_net_[29] ) );
  AND U155 ( .A(B[8]), .B(A[20]), .Z(\_38_net_[28] ) );
  AND U156 ( .A(B[7]), .B(A[20]), .Z(\_38_net_[27] ) );
  AND U157 ( .A(B[6]), .B(A[20]), .Z(\_38_net_[26] ) );
  AND U158 ( .A(B[5]), .B(A[20]), .Z(\_38_net_[25] ) );
  AND U159 ( .A(B[4]), .B(A[20]), .Z(\_38_net_[24] ) );
  AND U160 ( .A(B[3]), .B(A[20]), .Z(\_38_net_[23] ) );
  AND U161 ( .A(B[2]), .B(A[20]), .Z(\_38_net_[22] ) );
  AND U162 ( .A(B[1]), .B(A[20]), .Z(\_38_net_[21] ) );
  AND U163 ( .A(A[20]), .B(B[0]), .Z(\_38_net_[20] ) );
  AND U164 ( .A(B[12]), .B(A[19]), .Z(\_36_net_[31] ) );
  AND U165 ( .A(B[11]), .B(A[19]), .Z(\_36_net_[30] ) );
  AND U166 ( .A(B[10]), .B(A[19]), .Z(\_36_net_[29] ) );
  AND U167 ( .A(B[9]), .B(A[19]), .Z(\_36_net_[28] ) );
  AND U168 ( .A(B[8]), .B(A[19]), .Z(\_36_net_[27] ) );
  AND U169 ( .A(B[7]), .B(A[19]), .Z(\_36_net_[26] ) );
  AND U170 ( .A(B[6]), .B(A[19]), .Z(\_36_net_[25] ) );
  AND U171 ( .A(B[5]), .B(A[19]), .Z(\_36_net_[24] ) );
  AND U172 ( .A(B[4]), .B(A[19]), .Z(\_36_net_[23] ) );
  AND U173 ( .A(B[3]), .B(A[19]), .Z(\_36_net_[22] ) );
  AND U174 ( .A(B[2]), .B(A[19]), .Z(\_36_net_[21] ) );
  AND U175 ( .A(B[1]), .B(A[19]), .Z(\_36_net_[20] ) );
  AND U176 ( .A(A[19]), .B(B[0]), .Z(\_36_net_[19] ) );
  AND U177 ( .A(B[13]), .B(A[18]), .Z(\_34_net_[31] ) );
  AND U178 ( .A(B[12]), .B(A[18]), .Z(\_34_net_[30] ) );
  AND U179 ( .A(B[11]), .B(A[18]), .Z(\_34_net_[29] ) );
  AND U180 ( .A(B[10]), .B(A[18]), .Z(\_34_net_[28] ) );
  AND U181 ( .A(B[9]), .B(A[18]), .Z(\_34_net_[27] ) );
  AND U182 ( .A(B[8]), .B(A[18]), .Z(\_34_net_[26] ) );
  AND U183 ( .A(B[7]), .B(A[18]), .Z(\_34_net_[25] ) );
  AND U184 ( .A(B[6]), .B(A[18]), .Z(\_34_net_[24] ) );
  AND U185 ( .A(B[5]), .B(A[18]), .Z(\_34_net_[23] ) );
  AND U186 ( .A(B[4]), .B(A[18]), .Z(\_34_net_[22] ) );
  AND U187 ( .A(B[3]), .B(A[18]), .Z(\_34_net_[21] ) );
  AND U188 ( .A(B[2]), .B(A[18]), .Z(\_34_net_[20] ) );
  AND U189 ( .A(B[1]), .B(A[18]), .Z(\_34_net_[19] ) );
  AND U190 ( .A(A[18]), .B(B[0]), .Z(\_34_net_[18] ) );
  AND U191 ( .A(B[14]), .B(A[17]), .Z(\_32_net_[31] ) );
  AND U192 ( .A(B[13]), .B(A[17]), .Z(\_32_net_[30] ) );
  AND U193 ( .A(B[12]), .B(A[17]), .Z(\_32_net_[29] ) );
  AND U194 ( .A(B[11]), .B(A[17]), .Z(\_32_net_[28] ) );
  AND U195 ( .A(B[10]), .B(A[17]), .Z(\_32_net_[27] ) );
  AND U196 ( .A(B[9]), .B(A[17]), .Z(\_32_net_[26] ) );
  AND U197 ( .A(B[8]), .B(A[17]), .Z(\_32_net_[25] ) );
  AND U198 ( .A(B[7]), .B(A[17]), .Z(\_32_net_[24] ) );
  AND U199 ( .A(B[6]), .B(A[17]), .Z(\_32_net_[23] ) );
  AND U200 ( .A(B[5]), .B(A[17]), .Z(\_32_net_[22] ) );
  AND U201 ( .A(B[4]), .B(A[17]), .Z(\_32_net_[21] ) );
  AND U202 ( .A(B[3]), .B(A[17]), .Z(\_32_net_[20] ) );
  AND U203 ( .A(B[2]), .B(A[17]), .Z(\_32_net_[19] ) );
  AND U204 ( .A(B[1]), .B(A[17]), .Z(\_32_net_[18] ) );
  AND U205 ( .A(A[17]), .B(B[0]), .Z(\_32_net_[17] ) );
  AND U206 ( .A(B[15]), .B(A[16]), .Z(\_30_net_[31] ) );
  AND U207 ( .A(B[14]), .B(A[16]), .Z(\_30_net_[30] ) );
  AND U208 ( .A(B[13]), .B(A[16]), .Z(\_30_net_[29] ) );
  AND U209 ( .A(B[12]), .B(A[16]), .Z(\_30_net_[28] ) );
  AND U210 ( .A(B[11]), .B(A[16]), .Z(\_30_net_[27] ) );
  AND U211 ( .A(B[10]), .B(A[16]), .Z(\_30_net_[26] ) );
  AND U212 ( .A(B[9]), .B(A[16]), .Z(\_30_net_[25] ) );
  AND U213 ( .A(B[8]), .B(A[16]), .Z(\_30_net_[24] ) );
  AND U214 ( .A(B[7]), .B(A[16]), .Z(\_30_net_[23] ) );
  AND U215 ( .A(B[6]), .B(A[16]), .Z(\_30_net_[22] ) );
  AND U216 ( .A(B[5]), .B(A[16]), .Z(\_30_net_[21] ) );
  AND U217 ( .A(B[4]), .B(A[16]), .Z(\_30_net_[20] ) );
  AND U218 ( .A(B[3]), .B(A[16]), .Z(\_30_net_[19] ) );
  AND U219 ( .A(B[2]), .B(A[16]), .Z(\_30_net_[18] ) );
  AND U220 ( .A(B[1]), .B(A[16]), .Z(\_30_net_[17] ) );
  AND U221 ( .A(A[16]), .B(B[0]), .Z(\_30_net_[16] ) );
  AND U222 ( .A(B[7]), .B(A[2]), .Z(\_2_net_[9] ) );
  AND U223 ( .A(B[6]), .B(A[2]), .Z(\_2_net_[8] ) );
  AND U224 ( .A(B[5]), .B(A[2]), .Z(\_2_net_[7] ) );
  AND U225 ( .A(B[4]), .B(A[2]), .Z(\_2_net_[6] ) );
  AND U226 ( .A(B[3]), .B(A[2]), .Z(\_2_net_[5] ) );
  AND U227 ( .A(B[2]), .B(A[2]), .Z(\_2_net_[4] ) );
  AND U228 ( .A(B[1]), .B(A[2]), .Z(\_2_net_[3] ) );
  AND U229 ( .A(A[2]), .B(B[29]), .Z(\_2_net_[31] ) );
  AND U230 ( .A(B[28]), .B(A[2]), .Z(\_2_net_[30] ) );
  AND U231 ( .A(B[0]), .B(A[2]), .Z(\_2_net_[2] ) );
  AND U232 ( .A(B[27]), .B(A[2]), .Z(\_2_net_[29] ) );
  AND U233 ( .A(B[26]), .B(A[2]), .Z(\_2_net_[28] ) );
  AND U234 ( .A(B[25]), .B(A[2]), .Z(\_2_net_[27] ) );
  AND U235 ( .A(B[24]), .B(A[2]), .Z(\_2_net_[26] ) );
  AND U236 ( .A(B[23]), .B(A[2]), .Z(\_2_net_[25] ) );
  AND U237 ( .A(B[22]), .B(A[2]), .Z(\_2_net_[24] ) );
  AND U238 ( .A(B[21]), .B(A[2]), .Z(\_2_net_[23] ) );
  AND U239 ( .A(B[20]), .B(A[2]), .Z(\_2_net_[22] ) );
  AND U240 ( .A(B[19]), .B(A[2]), .Z(\_2_net_[21] ) );
  AND U241 ( .A(B[18]), .B(A[2]), .Z(\_2_net_[20] ) );
  AND U242 ( .A(B[17]), .B(A[2]), .Z(\_2_net_[19] ) );
  AND U243 ( .A(B[16]), .B(A[2]), .Z(\_2_net_[18] ) );
  AND U244 ( .A(B[15]), .B(A[2]), .Z(\_2_net_[17] ) );
  AND U245 ( .A(B[14]), .B(A[2]), .Z(\_2_net_[16] ) );
  AND U246 ( .A(B[13]), .B(A[2]), .Z(\_2_net_[15] ) );
  AND U247 ( .A(B[12]), .B(A[2]), .Z(\_2_net_[14] ) );
  AND U248 ( .A(B[11]), .B(A[2]), .Z(\_2_net_[13] ) );
  AND U249 ( .A(B[10]), .B(A[2]), .Z(\_2_net_[12] ) );
  AND U250 ( .A(B[9]), .B(A[2]), .Z(\_2_net_[11] ) );
  AND U251 ( .A(B[8]), .B(A[2]), .Z(\_2_net_[10] ) );
  AND U252 ( .A(B[16]), .B(A[15]), .Z(\_28_net_[31] ) );
  AND U253 ( .A(B[15]), .B(A[15]), .Z(\_28_net_[30] ) );
  AND U254 ( .A(B[14]), .B(A[15]), .Z(\_28_net_[29] ) );
  AND U255 ( .A(B[13]), .B(A[15]), .Z(\_28_net_[28] ) );
  AND U256 ( .A(B[12]), .B(A[15]), .Z(\_28_net_[27] ) );
  AND U257 ( .A(B[11]), .B(A[15]), .Z(\_28_net_[26] ) );
  AND U258 ( .A(B[10]), .B(A[15]), .Z(\_28_net_[25] ) );
  AND U259 ( .A(B[9]), .B(A[15]), .Z(\_28_net_[24] ) );
  AND U260 ( .A(B[8]), .B(A[15]), .Z(\_28_net_[23] ) );
  AND U261 ( .A(B[7]), .B(A[15]), .Z(\_28_net_[22] ) );
  AND U262 ( .A(B[6]), .B(A[15]), .Z(\_28_net_[21] ) );
  AND U263 ( .A(B[5]), .B(A[15]), .Z(\_28_net_[20] ) );
  AND U264 ( .A(B[4]), .B(A[15]), .Z(\_28_net_[19] ) );
  AND U265 ( .A(B[3]), .B(A[15]), .Z(\_28_net_[18] ) );
  AND U266 ( .A(B[2]), .B(A[15]), .Z(\_28_net_[17] ) );
  AND U267 ( .A(B[1]), .B(A[15]), .Z(\_28_net_[16] ) );
  AND U268 ( .A(A[15]), .B(B[0]), .Z(\_28_net_[15] ) );
  AND U269 ( .A(B[17]), .B(A[14]), .Z(\_26_net_[31] ) );
  AND U270 ( .A(B[16]), .B(A[14]), .Z(\_26_net_[30] ) );
  AND U271 ( .A(B[15]), .B(A[14]), .Z(\_26_net_[29] ) );
  AND U272 ( .A(B[14]), .B(A[14]), .Z(\_26_net_[28] ) );
  AND U273 ( .A(B[13]), .B(A[14]), .Z(\_26_net_[27] ) );
  AND U274 ( .A(B[12]), .B(A[14]), .Z(\_26_net_[26] ) );
  AND U275 ( .A(B[11]), .B(A[14]), .Z(\_26_net_[25] ) );
  AND U276 ( .A(B[10]), .B(A[14]), .Z(\_26_net_[24] ) );
  AND U277 ( .A(B[9]), .B(A[14]), .Z(\_26_net_[23] ) );
  AND U278 ( .A(B[8]), .B(A[14]), .Z(\_26_net_[22] ) );
  AND U279 ( .A(B[7]), .B(A[14]), .Z(\_26_net_[21] ) );
  AND U280 ( .A(B[6]), .B(A[14]), .Z(\_26_net_[20] ) );
  AND U281 ( .A(B[5]), .B(A[14]), .Z(\_26_net_[19] ) );
  AND U282 ( .A(B[4]), .B(A[14]), .Z(\_26_net_[18] ) );
  AND U283 ( .A(B[3]), .B(A[14]), .Z(\_26_net_[17] ) );
  AND U284 ( .A(B[2]), .B(A[14]), .Z(\_26_net_[16] ) );
  AND U285 ( .A(B[1]), .B(A[14]), .Z(\_26_net_[15] ) );
  AND U286 ( .A(A[14]), .B(B[0]), .Z(\_26_net_[14] ) );
  AND U287 ( .A(B[18]), .B(A[13]), .Z(\_24_net_[31] ) );
  AND U288 ( .A(B[17]), .B(A[13]), .Z(\_24_net_[30] ) );
  AND U289 ( .A(B[16]), .B(A[13]), .Z(\_24_net_[29] ) );
  AND U290 ( .A(B[15]), .B(A[13]), .Z(\_24_net_[28] ) );
  AND U291 ( .A(B[14]), .B(A[13]), .Z(\_24_net_[27] ) );
  AND U292 ( .A(B[13]), .B(A[13]), .Z(\_24_net_[26] ) );
  AND U293 ( .A(B[12]), .B(A[13]), .Z(\_24_net_[25] ) );
  AND U294 ( .A(B[11]), .B(A[13]), .Z(\_24_net_[24] ) );
  AND U295 ( .A(B[10]), .B(A[13]), .Z(\_24_net_[23] ) );
  AND U296 ( .A(B[9]), .B(A[13]), .Z(\_24_net_[22] ) );
  AND U297 ( .A(B[8]), .B(A[13]), .Z(\_24_net_[21] ) );
  AND U298 ( .A(B[7]), .B(A[13]), .Z(\_24_net_[20] ) );
  AND U299 ( .A(B[6]), .B(A[13]), .Z(\_24_net_[19] ) );
  AND U300 ( .A(B[5]), .B(A[13]), .Z(\_24_net_[18] ) );
  AND U301 ( .A(B[4]), .B(A[13]), .Z(\_24_net_[17] ) );
  AND U302 ( .A(B[3]), .B(A[13]), .Z(\_24_net_[16] ) );
  AND U303 ( .A(B[2]), .B(A[13]), .Z(\_24_net_[15] ) );
  AND U304 ( .A(B[1]), .B(A[13]), .Z(\_24_net_[14] ) );
  AND U305 ( .A(A[13]), .B(B[0]), .Z(\_24_net_[13] ) );
  AND U306 ( .A(B[19]), .B(A[12]), .Z(\_22_net_[31] ) );
  AND U307 ( .A(B[18]), .B(A[12]), .Z(\_22_net_[30] ) );
  AND U308 ( .A(B[17]), .B(A[12]), .Z(\_22_net_[29] ) );
  AND U309 ( .A(B[16]), .B(A[12]), .Z(\_22_net_[28] ) );
  AND U310 ( .A(B[15]), .B(A[12]), .Z(\_22_net_[27] ) );
  AND U311 ( .A(B[14]), .B(A[12]), .Z(\_22_net_[26] ) );
  AND U312 ( .A(B[13]), .B(A[12]), .Z(\_22_net_[25] ) );
  AND U313 ( .A(B[12]), .B(A[12]), .Z(\_22_net_[24] ) );
  AND U314 ( .A(B[11]), .B(A[12]), .Z(\_22_net_[23] ) );
  AND U315 ( .A(B[10]), .B(A[12]), .Z(\_22_net_[22] ) );
  AND U316 ( .A(B[9]), .B(A[12]), .Z(\_22_net_[21] ) );
  AND U317 ( .A(B[8]), .B(A[12]), .Z(\_22_net_[20] ) );
  AND U318 ( .A(B[7]), .B(A[12]), .Z(\_22_net_[19] ) );
  AND U319 ( .A(B[6]), .B(A[12]), .Z(\_22_net_[18] ) );
  AND U320 ( .A(B[5]), .B(A[12]), .Z(\_22_net_[17] ) );
  AND U321 ( .A(B[4]), .B(A[12]), .Z(\_22_net_[16] ) );
  AND U322 ( .A(B[3]), .B(A[12]), .Z(\_22_net_[15] ) );
  AND U323 ( .A(B[2]), .B(A[12]), .Z(\_22_net_[14] ) );
  AND U324 ( .A(B[1]), .B(A[12]), .Z(\_22_net_[13] ) );
  AND U325 ( .A(A[12]), .B(B[0]), .Z(\_22_net_[12] ) );
  AND U326 ( .A(B[20]), .B(A[11]), .Z(\_20_net_[31] ) );
  AND U327 ( .A(B[19]), .B(A[11]), .Z(\_20_net_[30] ) );
  AND U328 ( .A(B[18]), .B(A[11]), .Z(\_20_net_[29] ) );
  AND U329 ( .A(B[17]), .B(A[11]), .Z(\_20_net_[28] ) );
  AND U330 ( .A(B[16]), .B(A[11]), .Z(\_20_net_[27] ) );
  AND U331 ( .A(B[15]), .B(A[11]), .Z(\_20_net_[26] ) );
  AND U332 ( .A(B[14]), .B(A[11]), .Z(\_20_net_[25] ) );
  AND U333 ( .A(B[13]), .B(A[11]), .Z(\_20_net_[24] ) );
  AND U334 ( .A(B[12]), .B(A[11]), .Z(\_20_net_[23] ) );
  AND U335 ( .A(B[11]), .B(A[11]), .Z(\_20_net_[22] ) );
  AND U336 ( .A(B[10]), .B(A[11]), .Z(\_20_net_[21] ) );
  AND U337 ( .A(B[9]), .B(A[11]), .Z(\_20_net_[20] ) );
  AND U338 ( .A(B[8]), .B(A[11]), .Z(\_20_net_[19] ) );
  AND U339 ( .A(B[7]), .B(A[11]), .Z(\_20_net_[18] ) );
  AND U340 ( .A(B[6]), .B(A[11]), .Z(\_20_net_[17] ) );
  AND U341 ( .A(B[5]), .B(A[11]), .Z(\_20_net_[16] ) );
  AND U342 ( .A(B[4]), .B(A[11]), .Z(\_20_net_[15] ) );
  AND U343 ( .A(B[3]), .B(A[11]), .Z(\_20_net_[14] ) );
  AND U344 ( .A(B[2]), .B(A[11]), .Z(\_20_net_[13] ) );
  AND U345 ( .A(B[1]), .B(A[11]), .Z(\_20_net_[12] ) );
  AND U346 ( .A(A[11]), .B(B[0]), .Z(\_20_net_[11] ) );
  AND U347 ( .A(B[21]), .B(A[10]), .Z(\_18_net_[31] ) );
  AND U348 ( .A(B[20]), .B(A[10]), .Z(\_18_net_[30] ) );
  AND U349 ( .A(B[19]), .B(A[10]), .Z(\_18_net_[29] ) );
  AND U350 ( .A(B[18]), .B(A[10]), .Z(\_18_net_[28] ) );
  AND U351 ( .A(B[17]), .B(A[10]), .Z(\_18_net_[27] ) );
  AND U352 ( .A(B[16]), .B(A[10]), .Z(\_18_net_[26] ) );
  AND U353 ( .A(B[15]), .B(A[10]), .Z(\_18_net_[25] ) );
  AND U354 ( .A(B[14]), .B(A[10]), .Z(\_18_net_[24] ) );
  AND U355 ( .A(B[13]), .B(A[10]), .Z(\_18_net_[23] ) );
  AND U356 ( .A(B[12]), .B(A[10]), .Z(\_18_net_[22] ) );
  AND U357 ( .A(B[11]), .B(A[10]), .Z(\_18_net_[21] ) );
  AND U358 ( .A(B[10]), .B(A[10]), .Z(\_18_net_[20] ) );
  AND U359 ( .A(B[9]), .B(A[10]), .Z(\_18_net_[19] ) );
  AND U360 ( .A(B[8]), .B(A[10]), .Z(\_18_net_[18] ) );
  AND U361 ( .A(B[7]), .B(A[10]), .Z(\_18_net_[17] ) );
  AND U362 ( .A(B[6]), .B(A[10]), .Z(\_18_net_[16] ) );
  AND U363 ( .A(B[5]), .B(A[10]), .Z(\_18_net_[15] ) );
  AND U364 ( .A(B[4]), .B(A[10]), .Z(\_18_net_[14] ) );
  AND U365 ( .A(B[3]), .B(A[10]), .Z(\_18_net_[13] ) );
  AND U366 ( .A(B[2]), .B(A[10]), .Z(\_18_net_[12] ) );
  AND U367 ( .A(B[1]), .B(A[10]), .Z(\_18_net_[11] ) );
  AND U368 ( .A(A[10]), .B(B[0]), .Z(\_18_net_[10] ) );
  AND U369 ( .A(B[0]), .B(A[9]), .Z(\_16_net_[9] ) );
  AND U370 ( .A(B[22]), .B(A[9]), .Z(\_16_net_[31] ) );
  AND U371 ( .A(B[21]), .B(A[9]), .Z(\_16_net_[30] ) );
  AND U372 ( .A(B[20]), .B(A[9]), .Z(\_16_net_[29] ) );
  AND U373 ( .A(B[19]), .B(A[9]), .Z(\_16_net_[28] ) );
  AND U374 ( .A(B[18]), .B(A[9]), .Z(\_16_net_[27] ) );
  AND U375 ( .A(B[17]), .B(A[9]), .Z(\_16_net_[26] ) );
  AND U376 ( .A(B[16]), .B(A[9]), .Z(\_16_net_[25] ) );
  AND U377 ( .A(B[15]), .B(A[9]), .Z(\_16_net_[24] ) );
  AND U378 ( .A(B[14]), .B(A[9]), .Z(\_16_net_[23] ) );
  AND U379 ( .A(B[13]), .B(A[9]), .Z(\_16_net_[22] ) );
  AND U380 ( .A(B[12]), .B(A[9]), .Z(\_16_net_[21] ) );
  AND U381 ( .A(B[11]), .B(A[9]), .Z(\_16_net_[20] ) );
  AND U382 ( .A(B[10]), .B(A[9]), .Z(\_16_net_[19] ) );
  AND U383 ( .A(B[9]), .B(A[9]), .Z(\_16_net_[18] ) );
  AND U384 ( .A(B[8]), .B(A[9]), .Z(\_16_net_[17] ) );
  AND U385 ( .A(B[7]), .B(A[9]), .Z(\_16_net_[16] ) );
  AND U386 ( .A(B[6]), .B(A[9]), .Z(\_16_net_[15] ) );
  AND U387 ( .A(B[5]), .B(A[9]), .Z(\_16_net_[14] ) );
  AND U388 ( .A(B[4]), .B(A[9]), .Z(\_16_net_[13] ) );
  AND U389 ( .A(B[3]), .B(A[9]), .Z(\_16_net_[12] ) );
  AND U390 ( .A(B[2]), .B(A[9]), .Z(\_16_net_[11] ) );
  AND U391 ( .A(A[9]), .B(B[1]), .Z(\_16_net_[10] ) );
  AND U392 ( .A(B[1]), .B(A[8]), .Z(\_14_net_[9] ) );
  AND U393 ( .A(B[0]), .B(A[8]), .Z(\_14_net_[8] ) );
  AND U394 ( .A(B[23]), .B(A[8]), .Z(\_14_net_[31] ) );
  AND U395 ( .A(B[22]), .B(A[8]), .Z(\_14_net_[30] ) );
  AND U396 ( .A(B[21]), .B(A[8]), .Z(\_14_net_[29] ) );
  AND U397 ( .A(B[20]), .B(A[8]), .Z(\_14_net_[28] ) );
  AND U398 ( .A(B[19]), .B(A[8]), .Z(\_14_net_[27] ) );
  AND U399 ( .A(B[18]), .B(A[8]), .Z(\_14_net_[26] ) );
  AND U400 ( .A(B[17]), .B(A[8]), .Z(\_14_net_[25] ) );
  AND U401 ( .A(B[16]), .B(A[8]), .Z(\_14_net_[24] ) );
  AND U402 ( .A(B[15]), .B(A[8]), .Z(\_14_net_[23] ) );
  AND U403 ( .A(B[14]), .B(A[8]), .Z(\_14_net_[22] ) );
  AND U404 ( .A(B[13]), .B(A[8]), .Z(\_14_net_[21] ) );
  AND U405 ( .A(B[12]), .B(A[8]), .Z(\_14_net_[20] ) );
  AND U406 ( .A(B[11]), .B(A[8]), .Z(\_14_net_[19] ) );
  AND U407 ( .A(B[10]), .B(A[8]), .Z(\_14_net_[18] ) );
  AND U408 ( .A(B[9]), .B(A[8]), .Z(\_14_net_[17] ) );
  AND U409 ( .A(B[8]), .B(A[8]), .Z(\_14_net_[16] ) );
  AND U410 ( .A(B[7]), .B(A[8]), .Z(\_14_net_[15] ) );
  AND U411 ( .A(B[6]), .B(A[8]), .Z(\_14_net_[14] ) );
  AND U412 ( .A(B[5]), .B(A[8]), .Z(\_14_net_[13] ) );
  AND U413 ( .A(B[4]), .B(A[8]), .Z(\_14_net_[12] ) );
  AND U414 ( .A(B[3]), .B(A[8]), .Z(\_14_net_[11] ) );
  AND U415 ( .A(A[8]), .B(B[2]), .Z(\_14_net_[10] ) );
  AND U416 ( .A(B[2]), .B(A[7]), .Z(\_12_net_[9] ) );
  AND U417 ( .A(B[1]), .B(A[7]), .Z(\_12_net_[8] ) );
  AND U418 ( .A(B[0]), .B(A[7]), .Z(\_12_net_[7] ) );
  AND U419 ( .A(B[24]), .B(A[7]), .Z(\_12_net_[31] ) );
  AND U420 ( .A(B[23]), .B(A[7]), .Z(\_12_net_[30] ) );
  AND U421 ( .A(B[22]), .B(A[7]), .Z(\_12_net_[29] ) );
  AND U422 ( .A(B[21]), .B(A[7]), .Z(\_12_net_[28] ) );
  AND U423 ( .A(B[20]), .B(A[7]), .Z(\_12_net_[27] ) );
  AND U424 ( .A(B[19]), .B(A[7]), .Z(\_12_net_[26] ) );
  AND U425 ( .A(B[18]), .B(A[7]), .Z(\_12_net_[25] ) );
  AND U426 ( .A(B[17]), .B(A[7]), .Z(\_12_net_[24] ) );
  AND U427 ( .A(B[16]), .B(A[7]), .Z(\_12_net_[23] ) );
  AND U428 ( .A(B[15]), .B(A[7]), .Z(\_12_net_[22] ) );
  AND U429 ( .A(B[14]), .B(A[7]), .Z(\_12_net_[21] ) );
  AND U430 ( .A(B[13]), .B(A[7]), .Z(\_12_net_[20] ) );
  AND U431 ( .A(B[12]), .B(A[7]), .Z(\_12_net_[19] ) );
  AND U432 ( .A(B[11]), .B(A[7]), .Z(\_12_net_[18] ) );
  AND U433 ( .A(B[10]), .B(A[7]), .Z(\_12_net_[17] ) );
  AND U434 ( .A(B[9]), .B(A[7]), .Z(\_12_net_[16] ) );
  AND U435 ( .A(B[8]), .B(A[7]), .Z(\_12_net_[15] ) );
  AND U436 ( .A(B[7]), .B(A[7]), .Z(\_12_net_[14] ) );
  AND U437 ( .A(B[6]), .B(A[7]), .Z(\_12_net_[13] ) );
  AND U438 ( .A(B[5]), .B(A[7]), .Z(\_12_net_[12] ) );
  AND U439 ( .A(B[4]), .B(A[7]), .Z(\_12_net_[11] ) );
  AND U440 ( .A(A[7]), .B(B[3]), .Z(\_12_net_[10] ) );
  AND U441 ( .A(B[3]), .B(A[6]), .Z(\_10_net_[9] ) );
  AND U442 ( .A(B[2]), .B(A[6]), .Z(\_10_net_[8] ) );
  AND U443 ( .A(B[1]), .B(A[6]), .Z(\_10_net_[7] ) );
  AND U444 ( .A(B[0]), .B(A[6]), .Z(\_10_net_[6] ) );
  AND U445 ( .A(B[25]), .B(A[6]), .Z(\_10_net_[31] ) );
  AND U446 ( .A(B[24]), .B(A[6]), .Z(\_10_net_[30] ) );
  AND U447 ( .A(B[23]), .B(A[6]), .Z(\_10_net_[29] ) );
  AND U448 ( .A(B[22]), .B(A[6]), .Z(\_10_net_[28] ) );
  AND U449 ( .A(B[21]), .B(A[6]), .Z(\_10_net_[27] ) );
  AND U450 ( .A(B[20]), .B(A[6]), .Z(\_10_net_[26] ) );
  AND U451 ( .A(B[19]), .B(A[6]), .Z(\_10_net_[25] ) );
  AND U452 ( .A(B[18]), .B(A[6]), .Z(\_10_net_[24] ) );
  AND U453 ( .A(B[17]), .B(A[6]), .Z(\_10_net_[23] ) );
  AND U454 ( .A(B[16]), .B(A[6]), .Z(\_10_net_[22] ) );
  AND U455 ( .A(B[15]), .B(A[6]), .Z(\_10_net_[21] ) );
  AND U456 ( .A(B[14]), .B(A[6]), .Z(\_10_net_[20] ) );
  AND U457 ( .A(B[13]), .B(A[6]), .Z(\_10_net_[19] ) );
  AND U458 ( .A(B[12]), .B(A[6]), .Z(\_10_net_[18] ) );
  AND U459 ( .A(B[11]), .B(A[6]), .Z(\_10_net_[17] ) );
  AND U460 ( .A(B[10]), .B(A[6]), .Z(\_10_net_[16] ) );
  AND U461 ( .A(B[9]), .B(A[6]), .Z(\_10_net_[15] ) );
  AND U462 ( .A(B[8]), .B(A[6]), .Z(\_10_net_[14] ) );
  AND U463 ( .A(B[7]), .B(A[6]), .Z(\_10_net_[13] ) );
  AND U464 ( .A(B[6]), .B(A[6]), .Z(\_10_net_[12] ) );
  AND U465 ( .A(B[5]), .B(A[6]), .Z(\_10_net_[11] ) );
  AND U466 ( .A(A[6]), .B(B[4]), .Z(\_10_net_[10] ) );
  AND U467 ( .A(B[8]), .B(A[1]), .Z(\_0_net_[9] ) );
  AND U468 ( .A(B[7]), .B(A[1]), .Z(\_0_net_[8] ) );
  AND U469 ( .A(B[6]), .B(A[1]), .Z(\_0_net_[7] ) );
  AND U470 ( .A(B[5]), .B(A[1]), .Z(\_0_net_[6] ) );
  AND U471 ( .A(B[4]), .B(A[1]), .Z(\_0_net_[5] ) );
  AND U472 ( .A(B[3]), .B(A[1]), .Z(\_0_net_[4] ) );
  AND U473 ( .A(B[2]), .B(A[1]), .Z(\_0_net_[3] ) );
  AND U474 ( .A(B[30]), .B(A[1]), .Z(\_0_net_[31] ) );
  AND U475 ( .A(B[29]), .B(A[1]), .Z(\_0_net_[30] ) );
  AND U476 ( .A(B[1]), .B(A[1]), .Z(\_0_net_[2] ) );
  AND U477 ( .A(B[28]), .B(A[1]), .Z(\_0_net_[29] ) );
  AND U478 ( .A(B[27]), .B(A[1]), .Z(\_0_net_[28] ) );
  AND U479 ( .A(B[26]), .B(A[1]), .Z(\_0_net_[27] ) );
  AND U480 ( .A(B[25]), .B(A[1]), .Z(\_0_net_[26] ) );
  AND U481 ( .A(B[24]), .B(A[1]), .Z(\_0_net_[25] ) );
  AND U482 ( .A(B[23]), .B(A[1]), .Z(\_0_net_[24] ) );
  AND U483 ( .A(B[22]), .B(A[1]), .Z(\_0_net_[23] ) );
  AND U484 ( .A(B[21]), .B(A[1]), .Z(\_0_net_[22] ) );
  AND U485 ( .A(B[20]), .B(A[1]), .Z(\_0_net_[21] ) );
  AND U486 ( .A(B[19]), .B(A[1]), .Z(\_0_net_[20] ) );
  AND U487 ( .A(B[0]), .B(A[1]), .Z(\_0_net_[1] ) );
  AND U488 ( .A(B[18]), .B(A[1]), .Z(\_0_net_[19] ) );
  AND U489 ( .A(B[17]), .B(A[1]), .Z(\_0_net_[18] ) );
  AND U490 ( .A(B[16]), .B(A[1]), .Z(\_0_net_[17] ) );
  AND U491 ( .A(B[15]), .B(A[1]), .Z(\_0_net_[16] ) );
  AND U492 ( .A(B[14]), .B(A[1]), .Z(\_0_net_[15] ) );
  AND U493 ( .A(B[13]), .B(A[1]), .Z(\_0_net_[14] ) );
  AND U494 ( .A(B[12]), .B(A[1]), .Z(\_0_net_[13] ) );
  AND U495 ( .A(B[11]), .B(A[1]), .Z(\_0_net_[12] ) );
  AND U496 ( .A(B[10]), .B(A[1]), .Z(\_0_net_[11] ) );
  AND U497 ( .A(A[1]), .B(B[9]), .Z(\_0_net_[10] ) );
endmodule


module FA_3969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(A), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(B), .Z(n1) );
endmodule


module FA_3970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_3999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N32_96 ( A, B, CI, S, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input CI;
  output CO;

  wire   [31:1] C;

  FA_3999 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_3998 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_3997 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_3996 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_3995 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_3994 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_3993 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_3992 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_3991 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_3990 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_3989 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_3988 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_3987 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_3986 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_3985 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_3984 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_3983 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_3982 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_3981 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_3980 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_3979 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_3978 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_3977 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_3976 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_3975 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_3974 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_3973 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_3972 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_3971 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_3970 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_3969 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]) );
endmodule


module matrixMult_N_M_3_N16_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;

  wire   [31:0] xy;
  wire   [31:0] oi;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign o[0] = 1'b0;

  MULT_N32_3 MULT_ ( .A({x[31:1], 1'b0}), .B({1'b0, y[30:0]}), .O({xy[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  ADD_N32_96 ADD_ ( .A({xy[31:1], 1'b0}), .B({o[31:1], 1'b0}), .CI(1'b0), .S({
        oi[31:1], SYNOPSYS_UNCONNECTED__1}) );
  DFF \o_reg[1]  ( .D(oi[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(oi[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(oi[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(oi[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(oi[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(oi[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(oi[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(oi[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(oi[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(oi[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10]) );
  DFF \o_reg[11]  ( .D(oi[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11]) );
  DFF \o_reg[12]  ( .D(oi[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12]) );
  DFF \o_reg[13]  ( .D(oi[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13]) );
  DFF \o_reg[14]  ( .D(oi[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14]) );
  DFF \o_reg[15]  ( .D(oi[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15]) );
  DFF \o_reg[16]  ( .D(oi[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16]) );
  DFF \o_reg[17]  ( .D(oi[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17]) );
  DFF \o_reg[18]  ( .D(oi[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18]) );
  DFF \o_reg[19]  ( .D(oi[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19]) );
  DFF \o_reg[20]  ( .D(oi[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20]) );
  DFF \o_reg[21]  ( .D(oi[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21]) );
  DFF \o_reg[22]  ( .D(oi[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22]) );
  DFF \o_reg[23]  ( .D(oi[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23]) );
  DFF \o_reg[24]  ( .D(oi[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24]) );
  DFF \o_reg[25]  ( .D(oi[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25]) );
  DFF \o_reg[26]  ( .D(oi[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26]) );
  DFF \o_reg[27]  ( .D(oi[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27]) );
  DFF \o_reg[28]  ( .D(oi[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28]) );
  DFF \o_reg[29]  ( .D(oi[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29]) );
  DFF \o_reg[30]  ( .D(oi[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30]) );
  DFF \o_reg[31]  ( .D(oi[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31]) );
endmodule

