
module mult_N128_CC8 ( clk, rst, a, b, c );
  input [127:0] a;
  input [15:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165;
  wire   [255:0] sreg;

  DFF \sreg_reg[239]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[118]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[117]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[116]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[115]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[114]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[113]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[112]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U19 ( .A(n689), .B(n688), .Z(n1) );
  NANDN U20 ( .A(n686), .B(n687), .Z(n2) );
  NAND U21 ( .A(n1), .B(n2), .Z(n797) );
  NANDN U22 ( .A(n855), .B(n856), .Z(n3) );
  NANDN U23 ( .A(n854), .B(n853), .Z(n4) );
  NAND U24 ( .A(n3), .B(n4), .Z(n888) );
  NAND U25 ( .A(n9485), .B(n646), .Z(n5) );
  NAND U26 ( .A(n73), .B(n92), .Z(n6) );
  NAND U27 ( .A(n6), .B(n5), .Z(n7) );
  NAND U28 ( .A(n7), .B(b[3]), .Z(n119) );
  OR U29 ( .A(n10008), .B(n10009), .Z(n8) );
  NANDN U30 ( .A(n10011), .B(n10010), .Z(n9) );
  AND U31 ( .A(n8), .B(n9), .Z(n10054) );
  NANDN U32 ( .A(n889), .B(n890), .Z(n10) );
  NANDN U33 ( .A(n888), .B(n887), .Z(n11) );
  NAND U34 ( .A(n10), .B(n11), .Z(n1025) );
  NANDN U35 ( .A(n817), .B(n818), .Z(n12) );
  NANDN U36 ( .A(n816), .B(n815), .Z(n13) );
  NAND U37 ( .A(n12), .B(n13), .Z(n881) );
  NANDN U38 ( .A(n10043), .B(n10044), .Z(n14) );
  NANDN U39 ( .A(n10042), .B(n10080), .Z(n15) );
  NAND U40 ( .A(n14), .B(n15), .Z(n10064) );
  XOR U41 ( .A(n126), .B(n125), .Z(n16) );
  NANDN U42 ( .A(n124), .B(n16), .Z(n17) );
  NAND U43 ( .A(n126), .B(n125), .Z(n18) );
  AND U44 ( .A(n17), .B(n18), .Z(n155) );
  NANDN U45 ( .A(n9719), .B(n9718), .Z(n19) );
  NANDN U46 ( .A(n9720), .B(n9721), .Z(n20) );
  AND U47 ( .A(n19), .B(n20), .Z(n9725) );
  XNOR U48 ( .A(n9894), .B(n9895), .Z(n9900) );
  XOR U49 ( .A(n9597), .B(n9596), .Z(n21) );
  NANDN U50 ( .A(n9595), .B(n21), .Z(n22) );
  NAND U51 ( .A(n9597), .B(n9596), .Z(n23) );
  AND U52 ( .A(n22), .B(n23), .Z(n9661) );
  XOR U53 ( .A(n10035), .B(n10034), .Z(n24) );
  NANDN U54 ( .A(n10033), .B(n24), .Z(n25) );
  NAND U55 ( .A(n10035), .B(n10034), .Z(n26) );
  AND U56 ( .A(n25), .B(n26), .Z(n10063) );
  NANDN U57 ( .A(n859), .B(n860), .Z(n27) );
  NANDN U58 ( .A(n858), .B(n857), .Z(n28) );
  NAND U59 ( .A(n27), .B(n28), .Z(n937) );
  NAND U60 ( .A(n2417), .B(n2416), .Z(n29) );
  NANDN U61 ( .A(n2414), .B(n2415), .Z(n30) );
  NAND U62 ( .A(n29), .B(n30), .Z(n2442) );
  NAND U63 ( .A(n7151), .B(n7150), .Z(n31) );
  NANDN U64 ( .A(n7148), .B(n7149), .Z(n32) );
  NAND U65 ( .A(n31), .B(n32), .Z(n7198) );
  XOR U66 ( .A(n9250), .B(n9251), .Z(n9253) );
  OR U67 ( .A(b[0]), .B(n10049), .Z(n33) );
  AND U68 ( .A(b[1]), .B(n33), .Z(n9494) );
  NANDN U69 ( .A(n603), .B(n604), .Z(n34) );
  NANDN U70 ( .A(n602), .B(n601), .Z(n35) );
  NAND U71 ( .A(n34), .B(n35), .Z(n680) );
  XNOR U72 ( .A(n585), .B(n586), .Z(n580) );
  NANDN U73 ( .A(n730), .B(n729), .Z(n36) );
  NANDN U74 ( .A(n731), .B(n732), .Z(n37) );
  AND U75 ( .A(n36), .B(n37), .Z(n739) );
  OR U76 ( .A(n795), .B(n794), .Z(n38) );
  NANDN U77 ( .A(n797), .B(n796), .Z(n39) );
  NAND U78 ( .A(n38), .B(n39), .Z(n815) );
  NANDN U79 ( .A(n9329), .B(n9330), .Z(n40) );
  NANDN U80 ( .A(n9328), .B(n9327), .Z(n41) );
  NAND U81 ( .A(n40), .B(n41), .Z(n9380) );
  XOR U82 ( .A(n9407), .B(n9408), .Z(n9410) );
  XNOR U83 ( .A(n9534), .B(n9535), .Z(n9530) );
  NANDN U84 ( .A(n194), .B(n195), .Z(n42) );
  NANDN U85 ( .A(n193), .B(n192), .Z(n43) );
  NAND U86 ( .A(n42), .B(n43), .Z(n231) );
  OR U87 ( .A(n473), .B(n472), .Z(n44) );
  NANDN U88 ( .A(n475), .B(n474), .Z(n45) );
  NAND U89 ( .A(n44), .B(n45), .Z(n536) );
  XOR U90 ( .A(n9652), .B(n9653), .Z(n9647) );
  NANDN U91 ( .A(n9765), .B(n9792), .Z(n46) );
  NANDN U92 ( .A(n9766), .B(n9767), .Z(n47) );
  AND U93 ( .A(n46), .B(n47), .Z(n9781) );
  XNOR U94 ( .A(n10080), .B(n10081), .Z(n10085) );
  NANDN U95 ( .A(n959), .B(n960), .Z(n48) );
  NANDN U96 ( .A(n958), .B(n957), .Z(n49) );
  NAND U97 ( .A(n48), .B(n49), .Z(n1036) );
  OR U98 ( .A(n9730), .B(n9731), .Z(n50) );
  NAND U99 ( .A(n9733), .B(n9732), .Z(n51) );
  NAND U100 ( .A(n50), .B(n51), .Z(n9831) );
  NAND U101 ( .A(n9789), .B(n9788), .Z(n52) );
  NANDN U102 ( .A(n9786), .B(n9787), .Z(n53) );
  NAND U103 ( .A(n52), .B(n53), .Z(n9841) );
  XOR U104 ( .A(n10050), .B(b[14]), .Z(n10106) );
  XOR U105 ( .A(n120), .B(n119), .Z(n54) );
  NANDN U106 ( .A(n118), .B(n54), .Z(n55) );
  NAND U107 ( .A(n120), .B(n119), .Z(n56) );
  AND U108 ( .A(n55), .B(n56), .Z(n126) );
  NANDN U109 ( .A(n311), .B(n312), .Z(n57) );
  NANDN U110 ( .A(n310), .B(n309), .Z(n58) );
  NAND U111 ( .A(n57), .B(n58), .Z(n351) );
  NANDN U112 ( .A(n670), .B(n671), .Z(n59) );
  NANDN U113 ( .A(n672), .B(n673), .Z(n60) );
  NAND U114 ( .A(n59), .B(n60), .Z(n736) );
  NANDN U115 ( .A(n9371), .B(n9372), .Z(n61) );
  NANDN U116 ( .A(n9370), .B(n9369), .Z(n62) );
  NAND U117 ( .A(n61), .B(n62), .Z(n9447) );
  NAND U118 ( .A(n9661), .B(n9659), .Z(n63) );
  XOR U119 ( .A(n9659), .B(n9661), .Z(n64) );
  NAND U120 ( .A(n64), .B(n9660), .Z(n65) );
  NAND U121 ( .A(n63), .B(n65), .Z(n9726) );
  NAND U122 ( .A(n9948), .B(n9946), .Z(n66) );
  XOR U123 ( .A(n9946), .B(n9948), .Z(n67) );
  NANDN U124 ( .A(n9947), .B(n67), .Z(n68) );
  NAND U125 ( .A(n66), .B(n68), .Z(n9992) );
  NAND U126 ( .A(n10063), .B(n10062), .Z(n69) );
  XOR U127 ( .A(n10062), .B(n10063), .Z(n70) );
  NAND U128 ( .A(n70), .B(n10061), .Z(n71) );
  NAND U129 ( .A(n69), .B(n71), .Z(n10096) );
  IV U130 ( .A(b[0]), .Z(n72) );
  IV U131 ( .A(b[1]), .Z(n73) );
  IV U132 ( .A(b[3]), .Z(n74) );
  IV U133 ( .A(b[15]), .Z(n75) );
  NAND U134 ( .A(b[0]), .B(a[0]), .Z(n77) );
  XNOR U135 ( .A(n77), .B(sreg[112]), .Z(c[112]) );
  NAND U136 ( .A(b[0]), .B(a[1]), .Z(n82) );
  NAND U137 ( .A(b[1]), .B(a[0]), .Z(n76) );
  XOR U138 ( .A(n82), .B(n76), .Z(n85) );
  XNOR U139 ( .A(sreg[113]), .B(n85), .Z(n87) );
  NANDN U140 ( .A(n77), .B(sreg[112]), .Z(n86) );
  XOR U141 ( .A(n87), .B(n86), .Z(c[113]) );
  NAND U142 ( .A(b[0]), .B(a[2]), .Z(n78) );
  XNOR U143 ( .A(b[1]), .B(n78), .Z(n80) );
  NAND U144 ( .A(a[1]), .B(n72), .Z(n79) );
  AND U145 ( .A(n80), .B(n79), .Z(n90) );
  NAND U146 ( .A(b[2]), .B(a[0]), .Z(n81) );
  XNOR U147 ( .A(b[1]), .B(n81), .Z(n84) );
  IV U148 ( .A(a[0]), .Z(n646) );
  NANDN U149 ( .A(n82), .B(n646), .Z(n83) );
  AND U150 ( .A(n84), .B(n83), .Z(n91) );
  XOR U151 ( .A(n90), .B(n91), .Z(n103) );
  NAND U152 ( .A(n85), .B(sreg[113]), .Z(n89) );
  OR U153 ( .A(n87), .B(n86), .Z(n88) );
  NAND U154 ( .A(n89), .B(n88), .Z(n102) );
  XNOR U155 ( .A(n102), .B(sreg[114]), .Z(n104) );
  XNOR U156 ( .A(n103), .B(n104), .Z(c[114]) );
  NAND U157 ( .A(n91), .B(n90), .Z(n120) );
  IV U158 ( .A(b[2]), .Z(n92) );
  XNOR U159 ( .A(b[1]), .B(n92), .Z(n9485) );
  XOR U160 ( .A(b[3]), .B(b[1]), .Z(n94) );
  XOR U161 ( .A(b[3]), .B(b[2]), .Z(n93) );
  AND U162 ( .A(n94), .B(n93), .Z(n9484) );
  XOR U163 ( .A(b[3]), .B(a[0]), .Z(n95) );
  AND U164 ( .A(n9484), .B(n95), .Z(n97) );
  XNOR U165 ( .A(b[3]), .B(a[1]), .Z(n115) );
  NANDN U166 ( .A(n115), .B(n9485), .Z(n96) );
  NANDN U167 ( .A(n97), .B(n96), .Z(n121) );
  NAND U168 ( .A(b[0]), .B(a[3]), .Z(n98) );
  XNOR U169 ( .A(b[1]), .B(n98), .Z(n100) );
  NAND U170 ( .A(a[2]), .B(n72), .Z(n99) );
  NAND U171 ( .A(n100), .B(n99), .Z(n122) );
  XNOR U172 ( .A(n121), .B(n122), .Z(n118) );
  XNOR U173 ( .A(n119), .B(n118), .Z(n101) );
  XNOR U174 ( .A(n120), .B(n101), .Z(n107) );
  XNOR U175 ( .A(sreg[115]), .B(n107), .Z(n109) );
  NAND U176 ( .A(n102), .B(sreg[114]), .Z(n106) );
  NANDN U177 ( .A(n104), .B(n103), .Z(n105) );
  AND U178 ( .A(n106), .B(n105), .Z(n108) );
  XOR U179 ( .A(n109), .B(n108), .Z(c[115]) );
  NAND U180 ( .A(sreg[115]), .B(n107), .Z(n111) );
  OR U181 ( .A(n109), .B(n108), .Z(n110) );
  NAND U182 ( .A(n111), .B(n110), .Z(n147) );
  XNOR U183 ( .A(n147), .B(sreg[116]), .Z(n149) );
  XNOR U184 ( .A(b[3]), .B(b[4]), .Z(n9623) );
  ANDN U185 ( .B(a[0]), .A(n9623), .Z(n144) );
  NAND U186 ( .A(b[0]), .B(a[4]), .Z(n112) );
  XNOR U187 ( .A(b[1]), .B(n112), .Z(n114) );
  NAND U188 ( .A(a[3]), .B(n72), .Z(n113) );
  AND U189 ( .A(n114), .B(n113), .Z(n142) );
  NANDN U190 ( .A(n115), .B(n9484), .Z(n117) );
  IV U191 ( .A(a[2]), .Z(n705) );
  XNOR U192 ( .A(b[3]), .B(n705), .Z(n138) );
  NAND U193 ( .A(n138), .B(n9485), .Z(n116) );
  AND U194 ( .A(n117), .B(n116), .Z(n141) );
  XNOR U195 ( .A(n142), .B(n141), .Z(n143) );
  XOR U196 ( .A(n144), .B(n143), .Z(n125) );
  NANDN U197 ( .A(n122), .B(n121), .Z(n124) );
  XOR U198 ( .A(n126), .B(n124), .Z(n123) );
  XOR U199 ( .A(n125), .B(n123), .Z(n148) );
  XOR U200 ( .A(n149), .B(n148), .Z(c[116]) );
  NAND U201 ( .A(b[0]), .B(a[5]), .Z(n127) );
  XNOR U202 ( .A(b[1]), .B(n127), .Z(n129) );
  NAND U203 ( .A(a[4]), .B(n72), .Z(n128) );
  AND U204 ( .A(n129), .B(n128), .Z(n158) );
  IV U205 ( .A(a[1]), .Z(n628) );
  XNOR U206 ( .A(b[5]), .B(n628), .Z(n166) );
  ANDN U207 ( .B(n166), .A(n9623), .Z(n134) );
  XOR U208 ( .A(b[5]), .B(a[0]), .Z(n132) );
  XOR U209 ( .A(b[5]), .B(b[3]), .Z(n131) );
  XOR U210 ( .A(b[5]), .B(b[4]), .Z(n130) );
  AND U211 ( .A(n131), .B(n130), .Z(n9680) );
  NAND U212 ( .A(n132), .B(n9680), .Z(n133) );
  NANDN U213 ( .A(n134), .B(n133), .Z(n159) );
  XNOR U214 ( .A(n158), .B(n159), .Z(n172) );
  ANDN U215 ( .B(n74), .A(b[4]), .Z(n135) );
  NAND U216 ( .A(b[5]), .B(n135), .Z(n137) );
  IV U217 ( .A(b[5]), .Z(n9622) );
  NOR U218 ( .A(n9622), .B(n9623), .Z(n9683) );
  NAND U219 ( .A(n646), .B(n9683), .Z(n136) );
  NAND U220 ( .A(n137), .B(n136), .Z(n170) );
  NAND U221 ( .A(n9484), .B(n138), .Z(n140) );
  XOR U222 ( .A(b[3]), .B(a[3]), .Z(n160) );
  NAND U223 ( .A(n160), .B(n9485), .Z(n139) );
  AND U224 ( .A(n140), .B(n139), .Z(n169) );
  XNOR U225 ( .A(n170), .B(n169), .Z(n171) );
  XOR U226 ( .A(n172), .B(n171), .Z(n152) );
  NANDN U227 ( .A(n142), .B(n141), .Z(n146) );
  NANDN U228 ( .A(n144), .B(n143), .Z(n145) );
  NAND U229 ( .A(n146), .B(n145), .Z(n153) );
  XOR U230 ( .A(n152), .B(n153), .Z(n154) );
  XNOR U231 ( .A(n155), .B(n154), .Z(n175) );
  XNOR U232 ( .A(sreg[117]), .B(n175), .Z(n177) );
  NAND U233 ( .A(n147), .B(sreg[116]), .Z(n151) );
  OR U234 ( .A(n149), .B(n148), .Z(n150) );
  AND U235 ( .A(n151), .B(n150), .Z(n176) );
  XOR U236 ( .A(n177), .B(n176), .Z(c[117]) );
  OR U237 ( .A(n153), .B(n152), .Z(n157) );
  NANDN U238 ( .A(n155), .B(n154), .Z(n156) );
  NAND U239 ( .A(n157), .B(n156), .Z(n183) );
  AND U240 ( .A(n159), .B(n158), .Z(n189) );
  IV U241 ( .A(a[4]), .Z(n834) );
  XNOR U242 ( .A(b[3]), .B(n834), .Z(n196) );
  NAND U243 ( .A(n196), .B(n9485), .Z(n162) );
  NAND U244 ( .A(n160), .B(n9484), .Z(n161) );
  NAND U245 ( .A(n162), .B(n161), .Z(n195) );
  NAND U246 ( .A(b[0]), .B(a[6]), .Z(n163) );
  XNOR U247 ( .A(b[1]), .B(n163), .Z(n165) );
  NAND U248 ( .A(a[5]), .B(n72), .Z(n164) );
  AND U249 ( .A(n165), .B(n164), .Z(n192) );
  XOR U250 ( .A(b[5]), .B(b[6]), .Z(n9746) );
  NAND U251 ( .A(a[0]), .B(n9746), .Z(n193) );
  XOR U252 ( .A(n192), .B(n193), .Z(n194) );
  XOR U253 ( .A(n195), .B(n194), .Z(n186) );
  NAND U254 ( .A(n9680), .B(n166), .Z(n168) );
  XOR U255 ( .A(b[5]), .B(a[2]), .Z(n199) );
  NANDN U256 ( .A(n9623), .B(n199), .Z(n167) );
  NAND U257 ( .A(n168), .B(n167), .Z(n187) );
  XNOR U258 ( .A(n186), .B(n187), .Z(n188) );
  XOR U259 ( .A(n189), .B(n188), .Z(n180) );
  NANDN U260 ( .A(n170), .B(n169), .Z(n174) );
  NAND U261 ( .A(n172), .B(n171), .Z(n173) );
  NAND U262 ( .A(n174), .B(n173), .Z(n181) );
  XNOR U263 ( .A(n180), .B(n181), .Z(n182) );
  XNOR U264 ( .A(n183), .B(n182), .Z(n216) );
  NAND U265 ( .A(sreg[117]), .B(n175), .Z(n179) );
  OR U266 ( .A(n177), .B(n176), .Z(n178) );
  NAND U267 ( .A(n179), .B(n178), .Z(n214) );
  XNOR U268 ( .A(n214), .B(sreg[118]), .Z(n215) );
  XOR U269 ( .A(n216), .B(n215), .Z(c[118]) );
  NANDN U270 ( .A(n181), .B(n180), .Z(n185) );
  NAND U271 ( .A(n183), .B(n182), .Z(n184) );
  NAND U272 ( .A(n185), .B(n184), .Z(n227) );
  NANDN U273 ( .A(n187), .B(n186), .Z(n191) );
  NANDN U274 ( .A(n189), .B(n188), .Z(n190) );
  NAND U275 ( .A(n191), .B(n190), .Z(n225) );
  NAND U276 ( .A(n9484), .B(n196), .Z(n198) );
  XOR U277 ( .A(b[3]), .B(a[5]), .Z(n245) );
  NAND U278 ( .A(n245), .B(n9485), .Z(n197) );
  AND U279 ( .A(n198), .B(n197), .Z(n230) );
  XNOR U280 ( .A(n231), .B(n230), .Z(n232) );
  IV U281 ( .A(a[3]), .Z(n754) );
  XNOR U282 ( .A(n9622), .B(n754), .Z(n253) );
  OR U283 ( .A(n253), .B(n9623), .Z(n201) );
  NAND U284 ( .A(n199), .B(n9680), .Z(n200) );
  NAND U285 ( .A(n201), .B(n200), .Z(n248) );
  XOR U286 ( .A(b[7]), .B(a[0]), .Z(n204) );
  XOR U287 ( .A(b[7]), .B(b[5]), .Z(n203) );
  XOR U288 ( .A(b[7]), .B(b[6]), .Z(n202) );
  AND U289 ( .A(n203), .B(n202), .Z(n9747) );
  NAND U290 ( .A(n204), .B(n9747), .Z(n206) );
  XOR U291 ( .A(b[7]), .B(a[1]), .Z(n242) );
  NAND U292 ( .A(n242), .B(n9746), .Z(n205) );
  NAND U293 ( .A(n206), .B(n205), .Z(n249) );
  XNOR U294 ( .A(n248), .B(n249), .Z(n239) );
  AND U295 ( .A(a[0]), .B(b[5]), .Z(n210) );
  NAND U296 ( .A(n646), .B(n9622), .Z(n207) );
  NAND U297 ( .A(n207), .B(b[6]), .Z(n208) );
  AND U298 ( .A(n208), .B(b[7]), .Z(n209) );
  NANDN U299 ( .A(n210), .B(n209), .Z(n236) );
  NAND U300 ( .A(b[0]), .B(a[7]), .Z(n211) );
  XNOR U301 ( .A(b[1]), .B(n211), .Z(n213) );
  NAND U302 ( .A(a[6]), .B(n72), .Z(n212) );
  AND U303 ( .A(n213), .B(n212), .Z(n237) );
  XNOR U304 ( .A(n236), .B(n237), .Z(n238) );
  XOR U305 ( .A(n239), .B(n238), .Z(n233) );
  XOR U306 ( .A(n232), .B(n233), .Z(n224) );
  XNOR U307 ( .A(n225), .B(n224), .Z(n226) );
  XNOR U308 ( .A(n227), .B(n226), .Z(n219) );
  XNOR U309 ( .A(n219), .B(sreg[119]), .Z(n221) );
  NAND U310 ( .A(n214), .B(sreg[118]), .Z(n218) );
  OR U311 ( .A(n216), .B(n215), .Z(n217) );
  AND U312 ( .A(n218), .B(n217), .Z(n220) );
  XOR U313 ( .A(n221), .B(n220), .Z(c[119]) );
  NAND U314 ( .A(n219), .B(sreg[119]), .Z(n223) );
  OR U315 ( .A(n221), .B(n220), .Z(n222) );
  NAND U316 ( .A(n223), .B(n222), .Z(n299) );
  XNOR U317 ( .A(n299), .B(sreg[120]), .Z(n301) );
  NAND U318 ( .A(n225), .B(n224), .Z(n229) );
  OR U319 ( .A(n227), .B(n226), .Z(n228) );
  NAND U320 ( .A(n229), .B(n228), .Z(n259) );
  NANDN U321 ( .A(n231), .B(n230), .Z(n235) );
  NAND U322 ( .A(n233), .B(n232), .Z(n234) );
  NAND U323 ( .A(n235), .B(n234), .Z(n256) );
  NANDN U324 ( .A(n237), .B(n236), .Z(n241) );
  NAND U325 ( .A(n239), .B(n238), .Z(n240) );
  NAND U326 ( .A(n241), .B(n240), .Z(n296) );
  IV U327 ( .A(b[7]), .Z(n9872) );
  XNOR U328 ( .A(n9872), .B(n705), .Z(n268) );
  NANDN U329 ( .A(n268), .B(n9746), .Z(n244) );
  NAND U330 ( .A(n242), .B(n9747), .Z(n243) );
  NAND U331 ( .A(n244), .B(n243), .Z(n281) );
  IV U332 ( .A(a[6]), .Z(n970) );
  XNOR U333 ( .A(b[3]), .B(n970), .Z(n265) );
  NAND U334 ( .A(n265), .B(n9485), .Z(n247) );
  NAND U335 ( .A(n245), .B(n9484), .Z(n246) );
  AND U336 ( .A(n247), .B(n246), .Z(n282) );
  XNOR U337 ( .A(n281), .B(n282), .Z(n283) );
  NAND U338 ( .A(n249), .B(n248), .Z(n284) );
  XOR U339 ( .A(n283), .B(n284), .Z(n293) );
  XOR U340 ( .A(b[7]), .B(b[8]), .Z(n9865) );
  NANDN U341 ( .A(n646), .B(n9865), .Z(n290) );
  NAND U342 ( .A(b[0]), .B(a[8]), .Z(n250) );
  XNOR U343 ( .A(b[1]), .B(n250), .Z(n252) );
  NAND U344 ( .A(a[7]), .B(n72), .Z(n251) );
  AND U345 ( .A(n252), .B(n251), .Z(n288) );
  NANDN U346 ( .A(n253), .B(n9680), .Z(n255) );
  XOR U347 ( .A(b[5]), .B(a[4]), .Z(n278) );
  NANDN U348 ( .A(n9623), .B(n278), .Z(n254) );
  AND U349 ( .A(n255), .B(n254), .Z(n287) );
  XNOR U350 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U351 ( .A(n290), .B(n289), .Z(n294) );
  XNOR U352 ( .A(n293), .B(n294), .Z(n295) );
  XNOR U353 ( .A(n296), .B(n295), .Z(n257) );
  XNOR U354 ( .A(n256), .B(n257), .Z(n258) );
  XOR U355 ( .A(n259), .B(n258), .Z(n300) );
  XOR U356 ( .A(n301), .B(n300), .Z(c[120]) );
  NANDN U357 ( .A(n257), .B(n256), .Z(n261) );
  NAND U358 ( .A(n259), .B(n258), .Z(n260) );
  NAND U359 ( .A(n261), .B(n260), .Z(n312) );
  NAND U360 ( .A(b[0]), .B(a[9]), .Z(n262) );
  XNOR U361 ( .A(b[1]), .B(n262), .Z(n264) );
  NAND U362 ( .A(a[8]), .B(n72), .Z(n263) );
  AND U363 ( .A(n264), .B(n263), .Z(n326) );
  NAND U364 ( .A(n9484), .B(n265), .Z(n267) );
  IV U365 ( .A(a[7]), .Z(n1075) );
  XNOR U366 ( .A(b[3]), .B(n1075), .Z(n339) );
  NAND U367 ( .A(n339), .B(n9485), .Z(n266) );
  AND U368 ( .A(n267), .B(n266), .Z(n325) );
  XNOR U369 ( .A(n326), .B(n325), .Z(n327) );
  XOR U370 ( .A(b[7]), .B(a[3]), .Z(n345) );
  NAND U371 ( .A(n345), .B(n9746), .Z(n270) );
  NANDN U372 ( .A(n268), .B(n9747), .Z(n269) );
  NAND U373 ( .A(n270), .B(n269), .Z(n331) );
  XNOR U374 ( .A(b[9]), .B(n628), .Z(n333) );
  NAND U375 ( .A(n9865), .B(n333), .Z(n274) );
  XOR U376 ( .A(b[9]), .B(a[0]), .Z(n391) );
  XOR U377 ( .A(b[9]), .B(b[7]), .Z(n272) );
  XOR U378 ( .A(b[9]), .B(b[8]), .Z(n271) );
  AND U379 ( .A(n272), .B(n271), .Z(n9930) );
  NAND U380 ( .A(n391), .B(n9930), .Z(n273) );
  AND U381 ( .A(n274), .B(n273), .Z(n332) );
  XNOR U382 ( .A(n331), .B(n332), .Z(n322) );
  ANDN U383 ( .B(n9872), .A(b[8]), .Z(n275) );
  NAND U384 ( .A(b[9]), .B(n275), .Z(n277) );
  AND U385 ( .A(n9865), .B(b[9]), .Z(n9932) );
  NAND U386 ( .A(n646), .B(n9932), .Z(n276) );
  NAND U387 ( .A(n277), .B(n276), .Z(n320) );
  IV U388 ( .A(a[5]), .Z(n894) );
  XNOR U389 ( .A(b[5]), .B(n894), .Z(n336) );
  NANDN U390 ( .A(n9623), .B(n336), .Z(n280) );
  NAND U391 ( .A(n278), .B(n9680), .Z(n279) );
  NAND U392 ( .A(n280), .B(n279), .Z(n319) );
  XOR U393 ( .A(n320), .B(n319), .Z(n321) );
  XOR U394 ( .A(n322), .B(n321), .Z(n328) );
  XOR U395 ( .A(n327), .B(n328), .Z(n316) );
  NANDN U396 ( .A(n282), .B(n281), .Z(n286) );
  NANDN U397 ( .A(n284), .B(n283), .Z(n285) );
  NAND U398 ( .A(n286), .B(n285), .Z(n313) );
  NANDN U399 ( .A(n288), .B(n287), .Z(n292) );
  NAND U400 ( .A(n290), .B(n289), .Z(n291) );
  NAND U401 ( .A(n292), .B(n291), .Z(n314) );
  XNOR U402 ( .A(n313), .B(n314), .Z(n315) );
  XNOR U403 ( .A(n316), .B(n315), .Z(n309) );
  NANDN U404 ( .A(n294), .B(n293), .Z(n298) );
  NAND U405 ( .A(n296), .B(n295), .Z(n297) );
  AND U406 ( .A(n298), .B(n297), .Z(n310) );
  XOR U407 ( .A(n309), .B(n310), .Z(n311) );
  XOR U408 ( .A(n312), .B(n311), .Z(n304) );
  XNOR U409 ( .A(n304), .B(sreg[121]), .Z(n306) );
  NAND U410 ( .A(n299), .B(sreg[120]), .Z(n303) );
  OR U411 ( .A(n301), .B(n300), .Z(n302) );
  AND U412 ( .A(n303), .B(n302), .Z(n305) );
  XOR U413 ( .A(n306), .B(n305), .Z(c[121]) );
  NAND U414 ( .A(n304), .B(sreg[121]), .Z(n308) );
  OR U415 ( .A(n306), .B(n305), .Z(n307) );
  NAND U416 ( .A(n308), .B(n307), .Z(n400) );
  XNOR U417 ( .A(n400), .B(sreg[122]), .Z(n402) );
  NANDN U418 ( .A(n314), .B(n313), .Z(n318) );
  NAND U419 ( .A(n316), .B(n315), .Z(n317) );
  NAND U420 ( .A(n318), .B(n317), .Z(n349) );
  OR U421 ( .A(n320), .B(n319), .Z(n324) );
  NANDN U422 ( .A(n322), .B(n321), .Z(n323) );
  NAND U423 ( .A(n324), .B(n323), .Z(n356) );
  NANDN U424 ( .A(n326), .B(n325), .Z(n330) );
  NANDN U425 ( .A(n328), .B(n327), .Z(n329) );
  NAND U426 ( .A(n330), .B(n329), .Z(n355) );
  NANDN U427 ( .A(n332), .B(n331), .Z(n375) );
  NAND U428 ( .A(n9930), .B(n333), .Z(n335) );
  XOR U429 ( .A(b[9]), .B(a[2]), .Z(n386) );
  NAND U430 ( .A(n9865), .B(n386), .Z(n334) );
  NAND U431 ( .A(n335), .B(n334), .Z(n373) );
  NAND U432 ( .A(n9680), .B(n336), .Z(n338) );
  XNOR U433 ( .A(b[5]), .B(n970), .Z(n397) );
  NANDN U434 ( .A(n9623), .B(n397), .Z(n337) );
  AND U435 ( .A(n338), .B(n337), .Z(n372) );
  XNOR U436 ( .A(n373), .B(n372), .Z(n374) );
  XNOR U437 ( .A(n375), .B(n374), .Z(n361) );
  NAND U438 ( .A(n9484), .B(n339), .Z(n341) );
  XOR U439 ( .A(b[3]), .B(a[8]), .Z(n383) );
  NAND U440 ( .A(n383), .B(n9485), .Z(n340) );
  AND U441 ( .A(n341), .B(n340), .Z(n360) );
  XNOR U442 ( .A(n361), .B(n360), .Z(n362) );
  XNOR U443 ( .A(b[9]), .B(b[10]), .Z(n10020) );
  ANDN U444 ( .B(a[0]), .A(n10020), .Z(n369) );
  NAND U445 ( .A(b[0]), .B(a[10]), .Z(n342) );
  XNOR U446 ( .A(b[1]), .B(n342), .Z(n344) );
  NAND U447 ( .A(a[9]), .B(n72), .Z(n343) );
  AND U448 ( .A(n344), .B(n343), .Z(n367) );
  XNOR U449 ( .A(n9872), .B(n834), .Z(n378) );
  NANDN U450 ( .A(n378), .B(n9746), .Z(n347) );
  NAND U451 ( .A(n345), .B(n9747), .Z(n346) );
  AND U452 ( .A(n347), .B(n346), .Z(n366) );
  XNOR U453 ( .A(n367), .B(n366), .Z(n368) );
  XOR U454 ( .A(n369), .B(n368), .Z(n363) );
  XNOR U455 ( .A(n362), .B(n363), .Z(n354) );
  XNOR U456 ( .A(n355), .B(n354), .Z(n357) );
  XNOR U457 ( .A(n356), .B(n357), .Z(n348) );
  XNOR U458 ( .A(n349), .B(n348), .Z(n350) );
  XOR U459 ( .A(n351), .B(n350), .Z(n401) );
  XOR U460 ( .A(n402), .B(n401), .Z(c[122]) );
  NANDN U461 ( .A(n349), .B(n348), .Z(n353) );
  NAND U462 ( .A(n351), .B(n350), .Z(n352) );
  NAND U463 ( .A(n353), .B(n352), .Z(n413) );
  NAND U464 ( .A(n355), .B(n354), .Z(n359) );
  NANDN U465 ( .A(n357), .B(n356), .Z(n358) );
  NAND U466 ( .A(n359), .B(n358), .Z(n411) );
  NANDN U467 ( .A(n361), .B(n360), .Z(n365) );
  NANDN U468 ( .A(n363), .B(n362), .Z(n364) );
  NAND U469 ( .A(n365), .B(n364), .Z(n418) );
  NANDN U470 ( .A(n367), .B(n366), .Z(n371) );
  NANDN U471 ( .A(n369), .B(n368), .Z(n370) );
  NAND U472 ( .A(n371), .B(n370), .Z(n417) );
  NANDN U473 ( .A(n373), .B(n372), .Z(n377) );
  NAND U474 ( .A(n375), .B(n374), .Z(n376) );
  NAND U475 ( .A(n377), .B(n376), .Z(n454) );
  XNOR U476 ( .A(n9872), .B(n894), .Z(n436) );
  NANDN U477 ( .A(n436), .B(n9746), .Z(n380) );
  NANDN U478 ( .A(n378), .B(n9747), .Z(n379) );
  NAND U479 ( .A(n380), .B(n379), .Z(n425) );
  IV U480 ( .A(b[9]), .Z(n9984) );
  ANDN U481 ( .B(n9984), .A(b[10]), .Z(n381) );
  NANDN U482 ( .A(n381), .B(a[0]), .Z(n382) );
  NAND U483 ( .A(b[9]), .B(b[10]), .Z(n10018) );
  IV U484 ( .A(b[11]), .Z(n9967) );
  ANDN U485 ( .B(n10018), .A(n9967), .Z(n10078) );
  NAND U486 ( .A(n382), .B(n10078), .Z(n422) );
  IV U487 ( .A(a[9]), .Z(n1204) );
  XNOR U488 ( .A(b[3]), .B(n1204), .Z(n439) );
  NAND U489 ( .A(n439), .B(n9485), .Z(n385) );
  NAND U490 ( .A(n383), .B(n9484), .Z(n384) );
  NAND U491 ( .A(n385), .B(n384), .Z(n423) );
  XOR U492 ( .A(n422), .B(n423), .Z(n424) );
  XNOR U493 ( .A(n425), .B(n424), .Z(n455) );
  XNOR U494 ( .A(n454), .B(n455), .Z(n456) );
  XNOR U495 ( .A(n9984), .B(n754), .Z(n445) );
  NANDN U496 ( .A(n445), .B(n9865), .Z(n388) );
  NAND U497 ( .A(n386), .B(n9930), .Z(n387) );
  NAND U498 ( .A(n388), .B(n387), .Z(n435) );
  XOR U499 ( .A(b[11]), .B(b[9]), .Z(n390) );
  XOR U500 ( .A(b[11]), .B(b[10]), .Z(n389) );
  AND U501 ( .A(n390), .B(n389), .Z(n9968) );
  NANDN U502 ( .A(n391), .B(n9968), .Z(n393) );
  XNOR U503 ( .A(n9967), .B(n628), .Z(n431) );
  OR U504 ( .A(n431), .B(n10020), .Z(n392) );
  NAND U505 ( .A(n393), .B(n392), .Z(n434) );
  XNOR U506 ( .A(n435), .B(n434), .Z(n451) );
  NAND U507 ( .A(b[0]), .B(a[11]), .Z(n394) );
  XNOR U508 ( .A(b[1]), .B(n394), .Z(n396) );
  NAND U509 ( .A(a[10]), .B(n72), .Z(n395) );
  AND U510 ( .A(n396), .B(n395), .Z(n449) );
  NAND U511 ( .A(n9680), .B(n397), .Z(n399) );
  XNOR U512 ( .A(b[5]), .B(n1075), .Z(n428) );
  NANDN U513 ( .A(n9623), .B(n428), .Z(n398) );
  AND U514 ( .A(n399), .B(n398), .Z(n448) );
  XNOR U515 ( .A(n449), .B(n448), .Z(n450) );
  XOR U516 ( .A(n451), .B(n450), .Z(n457) );
  XOR U517 ( .A(n456), .B(n457), .Z(n416) );
  XNOR U518 ( .A(n417), .B(n416), .Z(n419) );
  XNOR U519 ( .A(n418), .B(n419), .Z(n410) );
  XOR U520 ( .A(n411), .B(n410), .Z(n412) );
  XNOR U521 ( .A(n413), .B(n412), .Z(n405) );
  XNOR U522 ( .A(n405), .B(sreg[123]), .Z(n407) );
  NAND U523 ( .A(n400), .B(sreg[122]), .Z(n404) );
  OR U524 ( .A(n402), .B(n401), .Z(n403) );
  AND U525 ( .A(n404), .B(n403), .Z(n406) );
  XOR U526 ( .A(n407), .B(n406), .Z(c[123]) );
  NAND U527 ( .A(n405), .B(sreg[123]), .Z(n409) );
  OR U528 ( .A(n407), .B(n406), .Z(n408) );
  NAND U529 ( .A(n409), .B(n408), .Z(n520) );
  XNOR U530 ( .A(n520), .B(sreg[124]), .Z(n522) );
  NAND U531 ( .A(n411), .B(n410), .Z(n415) );
  NAND U532 ( .A(n413), .B(n412), .Z(n414) );
  NAND U533 ( .A(n415), .B(n414), .Z(n463) );
  NAND U534 ( .A(n417), .B(n416), .Z(n421) );
  NANDN U535 ( .A(n419), .B(n418), .Z(n420) );
  NAND U536 ( .A(n421), .B(n420), .Z(n460) );
  NANDN U537 ( .A(n423), .B(n422), .Z(n427) );
  OR U538 ( .A(n425), .B(n424), .Z(n426) );
  NAND U539 ( .A(n427), .B(n426), .Z(n469) );
  NAND U540 ( .A(n9680), .B(n428), .Z(n430) );
  IV U541 ( .A(a[8]), .Z(n1126) );
  XNOR U542 ( .A(b[5]), .B(n1126), .Z(n503) );
  NANDN U543 ( .A(n9623), .B(n503), .Z(n429) );
  NAND U544 ( .A(n430), .B(n429), .Z(n473) );
  XNOR U545 ( .A(n9967), .B(n705), .Z(n506) );
  OR U546 ( .A(n506), .B(n10020), .Z(n433) );
  NANDN U547 ( .A(n431), .B(n9968), .Z(n432) );
  NAND U548 ( .A(n433), .B(n432), .Z(n472) );
  XOR U549 ( .A(n473), .B(n472), .Z(n474) );
  NAND U550 ( .A(n435), .B(n434), .Z(n485) );
  XNOR U551 ( .A(n9872), .B(n970), .Z(n517) );
  NANDN U552 ( .A(n517), .B(n9746), .Z(n438) );
  NANDN U553 ( .A(n436), .B(n9747), .Z(n437) );
  NAND U554 ( .A(n438), .B(n437), .Z(n483) );
  NAND U555 ( .A(n9484), .B(n439), .Z(n441) );
  XOR U556 ( .A(b[3]), .B(a[10]), .Z(n497) );
  NAND U557 ( .A(n497), .B(n9485), .Z(n440) );
  AND U558 ( .A(n441), .B(n440), .Z(n482) );
  XNOR U559 ( .A(n483), .B(n482), .Z(n484) );
  XNOR U560 ( .A(n485), .B(n484), .Z(n475) );
  XNOR U561 ( .A(n474), .B(n475), .Z(n478) );
  XOR U562 ( .A(n9967), .B(b[12]), .Z(n10051) );
  ANDN U563 ( .B(a[0]), .A(n10051), .Z(n491) );
  NAND U564 ( .A(b[0]), .B(a[12]), .Z(n442) );
  XNOR U565 ( .A(b[1]), .B(n442), .Z(n444) );
  NAND U566 ( .A(a[11]), .B(n72), .Z(n443) );
  AND U567 ( .A(n444), .B(n443), .Z(n489) );
  NANDN U568 ( .A(n445), .B(n9930), .Z(n447) );
  XOR U569 ( .A(b[9]), .B(a[4]), .Z(n500) );
  NAND U570 ( .A(n9865), .B(n500), .Z(n446) );
  AND U571 ( .A(n447), .B(n446), .Z(n488) );
  XNOR U572 ( .A(n489), .B(n488), .Z(n490) );
  XOR U573 ( .A(n491), .B(n490), .Z(n476) );
  NANDN U574 ( .A(n449), .B(n448), .Z(n453) );
  NAND U575 ( .A(n451), .B(n450), .Z(n452) );
  NAND U576 ( .A(n453), .B(n452), .Z(n477) );
  XOR U577 ( .A(n476), .B(n477), .Z(n479) );
  XOR U578 ( .A(n478), .B(n479), .Z(n467) );
  NANDN U579 ( .A(n455), .B(n454), .Z(n459) );
  NAND U580 ( .A(n457), .B(n456), .Z(n458) );
  AND U581 ( .A(n459), .B(n458), .Z(n466) );
  XOR U582 ( .A(n467), .B(n466), .Z(n468) );
  XNOR U583 ( .A(n469), .B(n468), .Z(n461) );
  XNOR U584 ( .A(n460), .B(n461), .Z(n462) );
  XOR U585 ( .A(n463), .B(n462), .Z(n521) );
  XOR U586 ( .A(n522), .B(n521), .Z(c[124]) );
  NANDN U587 ( .A(n461), .B(n460), .Z(n465) );
  NAND U588 ( .A(n463), .B(n462), .Z(n464) );
  NAND U589 ( .A(n465), .B(n464), .Z(n533) );
  OR U590 ( .A(n467), .B(n466), .Z(n471) );
  NAND U591 ( .A(n469), .B(n468), .Z(n470) );
  NAND U592 ( .A(n471), .B(n470), .Z(n531) );
  NANDN U593 ( .A(n477), .B(n476), .Z(n481) );
  OR U594 ( .A(n479), .B(n478), .Z(n480) );
  NAND U595 ( .A(n481), .B(n480), .Z(n537) );
  XNOR U596 ( .A(n536), .B(n537), .Z(n538) );
  NANDN U597 ( .A(n483), .B(n482), .Z(n487) );
  NAND U598 ( .A(n485), .B(n484), .Z(n486) );
  NAND U599 ( .A(n487), .B(n486), .Z(n577) );
  NANDN U600 ( .A(n489), .B(n488), .Z(n493) );
  NANDN U601 ( .A(n491), .B(n490), .Z(n492) );
  AND U602 ( .A(n493), .B(n492), .Z(n578) );
  XNOR U603 ( .A(n577), .B(n578), .Z(n579) );
  NOR U604 ( .A(b[11]), .B(b[12]), .Z(n494) );
  NAND U605 ( .A(b[13]), .B(n494), .Z(n496) );
  IV U606 ( .A(b[13]), .Z(n10050) );
  NOR U607 ( .A(n10050), .B(n10051), .Z(n10073) );
  NAND U608 ( .A(n646), .B(n10073), .Z(n495) );
  NAND U609 ( .A(n496), .B(n495), .Z(n558) );
  IV U610 ( .A(a[11]), .Z(n1360) );
  XNOR U611 ( .A(n74), .B(n1360), .Z(n574) );
  NANDN U612 ( .A(n574), .B(n9485), .Z(n499) );
  NAND U613 ( .A(n497), .B(n9484), .Z(n498) );
  NAND U614 ( .A(n499), .B(n498), .Z(n556) );
  XNOR U615 ( .A(b[9]), .B(n894), .Z(n544) );
  NAND U616 ( .A(n9865), .B(n544), .Z(n502) );
  NAND U617 ( .A(n500), .B(n9930), .Z(n501) );
  AND U618 ( .A(n502), .B(n501), .Z(n557) );
  XNOR U619 ( .A(n556), .B(n557), .Z(n559) );
  XOR U620 ( .A(n558), .B(n559), .Z(n583) );
  NAND U621 ( .A(n9680), .B(n503), .Z(n505) );
  XOR U622 ( .A(b[5]), .B(a[9]), .Z(n568) );
  NANDN U623 ( .A(n9623), .B(n568), .Z(n504) );
  NAND U624 ( .A(n505), .B(n504), .Z(n584) );
  XNOR U625 ( .A(n583), .B(n584), .Z(n586) );
  XOR U626 ( .A(b[11]), .B(a[3]), .Z(n565) );
  NANDN U627 ( .A(n10020), .B(n565), .Z(n508) );
  NANDN U628 ( .A(n506), .B(n9968), .Z(n507) );
  NAND U629 ( .A(n508), .B(n507), .Z(n543) );
  XNOR U630 ( .A(b[13]), .B(n628), .Z(n547) );
  ANDN U631 ( .B(n547), .A(n10051), .Z(n513) );
  XOR U632 ( .A(b[13]), .B(a[0]), .Z(n511) );
  XOR U633 ( .A(b[13]), .B(b[11]), .Z(n510) );
  XOR U634 ( .A(b[13]), .B(b[12]), .Z(n509) );
  AND U635 ( .A(n510), .B(n509), .Z(n10070) );
  NAND U636 ( .A(n511), .B(n10070), .Z(n512) );
  NANDN U637 ( .A(n513), .B(n512), .Z(n542) );
  XNOR U638 ( .A(n543), .B(n542), .Z(n553) );
  NAND U639 ( .A(b[0]), .B(a[13]), .Z(n514) );
  XNOR U640 ( .A(b[1]), .B(n514), .Z(n516) );
  NAND U641 ( .A(a[12]), .B(n72), .Z(n515) );
  AND U642 ( .A(n516), .B(n515), .Z(n551) );
  XOR U643 ( .A(b[7]), .B(a[7]), .Z(n571) );
  NAND U644 ( .A(n571), .B(n9746), .Z(n519) );
  NANDN U645 ( .A(n517), .B(n9747), .Z(n518) );
  AND U646 ( .A(n519), .B(n518), .Z(n550) );
  XNOR U647 ( .A(n551), .B(n550), .Z(n552) );
  XOR U648 ( .A(n553), .B(n552), .Z(n585) );
  XOR U649 ( .A(n579), .B(n580), .Z(n539) );
  XOR U650 ( .A(n538), .B(n539), .Z(n530) );
  XOR U651 ( .A(n531), .B(n530), .Z(n532) );
  XNOR U652 ( .A(n533), .B(n532), .Z(n525) );
  XNOR U653 ( .A(n525), .B(sreg[125]), .Z(n527) );
  NAND U654 ( .A(n520), .B(sreg[124]), .Z(n524) );
  OR U655 ( .A(n522), .B(n521), .Z(n523) );
  AND U656 ( .A(n524), .B(n523), .Z(n526) );
  XOR U657 ( .A(n527), .B(n526), .Z(c[125]) );
  NAND U658 ( .A(n525), .B(sreg[125]), .Z(n529) );
  OR U659 ( .A(n527), .B(n526), .Z(n528) );
  NAND U660 ( .A(n529), .B(n528), .Z(n660) );
  XNOR U661 ( .A(n660), .B(sreg[126]), .Z(n662) );
  NAND U662 ( .A(n531), .B(n530), .Z(n535) );
  NAND U663 ( .A(n533), .B(n532), .Z(n534) );
  NAND U664 ( .A(n535), .B(n534), .Z(n592) );
  NANDN U665 ( .A(n537), .B(n536), .Z(n541) );
  NAND U666 ( .A(n539), .B(n538), .Z(n540) );
  NAND U667 ( .A(n541), .B(n540), .Z(n589) );
  AND U668 ( .A(n543), .B(n542), .Z(n603) );
  NAND U669 ( .A(n9930), .B(n544), .Z(n546) );
  XNOR U670 ( .A(b[9]), .B(n970), .Z(n634) );
  NAND U671 ( .A(n9865), .B(n634), .Z(n545) );
  NAND U672 ( .A(n546), .B(n545), .Z(n602) );
  NAND U673 ( .A(n10070), .B(n547), .Z(n549) );
  XOR U674 ( .A(b[13]), .B(a[2]), .Z(n623) );
  NANDN U675 ( .A(n10051), .B(n623), .Z(n548) );
  AND U676 ( .A(n549), .B(n548), .Z(n601) );
  XNOR U677 ( .A(n602), .B(n601), .Z(n604) );
  XOR U678 ( .A(n603), .B(n604), .Z(n654) );
  NANDN U679 ( .A(n551), .B(n550), .Z(n555) );
  NAND U680 ( .A(n553), .B(n552), .Z(n554) );
  NAND U681 ( .A(n555), .B(n554), .Z(n655) );
  XOR U682 ( .A(n654), .B(n655), .Z(n657) );
  NANDN U683 ( .A(n557), .B(n556), .Z(n561) );
  NAND U684 ( .A(n559), .B(n558), .Z(n560) );
  NAND U685 ( .A(n561), .B(n560), .Z(n614) );
  ANDN U686 ( .B(a[0]), .A(n10106), .Z(n608) );
  NAND U687 ( .A(b[0]), .B(a[14]), .Z(n562) );
  XNOR U688 ( .A(b[1]), .B(n562), .Z(n564) );
  NAND U689 ( .A(a[13]), .B(n72), .Z(n563) );
  AND U690 ( .A(n564), .B(n563), .Z(n606) );
  XNOR U691 ( .A(n9967), .B(n834), .Z(n637) );
  OR U692 ( .A(n637), .B(n10020), .Z(n567) );
  NAND U693 ( .A(n565), .B(n9968), .Z(n566) );
  AND U694 ( .A(n567), .B(n566), .Z(n605) );
  XNOR U695 ( .A(n606), .B(n605), .Z(n607) );
  XOR U696 ( .A(n608), .B(n607), .Z(n611) );
  IV U697 ( .A(a[10]), .Z(n1282) );
  XNOR U698 ( .A(b[5]), .B(n1282), .Z(n640) );
  NANDN U699 ( .A(n9623), .B(n640), .Z(n570) );
  NAND U700 ( .A(n568), .B(n9680), .Z(n569) );
  NAND U701 ( .A(n570), .B(n569), .Z(n620) );
  XNOR U702 ( .A(n9872), .B(n1126), .Z(n651) );
  NANDN U703 ( .A(n651), .B(n9746), .Z(n573) );
  NAND U704 ( .A(n571), .B(n9747), .Z(n572) );
  NAND U705 ( .A(n573), .B(n572), .Z(n617) );
  IV U706 ( .A(a[12]), .Z(n1438) );
  XNOR U707 ( .A(b[3]), .B(n1438), .Z(n643) );
  NAND U708 ( .A(n643), .B(n9485), .Z(n576) );
  NANDN U709 ( .A(n574), .B(n9484), .Z(n575) );
  AND U710 ( .A(n576), .B(n575), .Z(n618) );
  XNOR U711 ( .A(n617), .B(n618), .Z(n619) );
  XNOR U712 ( .A(n620), .B(n619), .Z(n612) );
  XNOR U713 ( .A(n611), .B(n612), .Z(n613) );
  XNOR U714 ( .A(n614), .B(n613), .Z(n656) );
  XNOR U715 ( .A(n657), .B(n656), .Z(n598) );
  NANDN U716 ( .A(n578), .B(n577), .Z(n582) );
  NAND U717 ( .A(n580), .B(n579), .Z(n581) );
  NAND U718 ( .A(n582), .B(n581), .Z(n595) );
  OR U719 ( .A(n584), .B(n583), .Z(n588) );
  NANDN U720 ( .A(n586), .B(n585), .Z(n587) );
  AND U721 ( .A(n588), .B(n587), .Z(n596) );
  XNOR U722 ( .A(n595), .B(n596), .Z(n597) );
  XNOR U723 ( .A(n598), .B(n597), .Z(n590) );
  XNOR U724 ( .A(n589), .B(n590), .Z(n591) );
  XOR U725 ( .A(n592), .B(n591), .Z(n661) );
  XOR U726 ( .A(n662), .B(n661), .Z(c[126]) );
  NANDN U727 ( .A(n590), .B(n589), .Z(n594) );
  NAND U728 ( .A(n592), .B(n591), .Z(n593) );
  NAND U729 ( .A(n594), .B(n593), .Z(n673) );
  NANDN U730 ( .A(n596), .B(n595), .Z(n600) );
  NAND U731 ( .A(n598), .B(n597), .Z(n599) );
  NAND U732 ( .A(n600), .B(n599), .Z(n671) );
  NANDN U733 ( .A(n606), .B(n605), .Z(n610) );
  NANDN U734 ( .A(n608), .B(n607), .Z(n609) );
  AND U735 ( .A(n610), .B(n609), .Z(n681) );
  XNOR U736 ( .A(n680), .B(n681), .Z(n682) );
  NANDN U737 ( .A(n612), .B(n611), .Z(n616) );
  NAND U738 ( .A(n614), .B(n613), .Z(n615) );
  AND U739 ( .A(n616), .B(n615), .Z(n683) );
  XNOR U740 ( .A(n682), .B(n683), .Z(n677) );
  NANDN U741 ( .A(n618), .B(n617), .Z(n622) );
  NAND U742 ( .A(n620), .B(n619), .Z(n621) );
  NAND U743 ( .A(n622), .B(n621), .Z(n730) );
  XNOR U744 ( .A(n10050), .B(n754), .Z(n696) );
  OR U745 ( .A(n696), .B(n10051), .Z(n625) );
  NAND U746 ( .A(n623), .B(n10070), .Z(n624) );
  NAND U747 ( .A(n625), .B(n624), .Z(n716) );
  XOR U748 ( .A(b[15]), .B(a[0]), .Z(n627) );
  XOR U749 ( .A(b[15]), .B(b[13]), .Z(n10142) );
  XOR U750 ( .A(b[15]), .B(b[14]), .Z(n626) );
  AND U751 ( .A(n10142), .B(n626), .Z(n10107) );
  NAND U752 ( .A(n627), .B(n10107), .Z(n630) );
  XNOR U753 ( .A(n75), .B(n628), .Z(n706) );
  OR U754 ( .A(n706), .B(n10106), .Z(n629) );
  NAND U755 ( .A(n630), .B(n629), .Z(n715) );
  XNOR U756 ( .A(n716), .B(n715), .Z(n693) );
  NAND U757 ( .A(b[0]), .B(a[15]), .Z(n631) );
  XNOR U758 ( .A(b[1]), .B(n631), .Z(n633) );
  NAND U759 ( .A(a[14]), .B(n72), .Z(n632) );
  AND U760 ( .A(n633), .B(n632), .Z(n691) );
  NAND U761 ( .A(n9930), .B(n634), .Z(n636) );
  XNOR U762 ( .A(b[9]), .B(n1075), .Z(n720) );
  NAND U763 ( .A(n9865), .B(n720), .Z(n635) );
  AND U764 ( .A(n636), .B(n635), .Z(n690) );
  XNOR U765 ( .A(n691), .B(n690), .Z(n692) );
  XOR U766 ( .A(n693), .B(n692), .Z(n729) );
  XOR U767 ( .A(n730), .B(n729), .Z(n731) );
  XOR U768 ( .A(b[11]), .B(a[5]), .Z(n702) );
  NANDN U769 ( .A(n10020), .B(n702), .Z(n639) );
  NANDN U770 ( .A(n637), .B(n9968), .Z(n638) );
  NAND U771 ( .A(n639), .B(n638), .Z(n688) );
  NAND U772 ( .A(n9680), .B(n640), .Z(n642) );
  XOR U773 ( .A(b[5]), .B(a[11]), .Z(n709) );
  NANDN U774 ( .A(n9623), .B(n709), .Z(n641) );
  AND U775 ( .A(n642), .B(n641), .Z(n686) );
  NAND U776 ( .A(n9484), .B(n643), .Z(n645) );
  IV U777 ( .A(a[13]), .Z(n1516) );
  XNOR U778 ( .A(b[3]), .B(n1516), .Z(n717) );
  NAND U779 ( .A(n717), .B(n9485), .Z(n644) );
  NAND U780 ( .A(n645), .B(n644), .Z(n687) );
  XOR U781 ( .A(n686), .B(n687), .Z(n689) );
  XOR U782 ( .A(n688), .B(n689), .Z(n726) );
  AND U783 ( .A(a[0]), .B(b[13]), .Z(n650) );
  NAND U784 ( .A(n646), .B(n10050), .Z(n647) );
  NAND U785 ( .A(b[14]), .B(n647), .Z(n648) );
  AND U786 ( .A(n648), .B(b[15]), .Z(n649) );
  NANDN U787 ( .A(n650), .B(n649), .Z(n723) );
  XNOR U788 ( .A(n9872), .B(n1204), .Z(n712) );
  NANDN U789 ( .A(n712), .B(n9746), .Z(n653) );
  NANDN U790 ( .A(n651), .B(n9747), .Z(n652) );
  NAND U791 ( .A(n653), .B(n652), .Z(n724) );
  XNOR U792 ( .A(n723), .B(n724), .Z(n725) );
  XOR U793 ( .A(n726), .B(n725), .Z(n732) );
  XNOR U794 ( .A(n731), .B(n732), .Z(n674) );
  NANDN U795 ( .A(n655), .B(n654), .Z(n659) );
  OR U796 ( .A(n657), .B(n656), .Z(n658) );
  AND U797 ( .A(n659), .B(n658), .Z(n675) );
  XOR U798 ( .A(n674), .B(n675), .Z(n676) );
  XOR U799 ( .A(n677), .B(n676), .Z(n670) );
  XOR U800 ( .A(n671), .B(n670), .Z(n672) );
  XOR U801 ( .A(n673), .B(n672), .Z(n665) );
  XNOR U802 ( .A(n665), .B(sreg[127]), .Z(n667) );
  NAND U803 ( .A(n660), .B(sreg[126]), .Z(n664) );
  OR U804 ( .A(n662), .B(n661), .Z(n663) );
  AND U805 ( .A(n664), .B(n663), .Z(n666) );
  XOR U806 ( .A(n667), .B(n666), .Z(c[127]) );
  NAND U807 ( .A(n665), .B(sreg[127]), .Z(n669) );
  OR U808 ( .A(n667), .B(n666), .Z(n668) );
  NAND U809 ( .A(n669), .B(n668), .Z(n804) );
  XNOR U810 ( .A(n804), .B(sreg[128]), .Z(n806) );
  NAND U811 ( .A(n675), .B(n674), .Z(n679) );
  NANDN U812 ( .A(n677), .B(n676), .Z(n678) );
  NAND U813 ( .A(n679), .B(n678), .Z(n733) );
  NANDN U814 ( .A(n681), .B(n680), .Z(n685) );
  NAND U815 ( .A(n683), .B(n682), .Z(n684) );
  NAND U816 ( .A(n685), .B(n684), .Z(n742) );
  NANDN U817 ( .A(n691), .B(n690), .Z(n695) );
  NAND U818 ( .A(n693), .B(n692), .Z(n694) );
  AND U819 ( .A(n695), .B(n694), .Z(n794) );
  XNOR U820 ( .A(n10050), .B(n834), .Z(n782) );
  OR U821 ( .A(n782), .B(n10051), .Z(n698) );
  NANDN U822 ( .A(n696), .B(n10070), .Z(n697) );
  NAND U823 ( .A(n698), .B(n697), .Z(n791) );
  NAND U824 ( .A(b[0]), .B(a[16]), .Z(n699) );
  XNOR U825 ( .A(b[1]), .B(n699), .Z(n701) );
  NAND U826 ( .A(a[15]), .B(n72), .Z(n700) );
  AND U827 ( .A(n701), .B(n700), .Z(n788) );
  NAND U828 ( .A(b[15]), .B(a[0]), .Z(n789) );
  XNOR U829 ( .A(n788), .B(n789), .Z(n790) );
  XOR U830 ( .A(n791), .B(n790), .Z(n795) );
  XOR U831 ( .A(n794), .B(n795), .Z(n796) );
  XNOR U832 ( .A(n797), .B(n796), .Z(n801) );
  XNOR U833 ( .A(n9967), .B(n970), .Z(n751) );
  OR U834 ( .A(n751), .B(n10020), .Z(n704) );
  NAND U835 ( .A(n702), .B(n9968), .Z(n703) );
  NAND U836 ( .A(n704), .B(n703), .Z(n764) );
  XNOR U837 ( .A(n75), .B(n705), .Z(n755) );
  OR U838 ( .A(n755), .B(n10106), .Z(n708) );
  NANDN U839 ( .A(n706), .B(n10107), .Z(n707) );
  NAND U840 ( .A(n708), .B(n707), .Z(n761) );
  XNOR U841 ( .A(n9622), .B(n1438), .Z(n773) );
  OR U842 ( .A(n773), .B(n9623), .Z(n711) );
  NAND U843 ( .A(n709), .B(n9680), .Z(n710) );
  AND U844 ( .A(n711), .B(n710), .Z(n762) );
  XNOR U845 ( .A(n761), .B(n762), .Z(n763) );
  XNOR U846 ( .A(n764), .B(n763), .Z(n767) );
  XOR U847 ( .A(b[7]), .B(a[10]), .Z(n776) );
  NAND U848 ( .A(n776), .B(n9746), .Z(n714) );
  NANDN U849 ( .A(n712), .B(n9747), .Z(n713) );
  NAND U850 ( .A(n714), .B(n713), .Z(n768) );
  XOR U851 ( .A(n767), .B(n768), .Z(n770) );
  NAND U852 ( .A(n716), .B(n715), .Z(n748) );
  NAND U853 ( .A(n9484), .B(n717), .Z(n719) );
  XOR U854 ( .A(b[3]), .B(a[14]), .Z(n779) );
  NAND U855 ( .A(n779), .B(n9485), .Z(n718) );
  NAND U856 ( .A(n719), .B(n718), .Z(n746) );
  NAND U857 ( .A(n9930), .B(n720), .Z(n722) );
  XOR U858 ( .A(b[9]), .B(a[8]), .Z(n758) );
  NAND U859 ( .A(n9865), .B(n758), .Z(n721) );
  AND U860 ( .A(n722), .B(n721), .Z(n745) );
  XNOR U861 ( .A(n746), .B(n745), .Z(n747) );
  XNOR U862 ( .A(n748), .B(n747), .Z(n769) );
  XNOR U863 ( .A(n770), .B(n769), .Z(n798) );
  NANDN U864 ( .A(n724), .B(n723), .Z(n728) );
  NAND U865 ( .A(n726), .B(n725), .Z(n727) );
  NAND U866 ( .A(n728), .B(n727), .Z(n799) );
  XNOR U867 ( .A(n798), .B(n799), .Z(n800) );
  XNOR U868 ( .A(n801), .B(n800), .Z(n740) );
  XOR U869 ( .A(n740), .B(n739), .Z(n741) );
  XNOR U870 ( .A(n742), .B(n741), .Z(n734) );
  XNOR U871 ( .A(n733), .B(n734), .Z(n735) );
  XOR U872 ( .A(n736), .B(n735), .Z(n805) );
  XOR U873 ( .A(n806), .B(n805), .Z(c[128]) );
  NANDN U874 ( .A(n734), .B(n733), .Z(n738) );
  NAND U875 ( .A(n736), .B(n735), .Z(n737) );
  NAND U876 ( .A(n738), .B(n737), .Z(n812) );
  OR U877 ( .A(n740), .B(n739), .Z(n744) );
  NAND U878 ( .A(n742), .B(n741), .Z(n743) );
  NAND U879 ( .A(n744), .B(n743), .Z(n810) );
  NANDN U880 ( .A(n746), .B(n745), .Z(n750) );
  NAND U881 ( .A(n748), .B(n747), .Z(n749) );
  NAND U882 ( .A(n750), .B(n749), .Z(n825) );
  XNOR U883 ( .A(n9967), .B(n1075), .Z(n831) );
  OR U884 ( .A(n831), .B(n10020), .Z(n753) );
  NANDN U885 ( .A(n751), .B(n9968), .Z(n752) );
  NAND U886 ( .A(n753), .B(n752), .Z(n844) );
  XNOR U887 ( .A(n75), .B(n754), .Z(n835) );
  OR U888 ( .A(n835), .B(n10106), .Z(n757) );
  NANDN U889 ( .A(n755), .B(n10107), .Z(n756) );
  NAND U890 ( .A(n757), .B(n756), .Z(n841) );
  XNOR U891 ( .A(n9984), .B(n1204), .Z(n838) );
  NANDN U892 ( .A(n838), .B(n9865), .Z(n760) );
  NAND U893 ( .A(n758), .B(n9930), .Z(n759) );
  AND U894 ( .A(n760), .B(n759), .Z(n842) );
  XNOR U895 ( .A(n841), .B(n842), .Z(n843) );
  XOR U896 ( .A(n844), .B(n843), .Z(n826) );
  XNOR U897 ( .A(n825), .B(n826), .Z(n827) );
  NANDN U898 ( .A(n762), .B(n761), .Z(n766) );
  NAND U899 ( .A(n764), .B(n763), .Z(n765) );
  AND U900 ( .A(n766), .B(n765), .Z(n828) );
  XNOR U901 ( .A(n827), .B(n828), .Z(n822) );
  NANDN U902 ( .A(n768), .B(n767), .Z(n772) );
  OR U903 ( .A(n770), .B(n769), .Z(n771) );
  NAND U904 ( .A(n772), .B(n771), .Z(n820) );
  XNOR U905 ( .A(n9622), .B(n1516), .Z(n867) );
  OR U906 ( .A(n867), .B(n9623), .Z(n775) );
  NANDN U907 ( .A(n773), .B(n9680), .Z(n774) );
  NAND U908 ( .A(n775), .B(n774), .Z(n850) );
  XNOR U909 ( .A(n9872), .B(n1360), .Z(n870) );
  NANDN U910 ( .A(n870), .B(n9746), .Z(n778) );
  NAND U911 ( .A(n776), .B(n9747), .Z(n777) );
  NAND U912 ( .A(n778), .B(n777), .Z(n847) );
  IV U913 ( .A(a[15]), .Z(n1672) );
  XNOR U914 ( .A(n74), .B(n1672), .Z(n873) );
  NANDN U915 ( .A(n873), .B(n9485), .Z(n781) );
  NAND U916 ( .A(n779), .B(n9484), .Z(n780) );
  AND U917 ( .A(n781), .B(n780), .Z(n848) );
  XNOR U918 ( .A(n847), .B(n848), .Z(n849) );
  XNOR U919 ( .A(n850), .B(n849), .Z(n856) );
  XNOR U920 ( .A(n10050), .B(n894), .Z(n864) );
  OR U921 ( .A(n864), .B(n10051), .Z(n784) );
  NANDN U922 ( .A(n782), .B(n10070), .Z(n783) );
  NAND U923 ( .A(n784), .B(n783), .Z(n860) );
  NAND U924 ( .A(b[0]), .B(a[17]), .Z(n785) );
  XNOR U925 ( .A(b[1]), .B(n785), .Z(n787) );
  NAND U926 ( .A(a[16]), .B(n72), .Z(n786) );
  AND U927 ( .A(n787), .B(n786), .Z(n857) );
  NAND U928 ( .A(b[15]), .B(a[1]), .Z(n858) );
  XOR U929 ( .A(n857), .B(n858), .Z(n859) );
  XOR U930 ( .A(n860), .B(n859), .Z(n853) );
  NANDN U931 ( .A(n789), .B(n788), .Z(n793) );
  NAND U932 ( .A(n791), .B(n790), .Z(n792) );
  NAND U933 ( .A(n793), .B(n792), .Z(n854) );
  XOR U934 ( .A(n853), .B(n854), .Z(n855) );
  XNOR U935 ( .A(n856), .B(n855), .Z(n819) );
  XOR U936 ( .A(n820), .B(n819), .Z(n821) );
  XOR U937 ( .A(n822), .B(n821), .Z(n817) );
  NANDN U938 ( .A(n799), .B(n798), .Z(n803) );
  NANDN U939 ( .A(n801), .B(n800), .Z(n802) );
  NAND U940 ( .A(n803), .B(n802), .Z(n816) );
  XNOR U941 ( .A(n815), .B(n816), .Z(n818) );
  XNOR U942 ( .A(n817), .B(n818), .Z(n809) );
  XOR U943 ( .A(n810), .B(n809), .Z(n811) );
  XNOR U944 ( .A(n812), .B(n811), .Z(n876) );
  XNOR U945 ( .A(n876), .B(sreg[129]), .Z(n878) );
  NAND U946 ( .A(n804), .B(sreg[128]), .Z(n808) );
  OR U947 ( .A(n806), .B(n805), .Z(n807) );
  AND U948 ( .A(n808), .B(n807), .Z(n877) );
  XOR U949 ( .A(n878), .B(n877), .Z(c[129]) );
  NAND U950 ( .A(n810), .B(n809), .Z(n814) );
  NAND U951 ( .A(n812), .B(n811), .Z(n813) );
  NAND U952 ( .A(n814), .B(n813), .Z(n884) );
  NAND U953 ( .A(n820), .B(n819), .Z(n824) );
  NANDN U954 ( .A(n822), .B(n821), .Z(n823) );
  NAND U955 ( .A(n824), .B(n823), .Z(n949) );
  NANDN U956 ( .A(n826), .B(n825), .Z(n830) );
  NAND U957 ( .A(n828), .B(n827), .Z(n829) );
  NAND U958 ( .A(n830), .B(n829), .Z(n946) );
  XNOR U959 ( .A(n9967), .B(n1126), .Z(n891) );
  OR U960 ( .A(n891), .B(n10020), .Z(n833) );
  NANDN U961 ( .A(n831), .B(n9968), .Z(n832) );
  NAND U962 ( .A(n833), .B(n832), .Z(n904) );
  XNOR U963 ( .A(n75), .B(n834), .Z(n895) );
  OR U964 ( .A(n895), .B(n10106), .Z(n837) );
  NANDN U965 ( .A(n835), .B(n10107), .Z(n836) );
  NAND U966 ( .A(n837), .B(n836), .Z(n901) );
  XNOR U967 ( .A(n9984), .B(n1282), .Z(n898) );
  NANDN U968 ( .A(n898), .B(n9865), .Z(n840) );
  NANDN U969 ( .A(n838), .B(n9930), .Z(n839) );
  AND U970 ( .A(n840), .B(n839), .Z(n902) );
  XNOR U971 ( .A(n901), .B(n902), .Z(n903) );
  XNOR U972 ( .A(n904), .B(n903), .Z(n940) );
  NANDN U973 ( .A(n842), .B(n841), .Z(n846) );
  NAND U974 ( .A(n844), .B(n843), .Z(n845) );
  NAND U975 ( .A(n846), .B(n845), .Z(n941) );
  XOR U976 ( .A(n940), .B(n941), .Z(n943) );
  NANDN U977 ( .A(n848), .B(n847), .Z(n852) );
  NAND U978 ( .A(n850), .B(n849), .Z(n851) );
  NAND U979 ( .A(n852), .B(n851), .Z(n942) );
  XNOR U980 ( .A(n943), .B(n942), .Z(n890) );
  NAND U981 ( .A(b[0]), .B(a[18]), .Z(n861) );
  XNOR U982 ( .A(b[1]), .B(n861), .Z(n863) );
  NAND U983 ( .A(a[17]), .B(n72), .Z(n862) );
  AND U984 ( .A(n863), .B(n862), .Z(n913) );
  XNOR U985 ( .A(n10050), .B(n970), .Z(n922) );
  OR U986 ( .A(n922), .B(n10051), .Z(n866) );
  NANDN U987 ( .A(n864), .B(n10070), .Z(n865) );
  AND U988 ( .A(n866), .B(n865), .Z(n914) );
  XOR U989 ( .A(n913), .B(n914), .Z(n916) );
  NAND U990 ( .A(a[2]), .B(b[15]), .Z(n915) );
  XOR U991 ( .A(n916), .B(n915), .Z(n934) );
  IV U992 ( .A(a[14]), .Z(n1621) );
  XNOR U993 ( .A(n9622), .B(n1621), .Z(n925) );
  OR U994 ( .A(n925), .B(n9623), .Z(n869) );
  NANDN U995 ( .A(n867), .B(n9680), .Z(n868) );
  NAND U996 ( .A(n869), .B(n868), .Z(n910) );
  XNOR U997 ( .A(n9872), .B(n1438), .Z(n928) );
  NANDN U998 ( .A(n928), .B(n9746), .Z(n872) );
  NANDN U999 ( .A(n870), .B(n9747), .Z(n871) );
  NAND U1000 ( .A(n872), .B(n871), .Z(n907) );
  IV U1001 ( .A(a[16]), .Z(n1750) );
  XNOR U1002 ( .A(n74), .B(n1750), .Z(n931) );
  NANDN U1003 ( .A(n931), .B(n9485), .Z(n875) );
  NANDN U1004 ( .A(n873), .B(n9484), .Z(n874) );
  AND U1005 ( .A(n875), .B(n874), .Z(n908) );
  XNOR U1006 ( .A(n907), .B(n908), .Z(n909) );
  XOR U1007 ( .A(n910), .B(n909), .Z(n935) );
  XOR U1008 ( .A(n934), .B(n935), .Z(n936) );
  XOR U1009 ( .A(n937), .B(n936), .Z(n887) );
  XOR U1010 ( .A(n888), .B(n887), .Z(n889) );
  XOR U1011 ( .A(n890), .B(n889), .Z(n947) );
  XOR U1012 ( .A(n946), .B(n947), .Z(n948) );
  XNOR U1013 ( .A(n949), .B(n948), .Z(n882) );
  XNOR U1014 ( .A(n881), .B(n882), .Z(n883) );
  XNOR U1015 ( .A(n884), .B(n883), .Z(n952) );
  XNOR U1016 ( .A(n952), .B(sreg[130]), .Z(n954) );
  NAND U1017 ( .A(n876), .B(sreg[129]), .Z(n880) );
  OR U1018 ( .A(n878), .B(n877), .Z(n879) );
  AND U1019 ( .A(n880), .B(n879), .Z(n953) );
  XOR U1020 ( .A(n954), .B(n953), .Z(c[130]) );
  NANDN U1021 ( .A(n882), .B(n881), .Z(n886) );
  NAND U1022 ( .A(n884), .B(n883), .Z(n885) );
  NAND U1023 ( .A(n886), .B(n885), .Z(n960) );
  XNOR U1024 ( .A(n9967), .B(n1204), .Z(n967) );
  OR U1025 ( .A(n967), .B(n10020), .Z(n893) );
  NANDN U1026 ( .A(n891), .B(n9968), .Z(n892) );
  NAND U1027 ( .A(n893), .B(n892), .Z(n980) );
  XNOR U1028 ( .A(n75), .B(n894), .Z(n971) );
  OR U1029 ( .A(n971), .B(n10106), .Z(n897) );
  NANDN U1030 ( .A(n895), .B(n10107), .Z(n896) );
  NAND U1031 ( .A(n897), .B(n896), .Z(n977) );
  XNOR U1032 ( .A(n9984), .B(n1360), .Z(n974) );
  NANDN U1033 ( .A(n974), .B(n9865), .Z(n900) );
  NANDN U1034 ( .A(n898), .B(n9930), .Z(n899) );
  AND U1035 ( .A(n900), .B(n899), .Z(n978) );
  XNOR U1036 ( .A(n977), .B(n978), .Z(n979) );
  XNOR U1037 ( .A(n980), .B(n979), .Z(n1016) );
  NANDN U1038 ( .A(n902), .B(n901), .Z(n906) );
  NAND U1039 ( .A(n904), .B(n903), .Z(n905) );
  NAND U1040 ( .A(n906), .B(n905), .Z(n1017) );
  XNOR U1041 ( .A(n1016), .B(n1017), .Z(n1018) );
  NANDN U1042 ( .A(n908), .B(n907), .Z(n912) );
  NAND U1043 ( .A(n910), .B(n909), .Z(n911) );
  AND U1044 ( .A(n912), .B(n911), .Z(n1019) );
  XNOR U1045 ( .A(n1018), .B(n1019), .Z(n963) );
  NANDN U1046 ( .A(n914), .B(n913), .Z(n918) );
  OR U1047 ( .A(n916), .B(n915), .Z(n917) );
  NAND U1048 ( .A(n918), .B(n917), .Z(n1013) );
  NAND U1049 ( .A(b[0]), .B(a[19]), .Z(n919) );
  XNOR U1050 ( .A(b[1]), .B(n919), .Z(n921) );
  NAND U1051 ( .A(a[18]), .B(n72), .Z(n920) );
  AND U1052 ( .A(n921), .B(n920), .Z(n989) );
  XNOR U1053 ( .A(n10050), .B(n1075), .Z(n998) );
  OR U1054 ( .A(n998), .B(n10051), .Z(n924) );
  NANDN U1055 ( .A(n922), .B(n10070), .Z(n923) );
  AND U1056 ( .A(n924), .B(n923), .Z(n990) );
  XOR U1057 ( .A(n989), .B(n990), .Z(n992) );
  NAND U1058 ( .A(a[3]), .B(b[15]), .Z(n991) );
  XOR U1059 ( .A(n992), .B(n991), .Z(n1010) );
  XNOR U1060 ( .A(n9622), .B(n1672), .Z(n1001) );
  OR U1061 ( .A(n1001), .B(n9623), .Z(n927) );
  NANDN U1062 ( .A(n925), .B(n9680), .Z(n926) );
  NAND U1063 ( .A(n927), .B(n926), .Z(n986) );
  XNOR U1064 ( .A(n9872), .B(n1516), .Z(n1004) );
  NANDN U1065 ( .A(n1004), .B(n9746), .Z(n930) );
  NANDN U1066 ( .A(n928), .B(n9747), .Z(n929) );
  NAND U1067 ( .A(n930), .B(n929), .Z(n983) );
  IV U1068 ( .A(a[17]), .Z(n1828) );
  XNOR U1069 ( .A(n74), .B(n1828), .Z(n1007) );
  NANDN U1070 ( .A(n1007), .B(n9485), .Z(n933) );
  NANDN U1071 ( .A(n931), .B(n9484), .Z(n932) );
  AND U1072 ( .A(n933), .B(n932), .Z(n984) );
  XNOR U1073 ( .A(n983), .B(n984), .Z(n985) );
  XOR U1074 ( .A(n986), .B(n985), .Z(n1011) );
  XOR U1075 ( .A(n1010), .B(n1011), .Z(n1012) );
  XNOR U1076 ( .A(n1013), .B(n1012), .Z(n961) );
  NAND U1077 ( .A(n935), .B(n934), .Z(n939) );
  NAND U1078 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1079 ( .A(n939), .B(n938), .Z(n962) );
  XOR U1080 ( .A(n961), .B(n962), .Z(n964) );
  XNOR U1081 ( .A(n963), .B(n964), .Z(n1022) );
  NANDN U1082 ( .A(n941), .B(n940), .Z(n945) );
  OR U1083 ( .A(n943), .B(n942), .Z(n944) );
  NAND U1084 ( .A(n945), .B(n944), .Z(n1023) );
  XNOR U1085 ( .A(n1022), .B(n1023), .Z(n1024) );
  XNOR U1086 ( .A(n1025), .B(n1024), .Z(n957) );
  OR U1087 ( .A(n947), .B(n946), .Z(n951) );
  NANDN U1088 ( .A(n949), .B(n948), .Z(n950) );
  NAND U1089 ( .A(n951), .B(n950), .Z(n958) );
  XOR U1090 ( .A(n957), .B(n958), .Z(n959) );
  XOR U1091 ( .A(n960), .B(n959), .Z(n1028) );
  XNOR U1092 ( .A(n1028), .B(sreg[131]), .Z(n1030) );
  NAND U1093 ( .A(n952), .B(sreg[130]), .Z(n956) );
  OR U1094 ( .A(n954), .B(n953), .Z(n955) );
  AND U1095 ( .A(n956), .B(n955), .Z(n1029) );
  XOR U1096 ( .A(n1030), .B(n1029), .Z(c[131]) );
  NANDN U1097 ( .A(n962), .B(n961), .Z(n966) );
  OR U1098 ( .A(n964), .B(n963), .Z(n965) );
  NAND U1099 ( .A(n966), .B(n965), .Z(n1103) );
  XNOR U1100 ( .A(n9967), .B(n1282), .Z(n1072) );
  OR U1101 ( .A(n1072), .B(n10020), .Z(n969) );
  NANDN U1102 ( .A(n967), .B(n9968), .Z(n968) );
  NAND U1103 ( .A(n969), .B(n968), .Z(n1085) );
  XNOR U1104 ( .A(n75), .B(n970), .Z(n1076) );
  OR U1105 ( .A(n1076), .B(n10106), .Z(n973) );
  NANDN U1106 ( .A(n971), .B(n10107), .Z(n972) );
  NAND U1107 ( .A(n973), .B(n972), .Z(n1082) );
  XNOR U1108 ( .A(n9984), .B(n1438), .Z(n1079) );
  NANDN U1109 ( .A(n1079), .B(n9865), .Z(n976) );
  NANDN U1110 ( .A(n974), .B(n9930), .Z(n975) );
  AND U1111 ( .A(n976), .B(n975), .Z(n1083) );
  XNOR U1112 ( .A(n1082), .B(n1083), .Z(n1084) );
  XNOR U1113 ( .A(n1085), .B(n1084), .Z(n1094) );
  NANDN U1114 ( .A(n978), .B(n977), .Z(n982) );
  NAND U1115 ( .A(n980), .B(n979), .Z(n981) );
  NAND U1116 ( .A(n982), .B(n981), .Z(n1095) );
  XNOR U1117 ( .A(n1094), .B(n1095), .Z(n1096) );
  NANDN U1118 ( .A(n984), .B(n983), .Z(n988) );
  NAND U1119 ( .A(n986), .B(n985), .Z(n987) );
  AND U1120 ( .A(n988), .B(n987), .Z(n1097) );
  XNOR U1121 ( .A(n1096), .B(n1097), .Z(n1041) );
  NANDN U1122 ( .A(n990), .B(n989), .Z(n994) );
  OR U1123 ( .A(n992), .B(n991), .Z(n993) );
  NAND U1124 ( .A(n994), .B(n993), .Z(n1069) );
  NAND U1125 ( .A(b[0]), .B(a[20]), .Z(n995) );
  XNOR U1126 ( .A(b[1]), .B(n995), .Z(n997) );
  NAND U1127 ( .A(a[19]), .B(n72), .Z(n996) );
  AND U1128 ( .A(n997), .B(n996), .Z(n1045) );
  XNOR U1129 ( .A(n10050), .B(n1126), .Z(n1054) );
  OR U1130 ( .A(n1054), .B(n10051), .Z(n1000) );
  NANDN U1131 ( .A(n998), .B(n10070), .Z(n999) );
  AND U1132 ( .A(n1000), .B(n999), .Z(n1046) );
  XOR U1133 ( .A(n1045), .B(n1046), .Z(n1048) );
  NAND U1134 ( .A(a[4]), .B(b[15]), .Z(n1047) );
  XOR U1135 ( .A(n1048), .B(n1047), .Z(n1066) );
  XNOR U1136 ( .A(n9622), .B(n1750), .Z(n1057) );
  OR U1137 ( .A(n1057), .B(n9623), .Z(n1003) );
  NANDN U1138 ( .A(n1001), .B(n9680), .Z(n1002) );
  NAND U1139 ( .A(n1003), .B(n1002), .Z(n1091) );
  XNOR U1140 ( .A(n9872), .B(n1621), .Z(n1060) );
  NANDN U1141 ( .A(n1060), .B(n9746), .Z(n1006) );
  NANDN U1142 ( .A(n1004), .B(n9747), .Z(n1005) );
  NAND U1143 ( .A(n1006), .B(n1005), .Z(n1088) );
  IV U1144 ( .A(a[18]), .Z(n1906) );
  XNOR U1145 ( .A(n74), .B(n1906), .Z(n1063) );
  NANDN U1146 ( .A(n1063), .B(n9485), .Z(n1009) );
  NANDN U1147 ( .A(n1007), .B(n9484), .Z(n1008) );
  AND U1148 ( .A(n1009), .B(n1008), .Z(n1089) );
  XNOR U1149 ( .A(n1088), .B(n1089), .Z(n1090) );
  XOR U1150 ( .A(n1091), .B(n1090), .Z(n1067) );
  XOR U1151 ( .A(n1066), .B(n1067), .Z(n1068) );
  XNOR U1152 ( .A(n1069), .B(n1068), .Z(n1039) );
  NAND U1153 ( .A(n1011), .B(n1010), .Z(n1015) );
  NAND U1154 ( .A(n1013), .B(n1012), .Z(n1014) );
  NAND U1155 ( .A(n1015), .B(n1014), .Z(n1040) );
  XOR U1156 ( .A(n1039), .B(n1040), .Z(n1042) );
  XNOR U1157 ( .A(n1041), .B(n1042), .Z(n1100) );
  NANDN U1158 ( .A(n1017), .B(n1016), .Z(n1021) );
  NAND U1159 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U1160 ( .A(n1021), .B(n1020), .Z(n1101) );
  XNOR U1161 ( .A(n1100), .B(n1101), .Z(n1102) );
  XOR U1162 ( .A(n1103), .B(n1102), .Z(n1033) );
  NANDN U1163 ( .A(n1023), .B(n1022), .Z(n1027) );
  NAND U1164 ( .A(n1025), .B(n1024), .Z(n1026) );
  NAND U1165 ( .A(n1027), .B(n1026), .Z(n1034) );
  XNOR U1166 ( .A(n1033), .B(n1034), .Z(n1035) );
  XNOR U1167 ( .A(n1036), .B(n1035), .Z(n1106) );
  XNOR U1168 ( .A(n1106), .B(sreg[132]), .Z(n1108) );
  NAND U1169 ( .A(n1028), .B(sreg[131]), .Z(n1032) );
  OR U1170 ( .A(n1030), .B(n1029), .Z(n1031) );
  AND U1171 ( .A(n1032), .B(n1031), .Z(n1107) );
  XOR U1172 ( .A(n1108), .B(n1107), .Z(c[132]) );
  NANDN U1173 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U1174 ( .A(n1036), .B(n1035), .Z(n1037) );
  NAND U1175 ( .A(n1038), .B(n1037), .Z(n1114) );
  NANDN U1176 ( .A(n1040), .B(n1039), .Z(n1044) );
  OR U1177 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1178 ( .A(n1044), .B(n1043), .Z(n1181) );
  NANDN U1179 ( .A(n1046), .B(n1045), .Z(n1050) );
  OR U1180 ( .A(n1048), .B(n1047), .Z(n1049) );
  NAND U1181 ( .A(n1050), .B(n1049), .Z(n1169) );
  NAND U1182 ( .A(b[0]), .B(a[21]), .Z(n1051) );
  XNOR U1183 ( .A(b[1]), .B(n1051), .Z(n1053) );
  NAND U1184 ( .A(a[20]), .B(n72), .Z(n1052) );
  AND U1185 ( .A(n1053), .B(n1052), .Z(n1145) );
  XNOR U1186 ( .A(n10050), .B(n1204), .Z(n1154) );
  OR U1187 ( .A(n1154), .B(n10051), .Z(n1056) );
  NANDN U1188 ( .A(n1054), .B(n10070), .Z(n1055) );
  AND U1189 ( .A(n1056), .B(n1055), .Z(n1146) );
  XOR U1190 ( .A(n1145), .B(n1146), .Z(n1148) );
  NAND U1191 ( .A(a[5]), .B(b[15]), .Z(n1147) );
  XOR U1192 ( .A(n1148), .B(n1147), .Z(n1166) );
  XNOR U1193 ( .A(n9622), .B(n1828), .Z(n1157) );
  OR U1194 ( .A(n1157), .B(n9623), .Z(n1059) );
  NANDN U1195 ( .A(n1057), .B(n9680), .Z(n1058) );
  NAND U1196 ( .A(n1059), .B(n1058), .Z(n1142) );
  XNOR U1197 ( .A(n9872), .B(n1672), .Z(n1160) );
  NANDN U1198 ( .A(n1160), .B(n9746), .Z(n1062) );
  NANDN U1199 ( .A(n1060), .B(n9747), .Z(n1061) );
  NAND U1200 ( .A(n1062), .B(n1061), .Z(n1139) );
  IV U1201 ( .A(a[19]), .Z(n1984) );
  XNOR U1202 ( .A(n74), .B(n1984), .Z(n1163) );
  NANDN U1203 ( .A(n1163), .B(n9485), .Z(n1065) );
  NANDN U1204 ( .A(n1063), .B(n9484), .Z(n1064) );
  AND U1205 ( .A(n1065), .B(n1064), .Z(n1140) );
  XNOR U1206 ( .A(n1139), .B(n1140), .Z(n1141) );
  XOR U1207 ( .A(n1142), .B(n1141), .Z(n1167) );
  XOR U1208 ( .A(n1166), .B(n1167), .Z(n1168) );
  XNOR U1209 ( .A(n1169), .B(n1168), .Z(n1117) );
  NAND U1210 ( .A(n1067), .B(n1066), .Z(n1071) );
  NAND U1211 ( .A(n1069), .B(n1068), .Z(n1070) );
  NAND U1212 ( .A(n1071), .B(n1070), .Z(n1118) );
  XOR U1213 ( .A(n1117), .B(n1118), .Z(n1120) );
  XNOR U1214 ( .A(n9967), .B(n1360), .Z(n1123) );
  OR U1215 ( .A(n1123), .B(n10020), .Z(n1074) );
  NANDN U1216 ( .A(n1072), .B(n9968), .Z(n1073) );
  NAND U1217 ( .A(n1074), .B(n1073), .Z(n1136) );
  XNOR U1218 ( .A(n75), .B(n1075), .Z(n1127) );
  OR U1219 ( .A(n1127), .B(n10106), .Z(n1078) );
  NANDN U1220 ( .A(n1076), .B(n10107), .Z(n1077) );
  NAND U1221 ( .A(n1078), .B(n1077), .Z(n1133) );
  XNOR U1222 ( .A(n9984), .B(n1516), .Z(n1130) );
  NANDN U1223 ( .A(n1130), .B(n9865), .Z(n1081) );
  NANDN U1224 ( .A(n1079), .B(n9930), .Z(n1080) );
  AND U1225 ( .A(n1081), .B(n1080), .Z(n1134) );
  XNOR U1226 ( .A(n1133), .B(n1134), .Z(n1135) );
  XNOR U1227 ( .A(n1136), .B(n1135), .Z(n1172) );
  NANDN U1228 ( .A(n1083), .B(n1082), .Z(n1087) );
  NAND U1229 ( .A(n1085), .B(n1084), .Z(n1086) );
  NAND U1230 ( .A(n1087), .B(n1086), .Z(n1173) );
  XNOR U1231 ( .A(n1172), .B(n1173), .Z(n1174) );
  NANDN U1232 ( .A(n1089), .B(n1088), .Z(n1093) );
  NAND U1233 ( .A(n1091), .B(n1090), .Z(n1092) );
  AND U1234 ( .A(n1093), .B(n1092), .Z(n1175) );
  XNOR U1235 ( .A(n1174), .B(n1175), .Z(n1119) );
  XNOR U1236 ( .A(n1120), .B(n1119), .Z(n1178) );
  NANDN U1237 ( .A(n1095), .B(n1094), .Z(n1099) );
  NAND U1238 ( .A(n1097), .B(n1096), .Z(n1098) );
  NAND U1239 ( .A(n1099), .B(n1098), .Z(n1179) );
  XNOR U1240 ( .A(n1178), .B(n1179), .Z(n1180) );
  XOR U1241 ( .A(n1181), .B(n1180), .Z(n1111) );
  NANDN U1242 ( .A(n1101), .B(n1100), .Z(n1105) );
  NANDN U1243 ( .A(n1103), .B(n1102), .Z(n1104) );
  NAND U1244 ( .A(n1105), .B(n1104), .Z(n1112) );
  XNOR U1245 ( .A(n1111), .B(n1112), .Z(n1113) );
  XNOR U1246 ( .A(n1114), .B(n1113), .Z(n1184) );
  XNOR U1247 ( .A(n1184), .B(sreg[133]), .Z(n1186) );
  NAND U1248 ( .A(n1106), .B(sreg[132]), .Z(n1110) );
  OR U1249 ( .A(n1108), .B(n1107), .Z(n1109) );
  AND U1250 ( .A(n1110), .B(n1109), .Z(n1185) );
  XOR U1251 ( .A(n1186), .B(n1185), .Z(c[133]) );
  NANDN U1252 ( .A(n1112), .B(n1111), .Z(n1116) );
  NAND U1253 ( .A(n1114), .B(n1113), .Z(n1115) );
  NAND U1254 ( .A(n1116), .B(n1115), .Z(n1192) );
  NANDN U1255 ( .A(n1118), .B(n1117), .Z(n1122) );
  OR U1256 ( .A(n1120), .B(n1119), .Z(n1121) );
  NAND U1257 ( .A(n1122), .B(n1121), .Z(n1259) );
  XNOR U1258 ( .A(n9967), .B(n1438), .Z(n1201) );
  OR U1259 ( .A(n1201), .B(n10020), .Z(n1125) );
  NANDN U1260 ( .A(n1123), .B(n9968), .Z(n1124) );
  NAND U1261 ( .A(n1125), .B(n1124), .Z(n1214) );
  XNOR U1262 ( .A(n75), .B(n1126), .Z(n1205) );
  OR U1263 ( .A(n1205), .B(n10106), .Z(n1129) );
  NANDN U1264 ( .A(n1127), .B(n10107), .Z(n1128) );
  NAND U1265 ( .A(n1129), .B(n1128), .Z(n1211) );
  XNOR U1266 ( .A(n9984), .B(n1621), .Z(n1208) );
  NANDN U1267 ( .A(n1208), .B(n9865), .Z(n1132) );
  NANDN U1268 ( .A(n1130), .B(n9930), .Z(n1131) );
  AND U1269 ( .A(n1132), .B(n1131), .Z(n1212) );
  XNOR U1270 ( .A(n1211), .B(n1212), .Z(n1213) );
  XNOR U1271 ( .A(n1214), .B(n1213), .Z(n1250) );
  NANDN U1272 ( .A(n1134), .B(n1133), .Z(n1138) );
  NAND U1273 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1274 ( .A(n1138), .B(n1137), .Z(n1251) );
  XNOR U1275 ( .A(n1250), .B(n1251), .Z(n1252) );
  NANDN U1276 ( .A(n1140), .B(n1139), .Z(n1144) );
  NAND U1277 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U1278 ( .A(n1144), .B(n1143), .Z(n1253) );
  XNOR U1279 ( .A(n1252), .B(n1253), .Z(n1197) );
  NANDN U1280 ( .A(n1146), .B(n1145), .Z(n1150) );
  OR U1281 ( .A(n1148), .B(n1147), .Z(n1149) );
  NAND U1282 ( .A(n1150), .B(n1149), .Z(n1247) );
  NAND U1283 ( .A(b[0]), .B(a[22]), .Z(n1151) );
  XNOR U1284 ( .A(b[1]), .B(n1151), .Z(n1153) );
  NAND U1285 ( .A(a[21]), .B(n72), .Z(n1152) );
  AND U1286 ( .A(n1153), .B(n1152), .Z(n1223) );
  XNOR U1287 ( .A(n10050), .B(n1282), .Z(n1232) );
  OR U1288 ( .A(n1232), .B(n10051), .Z(n1156) );
  NANDN U1289 ( .A(n1154), .B(n10070), .Z(n1155) );
  AND U1290 ( .A(n1156), .B(n1155), .Z(n1224) );
  XOR U1291 ( .A(n1223), .B(n1224), .Z(n1226) );
  NAND U1292 ( .A(a[6]), .B(b[15]), .Z(n1225) );
  XOR U1293 ( .A(n1226), .B(n1225), .Z(n1244) );
  XNOR U1294 ( .A(n9622), .B(n1906), .Z(n1235) );
  OR U1295 ( .A(n1235), .B(n9623), .Z(n1159) );
  NANDN U1296 ( .A(n1157), .B(n9680), .Z(n1158) );
  NAND U1297 ( .A(n1159), .B(n1158), .Z(n1220) );
  XNOR U1298 ( .A(n9872), .B(n1750), .Z(n1238) );
  NANDN U1299 ( .A(n1238), .B(n9746), .Z(n1162) );
  NANDN U1300 ( .A(n1160), .B(n9747), .Z(n1161) );
  NAND U1301 ( .A(n1162), .B(n1161), .Z(n1217) );
  IV U1302 ( .A(a[20]), .Z(n2062) );
  XNOR U1303 ( .A(n74), .B(n2062), .Z(n1241) );
  NANDN U1304 ( .A(n1241), .B(n9485), .Z(n1165) );
  NANDN U1305 ( .A(n1163), .B(n9484), .Z(n1164) );
  AND U1306 ( .A(n1165), .B(n1164), .Z(n1218) );
  XNOR U1307 ( .A(n1217), .B(n1218), .Z(n1219) );
  XOR U1308 ( .A(n1220), .B(n1219), .Z(n1245) );
  XOR U1309 ( .A(n1244), .B(n1245), .Z(n1246) );
  XNOR U1310 ( .A(n1247), .B(n1246), .Z(n1195) );
  NAND U1311 ( .A(n1167), .B(n1166), .Z(n1171) );
  NAND U1312 ( .A(n1169), .B(n1168), .Z(n1170) );
  NAND U1313 ( .A(n1171), .B(n1170), .Z(n1196) );
  XOR U1314 ( .A(n1195), .B(n1196), .Z(n1198) );
  XNOR U1315 ( .A(n1197), .B(n1198), .Z(n1256) );
  NANDN U1316 ( .A(n1173), .B(n1172), .Z(n1177) );
  NAND U1317 ( .A(n1175), .B(n1174), .Z(n1176) );
  NAND U1318 ( .A(n1177), .B(n1176), .Z(n1257) );
  XNOR U1319 ( .A(n1256), .B(n1257), .Z(n1258) );
  XOR U1320 ( .A(n1259), .B(n1258), .Z(n1189) );
  NANDN U1321 ( .A(n1179), .B(n1178), .Z(n1183) );
  NANDN U1322 ( .A(n1181), .B(n1180), .Z(n1182) );
  NAND U1323 ( .A(n1183), .B(n1182), .Z(n1190) );
  XNOR U1324 ( .A(n1189), .B(n1190), .Z(n1191) );
  XNOR U1325 ( .A(n1192), .B(n1191), .Z(n1262) );
  XNOR U1326 ( .A(n1262), .B(sreg[134]), .Z(n1264) );
  NAND U1327 ( .A(n1184), .B(sreg[133]), .Z(n1188) );
  OR U1328 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1329 ( .A(n1188), .B(n1187), .Z(n1263) );
  XOR U1330 ( .A(n1264), .B(n1263), .Z(c[134]) );
  NANDN U1331 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U1332 ( .A(n1192), .B(n1191), .Z(n1193) );
  NAND U1333 ( .A(n1194), .B(n1193), .Z(n1270) );
  NANDN U1334 ( .A(n1196), .B(n1195), .Z(n1200) );
  OR U1335 ( .A(n1198), .B(n1197), .Z(n1199) );
  NAND U1336 ( .A(n1200), .B(n1199), .Z(n1337) );
  XNOR U1337 ( .A(n9967), .B(n1516), .Z(n1279) );
  OR U1338 ( .A(n1279), .B(n10020), .Z(n1203) );
  NANDN U1339 ( .A(n1201), .B(n9968), .Z(n1202) );
  NAND U1340 ( .A(n1203), .B(n1202), .Z(n1292) );
  XNOR U1341 ( .A(n75), .B(n1204), .Z(n1283) );
  OR U1342 ( .A(n1283), .B(n10106), .Z(n1207) );
  NANDN U1343 ( .A(n1205), .B(n10107), .Z(n1206) );
  NAND U1344 ( .A(n1207), .B(n1206), .Z(n1289) );
  XNOR U1345 ( .A(n9984), .B(n1672), .Z(n1286) );
  NANDN U1346 ( .A(n1286), .B(n9865), .Z(n1210) );
  NANDN U1347 ( .A(n1208), .B(n9930), .Z(n1209) );
  AND U1348 ( .A(n1210), .B(n1209), .Z(n1290) );
  XNOR U1349 ( .A(n1289), .B(n1290), .Z(n1291) );
  XNOR U1350 ( .A(n1292), .B(n1291), .Z(n1328) );
  NANDN U1351 ( .A(n1212), .B(n1211), .Z(n1216) );
  NAND U1352 ( .A(n1214), .B(n1213), .Z(n1215) );
  NAND U1353 ( .A(n1216), .B(n1215), .Z(n1329) );
  XNOR U1354 ( .A(n1328), .B(n1329), .Z(n1330) );
  NANDN U1355 ( .A(n1218), .B(n1217), .Z(n1222) );
  NAND U1356 ( .A(n1220), .B(n1219), .Z(n1221) );
  AND U1357 ( .A(n1222), .B(n1221), .Z(n1331) );
  XNOR U1358 ( .A(n1330), .B(n1331), .Z(n1275) );
  NANDN U1359 ( .A(n1224), .B(n1223), .Z(n1228) );
  OR U1360 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1361 ( .A(n1228), .B(n1227), .Z(n1325) );
  NAND U1362 ( .A(b[0]), .B(a[23]), .Z(n1229) );
  XNOR U1363 ( .A(b[1]), .B(n1229), .Z(n1231) );
  NAND U1364 ( .A(a[22]), .B(n72), .Z(n1230) );
  AND U1365 ( .A(n1231), .B(n1230), .Z(n1301) );
  XNOR U1366 ( .A(n10050), .B(n1360), .Z(n1310) );
  OR U1367 ( .A(n1310), .B(n10051), .Z(n1234) );
  NANDN U1368 ( .A(n1232), .B(n10070), .Z(n1233) );
  AND U1369 ( .A(n1234), .B(n1233), .Z(n1302) );
  XOR U1370 ( .A(n1301), .B(n1302), .Z(n1304) );
  NAND U1371 ( .A(a[7]), .B(b[15]), .Z(n1303) );
  XOR U1372 ( .A(n1304), .B(n1303), .Z(n1322) );
  XNOR U1373 ( .A(n9622), .B(n1984), .Z(n1313) );
  OR U1374 ( .A(n1313), .B(n9623), .Z(n1237) );
  NANDN U1375 ( .A(n1235), .B(n9680), .Z(n1236) );
  NAND U1376 ( .A(n1237), .B(n1236), .Z(n1298) );
  XNOR U1377 ( .A(n9872), .B(n1828), .Z(n1316) );
  NANDN U1378 ( .A(n1316), .B(n9746), .Z(n1240) );
  NANDN U1379 ( .A(n1238), .B(n9747), .Z(n1239) );
  NAND U1380 ( .A(n1240), .B(n1239), .Z(n1295) );
  IV U1381 ( .A(a[21]), .Z(n2167) );
  XNOR U1382 ( .A(n74), .B(n2167), .Z(n1319) );
  NANDN U1383 ( .A(n1319), .B(n9485), .Z(n1243) );
  NANDN U1384 ( .A(n1241), .B(n9484), .Z(n1242) );
  AND U1385 ( .A(n1243), .B(n1242), .Z(n1296) );
  XNOR U1386 ( .A(n1295), .B(n1296), .Z(n1297) );
  XOR U1387 ( .A(n1298), .B(n1297), .Z(n1323) );
  XOR U1388 ( .A(n1322), .B(n1323), .Z(n1324) );
  XNOR U1389 ( .A(n1325), .B(n1324), .Z(n1273) );
  NAND U1390 ( .A(n1245), .B(n1244), .Z(n1249) );
  NAND U1391 ( .A(n1247), .B(n1246), .Z(n1248) );
  NAND U1392 ( .A(n1249), .B(n1248), .Z(n1274) );
  XOR U1393 ( .A(n1273), .B(n1274), .Z(n1276) );
  XNOR U1394 ( .A(n1275), .B(n1276), .Z(n1334) );
  NANDN U1395 ( .A(n1251), .B(n1250), .Z(n1255) );
  NAND U1396 ( .A(n1253), .B(n1252), .Z(n1254) );
  NAND U1397 ( .A(n1255), .B(n1254), .Z(n1335) );
  XNOR U1398 ( .A(n1334), .B(n1335), .Z(n1336) );
  XOR U1399 ( .A(n1337), .B(n1336), .Z(n1267) );
  NANDN U1400 ( .A(n1257), .B(n1256), .Z(n1261) );
  NANDN U1401 ( .A(n1259), .B(n1258), .Z(n1260) );
  NAND U1402 ( .A(n1261), .B(n1260), .Z(n1268) );
  XNOR U1403 ( .A(n1267), .B(n1268), .Z(n1269) );
  XNOR U1404 ( .A(n1270), .B(n1269), .Z(n1340) );
  XNOR U1405 ( .A(n1340), .B(sreg[135]), .Z(n1342) );
  NAND U1406 ( .A(n1262), .B(sreg[134]), .Z(n1266) );
  OR U1407 ( .A(n1264), .B(n1263), .Z(n1265) );
  AND U1408 ( .A(n1266), .B(n1265), .Z(n1341) );
  XOR U1409 ( .A(n1342), .B(n1341), .Z(c[135]) );
  NANDN U1410 ( .A(n1268), .B(n1267), .Z(n1272) );
  NAND U1411 ( .A(n1270), .B(n1269), .Z(n1271) );
  NAND U1412 ( .A(n1272), .B(n1271), .Z(n1348) );
  NANDN U1413 ( .A(n1274), .B(n1273), .Z(n1278) );
  OR U1414 ( .A(n1276), .B(n1275), .Z(n1277) );
  NAND U1415 ( .A(n1278), .B(n1277), .Z(n1415) );
  XNOR U1416 ( .A(n9967), .B(n1621), .Z(n1357) );
  OR U1417 ( .A(n1357), .B(n10020), .Z(n1281) );
  NANDN U1418 ( .A(n1279), .B(n9968), .Z(n1280) );
  NAND U1419 ( .A(n1281), .B(n1280), .Z(n1370) );
  XNOR U1420 ( .A(n75), .B(n1282), .Z(n1361) );
  OR U1421 ( .A(n1361), .B(n10106), .Z(n1285) );
  NANDN U1422 ( .A(n1283), .B(n10107), .Z(n1284) );
  NAND U1423 ( .A(n1285), .B(n1284), .Z(n1367) );
  XNOR U1424 ( .A(n9984), .B(n1750), .Z(n1364) );
  NANDN U1425 ( .A(n1364), .B(n9865), .Z(n1288) );
  NANDN U1426 ( .A(n1286), .B(n9930), .Z(n1287) );
  AND U1427 ( .A(n1288), .B(n1287), .Z(n1368) );
  XNOR U1428 ( .A(n1367), .B(n1368), .Z(n1369) );
  XNOR U1429 ( .A(n1370), .B(n1369), .Z(n1406) );
  NANDN U1430 ( .A(n1290), .B(n1289), .Z(n1294) );
  NAND U1431 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U1432 ( .A(n1294), .B(n1293), .Z(n1407) );
  XNOR U1433 ( .A(n1406), .B(n1407), .Z(n1408) );
  NANDN U1434 ( .A(n1296), .B(n1295), .Z(n1300) );
  NAND U1435 ( .A(n1298), .B(n1297), .Z(n1299) );
  AND U1436 ( .A(n1300), .B(n1299), .Z(n1409) );
  XNOR U1437 ( .A(n1408), .B(n1409), .Z(n1353) );
  NANDN U1438 ( .A(n1302), .B(n1301), .Z(n1306) );
  OR U1439 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1440 ( .A(n1306), .B(n1305), .Z(n1403) );
  NAND U1441 ( .A(b[0]), .B(a[24]), .Z(n1307) );
  XNOR U1442 ( .A(b[1]), .B(n1307), .Z(n1309) );
  NAND U1443 ( .A(a[23]), .B(n72), .Z(n1308) );
  AND U1444 ( .A(n1309), .B(n1308), .Z(n1379) );
  XNOR U1445 ( .A(n10050), .B(n1438), .Z(n1388) );
  OR U1446 ( .A(n1388), .B(n10051), .Z(n1312) );
  NANDN U1447 ( .A(n1310), .B(n10070), .Z(n1311) );
  AND U1448 ( .A(n1312), .B(n1311), .Z(n1380) );
  XOR U1449 ( .A(n1379), .B(n1380), .Z(n1382) );
  NAND U1450 ( .A(a[8]), .B(b[15]), .Z(n1381) );
  XOR U1451 ( .A(n1382), .B(n1381), .Z(n1400) );
  XNOR U1452 ( .A(n9622), .B(n2062), .Z(n1391) );
  OR U1453 ( .A(n1391), .B(n9623), .Z(n1315) );
  NANDN U1454 ( .A(n1313), .B(n9680), .Z(n1314) );
  NAND U1455 ( .A(n1315), .B(n1314), .Z(n1376) );
  XNOR U1456 ( .A(n9872), .B(n1906), .Z(n1394) );
  NANDN U1457 ( .A(n1394), .B(n9746), .Z(n1318) );
  NANDN U1458 ( .A(n1316), .B(n9747), .Z(n1317) );
  NAND U1459 ( .A(n1318), .B(n1317), .Z(n1373) );
  IV U1460 ( .A(a[22]), .Z(n2245) );
  XNOR U1461 ( .A(n74), .B(n2245), .Z(n1397) );
  NANDN U1462 ( .A(n1397), .B(n9485), .Z(n1321) );
  NANDN U1463 ( .A(n1319), .B(n9484), .Z(n1320) );
  AND U1464 ( .A(n1321), .B(n1320), .Z(n1374) );
  XNOR U1465 ( .A(n1373), .B(n1374), .Z(n1375) );
  XOR U1466 ( .A(n1376), .B(n1375), .Z(n1401) );
  XOR U1467 ( .A(n1400), .B(n1401), .Z(n1402) );
  XNOR U1468 ( .A(n1403), .B(n1402), .Z(n1351) );
  NAND U1469 ( .A(n1323), .B(n1322), .Z(n1327) );
  NAND U1470 ( .A(n1325), .B(n1324), .Z(n1326) );
  NAND U1471 ( .A(n1327), .B(n1326), .Z(n1352) );
  XOR U1472 ( .A(n1351), .B(n1352), .Z(n1354) );
  XNOR U1473 ( .A(n1353), .B(n1354), .Z(n1412) );
  NANDN U1474 ( .A(n1329), .B(n1328), .Z(n1333) );
  NAND U1475 ( .A(n1331), .B(n1330), .Z(n1332) );
  NAND U1476 ( .A(n1333), .B(n1332), .Z(n1413) );
  XNOR U1477 ( .A(n1412), .B(n1413), .Z(n1414) );
  XOR U1478 ( .A(n1415), .B(n1414), .Z(n1345) );
  NANDN U1479 ( .A(n1335), .B(n1334), .Z(n1339) );
  NANDN U1480 ( .A(n1337), .B(n1336), .Z(n1338) );
  NAND U1481 ( .A(n1339), .B(n1338), .Z(n1346) );
  XNOR U1482 ( .A(n1345), .B(n1346), .Z(n1347) );
  XNOR U1483 ( .A(n1348), .B(n1347), .Z(n1418) );
  XNOR U1484 ( .A(n1418), .B(sreg[136]), .Z(n1420) );
  NAND U1485 ( .A(n1340), .B(sreg[135]), .Z(n1344) );
  OR U1486 ( .A(n1342), .B(n1341), .Z(n1343) );
  AND U1487 ( .A(n1344), .B(n1343), .Z(n1419) );
  XOR U1488 ( .A(n1420), .B(n1419), .Z(c[136]) );
  NANDN U1489 ( .A(n1346), .B(n1345), .Z(n1350) );
  NAND U1490 ( .A(n1348), .B(n1347), .Z(n1349) );
  NAND U1491 ( .A(n1350), .B(n1349), .Z(n1426) );
  NANDN U1492 ( .A(n1352), .B(n1351), .Z(n1356) );
  OR U1493 ( .A(n1354), .B(n1353), .Z(n1355) );
  NAND U1494 ( .A(n1356), .B(n1355), .Z(n1493) );
  XNOR U1495 ( .A(n9967), .B(n1672), .Z(n1435) );
  OR U1496 ( .A(n1435), .B(n10020), .Z(n1359) );
  NANDN U1497 ( .A(n1357), .B(n9968), .Z(n1358) );
  NAND U1498 ( .A(n1359), .B(n1358), .Z(n1448) );
  XNOR U1499 ( .A(n75), .B(n1360), .Z(n1439) );
  OR U1500 ( .A(n1439), .B(n10106), .Z(n1363) );
  NANDN U1501 ( .A(n1361), .B(n10107), .Z(n1362) );
  NAND U1502 ( .A(n1363), .B(n1362), .Z(n1445) );
  XNOR U1503 ( .A(n9984), .B(n1828), .Z(n1442) );
  NANDN U1504 ( .A(n1442), .B(n9865), .Z(n1366) );
  NANDN U1505 ( .A(n1364), .B(n9930), .Z(n1365) );
  AND U1506 ( .A(n1366), .B(n1365), .Z(n1446) );
  XNOR U1507 ( .A(n1445), .B(n1446), .Z(n1447) );
  XNOR U1508 ( .A(n1448), .B(n1447), .Z(n1484) );
  NANDN U1509 ( .A(n1368), .B(n1367), .Z(n1372) );
  NAND U1510 ( .A(n1370), .B(n1369), .Z(n1371) );
  NAND U1511 ( .A(n1372), .B(n1371), .Z(n1485) );
  XNOR U1512 ( .A(n1484), .B(n1485), .Z(n1486) );
  NANDN U1513 ( .A(n1374), .B(n1373), .Z(n1378) );
  NAND U1514 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U1515 ( .A(n1378), .B(n1377), .Z(n1487) );
  XNOR U1516 ( .A(n1486), .B(n1487), .Z(n1431) );
  NANDN U1517 ( .A(n1380), .B(n1379), .Z(n1384) );
  OR U1518 ( .A(n1382), .B(n1381), .Z(n1383) );
  NAND U1519 ( .A(n1384), .B(n1383), .Z(n1481) );
  NAND U1520 ( .A(b[0]), .B(a[25]), .Z(n1385) );
  XNOR U1521 ( .A(b[1]), .B(n1385), .Z(n1387) );
  NAND U1522 ( .A(a[24]), .B(n72), .Z(n1386) );
  AND U1523 ( .A(n1387), .B(n1386), .Z(n1457) );
  XNOR U1524 ( .A(n10050), .B(n1516), .Z(n1463) );
  OR U1525 ( .A(n1463), .B(n10051), .Z(n1390) );
  NANDN U1526 ( .A(n1388), .B(n10070), .Z(n1389) );
  AND U1527 ( .A(n1390), .B(n1389), .Z(n1458) );
  XOR U1528 ( .A(n1457), .B(n1458), .Z(n1460) );
  NAND U1529 ( .A(a[9]), .B(b[15]), .Z(n1459) );
  XOR U1530 ( .A(n1460), .B(n1459), .Z(n1478) );
  XNOR U1531 ( .A(n9622), .B(n2167), .Z(n1469) );
  OR U1532 ( .A(n1469), .B(n9623), .Z(n1393) );
  NANDN U1533 ( .A(n1391), .B(n9680), .Z(n1392) );
  NAND U1534 ( .A(n1393), .B(n1392), .Z(n1454) );
  XNOR U1535 ( .A(n9872), .B(n1984), .Z(n1472) );
  NANDN U1536 ( .A(n1472), .B(n9746), .Z(n1396) );
  NANDN U1537 ( .A(n1394), .B(n9747), .Z(n1395) );
  NAND U1538 ( .A(n1396), .B(n1395), .Z(n1451) );
  IV U1539 ( .A(a[23]), .Z(n2323) );
  XNOR U1540 ( .A(n74), .B(n2323), .Z(n1475) );
  NANDN U1541 ( .A(n1475), .B(n9485), .Z(n1399) );
  NANDN U1542 ( .A(n1397), .B(n9484), .Z(n1398) );
  AND U1543 ( .A(n1399), .B(n1398), .Z(n1452) );
  XNOR U1544 ( .A(n1451), .B(n1452), .Z(n1453) );
  XOR U1545 ( .A(n1454), .B(n1453), .Z(n1479) );
  XOR U1546 ( .A(n1478), .B(n1479), .Z(n1480) );
  XNOR U1547 ( .A(n1481), .B(n1480), .Z(n1429) );
  NAND U1548 ( .A(n1401), .B(n1400), .Z(n1405) );
  NAND U1549 ( .A(n1403), .B(n1402), .Z(n1404) );
  NAND U1550 ( .A(n1405), .B(n1404), .Z(n1430) );
  XOR U1551 ( .A(n1429), .B(n1430), .Z(n1432) );
  XNOR U1552 ( .A(n1431), .B(n1432), .Z(n1490) );
  NANDN U1553 ( .A(n1407), .B(n1406), .Z(n1411) );
  NAND U1554 ( .A(n1409), .B(n1408), .Z(n1410) );
  NAND U1555 ( .A(n1411), .B(n1410), .Z(n1491) );
  XNOR U1556 ( .A(n1490), .B(n1491), .Z(n1492) );
  XOR U1557 ( .A(n1493), .B(n1492), .Z(n1423) );
  NANDN U1558 ( .A(n1413), .B(n1412), .Z(n1417) );
  NANDN U1559 ( .A(n1415), .B(n1414), .Z(n1416) );
  NAND U1560 ( .A(n1417), .B(n1416), .Z(n1424) );
  XNOR U1561 ( .A(n1423), .B(n1424), .Z(n1425) );
  XNOR U1562 ( .A(n1426), .B(n1425), .Z(n1496) );
  XNOR U1563 ( .A(n1496), .B(sreg[137]), .Z(n1498) );
  NAND U1564 ( .A(n1418), .B(sreg[136]), .Z(n1422) );
  OR U1565 ( .A(n1420), .B(n1419), .Z(n1421) );
  AND U1566 ( .A(n1422), .B(n1421), .Z(n1497) );
  XOR U1567 ( .A(n1498), .B(n1497), .Z(c[137]) );
  NANDN U1568 ( .A(n1424), .B(n1423), .Z(n1428) );
  NAND U1569 ( .A(n1426), .B(n1425), .Z(n1427) );
  NAND U1570 ( .A(n1428), .B(n1427), .Z(n1504) );
  NANDN U1571 ( .A(n1430), .B(n1429), .Z(n1434) );
  OR U1572 ( .A(n1432), .B(n1431), .Z(n1433) );
  NAND U1573 ( .A(n1434), .B(n1433), .Z(n1571) );
  XNOR U1574 ( .A(n9967), .B(n1750), .Z(n1513) );
  OR U1575 ( .A(n1513), .B(n10020), .Z(n1437) );
  NANDN U1576 ( .A(n1435), .B(n9968), .Z(n1436) );
  NAND U1577 ( .A(n1437), .B(n1436), .Z(n1526) );
  XNOR U1578 ( .A(n75), .B(n1438), .Z(n1517) );
  OR U1579 ( .A(n1517), .B(n10106), .Z(n1441) );
  NANDN U1580 ( .A(n1439), .B(n10107), .Z(n1440) );
  NAND U1581 ( .A(n1441), .B(n1440), .Z(n1523) );
  XNOR U1582 ( .A(n9984), .B(n1906), .Z(n1520) );
  NANDN U1583 ( .A(n1520), .B(n9865), .Z(n1444) );
  NANDN U1584 ( .A(n1442), .B(n9930), .Z(n1443) );
  AND U1585 ( .A(n1444), .B(n1443), .Z(n1524) );
  XNOR U1586 ( .A(n1523), .B(n1524), .Z(n1525) );
  XNOR U1587 ( .A(n1526), .B(n1525), .Z(n1562) );
  NANDN U1588 ( .A(n1446), .B(n1445), .Z(n1450) );
  NAND U1589 ( .A(n1448), .B(n1447), .Z(n1449) );
  NAND U1590 ( .A(n1450), .B(n1449), .Z(n1563) );
  XNOR U1591 ( .A(n1562), .B(n1563), .Z(n1564) );
  NANDN U1592 ( .A(n1452), .B(n1451), .Z(n1456) );
  NAND U1593 ( .A(n1454), .B(n1453), .Z(n1455) );
  AND U1594 ( .A(n1456), .B(n1455), .Z(n1565) );
  XNOR U1595 ( .A(n1564), .B(n1565), .Z(n1509) );
  NANDN U1596 ( .A(n1458), .B(n1457), .Z(n1462) );
  OR U1597 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1598 ( .A(n1462), .B(n1461), .Z(n1559) );
  XNOR U1599 ( .A(n10050), .B(n1621), .Z(n1544) );
  OR U1600 ( .A(n1544), .B(n10051), .Z(n1465) );
  NANDN U1601 ( .A(n1463), .B(n10070), .Z(n1464) );
  AND U1602 ( .A(n1465), .B(n1464), .Z(n1536) );
  NAND U1603 ( .A(b[0]), .B(a[26]), .Z(n1466) );
  XNOR U1604 ( .A(b[1]), .B(n1466), .Z(n1468) );
  NAND U1605 ( .A(a[25]), .B(n72), .Z(n1467) );
  AND U1606 ( .A(n1468), .B(n1467), .Z(n1535) );
  XOR U1607 ( .A(n1536), .B(n1535), .Z(n1538) );
  NAND U1608 ( .A(a[10]), .B(b[15]), .Z(n1537) );
  XOR U1609 ( .A(n1538), .B(n1537), .Z(n1556) );
  XNOR U1610 ( .A(n9622), .B(n2245), .Z(n1547) );
  OR U1611 ( .A(n1547), .B(n9623), .Z(n1471) );
  NANDN U1612 ( .A(n1469), .B(n9680), .Z(n1470) );
  NAND U1613 ( .A(n1471), .B(n1470), .Z(n1532) );
  XNOR U1614 ( .A(n9872), .B(n2062), .Z(n1550) );
  NANDN U1615 ( .A(n1550), .B(n9746), .Z(n1474) );
  NANDN U1616 ( .A(n1472), .B(n9747), .Z(n1473) );
  NAND U1617 ( .A(n1474), .B(n1473), .Z(n1529) );
  IV U1618 ( .A(a[24]), .Z(n2374) );
  XNOR U1619 ( .A(n74), .B(n2374), .Z(n1553) );
  NANDN U1620 ( .A(n1553), .B(n9485), .Z(n1477) );
  NANDN U1621 ( .A(n1475), .B(n9484), .Z(n1476) );
  AND U1622 ( .A(n1477), .B(n1476), .Z(n1530) );
  XNOR U1623 ( .A(n1529), .B(n1530), .Z(n1531) );
  XOR U1624 ( .A(n1532), .B(n1531), .Z(n1557) );
  XOR U1625 ( .A(n1556), .B(n1557), .Z(n1558) );
  XNOR U1626 ( .A(n1559), .B(n1558), .Z(n1507) );
  NAND U1627 ( .A(n1479), .B(n1478), .Z(n1483) );
  NAND U1628 ( .A(n1481), .B(n1480), .Z(n1482) );
  NAND U1629 ( .A(n1483), .B(n1482), .Z(n1508) );
  XOR U1630 ( .A(n1507), .B(n1508), .Z(n1510) );
  XNOR U1631 ( .A(n1509), .B(n1510), .Z(n1568) );
  NANDN U1632 ( .A(n1485), .B(n1484), .Z(n1489) );
  NAND U1633 ( .A(n1487), .B(n1486), .Z(n1488) );
  NAND U1634 ( .A(n1489), .B(n1488), .Z(n1569) );
  XNOR U1635 ( .A(n1568), .B(n1569), .Z(n1570) );
  XOR U1636 ( .A(n1571), .B(n1570), .Z(n1501) );
  NANDN U1637 ( .A(n1491), .B(n1490), .Z(n1495) );
  NANDN U1638 ( .A(n1493), .B(n1492), .Z(n1494) );
  NAND U1639 ( .A(n1495), .B(n1494), .Z(n1502) );
  XNOR U1640 ( .A(n1501), .B(n1502), .Z(n1503) );
  XNOR U1641 ( .A(n1504), .B(n1503), .Z(n1574) );
  XNOR U1642 ( .A(n1574), .B(sreg[138]), .Z(n1576) );
  NAND U1643 ( .A(n1496), .B(sreg[137]), .Z(n1500) );
  OR U1644 ( .A(n1498), .B(n1497), .Z(n1499) );
  AND U1645 ( .A(n1500), .B(n1499), .Z(n1575) );
  XOR U1646 ( .A(n1576), .B(n1575), .Z(c[138]) );
  NANDN U1647 ( .A(n1502), .B(n1501), .Z(n1506) );
  NAND U1648 ( .A(n1504), .B(n1503), .Z(n1505) );
  NAND U1649 ( .A(n1506), .B(n1505), .Z(n1582) );
  NANDN U1650 ( .A(n1508), .B(n1507), .Z(n1512) );
  OR U1651 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U1652 ( .A(n1512), .B(n1511), .Z(n1649) );
  XNOR U1653 ( .A(n9967), .B(n1828), .Z(n1618) );
  OR U1654 ( .A(n1618), .B(n10020), .Z(n1515) );
  NANDN U1655 ( .A(n1513), .B(n9968), .Z(n1514) );
  NAND U1656 ( .A(n1515), .B(n1514), .Z(n1631) );
  XNOR U1657 ( .A(n75), .B(n1516), .Z(n1622) );
  OR U1658 ( .A(n1622), .B(n10106), .Z(n1519) );
  NANDN U1659 ( .A(n1517), .B(n10107), .Z(n1518) );
  NAND U1660 ( .A(n1519), .B(n1518), .Z(n1628) );
  XNOR U1661 ( .A(n9984), .B(n1984), .Z(n1625) );
  NANDN U1662 ( .A(n1625), .B(n9865), .Z(n1522) );
  NANDN U1663 ( .A(n1520), .B(n9930), .Z(n1521) );
  AND U1664 ( .A(n1522), .B(n1521), .Z(n1629) );
  XNOR U1665 ( .A(n1628), .B(n1629), .Z(n1630) );
  XNOR U1666 ( .A(n1631), .B(n1630), .Z(n1640) );
  NANDN U1667 ( .A(n1524), .B(n1523), .Z(n1528) );
  NAND U1668 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1669 ( .A(n1528), .B(n1527), .Z(n1641) );
  XNOR U1670 ( .A(n1640), .B(n1641), .Z(n1642) );
  NANDN U1671 ( .A(n1530), .B(n1529), .Z(n1534) );
  NAND U1672 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1673 ( .A(n1534), .B(n1533), .Z(n1643) );
  XNOR U1674 ( .A(n1642), .B(n1643), .Z(n1587) );
  NANDN U1675 ( .A(n1536), .B(n1535), .Z(n1540) );
  OR U1676 ( .A(n1538), .B(n1537), .Z(n1539) );
  NAND U1677 ( .A(n1540), .B(n1539), .Z(n1615) );
  NAND U1678 ( .A(b[0]), .B(a[27]), .Z(n1541) );
  XNOR U1679 ( .A(b[1]), .B(n1541), .Z(n1543) );
  NAND U1680 ( .A(a[26]), .B(n72), .Z(n1542) );
  AND U1681 ( .A(n1543), .B(n1542), .Z(n1591) );
  XNOR U1682 ( .A(n10050), .B(n1672), .Z(n1600) );
  OR U1683 ( .A(n1600), .B(n10051), .Z(n1546) );
  NANDN U1684 ( .A(n1544), .B(n10070), .Z(n1545) );
  AND U1685 ( .A(n1546), .B(n1545), .Z(n1592) );
  XOR U1686 ( .A(n1591), .B(n1592), .Z(n1594) );
  NAND U1687 ( .A(a[11]), .B(b[15]), .Z(n1593) );
  XOR U1688 ( .A(n1594), .B(n1593), .Z(n1612) );
  XNOR U1689 ( .A(n9622), .B(n2323), .Z(n1603) );
  OR U1690 ( .A(n1603), .B(n9623), .Z(n1549) );
  NANDN U1691 ( .A(n1547), .B(n9680), .Z(n1548) );
  NAND U1692 ( .A(n1549), .B(n1548), .Z(n1637) );
  XNOR U1693 ( .A(n9872), .B(n2167), .Z(n1606) );
  NANDN U1694 ( .A(n1606), .B(n9746), .Z(n1552) );
  NANDN U1695 ( .A(n1550), .B(n9747), .Z(n1551) );
  NAND U1696 ( .A(n1552), .B(n1551), .Z(n1634) );
  IV U1697 ( .A(a[25]), .Z(n2450) );
  XNOR U1698 ( .A(n74), .B(n2450), .Z(n1609) );
  NANDN U1699 ( .A(n1609), .B(n9485), .Z(n1555) );
  NANDN U1700 ( .A(n1553), .B(n9484), .Z(n1554) );
  AND U1701 ( .A(n1555), .B(n1554), .Z(n1635) );
  XNOR U1702 ( .A(n1634), .B(n1635), .Z(n1636) );
  XOR U1703 ( .A(n1637), .B(n1636), .Z(n1613) );
  XOR U1704 ( .A(n1612), .B(n1613), .Z(n1614) );
  XNOR U1705 ( .A(n1615), .B(n1614), .Z(n1585) );
  NAND U1706 ( .A(n1557), .B(n1556), .Z(n1561) );
  NAND U1707 ( .A(n1559), .B(n1558), .Z(n1560) );
  NAND U1708 ( .A(n1561), .B(n1560), .Z(n1586) );
  XOR U1709 ( .A(n1585), .B(n1586), .Z(n1588) );
  XNOR U1710 ( .A(n1587), .B(n1588), .Z(n1646) );
  NANDN U1711 ( .A(n1563), .B(n1562), .Z(n1567) );
  NAND U1712 ( .A(n1565), .B(n1564), .Z(n1566) );
  NAND U1713 ( .A(n1567), .B(n1566), .Z(n1647) );
  XNOR U1714 ( .A(n1646), .B(n1647), .Z(n1648) );
  XOR U1715 ( .A(n1649), .B(n1648), .Z(n1579) );
  NANDN U1716 ( .A(n1569), .B(n1568), .Z(n1573) );
  NANDN U1717 ( .A(n1571), .B(n1570), .Z(n1572) );
  NAND U1718 ( .A(n1573), .B(n1572), .Z(n1580) );
  XNOR U1719 ( .A(n1579), .B(n1580), .Z(n1581) );
  XNOR U1720 ( .A(n1582), .B(n1581), .Z(n1652) );
  XNOR U1721 ( .A(n1652), .B(sreg[139]), .Z(n1654) );
  NAND U1722 ( .A(n1574), .B(sreg[138]), .Z(n1578) );
  OR U1723 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U1724 ( .A(n1578), .B(n1577), .Z(n1653) );
  XOR U1725 ( .A(n1654), .B(n1653), .Z(c[139]) );
  NANDN U1726 ( .A(n1580), .B(n1579), .Z(n1584) );
  NAND U1727 ( .A(n1582), .B(n1581), .Z(n1583) );
  NAND U1728 ( .A(n1584), .B(n1583), .Z(n1660) );
  NANDN U1729 ( .A(n1586), .B(n1585), .Z(n1590) );
  OR U1730 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U1731 ( .A(n1590), .B(n1589), .Z(n1727) );
  NANDN U1732 ( .A(n1592), .B(n1591), .Z(n1596) );
  OR U1733 ( .A(n1594), .B(n1593), .Z(n1595) );
  NAND U1734 ( .A(n1596), .B(n1595), .Z(n1715) );
  NAND U1735 ( .A(b[0]), .B(a[28]), .Z(n1597) );
  XNOR U1736 ( .A(b[1]), .B(n1597), .Z(n1599) );
  NAND U1737 ( .A(a[27]), .B(n72), .Z(n1598) );
  AND U1738 ( .A(n1599), .B(n1598), .Z(n1691) );
  XNOR U1739 ( .A(n10050), .B(n1750), .Z(n1700) );
  OR U1740 ( .A(n1700), .B(n10051), .Z(n1602) );
  NANDN U1741 ( .A(n1600), .B(n10070), .Z(n1601) );
  AND U1742 ( .A(n1602), .B(n1601), .Z(n1692) );
  XOR U1743 ( .A(n1691), .B(n1692), .Z(n1694) );
  NAND U1744 ( .A(a[12]), .B(b[15]), .Z(n1693) );
  XOR U1745 ( .A(n1694), .B(n1693), .Z(n1712) );
  XNOR U1746 ( .A(n9622), .B(n2374), .Z(n1703) );
  OR U1747 ( .A(n1703), .B(n9623), .Z(n1605) );
  NANDN U1748 ( .A(n1603), .B(n9680), .Z(n1604) );
  NAND U1749 ( .A(n1605), .B(n1604), .Z(n1688) );
  XNOR U1750 ( .A(n9872), .B(n2245), .Z(n1706) );
  NANDN U1751 ( .A(n1706), .B(n9746), .Z(n1608) );
  NANDN U1752 ( .A(n1606), .B(n9747), .Z(n1607) );
  NAND U1753 ( .A(n1608), .B(n1607), .Z(n1685) );
  IV U1754 ( .A(a[26]), .Z(n2555) );
  XNOR U1755 ( .A(n74), .B(n2555), .Z(n1709) );
  NANDN U1756 ( .A(n1709), .B(n9485), .Z(n1611) );
  NANDN U1757 ( .A(n1609), .B(n9484), .Z(n1610) );
  AND U1758 ( .A(n1611), .B(n1610), .Z(n1686) );
  XNOR U1759 ( .A(n1685), .B(n1686), .Z(n1687) );
  XOR U1760 ( .A(n1688), .B(n1687), .Z(n1713) );
  XOR U1761 ( .A(n1712), .B(n1713), .Z(n1714) );
  XNOR U1762 ( .A(n1715), .B(n1714), .Z(n1663) );
  NAND U1763 ( .A(n1613), .B(n1612), .Z(n1617) );
  NAND U1764 ( .A(n1615), .B(n1614), .Z(n1616) );
  NAND U1765 ( .A(n1617), .B(n1616), .Z(n1664) );
  XOR U1766 ( .A(n1663), .B(n1664), .Z(n1666) );
  XNOR U1767 ( .A(n9967), .B(n1906), .Z(n1669) );
  OR U1768 ( .A(n1669), .B(n10020), .Z(n1620) );
  NANDN U1769 ( .A(n1618), .B(n9968), .Z(n1619) );
  NAND U1770 ( .A(n1620), .B(n1619), .Z(n1682) );
  XNOR U1771 ( .A(n75), .B(n1621), .Z(n1673) );
  OR U1772 ( .A(n1673), .B(n10106), .Z(n1624) );
  NANDN U1773 ( .A(n1622), .B(n10107), .Z(n1623) );
  NAND U1774 ( .A(n1624), .B(n1623), .Z(n1679) );
  XNOR U1775 ( .A(n9984), .B(n2062), .Z(n1676) );
  NANDN U1776 ( .A(n1676), .B(n9865), .Z(n1627) );
  NANDN U1777 ( .A(n1625), .B(n9930), .Z(n1626) );
  AND U1778 ( .A(n1627), .B(n1626), .Z(n1680) );
  XNOR U1779 ( .A(n1679), .B(n1680), .Z(n1681) );
  XNOR U1780 ( .A(n1682), .B(n1681), .Z(n1718) );
  NANDN U1781 ( .A(n1629), .B(n1628), .Z(n1633) );
  NAND U1782 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U1783 ( .A(n1633), .B(n1632), .Z(n1719) );
  XNOR U1784 ( .A(n1718), .B(n1719), .Z(n1720) );
  NANDN U1785 ( .A(n1635), .B(n1634), .Z(n1639) );
  NAND U1786 ( .A(n1637), .B(n1636), .Z(n1638) );
  AND U1787 ( .A(n1639), .B(n1638), .Z(n1721) );
  XNOR U1788 ( .A(n1720), .B(n1721), .Z(n1665) );
  XNOR U1789 ( .A(n1666), .B(n1665), .Z(n1724) );
  NANDN U1790 ( .A(n1641), .B(n1640), .Z(n1645) );
  NAND U1791 ( .A(n1643), .B(n1642), .Z(n1644) );
  NAND U1792 ( .A(n1645), .B(n1644), .Z(n1725) );
  XNOR U1793 ( .A(n1724), .B(n1725), .Z(n1726) );
  XOR U1794 ( .A(n1727), .B(n1726), .Z(n1657) );
  NANDN U1795 ( .A(n1647), .B(n1646), .Z(n1651) );
  NANDN U1796 ( .A(n1649), .B(n1648), .Z(n1650) );
  NAND U1797 ( .A(n1651), .B(n1650), .Z(n1658) );
  XNOR U1798 ( .A(n1657), .B(n1658), .Z(n1659) );
  XNOR U1799 ( .A(n1660), .B(n1659), .Z(n1730) );
  XNOR U1800 ( .A(n1730), .B(sreg[140]), .Z(n1732) );
  NAND U1801 ( .A(n1652), .B(sreg[139]), .Z(n1656) );
  OR U1802 ( .A(n1654), .B(n1653), .Z(n1655) );
  AND U1803 ( .A(n1656), .B(n1655), .Z(n1731) );
  XOR U1804 ( .A(n1732), .B(n1731), .Z(c[140]) );
  NANDN U1805 ( .A(n1658), .B(n1657), .Z(n1662) );
  NAND U1806 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U1807 ( .A(n1662), .B(n1661), .Z(n1738) );
  NANDN U1808 ( .A(n1664), .B(n1663), .Z(n1668) );
  OR U1809 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U1810 ( .A(n1668), .B(n1667), .Z(n1805) );
  XNOR U1811 ( .A(n9967), .B(n1984), .Z(n1747) );
  OR U1812 ( .A(n1747), .B(n10020), .Z(n1671) );
  NANDN U1813 ( .A(n1669), .B(n9968), .Z(n1670) );
  NAND U1814 ( .A(n1671), .B(n1670), .Z(n1760) );
  XNOR U1815 ( .A(n75), .B(n1672), .Z(n1751) );
  OR U1816 ( .A(n1751), .B(n10106), .Z(n1675) );
  NANDN U1817 ( .A(n1673), .B(n10107), .Z(n1674) );
  NAND U1818 ( .A(n1675), .B(n1674), .Z(n1757) );
  XNOR U1819 ( .A(n9984), .B(n2167), .Z(n1754) );
  NANDN U1820 ( .A(n1754), .B(n9865), .Z(n1678) );
  NANDN U1821 ( .A(n1676), .B(n9930), .Z(n1677) );
  AND U1822 ( .A(n1678), .B(n1677), .Z(n1758) );
  XNOR U1823 ( .A(n1757), .B(n1758), .Z(n1759) );
  XNOR U1824 ( .A(n1760), .B(n1759), .Z(n1796) );
  NANDN U1825 ( .A(n1680), .B(n1679), .Z(n1684) );
  NAND U1826 ( .A(n1682), .B(n1681), .Z(n1683) );
  NAND U1827 ( .A(n1684), .B(n1683), .Z(n1797) );
  XNOR U1828 ( .A(n1796), .B(n1797), .Z(n1798) );
  NANDN U1829 ( .A(n1686), .B(n1685), .Z(n1690) );
  NAND U1830 ( .A(n1688), .B(n1687), .Z(n1689) );
  AND U1831 ( .A(n1690), .B(n1689), .Z(n1799) );
  XNOR U1832 ( .A(n1798), .B(n1799), .Z(n1743) );
  NANDN U1833 ( .A(n1692), .B(n1691), .Z(n1696) );
  OR U1834 ( .A(n1694), .B(n1693), .Z(n1695) );
  NAND U1835 ( .A(n1696), .B(n1695), .Z(n1793) );
  NAND U1836 ( .A(b[0]), .B(a[29]), .Z(n1697) );
  XNOR U1837 ( .A(b[1]), .B(n1697), .Z(n1699) );
  NAND U1838 ( .A(a[28]), .B(n72), .Z(n1698) );
  AND U1839 ( .A(n1699), .B(n1698), .Z(n1769) );
  XNOR U1840 ( .A(n10050), .B(n1828), .Z(n1778) );
  OR U1841 ( .A(n1778), .B(n10051), .Z(n1702) );
  NANDN U1842 ( .A(n1700), .B(n10070), .Z(n1701) );
  AND U1843 ( .A(n1702), .B(n1701), .Z(n1770) );
  XOR U1844 ( .A(n1769), .B(n1770), .Z(n1772) );
  NAND U1845 ( .A(a[13]), .B(b[15]), .Z(n1771) );
  XOR U1846 ( .A(n1772), .B(n1771), .Z(n1790) );
  XNOR U1847 ( .A(n9622), .B(n2450), .Z(n1781) );
  OR U1848 ( .A(n1781), .B(n9623), .Z(n1705) );
  NANDN U1849 ( .A(n1703), .B(n9680), .Z(n1704) );
  NAND U1850 ( .A(n1705), .B(n1704), .Z(n1766) );
  XNOR U1851 ( .A(n9872), .B(n2323), .Z(n1784) );
  NANDN U1852 ( .A(n1784), .B(n9746), .Z(n1708) );
  NANDN U1853 ( .A(n1706), .B(n9747), .Z(n1707) );
  NAND U1854 ( .A(n1708), .B(n1707), .Z(n1763) );
  IV U1855 ( .A(a[27]), .Z(n2606) );
  XNOR U1856 ( .A(n74), .B(n2606), .Z(n1787) );
  NANDN U1857 ( .A(n1787), .B(n9485), .Z(n1711) );
  NANDN U1858 ( .A(n1709), .B(n9484), .Z(n1710) );
  AND U1859 ( .A(n1711), .B(n1710), .Z(n1764) );
  XNOR U1860 ( .A(n1763), .B(n1764), .Z(n1765) );
  XOR U1861 ( .A(n1766), .B(n1765), .Z(n1791) );
  XOR U1862 ( .A(n1790), .B(n1791), .Z(n1792) );
  XNOR U1863 ( .A(n1793), .B(n1792), .Z(n1741) );
  NAND U1864 ( .A(n1713), .B(n1712), .Z(n1717) );
  NAND U1865 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U1866 ( .A(n1717), .B(n1716), .Z(n1742) );
  XOR U1867 ( .A(n1741), .B(n1742), .Z(n1744) );
  XNOR U1868 ( .A(n1743), .B(n1744), .Z(n1802) );
  NANDN U1869 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U1870 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U1871 ( .A(n1723), .B(n1722), .Z(n1803) );
  XNOR U1872 ( .A(n1802), .B(n1803), .Z(n1804) );
  XOR U1873 ( .A(n1805), .B(n1804), .Z(n1735) );
  NANDN U1874 ( .A(n1725), .B(n1724), .Z(n1729) );
  NANDN U1875 ( .A(n1727), .B(n1726), .Z(n1728) );
  NAND U1876 ( .A(n1729), .B(n1728), .Z(n1736) );
  XNOR U1877 ( .A(n1735), .B(n1736), .Z(n1737) );
  XNOR U1878 ( .A(n1738), .B(n1737), .Z(n1808) );
  XNOR U1879 ( .A(n1808), .B(sreg[141]), .Z(n1810) );
  NAND U1880 ( .A(n1730), .B(sreg[140]), .Z(n1734) );
  OR U1881 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U1882 ( .A(n1734), .B(n1733), .Z(n1809) );
  XOR U1883 ( .A(n1810), .B(n1809), .Z(c[141]) );
  NANDN U1884 ( .A(n1736), .B(n1735), .Z(n1740) );
  NAND U1885 ( .A(n1738), .B(n1737), .Z(n1739) );
  NAND U1886 ( .A(n1740), .B(n1739), .Z(n1816) );
  NANDN U1887 ( .A(n1742), .B(n1741), .Z(n1746) );
  OR U1888 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U1889 ( .A(n1746), .B(n1745), .Z(n1883) );
  XNOR U1890 ( .A(n9967), .B(n2062), .Z(n1825) );
  OR U1891 ( .A(n1825), .B(n10020), .Z(n1749) );
  NANDN U1892 ( .A(n1747), .B(n9968), .Z(n1748) );
  NAND U1893 ( .A(n1749), .B(n1748), .Z(n1838) );
  XNOR U1894 ( .A(n75), .B(n1750), .Z(n1829) );
  OR U1895 ( .A(n1829), .B(n10106), .Z(n1753) );
  NANDN U1896 ( .A(n1751), .B(n10107), .Z(n1752) );
  NAND U1897 ( .A(n1753), .B(n1752), .Z(n1835) );
  XNOR U1898 ( .A(n9984), .B(n2245), .Z(n1832) );
  NANDN U1899 ( .A(n1832), .B(n9865), .Z(n1756) );
  NANDN U1900 ( .A(n1754), .B(n9930), .Z(n1755) );
  AND U1901 ( .A(n1756), .B(n1755), .Z(n1836) );
  XNOR U1902 ( .A(n1835), .B(n1836), .Z(n1837) );
  XNOR U1903 ( .A(n1838), .B(n1837), .Z(n1874) );
  NANDN U1904 ( .A(n1758), .B(n1757), .Z(n1762) );
  NAND U1905 ( .A(n1760), .B(n1759), .Z(n1761) );
  NAND U1906 ( .A(n1762), .B(n1761), .Z(n1875) );
  XNOR U1907 ( .A(n1874), .B(n1875), .Z(n1876) );
  NANDN U1908 ( .A(n1764), .B(n1763), .Z(n1768) );
  NAND U1909 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U1910 ( .A(n1768), .B(n1767), .Z(n1877) );
  XNOR U1911 ( .A(n1876), .B(n1877), .Z(n1821) );
  NANDN U1912 ( .A(n1770), .B(n1769), .Z(n1774) );
  OR U1913 ( .A(n1772), .B(n1771), .Z(n1773) );
  NAND U1914 ( .A(n1774), .B(n1773), .Z(n1871) );
  NAND U1915 ( .A(b[0]), .B(a[30]), .Z(n1775) );
  XNOR U1916 ( .A(b[1]), .B(n1775), .Z(n1777) );
  NAND U1917 ( .A(a[29]), .B(n72), .Z(n1776) );
  AND U1918 ( .A(n1777), .B(n1776), .Z(n1847) );
  XNOR U1919 ( .A(n10050), .B(n1906), .Z(n1856) );
  OR U1920 ( .A(n1856), .B(n10051), .Z(n1780) );
  NANDN U1921 ( .A(n1778), .B(n10070), .Z(n1779) );
  AND U1922 ( .A(n1780), .B(n1779), .Z(n1848) );
  XOR U1923 ( .A(n1847), .B(n1848), .Z(n1850) );
  NAND U1924 ( .A(a[14]), .B(b[15]), .Z(n1849) );
  XOR U1925 ( .A(n1850), .B(n1849), .Z(n1868) );
  XNOR U1926 ( .A(n9622), .B(n2555), .Z(n1859) );
  OR U1927 ( .A(n1859), .B(n9623), .Z(n1783) );
  NANDN U1928 ( .A(n1781), .B(n9680), .Z(n1782) );
  NAND U1929 ( .A(n1783), .B(n1782), .Z(n1844) );
  XNOR U1930 ( .A(n9872), .B(n2374), .Z(n1862) );
  NANDN U1931 ( .A(n1862), .B(n9746), .Z(n1786) );
  NANDN U1932 ( .A(n1784), .B(n9747), .Z(n1785) );
  NAND U1933 ( .A(n1786), .B(n1785), .Z(n1841) );
  IV U1934 ( .A(a[28]), .Z(n2711) );
  XNOR U1935 ( .A(n74), .B(n2711), .Z(n1865) );
  NANDN U1936 ( .A(n1865), .B(n9485), .Z(n1789) );
  NANDN U1937 ( .A(n1787), .B(n9484), .Z(n1788) );
  AND U1938 ( .A(n1789), .B(n1788), .Z(n1842) );
  XNOR U1939 ( .A(n1841), .B(n1842), .Z(n1843) );
  XOR U1940 ( .A(n1844), .B(n1843), .Z(n1869) );
  XOR U1941 ( .A(n1868), .B(n1869), .Z(n1870) );
  XNOR U1942 ( .A(n1871), .B(n1870), .Z(n1819) );
  NAND U1943 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U1944 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U1945 ( .A(n1795), .B(n1794), .Z(n1820) );
  XOR U1946 ( .A(n1819), .B(n1820), .Z(n1822) );
  XNOR U1947 ( .A(n1821), .B(n1822), .Z(n1880) );
  NANDN U1948 ( .A(n1797), .B(n1796), .Z(n1801) );
  NAND U1949 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U1950 ( .A(n1801), .B(n1800), .Z(n1881) );
  XNOR U1951 ( .A(n1880), .B(n1881), .Z(n1882) );
  XOR U1952 ( .A(n1883), .B(n1882), .Z(n1813) );
  NANDN U1953 ( .A(n1803), .B(n1802), .Z(n1807) );
  NANDN U1954 ( .A(n1805), .B(n1804), .Z(n1806) );
  NAND U1955 ( .A(n1807), .B(n1806), .Z(n1814) );
  XNOR U1956 ( .A(n1813), .B(n1814), .Z(n1815) );
  XNOR U1957 ( .A(n1816), .B(n1815), .Z(n1886) );
  XNOR U1958 ( .A(n1886), .B(sreg[142]), .Z(n1888) );
  NAND U1959 ( .A(n1808), .B(sreg[141]), .Z(n1812) );
  OR U1960 ( .A(n1810), .B(n1809), .Z(n1811) );
  AND U1961 ( .A(n1812), .B(n1811), .Z(n1887) );
  XOR U1962 ( .A(n1888), .B(n1887), .Z(c[142]) );
  NANDN U1963 ( .A(n1814), .B(n1813), .Z(n1818) );
  NAND U1964 ( .A(n1816), .B(n1815), .Z(n1817) );
  NAND U1965 ( .A(n1818), .B(n1817), .Z(n1894) );
  NANDN U1966 ( .A(n1820), .B(n1819), .Z(n1824) );
  OR U1967 ( .A(n1822), .B(n1821), .Z(n1823) );
  NAND U1968 ( .A(n1824), .B(n1823), .Z(n1961) );
  XNOR U1969 ( .A(n9967), .B(n2167), .Z(n1903) );
  OR U1970 ( .A(n1903), .B(n10020), .Z(n1827) );
  NANDN U1971 ( .A(n1825), .B(n9968), .Z(n1826) );
  NAND U1972 ( .A(n1827), .B(n1826), .Z(n1916) );
  XNOR U1973 ( .A(n75), .B(n1828), .Z(n1907) );
  OR U1974 ( .A(n1907), .B(n10106), .Z(n1831) );
  NANDN U1975 ( .A(n1829), .B(n10107), .Z(n1830) );
  NAND U1976 ( .A(n1831), .B(n1830), .Z(n1913) );
  XNOR U1977 ( .A(n9984), .B(n2323), .Z(n1910) );
  NANDN U1978 ( .A(n1910), .B(n9865), .Z(n1834) );
  NANDN U1979 ( .A(n1832), .B(n9930), .Z(n1833) );
  AND U1980 ( .A(n1834), .B(n1833), .Z(n1914) );
  XNOR U1981 ( .A(n1913), .B(n1914), .Z(n1915) );
  XNOR U1982 ( .A(n1916), .B(n1915), .Z(n1952) );
  NANDN U1983 ( .A(n1836), .B(n1835), .Z(n1840) );
  NAND U1984 ( .A(n1838), .B(n1837), .Z(n1839) );
  NAND U1985 ( .A(n1840), .B(n1839), .Z(n1953) );
  XNOR U1986 ( .A(n1952), .B(n1953), .Z(n1954) );
  NANDN U1987 ( .A(n1842), .B(n1841), .Z(n1846) );
  NAND U1988 ( .A(n1844), .B(n1843), .Z(n1845) );
  AND U1989 ( .A(n1846), .B(n1845), .Z(n1955) );
  XNOR U1990 ( .A(n1954), .B(n1955), .Z(n1899) );
  NANDN U1991 ( .A(n1848), .B(n1847), .Z(n1852) );
  OR U1992 ( .A(n1850), .B(n1849), .Z(n1851) );
  NAND U1993 ( .A(n1852), .B(n1851), .Z(n1949) );
  NAND U1994 ( .A(b[0]), .B(a[31]), .Z(n1853) );
  XNOR U1995 ( .A(b[1]), .B(n1853), .Z(n1855) );
  NAND U1996 ( .A(a[30]), .B(n72), .Z(n1854) );
  AND U1997 ( .A(n1855), .B(n1854), .Z(n1925) );
  XNOR U1998 ( .A(n10050), .B(n1984), .Z(n1934) );
  OR U1999 ( .A(n1934), .B(n10051), .Z(n1858) );
  NANDN U2000 ( .A(n1856), .B(n10070), .Z(n1857) );
  AND U2001 ( .A(n1858), .B(n1857), .Z(n1926) );
  XOR U2002 ( .A(n1925), .B(n1926), .Z(n1928) );
  NAND U2003 ( .A(a[15]), .B(b[15]), .Z(n1927) );
  XOR U2004 ( .A(n1928), .B(n1927), .Z(n1946) );
  XNOR U2005 ( .A(n9622), .B(n2606), .Z(n1937) );
  OR U2006 ( .A(n1937), .B(n9623), .Z(n1861) );
  NANDN U2007 ( .A(n1859), .B(n9680), .Z(n1860) );
  NAND U2008 ( .A(n1861), .B(n1860), .Z(n1922) );
  XNOR U2009 ( .A(n9872), .B(n2450), .Z(n1940) );
  NANDN U2010 ( .A(n1940), .B(n9746), .Z(n1864) );
  NANDN U2011 ( .A(n1862), .B(n9747), .Z(n1863) );
  NAND U2012 ( .A(n1864), .B(n1863), .Z(n1919) );
  IV U2013 ( .A(a[29]), .Z(n2762) );
  XNOR U2014 ( .A(n74), .B(n2762), .Z(n1943) );
  NANDN U2015 ( .A(n1943), .B(n9485), .Z(n1867) );
  NANDN U2016 ( .A(n1865), .B(n9484), .Z(n1866) );
  AND U2017 ( .A(n1867), .B(n1866), .Z(n1920) );
  XNOR U2018 ( .A(n1919), .B(n1920), .Z(n1921) );
  XOR U2019 ( .A(n1922), .B(n1921), .Z(n1947) );
  XOR U2020 ( .A(n1946), .B(n1947), .Z(n1948) );
  XNOR U2021 ( .A(n1949), .B(n1948), .Z(n1897) );
  NAND U2022 ( .A(n1869), .B(n1868), .Z(n1873) );
  NAND U2023 ( .A(n1871), .B(n1870), .Z(n1872) );
  NAND U2024 ( .A(n1873), .B(n1872), .Z(n1898) );
  XOR U2025 ( .A(n1897), .B(n1898), .Z(n1900) );
  XNOR U2026 ( .A(n1899), .B(n1900), .Z(n1958) );
  NANDN U2027 ( .A(n1875), .B(n1874), .Z(n1879) );
  NAND U2028 ( .A(n1877), .B(n1876), .Z(n1878) );
  NAND U2029 ( .A(n1879), .B(n1878), .Z(n1959) );
  XNOR U2030 ( .A(n1958), .B(n1959), .Z(n1960) );
  XOR U2031 ( .A(n1961), .B(n1960), .Z(n1891) );
  NANDN U2032 ( .A(n1881), .B(n1880), .Z(n1885) );
  NANDN U2033 ( .A(n1883), .B(n1882), .Z(n1884) );
  NAND U2034 ( .A(n1885), .B(n1884), .Z(n1892) );
  XNOR U2035 ( .A(n1891), .B(n1892), .Z(n1893) );
  XNOR U2036 ( .A(n1894), .B(n1893), .Z(n1964) );
  XNOR U2037 ( .A(n1964), .B(sreg[143]), .Z(n1966) );
  NAND U2038 ( .A(n1886), .B(sreg[142]), .Z(n1890) );
  OR U2039 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U2040 ( .A(n1890), .B(n1889), .Z(n1965) );
  XOR U2041 ( .A(n1966), .B(n1965), .Z(c[143]) );
  NANDN U2042 ( .A(n1892), .B(n1891), .Z(n1896) );
  NAND U2043 ( .A(n1894), .B(n1893), .Z(n1895) );
  NAND U2044 ( .A(n1896), .B(n1895), .Z(n1972) );
  NANDN U2045 ( .A(n1898), .B(n1897), .Z(n1902) );
  OR U2046 ( .A(n1900), .B(n1899), .Z(n1901) );
  NAND U2047 ( .A(n1902), .B(n1901), .Z(n2039) );
  XNOR U2048 ( .A(n9967), .B(n2245), .Z(n1981) );
  OR U2049 ( .A(n1981), .B(n10020), .Z(n1905) );
  NANDN U2050 ( .A(n1903), .B(n9968), .Z(n1904) );
  NAND U2051 ( .A(n1905), .B(n1904), .Z(n1994) );
  XNOR U2052 ( .A(n75), .B(n1906), .Z(n1985) );
  OR U2053 ( .A(n1985), .B(n10106), .Z(n1909) );
  NANDN U2054 ( .A(n1907), .B(n10107), .Z(n1908) );
  NAND U2055 ( .A(n1909), .B(n1908), .Z(n1991) );
  XNOR U2056 ( .A(n9984), .B(n2374), .Z(n1988) );
  NANDN U2057 ( .A(n1988), .B(n9865), .Z(n1912) );
  NANDN U2058 ( .A(n1910), .B(n9930), .Z(n1911) );
  AND U2059 ( .A(n1912), .B(n1911), .Z(n1992) );
  XNOR U2060 ( .A(n1991), .B(n1992), .Z(n1993) );
  XNOR U2061 ( .A(n1994), .B(n1993), .Z(n2030) );
  NANDN U2062 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2063 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2064 ( .A(n1918), .B(n1917), .Z(n2031) );
  XNOR U2065 ( .A(n2030), .B(n2031), .Z(n2032) );
  NANDN U2066 ( .A(n1920), .B(n1919), .Z(n1924) );
  NAND U2067 ( .A(n1922), .B(n1921), .Z(n1923) );
  AND U2068 ( .A(n1924), .B(n1923), .Z(n2033) );
  XNOR U2069 ( .A(n2032), .B(n2033), .Z(n1977) );
  NANDN U2070 ( .A(n1926), .B(n1925), .Z(n1930) );
  OR U2071 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2072 ( .A(n1930), .B(n1929), .Z(n2027) );
  NAND U2073 ( .A(b[0]), .B(a[32]), .Z(n1931) );
  XNOR U2074 ( .A(b[1]), .B(n1931), .Z(n1933) );
  NAND U2075 ( .A(a[31]), .B(n72), .Z(n1932) );
  AND U2076 ( .A(n1933), .B(n1932), .Z(n2003) );
  XNOR U2077 ( .A(n10050), .B(n2062), .Z(n2012) );
  OR U2078 ( .A(n2012), .B(n10051), .Z(n1936) );
  NANDN U2079 ( .A(n1934), .B(n10070), .Z(n1935) );
  AND U2080 ( .A(n1936), .B(n1935), .Z(n2004) );
  XOR U2081 ( .A(n2003), .B(n2004), .Z(n2006) );
  NAND U2082 ( .A(a[16]), .B(b[15]), .Z(n2005) );
  XOR U2083 ( .A(n2006), .B(n2005), .Z(n2024) );
  XNOR U2084 ( .A(n9622), .B(n2711), .Z(n2015) );
  OR U2085 ( .A(n2015), .B(n9623), .Z(n1939) );
  NANDN U2086 ( .A(n1937), .B(n9680), .Z(n1938) );
  NAND U2087 ( .A(n1939), .B(n1938), .Z(n2000) );
  XNOR U2088 ( .A(n9872), .B(n2555), .Z(n2018) );
  NANDN U2089 ( .A(n2018), .B(n9746), .Z(n1942) );
  NANDN U2090 ( .A(n1940), .B(n9747), .Z(n1941) );
  NAND U2091 ( .A(n1942), .B(n1941), .Z(n1997) );
  IV U2092 ( .A(a[30]), .Z(n2840) );
  XNOR U2093 ( .A(n74), .B(n2840), .Z(n2021) );
  NANDN U2094 ( .A(n2021), .B(n9485), .Z(n1945) );
  NANDN U2095 ( .A(n1943), .B(n9484), .Z(n1944) );
  AND U2096 ( .A(n1945), .B(n1944), .Z(n1998) );
  XNOR U2097 ( .A(n1997), .B(n1998), .Z(n1999) );
  XOR U2098 ( .A(n2000), .B(n1999), .Z(n2025) );
  XOR U2099 ( .A(n2024), .B(n2025), .Z(n2026) );
  XNOR U2100 ( .A(n2027), .B(n2026), .Z(n1975) );
  NAND U2101 ( .A(n1947), .B(n1946), .Z(n1951) );
  NAND U2102 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U2103 ( .A(n1951), .B(n1950), .Z(n1976) );
  XOR U2104 ( .A(n1975), .B(n1976), .Z(n1978) );
  XNOR U2105 ( .A(n1977), .B(n1978), .Z(n2036) );
  NANDN U2106 ( .A(n1953), .B(n1952), .Z(n1957) );
  NAND U2107 ( .A(n1955), .B(n1954), .Z(n1956) );
  NAND U2108 ( .A(n1957), .B(n1956), .Z(n2037) );
  XNOR U2109 ( .A(n2036), .B(n2037), .Z(n2038) );
  XOR U2110 ( .A(n2039), .B(n2038), .Z(n1969) );
  NANDN U2111 ( .A(n1959), .B(n1958), .Z(n1963) );
  NANDN U2112 ( .A(n1961), .B(n1960), .Z(n1962) );
  NAND U2113 ( .A(n1963), .B(n1962), .Z(n1970) );
  XNOR U2114 ( .A(n1969), .B(n1970), .Z(n1971) );
  XNOR U2115 ( .A(n1972), .B(n1971), .Z(n2042) );
  XNOR U2116 ( .A(n2042), .B(sreg[144]), .Z(n2044) );
  NAND U2117 ( .A(n1964), .B(sreg[143]), .Z(n1968) );
  OR U2118 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2119 ( .A(n1968), .B(n1967), .Z(n2043) );
  XOR U2120 ( .A(n2044), .B(n2043), .Z(c[144]) );
  NANDN U2121 ( .A(n1970), .B(n1969), .Z(n1974) );
  NAND U2122 ( .A(n1972), .B(n1971), .Z(n1973) );
  NAND U2123 ( .A(n1974), .B(n1973), .Z(n2050) );
  NANDN U2124 ( .A(n1976), .B(n1975), .Z(n1980) );
  OR U2125 ( .A(n1978), .B(n1977), .Z(n1979) );
  NAND U2126 ( .A(n1980), .B(n1979), .Z(n2117) );
  XNOR U2127 ( .A(n9967), .B(n2323), .Z(n2059) );
  OR U2128 ( .A(n2059), .B(n10020), .Z(n1983) );
  NANDN U2129 ( .A(n1981), .B(n9968), .Z(n1982) );
  NAND U2130 ( .A(n1983), .B(n1982), .Z(n2072) );
  XNOR U2131 ( .A(n75), .B(n1984), .Z(n2063) );
  OR U2132 ( .A(n2063), .B(n10106), .Z(n1987) );
  NANDN U2133 ( .A(n1985), .B(n10107), .Z(n1986) );
  NAND U2134 ( .A(n1987), .B(n1986), .Z(n2069) );
  XNOR U2135 ( .A(n9984), .B(n2450), .Z(n2066) );
  NANDN U2136 ( .A(n2066), .B(n9865), .Z(n1990) );
  NANDN U2137 ( .A(n1988), .B(n9930), .Z(n1989) );
  AND U2138 ( .A(n1990), .B(n1989), .Z(n2070) );
  XNOR U2139 ( .A(n2069), .B(n2070), .Z(n2071) );
  XNOR U2140 ( .A(n2072), .B(n2071), .Z(n2108) );
  NANDN U2141 ( .A(n1992), .B(n1991), .Z(n1996) );
  NAND U2142 ( .A(n1994), .B(n1993), .Z(n1995) );
  NAND U2143 ( .A(n1996), .B(n1995), .Z(n2109) );
  XNOR U2144 ( .A(n2108), .B(n2109), .Z(n2110) );
  NANDN U2145 ( .A(n1998), .B(n1997), .Z(n2002) );
  NAND U2146 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2147 ( .A(n2002), .B(n2001), .Z(n2111) );
  XNOR U2148 ( .A(n2110), .B(n2111), .Z(n2055) );
  NANDN U2149 ( .A(n2004), .B(n2003), .Z(n2008) );
  OR U2150 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2151 ( .A(n2008), .B(n2007), .Z(n2105) );
  NAND U2152 ( .A(b[0]), .B(a[33]), .Z(n2009) );
  XNOR U2153 ( .A(b[1]), .B(n2009), .Z(n2011) );
  NAND U2154 ( .A(a[32]), .B(n72), .Z(n2010) );
  AND U2155 ( .A(n2011), .B(n2010), .Z(n2081) );
  XNOR U2156 ( .A(n10050), .B(n2167), .Z(n2087) );
  OR U2157 ( .A(n2087), .B(n10051), .Z(n2014) );
  NANDN U2158 ( .A(n2012), .B(n10070), .Z(n2013) );
  AND U2159 ( .A(n2014), .B(n2013), .Z(n2082) );
  XOR U2160 ( .A(n2081), .B(n2082), .Z(n2084) );
  NAND U2161 ( .A(a[17]), .B(b[15]), .Z(n2083) );
  XOR U2162 ( .A(n2084), .B(n2083), .Z(n2102) );
  XNOR U2163 ( .A(n9622), .B(n2762), .Z(n2093) );
  OR U2164 ( .A(n2093), .B(n9623), .Z(n2017) );
  NANDN U2165 ( .A(n2015), .B(n9680), .Z(n2016) );
  NAND U2166 ( .A(n2017), .B(n2016), .Z(n2078) );
  XNOR U2167 ( .A(n9872), .B(n2606), .Z(n2096) );
  NANDN U2168 ( .A(n2096), .B(n9746), .Z(n2020) );
  NANDN U2169 ( .A(n2018), .B(n9747), .Z(n2019) );
  NAND U2170 ( .A(n2020), .B(n2019), .Z(n2075) );
  IV U2171 ( .A(a[31]), .Z(n2918) );
  XNOR U2172 ( .A(n74), .B(n2918), .Z(n2099) );
  NANDN U2173 ( .A(n2099), .B(n9485), .Z(n2023) );
  NANDN U2174 ( .A(n2021), .B(n9484), .Z(n2022) );
  AND U2175 ( .A(n2023), .B(n2022), .Z(n2076) );
  XNOR U2176 ( .A(n2075), .B(n2076), .Z(n2077) );
  XOR U2177 ( .A(n2078), .B(n2077), .Z(n2103) );
  XOR U2178 ( .A(n2102), .B(n2103), .Z(n2104) );
  XNOR U2179 ( .A(n2105), .B(n2104), .Z(n2053) );
  NAND U2180 ( .A(n2025), .B(n2024), .Z(n2029) );
  NAND U2181 ( .A(n2027), .B(n2026), .Z(n2028) );
  NAND U2182 ( .A(n2029), .B(n2028), .Z(n2054) );
  XOR U2183 ( .A(n2053), .B(n2054), .Z(n2056) );
  XNOR U2184 ( .A(n2055), .B(n2056), .Z(n2114) );
  NANDN U2185 ( .A(n2031), .B(n2030), .Z(n2035) );
  NAND U2186 ( .A(n2033), .B(n2032), .Z(n2034) );
  NAND U2187 ( .A(n2035), .B(n2034), .Z(n2115) );
  XNOR U2188 ( .A(n2114), .B(n2115), .Z(n2116) );
  XOR U2189 ( .A(n2117), .B(n2116), .Z(n2047) );
  NANDN U2190 ( .A(n2037), .B(n2036), .Z(n2041) );
  NANDN U2191 ( .A(n2039), .B(n2038), .Z(n2040) );
  NAND U2192 ( .A(n2041), .B(n2040), .Z(n2048) );
  XNOR U2193 ( .A(n2047), .B(n2048), .Z(n2049) );
  XNOR U2194 ( .A(n2050), .B(n2049), .Z(n2120) );
  XNOR U2195 ( .A(n2120), .B(sreg[145]), .Z(n2122) );
  NAND U2196 ( .A(n2042), .B(sreg[144]), .Z(n2046) );
  OR U2197 ( .A(n2044), .B(n2043), .Z(n2045) );
  AND U2198 ( .A(n2046), .B(n2045), .Z(n2121) );
  XOR U2199 ( .A(n2122), .B(n2121), .Z(c[145]) );
  NANDN U2200 ( .A(n2048), .B(n2047), .Z(n2052) );
  NAND U2201 ( .A(n2050), .B(n2049), .Z(n2051) );
  NAND U2202 ( .A(n2052), .B(n2051), .Z(n2128) );
  NANDN U2203 ( .A(n2054), .B(n2053), .Z(n2058) );
  OR U2204 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U2205 ( .A(n2058), .B(n2057), .Z(n2195) );
  XNOR U2206 ( .A(n9967), .B(n2374), .Z(n2164) );
  OR U2207 ( .A(n2164), .B(n10020), .Z(n2061) );
  NANDN U2208 ( .A(n2059), .B(n9968), .Z(n2060) );
  NAND U2209 ( .A(n2061), .B(n2060), .Z(n2177) );
  XNOR U2210 ( .A(n75), .B(n2062), .Z(n2168) );
  OR U2211 ( .A(n2168), .B(n10106), .Z(n2065) );
  NANDN U2212 ( .A(n2063), .B(n10107), .Z(n2064) );
  NAND U2213 ( .A(n2065), .B(n2064), .Z(n2174) );
  XNOR U2214 ( .A(n9984), .B(n2555), .Z(n2171) );
  NANDN U2215 ( .A(n2171), .B(n9865), .Z(n2068) );
  NANDN U2216 ( .A(n2066), .B(n9930), .Z(n2067) );
  AND U2217 ( .A(n2068), .B(n2067), .Z(n2175) );
  XNOR U2218 ( .A(n2174), .B(n2175), .Z(n2176) );
  XNOR U2219 ( .A(n2177), .B(n2176), .Z(n2186) );
  NANDN U2220 ( .A(n2070), .B(n2069), .Z(n2074) );
  NAND U2221 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U2222 ( .A(n2074), .B(n2073), .Z(n2187) );
  XNOR U2223 ( .A(n2186), .B(n2187), .Z(n2188) );
  NANDN U2224 ( .A(n2076), .B(n2075), .Z(n2080) );
  NAND U2225 ( .A(n2078), .B(n2077), .Z(n2079) );
  AND U2226 ( .A(n2080), .B(n2079), .Z(n2189) );
  XNOR U2227 ( .A(n2188), .B(n2189), .Z(n2133) );
  NANDN U2228 ( .A(n2082), .B(n2081), .Z(n2086) );
  OR U2229 ( .A(n2084), .B(n2083), .Z(n2085) );
  NAND U2230 ( .A(n2086), .B(n2085), .Z(n2161) );
  XNOR U2231 ( .A(n10050), .B(n2245), .Z(n2146) );
  OR U2232 ( .A(n2146), .B(n10051), .Z(n2089) );
  NANDN U2233 ( .A(n2087), .B(n10070), .Z(n2088) );
  AND U2234 ( .A(n2089), .B(n2088), .Z(n2138) );
  NAND U2235 ( .A(b[0]), .B(a[34]), .Z(n2090) );
  XNOR U2236 ( .A(b[1]), .B(n2090), .Z(n2092) );
  NAND U2237 ( .A(a[33]), .B(n72), .Z(n2091) );
  AND U2238 ( .A(n2092), .B(n2091), .Z(n2137) );
  XOR U2239 ( .A(n2138), .B(n2137), .Z(n2140) );
  NAND U2240 ( .A(a[18]), .B(b[15]), .Z(n2139) );
  XOR U2241 ( .A(n2140), .B(n2139), .Z(n2158) );
  XNOR U2242 ( .A(n9622), .B(n2840), .Z(n2149) );
  OR U2243 ( .A(n2149), .B(n9623), .Z(n2095) );
  NANDN U2244 ( .A(n2093), .B(n9680), .Z(n2094) );
  NAND U2245 ( .A(n2095), .B(n2094), .Z(n2183) );
  XNOR U2246 ( .A(n9872), .B(n2711), .Z(n2152) );
  NANDN U2247 ( .A(n2152), .B(n9746), .Z(n2098) );
  NANDN U2248 ( .A(n2096), .B(n9747), .Z(n2097) );
  NAND U2249 ( .A(n2098), .B(n2097), .Z(n2180) );
  IV U2250 ( .A(a[32]), .Z(n2996) );
  XNOR U2251 ( .A(n74), .B(n2996), .Z(n2155) );
  NANDN U2252 ( .A(n2155), .B(n9485), .Z(n2101) );
  NANDN U2253 ( .A(n2099), .B(n9484), .Z(n2100) );
  AND U2254 ( .A(n2101), .B(n2100), .Z(n2181) );
  XNOR U2255 ( .A(n2180), .B(n2181), .Z(n2182) );
  XOR U2256 ( .A(n2183), .B(n2182), .Z(n2159) );
  XOR U2257 ( .A(n2158), .B(n2159), .Z(n2160) );
  XNOR U2258 ( .A(n2161), .B(n2160), .Z(n2131) );
  NAND U2259 ( .A(n2103), .B(n2102), .Z(n2107) );
  NAND U2260 ( .A(n2105), .B(n2104), .Z(n2106) );
  NAND U2261 ( .A(n2107), .B(n2106), .Z(n2132) );
  XOR U2262 ( .A(n2131), .B(n2132), .Z(n2134) );
  XNOR U2263 ( .A(n2133), .B(n2134), .Z(n2192) );
  NANDN U2264 ( .A(n2109), .B(n2108), .Z(n2113) );
  NAND U2265 ( .A(n2111), .B(n2110), .Z(n2112) );
  NAND U2266 ( .A(n2113), .B(n2112), .Z(n2193) );
  XNOR U2267 ( .A(n2192), .B(n2193), .Z(n2194) );
  XOR U2268 ( .A(n2195), .B(n2194), .Z(n2125) );
  NANDN U2269 ( .A(n2115), .B(n2114), .Z(n2119) );
  NANDN U2270 ( .A(n2117), .B(n2116), .Z(n2118) );
  NAND U2271 ( .A(n2119), .B(n2118), .Z(n2126) );
  XNOR U2272 ( .A(n2125), .B(n2126), .Z(n2127) );
  XNOR U2273 ( .A(n2128), .B(n2127), .Z(n2198) );
  XNOR U2274 ( .A(n2198), .B(sreg[146]), .Z(n2200) );
  NAND U2275 ( .A(n2120), .B(sreg[145]), .Z(n2124) );
  OR U2276 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U2277 ( .A(n2124), .B(n2123), .Z(n2199) );
  XOR U2278 ( .A(n2200), .B(n2199), .Z(c[146]) );
  NANDN U2279 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U2280 ( .A(n2128), .B(n2127), .Z(n2129) );
  NAND U2281 ( .A(n2130), .B(n2129), .Z(n2206) );
  NANDN U2282 ( .A(n2132), .B(n2131), .Z(n2136) );
  OR U2283 ( .A(n2134), .B(n2133), .Z(n2135) );
  NAND U2284 ( .A(n2136), .B(n2135), .Z(n2273) );
  NANDN U2285 ( .A(n2138), .B(n2137), .Z(n2142) );
  OR U2286 ( .A(n2140), .B(n2139), .Z(n2141) );
  NAND U2287 ( .A(n2142), .B(n2141), .Z(n2239) );
  NAND U2288 ( .A(b[0]), .B(a[35]), .Z(n2143) );
  XNOR U2289 ( .A(b[1]), .B(n2143), .Z(n2145) );
  NAND U2290 ( .A(a[34]), .B(n72), .Z(n2144) );
  AND U2291 ( .A(n2145), .B(n2144), .Z(n2215) );
  XNOR U2292 ( .A(n10050), .B(n2323), .Z(n2221) );
  OR U2293 ( .A(n2221), .B(n10051), .Z(n2148) );
  NANDN U2294 ( .A(n2146), .B(n10070), .Z(n2147) );
  AND U2295 ( .A(n2148), .B(n2147), .Z(n2216) );
  XOR U2296 ( .A(n2215), .B(n2216), .Z(n2218) );
  NAND U2297 ( .A(a[19]), .B(b[15]), .Z(n2217) );
  XOR U2298 ( .A(n2218), .B(n2217), .Z(n2236) );
  XNOR U2299 ( .A(n9622), .B(n2918), .Z(n2227) );
  OR U2300 ( .A(n2227), .B(n9623), .Z(n2151) );
  NANDN U2301 ( .A(n2149), .B(n9680), .Z(n2150) );
  NAND U2302 ( .A(n2151), .B(n2150), .Z(n2261) );
  XNOR U2303 ( .A(n9872), .B(n2762), .Z(n2230) );
  NANDN U2304 ( .A(n2230), .B(n9746), .Z(n2154) );
  NANDN U2305 ( .A(n2152), .B(n9747), .Z(n2153) );
  NAND U2306 ( .A(n2154), .B(n2153), .Z(n2258) );
  IV U2307 ( .A(a[33]), .Z(n3074) );
  XNOR U2308 ( .A(n74), .B(n3074), .Z(n2233) );
  NANDN U2309 ( .A(n2233), .B(n9485), .Z(n2157) );
  NANDN U2310 ( .A(n2155), .B(n9484), .Z(n2156) );
  AND U2311 ( .A(n2157), .B(n2156), .Z(n2259) );
  XNOR U2312 ( .A(n2258), .B(n2259), .Z(n2260) );
  XOR U2313 ( .A(n2261), .B(n2260), .Z(n2237) );
  XOR U2314 ( .A(n2236), .B(n2237), .Z(n2238) );
  XNOR U2315 ( .A(n2239), .B(n2238), .Z(n2209) );
  NAND U2316 ( .A(n2159), .B(n2158), .Z(n2163) );
  NAND U2317 ( .A(n2161), .B(n2160), .Z(n2162) );
  NAND U2318 ( .A(n2163), .B(n2162), .Z(n2210) );
  XOR U2319 ( .A(n2209), .B(n2210), .Z(n2212) );
  XNOR U2320 ( .A(n9967), .B(n2450), .Z(n2242) );
  OR U2321 ( .A(n2242), .B(n10020), .Z(n2166) );
  NANDN U2322 ( .A(n2164), .B(n9968), .Z(n2165) );
  NAND U2323 ( .A(n2166), .B(n2165), .Z(n2255) );
  XNOR U2324 ( .A(n75), .B(n2167), .Z(n2246) );
  OR U2325 ( .A(n2246), .B(n10106), .Z(n2170) );
  NANDN U2326 ( .A(n2168), .B(n10107), .Z(n2169) );
  NAND U2327 ( .A(n2170), .B(n2169), .Z(n2252) );
  XNOR U2328 ( .A(n9984), .B(n2606), .Z(n2249) );
  NANDN U2329 ( .A(n2249), .B(n9865), .Z(n2173) );
  NANDN U2330 ( .A(n2171), .B(n9930), .Z(n2172) );
  AND U2331 ( .A(n2173), .B(n2172), .Z(n2253) );
  XNOR U2332 ( .A(n2252), .B(n2253), .Z(n2254) );
  XNOR U2333 ( .A(n2255), .B(n2254), .Z(n2264) );
  NANDN U2334 ( .A(n2175), .B(n2174), .Z(n2179) );
  NAND U2335 ( .A(n2177), .B(n2176), .Z(n2178) );
  NAND U2336 ( .A(n2179), .B(n2178), .Z(n2265) );
  XNOR U2337 ( .A(n2264), .B(n2265), .Z(n2266) );
  NANDN U2338 ( .A(n2181), .B(n2180), .Z(n2185) );
  NAND U2339 ( .A(n2183), .B(n2182), .Z(n2184) );
  AND U2340 ( .A(n2185), .B(n2184), .Z(n2267) );
  XNOR U2341 ( .A(n2266), .B(n2267), .Z(n2211) );
  XNOR U2342 ( .A(n2212), .B(n2211), .Z(n2270) );
  NANDN U2343 ( .A(n2187), .B(n2186), .Z(n2191) );
  NAND U2344 ( .A(n2189), .B(n2188), .Z(n2190) );
  NAND U2345 ( .A(n2191), .B(n2190), .Z(n2271) );
  XNOR U2346 ( .A(n2270), .B(n2271), .Z(n2272) );
  XOR U2347 ( .A(n2273), .B(n2272), .Z(n2203) );
  NANDN U2348 ( .A(n2193), .B(n2192), .Z(n2197) );
  NANDN U2349 ( .A(n2195), .B(n2194), .Z(n2196) );
  NAND U2350 ( .A(n2197), .B(n2196), .Z(n2204) );
  XNOR U2351 ( .A(n2203), .B(n2204), .Z(n2205) );
  XNOR U2352 ( .A(n2206), .B(n2205), .Z(n2276) );
  XNOR U2353 ( .A(n2276), .B(sreg[147]), .Z(n2278) );
  NAND U2354 ( .A(n2198), .B(sreg[146]), .Z(n2202) );
  OR U2355 ( .A(n2200), .B(n2199), .Z(n2201) );
  AND U2356 ( .A(n2202), .B(n2201), .Z(n2277) );
  XOR U2357 ( .A(n2278), .B(n2277), .Z(c[147]) );
  NANDN U2358 ( .A(n2204), .B(n2203), .Z(n2208) );
  NAND U2359 ( .A(n2206), .B(n2205), .Z(n2207) );
  NAND U2360 ( .A(n2208), .B(n2207), .Z(n2284) );
  NANDN U2361 ( .A(n2210), .B(n2209), .Z(n2214) );
  OR U2362 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U2363 ( .A(n2214), .B(n2213), .Z(n2351) );
  NANDN U2364 ( .A(n2216), .B(n2215), .Z(n2220) );
  OR U2365 ( .A(n2218), .B(n2217), .Z(n2219) );
  NAND U2366 ( .A(n2220), .B(n2219), .Z(n2317) );
  XNOR U2367 ( .A(n10050), .B(n2374), .Z(n2299) );
  OR U2368 ( .A(n2299), .B(n10051), .Z(n2223) );
  NANDN U2369 ( .A(n2221), .B(n10070), .Z(n2222) );
  AND U2370 ( .A(n2223), .B(n2222), .Z(n2294) );
  NAND U2371 ( .A(b[0]), .B(a[36]), .Z(n2224) );
  XNOR U2372 ( .A(b[1]), .B(n2224), .Z(n2226) );
  NAND U2373 ( .A(a[35]), .B(n72), .Z(n2225) );
  AND U2374 ( .A(n2226), .B(n2225), .Z(n2293) );
  XOR U2375 ( .A(n2294), .B(n2293), .Z(n2296) );
  NAND U2376 ( .A(a[20]), .B(b[15]), .Z(n2295) );
  XOR U2377 ( .A(n2296), .B(n2295), .Z(n2314) );
  XNOR U2378 ( .A(n9622), .B(n2996), .Z(n2305) );
  OR U2379 ( .A(n2305), .B(n9623), .Z(n2229) );
  NANDN U2380 ( .A(n2227), .B(n9680), .Z(n2228) );
  NAND U2381 ( .A(n2229), .B(n2228), .Z(n2339) );
  XNOR U2382 ( .A(n9872), .B(n2840), .Z(n2308) );
  NANDN U2383 ( .A(n2308), .B(n9746), .Z(n2232) );
  NANDN U2384 ( .A(n2230), .B(n9747), .Z(n2231) );
  NAND U2385 ( .A(n2232), .B(n2231), .Z(n2336) );
  IV U2386 ( .A(a[34]), .Z(n3179) );
  XNOR U2387 ( .A(n74), .B(n3179), .Z(n2311) );
  NANDN U2388 ( .A(n2311), .B(n9485), .Z(n2235) );
  NANDN U2389 ( .A(n2233), .B(n9484), .Z(n2234) );
  AND U2390 ( .A(n2235), .B(n2234), .Z(n2337) );
  XNOR U2391 ( .A(n2336), .B(n2337), .Z(n2338) );
  XOR U2392 ( .A(n2339), .B(n2338), .Z(n2315) );
  XOR U2393 ( .A(n2314), .B(n2315), .Z(n2316) );
  XNOR U2394 ( .A(n2317), .B(n2316), .Z(n2287) );
  NAND U2395 ( .A(n2237), .B(n2236), .Z(n2241) );
  NAND U2396 ( .A(n2239), .B(n2238), .Z(n2240) );
  NAND U2397 ( .A(n2241), .B(n2240), .Z(n2288) );
  XOR U2398 ( .A(n2287), .B(n2288), .Z(n2290) );
  XNOR U2399 ( .A(n9967), .B(n2555), .Z(n2320) );
  OR U2400 ( .A(n2320), .B(n10020), .Z(n2244) );
  NANDN U2401 ( .A(n2242), .B(n9968), .Z(n2243) );
  NAND U2402 ( .A(n2244), .B(n2243), .Z(n2333) );
  XNOR U2403 ( .A(n75), .B(n2245), .Z(n2324) );
  OR U2404 ( .A(n2324), .B(n10106), .Z(n2248) );
  NANDN U2405 ( .A(n2246), .B(n10107), .Z(n2247) );
  NAND U2406 ( .A(n2248), .B(n2247), .Z(n2330) );
  XNOR U2407 ( .A(n9984), .B(n2711), .Z(n2327) );
  NANDN U2408 ( .A(n2327), .B(n9865), .Z(n2251) );
  NANDN U2409 ( .A(n2249), .B(n9930), .Z(n2250) );
  AND U2410 ( .A(n2251), .B(n2250), .Z(n2331) );
  XNOR U2411 ( .A(n2330), .B(n2331), .Z(n2332) );
  XNOR U2412 ( .A(n2333), .B(n2332), .Z(n2342) );
  NANDN U2413 ( .A(n2253), .B(n2252), .Z(n2257) );
  NAND U2414 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2415 ( .A(n2257), .B(n2256), .Z(n2343) );
  XNOR U2416 ( .A(n2342), .B(n2343), .Z(n2344) );
  NANDN U2417 ( .A(n2259), .B(n2258), .Z(n2263) );
  NAND U2418 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U2419 ( .A(n2263), .B(n2262), .Z(n2345) );
  XNOR U2420 ( .A(n2344), .B(n2345), .Z(n2289) );
  XNOR U2421 ( .A(n2290), .B(n2289), .Z(n2348) );
  NANDN U2422 ( .A(n2265), .B(n2264), .Z(n2269) );
  NAND U2423 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U2424 ( .A(n2269), .B(n2268), .Z(n2349) );
  XNOR U2425 ( .A(n2348), .B(n2349), .Z(n2350) );
  XOR U2426 ( .A(n2351), .B(n2350), .Z(n2281) );
  NANDN U2427 ( .A(n2271), .B(n2270), .Z(n2275) );
  NANDN U2428 ( .A(n2273), .B(n2272), .Z(n2274) );
  NAND U2429 ( .A(n2275), .B(n2274), .Z(n2282) );
  XNOR U2430 ( .A(n2281), .B(n2282), .Z(n2283) );
  XNOR U2431 ( .A(n2284), .B(n2283), .Z(n2354) );
  XNOR U2432 ( .A(n2354), .B(sreg[148]), .Z(n2356) );
  NAND U2433 ( .A(n2276), .B(sreg[147]), .Z(n2280) );
  OR U2434 ( .A(n2278), .B(n2277), .Z(n2279) );
  AND U2435 ( .A(n2280), .B(n2279), .Z(n2355) );
  XOR U2436 ( .A(n2356), .B(n2355), .Z(c[148]) );
  NANDN U2437 ( .A(n2282), .B(n2281), .Z(n2286) );
  NAND U2438 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U2439 ( .A(n2286), .B(n2285), .Z(n2362) );
  NANDN U2440 ( .A(n2288), .B(n2287), .Z(n2292) );
  OR U2441 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U2442 ( .A(n2292), .B(n2291), .Z(n2427) );
  NANDN U2443 ( .A(n2294), .B(n2293), .Z(n2298) );
  OR U2444 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2445 ( .A(n2298), .B(n2297), .Z(n2417) );
  XNOR U2446 ( .A(n10050), .B(n2450), .Z(n2402) );
  OR U2447 ( .A(n2402), .B(n10051), .Z(n2301) );
  NANDN U2448 ( .A(n2299), .B(n10070), .Z(n2300) );
  NAND U2449 ( .A(n2301), .B(n2300), .Z(n2393) );
  AND U2450 ( .A(a[37]), .B(b[0]), .Z(n2302) );
  XOR U2451 ( .A(b[1]), .B(n2302), .Z(n2304) );
  NAND U2452 ( .A(a[36]), .B(n72), .Z(n2303) );
  NAND U2453 ( .A(n2304), .B(n2303), .Z(n2394) );
  XNOR U2454 ( .A(n2393), .B(n2394), .Z(n2395) );
  NAND U2455 ( .A(a[21]), .B(b[15]), .Z(n2396) );
  XOR U2456 ( .A(n2395), .B(n2396), .Z(n2414) );
  XNOR U2457 ( .A(n9622), .B(n3074), .Z(n2405) );
  OR U2458 ( .A(n2405), .B(n9623), .Z(n2307) );
  NANDN U2459 ( .A(n2305), .B(n9680), .Z(n2306) );
  NAND U2460 ( .A(n2307), .B(n2306), .Z(n2390) );
  XNOR U2461 ( .A(n9872), .B(n2918), .Z(n2408) );
  NANDN U2462 ( .A(n2408), .B(n9746), .Z(n2310) );
  NANDN U2463 ( .A(n2308), .B(n9747), .Z(n2309) );
  NAND U2464 ( .A(n2310), .B(n2309), .Z(n2387) );
  IV U2465 ( .A(a[35]), .Z(n3257) );
  XNOR U2466 ( .A(n74), .B(n3257), .Z(n2411) );
  NANDN U2467 ( .A(n2411), .B(n9485), .Z(n2313) );
  NANDN U2468 ( .A(n2311), .B(n9484), .Z(n2312) );
  AND U2469 ( .A(n2313), .B(n2312), .Z(n2388) );
  XNOR U2470 ( .A(n2387), .B(n2388), .Z(n2389) );
  XOR U2471 ( .A(n2390), .B(n2389), .Z(n2415) );
  XNOR U2472 ( .A(n2414), .B(n2415), .Z(n2416) );
  XNOR U2473 ( .A(n2417), .B(n2416), .Z(n2365) );
  NAND U2474 ( .A(n2315), .B(n2314), .Z(n2319) );
  NAND U2475 ( .A(n2317), .B(n2316), .Z(n2318) );
  NAND U2476 ( .A(n2319), .B(n2318), .Z(n2366) );
  XOR U2477 ( .A(n2365), .B(n2366), .Z(n2368) );
  XNOR U2478 ( .A(n9967), .B(n2606), .Z(n2371) );
  OR U2479 ( .A(n2371), .B(n10020), .Z(n2322) );
  NANDN U2480 ( .A(n2320), .B(n9968), .Z(n2321) );
  NAND U2481 ( .A(n2322), .B(n2321), .Z(n2384) );
  XNOR U2482 ( .A(n75), .B(n2323), .Z(n2375) );
  OR U2483 ( .A(n2375), .B(n10106), .Z(n2326) );
  NANDN U2484 ( .A(n2324), .B(n10107), .Z(n2325) );
  NAND U2485 ( .A(n2326), .B(n2325), .Z(n2381) );
  XNOR U2486 ( .A(n9984), .B(n2762), .Z(n2378) );
  NANDN U2487 ( .A(n2378), .B(n9865), .Z(n2329) );
  NANDN U2488 ( .A(n2327), .B(n9930), .Z(n2328) );
  AND U2489 ( .A(n2329), .B(n2328), .Z(n2382) );
  XNOR U2490 ( .A(n2381), .B(n2382), .Z(n2383) );
  XNOR U2491 ( .A(n2384), .B(n2383), .Z(n2418) );
  NANDN U2492 ( .A(n2331), .B(n2330), .Z(n2335) );
  NAND U2493 ( .A(n2333), .B(n2332), .Z(n2334) );
  NAND U2494 ( .A(n2335), .B(n2334), .Z(n2419) );
  XNOR U2495 ( .A(n2418), .B(n2419), .Z(n2420) );
  NANDN U2496 ( .A(n2337), .B(n2336), .Z(n2341) );
  NAND U2497 ( .A(n2339), .B(n2338), .Z(n2340) );
  AND U2498 ( .A(n2341), .B(n2340), .Z(n2421) );
  XNOR U2499 ( .A(n2420), .B(n2421), .Z(n2367) );
  XNOR U2500 ( .A(n2368), .B(n2367), .Z(n2424) );
  NANDN U2501 ( .A(n2343), .B(n2342), .Z(n2347) );
  NAND U2502 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U2503 ( .A(n2347), .B(n2346), .Z(n2425) );
  XNOR U2504 ( .A(n2424), .B(n2425), .Z(n2426) );
  XOR U2505 ( .A(n2427), .B(n2426), .Z(n2359) );
  NANDN U2506 ( .A(n2349), .B(n2348), .Z(n2353) );
  NANDN U2507 ( .A(n2351), .B(n2350), .Z(n2352) );
  NAND U2508 ( .A(n2353), .B(n2352), .Z(n2360) );
  XNOR U2509 ( .A(n2359), .B(n2360), .Z(n2361) );
  XNOR U2510 ( .A(n2362), .B(n2361), .Z(n2430) );
  XNOR U2511 ( .A(n2430), .B(sreg[149]), .Z(n2432) );
  NAND U2512 ( .A(n2354), .B(sreg[148]), .Z(n2358) );
  OR U2513 ( .A(n2356), .B(n2355), .Z(n2357) );
  AND U2514 ( .A(n2358), .B(n2357), .Z(n2431) );
  XOR U2515 ( .A(n2432), .B(n2431), .Z(c[149]) );
  NANDN U2516 ( .A(n2360), .B(n2359), .Z(n2364) );
  NAND U2517 ( .A(n2362), .B(n2361), .Z(n2363) );
  NAND U2518 ( .A(n2364), .B(n2363), .Z(n2438) );
  NANDN U2519 ( .A(n2366), .B(n2365), .Z(n2370) );
  OR U2520 ( .A(n2368), .B(n2367), .Z(n2369) );
  NAND U2521 ( .A(n2370), .B(n2369), .Z(n2505) );
  XNOR U2522 ( .A(n9967), .B(n2711), .Z(n2447) );
  OR U2523 ( .A(n2447), .B(n10020), .Z(n2373) );
  NANDN U2524 ( .A(n2371), .B(n9968), .Z(n2372) );
  NAND U2525 ( .A(n2373), .B(n2372), .Z(n2460) );
  XNOR U2526 ( .A(n75), .B(n2374), .Z(n2451) );
  OR U2527 ( .A(n2451), .B(n10106), .Z(n2377) );
  NANDN U2528 ( .A(n2375), .B(n10107), .Z(n2376) );
  NAND U2529 ( .A(n2377), .B(n2376), .Z(n2457) );
  XNOR U2530 ( .A(n9984), .B(n2840), .Z(n2454) );
  NANDN U2531 ( .A(n2454), .B(n9865), .Z(n2380) );
  NANDN U2532 ( .A(n2378), .B(n9930), .Z(n2379) );
  AND U2533 ( .A(n2380), .B(n2379), .Z(n2458) );
  XNOR U2534 ( .A(n2457), .B(n2458), .Z(n2459) );
  XNOR U2535 ( .A(n2460), .B(n2459), .Z(n2496) );
  NANDN U2536 ( .A(n2382), .B(n2381), .Z(n2386) );
  NAND U2537 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U2538 ( .A(n2386), .B(n2385), .Z(n2497) );
  XNOR U2539 ( .A(n2496), .B(n2497), .Z(n2498) );
  NANDN U2540 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U2541 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U2542 ( .A(n2392), .B(n2391), .Z(n2499) );
  XNOR U2543 ( .A(n2498), .B(n2499), .Z(n2443) );
  NANDN U2544 ( .A(n2394), .B(n2393), .Z(n2398) );
  NANDN U2545 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U2546 ( .A(n2398), .B(n2397), .Z(n2493) );
  NAND U2547 ( .A(b[0]), .B(a[38]), .Z(n2399) );
  XNOR U2548 ( .A(b[1]), .B(n2399), .Z(n2401) );
  NAND U2549 ( .A(a[37]), .B(n72), .Z(n2400) );
  AND U2550 ( .A(n2401), .B(n2400), .Z(n2469) );
  XNOR U2551 ( .A(n10050), .B(n2555), .Z(n2478) );
  OR U2552 ( .A(n2478), .B(n10051), .Z(n2404) );
  NANDN U2553 ( .A(n2402), .B(n10070), .Z(n2403) );
  AND U2554 ( .A(n2404), .B(n2403), .Z(n2470) );
  XOR U2555 ( .A(n2469), .B(n2470), .Z(n2472) );
  NAND U2556 ( .A(a[22]), .B(b[15]), .Z(n2471) );
  XOR U2557 ( .A(n2472), .B(n2471), .Z(n2490) );
  XNOR U2558 ( .A(n9622), .B(n3179), .Z(n2481) );
  OR U2559 ( .A(n2481), .B(n9623), .Z(n2407) );
  NANDN U2560 ( .A(n2405), .B(n9680), .Z(n2406) );
  NAND U2561 ( .A(n2407), .B(n2406), .Z(n2466) );
  XNOR U2562 ( .A(n9872), .B(n2996), .Z(n2484) );
  NANDN U2563 ( .A(n2484), .B(n9746), .Z(n2410) );
  NANDN U2564 ( .A(n2408), .B(n9747), .Z(n2409) );
  NAND U2565 ( .A(n2410), .B(n2409), .Z(n2463) );
  IV U2566 ( .A(a[36]), .Z(n3308) );
  XNOR U2567 ( .A(n74), .B(n3308), .Z(n2487) );
  NANDN U2568 ( .A(n2487), .B(n9485), .Z(n2413) );
  NANDN U2569 ( .A(n2411), .B(n9484), .Z(n2412) );
  AND U2570 ( .A(n2413), .B(n2412), .Z(n2464) );
  XNOR U2571 ( .A(n2463), .B(n2464), .Z(n2465) );
  XOR U2572 ( .A(n2466), .B(n2465), .Z(n2491) );
  XOR U2573 ( .A(n2490), .B(n2491), .Z(n2492) );
  XNOR U2574 ( .A(n2493), .B(n2492), .Z(n2441) );
  XOR U2575 ( .A(n2441), .B(n2442), .Z(n2444) );
  XNOR U2576 ( .A(n2443), .B(n2444), .Z(n2502) );
  NANDN U2577 ( .A(n2419), .B(n2418), .Z(n2423) );
  NAND U2578 ( .A(n2421), .B(n2420), .Z(n2422) );
  NAND U2579 ( .A(n2423), .B(n2422), .Z(n2503) );
  XNOR U2580 ( .A(n2502), .B(n2503), .Z(n2504) );
  XOR U2581 ( .A(n2505), .B(n2504), .Z(n2435) );
  NANDN U2582 ( .A(n2425), .B(n2424), .Z(n2429) );
  NANDN U2583 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U2584 ( .A(n2429), .B(n2428), .Z(n2436) );
  XNOR U2585 ( .A(n2435), .B(n2436), .Z(n2437) );
  XNOR U2586 ( .A(n2438), .B(n2437), .Z(n2508) );
  XNOR U2587 ( .A(n2508), .B(sreg[150]), .Z(n2510) );
  NAND U2588 ( .A(n2430), .B(sreg[149]), .Z(n2434) );
  OR U2589 ( .A(n2432), .B(n2431), .Z(n2433) );
  AND U2590 ( .A(n2434), .B(n2433), .Z(n2509) );
  XOR U2591 ( .A(n2510), .B(n2509), .Z(c[150]) );
  NANDN U2592 ( .A(n2436), .B(n2435), .Z(n2440) );
  NAND U2593 ( .A(n2438), .B(n2437), .Z(n2439) );
  NAND U2594 ( .A(n2440), .B(n2439), .Z(n2516) );
  NANDN U2595 ( .A(n2442), .B(n2441), .Z(n2446) );
  OR U2596 ( .A(n2444), .B(n2443), .Z(n2445) );
  NAND U2597 ( .A(n2446), .B(n2445), .Z(n2583) );
  XNOR U2598 ( .A(n9967), .B(n2762), .Z(n2552) );
  OR U2599 ( .A(n2552), .B(n10020), .Z(n2449) );
  NANDN U2600 ( .A(n2447), .B(n9968), .Z(n2448) );
  NAND U2601 ( .A(n2449), .B(n2448), .Z(n2565) );
  XNOR U2602 ( .A(n75), .B(n2450), .Z(n2556) );
  OR U2603 ( .A(n2556), .B(n10106), .Z(n2453) );
  NANDN U2604 ( .A(n2451), .B(n10107), .Z(n2452) );
  NAND U2605 ( .A(n2453), .B(n2452), .Z(n2562) );
  XNOR U2606 ( .A(n9984), .B(n2918), .Z(n2559) );
  NANDN U2607 ( .A(n2559), .B(n9865), .Z(n2456) );
  NANDN U2608 ( .A(n2454), .B(n9930), .Z(n2455) );
  AND U2609 ( .A(n2456), .B(n2455), .Z(n2563) );
  XNOR U2610 ( .A(n2562), .B(n2563), .Z(n2564) );
  XNOR U2611 ( .A(n2565), .B(n2564), .Z(n2574) );
  NANDN U2612 ( .A(n2458), .B(n2457), .Z(n2462) );
  NAND U2613 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U2614 ( .A(n2462), .B(n2461), .Z(n2575) );
  XNOR U2615 ( .A(n2574), .B(n2575), .Z(n2576) );
  NANDN U2616 ( .A(n2464), .B(n2463), .Z(n2468) );
  NAND U2617 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2618 ( .A(n2468), .B(n2467), .Z(n2577) );
  XNOR U2619 ( .A(n2576), .B(n2577), .Z(n2521) );
  NANDN U2620 ( .A(n2470), .B(n2469), .Z(n2474) );
  OR U2621 ( .A(n2472), .B(n2471), .Z(n2473) );
  NAND U2622 ( .A(n2474), .B(n2473), .Z(n2549) );
  NAND U2623 ( .A(b[0]), .B(a[39]), .Z(n2475) );
  XNOR U2624 ( .A(b[1]), .B(n2475), .Z(n2477) );
  NAND U2625 ( .A(a[38]), .B(n72), .Z(n2476) );
  AND U2626 ( .A(n2477), .B(n2476), .Z(n2525) );
  XNOR U2627 ( .A(n10050), .B(n2606), .Z(n2534) );
  OR U2628 ( .A(n2534), .B(n10051), .Z(n2480) );
  NANDN U2629 ( .A(n2478), .B(n10070), .Z(n2479) );
  AND U2630 ( .A(n2480), .B(n2479), .Z(n2526) );
  XOR U2631 ( .A(n2525), .B(n2526), .Z(n2528) );
  NAND U2632 ( .A(a[23]), .B(b[15]), .Z(n2527) );
  XOR U2633 ( .A(n2528), .B(n2527), .Z(n2546) );
  XNOR U2634 ( .A(n9622), .B(n3257), .Z(n2537) );
  OR U2635 ( .A(n2537), .B(n9623), .Z(n2483) );
  NANDN U2636 ( .A(n2481), .B(n9680), .Z(n2482) );
  NAND U2637 ( .A(n2483), .B(n2482), .Z(n2571) );
  XNOR U2638 ( .A(n9872), .B(n3074), .Z(n2540) );
  NANDN U2639 ( .A(n2540), .B(n9746), .Z(n2486) );
  NANDN U2640 ( .A(n2484), .B(n9747), .Z(n2485) );
  NAND U2641 ( .A(n2486), .B(n2485), .Z(n2568) );
  IV U2642 ( .A(a[37]), .Z(n3386) );
  XNOR U2643 ( .A(n74), .B(n3386), .Z(n2543) );
  NANDN U2644 ( .A(n2543), .B(n9485), .Z(n2489) );
  NANDN U2645 ( .A(n2487), .B(n9484), .Z(n2488) );
  AND U2646 ( .A(n2489), .B(n2488), .Z(n2569) );
  XNOR U2647 ( .A(n2568), .B(n2569), .Z(n2570) );
  XOR U2648 ( .A(n2571), .B(n2570), .Z(n2547) );
  XOR U2649 ( .A(n2546), .B(n2547), .Z(n2548) );
  XNOR U2650 ( .A(n2549), .B(n2548), .Z(n2519) );
  NAND U2651 ( .A(n2491), .B(n2490), .Z(n2495) );
  NAND U2652 ( .A(n2493), .B(n2492), .Z(n2494) );
  NAND U2653 ( .A(n2495), .B(n2494), .Z(n2520) );
  XOR U2654 ( .A(n2519), .B(n2520), .Z(n2522) );
  XNOR U2655 ( .A(n2521), .B(n2522), .Z(n2580) );
  NANDN U2656 ( .A(n2497), .B(n2496), .Z(n2501) );
  NAND U2657 ( .A(n2499), .B(n2498), .Z(n2500) );
  NAND U2658 ( .A(n2501), .B(n2500), .Z(n2581) );
  XNOR U2659 ( .A(n2580), .B(n2581), .Z(n2582) );
  XOR U2660 ( .A(n2583), .B(n2582), .Z(n2513) );
  NANDN U2661 ( .A(n2503), .B(n2502), .Z(n2507) );
  NANDN U2662 ( .A(n2505), .B(n2504), .Z(n2506) );
  NAND U2663 ( .A(n2507), .B(n2506), .Z(n2514) );
  XNOR U2664 ( .A(n2513), .B(n2514), .Z(n2515) );
  XNOR U2665 ( .A(n2516), .B(n2515), .Z(n2586) );
  XNOR U2666 ( .A(n2586), .B(sreg[151]), .Z(n2588) );
  NAND U2667 ( .A(n2508), .B(sreg[150]), .Z(n2512) );
  OR U2668 ( .A(n2510), .B(n2509), .Z(n2511) );
  AND U2669 ( .A(n2512), .B(n2511), .Z(n2587) );
  XOR U2670 ( .A(n2588), .B(n2587), .Z(c[151]) );
  NANDN U2671 ( .A(n2514), .B(n2513), .Z(n2518) );
  NAND U2672 ( .A(n2516), .B(n2515), .Z(n2517) );
  NAND U2673 ( .A(n2518), .B(n2517), .Z(n2594) );
  NANDN U2674 ( .A(n2520), .B(n2519), .Z(n2524) );
  OR U2675 ( .A(n2522), .B(n2521), .Z(n2523) );
  NAND U2676 ( .A(n2524), .B(n2523), .Z(n2661) );
  NANDN U2677 ( .A(n2526), .B(n2525), .Z(n2530) );
  OR U2678 ( .A(n2528), .B(n2527), .Z(n2529) );
  NAND U2679 ( .A(n2530), .B(n2529), .Z(n2649) );
  NAND U2680 ( .A(b[0]), .B(a[40]), .Z(n2531) );
  XNOR U2681 ( .A(b[1]), .B(n2531), .Z(n2533) );
  NAND U2682 ( .A(a[39]), .B(n72), .Z(n2532) );
  AND U2683 ( .A(n2533), .B(n2532), .Z(n2625) );
  XNOR U2684 ( .A(n10050), .B(n2711), .Z(n2631) );
  OR U2685 ( .A(n2631), .B(n10051), .Z(n2536) );
  NANDN U2686 ( .A(n2534), .B(n10070), .Z(n2535) );
  AND U2687 ( .A(n2536), .B(n2535), .Z(n2626) );
  XOR U2688 ( .A(n2625), .B(n2626), .Z(n2628) );
  NAND U2689 ( .A(a[24]), .B(b[15]), .Z(n2627) );
  XOR U2690 ( .A(n2628), .B(n2627), .Z(n2646) );
  XNOR U2691 ( .A(n9622), .B(n3308), .Z(n2637) );
  OR U2692 ( .A(n2637), .B(n9623), .Z(n2539) );
  NANDN U2693 ( .A(n2537), .B(n9680), .Z(n2538) );
  NAND U2694 ( .A(n2539), .B(n2538), .Z(n2622) );
  XNOR U2695 ( .A(n9872), .B(n3179), .Z(n2640) );
  NANDN U2696 ( .A(n2640), .B(n9746), .Z(n2542) );
  NANDN U2697 ( .A(n2540), .B(n9747), .Z(n2541) );
  NAND U2698 ( .A(n2542), .B(n2541), .Z(n2619) );
  IV U2699 ( .A(a[38]), .Z(n3464) );
  XNOR U2700 ( .A(n74), .B(n3464), .Z(n2643) );
  NANDN U2701 ( .A(n2643), .B(n9485), .Z(n2545) );
  NANDN U2702 ( .A(n2543), .B(n9484), .Z(n2544) );
  AND U2703 ( .A(n2545), .B(n2544), .Z(n2620) );
  XNOR U2704 ( .A(n2619), .B(n2620), .Z(n2621) );
  XOR U2705 ( .A(n2622), .B(n2621), .Z(n2647) );
  XOR U2706 ( .A(n2646), .B(n2647), .Z(n2648) );
  XNOR U2707 ( .A(n2649), .B(n2648), .Z(n2597) );
  NAND U2708 ( .A(n2547), .B(n2546), .Z(n2551) );
  NAND U2709 ( .A(n2549), .B(n2548), .Z(n2550) );
  NAND U2710 ( .A(n2551), .B(n2550), .Z(n2598) );
  XOR U2711 ( .A(n2597), .B(n2598), .Z(n2600) );
  XNOR U2712 ( .A(n9967), .B(n2840), .Z(n2603) );
  OR U2713 ( .A(n2603), .B(n10020), .Z(n2554) );
  NANDN U2714 ( .A(n2552), .B(n9968), .Z(n2553) );
  NAND U2715 ( .A(n2554), .B(n2553), .Z(n2616) );
  XNOR U2716 ( .A(n75), .B(n2555), .Z(n2607) );
  OR U2717 ( .A(n2607), .B(n10106), .Z(n2558) );
  NANDN U2718 ( .A(n2556), .B(n10107), .Z(n2557) );
  NAND U2719 ( .A(n2558), .B(n2557), .Z(n2613) );
  XNOR U2720 ( .A(n9984), .B(n2996), .Z(n2610) );
  NANDN U2721 ( .A(n2610), .B(n9865), .Z(n2561) );
  NANDN U2722 ( .A(n2559), .B(n9930), .Z(n2560) );
  AND U2723 ( .A(n2561), .B(n2560), .Z(n2614) );
  XNOR U2724 ( .A(n2613), .B(n2614), .Z(n2615) );
  XNOR U2725 ( .A(n2616), .B(n2615), .Z(n2652) );
  NANDN U2726 ( .A(n2563), .B(n2562), .Z(n2567) );
  NAND U2727 ( .A(n2565), .B(n2564), .Z(n2566) );
  NAND U2728 ( .A(n2567), .B(n2566), .Z(n2653) );
  XNOR U2729 ( .A(n2652), .B(n2653), .Z(n2654) );
  NANDN U2730 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U2731 ( .A(n2571), .B(n2570), .Z(n2572) );
  AND U2732 ( .A(n2573), .B(n2572), .Z(n2655) );
  XNOR U2733 ( .A(n2654), .B(n2655), .Z(n2599) );
  XNOR U2734 ( .A(n2600), .B(n2599), .Z(n2658) );
  NANDN U2735 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U2736 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U2737 ( .A(n2579), .B(n2578), .Z(n2659) );
  XNOR U2738 ( .A(n2658), .B(n2659), .Z(n2660) );
  XOR U2739 ( .A(n2661), .B(n2660), .Z(n2591) );
  NANDN U2740 ( .A(n2581), .B(n2580), .Z(n2585) );
  NANDN U2741 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U2742 ( .A(n2585), .B(n2584), .Z(n2592) );
  XNOR U2743 ( .A(n2591), .B(n2592), .Z(n2593) );
  XNOR U2744 ( .A(n2594), .B(n2593), .Z(n2664) );
  XNOR U2745 ( .A(n2664), .B(sreg[152]), .Z(n2666) );
  NAND U2746 ( .A(n2586), .B(sreg[151]), .Z(n2590) );
  OR U2747 ( .A(n2588), .B(n2587), .Z(n2589) );
  AND U2748 ( .A(n2590), .B(n2589), .Z(n2665) );
  XOR U2749 ( .A(n2666), .B(n2665), .Z(c[152]) );
  NANDN U2750 ( .A(n2592), .B(n2591), .Z(n2596) );
  NAND U2751 ( .A(n2594), .B(n2593), .Z(n2595) );
  NAND U2752 ( .A(n2596), .B(n2595), .Z(n2672) );
  NANDN U2753 ( .A(n2598), .B(n2597), .Z(n2602) );
  OR U2754 ( .A(n2600), .B(n2599), .Z(n2601) );
  NAND U2755 ( .A(n2602), .B(n2601), .Z(n2739) );
  XNOR U2756 ( .A(n9967), .B(n2918), .Z(n2708) );
  OR U2757 ( .A(n2708), .B(n10020), .Z(n2605) );
  NANDN U2758 ( .A(n2603), .B(n9968), .Z(n2604) );
  NAND U2759 ( .A(n2605), .B(n2604), .Z(n2721) );
  XNOR U2760 ( .A(n75), .B(n2606), .Z(n2712) );
  OR U2761 ( .A(n2712), .B(n10106), .Z(n2609) );
  NANDN U2762 ( .A(n2607), .B(n10107), .Z(n2608) );
  NAND U2763 ( .A(n2609), .B(n2608), .Z(n2718) );
  XNOR U2764 ( .A(n9984), .B(n3074), .Z(n2715) );
  NANDN U2765 ( .A(n2715), .B(n9865), .Z(n2612) );
  NANDN U2766 ( .A(n2610), .B(n9930), .Z(n2611) );
  AND U2767 ( .A(n2612), .B(n2611), .Z(n2719) );
  XNOR U2768 ( .A(n2718), .B(n2719), .Z(n2720) );
  XNOR U2769 ( .A(n2721), .B(n2720), .Z(n2730) );
  NANDN U2770 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U2771 ( .A(n2616), .B(n2615), .Z(n2617) );
  NAND U2772 ( .A(n2618), .B(n2617), .Z(n2731) );
  XNOR U2773 ( .A(n2730), .B(n2731), .Z(n2732) );
  NANDN U2774 ( .A(n2620), .B(n2619), .Z(n2624) );
  NAND U2775 ( .A(n2622), .B(n2621), .Z(n2623) );
  AND U2776 ( .A(n2624), .B(n2623), .Z(n2733) );
  XNOR U2777 ( .A(n2732), .B(n2733), .Z(n2677) );
  NANDN U2778 ( .A(n2626), .B(n2625), .Z(n2630) );
  OR U2779 ( .A(n2628), .B(n2627), .Z(n2629) );
  NAND U2780 ( .A(n2630), .B(n2629), .Z(n2705) );
  XNOR U2781 ( .A(n10050), .B(n2762), .Z(n2687) );
  OR U2782 ( .A(n2687), .B(n10051), .Z(n2633) );
  NANDN U2783 ( .A(n2631), .B(n10070), .Z(n2632) );
  AND U2784 ( .A(n2633), .B(n2632), .Z(n2682) );
  NAND U2785 ( .A(b[0]), .B(a[41]), .Z(n2634) );
  XNOR U2786 ( .A(b[1]), .B(n2634), .Z(n2636) );
  NAND U2787 ( .A(a[40]), .B(n72), .Z(n2635) );
  AND U2788 ( .A(n2636), .B(n2635), .Z(n2681) );
  XOR U2789 ( .A(n2682), .B(n2681), .Z(n2684) );
  NAND U2790 ( .A(a[25]), .B(b[15]), .Z(n2683) );
  XOR U2791 ( .A(n2684), .B(n2683), .Z(n2702) );
  XNOR U2792 ( .A(n9622), .B(n3386), .Z(n2693) );
  OR U2793 ( .A(n2693), .B(n9623), .Z(n2639) );
  NANDN U2794 ( .A(n2637), .B(n9680), .Z(n2638) );
  NAND U2795 ( .A(n2639), .B(n2638), .Z(n2727) );
  XNOR U2796 ( .A(n9872), .B(n3257), .Z(n2696) );
  NANDN U2797 ( .A(n2696), .B(n9746), .Z(n2642) );
  NANDN U2798 ( .A(n2640), .B(n9747), .Z(n2641) );
  NAND U2799 ( .A(n2642), .B(n2641), .Z(n2724) );
  IV U2800 ( .A(a[39]), .Z(n3542) );
  XNOR U2801 ( .A(n74), .B(n3542), .Z(n2699) );
  NANDN U2802 ( .A(n2699), .B(n9485), .Z(n2645) );
  NANDN U2803 ( .A(n2643), .B(n9484), .Z(n2644) );
  AND U2804 ( .A(n2645), .B(n2644), .Z(n2725) );
  XNOR U2805 ( .A(n2724), .B(n2725), .Z(n2726) );
  XOR U2806 ( .A(n2727), .B(n2726), .Z(n2703) );
  XOR U2807 ( .A(n2702), .B(n2703), .Z(n2704) );
  XNOR U2808 ( .A(n2705), .B(n2704), .Z(n2675) );
  NAND U2809 ( .A(n2647), .B(n2646), .Z(n2651) );
  NAND U2810 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U2811 ( .A(n2651), .B(n2650), .Z(n2676) );
  XOR U2812 ( .A(n2675), .B(n2676), .Z(n2678) );
  XNOR U2813 ( .A(n2677), .B(n2678), .Z(n2736) );
  NANDN U2814 ( .A(n2653), .B(n2652), .Z(n2657) );
  NAND U2815 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U2816 ( .A(n2657), .B(n2656), .Z(n2737) );
  XNOR U2817 ( .A(n2736), .B(n2737), .Z(n2738) );
  XOR U2818 ( .A(n2739), .B(n2738), .Z(n2669) );
  NANDN U2819 ( .A(n2659), .B(n2658), .Z(n2663) );
  NANDN U2820 ( .A(n2661), .B(n2660), .Z(n2662) );
  NAND U2821 ( .A(n2663), .B(n2662), .Z(n2670) );
  XNOR U2822 ( .A(n2669), .B(n2670), .Z(n2671) );
  XNOR U2823 ( .A(n2672), .B(n2671), .Z(n2742) );
  XNOR U2824 ( .A(n2742), .B(sreg[153]), .Z(n2744) );
  NAND U2825 ( .A(n2664), .B(sreg[152]), .Z(n2668) );
  OR U2826 ( .A(n2666), .B(n2665), .Z(n2667) );
  AND U2827 ( .A(n2668), .B(n2667), .Z(n2743) );
  XOR U2828 ( .A(n2744), .B(n2743), .Z(c[153]) );
  NANDN U2829 ( .A(n2670), .B(n2669), .Z(n2674) );
  NAND U2830 ( .A(n2672), .B(n2671), .Z(n2673) );
  NAND U2831 ( .A(n2674), .B(n2673), .Z(n2750) );
  NANDN U2832 ( .A(n2676), .B(n2675), .Z(n2680) );
  OR U2833 ( .A(n2678), .B(n2677), .Z(n2679) );
  NAND U2834 ( .A(n2680), .B(n2679), .Z(n2817) );
  NANDN U2835 ( .A(n2682), .B(n2681), .Z(n2686) );
  OR U2836 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U2837 ( .A(n2686), .B(n2685), .Z(n2805) );
  XNOR U2838 ( .A(n10050), .B(n2840), .Z(n2790) );
  OR U2839 ( .A(n2790), .B(n10051), .Z(n2689) );
  NANDN U2840 ( .A(n2687), .B(n10070), .Z(n2688) );
  AND U2841 ( .A(n2689), .B(n2688), .Z(n2782) );
  NAND U2842 ( .A(b[0]), .B(a[42]), .Z(n2690) );
  XNOR U2843 ( .A(b[1]), .B(n2690), .Z(n2692) );
  NAND U2844 ( .A(a[41]), .B(n72), .Z(n2691) );
  AND U2845 ( .A(n2692), .B(n2691), .Z(n2781) );
  XOR U2846 ( .A(n2782), .B(n2781), .Z(n2784) );
  NAND U2847 ( .A(a[26]), .B(b[15]), .Z(n2783) );
  XOR U2848 ( .A(n2784), .B(n2783), .Z(n2802) );
  XNOR U2849 ( .A(n9622), .B(n3464), .Z(n2793) );
  OR U2850 ( .A(n2793), .B(n9623), .Z(n2695) );
  NANDN U2851 ( .A(n2693), .B(n9680), .Z(n2694) );
  NAND U2852 ( .A(n2695), .B(n2694), .Z(n2778) );
  XNOR U2853 ( .A(n9872), .B(n3308), .Z(n2796) );
  NANDN U2854 ( .A(n2796), .B(n9746), .Z(n2698) );
  NANDN U2855 ( .A(n2696), .B(n9747), .Z(n2697) );
  NAND U2856 ( .A(n2698), .B(n2697), .Z(n2775) );
  IV U2857 ( .A(a[40]), .Z(n3647) );
  XNOR U2858 ( .A(n74), .B(n3647), .Z(n2799) );
  NANDN U2859 ( .A(n2799), .B(n9485), .Z(n2701) );
  NANDN U2860 ( .A(n2699), .B(n9484), .Z(n2700) );
  AND U2861 ( .A(n2701), .B(n2700), .Z(n2776) );
  XNOR U2862 ( .A(n2775), .B(n2776), .Z(n2777) );
  XOR U2863 ( .A(n2778), .B(n2777), .Z(n2803) );
  XOR U2864 ( .A(n2802), .B(n2803), .Z(n2804) );
  XNOR U2865 ( .A(n2805), .B(n2804), .Z(n2753) );
  NAND U2866 ( .A(n2703), .B(n2702), .Z(n2707) );
  NAND U2867 ( .A(n2705), .B(n2704), .Z(n2706) );
  NAND U2868 ( .A(n2707), .B(n2706), .Z(n2754) );
  XOR U2869 ( .A(n2753), .B(n2754), .Z(n2756) );
  XNOR U2870 ( .A(n9967), .B(n2996), .Z(n2759) );
  OR U2871 ( .A(n2759), .B(n10020), .Z(n2710) );
  NANDN U2872 ( .A(n2708), .B(n9968), .Z(n2709) );
  NAND U2873 ( .A(n2710), .B(n2709), .Z(n2772) );
  XNOR U2874 ( .A(n75), .B(n2711), .Z(n2763) );
  OR U2875 ( .A(n2763), .B(n10106), .Z(n2714) );
  NANDN U2876 ( .A(n2712), .B(n10107), .Z(n2713) );
  NAND U2877 ( .A(n2714), .B(n2713), .Z(n2769) );
  XNOR U2878 ( .A(n9984), .B(n3179), .Z(n2766) );
  NANDN U2879 ( .A(n2766), .B(n9865), .Z(n2717) );
  NANDN U2880 ( .A(n2715), .B(n9930), .Z(n2716) );
  AND U2881 ( .A(n2717), .B(n2716), .Z(n2770) );
  XNOR U2882 ( .A(n2769), .B(n2770), .Z(n2771) );
  XNOR U2883 ( .A(n2772), .B(n2771), .Z(n2808) );
  NANDN U2884 ( .A(n2719), .B(n2718), .Z(n2723) );
  NAND U2885 ( .A(n2721), .B(n2720), .Z(n2722) );
  NAND U2886 ( .A(n2723), .B(n2722), .Z(n2809) );
  XNOR U2887 ( .A(n2808), .B(n2809), .Z(n2810) );
  NANDN U2888 ( .A(n2725), .B(n2724), .Z(n2729) );
  NAND U2889 ( .A(n2727), .B(n2726), .Z(n2728) );
  AND U2890 ( .A(n2729), .B(n2728), .Z(n2811) );
  XNOR U2891 ( .A(n2810), .B(n2811), .Z(n2755) );
  XNOR U2892 ( .A(n2756), .B(n2755), .Z(n2814) );
  NANDN U2893 ( .A(n2731), .B(n2730), .Z(n2735) );
  NAND U2894 ( .A(n2733), .B(n2732), .Z(n2734) );
  NAND U2895 ( .A(n2735), .B(n2734), .Z(n2815) );
  XNOR U2896 ( .A(n2814), .B(n2815), .Z(n2816) );
  XOR U2897 ( .A(n2817), .B(n2816), .Z(n2747) );
  NANDN U2898 ( .A(n2737), .B(n2736), .Z(n2741) );
  NANDN U2899 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U2900 ( .A(n2741), .B(n2740), .Z(n2748) );
  XNOR U2901 ( .A(n2747), .B(n2748), .Z(n2749) );
  XNOR U2902 ( .A(n2750), .B(n2749), .Z(n2820) );
  XNOR U2903 ( .A(n2820), .B(sreg[154]), .Z(n2822) );
  NAND U2904 ( .A(n2742), .B(sreg[153]), .Z(n2746) );
  OR U2905 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U2906 ( .A(n2746), .B(n2745), .Z(n2821) );
  XOR U2907 ( .A(n2822), .B(n2821), .Z(c[154]) );
  NANDN U2908 ( .A(n2748), .B(n2747), .Z(n2752) );
  NAND U2909 ( .A(n2750), .B(n2749), .Z(n2751) );
  NAND U2910 ( .A(n2752), .B(n2751), .Z(n2828) );
  NANDN U2911 ( .A(n2754), .B(n2753), .Z(n2758) );
  OR U2912 ( .A(n2756), .B(n2755), .Z(n2757) );
  NAND U2913 ( .A(n2758), .B(n2757), .Z(n2895) );
  XNOR U2914 ( .A(n9967), .B(n3074), .Z(n2837) );
  OR U2915 ( .A(n2837), .B(n10020), .Z(n2761) );
  NANDN U2916 ( .A(n2759), .B(n9968), .Z(n2760) );
  NAND U2917 ( .A(n2761), .B(n2760), .Z(n2850) );
  XNOR U2918 ( .A(n75), .B(n2762), .Z(n2841) );
  OR U2919 ( .A(n2841), .B(n10106), .Z(n2765) );
  NANDN U2920 ( .A(n2763), .B(n10107), .Z(n2764) );
  NAND U2921 ( .A(n2765), .B(n2764), .Z(n2847) );
  XNOR U2922 ( .A(n9984), .B(n3257), .Z(n2844) );
  NANDN U2923 ( .A(n2844), .B(n9865), .Z(n2768) );
  NANDN U2924 ( .A(n2766), .B(n9930), .Z(n2767) );
  AND U2925 ( .A(n2768), .B(n2767), .Z(n2848) );
  XNOR U2926 ( .A(n2847), .B(n2848), .Z(n2849) );
  XNOR U2927 ( .A(n2850), .B(n2849), .Z(n2886) );
  NANDN U2928 ( .A(n2770), .B(n2769), .Z(n2774) );
  NAND U2929 ( .A(n2772), .B(n2771), .Z(n2773) );
  NAND U2930 ( .A(n2774), .B(n2773), .Z(n2887) );
  XNOR U2931 ( .A(n2886), .B(n2887), .Z(n2888) );
  NANDN U2932 ( .A(n2776), .B(n2775), .Z(n2780) );
  NAND U2933 ( .A(n2778), .B(n2777), .Z(n2779) );
  AND U2934 ( .A(n2780), .B(n2779), .Z(n2889) );
  XNOR U2935 ( .A(n2888), .B(n2889), .Z(n2833) );
  NANDN U2936 ( .A(n2782), .B(n2781), .Z(n2786) );
  OR U2937 ( .A(n2784), .B(n2783), .Z(n2785) );
  NAND U2938 ( .A(n2786), .B(n2785), .Z(n2883) );
  NAND U2939 ( .A(b[0]), .B(a[43]), .Z(n2787) );
  XNOR U2940 ( .A(b[1]), .B(n2787), .Z(n2789) );
  NAND U2941 ( .A(a[42]), .B(n72), .Z(n2788) );
  AND U2942 ( .A(n2789), .B(n2788), .Z(n2859) );
  XNOR U2943 ( .A(n10050), .B(n2918), .Z(n2868) );
  OR U2944 ( .A(n2868), .B(n10051), .Z(n2792) );
  NANDN U2945 ( .A(n2790), .B(n10070), .Z(n2791) );
  AND U2946 ( .A(n2792), .B(n2791), .Z(n2860) );
  XOR U2947 ( .A(n2859), .B(n2860), .Z(n2862) );
  NAND U2948 ( .A(a[27]), .B(b[15]), .Z(n2861) );
  XOR U2949 ( .A(n2862), .B(n2861), .Z(n2880) );
  XNOR U2950 ( .A(n9622), .B(n3542), .Z(n2871) );
  OR U2951 ( .A(n2871), .B(n9623), .Z(n2795) );
  NANDN U2952 ( .A(n2793), .B(n9680), .Z(n2794) );
  NAND U2953 ( .A(n2795), .B(n2794), .Z(n2856) );
  XNOR U2954 ( .A(n9872), .B(n3386), .Z(n2874) );
  NANDN U2955 ( .A(n2874), .B(n9746), .Z(n2798) );
  NANDN U2956 ( .A(n2796), .B(n9747), .Z(n2797) );
  NAND U2957 ( .A(n2798), .B(n2797), .Z(n2853) );
  IV U2958 ( .A(a[41]), .Z(n3725) );
  XNOR U2959 ( .A(n74), .B(n3725), .Z(n2877) );
  NANDN U2960 ( .A(n2877), .B(n9485), .Z(n2801) );
  NANDN U2961 ( .A(n2799), .B(n9484), .Z(n2800) );
  AND U2962 ( .A(n2801), .B(n2800), .Z(n2854) );
  XNOR U2963 ( .A(n2853), .B(n2854), .Z(n2855) );
  XOR U2964 ( .A(n2856), .B(n2855), .Z(n2881) );
  XOR U2965 ( .A(n2880), .B(n2881), .Z(n2882) );
  XNOR U2966 ( .A(n2883), .B(n2882), .Z(n2831) );
  NAND U2967 ( .A(n2803), .B(n2802), .Z(n2807) );
  NAND U2968 ( .A(n2805), .B(n2804), .Z(n2806) );
  NAND U2969 ( .A(n2807), .B(n2806), .Z(n2832) );
  XOR U2970 ( .A(n2831), .B(n2832), .Z(n2834) );
  XNOR U2971 ( .A(n2833), .B(n2834), .Z(n2892) );
  NANDN U2972 ( .A(n2809), .B(n2808), .Z(n2813) );
  NAND U2973 ( .A(n2811), .B(n2810), .Z(n2812) );
  NAND U2974 ( .A(n2813), .B(n2812), .Z(n2893) );
  XNOR U2975 ( .A(n2892), .B(n2893), .Z(n2894) );
  XOR U2976 ( .A(n2895), .B(n2894), .Z(n2825) );
  NANDN U2977 ( .A(n2815), .B(n2814), .Z(n2819) );
  NANDN U2978 ( .A(n2817), .B(n2816), .Z(n2818) );
  NAND U2979 ( .A(n2819), .B(n2818), .Z(n2826) );
  XNOR U2980 ( .A(n2825), .B(n2826), .Z(n2827) );
  XNOR U2981 ( .A(n2828), .B(n2827), .Z(n2898) );
  XNOR U2982 ( .A(n2898), .B(sreg[155]), .Z(n2900) );
  NAND U2983 ( .A(n2820), .B(sreg[154]), .Z(n2824) );
  OR U2984 ( .A(n2822), .B(n2821), .Z(n2823) );
  AND U2985 ( .A(n2824), .B(n2823), .Z(n2899) );
  XOR U2986 ( .A(n2900), .B(n2899), .Z(c[155]) );
  NANDN U2987 ( .A(n2826), .B(n2825), .Z(n2830) );
  NAND U2988 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U2989 ( .A(n2830), .B(n2829), .Z(n2906) );
  NANDN U2990 ( .A(n2832), .B(n2831), .Z(n2836) );
  OR U2991 ( .A(n2834), .B(n2833), .Z(n2835) );
  NAND U2992 ( .A(n2836), .B(n2835), .Z(n2973) );
  XNOR U2993 ( .A(n9967), .B(n3179), .Z(n2915) );
  OR U2994 ( .A(n2915), .B(n10020), .Z(n2839) );
  NANDN U2995 ( .A(n2837), .B(n9968), .Z(n2838) );
  NAND U2996 ( .A(n2839), .B(n2838), .Z(n2928) );
  XNOR U2997 ( .A(n75), .B(n2840), .Z(n2919) );
  OR U2998 ( .A(n2919), .B(n10106), .Z(n2843) );
  NANDN U2999 ( .A(n2841), .B(n10107), .Z(n2842) );
  NAND U3000 ( .A(n2843), .B(n2842), .Z(n2925) );
  XNOR U3001 ( .A(n9984), .B(n3308), .Z(n2922) );
  NANDN U3002 ( .A(n2922), .B(n9865), .Z(n2846) );
  NANDN U3003 ( .A(n2844), .B(n9930), .Z(n2845) );
  AND U3004 ( .A(n2846), .B(n2845), .Z(n2926) );
  XNOR U3005 ( .A(n2925), .B(n2926), .Z(n2927) );
  XNOR U3006 ( .A(n2928), .B(n2927), .Z(n2964) );
  NANDN U3007 ( .A(n2848), .B(n2847), .Z(n2852) );
  NAND U3008 ( .A(n2850), .B(n2849), .Z(n2851) );
  NAND U3009 ( .A(n2852), .B(n2851), .Z(n2965) );
  XNOR U3010 ( .A(n2964), .B(n2965), .Z(n2966) );
  NANDN U3011 ( .A(n2854), .B(n2853), .Z(n2858) );
  NAND U3012 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U3013 ( .A(n2858), .B(n2857), .Z(n2967) );
  XNOR U3014 ( .A(n2966), .B(n2967), .Z(n2911) );
  NANDN U3015 ( .A(n2860), .B(n2859), .Z(n2864) );
  OR U3016 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U3017 ( .A(n2864), .B(n2863), .Z(n2961) );
  NAND U3018 ( .A(b[0]), .B(a[44]), .Z(n2865) );
  XNOR U3019 ( .A(b[1]), .B(n2865), .Z(n2867) );
  NAND U3020 ( .A(a[43]), .B(n72), .Z(n2866) );
  AND U3021 ( .A(n2867), .B(n2866), .Z(n2937) );
  XNOR U3022 ( .A(n10050), .B(n2996), .Z(n2946) );
  OR U3023 ( .A(n2946), .B(n10051), .Z(n2870) );
  NANDN U3024 ( .A(n2868), .B(n10070), .Z(n2869) );
  AND U3025 ( .A(n2870), .B(n2869), .Z(n2938) );
  XOR U3026 ( .A(n2937), .B(n2938), .Z(n2940) );
  NAND U3027 ( .A(a[28]), .B(b[15]), .Z(n2939) );
  XOR U3028 ( .A(n2940), .B(n2939), .Z(n2958) );
  XNOR U3029 ( .A(n9622), .B(n3647), .Z(n2949) );
  OR U3030 ( .A(n2949), .B(n9623), .Z(n2873) );
  NANDN U3031 ( .A(n2871), .B(n9680), .Z(n2872) );
  NAND U3032 ( .A(n2873), .B(n2872), .Z(n2934) );
  XNOR U3033 ( .A(n9872), .B(n3464), .Z(n2952) );
  NANDN U3034 ( .A(n2952), .B(n9746), .Z(n2876) );
  NANDN U3035 ( .A(n2874), .B(n9747), .Z(n2875) );
  NAND U3036 ( .A(n2876), .B(n2875), .Z(n2931) );
  IV U3037 ( .A(a[42]), .Z(n3776) );
  XNOR U3038 ( .A(n74), .B(n3776), .Z(n2955) );
  NANDN U3039 ( .A(n2955), .B(n9485), .Z(n2879) );
  NANDN U3040 ( .A(n2877), .B(n9484), .Z(n2878) );
  AND U3041 ( .A(n2879), .B(n2878), .Z(n2932) );
  XNOR U3042 ( .A(n2931), .B(n2932), .Z(n2933) );
  XOR U3043 ( .A(n2934), .B(n2933), .Z(n2959) );
  XOR U3044 ( .A(n2958), .B(n2959), .Z(n2960) );
  XNOR U3045 ( .A(n2961), .B(n2960), .Z(n2909) );
  NAND U3046 ( .A(n2881), .B(n2880), .Z(n2885) );
  NAND U3047 ( .A(n2883), .B(n2882), .Z(n2884) );
  NAND U3048 ( .A(n2885), .B(n2884), .Z(n2910) );
  XOR U3049 ( .A(n2909), .B(n2910), .Z(n2912) );
  XNOR U3050 ( .A(n2911), .B(n2912), .Z(n2970) );
  NANDN U3051 ( .A(n2887), .B(n2886), .Z(n2891) );
  NAND U3052 ( .A(n2889), .B(n2888), .Z(n2890) );
  NAND U3053 ( .A(n2891), .B(n2890), .Z(n2971) );
  XNOR U3054 ( .A(n2970), .B(n2971), .Z(n2972) );
  XOR U3055 ( .A(n2973), .B(n2972), .Z(n2903) );
  NANDN U3056 ( .A(n2893), .B(n2892), .Z(n2897) );
  NANDN U3057 ( .A(n2895), .B(n2894), .Z(n2896) );
  NAND U3058 ( .A(n2897), .B(n2896), .Z(n2904) );
  XNOR U3059 ( .A(n2903), .B(n2904), .Z(n2905) );
  XNOR U3060 ( .A(n2906), .B(n2905), .Z(n2976) );
  XNOR U3061 ( .A(n2976), .B(sreg[156]), .Z(n2978) );
  NAND U3062 ( .A(n2898), .B(sreg[155]), .Z(n2902) );
  OR U3063 ( .A(n2900), .B(n2899), .Z(n2901) );
  AND U3064 ( .A(n2902), .B(n2901), .Z(n2977) );
  XOR U3065 ( .A(n2978), .B(n2977), .Z(c[156]) );
  NANDN U3066 ( .A(n2904), .B(n2903), .Z(n2908) );
  NAND U3067 ( .A(n2906), .B(n2905), .Z(n2907) );
  NAND U3068 ( .A(n2908), .B(n2907), .Z(n2984) );
  NANDN U3069 ( .A(n2910), .B(n2909), .Z(n2914) );
  OR U3070 ( .A(n2912), .B(n2911), .Z(n2913) );
  NAND U3071 ( .A(n2914), .B(n2913), .Z(n3051) );
  XNOR U3072 ( .A(n9967), .B(n3257), .Z(n2993) );
  OR U3073 ( .A(n2993), .B(n10020), .Z(n2917) );
  NANDN U3074 ( .A(n2915), .B(n9968), .Z(n2916) );
  NAND U3075 ( .A(n2917), .B(n2916), .Z(n3006) );
  XNOR U3076 ( .A(n75), .B(n2918), .Z(n2997) );
  OR U3077 ( .A(n2997), .B(n10106), .Z(n2921) );
  NANDN U3078 ( .A(n2919), .B(n10107), .Z(n2920) );
  NAND U3079 ( .A(n2921), .B(n2920), .Z(n3003) );
  XNOR U3080 ( .A(n9984), .B(n3386), .Z(n3000) );
  NANDN U3081 ( .A(n3000), .B(n9865), .Z(n2924) );
  NANDN U3082 ( .A(n2922), .B(n9930), .Z(n2923) );
  AND U3083 ( .A(n2924), .B(n2923), .Z(n3004) );
  XNOR U3084 ( .A(n3003), .B(n3004), .Z(n3005) );
  XNOR U3085 ( .A(n3006), .B(n3005), .Z(n3042) );
  NANDN U3086 ( .A(n2926), .B(n2925), .Z(n2930) );
  NAND U3087 ( .A(n2928), .B(n2927), .Z(n2929) );
  NAND U3088 ( .A(n2930), .B(n2929), .Z(n3043) );
  XNOR U3089 ( .A(n3042), .B(n3043), .Z(n3044) );
  NANDN U3090 ( .A(n2932), .B(n2931), .Z(n2936) );
  NAND U3091 ( .A(n2934), .B(n2933), .Z(n2935) );
  AND U3092 ( .A(n2936), .B(n2935), .Z(n3045) );
  XNOR U3093 ( .A(n3044), .B(n3045), .Z(n2989) );
  NANDN U3094 ( .A(n2938), .B(n2937), .Z(n2942) );
  OR U3095 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3096 ( .A(n2942), .B(n2941), .Z(n3039) );
  NAND U3097 ( .A(b[0]), .B(a[45]), .Z(n2943) );
  XNOR U3098 ( .A(b[1]), .B(n2943), .Z(n2945) );
  NAND U3099 ( .A(a[44]), .B(n72), .Z(n2944) );
  AND U3100 ( .A(n2945), .B(n2944), .Z(n3015) );
  XNOR U3101 ( .A(n10050), .B(n3074), .Z(n3021) );
  OR U3102 ( .A(n3021), .B(n10051), .Z(n2948) );
  NANDN U3103 ( .A(n2946), .B(n10070), .Z(n2947) );
  AND U3104 ( .A(n2948), .B(n2947), .Z(n3016) );
  XOR U3105 ( .A(n3015), .B(n3016), .Z(n3018) );
  NAND U3106 ( .A(a[29]), .B(b[15]), .Z(n3017) );
  XOR U3107 ( .A(n3018), .B(n3017), .Z(n3036) );
  XNOR U3108 ( .A(n9622), .B(n3725), .Z(n3027) );
  OR U3109 ( .A(n3027), .B(n9623), .Z(n2951) );
  NANDN U3110 ( .A(n2949), .B(n9680), .Z(n2950) );
  NAND U3111 ( .A(n2951), .B(n2950), .Z(n3012) );
  XNOR U3112 ( .A(n9872), .B(n3542), .Z(n3030) );
  NANDN U3113 ( .A(n3030), .B(n9746), .Z(n2954) );
  NANDN U3114 ( .A(n2952), .B(n9747), .Z(n2953) );
  NAND U3115 ( .A(n2954), .B(n2953), .Z(n3009) );
  IV U3116 ( .A(a[43]), .Z(n3881) );
  XNOR U3117 ( .A(n74), .B(n3881), .Z(n3033) );
  NANDN U3118 ( .A(n3033), .B(n9485), .Z(n2957) );
  NANDN U3119 ( .A(n2955), .B(n9484), .Z(n2956) );
  AND U3120 ( .A(n2957), .B(n2956), .Z(n3010) );
  XNOR U3121 ( .A(n3009), .B(n3010), .Z(n3011) );
  XOR U3122 ( .A(n3012), .B(n3011), .Z(n3037) );
  XOR U3123 ( .A(n3036), .B(n3037), .Z(n3038) );
  XNOR U3124 ( .A(n3039), .B(n3038), .Z(n2987) );
  NAND U3125 ( .A(n2959), .B(n2958), .Z(n2963) );
  NAND U3126 ( .A(n2961), .B(n2960), .Z(n2962) );
  NAND U3127 ( .A(n2963), .B(n2962), .Z(n2988) );
  XOR U3128 ( .A(n2987), .B(n2988), .Z(n2990) );
  XNOR U3129 ( .A(n2989), .B(n2990), .Z(n3048) );
  NANDN U3130 ( .A(n2965), .B(n2964), .Z(n2969) );
  NAND U3131 ( .A(n2967), .B(n2966), .Z(n2968) );
  NAND U3132 ( .A(n2969), .B(n2968), .Z(n3049) );
  XNOR U3133 ( .A(n3048), .B(n3049), .Z(n3050) );
  XOR U3134 ( .A(n3051), .B(n3050), .Z(n2981) );
  NANDN U3135 ( .A(n2971), .B(n2970), .Z(n2975) );
  NANDN U3136 ( .A(n2973), .B(n2972), .Z(n2974) );
  NAND U3137 ( .A(n2975), .B(n2974), .Z(n2982) );
  XNOR U3138 ( .A(n2981), .B(n2982), .Z(n2983) );
  XNOR U3139 ( .A(n2984), .B(n2983), .Z(n3054) );
  XNOR U3140 ( .A(n3054), .B(sreg[157]), .Z(n3056) );
  NAND U3141 ( .A(n2976), .B(sreg[156]), .Z(n2980) );
  OR U3142 ( .A(n2978), .B(n2977), .Z(n2979) );
  AND U3143 ( .A(n2980), .B(n2979), .Z(n3055) );
  XOR U3144 ( .A(n3056), .B(n3055), .Z(c[157]) );
  NANDN U3145 ( .A(n2982), .B(n2981), .Z(n2986) );
  NAND U3146 ( .A(n2984), .B(n2983), .Z(n2985) );
  NAND U3147 ( .A(n2986), .B(n2985), .Z(n3062) );
  NANDN U3148 ( .A(n2988), .B(n2987), .Z(n2992) );
  OR U3149 ( .A(n2990), .B(n2989), .Z(n2991) );
  NAND U3150 ( .A(n2992), .B(n2991), .Z(n3129) );
  XNOR U3151 ( .A(n9967), .B(n3308), .Z(n3071) );
  OR U3152 ( .A(n3071), .B(n10020), .Z(n2995) );
  NANDN U3153 ( .A(n2993), .B(n9968), .Z(n2994) );
  NAND U3154 ( .A(n2995), .B(n2994), .Z(n3084) );
  XNOR U3155 ( .A(n75), .B(n2996), .Z(n3075) );
  OR U3156 ( .A(n3075), .B(n10106), .Z(n2999) );
  NANDN U3157 ( .A(n2997), .B(n10107), .Z(n2998) );
  NAND U3158 ( .A(n2999), .B(n2998), .Z(n3081) );
  XNOR U3159 ( .A(n9984), .B(n3464), .Z(n3078) );
  NANDN U3160 ( .A(n3078), .B(n9865), .Z(n3002) );
  NANDN U3161 ( .A(n3000), .B(n9930), .Z(n3001) );
  AND U3162 ( .A(n3002), .B(n3001), .Z(n3082) );
  XNOR U3163 ( .A(n3081), .B(n3082), .Z(n3083) );
  XNOR U3164 ( .A(n3084), .B(n3083), .Z(n3120) );
  NANDN U3165 ( .A(n3004), .B(n3003), .Z(n3008) );
  NAND U3166 ( .A(n3006), .B(n3005), .Z(n3007) );
  NAND U3167 ( .A(n3008), .B(n3007), .Z(n3121) );
  XNOR U3168 ( .A(n3120), .B(n3121), .Z(n3122) );
  NANDN U3169 ( .A(n3010), .B(n3009), .Z(n3014) );
  NAND U3170 ( .A(n3012), .B(n3011), .Z(n3013) );
  AND U3171 ( .A(n3014), .B(n3013), .Z(n3123) );
  XNOR U3172 ( .A(n3122), .B(n3123), .Z(n3067) );
  NANDN U3173 ( .A(n3016), .B(n3015), .Z(n3020) );
  OR U3174 ( .A(n3018), .B(n3017), .Z(n3019) );
  NAND U3175 ( .A(n3020), .B(n3019), .Z(n3117) );
  XNOR U3176 ( .A(n10050), .B(n3179), .Z(n3102) );
  OR U3177 ( .A(n3102), .B(n10051), .Z(n3023) );
  NANDN U3178 ( .A(n3021), .B(n10070), .Z(n3022) );
  AND U3179 ( .A(n3023), .B(n3022), .Z(n3094) );
  NAND U3180 ( .A(b[0]), .B(a[46]), .Z(n3024) );
  XNOR U3181 ( .A(b[1]), .B(n3024), .Z(n3026) );
  NAND U3182 ( .A(a[45]), .B(n72), .Z(n3025) );
  AND U3183 ( .A(n3026), .B(n3025), .Z(n3093) );
  XOR U3184 ( .A(n3094), .B(n3093), .Z(n3096) );
  NAND U3185 ( .A(a[30]), .B(b[15]), .Z(n3095) );
  XOR U3186 ( .A(n3096), .B(n3095), .Z(n3114) );
  XNOR U3187 ( .A(n9622), .B(n3776), .Z(n3105) );
  OR U3188 ( .A(n3105), .B(n9623), .Z(n3029) );
  NANDN U3189 ( .A(n3027), .B(n9680), .Z(n3028) );
  NAND U3190 ( .A(n3029), .B(n3028), .Z(n3090) );
  XNOR U3191 ( .A(n9872), .B(n3647), .Z(n3108) );
  NANDN U3192 ( .A(n3108), .B(n9746), .Z(n3032) );
  NANDN U3193 ( .A(n3030), .B(n9747), .Z(n3031) );
  NAND U3194 ( .A(n3032), .B(n3031), .Z(n3087) );
  IV U3195 ( .A(a[44]), .Z(n3959) );
  XNOR U3196 ( .A(n74), .B(n3959), .Z(n3111) );
  NANDN U3197 ( .A(n3111), .B(n9485), .Z(n3035) );
  NANDN U3198 ( .A(n3033), .B(n9484), .Z(n3034) );
  AND U3199 ( .A(n3035), .B(n3034), .Z(n3088) );
  XNOR U3200 ( .A(n3087), .B(n3088), .Z(n3089) );
  XOR U3201 ( .A(n3090), .B(n3089), .Z(n3115) );
  XOR U3202 ( .A(n3114), .B(n3115), .Z(n3116) );
  XNOR U3203 ( .A(n3117), .B(n3116), .Z(n3065) );
  NAND U3204 ( .A(n3037), .B(n3036), .Z(n3041) );
  NAND U3205 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3206 ( .A(n3041), .B(n3040), .Z(n3066) );
  XOR U3207 ( .A(n3065), .B(n3066), .Z(n3068) );
  XNOR U3208 ( .A(n3067), .B(n3068), .Z(n3126) );
  NANDN U3209 ( .A(n3043), .B(n3042), .Z(n3047) );
  NAND U3210 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U3211 ( .A(n3047), .B(n3046), .Z(n3127) );
  XNOR U3212 ( .A(n3126), .B(n3127), .Z(n3128) );
  XOR U3213 ( .A(n3129), .B(n3128), .Z(n3059) );
  NANDN U3214 ( .A(n3049), .B(n3048), .Z(n3053) );
  NANDN U3215 ( .A(n3051), .B(n3050), .Z(n3052) );
  NAND U3216 ( .A(n3053), .B(n3052), .Z(n3060) );
  XNOR U3217 ( .A(n3059), .B(n3060), .Z(n3061) );
  XNOR U3218 ( .A(n3062), .B(n3061), .Z(n3132) );
  XNOR U3219 ( .A(n3132), .B(sreg[158]), .Z(n3134) );
  NAND U3220 ( .A(n3054), .B(sreg[157]), .Z(n3058) );
  OR U3221 ( .A(n3056), .B(n3055), .Z(n3057) );
  AND U3222 ( .A(n3058), .B(n3057), .Z(n3133) );
  XOR U3223 ( .A(n3134), .B(n3133), .Z(c[158]) );
  NANDN U3224 ( .A(n3060), .B(n3059), .Z(n3064) );
  NAND U3225 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3226 ( .A(n3064), .B(n3063), .Z(n3140) );
  NANDN U3227 ( .A(n3066), .B(n3065), .Z(n3070) );
  OR U3228 ( .A(n3068), .B(n3067), .Z(n3069) );
  NAND U3229 ( .A(n3070), .B(n3069), .Z(n3207) );
  XNOR U3230 ( .A(n9967), .B(n3386), .Z(n3176) );
  OR U3231 ( .A(n3176), .B(n10020), .Z(n3073) );
  NANDN U3232 ( .A(n3071), .B(n9968), .Z(n3072) );
  NAND U3233 ( .A(n3073), .B(n3072), .Z(n3189) );
  XNOR U3234 ( .A(n75), .B(n3074), .Z(n3180) );
  OR U3235 ( .A(n3180), .B(n10106), .Z(n3077) );
  NANDN U3236 ( .A(n3075), .B(n10107), .Z(n3076) );
  NAND U3237 ( .A(n3077), .B(n3076), .Z(n3186) );
  XNOR U3238 ( .A(n9984), .B(n3542), .Z(n3183) );
  NANDN U3239 ( .A(n3183), .B(n9865), .Z(n3080) );
  NANDN U3240 ( .A(n3078), .B(n9930), .Z(n3079) );
  AND U3241 ( .A(n3080), .B(n3079), .Z(n3187) );
  XNOR U3242 ( .A(n3186), .B(n3187), .Z(n3188) );
  XNOR U3243 ( .A(n3189), .B(n3188), .Z(n3198) );
  NANDN U3244 ( .A(n3082), .B(n3081), .Z(n3086) );
  NAND U3245 ( .A(n3084), .B(n3083), .Z(n3085) );
  NAND U3246 ( .A(n3086), .B(n3085), .Z(n3199) );
  XNOR U3247 ( .A(n3198), .B(n3199), .Z(n3200) );
  NANDN U3248 ( .A(n3088), .B(n3087), .Z(n3092) );
  NAND U3249 ( .A(n3090), .B(n3089), .Z(n3091) );
  AND U3250 ( .A(n3092), .B(n3091), .Z(n3201) );
  XNOR U3251 ( .A(n3200), .B(n3201), .Z(n3145) );
  NANDN U3252 ( .A(n3094), .B(n3093), .Z(n3098) );
  OR U3253 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U3254 ( .A(n3098), .B(n3097), .Z(n3173) );
  NAND U3255 ( .A(b[0]), .B(a[47]), .Z(n3099) );
  XNOR U3256 ( .A(b[1]), .B(n3099), .Z(n3101) );
  NAND U3257 ( .A(a[46]), .B(n72), .Z(n3100) );
  AND U3258 ( .A(n3101), .B(n3100), .Z(n3149) );
  XNOR U3259 ( .A(n10050), .B(n3257), .Z(n3158) );
  OR U3260 ( .A(n3158), .B(n10051), .Z(n3104) );
  NANDN U3261 ( .A(n3102), .B(n10070), .Z(n3103) );
  AND U3262 ( .A(n3104), .B(n3103), .Z(n3150) );
  XOR U3263 ( .A(n3149), .B(n3150), .Z(n3152) );
  NAND U3264 ( .A(a[31]), .B(b[15]), .Z(n3151) );
  XOR U3265 ( .A(n3152), .B(n3151), .Z(n3170) );
  XNOR U3266 ( .A(n9622), .B(n3881), .Z(n3161) );
  OR U3267 ( .A(n3161), .B(n9623), .Z(n3107) );
  NANDN U3268 ( .A(n3105), .B(n9680), .Z(n3106) );
  NAND U3269 ( .A(n3107), .B(n3106), .Z(n3195) );
  XNOR U3270 ( .A(n9872), .B(n3725), .Z(n3164) );
  NANDN U3271 ( .A(n3164), .B(n9746), .Z(n3110) );
  NANDN U3272 ( .A(n3108), .B(n9747), .Z(n3109) );
  NAND U3273 ( .A(n3110), .B(n3109), .Z(n3192) );
  IV U3274 ( .A(a[45]), .Z(n4037) );
  XNOR U3275 ( .A(n74), .B(n4037), .Z(n3167) );
  NANDN U3276 ( .A(n3167), .B(n9485), .Z(n3113) );
  NANDN U3277 ( .A(n3111), .B(n9484), .Z(n3112) );
  AND U3278 ( .A(n3113), .B(n3112), .Z(n3193) );
  XNOR U3279 ( .A(n3192), .B(n3193), .Z(n3194) );
  XOR U3280 ( .A(n3195), .B(n3194), .Z(n3171) );
  XOR U3281 ( .A(n3170), .B(n3171), .Z(n3172) );
  XNOR U3282 ( .A(n3173), .B(n3172), .Z(n3143) );
  NAND U3283 ( .A(n3115), .B(n3114), .Z(n3119) );
  NAND U3284 ( .A(n3117), .B(n3116), .Z(n3118) );
  NAND U3285 ( .A(n3119), .B(n3118), .Z(n3144) );
  XOR U3286 ( .A(n3143), .B(n3144), .Z(n3146) );
  XNOR U3287 ( .A(n3145), .B(n3146), .Z(n3204) );
  NANDN U3288 ( .A(n3121), .B(n3120), .Z(n3125) );
  NAND U3289 ( .A(n3123), .B(n3122), .Z(n3124) );
  NAND U3290 ( .A(n3125), .B(n3124), .Z(n3205) );
  XNOR U3291 ( .A(n3204), .B(n3205), .Z(n3206) );
  XOR U3292 ( .A(n3207), .B(n3206), .Z(n3137) );
  NANDN U3293 ( .A(n3127), .B(n3126), .Z(n3131) );
  NANDN U3294 ( .A(n3129), .B(n3128), .Z(n3130) );
  NAND U3295 ( .A(n3131), .B(n3130), .Z(n3138) );
  XNOR U3296 ( .A(n3137), .B(n3138), .Z(n3139) );
  XNOR U3297 ( .A(n3140), .B(n3139), .Z(n3210) );
  XNOR U3298 ( .A(n3210), .B(sreg[159]), .Z(n3212) );
  NAND U3299 ( .A(n3132), .B(sreg[158]), .Z(n3136) );
  OR U3300 ( .A(n3134), .B(n3133), .Z(n3135) );
  AND U3301 ( .A(n3136), .B(n3135), .Z(n3211) );
  XOR U3302 ( .A(n3212), .B(n3211), .Z(c[159]) );
  NANDN U3303 ( .A(n3138), .B(n3137), .Z(n3142) );
  NAND U3304 ( .A(n3140), .B(n3139), .Z(n3141) );
  NAND U3305 ( .A(n3142), .B(n3141), .Z(n3218) );
  NANDN U3306 ( .A(n3144), .B(n3143), .Z(n3148) );
  OR U3307 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3308 ( .A(n3148), .B(n3147), .Z(n3285) );
  NANDN U3309 ( .A(n3150), .B(n3149), .Z(n3154) );
  OR U3310 ( .A(n3152), .B(n3151), .Z(n3153) );
  NAND U3311 ( .A(n3154), .B(n3153), .Z(n3251) );
  NAND U3312 ( .A(b[0]), .B(a[48]), .Z(n3155) );
  XNOR U3313 ( .A(b[1]), .B(n3155), .Z(n3157) );
  NAND U3314 ( .A(a[47]), .B(n72), .Z(n3156) );
  AND U3315 ( .A(n3157), .B(n3156), .Z(n3227) );
  XNOR U3316 ( .A(n10050), .B(n3308), .Z(n3236) );
  OR U3317 ( .A(n3236), .B(n10051), .Z(n3160) );
  NANDN U3318 ( .A(n3158), .B(n10070), .Z(n3159) );
  AND U3319 ( .A(n3160), .B(n3159), .Z(n3228) );
  XOR U3320 ( .A(n3227), .B(n3228), .Z(n3230) );
  NAND U3321 ( .A(a[32]), .B(b[15]), .Z(n3229) );
  XOR U3322 ( .A(n3230), .B(n3229), .Z(n3248) );
  XNOR U3323 ( .A(n9622), .B(n3959), .Z(n3239) );
  OR U3324 ( .A(n3239), .B(n9623), .Z(n3163) );
  NANDN U3325 ( .A(n3161), .B(n9680), .Z(n3162) );
  NAND U3326 ( .A(n3163), .B(n3162), .Z(n3273) );
  XNOR U3327 ( .A(n9872), .B(n3776), .Z(n3242) );
  NANDN U3328 ( .A(n3242), .B(n9746), .Z(n3166) );
  NANDN U3329 ( .A(n3164), .B(n9747), .Z(n3165) );
  NAND U3330 ( .A(n3166), .B(n3165), .Z(n3270) );
  IV U3331 ( .A(a[46]), .Z(n4088) );
  XNOR U3332 ( .A(n74), .B(n4088), .Z(n3245) );
  NANDN U3333 ( .A(n3245), .B(n9485), .Z(n3169) );
  NANDN U3334 ( .A(n3167), .B(n9484), .Z(n3168) );
  AND U3335 ( .A(n3169), .B(n3168), .Z(n3271) );
  XNOR U3336 ( .A(n3270), .B(n3271), .Z(n3272) );
  XOR U3337 ( .A(n3273), .B(n3272), .Z(n3249) );
  XOR U3338 ( .A(n3248), .B(n3249), .Z(n3250) );
  XNOR U3339 ( .A(n3251), .B(n3250), .Z(n3221) );
  NAND U3340 ( .A(n3171), .B(n3170), .Z(n3175) );
  NAND U3341 ( .A(n3173), .B(n3172), .Z(n3174) );
  NAND U3342 ( .A(n3175), .B(n3174), .Z(n3222) );
  XOR U3343 ( .A(n3221), .B(n3222), .Z(n3224) );
  XNOR U3344 ( .A(n9967), .B(n3464), .Z(n3254) );
  OR U3345 ( .A(n3254), .B(n10020), .Z(n3178) );
  NANDN U3346 ( .A(n3176), .B(n9968), .Z(n3177) );
  NAND U3347 ( .A(n3178), .B(n3177), .Z(n3267) );
  XNOR U3348 ( .A(n75), .B(n3179), .Z(n3258) );
  OR U3349 ( .A(n3258), .B(n10106), .Z(n3182) );
  NANDN U3350 ( .A(n3180), .B(n10107), .Z(n3181) );
  NAND U3351 ( .A(n3182), .B(n3181), .Z(n3264) );
  XNOR U3352 ( .A(n9984), .B(n3647), .Z(n3261) );
  NANDN U3353 ( .A(n3261), .B(n9865), .Z(n3185) );
  NANDN U3354 ( .A(n3183), .B(n9930), .Z(n3184) );
  AND U3355 ( .A(n3185), .B(n3184), .Z(n3265) );
  XNOR U3356 ( .A(n3264), .B(n3265), .Z(n3266) );
  XNOR U3357 ( .A(n3267), .B(n3266), .Z(n3276) );
  NANDN U3358 ( .A(n3187), .B(n3186), .Z(n3191) );
  NAND U3359 ( .A(n3189), .B(n3188), .Z(n3190) );
  NAND U3360 ( .A(n3191), .B(n3190), .Z(n3277) );
  XNOR U3361 ( .A(n3276), .B(n3277), .Z(n3278) );
  NANDN U3362 ( .A(n3193), .B(n3192), .Z(n3197) );
  NAND U3363 ( .A(n3195), .B(n3194), .Z(n3196) );
  AND U3364 ( .A(n3197), .B(n3196), .Z(n3279) );
  XNOR U3365 ( .A(n3278), .B(n3279), .Z(n3223) );
  XNOR U3366 ( .A(n3224), .B(n3223), .Z(n3282) );
  NANDN U3367 ( .A(n3199), .B(n3198), .Z(n3203) );
  NAND U3368 ( .A(n3201), .B(n3200), .Z(n3202) );
  NAND U3369 ( .A(n3203), .B(n3202), .Z(n3283) );
  XNOR U3370 ( .A(n3282), .B(n3283), .Z(n3284) );
  XOR U3371 ( .A(n3285), .B(n3284), .Z(n3215) );
  NANDN U3372 ( .A(n3205), .B(n3204), .Z(n3209) );
  NANDN U3373 ( .A(n3207), .B(n3206), .Z(n3208) );
  NAND U3374 ( .A(n3209), .B(n3208), .Z(n3216) );
  XNOR U3375 ( .A(n3215), .B(n3216), .Z(n3217) );
  XNOR U3376 ( .A(n3218), .B(n3217), .Z(n3288) );
  XNOR U3377 ( .A(n3288), .B(sreg[160]), .Z(n3290) );
  NAND U3378 ( .A(n3210), .B(sreg[159]), .Z(n3214) );
  OR U3379 ( .A(n3212), .B(n3211), .Z(n3213) );
  AND U3380 ( .A(n3214), .B(n3213), .Z(n3289) );
  XOR U3381 ( .A(n3290), .B(n3289), .Z(c[160]) );
  NANDN U3382 ( .A(n3216), .B(n3215), .Z(n3220) );
  NAND U3383 ( .A(n3218), .B(n3217), .Z(n3219) );
  NAND U3384 ( .A(n3220), .B(n3219), .Z(n3296) );
  NANDN U3385 ( .A(n3222), .B(n3221), .Z(n3226) );
  OR U3386 ( .A(n3224), .B(n3223), .Z(n3225) );
  NAND U3387 ( .A(n3226), .B(n3225), .Z(n3363) );
  NANDN U3388 ( .A(n3228), .B(n3227), .Z(n3232) );
  OR U3389 ( .A(n3230), .B(n3229), .Z(n3231) );
  NAND U3390 ( .A(n3232), .B(n3231), .Z(n3351) );
  NAND U3391 ( .A(b[0]), .B(a[49]), .Z(n3233) );
  XNOR U3392 ( .A(b[1]), .B(n3233), .Z(n3235) );
  NAND U3393 ( .A(a[48]), .B(n72), .Z(n3234) );
  AND U3394 ( .A(n3235), .B(n3234), .Z(n3327) );
  XNOR U3395 ( .A(n10050), .B(n3386), .Z(n3336) );
  OR U3396 ( .A(n3336), .B(n10051), .Z(n3238) );
  NANDN U3397 ( .A(n3236), .B(n10070), .Z(n3237) );
  AND U3398 ( .A(n3238), .B(n3237), .Z(n3328) );
  XOR U3399 ( .A(n3327), .B(n3328), .Z(n3330) );
  NAND U3400 ( .A(a[33]), .B(b[15]), .Z(n3329) );
  XOR U3401 ( .A(n3330), .B(n3329), .Z(n3348) );
  XNOR U3402 ( .A(n9622), .B(n4037), .Z(n3339) );
  OR U3403 ( .A(n3339), .B(n9623), .Z(n3241) );
  NANDN U3404 ( .A(n3239), .B(n9680), .Z(n3240) );
  NAND U3405 ( .A(n3241), .B(n3240), .Z(n3324) );
  XNOR U3406 ( .A(n9872), .B(n3881), .Z(n3342) );
  NANDN U3407 ( .A(n3342), .B(n9746), .Z(n3244) );
  NANDN U3408 ( .A(n3242), .B(n9747), .Z(n3243) );
  NAND U3409 ( .A(n3244), .B(n3243), .Z(n3321) );
  IV U3410 ( .A(a[47]), .Z(n4166) );
  XNOR U3411 ( .A(n74), .B(n4166), .Z(n3345) );
  NANDN U3412 ( .A(n3345), .B(n9485), .Z(n3247) );
  NANDN U3413 ( .A(n3245), .B(n9484), .Z(n3246) );
  AND U3414 ( .A(n3247), .B(n3246), .Z(n3322) );
  XNOR U3415 ( .A(n3321), .B(n3322), .Z(n3323) );
  XOR U3416 ( .A(n3324), .B(n3323), .Z(n3349) );
  XOR U3417 ( .A(n3348), .B(n3349), .Z(n3350) );
  XNOR U3418 ( .A(n3351), .B(n3350), .Z(n3299) );
  NAND U3419 ( .A(n3249), .B(n3248), .Z(n3253) );
  NAND U3420 ( .A(n3251), .B(n3250), .Z(n3252) );
  NAND U3421 ( .A(n3253), .B(n3252), .Z(n3300) );
  XOR U3422 ( .A(n3299), .B(n3300), .Z(n3302) );
  XNOR U3423 ( .A(n9967), .B(n3542), .Z(n3305) );
  OR U3424 ( .A(n3305), .B(n10020), .Z(n3256) );
  NANDN U3425 ( .A(n3254), .B(n9968), .Z(n3255) );
  NAND U3426 ( .A(n3256), .B(n3255), .Z(n3318) );
  XNOR U3427 ( .A(n75), .B(n3257), .Z(n3309) );
  OR U3428 ( .A(n3309), .B(n10106), .Z(n3260) );
  NANDN U3429 ( .A(n3258), .B(n10107), .Z(n3259) );
  NAND U3430 ( .A(n3260), .B(n3259), .Z(n3315) );
  XNOR U3431 ( .A(n9984), .B(n3725), .Z(n3312) );
  NANDN U3432 ( .A(n3312), .B(n9865), .Z(n3263) );
  NANDN U3433 ( .A(n3261), .B(n9930), .Z(n3262) );
  AND U3434 ( .A(n3263), .B(n3262), .Z(n3316) );
  XNOR U3435 ( .A(n3315), .B(n3316), .Z(n3317) );
  XNOR U3436 ( .A(n3318), .B(n3317), .Z(n3354) );
  NANDN U3437 ( .A(n3265), .B(n3264), .Z(n3269) );
  NAND U3438 ( .A(n3267), .B(n3266), .Z(n3268) );
  NAND U3439 ( .A(n3269), .B(n3268), .Z(n3355) );
  XNOR U3440 ( .A(n3354), .B(n3355), .Z(n3356) );
  NANDN U3441 ( .A(n3271), .B(n3270), .Z(n3275) );
  NAND U3442 ( .A(n3273), .B(n3272), .Z(n3274) );
  AND U3443 ( .A(n3275), .B(n3274), .Z(n3357) );
  XNOR U3444 ( .A(n3356), .B(n3357), .Z(n3301) );
  XNOR U3445 ( .A(n3302), .B(n3301), .Z(n3360) );
  NANDN U3446 ( .A(n3277), .B(n3276), .Z(n3281) );
  NAND U3447 ( .A(n3279), .B(n3278), .Z(n3280) );
  NAND U3448 ( .A(n3281), .B(n3280), .Z(n3361) );
  XNOR U3449 ( .A(n3360), .B(n3361), .Z(n3362) );
  XOR U3450 ( .A(n3363), .B(n3362), .Z(n3293) );
  NANDN U3451 ( .A(n3283), .B(n3282), .Z(n3287) );
  NANDN U3452 ( .A(n3285), .B(n3284), .Z(n3286) );
  NAND U3453 ( .A(n3287), .B(n3286), .Z(n3294) );
  XNOR U3454 ( .A(n3293), .B(n3294), .Z(n3295) );
  XNOR U3455 ( .A(n3296), .B(n3295), .Z(n3366) );
  XNOR U3456 ( .A(n3366), .B(sreg[161]), .Z(n3368) );
  NAND U3457 ( .A(n3288), .B(sreg[160]), .Z(n3292) );
  OR U3458 ( .A(n3290), .B(n3289), .Z(n3291) );
  AND U3459 ( .A(n3292), .B(n3291), .Z(n3367) );
  XOR U3460 ( .A(n3368), .B(n3367), .Z(c[161]) );
  NANDN U3461 ( .A(n3294), .B(n3293), .Z(n3298) );
  NAND U3462 ( .A(n3296), .B(n3295), .Z(n3297) );
  NAND U3463 ( .A(n3298), .B(n3297), .Z(n3374) );
  NANDN U3464 ( .A(n3300), .B(n3299), .Z(n3304) );
  OR U3465 ( .A(n3302), .B(n3301), .Z(n3303) );
  NAND U3466 ( .A(n3304), .B(n3303), .Z(n3441) );
  XNOR U3467 ( .A(n9967), .B(n3647), .Z(n3383) );
  OR U3468 ( .A(n3383), .B(n10020), .Z(n3307) );
  NANDN U3469 ( .A(n3305), .B(n9968), .Z(n3306) );
  NAND U3470 ( .A(n3307), .B(n3306), .Z(n3396) );
  XNOR U3471 ( .A(n75), .B(n3308), .Z(n3387) );
  OR U3472 ( .A(n3387), .B(n10106), .Z(n3311) );
  NANDN U3473 ( .A(n3309), .B(n10107), .Z(n3310) );
  NAND U3474 ( .A(n3311), .B(n3310), .Z(n3393) );
  XNOR U3475 ( .A(n9984), .B(n3776), .Z(n3390) );
  NANDN U3476 ( .A(n3390), .B(n9865), .Z(n3314) );
  NANDN U3477 ( .A(n3312), .B(n9930), .Z(n3313) );
  AND U3478 ( .A(n3314), .B(n3313), .Z(n3394) );
  XNOR U3479 ( .A(n3393), .B(n3394), .Z(n3395) );
  XNOR U3480 ( .A(n3396), .B(n3395), .Z(n3432) );
  NANDN U3481 ( .A(n3316), .B(n3315), .Z(n3320) );
  NAND U3482 ( .A(n3318), .B(n3317), .Z(n3319) );
  NAND U3483 ( .A(n3320), .B(n3319), .Z(n3433) );
  XNOR U3484 ( .A(n3432), .B(n3433), .Z(n3434) );
  NANDN U3485 ( .A(n3322), .B(n3321), .Z(n3326) );
  NAND U3486 ( .A(n3324), .B(n3323), .Z(n3325) );
  AND U3487 ( .A(n3326), .B(n3325), .Z(n3435) );
  XNOR U3488 ( .A(n3434), .B(n3435), .Z(n3379) );
  NANDN U3489 ( .A(n3328), .B(n3327), .Z(n3332) );
  OR U3490 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND U3491 ( .A(n3332), .B(n3331), .Z(n3429) );
  NAND U3492 ( .A(b[0]), .B(a[50]), .Z(n3333) );
  XNOR U3493 ( .A(b[1]), .B(n3333), .Z(n3335) );
  NAND U3494 ( .A(a[49]), .B(n72), .Z(n3334) );
  AND U3495 ( .A(n3335), .B(n3334), .Z(n3405) );
  XNOR U3496 ( .A(n10050), .B(n3464), .Z(n3414) );
  OR U3497 ( .A(n3414), .B(n10051), .Z(n3338) );
  NANDN U3498 ( .A(n3336), .B(n10070), .Z(n3337) );
  AND U3499 ( .A(n3338), .B(n3337), .Z(n3406) );
  XOR U3500 ( .A(n3405), .B(n3406), .Z(n3408) );
  NAND U3501 ( .A(a[34]), .B(b[15]), .Z(n3407) );
  XOR U3502 ( .A(n3408), .B(n3407), .Z(n3426) );
  XNOR U3503 ( .A(n9622), .B(n4088), .Z(n3417) );
  OR U3504 ( .A(n3417), .B(n9623), .Z(n3341) );
  NANDN U3505 ( .A(n3339), .B(n9680), .Z(n3340) );
  NAND U3506 ( .A(n3341), .B(n3340), .Z(n3402) );
  XNOR U3507 ( .A(n9872), .B(n3959), .Z(n3420) );
  NANDN U3508 ( .A(n3420), .B(n9746), .Z(n3344) );
  NANDN U3509 ( .A(n3342), .B(n9747), .Z(n3343) );
  NAND U3510 ( .A(n3344), .B(n3343), .Z(n3399) );
  IV U3511 ( .A(a[48]), .Z(n4244) );
  XNOR U3512 ( .A(n74), .B(n4244), .Z(n3423) );
  NANDN U3513 ( .A(n3423), .B(n9485), .Z(n3347) );
  NANDN U3514 ( .A(n3345), .B(n9484), .Z(n3346) );
  AND U3515 ( .A(n3347), .B(n3346), .Z(n3400) );
  XNOR U3516 ( .A(n3399), .B(n3400), .Z(n3401) );
  XOR U3517 ( .A(n3402), .B(n3401), .Z(n3427) );
  XOR U3518 ( .A(n3426), .B(n3427), .Z(n3428) );
  XNOR U3519 ( .A(n3429), .B(n3428), .Z(n3377) );
  NAND U3520 ( .A(n3349), .B(n3348), .Z(n3353) );
  NAND U3521 ( .A(n3351), .B(n3350), .Z(n3352) );
  NAND U3522 ( .A(n3353), .B(n3352), .Z(n3378) );
  XOR U3523 ( .A(n3377), .B(n3378), .Z(n3380) );
  XNOR U3524 ( .A(n3379), .B(n3380), .Z(n3438) );
  NANDN U3525 ( .A(n3355), .B(n3354), .Z(n3359) );
  NAND U3526 ( .A(n3357), .B(n3356), .Z(n3358) );
  NAND U3527 ( .A(n3359), .B(n3358), .Z(n3439) );
  XNOR U3528 ( .A(n3438), .B(n3439), .Z(n3440) );
  XOR U3529 ( .A(n3441), .B(n3440), .Z(n3371) );
  NANDN U3530 ( .A(n3361), .B(n3360), .Z(n3365) );
  NANDN U3531 ( .A(n3363), .B(n3362), .Z(n3364) );
  NAND U3532 ( .A(n3365), .B(n3364), .Z(n3372) );
  XNOR U3533 ( .A(n3371), .B(n3372), .Z(n3373) );
  XNOR U3534 ( .A(n3374), .B(n3373), .Z(n3444) );
  XNOR U3535 ( .A(n3444), .B(sreg[162]), .Z(n3446) );
  NAND U3536 ( .A(n3366), .B(sreg[161]), .Z(n3370) );
  OR U3537 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3538 ( .A(n3370), .B(n3369), .Z(n3445) );
  XOR U3539 ( .A(n3446), .B(n3445), .Z(c[162]) );
  NANDN U3540 ( .A(n3372), .B(n3371), .Z(n3376) );
  NAND U3541 ( .A(n3374), .B(n3373), .Z(n3375) );
  NAND U3542 ( .A(n3376), .B(n3375), .Z(n3452) );
  NANDN U3543 ( .A(n3378), .B(n3377), .Z(n3382) );
  OR U3544 ( .A(n3380), .B(n3379), .Z(n3381) );
  NAND U3545 ( .A(n3382), .B(n3381), .Z(n3519) );
  XNOR U3546 ( .A(n9967), .B(n3725), .Z(n3461) );
  OR U3547 ( .A(n3461), .B(n10020), .Z(n3385) );
  NANDN U3548 ( .A(n3383), .B(n9968), .Z(n3384) );
  NAND U3549 ( .A(n3385), .B(n3384), .Z(n3474) );
  XNOR U3550 ( .A(n75), .B(n3386), .Z(n3465) );
  OR U3551 ( .A(n3465), .B(n10106), .Z(n3389) );
  NANDN U3552 ( .A(n3387), .B(n10107), .Z(n3388) );
  NAND U3553 ( .A(n3389), .B(n3388), .Z(n3471) );
  XNOR U3554 ( .A(n9984), .B(n3881), .Z(n3468) );
  NANDN U3555 ( .A(n3468), .B(n9865), .Z(n3392) );
  NANDN U3556 ( .A(n3390), .B(n9930), .Z(n3391) );
  AND U3557 ( .A(n3392), .B(n3391), .Z(n3472) );
  XNOR U3558 ( .A(n3471), .B(n3472), .Z(n3473) );
  XNOR U3559 ( .A(n3474), .B(n3473), .Z(n3510) );
  NANDN U3560 ( .A(n3394), .B(n3393), .Z(n3398) );
  NAND U3561 ( .A(n3396), .B(n3395), .Z(n3397) );
  NAND U3562 ( .A(n3398), .B(n3397), .Z(n3511) );
  XNOR U3563 ( .A(n3510), .B(n3511), .Z(n3512) );
  NANDN U3564 ( .A(n3400), .B(n3399), .Z(n3404) );
  NAND U3565 ( .A(n3402), .B(n3401), .Z(n3403) );
  AND U3566 ( .A(n3404), .B(n3403), .Z(n3513) );
  XNOR U3567 ( .A(n3512), .B(n3513), .Z(n3457) );
  NANDN U3568 ( .A(n3406), .B(n3405), .Z(n3410) );
  OR U3569 ( .A(n3408), .B(n3407), .Z(n3409) );
  NAND U3570 ( .A(n3410), .B(n3409), .Z(n3507) );
  NAND U3571 ( .A(b[0]), .B(a[51]), .Z(n3411) );
  XNOR U3572 ( .A(b[1]), .B(n3411), .Z(n3413) );
  NAND U3573 ( .A(a[50]), .B(n72), .Z(n3412) );
  AND U3574 ( .A(n3413), .B(n3412), .Z(n3483) );
  XNOR U3575 ( .A(n10050), .B(n3542), .Z(n3492) );
  OR U3576 ( .A(n3492), .B(n10051), .Z(n3416) );
  NANDN U3577 ( .A(n3414), .B(n10070), .Z(n3415) );
  AND U3578 ( .A(n3416), .B(n3415), .Z(n3484) );
  XOR U3579 ( .A(n3483), .B(n3484), .Z(n3486) );
  NAND U3580 ( .A(a[35]), .B(b[15]), .Z(n3485) );
  XOR U3581 ( .A(n3486), .B(n3485), .Z(n3504) );
  XNOR U3582 ( .A(n9622), .B(n4166), .Z(n3495) );
  OR U3583 ( .A(n3495), .B(n9623), .Z(n3419) );
  NANDN U3584 ( .A(n3417), .B(n9680), .Z(n3418) );
  NAND U3585 ( .A(n3419), .B(n3418), .Z(n3480) );
  XNOR U3586 ( .A(n9872), .B(n4037), .Z(n3498) );
  NANDN U3587 ( .A(n3498), .B(n9746), .Z(n3422) );
  NANDN U3588 ( .A(n3420), .B(n9747), .Z(n3421) );
  NAND U3589 ( .A(n3422), .B(n3421), .Z(n3477) );
  IV U3590 ( .A(a[49]), .Z(n4322) );
  XNOR U3591 ( .A(n74), .B(n4322), .Z(n3501) );
  NANDN U3592 ( .A(n3501), .B(n9485), .Z(n3425) );
  NANDN U3593 ( .A(n3423), .B(n9484), .Z(n3424) );
  AND U3594 ( .A(n3425), .B(n3424), .Z(n3478) );
  XNOR U3595 ( .A(n3477), .B(n3478), .Z(n3479) );
  XOR U3596 ( .A(n3480), .B(n3479), .Z(n3505) );
  XOR U3597 ( .A(n3504), .B(n3505), .Z(n3506) );
  XNOR U3598 ( .A(n3507), .B(n3506), .Z(n3455) );
  NAND U3599 ( .A(n3427), .B(n3426), .Z(n3431) );
  NAND U3600 ( .A(n3429), .B(n3428), .Z(n3430) );
  NAND U3601 ( .A(n3431), .B(n3430), .Z(n3456) );
  XOR U3602 ( .A(n3455), .B(n3456), .Z(n3458) );
  XNOR U3603 ( .A(n3457), .B(n3458), .Z(n3516) );
  NANDN U3604 ( .A(n3433), .B(n3432), .Z(n3437) );
  NAND U3605 ( .A(n3435), .B(n3434), .Z(n3436) );
  NAND U3606 ( .A(n3437), .B(n3436), .Z(n3517) );
  XNOR U3607 ( .A(n3516), .B(n3517), .Z(n3518) );
  XOR U3608 ( .A(n3519), .B(n3518), .Z(n3449) );
  NANDN U3609 ( .A(n3439), .B(n3438), .Z(n3443) );
  NANDN U3610 ( .A(n3441), .B(n3440), .Z(n3442) );
  NAND U3611 ( .A(n3443), .B(n3442), .Z(n3450) );
  XNOR U3612 ( .A(n3449), .B(n3450), .Z(n3451) );
  XNOR U3613 ( .A(n3452), .B(n3451), .Z(n3522) );
  XNOR U3614 ( .A(n3522), .B(sreg[163]), .Z(n3524) );
  NAND U3615 ( .A(n3444), .B(sreg[162]), .Z(n3448) );
  OR U3616 ( .A(n3446), .B(n3445), .Z(n3447) );
  AND U3617 ( .A(n3448), .B(n3447), .Z(n3523) );
  XOR U3618 ( .A(n3524), .B(n3523), .Z(c[163]) );
  NANDN U3619 ( .A(n3450), .B(n3449), .Z(n3454) );
  NAND U3620 ( .A(n3452), .B(n3451), .Z(n3453) );
  NAND U3621 ( .A(n3454), .B(n3453), .Z(n3530) );
  NANDN U3622 ( .A(n3456), .B(n3455), .Z(n3460) );
  OR U3623 ( .A(n3458), .B(n3457), .Z(n3459) );
  NAND U3624 ( .A(n3460), .B(n3459), .Z(n3597) );
  XNOR U3625 ( .A(n9967), .B(n3776), .Z(n3539) );
  OR U3626 ( .A(n3539), .B(n10020), .Z(n3463) );
  NANDN U3627 ( .A(n3461), .B(n9968), .Z(n3462) );
  NAND U3628 ( .A(n3463), .B(n3462), .Z(n3552) );
  XNOR U3629 ( .A(n75), .B(n3464), .Z(n3543) );
  OR U3630 ( .A(n3543), .B(n10106), .Z(n3467) );
  NANDN U3631 ( .A(n3465), .B(n10107), .Z(n3466) );
  NAND U3632 ( .A(n3467), .B(n3466), .Z(n3549) );
  XNOR U3633 ( .A(n9984), .B(n3959), .Z(n3546) );
  NANDN U3634 ( .A(n3546), .B(n9865), .Z(n3470) );
  NANDN U3635 ( .A(n3468), .B(n9930), .Z(n3469) );
  AND U3636 ( .A(n3470), .B(n3469), .Z(n3550) );
  XNOR U3637 ( .A(n3549), .B(n3550), .Z(n3551) );
  XNOR U3638 ( .A(n3552), .B(n3551), .Z(n3588) );
  NANDN U3639 ( .A(n3472), .B(n3471), .Z(n3476) );
  NAND U3640 ( .A(n3474), .B(n3473), .Z(n3475) );
  NAND U3641 ( .A(n3476), .B(n3475), .Z(n3589) );
  XNOR U3642 ( .A(n3588), .B(n3589), .Z(n3590) );
  NANDN U3643 ( .A(n3478), .B(n3477), .Z(n3482) );
  NAND U3644 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U3645 ( .A(n3482), .B(n3481), .Z(n3591) );
  XNOR U3646 ( .A(n3590), .B(n3591), .Z(n3535) );
  NANDN U3647 ( .A(n3484), .B(n3483), .Z(n3488) );
  OR U3648 ( .A(n3486), .B(n3485), .Z(n3487) );
  NAND U3649 ( .A(n3488), .B(n3487), .Z(n3585) );
  NAND U3650 ( .A(b[0]), .B(a[52]), .Z(n3489) );
  XNOR U3651 ( .A(b[1]), .B(n3489), .Z(n3491) );
  NAND U3652 ( .A(a[51]), .B(n72), .Z(n3490) );
  AND U3653 ( .A(n3491), .B(n3490), .Z(n3561) );
  XNOR U3654 ( .A(n10050), .B(n3647), .Z(n3567) );
  OR U3655 ( .A(n3567), .B(n10051), .Z(n3494) );
  NANDN U3656 ( .A(n3492), .B(n10070), .Z(n3493) );
  AND U3657 ( .A(n3494), .B(n3493), .Z(n3562) );
  XOR U3658 ( .A(n3561), .B(n3562), .Z(n3564) );
  NAND U3659 ( .A(a[36]), .B(b[15]), .Z(n3563) );
  XOR U3660 ( .A(n3564), .B(n3563), .Z(n3582) );
  XNOR U3661 ( .A(n9622), .B(n4244), .Z(n3573) );
  OR U3662 ( .A(n3573), .B(n9623), .Z(n3497) );
  NANDN U3663 ( .A(n3495), .B(n9680), .Z(n3496) );
  NAND U3664 ( .A(n3497), .B(n3496), .Z(n3558) );
  XNOR U3665 ( .A(n9872), .B(n4088), .Z(n3576) );
  NANDN U3666 ( .A(n3576), .B(n9746), .Z(n3500) );
  NANDN U3667 ( .A(n3498), .B(n9747), .Z(n3499) );
  NAND U3668 ( .A(n3500), .B(n3499), .Z(n3555) );
  IV U3669 ( .A(a[50]), .Z(n4427) );
  XNOR U3670 ( .A(n74), .B(n4427), .Z(n3579) );
  NANDN U3671 ( .A(n3579), .B(n9485), .Z(n3503) );
  NANDN U3672 ( .A(n3501), .B(n9484), .Z(n3502) );
  AND U3673 ( .A(n3503), .B(n3502), .Z(n3556) );
  XNOR U3674 ( .A(n3555), .B(n3556), .Z(n3557) );
  XOR U3675 ( .A(n3558), .B(n3557), .Z(n3583) );
  XOR U3676 ( .A(n3582), .B(n3583), .Z(n3584) );
  XNOR U3677 ( .A(n3585), .B(n3584), .Z(n3533) );
  NAND U3678 ( .A(n3505), .B(n3504), .Z(n3509) );
  NAND U3679 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U3680 ( .A(n3509), .B(n3508), .Z(n3534) );
  XOR U3681 ( .A(n3533), .B(n3534), .Z(n3536) );
  XNOR U3682 ( .A(n3535), .B(n3536), .Z(n3594) );
  NANDN U3683 ( .A(n3511), .B(n3510), .Z(n3515) );
  NAND U3684 ( .A(n3513), .B(n3512), .Z(n3514) );
  NAND U3685 ( .A(n3515), .B(n3514), .Z(n3595) );
  XNOR U3686 ( .A(n3594), .B(n3595), .Z(n3596) );
  XOR U3687 ( .A(n3597), .B(n3596), .Z(n3527) );
  NANDN U3688 ( .A(n3517), .B(n3516), .Z(n3521) );
  NANDN U3689 ( .A(n3519), .B(n3518), .Z(n3520) );
  NAND U3690 ( .A(n3521), .B(n3520), .Z(n3528) );
  XNOR U3691 ( .A(n3527), .B(n3528), .Z(n3529) );
  XNOR U3692 ( .A(n3530), .B(n3529), .Z(n3600) );
  XNOR U3693 ( .A(n3600), .B(sreg[164]), .Z(n3602) );
  NAND U3694 ( .A(n3522), .B(sreg[163]), .Z(n3526) );
  OR U3695 ( .A(n3524), .B(n3523), .Z(n3525) );
  AND U3696 ( .A(n3526), .B(n3525), .Z(n3601) );
  XOR U3697 ( .A(n3602), .B(n3601), .Z(c[164]) );
  NANDN U3698 ( .A(n3528), .B(n3527), .Z(n3532) );
  NAND U3699 ( .A(n3530), .B(n3529), .Z(n3531) );
  NAND U3700 ( .A(n3532), .B(n3531), .Z(n3608) );
  NANDN U3701 ( .A(n3534), .B(n3533), .Z(n3538) );
  OR U3702 ( .A(n3536), .B(n3535), .Z(n3537) );
  NAND U3703 ( .A(n3538), .B(n3537), .Z(n3675) );
  XNOR U3704 ( .A(n9967), .B(n3881), .Z(n3644) );
  OR U3705 ( .A(n3644), .B(n10020), .Z(n3541) );
  NANDN U3706 ( .A(n3539), .B(n9968), .Z(n3540) );
  NAND U3707 ( .A(n3541), .B(n3540), .Z(n3657) );
  XNOR U3708 ( .A(n75), .B(n3542), .Z(n3648) );
  OR U3709 ( .A(n3648), .B(n10106), .Z(n3545) );
  NANDN U3710 ( .A(n3543), .B(n10107), .Z(n3544) );
  NAND U3711 ( .A(n3545), .B(n3544), .Z(n3654) );
  XNOR U3712 ( .A(n9984), .B(n4037), .Z(n3651) );
  NANDN U3713 ( .A(n3651), .B(n9865), .Z(n3548) );
  NANDN U3714 ( .A(n3546), .B(n9930), .Z(n3547) );
  AND U3715 ( .A(n3548), .B(n3547), .Z(n3655) );
  XNOR U3716 ( .A(n3654), .B(n3655), .Z(n3656) );
  XNOR U3717 ( .A(n3657), .B(n3656), .Z(n3666) );
  NANDN U3718 ( .A(n3550), .B(n3549), .Z(n3554) );
  NAND U3719 ( .A(n3552), .B(n3551), .Z(n3553) );
  NAND U3720 ( .A(n3554), .B(n3553), .Z(n3667) );
  XNOR U3721 ( .A(n3666), .B(n3667), .Z(n3668) );
  NANDN U3722 ( .A(n3556), .B(n3555), .Z(n3560) );
  NAND U3723 ( .A(n3558), .B(n3557), .Z(n3559) );
  AND U3724 ( .A(n3560), .B(n3559), .Z(n3669) );
  XNOR U3725 ( .A(n3668), .B(n3669), .Z(n3613) );
  NANDN U3726 ( .A(n3562), .B(n3561), .Z(n3566) );
  OR U3727 ( .A(n3564), .B(n3563), .Z(n3565) );
  NAND U3728 ( .A(n3566), .B(n3565), .Z(n3641) );
  XNOR U3729 ( .A(n10050), .B(n3725), .Z(n3626) );
  OR U3730 ( .A(n3626), .B(n10051), .Z(n3569) );
  NANDN U3731 ( .A(n3567), .B(n10070), .Z(n3568) );
  AND U3732 ( .A(n3569), .B(n3568), .Z(n3618) );
  NAND U3733 ( .A(b[0]), .B(a[53]), .Z(n3570) );
  XNOR U3734 ( .A(b[1]), .B(n3570), .Z(n3572) );
  NAND U3735 ( .A(a[52]), .B(n72), .Z(n3571) );
  AND U3736 ( .A(n3572), .B(n3571), .Z(n3617) );
  XOR U3737 ( .A(n3618), .B(n3617), .Z(n3620) );
  NAND U3738 ( .A(a[37]), .B(b[15]), .Z(n3619) );
  XOR U3739 ( .A(n3620), .B(n3619), .Z(n3638) );
  XNOR U3740 ( .A(n9622), .B(n4322), .Z(n3629) );
  OR U3741 ( .A(n3629), .B(n9623), .Z(n3575) );
  NANDN U3742 ( .A(n3573), .B(n9680), .Z(n3574) );
  NAND U3743 ( .A(n3575), .B(n3574), .Z(n3663) );
  XNOR U3744 ( .A(n9872), .B(n4166), .Z(n3632) );
  NANDN U3745 ( .A(n3632), .B(n9746), .Z(n3578) );
  NANDN U3746 ( .A(n3576), .B(n9747), .Z(n3577) );
  NAND U3747 ( .A(n3578), .B(n3577), .Z(n3660) );
  IV U3748 ( .A(a[51]), .Z(n4478) );
  XNOR U3749 ( .A(n74), .B(n4478), .Z(n3635) );
  NANDN U3750 ( .A(n3635), .B(n9485), .Z(n3581) );
  NANDN U3751 ( .A(n3579), .B(n9484), .Z(n3580) );
  AND U3752 ( .A(n3581), .B(n3580), .Z(n3661) );
  XNOR U3753 ( .A(n3660), .B(n3661), .Z(n3662) );
  XOR U3754 ( .A(n3663), .B(n3662), .Z(n3639) );
  XOR U3755 ( .A(n3638), .B(n3639), .Z(n3640) );
  XNOR U3756 ( .A(n3641), .B(n3640), .Z(n3611) );
  NAND U3757 ( .A(n3583), .B(n3582), .Z(n3587) );
  NAND U3758 ( .A(n3585), .B(n3584), .Z(n3586) );
  NAND U3759 ( .A(n3587), .B(n3586), .Z(n3612) );
  XOR U3760 ( .A(n3611), .B(n3612), .Z(n3614) );
  XNOR U3761 ( .A(n3613), .B(n3614), .Z(n3672) );
  NANDN U3762 ( .A(n3589), .B(n3588), .Z(n3593) );
  NAND U3763 ( .A(n3591), .B(n3590), .Z(n3592) );
  NAND U3764 ( .A(n3593), .B(n3592), .Z(n3673) );
  XNOR U3765 ( .A(n3672), .B(n3673), .Z(n3674) );
  XOR U3766 ( .A(n3675), .B(n3674), .Z(n3605) );
  NANDN U3767 ( .A(n3595), .B(n3594), .Z(n3599) );
  NANDN U3768 ( .A(n3597), .B(n3596), .Z(n3598) );
  NAND U3769 ( .A(n3599), .B(n3598), .Z(n3606) );
  XNOR U3770 ( .A(n3605), .B(n3606), .Z(n3607) );
  XNOR U3771 ( .A(n3608), .B(n3607), .Z(n3678) );
  XNOR U3772 ( .A(n3678), .B(sreg[165]), .Z(n3680) );
  NAND U3773 ( .A(n3600), .B(sreg[164]), .Z(n3604) );
  OR U3774 ( .A(n3602), .B(n3601), .Z(n3603) );
  AND U3775 ( .A(n3604), .B(n3603), .Z(n3679) );
  XOR U3776 ( .A(n3680), .B(n3679), .Z(c[165]) );
  NANDN U3777 ( .A(n3606), .B(n3605), .Z(n3610) );
  NAND U3778 ( .A(n3608), .B(n3607), .Z(n3609) );
  NAND U3779 ( .A(n3610), .B(n3609), .Z(n3686) );
  NANDN U3780 ( .A(n3612), .B(n3611), .Z(n3616) );
  OR U3781 ( .A(n3614), .B(n3613), .Z(n3615) );
  NAND U3782 ( .A(n3616), .B(n3615), .Z(n3753) );
  NANDN U3783 ( .A(n3618), .B(n3617), .Z(n3622) );
  OR U3784 ( .A(n3620), .B(n3619), .Z(n3621) );
  NAND U3785 ( .A(n3622), .B(n3621), .Z(n3719) );
  NAND U3786 ( .A(b[0]), .B(a[54]), .Z(n3623) );
  XNOR U3787 ( .A(b[1]), .B(n3623), .Z(n3625) );
  NAND U3788 ( .A(a[53]), .B(n72), .Z(n3624) );
  AND U3789 ( .A(n3625), .B(n3624), .Z(n3695) );
  XNOR U3790 ( .A(n10050), .B(n3776), .Z(n3701) );
  OR U3791 ( .A(n3701), .B(n10051), .Z(n3628) );
  NANDN U3792 ( .A(n3626), .B(n10070), .Z(n3627) );
  AND U3793 ( .A(n3628), .B(n3627), .Z(n3696) );
  XOR U3794 ( .A(n3695), .B(n3696), .Z(n3698) );
  NAND U3795 ( .A(a[38]), .B(b[15]), .Z(n3697) );
  XOR U3796 ( .A(n3698), .B(n3697), .Z(n3716) );
  XNOR U3797 ( .A(n9622), .B(n4427), .Z(n3707) );
  OR U3798 ( .A(n3707), .B(n9623), .Z(n3631) );
  NANDN U3799 ( .A(n3629), .B(n9680), .Z(n3630) );
  NAND U3800 ( .A(n3631), .B(n3630), .Z(n3741) );
  XNOR U3801 ( .A(n9872), .B(n4244), .Z(n3710) );
  NANDN U3802 ( .A(n3710), .B(n9746), .Z(n3634) );
  NANDN U3803 ( .A(n3632), .B(n9747), .Z(n3633) );
  NAND U3804 ( .A(n3634), .B(n3633), .Z(n3738) );
  IV U3805 ( .A(a[52]), .Z(n4556) );
  XNOR U3806 ( .A(n74), .B(n4556), .Z(n3713) );
  NANDN U3807 ( .A(n3713), .B(n9485), .Z(n3637) );
  NANDN U3808 ( .A(n3635), .B(n9484), .Z(n3636) );
  AND U3809 ( .A(n3637), .B(n3636), .Z(n3739) );
  XNOR U3810 ( .A(n3738), .B(n3739), .Z(n3740) );
  XOR U3811 ( .A(n3741), .B(n3740), .Z(n3717) );
  XOR U3812 ( .A(n3716), .B(n3717), .Z(n3718) );
  XNOR U3813 ( .A(n3719), .B(n3718), .Z(n3689) );
  NAND U3814 ( .A(n3639), .B(n3638), .Z(n3643) );
  NAND U3815 ( .A(n3641), .B(n3640), .Z(n3642) );
  NAND U3816 ( .A(n3643), .B(n3642), .Z(n3690) );
  XOR U3817 ( .A(n3689), .B(n3690), .Z(n3692) );
  XNOR U3818 ( .A(n9967), .B(n3959), .Z(n3722) );
  OR U3819 ( .A(n3722), .B(n10020), .Z(n3646) );
  NANDN U3820 ( .A(n3644), .B(n9968), .Z(n3645) );
  NAND U3821 ( .A(n3646), .B(n3645), .Z(n3735) );
  XNOR U3822 ( .A(n75), .B(n3647), .Z(n3726) );
  OR U3823 ( .A(n3726), .B(n10106), .Z(n3650) );
  NANDN U3824 ( .A(n3648), .B(n10107), .Z(n3649) );
  NAND U3825 ( .A(n3650), .B(n3649), .Z(n3732) );
  XNOR U3826 ( .A(n9984), .B(n4088), .Z(n3729) );
  NANDN U3827 ( .A(n3729), .B(n9865), .Z(n3653) );
  NANDN U3828 ( .A(n3651), .B(n9930), .Z(n3652) );
  AND U3829 ( .A(n3653), .B(n3652), .Z(n3733) );
  XNOR U3830 ( .A(n3732), .B(n3733), .Z(n3734) );
  XNOR U3831 ( .A(n3735), .B(n3734), .Z(n3744) );
  NANDN U3832 ( .A(n3655), .B(n3654), .Z(n3659) );
  NAND U3833 ( .A(n3657), .B(n3656), .Z(n3658) );
  NAND U3834 ( .A(n3659), .B(n3658), .Z(n3745) );
  XNOR U3835 ( .A(n3744), .B(n3745), .Z(n3746) );
  NANDN U3836 ( .A(n3661), .B(n3660), .Z(n3665) );
  NAND U3837 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U3838 ( .A(n3665), .B(n3664), .Z(n3747) );
  XNOR U3839 ( .A(n3746), .B(n3747), .Z(n3691) );
  XNOR U3840 ( .A(n3692), .B(n3691), .Z(n3750) );
  NANDN U3841 ( .A(n3667), .B(n3666), .Z(n3671) );
  NAND U3842 ( .A(n3669), .B(n3668), .Z(n3670) );
  NAND U3843 ( .A(n3671), .B(n3670), .Z(n3751) );
  XNOR U3844 ( .A(n3750), .B(n3751), .Z(n3752) );
  XOR U3845 ( .A(n3753), .B(n3752), .Z(n3683) );
  NANDN U3846 ( .A(n3673), .B(n3672), .Z(n3677) );
  NANDN U3847 ( .A(n3675), .B(n3674), .Z(n3676) );
  NAND U3848 ( .A(n3677), .B(n3676), .Z(n3684) );
  XNOR U3849 ( .A(n3683), .B(n3684), .Z(n3685) );
  XNOR U3850 ( .A(n3686), .B(n3685), .Z(n3756) );
  XNOR U3851 ( .A(n3756), .B(sreg[166]), .Z(n3758) );
  NAND U3852 ( .A(n3678), .B(sreg[165]), .Z(n3682) );
  OR U3853 ( .A(n3680), .B(n3679), .Z(n3681) );
  AND U3854 ( .A(n3682), .B(n3681), .Z(n3757) );
  XOR U3855 ( .A(n3758), .B(n3757), .Z(c[166]) );
  NANDN U3856 ( .A(n3684), .B(n3683), .Z(n3688) );
  NAND U3857 ( .A(n3686), .B(n3685), .Z(n3687) );
  NAND U3858 ( .A(n3688), .B(n3687), .Z(n3764) );
  NANDN U3859 ( .A(n3690), .B(n3689), .Z(n3694) );
  OR U3860 ( .A(n3692), .B(n3691), .Z(n3693) );
  NAND U3861 ( .A(n3694), .B(n3693), .Z(n3831) );
  NANDN U3862 ( .A(n3696), .B(n3695), .Z(n3700) );
  OR U3863 ( .A(n3698), .B(n3697), .Z(n3699) );
  NAND U3864 ( .A(n3700), .B(n3699), .Z(n3819) );
  XNOR U3865 ( .A(n10050), .B(n3881), .Z(n3804) );
  OR U3866 ( .A(n3804), .B(n10051), .Z(n3703) );
  NANDN U3867 ( .A(n3701), .B(n10070), .Z(n3702) );
  AND U3868 ( .A(n3703), .B(n3702), .Z(n3796) );
  NAND U3869 ( .A(b[0]), .B(a[55]), .Z(n3704) );
  XNOR U3870 ( .A(b[1]), .B(n3704), .Z(n3706) );
  NAND U3871 ( .A(a[54]), .B(n72), .Z(n3705) );
  AND U3872 ( .A(n3706), .B(n3705), .Z(n3795) );
  XOR U3873 ( .A(n3796), .B(n3795), .Z(n3798) );
  NAND U3874 ( .A(a[39]), .B(b[15]), .Z(n3797) );
  XOR U3875 ( .A(n3798), .B(n3797), .Z(n3816) );
  XNOR U3876 ( .A(n9622), .B(n4478), .Z(n3807) );
  OR U3877 ( .A(n3807), .B(n9623), .Z(n3709) );
  NANDN U3878 ( .A(n3707), .B(n9680), .Z(n3708) );
  NAND U3879 ( .A(n3709), .B(n3708), .Z(n3792) );
  XNOR U3880 ( .A(n9872), .B(n4322), .Z(n3810) );
  NANDN U3881 ( .A(n3810), .B(n9746), .Z(n3712) );
  NANDN U3882 ( .A(n3710), .B(n9747), .Z(n3711) );
  NAND U3883 ( .A(n3712), .B(n3711), .Z(n3789) );
  IV U3884 ( .A(a[53]), .Z(n4661) );
  XNOR U3885 ( .A(n74), .B(n4661), .Z(n3813) );
  NANDN U3886 ( .A(n3813), .B(n9485), .Z(n3715) );
  NANDN U3887 ( .A(n3713), .B(n9484), .Z(n3714) );
  AND U3888 ( .A(n3715), .B(n3714), .Z(n3790) );
  XNOR U3889 ( .A(n3789), .B(n3790), .Z(n3791) );
  XOR U3890 ( .A(n3792), .B(n3791), .Z(n3817) );
  XOR U3891 ( .A(n3816), .B(n3817), .Z(n3818) );
  XNOR U3892 ( .A(n3819), .B(n3818), .Z(n3767) );
  NAND U3893 ( .A(n3717), .B(n3716), .Z(n3721) );
  NAND U3894 ( .A(n3719), .B(n3718), .Z(n3720) );
  NAND U3895 ( .A(n3721), .B(n3720), .Z(n3768) );
  XOR U3896 ( .A(n3767), .B(n3768), .Z(n3770) );
  XNOR U3897 ( .A(n9967), .B(n4037), .Z(n3773) );
  OR U3898 ( .A(n3773), .B(n10020), .Z(n3724) );
  NANDN U3899 ( .A(n3722), .B(n9968), .Z(n3723) );
  NAND U3900 ( .A(n3724), .B(n3723), .Z(n3786) );
  XNOR U3901 ( .A(n75), .B(n3725), .Z(n3777) );
  OR U3902 ( .A(n3777), .B(n10106), .Z(n3728) );
  NANDN U3903 ( .A(n3726), .B(n10107), .Z(n3727) );
  NAND U3904 ( .A(n3728), .B(n3727), .Z(n3783) );
  XNOR U3905 ( .A(n9984), .B(n4166), .Z(n3780) );
  NANDN U3906 ( .A(n3780), .B(n9865), .Z(n3731) );
  NANDN U3907 ( .A(n3729), .B(n9930), .Z(n3730) );
  AND U3908 ( .A(n3731), .B(n3730), .Z(n3784) );
  XNOR U3909 ( .A(n3783), .B(n3784), .Z(n3785) );
  XNOR U3910 ( .A(n3786), .B(n3785), .Z(n3822) );
  NANDN U3911 ( .A(n3733), .B(n3732), .Z(n3737) );
  NAND U3912 ( .A(n3735), .B(n3734), .Z(n3736) );
  NAND U3913 ( .A(n3737), .B(n3736), .Z(n3823) );
  XNOR U3914 ( .A(n3822), .B(n3823), .Z(n3824) );
  NANDN U3915 ( .A(n3739), .B(n3738), .Z(n3743) );
  NAND U3916 ( .A(n3741), .B(n3740), .Z(n3742) );
  AND U3917 ( .A(n3743), .B(n3742), .Z(n3825) );
  XNOR U3918 ( .A(n3824), .B(n3825), .Z(n3769) );
  XNOR U3919 ( .A(n3770), .B(n3769), .Z(n3828) );
  NANDN U3920 ( .A(n3745), .B(n3744), .Z(n3749) );
  NAND U3921 ( .A(n3747), .B(n3746), .Z(n3748) );
  NAND U3922 ( .A(n3749), .B(n3748), .Z(n3829) );
  XNOR U3923 ( .A(n3828), .B(n3829), .Z(n3830) );
  XOR U3924 ( .A(n3831), .B(n3830), .Z(n3761) );
  NANDN U3925 ( .A(n3751), .B(n3750), .Z(n3755) );
  NANDN U3926 ( .A(n3753), .B(n3752), .Z(n3754) );
  NAND U3927 ( .A(n3755), .B(n3754), .Z(n3762) );
  XNOR U3928 ( .A(n3761), .B(n3762), .Z(n3763) );
  XNOR U3929 ( .A(n3764), .B(n3763), .Z(n3834) );
  XNOR U3930 ( .A(n3834), .B(sreg[167]), .Z(n3836) );
  NAND U3931 ( .A(n3756), .B(sreg[166]), .Z(n3760) );
  OR U3932 ( .A(n3758), .B(n3757), .Z(n3759) );
  AND U3933 ( .A(n3760), .B(n3759), .Z(n3835) );
  XOR U3934 ( .A(n3836), .B(n3835), .Z(c[167]) );
  NANDN U3935 ( .A(n3762), .B(n3761), .Z(n3766) );
  NAND U3936 ( .A(n3764), .B(n3763), .Z(n3765) );
  NAND U3937 ( .A(n3766), .B(n3765), .Z(n3842) );
  NANDN U3938 ( .A(n3768), .B(n3767), .Z(n3772) );
  OR U3939 ( .A(n3770), .B(n3769), .Z(n3771) );
  NAND U3940 ( .A(n3772), .B(n3771), .Z(n3909) );
  XNOR U3941 ( .A(n9967), .B(n4088), .Z(n3878) );
  OR U3942 ( .A(n3878), .B(n10020), .Z(n3775) );
  NANDN U3943 ( .A(n3773), .B(n9968), .Z(n3774) );
  NAND U3944 ( .A(n3775), .B(n3774), .Z(n3891) );
  XNOR U3945 ( .A(n75), .B(n3776), .Z(n3882) );
  OR U3946 ( .A(n3882), .B(n10106), .Z(n3779) );
  NANDN U3947 ( .A(n3777), .B(n10107), .Z(n3778) );
  NAND U3948 ( .A(n3779), .B(n3778), .Z(n3888) );
  XNOR U3949 ( .A(n9984), .B(n4244), .Z(n3885) );
  NANDN U3950 ( .A(n3885), .B(n9865), .Z(n3782) );
  NANDN U3951 ( .A(n3780), .B(n9930), .Z(n3781) );
  AND U3952 ( .A(n3782), .B(n3781), .Z(n3889) );
  XNOR U3953 ( .A(n3888), .B(n3889), .Z(n3890) );
  XNOR U3954 ( .A(n3891), .B(n3890), .Z(n3900) );
  NANDN U3955 ( .A(n3784), .B(n3783), .Z(n3788) );
  NAND U3956 ( .A(n3786), .B(n3785), .Z(n3787) );
  NAND U3957 ( .A(n3788), .B(n3787), .Z(n3901) );
  XNOR U3958 ( .A(n3900), .B(n3901), .Z(n3902) );
  NANDN U3959 ( .A(n3790), .B(n3789), .Z(n3794) );
  NAND U3960 ( .A(n3792), .B(n3791), .Z(n3793) );
  AND U3961 ( .A(n3794), .B(n3793), .Z(n3903) );
  XNOR U3962 ( .A(n3902), .B(n3903), .Z(n3847) );
  NANDN U3963 ( .A(n3796), .B(n3795), .Z(n3800) );
  OR U3964 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U3965 ( .A(n3800), .B(n3799), .Z(n3875) );
  NAND U3966 ( .A(b[0]), .B(a[56]), .Z(n3801) );
  XNOR U3967 ( .A(b[1]), .B(n3801), .Z(n3803) );
  NAND U3968 ( .A(a[55]), .B(n72), .Z(n3802) );
  AND U3969 ( .A(n3803), .B(n3802), .Z(n3851) );
  XNOR U3970 ( .A(n10050), .B(n3959), .Z(n3860) );
  OR U3971 ( .A(n3860), .B(n10051), .Z(n3806) );
  NANDN U3972 ( .A(n3804), .B(n10070), .Z(n3805) );
  AND U3973 ( .A(n3806), .B(n3805), .Z(n3852) );
  XOR U3974 ( .A(n3851), .B(n3852), .Z(n3854) );
  NAND U3975 ( .A(a[40]), .B(b[15]), .Z(n3853) );
  XOR U3976 ( .A(n3854), .B(n3853), .Z(n3872) );
  XNOR U3977 ( .A(n9622), .B(n4556), .Z(n3863) );
  OR U3978 ( .A(n3863), .B(n9623), .Z(n3809) );
  NANDN U3979 ( .A(n3807), .B(n9680), .Z(n3808) );
  NAND U3980 ( .A(n3809), .B(n3808), .Z(n3897) );
  XNOR U3981 ( .A(n9872), .B(n4427), .Z(n3866) );
  NANDN U3982 ( .A(n3866), .B(n9746), .Z(n3812) );
  NANDN U3983 ( .A(n3810), .B(n9747), .Z(n3811) );
  NAND U3984 ( .A(n3812), .B(n3811), .Z(n3894) );
  IV U3985 ( .A(a[54]), .Z(n4712) );
  XNOR U3986 ( .A(n74), .B(n4712), .Z(n3869) );
  NANDN U3987 ( .A(n3869), .B(n9485), .Z(n3815) );
  NANDN U3988 ( .A(n3813), .B(n9484), .Z(n3814) );
  AND U3989 ( .A(n3815), .B(n3814), .Z(n3895) );
  XNOR U3990 ( .A(n3894), .B(n3895), .Z(n3896) );
  XOR U3991 ( .A(n3897), .B(n3896), .Z(n3873) );
  XOR U3992 ( .A(n3872), .B(n3873), .Z(n3874) );
  XNOR U3993 ( .A(n3875), .B(n3874), .Z(n3845) );
  NAND U3994 ( .A(n3817), .B(n3816), .Z(n3821) );
  NAND U3995 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U3996 ( .A(n3821), .B(n3820), .Z(n3846) );
  XOR U3997 ( .A(n3845), .B(n3846), .Z(n3848) );
  XNOR U3998 ( .A(n3847), .B(n3848), .Z(n3906) );
  NANDN U3999 ( .A(n3823), .B(n3822), .Z(n3827) );
  NAND U4000 ( .A(n3825), .B(n3824), .Z(n3826) );
  NAND U4001 ( .A(n3827), .B(n3826), .Z(n3907) );
  XNOR U4002 ( .A(n3906), .B(n3907), .Z(n3908) );
  XOR U4003 ( .A(n3909), .B(n3908), .Z(n3839) );
  NANDN U4004 ( .A(n3829), .B(n3828), .Z(n3833) );
  NANDN U4005 ( .A(n3831), .B(n3830), .Z(n3832) );
  NAND U4006 ( .A(n3833), .B(n3832), .Z(n3840) );
  XNOR U4007 ( .A(n3839), .B(n3840), .Z(n3841) );
  XNOR U4008 ( .A(n3842), .B(n3841), .Z(n3912) );
  XNOR U4009 ( .A(n3912), .B(sreg[168]), .Z(n3914) );
  NAND U4010 ( .A(n3834), .B(sreg[167]), .Z(n3838) );
  OR U4011 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U4012 ( .A(n3838), .B(n3837), .Z(n3913) );
  XOR U4013 ( .A(n3914), .B(n3913), .Z(c[168]) );
  NANDN U4014 ( .A(n3840), .B(n3839), .Z(n3844) );
  NAND U4015 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4016 ( .A(n3844), .B(n3843), .Z(n3920) );
  NANDN U4017 ( .A(n3846), .B(n3845), .Z(n3850) );
  OR U4018 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U4019 ( .A(n3850), .B(n3849), .Z(n3987) );
  NANDN U4020 ( .A(n3852), .B(n3851), .Z(n3856) );
  OR U4021 ( .A(n3854), .B(n3853), .Z(n3855) );
  NAND U4022 ( .A(n3856), .B(n3855), .Z(n3953) );
  NAND U4023 ( .A(b[0]), .B(a[57]), .Z(n3857) );
  XNOR U4024 ( .A(b[1]), .B(n3857), .Z(n3859) );
  NAND U4025 ( .A(a[56]), .B(n72), .Z(n3858) );
  AND U4026 ( .A(n3859), .B(n3858), .Z(n3929) );
  XNOR U4027 ( .A(n10050), .B(n4037), .Z(n3935) );
  OR U4028 ( .A(n3935), .B(n10051), .Z(n3862) );
  NANDN U4029 ( .A(n3860), .B(n10070), .Z(n3861) );
  AND U4030 ( .A(n3862), .B(n3861), .Z(n3930) );
  XOR U4031 ( .A(n3929), .B(n3930), .Z(n3932) );
  NAND U4032 ( .A(a[41]), .B(b[15]), .Z(n3931) );
  XOR U4033 ( .A(n3932), .B(n3931), .Z(n3950) );
  XNOR U4034 ( .A(n9622), .B(n4661), .Z(n3941) );
  OR U4035 ( .A(n3941), .B(n9623), .Z(n3865) );
  NANDN U4036 ( .A(n3863), .B(n9680), .Z(n3864) );
  NAND U4037 ( .A(n3865), .B(n3864), .Z(n3975) );
  XNOR U4038 ( .A(n9872), .B(n4478), .Z(n3944) );
  NANDN U4039 ( .A(n3944), .B(n9746), .Z(n3868) );
  NANDN U4040 ( .A(n3866), .B(n9747), .Z(n3867) );
  NAND U4041 ( .A(n3868), .B(n3867), .Z(n3972) );
  IV U4042 ( .A(a[55]), .Z(n4790) );
  XNOR U4043 ( .A(n74), .B(n4790), .Z(n3947) );
  NANDN U4044 ( .A(n3947), .B(n9485), .Z(n3871) );
  NANDN U4045 ( .A(n3869), .B(n9484), .Z(n3870) );
  AND U4046 ( .A(n3871), .B(n3870), .Z(n3973) );
  XNOR U4047 ( .A(n3972), .B(n3973), .Z(n3974) );
  XOR U4048 ( .A(n3975), .B(n3974), .Z(n3951) );
  XOR U4049 ( .A(n3950), .B(n3951), .Z(n3952) );
  XNOR U4050 ( .A(n3953), .B(n3952), .Z(n3923) );
  NAND U4051 ( .A(n3873), .B(n3872), .Z(n3877) );
  NAND U4052 ( .A(n3875), .B(n3874), .Z(n3876) );
  NAND U4053 ( .A(n3877), .B(n3876), .Z(n3924) );
  XOR U4054 ( .A(n3923), .B(n3924), .Z(n3926) );
  XNOR U4055 ( .A(n9967), .B(n4166), .Z(n3956) );
  OR U4056 ( .A(n3956), .B(n10020), .Z(n3880) );
  NANDN U4057 ( .A(n3878), .B(n9968), .Z(n3879) );
  NAND U4058 ( .A(n3880), .B(n3879), .Z(n3969) );
  XNOR U4059 ( .A(n75), .B(n3881), .Z(n3960) );
  OR U4060 ( .A(n3960), .B(n10106), .Z(n3884) );
  NANDN U4061 ( .A(n3882), .B(n10107), .Z(n3883) );
  NAND U4062 ( .A(n3884), .B(n3883), .Z(n3966) );
  XNOR U4063 ( .A(n9984), .B(n4322), .Z(n3963) );
  NANDN U4064 ( .A(n3963), .B(n9865), .Z(n3887) );
  NANDN U4065 ( .A(n3885), .B(n9930), .Z(n3886) );
  AND U4066 ( .A(n3887), .B(n3886), .Z(n3967) );
  XNOR U4067 ( .A(n3966), .B(n3967), .Z(n3968) );
  XNOR U4068 ( .A(n3969), .B(n3968), .Z(n3978) );
  NANDN U4069 ( .A(n3889), .B(n3888), .Z(n3893) );
  NAND U4070 ( .A(n3891), .B(n3890), .Z(n3892) );
  NAND U4071 ( .A(n3893), .B(n3892), .Z(n3979) );
  XNOR U4072 ( .A(n3978), .B(n3979), .Z(n3980) );
  NANDN U4073 ( .A(n3895), .B(n3894), .Z(n3899) );
  NAND U4074 ( .A(n3897), .B(n3896), .Z(n3898) );
  AND U4075 ( .A(n3899), .B(n3898), .Z(n3981) );
  XNOR U4076 ( .A(n3980), .B(n3981), .Z(n3925) );
  XNOR U4077 ( .A(n3926), .B(n3925), .Z(n3984) );
  NANDN U4078 ( .A(n3901), .B(n3900), .Z(n3905) );
  NAND U4079 ( .A(n3903), .B(n3902), .Z(n3904) );
  NAND U4080 ( .A(n3905), .B(n3904), .Z(n3985) );
  XNOR U4081 ( .A(n3984), .B(n3985), .Z(n3986) );
  XOR U4082 ( .A(n3987), .B(n3986), .Z(n3917) );
  NANDN U4083 ( .A(n3907), .B(n3906), .Z(n3911) );
  NANDN U4084 ( .A(n3909), .B(n3908), .Z(n3910) );
  NAND U4085 ( .A(n3911), .B(n3910), .Z(n3918) );
  XNOR U4086 ( .A(n3917), .B(n3918), .Z(n3919) );
  XNOR U4087 ( .A(n3920), .B(n3919), .Z(n3990) );
  XNOR U4088 ( .A(n3990), .B(sreg[169]), .Z(n3992) );
  NAND U4089 ( .A(n3912), .B(sreg[168]), .Z(n3916) );
  OR U4090 ( .A(n3914), .B(n3913), .Z(n3915) );
  AND U4091 ( .A(n3916), .B(n3915), .Z(n3991) );
  XOR U4092 ( .A(n3992), .B(n3991), .Z(c[169]) );
  NANDN U4093 ( .A(n3918), .B(n3917), .Z(n3922) );
  NAND U4094 ( .A(n3920), .B(n3919), .Z(n3921) );
  NAND U4095 ( .A(n3922), .B(n3921), .Z(n3998) );
  NANDN U4096 ( .A(n3924), .B(n3923), .Z(n3928) );
  OR U4097 ( .A(n3926), .B(n3925), .Z(n3927) );
  NAND U4098 ( .A(n3928), .B(n3927), .Z(n4065) );
  NANDN U4099 ( .A(n3930), .B(n3929), .Z(n3934) );
  OR U4100 ( .A(n3932), .B(n3931), .Z(n3933) );
  NAND U4101 ( .A(n3934), .B(n3933), .Z(n4031) );
  XNOR U4102 ( .A(n10050), .B(n4088), .Z(n4016) );
  OR U4103 ( .A(n4016), .B(n10051), .Z(n3937) );
  NANDN U4104 ( .A(n3935), .B(n10070), .Z(n3936) );
  AND U4105 ( .A(n3937), .B(n3936), .Z(n4008) );
  NAND U4106 ( .A(b[0]), .B(a[58]), .Z(n3938) );
  XNOR U4107 ( .A(b[1]), .B(n3938), .Z(n3940) );
  NAND U4108 ( .A(a[57]), .B(n72), .Z(n3939) );
  AND U4109 ( .A(n3940), .B(n3939), .Z(n4007) );
  XOR U4110 ( .A(n4008), .B(n4007), .Z(n4010) );
  NAND U4111 ( .A(a[42]), .B(b[15]), .Z(n4009) );
  XOR U4112 ( .A(n4010), .B(n4009), .Z(n4028) );
  XNOR U4113 ( .A(n9622), .B(n4712), .Z(n4019) );
  OR U4114 ( .A(n4019), .B(n9623), .Z(n3943) );
  NANDN U4115 ( .A(n3941), .B(n9680), .Z(n3942) );
  NAND U4116 ( .A(n3943), .B(n3942), .Z(n4053) );
  XNOR U4117 ( .A(n9872), .B(n4556), .Z(n4022) );
  NANDN U4118 ( .A(n4022), .B(n9746), .Z(n3946) );
  NANDN U4119 ( .A(n3944), .B(n9747), .Z(n3945) );
  NAND U4120 ( .A(n3946), .B(n3945), .Z(n4050) );
  IV U4121 ( .A(a[56]), .Z(n4868) );
  XNOR U4122 ( .A(n74), .B(n4868), .Z(n4025) );
  NANDN U4123 ( .A(n4025), .B(n9485), .Z(n3949) );
  NANDN U4124 ( .A(n3947), .B(n9484), .Z(n3948) );
  AND U4125 ( .A(n3949), .B(n3948), .Z(n4051) );
  XNOR U4126 ( .A(n4050), .B(n4051), .Z(n4052) );
  XOR U4127 ( .A(n4053), .B(n4052), .Z(n4029) );
  XOR U4128 ( .A(n4028), .B(n4029), .Z(n4030) );
  XNOR U4129 ( .A(n4031), .B(n4030), .Z(n4001) );
  NAND U4130 ( .A(n3951), .B(n3950), .Z(n3955) );
  NAND U4131 ( .A(n3953), .B(n3952), .Z(n3954) );
  NAND U4132 ( .A(n3955), .B(n3954), .Z(n4002) );
  XOR U4133 ( .A(n4001), .B(n4002), .Z(n4004) );
  XNOR U4134 ( .A(n9967), .B(n4244), .Z(n4034) );
  OR U4135 ( .A(n4034), .B(n10020), .Z(n3958) );
  NANDN U4136 ( .A(n3956), .B(n9968), .Z(n3957) );
  NAND U4137 ( .A(n3958), .B(n3957), .Z(n4047) );
  XNOR U4138 ( .A(n75), .B(n3959), .Z(n4038) );
  OR U4139 ( .A(n4038), .B(n10106), .Z(n3962) );
  NANDN U4140 ( .A(n3960), .B(n10107), .Z(n3961) );
  NAND U4141 ( .A(n3962), .B(n3961), .Z(n4044) );
  XNOR U4142 ( .A(n9984), .B(n4427), .Z(n4041) );
  NANDN U4143 ( .A(n4041), .B(n9865), .Z(n3965) );
  NANDN U4144 ( .A(n3963), .B(n9930), .Z(n3964) );
  AND U4145 ( .A(n3965), .B(n3964), .Z(n4045) );
  XNOR U4146 ( .A(n4044), .B(n4045), .Z(n4046) );
  XNOR U4147 ( .A(n4047), .B(n4046), .Z(n4056) );
  NANDN U4148 ( .A(n3967), .B(n3966), .Z(n3971) );
  NAND U4149 ( .A(n3969), .B(n3968), .Z(n3970) );
  NAND U4150 ( .A(n3971), .B(n3970), .Z(n4057) );
  XNOR U4151 ( .A(n4056), .B(n4057), .Z(n4058) );
  NANDN U4152 ( .A(n3973), .B(n3972), .Z(n3977) );
  NAND U4153 ( .A(n3975), .B(n3974), .Z(n3976) );
  AND U4154 ( .A(n3977), .B(n3976), .Z(n4059) );
  XNOR U4155 ( .A(n4058), .B(n4059), .Z(n4003) );
  XNOR U4156 ( .A(n4004), .B(n4003), .Z(n4062) );
  NANDN U4157 ( .A(n3979), .B(n3978), .Z(n3983) );
  NAND U4158 ( .A(n3981), .B(n3980), .Z(n3982) );
  NAND U4159 ( .A(n3983), .B(n3982), .Z(n4063) );
  XNOR U4160 ( .A(n4062), .B(n4063), .Z(n4064) );
  XOR U4161 ( .A(n4065), .B(n4064), .Z(n3995) );
  NANDN U4162 ( .A(n3985), .B(n3984), .Z(n3989) );
  NANDN U4163 ( .A(n3987), .B(n3986), .Z(n3988) );
  NAND U4164 ( .A(n3989), .B(n3988), .Z(n3996) );
  XNOR U4165 ( .A(n3995), .B(n3996), .Z(n3997) );
  XNOR U4166 ( .A(n3998), .B(n3997), .Z(n4068) );
  XNOR U4167 ( .A(n4068), .B(sreg[170]), .Z(n4070) );
  NAND U4168 ( .A(n3990), .B(sreg[169]), .Z(n3994) );
  OR U4169 ( .A(n3992), .B(n3991), .Z(n3993) );
  AND U4170 ( .A(n3994), .B(n3993), .Z(n4069) );
  XOR U4171 ( .A(n4070), .B(n4069), .Z(c[170]) );
  NANDN U4172 ( .A(n3996), .B(n3995), .Z(n4000) );
  NAND U4173 ( .A(n3998), .B(n3997), .Z(n3999) );
  NAND U4174 ( .A(n4000), .B(n3999), .Z(n4076) );
  NANDN U4175 ( .A(n4002), .B(n4001), .Z(n4006) );
  OR U4176 ( .A(n4004), .B(n4003), .Z(n4005) );
  NAND U4177 ( .A(n4006), .B(n4005), .Z(n4143) );
  NANDN U4178 ( .A(n4008), .B(n4007), .Z(n4012) );
  OR U4179 ( .A(n4010), .B(n4009), .Z(n4011) );
  NAND U4180 ( .A(n4012), .B(n4011), .Z(n4131) );
  NAND U4181 ( .A(b[0]), .B(a[59]), .Z(n4013) );
  XNOR U4182 ( .A(b[1]), .B(n4013), .Z(n4015) );
  NAND U4183 ( .A(a[58]), .B(n72), .Z(n4014) );
  AND U4184 ( .A(n4015), .B(n4014), .Z(n4107) );
  XNOR U4185 ( .A(n10050), .B(n4166), .Z(n4113) );
  OR U4186 ( .A(n4113), .B(n10051), .Z(n4018) );
  NANDN U4187 ( .A(n4016), .B(n10070), .Z(n4017) );
  AND U4188 ( .A(n4018), .B(n4017), .Z(n4108) );
  XOR U4189 ( .A(n4107), .B(n4108), .Z(n4110) );
  NAND U4190 ( .A(a[43]), .B(b[15]), .Z(n4109) );
  XOR U4191 ( .A(n4110), .B(n4109), .Z(n4128) );
  XNOR U4192 ( .A(n9622), .B(n4790), .Z(n4119) );
  OR U4193 ( .A(n4119), .B(n9623), .Z(n4021) );
  NANDN U4194 ( .A(n4019), .B(n9680), .Z(n4020) );
  NAND U4195 ( .A(n4021), .B(n4020), .Z(n4104) );
  XNOR U4196 ( .A(n9872), .B(n4661), .Z(n4122) );
  NANDN U4197 ( .A(n4122), .B(n9746), .Z(n4024) );
  NANDN U4198 ( .A(n4022), .B(n9747), .Z(n4023) );
  NAND U4199 ( .A(n4024), .B(n4023), .Z(n4101) );
  IV U4200 ( .A(a[57]), .Z(n4973) );
  XNOR U4201 ( .A(n74), .B(n4973), .Z(n4125) );
  NANDN U4202 ( .A(n4125), .B(n9485), .Z(n4027) );
  NANDN U4203 ( .A(n4025), .B(n9484), .Z(n4026) );
  AND U4204 ( .A(n4027), .B(n4026), .Z(n4102) );
  XNOR U4205 ( .A(n4101), .B(n4102), .Z(n4103) );
  XOR U4206 ( .A(n4104), .B(n4103), .Z(n4129) );
  XOR U4207 ( .A(n4128), .B(n4129), .Z(n4130) );
  XNOR U4208 ( .A(n4131), .B(n4130), .Z(n4079) );
  NAND U4209 ( .A(n4029), .B(n4028), .Z(n4033) );
  NAND U4210 ( .A(n4031), .B(n4030), .Z(n4032) );
  NAND U4211 ( .A(n4033), .B(n4032), .Z(n4080) );
  XOR U4212 ( .A(n4079), .B(n4080), .Z(n4082) );
  XNOR U4213 ( .A(n9967), .B(n4322), .Z(n4085) );
  OR U4214 ( .A(n4085), .B(n10020), .Z(n4036) );
  NANDN U4215 ( .A(n4034), .B(n9968), .Z(n4035) );
  NAND U4216 ( .A(n4036), .B(n4035), .Z(n4098) );
  XNOR U4217 ( .A(n75), .B(n4037), .Z(n4089) );
  OR U4218 ( .A(n4089), .B(n10106), .Z(n4040) );
  NANDN U4219 ( .A(n4038), .B(n10107), .Z(n4039) );
  NAND U4220 ( .A(n4040), .B(n4039), .Z(n4095) );
  XNOR U4221 ( .A(n9984), .B(n4478), .Z(n4092) );
  NANDN U4222 ( .A(n4092), .B(n9865), .Z(n4043) );
  NANDN U4223 ( .A(n4041), .B(n9930), .Z(n4042) );
  AND U4224 ( .A(n4043), .B(n4042), .Z(n4096) );
  XNOR U4225 ( .A(n4095), .B(n4096), .Z(n4097) );
  XNOR U4226 ( .A(n4098), .B(n4097), .Z(n4134) );
  NANDN U4227 ( .A(n4045), .B(n4044), .Z(n4049) );
  NAND U4228 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4229 ( .A(n4049), .B(n4048), .Z(n4135) );
  XNOR U4230 ( .A(n4134), .B(n4135), .Z(n4136) );
  NANDN U4231 ( .A(n4051), .B(n4050), .Z(n4055) );
  NAND U4232 ( .A(n4053), .B(n4052), .Z(n4054) );
  AND U4233 ( .A(n4055), .B(n4054), .Z(n4137) );
  XNOR U4234 ( .A(n4136), .B(n4137), .Z(n4081) );
  XNOR U4235 ( .A(n4082), .B(n4081), .Z(n4140) );
  NANDN U4236 ( .A(n4057), .B(n4056), .Z(n4061) );
  NAND U4237 ( .A(n4059), .B(n4058), .Z(n4060) );
  NAND U4238 ( .A(n4061), .B(n4060), .Z(n4141) );
  XNOR U4239 ( .A(n4140), .B(n4141), .Z(n4142) );
  XOR U4240 ( .A(n4143), .B(n4142), .Z(n4073) );
  NANDN U4241 ( .A(n4063), .B(n4062), .Z(n4067) );
  NANDN U4242 ( .A(n4065), .B(n4064), .Z(n4066) );
  NAND U4243 ( .A(n4067), .B(n4066), .Z(n4074) );
  XNOR U4244 ( .A(n4073), .B(n4074), .Z(n4075) );
  XNOR U4245 ( .A(n4076), .B(n4075), .Z(n4146) );
  XNOR U4246 ( .A(n4146), .B(sreg[171]), .Z(n4148) );
  NAND U4247 ( .A(n4068), .B(sreg[170]), .Z(n4072) );
  OR U4248 ( .A(n4070), .B(n4069), .Z(n4071) );
  AND U4249 ( .A(n4072), .B(n4071), .Z(n4147) );
  XOR U4250 ( .A(n4148), .B(n4147), .Z(c[171]) );
  NANDN U4251 ( .A(n4074), .B(n4073), .Z(n4078) );
  NAND U4252 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U4253 ( .A(n4078), .B(n4077), .Z(n4154) );
  NANDN U4254 ( .A(n4080), .B(n4079), .Z(n4084) );
  OR U4255 ( .A(n4082), .B(n4081), .Z(n4083) );
  NAND U4256 ( .A(n4084), .B(n4083), .Z(n4221) );
  XNOR U4257 ( .A(n9967), .B(n4427), .Z(n4163) );
  OR U4258 ( .A(n4163), .B(n10020), .Z(n4087) );
  NANDN U4259 ( .A(n4085), .B(n9968), .Z(n4086) );
  NAND U4260 ( .A(n4087), .B(n4086), .Z(n4176) );
  XNOR U4261 ( .A(n75), .B(n4088), .Z(n4167) );
  OR U4262 ( .A(n4167), .B(n10106), .Z(n4091) );
  NANDN U4263 ( .A(n4089), .B(n10107), .Z(n4090) );
  NAND U4264 ( .A(n4091), .B(n4090), .Z(n4173) );
  XNOR U4265 ( .A(n9984), .B(n4556), .Z(n4170) );
  NANDN U4266 ( .A(n4170), .B(n9865), .Z(n4094) );
  NANDN U4267 ( .A(n4092), .B(n9930), .Z(n4093) );
  AND U4268 ( .A(n4094), .B(n4093), .Z(n4174) );
  XNOR U4269 ( .A(n4173), .B(n4174), .Z(n4175) );
  XNOR U4270 ( .A(n4176), .B(n4175), .Z(n4212) );
  NANDN U4271 ( .A(n4096), .B(n4095), .Z(n4100) );
  NAND U4272 ( .A(n4098), .B(n4097), .Z(n4099) );
  NAND U4273 ( .A(n4100), .B(n4099), .Z(n4213) );
  XNOR U4274 ( .A(n4212), .B(n4213), .Z(n4214) );
  NANDN U4275 ( .A(n4102), .B(n4101), .Z(n4106) );
  NAND U4276 ( .A(n4104), .B(n4103), .Z(n4105) );
  AND U4277 ( .A(n4106), .B(n4105), .Z(n4215) );
  XNOR U4278 ( .A(n4214), .B(n4215), .Z(n4159) );
  NANDN U4279 ( .A(n4108), .B(n4107), .Z(n4112) );
  OR U4280 ( .A(n4110), .B(n4109), .Z(n4111) );
  NAND U4281 ( .A(n4112), .B(n4111), .Z(n4209) );
  XNOR U4282 ( .A(n10050), .B(n4244), .Z(n4194) );
  OR U4283 ( .A(n4194), .B(n10051), .Z(n4115) );
  NANDN U4284 ( .A(n4113), .B(n10070), .Z(n4114) );
  AND U4285 ( .A(n4115), .B(n4114), .Z(n4186) );
  NAND U4286 ( .A(b[0]), .B(a[60]), .Z(n4116) );
  XNOR U4287 ( .A(b[1]), .B(n4116), .Z(n4118) );
  NAND U4288 ( .A(a[59]), .B(n72), .Z(n4117) );
  AND U4289 ( .A(n4118), .B(n4117), .Z(n4185) );
  XOR U4290 ( .A(n4186), .B(n4185), .Z(n4188) );
  NAND U4291 ( .A(a[44]), .B(b[15]), .Z(n4187) );
  XOR U4292 ( .A(n4188), .B(n4187), .Z(n4206) );
  XNOR U4293 ( .A(n9622), .B(n4868), .Z(n4197) );
  OR U4294 ( .A(n4197), .B(n9623), .Z(n4121) );
  NANDN U4295 ( .A(n4119), .B(n9680), .Z(n4120) );
  NAND U4296 ( .A(n4121), .B(n4120), .Z(n4182) );
  XNOR U4297 ( .A(n9872), .B(n4712), .Z(n4200) );
  NANDN U4298 ( .A(n4200), .B(n9746), .Z(n4124) );
  NANDN U4299 ( .A(n4122), .B(n9747), .Z(n4123) );
  NAND U4300 ( .A(n4124), .B(n4123), .Z(n4179) );
  IV U4301 ( .A(a[58]), .Z(n5051) );
  XNOR U4302 ( .A(n74), .B(n5051), .Z(n4203) );
  NANDN U4303 ( .A(n4203), .B(n9485), .Z(n4127) );
  NANDN U4304 ( .A(n4125), .B(n9484), .Z(n4126) );
  AND U4305 ( .A(n4127), .B(n4126), .Z(n4180) );
  XNOR U4306 ( .A(n4179), .B(n4180), .Z(n4181) );
  XOR U4307 ( .A(n4182), .B(n4181), .Z(n4207) );
  XOR U4308 ( .A(n4206), .B(n4207), .Z(n4208) );
  XNOR U4309 ( .A(n4209), .B(n4208), .Z(n4157) );
  NAND U4310 ( .A(n4129), .B(n4128), .Z(n4133) );
  NAND U4311 ( .A(n4131), .B(n4130), .Z(n4132) );
  NAND U4312 ( .A(n4133), .B(n4132), .Z(n4158) );
  XOR U4313 ( .A(n4157), .B(n4158), .Z(n4160) );
  XNOR U4314 ( .A(n4159), .B(n4160), .Z(n4218) );
  NANDN U4315 ( .A(n4135), .B(n4134), .Z(n4139) );
  NAND U4316 ( .A(n4137), .B(n4136), .Z(n4138) );
  NAND U4317 ( .A(n4139), .B(n4138), .Z(n4219) );
  XNOR U4318 ( .A(n4218), .B(n4219), .Z(n4220) );
  XOR U4319 ( .A(n4221), .B(n4220), .Z(n4151) );
  NANDN U4320 ( .A(n4141), .B(n4140), .Z(n4145) );
  NANDN U4321 ( .A(n4143), .B(n4142), .Z(n4144) );
  NAND U4322 ( .A(n4145), .B(n4144), .Z(n4152) );
  XNOR U4323 ( .A(n4151), .B(n4152), .Z(n4153) );
  XNOR U4324 ( .A(n4154), .B(n4153), .Z(n4224) );
  XNOR U4325 ( .A(n4224), .B(sreg[172]), .Z(n4226) );
  NAND U4326 ( .A(n4146), .B(sreg[171]), .Z(n4150) );
  OR U4327 ( .A(n4148), .B(n4147), .Z(n4149) );
  AND U4328 ( .A(n4150), .B(n4149), .Z(n4225) );
  XOR U4329 ( .A(n4226), .B(n4225), .Z(c[172]) );
  NANDN U4330 ( .A(n4152), .B(n4151), .Z(n4156) );
  NAND U4331 ( .A(n4154), .B(n4153), .Z(n4155) );
  NAND U4332 ( .A(n4156), .B(n4155), .Z(n4232) );
  NANDN U4333 ( .A(n4158), .B(n4157), .Z(n4162) );
  OR U4334 ( .A(n4160), .B(n4159), .Z(n4161) );
  NAND U4335 ( .A(n4162), .B(n4161), .Z(n4299) );
  XNOR U4336 ( .A(n9967), .B(n4478), .Z(n4241) );
  OR U4337 ( .A(n4241), .B(n10020), .Z(n4165) );
  NANDN U4338 ( .A(n4163), .B(n9968), .Z(n4164) );
  NAND U4339 ( .A(n4165), .B(n4164), .Z(n4254) );
  XNOR U4340 ( .A(n75), .B(n4166), .Z(n4245) );
  OR U4341 ( .A(n4245), .B(n10106), .Z(n4169) );
  NANDN U4342 ( .A(n4167), .B(n10107), .Z(n4168) );
  NAND U4343 ( .A(n4169), .B(n4168), .Z(n4251) );
  XNOR U4344 ( .A(n9984), .B(n4661), .Z(n4248) );
  NANDN U4345 ( .A(n4248), .B(n9865), .Z(n4172) );
  NANDN U4346 ( .A(n4170), .B(n9930), .Z(n4171) );
  AND U4347 ( .A(n4172), .B(n4171), .Z(n4252) );
  XNOR U4348 ( .A(n4251), .B(n4252), .Z(n4253) );
  XNOR U4349 ( .A(n4254), .B(n4253), .Z(n4290) );
  NANDN U4350 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U4351 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U4352 ( .A(n4178), .B(n4177), .Z(n4291) );
  XNOR U4353 ( .A(n4290), .B(n4291), .Z(n4292) );
  NANDN U4354 ( .A(n4180), .B(n4179), .Z(n4184) );
  NAND U4355 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U4356 ( .A(n4184), .B(n4183), .Z(n4293) );
  XNOR U4357 ( .A(n4292), .B(n4293), .Z(n4237) );
  NANDN U4358 ( .A(n4186), .B(n4185), .Z(n4190) );
  OR U4359 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4360 ( .A(n4190), .B(n4189), .Z(n4287) );
  NAND U4361 ( .A(b[0]), .B(a[61]), .Z(n4191) );
  XNOR U4362 ( .A(b[1]), .B(n4191), .Z(n4193) );
  NAND U4363 ( .A(a[60]), .B(n72), .Z(n4192) );
  AND U4364 ( .A(n4193), .B(n4192), .Z(n4263) );
  XNOR U4365 ( .A(n10050), .B(n4322), .Z(n4272) );
  OR U4366 ( .A(n4272), .B(n10051), .Z(n4196) );
  NANDN U4367 ( .A(n4194), .B(n10070), .Z(n4195) );
  AND U4368 ( .A(n4196), .B(n4195), .Z(n4264) );
  XOR U4369 ( .A(n4263), .B(n4264), .Z(n4266) );
  NAND U4370 ( .A(a[45]), .B(b[15]), .Z(n4265) );
  XOR U4371 ( .A(n4266), .B(n4265), .Z(n4284) );
  XNOR U4372 ( .A(n9622), .B(n4973), .Z(n4275) );
  OR U4373 ( .A(n4275), .B(n9623), .Z(n4199) );
  NANDN U4374 ( .A(n4197), .B(n9680), .Z(n4198) );
  NAND U4375 ( .A(n4199), .B(n4198), .Z(n4260) );
  XNOR U4376 ( .A(n9872), .B(n4790), .Z(n4278) );
  NANDN U4377 ( .A(n4278), .B(n9746), .Z(n4202) );
  NANDN U4378 ( .A(n4200), .B(n9747), .Z(n4201) );
  NAND U4379 ( .A(n4202), .B(n4201), .Z(n4257) );
  IV U4380 ( .A(a[59]), .Z(n5102) );
  XNOR U4381 ( .A(n74), .B(n5102), .Z(n4281) );
  NANDN U4382 ( .A(n4281), .B(n9485), .Z(n4205) );
  NANDN U4383 ( .A(n4203), .B(n9484), .Z(n4204) );
  AND U4384 ( .A(n4205), .B(n4204), .Z(n4258) );
  XNOR U4385 ( .A(n4257), .B(n4258), .Z(n4259) );
  XOR U4386 ( .A(n4260), .B(n4259), .Z(n4285) );
  XOR U4387 ( .A(n4284), .B(n4285), .Z(n4286) );
  XNOR U4388 ( .A(n4287), .B(n4286), .Z(n4235) );
  NAND U4389 ( .A(n4207), .B(n4206), .Z(n4211) );
  NAND U4390 ( .A(n4209), .B(n4208), .Z(n4210) );
  NAND U4391 ( .A(n4211), .B(n4210), .Z(n4236) );
  XOR U4392 ( .A(n4235), .B(n4236), .Z(n4238) );
  XNOR U4393 ( .A(n4237), .B(n4238), .Z(n4296) );
  NANDN U4394 ( .A(n4213), .B(n4212), .Z(n4217) );
  NAND U4395 ( .A(n4215), .B(n4214), .Z(n4216) );
  NAND U4396 ( .A(n4217), .B(n4216), .Z(n4297) );
  XNOR U4397 ( .A(n4296), .B(n4297), .Z(n4298) );
  XOR U4398 ( .A(n4299), .B(n4298), .Z(n4229) );
  NANDN U4399 ( .A(n4219), .B(n4218), .Z(n4223) );
  NANDN U4400 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U4401 ( .A(n4223), .B(n4222), .Z(n4230) );
  XNOR U4402 ( .A(n4229), .B(n4230), .Z(n4231) );
  XNOR U4403 ( .A(n4232), .B(n4231), .Z(n4302) );
  XNOR U4404 ( .A(n4302), .B(sreg[173]), .Z(n4304) );
  NAND U4405 ( .A(n4224), .B(sreg[172]), .Z(n4228) );
  OR U4406 ( .A(n4226), .B(n4225), .Z(n4227) );
  AND U4407 ( .A(n4228), .B(n4227), .Z(n4303) );
  XOR U4408 ( .A(n4304), .B(n4303), .Z(c[173]) );
  NANDN U4409 ( .A(n4230), .B(n4229), .Z(n4234) );
  NAND U4410 ( .A(n4232), .B(n4231), .Z(n4233) );
  NAND U4411 ( .A(n4234), .B(n4233), .Z(n4310) );
  NANDN U4412 ( .A(n4236), .B(n4235), .Z(n4240) );
  OR U4413 ( .A(n4238), .B(n4237), .Z(n4239) );
  NAND U4414 ( .A(n4240), .B(n4239), .Z(n4377) );
  XNOR U4415 ( .A(n9967), .B(n4556), .Z(n4319) );
  OR U4416 ( .A(n4319), .B(n10020), .Z(n4243) );
  NANDN U4417 ( .A(n4241), .B(n9968), .Z(n4242) );
  NAND U4418 ( .A(n4243), .B(n4242), .Z(n4332) );
  XNOR U4419 ( .A(n75), .B(n4244), .Z(n4323) );
  OR U4420 ( .A(n4323), .B(n10106), .Z(n4247) );
  NANDN U4421 ( .A(n4245), .B(n10107), .Z(n4246) );
  NAND U4422 ( .A(n4247), .B(n4246), .Z(n4329) );
  XNOR U4423 ( .A(n9984), .B(n4712), .Z(n4326) );
  NANDN U4424 ( .A(n4326), .B(n9865), .Z(n4250) );
  NANDN U4425 ( .A(n4248), .B(n9930), .Z(n4249) );
  AND U4426 ( .A(n4250), .B(n4249), .Z(n4330) );
  XNOR U4427 ( .A(n4329), .B(n4330), .Z(n4331) );
  XNOR U4428 ( .A(n4332), .B(n4331), .Z(n4368) );
  NANDN U4429 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U4430 ( .A(n4254), .B(n4253), .Z(n4255) );
  NAND U4431 ( .A(n4256), .B(n4255), .Z(n4369) );
  XNOR U4432 ( .A(n4368), .B(n4369), .Z(n4370) );
  NANDN U4433 ( .A(n4258), .B(n4257), .Z(n4262) );
  NAND U4434 ( .A(n4260), .B(n4259), .Z(n4261) );
  AND U4435 ( .A(n4262), .B(n4261), .Z(n4371) );
  XNOR U4436 ( .A(n4370), .B(n4371), .Z(n4315) );
  NANDN U4437 ( .A(n4264), .B(n4263), .Z(n4268) );
  OR U4438 ( .A(n4266), .B(n4265), .Z(n4267) );
  NAND U4439 ( .A(n4268), .B(n4267), .Z(n4365) );
  NAND U4440 ( .A(b[0]), .B(a[62]), .Z(n4269) );
  XNOR U4441 ( .A(b[1]), .B(n4269), .Z(n4271) );
  NAND U4442 ( .A(a[61]), .B(n72), .Z(n4270) );
  AND U4443 ( .A(n4271), .B(n4270), .Z(n4341) );
  XNOR U4444 ( .A(n10050), .B(n4427), .Z(n4350) );
  OR U4445 ( .A(n4350), .B(n10051), .Z(n4274) );
  NANDN U4446 ( .A(n4272), .B(n10070), .Z(n4273) );
  AND U4447 ( .A(n4274), .B(n4273), .Z(n4342) );
  XOR U4448 ( .A(n4341), .B(n4342), .Z(n4344) );
  NAND U4449 ( .A(a[46]), .B(b[15]), .Z(n4343) );
  XOR U4450 ( .A(n4344), .B(n4343), .Z(n4362) );
  XNOR U4451 ( .A(n9622), .B(n5051), .Z(n4353) );
  OR U4452 ( .A(n4353), .B(n9623), .Z(n4277) );
  NANDN U4453 ( .A(n4275), .B(n9680), .Z(n4276) );
  NAND U4454 ( .A(n4277), .B(n4276), .Z(n4338) );
  XNOR U4455 ( .A(n9872), .B(n4868), .Z(n4356) );
  NANDN U4456 ( .A(n4356), .B(n9746), .Z(n4280) );
  NANDN U4457 ( .A(n4278), .B(n9747), .Z(n4279) );
  NAND U4458 ( .A(n4280), .B(n4279), .Z(n4335) );
  IV U4459 ( .A(a[60]), .Z(n5180) );
  XNOR U4460 ( .A(n74), .B(n5180), .Z(n4359) );
  NANDN U4461 ( .A(n4359), .B(n9485), .Z(n4283) );
  NANDN U4462 ( .A(n4281), .B(n9484), .Z(n4282) );
  AND U4463 ( .A(n4283), .B(n4282), .Z(n4336) );
  XNOR U4464 ( .A(n4335), .B(n4336), .Z(n4337) );
  XOR U4465 ( .A(n4338), .B(n4337), .Z(n4363) );
  XOR U4466 ( .A(n4362), .B(n4363), .Z(n4364) );
  XNOR U4467 ( .A(n4365), .B(n4364), .Z(n4313) );
  NAND U4468 ( .A(n4285), .B(n4284), .Z(n4289) );
  NAND U4469 ( .A(n4287), .B(n4286), .Z(n4288) );
  NAND U4470 ( .A(n4289), .B(n4288), .Z(n4314) );
  XOR U4471 ( .A(n4313), .B(n4314), .Z(n4316) );
  XNOR U4472 ( .A(n4315), .B(n4316), .Z(n4374) );
  NANDN U4473 ( .A(n4291), .B(n4290), .Z(n4295) );
  NAND U4474 ( .A(n4293), .B(n4292), .Z(n4294) );
  NAND U4475 ( .A(n4295), .B(n4294), .Z(n4375) );
  XNOR U4476 ( .A(n4374), .B(n4375), .Z(n4376) );
  XOR U4477 ( .A(n4377), .B(n4376), .Z(n4307) );
  NANDN U4478 ( .A(n4297), .B(n4296), .Z(n4301) );
  NANDN U4479 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U4480 ( .A(n4301), .B(n4300), .Z(n4308) );
  XNOR U4481 ( .A(n4307), .B(n4308), .Z(n4309) );
  XNOR U4482 ( .A(n4310), .B(n4309), .Z(n4380) );
  XNOR U4483 ( .A(n4380), .B(sreg[174]), .Z(n4382) );
  NAND U4484 ( .A(n4302), .B(sreg[173]), .Z(n4306) );
  OR U4485 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4486 ( .A(n4306), .B(n4305), .Z(n4381) );
  XOR U4487 ( .A(n4382), .B(n4381), .Z(c[174]) );
  NANDN U4488 ( .A(n4308), .B(n4307), .Z(n4312) );
  NAND U4489 ( .A(n4310), .B(n4309), .Z(n4311) );
  NAND U4490 ( .A(n4312), .B(n4311), .Z(n4388) );
  NANDN U4491 ( .A(n4314), .B(n4313), .Z(n4318) );
  OR U4492 ( .A(n4316), .B(n4315), .Z(n4317) );
  NAND U4493 ( .A(n4318), .B(n4317), .Z(n4455) );
  XNOR U4494 ( .A(n9967), .B(n4661), .Z(n4424) );
  OR U4495 ( .A(n4424), .B(n10020), .Z(n4321) );
  NANDN U4496 ( .A(n4319), .B(n9968), .Z(n4320) );
  NAND U4497 ( .A(n4321), .B(n4320), .Z(n4437) );
  XNOR U4498 ( .A(n75), .B(n4322), .Z(n4428) );
  OR U4499 ( .A(n4428), .B(n10106), .Z(n4325) );
  NANDN U4500 ( .A(n4323), .B(n10107), .Z(n4324) );
  NAND U4501 ( .A(n4325), .B(n4324), .Z(n4434) );
  XNOR U4502 ( .A(n9984), .B(n4790), .Z(n4431) );
  NANDN U4503 ( .A(n4431), .B(n9865), .Z(n4328) );
  NANDN U4504 ( .A(n4326), .B(n9930), .Z(n4327) );
  AND U4505 ( .A(n4328), .B(n4327), .Z(n4435) );
  XNOR U4506 ( .A(n4434), .B(n4435), .Z(n4436) );
  XNOR U4507 ( .A(n4437), .B(n4436), .Z(n4446) );
  NANDN U4508 ( .A(n4330), .B(n4329), .Z(n4334) );
  NAND U4509 ( .A(n4332), .B(n4331), .Z(n4333) );
  NAND U4510 ( .A(n4334), .B(n4333), .Z(n4447) );
  XNOR U4511 ( .A(n4446), .B(n4447), .Z(n4448) );
  NANDN U4512 ( .A(n4336), .B(n4335), .Z(n4340) );
  NAND U4513 ( .A(n4338), .B(n4337), .Z(n4339) );
  AND U4514 ( .A(n4340), .B(n4339), .Z(n4449) );
  XNOR U4515 ( .A(n4448), .B(n4449), .Z(n4393) );
  NANDN U4516 ( .A(n4342), .B(n4341), .Z(n4346) );
  OR U4517 ( .A(n4344), .B(n4343), .Z(n4345) );
  NAND U4518 ( .A(n4346), .B(n4345), .Z(n4421) );
  NAND U4519 ( .A(b[0]), .B(a[63]), .Z(n4347) );
  XNOR U4520 ( .A(b[1]), .B(n4347), .Z(n4349) );
  NAND U4521 ( .A(a[62]), .B(n72), .Z(n4348) );
  AND U4522 ( .A(n4349), .B(n4348), .Z(n4397) );
  XNOR U4523 ( .A(n10050), .B(n4478), .Z(n4406) );
  OR U4524 ( .A(n4406), .B(n10051), .Z(n4352) );
  NANDN U4525 ( .A(n4350), .B(n10070), .Z(n4351) );
  AND U4526 ( .A(n4352), .B(n4351), .Z(n4398) );
  XOR U4527 ( .A(n4397), .B(n4398), .Z(n4400) );
  NAND U4528 ( .A(a[47]), .B(b[15]), .Z(n4399) );
  XOR U4529 ( .A(n4400), .B(n4399), .Z(n4418) );
  XNOR U4530 ( .A(n9622), .B(n5102), .Z(n4409) );
  OR U4531 ( .A(n4409), .B(n9623), .Z(n4355) );
  NANDN U4532 ( .A(n4353), .B(n9680), .Z(n4354) );
  NAND U4533 ( .A(n4355), .B(n4354), .Z(n4443) );
  XNOR U4534 ( .A(n9872), .B(n4973), .Z(n4412) );
  NANDN U4535 ( .A(n4412), .B(n9746), .Z(n4358) );
  NANDN U4536 ( .A(n4356), .B(n9747), .Z(n4357) );
  NAND U4537 ( .A(n4358), .B(n4357), .Z(n4440) );
  IV U4538 ( .A(a[61]), .Z(n5258) );
  XNOR U4539 ( .A(n74), .B(n5258), .Z(n4415) );
  NANDN U4540 ( .A(n4415), .B(n9485), .Z(n4361) );
  NANDN U4541 ( .A(n4359), .B(n9484), .Z(n4360) );
  AND U4542 ( .A(n4361), .B(n4360), .Z(n4441) );
  XNOR U4543 ( .A(n4440), .B(n4441), .Z(n4442) );
  XOR U4544 ( .A(n4443), .B(n4442), .Z(n4419) );
  XOR U4545 ( .A(n4418), .B(n4419), .Z(n4420) );
  XNOR U4546 ( .A(n4421), .B(n4420), .Z(n4391) );
  NAND U4547 ( .A(n4363), .B(n4362), .Z(n4367) );
  NAND U4548 ( .A(n4365), .B(n4364), .Z(n4366) );
  NAND U4549 ( .A(n4367), .B(n4366), .Z(n4392) );
  XOR U4550 ( .A(n4391), .B(n4392), .Z(n4394) );
  XNOR U4551 ( .A(n4393), .B(n4394), .Z(n4452) );
  NANDN U4552 ( .A(n4369), .B(n4368), .Z(n4373) );
  NAND U4553 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U4554 ( .A(n4373), .B(n4372), .Z(n4453) );
  XNOR U4555 ( .A(n4452), .B(n4453), .Z(n4454) );
  XOR U4556 ( .A(n4455), .B(n4454), .Z(n4385) );
  NANDN U4557 ( .A(n4375), .B(n4374), .Z(n4379) );
  NANDN U4558 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U4559 ( .A(n4379), .B(n4378), .Z(n4386) );
  XNOR U4560 ( .A(n4385), .B(n4386), .Z(n4387) );
  XNOR U4561 ( .A(n4388), .B(n4387), .Z(n4458) );
  XNOR U4562 ( .A(n4458), .B(sreg[175]), .Z(n4460) );
  NAND U4563 ( .A(n4380), .B(sreg[174]), .Z(n4384) );
  OR U4564 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U4565 ( .A(n4384), .B(n4383), .Z(n4459) );
  XOR U4566 ( .A(n4460), .B(n4459), .Z(c[175]) );
  NANDN U4567 ( .A(n4386), .B(n4385), .Z(n4390) );
  NAND U4568 ( .A(n4388), .B(n4387), .Z(n4389) );
  NAND U4569 ( .A(n4390), .B(n4389), .Z(n4466) );
  NANDN U4570 ( .A(n4392), .B(n4391), .Z(n4396) );
  OR U4571 ( .A(n4394), .B(n4393), .Z(n4395) );
  NAND U4572 ( .A(n4396), .B(n4395), .Z(n4533) );
  NANDN U4573 ( .A(n4398), .B(n4397), .Z(n4402) );
  OR U4574 ( .A(n4400), .B(n4399), .Z(n4401) );
  NAND U4575 ( .A(n4402), .B(n4401), .Z(n4521) );
  NAND U4576 ( .A(b[0]), .B(a[64]), .Z(n4403) );
  XNOR U4577 ( .A(b[1]), .B(n4403), .Z(n4405) );
  NAND U4578 ( .A(a[63]), .B(n72), .Z(n4404) );
  AND U4579 ( .A(n4405), .B(n4404), .Z(n4497) );
  XNOR U4580 ( .A(n10050), .B(n4556), .Z(n4506) );
  OR U4581 ( .A(n4506), .B(n10051), .Z(n4408) );
  NANDN U4582 ( .A(n4406), .B(n10070), .Z(n4407) );
  AND U4583 ( .A(n4408), .B(n4407), .Z(n4498) );
  XOR U4584 ( .A(n4497), .B(n4498), .Z(n4500) );
  NAND U4585 ( .A(a[48]), .B(b[15]), .Z(n4499) );
  XOR U4586 ( .A(n4500), .B(n4499), .Z(n4518) );
  XNOR U4587 ( .A(n9622), .B(n5180), .Z(n4509) );
  OR U4588 ( .A(n4509), .B(n9623), .Z(n4411) );
  NANDN U4589 ( .A(n4409), .B(n9680), .Z(n4410) );
  NAND U4590 ( .A(n4411), .B(n4410), .Z(n4494) );
  XNOR U4591 ( .A(n9872), .B(n5051), .Z(n4512) );
  NANDN U4592 ( .A(n4512), .B(n9746), .Z(n4414) );
  NANDN U4593 ( .A(n4412), .B(n9747), .Z(n4413) );
  NAND U4594 ( .A(n4414), .B(n4413), .Z(n4491) );
  IV U4595 ( .A(a[62]), .Z(n5336) );
  XNOR U4596 ( .A(n74), .B(n5336), .Z(n4515) );
  NANDN U4597 ( .A(n4515), .B(n9485), .Z(n4417) );
  NANDN U4598 ( .A(n4415), .B(n9484), .Z(n4416) );
  AND U4599 ( .A(n4417), .B(n4416), .Z(n4492) );
  XNOR U4600 ( .A(n4491), .B(n4492), .Z(n4493) );
  XOR U4601 ( .A(n4494), .B(n4493), .Z(n4519) );
  XOR U4602 ( .A(n4518), .B(n4519), .Z(n4520) );
  XNOR U4603 ( .A(n4521), .B(n4520), .Z(n4469) );
  NAND U4604 ( .A(n4419), .B(n4418), .Z(n4423) );
  NAND U4605 ( .A(n4421), .B(n4420), .Z(n4422) );
  NAND U4606 ( .A(n4423), .B(n4422), .Z(n4470) );
  XOR U4607 ( .A(n4469), .B(n4470), .Z(n4472) );
  XNOR U4608 ( .A(n9967), .B(n4712), .Z(n4475) );
  OR U4609 ( .A(n4475), .B(n10020), .Z(n4426) );
  NANDN U4610 ( .A(n4424), .B(n9968), .Z(n4425) );
  NAND U4611 ( .A(n4426), .B(n4425), .Z(n4488) );
  XNOR U4612 ( .A(n75), .B(n4427), .Z(n4479) );
  OR U4613 ( .A(n4479), .B(n10106), .Z(n4430) );
  NANDN U4614 ( .A(n4428), .B(n10107), .Z(n4429) );
  NAND U4615 ( .A(n4430), .B(n4429), .Z(n4485) );
  XNOR U4616 ( .A(n9984), .B(n4868), .Z(n4482) );
  NANDN U4617 ( .A(n4482), .B(n9865), .Z(n4433) );
  NANDN U4618 ( .A(n4431), .B(n9930), .Z(n4432) );
  AND U4619 ( .A(n4433), .B(n4432), .Z(n4486) );
  XNOR U4620 ( .A(n4485), .B(n4486), .Z(n4487) );
  XNOR U4621 ( .A(n4488), .B(n4487), .Z(n4524) );
  NANDN U4622 ( .A(n4435), .B(n4434), .Z(n4439) );
  NAND U4623 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U4624 ( .A(n4439), .B(n4438), .Z(n4525) );
  XNOR U4625 ( .A(n4524), .B(n4525), .Z(n4526) );
  NANDN U4626 ( .A(n4441), .B(n4440), .Z(n4445) );
  NAND U4627 ( .A(n4443), .B(n4442), .Z(n4444) );
  AND U4628 ( .A(n4445), .B(n4444), .Z(n4527) );
  XNOR U4629 ( .A(n4526), .B(n4527), .Z(n4471) );
  XNOR U4630 ( .A(n4472), .B(n4471), .Z(n4530) );
  NANDN U4631 ( .A(n4447), .B(n4446), .Z(n4451) );
  NAND U4632 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U4633 ( .A(n4451), .B(n4450), .Z(n4531) );
  XNOR U4634 ( .A(n4530), .B(n4531), .Z(n4532) );
  XOR U4635 ( .A(n4533), .B(n4532), .Z(n4463) );
  NANDN U4636 ( .A(n4453), .B(n4452), .Z(n4457) );
  NANDN U4637 ( .A(n4455), .B(n4454), .Z(n4456) );
  NAND U4638 ( .A(n4457), .B(n4456), .Z(n4464) );
  XNOR U4639 ( .A(n4463), .B(n4464), .Z(n4465) );
  XNOR U4640 ( .A(n4466), .B(n4465), .Z(n4536) );
  XNOR U4641 ( .A(n4536), .B(sreg[176]), .Z(n4538) );
  NAND U4642 ( .A(n4458), .B(sreg[175]), .Z(n4462) );
  OR U4643 ( .A(n4460), .B(n4459), .Z(n4461) );
  AND U4644 ( .A(n4462), .B(n4461), .Z(n4537) );
  XOR U4645 ( .A(n4538), .B(n4537), .Z(c[176]) );
  NANDN U4646 ( .A(n4464), .B(n4463), .Z(n4468) );
  NAND U4647 ( .A(n4466), .B(n4465), .Z(n4467) );
  NAND U4648 ( .A(n4468), .B(n4467), .Z(n4544) );
  NANDN U4649 ( .A(n4470), .B(n4469), .Z(n4474) );
  OR U4650 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U4651 ( .A(n4474), .B(n4473), .Z(n4611) );
  XNOR U4652 ( .A(n9967), .B(n4790), .Z(n4553) );
  OR U4653 ( .A(n4553), .B(n10020), .Z(n4477) );
  NANDN U4654 ( .A(n4475), .B(n9968), .Z(n4476) );
  NAND U4655 ( .A(n4477), .B(n4476), .Z(n4566) );
  XNOR U4656 ( .A(n75), .B(n4478), .Z(n4557) );
  OR U4657 ( .A(n4557), .B(n10106), .Z(n4481) );
  NANDN U4658 ( .A(n4479), .B(n10107), .Z(n4480) );
  NAND U4659 ( .A(n4481), .B(n4480), .Z(n4563) );
  XNOR U4660 ( .A(n9984), .B(n4973), .Z(n4560) );
  NANDN U4661 ( .A(n4560), .B(n9865), .Z(n4484) );
  NANDN U4662 ( .A(n4482), .B(n9930), .Z(n4483) );
  AND U4663 ( .A(n4484), .B(n4483), .Z(n4564) );
  XNOR U4664 ( .A(n4563), .B(n4564), .Z(n4565) );
  XNOR U4665 ( .A(n4566), .B(n4565), .Z(n4602) );
  NANDN U4666 ( .A(n4486), .B(n4485), .Z(n4490) );
  NAND U4667 ( .A(n4488), .B(n4487), .Z(n4489) );
  NAND U4668 ( .A(n4490), .B(n4489), .Z(n4603) );
  XNOR U4669 ( .A(n4602), .B(n4603), .Z(n4604) );
  NANDN U4670 ( .A(n4492), .B(n4491), .Z(n4496) );
  NAND U4671 ( .A(n4494), .B(n4493), .Z(n4495) );
  AND U4672 ( .A(n4496), .B(n4495), .Z(n4605) );
  XNOR U4673 ( .A(n4604), .B(n4605), .Z(n4549) );
  NANDN U4674 ( .A(n4498), .B(n4497), .Z(n4502) );
  OR U4675 ( .A(n4500), .B(n4499), .Z(n4501) );
  NAND U4676 ( .A(n4502), .B(n4501), .Z(n4599) );
  NAND U4677 ( .A(b[0]), .B(a[65]), .Z(n4503) );
  XNOR U4678 ( .A(b[1]), .B(n4503), .Z(n4505) );
  NAND U4679 ( .A(a[64]), .B(n72), .Z(n4504) );
  AND U4680 ( .A(n4505), .B(n4504), .Z(n4575) );
  XNOR U4681 ( .A(n10050), .B(n4661), .Z(n4584) );
  OR U4682 ( .A(n4584), .B(n10051), .Z(n4508) );
  NANDN U4683 ( .A(n4506), .B(n10070), .Z(n4507) );
  AND U4684 ( .A(n4508), .B(n4507), .Z(n4576) );
  XOR U4685 ( .A(n4575), .B(n4576), .Z(n4578) );
  NAND U4686 ( .A(a[49]), .B(b[15]), .Z(n4577) );
  XOR U4687 ( .A(n4578), .B(n4577), .Z(n4596) );
  XNOR U4688 ( .A(n9622), .B(n5258), .Z(n4587) );
  OR U4689 ( .A(n4587), .B(n9623), .Z(n4511) );
  NANDN U4690 ( .A(n4509), .B(n9680), .Z(n4510) );
  NAND U4691 ( .A(n4511), .B(n4510), .Z(n4572) );
  XNOR U4692 ( .A(n9872), .B(n5102), .Z(n4590) );
  NANDN U4693 ( .A(n4590), .B(n9746), .Z(n4514) );
  NANDN U4694 ( .A(n4512), .B(n9747), .Z(n4513) );
  NAND U4695 ( .A(n4514), .B(n4513), .Z(n4569) );
  IV U4696 ( .A(a[63]), .Z(n5414) );
  XNOR U4697 ( .A(n74), .B(n5414), .Z(n4593) );
  NANDN U4698 ( .A(n4593), .B(n9485), .Z(n4517) );
  NANDN U4699 ( .A(n4515), .B(n9484), .Z(n4516) );
  AND U4700 ( .A(n4517), .B(n4516), .Z(n4570) );
  XNOR U4701 ( .A(n4569), .B(n4570), .Z(n4571) );
  XOR U4702 ( .A(n4572), .B(n4571), .Z(n4597) );
  XOR U4703 ( .A(n4596), .B(n4597), .Z(n4598) );
  XNOR U4704 ( .A(n4599), .B(n4598), .Z(n4547) );
  NAND U4705 ( .A(n4519), .B(n4518), .Z(n4523) );
  NAND U4706 ( .A(n4521), .B(n4520), .Z(n4522) );
  NAND U4707 ( .A(n4523), .B(n4522), .Z(n4548) );
  XOR U4708 ( .A(n4547), .B(n4548), .Z(n4550) );
  XNOR U4709 ( .A(n4549), .B(n4550), .Z(n4608) );
  NANDN U4710 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U4711 ( .A(n4527), .B(n4526), .Z(n4528) );
  NAND U4712 ( .A(n4529), .B(n4528), .Z(n4609) );
  XNOR U4713 ( .A(n4608), .B(n4609), .Z(n4610) );
  XOR U4714 ( .A(n4611), .B(n4610), .Z(n4541) );
  NANDN U4715 ( .A(n4531), .B(n4530), .Z(n4535) );
  NANDN U4716 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U4717 ( .A(n4535), .B(n4534), .Z(n4542) );
  XNOR U4718 ( .A(n4541), .B(n4542), .Z(n4543) );
  XNOR U4719 ( .A(n4544), .B(n4543), .Z(n4614) );
  XNOR U4720 ( .A(n4614), .B(sreg[177]), .Z(n4616) );
  NAND U4721 ( .A(n4536), .B(sreg[176]), .Z(n4540) );
  OR U4722 ( .A(n4538), .B(n4537), .Z(n4539) );
  AND U4723 ( .A(n4540), .B(n4539), .Z(n4615) );
  XOR U4724 ( .A(n4616), .B(n4615), .Z(c[177]) );
  NANDN U4725 ( .A(n4542), .B(n4541), .Z(n4546) );
  NAND U4726 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U4727 ( .A(n4546), .B(n4545), .Z(n4622) );
  NANDN U4728 ( .A(n4548), .B(n4547), .Z(n4552) );
  OR U4729 ( .A(n4550), .B(n4549), .Z(n4551) );
  NAND U4730 ( .A(n4552), .B(n4551), .Z(n4689) );
  XNOR U4731 ( .A(n9967), .B(n4868), .Z(n4658) );
  OR U4732 ( .A(n4658), .B(n10020), .Z(n4555) );
  NANDN U4733 ( .A(n4553), .B(n9968), .Z(n4554) );
  NAND U4734 ( .A(n4555), .B(n4554), .Z(n4671) );
  XNOR U4735 ( .A(n75), .B(n4556), .Z(n4662) );
  OR U4736 ( .A(n4662), .B(n10106), .Z(n4559) );
  NANDN U4737 ( .A(n4557), .B(n10107), .Z(n4558) );
  NAND U4738 ( .A(n4559), .B(n4558), .Z(n4668) );
  XNOR U4739 ( .A(n9984), .B(n5051), .Z(n4665) );
  NANDN U4740 ( .A(n4665), .B(n9865), .Z(n4562) );
  NANDN U4741 ( .A(n4560), .B(n9930), .Z(n4561) );
  AND U4742 ( .A(n4562), .B(n4561), .Z(n4669) );
  XNOR U4743 ( .A(n4668), .B(n4669), .Z(n4670) );
  XNOR U4744 ( .A(n4671), .B(n4670), .Z(n4680) );
  NANDN U4745 ( .A(n4564), .B(n4563), .Z(n4568) );
  NAND U4746 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U4747 ( .A(n4568), .B(n4567), .Z(n4681) );
  XNOR U4748 ( .A(n4680), .B(n4681), .Z(n4682) );
  NANDN U4749 ( .A(n4570), .B(n4569), .Z(n4574) );
  NAND U4750 ( .A(n4572), .B(n4571), .Z(n4573) );
  AND U4751 ( .A(n4574), .B(n4573), .Z(n4683) );
  XNOR U4752 ( .A(n4682), .B(n4683), .Z(n4627) );
  NANDN U4753 ( .A(n4576), .B(n4575), .Z(n4580) );
  OR U4754 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U4755 ( .A(n4580), .B(n4579), .Z(n4655) );
  NAND U4756 ( .A(b[0]), .B(a[66]), .Z(n4581) );
  XNOR U4757 ( .A(b[1]), .B(n4581), .Z(n4583) );
  NAND U4758 ( .A(a[65]), .B(n72), .Z(n4582) );
  AND U4759 ( .A(n4583), .B(n4582), .Z(n4631) );
  XNOR U4760 ( .A(n10050), .B(n4712), .Z(n4637) );
  OR U4761 ( .A(n4637), .B(n10051), .Z(n4586) );
  NANDN U4762 ( .A(n4584), .B(n10070), .Z(n4585) );
  AND U4763 ( .A(n4586), .B(n4585), .Z(n4632) );
  XOR U4764 ( .A(n4631), .B(n4632), .Z(n4634) );
  NAND U4765 ( .A(a[50]), .B(b[15]), .Z(n4633) );
  XOR U4766 ( .A(n4634), .B(n4633), .Z(n4652) );
  XNOR U4767 ( .A(n9622), .B(n5336), .Z(n4643) );
  OR U4768 ( .A(n4643), .B(n9623), .Z(n4589) );
  NANDN U4769 ( .A(n4587), .B(n9680), .Z(n4588) );
  NAND U4770 ( .A(n4589), .B(n4588), .Z(n4677) );
  XNOR U4771 ( .A(n9872), .B(n5180), .Z(n4646) );
  NANDN U4772 ( .A(n4646), .B(n9746), .Z(n4592) );
  NANDN U4773 ( .A(n4590), .B(n9747), .Z(n4591) );
  NAND U4774 ( .A(n4592), .B(n4591), .Z(n4674) );
  IV U4775 ( .A(a[64]), .Z(n5492) );
  XNOR U4776 ( .A(n74), .B(n5492), .Z(n4649) );
  NANDN U4777 ( .A(n4649), .B(n9485), .Z(n4595) );
  NANDN U4778 ( .A(n4593), .B(n9484), .Z(n4594) );
  AND U4779 ( .A(n4595), .B(n4594), .Z(n4675) );
  XNOR U4780 ( .A(n4674), .B(n4675), .Z(n4676) );
  XOR U4781 ( .A(n4677), .B(n4676), .Z(n4653) );
  XOR U4782 ( .A(n4652), .B(n4653), .Z(n4654) );
  XNOR U4783 ( .A(n4655), .B(n4654), .Z(n4625) );
  NAND U4784 ( .A(n4597), .B(n4596), .Z(n4601) );
  NAND U4785 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U4786 ( .A(n4601), .B(n4600), .Z(n4626) );
  XOR U4787 ( .A(n4625), .B(n4626), .Z(n4628) );
  XNOR U4788 ( .A(n4627), .B(n4628), .Z(n4686) );
  NANDN U4789 ( .A(n4603), .B(n4602), .Z(n4607) );
  NAND U4790 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U4791 ( .A(n4607), .B(n4606), .Z(n4687) );
  XNOR U4792 ( .A(n4686), .B(n4687), .Z(n4688) );
  XOR U4793 ( .A(n4689), .B(n4688), .Z(n4619) );
  NANDN U4794 ( .A(n4609), .B(n4608), .Z(n4613) );
  NANDN U4795 ( .A(n4611), .B(n4610), .Z(n4612) );
  NAND U4796 ( .A(n4613), .B(n4612), .Z(n4620) );
  XNOR U4797 ( .A(n4619), .B(n4620), .Z(n4621) );
  XNOR U4798 ( .A(n4622), .B(n4621), .Z(n4692) );
  XNOR U4799 ( .A(n4692), .B(sreg[178]), .Z(n4694) );
  NAND U4800 ( .A(n4614), .B(sreg[177]), .Z(n4618) );
  OR U4801 ( .A(n4616), .B(n4615), .Z(n4617) );
  AND U4802 ( .A(n4618), .B(n4617), .Z(n4693) );
  XOR U4803 ( .A(n4694), .B(n4693), .Z(c[178]) );
  NANDN U4804 ( .A(n4620), .B(n4619), .Z(n4624) );
  NAND U4805 ( .A(n4622), .B(n4621), .Z(n4623) );
  NAND U4806 ( .A(n4624), .B(n4623), .Z(n4700) );
  NANDN U4807 ( .A(n4626), .B(n4625), .Z(n4630) );
  OR U4808 ( .A(n4628), .B(n4627), .Z(n4629) );
  NAND U4809 ( .A(n4630), .B(n4629), .Z(n4767) );
  NANDN U4810 ( .A(n4632), .B(n4631), .Z(n4636) );
  OR U4811 ( .A(n4634), .B(n4633), .Z(n4635) );
  NAND U4812 ( .A(n4636), .B(n4635), .Z(n4755) );
  XNOR U4813 ( .A(n10050), .B(n4790), .Z(n4740) );
  OR U4814 ( .A(n4740), .B(n10051), .Z(n4639) );
  NANDN U4815 ( .A(n4637), .B(n10070), .Z(n4638) );
  AND U4816 ( .A(n4639), .B(n4638), .Z(n4732) );
  NAND U4817 ( .A(b[0]), .B(a[67]), .Z(n4640) );
  XNOR U4818 ( .A(b[1]), .B(n4640), .Z(n4642) );
  NAND U4819 ( .A(a[66]), .B(n72), .Z(n4641) );
  AND U4820 ( .A(n4642), .B(n4641), .Z(n4731) );
  XOR U4821 ( .A(n4732), .B(n4731), .Z(n4734) );
  NAND U4822 ( .A(a[51]), .B(b[15]), .Z(n4733) );
  XOR U4823 ( .A(n4734), .B(n4733), .Z(n4752) );
  XNOR U4824 ( .A(n9622), .B(n5414), .Z(n4743) );
  OR U4825 ( .A(n4743), .B(n9623), .Z(n4645) );
  NANDN U4826 ( .A(n4643), .B(n9680), .Z(n4644) );
  NAND U4827 ( .A(n4645), .B(n4644), .Z(n4728) );
  XNOR U4828 ( .A(n9872), .B(n5258), .Z(n4746) );
  NANDN U4829 ( .A(n4746), .B(n9746), .Z(n4648) );
  NANDN U4830 ( .A(n4646), .B(n9747), .Z(n4647) );
  NAND U4831 ( .A(n4648), .B(n4647), .Z(n4725) );
  IV U4832 ( .A(a[65]), .Z(n5570) );
  XNOR U4833 ( .A(n74), .B(n5570), .Z(n4749) );
  NANDN U4834 ( .A(n4749), .B(n9485), .Z(n4651) );
  NANDN U4835 ( .A(n4649), .B(n9484), .Z(n4650) );
  AND U4836 ( .A(n4651), .B(n4650), .Z(n4726) );
  XNOR U4837 ( .A(n4725), .B(n4726), .Z(n4727) );
  XOR U4838 ( .A(n4728), .B(n4727), .Z(n4753) );
  XOR U4839 ( .A(n4752), .B(n4753), .Z(n4754) );
  XNOR U4840 ( .A(n4755), .B(n4754), .Z(n4703) );
  NAND U4841 ( .A(n4653), .B(n4652), .Z(n4657) );
  NAND U4842 ( .A(n4655), .B(n4654), .Z(n4656) );
  NAND U4843 ( .A(n4657), .B(n4656), .Z(n4704) );
  XOR U4844 ( .A(n4703), .B(n4704), .Z(n4706) );
  XNOR U4845 ( .A(n9967), .B(n4973), .Z(n4709) );
  OR U4846 ( .A(n4709), .B(n10020), .Z(n4660) );
  NANDN U4847 ( .A(n4658), .B(n9968), .Z(n4659) );
  NAND U4848 ( .A(n4660), .B(n4659), .Z(n4722) );
  XNOR U4849 ( .A(n75), .B(n4661), .Z(n4713) );
  OR U4850 ( .A(n4713), .B(n10106), .Z(n4664) );
  NANDN U4851 ( .A(n4662), .B(n10107), .Z(n4663) );
  NAND U4852 ( .A(n4664), .B(n4663), .Z(n4719) );
  XNOR U4853 ( .A(n9984), .B(n5102), .Z(n4716) );
  NANDN U4854 ( .A(n4716), .B(n9865), .Z(n4667) );
  NANDN U4855 ( .A(n4665), .B(n9930), .Z(n4666) );
  AND U4856 ( .A(n4667), .B(n4666), .Z(n4720) );
  XNOR U4857 ( .A(n4719), .B(n4720), .Z(n4721) );
  XNOR U4858 ( .A(n4722), .B(n4721), .Z(n4758) );
  NANDN U4859 ( .A(n4669), .B(n4668), .Z(n4673) );
  NAND U4860 ( .A(n4671), .B(n4670), .Z(n4672) );
  NAND U4861 ( .A(n4673), .B(n4672), .Z(n4759) );
  XNOR U4862 ( .A(n4758), .B(n4759), .Z(n4760) );
  NANDN U4863 ( .A(n4675), .B(n4674), .Z(n4679) );
  NAND U4864 ( .A(n4677), .B(n4676), .Z(n4678) );
  AND U4865 ( .A(n4679), .B(n4678), .Z(n4761) );
  XNOR U4866 ( .A(n4760), .B(n4761), .Z(n4705) );
  XNOR U4867 ( .A(n4706), .B(n4705), .Z(n4764) );
  NANDN U4868 ( .A(n4681), .B(n4680), .Z(n4685) );
  NAND U4869 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U4870 ( .A(n4685), .B(n4684), .Z(n4765) );
  XNOR U4871 ( .A(n4764), .B(n4765), .Z(n4766) );
  XOR U4872 ( .A(n4767), .B(n4766), .Z(n4697) );
  NANDN U4873 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U4874 ( .A(n4689), .B(n4688), .Z(n4690) );
  NAND U4875 ( .A(n4691), .B(n4690), .Z(n4698) );
  XNOR U4876 ( .A(n4697), .B(n4698), .Z(n4699) );
  XNOR U4877 ( .A(n4700), .B(n4699), .Z(n4770) );
  XNOR U4878 ( .A(n4770), .B(sreg[179]), .Z(n4772) );
  NAND U4879 ( .A(n4692), .B(sreg[178]), .Z(n4696) );
  OR U4880 ( .A(n4694), .B(n4693), .Z(n4695) );
  AND U4881 ( .A(n4696), .B(n4695), .Z(n4771) );
  XOR U4882 ( .A(n4772), .B(n4771), .Z(c[179]) );
  NANDN U4883 ( .A(n4698), .B(n4697), .Z(n4702) );
  NAND U4884 ( .A(n4700), .B(n4699), .Z(n4701) );
  NAND U4885 ( .A(n4702), .B(n4701), .Z(n4778) );
  NANDN U4886 ( .A(n4704), .B(n4703), .Z(n4708) );
  OR U4887 ( .A(n4706), .B(n4705), .Z(n4707) );
  NAND U4888 ( .A(n4708), .B(n4707), .Z(n4845) );
  XNOR U4889 ( .A(n9967), .B(n5051), .Z(n4787) );
  OR U4890 ( .A(n4787), .B(n10020), .Z(n4711) );
  NANDN U4891 ( .A(n4709), .B(n9968), .Z(n4710) );
  NAND U4892 ( .A(n4711), .B(n4710), .Z(n4800) );
  XNOR U4893 ( .A(n75), .B(n4712), .Z(n4791) );
  OR U4894 ( .A(n4791), .B(n10106), .Z(n4715) );
  NANDN U4895 ( .A(n4713), .B(n10107), .Z(n4714) );
  NAND U4896 ( .A(n4715), .B(n4714), .Z(n4797) );
  XNOR U4897 ( .A(n9984), .B(n5180), .Z(n4794) );
  NANDN U4898 ( .A(n4794), .B(n9865), .Z(n4718) );
  NANDN U4899 ( .A(n4716), .B(n9930), .Z(n4717) );
  AND U4900 ( .A(n4718), .B(n4717), .Z(n4798) );
  XNOR U4901 ( .A(n4797), .B(n4798), .Z(n4799) );
  XNOR U4902 ( .A(n4800), .B(n4799), .Z(n4836) );
  NANDN U4903 ( .A(n4720), .B(n4719), .Z(n4724) );
  NAND U4904 ( .A(n4722), .B(n4721), .Z(n4723) );
  NAND U4905 ( .A(n4724), .B(n4723), .Z(n4837) );
  XNOR U4906 ( .A(n4836), .B(n4837), .Z(n4838) );
  NANDN U4907 ( .A(n4726), .B(n4725), .Z(n4730) );
  NAND U4908 ( .A(n4728), .B(n4727), .Z(n4729) );
  AND U4909 ( .A(n4730), .B(n4729), .Z(n4839) );
  XNOR U4910 ( .A(n4838), .B(n4839), .Z(n4783) );
  NANDN U4911 ( .A(n4732), .B(n4731), .Z(n4736) );
  OR U4912 ( .A(n4734), .B(n4733), .Z(n4735) );
  NAND U4913 ( .A(n4736), .B(n4735), .Z(n4833) );
  NAND U4914 ( .A(b[0]), .B(a[68]), .Z(n4737) );
  XNOR U4915 ( .A(b[1]), .B(n4737), .Z(n4739) );
  NAND U4916 ( .A(a[67]), .B(n72), .Z(n4738) );
  AND U4917 ( .A(n4739), .B(n4738), .Z(n4809) );
  XNOR U4918 ( .A(n10050), .B(n4868), .Z(n4818) );
  OR U4919 ( .A(n4818), .B(n10051), .Z(n4742) );
  NANDN U4920 ( .A(n4740), .B(n10070), .Z(n4741) );
  AND U4921 ( .A(n4742), .B(n4741), .Z(n4810) );
  XOR U4922 ( .A(n4809), .B(n4810), .Z(n4812) );
  NAND U4923 ( .A(a[52]), .B(b[15]), .Z(n4811) );
  XOR U4924 ( .A(n4812), .B(n4811), .Z(n4830) );
  XNOR U4925 ( .A(n9622), .B(n5492), .Z(n4821) );
  OR U4926 ( .A(n4821), .B(n9623), .Z(n4745) );
  NANDN U4927 ( .A(n4743), .B(n9680), .Z(n4744) );
  NAND U4928 ( .A(n4745), .B(n4744), .Z(n4806) );
  XNOR U4929 ( .A(n9872), .B(n5336), .Z(n4824) );
  NANDN U4930 ( .A(n4824), .B(n9746), .Z(n4748) );
  NANDN U4931 ( .A(n4746), .B(n9747), .Z(n4747) );
  NAND U4932 ( .A(n4748), .B(n4747), .Z(n4803) );
  IV U4933 ( .A(a[66]), .Z(n5675) );
  XNOR U4934 ( .A(n74), .B(n5675), .Z(n4827) );
  NANDN U4935 ( .A(n4827), .B(n9485), .Z(n4751) );
  NANDN U4936 ( .A(n4749), .B(n9484), .Z(n4750) );
  AND U4937 ( .A(n4751), .B(n4750), .Z(n4804) );
  XNOR U4938 ( .A(n4803), .B(n4804), .Z(n4805) );
  XOR U4939 ( .A(n4806), .B(n4805), .Z(n4831) );
  XOR U4940 ( .A(n4830), .B(n4831), .Z(n4832) );
  XNOR U4941 ( .A(n4833), .B(n4832), .Z(n4781) );
  NAND U4942 ( .A(n4753), .B(n4752), .Z(n4757) );
  NAND U4943 ( .A(n4755), .B(n4754), .Z(n4756) );
  NAND U4944 ( .A(n4757), .B(n4756), .Z(n4782) );
  XOR U4945 ( .A(n4781), .B(n4782), .Z(n4784) );
  XNOR U4946 ( .A(n4783), .B(n4784), .Z(n4842) );
  NANDN U4947 ( .A(n4759), .B(n4758), .Z(n4763) );
  NAND U4948 ( .A(n4761), .B(n4760), .Z(n4762) );
  NAND U4949 ( .A(n4763), .B(n4762), .Z(n4843) );
  XNOR U4950 ( .A(n4842), .B(n4843), .Z(n4844) );
  XOR U4951 ( .A(n4845), .B(n4844), .Z(n4775) );
  NANDN U4952 ( .A(n4765), .B(n4764), .Z(n4769) );
  NANDN U4953 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U4954 ( .A(n4769), .B(n4768), .Z(n4776) );
  XNOR U4955 ( .A(n4775), .B(n4776), .Z(n4777) );
  XNOR U4956 ( .A(n4778), .B(n4777), .Z(n4848) );
  XNOR U4957 ( .A(n4848), .B(sreg[180]), .Z(n4850) );
  NAND U4958 ( .A(n4770), .B(sreg[179]), .Z(n4774) );
  OR U4959 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U4960 ( .A(n4774), .B(n4773), .Z(n4849) );
  XOR U4961 ( .A(n4850), .B(n4849), .Z(c[180]) );
  NANDN U4962 ( .A(n4776), .B(n4775), .Z(n4780) );
  NAND U4963 ( .A(n4778), .B(n4777), .Z(n4779) );
  NAND U4964 ( .A(n4780), .B(n4779), .Z(n4856) );
  NANDN U4965 ( .A(n4782), .B(n4781), .Z(n4786) );
  OR U4966 ( .A(n4784), .B(n4783), .Z(n4785) );
  NAND U4967 ( .A(n4786), .B(n4785), .Z(n4923) );
  XNOR U4968 ( .A(n9967), .B(n5102), .Z(n4865) );
  OR U4969 ( .A(n4865), .B(n10020), .Z(n4789) );
  NANDN U4970 ( .A(n4787), .B(n9968), .Z(n4788) );
  NAND U4971 ( .A(n4789), .B(n4788), .Z(n4878) );
  XNOR U4972 ( .A(n75), .B(n4790), .Z(n4869) );
  OR U4973 ( .A(n4869), .B(n10106), .Z(n4793) );
  NANDN U4974 ( .A(n4791), .B(n10107), .Z(n4792) );
  NAND U4975 ( .A(n4793), .B(n4792), .Z(n4875) );
  XNOR U4976 ( .A(n9984), .B(n5258), .Z(n4872) );
  NANDN U4977 ( .A(n4872), .B(n9865), .Z(n4796) );
  NANDN U4978 ( .A(n4794), .B(n9930), .Z(n4795) );
  AND U4979 ( .A(n4796), .B(n4795), .Z(n4876) );
  XNOR U4980 ( .A(n4875), .B(n4876), .Z(n4877) );
  XNOR U4981 ( .A(n4878), .B(n4877), .Z(n4914) );
  NANDN U4982 ( .A(n4798), .B(n4797), .Z(n4802) );
  NAND U4983 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U4984 ( .A(n4802), .B(n4801), .Z(n4915) );
  XNOR U4985 ( .A(n4914), .B(n4915), .Z(n4916) );
  NANDN U4986 ( .A(n4804), .B(n4803), .Z(n4808) );
  NAND U4987 ( .A(n4806), .B(n4805), .Z(n4807) );
  AND U4988 ( .A(n4808), .B(n4807), .Z(n4917) );
  XNOR U4989 ( .A(n4916), .B(n4917), .Z(n4861) );
  NANDN U4990 ( .A(n4810), .B(n4809), .Z(n4814) );
  OR U4991 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U4992 ( .A(n4814), .B(n4813), .Z(n4911) );
  NAND U4993 ( .A(b[0]), .B(a[69]), .Z(n4815) );
  XNOR U4994 ( .A(b[1]), .B(n4815), .Z(n4817) );
  NAND U4995 ( .A(a[68]), .B(n72), .Z(n4816) );
  AND U4996 ( .A(n4817), .B(n4816), .Z(n4887) );
  XNOR U4997 ( .A(n10050), .B(n4973), .Z(n4893) );
  OR U4998 ( .A(n4893), .B(n10051), .Z(n4820) );
  NANDN U4999 ( .A(n4818), .B(n10070), .Z(n4819) );
  AND U5000 ( .A(n4820), .B(n4819), .Z(n4888) );
  XOR U5001 ( .A(n4887), .B(n4888), .Z(n4890) );
  NAND U5002 ( .A(a[53]), .B(b[15]), .Z(n4889) );
  XOR U5003 ( .A(n4890), .B(n4889), .Z(n4908) );
  XNOR U5004 ( .A(n9622), .B(n5570), .Z(n4899) );
  OR U5005 ( .A(n4899), .B(n9623), .Z(n4823) );
  NANDN U5006 ( .A(n4821), .B(n9680), .Z(n4822) );
  NAND U5007 ( .A(n4823), .B(n4822), .Z(n4884) );
  XNOR U5008 ( .A(n9872), .B(n5414), .Z(n4902) );
  NANDN U5009 ( .A(n4902), .B(n9746), .Z(n4826) );
  NANDN U5010 ( .A(n4824), .B(n9747), .Z(n4825) );
  NAND U5011 ( .A(n4826), .B(n4825), .Z(n4881) );
  IV U5012 ( .A(a[67]), .Z(n5726) );
  XNOR U5013 ( .A(n74), .B(n5726), .Z(n4905) );
  NANDN U5014 ( .A(n4905), .B(n9485), .Z(n4829) );
  NANDN U5015 ( .A(n4827), .B(n9484), .Z(n4828) );
  AND U5016 ( .A(n4829), .B(n4828), .Z(n4882) );
  XNOR U5017 ( .A(n4881), .B(n4882), .Z(n4883) );
  XOR U5018 ( .A(n4884), .B(n4883), .Z(n4909) );
  XOR U5019 ( .A(n4908), .B(n4909), .Z(n4910) );
  XNOR U5020 ( .A(n4911), .B(n4910), .Z(n4859) );
  NAND U5021 ( .A(n4831), .B(n4830), .Z(n4835) );
  NAND U5022 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5023 ( .A(n4835), .B(n4834), .Z(n4860) );
  XOR U5024 ( .A(n4859), .B(n4860), .Z(n4862) );
  XNOR U5025 ( .A(n4861), .B(n4862), .Z(n4920) );
  NANDN U5026 ( .A(n4837), .B(n4836), .Z(n4841) );
  NAND U5027 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5028 ( .A(n4841), .B(n4840), .Z(n4921) );
  XNOR U5029 ( .A(n4920), .B(n4921), .Z(n4922) );
  XOR U5030 ( .A(n4923), .B(n4922), .Z(n4853) );
  NANDN U5031 ( .A(n4843), .B(n4842), .Z(n4847) );
  NANDN U5032 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5033 ( .A(n4847), .B(n4846), .Z(n4854) );
  XNOR U5034 ( .A(n4853), .B(n4854), .Z(n4855) );
  XNOR U5035 ( .A(n4856), .B(n4855), .Z(n4926) );
  XNOR U5036 ( .A(n4926), .B(sreg[181]), .Z(n4928) );
  NAND U5037 ( .A(n4848), .B(sreg[180]), .Z(n4852) );
  OR U5038 ( .A(n4850), .B(n4849), .Z(n4851) );
  AND U5039 ( .A(n4852), .B(n4851), .Z(n4927) );
  XOR U5040 ( .A(n4928), .B(n4927), .Z(c[181]) );
  NANDN U5041 ( .A(n4854), .B(n4853), .Z(n4858) );
  NAND U5042 ( .A(n4856), .B(n4855), .Z(n4857) );
  NAND U5043 ( .A(n4858), .B(n4857), .Z(n4934) );
  NANDN U5044 ( .A(n4860), .B(n4859), .Z(n4864) );
  OR U5045 ( .A(n4862), .B(n4861), .Z(n4863) );
  NAND U5046 ( .A(n4864), .B(n4863), .Z(n5001) );
  XNOR U5047 ( .A(n9967), .B(n5180), .Z(n4970) );
  OR U5048 ( .A(n4970), .B(n10020), .Z(n4867) );
  NANDN U5049 ( .A(n4865), .B(n9968), .Z(n4866) );
  NAND U5050 ( .A(n4867), .B(n4866), .Z(n4983) );
  XNOR U5051 ( .A(n75), .B(n4868), .Z(n4974) );
  OR U5052 ( .A(n4974), .B(n10106), .Z(n4871) );
  NANDN U5053 ( .A(n4869), .B(n10107), .Z(n4870) );
  NAND U5054 ( .A(n4871), .B(n4870), .Z(n4980) );
  XNOR U5055 ( .A(n9984), .B(n5336), .Z(n4977) );
  NANDN U5056 ( .A(n4977), .B(n9865), .Z(n4874) );
  NANDN U5057 ( .A(n4872), .B(n9930), .Z(n4873) );
  AND U5058 ( .A(n4874), .B(n4873), .Z(n4981) );
  XNOR U5059 ( .A(n4980), .B(n4981), .Z(n4982) );
  XNOR U5060 ( .A(n4983), .B(n4982), .Z(n4992) );
  NANDN U5061 ( .A(n4876), .B(n4875), .Z(n4880) );
  NAND U5062 ( .A(n4878), .B(n4877), .Z(n4879) );
  NAND U5063 ( .A(n4880), .B(n4879), .Z(n4993) );
  XNOR U5064 ( .A(n4992), .B(n4993), .Z(n4994) );
  NANDN U5065 ( .A(n4882), .B(n4881), .Z(n4886) );
  NAND U5066 ( .A(n4884), .B(n4883), .Z(n4885) );
  AND U5067 ( .A(n4886), .B(n4885), .Z(n4995) );
  XNOR U5068 ( .A(n4994), .B(n4995), .Z(n4939) );
  NANDN U5069 ( .A(n4888), .B(n4887), .Z(n4892) );
  OR U5070 ( .A(n4890), .B(n4889), .Z(n4891) );
  NAND U5071 ( .A(n4892), .B(n4891), .Z(n4967) );
  XNOR U5072 ( .A(n10050), .B(n5051), .Z(n4952) );
  OR U5073 ( .A(n4952), .B(n10051), .Z(n4895) );
  NANDN U5074 ( .A(n4893), .B(n10070), .Z(n4894) );
  AND U5075 ( .A(n4895), .B(n4894), .Z(n4944) );
  NAND U5076 ( .A(b[0]), .B(a[70]), .Z(n4896) );
  XNOR U5077 ( .A(b[1]), .B(n4896), .Z(n4898) );
  NAND U5078 ( .A(a[69]), .B(n72), .Z(n4897) );
  AND U5079 ( .A(n4898), .B(n4897), .Z(n4943) );
  XOR U5080 ( .A(n4944), .B(n4943), .Z(n4946) );
  NAND U5081 ( .A(a[54]), .B(b[15]), .Z(n4945) );
  XOR U5082 ( .A(n4946), .B(n4945), .Z(n4964) );
  XNOR U5083 ( .A(n9622), .B(n5675), .Z(n4955) );
  OR U5084 ( .A(n4955), .B(n9623), .Z(n4901) );
  NANDN U5085 ( .A(n4899), .B(n9680), .Z(n4900) );
  NAND U5086 ( .A(n4901), .B(n4900), .Z(n4989) );
  XNOR U5087 ( .A(n9872), .B(n5492), .Z(n4958) );
  NANDN U5088 ( .A(n4958), .B(n9746), .Z(n4904) );
  NANDN U5089 ( .A(n4902), .B(n9747), .Z(n4903) );
  NAND U5090 ( .A(n4904), .B(n4903), .Z(n4986) );
  IV U5091 ( .A(a[68]), .Z(n5804) );
  XNOR U5092 ( .A(n74), .B(n5804), .Z(n4961) );
  NANDN U5093 ( .A(n4961), .B(n9485), .Z(n4907) );
  NANDN U5094 ( .A(n4905), .B(n9484), .Z(n4906) );
  AND U5095 ( .A(n4907), .B(n4906), .Z(n4987) );
  XNOR U5096 ( .A(n4986), .B(n4987), .Z(n4988) );
  XOR U5097 ( .A(n4989), .B(n4988), .Z(n4965) );
  XOR U5098 ( .A(n4964), .B(n4965), .Z(n4966) );
  XNOR U5099 ( .A(n4967), .B(n4966), .Z(n4937) );
  NAND U5100 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U5101 ( .A(n4911), .B(n4910), .Z(n4912) );
  NAND U5102 ( .A(n4913), .B(n4912), .Z(n4938) );
  XOR U5103 ( .A(n4937), .B(n4938), .Z(n4940) );
  XNOR U5104 ( .A(n4939), .B(n4940), .Z(n4998) );
  NANDN U5105 ( .A(n4915), .B(n4914), .Z(n4919) );
  NAND U5106 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U5107 ( .A(n4919), .B(n4918), .Z(n4999) );
  XNOR U5108 ( .A(n4998), .B(n4999), .Z(n5000) );
  XOR U5109 ( .A(n5001), .B(n5000), .Z(n4931) );
  NANDN U5110 ( .A(n4921), .B(n4920), .Z(n4925) );
  NANDN U5111 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U5112 ( .A(n4925), .B(n4924), .Z(n4932) );
  XNOR U5113 ( .A(n4931), .B(n4932), .Z(n4933) );
  XNOR U5114 ( .A(n4934), .B(n4933), .Z(n5004) );
  XNOR U5115 ( .A(n5004), .B(sreg[182]), .Z(n5006) );
  NAND U5116 ( .A(n4926), .B(sreg[181]), .Z(n4930) );
  OR U5117 ( .A(n4928), .B(n4927), .Z(n4929) );
  AND U5118 ( .A(n4930), .B(n4929), .Z(n5005) );
  XOR U5119 ( .A(n5006), .B(n5005), .Z(c[182]) );
  NANDN U5120 ( .A(n4932), .B(n4931), .Z(n4936) );
  NAND U5121 ( .A(n4934), .B(n4933), .Z(n4935) );
  NAND U5122 ( .A(n4936), .B(n4935), .Z(n5012) );
  NANDN U5123 ( .A(n4938), .B(n4937), .Z(n4942) );
  OR U5124 ( .A(n4940), .B(n4939), .Z(n4941) );
  NAND U5125 ( .A(n4942), .B(n4941), .Z(n5079) );
  NANDN U5126 ( .A(n4944), .B(n4943), .Z(n4948) );
  OR U5127 ( .A(n4946), .B(n4945), .Z(n4947) );
  NAND U5128 ( .A(n4948), .B(n4947), .Z(n5045) );
  NAND U5129 ( .A(b[0]), .B(a[71]), .Z(n4949) );
  XNOR U5130 ( .A(b[1]), .B(n4949), .Z(n4951) );
  NAND U5131 ( .A(a[70]), .B(n72), .Z(n4950) );
  AND U5132 ( .A(n4951), .B(n4950), .Z(n5021) );
  XNOR U5133 ( .A(n10050), .B(n5102), .Z(n5030) );
  OR U5134 ( .A(n5030), .B(n10051), .Z(n4954) );
  NANDN U5135 ( .A(n4952), .B(n10070), .Z(n4953) );
  AND U5136 ( .A(n4954), .B(n4953), .Z(n5022) );
  XOR U5137 ( .A(n5021), .B(n5022), .Z(n5024) );
  NAND U5138 ( .A(a[55]), .B(b[15]), .Z(n5023) );
  XOR U5139 ( .A(n5024), .B(n5023), .Z(n5042) );
  XNOR U5140 ( .A(n9622), .B(n5726), .Z(n5033) );
  OR U5141 ( .A(n5033), .B(n9623), .Z(n4957) );
  NANDN U5142 ( .A(n4955), .B(n9680), .Z(n4956) );
  NAND U5143 ( .A(n4957), .B(n4956), .Z(n5067) );
  XNOR U5144 ( .A(n9872), .B(n5570), .Z(n5036) );
  NANDN U5145 ( .A(n5036), .B(n9746), .Z(n4960) );
  NANDN U5146 ( .A(n4958), .B(n9747), .Z(n4959) );
  NAND U5147 ( .A(n4960), .B(n4959), .Z(n5064) );
  IV U5148 ( .A(a[69]), .Z(n5882) );
  XNOR U5149 ( .A(n74), .B(n5882), .Z(n5039) );
  NANDN U5150 ( .A(n5039), .B(n9485), .Z(n4963) );
  NANDN U5151 ( .A(n4961), .B(n9484), .Z(n4962) );
  AND U5152 ( .A(n4963), .B(n4962), .Z(n5065) );
  XNOR U5153 ( .A(n5064), .B(n5065), .Z(n5066) );
  XOR U5154 ( .A(n5067), .B(n5066), .Z(n5043) );
  XOR U5155 ( .A(n5042), .B(n5043), .Z(n5044) );
  XNOR U5156 ( .A(n5045), .B(n5044), .Z(n5015) );
  NAND U5157 ( .A(n4965), .B(n4964), .Z(n4969) );
  NAND U5158 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U5159 ( .A(n4969), .B(n4968), .Z(n5016) );
  XOR U5160 ( .A(n5015), .B(n5016), .Z(n5018) );
  XNOR U5161 ( .A(n9967), .B(n5258), .Z(n5048) );
  OR U5162 ( .A(n5048), .B(n10020), .Z(n4972) );
  NANDN U5163 ( .A(n4970), .B(n9968), .Z(n4971) );
  NAND U5164 ( .A(n4972), .B(n4971), .Z(n5061) );
  XNOR U5165 ( .A(n75), .B(n4973), .Z(n5052) );
  OR U5166 ( .A(n5052), .B(n10106), .Z(n4976) );
  NANDN U5167 ( .A(n4974), .B(n10107), .Z(n4975) );
  NAND U5168 ( .A(n4976), .B(n4975), .Z(n5058) );
  XNOR U5169 ( .A(n9984), .B(n5414), .Z(n5055) );
  NANDN U5170 ( .A(n5055), .B(n9865), .Z(n4979) );
  NANDN U5171 ( .A(n4977), .B(n9930), .Z(n4978) );
  AND U5172 ( .A(n4979), .B(n4978), .Z(n5059) );
  XNOR U5173 ( .A(n5058), .B(n5059), .Z(n5060) );
  XNOR U5174 ( .A(n5061), .B(n5060), .Z(n5070) );
  NANDN U5175 ( .A(n4981), .B(n4980), .Z(n4985) );
  NAND U5176 ( .A(n4983), .B(n4982), .Z(n4984) );
  NAND U5177 ( .A(n4985), .B(n4984), .Z(n5071) );
  XNOR U5178 ( .A(n5070), .B(n5071), .Z(n5072) );
  NANDN U5179 ( .A(n4987), .B(n4986), .Z(n4991) );
  NAND U5180 ( .A(n4989), .B(n4988), .Z(n4990) );
  AND U5181 ( .A(n4991), .B(n4990), .Z(n5073) );
  XNOR U5182 ( .A(n5072), .B(n5073), .Z(n5017) );
  XNOR U5183 ( .A(n5018), .B(n5017), .Z(n5076) );
  NANDN U5184 ( .A(n4993), .B(n4992), .Z(n4997) );
  NAND U5185 ( .A(n4995), .B(n4994), .Z(n4996) );
  NAND U5186 ( .A(n4997), .B(n4996), .Z(n5077) );
  XNOR U5187 ( .A(n5076), .B(n5077), .Z(n5078) );
  XOR U5188 ( .A(n5079), .B(n5078), .Z(n5009) );
  NANDN U5189 ( .A(n4999), .B(n4998), .Z(n5003) );
  NANDN U5190 ( .A(n5001), .B(n5000), .Z(n5002) );
  NAND U5191 ( .A(n5003), .B(n5002), .Z(n5010) );
  XNOR U5192 ( .A(n5009), .B(n5010), .Z(n5011) );
  XNOR U5193 ( .A(n5012), .B(n5011), .Z(n5082) );
  XNOR U5194 ( .A(n5082), .B(sreg[183]), .Z(n5084) );
  NAND U5195 ( .A(n5004), .B(sreg[182]), .Z(n5008) );
  OR U5196 ( .A(n5006), .B(n5005), .Z(n5007) );
  AND U5197 ( .A(n5008), .B(n5007), .Z(n5083) );
  XOR U5198 ( .A(n5084), .B(n5083), .Z(c[183]) );
  NANDN U5199 ( .A(n5010), .B(n5009), .Z(n5014) );
  NAND U5200 ( .A(n5012), .B(n5011), .Z(n5013) );
  NAND U5201 ( .A(n5014), .B(n5013), .Z(n5090) );
  NANDN U5202 ( .A(n5016), .B(n5015), .Z(n5020) );
  OR U5203 ( .A(n5018), .B(n5017), .Z(n5019) );
  NAND U5204 ( .A(n5020), .B(n5019), .Z(n5157) );
  NANDN U5205 ( .A(n5022), .B(n5021), .Z(n5026) );
  OR U5206 ( .A(n5024), .B(n5023), .Z(n5025) );
  NAND U5207 ( .A(n5026), .B(n5025), .Z(n5145) );
  NAND U5208 ( .A(b[0]), .B(a[72]), .Z(n5027) );
  XNOR U5209 ( .A(b[1]), .B(n5027), .Z(n5029) );
  NAND U5210 ( .A(a[71]), .B(n72), .Z(n5028) );
  AND U5211 ( .A(n5029), .B(n5028), .Z(n5121) );
  XNOR U5212 ( .A(n10050), .B(n5180), .Z(n5130) );
  OR U5213 ( .A(n5130), .B(n10051), .Z(n5032) );
  NANDN U5214 ( .A(n5030), .B(n10070), .Z(n5031) );
  AND U5215 ( .A(n5032), .B(n5031), .Z(n5122) );
  XOR U5216 ( .A(n5121), .B(n5122), .Z(n5124) );
  NAND U5217 ( .A(a[56]), .B(b[15]), .Z(n5123) );
  XOR U5218 ( .A(n5124), .B(n5123), .Z(n5142) );
  XNOR U5219 ( .A(n9622), .B(n5804), .Z(n5133) );
  OR U5220 ( .A(n5133), .B(n9623), .Z(n5035) );
  NANDN U5221 ( .A(n5033), .B(n9680), .Z(n5034) );
  NAND U5222 ( .A(n5035), .B(n5034), .Z(n5118) );
  XNOR U5223 ( .A(n9872), .B(n5675), .Z(n5136) );
  NANDN U5224 ( .A(n5136), .B(n9746), .Z(n5038) );
  NANDN U5225 ( .A(n5036), .B(n9747), .Z(n5037) );
  NAND U5226 ( .A(n5038), .B(n5037), .Z(n5115) );
  IV U5227 ( .A(a[70]), .Z(n5960) );
  XNOR U5228 ( .A(n74), .B(n5960), .Z(n5139) );
  NANDN U5229 ( .A(n5139), .B(n9485), .Z(n5041) );
  NANDN U5230 ( .A(n5039), .B(n9484), .Z(n5040) );
  AND U5231 ( .A(n5041), .B(n5040), .Z(n5116) );
  XNOR U5232 ( .A(n5115), .B(n5116), .Z(n5117) );
  XOR U5233 ( .A(n5118), .B(n5117), .Z(n5143) );
  XOR U5234 ( .A(n5142), .B(n5143), .Z(n5144) );
  XNOR U5235 ( .A(n5145), .B(n5144), .Z(n5093) );
  NAND U5236 ( .A(n5043), .B(n5042), .Z(n5047) );
  NAND U5237 ( .A(n5045), .B(n5044), .Z(n5046) );
  NAND U5238 ( .A(n5047), .B(n5046), .Z(n5094) );
  XOR U5239 ( .A(n5093), .B(n5094), .Z(n5096) );
  XNOR U5240 ( .A(n9967), .B(n5336), .Z(n5099) );
  OR U5241 ( .A(n5099), .B(n10020), .Z(n5050) );
  NANDN U5242 ( .A(n5048), .B(n9968), .Z(n5049) );
  NAND U5243 ( .A(n5050), .B(n5049), .Z(n5112) );
  XNOR U5244 ( .A(n75), .B(n5051), .Z(n5103) );
  OR U5245 ( .A(n5103), .B(n10106), .Z(n5054) );
  NANDN U5246 ( .A(n5052), .B(n10107), .Z(n5053) );
  NAND U5247 ( .A(n5054), .B(n5053), .Z(n5109) );
  XNOR U5248 ( .A(n9984), .B(n5492), .Z(n5106) );
  NANDN U5249 ( .A(n5106), .B(n9865), .Z(n5057) );
  NANDN U5250 ( .A(n5055), .B(n9930), .Z(n5056) );
  AND U5251 ( .A(n5057), .B(n5056), .Z(n5110) );
  XNOR U5252 ( .A(n5109), .B(n5110), .Z(n5111) );
  XNOR U5253 ( .A(n5112), .B(n5111), .Z(n5148) );
  NANDN U5254 ( .A(n5059), .B(n5058), .Z(n5063) );
  NAND U5255 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U5256 ( .A(n5063), .B(n5062), .Z(n5149) );
  XNOR U5257 ( .A(n5148), .B(n5149), .Z(n5150) );
  NANDN U5258 ( .A(n5065), .B(n5064), .Z(n5069) );
  NAND U5259 ( .A(n5067), .B(n5066), .Z(n5068) );
  AND U5260 ( .A(n5069), .B(n5068), .Z(n5151) );
  XNOR U5261 ( .A(n5150), .B(n5151), .Z(n5095) );
  XNOR U5262 ( .A(n5096), .B(n5095), .Z(n5154) );
  NANDN U5263 ( .A(n5071), .B(n5070), .Z(n5075) );
  NAND U5264 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U5265 ( .A(n5075), .B(n5074), .Z(n5155) );
  XNOR U5266 ( .A(n5154), .B(n5155), .Z(n5156) );
  XOR U5267 ( .A(n5157), .B(n5156), .Z(n5087) );
  NANDN U5268 ( .A(n5077), .B(n5076), .Z(n5081) );
  NANDN U5269 ( .A(n5079), .B(n5078), .Z(n5080) );
  NAND U5270 ( .A(n5081), .B(n5080), .Z(n5088) );
  XNOR U5271 ( .A(n5087), .B(n5088), .Z(n5089) );
  XNOR U5272 ( .A(n5090), .B(n5089), .Z(n5160) );
  XNOR U5273 ( .A(n5160), .B(sreg[184]), .Z(n5162) );
  NAND U5274 ( .A(n5082), .B(sreg[183]), .Z(n5086) );
  OR U5275 ( .A(n5084), .B(n5083), .Z(n5085) );
  AND U5276 ( .A(n5086), .B(n5085), .Z(n5161) );
  XOR U5277 ( .A(n5162), .B(n5161), .Z(c[184]) );
  NANDN U5278 ( .A(n5088), .B(n5087), .Z(n5092) );
  NAND U5279 ( .A(n5090), .B(n5089), .Z(n5091) );
  NAND U5280 ( .A(n5092), .B(n5091), .Z(n5168) );
  NANDN U5281 ( .A(n5094), .B(n5093), .Z(n5098) );
  OR U5282 ( .A(n5096), .B(n5095), .Z(n5097) );
  NAND U5283 ( .A(n5098), .B(n5097), .Z(n5235) );
  XNOR U5284 ( .A(n9967), .B(n5414), .Z(n5177) );
  OR U5285 ( .A(n5177), .B(n10020), .Z(n5101) );
  NANDN U5286 ( .A(n5099), .B(n9968), .Z(n5100) );
  NAND U5287 ( .A(n5101), .B(n5100), .Z(n5190) );
  XNOR U5288 ( .A(n75), .B(n5102), .Z(n5181) );
  OR U5289 ( .A(n5181), .B(n10106), .Z(n5105) );
  NANDN U5290 ( .A(n5103), .B(n10107), .Z(n5104) );
  NAND U5291 ( .A(n5105), .B(n5104), .Z(n5187) );
  XNOR U5292 ( .A(n9984), .B(n5570), .Z(n5184) );
  NANDN U5293 ( .A(n5184), .B(n9865), .Z(n5108) );
  NANDN U5294 ( .A(n5106), .B(n9930), .Z(n5107) );
  AND U5295 ( .A(n5108), .B(n5107), .Z(n5188) );
  XNOR U5296 ( .A(n5187), .B(n5188), .Z(n5189) );
  XNOR U5297 ( .A(n5190), .B(n5189), .Z(n5226) );
  NANDN U5298 ( .A(n5110), .B(n5109), .Z(n5114) );
  NAND U5299 ( .A(n5112), .B(n5111), .Z(n5113) );
  NAND U5300 ( .A(n5114), .B(n5113), .Z(n5227) );
  XNOR U5301 ( .A(n5226), .B(n5227), .Z(n5228) );
  NANDN U5302 ( .A(n5116), .B(n5115), .Z(n5120) );
  NAND U5303 ( .A(n5118), .B(n5117), .Z(n5119) );
  AND U5304 ( .A(n5120), .B(n5119), .Z(n5229) );
  XNOR U5305 ( .A(n5228), .B(n5229), .Z(n5173) );
  NANDN U5306 ( .A(n5122), .B(n5121), .Z(n5126) );
  OR U5307 ( .A(n5124), .B(n5123), .Z(n5125) );
  NAND U5308 ( .A(n5126), .B(n5125), .Z(n5223) );
  NAND U5309 ( .A(b[0]), .B(a[73]), .Z(n5127) );
  XNOR U5310 ( .A(b[1]), .B(n5127), .Z(n5129) );
  NAND U5311 ( .A(a[72]), .B(n72), .Z(n5128) );
  AND U5312 ( .A(n5129), .B(n5128), .Z(n5199) );
  XNOR U5313 ( .A(n10050), .B(n5258), .Z(n5208) );
  OR U5314 ( .A(n5208), .B(n10051), .Z(n5132) );
  NANDN U5315 ( .A(n5130), .B(n10070), .Z(n5131) );
  AND U5316 ( .A(n5132), .B(n5131), .Z(n5200) );
  XOR U5317 ( .A(n5199), .B(n5200), .Z(n5202) );
  NAND U5318 ( .A(a[57]), .B(b[15]), .Z(n5201) );
  XOR U5319 ( .A(n5202), .B(n5201), .Z(n5220) );
  XNOR U5320 ( .A(n9622), .B(n5882), .Z(n5211) );
  OR U5321 ( .A(n5211), .B(n9623), .Z(n5135) );
  NANDN U5322 ( .A(n5133), .B(n9680), .Z(n5134) );
  NAND U5323 ( .A(n5135), .B(n5134), .Z(n5196) );
  XNOR U5324 ( .A(n9872), .B(n5726), .Z(n5214) );
  NANDN U5325 ( .A(n5214), .B(n9746), .Z(n5138) );
  NANDN U5326 ( .A(n5136), .B(n9747), .Z(n5137) );
  NAND U5327 ( .A(n5138), .B(n5137), .Z(n5193) );
  IV U5328 ( .A(a[71]), .Z(n6038) );
  XNOR U5329 ( .A(n74), .B(n6038), .Z(n5217) );
  NANDN U5330 ( .A(n5217), .B(n9485), .Z(n5141) );
  NANDN U5331 ( .A(n5139), .B(n9484), .Z(n5140) );
  AND U5332 ( .A(n5141), .B(n5140), .Z(n5194) );
  XNOR U5333 ( .A(n5193), .B(n5194), .Z(n5195) );
  XOR U5334 ( .A(n5196), .B(n5195), .Z(n5221) );
  XOR U5335 ( .A(n5220), .B(n5221), .Z(n5222) );
  XNOR U5336 ( .A(n5223), .B(n5222), .Z(n5171) );
  NAND U5337 ( .A(n5143), .B(n5142), .Z(n5147) );
  NAND U5338 ( .A(n5145), .B(n5144), .Z(n5146) );
  NAND U5339 ( .A(n5147), .B(n5146), .Z(n5172) );
  XOR U5340 ( .A(n5171), .B(n5172), .Z(n5174) );
  XNOR U5341 ( .A(n5173), .B(n5174), .Z(n5232) );
  NANDN U5342 ( .A(n5149), .B(n5148), .Z(n5153) );
  NAND U5343 ( .A(n5151), .B(n5150), .Z(n5152) );
  NAND U5344 ( .A(n5153), .B(n5152), .Z(n5233) );
  XNOR U5345 ( .A(n5232), .B(n5233), .Z(n5234) );
  XOR U5346 ( .A(n5235), .B(n5234), .Z(n5165) );
  NANDN U5347 ( .A(n5155), .B(n5154), .Z(n5159) );
  NANDN U5348 ( .A(n5157), .B(n5156), .Z(n5158) );
  NAND U5349 ( .A(n5159), .B(n5158), .Z(n5166) );
  XNOR U5350 ( .A(n5165), .B(n5166), .Z(n5167) );
  XNOR U5351 ( .A(n5168), .B(n5167), .Z(n5238) );
  XNOR U5352 ( .A(n5238), .B(sreg[185]), .Z(n5240) );
  NAND U5353 ( .A(n5160), .B(sreg[184]), .Z(n5164) );
  OR U5354 ( .A(n5162), .B(n5161), .Z(n5163) );
  AND U5355 ( .A(n5164), .B(n5163), .Z(n5239) );
  XOR U5356 ( .A(n5240), .B(n5239), .Z(c[185]) );
  NANDN U5357 ( .A(n5166), .B(n5165), .Z(n5170) );
  NAND U5358 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U5359 ( .A(n5170), .B(n5169), .Z(n5246) );
  NANDN U5360 ( .A(n5172), .B(n5171), .Z(n5176) );
  OR U5361 ( .A(n5174), .B(n5173), .Z(n5175) );
  NAND U5362 ( .A(n5176), .B(n5175), .Z(n5313) );
  XNOR U5363 ( .A(n9967), .B(n5492), .Z(n5255) );
  OR U5364 ( .A(n5255), .B(n10020), .Z(n5179) );
  NANDN U5365 ( .A(n5177), .B(n9968), .Z(n5178) );
  NAND U5366 ( .A(n5179), .B(n5178), .Z(n5268) );
  XNOR U5367 ( .A(n75), .B(n5180), .Z(n5259) );
  OR U5368 ( .A(n5259), .B(n10106), .Z(n5183) );
  NANDN U5369 ( .A(n5181), .B(n10107), .Z(n5182) );
  NAND U5370 ( .A(n5183), .B(n5182), .Z(n5265) );
  XNOR U5371 ( .A(n9984), .B(n5675), .Z(n5262) );
  NANDN U5372 ( .A(n5262), .B(n9865), .Z(n5186) );
  NANDN U5373 ( .A(n5184), .B(n9930), .Z(n5185) );
  AND U5374 ( .A(n5186), .B(n5185), .Z(n5266) );
  XNOR U5375 ( .A(n5265), .B(n5266), .Z(n5267) );
  XNOR U5376 ( .A(n5268), .B(n5267), .Z(n5304) );
  NANDN U5377 ( .A(n5188), .B(n5187), .Z(n5192) );
  NAND U5378 ( .A(n5190), .B(n5189), .Z(n5191) );
  NAND U5379 ( .A(n5192), .B(n5191), .Z(n5305) );
  XNOR U5380 ( .A(n5304), .B(n5305), .Z(n5306) );
  NANDN U5381 ( .A(n5194), .B(n5193), .Z(n5198) );
  NAND U5382 ( .A(n5196), .B(n5195), .Z(n5197) );
  AND U5383 ( .A(n5198), .B(n5197), .Z(n5307) );
  XNOR U5384 ( .A(n5306), .B(n5307), .Z(n5251) );
  NANDN U5385 ( .A(n5200), .B(n5199), .Z(n5204) );
  OR U5386 ( .A(n5202), .B(n5201), .Z(n5203) );
  NAND U5387 ( .A(n5204), .B(n5203), .Z(n5301) );
  NAND U5388 ( .A(b[0]), .B(a[74]), .Z(n5205) );
  XNOR U5389 ( .A(b[1]), .B(n5205), .Z(n5207) );
  NAND U5390 ( .A(a[73]), .B(n72), .Z(n5206) );
  AND U5391 ( .A(n5207), .B(n5206), .Z(n5277) );
  XNOR U5392 ( .A(n10050), .B(n5336), .Z(n5286) );
  OR U5393 ( .A(n5286), .B(n10051), .Z(n5210) );
  NANDN U5394 ( .A(n5208), .B(n10070), .Z(n5209) );
  AND U5395 ( .A(n5210), .B(n5209), .Z(n5278) );
  XOR U5396 ( .A(n5277), .B(n5278), .Z(n5280) );
  NAND U5397 ( .A(a[58]), .B(b[15]), .Z(n5279) );
  XOR U5398 ( .A(n5280), .B(n5279), .Z(n5298) );
  XNOR U5399 ( .A(n9622), .B(n5960), .Z(n5289) );
  OR U5400 ( .A(n5289), .B(n9623), .Z(n5213) );
  NANDN U5401 ( .A(n5211), .B(n9680), .Z(n5212) );
  NAND U5402 ( .A(n5213), .B(n5212), .Z(n5274) );
  XNOR U5403 ( .A(n9872), .B(n5804), .Z(n5292) );
  NANDN U5404 ( .A(n5292), .B(n9746), .Z(n5216) );
  NANDN U5405 ( .A(n5214), .B(n9747), .Z(n5215) );
  NAND U5406 ( .A(n5216), .B(n5215), .Z(n5271) );
  IV U5407 ( .A(a[72]), .Z(n6143) );
  XNOR U5408 ( .A(n74), .B(n6143), .Z(n5295) );
  NANDN U5409 ( .A(n5295), .B(n9485), .Z(n5219) );
  NANDN U5410 ( .A(n5217), .B(n9484), .Z(n5218) );
  AND U5411 ( .A(n5219), .B(n5218), .Z(n5272) );
  XNOR U5412 ( .A(n5271), .B(n5272), .Z(n5273) );
  XOR U5413 ( .A(n5274), .B(n5273), .Z(n5299) );
  XOR U5414 ( .A(n5298), .B(n5299), .Z(n5300) );
  XNOR U5415 ( .A(n5301), .B(n5300), .Z(n5249) );
  NAND U5416 ( .A(n5221), .B(n5220), .Z(n5225) );
  NAND U5417 ( .A(n5223), .B(n5222), .Z(n5224) );
  NAND U5418 ( .A(n5225), .B(n5224), .Z(n5250) );
  XOR U5419 ( .A(n5249), .B(n5250), .Z(n5252) );
  XNOR U5420 ( .A(n5251), .B(n5252), .Z(n5310) );
  NANDN U5421 ( .A(n5227), .B(n5226), .Z(n5231) );
  NAND U5422 ( .A(n5229), .B(n5228), .Z(n5230) );
  NAND U5423 ( .A(n5231), .B(n5230), .Z(n5311) );
  XNOR U5424 ( .A(n5310), .B(n5311), .Z(n5312) );
  XOR U5425 ( .A(n5313), .B(n5312), .Z(n5243) );
  NANDN U5426 ( .A(n5233), .B(n5232), .Z(n5237) );
  NANDN U5427 ( .A(n5235), .B(n5234), .Z(n5236) );
  NAND U5428 ( .A(n5237), .B(n5236), .Z(n5244) );
  XNOR U5429 ( .A(n5243), .B(n5244), .Z(n5245) );
  XNOR U5430 ( .A(n5246), .B(n5245), .Z(n5316) );
  XNOR U5431 ( .A(n5316), .B(sreg[186]), .Z(n5318) );
  NAND U5432 ( .A(n5238), .B(sreg[185]), .Z(n5242) );
  OR U5433 ( .A(n5240), .B(n5239), .Z(n5241) );
  AND U5434 ( .A(n5242), .B(n5241), .Z(n5317) );
  XOR U5435 ( .A(n5318), .B(n5317), .Z(c[186]) );
  NANDN U5436 ( .A(n5244), .B(n5243), .Z(n5248) );
  NAND U5437 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U5438 ( .A(n5248), .B(n5247), .Z(n5324) );
  NANDN U5439 ( .A(n5250), .B(n5249), .Z(n5254) );
  OR U5440 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U5441 ( .A(n5254), .B(n5253), .Z(n5391) );
  XNOR U5442 ( .A(n9967), .B(n5570), .Z(n5333) );
  OR U5443 ( .A(n5333), .B(n10020), .Z(n5257) );
  NANDN U5444 ( .A(n5255), .B(n9968), .Z(n5256) );
  NAND U5445 ( .A(n5257), .B(n5256), .Z(n5346) );
  XNOR U5446 ( .A(n75), .B(n5258), .Z(n5337) );
  OR U5447 ( .A(n5337), .B(n10106), .Z(n5261) );
  NANDN U5448 ( .A(n5259), .B(n10107), .Z(n5260) );
  NAND U5449 ( .A(n5261), .B(n5260), .Z(n5343) );
  XNOR U5450 ( .A(n9984), .B(n5726), .Z(n5340) );
  NANDN U5451 ( .A(n5340), .B(n9865), .Z(n5264) );
  NANDN U5452 ( .A(n5262), .B(n9930), .Z(n5263) );
  AND U5453 ( .A(n5264), .B(n5263), .Z(n5344) );
  XNOR U5454 ( .A(n5343), .B(n5344), .Z(n5345) );
  XNOR U5455 ( .A(n5346), .B(n5345), .Z(n5382) );
  NANDN U5456 ( .A(n5266), .B(n5265), .Z(n5270) );
  NAND U5457 ( .A(n5268), .B(n5267), .Z(n5269) );
  NAND U5458 ( .A(n5270), .B(n5269), .Z(n5383) );
  XNOR U5459 ( .A(n5382), .B(n5383), .Z(n5384) );
  NANDN U5460 ( .A(n5272), .B(n5271), .Z(n5276) );
  NAND U5461 ( .A(n5274), .B(n5273), .Z(n5275) );
  AND U5462 ( .A(n5276), .B(n5275), .Z(n5385) );
  XNOR U5463 ( .A(n5384), .B(n5385), .Z(n5329) );
  NANDN U5464 ( .A(n5278), .B(n5277), .Z(n5282) );
  OR U5465 ( .A(n5280), .B(n5279), .Z(n5281) );
  NAND U5466 ( .A(n5282), .B(n5281), .Z(n5379) );
  NAND U5467 ( .A(b[0]), .B(a[75]), .Z(n5283) );
  XNOR U5468 ( .A(b[1]), .B(n5283), .Z(n5285) );
  NAND U5469 ( .A(a[74]), .B(n72), .Z(n5284) );
  AND U5470 ( .A(n5285), .B(n5284), .Z(n5355) );
  XNOR U5471 ( .A(n10050), .B(n5414), .Z(n5364) );
  OR U5472 ( .A(n5364), .B(n10051), .Z(n5288) );
  NANDN U5473 ( .A(n5286), .B(n10070), .Z(n5287) );
  AND U5474 ( .A(n5288), .B(n5287), .Z(n5356) );
  XOR U5475 ( .A(n5355), .B(n5356), .Z(n5358) );
  NAND U5476 ( .A(a[59]), .B(b[15]), .Z(n5357) );
  XOR U5477 ( .A(n5358), .B(n5357), .Z(n5376) );
  XNOR U5478 ( .A(n9622), .B(n6038), .Z(n5367) );
  OR U5479 ( .A(n5367), .B(n9623), .Z(n5291) );
  NANDN U5480 ( .A(n5289), .B(n9680), .Z(n5290) );
  NAND U5481 ( .A(n5291), .B(n5290), .Z(n5352) );
  XNOR U5482 ( .A(n9872), .B(n5882), .Z(n5370) );
  NANDN U5483 ( .A(n5370), .B(n9746), .Z(n5294) );
  NANDN U5484 ( .A(n5292), .B(n9747), .Z(n5293) );
  NAND U5485 ( .A(n5294), .B(n5293), .Z(n5349) );
  IV U5486 ( .A(a[73]), .Z(n6194) );
  XNOR U5487 ( .A(n74), .B(n6194), .Z(n5373) );
  NANDN U5488 ( .A(n5373), .B(n9485), .Z(n5297) );
  NANDN U5489 ( .A(n5295), .B(n9484), .Z(n5296) );
  AND U5490 ( .A(n5297), .B(n5296), .Z(n5350) );
  XNOR U5491 ( .A(n5349), .B(n5350), .Z(n5351) );
  XOR U5492 ( .A(n5352), .B(n5351), .Z(n5377) );
  XOR U5493 ( .A(n5376), .B(n5377), .Z(n5378) );
  XNOR U5494 ( .A(n5379), .B(n5378), .Z(n5327) );
  NAND U5495 ( .A(n5299), .B(n5298), .Z(n5303) );
  NAND U5496 ( .A(n5301), .B(n5300), .Z(n5302) );
  NAND U5497 ( .A(n5303), .B(n5302), .Z(n5328) );
  XOR U5498 ( .A(n5327), .B(n5328), .Z(n5330) );
  XNOR U5499 ( .A(n5329), .B(n5330), .Z(n5388) );
  NANDN U5500 ( .A(n5305), .B(n5304), .Z(n5309) );
  NAND U5501 ( .A(n5307), .B(n5306), .Z(n5308) );
  NAND U5502 ( .A(n5309), .B(n5308), .Z(n5389) );
  XNOR U5503 ( .A(n5388), .B(n5389), .Z(n5390) );
  XOR U5504 ( .A(n5391), .B(n5390), .Z(n5321) );
  NANDN U5505 ( .A(n5311), .B(n5310), .Z(n5315) );
  NANDN U5506 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U5507 ( .A(n5315), .B(n5314), .Z(n5322) );
  XNOR U5508 ( .A(n5321), .B(n5322), .Z(n5323) );
  XNOR U5509 ( .A(n5324), .B(n5323), .Z(n5394) );
  XNOR U5510 ( .A(n5394), .B(sreg[187]), .Z(n5396) );
  NAND U5511 ( .A(n5316), .B(sreg[186]), .Z(n5320) );
  OR U5512 ( .A(n5318), .B(n5317), .Z(n5319) );
  AND U5513 ( .A(n5320), .B(n5319), .Z(n5395) );
  XOR U5514 ( .A(n5396), .B(n5395), .Z(c[187]) );
  NANDN U5515 ( .A(n5322), .B(n5321), .Z(n5326) );
  NAND U5516 ( .A(n5324), .B(n5323), .Z(n5325) );
  NAND U5517 ( .A(n5326), .B(n5325), .Z(n5402) );
  NANDN U5518 ( .A(n5328), .B(n5327), .Z(n5332) );
  OR U5519 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U5520 ( .A(n5332), .B(n5331), .Z(n5469) );
  XNOR U5521 ( .A(n9967), .B(n5675), .Z(n5411) );
  OR U5522 ( .A(n5411), .B(n10020), .Z(n5335) );
  NANDN U5523 ( .A(n5333), .B(n9968), .Z(n5334) );
  NAND U5524 ( .A(n5335), .B(n5334), .Z(n5424) );
  XNOR U5525 ( .A(n75), .B(n5336), .Z(n5415) );
  OR U5526 ( .A(n5415), .B(n10106), .Z(n5339) );
  NANDN U5527 ( .A(n5337), .B(n10107), .Z(n5338) );
  NAND U5528 ( .A(n5339), .B(n5338), .Z(n5421) );
  XNOR U5529 ( .A(n9984), .B(n5804), .Z(n5418) );
  NANDN U5530 ( .A(n5418), .B(n9865), .Z(n5342) );
  NANDN U5531 ( .A(n5340), .B(n9930), .Z(n5341) );
  AND U5532 ( .A(n5342), .B(n5341), .Z(n5422) );
  XNOR U5533 ( .A(n5421), .B(n5422), .Z(n5423) );
  XNOR U5534 ( .A(n5424), .B(n5423), .Z(n5460) );
  NANDN U5535 ( .A(n5344), .B(n5343), .Z(n5348) );
  NAND U5536 ( .A(n5346), .B(n5345), .Z(n5347) );
  NAND U5537 ( .A(n5348), .B(n5347), .Z(n5461) );
  XNOR U5538 ( .A(n5460), .B(n5461), .Z(n5462) );
  NANDN U5539 ( .A(n5350), .B(n5349), .Z(n5354) );
  NAND U5540 ( .A(n5352), .B(n5351), .Z(n5353) );
  AND U5541 ( .A(n5354), .B(n5353), .Z(n5463) );
  XNOR U5542 ( .A(n5462), .B(n5463), .Z(n5407) );
  NANDN U5543 ( .A(n5356), .B(n5355), .Z(n5360) );
  OR U5544 ( .A(n5358), .B(n5357), .Z(n5359) );
  NAND U5545 ( .A(n5360), .B(n5359), .Z(n5457) );
  NAND U5546 ( .A(b[0]), .B(a[76]), .Z(n5361) );
  XNOR U5547 ( .A(b[1]), .B(n5361), .Z(n5363) );
  NAND U5548 ( .A(a[75]), .B(n72), .Z(n5362) );
  AND U5549 ( .A(n5363), .B(n5362), .Z(n5433) );
  XNOR U5550 ( .A(n10050), .B(n5492), .Z(n5442) );
  OR U5551 ( .A(n5442), .B(n10051), .Z(n5366) );
  NANDN U5552 ( .A(n5364), .B(n10070), .Z(n5365) );
  AND U5553 ( .A(n5366), .B(n5365), .Z(n5434) );
  XOR U5554 ( .A(n5433), .B(n5434), .Z(n5436) );
  NAND U5555 ( .A(a[60]), .B(b[15]), .Z(n5435) );
  XOR U5556 ( .A(n5436), .B(n5435), .Z(n5454) );
  XNOR U5557 ( .A(n9622), .B(n6143), .Z(n5445) );
  OR U5558 ( .A(n5445), .B(n9623), .Z(n5369) );
  NANDN U5559 ( .A(n5367), .B(n9680), .Z(n5368) );
  NAND U5560 ( .A(n5369), .B(n5368), .Z(n5430) );
  XNOR U5561 ( .A(n9872), .B(n5960), .Z(n5448) );
  NANDN U5562 ( .A(n5448), .B(n9746), .Z(n5372) );
  NANDN U5563 ( .A(n5370), .B(n9747), .Z(n5371) );
  NAND U5564 ( .A(n5372), .B(n5371), .Z(n5427) );
  IV U5565 ( .A(a[74]), .Z(n6272) );
  XNOR U5566 ( .A(n74), .B(n6272), .Z(n5451) );
  NANDN U5567 ( .A(n5451), .B(n9485), .Z(n5375) );
  NANDN U5568 ( .A(n5373), .B(n9484), .Z(n5374) );
  AND U5569 ( .A(n5375), .B(n5374), .Z(n5428) );
  XNOR U5570 ( .A(n5427), .B(n5428), .Z(n5429) );
  XOR U5571 ( .A(n5430), .B(n5429), .Z(n5455) );
  XOR U5572 ( .A(n5454), .B(n5455), .Z(n5456) );
  XNOR U5573 ( .A(n5457), .B(n5456), .Z(n5405) );
  NAND U5574 ( .A(n5377), .B(n5376), .Z(n5381) );
  NAND U5575 ( .A(n5379), .B(n5378), .Z(n5380) );
  NAND U5576 ( .A(n5381), .B(n5380), .Z(n5406) );
  XOR U5577 ( .A(n5405), .B(n5406), .Z(n5408) );
  XNOR U5578 ( .A(n5407), .B(n5408), .Z(n5466) );
  NANDN U5579 ( .A(n5383), .B(n5382), .Z(n5387) );
  NAND U5580 ( .A(n5385), .B(n5384), .Z(n5386) );
  NAND U5581 ( .A(n5387), .B(n5386), .Z(n5467) );
  XNOR U5582 ( .A(n5466), .B(n5467), .Z(n5468) );
  XOR U5583 ( .A(n5469), .B(n5468), .Z(n5399) );
  NANDN U5584 ( .A(n5389), .B(n5388), .Z(n5393) );
  NANDN U5585 ( .A(n5391), .B(n5390), .Z(n5392) );
  NAND U5586 ( .A(n5393), .B(n5392), .Z(n5400) );
  XNOR U5587 ( .A(n5399), .B(n5400), .Z(n5401) );
  XNOR U5588 ( .A(n5402), .B(n5401), .Z(n5472) );
  XNOR U5589 ( .A(n5472), .B(sreg[188]), .Z(n5474) );
  NAND U5590 ( .A(n5394), .B(sreg[187]), .Z(n5398) );
  OR U5591 ( .A(n5396), .B(n5395), .Z(n5397) );
  AND U5592 ( .A(n5398), .B(n5397), .Z(n5473) );
  XOR U5593 ( .A(n5474), .B(n5473), .Z(c[188]) );
  NANDN U5594 ( .A(n5400), .B(n5399), .Z(n5404) );
  NAND U5595 ( .A(n5402), .B(n5401), .Z(n5403) );
  NAND U5596 ( .A(n5404), .B(n5403), .Z(n5480) );
  NANDN U5597 ( .A(n5406), .B(n5405), .Z(n5410) );
  OR U5598 ( .A(n5408), .B(n5407), .Z(n5409) );
  NAND U5599 ( .A(n5410), .B(n5409), .Z(n5547) );
  XNOR U5600 ( .A(n9967), .B(n5726), .Z(n5489) );
  OR U5601 ( .A(n5489), .B(n10020), .Z(n5413) );
  NANDN U5602 ( .A(n5411), .B(n9968), .Z(n5412) );
  NAND U5603 ( .A(n5413), .B(n5412), .Z(n5502) );
  XNOR U5604 ( .A(n75), .B(n5414), .Z(n5493) );
  OR U5605 ( .A(n5493), .B(n10106), .Z(n5417) );
  NANDN U5606 ( .A(n5415), .B(n10107), .Z(n5416) );
  NAND U5607 ( .A(n5417), .B(n5416), .Z(n5499) );
  XNOR U5608 ( .A(n9984), .B(n5882), .Z(n5496) );
  NANDN U5609 ( .A(n5496), .B(n9865), .Z(n5420) );
  NANDN U5610 ( .A(n5418), .B(n9930), .Z(n5419) );
  AND U5611 ( .A(n5420), .B(n5419), .Z(n5500) );
  XNOR U5612 ( .A(n5499), .B(n5500), .Z(n5501) );
  XNOR U5613 ( .A(n5502), .B(n5501), .Z(n5538) );
  NANDN U5614 ( .A(n5422), .B(n5421), .Z(n5426) );
  NAND U5615 ( .A(n5424), .B(n5423), .Z(n5425) );
  NAND U5616 ( .A(n5426), .B(n5425), .Z(n5539) );
  XNOR U5617 ( .A(n5538), .B(n5539), .Z(n5540) );
  NANDN U5618 ( .A(n5428), .B(n5427), .Z(n5432) );
  NAND U5619 ( .A(n5430), .B(n5429), .Z(n5431) );
  AND U5620 ( .A(n5432), .B(n5431), .Z(n5541) );
  XNOR U5621 ( .A(n5540), .B(n5541), .Z(n5485) );
  NANDN U5622 ( .A(n5434), .B(n5433), .Z(n5438) );
  OR U5623 ( .A(n5436), .B(n5435), .Z(n5437) );
  NAND U5624 ( .A(n5438), .B(n5437), .Z(n5535) );
  NAND U5625 ( .A(b[0]), .B(a[77]), .Z(n5439) );
  XNOR U5626 ( .A(b[1]), .B(n5439), .Z(n5441) );
  NAND U5627 ( .A(a[76]), .B(n72), .Z(n5440) );
  AND U5628 ( .A(n5441), .B(n5440), .Z(n5511) );
  XNOR U5629 ( .A(n10050), .B(n5570), .Z(n5517) );
  OR U5630 ( .A(n5517), .B(n10051), .Z(n5444) );
  NANDN U5631 ( .A(n5442), .B(n10070), .Z(n5443) );
  AND U5632 ( .A(n5444), .B(n5443), .Z(n5512) );
  XOR U5633 ( .A(n5511), .B(n5512), .Z(n5514) );
  NAND U5634 ( .A(a[61]), .B(b[15]), .Z(n5513) );
  XOR U5635 ( .A(n5514), .B(n5513), .Z(n5532) );
  XNOR U5636 ( .A(n9622), .B(n6194), .Z(n5523) );
  OR U5637 ( .A(n5523), .B(n9623), .Z(n5447) );
  NANDN U5638 ( .A(n5445), .B(n9680), .Z(n5446) );
  NAND U5639 ( .A(n5447), .B(n5446), .Z(n5508) );
  XNOR U5640 ( .A(n9872), .B(n6038), .Z(n5526) );
  NANDN U5641 ( .A(n5526), .B(n9746), .Z(n5450) );
  NANDN U5642 ( .A(n5448), .B(n9747), .Z(n5449) );
  NAND U5643 ( .A(n5450), .B(n5449), .Z(n5505) );
  IV U5644 ( .A(a[75]), .Z(n6377) );
  XNOR U5645 ( .A(n74), .B(n6377), .Z(n5529) );
  NANDN U5646 ( .A(n5529), .B(n9485), .Z(n5453) );
  NANDN U5647 ( .A(n5451), .B(n9484), .Z(n5452) );
  AND U5648 ( .A(n5453), .B(n5452), .Z(n5506) );
  XNOR U5649 ( .A(n5505), .B(n5506), .Z(n5507) );
  XOR U5650 ( .A(n5508), .B(n5507), .Z(n5533) );
  XOR U5651 ( .A(n5532), .B(n5533), .Z(n5534) );
  XNOR U5652 ( .A(n5535), .B(n5534), .Z(n5483) );
  NAND U5653 ( .A(n5455), .B(n5454), .Z(n5459) );
  NAND U5654 ( .A(n5457), .B(n5456), .Z(n5458) );
  NAND U5655 ( .A(n5459), .B(n5458), .Z(n5484) );
  XOR U5656 ( .A(n5483), .B(n5484), .Z(n5486) );
  XNOR U5657 ( .A(n5485), .B(n5486), .Z(n5544) );
  NANDN U5658 ( .A(n5461), .B(n5460), .Z(n5465) );
  NAND U5659 ( .A(n5463), .B(n5462), .Z(n5464) );
  NAND U5660 ( .A(n5465), .B(n5464), .Z(n5545) );
  XNOR U5661 ( .A(n5544), .B(n5545), .Z(n5546) );
  XOR U5662 ( .A(n5547), .B(n5546), .Z(n5477) );
  NANDN U5663 ( .A(n5467), .B(n5466), .Z(n5471) );
  NANDN U5664 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U5665 ( .A(n5471), .B(n5470), .Z(n5478) );
  XNOR U5666 ( .A(n5477), .B(n5478), .Z(n5479) );
  XNOR U5667 ( .A(n5480), .B(n5479), .Z(n5550) );
  XNOR U5668 ( .A(n5550), .B(sreg[189]), .Z(n5552) );
  NAND U5669 ( .A(n5472), .B(sreg[188]), .Z(n5476) );
  OR U5670 ( .A(n5474), .B(n5473), .Z(n5475) );
  AND U5671 ( .A(n5476), .B(n5475), .Z(n5551) );
  XOR U5672 ( .A(n5552), .B(n5551), .Z(c[189]) );
  NANDN U5673 ( .A(n5478), .B(n5477), .Z(n5482) );
  NAND U5674 ( .A(n5480), .B(n5479), .Z(n5481) );
  NAND U5675 ( .A(n5482), .B(n5481), .Z(n5558) );
  NANDN U5676 ( .A(n5484), .B(n5483), .Z(n5488) );
  OR U5677 ( .A(n5486), .B(n5485), .Z(n5487) );
  NAND U5678 ( .A(n5488), .B(n5487), .Z(n5625) );
  XNOR U5679 ( .A(n9967), .B(n5804), .Z(n5567) );
  OR U5680 ( .A(n5567), .B(n10020), .Z(n5491) );
  NANDN U5681 ( .A(n5489), .B(n9968), .Z(n5490) );
  NAND U5682 ( .A(n5491), .B(n5490), .Z(n5580) );
  XNOR U5683 ( .A(n75), .B(n5492), .Z(n5571) );
  OR U5684 ( .A(n5571), .B(n10106), .Z(n5495) );
  NANDN U5685 ( .A(n5493), .B(n10107), .Z(n5494) );
  NAND U5686 ( .A(n5495), .B(n5494), .Z(n5577) );
  XNOR U5687 ( .A(n9984), .B(n5960), .Z(n5574) );
  NANDN U5688 ( .A(n5574), .B(n9865), .Z(n5498) );
  NANDN U5689 ( .A(n5496), .B(n9930), .Z(n5497) );
  AND U5690 ( .A(n5498), .B(n5497), .Z(n5578) );
  XNOR U5691 ( .A(n5577), .B(n5578), .Z(n5579) );
  XNOR U5692 ( .A(n5580), .B(n5579), .Z(n5616) );
  NANDN U5693 ( .A(n5500), .B(n5499), .Z(n5504) );
  NAND U5694 ( .A(n5502), .B(n5501), .Z(n5503) );
  NAND U5695 ( .A(n5504), .B(n5503), .Z(n5617) );
  XNOR U5696 ( .A(n5616), .B(n5617), .Z(n5618) );
  NANDN U5697 ( .A(n5506), .B(n5505), .Z(n5510) );
  NAND U5698 ( .A(n5508), .B(n5507), .Z(n5509) );
  AND U5699 ( .A(n5510), .B(n5509), .Z(n5619) );
  XNOR U5700 ( .A(n5618), .B(n5619), .Z(n5563) );
  NANDN U5701 ( .A(n5512), .B(n5511), .Z(n5516) );
  OR U5702 ( .A(n5514), .B(n5513), .Z(n5515) );
  NAND U5703 ( .A(n5516), .B(n5515), .Z(n5613) );
  XNOR U5704 ( .A(n10050), .B(n5675), .Z(n5598) );
  OR U5705 ( .A(n5598), .B(n10051), .Z(n5519) );
  NANDN U5706 ( .A(n5517), .B(n10070), .Z(n5518) );
  AND U5707 ( .A(n5519), .B(n5518), .Z(n5590) );
  NAND U5708 ( .A(b[0]), .B(a[78]), .Z(n5520) );
  XNOR U5709 ( .A(b[1]), .B(n5520), .Z(n5522) );
  NAND U5710 ( .A(a[77]), .B(n72), .Z(n5521) );
  AND U5711 ( .A(n5522), .B(n5521), .Z(n5589) );
  XOR U5712 ( .A(n5590), .B(n5589), .Z(n5592) );
  NAND U5713 ( .A(a[62]), .B(b[15]), .Z(n5591) );
  XOR U5714 ( .A(n5592), .B(n5591), .Z(n5610) );
  XNOR U5715 ( .A(n9622), .B(n6272), .Z(n5601) );
  OR U5716 ( .A(n5601), .B(n9623), .Z(n5525) );
  NANDN U5717 ( .A(n5523), .B(n9680), .Z(n5524) );
  NAND U5718 ( .A(n5525), .B(n5524), .Z(n5586) );
  XNOR U5719 ( .A(n9872), .B(n6143), .Z(n5604) );
  NANDN U5720 ( .A(n5604), .B(n9746), .Z(n5528) );
  NANDN U5721 ( .A(n5526), .B(n9747), .Z(n5527) );
  NAND U5722 ( .A(n5528), .B(n5527), .Z(n5583) );
  IV U5723 ( .A(a[76]), .Z(n6428) );
  XNOR U5724 ( .A(n74), .B(n6428), .Z(n5607) );
  NANDN U5725 ( .A(n5607), .B(n9485), .Z(n5531) );
  NANDN U5726 ( .A(n5529), .B(n9484), .Z(n5530) );
  AND U5727 ( .A(n5531), .B(n5530), .Z(n5584) );
  XNOR U5728 ( .A(n5583), .B(n5584), .Z(n5585) );
  XOR U5729 ( .A(n5586), .B(n5585), .Z(n5611) );
  XOR U5730 ( .A(n5610), .B(n5611), .Z(n5612) );
  XNOR U5731 ( .A(n5613), .B(n5612), .Z(n5561) );
  NAND U5732 ( .A(n5533), .B(n5532), .Z(n5537) );
  NAND U5733 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U5734 ( .A(n5537), .B(n5536), .Z(n5562) );
  XOR U5735 ( .A(n5561), .B(n5562), .Z(n5564) );
  XNOR U5736 ( .A(n5563), .B(n5564), .Z(n5622) );
  NANDN U5737 ( .A(n5539), .B(n5538), .Z(n5543) );
  NAND U5738 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U5739 ( .A(n5543), .B(n5542), .Z(n5623) );
  XNOR U5740 ( .A(n5622), .B(n5623), .Z(n5624) );
  XOR U5741 ( .A(n5625), .B(n5624), .Z(n5555) );
  NANDN U5742 ( .A(n5545), .B(n5544), .Z(n5549) );
  NANDN U5743 ( .A(n5547), .B(n5546), .Z(n5548) );
  NAND U5744 ( .A(n5549), .B(n5548), .Z(n5556) );
  XNOR U5745 ( .A(n5555), .B(n5556), .Z(n5557) );
  XNOR U5746 ( .A(n5558), .B(n5557), .Z(n5628) );
  XNOR U5747 ( .A(n5628), .B(sreg[190]), .Z(n5630) );
  NAND U5748 ( .A(n5550), .B(sreg[189]), .Z(n5554) );
  OR U5749 ( .A(n5552), .B(n5551), .Z(n5553) );
  AND U5750 ( .A(n5554), .B(n5553), .Z(n5629) );
  XOR U5751 ( .A(n5630), .B(n5629), .Z(c[190]) );
  NANDN U5752 ( .A(n5556), .B(n5555), .Z(n5560) );
  NAND U5753 ( .A(n5558), .B(n5557), .Z(n5559) );
  NAND U5754 ( .A(n5560), .B(n5559), .Z(n5636) );
  NANDN U5755 ( .A(n5562), .B(n5561), .Z(n5566) );
  OR U5756 ( .A(n5564), .B(n5563), .Z(n5565) );
  NAND U5757 ( .A(n5566), .B(n5565), .Z(n5703) );
  XNOR U5758 ( .A(n9967), .B(n5882), .Z(n5672) );
  OR U5759 ( .A(n5672), .B(n10020), .Z(n5569) );
  NANDN U5760 ( .A(n5567), .B(n9968), .Z(n5568) );
  NAND U5761 ( .A(n5569), .B(n5568), .Z(n5685) );
  XNOR U5762 ( .A(n75), .B(n5570), .Z(n5676) );
  OR U5763 ( .A(n5676), .B(n10106), .Z(n5573) );
  NANDN U5764 ( .A(n5571), .B(n10107), .Z(n5572) );
  NAND U5765 ( .A(n5573), .B(n5572), .Z(n5682) );
  XNOR U5766 ( .A(n9984), .B(n6038), .Z(n5679) );
  NANDN U5767 ( .A(n5679), .B(n9865), .Z(n5576) );
  NANDN U5768 ( .A(n5574), .B(n9930), .Z(n5575) );
  AND U5769 ( .A(n5576), .B(n5575), .Z(n5683) );
  XNOR U5770 ( .A(n5682), .B(n5683), .Z(n5684) );
  XNOR U5771 ( .A(n5685), .B(n5684), .Z(n5694) );
  NANDN U5772 ( .A(n5578), .B(n5577), .Z(n5582) );
  NAND U5773 ( .A(n5580), .B(n5579), .Z(n5581) );
  NAND U5774 ( .A(n5582), .B(n5581), .Z(n5695) );
  XNOR U5775 ( .A(n5694), .B(n5695), .Z(n5696) );
  NANDN U5776 ( .A(n5584), .B(n5583), .Z(n5588) );
  NAND U5777 ( .A(n5586), .B(n5585), .Z(n5587) );
  AND U5778 ( .A(n5588), .B(n5587), .Z(n5697) );
  XNOR U5779 ( .A(n5696), .B(n5697), .Z(n5641) );
  NANDN U5780 ( .A(n5590), .B(n5589), .Z(n5594) );
  OR U5781 ( .A(n5592), .B(n5591), .Z(n5593) );
  NAND U5782 ( .A(n5594), .B(n5593), .Z(n5669) );
  NAND U5783 ( .A(b[0]), .B(a[79]), .Z(n5595) );
  XNOR U5784 ( .A(b[1]), .B(n5595), .Z(n5597) );
  NAND U5785 ( .A(a[78]), .B(n72), .Z(n5596) );
  AND U5786 ( .A(n5597), .B(n5596), .Z(n5645) );
  XNOR U5787 ( .A(n10050), .B(n5726), .Z(n5654) );
  OR U5788 ( .A(n5654), .B(n10051), .Z(n5600) );
  NANDN U5789 ( .A(n5598), .B(n10070), .Z(n5599) );
  AND U5790 ( .A(n5600), .B(n5599), .Z(n5646) );
  XOR U5791 ( .A(n5645), .B(n5646), .Z(n5648) );
  NAND U5792 ( .A(a[63]), .B(b[15]), .Z(n5647) );
  XOR U5793 ( .A(n5648), .B(n5647), .Z(n5666) );
  XNOR U5794 ( .A(n9622), .B(n6377), .Z(n5657) );
  OR U5795 ( .A(n5657), .B(n9623), .Z(n5603) );
  NANDN U5796 ( .A(n5601), .B(n9680), .Z(n5602) );
  NAND U5797 ( .A(n5603), .B(n5602), .Z(n5691) );
  XNOR U5798 ( .A(n9872), .B(n6194), .Z(n5660) );
  NANDN U5799 ( .A(n5660), .B(n9746), .Z(n5606) );
  NANDN U5800 ( .A(n5604), .B(n9747), .Z(n5605) );
  NAND U5801 ( .A(n5606), .B(n5605), .Z(n5688) );
  IV U5802 ( .A(a[77]), .Z(n6533) );
  XNOR U5803 ( .A(n74), .B(n6533), .Z(n5663) );
  NANDN U5804 ( .A(n5663), .B(n9485), .Z(n5609) );
  NANDN U5805 ( .A(n5607), .B(n9484), .Z(n5608) );
  AND U5806 ( .A(n5609), .B(n5608), .Z(n5689) );
  XNOR U5807 ( .A(n5688), .B(n5689), .Z(n5690) );
  XOR U5808 ( .A(n5691), .B(n5690), .Z(n5667) );
  XOR U5809 ( .A(n5666), .B(n5667), .Z(n5668) );
  XNOR U5810 ( .A(n5669), .B(n5668), .Z(n5639) );
  NAND U5811 ( .A(n5611), .B(n5610), .Z(n5615) );
  NAND U5812 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U5813 ( .A(n5615), .B(n5614), .Z(n5640) );
  XOR U5814 ( .A(n5639), .B(n5640), .Z(n5642) );
  XNOR U5815 ( .A(n5641), .B(n5642), .Z(n5700) );
  NANDN U5816 ( .A(n5617), .B(n5616), .Z(n5621) );
  NAND U5817 ( .A(n5619), .B(n5618), .Z(n5620) );
  NAND U5818 ( .A(n5621), .B(n5620), .Z(n5701) );
  XNOR U5819 ( .A(n5700), .B(n5701), .Z(n5702) );
  XOR U5820 ( .A(n5703), .B(n5702), .Z(n5633) );
  NANDN U5821 ( .A(n5623), .B(n5622), .Z(n5627) );
  NANDN U5822 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U5823 ( .A(n5627), .B(n5626), .Z(n5634) );
  XNOR U5824 ( .A(n5633), .B(n5634), .Z(n5635) );
  XNOR U5825 ( .A(n5636), .B(n5635), .Z(n5706) );
  XNOR U5826 ( .A(n5706), .B(sreg[191]), .Z(n5708) );
  NAND U5827 ( .A(n5628), .B(sreg[190]), .Z(n5632) );
  OR U5828 ( .A(n5630), .B(n5629), .Z(n5631) );
  AND U5829 ( .A(n5632), .B(n5631), .Z(n5707) );
  XOR U5830 ( .A(n5708), .B(n5707), .Z(c[191]) );
  NANDN U5831 ( .A(n5634), .B(n5633), .Z(n5638) );
  NAND U5832 ( .A(n5636), .B(n5635), .Z(n5637) );
  NAND U5833 ( .A(n5638), .B(n5637), .Z(n5714) );
  NANDN U5834 ( .A(n5640), .B(n5639), .Z(n5644) );
  OR U5835 ( .A(n5642), .B(n5641), .Z(n5643) );
  NAND U5836 ( .A(n5644), .B(n5643), .Z(n5781) );
  NANDN U5837 ( .A(n5646), .B(n5645), .Z(n5650) );
  OR U5838 ( .A(n5648), .B(n5647), .Z(n5649) );
  NAND U5839 ( .A(n5650), .B(n5649), .Z(n5769) );
  NAND U5840 ( .A(b[0]), .B(a[80]), .Z(n5651) );
  XNOR U5841 ( .A(b[1]), .B(n5651), .Z(n5653) );
  NAND U5842 ( .A(a[79]), .B(n72), .Z(n5652) );
  AND U5843 ( .A(n5653), .B(n5652), .Z(n5745) );
  XNOR U5844 ( .A(n10050), .B(n5804), .Z(n5751) );
  OR U5845 ( .A(n5751), .B(n10051), .Z(n5656) );
  NANDN U5846 ( .A(n5654), .B(n10070), .Z(n5655) );
  AND U5847 ( .A(n5656), .B(n5655), .Z(n5746) );
  XOR U5848 ( .A(n5745), .B(n5746), .Z(n5748) );
  NAND U5849 ( .A(a[64]), .B(b[15]), .Z(n5747) );
  XOR U5850 ( .A(n5748), .B(n5747), .Z(n5766) );
  XNOR U5851 ( .A(n9622), .B(n6428), .Z(n5757) );
  OR U5852 ( .A(n5757), .B(n9623), .Z(n5659) );
  NANDN U5853 ( .A(n5657), .B(n9680), .Z(n5658) );
  NAND U5854 ( .A(n5659), .B(n5658), .Z(n5742) );
  XNOR U5855 ( .A(n9872), .B(n6272), .Z(n5760) );
  NANDN U5856 ( .A(n5760), .B(n9746), .Z(n5662) );
  NANDN U5857 ( .A(n5660), .B(n9747), .Z(n5661) );
  NAND U5858 ( .A(n5662), .B(n5661), .Z(n5739) );
  IV U5859 ( .A(a[78]), .Z(n6584) );
  XNOR U5860 ( .A(n74), .B(n6584), .Z(n5763) );
  NANDN U5861 ( .A(n5763), .B(n9485), .Z(n5665) );
  NANDN U5862 ( .A(n5663), .B(n9484), .Z(n5664) );
  AND U5863 ( .A(n5665), .B(n5664), .Z(n5740) );
  XNOR U5864 ( .A(n5739), .B(n5740), .Z(n5741) );
  XOR U5865 ( .A(n5742), .B(n5741), .Z(n5767) );
  XOR U5866 ( .A(n5766), .B(n5767), .Z(n5768) );
  XNOR U5867 ( .A(n5769), .B(n5768), .Z(n5717) );
  NAND U5868 ( .A(n5667), .B(n5666), .Z(n5671) );
  NAND U5869 ( .A(n5669), .B(n5668), .Z(n5670) );
  NAND U5870 ( .A(n5671), .B(n5670), .Z(n5718) );
  XOR U5871 ( .A(n5717), .B(n5718), .Z(n5720) );
  XNOR U5872 ( .A(n9967), .B(n5960), .Z(n5723) );
  OR U5873 ( .A(n5723), .B(n10020), .Z(n5674) );
  NANDN U5874 ( .A(n5672), .B(n9968), .Z(n5673) );
  NAND U5875 ( .A(n5674), .B(n5673), .Z(n5736) );
  XNOR U5876 ( .A(n75), .B(n5675), .Z(n5727) );
  OR U5877 ( .A(n5727), .B(n10106), .Z(n5678) );
  NANDN U5878 ( .A(n5676), .B(n10107), .Z(n5677) );
  NAND U5879 ( .A(n5678), .B(n5677), .Z(n5733) );
  XNOR U5880 ( .A(n9984), .B(n6143), .Z(n5730) );
  NANDN U5881 ( .A(n5730), .B(n9865), .Z(n5681) );
  NANDN U5882 ( .A(n5679), .B(n9930), .Z(n5680) );
  AND U5883 ( .A(n5681), .B(n5680), .Z(n5734) );
  XNOR U5884 ( .A(n5733), .B(n5734), .Z(n5735) );
  XNOR U5885 ( .A(n5736), .B(n5735), .Z(n5772) );
  NANDN U5886 ( .A(n5683), .B(n5682), .Z(n5687) );
  NAND U5887 ( .A(n5685), .B(n5684), .Z(n5686) );
  NAND U5888 ( .A(n5687), .B(n5686), .Z(n5773) );
  XNOR U5889 ( .A(n5772), .B(n5773), .Z(n5774) );
  NANDN U5890 ( .A(n5689), .B(n5688), .Z(n5693) );
  NAND U5891 ( .A(n5691), .B(n5690), .Z(n5692) );
  AND U5892 ( .A(n5693), .B(n5692), .Z(n5775) );
  XNOR U5893 ( .A(n5774), .B(n5775), .Z(n5719) );
  XNOR U5894 ( .A(n5720), .B(n5719), .Z(n5778) );
  NANDN U5895 ( .A(n5695), .B(n5694), .Z(n5699) );
  NAND U5896 ( .A(n5697), .B(n5696), .Z(n5698) );
  NAND U5897 ( .A(n5699), .B(n5698), .Z(n5779) );
  XNOR U5898 ( .A(n5778), .B(n5779), .Z(n5780) );
  XOR U5899 ( .A(n5781), .B(n5780), .Z(n5711) );
  NANDN U5900 ( .A(n5701), .B(n5700), .Z(n5705) );
  NANDN U5901 ( .A(n5703), .B(n5702), .Z(n5704) );
  NAND U5902 ( .A(n5705), .B(n5704), .Z(n5712) );
  XNOR U5903 ( .A(n5711), .B(n5712), .Z(n5713) );
  XNOR U5904 ( .A(n5714), .B(n5713), .Z(n5784) );
  XNOR U5905 ( .A(n5784), .B(sreg[192]), .Z(n5786) );
  NAND U5906 ( .A(n5706), .B(sreg[191]), .Z(n5710) );
  OR U5907 ( .A(n5708), .B(n5707), .Z(n5709) );
  AND U5908 ( .A(n5710), .B(n5709), .Z(n5785) );
  XOR U5909 ( .A(n5786), .B(n5785), .Z(c[192]) );
  NANDN U5910 ( .A(n5712), .B(n5711), .Z(n5716) );
  NAND U5911 ( .A(n5714), .B(n5713), .Z(n5715) );
  NAND U5912 ( .A(n5716), .B(n5715), .Z(n5792) );
  NANDN U5913 ( .A(n5718), .B(n5717), .Z(n5722) );
  OR U5914 ( .A(n5720), .B(n5719), .Z(n5721) );
  NAND U5915 ( .A(n5722), .B(n5721), .Z(n5859) );
  XNOR U5916 ( .A(n9967), .B(n6038), .Z(n5801) );
  OR U5917 ( .A(n5801), .B(n10020), .Z(n5725) );
  NANDN U5918 ( .A(n5723), .B(n9968), .Z(n5724) );
  NAND U5919 ( .A(n5725), .B(n5724), .Z(n5814) );
  XNOR U5920 ( .A(n75), .B(n5726), .Z(n5805) );
  OR U5921 ( .A(n5805), .B(n10106), .Z(n5729) );
  NANDN U5922 ( .A(n5727), .B(n10107), .Z(n5728) );
  NAND U5923 ( .A(n5729), .B(n5728), .Z(n5811) );
  XNOR U5924 ( .A(n9984), .B(n6194), .Z(n5808) );
  NANDN U5925 ( .A(n5808), .B(n9865), .Z(n5732) );
  NANDN U5926 ( .A(n5730), .B(n9930), .Z(n5731) );
  AND U5927 ( .A(n5732), .B(n5731), .Z(n5812) );
  XNOR U5928 ( .A(n5811), .B(n5812), .Z(n5813) );
  XNOR U5929 ( .A(n5814), .B(n5813), .Z(n5850) );
  NANDN U5930 ( .A(n5734), .B(n5733), .Z(n5738) );
  NAND U5931 ( .A(n5736), .B(n5735), .Z(n5737) );
  NAND U5932 ( .A(n5738), .B(n5737), .Z(n5851) );
  XNOR U5933 ( .A(n5850), .B(n5851), .Z(n5852) );
  NANDN U5934 ( .A(n5740), .B(n5739), .Z(n5744) );
  NAND U5935 ( .A(n5742), .B(n5741), .Z(n5743) );
  AND U5936 ( .A(n5744), .B(n5743), .Z(n5853) );
  XNOR U5937 ( .A(n5852), .B(n5853), .Z(n5797) );
  NANDN U5938 ( .A(n5746), .B(n5745), .Z(n5750) );
  OR U5939 ( .A(n5748), .B(n5747), .Z(n5749) );
  NAND U5940 ( .A(n5750), .B(n5749), .Z(n5847) );
  XNOR U5941 ( .A(n10050), .B(n5882), .Z(n5832) );
  OR U5942 ( .A(n5832), .B(n10051), .Z(n5753) );
  NANDN U5943 ( .A(n5751), .B(n10070), .Z(n5752) );
  AND U5944 ( .A(n5753), .B(n5752), .Z(n5824) );
  NAND U5945 ( .A(b[0]), .B(a[81]), .Z(n5754) );
  XNOR U5946 ( .A(b[1]), .B(n5754), .Z(n5756) );
  NAND U5947 ( .A(a[80]), .B(n72), .Z(n5755) );
  AND U5948 ( .A(n5756), .B(n5755), .Z(n5823) );
  XOR U5949 ( .A(n5824), .B(n5823), .Z(n5826) );
  NAND U5950 ( .A(a[65]), .B(b[15]), .Z(n5825) );
  XOR U5951 ( .A(n5826), .B(n5825), .Z(n5844) );
  XNOR U5952 ( .A(n9622), .B(n6533), .Z(n5835) );
  OR U5953 ( .A(n5835), .B(n9623), .Z(n5759) );
  NANDN U5954 ( .A(n5757), .B(n9680), .Z(n5758) );
  NAND U5955 ( .A(n5759), .B(n5758), .Z(n5820) );
  XNOR U5956 ( .A(n9872), .B(n6377), .Z(n5838) );
  NANDN U5957 ( .A(n5838), .B(n9746), .Z(n5762) );
  NANDN U5958 ( .A(n5760), .B(n9747), .Z(n5761) );
  NAND U5959 ( .A(n5762), .B(n5761), .Z(n5817) );
  IV U5960 ( .A(a[79]), .Z(n6662) );
  XNOR U5961 ( .A(n74), .B(n6662), .Z(n5841) );
  NANDN U5962 ( .A(n5841), .B(n9485), .Z(n5765) );
  NANDN U5963 ( .A(n5763), .B(n9484), .Z(n5764) );
  AND U5964 ( .A(n5765), .B(n5764), .Z(n5818) );
  XNOR U5965 ( .A(n5817), .B(n5818), .Z(n5819) );
  XOR U5966 ( .A(n5820), .B(n5819), .Z(n5845) );
  XOR U5967 ( .A(n5844), .B(n5845), .Z(n5846) );
  XNOR U5968 ( .A(n5847), .B(n5846), .Z(n5795) );
  NAND U5969 ( .A(n5767), .B(n5766), .Z(n5771) );
  NAND U5970 ( .A(n5769), .B(n5768), .Z(n5770) );
  NAND U5971 ( .A(n5771), .B(n5770), .Z(n5796) );
  XOR U5972 ( .A(n5795), .B(n5796), .Z(n5798) );
  XNOR U5973 ( .A(n5797), .B(n5798), .Z(n5856) );
  NANDN U5974 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U5975 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U5976 ( .A(n5777), .B(n5776), .Z(n5857) );
  XNOR U5977 ( .A(n5856), .B(n5857), .Z(n5858) );
  XOR U5978 ( .A(n5859), .B(n5858), .Z(n5789) );
  NANDN U5979 ( .A(n5779), .B(n5778), .Z(n5783) );
  NANDN U5980 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U5981 ( .A(n5783), .B(n5782), .Z(n5790) );
  XNOR U5982 ( .A(n5789), .B(n5790), .Z(n5791) );
  XNOR U5983 ( .A(n5792), .B(n5791), .Z(n5862) );
  XNOR U5984 ( .A(n5862), .B(sreg[193]), .Z(n5864) );
  NAND U5985 ( .A(n5784), .B(sreg[192]), .Z(n5788) );
  OR U5986 ( .A(n5786), .B(n5785), .Z(n5787) );
  AND U5987 ( .A(n5788), .B(n5787), .Z(n5863) );
  XOR U5988 ( .A(n5864), .B(n5863), .Z(c[193]) );
  NANDN U5989 ( .A(n5790), .B(n5789), .Z(n5794) );
  NAND U5990 ( .A(n5792), .B(n5791), .Z(n5793) );
  NAND U5991 ( .A(n5794), .B(n5793), .Z(n5870) );
  NANDN U5992 ( .A(n5796), .B(n5795), .Z(n5800) );
  OR U5993 ( .A(n5798), .B(n5797), .Z(n5799) );
  NAND U5994 ( .A(n5800), .B(n5799), .Z(n5937) );
  XNOR U5995 ( .A(n9967), .B(n6143), .Z(n5879) );
  OR U5996 ( .A(n5879), .B(n10020), .Z(n5803) );
  NANDN U5997 ( .A(n5801), .B(n9968), .Z(n5802) );
  NAND U5998 ( .A(n5803), .B(n5802), .Z(n5892) );
  XNOR U5999 ( .A(n75), .B(n5804), .Z(n5883) );
  OR U6000 ( .A(n5883), .B(n10106), .Z(n5807) );
  NANDN U6001 ( .A(n5805), .B(n10107), .Z(n5806) );
  NAND U6002 ( .A(n5807), .B(n5806), .Z(n5889) );
  XNOR U6003 ( .A(n9984), .B(n6272), .Z(n5886) );
  NANDN U6004 ( .A(n5886), .B(n9865), .Z(n5810) );
  NANDN U6005 ( .A(n5808), .B(n9930), .Z(n5809) );
  AND U6006 ( .A(n5810), .B(n5809), .Z(n5890) );
  XNOR U6007 ( .A(n5889), .B(n5890), .Z(n5891) );
  XNOR U6008 ( .A(n5892), .B(n5891), .Z(n5928) );
  NANDN U6009 ( .A(n5812), .B(n5811), .Z(n5816) );
  NAND U6010 ( .A(n5814), .B(n5813), .Z(n5815) );
  NAND U6011 ( .A(n5816), .B(n5815), .Z(n5929) );
  XNOR U6012 ( .A(n5928), .B(n5929), .Z(n5930) );
  NANDN U6013 ( .A(n5818), .B(n5817), .Z(n5822) );
  NAND U6014 ( .A(n5820), .B(n5819), .Z(n5821) );
  AND U6015 ( .A(n5822), .B(n5821), .Z(n5931) );
  XNOR U6016 ( .A(n5930), .B(n5931), .Z(n5875) );
  NANDN U6017 ( .A(n5824), .B(n5823), .Z(n5828) );
  OR U6018 ( .A(n5826), .B(n5825), .Z(n5827) );
  NAND U6019 ( .A(n5828), .B(n5827), .Z(n5925) );
  NAND U6020 ( .A(b[0]), .B(a[82]), .Z(n5829) );
  XNOR U6021 ( .A(b[1]), .B(n5829), .Z(n5831) );
  NAND U6022 ( .A(a[81]), .B(n72), .Z(n5830) );
  AND U6023 ( .A(n5831), .B(n5830), .Z(n5901) );
  XNOR U6024 ( .A(n10050), .B(n5960), .Z(n5907) );
  OR U6025 ( .A(n5907), .B(n10051), .Z(n5834) );
  NANDN U6026 ( .A(n5832), .B(n10070), .Z(n5833) );
  AND U6027 ( .A(n5834), .B(n5833), .Z(n5902) );
  XOR U6028 ( .A(n5901), .B(n5902), .Z(n5904) );
  NAND U6029 ( .A(a[66]), .B(b[15]), .Z(n5903) );
  XOR U6030 ( .A(n5904), .B(n5903), .Z(n5922) );
  XNOR U6031 ( .A(n9622), .B(n6584), .Z(n5913) );
  OR U6032 ( .A(n5913), .B(n9623), .Z(n5837) );
  NANDN U6033 ( .A(n5835), .B(n9680), .Z(n5836) );
  NAND U6034 ( .A(n5837), .B(n5836), .Z(n5898) );
  XNOR U6035 ( .A(n9872), .B(n6428), .Z(n5916) );
  NANDN U6036 ( .A(n5916), .B(n9746), .Z(n5840) );
  NANDN U6037 ( .A(n5838), .B(n9747), .Z(n5839) );
  NAND U6038 ( .A(n5840), .B(n5839), .Z(n5895) );
  IV U6039 ( .A(a[80]), .Z(n6740) );
  XNOR U6040 ( .A(n74), .B(n6740), .Z(n5919) );
  NANDN U6041 ( .A(n5919), .B(n9485), .Z(n5843) );
  NANDN U6042 ( .A(n5841), .B(n9484), .Z(n5842) );
  AND U6043 ( .A(n5843), .B(n5842), .Z(n5896) );
  XNOR U6044 ( .A(n5895), .B(n5896), .Z(n5897) );
  XOR U6045 ( .A(n5898), .B(n5897), .Z(n5923) );
  XOR U6046 ( .A(n5922), .B(n5923), .Z(n5924) );
  XNOR U6047 ( .A(n5925), .B(n5924), .Z(n5873) );
  NAND U6048 ( .A(n5845), .B(n5844), .Z(n5849) );
  NAND U6049 ( .A(n5847), .B(n5846), .Z(n5848) );
  NAND U6050 ( .A(n5849), .B(n5848), .Z(n5874) );
  XOR U6051 ( .A(n5873), .B(n5874), .Z(n5876) );
  XNOR U6052 ( .A(n5875), .B(n5876), .Z(n5934) );
  NANDN U6053 ( .A(n5851), .B(n5850), .Z(n5855) );
  NAND U6054 ( .A(n5853), .B(n5852), .Z(n5854) );
  NAND U6055 ( .A(n5855), .B(n5854), .Z(n5935) );
  XNOR U6056 ( .A(n5934), .B(n5935), .Z(n5936) );
  XOR U6057 ( .A(n5937), .B(n5936), .Z(n5867) );
  NANDN U6058 ( .A(n5857), .B(n5856), .Z(n5861) );
  NANDN U6059 ( .A(n5859), .B(n5858), .Z(n5860) );
  NAND U6060 ( .A(n5861), .B(n5860), .Z(n5868) );
  XNOR U6061 ( .A(n5867), .B(n5868), .Z(n5869) );
  XNOR U6062 ( .A(n5870), .B(n5869), .Z(n5940) );
  XNOR U6063 ( .A(n5940), .B(sreg[194]), .Z(n5942) );
  NAND U6064 ( .A(n5862), .B(sreg[193]), .Z(n5866) );
  OR U6065 ( .A(n5864), .B(n5863), .Z(n5865) );
  AND U6066 ( .A(n5866), .B(n5865), .Z(n5941) );
  XOR U6067 ( .A(n5942), .B(n5941), .Z(c[194]) );
  NANDN U6068 ( .A(n5868), .B(n5867), .Z(n5872) );
  NAND U6069 ( .A(n5870), .B(n5869), .Z(n5871) );
  NAND U6070 ( .A(n5872), .B(n5871), .Z(n5948) );
  NANDN U6071 ( .A(n5874), .B(n5873), .Z(n5878) );
  OR U6072 ( .A(n5876), .B(n5875), .Z(n5877) );
  NAND U6073 ( .A(n5878), .B(n5877), .Z(n6015) );
  XNOR U6074 ( .A(n9967), .B(n6194), .Z(n5957) );
  OR U6075 ( .A(n5957), .B(n10020), .Z(n5881) );
  NANDN U6076 ( .A(n5879), .B(n9968), .Z(n5880) );
  NAND U6077 ( .A(n5881), .B(n5880), .Z(n5970) );
  XNOR U6078 ( .A(n75), .B(n5882), .Z(n5961) );
  OR U6079 ( .A(n5961), .B(n10106), .Z(n5885) );
  NANDN U6080 ( .A(n5883), .B(n10107), .Z(n5884) );
  NAND U6081 ( .A(n5885), .B(n5884), .Z(n5967) );
  XNOR U6082 ( .A(n9984), .B(n6377), .Z(n5964) );
  NANDN U6083 ( .A(n5964), .B(n9865), .Z(n5888) );
  NANDN U6084 ( .A(n5886), .B(n9930), .Z(n5887) );
  AND U6085 ( .A(n5888), .B(n5887), .Z(n5968) );
  XNOR U6086 ( .A(n5967), .B(n5968), .Z(n5969) );
  XNOR U6087 ( .A(n5970), .B(n5969), .Z(n6006) );
  NANDN U6088 ( .A(n5890), .B(n5889), .Z(n5894) );
  NAND U6089 ( .A(n5892), .B(n5891), .Z(n5893) );
  NAND U6090 ( .A(n5894), .B(n5893), .Z(n6007) );
  XNOR U6091 ( .A(n6006), .B(n6007), .Z(n6008) );
  NANDN U6092 ( .A(n5896), .B(n5895), .Z(n5900) );
  NAND U6093 ( .A(n5898), .B(n5897), .Z(n5899) );
  AND U6094 ( .A(n5900), .B(n5899), .Z(n6009) );
  XNOR U6095 ( .A(n6008), .B(n6009), .Z(n5953) );
  NANDN U6096 ( .A(n5902), .B(n5901), .Z(n5906) );
  OR U6097 ( .A(n5904), .B(n5903), .Z(n5905) );
  NAND U6098 ( .A(n5906), .B(n5905), .Z(n6003) );
  XNOR U6099 ( .A(n10050), .B(n6038), .Z(n5988) );
  OR U6100 ( .A(n5988), .B(n10051), .Z(n5909) );
  NANDN U6101 ( .A(n5907), .B(n10070), .Z(n5908) );
  AND U6102 ( .A(n5909), .B(n5908), .Z(n5980) );
  NAND U6103 ( .A(b[0]), .B(a[83]), .Z(n5910) );
  XNOR U6104 ( .A(b[1]), .B(n5910), .Z(n5912) );
  NAND U6105 ( .A(a[82]), .B(n72), .Z(n5911) );
  AND U6106 ( .A(n5912), .B(n5911), .Z(n5979) );
  XOR U6107 ( .A(n5980), .B(n5979), .Z(n5982) );
  NAND U6108 ( .A(a[67]), .B(b[15]), .Z(n5981) );
  XOR U6109 ( .A(n5982), .B(n5981), .Z(n6000) );
  XNOR U6110 ( .A(n9622), .B(n6662), .Z(n5991) );
  OR U6111 ( .A(n5991), .B(n9623), .Z(n5915) );
  NANDN U6112 ( .A(n5913), .B(n9680), .Z(n5914) );
  NAND U6113 ( .A(n5915), .B(n5914), .Z(n5976) );
  XNOR U6114 ( .A(n9872), .B(n6533), .Z(n5994) );
  NANDN U6115 ( .A(n5994), .B(n9746), .Z(n5918) );
  NANDN U6116 ( .A(n5916), .B(n9747), .Z(n5917) );
  NAND U6117 ( .A(n5918), .B(n5917), .Z(n5973) );
  IV U6118 ( .A(a[81]), .Z(n6845) );
  XNOR U6119 ( .A(n74), .B(n6845), .Z(n5997) );
  NANDN U6120 ( .A(n5997), .B(n9485), .Z(n5921) );
  NANDN U6121 ( .A(n5919), .B(n9484), .Z(n5920) );
  AND U6122 ( .A(n5921), .B(n5920), .Z(n5974) );
  XNOR U6123 ( .A(n5973), .B(n5974), .Z(n5975) );
  XOR U6124 ( .A(n5976), .B(n5975), .Z(n6001) );
  XOR U6125 ( .A(n6000), .B(n6001), .Z(n6002) );
  XNOR U6126 ( .A(n6003), .B(n6002), .Z(n5951) );
  NAND U6127 ( .A(n5923), .B(n5922), .Z(n5927) );
  NAND U6128 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U6129 ( .A(n5927), .B(n5926), .Z(n5952) );
  XOR U6130 ( .A(n5951), .B(n5952), .Z(n5954) );
  XNOR U6131 ( .A(n5953), .B(n5954), .Z(n6012) );
  NANDN U6132 ( .A(n5929), .B(n5928), .Z(n5933) );
  NAND U6133 ( .A(n5931), .B(n5930), .Z(n5932) );
  NAND U6134 ( .A(n5933), .B(n5932), .Z(n6013) );
  XNOR U6135 ( .A(n6012), .B(n6013), .Z(n6014) );
  XOR U6136 ( .A(n6015), .B(n6014), .Z(n5945) );
  NANDN U6137 ( .A(n5935), .B(n5934), .Z(n5939) );
  NANDN U6138 ( .A(n5937), .B(n5936), .Z(n5938) );
  NAND U6139 ( .A(n5939), .B(n5938), .Z(n5946) );
  XNOR U6140 ( .A(n5945), .B(n5946), .Z(n5947) );
  XNOR U6141 ( .A(n5948), .B(n5947), .Z(n6018) );
  XNOR U6142 ( .A(n6018), .B(sreg[195]), .Z(n6020) );
  NAND U6143 ( .A(n5940), .B(sreg[194]), .Z(n5944) );
  OR U6144 ( .A(n5942), .B(n5941), .Z(n5943) );
  AND U6145 ( .A(n5944), .B(n5943), .Z(n6019) );
  XOR U6146 ( .A(n6020), .B(n6019), .Z(c[195]) );
  NANDN U6147 ( .A(n5946), .B(n5945), .Z(n5950) );
  NAND U6148 ( .A(n5948), .B(n5947), .Z(n5949) );
  NAND U6149 ( .A(n5950), .B(n5949), .Z(n6026) );
  NANDN U6150 ( .A(n5952), .B(n5951), .Z(n5956) );
  OR U6151 ( .A(n5954), .B(n5953), .Z(n5955) );
  NAND U6152 ( .A(n5956), .B(n5955), .Z(n6093) );
  XNOR U6153 ( .A(n9967), .B(n6272), .Z(n6035) );
  OR U6154 ( .A(n6035), .B(n10020), .Z(n5959) );
  NANDN U6155 ( .A(n5957), .B(n9968), .Z(n5958) );
  NAND U6156 ( .A(n5959), .B(n5958), .Z(n6048) );
  XNOR U6157 ( .A(n75), .B(n5960), .Z(n6039) );
  OR U6158 ( .A(n6039), .B(n10106), .Z(n5963) );
  NANDN U6159 ( .A(n5961), .B(n10107), .Z(n5962) );
  NAND U6160 ( .A(n5963), .B(n5962), .Z(n6045) );
  XNOR U6161 ( .A(n9984), .B(n6428), .Z(n6042) );
  NANDN U6162 ( .A(n6042), .B(n9865), .Z(n5966) );
  NANDN U6163 ( .A(n5964), .B(n9930), .Z(n5965) );
  AND U6164 ( .A(n5966), .B(n5965), .Z(n6046) );
  XNOR U6165 ( .A(n6045), .B(n6046), .Z(n6047) );
  XNOR U6166 ( .A(n6048), .B(n6047), .Z(n6084) );
  NANDN U6167 ( .A(n5968), .B(n5967), .Z(n5972) );
  NAND U6168 ( .A(n5970), .B(n5969), .Z(n5971) );
  NAND U6169 ( .A(n5972), .B(n5971), .Z(n6085) );
  XNOR U6170 ( .A(n6084), .B(n6085), .Z(n6086) );
  NANDN U6171 ( .A(n5974), .B(n5973), .Z(n5978) );
  NAND U6172 ( .A(n5976), .B(n5975), .Z(n5977) );
  AND U6173 ( .A(n5978), .B(n5977), .Z(n6087) );
  XNOR U6174 ( .A(n6086), .B(n6087), .Z(n6031) );
  NANDN U6175 ( .A(n5980), .B(n5979), .Z(n5984) );
  OR U6176 ( .A(n5982), .B(n5981), .Z(n5983) );
  NAND U6177 ( .A(n5984), .B(n5983), .Z(n6081) );
  NAND U6178 ( .A(b[0]), .B(a[84]), .Z(n5985) );
  XNOR U6179 ( .A(b[1]), .B(n5985), .Z(n5987) );
  NAND U6180 ( .A(a[83]), .B(n72), .Z(n5986) );
  AND U6181 ( .A(n5987), .B(n5986), .Z(n6057) );
  XNOR U6182 ( .A(n10050), .B(n6143), .Z(n6066) );
  OR U6183 ( .A(n6066), .B(n10051), .Z(n5990) );
  NANDN U6184 ( .A(n5988), .B(n10070), .Z(n5989) );
  AND U6185 ( .A(n5990), .B(n5989), .Z(n6058) );
  XOR U6186 ( .A(n6057), .B(n6058), .Z(n6060) );
  NAND U6187 ( .A(a[68]), .B(b[15]), .Z(n6059) );
  XOR U6188 ( .A(n6060), .B(n6059), .Z(n6078) );
  XNOR U6189 ( .A(n9622), .B(n6740), .Z(n6069) );
  OR U6190 ( .A(n6069), .B(n9623), .Z(n5993) );
  NANDN U6191 ( .A(n5991), .B(n9680), .Z(n5992) );
  NAND U6192 ( .A(n5993), .B(n5992), .Z(n6054) );
  XNOR U6193 ( .A(n9872), .B(n6584), .Z(n6072) );
  NANDN U6194 ( .A(n6072), .B(n9746), .Z(n5996) );
  NANDN U6195 ( .A(n5994), .B(n9747), .Z(n5995) );
  NAND U6196 ( .A(n5996), .B(n5995), .Z(n6051) );
  IV U6197 ( .A(a[82]), .Z(n6896) );
  XNOR U6198 ( .A(n74), .B(n6896), .Z(n6075) );
  NANDN U6199 ( .A(n6075), .B(n9485), .Z(n5999) );
  NANDN U6200 ( .A(n5997), .B(n9484), .Z(n5998) );
  AND U6201 ( .A(n5999), .B(n5998), .Z(n6052) );
  XNOR U6202 ( .A(n6051), .B(n6052), .Z(n6053) );
  XOR U6203 ( .A(n6054), .B(n6053), .Z(n6079) );
  XOR U6204 ( .A(n6078), .B(n6079), .Z(n6080) );
  XNOR U6205 ( .A(n6081), .B(n6080), .Z(n6029) );
  NAND U6206 ( .A(n6001), .B(n6000), .Z(n6005) );
  NAND U6207 ( .A(n6003), .B(n6002), .Z(n6004) );
  NAND U6208 ( .A(n6005), .B(n6004), .Z(n6030) );
  XOR U6209 ( .A(n6029), .B(n6030), .Z(n6032) );
  XNOR U6210 ( .A(n6031), .B(n6032), .Z(n6090) );
  NANDN U6211 ( .A(n6007), .B(n6006), .Z(n6011) );
  NAND U6212 ( .A(n6009), .B(n6008), .Z(n6010) );
  NAND U6213 ( .A(n6011), .B(n6010), .Z(n6091) );
  XNOR U6214 ( .A(n6090), .B(n6091), .Z(n6092) );
  XOR U6215 ( .A(n6093), .B(n6092), .Z(n6023) );
  NANDN U6216 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U6217 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U6218 ( .A(n6017), .B(n6016), .Z(n6024) );
  XNOR U6219 ( .A(n6023), .B(n6024), .Z(n6025) );
  XNOR U6220 ( .A(n6026), .B(n6025), .Z(n6096) );
  XNOR U6221 ( .A(n6096), .B(sreg[196]), .Z(n6098) );
  NAND U6222 ( .A(n6018), .B(sreg[195]), .Z(n6022) );
  OR U6223 ( .A(n6020), .B(n6019), .Z(n6021) );
  AND U6224 ( .A(n6022), .B(n6021), .Z(n6097) );
  XOR U6225 ( .A(n6098), .B(n6097), .Z(c[196]) );
  NANDN U6226 ( .A(n6024), .B(n6023), .Z(n6028) );
  NAND U6227 ( .A(n6026), .B(n6025), .Z(n6027) );
  NAND U6228 ( .A(n6028), .B(n6027), .Z(n6104) );
  NANDN U6229 ( .A(n6030), .B(n6029), .Z(n6034) );
  OR U6230 ( .A(n6032), .B(n6031), .Z(n6033) );
  NAND U6231 ( .A(n6034), .B(n6033), .Z(n6171) );
  XNOR U6232 ( .A(n9967), .B(n6377), .Z(n6140) );
  OR U6233 ( .A(n6140), .B(n10020), .Z(n6037) );
  NANDN U6234 ( .A(n6035), .B(n9968), .Z(n6036) );
  NAND U6235 ( .A(n6037), .B(n6036), .Z(n6153) );
  XNOR U6236 ( .A(n75), .B(n6038), .Z(n6144) );
  OR U6237 ( .A(n6144), .B(n10106), .Z(n6041) );
  NANDN U6238 ( .A(n6039), .B(n10107), .Z(n6040) );
  NAND U6239 ( .A(n6041), .B(n6040), .Z(n6150) );
  XNOR U6240 ( .A(n9984), .B(n6533), .Z(n6147) );
  NANDN U6241 ( .A(n6147), .B(n9865), .Z(n6044) );
  NANDN U6242 ( .A(n6042), .B(n9930), .Z(n6043) );
  AND U6243 ( .A(n6044), .B(n6043), .Z(n6151) );
  XNOR U6244 ( .A(n6150), .B(n6151), .Z(n6152) );
  XNOR U6245 ( .A(n6153), .B(n6152), .Z(n6162) );
  NANDN U6246 ( .A(n6046), .B(n6045), .Z(n6050) );
  NAND U6247 ( .A(n6048), .B(n6047), .Z(n6049) );
  NAND U6248 ( .A(n6050), .B(n6049), .Z(n6163) );
  XNOR U6249 ( .A(n6162), .B(n6163), .Z(n6164) );
  NANDN U6250 ( .A(n6052), .B(n6051), .Z(n6056) );
  NAND U6251 ( .A(n6054), .B(n6053), .Z(n6055) );
  AND U6252 ( .A(n6056), .B(n6055), .Z(n6165) );
  XNOR U6253 ( .A(n6164), .B(n6165), .Z(n6109) );
  NANDN U6254 ( .A(n6058), .B(n6057), .Z(n6062) );
  OR U6255 ( .A(n6060), .B(n6059), .Z(n6061) );
  NAND U6256 ( .A(n6062), .B(n6061), .Z(n6137) );
  NAND U6257 ( .A(b[0]), .B(a[85]), .Z(n6063) );
  XNOR U6258 ( .A(b[1]), .B(n6063), .Z(n6065) );
  NAND U6259 ( .A(a[84]), .B(n72), .Z(n6064) );
  AND U6260 ( .A(n6065), .B(n6064), .Z(n6113) );
  XNOR U6261 ( .A(n10050), .B(n6194), .Z(n6122) );
  OR U6262 ( .A(n6122), .B(n10051), .Z(n6068) );
  NANDN U6263 ( .A(n6066), .B(n10070), .Z(n6067) );
  AND U6264 ( .A(n6068), .B(n6067), .Z(n6114) );
  XOR U6265 ( .A(n6113), .B(n6114), .Z(n6116) );
  NAND U6266 ( .A(a[69]), .B(b[15]), .Z(n6115) );
  XOR U6267 ( .A(n6116), .B(n6115), .Z(n6134) );
  XNOR U6268 ( .A(n9622), .B(n6845), .Z(n6125) );
  OR U6269 ( .A(n6125), .B(n9623), .Z(n6071) );
  NANDN U6270 ( .A(n6069), .B(n9680), .Z(n6070) );
  NAND U6271 ( .A(n6071), .B(n6070), .Z(n6159) );
  XNOR U6272 ( .A(n9872), .B(n6662), .Z(n6128) );
  NANDN U6273 ( .A(n6128), .B(n9746), .Z(n6074) );
  NANDN U6274 ( .A(n6072), .B(n9747), .Z(n6073) );
  NAND U6275 ( .A(n6074), .B(n6073), .Z(n6156) );
  IV U6276 ( .A(a[83]), .Z(n7001) );
  XNOR U6277 ( .A(n74), .B(n7001), .Z(n6131) );
  NANDN U6278 ( .A(n6131), .B(n9485), .Z(n6077) );
  NANDN U6279 ( .A(n6075), .B(n9484), .Z(n6076) );
  AND U6280 ( .A(n6077), .B(n6076), .Z(n6157) );
  XNOR U6281 ( .A(n6156), .B(n6157), .Z(n6158) );
  XOR U6282 ( .A(n6159), .B(n6158), .Z(n6135) );
  XOR U6283 ( .A(n6134), .B(n6135), .Z(n6136) );
  XNOR U6284 ( .A(n6137), .B(n6136), .Z(n6107) );
  NAND U6285 ( .A(n6079), .B(n6078), .Z(n6083) );
  NAND U6286 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U6287 ( .A(n6083), .B(n6082), .Z(n6108) );
  XOR U6288 ( .A(n6107), .B(n6108), .Z(n6110) );
  XNOR U6289 ( .A(n6109), .B(n6110), .Z(n6168) );
  NANDN U6290 ( .A(n6085), .B(n6084), .Z(n6089) );
  NAND U6291 ( .A(n6087), .B(n6086), .Z(n6088) );
  NAND U6292 ( .A(n6089), .B(n6088), .Z(n6169) );
  XNOR U6293 ( .A(n6168), .B(n6169), .Z(n6170) );
  XOR U6294 ( .A(n6171), .B(n6170), .Z(n6101) );
  NANDN U6295 ( .A(n6091), .B(n6090), .Z(n6095) );
  NANDN U6296 ( .A(n6093), .B(n6092), .Z(n6094) );
  NAND U6297 ( .A(n6095), .B(n6094), .Z(n6102) );
  XNOR U6298 ( .A(n6101), .B(n6102), .Z(n6103) );
  XNOR U6299 ( .A(n6104), .B(n6103), .Z(n6174) );
  XNOR U6300 ( .A(n6174), .B(sreg[197]), .Z(n6176) );
  NAND U6301 ( .A(n6096), .B(sreg[196]), .Z(n6100) );
  OR U6302 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U6303 ( .A(n6100), .B(n6099), .Z(n6175) );
  XOR U6304 ( .A(n6176), .B(n6175), .Z(c[197]) );
  NANDN U6305 ( .A(n6102), .B(n6101), .Z(n6106) );
  NAND U6306 ( .A(n6104), .B(n6103), .Z(n6105) );
  NAND U6307 ( .A(n6106), .B(n6105), .Z(n6182) );
  NANDN U6308 ( .A(n6108), .B(n6107), .Z(n6112) );
  OR U6309 ( .A(n6110), .B(n6109), .Z(n6111) );
  NAND U6310 ( .A(n6112), .B(n6111), .Z(n6249) );
  NANDN U6311 ( .A(n6114), .B(n6113), .Z(n6118) );
  OR U6312 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6313 ( .A(n6118), .B(n6117), .Z(n6237) );
  NAND U6314 ( .A(b[0]), .B(a[86]), .Z(n6119) );
  XNOR U6315 ( .A(b[1]), .B(n6119), .Z(n6121) );
  NAND U6316 ( .A(a[85]), .B(n72), .Z(n6120) );
  AND U6317 ( .A(n6121), .B(n6120), .Z(n6213) );
  XNOR U6318 ( .A(n10050), .B(n6272), .Z(n6219) );
  OR U6319 ( .A(n6219), .B(n10051), .Z(n6124) );
  NANDN U6320 ( .A(n6122), .B(n10070), .Z(n6123) );
  AND U6321 ( .A(n6124), .B(n6123), .Z(n6214) );
  XOR U6322 ( .A(n6213), .B(n6214), .Z(n6216) );
  NAND U6323 ( .A(a[70]), .B(b[15]), .Z(n6215) );
  XOR U6324 ( .A(n6216), .B(n6215), .Z(n6234) );
  XNOR U6325 ( .A(n9622), .B(n6896), .Z(n6225) );
  OR U6326 ( .A(n6225), .B(n9623), .Z(n6127) );
  NANDN U6327 ( .A(n6125), .B(n9680), .Z(n6126) );
  NAND U6328 ( .A(n6127), .B(n6126), .Z(n6210) );
  XNOR U6329 ( .A(n9872), .B(n6740), .Z(n6228) );
  NANDN U6330 ( .A(n6228), .B(n9746), .Z(n6130) );
  NANDN U6331 ( .A(n6128), .B(n9747), .Z(n6129) );
  NAND U6332 ( .A(n6130), .B(n6129), .Z(n6207) );
  IV U6333 ( .A(a[84]), .Z(n7079) );
  XNOR U6334 ( .A(n74), .B(n7079), .Z(n6231) );
  NANDN U6335 ( .A(n6231), .B(n9485), .Z(n6133) );
  NANDN U6336 ( .A(n6131), .B(n9484), .Z(n6132) );
  AND U6337 ( .A(n6133), .B(n6132), .Z(n6208) );
  XNOR U6338 ( .A(n6207), .B(n6208), .Z(n6209) );
  XOR U6339 ( .A(n6210), .B(n6209), .Z(n6235) );
  XOR U6340 ( .A(n6234), .B(n6235), .Z(n6236) );
  XNOR U6341 ( .A(n6237), .B(n6236), .Z(n6185) );
  NAND U6342 ( .A(n6135), .B(n6134), .Z(n6139) );
  NAND U6343 ( .A(n6137), .B(n6136), .Z(n6138) );
  NAND U6344 ( .A(n6139), .B(n6138), .Z(n6186) );
  XOR U6345 ( .A(n6185), .B(n6186), .Z(n6188) );
  XNOR U6346 ( .A(n9967), .B(n6428), .Z(n6191) );
  OR U6347 ( .A(n6191), .B(n10020), .Z(n6142) );
  NANDN U6348 ( .A(n6140), .B(n9968), .Z(n6141) );
  NAND U6349 ( .A(n6142), .B(n6141), .Z(n6204) );
  XNOR U6350 ( .A(n75), .B(n6143), .Z(n6195) );
  OR U6351 ( .A(n6195), .B(n10106), .Z(n6146) );
  NANDN U6352 ( .A(n6144), .B(n10107), .Z(n6145) );
  NAND U6353 ( .A(n6146), .B(n6145), .Z(n6201) );
  XNOR U6354 ( .A(n9984), .B(n6584), .Z(n6198) );
  NANDN U6355 ( .A(n6198), .B(n9865), .Z(n6149) );
  NANDN U6356 ( .A(n6147), .B(n9930), .Z(n6148) );
  AND U6357 ( .A(n6149), .B(n6148), .Z(n6202) );
  XNOR U6358 ( .A(n6201), .B(n6202), .Z(n6203) );
  XNOR U6359 ( .A(n6204), .B(n6203), .Z(n6240) );
  NANDN U6360 ( .A(n6151), .B(n6150), .Z(n6155) );
  NAND U6361 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6362 ( .A(n6155), .B(n6154), .Z(n6241) );
  XNOR U6363 ( .A(n6240), .B(n6241), .Z(n6242) );
  NANDN U6364 ( .A(n6157), .B(n6156), .Z(n6161) );
  NAND U6365 ( .A(n6159), .B(n6158), .Z(n6160) );
  AND U6366 ( .A(n6161), .B(n6160), .Z(n6243) );
  XNOR U6367 ( .A(n6242), .B(n6243), .Z(n6187) );
  XNOR U6368 ( .A(n6188), .B(n6187), .Z(n6246) );
  NANDN U6369 ( .A(n6163), .B(n6162), .Z(n6167) );
  NAND U6370 ( .A(n6165), .B(n6164), .Z(n6166) );
  NAND U6371 ( .A(n6167), .B(n6166), .Z(n6247) );
  XNOR U6372 ( .A(n6246), .B(n6247), .Z(n6248) );
  XOR U6373 ( .A(n6249), .B(n6248), .Z(n6179) );
  NANDN U6374 ( .A(n6169), .B(n6168), .Z(n6173) );
  NANDN U6375 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U6376 ( .A(n6173), .B(n6172), .Z(n6180) );
  XNOR U6377 ( .A(n6179), .B(n6180), .Z(n6181) );
  XNOR U6378 ( .A(n6182), .B(n6181), .Z(n6252) );
  XNOR U6379 ( .A(n6252), .B(sreg[198]), .Z(n6254) );
  NAND U6380 ( .A(n6174), .B(sreg[197]), .Z(n6178) );
  OR U6381 ( .A(n6176), .B(n6175), .Z(n6177) );
  AND U6382 ( .A(n6178), .B(n6177), .Z(n6253) );
  XOR U6383 ( .A(n6254), .B(n6253), .Z(c[198]) );
  NANDN U6384 ( .A(n6180), .B(n6179), .Z(n6184) );
  NAND U6385 ( .A(n6182), .B(n6181), .Z(n6183) );
  NAND U6386 ( .A(n6184), .B(n6183), .Z(n6260) );
  NANDN U6387 ( .A(n6186), .B(n6185), .Z(n6190) );
  OR U6388 ( .A(n6188), .B(n6187), .Z(n6189) );
  NAND U6389 ( .A(n6190), .B(n6189), .Z(n6327) );
  XNOR U6390 ( .A(n9967), .B(n6533), .Z(n6269) );
  OR U6391 ( .A(n6269), .B(n10020), .Z(n6193) );
  NANDN U6392 ( .A(n6191), .B(n9968), .Z(n6192) );
  NAND U6393 ( .A(n6193), .B(n6192), .Z(n6282) );
  XNOR U6394 ( .A(n75), .B(n6194), .Z(n6273) );
  OR U6395 ( .A(n6273), .B(n10106), .Z(n6197) );
  NANDN U6396 ( .A(n6195), .B(n10107), .Z(n6196) );
  NAND U6397 ( .A(n6197), .B(n6196), .Z(n6279) );
  XNOR U6398 ( .A(n9984), .B(n6662), .Z(n6276) );
  NANDN U6399 ( .A(n6276), .B(n9865), .Z(n6200) );
  NANDN U6400 ( .A(n6198), .B(n9930), .Z(n6199) );
  AND U6401 ( .A(n6200), .B(n6199), .Z(n6280) );
  XNOR U6402 ( .A(n6279), .B(n6280), .Z(n6281) );
  XNOR U6403 ( .A(n6282), .B(n6281), .Z(n6318) );
  NANDN U6404 ( .A(n6202), .B(n6201), .Z(n6206) );
  NAND U6405 ( .A(n6204), .B(n6203), .Z(n6205) );
  NAND U6406 ( .A(n6206), .B(n6205), .Z(n6319) );
  XNOR U6407 ( .A(n6318), .B(n6319), .Z(n6320) );
  NANDN U6408 ( .A(n6208), .B(n6207), .Z(n6212) );
  NAND U6409 ( .A(n6210), .B(n6209), .Z(n6211) );
  AND U6410 ( .A(n6212), .B(n6211), .Z(n6321) );
  XNOR U6411 ( .A(n6320), .B(n6321), .Z(n6265) );
  NANDN U6412 ( .A(n6214), .B(n6213), .Z(n6218) );
  OR U6413 ( .A(n6216), .B(n6215), .Z(n6217) );
  NAND U6414 ( .A(n6218), .B(n6217), .Z(n6315) );
  XNOR U6415 ( .A(n10050), .B(n6377), .Z(n6300) );
  OR U6416 ( .A(n6300), .B(n10051), .Z(n6221) );
  NANDN U6417 ( .A(n6219), .B(n10070), .Z(n6220) );
  AND U6418 ( .A(n6221), .B(n6220), .Z(n6292) );
  NAND U6419 ( .A(b[0]), .B(a[87]), .Z(n6222) );
  XNOR U6420 ( .A(b[1]), .B(n6222), .Z(n6224) );
  NAND U6421 ( .A(a[86]), .B(n72), .Z(n6223) );
  AND U6422 ( .A(n6224), .B(n6223), .Z(n6291) );
  XOR U6423 ( .A(n6292), .B(n6291), .Z(n6294) );
  NAND U6424 ( .A(a[71]), .B(b[15]), .Z(n6293) );
  XOR U6425 ( .A(n6294), .B(n6293), .Z(n6312) );
  XNOR U6426 ( .A(n9622), .B(n7001), .Z(n6303) );
  OR U6427 ( .A(n6303), .B(n9623), .Z(n6227) );
  NANDN U6428 ( .A(n6225), .B(n9680), .Z(n6226) );
  NAND U6429 ( .A(n6227), .B(n6226), .Z(n6288) );
  XNOR U6430 ( .A(n9872), .B(n6845), .Z(n6306) );
  NANDN U6431 ( .A(n6306), .B(n9746), .Z(n6230) );
  NANDN U6432 ( .A(n6228), .B(n9747), .Z(n6229) );
  NAND U6433 ( .A(n6230), .B(n6229), .Z(n6285) );
  IV U6434 ( .A(a[85]), .Z(n7155) );
  XNOR U6435 ( .A(n74), .B(n7155), .Z(n6309) );
  NANDN U6436 ( .A(n6309), .B(n9485), .Z(n6233) );
  NANDN U6437 ( .A(n6231), .B(n9484), .Z(n6232) );
  AND U6438 ( .A(n6233), .B(n6232), .Z(n6286) );
  XNOR U6439 ( .A(n6285), .B(n6286), .Z(n6287) );
  XOR U6440 ( .A(n6288), .B(n6287), .Z(n6313) );
  XOR U6441 ( .A(n6312), .B(n6313), .Z(n6314) );
  XNOR U6442 ( .A(n6315), .B(n6314), .Z(n6263) );
  NAND U6443 ( .A(n6235), .B(n6234), .Z(n6239) );
  NAND U6444 ( .A(n6237), .B(n6236), .Z(n6238) );
  NAND U6445 ( .A(n6239), .B(n6238), .Z(n6264) );
  XOR U6446 ( .A(n6263), .B(n6264), .Z(n6266) );
  XNOR U6447 ( .A(n6265), .B(n6266), .Z(n6324) );
  NANDN U6448 ( .A(n6241), .B(n6240), .Z(n6245) );
  NAND U6449 ( .A(n6243), .B(n6242), .Z(n6244) );
  NAND U6450 ( .A(n6245), .B(n6244), .Z(n6325) );
  XNOR U6451 ( .A(n6324), .B(n6325), .Z(n6326) );
  XOR U6452 ( .A(n6327), .B(n6326), .Z(n6257) );
  NANDN U6453 ( .A(n6247), .B(n6246), .Z(n6251) );
  NANDN U6454 ( .A(n6249), .B(n6248), .Z(n6250) );
  NAND U6455 ( .A(n6251), .B(n6250), .Z(n6258) );
  XNOR U6456 ( .A(n6257), .B(n6258), .Z(n6259) );
  XNOR U6457 ( .A(n6260), .B(n6259), .Z(n6330) );
  XNOR U6458 ( .A(n6330), .B(sreg[199]), .Z(n6332) );
  NAND U6459 ( .A(n6252), .B(sreg[198]), .Z(n6256) );
  OR U6460 ( .A(n6254), .B(n6253), .Z(n6255) );
  AND U6461 ( .A(n6256), .B(n6255), .Z(n6331) );
  XOR U6462 ( .A(n6332), .B(n6331), .Z(c[199]) );
  NANDN U6463 ( .A(n6258), .B(n6257), .Z(n6262) );
  NAND U6464 ( .A(n6260), .B(n6259), .Z(n6261) );
  NAND U6465 ( .A(n6262), .B(n6261), .Z(n6338) );
  NANDN U6466 ( .A(n6264), .B(n6263), .Z(n6268) );
  OR U6467 ( .A(n6266), .B(n6265), .Z(n6267) );
  NAND U6468 ( .A(n6268), .B(n6267), .Z(n6405) );
  XNOR U6469 ( .A(n9967), .B(n6584), .Z(n6374) );
  OR U6470 ( .A(n6374), .B(n10020), .Z(n6271) );
  NANDN U6471 ( .A(n6269), .B(n9968), .Z(n6270) );
  NAND U6472 ( .A(n6271), .B(n6270), .Z(n6387) );
  XNOR U6473 ( .A(n75), .B(n6272), .Z(n6378) );
  OR U6474 ( .A(n6378), .B(n10106), .Z(n6275) );
  NANDN U6475 ( .A(n6273), .B(n10107), .Z(n6274) );
  NAND U6476 ( .A(n6275), .B(n6274), .Z(n6384) );
  XNOR U6477 ( .A(n9984), .B(n6740), .Z(n6381) );
  NANDN U6478 ( .A(n6381), .B(n9865), .Z(n6278) );
  NANDN U6479 ( .A(n6276), .B(n9930), .Z(n6277) );
  AND U6480 ( .A(n6278), .B(n6277), .Z(n6385) );
  XNOR U6481 ( .A(n6384), .B(n6385), .Z(n6386) );
  XNOR U6482 ( .A(n6387), .B(n6386), .Z(n6396) );
  NANDN U6483 ( .A(n6280), .B(n6279), .Z(n6284) );
  NAND U6484 ( .A(n6282), .B(n6281), .Z(n6283) );
  NAND U6485 ( .A(n6284), .B(n6283), .Z(n6397) );
  XNOR U6486 ( .A(n6396), .B(n6397), .Z(n6398) );
  NANDN U6487 ( .A(n6286), .B(n6285), .Z(n6290) );
  NAND U6488 ( .A(n6288), .B(n6287), .Z(n6289) );
  AND U6489 ( .A(n6290), .B(n6289), .Z(n6399) );
  XNOR U6490 ( .A(n6398), .B(n6399), .Z(n6343) );
  NANDN U6491 ( .A(n6292), .B(n6291), .Z(n6296) );
  OR U6492 ( .A(n6294), .B(n6293), .Z(n6295) );
  NAND U6493 ( .A(n6296), .B(n6295), .Z(n6371) );
  NAND U6494 ( .A(b[0]), .B(a[88]), .Z(n6297) );
  XNOR U6495 ( .A(b[1]), .B(n6297), .Z(n6299) );
  NAND U6496 ( .A(a[87]), .B(n72), .Z(n6298) );
  AND U6497 ( .A(n6299), .B(n6298), .Z(n6347) );
  XNOR U6498 ( .A(n10050), .B(n6428), .Z(n6356) );
  OR U6499 ( .A(n6356), .B(n10051), .Z(n6302) );
  NANDN U6500 ( .A(n6300), .B(n10070), .Z(n6301) );
  AND U6501 ( .A(n6302), .B(n6301), .Z(n6348) );
  XOR U6502 ( .A(n6347), .B(n6348), .Z(n6350) );
  NAND U6503 ( .A(a[72]), .B(b[15]), .Z(n6349) );
  XOR U6504 ( .A(n6350), .B(n6349), .Z(n6368) );
  XNOR U6505 ( .A(n9622), .B(n7079), .Z(n6359) );
  OR U6506 ( .A(n6359), .B(n9623), .Z(n6305) );
  NANDN U6507 ( .A(n6303), .B(n9680), .Z(n6304) );
  NAND U6508 ( .A(n6305), .B(n6304), .Z(n6393) );
  XNOR U6509 ( .A(n9872), .B(n6896), .Z(n6362) );
  NANDN U6510 ( .A(n6362), .B(n9746), .Z(n6308) );
  NANDN U6511 ( .A(n6306), .B(n9747), .Z(n6307) );
  NAND U6512 ( .A(n6308), .B(n6307), .Z(n6390) );
  IV U6513 ( .A(a[86]), .Z(n7233) );
  XNOR U6514 ( .A(n74), .B(n7233), .Z(n6365) );
  NANDN U6515 ( .A(n6365), .B(n9485), .Z(n6311) );
  NANDN U6516 ( .A(n6309), .B(n9484), .Z(n6310) );
  AND U6517 ( .A(n6311), .B(n6310), .Z(n6391) );
  XNOR U6518 ( .A(n6390), .B(n6391), .Z(n6392) );
  XOR U6519 ( .A(n6393), .B(n6392), .Z(n6369) );
  XOR U6520 ( .A(n6368), .B(n6369), .Z(n6370) );
  XNOR U6521 ( .A(n6371), .B(n6370), .Z(n6341) );
  NAND U6522 ( .A(n6313), .B(n6312), .Z(n6317) );
  NAND U6523 ( .A(n6315), .B(n6314), .Z(n6316) );
  NAND U6524 ( .A(n6317), .B(n6316), .Z(n6342) );
  XOR U6525 ( .A(n6341), .B(n6342), .Z(n6344) );
  XNOR U6526 ( .A(n6343), .B(n6344), .Z(n6402) );
  NANDN U6527 ( .A(n6319), .B(n6318), .Z(n6323) );
  NAND U6528 ( .A(n6321), .B(n6320), .Z(n6322) );
  NAND U6529 ( .A(n6323), .B(n6322), .Z(n6403) );
  XNOR U6530 ( .A(n6402), .B(n6403), .Z(n6404) );
  XOR U6531 ( .A(n6405), .B(n6404), .Z(n6335) );
  NANDN U6532 ( .A(n6325), .B(n6324), .Z(n6329) );
  NANDN U6533 ( .A(n6327), .B(n6326), .Z(n6328) );
  NAND U6534 ( .A(n6329), .B(n6328), .Z(n6336) );
  XNOR U6535 ( .A(n6335), .B(n6336), .Z(n6337) );
  XNOR U6536 ( .A(n6338), .B(n6337), .Z(n6408) );
  XNOR U6537 ( .A(n6408), .B(sreg[200]), .Z(n6410) );
  NAND U6538 ( .A(n6330), .B(sreg[199]), .Z(n6334) );
  OR U6539 ( .A(n6332), .B(n6331), .Z(n6333) );
  AND U6540 ( .A(n6334), .B(n6333), .Z(n6409) );
  XOR U6541 ( .A(n6410), .B(n6409), .Z(c[200]) );
  NANDN U6542 ( .A(n6336), .B(n6335), .Z(n6340) );
  NAND U6543 ( .A(n6338), .B(n6337), .Z(n6339) );
  NAND U6544 ( .A(n6340), .B(n6339), .Z(n6416) );
  NANDN U6545 ( .A(n6342), .B(n6341), .Z(n6346) );
  OR U6546 ( .A(n6344), .B(n6343), .Z(n6345) );
  NAND U6547 ( .A(n6346), .B(n6345), .Z(n6483) );
  NANDN U6548 ( .A(n6348), .B(n6347), .Z(n6352) );
  OR U6549 ( .A(n6350), .B(n6349), .Z(n6351) );
  NAND U6550 ( .A(n6352), .B(n6351), .Z(n6471) );
  NAND U6551 ( .A(b[0]), .B(a[89]), .Z(n6353) );
  XNOR U6552 ( .A(b[1]), .B(n6353), .Z(n6355) );
  NAND U6553 ( .A(a[88]), .B(n72), .Z(n6354) );
  AND U6554 ( .A(n6355), .B(n6354), .Z(n6447) );
  XNOR U6555 ( .A(n10050), .B(n6533), .Z(n6453) );
  OR U6556 ( .A(n6453), .B(n10051), .Z(n6358) );
  NANDN U6557 ( .A(n6356), .B(n10070), .Z(n6357) );
  AND U6558 ( .A(n6358), .B(n6357), .Z(n6448) );
  XOR U6559 ( .A(n6447), .B(n6448), .Z(n6450) );
  NAND U6560 ( .A(a[73]), .B(b[15]), .Z(n6449) );
  XOR U6561 ( .A(n6450), .B(n6449), .Z(n6468) );
  XNOR U6562 ( .A(n9622), .B(n7155), .Z(n6459) );
  OR U6563 ( .A(n6459), .B(n9623), .Z(n6361) );
  NANDN U6564 ( .A(n6359), .B(n9680), .Z(n6360) );
  NAND U6565 ( .A(n6361), .B(n6360), .Z(n6444) );
  XNOR U6566 ( .A(n9872), .B(n7001), .Z(n6462) );
  NANDN U6567 ( .A(n6462), .B(n9746), .Z(n6364) );
  NANDN U6568 ( .A(n6362), .B(n9747), .Z(n6363) );
  NAND U6569 ( .A(n6364), .B(n6363), .Z(n6441) );
  IV U6570 ( .A(a[87]), .Z(n7284) );
  XNOR U6571 ( .A(n74), .B(n7284), .Z(n6465) );
  NANDN U6572 ( .A(n6465), .B(n9485), .Z(n6367) );
  NANDN U6573 ( .A(n6365), .B(n9484), .Z(n6366) );
  AND U6574 ( .A(n6367), .B(n6366), .Z(n6442) );
  XNOR U6575 ( .A(n6441), .B(n6442), .Z(n6443) );
  XOR U6576 ( .A(n6444), .B(n6443), .Z(n6469) );
  XOR U6577 ( .A(n6468), .B(n6469), .Z(n6470) );
  XNOR U6578 ( .A(n6471), .B(n6470), .Z(n6419) );
  NAND U6579 ( .A(n6369), .B(n6368), .Z(n6373) );
  NAND U6580 ( .A(n6371), .B(n6370), .Z(n6372) );
  NAND U6581 ( .A(n6373), .B(n6372), .Z(n6420) );
  XOR U6582 ( .A(n6419), .B(n6420), .Z(n6422) );
  XNOR U6583 ( .A(n9967), .B(n6662), .Z(n6425) );
  OR U6584 ( .A(n6425), .B(n10020), .Z(n6376) );
  NANDN U6585 ( .A(n6374), .B(n9968), .Z(n6375) );
  NAND U6586 ( .A(n6376), .B(n6375), .Z(n6438) );
  XNOR U6587 ( .A(n75), .B(n6377), .Z(n6429) );
  OR U6588 ( .A(n6429), .B(n10106), .Z(n6380) );
  NANDN U6589 ( .A(n6378), .B(n10107), .Z(n6379) );
  NAND U6590 ( .A(n6380), .B(n6379), .Z(n6435) );
  XNOR U6591 ( .A(n9984), .B(n6845), .Z(n6432) );
  NANDN U6592 ( .A(n6432), .B(n9865), .Z(n6383) );
  NANDN U6593 ( .A(n6381), .B(n9930), .Z(n6382) );
  AND U6594 ( .A(n6383), .B(n6382), .Z(n6436) );
  XNOR U6595 ( .A(n6435), .B(n6436), .Z(n6437) );
  XNOR U6596 ( .A(n6438), .B(n6437), .Z(n6474) );
  NANDN U6597 ( .A(n6385), .B(n6384), .Z(n6389) );
  NAND U6598 ( .A(n6387), .B(n6386), .Z(n6388) );
  NAND U6599 ( .A(n6389), .B(n6388), .Z(n6475) );
  XNOR U6600 ( .A(n6474), .B(n6475), .Z(n6476) );
  NANDN U6601 ( .A(n6391), .B(n6390), .Z(n6395) );
  NAND U6602 ( .A(n6393), .B(n6392), .Z(n6394) );
  AND U6603 ( .A(n6395), .B(n6394), .Z(n6477) );
  XNOR U6604 ( .A(n6476), .B(n6477), .Z(n6421) );
  XNOR U6605 ( .A(n6422), .B(n6421), .Z(n6480) );
  NANDN U6606 ( .A(n6397), .B(n6396), .Z(n6401) );
  NAND U6607 ( .A(n6399), .B(n6398), .Z(n6400) );
  NAND U6608 ( .A(n6401), .B(n6400), .Z(n6481) );
  XNOR U6609 ( .A(n6480), .B(n6481), .Z(n6482) );
  XOR U6610 ( .A(n6483), .B(n6482), .Z(n6413) );
  NANDN U6611 ( .A(n6403), .B(n6402), .Z(n6407) );
  NANDN U6612 ( .A(n6405), .B(n6404), .Z(n6406) );
  NAND U6613 ( .A(n6407), .B(n6406), .Z(n6414) );
  XNOR U6614 ( .A(n6413), .B(n6414), .Z(n6415) );
  XNOR U6615 ( .A(n6416), .B(n6415), .Z(n6486) );
  XNOR U6616 ( .A(n6486), .B(sreg[201]), .Z(n6488) );
  NAND U6617 ( .A(n6408), .B(sreg[200]), .Z(n6412) );
  OR U6618 ( .A(n6410), .B(n6409), .Z(n6411) );
  AND U6619 ( .A(n6412), .B(n6411), .Z(n6487) );
  XOR U6620 ( .A(n6488), .B(n6487), .Z(c[201]) );
  NANDN U6621 ( .A(n6414), .B(n6413), .Z(n6418) );
  NAND U6622 ( .A(n6416), .B(n6415), .Z(n6417) );
  NAND U6623 ( .A(n6418), .B(n6417), .Z(n6494) );
  NANDN U6624 ( .A(n6420), .B(n6419), .Z(n6424) );
  OR U6625 ( .A(n6422), .B(n6421), .Z(n6423) );
  NAND U6626 ( .A(n6424), .B(n6423), .Z(n6561) );
  XNOR U6627 ( .A(n9967), .B(n6740), .Z(n6530) );
  OR U6628 ( .A(n6530), .B(n10020), .Z(n6427) );
  NANDN U6629 ( .A(n6425), .B(n9968), .Z(n6426) );
  NAND U6630 ( .A(n6427), .B(n6426), .Z(n6543) );
  XNOR U6631 ( .A(n75), .B(n6428), .Z(n6534) );
  OR U6632 ( .A(n6534), .B(n10106), .Z(n6431) );
  NANDN U6633 ( .A(n6429), .B(n10107), .Z(n6430) );
  NAND U6634 ( .A(n6431), .B(n6430), .Z(n6540) );
  XNOR U6635 ( .A(n9984), .B(n6896), .Z(n6537) );
  NANDN U6636 ( .A(n6537), .B(n9865), .Z(n6434) );
  NANDN U6637 ( .A(n6432), .B(n9930), .Z(n6433) );
  AND U6638 ( .A(n6434), .B(n6433), .Z(n6541) );
  XNOR U6639 ( .A(n6540), .B(n6541), .Z(n6542) );
  XNOR U6640 ( .A(n6543), .B(n6542), .Z(n6552) );
  NANDN U6641 ( .A(n6436), .B(n6435), .Z(n6440) );
  NAND U6642 ( .A(n6438), .B(n6437), .Z(n6439) );
  NAND U6643 ( .A(n6440), .B(n6439), .Z(n6553) );
  XNOR U6644 ( .A(n6552), .B(n6553), .Z(n6554) );
  NANDN U6645 ( .A(n6442), .B(n6441), .Z(n6446) );
  NAND U6646 ( .A(n6444), .B(n6443), .Z(n6445) );
  AND U6647 ( .A(n6446), .B(n6445), .Z(n6555) );
  XNOR U6648 ( .A(n6554), .B(n6555), .Z(n6499) );
  NANDN U6649 ( .A(n6448), .B(n6447), .Z(n6452) );
  OR U6650 ( .A(n6450), .B(n6449), .Z(n6451) );
  NAND U6651 ( .A(n6452), .B(n6451), .Z(n6527) );
  XNOR U6652 ( .A(n10050), .B(n6584), .Z(n6512) );
  OR U6653 ( .A(n6512), .B(n10051), .Z(n6455) );
  NANDN U6654 ( .A(n6453), .B(n10070), .Z(n6454) );
  AND U6655 ( .A(n6455), .B(n6454), .Z(n6504) );
  NAND U6656 ( .A(b[0]), .B(a[90]), .Z(n6456) );
  XNOR U6657 ( .A(b[1]), .B(n6456), .Z(n6458) );
  NAND U6658 ( .A(a[89]), .B(n72), .Z(n6457) );
  AND U6659 ( .A(n6458), .B(n6457), .Z(n6503) );
  XOR U6660 ( .A(n6504), .B(n6503), .Z(n6506) );
  NAND U6661 ( .A(a[74]), .B(b[15]), .Z(n6505) );
  XOR U6662 ( .A(n6506), .B(n6505), .Z(n6524) );
  XNOR U6663 ( .A(n9622), .B(n7233), .Z(n6515) );
  OR U6664 ( .A(n6515), .B(n9623), .Z(n6461) );
  NANDN U6665 ( .A(n6459), .B(n9680), .Z(n6460) );
  NAND U6666 ( .A(n6461), .B(n6460), .Z(n6549) );
  XNOR U6667 ( .A(n9872), .B(n7079), .Z(n6518) );
  NANDN U6668 ( .A(n6518), .B(n9746), .Z(n6464) );
  NANDN U6669 ( .A(n6462), .B(n9747), .Z(n6463) );
  NAND U6670 ( .A(n6464), .B(n6463), .Z(n6546) );
  IV U6671 ( .A(a[88]), .Z(n7389) );
  XNOR U6672 ( .A(n74), .B(n7389), .Z(n6521) );
  NANDN U6673 ( .A(n6521), .B(n9485), .Z(n6467) );
  NANDN U6674 ( .A(n6465), .B(n9484), .Z(n6466) );
  AND U6675 ( .A(n6467), .B(n6466), .Z(n6547) );
  XNOR U6676 ( .A(n6546), .B(n6547), .Z(n6548) );
  XOR U6677 ( .A(n6549), .B(n6548), .Z(n6525) );
  XOR U6678 ( .A(n6524), .B(n6525), .Z(n6526) );
  XNOR U6679 ( .A(n6527), .B(n6526), .Z(n6497) );
  NAND U6680 ( .A(n6469), .B(n6468), .Z(n6473) );
  NAND U6681 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U6682 ( .A(n6473), .B(n6472), .Z(n6498) );
  XOR U6683 ( .A(n6497), .B(n6498), .Z(n6500) );
  XNOR U6684 ( .A(n6499), .B(n6500), .Z(n6558) );
  NANDN U6685 ( .A(n6475), .B(n6474), .Z(n6479) );
  NAND U6686 ( .A(n6477), .B(n6476), .Z(n6478) );
  NAND U6687 ( .A(n6479), .B(n6478), .Z(n6559) );
  XNOR U6688 ( .A(n6558), .B(n6559), .Z(n6560) );
  XOR U6689 ( .A(n6561), .B(n6560), .Z(n6491) );
  NANDN U6690 ( .A(n6481), .B(n6480), .Z(n6485) );
  NANDN U6691 ( .A(n6483), .B(n6482), .Z(n6484) );
  NAND U6692 ( .A(n6485), .B(n6484), .Z(n6492) );
  XNOR U6693 ( .A(n6491), .B(n6492), .Z(n6493) );
  XNOR U6694 ( .A(n6494), .B(n6493), .Z(n6564) );
  XNOR U6695 ( .A(n6564), .B(sreg[202]), .Z(n6566) );
  NAND U6696 ( .A(n6486), .B(sreg[201]), .Z(n6490) );
  OR U6697 ( .A(n6488), .B(n6487), .Z(n6489) );
  AND U6698 ( .A(n6490), .B(n6489), .Z(n6565) );
  XOR U6699 ( .A(n6566), .B(n6565), .Z(c[202]) );
  NANDN U6700 ( .A(n6492), .B(n6491), .Z(n6496) );
  NAND U6701 ( .A(n6494), .B(n6493), .Z(n6495) );
  NAND U6702 ( .A(n6496), .B(n6495), .Z(n6572) );
  NANDN U6703 ( .A(n6498), .B(n6497), .Z(n6502) );
  OR U6704 ( .A(n6500), .B(n6499), .Z(n6501) );
  NAND U6705 ( .A(n6502), .B(n6501), .Z(n6639) );
  NANDN U6706 ( .A(n6504), .B(n6503), .Z(n6508) );
  OR U6707 ( .A(n6506), .B(n6505), .Z(n6507) );
  NAND U6708 ( .A(n6508), .B(n6507), .Z(n6627) );
  NAND U6709 ( .A(b[0]), .B(a[91]), .Z(n6509) );
  XNOR U6710 ( .A(b[1]), .B(n6509), .Z(n6511) );
  NAND U6711 ( .A(a[90]), .B(n72), .Z(n6510) );
  AND U6712 ( .A(n6511), .B(n6510), .Z(n6603) );
  XNOR U6713 ( .A(n10050), .B(n6662), .Z(n6612) );
  OR U6714 ( .A(n6612), .B(n10051), .Z(n6514) );
  NANDN U6715 ( .A(n6512), .B(n10070), .Z(n6513) );
  AND U6716 ( .A(n6514), .B(n6513), .Z(n6604) );
  XOR U6717 ( .A(n6603), .B(n6604), .Z(n6606) );
  NAND U6718 ( .A(a[75]), .B(b[15]), .Z(n6605) );
  XOR U6719 ( .A(n6606), .B(n6605), .Z(n6624) );
  XNOR U6720 ( .A(n9622), .B(n7284), .Z(n6615) );
  OR U6721 ( .A(n6615), .B(n9623), .Z(n6517) );
  NANDN U6722 ( .A(n6515), .B(n9680), .Z(n6516) );
  NAND U6723 ( .A(n6517), .B(n6516), .Z(n6600) );
  XNOR U6724 ( .A(n9872), .B(n7155), .Z(n6618) );
  NANDN U6725 ( .A(n6618), .B(n9746), .Z(n6520) );
  NANDN U6726 ( .A(n6518), .B(n9747), .Z(n6519) );
  NAND U6727 ( .A(n6520), .B(n6519), .Z(n6597) );
  IV U6728 ( .A(a[89]), .Z(n7467) );
  XNOR U6729 ( .A(n74), .B(n7467), .Z(n6621) );
  NANDN U6730 ( .A(n6621), .B(n9485), .Z(n6523) );
  NANDN U6731 ( .A(n6521), .B(n9484), .Z(n6522) );
  AND U6732 ( .A(n6523), .B(n6522), .Z(n6598) );
  XNOR U6733 ( .A(n6597), .B(n6598), .Z(n6599) );
  XOR U6734 ( .A(n6600), .B(n6599), .Z(n6625) );
  XOR U6735 ( .A(n6624), .B(n6625), .Z(n6626) );
  XNOR U6736 ( .A(n6627), .B(n6626), .Z(n6575) );
  NAND U6737 ( .A(n6525), .B(n6524), .Z(n6529) );
  NAND U6738 ( .A(n6527), .B(n6526), .Z(n6528) );
  NAND U6739 ( .A(n6529), .B(n6528), .Z(n6576) );
  XOR U6740 ( .A(n6575), .B(n6576), .Z(n6578) );
  XNOR U6741 ( .A(n9967), .B(n6845), .Z(n6581) );
  OR U6742 ( .A(n6581), .B(n10020), .Z(n6532) );
  NANDN U6743 ( .A(n6530), .B(n9968), .Z(n6531) );
  NAND U6744 ( .A(n6532), .B(n6531), .Z(n6594) );
  XNOR U6745 ( .A(n75), .B(n6533), .Z(n6585) );
  OR U6746 ( .A(n6585), .B(n10106), .Z(n6536) );
  NANDN U6747 ( .A(n6534), .B(n10107), .Z(n6535) );
  NAND U6748 ( .A(n6536), .B(n6535), .Z(n6591) );
  XNOR U6749 ( .A(n9984), .B(n7001), .Z(n6588) );
  NANDN U6750 ( .A(n6588), .B(n9865), .Z(n6539) );
  NANDN U6751 ( .A(n6537), .B(n9930), .Z(n6538) );
  AND U6752 ( .A(n6539), .B(n6538), .Z(n6592) );
  XNOR U6753 ( .A(n6591), .B(n6592), .Z(n6593) );
  XNOR U6754 ( .A(n6594), .B(n6593), .Z(n6630) );
  NANDN U6755 ( .A(n6541), .B(n6540), .Z(n6545) );
  NAND U6756 ( .A(n6543), .B(n6542), .Z(n6544) );
  NAND U6757 ( .A(n6545), .B(n6544), .Z(n6631) );
  XNOR U6758 ( .A(n6630), .B(n6631), .Z(n6632) );
  NANDN U6759 ( .A(n6547), .B(n6546), .Z(n6551) );
  NAND U6760 ( .A(n6549), .B(n6548), .Z(n6550) );
  AND U6761 ( .A(n6551), .B(n6550), .Z(n6633) );
  XNOR U6762 ( .A(n6632), .B(n6633), .Z(n6577) );
  XNOR U6763 ( .A(n6578), .B(n6577), .Z(n6636) );
  NANDN U6764 ( .A(n6553), .B(n6552), .Z(n6557) );
  NAND U6765 ( .A(n6555), .B(n6554), .Z(n6556) );
  NAND U6766 ( .A(n6557), .B(n6556), .Z(n6637) );
  XNOR U6767 ( .A(n6636), .B(n6637), .Z(n6638) );
  XOR U6768 ( .A(n6639), .B(n6638), .Z(n6569) );
  NANDN U6769 ( .A(n6559), .B(n6558), .Z(n6563) );
  NANDN U6770 ( .A(n6561), .B(n6560), .Z(n6562) );
  NAND U6771 ( .A(n6563), .B(n6562), .Z(n6570) );
  XNOR U6772 ( .A(n6569), .B(n6570), .Z(n6571) );
  XNOR U6773 ( .A(n6572), .B(n6571), .Z(n6642) );
  XNOR U6774 ( .A(n6642), .B(sreg[203]), .Z(n6644) );
  NAND U6775 ( .A(n6564), .B(sreg[202]), .Z(n6568) );
  OR U6776 ( .A(n6566), .B(n6565), .Z(n6567) );
  AND U6777 ( .A(n6568), .B(n6567), .Z(n6643) );
  XOR U6778 ( .A(n6644), .B(n6643), .Z(c[203]) );
  NANDN U6779 ( .A(n6570), .B(n6569), .Z(n6574) );
  NAND U6780 ( .A(n6572), .B(n6571), .Z(n6573) );
  NAND U6781 ( .A(n6574), .B(n6573), .Z(n6650) );
  NANDN U6782 ( .A(n6576), .B(n6575), .Z(n6580) );
  OR U6783 ( .A(n6578), .B(n6577), .Z(n6579) );
  NAND U6784 ( .A(n6580), .B(n6579), .Z(n6717) );
  XNOR U6785 ( .A(n9967), .B(n6896), .Z(n6659) );
  OR U6786 ( .A(n6659), .B(n10020), .Z(n6583) );
  NANDN U6787 ( .A(n6581), .B(n9968), .Z(n6582) );
  NAND U6788 ( .A(n6583), .B(n6582), .Z(n6672) );
  XNOR U6789 ( .A(n75), .B(n6584), .Z(n6663) );
  OR U6790 ( .A(n6663), .B(n10106), .Z(n6587) );
  NANDN U6791 ( .A(n6585), .B(n10107), .Z(n6586) );
  NAND U6792 ( .A(n6587), .B(n6586), .Z(n6669) );
  XNOR U6793 ( .A(n9984), .B(n7079), .Z(n6666) );
  NANDN U6794 ( .A(n6666), .B(n9865), .Z(n6590) );
  NANDN U6795 ( .A(n6588), .B(n9930), .Z(n6589) );
  AND U6796 ( .A(n6590), .B(n6589), .Z(n6670) );
  XNOR U6797 ( .A(n6669), .B(n6670), .Z(n6671) );
  XNOR U6798 ( .A(n6672), .B(n6671), .Z(n6708) );
  NANDN U6799 ( .A(n6592), .B(n6591), .Z(n6596) );
  NAND U6800 ( .A(n6594), .B(n6593), .Z(n6595) );
  NAND U6801 ( .A(n6596), .B(n6595), .Z(n6709) );
  XNOR U6802 ( .A(n6708), .B(n6709), .Z(n6710) );
  NANDN U6803 ( .A(n6598), .B(n6597), .Z(n6602) );
  NAND U6804 ( .A(n6600), .B(n6599), .Z(n6601) );
  AND U6805 ( .A(n6602), .B(n6601), .Z(n6711) );
  XNOR U6806 ( .A(n6710), .B(n6711), .Z(n6655) );
  NANDN U6807 ( .A(n6604), .B(n6603), .Z(n6608) );
  OR U6808 ( .A(n6606), .B(n6605), .Z(n6607) );
  NAND U6809 ( .A(n6608), .B(n6607), .Z(n6705) );
  NAND U6810 ( .A(b[0]), .B(a[92]), .Z(n6609) );
  XNOR U6811 ( .A(b[1]), .B(n6609), .Z(n6611) );
  NAND U6812 ( .A(a[91]), .B(n72), .Z(n6610) );
  AND U6813 ( .A(n6611), .B(n6610), .Z(n6681) );
  XNOR U6814 ( .A(n10050), .B(n6740), .Z(n6690) );
  OR U6815 ( .A(n6690), .B(n10051), .Z(n6614) );
  NANDN U6816 ( .A(n6612), .B(n10070), .Z(n6613) );
  AND U6817 ( .A(n6614), .B(n6613), .Z(n6682) );
  XOR U6818 ( .A(n6681), .B(n6682), .Z(n6684) );
  NAND U6819 ( .A(a[76]), .B(b[15]), .Z(n6683) );
  XOR U6820 ( .A(n6684), .B(n6683), .Z(n6702) );
  XNOR U6821 ( .A(n9622), .B(n7389), .Z(n6693) );
  OR U6822 ( .A(n6693), .B(n9623), .Z(n6617) );
  NANDN U6823 ( .A(n6615), .B(n9680), .Z(n6616) );
  NAND U6824 ( .A(n6617), .B(n6616), .Z(n6678) );
  XNOR U6825 ( .A(n9872), .B(n7233), .Z(n6696) );
  NANDN U6826 ( .A(n6696), .B(n9746), .Z(n6620) );
  NANDN U6827 ( .A(n6618), .B(n9747), .Z(n6619) );
  NAND U6828 ( .A(n6620), .B(n6619), .Z(n6675) );
  IV U6829 ( .A(a[90]), .Z(n7545) );
  XNOR U6830 ( .A(n74), .B(n7545), .Z(n6699) );
  NANDN U6831 ( .A(n6699), .B(n9485), .Z(n6623) );
  NANDN U6832 ( .A(n6621), .B(n9484), .Z(n6622) );
  AND U6833 ( .A(n6623), .B(n6622), .Z(n6676) );
  XNOR U6834 ( .A(n6675), .B(n6676), .Z(n6677) );
  XOR U6835 ( .A(n6678), .B(n6677), .Z(n6703) );
  XOR U6836 ( .A(n6702), .B(n6703), .Z(n6704) );
  XNOR U6837 ( .A(n6705), .B(n6704), .Z(n6653) );
  NAND U6838 ( .A(n6625), .B(n6624), .Z(n6629) );
  NAND U6839 ( .A(n6627), .B(n6626), .Z(n6628) );
  NAND U6840 ( .A(n6629), .B(n6628), .Z(n6654) );
  XOR U6841 ( .A(n6653), .B(n6654), .Z(n6656) );
  XNOR U6842 ( .A(n6655), .B(n6656), .Z(n6714) );
  NANDN U6843 ( .A(n6631), .B(n6630), .Z(n6635) );
  NAND U6844 ( .A(n6633), .B(n6632), .Z(n6634) );
  NAND U6845 ( .A(n6635), .B(n6634), .Z(n6715) );
  XNOR U6846 ( .A(n6714), .B(n6715), .Z(n6716) );
  XOR U6847 ( .A(n6717), .B(n6716), .Z(n6647) );
  NANDN U6848 ( .A(n6637), .B(n6636), .Z(n6641) );
  NANDN U6849 ( .A(n6639), .B(n6638), .Z(n6640) );
  NAND U6850 ( .A(n6641), .B(n6640), .Z(n6648) );
  XNOR U6851 ( .A(n6647), .B(n6648), .Z(n6649) );
  XNOR U6852 ( .A(n6650), .B(n6649), .Z(n6720) );
  XNOR U6853 ( .A(n6720), .B(sreg[204]), .Z(n6722) );
  NAND U6854 ( .A(n6642), .B(sreg[203]), .Z(n6646) );
  OR U6855 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U6856 ( .A(n6646), .B(n6645), .Z(n6721) );
  XOR U6857 ( .A(n6722), .B(n6721), .Z(c[204]) );
  NANDN U6858 ( .A(n6648), .B(n6647), .Z(n6652) );
  NAND U6859 ( .A(n6650), .B(n6649), .Z(n6651) );
  NAND U6860 ( .A(n6652), .B(n6651), .Z(n6728) );
  NANDN U6861 ( .A(n6654), .B(n6653), .Z(n6658) );
  OR U6862 ( .A(n6656), .B(n6655), .Z(n6657) );
  NAND U6863 ( .A(n6658), .B(n6657), .Z(n6795) );
  XNOR U6864 ( .A(n9967), .B(n7001), .Z(n6737) );
  OR U6865 ( .A(n6737), .B(n10020), .Z(n6661) );
  NANDN U6866 ( .A(n6659), .B(n9968), .Z(n6660) );
  NAND U6867 ( .A(n6661), .B(n6660), .Z(n6750) );
  XNOR U6868 ( .A(n75), .B(n6662), .Z(n6741) );
  OR U6869 ( .A(n6741), .B(n10106), .Z(n6665) );
  NANDN U6870 ( .A(n6663), .B(n10107), .Z(n6664) );
  NAND U6871 ( .A(n6665), .B(n6664), .Z(n6747) );
  XNOR U6872 ( .A(n9984), .B(n7155), .Z(n6744) );
  NANDN U6873 ( .A(n6744), .B(n9865), .Z(n6668) );
  NANDN U6874 ( .A(n6666), .B(n9930), .Z(n6667) );
  AND U6875 ( .A(n6668), .B(n6667), .Z(n6748) );
  XNOR U6876 ( .A(n6747), .B(n6748), .Z(n6749) );
  XNOR U6877 ( .A(n6750), .B(n6749), .Z(n6786) );
  NANDN U6878 ( .A(n6670), .B(n6669), .Z(n6674) );
  NAND U6879 ( .A(n6672), .B(n6671), .Z(n6673) );
  NAND U6880 ( .A(n6674), .B(n6673), .Z(n6787) );
  XNOR U6881 ( .A(n6786), .B(n6787), .Z(n6788) );
  NANDN U6882 ( .A(n6676), .B(n6675), .Z(n6680) );
  NAND U6883 ( .A(n6678), .B(n6677), .Z(n6679) );
  AND U6884 ( .A(n6680), .B(n6679), .Z(n6789) );
  XNOR U6885 ( .A(n6788), .B(n6789), .Z(n6733) );
  NANDN U6886 ( .A(n6682), .B(n6681), .Z(n6686) );
  OR U6887 ( .A(n6684), .B(n6683), .Z(n6685) );
  NAND U6888 ( .A(n6686), .B(n6685), .Z(n6783) );
  NAND U6889 ( .A(b[0]), .B(a[93]), .Z(n6687) );
  XNOR U6890 ( .A(b[1]), .B(n6687), .Z(n6689) );
  NAND U6891 ( .A(a[92]), .B(n72), .Z(n6688) );
  AND U6892 ( .A(n6689), .B(n6688), .Z(n6759) );
  XNOR U6893 ( .A(n10050), .B(n6845), .Z(n6768) );
  OR U6894 ( .A(n6768), .B(n10051), .Z(n6692) );
  NANDN U6895 ( .A(n6690), .B(n10070), .Z(n6691) );
  AND U6896 ( .A(n6692), .B(n6691), .Z(n6760) );
  XOR U6897 ( .A(n6759), .B(n6760), .Z(n6762) );
  NAND U6898 ( .A(a[77]), .B(b[15]), .Z(n6761) );
  XOR U6899 ( .A(n6762), .B(n6761), .Z(n6780) );
  XNOR U6900 ( .A(n9622), .B(n7467), .Z(n6771) );
  OR U6901 ( .A(n6771), .B(n9623), .Z(n6695) );
  NANDN U6902 ( .A(n6693), .B(n9680), .Z(n6694) );
  NAND U6903 ( .A(n6695), .B(n6694), .Z(n6756) );
  XNOR U6904 ( .A(n9872), .B(n7284), .Z(n6774) );
  NANDN U6905 ( .A(n6774), .B(n9746), .Z(n6698) );
  NANDN U6906 ( .A(n6696), .B(n9747), .Z(n6697) );
  NAND U6907 ( .A(n6698), .B(n6697), .Z(n6753) );
  IV U6908 ( .A(a[91]), .Z(n7623) );
  XNOR U6909 ( .A(n74), .B(n7623), .Z(n6777) );
  NANDN U6910 ( .A(n6777), .B(n9485), .Z(n6701) );
  NANDN U6911 ( .A(n6699), .B(n9484), .Z(n6700) );
  AND U6912 ( .A(n6701), .B(n6700), .Z(n6754) );
  XNOR U6913 ( .A(n6753), .B(n6754), .Z(n6755) );
  XOR U6914 ( .A(n6756), .B(n6755), .Z(n6781) );
  XOR U6915 ( .A(n6780), .B(n6781), .Z(n6782) );
  XNOR U6916 ( .A(n6783), .B(n6782), .Z(n6731) );
  NAND U6917 ( .A(n6703), .B(n6702), .Z(n6707) );
  NAND U6918 ( .A(n6705), .B(n6704), .Z(n6706) );
  NAND U6919 ( .A(n6707), .B(n6706), .Z(n6732) );
  XOR U6920 ( .A(n6731), .B(n6732), .Z(n6734) );
  XNOR U6921 ( .A(n6733), .B(n6734), .Z(n6792) );
  NANDN U6922 ( .A(n6709), .B(n6708), .Z(n6713) );
  NAND U6923 ( .A(n6711), .B(n6710), .Z(n6712) );
  NAND U6924 ( .A(n6713), .B(n6712), .Z(n6793) );
  XNOR U6925 ( .A(n6792), .B(n6793), .Z(n6794) );
  XOR U6926 ( .A(n6795), .B(n6794), .Z(n6725) );
  NANDN U6927 ( .A(n6715), .B(n6714), .Z(n6719) );
  NANDN U6928 ( .A(n6717), .B(n6716), .Z(n6718) );
  NAND U6929 ( .A(n6719), .B(n6718), .Z(n6726) );
  XNOR U6930 ( .A(n6725), .B(n6726), .Z(n6727) );
  XNOR U6931 ( .A(n6728), .B(n6727), .Z(n6798) );
  XNOR U6932 ( .A(n6798), .B(sreg[205]), .Z(n6800) );
  NAND U6933 ( .A(n6720), .B(sreg[204]), .Z(n6724) );
  OR U6934 ( .A(n6722), .B(n6721), .Z(n6723) );
  AND U6935 ( .A(n6724), .B(n6723), .Z(n6799) );
  XOR U6936 ( .A(n6800), .B(n6799), .Z(c[205]) );
  NANDN U6937 ( .A(n6726), .B(n6725), .Z(n6730) );
  NAND U6938 ( .A(n6728), .B(n6727), .Z(n6729) );
  NAND U6939 ( .A(n6730), .B(n6729), .Z(n6806) );
  NANDN U6940 ( .A(n6732), .B(n6731), .Z(n6736) );
  OR U6941 ( .A(n6734), .B(n6733), .Z(n6735) );
  NAND U6942 ( .A(n6736), .B(n6735), .Z(n6873) );
  XNOR U6943 ( .A(n9967), .B(n7079), .Z(n6842) );
  OR U6944 ( .A(n6842), .B(n10020), .Z(n6739) );
  NANDN U6945 ( .A(n6737), .B(n9968), .Z(n6738) );
  NAND U6946 ( .A(n6739), .B(n6738), .Z(n6855) );
  XNOR U6947 ( .A(n75), .B(n6740), .Z(n6846) );
  OR U6948 ( .A(n6846), .B(n10106), .Z(n6743) );
  NANDN U6949 ( .A(n6741), .B(n10107), .Z(n6742) );
  NAND U6950 ( .A(n6743), .B(n6742), .Z(n6852) );
  XNOR U6951 ( .A(n9984), .B(n7233), .Z(n6849) );
  NANDN U6952 ( .A(n6849), .B(n9865), .Z(n6746) );
  NANDN U6953 ( .A(n6744), .B(n9930), .Z(n6745) );
  AND U6954 ( .A(n6746), .B(n6745), .Z(n6853) );
  XNOR U6955 ( .A(n6852), .B(n6853), .Z(n6854) );
  XNOR U6956 ( .A(n6855), .B(n6854), .Z(n6864) );
  NANDN U6957 ( .A(n6748), .B(n6747), .Z(n6752) );
  NAND U6958 ( .A(n6750), .B(n6749), .Z(n6751) );
  NAND U6959 ( .A(n6752), .B(n6751), .Z(n6865) );
  XNOR U6960 ( .A(n6864), .B(n6865), .Z(n6866) );
  NANDN U6961 ( .A(n6754), .B(n6753), .Z(n6758) );
  NAND U6962 ( .A(n6756), .B(n6755), .Z(n6757) );
  AND U6963 ( .A(n6758), .B(n6757), .Z(n6867) );
  XNOR U6964 ( .A(n6866), .B(n6867), .Z(n6811) );
  NANDN U6965 ( .A(n6760), .B(n6759), .Z(n6764) );
  OR U6966 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U6967 ( .A(n6764), .B(n6763), .Z(n6839) );
  NAND U6968 ( .A(b[0]), .B(a[94]), .Z(n6765) );
  XNOR U6969 ( .A(b[1]), .B(n6765), .Z(n6767) );
  NAND U6970 ( .A(a[93]), .B(n72), .Z(n6766) );
  AND U6971 ( .A(n6767), .B(n6766), .Z(n6815) );
  XNOR U6972 ( .A(n10050), .B(n6896), .Z(n6824) );
  OR U6973 ( .A(n6824), .B(n10051), .Z(n6770) );
  NANDN U6974 ( .A(n6768), .B(n10070), .Z(n6769) );
  AND U6975 ( .A(n6770), .B(n6769), .Z(n6816) );
  XOR U6976 ( .A(n6815), .B(n6816), .Z(n6818) );
  NAND U6977 ( .A(a[78]), .B(b[15]), .Z(n6817) );
  XOR U6978 ( .A(n6818), .B(n6817), .Z(n6836) );
  XNOR U6979 ( .A(n9622), .B(n7545), .Z(n6827) );
  OR U6980 ( .A(n6827), .B(n9623), .Z(n6773) );
  NANDN U6981 ( .A(n6771), .B(n9680), .Z(n6772) );
  NAND U6982 ( .A(n6773), .B(n6772), .Z(n6861) );
  XNOR U6983 ( .A(n9872), .B(n7389), .Z(n6830) );
  NANDN U6984 ( .A(n6830), .B(n9746), .Z(n6776) );
  NANDN U6985 ( .A(n6774), .B(n9747), .Z(n6775) );
  NAND U6986 ( .A(n6776), .B(n6775), .Z(n6858) );
  IV U6987 ( .A(a[92]), .Z(n7674) );
  XNOR U6988 ( .A(n74), .B(n7674), .Z(n6833) );
  NANDN U6989 ( .A(n6833), .B(n9485), .Z(n6779) );
  NANDN U6990 ( .A(n6777), .B(n9484), .Z(n6778) );
  AND U6991 ( .A(n6779), .B(n6778), .Z(n6859) );
  XNOR U6992 ( .A(n6858), .B(n6859), .Z(n6860) );
  XOR U6993 ( .A(n6861), .B(n6860), .Z(n6837) );
  XOR U6994 ( .A(n6836), .B(n6837), .Z(n6838) );
  XNOR U6995 ( .A(n6839), .B(n6838), .Z(n6809) );
  NAND U6996 ( .A(n6781), .B(n6780), .Z(n6785) );
  NAND U6997 ( .A(n6783), .B(n6782), .Z(n6784) );
  NAND U6998 ( .A(n6785), .B(n6784), .Z(n6810) );
  XOR U6999 ( .A(n6809), .B(n6810), .Z(n6812) );
  XNOR U7000 ( .A(n6811), .B(n6812), .Z(n6870) );
  NANDN U7001 ( .A(n6787), .B(n6786), .Z(n6791) );
  NAND U7002 ( .A(n6789), .B(n6788), .Z(n6790) );
  NAND U7003 ( .A(n6791), .B(n6790), .Z(n6871) );
  XNOR U7004 ( .A(n6870), .B(n6871), .Z(n6872) );
  XOR U7005 ( .A(n6873), .B(n6872), .Z(n6803) );
  NANDN U7006 ( .A(n6793), .B(n6792), .Z(n6797) );
  NANDN U7007 ( .A(n6795), .B(n6794), .Z(n6796) );
  NAND U7008 ( .A(n6797), .B(n6796), .Z(n6804) );
  XNOR U7009 ( .A(n6803), .B(n6804), .Z(n6805) );
  XNOR U7010 ( .A(n6806), .B(n6805), .Z(n6876) );
  XNOR U7011 ( .A(n6876), .B(sreg[206]), .Z(n6878) );
  NAND U7012 ( .A(n6798), .B(sreg[205]), .Z(n6802) );
  OR U7013 ( .A(n6800), .B(n6799), .Z(n6801) );
  AND U7014 ( .A(n6802), .B(n6801), .Z(n6877) );
  XOR U7015 ( .A(n6878), .B(n6877), .Z(c[206]) );
  NANDN U7016 ( .A(n6804), .B(n6803), .Z(n6808) );
  NAND U7017 ( .A(n6806), .B(n6805), .Z(n6807) );
  NAND U7018 ( .A(n6808), .B(n6807), .Z(n6884) );
  NANDN U7019 ( .A(n6810), .B(n6809), .Z(n6814) );
  OR U7020 ( .A(n6812), .B(n6811), .Z(n6813) );
  NAND U7021 ( .A(n6814), .B(n6813), .Z(n6951) );
  NANDN U7022 ( .A(n6816), .B(n6815), .Z(n6820) );
  OR U7023 ( .A(n6818), .B(n6817), .Z(n6819) );
  NAND U7024 ( .A(n6820), .B(n6819), .Z(n6939) );
  NAND U7025 ( .A(b[0]), .B(a[95]), .Z(n6821) );
  XNOR U7026 ( .A(b[1]), .B(n6821), .Z(n6823) );
  NAND U7027 ( .A(a[94]), .B(n72), .Z(n6822) );
  AND U7028 ( .A(n6823), .B(n6822), .Z(n6915) );
  XNOR U7029 ( .A(n10050), .B(n7001), .Z(n6924) );
  OR U7030 ( .A(n6924), .B(n10051), .Z(n6826) );
  NANDN U7031 ( .A(n6824), .B(n10070), .Z(n6825) );
  AND U7032 ( .A(n6826), .B(n6825), .Z(n6916) );
  XOR U7033 ( .A(n6915), .B(n6916), .Z(n6918) );
  NAND U7034 ( .A(a[79]), .B(b[15]), .Z(n6917) );
  XOR U7035 ( .A(n6918), .B(n6917), .Z(n6936) );
  XNOR U7036 ( .A(n9622), .B(n7623), .Z(n6927) );
  OR U7037 ( .A(n6927), .B(n9623), .Z(n6829) );
  NANDN U7038 ( .A(n6827), .B(n9680), .Z(n6828) );
  NAND U7039 ( .A(n6829), .B(n6828), .Z(n6912) );
  XNOR U7040 ( .A(n9872), .B(n7467), .Z(n6930) );
  NANDN U7041 ( .A(n6930), .B(n9746), .Z(n6832) );
  NANDN U7042 ( .A(n6830), .B(n9747), .Z(n6831) );
  NAND U7043 ( .A(n6832), .B(n6831), .Z(n6909) );
  IV U7044 ( .A(a[93]), .Z(n7752) );
  XNOR U7045 ( .A(n74), .B(n7752), .Z(n6933) );
  NANDN U7046 ( .A(n6933), .B(n9485), .Z(n6835) );
  NANDN U7047 ( .A(n6833), .B(n9484), .Z(n6834) );
  AND U7048 ( .A(n6835), .B(n6834), .Z(n6910) );
  XNOR U7049 ( .A(n6909), .B(n6910), .Z(n6911) );
  XOR U7050 ( .A(n6912), .B(n6911), .Z(n6937) );
  XOR U7051 ( .A(n6936), .B(n6937), .Z(n6938) );
  XNOR U7052 ( .A(n6939), .B(n6938), .Z(n6887) );
  NAND U7053 ( .A(n6837), .B(n6836), .Z(n6841) );
  NAND U7054 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U7055 ( .A(n6841), .B(n6840), .Z(n6888) );
  XOR U7056 ( .A(n6887), .B(n6888), .Z(n6890) );
  XNOR U7057 ( .A(n9967), .B(n7155), .Z(n6893) );
  OR U7058 ( .A(n6893), .B(n10020), .Z(n6844) );
  NANDN U7059 ( .A(n6842), .B(n9968), .Z(n6843) );
  NAND U7060 ( .A(n6844), .B(n6843), .Z(n6906) );
  XNOR U7061 ( .A(n75), .B(n6845), .Z(n6897) );
  OR U7062 ( .A(n6897), .B(n10106), .Z(n6848) );
  NANDN U7063 ( .A(n6846), .B(n10107), .Z(n6847) );
  NAND U7064 ( .A(n6848), .B(n6847), .Z(n6903) );
  XNOR U7065 ( .A(n9984), .B(n7284), .Z(n6900) );
  NANDN U7066 ( .A(n6900), .B(n9865), .Z(n6851) );
  NANDN U7067 ( .A(n6849), .B(n9930), .Z(n6850) );
  AND U7068 ( .A(n6851), .B(n6850), .Z(n6904) );
  XNOR U7069 ( .A(n6903), .B(n6904), .Z(n6905) );
  XNOR U7070 ( .A(n6906), .B(n6905), .Z(n6942) );
  NANDN U7071 ( .A(n6853), .B(n6852), .Z(n6857) );
  NAND U7072 ( .A(n6855), .B(n6854), .Z(n6856) );
  NAND U7073 ( .A(n6857), .B(n6856), .Z(n6943) );
  XNOR U7074 ( .A(n6942), .B(n6943), .Z(n6944) );
  NANDN U7075 ( .A(n6859), .B(n6858), .Z(n6863) );
  NAND U7076 ( .A(n6861), .B(n6860), .Z(n6862) );
  AND U7077 ( .A(n6863), .B(n6862), .Z(n6945) );
  XNOR U7078 ( .A(n6944), .B(n6945), .Z(n6889) );
  XNOR U7079 ( .A(n6890), .B(n6889), .Z(n6948) );
  NANDN U7080 ( .A(n6865), .B(n6864), .Z(n6869) );
  NAND U7081 ( .A(n6867), .B(n6866), .Z(n6868) );
  NAND U7082 ( .A(n6869), .B(n6868), .Z(n6949) );
  XNOR U7083 ( .A(n6948), .B(n6949), .Z(n6950) );
  XOR U7084 ( .A(n6951), .B(n6950), .Z(n6881) );
  NANDN U7085 ( .A(n6871), .B(n6870), .Z(n6875) );
  NANDN U7086 ( .A(n6873), .B(n6872), .Z(n6874) );
  NAND U7087 ( .A(n6875), .B(n6874), .Z(n6882) );
  XNOR U7088 ( .A(n6881), .B(n6882), .Z(n6883) );
  XNOR U7089 ( .A(n6884), .B(n6883), .Z(n6954) );
  XNOR U7090 ( .A(n6954), .B(sreg[207]), .Z(n6956) );
  NAND U7091 ( .A(n6876), .B(sreg[206]), .Z(n6880) );
  OR U7092 ( .A(n6878), .B(n6877), .Z(n6879) );
  AND U7093 ( .A(n6880), .B(n6879), .Z(n6955) );
  XOR U7094 ( .A(n6956), .B(n6955), .Z(c[207]) );
  NANDN U7095 ( .A(n6882), .B(n6881), .Z(n6886) );
  NAND U7096 ( .A(n6884), .B(n6883), .Z(n6885) );
  NAND U7097 ( .A(n6886), .B(n6885), .Z(n6962) );
  NANDN U7098 ( .A(n6888), .B(n6887), .Z(n6892) );
  OR U7099 ( .A(n6890), .B(n6889), .Z(n6891) );
  NAND U7100 ( .A(n6892), .B(n6891), .Z(n7029) );
  XNOR U7101 ( .A(n9967), .B(n7233), .Z(n6998) );
  OR U7102 ( .A(n6998), .B(n10020), .Z(n6895) );
  NANDN U7103 ( .A(n6893), .B(n9968), .Z(n6894) );
  NAND U7104 ( .A(n6895), .B(n6894), .Z(n7011) );
  XNOR U7105 ( .A(n75), .B(n6896), .Z(n7002) );
  OR U7106 ( .A(n7002), .B(n10106), .Z(n6899) );
  NANDN U7107 ( .A(n6897), .B(n10107), .Z(n6898) );
  NAND U7108 ( .A(n6899), .B(n6898), .Z(n7008) );
  XNOR U7109 ( .A(n9984), .B(n7389), .Z(n7005) );
  NANDN U7110 ( .A(n7005), .B(n9865), .Z(n6902) );
  NANDN U7111 ( .A(n6900), .B(n9930), .Z(n6901) );
  AND U7112 ( .A(n6902), .B(n6901), .Z(n7009) );
  XNOR U7113 ( .A(n7008), .B(n7009), .Z(n7010) );
  XNOR U7114 ( .A(n7011), .B(n7010), .Z(n7020) );
  NANDN U7115 ( .A(n6904), .B(n6903), .Z(n6908) );
  NAND U7116 ( .A(n6906), .B(n6905), .Z(n6907) );
  NAND U7117 ( .A(n6908), .B(n6907), .Z(n7021) );
  XNOR U7118 ( .A(n7020), .B(n7021), .Z(n7022) );
  NANDN U7119 ( .A(n6910), .B(n6909), .Z(n6914) );
  NAND U7120 ( .A(n6912), .B(n6911), .Z(n6913) );
  AND U7121 ( .A(n6914), .B(n6913), .Z(n7023) );
  XNOR U7122 ( .A(n7022), .B(n7023), .Z(n6967) );
  NANDN U7123 ( .A(n6916), .B(n6915), .Z(n6920) );
  OR U7124 ( .A(n6918), .B(n6917), .Z(n6919) );
  NAND U7125 ( .A(n6920), .B(n6919), .Z(n6995) );
  NAND U7126 ( .A(b[0]), .B(a[96]), .Z(n6921) );
  XNOR U7127 ( .A(b[1]), .B(n6921), .Z(n6923) );
  NAND U7128 ( .A(a[95]), .B(n72), .Z(n6922) );
  AND U7129 ( .A(n6923), .B(n6922), .Z(n6971) );
  XNOR U7130 ( .A(n10050), .B(n7079), .Z(n6977) );
  OR U7131 ( .A(n6977), .B(n10051), .Z(n6926) );
  NANDN U7132 ( .A(n6924), .B(n10070), .Z(n6925) );
  AND U7133 ( .A(n6926), .B(n6925), .Z(n6972) );
  XOR U7134 ( .A(n6971), .B(n6972), .Z(n6974) );
  NAND U7135 ( .A(a[80]), .B(b[15]), .Z(n6973) );
  XOR U7136 ( .A(n6974), .B(n6973), .Z(n6992) );
  XNOR U7137 ( .A(n9622), .B(n7674), .Z(n6983) );
  OR U7138 ( .A(n6983), .B(n9623), .Z(n6929) );
  NANDN U7139 ( .A(n6927), .B(n9680), .Z(n6928) );
  NAND U7140 ( .A(n6929), .B(n6928), .Z(n7017) );
  XNOR U7141 ( .A(n9872), .B(n7545), .Z(n6986) );
  NANDN U7142 ( .A(n6986), .B(n9746), .Z(n6932) );
  NANDN U7143 ( .A(n6930), .B(n9747), .Z(n6931) );
  NAND U7144 ( .A(n6932), .B(n6931), .Z(n7014) );
  IV U7145 ( .A(a[94]), .Z(n7830) );
  XNOR U7146 ( .A(n74), .B(n7830), .Z(n6989) );
  NANDN U7147 ( .A(n6989), .B(n9485), .Z(n6935) );
  NANDN U7148 ( .A(n6933), .B(n9484), .Z(n6934) );
  AND U7149 ( .A(n6935), .B(n6934), .Z(n7015) );
  XNOR U7150 ( .A(n7014), .B(n7015), .Z(n7016) );
  XOR U7151 ( .A(n7017), .B(n7016), .Z(n6993) );
  XOR U7152 ( .A(n6992), .B(n6993), .Z(n6994) );
  XNOR U7153 ( .A(n6995), .B(n6994), .Z(n6965) );
  NAND U7154 ( .A(n6937), .B(n6936), .Z(n6941) );
  NAND U7155 ( .A(n6939), .B(n6938), .Z(n6940) );
  NAND U7156 ( .A(n6941), .B(n6940), .Z(n6966) );
  XOR U7157 ( .A(n6965), .B(n6966), .Z(n6968) );
  XNOR U7158 ( .A(n6967), .B(n6968), .Z(n7026) );
  NANDN U7159 ( .A(n6943), .B(n6942), .Z(n6947) );
  NAND U7160 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND U7161 ( .A(n6947), .B(n6946), .Z(n7027) );
  XNOR U7162 ( .A(n7026), .B(n7027), .Z(n7028) );
  XOR U7163 ( .A(n7029), .B(n7028), .Z(n6959) );
  NANDN U7164 ( .A(n6949), .B(n6948), .Z(n6953) );
  NANDN U7165 ( .A(n6951), .B(n6950), .Z(n6952) );
  NAND U7166 ( .A(n6953), .B(n6952), .Z(n6960) );
  XNOR U7167 ( .A(n6959), .B(n6960), .Z(n6961) );
  XNOR U7168 ( .A(n6962), .B(n6961), .Z(n7032) );
  XNOR U7169 ( .A(n7032), .B(sreg[208]), .Z(n7034) );
  NAND U7170 ( .A(n6954), .B(sreg[207]), .Z(n6958) );
  OR U7171 ( .A(n6956), .B(n6955), .Z(n6957) );
  AND U7172 ( .A(n6958), .B(n6957), .Z(n7033) );
  XOR U7173 ( .A(n7034), .B(n7033), .Z(c[208]) );
  NANDN U7174 ( .A(n6960), .B(n6959), .Z(n6964) );
  NAND U7175 ( .A(n6962), .B(n6961), .Z(n6963) );
  NAND U7176 ( .A(n6964), .B(n6963), .Z(n7040) );
  NANDN U7177 ( .A(n6966), .B(n6965), .Z(n6970) );
  OR U7178 ( .A(n6968), .B(n6967), .Z(n6969) );
  NAND U7179 ( .A(n6970), .B(n6969), .Z(n7107) );
  NANDN U7180 ( .A(n6972), .B(n6971), .Z(n6976) );
  OR U7181 ( .A(n6974), .B(n6973), .Z(n6975) );
  NAND U7182 ( .A(n6976), .B(n6975), .Z(n7073) );
  XNOR U7183 ( .A(n10050), .B(n7155), .Z(n7055) );
  OR U7184 ( .A(n7055), .B(n10051), .Z(n6979) );
  NANDN U7185 ( .A(n6977), .B(n10070), .Z(n6978) );
  AND U7186 ( .A(n6979), .B(n6978), .Z(n7050) );
  NAND U7187 ( .A(b[0]), .B(a[97]), .Z(n6980) );
  XNOR U7188 ( .A(b[1]), .B(n6980), .Z(n6982) );
  NAND U7189 ( .A(a[96]), .B(n72), .Z(n6981) );
  AND U7190 ( .A(n6982), .B(n6981), .Z(n7049) );
  XOR U7191 ( .A(n7050), .B(n7049), .Z(n7052) );
  NAND U7192 ( .A(a[81]), .B(b[15]), .Z(n7051) );
  XOR U7193 ( .A(n7052), .B(n7051), .Z(n7070) );
  XNOR U7194 ( .A(n9622), .B(n7752), .Z(n7061) );
  OR U7195 ( .A(n7061), .B(n9623), .Z(n6985) );
  NANDN U7196 ( .A(n6983), .B(n9680), .Z(n6984) );
  NAND U7197 ( .A(n6985), .B(n6984), .Z(n7095) );
  XNOR U7198 ( .A(n9872), .B(n7623), .Z(n7064) );
  NANDN U7199 ( .A(n7064), .B(n9746), .Z(n6988) );
  NANDN U7200 ( .A(n6986), .B(n9747), .Z(n6987) );
  NAND U7201 ( .A(n6988), .B(n6987), .Z(n7092) );
  IV U7202 ( .A(a[95]), .Z(n7908) );
  XNOR U7203 ( .A(n74), .B(n7908), .Z(n7067) );
  NANDN U7204 ( .A(n7067), .B(n9485), .Z(n6991) );
  NANDN U7205 ( .A(n6989), .B(n9484), .Z(n6990) );
  AND U7206 ( .A(n6991), .B(n6990), .Z(n7093) );
  XNOR U7207 ( .A(n7092), .B(n7093), .Z(n7094) );
  XOR U7208 ( .A(n7095), .B(n7094), .Z(n7071) );
  XOR U7209 ( .A(n7070), .B(n7071), .Z(n7072) );
  XNOR U7210 ( .A(n7073), .B(n7072), .Z(n7043) );
  NAND U7211 ( .A(n6993), .B(n6992), .Z(n6997) );
  NAND U7212 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U7213 ( .A(n6997), .B(n6996), .Z(n7044) );
  XOR U7214 ( .A(n7043), .B(n7044), .Z(n7046) );
  XNOR U7215 ( .A(n9967), .B(n7284), .Z(n7076) );
  OR U7216 ( .A(n7076), .B(n10020), .Z(n7000) );
  NANDN U7217 ( .A(n6998), .B(n9968), .Z(n6999) );
  NAND U7218 ( .A(n7000), .B(n6999), .Z(n7089) );
  XNOR U7219 ( .A(n75), .B(n7001), .Z(n7080) );
  OR U7220 ( .A(n7080), .B(n10106), .Z(n7004) );
  NANDN U7221 ( .A(n7002), .B(n10107), .Z(n7003) );
  NAND U7222 ( .A(n7004), .B(n7003), .Z(n7086) );
  XNOR U7223 ( .A(n9984), .B(n7467), .Z(n7083) );
  NANDN U7224 ( .A(n7083), .B(n9865), .Z(n7007) );
  NANDN U7225 ( .A(n7005), .B(n9930), .Z(n7006) );
  AND U7226 ( .A(n7007), .B(n7006), .Z(n7087) );
  XNOR U7227 ( .A(n7086), .B(n7087), .Z(n7088) );
  XNOR U7228 ( .A(n7089), .B(n7088), .Z(n7098) );
  NANDN U7229 ( .A(n7009), .B(n7008), .Z(n7013) );
  NAND U7230 ( .A(n7011), .B(n7010), .Z(n7012) );
  NAND U7231 ( .A(n7013), .B(n7012), .Z(n7099) );
  XNOR U7232 ( .A(n7098), .B(n7099), .Z(n7100) );
  NANDN U7233 ( .A(n7015), .B(n7014), .Z(n7019) );
  NAND U7234 ( .A(n7017), .B(n7016), .Z(n7018) );
  AND U7235 ( .A(n7019), .B(n7018), .Z(n7101) );
  XNOR U7236 ( .A(n7100), .B(n7101), .Z(n7045) );
  XNOR U7237 ( .A(n7046), .B(n7045), .Z(n7104) );
  NANDN U7238 ( .A(n7021), .B(n7020), .Z(n7025) );
  NAND U7239 ( .A(n7023), .B(n7022), .Z(n7024) );
  NAND U7240 ( .A(n7025), .B(n7024), .Z(n7105) );
  XNOR U7241 ( .A(n7104), .B(n7105), .Z(n7106) );
  XOR U7242 ( .A(n7107), .B(n7106), .Z(n7037) );
  NANDN U7243 ( .A(n7027), .B(n7026), .Z(n7031) );
  NANDN U7244 ( .A(n7029), .B(n7028), .Z(n7030) );
  NAND U7245 ( .A(n7031), .B(n7030), .Z(n7038) );
  XNOR U7246 ( .A(n7037), .B(n7038), .Z(n7039) );
  XNOR U7247 ( .A(n7040), .B(n7039), .Z(n7110) );
  XNOR U7248 ( .A(n7110), .B(sreg[209]), .Z(n7112) );
  NAND U7249 ( .A(n7032), .B(sreg[208]), .Z(n7036) );
  OR U7250 ( .A(n7034), .B(n7033), .Z(n7035) );
  AND U7251 ( .A(n7036), .B(n7035), .Z(n7111) );
  XOR U7252 ( .A(n7112), .B(n7111), .Z(c[209]) );
  NANDN U7253 ( .A(n7038), .B(n7037), .Z(n7042) );
  NAND U7254 ( .A(n7040), .B(n7039), .Z(n7041) );
  NAND U7255 ( .A(n7042), .B(n7041), .Z(n7118) );
  NANDN U7256 ( .A(n7044), .B(n7043), .Z(n7048) );
  OR U7257 ( .A(n7046), .B(n7045), .Z(n7047) );
  NAND U7258 ( .A(n7048), .B(n7047), .Z(n7183) );
  NANDN U7259 ( .A(n7050), .B(n7049), .Z(n7054) );
  OR U7260 ( .A(n7052), .B(n7051), .Z(n7053) );
  NAND U7261 ( .A(n7054), .B(n7053), .Z(n7151) );
  XNOR U7262 ( .A(n10050), .B(n7233), .Z(n7136) );
  OR U7263 ( .A(n7136), .B(n10051), .Z(n7057) );
  NANDN U7264 ( .A(n7055), .B(n10070), .Z(n7056) );
  NAND U7265 ( .A(n7057), .B(n7056), .Z(n7127) );
  AND U7266 ( .A(a[98]), .B(b[0]), .Z(n7058) );
  XOR U7267 ( .A(b[1]), .B(n7058), .Z(n7060) );
  NAND U7268 ( .A(a[97]), .B(n72), .Z(n7059) );
  NAND U7269 ( .A(n7060), .B(n7059), .Z(n7128) );
  XNOR U7270 ( .A(n7127), .B(n7128), .Z(n7129) );
  NAND U7271 ( .A(a[82]), .B(b[15]), .Z(n7130) );
  XOR U7272 ( .A(n7129), .B(n7130), .Z(n7148) );
  XNOR U7273 ( .A(n9622), .B(n7830), .Z(n7139) );
  OR U7274 ( .A(n7139), .B(n9623), .Z(n7063) );
  NANDN U7275 ( .A(n7061), .B(n9680), .Z(n7062) );
  NAND U7276 ( .A(n7063), .B(n7062), .Z(n7171) );
  XNOR U7277 ( .A(n9872), .B(n7674), .Z(n7142) );
  NANDN U7278 ( .A(n7142), .B(n9746), .Z(n7066) );
  NANDN U7279 ( .A(n7064), .B(n9747), .Z(n7065) );
  NAND U7280 ( .A(n7066), .B(n7065), .Z(n7168) );
  IV U7281 ( .A(a[96]), .Z(n7986) );
  XNOR U7282 ( .A(n74), .B(n7986), .Z(n7145) );
  NANDN U7283 ( .A(n7145), .B(n9485), .Z(n7069) );
  NANDN U7284 ( .A(n7067), .B(n9484), .Z(n7068) );
  AND U7285 ( .A(n7069), .B(n7068), .Z(n7169) );
  XNOR U7286 ( .A(n7168), .B(n7169), .Z(n7170) );
  XOR U7287 ( .A(n7171), .B(n7170), .Z(n7149) );
  XNOR U7288 ( .A(n7148), .B(n7149), .Z(n7150) );
  XNOR U7289 ( .A(n7151), .B(n7150), .Z(n7121) );
  NAND U7290 ( .A(n7071), .B(n7070), .Z(n7075) );
  NAND U7291 ( .A(n7073), .B(n7072), .Z(n7074) );
  NAND U7292 ( .A(n7075), .B(n7074), .Z(n7122) );
  XOR U7293 ( .A(n7121), .B(n7122), .Z(n7124) );
  XNOR U7294 ( .A(n9967), .B(n7389), .Z(n7152) );
  OR U7295 ( .A(n7152), .B(n10020), .Z(n7078) );
  NANDN U7296 ( .A(n7076), .B(n9968), .Z(n7077) );
  NAND U7297 ( .A(n7078), .B(n7077), .Z(n7165) );
  XNOR U7298 ( .A(n75), .B(n7079), .Z(n7156) );
  OR U7299 ( .A(n7156), .B(n10106), .Z(n7082) );
  NANDN U7300 ( .A(n7080), .B(n10107), .Z(n7081) );
  NAND U7301 ( .A(n7082), .B(n7081), .Z(n7162) );
  XNOR U7302 ( .A(n9984), .B(n7545), .Z(n7159) );
  NANDN U7303 ( .A(n7159), .B(n9865), .Z(n7085) );
  NANDN U7304 ( .A(n7083), .B(n9930), .Z(n7084) );
  AND U7305 ( .A(n7085), .B(n7084), .Z(n7163) );
  XNOR U7306 ( .A(n7162), .B(n7163), .Z(n7164) );
  XNOR U7307 ( .A(n7165), .B(n7164), .Z(n7174) );
  NANDN U7308 ( .A(n7087), .B(n7086), .Z(n7091) );
  NAND U7309 ( .A(n7089), .B(n7088), .Z(n7090) );
  NAND U7310 ( .A(n7091), .B(n7090), .Z(n7175) );
  XNOR U7311 ( .A(n7174), .B(n7175), .Z(n7176) );
  NANDN U7312 ( .A(n7093), .B(n7092), .Z(n7097) );
  NAND U7313 ( .A(n7095), .B(n7094), .Z(n7096) );
  AND U7314 ( .A(n7097), .B(n7096), .Z(n7177) );
  XNOR U7315 ( .A(n7176), .B(n7177), .Z(n7123) );
  XNOR U7316 ( .A(n7124), .B(n7123), .Z(n7180) );
  NANDN U7317 ( .A(n7099), .B(n7098), .Z(n7103) );
  NAND U7318 ( .A(n7101), .B(n7100), .Z(n7102) );
  NAND U7319 ( .A(n7103), .B(n7102), .Z(n7181) );
  XNOR U7320 ( .A(n7180), .B(n7181), .Z(n7182) );
  XOR U7321 ( .A(n7183), .B(n7182), .Z(n7115) );
  NANDN U7322 ( .A(n7105), .B(n7104), .Z(n7109) );
  NANDN U7323 ( .A(n7107), .B(n7106), .Z(n7108) );
  NAND U7324 ( .A(n7109), .B(n7108), .Z(n7116) );
  XNOR U7325 ( .A(n7115), .B(n7116), .Z(n7117) );
  XNOR U7326 ( .A(n7118), .B(n7117), .Z(n7186) );
  XNOR U7327 ( .A(n7186), .B(sreg[210]), .Z(n7188) );
  NAND U7328 ( .A(n7110), .B(sreg[209]), .Z(n7114) );
  OR U7329 ( .A(n7112), .B(n7111), .Z(n7113) );
  AND U7330 ( .A(n7114), .B(n7113), .Z(n7187) );
  XOR U7331 ( .A(n7188), .B(n7187), .Z(c[210]) );
  NANDN U7332 ( .A(n7116), .B(n7115), .Z(n7120) );
  NAND U7333 ( .A(n7118), .B(n7117), .Z(n7119) );
  NAND U7334 ( .A(n7120), .B(n7119), .Z(n7194) );
  NANDN U7335 ( .A(n7122), .B(n7121), .Z(n7126) );
  OR U7336 ( .A(n7124), .B(n7123), .Z(n7125) );
  NAND U7337 ( .A(n7126), .B(n7125), .Z(n7261) );
  NANDN U7338 ( .A(n7128), .B(n7127), .Z(n7132) );
  NANDN U7339 ( .A(n7130), .B(n7129), .Z(n7131) );
  NAND U7340 ( .A(n7132), .B(n7131), .Z(n7227) );
  NAND U7341 ( .A(b[0]), .B(a[99]), .Z(n7133) );
  XNOR U7342 ( .A(b[1]), .B(n7133), .Z(n7135) );
  NAND U7343 ( .A(a[98]), .B(n72), .Z(n7134) );
  AND U7344 ( .A(n7135), .B(n7134), .Z(n7203) );
  XNOR U7345 ( .A(n10050), .B(n7284), .Z(n7212) );
  OR U7346 ( .A(n7212), .B(n10051), .Z(n7138) );
  NANDN U7347 ( .A(n7136), .B(n10070), .Z(n7137) );
  AND U7348 ( .A(n7138), .B(n7137), .Z(n7204) );
  XOR U7349 ( .A(n7203), .B(n7204), .Z(n7206) );
  NAND U7350 ( .A(a[83]), .B(b[15]), .Z(n7205) );
  XOR U7351 ( .A(n7206), .B(n7205), .Z(n7224) );
  XNOR U7352 ( .A(n9622), .B(n7908), .Z(n7215) );
  OR U7353 ( .A(n7215), .B(n9623), .Z(n7141) );
  NANDN U7354 ( .A(n7139), .B(n9680), .Z(n7140) );
  NAND U7355 ( .A(n7141), .B(n7140), .Z(n7249) );
  XNOR U7356 ( .A(n9872), .B(n7752), .Z(n7218) );
  NANDN U7357 ( .A(n7218), .B(n9746), .Z(n7144) );
  NANDN U7358 ( .A(n7142), .B(n9747), .Z(n7143) );
  NAND U7359 ( .A(n7144), .B(n7143), .Z(n7246) );
  IV U7360 ( .A(a[97]), .Z(n8064) );
  XNOR U7361 ( .A(n74), .B(n8064), .Z(n7221) );
  NANDN U7362 ( .A(n7221), .B(n9485), .Z(n7147) );
  NANDN U7363 ( .A(n7145), .B(n9484), .Z(n7146) );
  AND U7364 ( .A(n7147), .B(n7146), .Z(n7247) );
  XNOR U7365 ( .A(n7246), .B(n7247), .Z(n7248) );
  XOR U7366 ( .A(n7249), .B(n7248), .Z(n7225) );
  XOR U7367 ( .A(n7224), .B(n7225), .Z(n7226) );
  XNOR U7368 ( .A(n7227), .B(n7226), .Z(n7197) );
  XOR U7369 ( .A(n7197), .B(n7198), .Z(n7200) );
  XNOR U7370 ( .A(n9967), .B(n7467), .Z(n7230) );
  OR U7371 ( .A(n7230), .B(n10020), .Z(n7154) );
  NANDN U7372 ( .A(n7152), .B(n9968), .Z(n7153) );
  NAND U7373 ( .A(n7154), .B(n7153), .Z(n7243) );
  XNOR U7374 ( .A(n75), .B(n7155), .Z(n7234) );
  OR U7375 ( .A(n7234), .B(n10106), .Z(n7158) );
  NANDN U7376 ( .A(n7156), .B(n10107), .Z(n7157) );
  NAND U7377 ( .A(n7158), .B(n7157), .Z(n7240) );
  XNOR U7378 ( .A(n9984), .B(n7623), .Z(n7237) );
  NANDN U7379 ( .A(n7237), .B(n9865), .Z(n7161) );
  NANDN U7380 ( .A(n7159), .B(n9930), .Z(n7160) );
  AND U7381 ( .A(n7161), .B(n7160), .Z(n7241) );
  XNOR U7382 ( .A(n7240), .B(n7241), .Z(n7242) );
  XNOR U7383 ( .A(n7243), .B(n7242), .Z(n7252) );
  NANDN U7384 ( .A(n7163), .B(n7162), .Z(n7167) );
  NAND U7385 ( .A(n7165), .B(n7164), .Z(n7166) );
  NAND U7386 ( .A(n7167), .B(n7166), .Z(n7253) );
  XNOR U7387 ( .A(n7252), .B(n7253), .Z(n7254) );
  NANDN U7388 ( .A(n7169), .B(n7168), .Z(n7173) );
  NAND U7389 ( .A(n7171), .B(n7170), .Z(n7172) );
  AND U7390 ( .A(n7173), .B(n7172), .Z(n7255) );
  XNOR U7391 ( .A(n7254), .B(n7255), .Z(n7199) );
  XNOR U7392 ( .A(n7200), .B(n7199), .Z(n7258) );
  NANDN U7393 ( .A(n7175), .B(n7174), .Z(n7179) );
  NAND U7394 ( .A(n7177), .B(n7176), .Z(n7178) );
  NAND U7395 ( .A(n7179), .B(n7178), .Z(n7259) );
  XNOR U7396 ( .A(n7258), .B(n7259), .Z(n7260) );
  XOR U7397 ( .A(n7261), .B(n7260), .Z(n7191) );
  NANDN U7398 ( .A(n7181), .B(n7180), .Z(n7185) );
  NANDN U7399 ( .A(n7183), .B(n7182), .Z(n7184) );
  NAND U7400 ( .A(n7185), .B(n7184), .Z(n7192) );
  XNOR U7401 ( .A(n7191), .B(n7192), .Z(n7193) );
  XNOR U7402 ( .A(n7194), .B(n7193), .Z(n7264) );
  XNOR U7403 ( .A(n7264), .B(sreg[211]), .Z(n7266) );
  NAND U7404 ( .A(n7186), .B(sreg[210]), .Z(n7190) );
  OR U7405 ( .A(n7188), .B(n7187), .Z(n7189) );
  AND U7406 ( .A(n7190), .B(n7189), .Z(n7265) );
  XOR U7407 ( .A(n7266), .B(n7265), .Z(c[211]) );
  NANDN U7408 ( .A(n7192), .B(n7191), .Z(n7196) );
  NAND U7409 ( .A(n7194), .B(n7193), .Z(n7195) );
  NAND U7410 ( .A(n7196), .B(n7195), .Z(n7272) );
  NANDN U7411 ( .A(n7198), .B(n7197), .Z(n7202) );
  OR U7412 ( .A(n7200), .B(n7199), .Z(n7201) );
  NAND U7413 ( .A(n7202), .B(n7201), .Z(n7339) );
  NANDN U7414 ( .A(n7204), .B(n7203), .Z(n7208) );
  OR U7415 ( .A(n7206), .B(n7205), .Z(n7207) );
  NAND U7416 ( .A(n7208), .B(n7207), .Z(n7327) );
  NAND U7417 ( .A(b[0]), .B(a[100]), .Z(n7209) );
  XNOR U7418 ( .A(b[1]), .B(n7209), .Z(n7211) );
  NAND U7419 ( .A(a[99]), .B(n72), .Z(n7210) );
  AND U7420 ( .A(n7211), .B(n7210), .Z(n7303) );
  XNOR U7421 ( .A(n10050), .B(n7389), .Z(n7312) );
  OR U7422 ( .A(n7312), .B(n10051), .Z(n7214) );
  NANDN U7423 ( .A(n7212), .B(n10070), .Z(n7213) );
  AND U7424 ( .A(n7214), .B(n7213), .Z(n7304) );
  XOR U7425 ( .A(n7303), .B(n7304), .Z(n7306) );
  NAND U7426 ( .A(a[84]), .B(b[15]), .Z(n7305) );
  XOR U7427 ( .A(n7306), .B(n7305), .Z(n7324) );
  XNOR U7428 ( .A(n9622), .B(n7986), .Z(n7315) );
  OR U7429 ( .A(n7315), .B(n9623), .Z(n7217) );
  NANDN U7430 ( .A(n7215), .B(n9680), .Z(n7216) );
  NAND U7431 ( .A(n7217), .B(n7216), .Z(n7300) );
  XNOR U7432 ( .A(n9872), .B(n7830), .Z(n7318) );
  NANDN U7433 ( .A(n7318), .B(n9746), .Z(n7220) );
  NANDN U7434 ( .A(n7218), .B(n9747), .Z(n7219) );
  NAND U7435 ( .A(n7220), .B(n7219), .Z(n7297) );
  IV U7436 ( .A(a[98]), .Z(n8169) );
  XNOR U7437 ( .A(n74), .B(n8169), .Z(n7321) );
  NANDN U7438 ( .A(n7321), .B(n9485), .Z(n7223) );
  NANDN U7439 ( .A(n7221), .B(n9484), .Z(n7222) );
  AND U7440 ( .A(n7223), .B(n7222), .Z(n7298) );
  XNOR U7441 ( .A(n7297), .B(n7298), .Z(n7299) );
  XOR U7442 ( .A(n7300), .B(n7299), .Z(n7325) );
  XOR U7443 ( .A(n7324), .B(n7325), .Z(n7326) );
  XNOR U7444 ( .A(n7327), .B(n7326), .Z(n7275) );
  NAND U7445 ( .A(n7225), .B(n7224), .Z(n7229) );
  NAND U7446 ( .A(n7227), .B(n7226), .Z(n7228) );
  NAND U7447 ( .A(n7229), .B(n7228), .Z(n7276) );
  XOR U7448 ( .A(n7275), .B(n7276), .Z(n7278) );
  XNOR U7449 ( .A(n9967), .B(n7545), .Z(n7281) );
  OR U7450 ( .A(n7281), .B(n10020), .Z(n7232) );
  NANDN U7451 ( .A(n7230), .B(n9968), .Z(n7231) );
  NAND U7452 ( .A(n7232), .B(n7231), .Z(n7294) );
  XNOR U7453 ( .A(n75), .B(n7233), .Z(n7285) );
  OR U7454 ( .A(n7285), .B(n10106), .Z(n7236) );
  NANDN U7455 ( .A(n7234), .B(n10107), .Z(n7235) );
  NAND U7456 ( .A(n7236), .B(n7235), .Z(n7291) );
  XNOR U7457 ( .A(n9984), .B(n7674), .Z(n7288) );
  NANDN U7458 ( .A(n7288), .B(n9865), .Z(n7239) );
  NANDN U7459 ( .A(n7237), .B(n9930), .Z(n7238) );
  AND U7460 ( .A(n7239), .B(n7238), .Z(n7292) );
  XNOR U7461 ( .A(n7291), .B(n7292), .Z(n7293) );
  XNOR U7462 ( .A(n7294), .B(n7293), .Z(n7330) );
  NANDN U7463 ( .A(n7241), .B(n7240), .Z(n7245) );
  NAND U7464 ( .A(n7243), .B(n7242), .Z(n7244) );
  NAND U7465 ( .A(n7245), .B(n7244), .Z(n7331) );
  XNOR U7466 ( .A(n7330), .B(n7331), .Z(n7332) );
  NANDN U7467 ( .A(n7247), .B(n7246), .Z(n7251) );
  NAND U7468 ( .A(n7249), .B(n7248), .Z(n7250) );
  AND U7469 ( .A(n7251), .B(n7250), .Z(n7333) );
  XNOR U7470 ( .A(n7332), .B(n7333), .Z(n7277) );
  XNOR U7471 ( .A(n7278), .B(n7277), .Z(n7336) );
  NANDN U7472 ( .A(n7253), .B(n7252), .Z(n7257) );
  NAND U7473 ( .A(n7255), .B(n7254), .Z(n7256) );
  NAND U7474 ( .A(n7257), .B(n7256), .Z(n7337) );
  XNOR U7475 ( .A(n7336), .B(n7337), .Z(n7338) );
  XOR U7476 ( .A(n7339), .B(n7338), .Z(n7269) );
  NANDN U7477 ( .A(n7259), .B(n7258), .Z(n7263) );
  NANDN U7478 ( .A(n7261), .B(n7260), .Z(n7262) );
  NAND U7479 ( .A(n7263), .B(n7262), .Z(n7270) );
  XNOR U7480 ( .A(n7269), .B(n7270), .Z(n7271) );
  XNOR U7481 ( .A(n7272), .B(n7271), .Z(n7342) );
  XNOR U7482 ( .A(n7342), .B(sreg[212]), .Z(n7344) );
  NAND U7483 ( .A(n7264), .B(sreg[211]), .Z(n7268) );
  OR U7484 ( .A(n7266), .B(n7265), .Z(n7267) );
  AND U7485 ( .A(n7268), .B(n7267), .Z(n7343) );
  XOR U7486 ( .A(n7344), .B(n7343), .Z(c[212]) );
  NANDN U7487 ( .A(n7270), .B(n7269), .Z(n7274) );
  NAND U7488 ( .A(n7272), .B(n7271), .Z(n7273) );
  NAND U7489 ( .A(n7274), .B(n7273), .Z(n7350) );
  NANDN U7490 ( .A(n7276), .B(n7275), .Z(n7280) );
  OR U7491 ( .A(n7278), .B(n7277), .Z(n7279) );
  NAND U7492 ( .A(n7280), .B(n7279), .Z(n7417) );
  XNOR U7493 ( .A(n9967), .B(n7623), .Z(n7386) );
  OR U7494 ( .A(n7386), .B(n10020), .Z(n7283) );
  NANDN U7495 ( .A(n7281), .B(n9968), .Z(n7282) );
  NAND U7496 ( .A(n7283), .B(n7282), .Z(n7399) );
  XNOR U7497 ( .A(n75), .B(n7284), .Z(n7390) );
  OR U7498 ( .A(n7390), .B(n10106), .Z(n7287) );
  NANDN U7499 ( .A(n7285), .B(n10107), .Z(n7286) );
  NAND U7500 ( .A(n7287), .B(n7286), .Z(n7396) );
  XNOR U7501 ( .A(n9984), .B(n7752), .Z(n7393) );
  NANDN U7502 ( .A(n7393), .B(n9865), .Z(n7290) );
  NANDN U7503 ( .A(n7288), .B(n9930), .Z(n7289) );
  AND U7504 ( .A(n7290), .B(n7289), .Z(n7397) );
  XNOR U7505 ( .A(n7396), .B(n7397), .Z(n7398) );
  XNOR U7506 ( .A(n7399), .B(n7398), .Z(n7408) );
  NANDN U7507 ( .A(n7292), .B(n7291), .Z(n7296) );
  NAND U7508 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U7509 ( .A(n7296), .B(n7295), .Z(n7409) );
  XNOR U7510 ( .A(n7408), .B(n7409), .Z(n7410) );
  NANDN U7511 ( .A(n7298), .B(n7297), .Z(n7302) );
  NAND U7512 ( .A(n7300), .B(n7299), .Z(n7301) );
  AND U7513 ( .A(n7302), .B(n7301), .Z(n7411) );
  XNOR U7514 ( .A(n7410), .B(n7411), .Z(n7355) );
  NANDN U7515 ( .A(n7304), .B(n7303), .Z(n7308) );
  OR U7516 ( .A(n7306), .B(n7305), .Z(n7307) );
  NAND U7517 ( .A(n7308), .B(n7307), .Z(n7383) );
  NAND U7518 ( .A(b[0]), .B(a[101]), .Z(n7309) );
  XNOR U7519 ( .A(b[1]), .B(n7309), .Z(n7311) );
  NAND U7520 ( .A(a[100]), .B(n72), .Z(n7310) );
  AND U7521 ( .A(n7311), .B(n7310), .Z(n7359) );
  XNOR U7522 ( .A(n10050), .B(n7467), .Z(n7365) );
  OR U7523 ( .A(n7365), .B(n10051), .Z(n7314) );
  NANDN U7524 ( .A(n7312), .B(n10070), .Z(n7313) );
  AND U7525 ( .A(n7314), .B(n7313), .Z(n7360) );
  XOR U7526 ( .A(n7359), .B(n7360), .Z(n7362) );
  NAND U7527 ( .A(a[85]), .B(b[15]), .Z(n7361) );
  XOR U7528 ( .A(n7362), .B(n7361), .Z(n7380) );
  XNOR U7529 ( .A(n9622), .B(n8064), .Z(n7371) );
  OR U7530 ( .A(n7371), .B(n9623), .Z(n7317) );
  NANDN U7531 ( .A(n7315), .B(n9680), .Z(n7316) );
  NAND U7532 ( .A(n7317), .B(n7316), .Z(n7405) );
  XNOR U7533 ( .A(n9872), .B(n7908), .Z(n7374) );
  NANDN U7534 ( .A(n7374), .B(n9746), .Z(n7320) );
  NANDN U7535 ( .A(n7318), .B(n9747), .Z(n7319) );
  NAND U7536 ( .A(n7320), .B(n7319), .Z(n7402) );
  IV U7537 ( .A(a[99]), .Z(n8220) );
  XNOR U7538 ( .A(n74), .B(n8220), .Z(n7377) );
  NANDN U7539 ( .A(n7377), .B(n9485), .Z(n7323) );
  NANDN U7540 ( .A(n7321), .B(n9484), .Z(n7322) );
  AND U7541 ( .A(n7323), .B(n7322), .Z(n7403) );
  XNOR U7542 ( .A(n7402), .B(n7403), .Z(n7404) );
  XOR U7543 ( .A(n7405), .B(n7404), .Z(n7381) );
  XOR U7544 ( .A(n7380), .B(n7381), .Z(n7382) );
  XNOR U7545 ( .A(n7383), .B(n7382), .Z(n7353) );
  NAND U7546 ( .A(n7325), .B(n7324), .Z(n7329) );
  NAND U7547 ( .A(n7327), .B(n7326), .Z(n7328) );
  NAND U7548 ( .A(n7329), .B(n7328), .Z(n7354) );
  XOR U7549 ( .A(n7353), .B(n7354), .Z(n7356) );
  XNOR U7550 ( .A(n7355), .B(n7356), .Z(n7414) );
  NANDN U7551 ( .A(n7331), .B(n7330), .Z(n7335) );
  NAND U7552 ( .A(n7333), .B(n7332), .Z(n7334) );
  NAND U7553 ( .A(n7335), .B(n7334), .Z(n7415) );
  XNOR U7554 ( .A(n7414), .B(n7415), .Z(n7416) );
  XOR U7555 ( .A(n7417), .B(n7416), .Z(n7347) );
  NANDN U7556 ( .A(n7337), .B(n7336), .Z(n7341) );
  NANDN U7557 ( .A(n7339), .B(n7338), .Z(n7340) );
  NAND U7558 ( .A(n7341), .B(n7340), .Z(n7348) );
  XNOR U7559 ( .A(n7347), .B(n7348), .Z(n7349) );
  XNOR U7560 ( .A(n7350), .B(n7349), .Z(n7420) );
  XNOR U7561 ( .A(n7420), .B(sreg[213]), .Z(n7422) );
  NAND U7562 ( .A(n7342), .B(sreg[212]), .Z(n7346) );
  OR U7563 ( .A(n7344), .B(n7343), .Z(n7345) );
  AND U7564 ( .A(n7346), .B(n7345), .Z(n7421) );
  XOR U7565 ( .A(n7422), .B(n7421), .Z(c[213]) );
  NANDN U7566 ( .A(n7348), .B(n7347), .Z(n7352) );
  NAND U7567 ( .A(n7350), .B(n7349), .Z(n7351) );
  NAND U7568 ( .A(n7352), .B(n7351), .Z(n7428) );
  NANDN U7569 ( .A(n7354), .B(n7353), .Z(n7358) );
  OR U7570 ( .A(n7356), .B(n7355), .Z(n7357) );
  NAND U7571 ( .A(n7358), .B(n7357), .Z(n7495) );
  NANDN U7572 ( .A(n7360), .B(n7359), .Z(n7364) );
  OR U7573 ( .A(n7362), .B(n7361), .Z(n7363) );
  NAND U7574 ( .A(n7364), .B(n7363), .Z(n7461) );
  XNOR U7575 ( .A(n10050), .B(n7545), .Z(n7446) );
  OR U7576 ( .A(n7446), .B(n10051), .Z(n7367) );
  NANDN U7577 ( .A(n7365), .B(n10070), .Z(n7366) );
  AND U7578 ( .A(n7367), .B(n7366), .Z(n7438) );
  NAND U7579 ( .A(b[0]), .B(a[102]), .Z(n7368) );
  XNOR U7580 ( .A(b[1]), .B(n7368), .Z(n7370) );
  NAND U7581 ( .A(a[101]), .B(n72), .Z(n7369) );
  AND U7582 ( .A(n7370), .B(n7369), .Z(n7437) );
  XOR U7583 ( .A(n7438), .B(n7437), .Z(n7440) );
  NAND U7584 ( .A(a[86]), .B(b[15]), .Z(n7439) );
  XOR U7585 ( .A(n7440), .B(n7439), .Z(n7458) );
  XNOR U7586 ( .A(n9622), .B(n8169), .Z(n7449) );
  OR U7587 ( .A(n7449), .B(n9623), .Z(n7373) );
  NANDN U7588 ( .A(n7371), .B(n9680), .Z(n7372) );
  NAND U7589 ( .A(n7373), .B(n7372), .Z(n7483) );
  XNOR U7590 ( .A(n9872), .B(n7986), .Z(n7452) );
  NANDN U7591 ( .A(n7452), .B(n9746), .Z(n7376) );
  NANDN U7592 ( .A(n7374), .B(n9747), .Z(n7375) );
  NAND U7593 ( .A(n7376), .B(n7375), .Z(n7480) );
  IV U7594 ( .A(a[100]), .Z(n8298) );
  XNOR U7595 ( .A(n74), .B(n8298), .Z(n7455) );
  NANDN U7596 ( .A(n7455), .B(n9485), .Z(n7379) );
  NANDN U7597 ( .A(n7377), .B(n9484), .Z(n7378) );
  AND U7598 ( .A(n7379), .B(n7378), .Z(n7481) );
  XNOR U7599 ( .A(n7480), .B(n7481), .Z(n7482) );
  XOR U7600 ( .A(n7483), .B(n7482), .Z(n7459) );
  XOR U7601 ( .A(n7458), .B(n7459), .Z(n7460) );
  XNOR U7602 ( .A(n7461), .B(n7460), .Z(n7431) );
  NAND U7603 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U7604 ( .A(n7383), .B(n7382), .Z(n7384) );
  NAND U7605 ( .A(n7385), .B(n7384), .Z(n7432) );
  XOR U7606 ( .A(n7431), .B(n7432), .Z(n7434) );
  XNOR U7607 ( .A(n9967), .B(n7674), .Z(n7464) );
  OR U7608 ( .A(n7464), .B(n10020), .Z(n7388) );
  NANDN U7609 ( .A(n7386), .B(n9968), .Z(n7387) );
  NAND U7610 ( .A(n7388), .B(n7387), .Z(n7477) );
  XNOR U7611 ( .A(n75), .B(n7389), .Z(n7468) );
  OR U7612 ( .A(n7468), .B(n10106), .Z(n7392) );
  NANDN U7613 ( .A(n7390), .B(n10107), .Z(n7391) );
  NAND U7614 ( .A(n7392), .B(n7391), .Z(n7474) );
  XNOR U7615 ( .A(n9984), .B(n7830), .Z(n7471) );
  NANDN U7616 ( .A(n7471), .B(n9865), .Z(n7395) );
  NANDN U7617 ( .A(n7393), .B(n9930), .Z(n7394) );
  AND U7618 ( .A(n7395), .B(n7394), .Z(n7475) );
  XNOR U7619 ( .A(n7474), .B(n7475), .Z(n7476) );
  XNOR U7620 ( .A(n7477), .B(n7476), .Z(n7486) );
  NANDN U7621 ( .A(n7397), .B(n7396), .Z(n7401) );
  NAND U7622 ( .A(n7399), .B(n7398), .Z(n7400) );
  NAND U7623 ( .A(n7401), .B(n7400), .Z(n7487) );
  XNOR U7624 ( .A(n7486), .B(n7487), .Z(n7488) );
  NANDN U7625 ( .A(n7403), .B(n7402), .Z(n7407) );
  NAND U7626 ( .A(n7405), .B(n7404), .Z(n7406) );
  AND U7627 ( .A(n7407), .B(n7406), .Z(n7489) );
  XNOR U7628 ( .A(n7488), .B(n7489), .Z(n7433) );
  XNOR U7629 ( .A(n7434), .B(n7433), .Z(n7492) );
  NANDN U7630 ( .A(n7409), .B(n7408), .Z(n7413) );
  NAND U7631 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U7632 ( .A(n7413), .B(n7412), .Z(n7493) );
  XNOR U7633 ( .A(n7492), .B(n7493), .Z(n7494) );
  XOR U7634 ( .A(n7495), .B(n7494), .Z(n7425) );
  NANDN U7635 ( .A(n7415), .B(n7414), .Z(n7419) );
  NANDN U7636 ( .A(n7417), .B(n7416), .Z(n7418) );
  NAND U7637 ( .A(n7419), .B(n7418), .Z(n7426) );
  XNOR U7638 ( .A(n7425), .B(n7426), .Z(n7427) );
  XNOR U7639 ( .A(n7428), .B(n7427), .Z(n7498) );
  XNOR U7640 ( .A(n7498), .B(sreg[214]), .Z(n7500) );
  NAND U7641 ( .A(n7420), .B(sreg[213]), .Z(n7424) );
  OR U7642 ( .A(n7422), .B(n7421), .Z(n7423) );
  AND U7643 ( .A(n7424), .B(n7423), .Z(n7499) );
  XOR U7644 ( .A(n7500), .B(n7499), .Z(c[214]) );
  NANDN U7645 ( .A(n7426), .B(n7425), .Z(n7430) );
  NAND U7646 ( .A(n7428), .B(n7427), .Z(n7429) );
  NAND U7647 ( .A(n7430), .B(n7429), .Z(n7506) );
  NANDN U7648 ( .A(n7432), .B(n7431), .Z(n7436) );
  OR U7649 ( .A(n7434), .B(n7433), .Z(n7435) );
  NAND U7650 ( .A(n7436), .B(n7435), .Z(n7573) );
  NANDN U7651 ( .A(n7438), .B(n7437), .Z(n7442) );
  OR U7652 ( .A(n7440), .B(n7439), .Z(n7441) );
  NAND U7653 ( .A(n7442), .B(n7441), .Z(n7539) );
  NAND U7654 ( .A(b[0]), .B(a[103]), .Z(n7443) );
  XNOR U7655 ( .A(b[1]), .B(n7443), .Z(n7445) );
  NAND U7656 ( .A(a[102]), .B(n72), .Z(n7444) );
  AND U7657 ( .A(n7445), .B(n7444), .Z(n7515) );
  XNOR U7658 ( .A(n10050), .B(n7623), .Z(n7524) );
  OR U7659 ( .A(n7524), .B(n10051), .Z(n7448) );
  NANDN U7660 ( .A(n7446), .B(n10070), .Z(n7447) );
  AND U7661 ( .A(n7448), .B(n7447), .Z(n7516) );
  XOR U7662 ( .A(n7515), .B(n7516), .Z(n7518) );
  NAND U7663 ( .A(a[87]), .B(b[15]), .Z(n7517) );
  XOR U7664 ( .A(n7518), .B(n7517), .Z(n7536) );
  XNOR U7665 ( .A(n9622), .B(n8220), .Z(n7527) );
  OR U7666 ( .A(n7527), .B(n9623), .Z(n7451) );
  NANDN U7667 ( .A(n7449), .B(n9680), .Z(n7450) );
  NAND U7668 ( .A(n7451), .B(n7450), .Z(n7561) );
  XNOR U7669 ( .A(n9872), .B(n8064), .Z(n7530) );
  NANDN U7670 ( .A(n7530), .B(n9746), .Z(n7454) );
  NANDN U7671 ( .A(n7452), .B(n9747), .Z(n7453) );
  NAND U7672 ( .A(n7454), .B(n7453), .Z(n7558) );
  IV U7673 ( .A(a[101]), .Z(n8376) );
  XNOR U7674 ( .A(n74), .B(n8376), .Z(n7533) );
  NANDN U7675 ( .A(n7533), .B(n9485), .Z(n7457) );
  NANDN U7676 ( .A(n7455), .B(n9484), .Z(n7456) );
  AND U7677 ( .A(n7457), .B(n7456), .Z(n7559) );
  XNOR U7678 ( .A(n7558), .B(n7559), .Z(n7560) );
  XOR U7679 ( .A(n7561), .B(n7560), .Z(n7537) );
  XOR U7680 ( .A(n7536), .B(n7537), .Z(n7538) );
  XNOR U7681 ( .A(n7539), .B(n7538), .Z(n7509) );
  NAND U7682 ( .A(n7459), .B(n7458), .Z(n7463) );
  NAND U7683 ( .A(n7461), .B(n7460), .Z(n7462) );
  NAND U7684 ( .A(n7463), .B(n7462), .Z(n7510) );
  XOR U7685 ( .A(n7509), .B(n7510), .Z(n7512) );
  XNOR U7686 ( .A(n9967), .B(n7752), .Z(n7542) );
  OR U7687 ( .A(n7542), .B(n10020), .Z(n7466) );
  NANDN U7688 ( .A(n7464), .B(n9968), .Z(n7465) );
  NAND U7689 ( .A(n7466), .B(n7465), .Z(n7555) );
  XNOR U7690 ( .A(n75), .B(n7467), .Z(n7546) );
  OR U7691 ( .A(n7546), .B(n10106), .Z(n7470) );
  NANDN U7692 ( .A(n7468), .B(n10107), .Z(n7469) );
  NAND U7693 ( .A(n7470), .B(n7469), .Z(n7552) );
  XNOR U7694 ( .A(n9984), .B(n7908), .Z(n7549) );
  NANDN U7695 ( .A(n7549), .B(n9865), .Z(n7473) );
  NANDN U7696 ( .A(n7471), .B(n9930), .Z(n7472) );
  AND U7697 ( .A(n7473), .B(n7472), .Z(n7553) );
  XNOR U7698 ( .A(n7552), .B(n7553), .Z(n7554) );
  XNOR U7699 ( .A(n7555), .B(n7554), .Z(n7564) );
  NANDN U7700 ( .A(n7475), .B(n7474), .Z(n7479) );
  NAND U7701 ( .A(n7477), .B(n7476), .Z(n7478) );
  NAND U7702 ( .A(n7479), .B(n7478), .Z(n7565) );
  XNOR U7703 ( .A(n7564), .B(n7565), .Z(n7566) );
  NANDN U7704 ( .A(n7481), .B(n7480), .Z(n7485) );
  NAND U7705 ( .A(n7483), .B(n7482), .Z(n7484) );
  AND U7706 ( .A(n7485), .B(n7484), .Z(n7567) );
  XNOR U7707 ( .A(n7566), .B(n7567), .Z(n7511) );
  XNOR U7708 ( .A(n7512), .B(n7511), .Z(n7570) );
  NANDN U7709 ( .A(n7487), .B(n7486), .Z(n7491) );
  NAND U7710 ( .A(n7489), .B(n7488), .Z(n7490) );
  NAND U7711 ( .A(n7491), .B(n7490), .Z(n7571) );
  XNOR U7712 ( .A(n7570), .B(n7571), .Z(n7572) );
  XOR U7713 ( .A(n7573), .B(n7572), .Z(n7503) );
  NANDN U7714 ( .A(n7493), .B(n7492), .Z(n7497) );
  NANDN U7715 ( .A(n7495), .B(n7494), .Z(n7496) );
  NAND U7716 ( .A(n7497), .B(n7496), .Z(n7504) );
  XNOR U7717 ( .A(n7503), .B(n7504), .Z(n7505) );
  XNOR U7718 ( .A(n7506), .B(n7505), .Z(n7576) );
  XNOR U7719 ( .A(n7576), .B(sreg[215]), .Z(n7578) );
  NAND U7720 ( .A(n7498), .B(sreg[214]), .Z(n7502) );
  OR U7721 ( .A(n7500), .B(n7499), .Z(n7501) );
  AND U7722 ( .A(n7502), .B(n7501), .Z(n7577) );
  XOR U7723 ( .A(n7578), .B(n7577), .Z(c[215]) );
  NANDN U7724 ( .A(n7504), .B(n7503), .Z(n7508) );
  NAND U7725 ( .A(n7506), .B(n7505), .Z(n7507) );
  NAND U7726 ( .A(n7508), .B(n7507), .Z(n7584) );
  NANDN U7727 ( .A(n7510), .B(n7509), .Z(n7514) );
  OR U7728 ( .A(n7512), .B(n7511), .Z(n7513) );
  NAND U7729 ( .A(n7514), .B(n7513), .Z(n7651) );
  NANDN U7730 ( .A(n7516), .B(n7515), .Z(n7520) );
  OR U7731 ( .A(n7518), .B(n7517), .Z(n7519) );
  NAND U7732 ( .A(n7520), .B(n7519), .Z(n7617) );
  NAND U7733 ( .A(b[0]), .B(a[104]), .Z(n7521) );
  XNOR U7734 ( .A(b[1]), .B(n7521), .Z(n7523) );
  NAND U7735 ( .A(a[103]), .B(n72), .Z(n7522) );
  AND U7736 ( .A(n7523), .B(n7522), .Z(n7593) );
  XNOR U7737 ( .A(n10050), .B(n7674), .Z(n7599) );
  OR U7738 ( .A(n7599), .B(n10051), .Z(n7526) );
  NANDN U7739 ( .A(n7524), .B(n10070), .Z(n7525) );
  AND U7740 ( .A(n7526), .B(n7525), .Z(n7594) );
  XOR U7741 ( .A(n7593), .B(n7594), .Z(n7596) );
  NAND U7742 ( .A(a[88]), .B(b[15]), .Z(n7595) );
  XOR U7743 ( .A(n7596), .B(n7595), .Z(n7614) );
  XNOR U7744 ( .A(n9622), .B(n8298), .Z(n7605) );
  OR U7745 ( .A(n7605), .B(n9623), .Z(n7529) );
  NANDN U7746 ( .A(n7527), .B(n9680), .Z(n7528) );
  NAND U7747 ( .A(n7529), .B(n7528), .Z(n7639) );
  XNOR U7748 ( .A(n9872), .B(n8169), .Z(n7608) );
  NANDN U7749 ( .A(n7608), .B(n9746), .Z(n7532) );
  NANDN U7750 ( .A(n7530), .B(n9747), .Z(n7531) );
  NAND U7751 ( .A(n7532), .B(n7531), .Z(n7636) );
  IV U7752 ( .A(a[102]), .Z(n8481) );
  XNOR U7753 ( .A(n74), .B(n8481), .Z(n7611) );
  NANDN U7754 ( .A(n7611), .B(n9485), .Z(n7535) );
  NANDN U7755 ( .A(n7533), .B(n9484), .Z(n7534) );
  AND U7756 ( .A(n7535), .B(n7534), .Z(n7637) );
  XNOR U7757 ( .A(n7636), .B(n7637), .Z(n7638) );
  XOR U7758 ( .A(n7639), .B(n7638), .Z(n7615) );
  XOR U7759 ( .A(n7614), .B(n7615), .Z(n7616) );
  XNOR U7760 ( .A(n7617), .B(n7616), .Z(n7587) );
  NAND U7761 ( .A(n7537), .B(n7536), .Z(n7541) );
  NAND U7762 ( .A(n7539), .B(n7538), .Z(n7540) );
  NAND U7763 ( .A(n7541), .B(n7540), .Z(n7588) );
  XOR U7764 ( .A(n7587), .B(n7588), .Z(n7590) );
  XNOR U7765 ( .A(n9967), .B(n7830), .Z(n7620) );
  OR U7766 ( .A(n7620), .B(n10020), .Z(n7544) );
  NANDN U7767 ( .A(n7542), .B(n9968), .Z(n7543) );
  NAND U7768 ( .A(n7544), .B(n7543), .Z(n7633) );
  XNOR U7769 ( .A(n75), .B(n7545), .Z(n7624) );
  OR U7770 ( .A(n7624), .B(n10106), .Z(n7548) );
  NANDN U7771 ( .A(n7546), .B(n10107), .Z(n7547) );
  NAND U7772 ( .A(n7548), .B(n7547), .Z(n7630) );
  XNOR U7773 ( .A(n9984), .B(n7986), .Z(n7627) );
  NANDN U7774 ( .A(n7627), .B(n9865), .Z(n7551) );
  NANDN U7775 ( .A(n7549), .B(n9930), .Z(n7550) );
  AND U7776 ( .A(n7551), .B(n7550), .Z(n7631) );
  XNOR U7777 ( .A(n7630), .B(n7631), .Z(n7632) );
  XNOR U7778 ( .A(n7633), .B(n7632), .Z(n7642) );
  NANDN U7779 ( .A(n7553), .B(n7552), .Z(n7557) );
  NAND U7780 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U7781 ( .A(n7557), .B(n7556), .Z(n7643) );
  XNOR U7782 ( .A(n7642), .B(n7643), .Z(n7644) );
  NANDN U7783 ( .A(n7559), .B(n7558), .Z(n7563) );
  NAND U7784 ( .A(n7561), .B(n7560), .Z(n7562) );
  AND U7785 ( .A(n7563), .B(n7562), .Z(n7645) );
  XNOR U7786 ( .A(n7644), .B(n7645), .Z(n7589) );
  XNOR U7787 ( .A(n7590), .B(n7589), .Z(n7648) );
  NANDN U7788 ( .A(n7565), .B(n7564), .Z(n7569) );
  NAND U7789 ( .A(n7567), .B(n7566), .Z(n7568) );
  NAND U7790 ( .A(n7569), .B(n7568), .Z(n7649) );
  XNOR U7791 ( .A(n7648), .B(n7649), .Z(n7650) );
  XOR U7792 ( .A(n7651), .B(n7650), .Z(n7581) );
  NANDN U7793 ( .A(n7571), .B(n7570), .Z(n7575) );
  NANDN U7794 ( .A(n7573), .B(n7572), .Z(n7574) );
  NAND U7795 ( .A(n7575), .B(n7574), .Z(n7582) );
  XNOR U7796 ( .A(n7581), .B(n7582), .Z(n7583) );
  XNOR U7797 ( .A(n7584), .B(n7583), .Z(n7654) );
  XNOR U7798 ( .A(n7654), .B(sreg[216]), .Z(n7656) );
  NAND U7799 ( .A(n7576), .B(sreg[215]), .Z(n7580) );
  OR U7800 ( .A(n7578), .B(n7577), .Z(n7579) );
  AND U7801 ( .A(n7580), .B(n7579), .Z(n7655) );
  XOR U7802 ( .A(n7656), .B(n7655), .Z(c[216]) );
  NANDN U7803 ( .A(n7582), .B(n7581), .Z(n7586) );
  NAND U7804 ( .A(n7584), .B(n7583), .Z(n7585) );
  NAND U7805 ( .A(n7586), .B(n7585), .Z(n7662) );
  NANDN U7806 ( .A(n7588), .B(n7587), .Z(n7592) );
  OR U7807 ( .A(n7590), .B(n7589), .Z(n7591) );
  NAND U7808 ( .A(n7592), .B(n7591), .Z(n7729) );
  NANDN U7809 ( .A(n7594), .B(n7593), .Z(n7598) );
  OR U7810 ( .A(n7596), .B(n7595), .Z(n7597) );
  NAND U7811 ( .A(n7598), .B(n7597), .Z(n7717) );
  XNOR U7812 ( .A(n10050), .B(n7752), .Z(n7702) );
  OR U7813 ( .A(n7702), .B(n10051), .Z(n7601) );
  NANDN U7814 ( .A(n7599), .B(n10070), .Z(n7600) );
  AND U7815 ( .A(n7601), .B(n7600), .Z(n7694) );
  NAND U7816 ( .A(b[0]), .B(a[105]), .Z(n7602) );
  XNOR U7817 ( .A(b[1]), .B(n7602), .Z(n7604) );
  NAND U7818 ( .A(a[104]), .B(n72), .Z(n7603) );
  AND U7819 ( .A(n7604), .B(n7603), .Z(n7693) );
  XOR U7820 ( .A(n7694), .B(n7693), .Z(n7696) );
  NAND U7821 ( .A(a[89]), .B(b[15]), .Z(n7695) );
  XOR U7822 ( .A(n7696), .B(n7695), .Z(n7714) );
  XNOR U7823 ( .A(n9622), .B(n8376), .Z(n7705) );
  OR U7824 ( .A(n7705), .B(n9623), .Z(n7607) );
  NANDN U7825 ( .A(n7605), .B(n9680), .Z(n7606) );
  NAND U7826 ( .A(n7607), .B(n7606), .Z(n7690) );
  XNOR U7827 ( .A(n9872), .B(n8220), .Z(n7708) );
  NANDN U7828 ( .A(n7708), .B(n9746), .Z(n7610) );
  NANDN U7829 ( .A(n7608), .B(n9747), .Z(n7609) );
  NAND U7830 ( .A(n7610), .B(n7609), .Z(n7687) );
  IV U7831 ( .A(a[103]), .Z(n8559) );
  XNOR U7832 ( .A(n74), .B(n8559), .Z(n7711) );
  NANDN U7833 ( .A(n7711), .B(n9485), .Z(n7613) );
  NANDN U7834 ( .A(n7611), .B(n9484), .Z(n7612) );
  AND U7835 ( .A(n7613), .B(n7612), .Z(n7688) );
  XNOR U7836 ( .A(n7687), .B(n7688), .Z(n7689) );
  XOR U7837 ( .A(n7690), .B(n7689), .Z(n7715) );
  XOR U7838 ( .A(n7714), .B(n7715), .Z(n7716) );
  XNOR U7839 ( .A(n7717), .B(n7716), .Z(n7665) );
  NAND U7840 ( .A(n7615), .B(n7614), .Z(n7619) );
  NAND U7841 ( .A(n7617), .B(n7616), .Z(n7618) );
  NAND U7842 ( .A(n7619), .B(n7618), .Z(n7666) );
  XOR U7843 ( .A(n7665), .B(n7666), .Z(n7668) );
  XNOR U7844 ( .A(n9967), .B(n7908), .Z(n7671) );
  OR U7845 ( .A(n7671), .B(n10020), .Z(n7622) );
  NANDN U7846 ( .A(n7620), .B(n9968), .Z(n7621) );
  NAND U7847 ( .A(n7622), .B(n7621), .Z(n7684) );
  XNOR U7848 ( .A(n75), .B(n7623), .Z(n7675) );
  OR U7849 ( .A(n7675), .B(n10106), .Z(n7626) );
  NANDN U7850 ( .A(n7624), .B(n10107), .Z(n7625) );
  NAND U7851 ( .A(n7626), .B(n7625), .Z(n7681) );
  XNOR U7852 ( .A(n9984), .B(n8064), .Z(n7678) );
  NANDN U7853 ( .A(n7678), .B(n9865), .Z(n7629) );
  NANDN U7854 ( .A(n7627), .B(n9930), .Z(n7628) );
  AND U7855 ( .A(n7629), .B(n7628), .Z(n7682) );
  XNOR U7856 ( .A(n7681), .B(n7682), .Z(n7683) );
  XNOR U7857 ( .A(n7684), .B(n7683), .Z(n7720) );
  NANDN U7858 ( .A(n7631), .B(n7630), .Z(n7635) );
  NAND U7859 ( .A(n7633), .B(n7632), .Z(n7634) );
  NAND U7860 ( .A(n7635), .B(n7634), .Z(n7721) );
  XNOR U7861 ( .A(n7720), .B(n7721), .Z(n7722) );
  NANDN U7862 ( .A(n7637), .B(n7636), .Z(n7641) );
  NAND U7863 ( .A(n7639), .B(n7638), .Z(n7640) );
  AND U7864 ( .A(n7641), .B(n7640), .Z(n7723) );
  XNOR U7865 ( .A(n7722), .B(n7723), .Z(n7667) );
  XNOR U7866 ( .A(n7668), .B(n7667), .Z(n7726) );
  NANDN U7867 ( .A(n7643), .B(n7642), .Z(n7647) );
  NAND U7868 ( .A(n7645), .B(n7644), .Z(n7646) );
  NAND U7869 ( .A(n7647), .B(n7646), .Z(n7727) );
  XNOR U7870 ( .A(n7726), .B(n7727), .Z(n7728) );
  XOR U7871 ( .A(n7729), .B(n7728), .Z(n7659) );
  NANDN U7872 ( .A(n7649), .B(n7648), .Z(n7653) );
  NANDN U7873 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U7874 ( .A(n7653), .B(n7652), .Z(n7660) );
  XNOR U7875 ( .A(n7659), .B(n7660), .Z(n7661) );
  XNOR U7876 ( .A(n7662), .B(n7661), .Z(n7732) );
  XNOR U7877 ( .A(n7732), .B(sreg[217]), .Z(n7734) );
  NAND U7878 ( .A(n7654), .B(sreg[216]), .Z(n7658) );
  OR U7879 ( .A(n7656), .B(n7655), .Z(n7657) );
  AND U7880 ( .A(n7658), .B(n7657), .Z(n7733) );
  XOR U7881 ( .A(n7734), .B(n7733), .Z(c[217]) );
  NANDN U7882 ( .A(n7660), .B(n7659), .Z(n7664) );
  NAND U7883 ( .A(n7662), .B(n7661), .Z(n7663) );
  NAND U7884 ( .A(n7664), .B(n7663), .Z(n7740) );
  NANDN U7885 ( .A(n7666), .B(n7665), .Z(n7670) );
  OR U7886 ( .A(n7668), .B(n7667), .Z(n7669) );
  NAND U7887 ( .A(n7670), .B(n7669), .Z(n7807) );
  XNOR U7888 ( .A(n9967), .B(n7986), .Z(n7749) );
  OR U7889 ( .A(n7749), .B(n10020), .Z(n7673) );
  NANDN U7890 ( .A(n7671), .B(n9968), .Z(n7672) );
  NAND U7891 ( .A(n7673), .B(n7672), .Z(n7762) );
  XNOR U7892 ( .A(n75), .B(n7674), .Z(n7753) );
  OR U7893 ( .A(n7753), .B(n10106), .Z(n7677) );
  NANDN U7894 ( .A(n7675), .B(n10107), .Z(n7676) );
  NAND U7895 ( .A(n7677), .B(n7676), .Z(n7759) );
  XNOR U7896 ( .A(n9984), .B(n8169), .Z(n7756) );
  NANDN U7897 ( .A(n7756), .B(n9865), .Z(n7680) );
  NANDN U7898 ( .A(n7678), .B(n9930), .Z(n7679) );
  AND U7899 ( .A(n7680), .B(n7679), .Z(n7760) );
  XNOR U7900 ( .A(n7759), .B(n7760), .Z(n7761) );
  XNOR U7901 ( .A(n7762), .B(n7761), .Z(n7798) );
  NANDN U7902 ( .A(n7682), .B(n7681), .Z(n7686) );
  NAND U7903 ( .A(n7684), .B(n7683), .Z(n7685) );
  NAND U7904 ( .A(n7686), .B(n7685), .Z(n7799) );
  XNOR U7905 ( .A(n7798), .B(n7799), .Z(n7800) );
  NANDN U7906 ( .A(n7688), .B(n7687), .Z(n7692) );
  NAND U7907 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U7908 ( .A(n7692), .B(n7691), .Z(n7801) );
  XNOR U7909 ( .A(n7800), .B(n7801), .Z(n7745) );
  NANDN U7910 ( .A(n7694), .B(n7693), .Z(n7698) );
  OR U7911 ( .A(n7696), .B(n7695), .Z(n7697) );
  NAND U7912 ( .A(n7698), .B(n7697), .Z(n7795) );
  NAND U7913 ( .A(b[0]), .B(a[106]), .Z(n7699) );
  XNOR U7914 ( .A(b[1]), .B(n7699), .Z(n7701) );
  NAND U7915 ( .A(a[105]), .B(n72), .Z(n7700) );
  AND U7916 ( .A(n7701), .B(n7700), .Z(n7771) );
  XNOR U7917 ( .A(n10050), .B(n7830), .Z(n7780) );
  OR U7918 ( .A(n7780), .B(n10051), .Z(n7704) );
  NANDN U7919 ( .A(n7702), .B(n10070), .Z(n7703) );
  AND U7920 ( .A(n7704), .B(n7703), .Z(n7772) );
  XOR U7921 ( .A(n7771), .B(n7772), .Z(n7774) );
  NAND U7922 ( .A(a[90]), .B(b[15]), .Z(n7773) );
  XOR U7923 ( .A(n7774), .B(n7773), .Z(n7792) );
  XNOR U7924 ( .A(n9622), .B(n8481), .Z(n7783) );
  OR U7925 ( .A(n7783), .B(n9623), .Z(n7707) );
  NANDN U7926 ( .A(n7705), .B(n9680), .Z(n7706) );
  NAND U7927 ( .A(n7707), .B(n7706), .Z(n7768) );
  XNOR U7928 ( .A(n9872), .B(n8298), .Z(n7786) );
  NANDN U7929 ( .A(n7786), .B(n9746), .Z(n7710) );
  NANDN U7930 ( .A(n7708), .B(n9747), .Z(n7709) );
  NAND U7931 ( .A(n7710), .B(n7709), .Z(n7765) );
  IV U7932 ( .A(a[104]), .Z(n8610) );
  XNOR U7933 ( .A(n74), .B(n8610), .Z(n7789) );
  NANDN U7934 ( .A(n7789), .B(n9485), .Z(n7713) );
  NANDN U7935 ( .A(n7711), .B(n9484), .Z(n7712) );
  AND U7936 ( .A(n7713), .B(n7712), .Z(n7766) );
  XNOR U7937 ( .A(n7765), .B(n7766), .Z(n7767) );
  XOR U7938 ( .A(n7768), .B(n7767), .Z(n7793) );
  XOR U7939 ( .A(n7792), .B(n7793), .Z(n7794) );
  XNOR U7940 ( .A(n7795), .B(n7794), .Z(n7743) );
  NAND U7941 ( .A(n7715), .B(n7714), .Z(n7719) );
  NAND U7942 ( .A(n7717), .B(n7716), .Z(n7718) );
  NAND U7943 ( .A(n7719), .B(n7718), .Z(n7744) );
  XOR U7944 ( .A(n7743), .B(n7744), .Z(n7746) );
  XNOR U7945 ( .A(n7745), .B(n7746), .Z(n7804) );
  NANDN U7946 ( .A(n7721), .B(n7720), .Z(n7725) );
  NAND U7947 ( .A(n7723), .B(n7722), .Z(n7724) );
  NAND U7948 ( .A(n7725), .B(n7724), .Z(n7805) );
  XNOR U7949 ( .A(n7804), .B(n7805), .Z(n7806) );
  XOR U7950 ( .A(n7807), .B(n7806), .Z(n7737) );
  NANDN U7951 ( .A(n7727), .B(n7726), .Z(n7731) );
  NANDN U7952 ( .A(n7729), .B(n7728), .Z(n7730) );
  NAND U7953 ( .A(n7731), .B(n7730), .Z(n7738) );
  XNOR U7954 ( .A(n7737), .B(n7738), .Z(n7739) );
  XNOR U7955 ( .A(n7740), .B(n7739), .Z(n7810) );
  XNOR U7956 ( .A(n7810), .B(sreg[218]), .Z(n7812) );
  NAND U7957 ( .A(n7732), .B(sreg[217]), .Z(n7736) );
  OR U7958 ( .A(n7734), .B(n7733), .Z(n7735) );
  AND U7959 ( .A(n7736), .B(n7735), .Z(n7811) );
  XOR U7960 ( .A(n7812), .B(n7811), .Z(c[218]) );
  NANDN U7961 ( .A(n7738), .B(n7737), .Z(n7742) );
  NAND U7962 ( .A(n7740), .B(n7739), .Z(n7741) );
  NAND U7963 ( .A(n7742), .B(n7741), .Z(n7818) );
  NANDN U7964 ( .A(n7744), .B(n7743), .Z(n7748) );
  OR U7965 ( .A(n7746), .B(n7745), .Z(n7747) );
  NAND U7966 ( .A(n7748), .B(n7747), .Z(n7885) );
  XNOR U7967 ( .A(n9967), .B(n8064), .Z(n7827) );
  OR U7968 ( .A(n7827), .B(n10020), .Z(n7751) );
  NANDN U7969 ( .A(n7749), .B(n9968), .Z(n7750) );
  NAND U7970 ( .A(n7751), .B(n7750), .Z(n7840) );
  XNOR U7971 ( .A(n75), .B(n7752), .Z(n7831) );
  OR U7972 ( .A(n7831), .B(n10106), .Z(n7755) );
  NANDN U7973 ( .A(n7753), .B(n10107), .Z(n7754) );
  NAND U7974 ( .A(n7755), .B(n7754), .Z(n7837) );
  XNOR U7975 ( .A(n9984), .B(n8220), .Z(n7834) );
  NANDN U7976 ( .A(n7834), .B(n9865), .Z(n7758) );
  NANDN U7977 ( .A(n7756), .B(n9930), .Z(n7757) );
  AND U7978 ( .A(n7758), .B(n7757), .Z(n7838) );
  XNOR U7979 ( .A(n7837), .B(n7838), .Z(n7839) );
  XNOR U7980 ( .A(n7840), .B(n7839), .Z(n7876) );
  NANDN U7981 ( .A(n7760), .B(n7759), .Z(n7764) );
  NAND U7982 ( .A(n7762), .B(n7761), .Z(n7763) );
  NAND U7983 ( .A(n7764), .B(n7763), .Z(n7877) );
  XNOR U7984 ( .A(n7876), .B(n7877), .Z(n7878) );
  NANDN U7985 ( .A(n7766), .B(n7765), .Z(n7770) );
  NAND U7986 ( .A(n7768), .B(n7767), .Z(n7769) );
  AND U7987 ( .A(n7770), .B(n7769), .Z(n7879) );
  XNOR U7988 ( .A(n7878), .B(n7879), .Z(n7823) );
  NANDN U7989 ( .A(n7772), .B(n7771), .Z(n7776) );
  OR U7990 ( .A(n7774), .B(n7773), .Z(n7775) );
  NAND U7991 ( .A(n7776), .B(n7775), .Z(n7873) );
  NAND U7992 ( .A(b[0]), .B(a[107]), .Z(n7777) );
  XNOR U7993 ( .A(b[1]), .B(n7777), .Z(n7779) );
  NAND U7994 ( .A(a[106]), .B(n72), .Z(n7778) );
  AND U7995 ( .A(n7779), .B(n7778), .Z(n7849) );
  XNOR U7996 ( .A(n10050), .B(n7908), .Z(n7855) );
  OR U7997 ( .A(n7855), .B(n10051), .Z(n7782) );
  NANDN U7998 ( .A(n7780), .B(n10070), .Z(n7781) );
  AND U7999 ( .A(n7782), .B(n7781), .Z(n7850) );
  XOR U8000 ( .A(n7849), .B(n7850), .Z(n7852) );
  NAND U8001 ( .A(a[91]), .B(b[15]), .Z(n7851) );
  XOR U8002 ( .A(n7852), .B(n7851), .Z(n7870) );
  XNOR U8003 ( .A(n9622), .B(n8559), .Z(n7861) );
  OR U8004 ( .A(n7861), .B(n9623), .Z(n7785) );
  NANDN U8005 ( .A(n7783), .B(n9680), .Z(n7784) );
  NAND U8006 ( .A(n7785), .B(n7784), .Z(n7846) );
  XNOR U8007 ( .A(n9872), .B(n8376), .Z(n7864) );
  NANDN U8008 ( .A(n7864), .B(n9746), .Z(n7788) );
  NANDN U8009 ( .A(n7786), .B(n9747), .Z(n7787) );
  NAND U8010 ( .A(n7788), .B(n7787), .Z(n7843) );
  IV U8011 ( .A(a[105]), .Z(n8688) );
  XNOR U8012 ( .A(n74), .B(n8688), .Z(n7867) );
  NANDN U8013 ( .A(n7867), .B(n9485), .Z(n7791) );
  NANDN U8014 ( .A(n7789), .B(n9484), .Z(n7790) );
  AND U8015 ( .A(n7791), .B(n7790), .Z(n7844) );
  XNOR U8016 ( .A(n7843), .B(n7844), .Z(n7845) );
  XOR U8017 ( .A(n7846), .B(n7845), .Z(n7871) );
  XOR U8018 ( .A(n7870), .B(n7871), .Z(n7872) );
  XNOR U8019 ( .A(n7873), .B(n7872), .Z(n7821) );
  NAND U8020 ( .A(n7793), .B(n7792), .Z(n7797) );
  NAND U8021 ( .A(n7795), .B(n7794), .Z(n7796) );
  NAND U8022 ( .A(n7797), .B(n7796), .Z(n7822) );
  XOR U8023 ( .A(n7821), .B(n7822), .Z(n7824) );
  XNOR U8024 ( .A(n7823), .B(n7824), .Z(n7882) );
  NANDN U8025 ( .A(n7799), .B(n7798), .Z(n7803) );
  NAND U8026 ( .A(n7801), .B(n7800), .Z(n7802) );
  NAND U8027 ( .A(n7803), .B(n7802), .Z(n7883) );
  XNOR U8028 ( .A(n7882), .B(n7883), .Z(n7884) );
  XOR U8029 ( .A(n7885), .B(n7884), .Z(n7815) );
  NANDN U8030 ( .A(n7805), .B(n7804), .Z(n7809) );
  NANDN U8031 ( .A(n7807), .B(n7806), .Z(n7808) );
  NAND U8032 ( .A(n7809), .B(n7808), .Z(n7816) );
  XNOR U8033 ( .A(n7815), .B(n7816), .Z(n7817) );
  XNOR U8034 ( .A(n7818), .B(n7817), .Z(n7888) );
  XNOR U8035 ( .A(n7888), .B(sreg[219]), .Z(n7890) );
  NAND U8036 ( .A(n7810), .B(sreg[218]), .Z(n7814) );
  OR U8037 ( .A(n7812), .B(n7811), .Z(n7813) );
  AND U8038 ( .A(n7814), .B(n7813), .Z(n7889) );
  XOR U8039 ( .A(n7890), .B(n7889), .Z(c[219]) );
  NANDN U8040 ( .A(n7816), .B(n7815), .Z(n7820) );
  NAND U8041 ( .A(n7818), .B(n7817), .Z(n7819) );
  NAND U8042 ( .A(n7820), .B(n7819), .Z(n7896) );
  NANDN U8043 ( .A(n7822), .B(n7821), .Z(n7826) );
  OR U8044 ( .A(n7824), .B(n7823), .Z(n7825) );
  NAND U8045 ( .A(n7826), .B(n7825), .Z(n7963) );
  XNOR U8046 ( .A(n9967), .B(n8169), .Z(n7905) );
  OR U8047 ( .A(n7905), .B(n10020), .Z(n7829) );
  NANDN U8048 ( .A(n7827), .B(n9968), .Z(n7828) );
  NAND U8049 ( .A(n7829), .B(n7828), .Z(n7918) );
  XNOR U8050 ( .A(n75), .B(n7830), .Z(n7909) );
  OR U8051 ( .A(n7909), .B(n10106), .Z(n7833) );
  NANDN U8052 ( .A(n7831), .B(n10107), .Z(n7832) );
  NAND U8053 ( .A(n7833), .B(n7832), .Z(n7915) );
  XNOR U8054 ( .A(n9984), .B(n8298), .Z(n7912) );
  NANDN U8055 ( .A(n7912), .B(n9865), .Z(n7836) );
  NANDN U8056 ( .A(n7834), .B(n9930), .Z(n7835) );
  AND U8057 ( .A(n7836), .B(n7835), .Z(n7916) );
  XNOR U8058 ( .A(n7915), .B(n7916), .Z(n7917) );
  XNOR U8059 ( .A(n7918), .B(n7917), .Z(n7954) );
  NANDN U8060 ( .A(n7838), .B(n7837), .Z(n7842) );
  NAND U8061 ( .A(n7840), .B(n7839), .Z(n7841) );
  NAND U8062 ( .A(n7842), .B(n7841), .Z(n7955) );
  XNOR U8063 ( .A(n7954), .B(n7955), .Z(n7956) );
  NANDN U8064 ( .A(n7844), .B(n7843), .Z(n7848) );
  NAND U8065 ( .A(n7846), .B(n7845), .Z(n7847) );
  AND U8066 ( .A(n7848), .B(n7847), .Z(n7957) );
  XNOR U8067 ( .A(n7956), .B(n7957), .Z(n7901) );
  NANDN U8068 ( .A(n7850), .B(n7849), .Z(n7854) );
  OR U8069 ( .A(n7852), .B(n7851), .Z(n7853) );
  NAND U8070 ( .A(n7854), .B(n7853), .Z(n7951) );
  XNOR U8071 ( .A(n10050), .B(n7986), .Z(n7936) );
  OR U8072 ( .A(n7936), .B(n10051), .Z(n7857) );
  NANDN U8073 ( .A(n7855), .B(n10070), .Z(n7856) );
  AND U8074 ( .A(n7857), .B(n7856), .Z(n7928) );
  NAND U8075 ( .A(b[0]), .B(a[108]), .Z(n7858) );
  XNOR U8076 ( .A(b[1]), .B(n7858), .Z(n7860) );
  NAND U8077 ( .A(a[107]), .B(n72), .Z(n7859) );
  AND U8078 ( .A(n7860), .B(n7859), .Z(n7927) );
  XOR U8079 ( .A(n7928), .B(n7927), .Z(n7930) );
  NAND U8080 ( .A(a[92]), .B(b[15]), .Z(n7929) );
  XOR U8081 ( .A(n7930), .B(n7929), .Z(n7948) );
  XNOR U8082 ( .A(n9622), .B(n8610), .Z(n7939) );
  OR U8083 ( .A(n7939), .B(n9623), .Z(n7863) );
  NANDN U8084 ( .A(n7861), .B(n9680), .Z(n7862) );
  NAND U8085 ( .A(n7863), .B(n7862), .Z(n7924) );
  XNOR U8086 ( .A(n9872), .B(n8481), .Z(n7942) );
  NANDN U8087 ( .A(n7942), .B(n9746), .Z(n7866) );
  NANDN U8088 ( .A(n7864), .B(n9747), .Z(n7865) );
  NAND U8089 ( .A(n7866), .B(n7865), .Z(n7921) );
  IV U8090 ( .A(a[106]), .Z(n8793) );
  XNOR U8091 ( .A(n74), .B(n8793), .Z(n7945) );
  NANDN U8092 ( .A(n7945), .B(n9485), .Z(n7869) );
  NANDN U8093 ( .A(n7867), .B(n9484), .Z(n7868) );
  AND U8094 ( .A(n7869), .B(n7868), .Z(n7922) );
  XNOR U8095 ( .A(n7921), .B(n7922), .Z(n7923) );
  XOR U8096 ( .A(n7924), .B(n7923), .Z(n7949) );
  XOR U8097 ( .A(n7948), .B(n7949), .Z(n7950) );
  XNOR U8098 ( .A(n7951), .B(n7950), .Z(n7899) );
  NAND U8099 ( .A(n7871), .B(n7870), .Z(n7875) );
  NAND U8100 ( .A(n7873), .B(n7872), .Z(n7874) );
  NAND U8101 ( .A(n7875), .B(n7874), .Z(n7900) );
  XOR U8102 ( .A(n7899), .B(n7900), .Z(n7902) );
  XNOR U8103 ( .A(n7901), .B(n7902), .Z(n7960) );
  NANDN U8104 ( .A(n7877), .B(n7876), .Z(n7881) );
  NAND U8105 ( .A(n7879), .B(n7878), .Z(n7880) );
  NAND U8106 ( .A(n7881), .B(n7880), .Z(n7961) );
  XNOR U8107 ( .A(n7960), .B(n7961), .Z(n7962) );
  XOR U8108 ( .A(n7963), .B(n7962), .Z(n7893) );
  NANDN U8109 ( .A(n7883), .B(n7882), .Z(n7887) );
  NANDN U8110 ( .A(n7885), .B(n7884), .Z(n7886) );
  NAND U8111 ( .A(n7887), .B(n7886), .Z(n7894) );
  XNOR U8112 ( .A(n7893), .B(n7894), .Z(n7895) );
  XNOR U8113 ( .A(n7896), .B(n7895), .Z(n7966) );
  XNOR U8114 ( .A(n7966), .B(sreg[220]), .Z(n7968) );
  NAND U8115 ( .A(n7888), .B(sreg[219]), .Z(n7892) );
  OR U8116 ( .A(n7890), .B(n7889), .Z(n7891) );
  AND U8117 ( .A(n7892), .B(n7891), .Z(n7967) );
  XOR U8118 ( .A(n7968), .B(n7967), .Z(c[220]) );
  NANDN U8119 ( .A(n7894), .B(n7893), .Z(n7898) );
  NAND U8120 ( .A(n7896), .B(n7895), .Z(n7897) );
  NAND U8121 ( .A(n7898), .B(n7897), .Z(n7974) );
  NANDN U8122 ( .A(n7900), .B(n7899), .Z(n7904) );
  OR U8123 ( .A(n7902), .B(n7901), .Z(n7903) );
  NAND U8124 ( .A(n7904), .B(n7903), .Z(n8041) );
  XNOR U8125 ( .A(n9967), .B(n8220), .Z(n7983) );
  OR U8126 ( .A(n7983), .B(n10020), .Z(n7907) );
  NANDN U8127 ( .A(n7905), .B(n9968), .Z(n7906) );
  NAND U8128 ( .A(n7907), .B(n7906), .Z(n7996) );
  XNOR U8129 ( .A(n75), .B(n7908), .Z(n7987) );
  OR U8130 ( .A(n7987), .B(n10106), .Z(n7911) );
  NANDN U8131 ( .A(n7909), .B(n10107), .Z(n7910) );
  NAND U8132 ( .A(n7911), .B(n7910), .Z(n7993) );
  XNOR U8133 ( .A(n9984), .B(n8376), .Z(n7990) );
  NANDN U8134 ( .A(n7990), .B(n9865), .Z(n7914) );
  NANDN U8135 ( .A(n7912), .B(n9930), .Z(n7913) );
  AND U8136 ( .A(n7914), .B(n7913), .Z(n7994) );
  XNOR U8137 ( .A(n7993), .B(n7994), .Z(n7995) );
  XNOR U8138 ( .A(n7996), .B(n7995), .Z(n8032) );
  NANDN U8139 ( .A(n7916), .B(n7915), .Z(n7920) );
  NAND U8140 ( .A(n7918), .B(n7917), .Z(n7919) );
  NAND U8141 ( .A(n7920), .B(n7919), .Z(n8033) );
  XNOR U8142 ( .A(n8032), .B(n8033), .Z(n8034) );
  NANDN U8143 ( .A(n7922), .B(n7921), .Z(n7926) );
  NAND U8144 ( .A(n7924), .B(n7923), .Z(n7925) );
  AND U8145 ( .A(n7926), .B(n7925), .Z(n8035) );
  XNOR U8146 ( .A(n8034), .B(n8035), .Z(n7979) );
  NANDN U8147 ( .A(n7928), .B(n7927), .Z(n7932) );
  OR U8148 ( .A(n7930), .B(n7929), .Z(n7931) );
  NAND U8149 ( .A(n7932), .B(n7931), .Z(n8029) );
  NAND U8150 ( .A(b[0]), .B(a[109]), .Z(n7933) );
  XNOR U8151 ( .A(b[1]), .B(n7933), .Z(n7935) );
  NAND U8152 ( .A(a[108]), .B(n72), .Z(n7934) );
  AND U8153 ( .A(n7935), .B(n7934), .Z(n8005) );
  XNOR U8154 ( .A(n10050), .B(n8064), .Z(n8011) );
  OR U8155 ( .A(n8011), .B(n10051), .Z(n7938) );
  NANDN U8156 ( .A(n7936), .B(n10070), .Z(n7937) );
  AND U8157 ( .A(n7938), .B(n7937), .Z(n8006) );
  XOR U8158 ( .A(n8005), .B(n8006), .Z(n8008) );
  NAND U8159 ( .A(a[93]), .B(b[15]), .Z(n8007) );
  XOR U8160 ( .A(n8008), .B(n8007), .Z(n8026) );
  XNOR U8161 ( .A(n9622), .B(n8688), .Z(n8017) );
  OR U8162 ( .A(n8017), .B(n9623), .Z(n7941) );
  NANDN U8163 ( .A(n7939), .B(n9680), .Z(n7940) );
  NAND U8164 ( .A(n7941), .B(n7940), .Z(n8002) );
  XNOR U8165 ( .A(n9872), .B(n8559), .Z(n8020) );
  NANDN U8166 ( .A(n8020), .B(n9746), .Z(n7944) );
  NANDN U8167 ( .A(n7942), .B(n9747), .Z(n7943) );
  NAND U8168 ( .A(n7944), .B(n7943), .Z(n7999) );
  IV U8169 ( .A(a[107]), .Z(n8844) );
  XNOR U8170 ( .A(n74), .B(n8844), .Z(n8023) );
  NANDN U8171 ( .A(n8023), .B(n9485), .Z(n7947) );
  NANDN U8172 ( .A(n7945), .B(n9484), .Z(n7946) );
  AND U8173 ( .A(n7947), .B(n7946), .Z(n8000) );
  XNOR U8174 ( .A(n7999), .B(n8000), .Z(n8001) );
  XOR U8175 ( .A(n8002), .B(n8001), .Z(n8027) );
  XOR U8176 ( .A(n8026), .B(n8027), .Z(n8028) );
  XNOR U8177 ( .A(n8029), .B(n8028), .Z(n7977) );
  NAND U8178 ( .A(n7949), .B(n7948), .Z(n7953) );
  NAND U8179 ( .A(n7951), .B(n7950), .Z(n7952) );
  NAND U8180 ( .A(n7953), .B(n7952), .Z(n7978) );
  XOR U8181 ( .A(n7977), .B(n7978), .Z(n7980) );
  XNOR U8182 ( .A(n7979), .B(n7980), .Z(n8038) );
  NANDN U8183 ( .A(n7955), .B(n7954), .Z(n7959) );
  NAND U8184 ( .A(n7957), .B(n7956), .Z(n7958) );
  NAND U8185 ( .A(n7959), .B(n7958), .Z(n8039) );
  XNOR U8186 ( .A(n8038), .B(n8039), .Z(n8040) );
  XOR U8187 ( .A(n8041), .B(n8040), .Z(n7971) );
  NANDN U8188 ( .A(n7961), .B(n7960), .Z(n7965) );
  NANDN U8189 ( .A(n7963), .B(n7962), .Z(n7964) );
  NAND U8190 ( .A(n7965), .B(n7964), .Z(n7972) );
  XNOR U8191 ( .A(n7971), .B(n7972), .Z(n7973) );
  XNOR U8192 ( .A(n7974), .B(n7973), .Z(n8044) );
  XNOR U8193 ( .A(n8044), .B(sreg[221]), .Z(n8046) );
  NAND U8194 ( .A(n7966), .B(sreg[220]), .Z(n7970) );
  OR U8195 ( .A(n7968), .B(n7967), .Z(n7969) );
  AND U8196 ( .A(n7970), .B(n7969), .Z(n8045) );
  XOR U8197 ( .A(n8046), .B(n8045), .Z(c[221]) );
  NANDN U8198 ( .A(n7972), .B(n7971), .Z(n7976) );
  NAND U8199 ( .A(n7974), .B(n7973), .Z(n7975) );
  NAND U8200 ( .A(n7976), .B(n7975), .Z(n8052) );
  NANDN U8201 ( .A(n7978), .B(n7977), .Z(n7982) );
  OR U8202 ( .A(n7980), .B(n7979), .Z(n7981) );
  NAND U8203 ( .A(n7982), .B(n7981), .Z(n8119) );
  XNOR U8204 ( .A(n9967), .B(n8298), .Z(n8061) );
  OR U8205 ( .A(n8061), .B(n10020), .Z(n7985) );
  NANDN U8206 ( .A(n7983), .B(n9968), .Z(n7984) );
  NAND U8207 ( .A(n7985), .B(n7984), .Z(n8074) );
  XNOR U8208 ( .A(n75), .B(n7986), .Z(n8065) );
  OR U8209 ( .A(n8065), .B(n10106), .Z(n7989) );
  NANDN U8210 ( .A(n7987), .B(n10107), .Z(n7988) );
  NAND U8211 ( .A(n7989), .B(n7988), .Z(n8071) );
  XNOR U8212 ( .A(n9984), .B(n8481), .Z(n8068) );
  NANDN U8213 ( .A(n8068), .B(n9865), .Z(n7992) );
  NANDN U8214 ( .A(n7990), .B(n9930), .Z(n7991) );
  AND U8215 ( .A(n7992), .B(n7991), .Z(n8072) );
  XNOR U8216 ( .A(n8071), .B(n8072), .Z(n8073) );
  XNOR U8217 ( .A(n8074), .B(n8073), .Z(n8110) );
  NANDN U8218 ( .A(n7994), .B(n7993), .Z(n7998) );
  NAND U8219 ( .A(n7996), .B(n7995), .Z(n7997) );
  NAND U8220 ( .A(n7998), .B(n7997), .Z(n8111) );
  XNOR U8221 ( .A(n8110), .B(n8111), .Z(n8112) );
  NANDN U8222 ( .A(n8000), .B(n7999), .Z(n8004) );
  NAND U8223 ( .A(n8002), .B(n8001), .Z(n8003) );
  AND U8224 ( .A(n8004), .B(n8003), .Z(n8113) );
  XNOR U8225 ( .A(n8112), .B(n8113), .Z(n8057) );
  NANDN U8226 ( .A(n8006), .B(n8005), .Z(n8010) );
  OR U8227 ( .A(n8008), .B(n8007), .Z(n8009) );
  NAND U8228 ( .A(n8010), .B(n8009), .Z(n8107) );
  XNOR U8229 ( .A(n10050), .B(n8169), .Z(n8089) );
  OR U8230 ( .A(n8089), .B(n10051), .Z(n8013) );
  NANDN U8231 ( .A(n8011), .B(n10070), .Z(n8012) );
  AND U8232 ( .A(n8013), .B(n8012), .Z(n8084) );
  NAND U8233 ( .A(b[0]), .B(a[110]), .Z(n8014) );
  XNOR U8234 ( .A(b[1]), .B(n8014), .Z(n8016) );
  NAND U8235 ( .A(n72), .B(a[109]), .Z(n8015) );
  AND U8236 ( .A(n8016), .B(n8015), .Z(n8083) );
  XOR U8237 ( .A(n8084), .B(n8083), .Z(n8086) );
  NAND U8238 ( .A(a[94]), .B(b[15]), .Z(n8085) );
  XOR U8239 ( .A(n8086), .B(n8085), .Z(n8104) );
  XNOR U8240 ( .A(n9622), .B(n8793), .Z(n8095) );
  OR U8241 ( .A(n8095), .B(n9623), .Z(n8019) );
  NANDN U8242 ( .A(n8017), .B(n9680), .Z(n8018) );
  NAND U8243 ( .A(n8019), .B(n8018), .Z(n8080) );
  XNOR U8244 ( .A(n9872), .B(n8610), .Z(n8098) );
  NANDN U8245 ( .A(n8098), .B(n9746), .Z(n8022) );
  NANDN U8246 ( .A(n8020), .B(n9747), .Z(n8021) );
  NAND U8247 ( .A(n8022), .B(n8021), .Z(n8077) );
  IV U8248 ( .A(a[108]), .Z(n8922) );
  XNOR U8249 ( .A(n74), .B(n8922), .Z(n8101) );
  NANDN U8250 ( .A(n8101), .B(n9485), .Z(n8025) );
  NANDN U8251 ( .A(n8023), .B(n9484), .Z(n8024) );
  AND U8252 ( .A(n8025), .B(n8024), .Z(n8078) );
  XNOR U8253 ( .A(n8077), .B(n8078), .Z(n8079) );
  XOR U8254 ( .A(n8080), .B(n8079), .Z(n8105) );
  XOR U8255 ( .A(n8104), .B(n8105), .Z(n8106) );
  XNOR U8256 ( .A(n8107), .B(n8106), .Z(n8055) );
  NAND U8257 ( .A(n8027), .B(n8026), .Z(n8031) );
  NAND U8258 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U8259 ( .A(n8031), .B(n8030), .Z(n8056) );
  XOR U8260 ( .A(n8055), .B(n8056), .Z(n8058) );
  XNOR U8261 ( .A(n8057), .B(n8058), .Z(n8116) );
  NANDN U8262 ( .A(n8033), .B(n8032), .Z(n8037) );
  NAND U8263 ( .A(n8035), .B(n8034), .Z(n8036) );
  NAND U8264 ( .A(n8037), .B(n8036), .Z(n8117) );
  XNOR U8265 ( .A(n8116), .B(n8117), .Z(n8118) );
  XOR U8266 ( .A(n8119), .B(n8118), .Z(n8049) );
  NANDN U8267 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U8268 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U8269 ( .A(n8043), .B(n8042), .Z(n8050) );
  XNOR U8270 ( .A(n8049), .B(n8050), .Z(n8051) );
  XNOR U8271 ( .A(n8052), .B(n8051), .Z(n8122) );
  XNOR U8272 ( .A(n8122), .B(sreg[222]), .Z(n8124) );
  NAND U8273 ( .A(n8044), .B(sreg[221]), .Z(n8048) );
  OR U8274 ( .A(n8046), .B(n8045), .Z(n8047) );
  AND U8275 ( .A(n8048), .B(n8047), .Z(n8123) );
  XOR U8276 ( .A(n8124), .B(n8123), .Z(c[222]) );
  NANDN U8277 ( .A(n8050), .B(n8049), .Z(n8054) );
  NAND U8278 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U8279 ( .A(n8054), .B(n8053), .Z(n8130) );
  NANDN U8280 ( .A(n8056), .B(n8055), .Z(n8060) );
  OR U8281 ( .A(n8058), .B(n8057), .Z(n8059) );
  NAND U8282 ( .A(n8060), .B(n8059), .Z(n8197) );
  XNOR U8283 ( .A(n9967), .B(n8376), .Z(n8166) );
  OR U8284 ( .A(n8166), .B(n10020), .Z(n8063) );
  NANDN U8285 ( .A(n8061), .B(n9968), .Z(n8062) );
  NAND U8286 ( .A(n8063), .B(n8062), .Z(n8179) );
  XNOR U8287 ( .A(n75), .B(n8064), .Z(n8170) );
  OR U8288 ( .A(n8170), .B(n10106), .Z(n8067) );
  NANDN U8289 ( .A(n8065), .B(n10107), .Z(n8066) );
  NAND U8290 ( .A(n8067), .B(n8066), .Z(n8176) );
  XNOR U8291 ( .A(n9984), .B(n8559), .Z(n8173) );
  NANDN U8292 ( .A(n8173), .B(n9865), .Z(n8070) );
  NANDN U8293 ( .A(n8068), .B(n9930), .Z(n8069) );
  AND U8294 ( .A(n8070), .B(n8069), .Z(n8177) );
  XNOR U8295 ( .A(n8176), .B(n8177), .Z(n8178) );
  XNOR U8296 ( .A(n8179), .B(n8178), .Z(n8188) );
  NANDN U8297 ( .A(n8072), .B(n8071), .Z(n8076) );
  NAND U8298 ( .A(n8074), .B(n8073), .Z(n8075) );
  NAND U8299 ( .A(n8076), .B(n8075), .Z(n8189) );
  XNOR U8300 ( .A(n8188), .B(n8189), .Z(n8190) );
  NANDN U8301 ( .A(n8078), .B(n8077), .Z(n8082) );
  NAND U8302 ( .A(n8080), .B(n8079), .Z(n8081) );
  AND U8303 ( .A(n8082), .B(n8081), .Z(n8191) );
  XNOR U8304 ( .A(n8190), .B(n8191), .Z(n8135) );
  NANDN U8305 ( .A(n8084), .B(n8083), .Z(n8088) );
  OR U8306 ( .A(n8086), .B(n8085), .Z(n8087) );
  NAND U8307 ( .A(n8088), .B(n8087), .Z(n8163) );
  XNOR U8308 ( .A(n10050), .B(n8220), .Z(n8148) );
  OR U8309 ( .A(n8148), .B(n10051), .Z(n8091) );
  NANDN U8310 ( .A(n8089), .B(n10070), .Z(n8090) );
  AND U8311 ( .A(n8091), .B(n8090), .Z(n8140) );
  NAND U8312 ( .A(b[0]), .B(a[111]), .Z(n8092) );
  XNOR U8313 ( .A(b[1]), .B(n8092), .Z(n8094) );
  NAND U8314 ( .A(a[110]), .B(n72), .Z(n8093) );
  AND U8315 ( .A(n8094), .B(n8093), .Z(n8139) );
  XOR U8316 ( .A(n8140), .B(n8139), .Z(n8142) );
  NAND U8317 ( .A(a[95]), .B(b[15]), .Z(n8141) );
  XOR U8318 ( .A(n8142), .B(n8141), .Z(n8160) );
  XNOR U8319 ( .A(n9622), .B(n8844), .Z(n8151) );
  OR U8320 ( .A(n8151), .B(n9623), .Z(n8097) );
  NANDN U8321 ( .A(n8095), .B(n9680), .Z(n8096) );
  NAND U8322 ( .A(n8097), .B(n8096), .Z(n8185) );
  XNOR U8323 ( .A(n9872), .B(n8688), .Z(n8154) );
  NANDN U8324 ( .A(n8154), .B(n9746), .Z(n8100) );
  NANDN U8325 ( .A(n8098), .B(n9747), .Z(n8099) );
  NAND U8326 ( .A(n8100), .B(n8099), .Z(n8182) );
  XOR U8327 ( .A(n74), .B(a[109]), .Z(n8157) );
  NANDN U8328 ( .A(n8157), .B(n9485), .Z(n8103) );
  NANDN U8329 ( .A(n8101), .B(n9484), .Z(n8102) );
  AND U8330 ( .A(n8103), .B(n8102), .Z(n8183) );
  XNOR U8331 ( .A(n8182), .B(n8183), .Z(n8184) );
  XOR U8332 ( .A(n8185), .B(n8184), .Z(n8161) );
  XOR U8333 ( .A(n8160), .B(n8161), .Z(n8162) );
  XNOR U8334 ( .A(n8163), .B(n8162), .Z(n8133) );
  NAND U8335 ( .A(n8105), .B(n8104), .Z(n8109) );
  NAND U8336 ( .A(n8107), .B(n8106), .Z(n8108) );
  NAND U8337 ( .A(n8109), .B(n8108), .Z(n8134) );
  XOR U8338 ( .A(n8133), .B(n8134), .Z(n8136) );
  XNOR U8339 ( .A(n8135), .B(n8136), .Z(n8194) );
  NANDN U8340 ( .A(n8111), .B(n8110), .Z(n8115) );
  NAND U8341 ( .A(n8113), .B(n8112), .Z(n8114) );
  NAND U8342 ( .A(n8115), .B(n8114), .Z(n8195) );
  XNOR U8343 ( .A(n8194), .B(n8195), .Z(n8196) );
  XOR U8344 ( .A(n8197), .B(n8196), .Z(n8127) );
  NANDN U8345 ( .A(n8117), .B(n8116), .Z(n8121) );
  NANDN U8346 ( .A(n8119), .B(n8118), .Z(n8120) );
  NAND U8347 ( .A(n8121), .B(n8120), .Z(n8128) );
  XNOR U8348 ( .A(n8127), .B(n8128), .Z(n8129) );
  XNOR U8349 ( .A(n8130), .B(n8129), .Z(n8200) );
  XNOR U8350 ( .A(n8200), .B(sreg[223]), .Z(n8202) );
  NAND U8351 ( .A(n8122), .B(sreg[222]), .Z(n8126) );
  OR U8352 ( .A(n8124), .B(n8123), .Z(n8125) );
  AND U8353 ( .A(n8126), .B(n8125), .Z(n8201) );
  XOR U8354 ( .A(n8202), .B(n8201), .Z(c[223]) );
  NANDN U8355 ( .A(n8128), .B(n8127), .Z(n8132) );
  NAND U8356 ( .A(n8130), .B(n8129), .Z(n8131) );
  NAND U8357 ( .A(n8132), .B(n8131), .Z(n8208) );
  NANDN U8358 ( .A(n8134), .B(n8133), .Z(n8138) );
  OR U8359 ( .A(n8136), .B(n8135), .Z(n8137) );
  NAND U8360 ( .A(n8138), .B(n8137), .Z(n8275) );
  NANDN U8361 ( .A(n8140), .B(n8139), .Z(n8144) );
  OR U8362 ( .A(n8142), .B(n8141), .Z(n8143) );
  NAND U8363 ( .A(n8144), .B(n8143), .Z(n8263) );
  NAND U8364 ( .A(b[0]), .B(a[112]), .Z(n8145) );
  XNOR U8365 ( .A(b[1]), .B(n8145), .Z(n8147) );
  NAND U8366 ( .A(n72), .B(a[111]), .Z(n8146) );
  AND U8367 ( .A(n8147), .B(n8146), .Z(n8239) );
  XNOR U8368 ( .A(n10050), .B(n8298), .Z(n8248) );
  OR U8369 ( .A(n8248), .B(n10051), .Z(n8150) );
  NANDN U8370 ( .A(n8148), .B(n10070), .Z(n8149) );
  AND U8371 ( .A(n8150), .B(n8149), .Z(n8240) );
  XOR U8372 ( .A(n8239), .B(n8240), .Z(n8242) );
  NAND U8373 ( .A(a[96]), .B(b[15]), .Z(n8241) );
  XOR U8374 ( .A(n8242), .B(n8241), .Z(n8260) );
  XNOR U8375 ( .A(n9622), .B(n8922), .Z(n8251) );
  OR U8376 ( .A(n8251), .B(n9623), .Z(n8153) );
  NANDN U8377 ( .A(n8151), .B(n9680), .Z(n8152) );
  NAND U8378 ( .A(n8153), .B(n8152), .Z(n8236) );
  XNOR U8379 ( .A(n9872), .B(n8793), .Z(n8254) );
  NANDN U8380 ( .A(n8254), .B(n9746), .Z(n8156) );
  NANDN U8381 ( .A(n8154), .B(n9747), .Z(n8155) );
  NAND U8382 ( .A(n8156), .B(n8155), .Z(n8233) );
  IV U8383 ( .A(a[110]), .Z(n9077) );
  XNOR U8384 ( .A(n74), .B(n9077), .Z(n8257) );
  NANDN U8385 ( .A(n8257), .B(n9485), .Z(n8159) );
  NANDN U8386 ( .A(n8157), .B(n9484), .Z(n8158) );
  AND U8387 ( .A(n8159), .B(n8158), .Z(n8234) );
  XNOR U8388 ( .A(n8233), .B(n8234), .Z(n8235) );
  XOR U8389 ( .A(n8236), .B(n8235), .Z(n8261) );
  XOR U8390 ( .A(n8260), .B(n8261), .Z(n8262) );
  XNOR U8391 ( .A(n8263), .B(n8262), .Z(n8211) );
  NAND U8392 ( .A(n8161), .B(n8160), .Z(n8165) );
  NAND U8393 ( .A(n8163), .B(n8162), .Z(n8164) );
  NAND U8394 ( .A(n8165), .B(n8164), .Z(n8212) );
  XOR U8395 ( .A(n8211), .B(n8212), .Z(n8214) );
  XNOR U8396 ( .A(n9967), .B(n8481), .Z(n8217) );
  OR U8397 ( .A(n8217), .B(n10020), .Z(n8168) );
  NANDN U8398 ( .A(n8166), .B(n9968), .Z(n8167) );
  NAND U8399 ( .A(n8168), .B(n8167), .Z(n8230) );
  XNOR U8400 ( .A(n75), .B(n8169), .Z(n8221) );
  OR U8401 ( .A(n8221), .B(n10106), .Z(n8172) );
  NANDN U8402 ( .A(n8170), .B(n10107), .Z(n8171) );
  NAND U8403 ( .A(n8172), .B(n8171), .Z(n8227) );
  XNOR U8404 ( .A(n9984), .B(n8610), .Z(n8224) );
  NANDN U8405 ( .A(n8224), .B(n9865), .Z(n8175) );
  NANDN U8406 ( .A(n8173), .B(n9930), .Z(n8174) );
  AND U8407 ( .A(n8175), .B(n8174), .Z(n8228) );
  XNOR U8408 ( .A(n8227), .B(n8228), .Z(n8229) );
  XNOR U8409 ( .A(n8230), .B(n8229), .Z(n8266) );
  NANDN U8410 ( .A(n8177), .B(n8176), .Z(n8181) );
  NAND U8411 ( .A(n8179), .B(n8178), .Z(n8180) );
  NAND U8412 ( .A(n8181), .B(n8180), .Z(n8267) );
  XNOR U8413 ( .A(n8266), .B(n8267), .Z(n8268) );
  NANDN U8414 ( .A(n8183), .B(n8182), .Z(n8187) );
  NAND U8415 ( .A(n8185), .B(n8184), .Z(n8186) );
  AND U8416 ( .A(n8187), .B(n8186), .Z(n8269) );
  XNOR U8417 ( .A(n8268), .B(n8269), .Z(n8213) );
  XNOR U8418 ( .A(n8214), .B(n8213), .Z(n8272) );
  NANDN U8419 ( .A(n8189), .B(n8188), .Z(n8193) );
  NAND U8420 ( .A(n8191), .B(n8190), .Z(n8192) );
  NAND U8421 ( .A(n8193), .B(n8192), .Z(n8273) );
  XNOR U8422 ( .A(n8272), .B(n8273), .Z(n8274) );
  XOR U8423 ( .A(n8275), .B(n8274), .Z(n8205) );
  NANDN U8424 ( .A(n8195), .B(n8194), .Z(n8199) );
  NANDN U8425 ( .A(n8197), .B(n8196), .Z(n8198) );
  NAND U8426 ( .A(n8199), .B(n8198), .Z(n8206) );
  XNOR U8427 ( .A(n8205), .B(n8206), .Z(n8207) );
  XNOR U8428 ( .A(n8208), .B(n8207), .Z(n8278) );
  XNOR U8429 ( .A(n8278), .B(sreg[224]), .Z(n8280) );
  NAND U8430 ( .A(n8200), .B(sreg[223]), .Z(n8204) );
  OR U8431 ( .A(n8202), .B(n8201), .Z(n8203) );
  AND U8432 ( .A(n8204), .B(n8203), .Z(n8279) );
  XOR U8433 ( .A(n8280), .B(n8279), .Z(c[224]) );
  NANDN U8434 ( .A(n8206), .B(n8205), .Z(n8210) );
  NAND U8435 ( .A(n8208), .B(n8207), .Z(n8209) );
  NAND U8436 ( .A(n8210), .B(n8209), .Z(n8286) );
  NANDN U8437 ( .A(n8212), .B(n8211), .Z(n8216) );
  OR U8438 ( .A(n8214), .B(n8213), .Z(n8215) );
  NAND U8439 ( .A(n8216), .B(n8215), .Z(n8353) );
  XNOR U8440 ( .A(n9967), .B(n8559), .Z(n8295) );
  OR U8441 ( .A(n8295), .B(n10020), .Z(n8219) );
  NANDN U8442 ( .A(n8217), .B(n9968), .Z(n8218) );
  NAND U8443 ( .A(n8219), .B(n8218), .Z(n8308) );
  XNOR U8444 ( .A(n75), .B(n8220), .Z(n8299) );
  OR U8445 ( .A(n8299), .B(n10106), .Z(n8223) );
  NANDN U8446 ( .A(n8221), .B(n10107), .Z(n8222) );
  NAND U8447 ( .A(n8223), .B(n8222), .Z(n8305) );
  XNOR U8448 ( .A(n9984), .B(n8688), .Z(n8302) );
  NANDN U8449 ( .A(n8302), .B(n9865), .Z(n8226) );
  NANDN U8450 ( .A(n8224), .B(n9930), .Z(n8225) );
  AND U8451 ( .A(n8226), .B(n8225), .Z(n8306) );
  XNOR U8452 ( .A(n8305), .B(n8306), .Z(n8307) );
  XNOR U8453 ( .A(n8308), .B(n8307), .Z(n8344) );
  NANDN U8454 ( .A(n8228), .B(n8227), .Z(n8232) );
  NAND U8455 ( .A(n8230), .B(n8229), .Z(n8231) );
  NAND U8456 ( .A(n8232), .B(n8231), .Z(n8345) );
  XNOR U8457 ( .A(n8344), .B(n8345), .Z(n8346) );
  NANDN U8458 ( .A(n8234), .B(n8233), .Z(n8238) );
  NAND U8459 ( .A(n8236), .B(n8235), .Z(n8237) );
  AND U8460 ( .A(n8238), .B(n8237), .Z(n8347) );
  XNOR U8461 ( .A(n8346), .B(n8347), .Z(n8291) );
  NANDN U8462 ( .A(n8240), .B(n8239), .Z(n8244) );
  OR U8463 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8464 ( .A(n8244), .B(n8243), .Z(n8341) );
  NAND U8465 ( .A(b[0]), .B(a[113]), .Z(n8245) );
  XNOR U8466 ( .A(b[1]), .B(n8245), .Z(n8247) );
  NAND U8467 ( .A(n72), .B(a[112]), .Z(n8246) );
  AND U8468 ( .A(n8247), .B(n8246), .Z(n8317) );
  XNOR U8469 ( .A(n10050), .B(n8376), .Z(n8326) );
  OR U8470 ( .A(n8326), .B(n10051), .Z(n8250) );
  NANDN U8471 ( .A(n8248), .B(n10070), .Z(n8249) );
  AND U8472 ( .A(n8250), .B(n8249), .Z(n8318) );
  XOR U8473 ( .A(n8317), .B(n8318), .Z(n8320) );
  NAND U8474 ( .A(a[97]), .B(b[15]), .Z(n8319) );
  XOR U8475 ( .A(n8320), .B(n8319), .Z(n8338) );
  XOR U8476 ( .A(n9622), .B(a[109]), .Z(n8329) );
  OR U8477 ( .A(n8329), .B(n9623), .Z(n8253) );
  NANDN U8478 ( .A(n8251), .B(n9680), .Z(n8252) );
  NAND U8479 ( .A(n8253), .B(n8252), .Z(n8314) );
  XNOR U8480 ( .A(n9872), .B(n8844), .Z(n8332) );
  NANDN U8481 ( .A(n8332), .B(n9746), .Z(n8256) );
  NANDN U8482 ( .A(n8254), .B(n9747), .Z(n8255) );
  NAND U8483 ( .A(n8256), .B(n8255), .Z(n8311) );
  XOR U8484 ( .A(n74), .B(a[111]), .Z(n8335) );
  NANDN U8485 ( .A(n8335), .B(n9485), .Z(n8259) );
  NANDN U8486 ( .A(n8257), .B(n9484), .Z(n8258) );
  AND U8487 ( .A(n8259), .B(n8258), .Z(n8312) );
  XNOR U8488 ( .A(n8311), .B(n8312), .Z(n8313) );
  XOR U8489 ( .A(n8314), .B(n8313), .Z(n8339) );
  XOR U8490 ( .A(n8338), .B(n8339), .Z(n8340) );
  XNOR U8491 ( .A(n8341), .B(n8340), .Z(n8289) );
  NAND U8492 ( .A(n8261), .B(n8260), .Z(n8265) );
  NAND U8493 ( .A(n8263), .B(n8262), .Z(n8264) );
  NAND U8494 ( .A(n8265), .B(n8264), .Z(n8290) );
  XOR U8495 ( .A(n8289), .B(n8290), .Z(n8292) );
  XNOR U8496 ( .A(n8291), .B(n8292), .Z(n8350) );
  NANDN U8497 ( .A(n8267), .B(n8266), .Z(n8271) );
  NAND U8498 ( .A(n8269), .B(n8268), .Z(n8270) );
  NAND U8499 ( .A(n8271), .B(n8270), .Z(n8351) );
  XNOR U8500 ( .A(n8350), .B(n8351), .Z(n8352) );
  XOR U8501 ( .A(n8353), .B(n8352), .Z(n8283) );
  NANDN U8502 ( .A(n8273), .B(n8272), .Z(n8277) );
  NANDN U8503 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U8504 ( .A(n8277), .B(n8276), .Z(n8284) );
  XNOR U8505 ( .A(n8283), .B(n8284), .Z(n8285) );
  XNOR U8506 ( .A(n8286), .B(n8285), .Z(n8356) );
  XNOR U8507 ( .A(n8356), .B(sreg[225]), .Z(n8358) );
  NAND U8508 ( .A(n8278), .B(sreg[224]), .Z(n8282) );
  OR U8509 ( .A(n8280), .B(n8279), .Z(n8281) );
  AND U8510 ( .A(n8282), .B(n8281), .Z(n8357) );
  XOR U8511 ( .A(n8358), .B(n8357), .Z(c[225]) );
  NANDN U8512 ( .A(n8284), .B(n8283), .Z(n8288) );
  NAND U8513 ( .A(n8286), .B(n8285), .Z(n8287) );
  NAND U8514 ( .A(n8288), .B(n8287), .Z(n8364) );
  NANDN U8515 ( .A(n8290), .B(n8289), .Z(n8294) );
  OR U8516 ( .A(n8292), .B(n8291), .Z(n8293) );
  NAND U8517 ( .A(n8294), .B(n8293), .Z(n8431) );
  XNOR U8518 ( .A(n9967), .B(n8610), .Z(n8373) );
  OR U8519 ( .A(n8373), .B(n10020), .Z(n8297) );
  NANDN U8520 ( .A(n8295), .B(n9968), .Z(n8296) );
  NAND U8521 ( .A(n8297), .B(n8296), .Z(n8386) );
  XNOR U8522 ( .A(n75), .B(n8298), .Z(n8377) );
  OR U8523 ( .A(n8377), .B(n10106), .Z(n8301) );
  NANDN U8524 ( .A(n8299), .B(n10107), .Z(n8300) );
  NAND U8525 ( .A(n8301), .B(n8300), .Z(n8383) );
  XNOR U8526 ( .A(n9984), .B(n8793), .Z(n8380) );
  NANDN U8527 ( .A(n8380), .B(n9865), .Z(n8304) );
  NANDN U8528 ( .A(n8302), .B(n9930), .Z(n8303) );
  AND U8529 ( .A(n8304), .B(n8303), .Z(n8384) );
  XNOR U8530 ( .A(n8383), .B(n8384), .Z(n8385) );
  XNOR U8531 ( .A(n8386), .B(n8385), .Z(n8422) );
  NANDN U8532 ( .A(n8306), .B(n8305), .Z(n8310) );
  NAND U8533 ( .A(n8308), .B(n8307), .Z(n8309) );
  NAND U8534 ( .A(n8310), .B(n8309), .Z(n8423) );
  XNOR U8535 ( .A(n8422), .B(n8423), .Z(n8424) );
  NANDN U8536 ( .A(n8312), .B(n8311), .Z(n8316) );
  NAND U8537 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U8538 ( .A(n8316), .B(n8315), .Z(n8425) );
  XNOR U8539 ( .A(n8424), .B(n8425), .Z(n8369) );
  NANDN U8540 ( .A(n8318), .B(n8317), .Z(n8322) );
  OR U8541 ( .A(n8320), .B(n8319), .Z(n8321) );
  NAND U8542 ( .A(n8322), .B(n8321), .Z(n8419) );
  NAND U8543 ( .A(b[0]), .B(a[114]), .Z(n8323) );
  XNOR U8544 ( .A(b[1]), .B(n8323), .Z(n8325) );
  NAND U8545 ( .A(n72), .B(a[113]), .Z(n8324) );
  AND U8546 ( .A(n8325), .B(n8324), .Z(n8395) );
  XNOR U8547 ( .A(n10050), .B(n8481), .Z(n8401) );
  OR U8548 ( .A(n8401), .B(n10051), .Z(n8328) );
  NANDN U8549 ( .A(n8326), .B(n10070), .Z(n8327) );
  AND U8550 ( .A(n8328), .B(n8327), .Z(n8396) );
  XOR U8551 ( .A(n8395), .B(n8396), .Z(n8398) );
  NAND U8552 ( .A(a[98]), .B(b[15]), .Z(n8397) );
  XOR U8553 ( .A(n8398), .B(n8397), .Z(n8416) );
  XNOR U8554 ( .A(n9622), .B(n9077), .Z(n8407) );
  OR U8555 ( .A(n8407), .B(n9623), .Z(n8331) );
  NANDN U8556 ( .A(n8329), .B(n9680), .Z(n8330) );
  NAND U8557 ( .A(n8331), .B(n8330), .Z(n8392) );
  XNOR U8558 ( .A(n9872), .B(n8922), .Z(n8410) );
  NANDN U8559 ( .A(n8410), .B(n9746), .Z(n8334) );
  NANDN U8560 ( .A(n8332), .B(n9747), .Z(n8333) );
  NAND U8561 ( .A(n8334), .B(n8333), .Z(n8389) );
  XOR U8562 ( .A(n74), .B(a[112]), .Z(n8413) );
  NANDN U8563 ( .A(n8413), .B(n9485), .Z(n8337) );
  NANDN U8564 ( .A(n8335), .B(n9484), .Z(n8336) );
  AND U8565 ( .A(n8337), .B(n8336), .Z(n8390) );
  XNOR U8566 ( .A(n8389), .B(n8390), .Z(n8391) );
  XOR U8567 ( .A(n8392), .B(n8391), .Z(n8417) );
  XOR U8568 ( .A(n8416), .B(n8417), .Z(n8418) );
  XNOR U8569 ( .A(n8419), .B(n8418), .Z(n8367) );
  NAND U8570 ( .A(n8339), .B(n8338), .Z(n8343) );
  NAND U8571 ( .A(n8341), .B(n8340), .Z(n8342) );
  NAND U8572 ( .A(n8343), .B(n8342), .Z(n8368) );
  XOR U8573 ( .A(n8367), .B(n8368), .Z(n8370) );
  XNOR U8574 ( .A(n8369), .B(n8370), .Z(n8428) );
  NANDN U8575 ( .A(n8345), .B(n8344), .Z(n8349) );
  NAND U8576 ( .A(n8347), .B(n8346), .Z(n8348) );
  NAND U8577 ( .A(n8349), .B(n8348), .Z(n8429) );
  XNOR U8578 ( .A(n8428), .B(n8429), .Z(n8430) );
  XOR U8579 ( .A(n8431), .B(n8430), .Z(n8361) );
  NANDN U8580 ( .A(n8351), .B(n8350), .Z(n8355) );
  NANDN U8581 ( .A(n8353), .B(n8352), .Z(n8354) );
  NAND U8582 ( .A(n8355), .B(n8354), .Z(n8362) );
  XNOR U8583 ( .A(n8361), .B(n8362), .Z(n8363) );
  XNOR U8584 ( .A(n8364), .B(n8363), .Z(n8434) );
  XNOR U8585 ( .A(n8434), .B(sreg[226]), .Z(n8436) );
  NAND U8586 ( .A(n8356), .B(sreg[225]), .Z(n8360) );
  OR U8587 ( .A(n8358), .B(n8357), .Z(n8359) );
  AND U8588 ( .A(n8360), .B(n8359), .Z(n8435) );
  XOR U8589 ( .A(n8436), .B(n8435), .Z(c[226]) );
  NANDN U8590 ( .A(n8362), .B(n8361), .Z(n8366) );
  NAND U8591 ( .A(n8364), .B(n8363), .Z(n8365) );
  NAND U8592 ( .A(n8366), .B(n8365), .Z(n8442) );
  NANDN U8593 ( .A(n8368), .B(n8367), .Z(n8372) );
  OR U8594 ( .A(n8370), .B(n8369), .Z(n8371) );
  NAND U8595 ( .A(n8372), .B(n8371), .Z(n8509) );
  XNOR U8596 ( .A(n9967), .B(n8688), .Z(n8478) );
  OR U8597 ( .A(n8478), .B(n10020), .Z(n8375) );
  NANDN U8598 ( .A(n8373), .B(n9968), .Z(n8374) );
  NAND U8599 ( .A(n8375), .B(n8374), .Z(n8491) );
  XNOR U8600 ( .A(n75), .B(n8376), .Z(n8482) );
  OR U8601 ( .A(n8482), .B(n10106), .Z(n8379) );
  NANDN U8602 ( .A(n8377), .B(n10107), .Z(n8378) );
  NAND U8603 ( .A(n8379), .B(n8378), .Z(n8488) );
  XNOR U8604 ( .A(n9984), .B(n8844), .Z(n8485) );
  NANDN U8605 ( .A(n8485), .B(n9865), .Z(n8382) );
  NANDN U8606 ( .A(n8380), .B(n9930), .Z(n8381) );
  AND U8607 ( .A(n8382), .B(n8381), .Z(n8489) );
  XNOR U8608 ( .A(n8488), .B(n8489), .Z(n8490) );
  XNOR U8609 ( .A(n8491), .B(n8490), .Z(n8500) );
  NANDN U8610 ( .A(n8384), .B(n8383), .Z(n8388) );
  NAND U8611 ( .A(n8386), .B(n8385), .Z(n8387) );
  NAND U8612 ( .A(n8388), .B(n8387), .Z(n8501) );
  XNOR U8613 ( .A(n8500), .B(n8501), .Z(n8502) );
  NANDN U8614 ( .A(n8390), .B(n8389), .Z(n8394) );
  NAND U8615 ( .A(n8392), .B(n8391), .Z(n8393) );
  AND U8616 ( .A(n8394), .B(n8393), .Z(n8503) );
  XNOR U8617 ( .A(n8502), .B(n8503), .Z(n8447) );
  NANDN U8618 ( .A(n8396), .B(n8395), .Z(n8400) );
  OR U8619 ( .A(n8398), .B(n8397), .Z(n8399) );
  NAND U8620 ( .A(n8400), .B(n8399), .Z(n8475) );
  XNOR U8621 ( .A(n10050), .B(n8559), .Z(n8457) );
  OR U8622 ( .A(n8457), .B(n10051), .Z(n8403) );
  NANDN U8623 ( .A(n8401), .B(n10070), .Z(n8402) );
  AND U8624 ( .A(n8403), .B(n8402), .Z(n8452) );
  NAND U8625 ( .A(b[0]), .B(a[115]), .Z(n8404) );
  XNOR U8626 ( .A(b[1]), .B(n8404), .Z(n8406) );
  NAND U8627 ( .A(a[114]), .B(n72), .Z(n8405) );
  AND U8628 ( .A(n8406), .B(n8405), .Z(n8451) );
  XOR U8629 ( .A(n8452), .B(n8451), .Z(n8454) );
  NAND U8630 ( .A(a[99]), .B(b[15]), .Z(n8453) );
  XOR U8631 ( .A(n8454), .B(n8453), .Z(n8472) );
  XOR U8632 ( .A(n9622), .B(a[111]), .Z(n8463) );
  OR U8633 ( .A(n8463), .B(n9623), .Z(n8409) );
  NANDN U8634 ( .A(n8407), .B(n9680), .Z(n8408) );
  NAND U8635 ( .A(n8409), .B(n8408), .Z(n8497) );
  XOR U8636 ( .A(n9872), .B(a[109]), .Z(n8466) );
  NANDN U8637 ( .A(n8466), .B(n9746), .Z(n8412) );
  NANDN U8638 ( .A(n8410), .B(n9747), .Z(n8411) );
  NAND U8639 ( .A(n8412), .B(n8411), .Z(n8494) );
  XOR U8640 ( .A(n74), .B(a[113]), .Z(n8469) );
  NANDN U8641 ( .A(n8469), .B(n9485), .Z(n8415) );
  NANDN U8642 ( .A(n8413), .B(n9484), .Z(n8414) );
  AND U8643 ( .A(n8415), .B(n8414), .Z(n8495) );
  XNOR U8644 ( .A(n8494), .B(n8495), .Z(n8496) );
  XOR U8645 ( .A(n8497), .B(n8496), .Z(n8473) );
  XOR U8646 ( .A(n8472), .B(n8473), .Z(n8474) );
  XNOR U8647 ( .A(n8475), .B(n8474), .Z(n8445) );
  NAND U8648 ( .A(n8417), .B(n8416), .Z(n8421) );
  NAND U8649 ( .A(n8419), .B(n8418), .Z(n8420) );
  NAND U8650 ( .A(n8421), .B(n8420), .Z(n8446) );
  XOR U8651 ( .A(n8445), .B(n8446), .Z(n8448) );
  XNOR U8652 ( .A(n8447), .B(n8448), .Z(n8506) );
  NANDN U8653 ( .A(n8423), .B(n8422), .Z(n8427) );
  NAND U8654 ( .A(n8425), .B(n8424), .Z(n8426) );
  NAND U8655 ( .A(n8427), .B(n8426), .Z(n8507) );
  XNOR U8656 ( .A(n8506), .B(n8507), .Z(n8508) );
  XOR U8657 ( .A(n8509), .B(n8508), .Z(n8439) );
  NANDN U8658 ( .A(n8429), .B(n8428), .Z(n8433) );
  NANDN U8659 ( .A(n8431), .B(n8430), .Z(n8432) );
  NAND U8660 ( .A(n8433), .B(n8432), .Z(n8440) );
  XNOR U8661 ( .A(n8439), .B(n8440), .Z(n8441) );
  XNOR U8662 ( .A(n8442), .B(n8441), .Z(n8512) );
  XNOR U8663 ( .A(n8512), .B(sreg[227]), .Z(n8514) );
  NAND U8664 ( .A(n8434), .B(sreg[226]), .Z(n8438) );
  OR U8665 ( .A(n8436), .B(n8435), .Z(n8437) );
  AND U8666 ( .A(n8438), .B(n8437), .Z(n8513) );
  XOR U8667 ( .A(n8514), .B(n8513), .Z(c[227]) );
  NANDN U8668 ( .A(n8440), .B(n8439), .Z(n8444) );
  NAND U8669 ( .A(n8442), .B(n8441), .Z(n8443) );
  NAND U8670 ( .A(n8444), .B(n8443), .Z(n8520) );
  NANDN U8671 ( .A(n8446), .B(n8445), .Z(n8450) );
  OR U8672 ( .A(n8448), .B(n8447), .Z(n8449) );
  NAND U8673 ( .A(n8450), .B(n8449), .Z(n8587) );
  NANDN U8674 ( .A(n8452), .B(n8451), .Z(n8456) );
  OR U8675 ( .A(n8454), .B(n8453), .Z(n8455) );
  NAND U8676 ( .A(n8456), .B(n8455), .Z(n8553) );
  XNOR U8677 ( .A(n10050), .B(n8610), .Z(n8538) );
  OR U8678 ( .A(n8538), .B(n10051), .Z(n8459) );
  NANDN U8679 ( .A(n8457), .B(n10070), .Z(n8458) );
  AND U8680 ( .A(n8459), .B(n8458), .Z(n8530) );
  NAND U8681 ( .A(b[0]), .B(a[116]), .Z(n8460) );
  XNOR U8682 ( .A(b[1]), .B(n8460), .Z(n8462) );
  NAND U8683 ( .A(n72), .B(a[115]), .Z(n8461) );
  AND U8684 ( .A(n8462), .B(n8461), .Z(n8529) );
  XOR U8685 ( .A(n8530), .B(n8529), .Z(n8532) );
  NAND U8686 ( .A(a[100]), .B(b[15]), .Z(n8531) );
  XOR U8687 ( .A(n8532), .B(n8531), .Z(n8550) );
  XOR U8688 ( .A(n9622), .B(a[112]), .Z(n8541) );
  OR U8689 ( .A(n8541), .B(n9623), .Z(n8465) );
  NANDN U8690 ( .A(n8463), .B(n9680), .Z(n8464) );
  NAND U8691 ( .A(n8465), .B(n8464), .Z(n8575) );
  XNOR U8692 ( .A(n9872), .B(n9077), .Z(n8544) );
  NANDN U8693 ( .A(n8544), .B(n9746), .Z(n8468) );
  NANDN U8694 ( .A(n8466), .B(n9747), .Z(n8467) );
  NAND U8695 ( .A(n8468), .B(n8467), .Z(n8572) );
  IV U8696 ( .A(a[114]), .Z(n9397) );
  XNOR U8697 ( .A(n74), .B(n9397), .Z(n8547) );
  NANDN U8698 ( .A(n8547), .B(n9485), .Z(n8471) );
  NANDN U8699 ( .A(n8469), .B(n9484), .Z(n8470) );
  AND U8700 ( .A(n8471), .B(n8470), .Z(n8573) );
  XNOR U8701 ( .A(n8572), .B(n8573), .Z(n8574) );
  XOR U8702 ( .A(n8575), .B(n8574), .Z(n8551) );
  XOR U8703 ( .A(n8550), .B(n8551), .Z(n8552) );
  XNOR U8704 ( .A(n8553), .B(n8552), .Z(n8523) );
  NAND U8705 ( .A(n8473), .B(n8472), .Z(n8477) );
  NAND U8706 ( .A(n8475), .B(n8474), .Z(n8476) );
  NAND U8707 ( .A(n8477), .B(n8476), .Z(n8524) );
  XOR U8708 ( .A(n8523), .B(n8524), .Z(n8526) );
  XNOR U8709 ( .A(n9967), .B(n8793), .Z(n8556) );
  OR U8710 ( .A(n8556), .B(n10020), .Z(n8480) );
  NANDN U8711 ( .A(n8478), .B(n9968), .Z(n8479) );
  NAND U8712 ( .A(n8480), .B(n8479), .Z(n8569) );
  XNOR U8713 ( .A(n75), .B(n8481), .Z(n8560) );
  OR U8714 ( .A(n8560), .B(n10106), .Z(n8484) );
  NANDN U8715 ( .A(n8482), .B(n10107), .Z(n8483) );
  NAND U8716 ( .A(n8484), .B(n8483), .Z(n8566) );
  XNOR U8717 ( .A(n9984), .B(n8922), .Z(n8563) );
  NANDN U8718 ( .A(n8563), .B(n9865), .Z(n8487) );
  NANDN U8719 ( .A(n8485), .B(n9930), .Z(n8486) );
  AND U8720 ( .A(n8487), .B(n8486), .Z(n8567) );
  XNOR U8721 ( .A(n8566), .B(n8567), .Z(n8568) );
  XNOR U8722 ( .A(n8569), .B(n8568), .Z(n8578) );
  NANDN U8723 ( .A(n8489), .B(n8488), .Z(n8493) );
  NAND U8724 ( .A(n8491), .B(n8490), .Z(n8492) );
  NAND U8725 ( .A(n8493), .B(n8492), .Z(n8579) );
  XNOR U8726 ( .A(n8578), .B(n8579), .Z(n8580) );
  NANDN U8727 ( .A(n8495), .B(n8494), .Z(n8499) );
  NAND U8728 ( .A(n8497), .B(n8496), .Z(n8498) );
  AND U8729 ( .A(n8499), .B(n8498), .Z(n8581) );
  XNOR U8730 ( .A(n8580), .B(n8581), .Z(n8525) );
  XNOR U8731 ( .A(n8526), .B(n8525), .Z(n8584) );
  NANDN U8732 ( .A(n8501), .B(n8500), .Z(n8505) );
  NAND U8733 ( .A(n8503), .B(n8502), .Z(n8504) );
  NAND U8734 ( .A(n8505), .B(n8504), .Z(n8585) );
  XNOR U8735 ( .A(n8584), .B(n8585), .Z(n8586) );
  XOR U8736 ( .A(n8587), .B(n8586), .Z(n8517) );
  NANDN U8737 ( .A(n8507), .B(n8506), .Z(n8511) );
  NANDN U8738 ( .A(n8509), .B(n8508), .Z(n8510) );
  NAND U8739 ( .A(n8511), .B(n8510), .Z(n8518) );
  XNOR U8740 ( .A(n8517), .B(n8518), .Z(n8519) );
  XNOR U8741 ( .A(n8520), .B(n8519), .Z(n8590) );
  XNOR U8742 ( .A(n8590), .B(sreg[228]), .Z(n8592) );
  NAND U8743 ( .A(n8512), .B(sreg[227]), .Z(n8516) );
  OR U8744 ( .A(n8514), .B(n8513), .Z(n8515) );
  AND U8745 ( .A(n8516), .B(n8515), .Z(n8591) );
  XOR U8746 ( .A(n8592), .B(n8591), .Z(c[228]) );
  NANDN U8747 ( .A(n8518), .B(n8517), .Z(n8522) );
  NAND U8748 ( .A(n8520), .B(n8519), .Z(n8521) );
  NAND U8749 ( .A(n8522), .B(n8521), .Z(n8598) );
  NANDN U8750 ( .A(n8524), .B(n8523), .Z(n8528) );
  OR U8751 ( .A(n8526), .B(n8525), .Z(n8527) );
  NAND U8752 ( .A(n8528), .B(n8527), .Z(n8665) );
  NANDN U8753 ( .A(n8530), .B(n8529), .Z(n8534) );
  OR U8754 ( .A(n8532), .B(n8531), .Z(n8533) );
  NAND U8755 ( .A(n8534), .B(n8533), .Z(n8653) );
  NAND U8756 ( .A(b[0]), .B(a[117]), .Z(n8535) );
  XNOR U8757 ( .A(b[1]), .B(n8535), .Z(n8537) );
  NAND U8758 ( .A(a[116]), .B(n72), .Z(n8536) );
  AND U8759 ( .A(n8537), .B(n8536), .Z(n8629) );
  XNOR U8760 ( .A(n10050), .B(n8688), .Z(n8638) );
  OR U8761 ( .A(n8638), .B(n10051), .Z(n8540) );
  NANDN U8762 ( .A(n8538), .B(n10070), .Z(n8539) );
  AND U8763 ( .A(n8540), .B(n8539), .Z(n8630) );
  XOR U8764 ( .A(n8629), .B(n8630), .Z(n8632) );
  NAND U8765 ( .A(a[101]), .B(b[15]), .Z(n8631) );
  XOR U8766 ( .A(n8632), .B(n8631), .Z(n8650) );
  XOR U8767 ( .A(n9622), .B(a[113]), .Z(n8641) );
  OR U8768 ( .A(n8641), .B(n9623), .Z(n8543) );
  NANDN U8769 ( .A(n8541), .B(n9680), .Z(n8542) );
  NAND U8770 ( .A(n8543), .B(n8542), .Z(n8626) );
  XOR U8771 ( .A(n9872), .B(a[111]), .Z(n8644) );
  NANDN U8772 ( .A(n8644), .B(n9746), .Z(n8546) );
  NANDN U8773 ( .A(n8544), .B(n9747), .Z(n8545) );
  NAND U8774 ( .A(n8546), .B(n8545), .Z(n8623) );
  XOR U8775 ( .A(n74), .B(a[115]), .Z(n8647) );
  NANDN U8776 ( .A(n8647), .B(n9485), .Z(n8549) );
  NANDN U8777 ( .A(n8547), .B(n9484), .Z(n8548) );
  AND U8778 ( .A(n8549), .B(n8548), .Z(n8624) );
  XNOR U8779 ( .A(n8623), .B(n8624), .Z(n8625) );
  XOR U8780 ( .A(n8626), .B(n8625), .Z(n8651) );
  XOR U8781 ( .A(n8650), .B(n8651), .Z(n8652) );
  XNOR U8782 ( .A(n8653), .B(n8652), .Z(n8601) );
  NAND U8783 ( .A(n8551), .B(n8550), .Z(n8555) );
  NAND U8784 ( .A(n8553), .B(n8552), .Z(n8554) );
  NAND U8785 ( .A(n8555), .B(n8554), .Z(n8602) );
  XOR U8786 ( .A(n8601), .B(n8602), .Z(n8604) );
  XNOR U8787 ( .A(n9967), .B(n8844), .Z(n8607) );
  OR U8788 ( .A(n8607), .B(n10020), .Z(n8558) );
  NANDN U8789 ( .A(n8556), .B(n9968), .Z(n8557) );
  NAND U8790 ( .A(n8558), .B(n8557), .Z(n8620) );
  XNOR U8791 ( .A(n75), .B(n8559), .Z(n8611) );
  OR U8792 ( .A(n8611), .B(n10106), .Z(n8562) );
  NANDN U8793 ( .A(n8560), .B(n10107), .Z(n8561) );
  NAND U8794 ( .A(n8562), .B(n8561), .Z(n8617) );
  XOR U8795 ( .A(n9984), .B(a[109]), .Z(n8614) );
  NANDN U8796 ( .A(n8614), .B(n9865), .Z(n8565) );
  NANDN U8797 ( .A(n8563), .B(n9930), .Z(n8564) );
  AND U8798 ( .A(n8565), .B(n8564), .Z(n8618) );
  XNOR U8799 ( .A(n8617), .B(n8618), .Z(n8619) );
  XNOR U8800 ( .A(n8620), .B(n8619), .Z(n8656) );
  NANDN U8801 ( .A(n8567), .B(n8566), .Z(n8571) );
  NAND U8802 ( .A(n8569), .B(n8568), .Z(n8570) );
  NAND U8803 ( .A(n8571), .B(n8570), .Z(n8657) );
  XNOR U8804 ( .A(n8656), .B(n8657), .Z(n8658) );
  NANDN U8805 ( .A(n8573), .B(n8572), .Z(n8577) );
  NAND U8806 ( .A(n8575), .B(n8574), .Z(n8576) );
  AND U8807 ( .A(n8577), .B(n8576), .Z(n8659) );
  XNOR U8808 ( .A(n8658), .B(n8659), .Z(n8603) );
  XNOR U8809 ( .A(n8604), .B(n8603), .Z(n8662) );
  NANDN U8810 ( .A(n8579), .B(n8578), .Z(n8583) );
  NAND U8811 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND U8812 ( .A(n8583), .B(n8582), .Z(n8663) );
  XNOR U8813 ( .A(n8662), .B(n8663), .Z(n8664) );
  XOR U8814 ( .A(n8665), .B(n8664), .Z(n8595) );
  NANDN U8815 ( .A(n8585), .B(n8584), .Z(n8589) );
  NANDN U8816 ( .A(n8587), .B(n8586), .Z(n8588) );
  NAND U8817 ( .A(n8589), .B(n8588), .Z(n8596) );
  XNOR U8818 ( .A(n8595), .B(n8596), .Z(n8597) );
  XNOR U8819 ( .A(n8598), .B(n8597), .Z(n8668) );
  XNOR U8820 ( .A(n8668), .B(sreg[229]), .Z(n8670) );
  NAND U8821 ( .A(n8590), .B(sreg[228]), .Z(n8594) );
  OR U8822 ( .A(n8592), .B(n8591), .Z(n8593) );
  AND U8823 ( .A(n8594), .B(n8593), .Z(n8669) );
  XOR U8824 ( .A(n8670), .B(n8669), .Z(c[229]) );
  NANDN U8825 ( .A(n8596), .B(n8595), .Z(n8600) );
  NAND U8826 ( .A(n8598), .B(n8597), .Z(n8599) );
  NAND U8827 ( .A(n8600), .B(n8599), .Z(n8676) );
  NANDN U8828 ( .A(n8602), .B(n8601), .Z(n8606) );
  OR U8829 ( .A(n8604), .B(n8603), .Z(n8605) );
  NAND U8830 ( .A(n8606), .B(n8605), .Z(n8743) );
  XNOR U8831 ( .A(n9967), .B(n8922), .Z(n8685) );
  OR U8832 ( .A(n8685), .B(n10020), .Z(n8609) );
  NANDN U8833 ( .A(n8607), .B(n9968), .Z(n8608) );
  NAND U8834 ( .A(n8609), .B(n8608), .Z(n8698) );
  XNOR U8835 ( .A(n75), .B(n8610), .Z(n8689) );
  OR U8836 ( .A(n8689), .B(n10106), .Z(n8613) );
  NANDN U8837 ( .A(n8611), .B(n10107), .Z(n8612) );
  NAND U8838 ( .A(n8613), .B(n8612), .Z(n8695) );
  XNOR U8839 ( .A(n9984), .B(n9077), .Z(n8692) );
  NANDN U8840 ( .A(n8692), .B(n9865), .Z(n8616) );
  NANDN U8841 ( .A(n8614), .B(n9930), .Z(n8615) );
  AND U8842 ( .A(n8616), .B(n8615), .Z(n8696) );
  XNOR U8843 ( .A(n8695), .B(n8696), .Z(n8697) );
  XNOR U8844 ( .A(n8698), .B(n8697), .Z(n8734) );
  NANDN U8845 ( .A(n8618), .B(n8617), .Z(n8622) );
  NAND U8846 ( .A(n8620), .B(n8619), .Z(n8621) );
  NAND U8847 ( .A(n8622), .B(n8621), .Z(n8735) );
  XNOR U8848 ( .A(n8734), .B(n8735), .Z(n8736) );
  NANDN U8849 ( .A(n8624), .B(n8623), .Z(n8628) );
  NAND U8850 ( .A(n8626), .B(n8625), .Z(n8627) );
  AND U8851 ( .A(n8628), .B(n8627), .Z(n8737) );
  XNOR U8852 ( .A(n8736), .B(n8737), .Z(n8681) );
  NANDN U8853 ( .A(n8630), .B(n8629), .Z(n8634) );
  OR U8854 ( .A(n8632), .B(n8631), .Z(n8633) );
  NAND U8855 ( .A(n8634), .B(n8633), .Z(n8731) );
  NAND U8856 ( .A(b[0]), .B(a[118]), .Z(n8635) );
  XNOR U8857 ( .A(b[1]), .B(n8635), .Z(n8637) );
  NAND U8858 ( .A(a[117]), .B(n72), .Z(n8636) );
  AND U8859 ( .A(n8637), .B(n8636), .Z(n8707) );
  XNOR U8860 ( .A(n10050), .B(n8793), .Z(n8713) );
  OR U8861 ( .A(n8713), .B(n10051), .Z(n8640) );
  NANDN U8862 ( .A(n8638), .B(n10070), .Z(n8639) );
  AND U8863 ( .A(n8640), .B(n8639), .Z(n8708) );
  XOR U8864 ( .A(n8707), .B(n8708), .Z(n8710) );
  NAND U8865 ( .A(a[102]), .B(b[15]), .Z(n8709) );
  XOR U8866 ( .A(n8710), .B(n8709), .Z(n8728) );
  XNOR U8867 ( .A(n9622), .B(n9397), .Z(n8719) );
  OR U8868 ( .A(n8719), .B(n9623), .Z(n8643) );
  NANDN U8869 ( .A(n8641), .B(n9680), .Z(n8642) );
  NAND U8870 ( .A(n8643), .B(n8642), .Z(n8704) );
  XOR U8871 ( .A(n9872), .B(a[112]), .Z(n8722) );
  NANDN U8872 ( .A(n8722), .B(n9746), .Z(n8646) );
  NANDN U8873 ( .A(n8644), .B(n9747), .Z(n8645) );
  NAND U8874 ( .A(n8646), .B(n8645), .Z(n8701) );
  IV U8875 ( .A(a[116]), .Z(n9542) );
  XNOR U8876 ( .A(n9542), .B(n74), .Z(n8725) );
  NANDN U8877 ( .A(n8725), .B(n9485), .Z(n8649) );
  NANDN U8878 ( .A(n8647), .B(n9484), .Z(n8648) );
  AND U8879 ( .A(n8649), .B(n8648), .Z(n8702) );
  XNOR U8880 ( .A(n8701), .B(n8702), .Z(n8703) );
  XOR U8881 ( .A(n8704), .B(n8703), .Z(n8729) );
  XOR U8882 ( .A(n8728), .B(n8729), .Z(n8730) );
  XNOR U8883 ( .A(n8731), .B(n8730), .Z(n8679) );
  NAND U8884 ( .A(n8651), .B(n8650), .Z(n8655) );
  NAND U8885 ( .A(n8653), .B(n8652), .Z(n8654) );
  NAND U8886 ( .A(n8655), .B(n8654), .Z(n8680) );
  XOR U8887 ( .A(n8679), .B(n8680), .Z(n8682) );
  XNOR U8888 ( .A(n8681), .B(n8682), .Z(n8740) );
  NANDN U8889 ( .A(n8657), .B(n8656), .Z(n8661) );
  NAND U8890 ( .A(n8659), .B(n8658), .Z(n8660) );
  NAND U8891 ( .A(n8661), .B(n8660), .Z(n8741) );
  XNOR U8892 ( .A(n8740), .B(n8741), .Z(n8742) );
  XOR U8893 ( .A(n8743), .B(n8742), .Z(n8673) );
  NANDN U8894 ( .A(n8663), .B(n8662), .Z(n8667) );
  NANDN U8895 ( .A(n8665), .B(n8664), .Z(n8666) );
  NAND U8896 ( .A(n8667), .B(n8666), .Z(n8674) );
  XNOR U8897 ( .A(n8673), .B(n8674), .Z(n8675) );
  XNOR U8898 ( .A(n8676), .B(n8675), .Z(n8746) );
  XNOR U8899 ( .A(n8746), .B(sreg[230]), .Z(n8748) );
  NAND U8900 ( .A(n8668), .B(sreg[229]), .Z(n8672) );
  OR U8901 ( .A(n8670), .B(n8669), .Z(n8671) );
  AND U8902 ( .A(n8672), .B(n8671), .Z(n8747) );
  XOR U8903 ( .A(n8748), .B(n8747), .Z(c[230]) );
  NANDN U8904 ( .A(n8674), .B(n8673), .Z(n8678) );
  NAND U8905 ( .A(n8676), .B(n8675), .Z(n8677) );
  NAND U8906 ( .A(n8678), .B(n8677), .Z(n8754) );
  NANDN U8907 ( .A(n8680), .B(n8679), .Z(n8684) );
  OR U8908 ( .A(n8682), .B(n8681), .Z(n8683) );
  NAND U8909 ( .A(n8684), .B(n8683), .Z(n8821) );
  XOR U8910 ( .A(n9967), .B(a[109]), .Z(n8790) );
  OR U8911 ( .A(n8790), .B(n10020), .Z(n8687) );
  NANDN U8912 ( .A(n8685), .B(n9968), .Z(n8686) );
  NAND U8913 ( .A(n8687), .B(n8686), .Z(n8803) );
  XNOR U8914 ( .A(n75), .B(n8688), .Z(n8794) );
  OR U8915 ( .A(n8794), .B(n10106), .Z(n8691) );
  NANDN U8916 ( .A(n8689), .B(n10107), .Z(n8690) );
  NAND U8917 ( .A(n8691), .B(n8690), .Z(n8800) );
  XOR U8918 ( .A(n9984), .B(a[111]), .Z(n8797) );
  NANDN U8919 ( .A(n8797), .B(n9865), .Z(n8694) );
  NANDN U8920 ( .A(n8692), .B(n9930), .Z(n8693) );
  AND U8921 ( .A(n8694), .B(n8693), .Z(n8801) );
  XNOR U8922 ( .A(n8800), .B(n8801), .Z(n8802) );
  XNOR U8923 ( .A(n8803), .B(n8802), .Z(n8812) );
  NANDN U8924 ( .A(n8696), .B(n8695), .Z(n8700) );
  NAND U8925 ( .A(n8698), .B(n8697), .Z(n8699) );
  NAND U8926 ( .A(n8700), .B(n8699), .Z(n8813) );
  XNOR U8927 ( .A(n8812), .B(n8813), .Z(n8814) );
  NANDN U8928 ( .A(n8702), .B(n8701), .Z(n8706) );
  NAND U8929 ( .A(n8704), .B(n8703), .Z(n8705) );
  AND U8930 ( .A(n8706), .B(n8705), .Z(n8815) );
  XNOR U8931 ( .A(n8814), .B(n8815), .Z(n8759) );
  NANDN U8932 ( .A(n8708), .B(n8707), .Z(n8712) );
  OR U8933 ( .A(n8710), .B(n8709), .Z(n8711) );
  NAND U8934 ( .A(n8712), .B(n8711), .Z(n8787) );
  XNOR U8935 ( .A(n10050), .B(n8844), .Z(n8772) );
  OR U8936 ( .A(n8772), .B(n10051), .Z(n8715) );
  NANDN U8937 ( .A(n8713), .B(n10070), .Z(n8714) );
  AND U8938 ( .A(n8715), .B(n8714), .Z(n8764) );
  NAND U8939 ( .A(b[0]), .B(a[119]), .Z(n8716) );
  XNOR U8940 ( .A(b[1]), .B(n8716), .Z(n8718) );
  NAND U8941 ( .A(a[118]), .B(n72), .Z(n8717) );
  AND U8942 ( .A(n8718), .B(n8717), .Z(n8763) );
  XOR U8943 ( .A(n8764), .B(n8763), .Z(n8766) );
  NAND U8944 ( .A(a[103]), .B(b[15]), .Z(n8765) );
  XOR U8945 ( .A(n8766), .B(n8765), .Z(n8784) );
  XOR U8946 ( .A(n9622), .B(a[115]), .Z(n8775) );
  OR U8947 ( .A(n8775), .B(n9623), .Z(n8721) );
  NANDN U8948 ( .A(n8719), .B(n9680), .Z(n8720) );
  NAND U8949 ( .A(n8721), .B(n8720), .Z(n8809) );
  XOR U8950 ( .A(n9872), .B(a[113]), .Z(n8778) );
  NANDN U8951 ( .A(n8778), .B(n9746), .Z(n8724) );
  NANDN U8952 ( .A(n8722), .B(n9747), .Z(n8723) );
  NAND U8953 ( .A(n8724), .B(n8723), .Z(n8806) );
  IV U8954 ( .A(a[117]), .Z(n9631) );
  XNOR U8955 ( .A(n74), .B(n9631), .Z(n8781) );
  NANDN U8956 ( .A(n8781), .B(n9485), .Z(n8727) );
  NANDN U8957 ( .A(n8725), .B(n9484), .Z(n8726) );
  AND U8958 ( .A(n8727), .B(n8726), .Z(n8807) );
  XNOR U8959 ( .A(n8806), .B(n8807), .Z(n8808) );
  XOR U8960 ( .A(n8809), .B(n8808), .Z(n8785) );
  XOR U8961 ( .A(n8784), .B(n8785), .Z(n8786) );
  XNOR U8962 ( .A(n8787), .B(n8786), .Z(n8757) );
  NAND U8963 ( .A(n8729), .B(n8728), .Z(n8733) );
  NAND U8964 ( .A(n8731), .B(n8730), .Z(n8732) );
  NAND U8965 ( .A(n8733), .B(n8732), .Z(n8758) );
  XOR U8966 ( .A(n8757), .B(n8758), .Z(n8760) );
  XNOR U8967 ( .A(n8759), .B(n8760), .Z(n8818) );
  NANDN U8968 ( .A(n8735), .B(n8734), .Z(n8739) );
  NAND U8969 ( .A(n8737), .B(n8736), .Z(n8738) );
  NAND U8970 ( .A(n8739), .B(n8738), .Z(n8819) );
  XNOR U8971 ( .A(n8818), .B(n8819), .Z(n8820) );
  XOR U8972 ( .A(n8821), .B(n8820), .Z(n8751) );
  NANDN U8973 ( .A(n8741), .B(n8740), .Z(n8745) );
  NANDN U8974 ( .A(n8743), .B(n8742), .Z(n8744) );
  NAND U8975 ( .A(n8745), .B(n8744), .Z(n8752) );
  XNOR U8976 ( .A(n8751), .B(n8752), .Z(n8753) );
  XNOR U8977 ( .A(n8754), .B(n8753), .Z(n8824) );
  XNOR U8978 ( .A(n8824), .B(sreg[231]), .Z(n8826) );
  NAND U8979 ( .A(n8746), .B(sreg[230]), .Z(n8750) );
  OR U8980 ( .A(n8748), .B(n8747), .Z(n8749) );
  AND U8981 ( .A(n8750), .B(n8749), .Z(n8825) );
  XOR U8982 ( .A(n8826), .B(n8825), .Z(c[231]) );
  NANDN U8983 ( .A(n8752), .B(n8751), .Z(n8756) );
  NAND U8984 ( .A(n8754), .B(n8753), .Z(n8755) );
  NAND U8985 ( .A(n8756), .B(n8755), .Z(n8832) );
  NANDN U8986 ( .A(n8758), .B(n8757), .Z(n8762) );
  OR U8987 ( .A(n8760), .B(n8759), .Z(n8761) );
  NAND U8988 ( .A(n8762), .B(n8761), .Z(n8899) );
  NANDN U8989 ( .A(n8764), .B(n8763), .Z(n8768) );
  OR U8990 ( .A(n8766), .B(n8765), .Z(n8767) );
  NAND U8991 ( .A(n8768), .B(n8767), .Z(n8887) );
  NAND U8992 ( .A(b[0]), .B(a[120]), .Z(n8769) );
  XNOR U8993 ( .A(b[1]), .B(n8769), .Z(n8771) );
  NAND U8994 ( .A(a[119]), .B(n72), .Z(n8770) );
  AND U8995 ( .A(n8771), .B(n8770), .Z(n8863) );
  XNOR U8996 ( .A(n10050), .B(n8922), .Z(n8872) );
  OR U8997 ( .A(n8872), .B(n10051), .Z(n8774) );
  NANDN U8998 ( .A(n8772), .B(n10070), .Z(n8773) );
  AND U8999 ( .A(n8774), .B(n8773), .Z(n8864) );
  XOR U9000 ( .A(n8863), .B(n8864), .Z(n8866) );
  NAND U9001 ( .A(a[104]), .B(b[15]), .Z(n8865) );
  XOR U9002 ( .A(n8866), .B(n8865), .Z(n8884) );
  XNOR U9003 ( .A(n9622), .B(n9542), .Z(n8875) );
  OR U9004 ( .A(n8875), .B(n9623), .Z(n8777) );
  NANDN U9005 ( .A(n8775), .B(n9680), .Z(n8776) );
  NAND U9006 ( .A(n8777), .B(n8776), .Z(n8860) );
  XNOR U9007 ( .A(n9872), .B(n9397), .Z(n8878) );
  NANDN U9008 ( .A(n8878), .B(n9746), .Z(n8780) );
  NANDN U9009 ( .A(n8778), .B(n9747), .Z(n8779) );
  NAND U9010 ( .A(n8780), .B(n8779), .Z(n8857) );
  IV U9011 ( .A(a[118]), .Z(n9684) );
  XNOR U9012 ( .A(n9684), .B(n74), .Z(n8881) );
  NANDN U9013 ( .A(n8881), .B(n9485), .Z(n8783) );
  NANDN U9014 ( .A(n8781), .B(n9484), .Z(n8782) );
  AND U9015 ( .A(n8783), .B(n8782), .Z(n8858) );
  XNOR U9016 ( .A(n8857), .B(n8858), .Z(n8859) );
  XOR U9017 ( .A(n8860), .B(n8859), .Z(n8885) );
  XOR U9018 ( .A(n8884), .B(n8885), .Z(n8886) );
  XNOR U9019 ( .A(n8887), .B(n8886), .Z(n8835) );
  NAND U9020 ( .A(n8785), .B(n8784), .Z(n8789) );
  NAND U9021 ( .A(n8787), .B(n8786), .Z(n8788) );
  NAND U9022 ( .A(n8789), .B(n8788), .Z(n8836) );
  XOR U9023 ( .A(n8835), .B(n8836), .Z(n8838) );
  XNOR U9024 ( .A(n9967), .B(n9077), .Z(n8841) );
  OR U9025 ( .A(n8841), .B(n10020), .Z(n8792) );
  NANDN U9026 ( .A(n8790), .B(n9968), .Z(n8791) );
  NAND U9027 ( .A(n8792), .B(n8791), .Z(n8854) );
  XNOR U9028 ( .A(n75), .B(n8793), .Z(n8845) );
  OR U9029 ( .A(n8845), .B(n10106), .Z(n8796) );
  NANDN U9030 ( .A(n8794), .B(n10107), .Z(n8795) );
  NAND U9031 ( .A(n8796), .B(n8795), .Z(n8851) );
  XOR U9032 ( .A(n9984), .B(a[112]), .Z(n8848) );
  NANDN U9033 ( .A(n8848), .B(n9865), .Z(n8799) );
  NANDN U9034 ( .A(n8797), .B(n9930), .Z(n8798) );
  AND U9035 ( .A(n8799), .B(n8798), .Z(n8852) );
  XNOR U9036 ( .A(n8851), .B(n8852), .Z(n8853) );
  XNOR U9037 ( .A(n8854), .B(n8853), .Z(n8890) );
  NANDN U9038 ( .A(n8801), .B(n8800), .Z(n8805) );
  NAND U9039 ( .A(n8803), .B(n8802), .Z(n8804) );
  NAND U9040 ( .A(n8805), .B(n8804), .Z(n8891) );
  XNOR U9041 ( .A(n8890), .B(n8891), .Z(n8892) );
  NANDN U9042 ( .A(n8807), .B(n8806), .Z(n8811) );
  NAND U9043 ( .A(n8809), .B(n8808), .Z(n8810) );
  AND U9044 ( .A(n8811), .B(n8810), .Z(n8893) );
  XNOR U9045 ( .A(n8892), .B(n8893), .Z(n8837) );
  XNOR U9046 ( .A(n8838), .B(n8837), .Z(n8896) );
  NANDN U9047 ( .A(n8813), .B(n8812), .Z(n8817) );
  NAND U9048 ( .A(n8815), .B(n8814), .Z(n8816) );
  NAND U9049 ( .A(n8817), .B(n8816), .Z(n8897) );
  XNOR U9050 ( .A(n8896), .B(n8897), .Z(n8898) );
  XOR U9051 ( .A(n8899), .B(n8898), .Z(n8829) );
  NANDN U9052 ( .A(n8819), .B(n8818), .Z(n8823) );
  NANDN U9053 ( .A(n8821), .B(n8820), .Z(n8822) );
  NAND U9054 ( .A(n8823), .B(n8822), .Z(n8830) );
  XNOR U9055 ( .A(n8829), .B(n8830), .Z(n8831) );
  XNOR U9056 ( .A(n8832), .B(n8831), .Z(n8902) );
  XNOR U9057 ( .A(n8902), .B(sreg[232]), .Z(n8904) );
  NAND U9058 ( .A(n8824), .B(sreg[231]), .Z(n8828) );
  OR U9059 ( .A(n8826), .B(n8825), .Z(n8827) );
  AND U9060 ( .A(n8828), .B(n8827), .Z(n8903) );
  XOR U9061 ( .A(n8904), .B(n8903), .Z(c[232]) );
  NANDN U9062 ( .A(n8830), .B(n8829), .Z(n8834) );
  NAND U9063 ( .A(n8832), .B(n8831), .Z(n8833) );
  NAND U9064 ( .A(n8834), .B(n8833), .Z(n8910) );
  NANDN U9065 ( .A(n8836), .B(n8835), .Z(n8840) );
  OR U9066 ( .A(n8838), .B(n8837), .Z(n8839) );
  NAND U9067 ( .A(n8840), .B(n8839), .Z(n8977) );
  XOR U9068 ( .A(n9967), .B(a[111]), .Z(n8919) );
  OR U9069 ( .A(n8919), .B(n10020), .Z(n8843) );
  NANDN U9070 ( .A(n8841), .B(n9968), .Z(n8842) );
  NAND U9071 ( .A(n8843), .B(n8842), .Z(n8932) );
  XNOR U9072 ( .A(n75), .B(n8844), .Z(n8923) );
  OR U9073 ( .A(n8923), .B(n10106), .Z(n8847) );
  NANDN U9074 ( .A(n8845), .B(n10107), .Z(n8846) );
  NAND U9075 ( .A(n8847), .B(n8846), .Z(n8929) );
  XOR U9076 ( .A(n9984), .B(a[113]), .Z(n8926) );
  NANDN U9077 ( .A(n8926), .B(n9865), .Z(n8850) );
  NANDN U9078 ( .A(n8848), .B(n9930), .Z(n8849) );
  AND U9079 ( .A(n8850), .B(n8849), .Z(n8930) );
  XNOR U9080 ( .A(n8929), .B(n8930), .Z(n8931) );
  XNOR U9081 ( .A(n8932), .B(n8931), .Z(n8968) );
  NANDN U9082 ( .A(n8852), .B(n8851), .Z(n8856) );
  NAND U9083 ( .A(n8854), .B(n8853), .Z(n8855) );
  NAND U9084 ( .A(n8856), .B(n8855), .Z(n8969) );
  XNOR U9085 ( .A(n8968), .B(n8969), .Z(n8970) );
  NANDN U9086 ( .A(n8858), .B(n8857), .Z(n8862) );
  NAND U9087 ( .A(n8860), .B(n8859), .Z(n8861) );
  AND U9088 ( .A(n8862), .B(n8861), .Z(n8971) );
  XNOR U9089 ( .A(n8970), .B(n8971), .Z(n8915) );
  NANDN U9090 ( .A(n8864), .B(n8863), .Z(n8868) );
  OR U9091 ( .A(n8866), .B(n8865), .Z(n8867) );
  NAND U9092 ( .A(n8868), .B(n8867), .Z(n8965) );
  NAND U9093 ( .A(b[0]), .B(a[121]), .Z(n8869) );
  XNOR U9094 ( .A(b[1]), .B(n8869), .Z(n8871) );
  NAND U9095 ( .A(a[120]), .B(n72), .Z(n8870) );
  AND U9096 ( .A(n8871), .B(n8870), .Z(n8941) );
  XOR U9097 ( .A(n10050), .B(a[109]), .Z(n8950) );
  OR U9098 ( .A(n8950), .B(n10051), .Z(n8874) );
  NANDN U9099 ( .A(n8872), .B(n10070), .Z(n8873) );
  AND U9100 ( .A(n8874), .B(n8873), .Z(n8942) );
  XOR U9101 ( .A(n8941), .B(n8942), .Z(n8944) );
  NAND U9102 ( .A(a[105]), .B(b[15]), .Z(n8943) );
  XOR U9103 ( .A(n8944), .B(n8943), .Z(n8962) );
  XNOR U9104 ( .A(n9622), .B(n9631), .Z(n8953) );
  OR U9105 ( .A(n8953), .B(n9623), .Z(n8877) );
  NANDN U9106 ( .A(n8875), .B(n9680), .Z(n8876) );
  NAND U9107 ( .A(n8877), .B(n8876), .Z(n8938) );
  XOR U9108 ( .A(n9872), .B(a[115]), .Z(n8956) );
  NANDN U9109 ( .A(n8956), .B(n9746), .Z(n8880) );
  NANDN U9110 ( .A(n8878), .B(n9747), .Z(n8879) );
  NAND U9111 ( .A(n8880), .B(n8879), .Z(n8935) );
  IV U9112 ( .A(a[119]), .Z(n9755) );
  XNOR U9113 ( .A(n9755), .B(n74), .Z(n8959) );
  NANDN U9114 ( .A(n8959), .B(n9485), .Z(n8883) );
  NANDN U9115 ( .A(n8881), .B(n9484), .Z(n8882) );
  AND U9116 ( .A(n8883), .B(n8882), .Z(n8936) );
  XNOR U9117 ( .A(n8935), .B(n8936), .Z(n8937) );
  XOR U9118 ( .A(n8938), .B(n8937), .Z(n8963) );
  XOR U9119 ( .A(n8962), .B(n8963), .Z(n8964) );
  XNOR U9120 ( .A(n8965), .B(n8964), .Z(n8913) );
  NAND U9121 ( .A(n8885), .B(n8884), .Z(n8889) );
  NAND U9122 ( .A(n8887), .B(n8886), .Z(n8888) );
  NAND U9123 ( .A(n8889), .B(n8888), .Z(n8914) );
  XOR U9124 ( .A(n8913), .B(n8914), .Z(n8916) );
  XNOR U9125 ( .A(n8915), .B(n8916), .Z(n8974) );
  NANDN U9126 ( .A(n8891), .B(n8890), .Z(n8895) );
  NAND U9127 ( .A(n8893), .B(n8892), .Z(n8894) );
  NAND U9128 ( .A(n8895), .B(n8894), .Z(n8975) );
  XNOR U9129 ( .A(n8974), .B(n8975), .Z(n8976) );
  XOR U9130 ( .A(n8977), .B(n8976), .Z(n8907) );
  NANDN U9131 ( .A(n8897), .B(n8896), .Z(n8901) );
  NANDN U9132 ( .A(n8899), .B(n8898), .Z(n8900) );
  NAND U9133 ( .A(n8901), .B(n8900), .Z(n8908) );
  XNOR U9134 ( .A(n8907), .B(n8908), .Z(n8909) );
  XNOR U9135 ( .A(n8910), .B(n8909), .Z(n8980) );
  XNOR U9136 ( .A(n8980), .B(sreg[233]), .Z(n8982) );
  NAND U9137 ( .A(n8902), .B(sreg[232]), .Z(n8906) );
  OR U9138 ( .A(n8904), .B(n8903), .Z(n8905) );
  AND U9139 ( .A(n8906), .B(n8905), .Z(n8981) );
  XOR U9140 ( .A(n8982), .B(n8981), .Z(c[233]) );
  NANDN U9141 ( .A(n8908), .B(n8907), .Z(n8912) );
  NAND U9142 ( .A(n8910), .B(n8909), .Z(n8911) );
  NAND U9143 ( .A(n8912), .B(n8911), .Z(n8988) );
  NANDN U9144 ( .A(n8914), .B(n8913), .Z(n8918) );
  OR U9145 ( .A(n8916), .B(n8915), .Z(n8917) );
  NAND U9146 ( .A(n8918), .B(n8917), .Z(n9054) );
  XOR U9147 ( .A(n9967), .B(a[112]), .Z(n9024) );
  OR U9148 ( .A(n9024), .B(n10020), .Z(n8921) );
  NANDN U9149 ( .A(n8919), .B(n9968), .Z(n8920) );
  NAND U9150 ( .A(n8921), .B(n8920), .Z(n9036) );
  XNOR U9151 ( .A(n75), .B(n8922), .Z(n9027) );
  OR U9152 ( .A(n9027), .B(n10106), .Z(n8925) );
  NANDN U9153 ( .A(n8923), .B(n10107), .Z(n8924) );
  NAND U9154 ( .A(n8925), .B(n8924), .Z(n9033) );
  XNOR U9155 ( .A(n9984), .B(n9397), .Z(n9030) );
  NANDN U9156 ( .A(n9030), .B(n9865), .Z(n8928) );
  NANDN U9157 ( .A(n8926), .B(n9930), .Z(n8927) );
  AND U9158 ( .A(n8928), .B(n8927), .Z(n9034) );
  XNOR U9159 ( .A(n9033), .B(n9034), .Z(n9035) );
  XNOR U9160 ( .A(n9036), .B(n9035), .Z(n9045) );
  NANDN U9161 ( .A(n8930), .B(n8929), .Z(n8934) );
  NAND U9162 ( .A(n8932), .B(n8931), .Z(n8933) );
  NAND U9163 ( .A(n8934), .B(n8933), .Z(n9046) );
  XNOR U9164 ( .A(n9045), .B(n9046), .Z(n9047) );
  NANDN U9165 ( .A(n8936), .B(n8935), .Z(n8940) );
  NAND U9166 ( .A(n8938), .B(n8937), .Z(n8939) );
  AND U9167 ( .A(n8940), .B(n8939), .Z(n9048) );
  XNOR U9168 ( .A(n9047), .B(n9048), .Z(n8993) );
  NANDN U9169 ( .A(n8942), .B(n8941), .Z(n8946) );
  OR U9170 ( .A(n8944), .B(n8943), .Z(n8945) );
  NAND U9171 ( .A(n8946), .B(n8945), .Z(n9021) );
  NAND U9172 ( .A(b[0]), .B(a[122]), .Z(n8947) );
  XNOR U9173 ( .A(b[1]), .B(n8947), .Z(n8949) );
  NAND U9174 ( .A(n72), .B(a[121]), .Z(n8948) );
  AND U9175 ( .A(n8949), .B(n8948), .Z(n8997) );
  XNOR U9176 ( .A(n10050), .B(n9077), .Z(n9006) );
  OR U9177 ( .A(n9006), .B(n10051), .Z(n8952) );
  NANDN U9178 ( .A(n8950), .B(n10070), .Z(n8951) );
  AND U9179 ( .A(n8952), .B(n8951), .Z(n8998) );
  XOR U9180 ( .A(n8997), .B(n8998), .Z(n9000) );
  NAND U9181 ( .A(a[106]), .B(b[15]), .Z(n8999) );
  XOR U9182 ( .A(n9000), .B(n8999), .Z(n9018) );
  XNOR U9183 ( .A(n9622), .B(n9684), .Z(n9009) );
  OR U9184 ( .A(n9009), .B(n9623), .Z(n8955) );
  NANDN U9185 ( .A(n8953), .B(n9680), .Z(n8954) );
  NAND U9186 ( .A(n8955), .B(n8954), .Z(n9042) );
  XNOR U9187 ( .A(n9872), .B(n9542), .Z(n9012) );
  NANDN U9188 ( .A(n9012), .B(n9746), .Z(n8958) );
  NANDN U9189 ( .A(n8956), .B(n9747), .Z(n8957) );
  NAND U9190 ( .A(n8958), .B(n8957), .Z(n9039) );
  IV U9191 ( .A(a[120]), .Z(n9815) );
  XNOR U9192 ( .A(n9815), .B(n74), .Z(n9015) );
  NANDN U9193 ( .A(n9015), .B(n9485), .Z(n8961) );
  NANDN U9194 ( .A(n8959), .B(n9484), .Z(n8960) );
  AND U9195 ( .A(n8961), .B(n8960), .Z(n9040) );
  XNOR U9196 ( .A(n9039), .B(n9040), .Z(n9041) );
  XOR U9197 ( .A(n9042), .B(n9041), .Z(n9019) );
  XOR U9198 ( .A(n9018), .B(n9019), .Z(n9020) );
  XNOR U9199 ( .A(n9021), .B(n9020), .Z(n8991) );
  NAND U9200 ( .A(n8963), .B(n8962), .Z(n8967) );
  NAND U9201 ( .A(n8965), .B(n8964), .Z(n8966) );
  NAND U9202 ( .A(n8967), .B(n8966), .Z(n8992) );
  XOR U9203 ( .A(n8991), .B(n8992), .Z(n8994) );
  XNOR U9204 ( .A(n8993), .B(n8994), .Z(n9051) );
  NANDN U9205 ( .A(n8969), .B(n8968), .Z(n8973) );
  NAND U9206 ( .A(n8971), .B(n8970), .Z(n8972) );
  NAND U9207 ( .A(n8973), .B(n8972), .Z(n9052) );
  XNOR U9208 ( .A(n9051), .B(n9052), .Z(n9053) );
  XOR U9209 ( .A(n9054), .B(n9053), .Z(n8985) );
  NANDN U9210 ( .A(n8975), .B(n8974), .Z(n8979) );
  NANDN U9211 ( .A(n8977), .B(n8976), .Z(n8978) );
  NAND U9212 ( .A(n8979), .B(n8978), .Z(n8986) );
  XNOR U9213 ( .A(n8985), .B(n8986), .Z(n8987) );
  XNOR U9214 ( .A(n8988), .B(n8987), .Z(n9057) );
  XNOR U9215 ( .A(n9057), .B(sreg[234]), .Z(n9059) );
  NAND U9216 ( .A(n8980), .B(sreg[233]), .Z(n8984) );
  OR U9217 ( .A(n8982), .B(n8981), .Z(n8983) );
  AND U9218 ( .A(n8984), .B(n8983), .Z(n9058) );
  XOR U9219 ( .A(n9059), .B(n9058), .Z(c[234]) );
  NANDN U9220 ( .A(n8986), .B(n8985), .Z(n8990) );
  NAND U9221 ( .A(n8988), .B(n8987), .Z(n8989) );
  NAND U9222 ( .A(n8990), .B(n8989), .Z(n9065) );
  NANDN U9223 ( .A(n8992), .B(n8991), .Z(n8996) );
  OR U9224 ( .A(n8994), .B(n8993), .Z(n8995) );
  NAND U9225 ( .A(n8996), .B(n8995), .Z(n9132) );
  NANDN U9226 ( .A(n8998), .B(n8997), .Z(n9002) );
  OR U9227 ( .A(n9000), .B(n8999), .Z(n9001) );
  NAND U9228 ( .A(n9002), .B(n9001), .Z(n9120) );
  NAND U9229 ( .A(b[0]), .B(a[123]), .Z(n9003) );
  XNOR U9230 ( .A(b[1]), .B(n9003), .Z(n9005) );
  NAND U9231 ( .A(a[122]), .B(n72), .Z(n9004) );
  AND U9232 ( .A(n9005), .B(n9004), .Z(n9096) );
  XOR U9233 ( .A(n10050), .B(a[111]), .Z(n9105) );
  OR U9234 ( .A(n9105), .B(n10051), .Z(n9008) );
  NANDN U9235 ( .A(n9006), .B(n10070), .Z(n9007) );
  AND U9236 ( .A(n9008), .B(n9007), .Z(n9097) );
  XOR U9237 ( .A(n9096), .B(n9097), .Z(n9099) );
  NAND U9238 ( .A(a[107]), .B(b[15]), .Z(n9098) );
  XOR U9239 ( .A(n9099), .B(n9098), .Z(n9117) );
  XNOR U9240 ( .A(n9622), .B(n9755), .Z(n9108) );
  OR U9241 ( .A(n9108), .B(n9623), .Z(n9011) );
  NANDN U9242 ( .A(n9009), .B(n9680), .Z(n9010) );
  NAND U9243 ( .A(n9011), .B(n9010), .Z(n9093) );
  XNOR U9244 ( .A(n9872), .B(n9631), .Z(n9111) );
  NANDN U9245 ( .A(n9111), .B(n9746), .Z(n9014) );
  NANDN U9246 ( .A(n9012), .B(n9747), .Z(n9013) );
  NAND U9247 ( .A(n9014), .B(n9013), .Z(n9090) );
  XOR U9248 ( .A(a[121]), .B(n74), .Z(n9114) );
  NANDN U9249 ( .A(n9114), .B(n9485), .Z(n9017) );
  NANDN U9250 ( .A(n9015), .B(n9484), .Z(n9016) );
  AND U9251 ( .A(n9017), .B(n9016), .Z(n9091) );
  XNOR U9252 ( .A(n9090), .B(n9091), .Z(n9092) );
  XOR U9253 ( .A(n9093), .B(n9092), .Z(n9118) );
  XOR U9254 ( .A(n9117), .B(n9118), .Z(n9119) );
  XNOR U9255 ( .A(n9120), .B(n9119), .Z(n9068) );
  NAND U9256 ( .A(n9019), .B(n9018), .Z(n9023) );
  NAND U9257 ( .A(n9021), .B(n9020), .Z(n9022) );
  NAND U9258 ( .A(n9023), .B(n9022), .Z(n9069) );
  XOR U9259 ( .A(n9068), .B(n9069), .Z(n9071) );
  XOR U9260 ( .A(n9967), .B(a[113]), .Z(n9074) );
  OR U9261 ( .A(n9074), .B(n10020), .Z(n9026) );
  NANDN U9262 ( .A(n9024), .B(n9968), .Z(n9025) );
  NAND U9263 ( .A(n9026), .B(n9025), .Z(n9087) );
  XOR U9264 ( .A(n75), .B(a[109]), .Z(n9078) );
  OR U9265 ( .A(n9078), .B(n10106), .Z(n9029) );
  NANDN U9266 ( .A(n9027), .B(n10107), .Z(n9028) );
  NAND U9267 ( .A(n9029), .B(n9028), .Z(n9084) );
  XOR U9268 ( .A(n9984), .B(a[115]), .Z(n9081) );
  NANDN U9269 ( .A(n9081), .B(n9865), .Z(n9032) );
  NANDN U9270 ( .A(n9030), .B(n9930), .Z(n9031) );
  AND U9271 ( .A(n9032), .B(n9031), .Z(n9085) );
  XNOR U9272 ( .A(n9084), .B(n9085), .Z(n9086) );
  XNOR U9273 ( .A(n9087), .B(n9086), .Z(n9123) );
  NANDN U9274 ( .A(n9034), .B(n9033), .Z(n9038) );
  NAND U9275 ( .A(n9036), .B(n9035), .Z(n9037) );
  NAND U9276 ( .A(n9038), .B(n9037), .Z(n9124) );
  XNOR U9277 ( .A(n9123), .B(n9124), .Z(n9125) );
  NANDN U9278 ( .A(n9040), .B(n9039), .Z(n9044) );
  NAND U9279 ( .A(n9042), .B(n9041), .Z(n9043) );
  AND U9280 ( .A(n9044), .B(n9043), .Z(n9126) );
  XNOR U9281 ( .A(n9125), .B(n9126), .Z(n9070) );
  XNOR U9282 ( .A(n9071), .B(n9070), .Z(n9129) );
  NANDN U9283 ( .A(n9046), .B(n9045), .Z(n9050) );
  NAND U9284 ( .A(n9048), .B(n9047), .Z(n9049) );
  NAND U9285 ( .A(n9050), .B(n9049), .Z(n9130) );
  XNOR U9286 ( .A(n9129), .B(n9130), .Z(n9131) );
  XOR U9287 ( .A(n9132), .B(n9131), .Z(n9062) );
  NANDN U9288 ( .A(n9052), .B(n9051), .Z(n9056) );
  NANDN U9289 ( .A(n9054), .B(n9053), .Z(n9055) );
  NAND U9290 ( .A(n9056), .B(n9055), .Z(n9063) );
  XNOR U9291 ( .A(n9062), .B(n9063), .Z(n9064) );
  XNOR U9292 ( .A(n9065), .B(n9064), .Z(n9135) );
  XNOR U9293 ( .A(n9135), .B(sreg[235]), .Z(n9137) );
  NAND U9294 ( .A(n9057), .B(sreg[234]), .Z(n9061) );
  OR U9295 ( .A(n9059), .B(n9058), .Z(n9060) );
  AND U9296 ( .A(n9061), .B(n9060), .Z(n9136) );
  XOR U9297 ( .A(n9137), .B(n9136), .Z(c[235]) );
  NANDN U9298 ( .A(n9063), .B(n9062), .Z(n9067) );
  NAND U9299 ( .A(n9065), .B(n9064), .Z(n9066) );
  NAND U9300 ( .A(n9067), .B(n9066), .Z(n9143) );
  NANDN U9301 ( .A(n9069), .B(n9068), .Z(n9073) );
  OR U9302 ( .A(n9071), .B(n9070), .Z(n9072) );
  NAND U9303 ( .A(n9073), .B(n9072), .Z(n9209) );
  XNOR U9304 ( .A(n9967), .B(n9397), .Z(n9155) );
  OR U9305 ( .A(n9155), .B(n10020), .Z(n9076) );
  NANDN U9306 ( .A(n9074), .B(n9968), .Z(n9075) );
  NAND U9307 ( .A(n9076), .B(n9075), .Z(n9164) );
  XNOR U9308 ( .A(n75), .B(n9077), .Z(n9158) );
  OR U9309 ( .A(n9158), .B(n10106), .Z(n9080) );
  NANDN U9310 ( .A(n9078), .B(n10107), .Z(n9079) );
  NAND U9311 ( .A(n9080), .B(n9079), .Z(n9161) );
  XNOR U9312 ( .A(n9984), .B(n9542), .Z(n9152) );
  NANDN U9313 ( .A(n9152), .B(n9865), .Z(n9083) );
  NANDN U9314 ( .A(n9081), .B(n9930), .Z(n9082) );
  AND U9315 ( .A(n9083), .B(n9082), .Z(n9162) );
  XNOR U9316 ( .A(n9161), .B(n9162), .Z(n9163) );
  XNOR U9317 ( .A(n9164), .B(n9163), .Z(n9200) );
  NANDN U9318 ( .A(n9085), .B(n9084), .Z(n9089) );
  NAND U9319 ( .A(n9087), .B(n9086), .Z(n9088) );
  NAND U9320 ( .A(n9089), .B(n9088), .Z(n9201) );
  XNOR U9321 ( .A(n9200), .B(n9201), .Z(n9202) );
  NANDN U9322 ( .A(n9091), .B(n9090), .Z(n9095) );
  NAND U9323 ( .A(n9093), .B(n9092), .Z(n9094) );
  AND U9324 ( .A(n9095), .B(n9094), .Z(n9203) );
  XNOR U9325 ( .A(n9202), .B(n9203), .Z(n9148) );
  NANDN U9326 ( .A(n9097), .B(n9096), .Z(n9101) );
  OR U9327 ( .A(n9099), .B(n9098), .Z(n9100) );
  NAND U9328 ( .A(n9101), .B(n9100), .Z(n9197) );
  NAND U9329 ( .A(b[0]), .B(a[124]), .Z(n9102) );
  XNOR U9330 ( .A(b[1]), .B(n9102), .Z(n9104) );
  NAND U9331 ( .A(n72), .B(a[123]), .Z(n9103) );
  AND U9332 ( .A(n9104), .B(n9103), .Z(n9173) );
  XOR U9333 ( .A(n10050), .B(a[112]), .Z(n9182) );
  OR U9334 ( .A(n9182), .B(n10051), .Z(n9107) );
  NANDN U9335 ( .A(n9105), .B(n10070), .Z(n9106) );
  AND U9336 ( .A(n9107), .B(n9106), .Z(n9174) );
  XOR U9337 ( .A(n9173), .B(n9174), .Z(n9176) );
  NAND U9338 ( .A(a[108]), .B(b[15]), .Z(n9175) );
  XOR U9339 ( .A(n9176), .B(n9175), .Z(n9194) );
  XNOR U9340 ( .A(n9815), .B(n9622), .Z(n9188) );
  OR U9341 ( .A(n9188), .B(n9623), .Z(n9110) );
  NANDN U9342 ( .A(n9108), .B(n9680), .Z(n9109) );
  NAND U9343 ( .A(n9110), .B(n9109), .Z(n9170) );
  XNOR U9344 ( .A(n9872), .B(n9684), .Z(n9191) );
  NANDN U9345 ( .A(n9191), .B(n9746), .Z(n9113) );
  NANDN U9346 ( .A(n9111), .B(n9747), .Z(n9112) );
  NAND U9347 ( .A(n9113), .B(n9112), .Z(n9167) );
  IV U9348 ( .A(a[122]), .Z(n10023) );
  XNOR U9349 ( .A(n10023), .B(n74), .Z(n9185) );
  NANDN U9350 ( .A(n9185), .B(n9485), .Z(n9116) );
  NANDN U9351 ( .A(n9114), .B(n9484), .Z(n9115) );
  AND U9352 ( .A(n9116), .B(n9115), .Z(n9168) );
  XNOR U9353 ( .A(n9167), .B(n9168), .Z(n9169) );
  XOR U9354 ( .A(n9170), .B(n9169), .Z(n9195) );
  XOR U9355 ( .A(n9194), .B(n9195), .Z(n9196) );
  XNOR U9356 ( .A(n9197), .B(n9196), .Z(n9146) );
  NAND U9357 ( .A(n9118), .B(n9117), .Z(n9122) );
  NAND U9358 ( .A(n9120), .B(n9119), .Z(n9121) );
  NAND U9359 ( .A(n9122), .B(n9121), .Z(n9147) );
  XOR U9360 ( .A(n9146), .B(n9147), .Z(n9149) );
  XNOR U9361 ( .A(n9148), .B(n9149), .Z(n9206) );
  NANDN U9362 ( .A(n9124), .B(n9123), .Z(n9128) );
  NAND U9363 ( .A(n9126), .B(n9125), .Z(n9127) );
  NAND U9364 ( .A(n9128), .B(n9127), .Z(n9207) );
  XNOR U9365 ( .A(n9206), .B(n9207), .Z(n9208) );
  XOR U9366 ( .A(n9209), .B(n9208), .Z(n9140) );
  NANDN U9367 ( .A(n9130), .B(n9129), .Z(n9134) );
  NANDN U9368 ( .A(n9132), .B(n9131), .Z(n9133) );
  NAND U9369 ( .A(n9134), .B(n9133), .Z(n9141) );
  XNOR U9370 ( .A(n9140), .B(n9141), .Z(n9142) );
  XNOR U9371 ( .A(n9143), .B(n9142), .Z(n9212) );
  XNOR U9372 ( .A(n9212), .B(sreg[236]), .Z(n9214) );
  NAND U9373 ( .A(n9135), .B(sreg[235]), .Z(n9139) );
  OR U9374 ( .A(n9137), .B(n9136), .Z(n9138) );
  AND U9375 ( .A(n9139), .B(n9138), .Z(n9213) );
  XOR U9376 ( .A(n9214), .B(n9213), .Z(c[236]) );
  NANDN U9377 ( .A(n9141), .B(n9140), .Z(n9145) );
  NAND U9378 ( .A(n9143), .B(n9142), .Z(n9144) );
  NAND U9379 ( .A(n9145), .B(n9144), .Z(n9220) );
  NANDN U9380 ( .A(n9147), .B(n9146), .Z(n9151) );
  OR U9381 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U9382 ( .A(n9151), .B(n9150), .Z(n9286) );
  XNOR U9383 ( .A(n9984), .B(n9631), .Z(n9262) );
  NANDN U9384 ( .A(n9262), .B(n9865), .Z(n9154) );
  NANDN U9385 ( .A(n9152), .B(n9930), .Z(n9153) );
  NAND U9386 ( .A(n9154), .B(n9153), .Z(n9259) );
  XOR U9387 ( .A(n9967), .B(a[115]), .Z(n9265) );
  OR U9388 ( .A(n9265), .B(n10020), .Z(n9157) );
  NANDN U9389 ( .A(n9155), .B(n9968), .Z(n9156) );
  NAND U9390 ( .A(n9157), .B(n9156), .Z(n9256) );
  XOR U9391 ( .A(n75), .B(a[111]), .Z(n9268) );
  OR U9392 ( .A(n9268), .B(n10106), .Z(n9160) );
  NANDN U9393 ( .A(n9158), .B(n10107), .Z(n9159) );
  AND U9394 ( .A(n9160), .B(n9159), .Z(n9257) );
  XNOR U9395 ( .A(n9256), .B(n9257), .Z(n9258) );
  XNOR U9396 ( .A(n9259), .B(n9258), .Z(n9277) );
  NANDN U9397 ( .A(n9162), .B(n9161), .Z(n9166) );
  NAND U9398 ( .A(n9164), .B(n9163), .Z(n9165) );
  NAND U9399 ( .A(n9166), .B(n9165), .Z(n9278) );
  XNOR U9400 ( .A(n9277), .B(n9278), .Z(n9279) );
  NANDN U9401 ( .A(n9168), .B(n9167), .Z(n9172) );
  NAND U9402 ( .A(n9170), .B(n9169), .Z(n9171) );
  AND U9403 ( .A(n9172), .B(n9171), .Z(n9280) );
  XNOR U9404 ( .A(n9279), .B(n9280), .Z(n9225) );
  NANDN U9405 ( .A(n9174), .B(n9173), .Z(n9178) );
  OR U9406 ( .A(n9176), .B(n9175), .Z(n9177) );
  NAND U9407 ( .A(n9178), .B(n9177), .Z(n9274) );
  NAND U9408 ( .A(b[0]), .B(a[125]), .Z(n9179) );
  XNOR U9409 ( .A(b[1]), .B(n9179), .Z(n9181) );
  NAND U9410 ( .A(a[124]), .B(n72), .Z(n9180) );
  AND U9411 ( .A(n9181), .B(n9180), .Z(n9231) );
  XOR U9412 ( .A(b[13]), .B(a[113]), .Z(n9238) );
  NANDN U9413 ( .A(n10051), .B(n9238), .Z(n9184) );
  NANDN U9414 ( .A(n9182), .B(n10070), .Z(n9183) );
  NAND U9415 ( .A(n9184), .B(n9183), .Z(n9229) );
  NAND U9416 ( .A(b[15]), .B(a[109]), .Z(n9230) );
  XNOR U9417 ( .A(n9229), .B(n9230), .Z(n9232) );
  XOR U9418 ( .A(n9231), .B(n9232), .Z(n9271) );
  XOR U9419 ( .A(a[123]), .B(n74), .Z(n9241) );
  NANDN U9420 ( .A(n9241), .B(n9485), .Z(n9187) );
  NANDN U9421 ( .A(n9185), .B(n9484), .Z(n9186) );
  NAND U9422 ( .A(n9187), .B(n9186), .Z(n9252) );
  XOR U9423 ( .A(a[121]), .B(n9622), .Z(n9244) );
  OR U9424 ( .A(n9244), .B(n9623), .Z(n9190) );
  NANDN U9425 ( .A(n9188), .B(n9680), .Z(n9189) );
  NAND U9426 ( .A(n9190), .B(n9189), .Z(n9250) );
  XNOR U9427 ( .A(n9872), .B(n9755), .Z(n9247) );
  NANDN U9428 ( .A(n9247), .B(n9746), .Z(n9193) );
  NANDN U9429 ( .A(n9191), .B(n9747), .Z(n9192) );
  AND U9430 ( .A(n9193), .B(n9192), .Z(n9251) );
  XOR U9431 ( .A(n9252), .B(n9253), .Z(n9272) );
  XNOR U9432 ( .A(n9271), .B(n9272), .Z(n9273) );
  XNOR U9433 ( .A(n9274), .B(n9273), .Z(n9223) );
  NAND U9434 ( .A(n9195), .B(n9194), .Z(n9199) );
  NAND U9435 ( .A(n9197), .B(n9196), .Z(n9198) );
  NAND U9436 ( .A(n9199), .B(n9198), .Z(n9224) );
  XOR U9437 ( .A(n9223), .B(n9224), .Z(n9226) );
  XNOR U9438 ( .A(n9225), .B(n9226), .Z(n9283) );
  NANDN U9439 ( .A(n9201), .B(n9200), .Z(n9205) );
  NAND U9440 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U9441 ( .A(n9205), .B(n9204), .Z(n9284) );
  XNOR U9442 ( .A(n9283), .B(n9284), .Z(n9285) );
  XOR U9443 ( .A(n9286), .B(n9285), .Z(n9217) );
  NANDN U9444 ( .A(n9207), .B(n9206), .Z(n9211) );
  NANDN U9445 ( .A(n9209), .B(n9208), .Z(n9210) );
  NAND U9446 ( .A(n9211), .B(n9210), .Z(n9218) );
  XNOR U9447 ( .A(n9217), .B(n9218), .Z(n9219) );
  XNOR U9448 ( .A(n9220), .B(n9219), .Z(n9289) );
  XNOR U9449 ( .A(n9289), .B(sreg[237]), .Z(n9291) );
  NAND U9450 ( .A(n9212), .B(sreg[236]), .Z(n9216) );
  OR U9451 ( .A(n9214), .B(n9213), .Z(n9215) );
  AND U9452 ( .A(n9216), .B(n9215), .Z(n9290) );
  XOR U9453 ( .A(n9291), .B(n9290), .Z(c[237]) );
  NANDN U9454 ( .A(n9218), .B(n9217), .Z(n9222) );
  NAND U9455 ( .A(n9220), .B(n9219), .Z(n9221) );
  NAND U9456 ( .A(n9222), .B(n9221), .Z(n9297) );
  NANDN U9457 ( .A(n9224), .B(n9223), .Z(n9228) );
  OR U9458 ( .A(n9226), .B(n9225), .Z(n9227) );
  NAND U9459 ( .A(n9228), .B(n9227), .Z(n9303) );
  NANDN U9460 ( .A(n9230), .B(n9229), .Z(n9234) );
  NAND U9461 ( .A(n9232), .B(n9231), .Z(n9233) );
  NAND U9462 ( .A(n9234), .B(n9233), .Z(n9330) );
  AND U9463 ( .A(b[15]), .B(a[110]), .Z(n9324) );
  NAND U9464 ( .A(a[126]), .B(b[0]), .Z(n9235) );
  XNOR U9465 ( .A(b[1]), .B(n9235), .Z(n9237) );
  NAND U9466 ( .A(a[125]), .B(n72), .Z(n9236) );
  AND U9467 ( .A(n9237), .B(n9236), .Z(n9322) );
  NAND U9468 ( .A(n10070), .B(n9238), .Z(n9240) );
  XOR U9469 ( .A(b[13]), .B(a[114]), .Z(n9309) );
  NANDN U9470 ( .A(n10051), .B(n9309), .Z(n9239) );
  AND U9471 ( .A(n9240), .B(n9239), .Z(n9321) );
  XNOR U9472 ( .A(n9322), .B(n9321), .Z(n9323) );
  XOR U9473 ( .A(n9324), .B(n9323), .Z(n9327) );
  IV U9474 ( .A(a[124]), .Z(n9920) );
  XNOR U9475 ( .A(n9920), .B(n74), .Z(n9312) );
  NANDN U9476 ( .A(n9312), .B(n9485), .Z(n9243) );
  NANDN U9477 ( .A(n9241), .B(n9484), .Z(n9242) );
  NAND U9478 ( .A(n9243), .B(n9242), .Z(n9349) );
  XNOR U9479 ( .A(n10023), .B(n9622), .Z(n9315) );
  OR U9480 ( .A(n9315), .B(n9623), .Z(n9246) );
  NANDN U9481 ( .A(n9244), .B(n9680), .Z(n9245) );
  NAND U9482 ( .A(n9246), .B(n9245), .Z(n9346) );
  XNOR U9483 ( .A(n9872), .B(n9815), .Z(n9318) );
  NANDN U9484 ( .A(n9318), .B(n9746), .Z(n9249) );
  NANDN U9485 ( .A(n9247), .B(n9747), .Z(n9248) );
  AND U9486 ( .A(n9249), .B(n9248), .Z(n9347) );
  XNOR U9487 ( .A(n9346), .B(n9347), .Z(n9348) );
  XNOR U9488 ( .A(n9349), .B(n9348), .Z(n9328) );
  XOR U9489 ( .A(n9327), .B(n9328), .Z(n9329) );
  XOR U9490 ( .A(n9330), .B(n9329), .Z(n9355) );
  NANDN U9491 ( .A(n9251), .B(n9250), .Z(n9255) );
  NANDN U9492 ( .A(n9253), .B(n9252), .Z(n9254) );
  NAND U9493 ( .A(n9255), .B(n9254), .Z(n9361) );
  NANDN U9494 ( .A(n9257), .B(n9256), .Z(n9261) );
  NAND U9495 ( .A(n9259), .B(n9258), .Z(n9260) );
  NAND U9496 ( .A(n9261), .B(n9260), .Z(n9359) );
  XNOR U9497 ( .A(n9984), .B(n9684), .Z(n9331) );
  NANDN U9498 ( .A(n9331), .B(n9865), .Z(n9264) );
  NANDN U9499 ( .A(n9262), .B(n9930), .Z(n9263) );
  NAND U9500 ( .A(n9264), .B(n9263), .Z(n9343) );
  XNOR U9501 ( .A(n9967), .B(n9542), .Z(n9334) );
  OR U9502 ( .A(n9334), .B(n10020), .Z(n9267) );
  NANDN U9503 ( .A(n9265), .B(n9968), .Z(n9266) );
  NAND U9504 ( .A(n9267), .B(n9266), .Z(n9340) );
  XOR U9505 ( .A(n75), .B(a[112]), .Z(n9337) );
  OR U9506 ( .A(n9337), .B(n10106), .Z(n9270) );
  NANDN U9507 ( .A(n9268), .B(n10107), .Z(n9269) );
  AND U9508 ( .A(n9270), .B(n9269), .Z(n9341) );
  XNOR U9509 ( .A(n9340), .B(n9341), .Z(n9342) );
  XOR U9510 ( .A(n9343), .B(n9342), .Z(n9358) );
  XNOR U9511 ( .A(n9359), .B(n9358), .Z(n9360) );
  XNOR U9512 ( .A(n9361), .B(n9360), .Z(n9353) );
  NANDN U9513 ( .A(n9272), .B(n9271), .Z(n9276) );
  NAND U9514 ( .A(n9274), .B(n9273), .Z(n9275) );
  AND U9515 ( .A(n9276), .B(n9275), .Z(n9352) );
  XNOR U9516 ( .A(n9353), .B(n9352), .Z(n9354) );
  XOR U9517 ( .A(n9355), .B(n9354), .Z(n9300) );
  NANDN U9518 ( .A(n9278), .B(n9277), .Z(n9282) );
  NAND U9519 ( .A(n9280), .B(n9279), .Z(n9281) );
  NAND U9520 ( .A(n9282), .B(n9281), .Z(n9301) );
  XOR U9521 ( .A(n9300), .B(n9301), .Z(n9302) );
  XOR U9522 ( .A(n9303), .B(n9302), .Z(n9294) );
  NANDN U9523 ( .A(n9284), .B(n9283), .Z(n9288) );
  NANDN U9524 ( .A(n9286), .B(n9285), .Z(n9287) );
  NAND U9525 ( .A(n9288), .B(n9287), .Z(n9295) );
  XNOR U9526 ( .A(n9294), .B(n9295), .Z(n9296) );
  XNOR U9527 ( .A(n9297), .B(n9296), .Z(n9364) );
  XNOR U9528 ( .A(n9364), .B(sreg[238]), .Z(n9366) );
  NAND U9529 ( .A(n9289), .B(sreg[237]), .Z(n9293) );
  OR U9530 ( .A(n9291), .B(n9290), .Z(n9292) );
  AND U9531 ( .A(n9293), .B(n9292), .Z(n9365) );
  XOR U9532 ( .A(n9366), .B(n9365), .Z(c[238]) );
  NANDN U9533 ( .A(n9295), .B(n9294), .Z(n9299) );
  NAND U9534 ( .A(n9297), .B(n9296), .Z(n9298) );
  NAND U9535 ( .A(n9299), .B(n9298), .Z(n9372) );
  OR U9536 ( .A(n9301), .B(n9300), .Z(n9305) );
  NANDN U9537 ( .A(n9303), .B(n9302), .Z(n9304) );
  NAND U9538 ( .A(n9305), .B(n9304), .Z(n9370) );
  NAND U9539 ( .A(b[0]), .B(a[127]), .Z(n9306) );
  XNOR U9540 ( .A(b[1]), .B(n9306), .Z(n9308) );
  NAND U9541 ( .A(a[126]), .B(n72), .Z(n9307) );
  AND U9542 ( .A(n9308), .B(n9307), .Z(n9421) );
  XOR U9543 ( .A(n10050), .B(a[115]), .Z(n9434) );
  OR U9544 ( .A(n9434), .B(n10051), .Z(n9311) );
  NAND U9545 ( .A(n9309), .B(n10070), .Z(n9310) );
  NAND U9546 ( .A(n9311), .B(n9310), .Z(n9419) );
  NAND U9547 ( .A(b[15]), .B(a[111]), .Z(n9420) );
  XNOR U9548 ( .A(n9419), .B(n9420), .Z(n9422) );
  XOR U9549 ( .A(n9421), .B(n9422), .Z(n9413) );
  IV U9550 ( .A(a[125]), .Z(n9978) );
  XNOR U9551 ( .A(n9978), .B(n74), .Z(n9425) );
  NANDN U9552 ( .A(n9425), .B(n9485), .Z(n9314) );
  NANDN U9553 ( .A(n9312), .B(n9484), .Z(n9313) );
  NAND U9554 ( .A(n9314), .B(n9313), .Z(n9409) );
  XOR U9555 ( .A(a[123]), .B(n9622), .Z(n9428) );
  OR U9556 ( .A(n9428), .B(n9623), .Z(n9317) );
  NANDN U9557 ( .A(n9315), .B(n9680), .Z(n9316) );
  NAND U9558 ( .A(n9317), .B(n9316), .Z(n9407) );
  XOR U9559 ( .A(n9872), .B(a[121]), .Z(n9431) );
  NANDN U9560 ( .A(n9431), .B(n9746), .Z(n9320) );
  NANDN U9561 ( .A(n9318), .B(n9747), .Z(n9319) );
  AND U9562 ( .A(n9320), .B(n9319), .Z(n9408) );
  XOR U9563 ( .A(n9409), .B(n9410), .Z(n9414) );
  XNOR U9564 ( .A(n9413), .B(n9414), .Z(n9415) );
  NANDN U9565 ( .A(n9322), .B(n9321), .Z(n9326) );
  NANDN U9566 ( .A(n9324), .B(n9323), .Z(n9325) );
  NAND U9567 ( .A(n9326), .B(n9325), .Z(n9416) );
  XOR U9568 ( .A(n9415), .B(n9416), .Z(n9379) );
  XNOR U9569 ( .A(n9379), .B(n9380), .Z(n9381) );
  XNOR U9570 ( .A(n9984), .B(n9755), .Z(n9391) );
  NANDN U9571 ( .A(n9391), .B(n9865), .Z(n9333) );
  NANDN U9572 ( .A(n9331), .B(n9930), .Z(n9332) );
  NAND U9573 ( .A(n9333), .B(n9332), .Z(n9404) );
  XNOR U9574 ( .A(n9967), .B(n9631), .Z(n9394) );
  OR U9575 ( .A(n9394), .B(n10020), .Z(n9336) );
  NANDN U9576 ( .A(n9334), .B(n9968), .Z(n9335) );
  NAND U9577 ( .A(n9336), .B(n9335), .Z(n9401) );
  XOR U9578 ( .A(n75), .B(a[113]), .Z(n9398) );
  OR U9579 ( .A(n9398), .B(n10106), .Z(n9339) );
  NANDN U9580 ( .A(n9337), .B(n10107), .Z(n9338) );
  AND U9581 ( .A(n9339), .B(n9338), .Z(n9402) );
  XNOR U9582 ( .A(n9401), .B(n9402), .Z(n9403) );
  XNOR U9583 ( .A(n9404), .B(n9403), .Z(n9388) );
  NANDN U9584 ( .A(n9341), .B(n9340), .Z(n9345) );
  NAND U9585 ( .A(n9343), .B(n9342), .Z(n9344) );
  NAND U9586 ( .A(n9345), .B(n9344), .Z(n9386) );
  NANDN U9587 ( .A(n9347), .B(n9346), .Z(n9351) );
  NAND U9588 ( .A(n9349), .B(n9348), .Z(n9350) );
  AND U9589 ( .A(n9351), .B(n9350), .Z(n9385) );
  XNOR U9590 ( .A(n9386), .B(n9385), .Z(n9387) );
  XOR U9591 ( .A(n9388), .B(n9387), .Z(n9382) );
  XOR U9592 ( .A(n9381), .B(n9382), .Z(n9375) );
  NANDN U9593 ( .A(n9353), .B(n9352), .Z(n9357) );
  NAND U9594 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U9595 ( .A(n9357), .B(n9356), .Z(n9373) );
  OR U9596 ( .A(n9359), .B(n9358), .Z(n9363) );
  OR U9597 ( .A(n9361), .B(n9360), .Z(n9362) );
  AND U9598 ( .A(n9363), .B(n9362), .Z(n9374) );
  XNOR U9599 ( .A(n9373), .B(n9374), .Z(n9376) );
  XOR U9600 ( .A(n9375), .B(n9376), .Z(n9369) );
  XOR U9601 ( .A(n9370), .B(n9369), .Z(n9371) );
  XOR U9602 ( .A(n9372), .B(n9371), .Z(n9437) );
  XNOR U9603 ( .A(n9437), .B(sreg[239]), .Z(n9439) );
  NAND U9604 ( .A(n9364), .B(sreg[238]), .Z(n9368) );
  OR U9605 ( .A(n9366), .B(n9365), .Z(n9367) );
  AND U9606 ( .A(n9368), .B(n9367), .Z(n9438) );
  XOR U9607 ( .A(n9439), .B(n9438), .Z(c[239]) );
  NANDN U9608 ( .A(n9374), .B(n9373), .Z(n9378) );
  NAND U9609 ( .A(n9376), .B(n9375), .Z(n9377) );
  NAND U9610 ( .A(n9378), .B(n9377), .Z(n9445) );
  NANDN U9611 ( .A(n9380), .B(n9379), .Z(n9384) );
  NAND U9612 ( .A(n9382), .B(n9381), .Z(n9383) );
  NAND U9613 ( .A(n9384), .B(n9383), .Z(n9452) );
  NANDN U9614 ( .A(n9386), .B(n9385), .Z(n9390) );
  NAND U9615 ( .A(n9388), .B(n9387), .Z(n9389) );
  NAND U9616 ( .A(n9390), .B(n9389), .Z(n9451) );
  XNOR U9617 ( .A(n9984), .B(n9815), .Z(n9465) );
  NANDN U9618 ( .A(n9465), .B(n9865), .Z(n9393) );
  NANDN U9619 ( .A(n9391), .B(n9930), .Z(n9392) );
  NAND U9620 ( .A(n9393), .B(n9392), .Z(n9474) );
  XNOR U9621 ( .A(n9967), .B(n9684), .Z(n9468) );
  OR U9622 ( .A(n9468), .B(n10020), .Z(n9396) );
  NANDN U9623 ( .A(n9394), .B(n9968), .Z(n9395) );
  NAND U9624 ( .A(n9396), .B(n9395), .Z(n9471) );
  XNOR U9625 ( .A(b[15]), .B(n9397), .Z(n9497) );
  NANDN U9626 ( .A(n10106), .B(n9497), .Z(n9400) );
  NANDN U9627 ( .A(n9398), .B(n10107), .Z(n9399) );
  AND U9628 ( .A(n9400), .B(n9399), .Z(n9472) );
  XNOR U9629 ( .A(n9471), .B(n9472), .Z(n9473) );
  XOR U9630 ( .A(n9474), .B(n9473), .Z(n9512) );
  NANDN U9631 ( .A(n9402), .B(n9401), .Z(n9406) );
  NAND U9632 ( .A(n9404), .B(n9403), .Z(n9405) );
  NAND U9633 ( .A(n9406), .B(n9405), .Z(n9510) );
  NANDN U9634 ( .A(n9408), .B(n9407), .Z(n9412) );
  NANDN U9635 ( .A(n9410), .B(n9409), .Z(n9411) );
  NAND U9636 ( .A(n9412), .B(n9411), .Z(n9509) );
  XOR U9637 ( .A(n9510), .B(n9509), .Z(n9511) );
  XOR U9638 ( .A(n9512), .B(n9511), .Z(n9504) );
  NANDN U9639 ( .A(n9414), .B(n9413), .Z(n9418) );
  NANDN U9640 ( .A(n9416), .B(n9415), .Z(n9417) );
  AND U9641 ( .A(n9418), .B(n9417), .Z(n9503) );
  XNOR U9642 ( .A(n9504), .B(n9503), .Z(n9505) );
  NANDN U9643 ( .A(n9420), .B(n9419), .Z(n9424) );
  NAND U9644 ( .A(n9422), .B(n9421), .Z(n9423) );
  NAND U9645 ( .A(n9424), .B(n9423), .Z(n9479) );
  XNOR U9646 ( .A(a[126]), .B(n74), .Z(n9483) );
  NAND U9647 ( .A(n9483), .B(n9485), .Z(n9427) );
  NANDN U9648 ( .A(n9425), .B(n9484), .Z(n9426) );
  NAND U9649 ( .A(n9427), .B(n9426), .Z(n9459) );
  XNOR U9650 ( .A(a[124]), .B(n9622), .Z(n9488) );
  NANDN U9651 ( .A(n9623), .B(n9488), .Z(n9430) );
  NANDN U9652 ( .A(n9428), .B(n9680), .Z(n9429) );
  NAND U9653 ( .A(n9430), .B(n9429), .Z(n9456) );
  XNOR U9654 ( .A(n10023), .B(n9872), .Z(n9462) );
  NANDN U9655 ( .A(n9462), .B(n9746), .Z(n9433) );
  NANDN U9656 ( .A(n9431), .B(n9747), .Z(n9432) );
  AND U9657 ( .A(n9433), .B(n9432), .Z(n9457) );
  XNOR U9658 ( .A(n9456), .B(n9457), .Z(n9458) );
  XNOR U9659 ( .A(n9459), .B(n9458), .Z(n9477) );
  IV U9660 ( .A(a[127]), .Z(n10049) );
  XNOR U9661 ( .A(n10050), .B(n9542), .Z(n9500) );
  OR U9662 ( .A(n9500), .B(n10051), .Z(n9436) );
  NANDN U9663 ( .A(n9434), .B(n10070), .Z(n9435) );
  NAND U9664 ( .A(n9436), .B(n9435), .Z(n9491) );
  NAND U9665 ( .A(b[15]), .B(a[112]), .Z(n9492) );
  XNOR U9666 ( .A(n9491), .B(n9492), .Z(n9493) );
  XOR U9667 ( .A(n9494), .B(n9493), .Z(n9478) );
  XOR U9668 ( .A(n9477), .B(n9478), .Z(n9480) );
  XOR U9669 ( .A(n9479), .B(n9480), .Z(n9506) );
  XOR U9670 ( .A(n9505), .B(n9506), .Z(n9450) );
  XNOR U9671 ( .A(n9451), .B(n9450), .Z(n9453) );
  XNOR U9672 ( .A(n9452), .B(n9453), .Z(n9444) );
  XOR U9673 ( .A(n9445), .B(n9444), .Z(n9446) );
  XOR U9674 ( .A(n9447), .B(n9446), .Z(n9443) );
  NAND U9675 ( .A(n9437), .B(sreg[239]), .Z(n9441) );
  OR U9676 ( .A(n9439), .B(n9438), .Z(n9440) );
  AND U9677 ( .A(n9441), .B(n9440), .Z(n9442) );
  XOR U9678 ( .A(n9443), .B(n9442), .Z(c[240]) );
  OR U9679 ( .A(n9443), .B(n9442), .Z(n9586) );
  NAND U9680 ( .A(n9445), .B(n9444), .Z(n9449) );
  NAND U9681 ( .A(n9447), .B(n9446), .Z(n9448) );
  NAND U9682 ( .A(n9449), .B(n9448), .Z(n9581) );
  NAND U9683 ( .A(n9451), .B(n9450), .Z(n9455) );
  NANDN U9684 ( .A(n9453), .B(n9452), .Z(n9454) );
  NAND U9685 ( .A(n9455), .B(n9454), .Z(n9579) );
  NANDN U9686 ( .A(n9457), .B(n9456), .Z(n9461) );
  NAND U9687 ( .A(n9459), .B(n9458), .Z(n9460) );
  NAND U9688 ( .A(n9461), .B(n9460), .Z(n9517) );
  XOR U9689 ( .A(a[123]), .B(n9872), .Z(n9552) );
  NANDN U9690 ( .A(n9552), .B(n9746), .Z(n9464) );
  NANDN U9691 ( .A(n9462), .B(n9747), .Z(n9463) );
  NAND U9692 ( .A(n9464), .B(n9463), .Z(n9569) );
  XOR U9693 ( .A(n9984), .B(a[121]), .Z(n9549) );
  NANDN U9694 ( .A(n9549), .B(n9865), .Z(n9467) );
  NANDN U9695 ( .A(n9465), .B(n9930), .Z(n9466) );
  NAND U9696 ( .A(n9467), .B(n9466), .Z(n9566) );
  XNOR U9697 ( .A(n9967), .B(n9755), .Z(n9546) );
  OR U9698 ( .A(n9546), .B(n10020), .Z(n9470) );
  NANDN U9699 ( .A(n9468), .B(n9968), .Z(n9469) );
  AND U9700 ( .A(n9470), .B(n9469), .Z(n9567) );
  XNOR U9701 ( .A(n9566), .B(n9567), .Z(n9568) );
  XNOR U9702 ( .A(n9569), .B(n9568), .Z(n9515) );
  NANDN U9703 ( .A(n9472), .B(n9471), .Z(n9476) );
  NAND U9704 ( .A(n9474), .B(n9473), .Z(n9475) );
  NAND U9705 ( .A(n9476), .B(n9475), .Z(n9516) );
  XOR U9706 ( .A(n9515), .B(n9516), .Z(n9518) );
  XOR U9707 ( .A(n9517), .B(n9518), .Z(n9523) );
  NANDN U9708 ( .A(n9478), .B(n9477), .Z(n9482) );
  OR U9709 ( .A(n9480), .B(n9479), .Z(n9481) );
  NAND U9710 ( .A(n9482), .B(n9481), .Z(n9522) );
  NAND U9711 ( .A(n9484), .B(n9483), .Z(n9487) );
  XOR U9712 ( .A(a[127]), .B(b[3]), .Z(n9539) );
  NAND U9713 ( .A(n9539), .B(n9485), .Z(n9486) );
  NAND U9714 ( .A(n9487), .B(n9486), .Z(n9563) );
  NAND U9715 ( .A(n9680), .B(n9488), .Z(n9490) );
  XOR U9716 ( .A(a[125]), .B(b[5]), .Z(n9555) );
  NANDN U9717 ( .A(n9623), .B(n9555), .Z(n9489) );
  NAND U9718 ( .A(n9490), .B(n9489), .Z(n9561) );
  XOR U9719 ( .A(n73), .B(n9561), .Z(n9562) );
  XOR U9720 ( .A(n9563), .B(n9562), .Z(n9528) );
  NANDN U9721 ( .A(n9492), .B(n9491), .Z(n9496) );
  NAND U9722 ( .A(n9494), .B(n9493), .Z(n9495) );
  AND U9723 ( .A(n9496), .B(n9495), .Z(n9527) );
  XNOR U9724 ( .A(n9528), .B(n9527), .Z(n9529) );
  XOR U9725 ( .A(n75), .B(a[115]), .Z(n9543) );
  OR U9726 ( .A(n9543), .B(n10106), .Z(n9499) );
  NAND U9727 ( .A(n10107), .B(n9497), .Z(n9498) );
  NAND U9728 ( .A(n9499), .B(n9498), .Z(n9535) );
  ANDN U9729 ( .B(a[113]), .A(n75), .Z(n9604) );
  IV U9730 ( .A(n9604), .Z(n9706) );
  NANDN U9731 ( .A(n9500), .B(n10070), .Z(n9502) );
  XNOR U9732 ( .A(b[13]), .B(n9631), .Z(n9558) );
  NANDN U9733 ( .A(n10051), .B(n9558), .Z(n9501) );
  NAND U9734 ( .A(n9502), .B(n9501), .Z(n9533) );
  XOR U9735 ( .A(n9706), .B(n9533), .Z(n9534) );
  XOR U9736 ( .A(n9529), .B(n9530), .Z(n9521) );
  XOR U9737 ( .A(n9522), .B(n9521), .Z(n9524) );
  XOR U9738 ( .A(n9523), .B(n9524), .Z(n9574) );
  NANDN U9739 ( .A(n9504), .B(n9503), .Z(n9508) );
  NAND U9740 ( .A(n9506), .B(n9505), .Z(n9507) );
  NAND U9741 ( .A(n9508), .B(n9507), .Z(n9572) );
  OR U9742 ( .A(n9510), .B(n9509), .Z(n9514) );
  NANDN U9743 ( .A(n9512), .B(n9511), .Z(n9513) );
  AND U9744 ( .A(n9514), .B(n9513), .Z(n9573) );
  XNOR U9745 ( .A(n9572), .B(n9573), .Z(n9575) );
  XOR U9746 ( .A(n9574), .B(n9575), .Z(n9578) );
  XOR U9747 ( .A(n9579), .B(n9578), .Z(n9580) );
  XOR U9748 ( .A(n9581), .B(n9580), .Z(n9585) );
  XOR U9749 ( .A(n9586), .B(n9585), .Z(c[241]) );
  NANDN U9750 ( .A(n9516), .B(n9515), .Z(n9520) );
  OR U9751 ( .A(n9518), .B(n9517), .Z(n9519) );
  NAND U9752 ( .A(n9520), .B(n9519), .Z(n9589) );
  NAND U9753 ( .A(n9522), .B(n9521), .Z(n9526) );
  NAND U9754 ( .A(n9524), .B(n9523), .Z(n9525) );
  AND U9755 ( .A(n9526), .B(n9525), .Z(n9590) );
  XNOR U9756 ( .A(n9589), .B(n9590), .Z(n9591) );
  NANDN U9757 ( .A(n9528), .B(n9527), .Z(n9532) );
  NAND U9758 ( .A(n9530), .B(n9529), .Z(n9531) );
  NAND U9759 ( .A(n9532), .B(n9531), .Z(n9644) );
  NANDN U9760 ( .A(n9533), .B(n9604), .Z(n9537) );
  NANDN U9761 ( .A(n9535), .B(n9534), .Z(n9536) );
  AND U9762 ( .A(n9537), .B(n9536), .Z(n9645) );
  XNOR U9763 ( .A(n9644), .B(n9645), .Z(n9646) );
  NAND U9764 ( .A(a[114]), .B(b[15]), .Z(n9607) );
  NAND U9765 ( .A(b[1]), .B(b[2]), .Z(n9630) );
  XNOR U9766 ( .A(b[3]), .B(n9630), .Z(n9541) );
  XNOR U9767 ( .A(b[2]), .B(b[1]), .Z(n9538) );
  NANDN U9768 ( .A(n9539), .B(n9538), .Z(n9540) );
  AND U9769 ( .A(n9541), .B(n9540), .Z(n9605) );
  XOR U9770 ( .A(n9706), .B(n9605), .Z(n9606) );
  XNOR U9771 ( .A(n9607), .B(n9606), .Z(n9613) );
  XNOR U9772 ( .A(n75), .B(n9542), .Z(n9632) );
  OR U9773 ( .A(n9632), .B(n10106), .Z(n9545) );
  NANDN U9774 ( .A(n9543), .B(n10107), .Z(n9544) );
  NAND U9775 ( .A(n9545), .B(n9544), .Z(n9610) );
  XNOR U9776 ( .A(n9967), .B(n9815), .Z(n9627) );
  OR U9777 ( .A(n9627), .B(n10020), .Z(n9548) );
  NANDN U9778 ( .A(n9546), .B(n9968), .Z(n9547) );
  AND U9779 ( .A(n9548), .B(n9547), .Z(n9611) );
  XNOR U9780 ( .A(n9610), .B(n9611), .Z(n9612) );
  XOR U9781 ( .A(n9613), .B(n9612), .Z(n9618) );
  XNOR U9782 ( .A(n9984), .B(n10023), .Z(n9638) );
  NANDN U9783 ( .A(n9638), .B(n9865), .Z(n9551) );
  NANDN U9784 ( .A(n9549), .B(n9930), .Z(n9550) );
  NAND U9785 ( .A(n9551), .B(n9550), .Z(n9601) );
  XNOR U9786 ( .A(n9920), .B(n9872), .Z(n9641) );
  NANDN U9787 ( .A(n9641), .B(n9746), .Z(n9554) );
  NANDN U9788 ( .A(n9552), .B(n9747), .Z(n9553) );
  NAND U9789 ( .A(n9554), .B(n9553), .Z(n9598) );
  IV U9790 ( .A(a[126]), .Z(n10074) );
  XNOR U9791 ( .A(n10074), .B(n9622), .Z(n9624) );
  OR U9792 ( .A(n9624), .B(n9623), .Z(n9557) );
  NAND U9793 ( .A(n9555), .B(n9680), .Z(n9556) );
  AND U9794 ( .A(n9557), .B(n9556), .Z(n9599) );
  XNOR U9795 ( .A(n9598), .B(n9599), .Z(n9600) );
  XNOR U9796 ( .A(n9601), .B(n9600), .Z(n9616) );
  NAND U9797 ( .A(n10070), .B(n9558), .Z(n9560) );
  XOR U9798 ( .A(b[13]), .B(a[118]), .Z(n9635) );
  NANDN U9799 ( .A(n10051), .B(n9635), .Z(n9559) );
  NAND U9800 ( .A(n9560), .B(n9559), .Z(n9617) );
  XOR U9801 ( .A(n9616), .B(n9617), .Z(n9619) );
  XOR U9802 ( .A(n9618), .B(n9619), .Z(n9652) );
  NANDN U9803 ( .A(n9561), .B(b[1]), .Z(n9565) );
  NANDN U9804 ( .A(n9563), .B(n9562), .Z(n9564) );
  AND U9805 ( .A(n9565), .B(n9564), .Z(n9650) );
  NANDN U9806 ( .A(n9567), .B(n9566), .Z(n9571) );
  NAND U9807 ( .A(n9569), .B(n9568), .Z(n9570) );
  NAND U9808 ( .A(n9571), .B(n9570), .Z(n9651) );
  XNOR U9809 ( .A(n9650), .B(n9651), .Z(n9653) );
  XNOR U9810 ( .A(n9646), .B(n9647), .Z(n9592) );
  XOR U9811 ( .A(n9591), .B(n9592), .Z(n9596) );
  NANDN U9812 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U9813 ( .A(n9575), .B(n9574), .Z(n9576) );
  AND U9814 ( .A(n9577), .B(n9576), .Z(n9595) );
  NAND U9815 ( .A(n9579), .B(n9578), .Z(n9583) );
  NAND U9816 ( .A(n9581), .B(n9580), .Z(n9582) );
  NAND U9817 ( .A(n9583), .B(n9582), .Z(n9597) );
  XOR U9818 ( .A(n9595), .B(n9597), .Z(n9584) );
  XOR U9819 ( .A(n9596), .B(n9584), .Z(n9587) );
  OR U9820 ( .A(n9586), .B(n9585), .Z(n9588) );
  XNOR U9821 ( .A(n9587), .B(n9588), .Z(c[242]) );
  NANDN U9822 ( .A(n9588), .B(n9587), .Z(n9658) );
  NANDN U9823 ( .A(n9590), .B(n9589), .Z(n9594) );
  NAND U9824 ( .A(n9592), .B(n9591), .Z(n9593) );
  AND U9825 ( .A(n9594), .B(n9593), .Z(n9659) );
  NANDN U9826 ( .A(n9599), .B(n9598), .Z(n9603) );
  NAND U9827 ( .A(n9601), .B(n9600), .Z(n9602) );
  NAND U9828 ( .A(n9603), .B(n9602), .Z(n9715) );
  NANDN U9829 ( .A(n9605), .B(n9604), .Z(n9609) );
  NAND U9830 ( .A(n9607), .B(n9606), .Z(n9608) );
  NAND U9831 ( .A(n9609), .B(n9608), .Z(n9712) );
  NANDN U9832 ( .A(n9611), .B(n9610), .Z(n9615) );
  NAND U9833 ( .A(n9613), .B(n9612), .Z(n9614) );
  NAND U9834 ( .A(n9615), .B(n9614), .Z(n9713) );
  XNOR U9835 ( .A(n9712), .B(n9713), .Z(n9714) );
  XOR U9836 ( .A(n9715), .B(n9714), .Z(n9662) );
  NANDN U9837 ( .A(n9617), .B(n9616), .Z(n9621) );
  OR U9838 ( .A(n9619), .B(n9618), .Z(n9620) );
  NAND U9839 ( .A(n9621), .B(n9620), .Z(n9663) );
  XNOR U9840 ( .A(n9662), .B(n9663), .Z(n9664) );
  XNOR U9841 ( .A(n10049), .B(n9622), .Z(n9681) );
  OR U9842 ( .A(n9681), .B(n9623), .Z(n9626) );
  NANDN U9843 ( .A(n9624), .B(n9680), .Z(n9625) );
  NAND U9844 ( .A(n9626), .B(n9625), .Z(n9700) );
  XOR U9845 ( .A(n9967), .B(a[121]), .Z(n9668) );
  OR U9846 ( .A(n9668), .B(n10020), .Z(n9629) );
  NANDN U9847 ( .A(n9627), .B(n9968), .Z(n9628) );
  AND U9848 ( .A(n9629), .B(n9628), .Z(n9701) );
  XNOR U9849 ( .A(n9700), .B(n9701), .Z(n9702) );
  NAND U9850 ( .A(b[15]), .B(a[115]), .Z(n9709) );
  ANDN U9851 ( .B(n9630), .A(n74), .Z(n9707) );
  XNOR U9852 ( .A(n9706), .B(n9707), .Z(n9708) );
  XOR U9853 ( .A(n9709), .B(n9708), .Z(n9703) );
  XOR U9854 ( .A(n9702), .B(n9703), .Z(n9690) );
  XNOR U9855 ( .A(b[15]), .B(n9631), .Z(n9685) );
  NANDN U9856 ( .A(n10106), .B(n9685), .Z(n9634) );
  NANDN U9857 ( .A(n9632), .B(n10107), .Z(n9633) );
  NAND U9858 ( .A(n9634), .B(n9633), .Z(n9688) );
  XNOR U9859 ( .A(b[13]), .B(n9755), .Z(n9677) );
  NANDN U9860 ( .A(n10051), .B(n9677), .Z(n9637) );
  NAND U9861 ( .A(n9635), .B(n10070), .Z(n9636) );
  NAND U9862 ( .A(n9637), .B(n9636), .Z(n9697) );
  XOR U9863 ( .A(n9984), .B(a[123]), .Z(n9671) );
  NANDN U9864 ( .A(n9671), .B(n9865), .Z(n9640) );
  NANDN U9865 ( .A(n9638), .B(n9930), .Z(n9639) );
  NAND U9866 ( .A(n9640), .B(n9639), .Z(n9694) );
  XNOR U9867 ( .A(n9978), .B(n9872), .Z(n9674) );
  NANDN U9868 ( .A(n9674), .B(n9746), .Z(n9643) );
  NANDN U9869 ( .A(n9641), .B(n9747), .Z(n9642) );
  AND U9870 ( .A(n9643), .B(n9642), .Z(n9695) );
  XNOR U9871 ( .A(n9694), .B(n9695), .Z(n9696) );
  XNOR U9872 ( .A(n9697), .B(n9696), .Z(n9689) );
  XNOR U9873 ( .A(n9688), .B(n9689), .Z(n9691) );
  XOR U9874 ( .A(n9690), .B(n9691), .Z(n9665) );
  XOR U9875 ( .A(n9664), .B(n9665), .Z(n9720) );
  NANDN U9876 ( .A(n9645), .B(n9644), .Z(n9649) );
  NANDN U9877 ( .A(n9647), .B(n9646), .Z(n9648) );
  NAND U9878 ( .A(n9649), .B(n9648), .Z(n9718) );
  OR U9879 ( .A(n9651), .B(n9650), .Z(n9655) );
  NANDN U9880 ( .A(n9653), .B(n9652), .Z(n9654) );
  AND U9881 ( .A(n9655), .B(n9654), .Z(n9719) );
  XNOR U9882 ( .A(n9718), .B(n9719), .Z(n9721) );
  XOR U9883 ( .A(n9720), .B(n9721), .Z(n9660) );
  XOR U9884 ( .A(n9661), .B(n9660), .Z(n9656) );
  XOR U9885 ( .A(n9659), .B(n9656), .Z(n9657) );
  XNOR U9886 ( .A(n9658), .B(n9657), .Z(c[243]) );
  NANDN U9887 ( .A(n9658), .B(n9657), .Z(n9723) );
  NANDN U9888 ( .A(n9663), .B(n9662), .Z(n9667) );
  NAND U9889 ( .A(n9665), .B(n9664), .Z(n9666) );
  NAND U9890 ( .A(n9667), .B(n9666), .Z(n9733) );
  XNOR U9891 ( .A(n9967), .B(n10023), .Z(n9751) );
  OR U9892 ( .A(n9751), .B(n10020), .Z(n9670) );
  NANDN U9893 ( .A(n9668), .B(n9968), .Z(n9669) );
  NAND U9894 ( .A(n9670), .B(n9669), .Z(n9743) );
  XNOR U9895 ( .A(n9920), .B(n9984), .Z(n9759) );
  NANDN U9896 ( .A(n9759), .B(n9865), .Z(n9673) );
  NANDN U9897 ( .A(n9671), .B(n9930), .Z(n9672) );
  NAND U9898 ( .A(n9673), .B(n9672), .Z(n9740) );
  XNOR U9899 ( .A(n10074), .B(n9872), .Z(n9748) );
  NANDN U9900 ( .A(n9748), .B(n9746), .Z(n9676) );
  NANDN U9901 ( .A(n9674), .B(n9747), .Z(n9675) );
  AND U9902 ( .A(n9676), .B(n9675), .Z(n9741) );
  XNOR U9903 ( .A(n9740), .B(n9741), .Z(n9742) );
  XNOR U9904 ( .A(n9743), .B(n9742), .Z(n9737) );
  NAND U9905 ( .A(n10070), .B(n9677), .Z(n9679) );
  XOR U9906 ( .A(b[13]), .B(a[120]), .Z(n9762) );
  NANDN U9907 ( .A(n10051), .B(n9762), .Z(n9678) );
  NAND U9908 ( .A(n9679), .B(n9678), .Z(n9734) );
  NANDN U9909 ( .A(n9681), .B(n9680), .Z(n9682) );
  NANDN U9910 ( .A(n9683), .B(n9682), .Z(n9765) );
  ANDN U9911 ( .B(a[116]), .A(n75), .Z(n9792) );
  XOR U9912 ( .A(n9765), .B(n9792), .Z(n9766) );
  XNOR U9913 ( .A(n75), .B(n9684), .Z(n9756) );
  OR U9914 ( .A(n9756), .B(n10106), .Z(n9687) );
  NAND U9915 ( .A(n10107), .B(n9685), .Z(n9686) );
  AND U9916 ( .A(n9687), .B(n9686), .Z(n9767) );
  XOR U9917 ( .A(n9766), .B(n9767), .Z(n9735) );
  XOR U9918 ( .A(n9734), .B(n9735), .Z(n9736) );
  XOR U9919 ( .A(n9737), .B(n9736), .Z(n9776) );
  NANDN U9920 ( .A(n9689), .B(n9688), .Z(n9693) );
  NAND U9921 ( .A(n9691), .B(n9690), .Z(n9692) );
  NAND U9922 ( .A(n9693), .B(n9692), .Z(n9774) );
  NANDN U9923 ( .A(n9695), .B(n9694), .Z(n9699) );
  NAND U9924 ( .A(n9697), .B(n9696), .Z(n9698) );
  NAND U9925 ( .A(n9699), .B(n9698), .Z(n9771) );
  NANDN U9926 ( .A(n9701), .B(n9700), .Z(n9705) );
  NAND U9927 ( .A(n9703), .B(n9702), .Z(n9704) );
  NAND U9928 ( .A(n9705), .B(n9704), .Z(n9769) );
  OR U9929 ( .A(n9707), .B(n9706), .Z(n9711) );
  OR U9930 ( .A(n9709), .B(n9708), .Z(n9710) );
  AND U9931 ( .A(n9711), .B(n9710), .Z(n9768) );
  XNOR U9932 ( .A(n9769), .B(n9768), .Z(n9770) );
  XOR U9933 ( .A(n9771), .B(n9770), .Z(n9775) );
  XOR U9934 ( .A(n9774), .B(n9775), .Z(n9777) );
  XOR U9935 ( .A(n9776), .B(n9777), .Z(n9730) );
  NANDN U9936 ( .A(n9713), .B(n9712), .Z(n9717) );
  NANDN U9937 ( .A(n9715), .B(n9714), .Z(n9716) );
  NAND U9938 ( .A(n9717), .B(n9716), .Z(n9731) );
  XOR U9939 ( .A(n9730), .B(n9731), .Z(n9732) );
  XNOR U9940 ( .A(n9733), .B(n9732), .Z(n9724) );
  XOR U9941 ( .A(n9724), .B(n9725), .Z(n9727) );
  XOR U9942 ( .A(n9726), .B(n9727), .Z(n9722) );
  XOR U9943 ( .A(n9723), .B(n9722), .Z(c[244]) );
  OR U9944 ( .A(n9723), .B(n9722), .Z(n9838) );
  NANDN U9945 ( .A(n9725), .B(n9724), .Z(n9729) );
  OR U9946 ( .A(n9727), .B(n9726), .Z(n9728) );
  NAND U9947 ( .A(n9729), .B(n9728), .Z(n9834) );
  OR U9948 ( .A(n9735), .B(n9734), .Z(n9739) );
  NAND U9949 ( .A(n9737), .B(n9736), .Z(n9738) );
  NAND U9950 ( .A(n9739), .B(n9738), .Z(n9783) );
  NANDN U9951 ( .A(n9741), .B(n9740), .Z(n9745) );
  NAND U9952 ( .A(n9743), .B(n9742), .Z(n9744) );
  NAND U9953 ( .A(n9745), .B(n9744), .Z(n9789) );
  XNOR U9954 ( .A(n10049), .B(n9872), .Z(n9811) );
  NANDN U9955 ( .A(n9811), .B(n9746), .Z(n9750) );
  NANDN U9956 ( .A(n9748), .B(n9747), .Z(n9749) );
  NAND U9957 ( .A(n9750), .B(n9749), .Z(n9819) );
  XOR U9958 ( .A(n9967), .B(a[123]), .Z(n9805) );
  OR U9959 ( .A(n9805), .B(n10020), .Z(n9753) );
  NANDN U9960 ( .A(n9751), .B(n9968), .Z(n9752) );
  AND U9961 ( .A(n9753), .B(n9752), .Z(n9820) );
  XNOR U9962 ( .A(n9819), .B(n9820), .Z(n9821) );
  NAND U9963 ( .A(b[3]), .B(b[4]), .Z(n9754) );
  NAND U9964 ( .A(b[5]), .B(n9754), .Z(n9791) );
  AND U9965 ( .A(b[15]), .B(a[117]), .Z(n9790) );
  XNOR U9966 ( .A(n9791), .B(n9790), .Z(n9793) );
  XOR U9967 ( .A(n9792), .B(n9793), .Z(n9822) );
  XOR U9968 ( .A(n9821), .B(n9822), .Z(n9786) );
  XNOR U9969 ( .A(b[15]), .B(n9755), .Z(n9816) );
  NANDN U9970 ( .A(n10106), .B(n9816), .Z(n9758) );
  NANDN U9971 ( .A(n9756), .B(n10107), .Z(n9757) );
  NAND U9972 ( .A(n9758), .B(n9757), .Z(n9799) );
  XNOR U9973 ( .A(n9978), .B(n9984), .Z(n9808) );
  NANDN U9974 ( .A(n9808), .B(n9865), .Z(n9761) );
  NANDN U9975 ( .A(n9759), .B(n9930), .Z(n9760) );
  NAND U9976 ( .A(n9761), .B(n9760), .Z(n9796) );
  XOR U9977 ( .A(n10050), .B(a[121]), .Z(n9802) );
  OR U9978 ( .A(n9802), .B(n10051), .Z(n9764) );
  NAND U9979 ( .A(n9762), .B(n10070), .Z(n9763) );
  AND U9980 ( .A(n9764), .B(n9763), .Z(n9797) );
  XNOR U9981 ( .A(n9796), .B(n9797), .Z(n9798) );
  XOR U9982 ( .A(n9799), .B(n9798), .Z(n9787) );
  XNOR U9983 ( .A(n9786), .B(n9787), .Z(n9788) );
  XNOR U9984 ( .A(n9789), .B(n9788), .Z(n9780) );
  XNOR U9985 ( .A(n9780), .B(n9781), .Z(n9782) );
  XNOR U9986 ( .A(n9783), .B(n9782), .Z(n9828) );
  NANDN U9987 ( .A(n9769), .B(n9768), .Z(n9773) );
  NANDN U9988 ( .A(n9771), .B(n9770), .Z(n9772) );
  NAND U9989 ( .A(n9773), .B(n9772), .Z(n9825) );
  OR U9990 ( .A(n9775), .B(n9774), .Z(n9779) );
  NAND U9991 ( .A(n9777), .B(n9776), .Z(n9778) );
  AND U9992 ( .A(n9779), .B(n9778), .Z(n9826) );
  XNOR U9993 ( .A(n9825), .B(n9826), .Z(n9827) );
  XOR U9994 ( .A(n9828), .B(n9827), .Z(n9832) );
  XOR U9995 ( .A(n9831), .B(n9832), .Z(n9833) );
  XOR U9996 ( .A(n9834), .B(n9833), .Z(n9837) );
  XOR U9997 ( .A(n9838), .B(n9837), .Z(c[245]) );
  NANDN U9998 ( .A(n9781), .B(n9780), .Z(n9785) );
  NAND U9999 ( .A(n9783), .B(n9782), .Z(n9784) );
  NAND U10000 ( .A(n9785), .B(n9784), .Z(n9844) );
  NAND U10001 ( .A(n9791), .B(n9790), .Z(n9795) );
  NANDN U10002 ( .A(n9793), .B(n9792), .Z(n9794) );
  NAND U10003 ( .A(n9795), .B(n9794), .Z(n9856) );
  NANDN U10004 ( .A(n9797), .B(n9796), .Z(n9801) );
  NAND U10005 ( .A(n9799), .B(n9798), .Z(n9800) );
  NAND U10006 ( .A(n9801), .B(n9800), .Z(n9850) );
  XNOR U10007 ( .A(n10050), .B(n10023), .Z(n9869) );
  OR U10008 ( .A(n9869), .B(n10051), .Z(n9804) );
  NANDN U10009 ( .A(n9802), .B(n10070), .Z(n9803) );
  NAND U10010 ( .A(n9804), .B(n9803), .Z(n9882) );
  XNOR U10011 ( .A(n9967), .B(n9920), .Z(n9862) );
  OR U10012 ( .A(n9862), .B(n10020), .Z(n9807) );
  NANDN U10013 ( .A(n9805), .B(n9968), .Z(n9806) );
  NAND U10014 ( .A(n9807), .B(n9806), .Z(n9879) );
  XNOR U10015 ( .A(n10074), .B(n9984), .Z(n9866) );
  NANDN U10016 ( .A(n9866), .B(n9865), .Z(n9810) );
  NANDN U10017 ( .A(n9808), .B(n9930), .Z(n9809) );
  AND U10018 ( .A(n9810), .B(n9809), .Z(n9880) );
  XNOR U10019 ( .A(n9879), .B(n9880), .Z(n9881) );
  XNOR U10020 ( .A(n9882), .B(n9881), .Z(n9847) );
  NAND U10021 ( .A(b[5]), .B(b[6]), .Z(n9873) );
  XNOR U10022 ( .A(b[7]), .B(n9873), .Z(n9814) );
  XNOR U10023 ( .A(b[6]), .B(b[5]), .Z(n9812) );
  NAND U10024 ( .A(n9812), .B(n9811), .Z(n9813) );
  AND U10025 ( .A(n9814), .B(n9813), .Z(n9874) );
  ANDN U10026 ( .B(a[118]), .A(n75), .Z(n9924) );
  XNOR U10027 ( .A(n9874), .B(n9924), .Z(n9875) );
  XNOR U10028 ( .A(n75), .B(n9815), .Z(n9859) );
  OR U10029 ( .A(n9859), .B(n10106), .Z(n9818) );
  NAND U10030 ( .A(n10107), .B(n9816), .Z(n9817) );
  AND U10031 ( .A(n9818), .B(n9817), .Z(n9876) );
  XNOR U10032 ( .A(n9875), .B(n9876), .Z(n9848) );
  XNOR U10033 ( .A(n9847), .B(n9848), .Z(n9849) );
  XOR U10034 ( .A(n9850), .B(n9849), .Z(n9853) );
  NANDN U10035 ( .A(n9820), .B(n9819), .Z(n9824) );
  NANDN U10036 ( .A(n9822), .B(n9821), .Z(n9823) );
  AND U10037 ( .A(n9824), .B(n9823), .Z(n9854) );
  XNOR U10038 ( .A(n9853), .B(n9854), .Z(n9855) );
  XNOR U10039 ( .A(n9856), .B(n9855), .Z(n9842) );
  XNOR U10040 ( .A(n9841), .B(n9842), .Z(n9843) );
  XNOR U10041 ( .A(n9844), .B(n9843), .Z(n9885) );
  NANDN U10042 ( .A(n9826), .B(n9825), .Z(n9830) );
  NANDN U10043 ( .A(n9828), .B(n9827), .Z(n9829) );
  AND U10044 ( .A(n9830), .B(n9829), .Z(n9886) );
  XNOR U10045 ( .A(n9885), .B(n9886), .Z(n9888) );
  OR U10046 ( .A(n9832), .B(n9831), .Z(n9836) );
  NAND U10047 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10048 ( .A(n9836), .B(n9835), .Z(n9887) );
  XNOR U10049 ( .A(n9888), .B(n9887), .Z(n9839) );
  OR U10050 ( .A(n9838), .B(n9837), .Z(n9840) );
  XNOR U10051 ( .A(n9839), .B(n9840), .Z(c[246]) );
  NANDN U10052 ( .A(n9840), .B(n9839), .Z(n9945) );
  NANDN U10053 ( .A(n9842), .B(n9841), .Z(n9846) );
  NANDN U10054 ( .A(n9844), .B(n9843), .Z(n9845) );
  NAND U10055 ( .A(n9846), .B(n9845), .Z(n9899) );
  NANDN U10056 ( .A(n9848), .B(n9847), .Z(n9852) );
  NANDN U10057 ( .A(n9850), .B(n9849), .Z(n9851) );
  AND U10058 ( .A(n9852), .B(n9851), .Z(n9892) );
  NANDN U10059 ( .A(n9854), .B(n9853), .Z(n9858) );
  NAND U10060 ( .A(n9856), .B(n9855), .Z(n9857) );
  NAND U10061 ( .A(n9858), .B(n9857), .Z(n9893) );
  XNOR U10062 ( .A(n9892), .B(n9893), .Z(n9895) );
  XOR U10063 ( .A(n75), .B(a[121]), .Z(n9934) );
  OR U10064 ( .A(n9934), .B(n10106), .Z(n9861) );
  NANDN U10065 ( .A(n9859), .B(n10107), .Z(n9860) );
  NAND U10066 ( .A(n9861), .B(n9860), .Z(n9940) );
  XNOR U10067 ( .A(n9967), .B(n9978), .Z(n9917) );
  OR U10068 ( .A(n9917), .B(n10020), .Z(n9864) );
  NANDN U10069 ( .A(n9862), .B(n9968), .Z(n9863) );
  NAND U10070 ( .A(n9864), .B(n9863), .Z(n9938) );
  XNOR U10071 ( .A(n10049), .B(n9984), .Z(n9931) );
  NANDN U10072 ( .A(n9931), .B(n9865), .Z(n9868) );
  NANDN U10073 ( .A(n9866), .B(n9930), .Z(n9867) );
  NAND U10074 ( .A(n9868), .B(n9867), .Z(n9911) );
  XOR U10075 ( .A(b[13]), .B(a[123]), .Z(n9921) );
  NANDN U10076 ( .A(n10051), .B(n9921), .Z(n9871) );
  NANDN U10077 ( .A(n9869), .B(n10070), .Z(n9870) );
  AND U10078 ( .A(n9871), .B(n9870), .Z(n9912) );
  XNOR U10079 ( .A(n9911), .B(n9912), .Z(n9913) );
  ANDN U10080 ( .B(n9873), .A(n9872), .Z(n9925) );
  XOR U10081 ( .A(n9925), .B(n9924), .Z(n9927) );
  NAND U10082 ( .A(a[119]), .B(b[15]), .Z(n9926) );
  XOR U10083 ( .A(n9927), .B(n9926), .Z(n9914) );
  XOR U10084 ( .A(n9913), .B(n9914), .Z(n9937) );
  XOR U10085 ( .A(n9938), .B(n9937), .Z(n9939) );
  XNOR U10086 ( .A(n9940), .B(n9939), .Z(n9908) );
  NANDN U10087 ( .A(n9874), .B(n9924), .Z(n9878) );
  NAND U10088 ( .A(n9876), .B(n9875), .Z(n9877) );
  NAND U10089 ( .A(n9878), .B(n9877), .Z(n9905) );
  NANDN U10090 ( .A(n9880), .B(n9879), .Z(n9884) );
  NAND U10091 ( .A(n9882), .B(n9881), .Z(n9883) );
  NAND U10092 ( .A(n9884), .B(n9883), .Z(n9906) );
  XNOR U10093 ( .A(n9905), .B(n9906), .Z(n9907) );
  XOR U10094 ( .A(n9908), .B(n9907), .Z(n9894) );
  IV U10095 ( .A(n9900), .Z(n9898) );
  NAND U10096 ( .A(n9886), .B(n9885), .Z(n9890) );
  NANDN U10097 ( .A(n9888), .B(n9887), .Z(n9889) );
  NAND U10098 ( .A(n9890), .B(n9889), .Z(n9901) );
  XNOR U10099 ( .A(n9898), .B(n9901), .Z(n9891) );
  XNOR U10100 ( .A(n9899), .B(n9891), .Z(n9944) );
  XNOR U10101 ( .A(n9945), .B(n9944), .Z(c[247]) );
  OR U10102 ( .A(n9893), .B(n9892), .Z(n9897) );
  NANDN U10103 ( .A(n9895), .B(n9894), .Z(n9896) );
  NAND U10104 ( .A(n9897), .B(n9896), .Z(n9948) );
  NAND U10105 ( .A(n9898), .B(n9899), .Z(n9904) );
  ANDN U10106 ( .B(n9900), .A(n9899), .Z(n9902) );
  NANDN U10107 ( .A(n9902), .B(n9901), .Z(n9903) );
  AND U10108 ( .A(n9904), .B(n9903), .Z(n9946) );
  NANDN U10109 ( .A(n9906), .B(n9905), .Z(n9910) );
  NAND U10110 ( .A(n9908), .B(n9907), .Z(n9909) );
  NAND U10111 ( .A(n9910), .B(n9909), .Z(n9952) );
  NANDN U10112 ( .A(n9912), .B(n9911), .Z(n9916) );
  NAND U10113 ( .A(n9914), .B(n9913), .Z(n9915) );
  NAND U10114 ( .A(n9916), .B(n9915), .Z(n9962) );
  XOR U10115 ( .A(a[126]), .B(b[11]), .Z(n9969) );
  NANDN U10116 ( .A(n10020), .B(n9969), .Z(n9919) );
  NANDN U10117 ( .A(n9917), .B(n9968), .Z(n9918) );
  AND U10118 ( .A(n9919), .B(n9918), .Z(n9955) );
  XNOR U10119 ( .A(b[13]), .B(n9920), .Z(n9977) );
  NANDN U10120 ( .A(n10051), .B(n9977), .Z(n9923) );
  NAND U10121 ( .A(n9921), .B(n10070), .Z(n9922) );
  AND U10122 ( .A(n9923), .B(n9922), .Z(n9956) );
  XNOR U10123 ( .A(n9955), .B(n9956), .Z(n9957) );
  NANDN U10124 ( .A(n9925), .B(n9924), .Z(n9929) );
  OR U10125 ( .A(n9927), .B(n9926), .Z(n9928) );
  AND U10126 ( .A(n9929), .B(n9928), .Z(n9958) );
  XOR U10127 ( .A(n9957), .B(n9958), .Z(n9961) );
  XNOR U10128 ( .A(n9962), .B(n9961), .Z(n9964) );
  NANDN U10129 ( .A(n9931), .B(n9930), .Z(n9933) );
  ANDN U10130 ( .B(n9933), .A(n9932), .Z(n9974) );
  ANDN U10131 ( .B(a[120]), .A(n75), .Z(n10014) );
  XNOR U10132 ( .A(b[15]), .B(n10023), .Z(n9981) );
  NANDN U10133 ( .A(n10106), .B(n9981), .Z(n9936) );
  NANDN U10134 ( .A(n9934), .B(n10107), .Z(n9935) );
  AND U10135 ( .A(n9936), .B(n9935), .Z(n9972) );
  XOR U10136 ( .A(n10014), .B(n9972), .Z(n9973) );
  XNOR U10137 ( .A(n9974), .B(n9973), .Z(n9963) );
  XOR U10138 ( .A(n9964), .B(n9963), .Z(n9949) );
  NAND U10139 ( .A(n9938), .B(n9937), .Z(n9942) );
  NAND U10140 ( .A(n9940), .B(n9939), .Z(n9941) );
  NAND U10141 ( .A(n9942), .B(n9941), .Z(n9950) );
  XNOR U10142 ( .A(n9949), .B(n9950), .Z(n9951) );
  XNOR U10143 ( .A(n9952), .B(n9951), .Z(n9947) );
  XOR U10144 ( .A(n9946), .B(n9947), .Z(n9943) );
  XOR U10145 ( .A(n9948), .B(n9943), .Z(n9986) );
  NANDN U10146 ( .A(n9945), .B(n9944), .Z(n9987) );
  XNOR U10147 ( .A(n9986), .B(n9987), .Z(c[248]) );
  NANDN U10148 ( .A(n9950), .B(n9949), .Z(n9954) );
  NAND U10149 ( .A(n9952), .B(n9951), .Z(n9953) );
  NAND U10150 ( .A(n9954), .B(n9953), .Z(n9991) );
  OR U10151 ( .A(n9956), .B(n9955), .Z(n9960) );
  OR U10152 ( .A(n9958), .B(n9957), .Z(n9959) );
  NAND U10153 ( .A(n9960), .B(n9959), .Z(n9998) );
  NAND U10154 ( .A(n9962), .B(n9961), .Z(n9966) );
  NANDN U10155 ( .A(n9964), .B(n9963), .Z(n9965) );
  NAND U10156 ( .A(n9966), .B(n9965), .Z(n9997) );
  XNOR U10157 ( .A(n9967), .B(n10049), .Z(n10019) );
  OR U10158 ( .A(n10019), .B(n10020), .Z(n9971) );
  NAND U10159 ( .A(n9969), .B(n9968), .Z(n9970) );
  NAND U10160 ( .A(n9971), .B(n9970), .Z(n10002) );
  OR U10161 ( .A(n10014), .B(n9972), .Z(n9976) );
  NANDN U10162 ( .A(n9974), .B(n9973), .Z(n9975) );
  AND U10163 ( .A(n9976), .B(n9975), .Z(n10003) );
  XNOR U10164 ( .A(n10002), .B(n10003), .Z(n10004) );
  NAND U10165 ( .A(n10070), .B(n9977), .Z(n9980) );
  XNOR U10166 ( .A(b[13]), .B(n9978), .Z(n10027) );
  NANDN U10167 ( .A(n10051), .B(n10027), .Z(n9979) );
  AND U10168 ( .A(n9980), .B(n9979), .Z(n10008) );
  XOR U10169 ( .A(b[15]), .B(a[123]), .Z(n10024) );
  NANDN U10170 ( .A(n10106), .B(n10024), .Z(n9983) );
  NAND U10171 ( .A(n9981), .B(n10107), .Z(n9982) );
  AND U10172 ( .A(n9983), .B(n9982), .Z(n10009) );
  XOR U10173 ( .A(n10008), .B(n10009), .Z(n10010) );
  NAND U10174 ( .A(b[7]), .B(b[8]), .Z(n9985) );
  ANDN U10175 ( .B(n9985), .A(n9984), .Z(n10012) );
  NAND U10176 ( .A(b[15]), .B(a[121]), .Z(n10013) );
  XOR U10177 ( .A(n10012), .B(n10013), .Z(n10015) );
  XNOR U10178 ( .A(n10014), .B(n10015), .Z(n10011) );
  XOR U10179 ( .A(n10010), .B(n10011), .Z(n10005) );
  XNOR U10180 ( .A(n10004), .B(n10005), .Z(n9996) );
  XNOR U10181 ( .A(n9997), .B(n9996), .Z(n9999) );
  XNOR U10182 ( .A(n9998), .B(n9999), .Z(n9990) );
  XOR U10183 ( .A(n9991), .B(n9990), .Z(n9993) );
  XOR U10184 ( .A(n9992), .B(n9993), .Z(n9988) );
  NANDN U10185 ( .A(n9987), .B(n9986), .Z(n9989) );
  XNOR U10186 ( .A(n9988), .B(n9989), .Z(c[249]) );
  NANDN U10187 ( .A(n9989), .B(n9988), .Z(n10032) );
  NANDN U10188 ( .A(n9991), .B(n9990), .Z(n9995) );
  OR U10189 ( .A(n9993), .B(n9992), .Z(n9994) );
  AND U10190 ( .A(n9995), .B(n9994), .Z(n10035) );
  NAND U10191 ( .A(n9997), .B(n9996), .Z(n10001) );
  NANDN U10192 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U10193 ( .A(n10001), .B(n10000), .Z(n10033) );
  NANDN U10194 ( .A(n10003), .B(n10002), .Z(n10007) );
  NANDN U10195 ( .A(n10005), .B(n10004), .Z(n10006) );
  NAND U10196 ( .A(n10007), .B(n10006), .Z(n10055) );
  XNOR U10197 ( .A(n10055), .B(n10054), .Z(n10056) );
  OR U10198 ( .A(n10013), .B(n10012), .Z(n10017) );
  NAND U10199 ( .A(n10015), .B(n10014), .Z(n10016) );
  NAND U10200 ( .A(n10017), .B(n10016), .Z(n10036) );
  XNOR U10201 ( .A(b[11]), .B(n10018), .Z(n10022) );
  NAND U10202 ( .A(n10020), .B(n10019), .Z(n10021) );
  AND U10203 ( .A(n10022), .B(n10021), .Z(n10042) );
  NOR U10204 ( .A(n10023), .B(n75), .Z(n10080) );
  XOR U10205 ( .A(n10042), .B(n10080), .Z(n10043) );
  XNOR U10206 ( .A(b[15]), .B(a[124]), .Z(n10045) );
  OR U10207 ( .A(n10045), .B(n10106), .Z(n10026) );
  NAND U10208 ( .A(n10107), .B(n10024), .Z(n10025) );
  AND U10209 ( .A(n10026), .B(n10025), .Z(n10044) );
  XOR U10210 ( .A(n10043), .B(n10044), .Z(n10037) );
  XOR U10211 ( .A(n10036), .B(n10037), .Z(n10038) );
  NAND U10212 ( .A(n10070), .B(n10027), .Z(n10029) );
  XNOR U10213 ( .A(a[126]), .B(n10050), .Z(n10048) );
  NANDN U10214 ( .A(n10051), .B(n10048), .Z(n10028) );
  AND U10215 ( .A(n10029), .B(n10028), .Z(n10039) );
  XOR U10216 ( .A(n10038), .B(n10039), .Z(n10057) );
  XOR U10217 ( .A(n10056), .B(n10057), .Z(n10034) );
  XOR U10218 ( .A(n10033), .B(n10034), .Z(n10030) );
  XNOR U10219 ( .A(n10035), .B(n10030), .Z(n10031) );
  XOR U10220 ( .A(n10032), .B(n10031), .Z(c[250]) );
  OR U10221 ( .A(n10032), .B(n10031), .Z(n10091) );
  OR U10222 ( .A(n10037), .B(n10036), .Z(n10041) );
  NAND U10223 ( .A(n10039), .B(n10038), .Z(n10040) );
  NAND U10224 ( .A(n10041), .B(n10040), .Z(n10067) );
  NAND U10225 ( .A(b[15]), .B(a[123]), .Z(n10079) );
  XNOR U10226 ( .A(n10078), .B(n10079), .Z(n10081) );
  XNOR U10227 ( .A(b[15]), .B(a[125]), .Z(n10075) );
  OR U10228 ( .A(n10075), .B(n10106), .Z(n10047) );
  NANDN U10229 ( .A(n10045), .B(n10107), .Z(n10046) );
  NAND U10230 ( .A(n10047), .B(n10046), .Z(n10084) );
  XOR U10231 ( .A(n10085), .B(n10084), .Z(n10086) );
  NAND U10232 ( .A(n10070), .B(n10048), .Z(n10053) );
  XNOR U10233 ( .A(n10050), .B(n10049), .Z(n10071) );
  OR U10234 ( .A(n10071), .B(n10051), .Z(n10052) );
  AND U10235 ( .A(n10053), .B(n10052), .Z(n10087) );
  XNOR U10236 ( .A(n10086), .B(n10087), .Z(n10065) );
  XNOR U10237 ( .A(n10064), .B(n10065), .Z(n10066) );
  XNOR U10238 ( .A(n10067), .B(n10066), .Z(n10061) );
  NANDN U10239 ( .A(n10055), .B(n10054), .Z(n10059) );
  NAND U10240 ( .A(n10057), .B(n10056), .Z(n10058) );
  AND U10241 ( .A(n10059), .B(n10058), .Z(n10062) );
  XOR U10242 ( .A(n10061), .B(n10062), .Z(n10060) );
  XOR U10243 ( .A(n10063), .B(n10060), .Z(n10090) );
  XNOR U10244 ( .A(n10091), .B(n10090), .Z(c[251]) );
  NANDN U10245 ( .A(n10065), .B(n10064), .Z(n10069) );
  NAND U10246 ( .A(n10067), .B(n10066), .Z(n10068) );
  NAND U10247 ( .A(n10069), .B(n10068), .Z(n10095) );
  NANDN U10248 ( .A(n10071), .B(n10070), .Z(n10072) );
  NANDN U10249 ( .A(n10073), .B(n10072), .Z(n10101) );
  ANDN U10250 ( .B(a[124]), .A(n75), .Z(n10126) );
  XOR U10251 ( .A(n10101), .B(n10126), .Z(n10103) );
  XNOR U10252 ( .A(n10074), .B(n75), .Z(n10108) );
  OR U10253 ( .A(n10108), .B(n10106), .Z(n10077) );
  NANDN U10254 ( .A(n10075), .B(n10107), .Z(n10076) );
  NAND U10255 ( .A(n10077), .B(n10076), .Z(n10102) );
  XNOR U10256 ( .A(n10103), .B(n10102), .Z(n10111) );
  OR U10257 ( .A(n10079), .B(n10078), .Z(n10083) );
  NANDN U10258 ( .A(n10081), .B(n10080), .Z(n10082) );
  AND U10259 ( .A(n10083), .B(n10082), .Z(n10112) );
  XNOR U10260 ( .A(n10111), .B(n10112), .Z(n10113) );
  OR U10261 ( .A(n10085), .B(n10084), .Z(n10089) );
  NAND U10262 ( .A(n10087), .B(n10086), .Z(n10088) );
  AND U10263 ( .A(n10089), .B(n10088), .Z(n10114) );
  XOR U10264 ( .A(n10113), .B(n10114), .Z(n10094) );
  XOR U10265 ( .A(n10095), .B(n10094), .Z(n10097) );
  XNOR U10266 ( .A(n10096), .B(n10097), .Z(n10092) );
  NANDN U10267 ( .A(n10091), .B(n10090), .Z(n10093) );
  XNOR U10268 ( .A(n10092), .B(n10093), .Z(c[252]) );
  NANDN U10269 ( .A(n10093), .B(n10092), .Z(n10118) );
  NANDN U10270 ( .A(n10095), .B(n10094), .Z(n10099) );
  NANDN U10271 ( .A(n10097), .B(n10096), .Z(n10098) );
  NAND U10272 ( .A(n10099), .B(n10098), .Z(n10133) );
  NAND U10273 ( .A(b[11]), .B(b[12]), .Z(n10100) );
  NAND U10274 ( .A(b[13]), .B(n10100), .Z(n10125) );
  AND U10275 ( .A(b[15]), .B(a[125]), .Z(n10124) );
  XNOR U10276 ( .A(n10125), .B(n10124), .Z(n10127) );
  XOR U10277 ( .A(n10126), .B(n10127), .Z(n10139) );
  NANDN U10278 ( .A(n10101), .B(n10126), .Z(n10105) );
  OR U10279 ( .A(n10103), .B(n10102), .Z(n10104) );
  NAND U10280 ( .A(n10105), .B(n10104), .Z(n10137) );
  XOR U10281 ( .A(n75), .B(a[127]), .Z(n10120) );
  OR U10282 ( .A(n10120), .B(n10106), .Z(n10110) );
  NANDN U10283 ( .A(n10108), .B(n10107), .Z(n10109) );
  NAND U10284 ( .A(n10110), .B(n10109), .Z(n10136) );
  XNOR U10285 ( .A(n10137), .B(n10136), .Z(n10138) );
  XOR U10286 ( .A(n10139), .B(n10138), .Z(n10130) );
  NANDN U10287 ( .A(n10112), .B(n10111), .Z(n10116) );
  NAND U10288 ( .A(n10114), .B(n10113), .Z(n10115) );
  NAND U10289 ( .A(n10116), .B(n10115), .Z(n10131) );
  XNOR U10290 ( .A(n10130), .B(n10131), .Z(n10132) );
  XNOR U10291 ( .A(n10133), .B(n10132), .Z(n10117) );
  XOR U10292 ( .A(n10118), .B(n10117), .Z(c[253]) );
  OR U10293 ( .A(n10118), .B(n10117), .Z(n10153) );
  NAND U10294 ( .A(b[13]), .B(b[14]), .Z(n10119) );
  XNOR U10295 ( .A(b[15]), .B(n10119), .Z(n10123) );
  XNOR U10296 ( .A(b[14]), .B(b[13]), .Z(n10121) );
  NAND U10297 ( .A(n10121), .B(n10120), .Z(n10122) );
  AND U10298 ( .A(n10123), .B(n10122), .Z(n10160) );
  NAND U10299 ( .A(a[126]), .B(b[15]), .Z(n10159) );
  NAND U10300 ( .A(n10125), .B(n10124), .Z(n10129) );
  NANDN U10301 ( .A(n10127), .B(n10126), .Z(n10128) );
  AND U10302 ( .A(n10129), .B(n10128), .Z(n10158) );
  XNOR U10303 ( .A(n10159), .B(n10158), .Z(n10161) );
  XNOR U10304 ( .A(n10160), .B(n10161), .Z(n10148) );
  NANDN U10305 ( .A(n10131), .B(n10130), .Z(n10135) );
  NANDN U10306 ( .A(n10133), .B(n10132), .Z(n10134) );
  NAND U10307 ( .A(n10135), .B(n10134), .Z(n10146) );
  NANDN U10308 ( .A(n10137), .B(n10136), .Z(n10141) );
  NANDN U10309 ( .A(n10139), .B(n10138), .Z(n10140) );
  AND U10310 ( .A(n10141), .B(n10140), .Z(n10147) );
  XOR U10311 ( .A(n10146), .B(n10147), .Z(n10149) );
  XOR U10312 ( .A(n10148), .B(n10149), .Z(n10152) );
  XOR U10313 ( .A(n10153), .B(n10152), .Z(c[254]) );
  NAND U10314 ( .A(b[15]), .B(b[13]), .Z(n10144) );
  NAND U10315 ( .A(b[14]), .B(n10142), .Z(n10143) );
  NAND U10316 ( .A(n10144), .B(n10143), .Z(n10145) );
  AND U10317 ( .A(n10145), .B(a[127]), .Z(n10157) );
  AND U10318 ( .A(n10147), .B(n10146), .Z(n10151) );
  AND U10319 ( .A(n10149), .B(n10148), .Z(n10150) );
  OR U10320 ( .A(n10151), .B(n10150), .Z(n10155) );
  OR U10321 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U10322 ( .A(n10155), .B(n10154), .Z(n10156) );
  XNOR U10323 ( .A(n10157), .B(n10156), .Z(n10165) );
  NOR U10324 ( .A(n10159), .B(n10158), .Z(n10163) );
  NOR U10325 ( .A(n10161), .B(n10160), .Z(n10162) );
  NOR U10326 ( .A(n10163), .B(n10162), .Z(n10164) );
  XNOR U10327 ( .A(n10165), .B(n10164), .Z(c[255]) );
endmodule

