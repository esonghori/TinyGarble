
module hamming_N160_CC1 ( clk, rst, x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222;

  XNOR U162 ( .A(n131), .B(n295), .Z(n133) );
  XNOR U163 ( .A(n398), .B(n749), .Z(n404) );
  XNOR U164 ( .A(n517), .B(n519), .Z(n538) );
  XNOR U165 ( .A(n594), .B(n596), .Z(n615) );
  XNOR U166 ( .A(n675), .B(n677), .Z(n696) );
  XNOR U167 ( .A(n161), .B(n163), .Z(n175) );
  XNOR U168 ( .A(n227), .B(n228), .Z(n240) );
  XNOR U169 ( .A(n446), .B(n448), .Z(n467) );
  XNOR U170 ( .A(n215), .B(n216), .Z(n223) );
  ANDN U171 ( .B(n1201), .A(n1200), .Z(n769) );
  XNOR U172 ( .A(n269), .B(n270), .Z(n282) );
  XNOR U173 ( .A(n369), .B(n370), .Z(n382) );
  XNOR U174 ( .A(n317), .B(n318), .Z(n330) );
  XNOR U175 ( .A(n555), .B(n927), .Z(n536) );
  XNOR U176 ( .A(n632), .B(n1011), .Z(n613) );
  XNOR U177 ( .A(n713), .B(n1095), .Z(n694) );
  XNOR U178 ( .A(n257), .B(n258), .Z(n265) );
  XNOR U179 ( .A(n305), .B(n306), .Z(n313) );
  XNOR U180 ( .A(n357), .B(n358), .Z(n365) );
  XNOR U181 ( .A(n133), .B(n134), .Z(n146) );
  XNOR U182 ( .A(n186), .B(n187), .Z(n199) );
  XNOR U183 ( .A(n855), .B(n854), .Z(n874) );
  XNOR U184 ( .A(n836), .B(n835), .Z(n833) );
  XNOR U185 ( .A(n174), .B(n175), .Z(n182) );
  XNOR U186 ( .A(n72), .B(n73), .Z(n85) );
  XNOR U187 ( .A(n239), .B(n462), .Z(n222) );
  XNOR U188 ( .A(n89), .B(n91), .Z(n103) );
  XNOR U189 ( .A(n1086), .B(n1085), .Z(n1083) );
  XNOR U190 ( .A(n1128), .B(n1127), .Z(n1125) );
  XNOR U191 ( .A(n1044), .B(n1043), .Z(n1041) );
  XNOR U192 ( .A(n918), .B(n917), .Z(n915) );
  XNOR U193 ( .A(n275), .B(n552), .Z(n281) );
  XNOR U194 ( .A(n299), .B(n591), .Z(n305) );
  XNOR U195 ( .A(n788), .B(n792), .Z(n790) );
  XNOR U196 ( .A(n329), .B(n610), .Z(n312) );
  XNOR U197 ( .A(n115), .B(n259), .Z(n121) );
  XNOR U198 ( .A(n184), .B(n394), .Z(n186) );
  XNOR U199 ( .A(n694), .B(n696), .Z(n734) );
  XNOR U200 ( .A(n209), .B(n443), .Z(n215) );
  XNOR U201 ( .A(n233), .B(n481), .Z(n239) );
  XNOR U202 ( .A(n364), .B(n365), .Z(n388) );
  XOR U203 ( .A(n145), .B(n283), .Z(n127) );
  XNOR U204 ( .A(n70), .B(n164), .Z(n72) );
  XNOR U205 ( .A(n96), .B(n217), .Z(n102) );
  XNOR U206 ( .A(n182), .B(n154), .Z(n336) );
  ANDN U207 ( .B(n989), .A(n597), .Z(n599) );
  ANDN U208 ( .B(n1203), .A(n793), .Z(n795) );
  NANDN U209 ( .A(n1221), .B(n1222), .Z(n1217) );
  XNOR U210 ( .A(n1191), .B(n1190), .Z(n1210) );
  XNOR U211 ( .A(n1170), .B(n1169), .Z(n1167) );
  XNOR U212 ( .A(n979), .B(n978), .Z(n996) );
  XNOR U213 ( .A(n960), .B(n959), .Z(n957) );
  XNOR U214 ( .A(n375), .B(n710), .Z(n381) );
  XNOR U215 ( .A(n323), .B(n629), .Z(n329) );
  XNOR U216 ( .A(n251), .B(n514), .Z(n257) );
  XNOR U217 ( .A(n351), .B(n672), .Z(n357) );
  XNOR U218 ( .A(n416), .B(n417), .Z(n429) );
  XNOR U219 ( .A(n752), .B(n754), .Z(n773) );
  XNOR U220 ( .A(n281), .B(n533), .Z(n264) );
  XNOR U221 ( .A(n404), .B(n405), .Z(n412) );
  XNOR U222 ( .A(n139), .B(n307), .Z(n145) );
  XNOR U223 ( .A(n108), .B(n110), .Z(n122) );
  XNOR U224 ( .A(n168), .B(n359), .Z(n174) );
  XNOR U225 ( .A(n878), .B(n877), .Z(n875) );
  XNOR U226 ( .A(n815), .B(n814), .Z(n832) );
  XOR U227 ( .A(n613), .B(n969), .Z(n575) );
  XNOR U228 ( .A(n203), .B(n204), .Z(n216) );
  XNOR U229 ( .A(n199), .B(n179), .Z(n383) );
  XOR U230 ( .A(n49), .B(n123), .Z(n54) );
  XNOR U231 ( .A(n85), .B(n65), .Z(n152) );
  XNOR U232 ( .A(n35), .B(n92), .Z(n37) );
  XNOR U233 ( .A(n465), .B(n467), .Z(n652) );
  ANDN U234 ( .B(n1159), .A(n755), .Z(n757) );
  ANDN U235 ( .B(n1033), .A(n635), .Z(n637) );
  ANDN U236 ( .B(n907), .A(n520), .Z(n522) );
  ANDN U237 ( .B(n949), .A(n558), .Z(n560) );
  ANDN U238 ( .B(n1117), .A(n716), .Z(n718) );
  ANDN U239 ( .B(n1075), .A(n678), .Z(n680) );
  XNOR U240 ( .A(n1065), .B(n1064), .Z(n1082) );
  XNOR U241 ( .A(n1105), .B(n1104), .Z(n1124) );
  XNOR U242 ( .A(n1149), .B(n1148), .Z(n1166) );
  XNOR U243 ( .A(n1021), .B(n1020), .Z(n1040) );
  XNOR U244 ( .A(n1000), .B(n999), .Z(n997) );
  XNOR U245 ( .A(n897), .B(n896), .Z(n914) );
  XNOR U246 ( .A(n937), .B(n936), .Z(n956) );
  ANDN U247 ( .B(n867), .A(n487), .Z(n489) );
  ANDN U248 ( .B(n825), .A(n449), .Z(n451) );
  XNOR U249 ( .A(n245), .B(n246), .Z(n258) );
  XNOR U250 ( .A(n345), .B(n346), .Z(n358) );
  XOR U251 ( .A(n422), .B(n787), .Z(n427) );
  XNOR U252 ( .A(n381), .B(n691), .Z(n364) );
  XOR U253 ( .A(n192), .B(n406), .Z(n197) );
  XOR U254 ( .A(n312), .B(n571), .Z(n287) );
  XNOR U255 ( .A(n41), .B(n111), .Z(n43) );
  XOR U256 ( .A(n78), .B(n176), .Z(n83) );
  XNOR U257 ( .A(n484), .B(n845), .Z(n465) );
  XOR U258 ( .A(n26), .B(n62), .Z(n31) );
  XOR U259 ( .A(n13), .B(n45), .Z(n14) );
  XNOR U260 ( .A(n648), .B(n658), .Z(n887) );
  XNOR U261 ( .A(n222), .B(n223), .Z(n335) );
  XNOR U262 ( .A(n102), .B(n103), .Z(n151) );
  XNOR U263 ( .A(n37), .B(n38), .Z(n61) );
  XOR U264 ( .A(n1), .B(n2), .Z(o[7]) );
  XOR U265 ( .A(n3), .B(n4), .Z(n2) );
  XOR U266 ( .A(n5), .B(n6), .Z(n1) );
  AND U267 ( .A(o[6]), .B(n3), .Z(n6) );
  AND U268 ( .A(n7), .B(n8), .Z(n5) );
  XNOR U269 ( .A(n9), .B(n10), .Z(n8) );
  XNOR U270 ( .A(n7), .B(n11), .Z(o[6]) );
  XNOR U271 ( .A(n3), .B(n9), .Z(n11) );
  XNOR U272 ( .A(n12), .B(n13), .Z(n9) );
  AND U273 ( .A(n14), .B(n15), .Z(n12) );
  XNOR U274 ( .A(n13), .B(n16), .Z(n15) );
  XOR U275 ( .A(n17), .B(n18), .Z(n3) );
  ANDN U276 ( .B(n19), .A(n20), .Z(n17) );
  XOR U277 ( .A(n18), .B(n21), .Z(n19) );
  XNOR U278 ( .A(n4), .B(n22), .Z(n7) );
  XNOR U279 ( .A(n23), .B(n24), .Z(n22) );
  ANDN U280 ( .B(n25), .A(n26), .Z(n23) );
  XNOR U281 ( .A(n27), .B(n28), .Z(n25) );
  IV U282 ( .A(n10), .Z(n4) );
  XOR U283 ( .A(n29), .B(n30), .Z(n10) );
  AND U284 ( .A(n31), .B(n32), .Z(n29) );
  XOR U285 ( .A(n33), .B(n30), .Z(n32) );
  XNOR U286 ( .A(n20), .B(n21), .Z(o[5]) );
  XNOR U287 ( .A(n34), .B(n35), .Z(n21) );
  ANDN U288 ( .B(n36), .A(n37), .Z(n34) );
  XOR U289 ( .A(n35), .B(n38), .Z(n36) );
  XOR U290 ( .A(n31), .B(n39), .Z(n20) );
  XOR U291 ( .A(n18), .B(n33), .Z(n39) );
  XNOR U292 ( .A(n14), .B(n16), .Z(n33) );
  XNOR U293 ( .A(n40), .B(n41), .Z(n16) );
  ANDN U294 ( .B(n42), .A(n43), .Z(n40) );
  XOR U295 ( .A(n41), .B(n44), .Z(n42) );
  XNOR U296 ( .A(n46), .B(n47), .Z(n45) );
  ANDN U297 ( .B(n48), .A(n49), .Z(n46) );
  XNOR U298 ( .A(n50), .B(n51), .Z(n48) );
  XOR U299 ( .A(n52), .B(n53), .Z(n13) );
  AND U300 ( .A(n54), .B(n55), .Z(n52) );
  XNOR U301 ( .A(n53), .B(n56), .Z(n55) );
  XOR U302 ( .A(n57), .B(n58), .Z(n18) );
  ANDN U303 ( .B(n59), .A(n60), .Z(n57) );
  XNOR U304 ( .A(n58), .B(n61), .Z(n59) );
  XNOR U305 ( .A(n27), .B(n63), .Z(n62) );
  IV U306 ( .A(n30), .Z(n63) );
  XOR U307 ( .A(n64), .B(n65), .Z(n30) );
  AND U308 ( .A(n66), .B(n67), .Z(n64) );
  XOR U309 ( .A(n68), .B(n65), .Z(n67) );
  XNOR U310 ( .A(n69), .B(n70), .Z(n27) );
  ANDN U311 ( .B(n71), .A(n72), .Z(n69) );
  XOR U312 ( .A(n70), .B(n73), .Z(n71) );
  XOR U313 ( .A(n24), .B(n74), .Z(n26) );
  XNOR U314 ( .A(n75), .B(n76), .Z(n74) );
  ANDN U315 ( .B(n77), .A(n78), .Z(n75) );
  XNOR U316 ( .A(n79), .B(n80), .Z(n77) );
  IV U317 ( .A(n28), .Z(n24) );
  XOR U318 ( .A(n81), .B(n82), .Z(n28) );
  AND U319 ( .A(n83), .B(n84), .Z(n81) );
  XOR U320 ( .A(n85), .B(n82), .Z(n84) );
  XOR U321 ( .A(n60), .B(n61), .Z(o[4]) );
  XNOR U322 ( .A(n86), .B(n87), .Z(n38) );
  ANDN U323 ( .B(n88), .A(n89), .Z(n86) );
  XOR U324 ( .A(n90), .B(n91), .Z(n88) );
  XNOR U325 ( .A(n93), .B(n94), .Z(n92) );
  ANDN U326 ( .B(n95), .A(n96), .Z(n93) );
  XNOR U327 ( .A(n97), .B(n98), .Z(n95) );
  XOR U328 ( .A(n99), .B(n100), .Z(n35) );
  ANDN U329 ( .B(n101), .A(n102), .Z(n99) );
  XOR U330 ( .A(n100), .B(n103), .Z(n101) );
  XOR U331 ( .A(n66), .B(n104), .Z(n60) );
  XOR U332 ( .A(n58), .B(n68), .Z(n104) );
  XNOR U333 ( .A(n54), .B(n56), .Z(n68) );
  XOR U334 ( .A(n43), .B(n44), .Z(n56) );
  XNOR U335 ( .A(n105), .B(n106), .Z(n44) );
  ANDN U336 ( .B(n107), .A(n108), .Z(n105) );
  XOR U337 ( .A(n109), .B(n110), .Z(n107) );
  XNOR U338 ( .A(n112), .B(n113), .Z(n111) );
  ANDN U339 ( .B(n114), .A(n115), .Z(n112) );
  XNOR U340 ( .A(n116), .B(n117), .Z(n114) );
  XOR U341 ( .A(n118), .B(n119), .Z(n41) );
  ANDN U342 ( .B(n120), .A(n121), .Z(n118) );
  XOR U343 ( .A(n119), .B(n122), .Z(n120) );
  XNOR U344 ( .A(n50), .B(n124), .Z(n123) );
  IV U345 ( .A(n53), .Z(n124) );
  XOR U346 ( .A(n125), .B(n126), .Z(n53) );
  AND U347 ( .A(n127), .B(n128), .Z(n125) );
  XNOR U348 ( .A(n126), .B(n129), .Z(n128) );
  XNOR U349 ( .A(n130), .B(n131), .Z(n50) );
  ANDN U350 ( .B(n132), .A(n133), .Z(n130) );
  XOR U351 ( .A(n131), .B(n134), .Z(n132) );
  XOR U352 ( .A(n47), .B(n135), .Z(n49) );
  XNOR U353 ( .A(n136), .B(n137), .Z(n135) );
  ANDN U354 ( .B(n138), .A(n139), .Z(n136) );
  XNOR U355 ( .A(n140), .B(n141), .Z(n138) );
  IV U356 ( .A(n51), .Z(n47) );
  XOR U357 ( .A(n142), .B(n143), .Z(n51) );
  ANDN U358 ( .B(n144), .A(n145), .Z(n142) );
  XOR U359 ( .A(n146), .B(n143), .Z(n144) );
  XOR U360 ( .A(n147), .B(n148), .Z(n58) );
  ANDN U361 ( .B(n149), .A(n150), .Z(n147) );
  XNOR U362 ( .A(n148), .B(n151), .Z(n149) );
  XNOR U363 ( .A(n83), .B(n152), .Z(n66) );
  XOR U364 ( .A(n153), .B(n154), .Z(n65) );
  AND U365 ( .A(n155), .B(n156), .Z(n153) );
  XOR U366 ( .A(n157), .B(n154), .Z(n156) );
  XNOR U367 ( .A(n158), .B(n159), .Z(n73) );
  ANDN U368 ( .B(n160), .A(n161), .Z(n158) );
  XOR U369 ( .A(n162), .B(n163), .Z(n160) );
  XNOR U370 ( .A(n165), .B(n166), .Z(n164) );
  ANDN U371 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U372 ( .A(n169), .B(n170), .Z(n167) );
  XOR U373 ( .A(n171), .B(n172), .Z(n70) );
  ANDN U374 ( .B(n173), .A(n174), .Z(n171) );
  XOR U375 ( .A(n172), .B(n175), .Z(n173) );
  XNOR U376 ( .A(n79), .B(n177), .Z(n176) );
  IV U377 ( .A(n82), .Z(n177) );
  XOR U378 ( .A(n178), .B(n179), .Z(n82) );
  AND U379 ( .A(n180), .B(n181), .Z(n178) );
  XOR U380 ( .A(n182), .B(n179), .Z(n181) );
  XNOR U381 ( .A(n183), .B(n184), .Z(n79) );
  ANDN U382 ( .B(n185), .A(n186), .Z(n183) );
  XOR U383 ( .A(n184), .B(n187), .Z(n185) );
  XOR U384 ( .A(n76), .B(n188), .Z(n78) );
  XNOR U385 ( .A(n189), .B(n190), .Z(n188) );
  ANDN U386 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U387 ( .A(n193), .B(n194), .Z(n191) );
  IV U388 ( .A(n80), .Z(n76) );
  XOR U389 ( .A(n195), .B(n196), .Z(n80) );
  AND U390 ( .A(n197), .B(n198), .Z(n195) );
  XOR U391 ( .A(n199), .B(n196), .Z(n198) );
  XOR U392 ( .A(n150), .B(n151), .Z(o[3]) );
  XNOR U393 ( .A(n200), .B(n201), .Z(n91) );
  ANDN U394 ( .B(n202), .A(n203), .Z(n200) );
  XNOR U395 ( .A(n201), .B(n204), .Z(n202) );
  XOR U396 ( .A(n87), .B(n205), .Z(n89) );
  XNOR U397 ( .A(n206), .B(n207), .Z(n205) );
  ANDN U398 ( .B(n208), .A(n209), .Z(n206) );
  XNOR U399 ( .A(n210), .B(n211), .Z(n208) );
  IV U400 ( .A(n90), .Z(n87) );
  XOR U401 ( .A(n212), .B(n213), .Z(n90) );
  ANDN U402 ( .B(n214), .A(n215), .Z(n212) );
  XOR U403 ( .A(n213), .B(n216), .Z(n214) );
  XNOR U404 ( .A(n97), .B(n218), .Z(n217) );
  IV U405 ( .A(n100), .Z(n218) );
  XOR U406 ( .A(n219), .B(n220), .Z(n100) );
  ANDN U407 ( .B(n221), .A(n222), .Z(n219) );
  XOR U408 ( .A(n220), .B(n223), .Z(n221) );
  XOR U409 ( .A(n224), .B(n225), .Z(n97) );
  ANDN U410 ( .B(n226), .A(n227), .Z(n224) );
  XNOR U411 ( .A(n225), .B(n228), .Z(n226) );
  XOR U412 ( .A(n94), .B(n229), .Z(n96) );
  XNOR U413 ( .A(n230), .B(n231), .Z(n229) );
  ANDN U414 ( .B(n232), .A(n233), .Z(n230) );
  XNOR U415 ( .A(n234), .B(n235), .Z(n232) );
  IV U416 ( .A(n98), .Z(n94) );
  XOR U417 ( .A(n236), .B(n237), .Z(n98) );
  ANDN U418 ( .B(n238), .A(n239), .Z(n236) );
  XOR U419 ( .A(n240), .B(n237), .Z(n238) );
  XOR U420 ( .A(n155), .B(n241), .Z(n150) );
  XOR U421 ( .A(n148), .B(n157), .Z(n241) );
  XNOR U422 ( .A(n127), .B(n129), .Z(n157) );
  XOR U423 ( .A(n121), .B(n122), .Z(n129) );
  XNOR U424 ( .A(n242), .B(n243), .Z(n110) );
  ANDN U425 ( .B(n244), .A(n245), .Z(n242) );
  XNOR U426 ( .A(n243), .B(n246), .Z(n244) );
  XOR U427 ( .A(n106), .B(n247), .Z(n108) );
  XNOR U428 ( .A(n248), .B(n249), .Z(n247) );
  ANDN U429 ( .B(n250), .A(n251), .Z(n248) );
  XNOR U430 ( .A(n252), .B(n253), .Z(n250) );
  IV U431 ( .A(n109), .Z(n106) );
  XOR U432 ( .A(n254), .B(n255), .Z(n109) );
  ANDN U433 ( .B(n256), .A(n257), .Z(n254) );
  XOR U434 ( .A(n255), .B(n258), .Z(n256) );
  XNOR U435 ( .A(n116), .B(n260), .Z(n259) );
  IV U436 ( .A(n119), .Z(n260) );
  XOR U437 ( .A(n261), .B(n262), .Z(n119) );
  ANDN U438 ( .B(n263), .A(n264), .Z(n261) );
  XOR U439 ( .A(n262), .B(n265), .Z(n263) );
  XOR U440 ( .A(n266), .B(n267), .Z(n116) );
  ANDN U441 ( .B(n268), .A(n269), .Z(n266) );
  XNOR U442 ( .A(n267), .B(n270), .Z(n268) );
  XOR U443 ( .A(n113), .B(n271), .Z(n115) );
  XNOR U444 ( .A(n272), .B(n273), .Z(n271) );
  ANDN U445 ( .B(n274), .A(n275), .Z(n272) );
  XNOR U446 ( .A(n276), .B(n277), .Z(n274) );
  IV U447 ( .A(n117), .Z(n113) );
  XOR U448 ( .A(n278), .B(n279), .Z(n117) );
  ANDN U449 ( .B(n280), .A(n281), .Z(n278) );
  XOR U450 ( .A(n282), .B(n279), .Z(n280) );
  XOR U451 ( .A(n146), .B(n284), .Z(n283) );
  IV U452 ( .A(n126), .Z(n284) );
  XOR U453 ( .A(n285), .B(n286), .Z(n126) );
  AND U454 ( .A(n287), .B(n288), .Z(n285) );
  XNOR U455 ( .A(n286), .B(n289), .Z(n288) );
  XNOR U456 ( .A(n290), .B(n291), .Z(n134) );
  ANDN U457 ( .B(n292), .A(n293), .Z(n290) );
  XNOR U458 ( .A(n291), .B(n294), .Z(n292) );
  XNOR U459 ( .A(n296), .B(n297), .Z(n295) );
  ANDN U460 ( .B(n298), .A(n299), .Z(n296) );
  XNOR U461 ( .A(n300), .B(n301), .Z(n298) );
  XOR U462 ( .A(n302), .B(n303), .Z(n131) );
  ANDN U463 ( .B(n304), .A(n305), .Z(n302) );
  XOR U464 ( .A(n303), .B(n306), .Z(n304) );
  XNOR U465 ( .A(n140), .B(n308), .Z(n307) );
  IV U466 ( .A(n143), .Z(n308) );
  XOR U467 ( .A(n309), .B(n310), .Z(n143) );
  ANDN U468 ( .B(n311), .A(n312), .Z(n309) );
  XOR U469 ( .A(n313), .B(n310), .Z(n311) );
  XOR U470 ( .A(n314), .B(n315), .Z(n140) );
  ANDN U471 ( .B(n316), .A(n317), .Z(n314) );
  XNOR U472 ( .A(n315), .B(n318), .Z(n316) );
  XOR U473 ( .A(n137), .B(n319), .Z(n139) );
  XNOR U474 ( .A(n320), .B(n321), .Z(n319) );
  ANDN U475 ( .B(n322), .A(n323), .Z(n320) );
  XNOR U476 ( .A(n324), .B(n325), .Z(n322) );
  IV U477 ( .A(n141), .Z(n137) );
  XOR U478 ( .A(n326), .B(n327), .Z(n141) );
  ANDN U479 ( .B(n328), .A(n329), .Z(n326) );
  XOR U480 ( .A(n330), .B(n327), .Z(n328) );
  XNOR U481 ( .A(n331), .B(n332), .Z(n148) );
  ANDN U482 ( .B(n333), .A(n334), .Z(n331) );
  XOR U483 ( .A(n332), .B(n335), .Z(n333) );
  XNOR U484 ( .A(n180), .B(n336), .Z(n155) );
  XOR U485 ( .A(n337), .B(n338), .Z(n154) );
  AND U486 ( .A(n339), .B(n340), .Z(n337) );
  XOR U487 ( .A(n341), .B(n338), .Z(n340) );
  XNOR U488 ( .A(n342), .B(n343), .Z(n163) );
  ANDN U489 ( .B(n344), .A(n345), .Z(n342) );
  XNOR U490 ( .A(n343), .B(n346), .Z(n344) );
  XOR U491 ( .A(n159), .B(n347), .Z(n161) );
  XNOR U492 ( .A(n348), .B(n349), .Z(n347) );
  ANDN U493 ( .B(n350), .A(n351), .Z(n348) );
  XNOR U494 ( .A(n352), .B(n353), .Z(n350) );
  IV U495 ( .A(n162), .Z(n159) );
  XOR U496 ( .A(n354), .B(n355), .Z(n162) );
  ANDN U497 ( .B(n356), .A(n357), .Z(n354) );
  XOR U498 ( .A(n355), .B(n358), .Z(n356) );
  XNOR U499 ( .A(n169), .B(n360), .Z(n359) );
  IV U500 ( .A(n172), .Z(n360) );
  XOR U501 ( .A(n361), .B(n362), .Z(n172) );
  ANDN U502 ( .B(n363), .A(n364), .Z(n361) );
  XOR U503 ( .A(n362), .B(n365), .Z(n363) );
  XOR U504 ( .A(n366), .B(n367), .Z(n169) );
  ANDN U505 ( .B(n368), .A(n369), .Z(n366) );
  XNOR U506 ( .A(n367), .B(n370), .Z(n368) );
  XOR U507 ( .A(n166), .B(n371), .Z(n168) );
  XNOR U508 ( .A(n372), .B(n373), .Z(n371) );
  ANDN U509 ( .B(n374), .A(n375), .Z(n372) );
  XNOR U510 ( .A(n376), .B(n377), .Z(n374) );
  IV U511 ( .A(n170), .Z(n166) );
  XOR U512 ( .A(n378), .B(n379), .Z(n170) );
  ANDN U513 ( .B(n380), .A(n381), .Z(n378) );
  XOR U514 ( .A(n382), .B(n379), .Z(n380) );
  XNOR U515 ( .A(n197), .B(n383), .Z(n180) );
  XOR U516 ( .A(n384), .B(n385), .Z(n179) );
  AND U517 ( .A(n386), .B(n387), .Z(n384) );
  XOR U518 ( .A(n388), .B(n385), .Z(n387) );
  XNOR U519 ( .A(n389), .B(n390), .Z(n187) );
  ANDN U520 ( .B(n391), .A(n392), .Z(n389) );
  XNOR U521 ( .A(n390), .B(n393), .Z(n391) );
  XNOR U522 ( .A(n395), .B(n396), .Z(n394) );
  ANDN U523 ( .B(n397), .A(n398), .Z(n395) );
  XNOR U524 ( .A(n399), .B(n400), .Z(n397) );
  XOR U525 ( .A(n401), .B(n402), .Z(n184) );
  ANDN U526 ( .B(n403), .A(n404), .Z(n401) );
  XOR U527 ( .A(n402), .B(n405), .Z(n403) );
  XNOR U528 ( .A(n193), .B(n407), .Z(n406) );
  IV U529 ( .A(n196), .Z(n407) );
  XOR U530 ( .A(n408), .B(n409), .Z(n196) );
  AND U531 ( .A(n410), .B(n411), .Z(n408) );
  XOR U532 ( .A(n412), .B(n409), .Z(n411) );
  XOR U533 ( .A(n413), .B(n414), .Z(n193) );
  ANDN U534 ( .B(n415), .A(n416), .Z(n413) );
  XNOR U535 ( .A(n414), .B(n417), .Z(n415) );
  XOR U536 ( .A(n190), .B(n418), .Z(n192) );
  XNOR U537 ( .A(n419), .B(n420), .Z(n418) );
  ANDN U538 ( .B(n421), .A(n422), .Z(n419) );
  XNOR U539 ( .A(n423), .B(n424), .Z(n421) );
  IV U540 ( .A(n194), .Z(n190) );
  XOR U541 ( .A(n425), .B(n426), .Z(n194) );
  AND U542 ( .A(n427), .B(n428), .Z(n425) );
  XOR U543 ( .A(n429), .B(n426), .Z(n428) );
  XOR U544 ( .A(n334), .B(n335), .Z(o[2]) );
  XNOR U545 ( .A(n430), .B(n431), .Z(n204) );
  NANDN U546 ( .A(n432), .B(n433), .Z(n431) );
  NANDN U547 ( .A(n434), .B(n430), .Z(n433) );
  XNOR U548 ( .A(n435), .B(n201), .Z(n203) );
  XNOR U549 ( .A(n436), .B(n437), .Z(n201) );
  NAND U550 ( .A(n438), .B(n439), .Z(n437) );
  XNOR U551 ( .A(n436), .B(n440), .Z(n438) );
  NOR U552 ( .A(n441), .B(n442), .Z(n435) );
  XOR U553 ( .A(n210), .B(n213), .Z(n443) );
  XNOR U554 ( .A(n444), .B(n445), .Z(n213) );
  NANDN U555 ( .A(n446), .B(n447), .Z(n445) );
  XOR U556 ( .A(n444), .B(n448), .Z(n447) );
  XNOR U557 ( .A(n449), .B(n450), .Z(n210) );
  NANDN U558 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U559 ( .A(n449), .B(n453), .Z(n452) );
  XOR U560 ( .A(n454), .B(n211), .Z(n209) );
  IV U561 ( .A(n207), .Z(n211) );
  XNOR U562 ( .A(n455), .B(n456), .Z(n207) );
  NAND U563 ( .A(n457), .B(n458), .Z(n456) );
  XOR U564 ( .A(n455), .B(n459), .Z(n457) );
  NOR U565 ( .A(n460), .B(n461), .Z(n454) );
  XNOR U566 ( .A(n240), .B(n220), .Z(n462) );
  XNOR U567 ( .A(n463), .B(n464), .Z(n220) );
  NANDN U568 ( .A(n465), .B(n466), .Z(n464) );
  XOR U569 ( .A(n463), .B(n467), .Z(n466) );
  XNOR U570 ( .A(n468), .B(n469), .Z(n228) );
  NANDN U571 ( .A(n470), .B(n471), .Z(n469) );
  NANDN U572 ( .A(n472), .B(n468), .Z(n471) );
  XNOR U573 ( .A(n473), .B(n225), .Z(n227) );
  XNOR U574 ( .A(n474), .B(n475), .Z(n225) );
  NAND U575 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U576 ( .A(n474), .B(n478), .Z(n476) );
  NOR U577 ( .A(n479), .B(n480), .Z(n473) );
  XOR U578 ( .A(n234), .B(n237), .Z(n481) );
  XNOR U579 ( .A(n482), .B(n483), .Z(n237) );
  NANDN U580 ( .A(n484), .B(n485), .Z(n483) );
  XNOR U581 ( .A(n482), .B(n486), .Z(n485) );
  XNOR U582 ( .A(n487), .B(n488), .Z(n234) );
  NANDN U583 ( .A(n489), .B(n490), .Z(n488) );
  NANDN U584 ( .A(n487), .B(n491), .Z(n490) );
  XOR U585 ( .A(n492), .B(n235), .Z(n233) );
  IV U586 ( .A(n231), .Z(n235) );
  XNOR U587 ( .A(n493), .B(n494), .Z(n231) );
  NAND U588 ( .A(n495), .B(n496), .Z(n494) );
  XOR U589 ( .A(n493), .B(n497), .Z(n495) );
  NOR U590 ( .A(n498), .B(n499), .Z(n492) );
  XOR U591 ( .A(n339), .B(n500), .Z(n334) );
  XNOR U592 ( .A(n332), .B(n341), .Z(n500) );
  XNOR U593 ( .A(n287), .B(n289), .Z(n341) );
  XOR U594 ( .A(n264), .B(n265), .Z(n289) );
  XNOR U595 ( .A(n501), .B(n502), .Z(n246) );
  NANDN U596 ( .A(n503), .B(n504), .Z(n502) );
  NANDN U597 ( .A(n505), .B(n501), .Z(n504) );
  XNOR U598 ( .A(n506), .B(n243), .Z(n245) );
  XNOR U599 ( .A(n507), .B(n508), .Z(n243) );
  NAND U600 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U601 ( .A(n507), .B(n511), .Z(n509) );
  NOR U602 ( .A(n512), .B(n513), .Z(n506) );
  XOR U603 ( .A(n252), .B(n255), .Z(n514) );
  XNOR U604 ( .A(n515), .B(n516), .Z(n255) );
  NANDN U605 ( .A(n517), .B(n518), .Z(n516) );
  XOR U606 ( .A(n515), .B(n519), .Z(n518) );
  XNOR U607 ( .A(n520), .B(n521), .Z(n252) );
  NANDN U608 ( .A(n522), .B(n523), .Z(n521) );
  NANDN U609 ( .A(n520), .B(n524), .Z(n523) );
  XOR U610 ( .A(n525), .B(n253), .Z(n251) );
  IV U611 ( .A(n249), .Z(n253) );
  XNOR U612 ( .A(n526), .B(n527), .Z(n249) );
  NAND U613 ( .A(n528), .B(n529), .Z(n527) );
  XOR U614 ( .A(n526), .B(n530), .Z(n528) );
  NOR U615 ( .A(n531), .B(n532), .Z(n525) );
  XNOR U616 ( .A(n282), .B(n262), .Z(n533) );
  XNOR U617 ( .A(n534), .B(n535), .Z(n262) );
  NANDN U618 ( .A(n536), .B(n537), .Z(n535) );
  XOR U619 ( .A(n534), .B(n538), .Z(n537) );
  XNOR U620 ( .A(n539), .B(n540), .Z(n270) );
  NANDN U621 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U622 ( .A(n543), .B(n539), .Z(n542) );
  XNOR U623 ( .A(n544), .B(n267), .Z(n269) );
  XNOR U624 ( .A(n545), .B(n546), .Z(n267) );
  NAND U625 ( .A(n547), .B(n548), .Z(n546) );
  XNOR U626 ( .A(n545), .B(n549), .Z(n547) );
  NOR U627 ( .A(n550), .B(n551), .Z(n544) );
  XOR U628 ( .A(n276), .B(n279), .Z(n552) );
  XNOR U629 ( .A(n553), .B(n554), .Z(n279) );
  NANDN U630 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U631 ( .A(n553), .B(n557), .Z(n556) );
  XNOR U632 ( .A(n558), .B(n559), .Z(n276) );
  NANDN U633 ( .A(n560), .B(n561), .Z(n559) );
  NANDN U634 ( .A(n558), .B(n562), .Z(n561) );
  XOR U635 ( .A(n563), .B(n277), .Z(n275) );
  IV U636 ( .A(n273), .Z(n277) );
  XNOR U637 ( .A(n564), .B(n565), .Z(n273) );
  NAND U638 ( .A(n566), .B(n567), .Z(n565) );
  XOR U639 ( .A(n564), .B(n568), .Z(n566) );
  NOR U640 ( .A(n569), .B(n570), .Z(n563) );
  XNOR U641 ( .A(n313), .B(n286), .Z(n571) );
  XNOR U642 ( .A(n572), .B(n573), .Z(n286) );
  NAND U643 ( .A(n574), .B(n575), .Z(n573) );
  XNOR U644 ( .A(n572), .B(n576), .Z(n574) );
  XOR U645 ( .A(n577), .B(n294), .Z(n306) );
  XNOR U646 ( .A(n578), .B(n579), .Z(n294) );
  NANDN U647 ( .A(n580), .B(n581), .Z(n579) );
  NANDN U648 ( .A(n582), .B(n578), .Z(n581) );
  IV U649 ( .A(n293), .Z(n577) );
  XNOR U650 ( .A(n583), .B(n291), .Z(n293) );
  XNOR U651 ( .A(n584), .B(n585), .Z(n291) );
  NAND U652 ( .A(n586), .B(n587), .Z(n585) );
  XNOR U653 ( .A(n584), .B(n588), .Z(n586) );
  NOR U654 ( .A(n589), .B(n590), .Z(n583) );
  XOR U655 ( .A(n300), .B(n303), .Z(n591) );
  XNOR U656 ( .A(n592), .B(n593), .Z(n303) );
  NANDN U657 ( .A(n594), .B(n595), .Z(n593) );
  XOR U658 ( .A(n592), .B(n596), .Z(n595) );
  XNOR U659 ( .A(n597), .B(n598), .Z(n300) );
  NANDN U660 ( .A(n599), .B(n600), .Z(n598) );
  NANDN U661 ( .A(n597), .B(n601), .Z(n600) );
  XOR U662 ( .A(n602), .B(n301), .Z(n299) );
  IV U663 ( .A(n297), .Z(n301) );
  XNOR U664 ( .A(n603), .B(n604), .Z(n297) );
  NAND U665 ( .A(n605), .B(n606), .Z(n604) );
  XOR U666 ( .A(n603), .B(n607), .Z(n605) );
  NOR U667 ( .A(n608), .B(n609), .Z(n602) );
  XNOR U668 ( .A(n330), .B(n310), .Z(n610) );
  XNOR U669 ( .A(n611), .B(n612), .Z(n310) );
  NANDN U670 ( .A(n613), .B(n614), .Z(n612) );
  XOR U671 ( .A(n611), .B(n615), .Z(n614) );
  XNOR U672 ( .A(n616), .B(n617), .Z(n318) );
  NANDN U673 ( .A(n618), .B(n619), .Z(n617) );
  NANDN U674 ( .A(n620), .B(n616), .Z(n619) );
  XNOR U675 ( .A(n621), .B(n315), .Z(n317) );
  XNOR U676 ( .A(n622), .B(n623), .Z(n315) );
  NAND U677 ( .A(n624), .B(n625), .Z(n623) );
  XNOR U678 ( .A(n622), .B(n626), .Z(n624) );
  NOR U679 ( .A(n627), .B(n628), .Z(n621) );
  XOR U680 ( .A(n324), .B(n327), .Z(n629) );
  XNOR U681 ( .A(n630), .B(n631), .Z(n327) );
  NANDN U682 ( .A(n632), .B(n633), .Z(n631) );
  XNOR U683 ( .A(n630), .B(n634), .Z(n633) );
  XNOR U684 ( .A(n635), .B(n636), .Z(n324) );
  NANDN U685 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U686 ( .A(n635), .B(n639), .Z(n638) );
  XOR U687 ( .A(n640), .B(n325), .Z(n323) );
  IV U688 ( .A(n321), .Z(n325) );
  XNOR U689 ( .A(n641), .B(n642), .Z(n321) );
  NAND U690 ( .A(n643), .B(n644), .Z(n642) );
  XOR U691 ( .A(n641), .B(n645), .Z(n643) );
  NOR U692 ( .A(n646), .B(n647), .Z(n640) );
  XNOR U693 ( .A(n648), .B(n649), .Z(n332) );
  NANDN U694 ( .A(n650), .B(n651), .Z(n649) );
  XOR U695 ( .A(n648), .B(n652), .Z(n651) );
  XNOR U696 ( .A(n386), .B(n653), .Z(n339) );
  XNOR U697 ( .A(n388), .B(n338), .Z(n653) );
  XNOR U698 ( .A(n654), .B(n655), .Z(n338) );
  NAND U699 ( .A(n656), .B(n657), .Z(n655) );
  XOR U700 ( .A(n654), .B(n658), .Z(n656) );
  XNOR U701 ( .A(n659), .B(n660), .Z(n346) );
  NANDN U702 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U703 ( .A(n663), .B(n659), .Z(n662) );
  XNOR U704 ( .A(n664), .B(n343), .Z(n345) );
  XNOR U705 ( .A(n665), .B(n666), .Z(n343) );
  NAND U706 ( .A(n667), .B(n668), .Z(n666) );
  XNOR U707 ( .A(n665), .B(n669), .Z(n667) );
  NOR U708 ( .A(n670), .B(n671), .Z(n664) );
  XOR U709 ( .A(n352), .B(n355), .Z(n672) );
  XNOR U710 ( .A(n673), .B(n674), .Z(n355) );
  NANDN U711 ( .A(n675), .B(n676), .Z(n674) );
  XOR U712 ( .A(n673), .B(n677), .Z(n676) );
  XNOR U713 ( .A(n678), .B(n679), .Z(n352) );
  NANDN U714 ( .A(n680), .B(n681), .Z(n679) );
  NANDN U715 ( .A(n678), .B(n682), .Z(n681) );
  XOR U716 ( .A(n683), .B(n353), .Z(n351) );
  IV U717 ( .A(n349), .Z(n353) );
  XNOR U718 ( .A(n684), .B(n685), .Z(n349) );
  NAND U719 ( .A(n686), .B(n687), .Z(n685) );
  XOR U720 ( .A(n684), .B(n688), .Z(n686) );
  NOR U721 ( .A(n689), .B(n690), .Z(n683) );
  XNOR U722 ( .A(n382), .B(n362), .Z(n691) );
  XNOR U723 ( .A(n692), .B(n693), .Z(n362) );
  NANDN U724 ( .A(n694), .B(n695), .Z(n693) );
  XOR U725 ( .A(n692), .B(n696), .Z(n695) );
  XNOR U726 ( .A(n697), .B(n698), .Z(n370) );
  NANDN U727 ( .A(n699), .B(n700), .Z(n698) );
  NANDN U728 ( .A(n701), .B(n697), .Z(n700) );
  XNOR U729 ( .A(n702), .B(n367), .Z(n369) );
  XNOR U730 ( .A(n703), .B(n704), .Z(n367) );
  NAND U731 ( .A(n705), .B(n706), .Z(n704) );
  XNOR U732 ( .A(n703), .B(n707), .Z(n705) );
  NOR U733 ( .A(n708), .B(n709), .Z(n702) );
  XOR U734 ( .A(n376), .B(n379), .Z(n710) );
  XNOR U735 ( .A(n711), .B(n712), .Z(n379) );
  NANDN U736 ( .A(n713), .B(n714), .Z(n712) );
  XNOR U737 ( .A(n711), .B(n715), .Z(n714) );
  XNOR U738 ( .A(n716), .B(n717), .Z(n376) );
  NANDN U739 ( .A(n718), .B(n719), .Z(n717) );
  NANDN U740 ( .A(n716), .B(n720), .Z(n719) );
  XOR U741 ( .A(n721), .B(n377), .Z(n375) );
  IV U742 ( .A(n373), .Z(n377) );
  XNOR U743 ( .A(n722), .B(n723), .Z(n373) );
  NAND U744 ( .A(n724), .B(n725), .Z(n723) );
  XOR U745 ( .A(n722), .B(n726), .Z(n724) );
  NOR U746 ( .A(n727), .B(n728), .Z(n721) );
  XNOR U747 ( .A(n410), .B(n729), .Z(n386) );
  XNOR U748 ( .A(n412), .B(n385), .Z(n729) );
  XOR U749 ( .A(n730), .B(n731), .Z(n385) );
  NAND U750 ( .A(n732), .B(n733), .Z(n731) );
  XNOR U751 ( .A(n730), .B(n734), .Z(n732) );
  XOR U752 ( .A(n735), .B(n393), .Z(n405) );
  XNOR U753 ( .A(n736), .B(n737), .Z(n393) );
  NANDN U754 ( .A(n738), .B(n739), .Z(n737) );
  NANDN U755 ( .A(n740), .B(n736), .Z(n739) );
  IV U756 ( .A(n392), .Z(n735) );
  XNOR U757 ( .A(n741), .B(n390), .Z(n392) );
  XNOR U758 ( .A(n742), .B(n743), .Z(n390) );
  NAND U759 ( .A(n744), .B(n745), .Z(n743) );
  XNOR U760 ( .A(n742), .B(n746), .Z(n744) );
  NOR U761 ( .A(n747), .B(n748), .Z(n741) );
  XOR U762 ( .A(n399), .B(n402), .Z(n749) );
  XNOR U763 ( .A(n750), .B(n751), .Z(n402) );
  NANDN U764 ( .A(n752), .B(n753), .Z(n751) );
  XOR U765 ( .A(n750), .B(n754), .Z(n753) );
  XNOR U766 ( .A(n755), .B(n756), .Z(n399) );
  NANDN U767 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U768 ( .A(n755), .B(n759), .Z(n758) );
  XOR U769 ( .A(n760), .B(n400), .Z(n398) );
  IV U770 ( .A(n396), .Z(n400) );
  XNOR U771 ( .A(n761), .B(n762), .Z(n396) );
  NAND U772 ( .A(n763), .B(n764), .Z(n762) );
  XOR U773 ( .A(n761), .B(n765), .Z(n763) );
  NOR U774 ( .A(n766), .B(n767), .Z(n760) );
  XNOR U775 ( .A(n427), .B(n768), .Z(n410) );
  XNOR U776 ( .A(n429), .B(n409), .Z(n768) );
  XOR U777 ( .A(n769), .B(n770), .Z(n409) );
  NAND U778 ( .A(n771), .B(n772), .Z(n770) );
  XNOR U779 ( .A(n769), .B(n773), .Z(n771) );
  XNOR U780 ( .A(n774), .B(n775), .Z(n417) );
  NANDN U781 ( .A(n776), .B(n777), .Z(n775) );
  NANDN U782 ( .A(n778), .B(n774), .Z(n777) );
  XNOR U783 ( .A(n779), .B(n414), .Z(n416) );
  XNOR U784 ( .A(n780), .B(n781), .Z(n414) );
  NAND U785 ( .A(n782), .B(n783), .Z(n781) );
  XNOR U786 ( .A(n780), .B(n784), .Z(n782) );
  NOR U787 ( .A(n785), .B(n786), .Z(n779) );
  XOR U788 ( .A(n423), .B(n426), .Z(n787) );
  XNOR U789 ( .A(n788), .B(n789), .Z(n426) );
  NAND U790 ( .A(n790), .B(n791), .Z(n789) );
  XNOR U791 ( .A(n793), .B(n794), .Z(n423) );
  NANDN U792 ( .A(n795), .B(n796), .Z(n794) );
  NANDN U793 ( .A(n793), .B(n797), .Z(n796) );
  XOR U794 ( .A(n798), .B(n424), .Z(n422) );
  IV U795 ( .A(n420), .Z(n424) );
  XNOR U796 ( .A(n799), .B(n800), .Z(n420) );
  NANDN U797 ( .A(n801), .B(n802), .Z(n800) );
  XOR U798 ( .A(n799), .B(n803), .Z(n802) );
  NOR U799 ( .A(n804), .B(n805), .Z(n798) );
  XOR U800 ( .A(n650), .B(n652), .Z(o[1]) );
  XOR U801 ( .A(n439), .B(n440), .Z(n448) );
  XOR U802 ( .A(n434), .B(n432), .Z(n440) );
  AND U803 ( .A(n806), .B(n430), .Z(n432) );
  OR U804 ( .A(n807), .B(n808), .Z(n430) );
  OR U805 ( .A(n809), .B(n810), .Z(n806) );
  NOR U806 ( .A(n811), .B(n812), .Z(n434) );
  XOR U807 ( .A(n441), .B(n813), .Z(n439) );
  XOR U808 ( .A(n442), .B(n436), .Z(n813) );
  NOR U809 ( .A(n814), .B(n815), .Z(n436) );
  OR U810 ( .A(n816), .B(n817), .Z(n442) );
  AND U811 ( .A(n818), .B(n819), .Z(n441) );
  OR U812 ( .A(n820), .B(n821), .Z(n819) );
  OR U813 ( .A(n822), .B(n823), .Z(n818) );
  XNOR U814 ( .A(n458), .B(n824), .Z(n446) );
  XNOR U815 ( .A(n444), .B(n459), .Z(n824) );
  XOR U816 ( .A(n453), .B(n451), .Z(n459) );
  NOR U817 ( .A(n826), .B(n827), .Z(n449) );
  OR U818 ( .A(n828), .B(n829), .Z(n825) );
  OR U819 ( .A(n830), .B(n831), .Z(n453) );
  OR U820 ( .A(n832), .B(n833), .Z(n444) );
  XOR U821 ( .A(n460), .B(n834), .Z(n458) );
  XOR U822 ( .A(n461), .B(n455), .Z(n834) );
  NOR U823 ( .A(n835), .B(n836), .Z(n455) );
  OR U824 ( .A(n837), .B(n838), .Z(n461) );
  AND U825 ( .A(n839), .B(n840), .Z(n460) );
  OR U826 ( .A(n841), .B(n842), .Z(n840) );
  OR U827 ( .A(n843), .B(n844), .Z(n839) );
  XOR U828 ( .A(n463), .B(n486), .Z(n845) );
  XNOR U829 ( .A(n477), .B(n478), .Z(n486) );
  XOR U830 ( .A(n472), .B(n470), .Z(n478) );
  AND U831 ( .A(n846), .B(n468), .Z(n470) );
  OR U832 ( .A(n847), .B(n848), .Z(n468) );
  OR U833 ( .A(n849), .B(n850), .Z(n846) );
  NOR U834 ( .A(n851), .B(n852), .Z(n472) );
  XOR U835 ( .A(n479), .B(n853), .Z(n477) );
  XOR U836 ( .A(n480), .B(n474), .Z(n853) );
  NOR U837 ( .A(n854), .B(n855), .Z(n474) );
  OR U838 ( .A(n856), .B(n857), .Z(n480) );
  AND U839 ( .A(n858), .B(n859), .Z(n479) );
  OR U840 ( .A(n860), .B(n861), .Z(n859) );
  OR U841 ( .A(n862), .B(n863), .Z(n858) );
  OR U842 ( .A(n864), .B(n865), .Z(n463) );
  XNOR U843 ( .A(n496), .B(n866), .Z(n484) );
  XNOR U844 ( .A(n482), .B(n497), .Z(n866) );
  XOR U845 ( .A(n491), .B(n489), .Z(n497) );
  NOR U846 ( .A(n868), .B(n869), .Z(n487) );
  OR U847 ( .A(n870), .B(n871), .Z(n867) );
  OR U848 ( .A(n872), .B(n873), .Z(n491) );
  OR U849 ( .A(n874), .B(n875), .Z(n482) );
  XOR U850 ( .A(n498), .B(n876), .Z(n496) );
  XOR U851 ( .A(n499), .B(n493), .Z(n876) );
  NOR U852 ( .A(n877), .B(n878), .Z(n493) );
  OR U853 ( .A(n879), .B(n880), .Z(n499) );
  AND U854 ( .A(n881), .B(n882), .Z(n498) );
  OR U855 ( .A(n883), .B(n884), .Z(n882) );
  OR U856 ( .A(n885), .B(n886), .Z(n881) );
  XOR U857 ( .A(n657), .B(n887), .Z(n650) );
  XNOR U858 ( .A(n575), .B(n576), .Z(n658) );
  XOR U859 ( .A(n536), .B(n538), .Z(n576) );
  XOR U860 ( .A(n510), .B(n511), .Z(n519) );
  XOR U861 ( .A(n505), .B(n503), .Z(n511) );
  AND U862 ( .A(n888), .B(n501), .Z(n503) );
  OR U863 ( .A(n889), .B(n890), .Z(n501) );
  OR U864 ( .A(n891), .B(n892), .Z(n888) );
  NOR U865 ( .A(n893), .B(n894), .Z(n505) );
  XOR U866 ( .A(n512), .B(n895), .Z(n510) );
  XOR U867 ( .A(n513), .B(n507), .Z(n895) );
  NOR U868 ( .A(n896), .B(n897), .Z(n507) );
  OR U869 ( .A(n898), .B(n899), .Z(n513) );
  AND U870 ( .A(n900), .B(n901), .Z(n512) );
  OR U871 ( .A(n902), .B(n903), .Z(n901) );
  OR U872 ( .A(n904), .B(n905), .Z(n900) );
  XNOR U873 ( .A(n529), .B(n906), .Z(n517) );
  XNOR U874 ( .A(n515), .B(n530), .Z(n906) );
  XOR U875 ( .A(n524), .B(n522), .Z(n530) );
  NOR U876 ( .A(n908), .B(n909), .Z(n520) );
  OR U877 ( .A(n910), .B(n911), .Z(n907) );
  OR U878 ( .A(n912), .B(n913), .Z(n524) );
  OR U879 ( .A(n914), .B(n915), .Z(n515) );
  XOR U880 ( .A(n531), .B(n916), .Z(n529) );
  XOR U881 ( .A(n532), .B(n526), .Z(n916) );
  NOR U882 ( .A(n917), .B(n918), .Z(n526) );
  OR U883 ( .A(n919), .B(n920), .Z(n532) );
  AND U884 ( .A(n921), .B(n922), .Z(n531) );
  OR U885 ( .A(n923), .B(n924), .Z(n922) );
  OR U886 ( .A(n925), .B(n926), .Z(n921) );
  XOR U887 ( .A(n534), .B(n557), .Z(n927) );
  XNOR U888 ( .A(n548), .B(n549), .Z(n557) );
  XOR U889 ( .A(n543), .B(n541), .Z(n549) );
  AND U890 ( .A(n928), .B(n539), .Z(n541) );
  OR U891 ( .A(n929), .B(n930), .Z(n539) );
  OR U892 ( .A(n931), .B(n932), .Z(n928) );
  NOR U893 ( .A(n933), .B(n934), .Z(n543) );
  XOR U894 ( .A(n550), .B(n935), .Z(n548) );
  XOR U895 ( .A(n551), .B(n545), .Z(n935) );
  NOR U896 ( .A(n936), .B(n937), .Z(n545) );
  OR U897 ( .A(n938), .B(n939), .Z(n551) );
  AND U898 ( .A(n940), .B(n941), .Z(n550) );
  OR U899 ( .A(n942), .B(n943), .Z(n941) );
  OR U900 ( .A(n944), .B(n945), .Z(n940) );
  OR U901 ( .A(n946), .B(n947), .Z(n534) );
  XNOR U902 ( .A(n567), .B(n948), .Z(n555) );
  XNOR U903 ( .A(n553), .B(n568), .Z(n948) );
  XOR U904 ( .A(n562), .B(n560), .Z(n568) );
  NOR U905 ( .A(n950), .B(n951), .Z(n558) );
  OR U906 ( .A(n952), .B(n953), .Z(n949) );
  OR U907 ( .A(n954), .B(n955), .Z(n562) );
  OR U908 ( .A(n956), .B(n957), .Z(n553) );
  XOR U909 ( .A(n569), .B(n958), .Z(n567) );
  XOR U910 ( .A(n570), .B(n564), .Z(n958) );
  NOR U911 ( .A(n959), .B(n960), .Z(n564) );
  OR U912 ( .A(n961), .B(n962), .Z(n570) );
  AND U913 ( .A(n963), .B(n964), .Z(n569) );
  OR U914 ( .A(n965), .B(n966), .Z(n964) );
  OR U915 ( .A(n967), .B(n968), .Z(n963) );
  XNOR U916 ( .A(n572), .B(n615), .Z(n969) );
  XOR U917 ( .A(n587), .B(n588), .Z(n596) );
  XOR U918 ( .A(n582), .B(n580), .Z(n588) );
  AND U919 ( .A(n970), .B(n578), .Z(n580) );
  OR U920 ( .A(n971), .B(n972), .Z(n578) );
  OR U921 ( .A(n973), .B(n974), .Z(n970) );
  NOR U922 ( .A(n975), .B(n976), .Z(n582) );
  XOR U923 ( .A(n589), .B(n977), .Z(n587) );
  XOR U924 ( .A(n590), .B(n584), .Z(n977) );
  NOR U925 ( .A(n978), .B(n979), .Z(n584) );
  OR U926 ( .A(n980), .B(n981), .Z(n590) );
  AND U927 ( .A(n982), .B(n983), .Z(n589) );
  OR U928 ( .A(n984), .B(n985), .Z(n983) );
  OR U929 ( .A(n986), .B(n987), .Z(n982) );
  XNOR U930 ( .A(n606), .B(n988), .Z(n594) );
  XNOR U931 ( .A(n592), .B(n607), .Z(n988) );
  XOR U932 ( .A(n601), .B(n599), .Z(n607) );
  NOR U933 ( .A(n990), .B(n991), .Z(n597) );
  OR U934 ( .A(n992), .B(n993), .Z(n989) );
  OR U935 ( .A(n994), .B(n995), .Z(n601) );
  OR U936 ( .A(n996), .B(n997), .Z(n592) );
  XOR U937 ( .A(n608), .B(n998), .Z(n606) );
  XOR U938 ( .A(n609), .B(n603), .Z(n998) );
  NOR U939 ( .A(n999), .B(n1000), .Z(n603) );
  OR U940 ( .A(n1001), .B(n1002), .Z(n609) );
  AND U941 ( .A(n1003), .B(n1004), .Z(n608) );
  OR U942 ( .A(n1005), .B(n1006), .Z(n1004) );
  OR U943 ( .A(n1007), .B(n1008), .Z(n1003) );
  OR U944 ( .A(n1009), .B(n1010), .Z(n572) );
  XOR U945 ( .A(n611), .B(n634), .Z(n1011) );
  XNOR U946 ( .A(n625), .B(n626), .Z(n634) );
  XOR U947 ( .A(n620), .B(n618), .Z(n626) );
  AND U948 ( .A(n1012), .B(n616), .Z(n618) );
  OR U949 ( .A(n1013), .B(n1014), .Z(n616) );
  OR U950 ( .A(n1015), .B(n1016), .Z(n1012) );
  NOR U951 ( .A(n1017), .B(n1018), .Z(n620) );
  XOR U952 ( .A(n627), .B(n1019), .Z(n625) );
  XOR U953 ( .A(n628), .B(n622), .Z(n1019) );
  NOR U954 ( .A(n1020), .B(n1021), .Z(n622) );
  OR U955 ( .A(n1022), .B(n1023), .Z(n628) );
  AND U956 ( .A(n1024), .B(n1025), .Z(n627) );
  OR U957 ( .A(n1026), .B(n1027), .Z(n1025) );
  OR U958 ( .A(n1028), .B(n1029), .Z(n1024) );
  OR U959 ( .A(n1030), .B(n1031), .Z(n611) );
  XNOR U960 ( .A(n644), .B(n1032), .Z(n632) );
  XNOR U961 ( .A(n630), .B(n645), .Z(n1032) );
  XOR U962 ( .A(n639), .B(n637), .Z(n645) );
  NOR U963 ( .A(n1034), .B(n1035), .Z(n635) );
  OR U964 ( .A(n1036), .B(n1037), .Z(n1033) );
  OR U965 ( .A(n1038), .B(n1039), .Z(n639) );
  OR U966 ( .A(n1040), .B(n1041), .Z(n630) );
  XOR U967 ( .A(n646), .B(n1042), .Z(n644) );
  XOR U968 ( .A(n647), .B(n641), .Z(n1042) );
  NOR U969 ( .A(n1043), .B(n1044), .Z(n641) );
  OR U970 ( .A(n1045), .B(n1046), .Z(n647) );
  AND U971 ( .A(n1047), .B(n1048), .Z(n646) );
  OR U972 ( .A(n1049), .B(n1050), .Z(n1048) );
  OR U973 ( .A(n1051), .B(n1052), .Z(n1047) );
  NANDN U974 ( .A(n1053), .B(n1054), .Z(n648) );
  XNOR U975 ( .A(n733), .B(n1055), .Z(n657) );
  XNOR U976 ( .A(n654), .B(n734), .Z(n1055) );
  XOR U977 ( .A(n668), .B(n669), .Z(n677) );
  XOR U978 ( .A(n663), .B(n661), .Z(n669) );
  AND U979 ( .A(n1056), .B(n659), .Z(n661) );
  OR U980 ( .A(n1057), .B(n1058), .Z(n659) );
  OR U981 ( .A(n1059), .B(n1060), .Z(n1056) );
  NOR U982 ( .A(n1061), .B(n1062), .Z(n663) );
  XOR U983 ( .A(n670), .B(n1063), .Z(n668) );
  XOR U984 ( .A(n671), .B(n665), .Z(n1063) );
  NOR U985 ( .A(n1064), .B(n1065), .Z(n665) );
  OR U986 ( .A(n1066), .B(n1067), .Z(n671) );
  AND U987 ( .A(n1068), .B(n1069), .Z(n670) );
  OR U988 ( .A(n1070), .B(n1071), .Z(n1069) );
  OR U989 ( .A(n1072), .B(n1073), .Z(n1068) );
  XNOR U990 ( .A(n687), .B(n1074), .Z(n675) );
  XNOR U991 ( .A(n673), .B(n688), .Z(n1074) );
  XOR U992 ( .A(n682), .B(n680), .Z(n688) );
  NOR U993 ( .A(n1076), .B(n1077), .Z(n678) );
  OR U994 ( .A(n1078), .B(n1079), .Z(n1075) );
  OR U995 ( .A(n1080), .B(n1081), .Z(n682) );
  OR U996 ( .A(n1082), .B(n1083), .Z(n673) );
  XOR U997 ( .A(n689), .B(n1084), .Z(n687) );
  XOR U998 ( .A(n690), .B(n684), .Z(n1084) );
  NOR U999 ( .A(n1085), .B(n1086), .Z(n684) );
  OR U1000 ( .A(n1087), .B(n1088), .Z(n690) );
  AND U1001 ( .A(n1089), .B(n1090), .Z(n689) );
  OR U1002 ( .A(n1091), .B(n1092), .Z(n1090) );
  OR U1003 ( .A(n1093), .B(n1094), .Z(n1089) );
  XOR U1004 ( .A(n692), .B(n715), .Z(n1095) );
  XNOR U1005 ( .A(n706), .B(n707), .Z(n715) );
  XOR U1006 ( .A(n701), .B(n699), .Z(n707) );
  AND U1007 ( .A(n1096), .B(n697), .Z(n699) );
  OR U1008 ( .A(n1097), .B(n1098), .Z(n697) );
  OR U1009 ( .A(n1099), .B(n1100), .Z(n1096) );
  NOR U1010 ( .A(n1101), .B(n1102), .Z(n701) );
  XOR U1011 ( .A(n708), .B(n1103), .Z(n706) );
  XOR U1012 ( .A(n709), .B(n703), .Z(n1103) );
  NOR U1013 ( .A(n1104), .B(n1105), .Z(n703) );
  OR U1014 ( .A(n1106), .B(n1107), .Z(n709) );
  AND U1015 ( .A(n1108), .B(n1109), .Z(n708) );
  OR U1016 ( .A(n1110), .B(n1111), .Z(n1109) );
  OR U1017 ( .A(n1112), .B(n1113), .Z(n1108) );
  OR U1018 ( .A(n1114), .B(n1115), .Z(n692) );
  XNOR U1019 ( .A(n725), .B(n1116), .Z(n713) );
  XNOR U1020 ( .A(n711), .B(n726), .Z(n1116) );
  XOR U1021 ( .A(n720), .B(n718), .Z(n726) );
  NOR U1022 ( .A(n1118), .B(n1119), .Z(n716) );
  OR U1023 ( .A(n1120), .B(n1121), .Z(n1117) );
  OR U1024 ( .A(n1122), .B(n1123), .Z(n720) );
  OR U1025 ( .A(n1124), .B(n1125), .Z(n711) );
  XOR U1026 ( .A(n727), .B(n1126), .Z(n725) );
  XOR U1027 ( .A(n728), .B(n722), .Z(n1126) );
  NOR U1028 ( .A(n1127), .B(n1128), .Z(n722) );
  OR U1029 ( .A(n1129), .B(n1130), .Z(n728) );
  AND U1030 ( .A(n1131), .B(n1132), .Z(n727) );
  OR U1031 ( .A(n1133), .B(n1134), .Z(n1132) );
  OR U1032 ( .A(n1135), .B(n1136), .Z(n1131) );
  NANDN U1033 ( .A(n1137), .B(n1138), .Z(n654) );
  XNOR U1034 ( .A(n772), .B(n1139), .Z(n733) );
  XOR U1035 ( .A(n730), .B(n773), .Z(n1139) );
  XOR U1036 ( .A(n745), .B(n746), .Z(n754) );
  XOR U1037 ( .A(n740), .B(n738), .Z(n746) );
  AND U1038 ( .A(n1140), .B(n736), .Z(n738) );
  OR U1039 ( .A(n1141), .B(n1142), .Z(n736) );
  OR U1040 ( .A(n1143), .B(n1144), .Z(n1140) );
  NOR U1041 ( .A(n1145), .B(n1146), .Z(n740) );
  XOR U1042 ( .A(n747), .B(n1147), .Z(n745) );
  XOR U1043 ( .A(n748), .B(n742), .Z(n1147) );
  NOR U1044 ( .A(n1148), .B(n1149), .Z(n742) );
  OR U1045 ( .A(n1150), .B(n1151), .Z(n748) );
  AND U1046 ( .A(n1152), .B(n1153), .Z(n747) );
  OR U1047 ( .A(n1154), .B(n1155), .Z(n1153) );
  OR U1048 ( .A(n1156), .B(n1157), .Z(n1152) );
  XNOR U1049 ( .A(n764), .B(n1158), .Z(n752) );
  XNOR U1050 ( .A(n750), .B(n765), .Z(n1158) );
  XOR U1051 ( .A(n759), .B(n757), .Z(n765) );
  NOR U1052 ( .A(n1160), .B(n1161), .Z(n755) );
  OR U1053 ( .A(n1162), .B(n1163), .Z(n1159) );
  OR U1054 ( .A(n1164), .B(n1165), .Z(n759) );
  OR U1055 ( .A(n1166), .B(n1167), .Z(n750) );
  XOR U1056 ( .A(n766), .B(n1168), .Z(n764) );
  XOR U1057 ( .A(n767), .B(n761), .Z(n1168) );
  NOR U1058 ( .A(n1169), .B(n1170), .Z(n761) );
  OR U1059 ( .A(n1171), .B(n1172), .Z(n767) );
  AND U1060 ( .A(n1173), .B(n1174), .Z(n766) );
  OR U1061 ( .A(n1175), .B(n1176), .Z(n1174) );
  OR U1062 ( .A(n1177), .B(n1178), .Z(n1173) );
  NOR U1063 ( .A(n1179), .B(n1180), .Z(n730) );
  XNOR U1064 ( .A(n791), .B(n1181), .Z(n772) );
  XNOR U1065 ( .A(n769), .B(n792), .Z(n1181) );
  XNOR U1066 ( .A(n783), .B(n784), .Z(n792) );
  XOR U1067 ( .A(n778), .B(n776), .Z(n784) );
  AND U1068 ( .A(n1182), .B(n774), .Z(n776) );
  OR U1069 ( .A(n1183), .B(n1184), .Z(n774) );
  OR U1070 ( .A(n1185), .B(n1186), .Z(n1182) );
  NOR U1071 ( .A(n1187), .B(n1188), .Z(n778) );
  XOR U1072 ( .A(n785), .B(n1189), .Z(n783) );
  XOR U1073 ( .A(n786), .B(n780), .Z(n1189) );
  NOR U1074 ( .A(n1190), .B(n1191), .Z(n780) );
  OR U1075 ( .A(n1192), .B(n1193), .Z(n786) );
  AND U1076 ( .A(n1194), .B(n1195), .Z(n785) );
  OR U1077 ( .A(n1196), .B(n1197), .Z(n1195) );
  OR U1078 ( .A(n1198), .B(n1199), .Z(n1194) );
  XNOR U1079 ( .A(n801), .B(n1202), .Z(n791) );
  XNOR U1080 ( .A(n788), .B(n803), .Z(n1202) );
  XOR U1081 ( .A(n797), .B(n795), .Z(n803) );
  NOR U1082 ( .A(n1204), .B(n1205), .Z(n793) );
  OR U1083 ( .A(n1206), .B(n1207), .Z(n1203) );
  OR U1084 ( .A(n1208), .B(n1209), .Z(n797) );
  NANDN U1085 ( .A(n1210), .B(n1211), .Z(n788) );
  XNOR U1086 ( .A(n804), .B(n1212), .Z(n801) );
  XOR U1087 ( .A(n805), .B(n799), .Z(n1212) );
  AND U1088 ( .A(n1213), .B(n1214), .Z(n799) );
  OR U1089 ( .A(n1215), .B(n1216), .Z(n805) );
  AND U1090 ( .A(n1217), .B(n1218), .Z(n804) );
  OR U1091 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR U1092 ( .A(n1053), .B(n1054), .Z(o[0]) );
  XOR U1093 ( .A(n865), .B(n864), .Z(n1054) );
  XNOR U1094 ( .A(n833), .B(n832), .Z(n864) );
  XNOR U1095 ( .A(n807), .B(n808), .Z(n814) );
  XNOR U1096 ( .A(n811), .B(n812), .Z(n808) );
  XNOR U1097 ( .A(y[159]), .B(x[159]), .Z(n812) );
  XNOR U1098 ( .A(y[158]), .B(x[158]), .Z(n811) );
  XNOR U1099 ( .A(n809), .B(n810), .Z(n807) );
  XNOR U1100 ( .A(y[157]), .B(x[157]), .Z(n810) );
  XNOR U1101 ( .A(y[156]), .B(x[156]), .Z(n809) );
  XNOR U1102 ( .A(n822), .B(n823), .Z(n815) );
  XNOR U1103 ( .A(n817), .B(n816), .Z(n823) );
  XNOR U1104 ( .A(y[155]), .B(x[155]), .Z(n816) );
  XNOR U1105 ( .A(y[154]), .B(x[154]), .Z(n817) );
  XNOR U1106 ( .A(n820), .B(n821), .Z(n822) );
  XNOR U1107 ( .A(y[153]), .B(x[153]), .Z(n821) );
  XNOR U1108 ( .A(y[152]), .B(x[152]), .Z(n820) );
  XNOR U1109 ( .A(n826), .B(n827), .Z(n835) );
  XNOR U1110 ( .A(n830), .B(n831), .Z(n827) );
  XNOR U1111 ( .A(y[151]), .B(x[151]), .Z(n831) );
  XNOR U1112 ( .A(y[150]), .B(x[150]), .Z(n830) );
  XNOR U1113 ( .A(n828), .B(n829), .Z(n826) );
  XNOR U1114 ( .A(y[149]), .B(x[149]), .Z(n829) );
  XNOR U1115 ( .A(y[148]), .B(x[148]), .Z(n828) );
  XNOR U1116 ( .A(n843), .B(n844), .Z(n836) );
  XNOR U1117 ( .A(n838), .B(n837), .Z(n844) );
  XNOR U1118 ( .A(y[147]), .B(x[147]), .Z(n837) );
  XNOR U1119 ( .A(y[146]), .B(x[146]), .Z(n838) );
  XNOR U1120 ( .A(n841), .B(n842), .Z(n843) );
  XNOR U1121 ( .A(y[145]), .B(x[145]), .Z(n842) );
  XNOR U1122 ( .A(y[144]), .B(x[144]), .Z(n841) );
  XNOR U1123 ( .A(n875), .B(n874), .Z(n865) );
  XNOR U1124 ( .A(n847), .B(n848), .Z(n854) );
  XNOR U1125 ( .A(n851), .B(n852), .Z(n848) );
  XNOR U1126 ( .A(y[143]), .B(x[143]), .Z(n852) );
  XNOR U1127 ( .A(y[142]), .B(x[142]), .Z(n851) );
  XNOR U1128 ( .A(n849), .B(n850), .Z(n847) );
  XNOR U1129 ( .A(y[141]), .B(x[141]), .Z(n850) );
  XNOR U1130 ( .A(y[140]), .B(x[140]), .Z(n849) );
  XNOR U1131 ( .A(n862), .B(n863), .Z(n855) );
  XNOR U1132 ( .A(n857), .B(n856), .Z(n863) );
  XNOR U1133 ( .A(y[139]), .B(x[139]), .Z(n856) );
  XNOR U1134 ( .A(y[138]), .B(x[138]), .Z(n857) );
  XNOR U1135 ( .A(n860), .B(n861), .Z(n862) );
  XNOR U1136 ( .A(y[137]), .B(x[137]), .Z(n861) );
  XNOR U1137 ( .A(y[136]), .B(x[136]), .Z(n860) );
  XNOR U1138 ( .A(n868), .B(n869), .Z(n877) );
  XNOR U1139 ( .A(n872), .B(n873), .Z(n869) );
  XNOR U1140 ( .A(y[135]), .B(x[135]), .Z(n873) );
  XNOR U1141 ( .A(y[134]), .B(x[134]), .Z(n872) );
  XNOR U1142 ( .A(n870), .B(n871), .Z(n868) );
  XNOR U1143 ( .A(y[133]), .B(x[133]), .Z(n871) );
  XNOR U1144 ( .A(y[132]), .B(x[132]), .Z(n870) );
  XNOR U1145 ( .A(n885), .B(n886), .Z(n878) );
  XNOR U1146 ( .A(n880), .B(n879), .Z(n886) );
  XNOR U1147 ( .A(y[131]), .B(x[131]), .Z(n879) );
  XNOR U1148 ( .A(y[130]), .B(x[130]), .Z(n880) );
  XNOR U1149 ( .A(n883), .B(n884), .Z(n885) );
  XNOR U1150 ( .A(y[129]), .B(x[129]), .Z(n884) );
  XNOR U1151 ( .A(y[128]), .B(x[128]), .Z(n883) );
  XOR U1152 ( .A(n1138), .B(n1137), .Z(n1053) );
  XNOR U1153 ( .A(n1010), .B(n1009), .Z(n1137) );
  XNOR U1154 ( .A(n947), .B(n946), .Z(n1009) );
  XNOR U1155 ( .A(n915), .B(n914), .Z(n946) );
  XNOR U1156 ( .A(n889), .B(n890), .Z(n896) );
  XNOR U1157 ( .A(n893), .B(n894), .Z(n890) );
  XNOR U1158 ( .A(y[127]), .B(x[127]), .Z(n894) );
  XNOR U1159 ( .A(y[126]), .B(x[126]), .Z(n893) );
  XNOR U1160 ( .A(n891), .B(n892), .Z(n889) );
  XNOR U1161 ( .A(y[125]), .B(x[125]), .Z(n892) );
  XNOR U1162 ( .A(y[124]), .B(x[124]), .Z(n891) );
  XNOR U1163 ( .A(n904), .B(n905), .Z(n897) );
  XNOR U1164 ( .A(n899), .B(n898), .Z(n905) );
  XNOR U1165 ( .A(y[123]), .B(x[123]), .Z(n898) );
  XNOR U1166 ( .A(y[122]), .B(x[122]), .Z(n899) );
  XNOR U1167 ( .A(n902), .B(n903), .Z(n904) );
  XNOR U1168 ( .A(y[121]), .B(x[121]), .Z(n903) );
  XNOR U1169 ( .A(y[120]), .B(x[120]), .Z(n902) );
  XNOR U1170 ( .A(n908), .B(n909), .Z(n917) );
  XNOR U1171 ( .A(n912), .B(n913), .Z(n909) );
  XNOR U1172 ( .A(y[119]), .B(x[119]), .Z(n913) );
  XNOR U1173 ( .A(y[118]), .B(x[118]), .Z(n912) );
  XNOR U1174 ( .A(n910), .B(n911), .Z(n908) );
  XNOR U1175 ( .A(y[117]), .B(x[117]), .Z(n911) );
  XNOR U1176 ( .A(y[116]), .B(x[116]), .Z(n910) );
  XNOR U1177 ( .A(n925), .B(n926), .Z(n918) );
  XNOR U1178 ( .A(n920), .B(n919), .Z(n926) );
  XNOR U1179 ( .A(y[115]), .B(x[115]), .Z(n919) );
  XNOR U1180 ( .A(y[114]), .B(x[114]), .Z(n920) );
  XNOR U1181 ( .A(n923), .B(n924), .Z(n925) );
  XNOR U1182 ( .A(y[113]), .B(x[113]), .Z(n924) );
  XNOR U1183 ( .A(y[112]), .B(x[112]), .Z(n923) );
  XNOR U1184 ( .A(n957), .B(n956), .Z(n947) );
  XNOR U1185 ( .A(n929), .B(n930), .Z(n936) );
  XNOR U1186 ( .A(n933), .B(n934), .Z(n930) );
  XNOR U1187 ( .A(y[111]), .B(x[111]), .Z(n934) );
  XNOR U1188 ( .A(y[110]), .B(x[110]), .Z(n933) );
  XNOR U1189 ( .A(n931), .B(n932), .Z(n929) );
  XNOR U1190 ( .A(y[109]), .B(x[109]), .Z(n932) );
  XNOR U1191 ( .A(y[108]), .B(x[108]), .Z(n931) );
  XNOR U1192 ( .A(n944), .B(n945), .Z(n937) );
  XNOR U1193 ( .A(n939), .B(n938), .Z(n945) );
  XNOR U1194 ( .A(y[107]), .B(x[107]), .Z(n938) );
  XNOR U1195 ( .A(y[106]), .B(x[106]), .Z(n939) );
  XNOR U1196 ( .A(n942), .B(n943), .Z(n944) );
  XNOR U1197 ( .A(y[105]), .B(x[105]), .Z(n943) );
  XNOR U1198 ( .A(y[104]), .B(x[104]), .Z(n942) );
  XNOR U1199 ( .A(n950), .B(n951), .Z(n959) );
  XNOR U1200 ( .A(n954), .B(n955), .Z(n951) );
  XNOR U1201 ( .A(y[103]), .B(x[103]), .Z(n955) );
  XNOR U1202 ( .A(y[102]), .B(x[102]), .Z(n954) );
  XNOR U1203 ( .A(n952), .B(n953), .Z(n950) );
  XNOR U1204 ( .A(y[101]), .B(x[101]), .Z(n953) );
  XNOR U1205 ( .A(y[100]), .B(x[100]), .Z(n952) );
  XNOR U1206 ( .A(n967), .B(n968), .Z(n960) );
  XNOR U1207 ( .A(n962), .B(n961), .Z(n968) );
  XNOR U1208 ( .A(y[99]), .B(x[99]), .Z(n961) );
  XNOR U1209 ( .A(y[98]), .B(x[98]), .Z(n962) );
  XNOR U1210 ( .A(n965), .B(n966), .Z(n967) );
  XNOR U1211 ( .A(y[97]), .B(x[97]), .Z(n966) );
  XNOR U1212 ( .A(y[96]), .B(x[96]), .Z(n965) );
  XNOR U1213 ( .A(n1031), .B(n1030), .Z(n1010) );
  XNOR U1214 ( .A(n997), .B(n996), .Z(n1030) );
  XNOR U1215 ( .A(n971), .B(n972), .Z(n978) );
  XNOR U1216 ( .A(n975), .B(n976), .Z(n972) );
  XNOR U1217 ( .A(y[95]), .B(x[95]), .Z(n976) );
  XNOR U1218 ( .A(y[94]), .B(x[94]), .Z(n975) );
  XNOR U1219 ( .A(n973), .B(n974), .Z(n971) );
  XNOR U1220 ( .A(y[93]), .B(x[93]), .Z(n974) );
  XNOR U1221 ( .A(y[92]), .B(x[92]), .Z(n973) );
  XNOR U1222 ( .A(n986), .B(n987), .Z(n979) );
  XNOR U1223 ( .A(n981), .B(n980), .Z(n987) );
  XNOR U1224 ( .A(y[91]), .B(x[91]), .Z(n980) );
  XNOR U1225 ( .A(y[90]), .B(x[90]), .Z(n981) );
  XNOR U1226 ( .A(n984), .B(n985), .Z(n986) );
  XNOR U1227 ( .A(y[89]), .B(x[89]), .Z(n985) );
  XNOR U1228 ( .A(y[88]), .B(x[88]), .Z(n984) );
  XNOR U1229 ( .A(n990), .B(n991), .Z(n999) );
  XNOR U1230 ( .A(n994), .B(n995), .Z(n991) );
  XNOR U1231 ( .A(y[87]), .B(x[87]), .Z(n995) );
  XNOR U1232 ( .A(y[86]), .B(x[86]), .Z(n994) );
  XNOR U1233 ( .A(n992), .B(n993), .Z(n990) );
  XNOR U1234 ( .A(y[85]), .B(x[85]), .Z(n993) );
  XNOR U1235 ( .A(y[84]), .B(x[84]), .Z(n992) );
  XNOR U1236 ( .A(n1007), .B(n1008), .Z(n1000) );
  XNOR U1237 ( .A(n1002), .B(n1001), .Z(n1008) );
  XNOR U1238 ( .A(y[83]), .B(x[83]), .Z(n1001) );
  XNOR U1239 ( .A(y[82]), .B(x[82]), .Z(n1002) );
  XNOR U1240 ( .A(n1005), .B(n1006), .Z(n1007) );
  XNOR U1241 ( .A(y[81]), .B(x[81]), .Z(n1006) );
  XNOR U1242 ( .A(y[80]), .B(x[80]), .Z(n1005) );
  XNOR U1243 ( .A(n1041), .B(n1040), .Z(n1031) );
  XNOR U1244 ( .A(n1013), .B(n1014), .Z(n1020) );
  XNOR U1245 ( .A(n1017), .B(n1018), .Z(n1014) );
  XNOR U1246 ( .A(y[79]), .B(x[79]), .Z(n1018) );
  XNOR U1247 ( .A(y[78]), .B(x[78]), .Z(n1017) );
  XNOR U1248 ( .A(n1015), .B(n1016), .Z(n1013) );
  XNOR U1249 ( .A(y[77]), .B(x[77]), .Z(n1016) );
  XNOR U1250 ( .A(y[76]), .B(x[76]), .Z(n1015) );
  XNOR U1251 ( .A(n1028), .B(n1029), .Z(n1021) );
  XNOR U1252 ( .A(n1023), .B(n1022), .Z(n1029) );
  XNOR U1253 ( .A(y[75]), .B(x[75]), .Z(n1022) );
  XNOR U1254 ( .A(y[74]), .B(x[74]), .Z(n1023) );
  XNOR U1255 ( .A(n1026), .B(n1027), .Z(n1028) );
  XNOR U1256 ( .A(y[73]), .B(x[73]), .Z(n1027) );
  XNOR U1257 ( .A(y[72]), .B(x[72]), .Z(n1026) );
  XNOR U1258 ( .A(n1034), .B(n1035), .Z(n1043) );
  XNOR U1259 ( .A(n1038), .B(n1039), .Z(n1035) );
  XNOR U1260 ( .A(y[71]), .B(x[71]), .Z(n1039) );
  XNOR U1261 ( .A(y[70]), .B(x[70]), .Z(n1038) );
  XNOR U1262 ( .A(n1036), .B(n1037), .Z(n1034) );
  XNOR U1263 ( .A(y[69]), .B(x[69]), .Z(n1037) );
  XNOR U1264 ( .A(y[68]), .B(x[68]), .Z(n1036) );
  XNOR U1265 ( .A(n1051), .B(n1052), .Z(n1044) );
  XNOR U1266 ( .A(n1046), .B(n1045), .Z(n1052) );
  XNOR U1267 ( .A(y[67]), .B(x[67]), .Z(n1045) );
  XNOR U1268 ( .A(y[66]), .B(x[66]), .Z(n1046) );
  XNOR U1269 ( .A(n1049), .B(n1050), .Z(n1051) );
  XNOR U1270 ( .A(y[65]), .B(x[65]), .Z(n1050) );
  XNOR U1271 ( .A(y[64]), .B(x[64]), .Z(n1049) );
  XOR U1272 ( .A(n1179), .B(n1180), .Z(n1138) );
  XNOR U1273 ( .A(n1115), .B(n1114), .Z(n1180) );
  XNOR U1274 ( .A(n1083), .B(n1082), .Z(n1114) );
  XNOR U1275 ( .A(n1057), .B(n1058), .Z(n1064) );
  XNOR U1276 ( .A(n1061), .B(n1062), .Z(n1058) );
  XNOR U1277 ( .A(y[63]), .B(x[63]), .Z(n1062) );
  XNOR U1278 ( .A(y[62]), .B(x[62]), .Z(n1061) );
  XNOR U1279 ( .A(n1059), .B(n1060), .Z(n1057) );
  XNOR U1280 ( .A(y[61]), .B(x[61]), .Z(n1060) );
  XNOR U1281 ( .A(y[60]), .B(x[60]), .Z(n1059) );
  XNOR U1282 ( .A(n1072), .B(n1073), .Z(n1065) );
  XNOR U1283 ( .A(n1067), .B(n1066), .Z(n1073) );
  XNOR U1284 ( .A(y[59]), .B(x[59]), .Z(n1066) );
  XNOR U1285 ( .A(y[58]), .B(x[58]), .Z(n1067) );
  XNOR U1286 ( .A(n1070), .B(n1071), .Z(n1072) );
  XNOR U1287 ( .A(y[57]), .B(x[57]), .Z(n1071) );
  XNOR U1288 ( .A(y[56]), .B(x[56]), .Z(n1070) );
  XNOR U1289 ( .A(n1076), .B(n1077), .Z(n1085) );
  XNOR U1290 ( .A(n1080), .B(n1081), .Z(n1077) );
  XNOR U1291 ( .A(y[55]), .B(x[55]), .Z(n1081) );
  XNOR U1292 ( .A(y[54]), .B(x[54]), .Z(n1080) );
  XNOR U1293 ( .A(n1078), .B(n1079), .Z(n1076) );
  XNOR U1294 ( .A(y[53]), .B(x[53]), .Z(n1079) );
  XNOR U1295 ( .A(y[52]), .B(x[52]), .Z(n1078) );
  XNOR U1296 ( .A(n1093), .B(n1094), .Z(n1086) );
  XNOR U1297 ( .A(n1088), .B(n1087), .Z(n1094) );
  XNOR U1298 ( .A(y[51]), .B(x[51]), .Z(n1087) );
  XNOR U1299 ( .A(y[50]), .B(x[50]), .Z(n1088) );
  XNOR U1300 ( .A(n1091), .B(n1092), .Z(n1093) );
  XNOR U1301 ( .A(y[49]), .B(x[49]), .Z(n1092) );
  XNOR U1302 ( .A(y[48]), .B(x[48]), .Z(n1091) );
  XNOR U1303 ( .A(n1125), .B(n1124), .Z(n1115) );
  XNOR U1304 ( .A(n1097), .B(n1098), .Z(n1104) );
  XNOR U1305 ( .A(n1101), .B(n1102), .Z(n1098) );
  XNOR U1306 ( .A(y[47]), .B(x[47]), .Z(n1102) );
  XNOR U1307 ( .A(y[46]), .B(x[46]), .Z(n1101) );
  XNOR U1308 ( .A(n1099), .B(n1100), .Z(n1097) );
  XNOR U1309 ( .A(y[45]), .B(x[45]), .Z(n1100) );
  XNOR U1310 ( .A(y[44]), .B(x[44]), .Z(n1099) );
  XNOR U1311 ( .A(n1112), .B(n1113), .Z(n1105) );
  XNOR U1312 ( .A(n1107), .B(n1106), .Z(n1113) );
  XNOR U1313 ( .A(y[43]), .B(x[43]), .Z(n1106) );
  XNOR U1314 ( .A(y[42]), .B(x[42]), .Z(n1107) );
  XNOR U1315 ( .A(n1110), .B(n1111), .Z(n1112) );
  XNOR U1316 ( .A(y[41]), .B(x[41]), .Z(n1111) );
  XNOR U1317 ( .A(y[40]), .B(x[40]), .Z(n1110) );
  XNOR U1318 ( .A(n1118), .B(n1119), .Z(n1127) );
  XNOR U1319 ( .A(n1122), .B(n1123), .Z(n1119) );
  XNOR U1320 ( .A(y[39]), .B(x[39]), .Z(n1123) );
  XNOR U1321 ( .A(y[38]), .B(x[38]), .Z(n1122) );
  XNOR U1322 ( .A(n1120), .B(n1121), .Z(n1118) );
  XNOR U1323 ( .A(y[37]), .B(x[37]), .Z(n1121) );
  XNOR U1324 ( .A(y[36]), .B(x[36]), .Z(n1120) );
  XNOR U1325 ( .A(n1135), .B(n1136), .Z(n1128) );
  XNOR U1326 ( .A(n1130), .B(n1129), .Z(n1136) );
  XNOR U1327 ( .A(y[35]), .B(x[35]), .Z(n1129) );
  XNOR U1328 ( .A(y[34]), .B(x[34]), .Z(n1130) );
  XNOR U1329 ( .A(n1133), .B(n1134), .Z(n1135) );
  XNOR U1330 ( .A(y[33]), .B(x[33]), .Z(n1134) );
  XNOR U1331 ( .A(y[32]), .B(x[32]), .Z(n1133) );
  XOR U1332 ( .A(n1201), .B(n1200), .Z(n1179) );
  XNOR U1333 ( .A(n1167), .B(n1166), .Z(n1200) );
  XNOR U1334 ( .A(n1141), .B(n1142), .Z(n1148) );
  XNOR U1335 ( .A(n1145), .B(n1146), .Z(n1142) );
  XNOR U1336 ( .A(y[31]), .B(x[31]), .Z(n1146) );
  XNOR U1337 ( .A(y[30]), .B(x[30]), .Z(n1145) );
  XNOR U1338 ( .A(n1143), .B(n1144), .Z(n1141) );
  XNOR U1339 ( .A(y[29]), .B(x[29]), .Z(n1144) );
  XNOR U1340 ( .A(y[28]), .B(x[28]), .Z(n1143) );
  XNOR U1341 ( .A(n1156), .B(n1157), .Z(n1149) );
  XNOR U1342 ( .A(n1151), .B(n1150), .Z(n1157) );
  XNOR U1343 ( .A(y[27]), .B(x[27]), .Z(n1150) );
  XNOR U1344 ( .A(y[26]), .B(x[26]), .Z(n1151) );
  XNOR U1345 ( .A(n1154), .B(n1155), .Z(n1156) );
  XNOR U1346 ( .A(y[25]), .B(x[25]), .Z(n1155) );
  XNOR U1347 ( .A(y[24]), .B(x[24]), .Z(n1154) );
  XNOR U1348 ( .A(n1160), .B(n1161), .Z(n1169) );
  XNOR U1349 ( .A(n1164), .B(n1165), .Z(n1161) );
  XNOR U1350 ( .A(y[23]), .B(x[23]), .Z(n1165) );
  XNOR U1351 ( .A(y[22]), .B(x[22]), .Z(n1164) );
  XNOR U1352 ( .A(n1162), .B(n1163), .Z(n1160) );
  XNOR U1353 ( .A(y[21]), .B(x[21]), .Z(n1163) );
  XNOR U1354 ( .A(y[20]), .B(x[20]), .Z(n1162) );
  XNOR U1355 ( .A(n1177), .B(n1178), .Z(n1170) );
  XNOR U1356 ( .A(n1172), .B(n1171), .Z(n1178) );
  XNOR U1357 ( .A(y[19]), .B(x[19]), .Z(n1171) );
  XNOR U1358 ( .A(y[18]), .B(x[18]), .Z(n1172) );
  XNOR U1359 ( .A(n1175), .B(n1176), .Z(n1177) );
  XNOR U1360 ( .A(y[17]), .B(x[17]), .Z(n1176) );
  XNOR U1361 ( .A(y[16]), .B(x[16]), .Z(n1175) );
  XNOR U1362 ( .A(n1211), .B(n1210), .Z(n1201) );
  XNOR U1363 ( .A(n1183), .B(n1184), .Z(n1190) );
  XNOR U1364 ( .A(n1187), .B(n1188), .Z(n1184) );
  XNOR U1365 ( .A(y[15]), .B(x[15]), .Z(n1188) );
  XNOR U1366 ( .A(y[14]), .B(x[14]), .Z(n1187) );
  XNOR U1367 ( .A(n1185), .B(n1186), .Z(n1183) );
  XNOR U1368 ( .A(y[13]), .B(x[13]), .Z(n1186) );
  XNOR U1369 ( .A(y[12]), .B(x[12]), .Z(n1185) );
  XNOR U1370 ( .A(n1198), .B(n1199), .Z(n1191) );
  XNOR U1371 ( .A(n1193), .B(n1192), .Z(n1199) );
  XNOR U1372 ( .A(y[11]), .B(x[11]), .Z(n1192) );
  XNOR U1373 ( .A(y[10]), .B(x[10]), .Z(n1193) );
  XNOR U1374 ( .A(n1196), .B(n1197), .Z(n1198) );
  XNOR U1375 ( .A(y[9]), .B(x[9]), .Z(n1197) );
  XNOR U1376 ( .A(y[8]), .B(x[8]), .Z(n1196) );
  XOR U1377 ( .A(n1213), .B(n1214), .Z(n1211) );
  XOR U1378 ( .A(n1204), .B(n1205), .Z(n1214) );
  XNOR U1379 ( .A(n1208), .B(n1209), .Z(n1205) );
  XNOR U1380 ( .A(y[7]), .B(x[7]), .Z(n1209) );
  XNOR U1381 ( .A(y[6]), .B(x[6]), .Z(n1208) );
  XNOR U1382 ( .A(n1206), .B(n1207), .Z(n1204) );
  XNOR U1383 ( .A(y[5]), .B(x[5]), .Z(n1207) );
  XNOR U1384 ( .A(y[4]), .B(x[4]), .Z(n1206) );
  XNOR U1385 ( .A(n1221), .B(n1222), .Z(n1213) );
  XOR U1386 ( .A(n1216), .B(n1215), .Z(n1222) );
  XNOR U1387 ( .A(y[3]), .B(x[3]), .Z(n1215) );
  XNOR U1388 ( .A(y[2]), .B(x[2]), .Z(n1216) );
  XNOR U1389 ( .A(n1219), .B(n1220), .Z(n1221) );
  XNOR U1390 ( .A(y[1]), .B(x[1]), .Z(n1220) );
  XNOR U1391 ( .A(y[0]), .B(x[0]), .Z(n1219) );
endmodule

